module top( \CM_rd0[0]_pad  , \CM_rd0[10]_pad  , \CM_rd0[11]_pad  , \CM_rd0[12]_pad  , \CM_rd0[13]_pad  , \CM_rd0[14]_pad  , \CM_rd0[15]_pad  , \CM_rd0[16]_pad  , \CM_rd0[17]_pad  , \CM_rd0[18]_pad  , \CM_rd0[19]_pad  , \CM_rd0[1]_pad  , \CM_rd0[20]_pad  , \CM_rd0[21]_pad  , \CM_rd0[22]_pad  , \CM_rd0[23]_pad  , \CM_rd0[2]_pad  , \CM_rd0[3]_pad  , \CM_rd0[4]_pad  , \CM_rd0[5]_pad  , \CM_rd0[6]_pad  , \CM_rd0[7]_pad  , \CM_rd0[8]_pad  , \CM_rd0[9]_pad  , \CM_rd1[0]_pad  , \CM_rd1[10]_pad  , \CM_rd1[11]_pad  , \CM_rd1[12]_pad  , \CM_rd1[13]_pad  , \CM_rd1[14]_pad  , \CM_rd1[15]_pad  , \CM_rd1[16]_pad  , \CM_rd1[17]_pad  , \CM_rd1[18]_pad  , \CM_rd1[19]_pad  , \CM_rd1[1]_pad  , \CM_rd1[20]_pad  , \CM_rd1[21]_pad  , \CM_rd1[22]_pad  , \CM_rd1[23]_pad  , \CM_rd1[2]_pad  , \CM_rd1[3]_pad  , \CM_rd1[4]_pad  , \CM_rd1[5]_pad  , \CM_rd1[6]_pad  , \CM_rd1[7]_pad  , \CM_rd1[8]_pad  , \CM_rd1[9]_pad  , \CM_rd2[0]_pad  , \CM_rd2[10]_pad  , \CM_rd2[11]_pad  , \CM_rd2[12]_pad  , \CM_rd2[13]_pad  , \CM_rd2[14]_pad  , \CM_rd2[15]_pad  , \CM_rd2[16]_pad  , \CM_rd2[17]_pad  , \CM_rd2[18]_pad  , \CM_rd2[19]_pad  , \CM_rd2[1]_pad  , \CM_rd2[20]_pad  , \CM_rd2[21]_pad  , \CM_rd2[22]_pad  , \CM_rd2[23]_pad  , \CM_rd2[2]_pad  , \CM_rd2[3]_pad  , \CM_rd2[4]_pad  , \CM_rd2[5]_pad  , \CM_rd2[6]_pad  , \CM_rd2[7]_pad  , \CM_rd2[8]_pad  , \CM_rd2[9]_pad  , \CM_rd3[0]_pad  , \CM_rd3[10]_pad  , \CM_rd3[11]_pad  , \CM_rd3[12]_pad  , \CM_rd3[13]_pad  , \CM_rd3[14]_pad  , \CM_rd3[15]_pad  , \CM_rd3[16]_pad  , \CM_rd3[17]_pad  , \CM_rd3[18]_pad  , \CM_rd3[19]_pad  , \CM_rd3[1]_pad  , \CM_rd3[20]_pad  , \CM_rd3[21]_pad  , \CM_rd3[22]_pad  , \CM_rd3[23]_pad  , \CM_rd3[2]_pad  , \CM_rd3[3]_pad  , \CM_rd3[4]_pad  , \CM_rd3[5]_pad  , \CM_rd3[6]_pad  , \CM_rd3[7]_pad  , \CM_rd3[8]_pad  , \CM_rd3[9]_pad  , \CM_rd4[0]_pad  , \CM_rd4[10]_pad  , \CM_rd4[11]_pad  , \CM_rd4[12]_pad  , \CM_rd4[13]_pad  , \CM_rd4[14]_pad  , \CM_rd4[15]_pad  , \CM_rd4[16]_pad  , \CM_rd4[17]_pad  , \CM_rd4[18]_pad  , \CM_rd4[19]_pad  , \CM_rd4[1]_pad  , \CM_rd4[20]_pad  , \CM_rd4[21]_pad  , \CM_rd4[22]_pad  , \CM_rd4[23]_pad  , \CM_rd4[2]_pad  , \CM_rd4[3]_pad  , \CM_rd4[4]_pad  , \CM_rd4[5]_pad  , \CM_rd4[6]_pad  , \CM_rd4[7]_pad  , \CM_rd4[8]_pad  , \CM_rd4[9]_pad  , \CM_rd5[0]_pad  , \CM_rd5[10]_pad  , \CM_rd5[11]_pad  , \CM_rd5[12]_pad  , \CM_rd5[13]_pad  , \CM_rd5[14]_pad  , \CM_rd5[15]_pad  , \CM_rd5[16]_pad  , \CM_rd5[17]_pad  , \CM_rd5[18]_pad  , \CM_rd5[19]_pad  , \CM_rd5[1]_pad  , \CM_rd5[20]_pad  , \CM_rd5[21]_pad  , \CM_rd5[22]_pad  , \CM_rd5[23]_pad  , \CM_rd5[2]_pad  , \CM_rd5[3]_pad  , \CM_rd5[4]_pad  , \CM_rd5[5]_pad  , \CM_rd5[6]_pad  , \CM_rd5[7]_pad  , \CM_rd5[8]_pad  , \CM_rd5[9]_pad  , \CM_rd6[0]_pad  , \CM_rd6[10]_pad  , \CM_rd6[11]_pad  , \CM_rd6[12]_pad  , \CM_rd6[13]_pad  , \CM_rd6[14]_pad  , \CM_rd6[15]_pad  , \CM_rd6[16]_pad  , \CM_rd6[17]_pad  , \CM_rd6[18]_pad  , \CM_rd6[19]_pad  , \CM_rd6[1]_pad  , \CM_rd6[20]_pad  , \CM_rd6[21]_pad  , \CM_rd6[22]_pad  , \CM_rd6[23]_pad  , \CM_rd6[2]_pad  , \CM_rd6[3]_pad  , \CM_rd6[4]_pad  , \CM_rd6[5]_pad  , \CM_rd6[6]_pad  , \CM_rd6[7]_pad  , \CM_rd6[8]_pad  , \CM_rd6[9]_pad  , \CM_rd7[0]_pad  , \CM_rd7[10]_pad  , \CM_rd7[11]_pad  , \CM_rd7[12]_pad  , \CM_rd7[13]_pad  , \CM_rd7[14]_pad  , \CM_rd7[15]_pad  , \CM_rd7[16]_pad  , \CM_rd7[17]_pad  , \CM_rd7[18]_pad  , \CM_rd7[19]_pad  , \CM_rd7[1]_pad  , \CM_rd7[20]_pad  , \CM_rd7[21]_pad  , \CM_rd7[22]_pad  , \CM_rd7[23]_pad  , \CM_rd7[2]_pad  , \CM_rd7[3]_pad  , \CM_rd7[4]_pad  , \CM_rd7[5]_pad  , \CM_rd7[6]_pad  , \CM_rd7[7]_pad  , \CM_rd7[8]_pad  , \CM_rd7[9]_pad  , \CM_rdm[0]_pad  , \CM_rdm[10]_pad  , \CM_rdm[11]_pad  , \CM_rdm[12]_pad  , \CM_rdm[13]_pad  , \CM_rdm[14]_pad  , \CM_rdm[15]_pad  , \CM_rdm[16]_pad  , \CM_rdm[17]_pad  , \CM_rdm[18]_pad  , \CM_rdm[19]_pad  , \CM_rdm[1]_pad  , \CM_rdm[20]_pad  , \CM_rdm[21]_pad  , \CM_rdm[22]_pad  , \CM_rdm[23]_pad  , \CM_rdm[2]_pad  , \CM_rdm[3]_pad  , \CM_rdm[4]_pad  , \CM_rdm[5]_pad  , \CM_rdm[6]_pad  , \CM_rdm[7]_pad  , \CM_rdm[8]_pad  , \CM_rdm[9]_pad  , \DM_rd0[0]_pad  , \DM_rd0[10]_pad  , \DM_rd0[11]_pad  , \DM_rd0[12]_pad  , \DM_rd0[13]_pad  , \DM_rd0[14]_pad  , \DM_rd0[15]_pad  , \DM_rd0[1]_pad  , \DM_rd0[2]_pad  , \DM_rd0[3]_pad  , \DM_rd0[4]_pad  , \DM_rd0[5]_pad  , \DM_rd0[6]_pad  , \DM_rd0[7]_pad  , \DM_rd0[8]_pad  , \DM_rd0[9]_pad  , \DM_rd1[0]_pad  , \DM_rd1[10]_pad  , \DM_rd1[11]_pad  , \DM_rd1[12]_pad  , \DM_rd1[13]_pad  , \DM_rd1[14]_pad  , \DM_rd1[15]_pad  , \DM_rd1[1]_pad  , \DM_rd1[2]_pad  , \DM_rd1[3]_pad  , \DM_rd1[4]_pad  , \DM_rd1[5]_pad  , \DM_rd1[6]_pad  , \DM_rd1[7]_pad  , \DM_rd1[8]_pad  , \DM_rd1[9]_pad  , \DM_rd2[0]_pad  , \DM_rd2[10]_pad  , \DM_rd2[11]_pad  , \DM_rd2[12]_pad  , \DM_rd2[13]_pad  , \DM_rd2[14]_pad  , \DM_rd2[15]_pad  , \DM_rd2[1]_pad  , \DM_rd2[2]_pad  , \DM_rd2[3]_pad  , \DM_rd2[4]_pad  , \DM_rd2[5]_pad  , \DM_rd2[6]_pad  , \DM_rd2[7]_pad  , \DM_rd2[8]_pad  , \DM_rd2[9]_pad  , \DM_rd3[0]_pad  , \DM_rd3[10]_pad  , \DM_rd3[11]_pad  , \DM_rd3[12]_pad  , \DM_rd3[13]_pad  , \DM_rd3[14]_pad  , \DM_rd3[15]_pad  , \DM_rd3[1]_pad  , \DM_rd3[2]_pad  , \DM_rd3[3]_pad  , \DM_rd3[4]_pad  , \DM_rd3[5]_pad  , \DM_rd3[6]_pad  , \DM_rd3[7]_pad  , \DM_rd3[8]_pad  , \DM_rd3[9]_pad  , \DM_rd4[0]_pad  , \DM_rd4[10]_pad  , \DM_rd4[11]_pad  , \DM_rd4[12]_pad  , \DM_rd4[13]_pad  , \DM_rd4[14]_pad  , \DM_rd4[15]_pad  , \DM_rd4[1]_pad  , \DM_rd4[2]_pad  , \DM_rd4[3]_pad  , \DM_rd4[4]_pad  , \DM_rd4[5]_pad  , \DM_rd4[6]_pad  , \DM_rd4[7]_pad  , \DM_rd4[8]_pad  , \DM_rd4[9]_pad  , \DM_rd5[0]_pad  , \DM_rd5[10]_pad  , \DM_rd5[11]_pad  , \DM_rd5[12]_pad  , \DM_rd5[13]_pad  , \DM_rd5[14]_pad  , \DM_rd5[15]_pad  , \DM_rd5[1]_pad  , \DM_rd5[2]_pad  , \DM_rd5[3]_pad  , \DM_rd5[4]_pad  , \DM_rd5[5]_pad  , \DM_rd5[6]_pad  , \DM_rd5[7]_pad  , \DM_rd5[8]_pad  , \DM_rd5[9]_pad  , \DM_rd6[0]_pad  , \DM_rd6[10]_pad  , \DM_rd6[11]_pad  , \DM_rd6[12]_pad  , \DM_rd6[13]_pad  , \DM_rd6[14]_pad  , \DM_rd6[15]_pad  , \DM_rd6[1]_pad  , \DM_rd6[2]_pad  , \DM_rd6[3]_pad  , \DM_rd6[4]_pad  , \DM_rd6[5]_pad  , \DM_rd6[6]_pad  , \DM_rd6[7]_pad  , \DM_rd6[8]_pad  , \DM_rd6[9]_pad  , \DM_rd7[0]_pad  , \DM_rd7[10]_pad  , \DM_rd7[11]_pad  , \DM_rd7[12]_pad  , \DM_rd7[13]_pad  , \DM_rd7[14]_pad  , \DM_rd7[15]_pad  , \DM_rd7[1]_pad  , \DM_rd7[2]_pad  , \DM_rd7[3]_pad  , \DM_rd7[4]_pad  , \DM_rd7[5]_pad  , \DM_rd7[6]_pad  , \DM_rd7[7]_pad  , \DM_rd7[8]_pad  , \DM_rd7[9]_pad  , \DM_rdm[0]_pad  , \DM_rdm[10]_pad  , \DM_rdm[11]_pad  , \DM_rdm[12]_pad  , \DM_rdm[13]_pad  , \DM_rdm[14]_pad  , \DM_rdm[15]_pad  , \DM_rdm[1]_pad  , \DM_rdm[2]_pad  , \DM_rdm[3]_pad  , \DM_rdm[4]_pad  , \DM_rdm[5]_pad  , \DM_rdm[6]_pad  , \DM_rdm[7]_pad  , \DM_rdm[8]_pad  , \DM_rdm[9]_pad  , IACKn_pad , \IRFS0_pad  , \IRFS1_pad  , \ISCLK0_pad  , \ISCLK1_pad  , \ITFS0_pad  , \ITFS1_pad  , \PIO_oe[0]_pad  , \PIO_oe[10]_pad  , \PIO_oe[11]_pad  , \PIO_oe[1]_pad  , \PIO_oe[2]_pad  , \PIO_oe[3]_pad  , \PIO_oe[4]_pad  , \PIO_oe[5]_pad  , \PIO_oe[6]_pad  , \PIO_oe[7]_pad  , \PIO_oe[8]_pad  , \PIO_oe[9]_pad  , \PIO_out[0]_pad  , \PIO_out[10]_pad  , \PIO_out[11]_pad  , \PIO_out[1]_pad  , \PIO_out[2]_pad  , \PIO_out[3]_pad  , \PIO_out[4]_pad  , \PIO_out[5]_pad  , \PIO_out[6]_pad  , \PIO_out[7]_pad  , \PIO_out[8]_pad  , \PIO_out[9]_pad  , PM_bdry_sel_pad , \PM_rd0[0]_pad  , \PM_rd0[10]_pad  , \PM_rd0[11]_pad  , \PM_rd0[12]_pad  , \PM_rd0[13]_pad  , \PM_rd0[14]_pad  , \PM_rd0[15]_pad  , \PM_rd0[1]_pad  , \PM_rd0[2]_pad  , \PM_rd0[3]_pad  , \PM_rd0[4]_pad  , \PM_rd0[5]_pad  , \PM_rd0[6]_pad  , \PM_rd0[7]_pad  , \PM_rd0[8]_pad  , \PM_rd0[9]_pad  , \PM_rd1[0]_pad  , \PM_rd1[10]_pad  , \PM_rd1[11]_pad  , \PM_rd1[12]_pad  , \PM_rd1[13]_pad  , \PM_rd1[14]_pad  , \PM_rd1[15]_pad  , \PM_rd1[1]_pad  , \PM_rd1[2]_pad  , \PM_rd1[3]_pad  , \PM_rd1[4]_pad  , \PM_rd1[5]_pad  , \PM_rd1[6]_pad  , \PM_rd1[7]_pad  , \PM_rd1[8]_pad  , \PM_rd1[9]_pad  , \PM_rd2[0]_pad  , \PM_rd2[10]_pad  , \PM_rd2[11]_pad  , \PM_rd2[12]_pad  , \PM_rd2[13]_pad  , \PM_rd2[14]_pad  , \PM_rd2[15]_pad  , \PM_rd2[1]_pad  , \PM_rd2[2]_pad  , \PM_rd2[3]_pad  , \PM_rd2[4]_pad  , \PM_rd2[5]_pad  , \PM_rd2[6]_pad  , \PM_rd2[7]_pad  , \PM_rd2[8]_pad  , \PM_rd2[9]_pad  , \PM_rd3[0]_pad  , \PM_rd3[10]_pad  , \PM_rd3[11]_pad  , \PM_rd3[12]_pad  , \PM_rd3[13]_pad  , \PM_rd3[14]_pad  , \PM_rd3[15]_pad  , \PM_rd3[1]_pad  , \PM_rd3[2]_pad  , \PM_rd3[3]_pad  , \PM_rd3[4]_pad  , \PM_rd3[5]_pad  , \PM_rd3[6]_pad  , \PM_rd3[7]_pad  , \PM_rd3[8]_pad  , \PM_rd3[9]_pad  , \PM_rd4[0]_pad  , \PM_rd4[10]_pad  , \PM_rd4[11]_pad  , \PM_rd4[12]_pad  , \PM_rd4[13]_pad  , \PM_rd4[14]_pad  , \PM_rd4[15]_pad  , \PM_rd4[1]_pad  , \PM_rd4[2]_pad  , \PM_rd4[3]_pad  , \PM_rd4[4]_pad  , \PM_rd4[5]_pad  , \PM_rd4[6]_pad  , \PM_rd4[7]_pad  , \PM_rd4[8]_pad  , \PM_rd4[9]_pad  , \PM_rd5[0]_pad  , \PM_rd5[10]_pad  , \PM_rd5[11]_pad  , \PM_rd5[12]_pad  , \PM_rd5[13]_pad  , \PM_rd5[14]_pad  , \PM_rd5[15]_pad  , \PM_rd5[1]_pad  , \PM_rd5[2]_pad  , \PM_rd5[3]_pad  , \PM_rd5[4]_pad  , \PM_rd5[5]_pad  , \PM_rd5[6]_pad  , \PM_rd5[7]_pad  , \PM_rd5[8]_pad  , \PM_rd5[9]_pad  , \PM_rd6[0]_pad  , \PM_rd6[10]_pad  , \PM_rd6[11]_pad  , \PM_rd6[12]_pad  , \PM_rd6[13]_pad  , \PM_rd6[14]_pad  , \PM_rd6[15]_pad  , \PM_rd6[1]_pad  , \PM_rd6[2]_pad  , \PM_rd6[3]_pad  , \PM_rd6[4]_pad  , \PM_rd6[5]_pad  , \PM_rd6[6]_pad  , \PM_rd6[7]_pad  , \PM_rd6[8]_pad  , \PM_rd6[9]_pad  , \PM_rd7[0]_pad  , \PM_rd7[10]_pad  , \PM_rd7[11]_pad  , \PM_rd7[12]_pad  , \PM_rd7[13]_pad  , \PM_rd7[14]_pad  , \PM_rd7[15]_pad  , \PM_rd7[1]_pad  , \PM_rd7[2]_pad  , \PM_rd7[3]_pad  , \PM_rd7[4]_pad  , \PM_rd7[5]_pad  , \PM_rd7[6]_pad  , \PM_rd7[7]_pad  , \PM_rd7[8]_pad  , \PM_rd7[9]_pad  , PWDACK_pad , T_BMODE_pad , T_BRn_pad , T_CLKI_OSC_pad , T_CLKI_PLL_pad , \T_ED[0]_pad  , \T_ED[10]_pad  , \T_ED[11]_pad  , \T_ED[12]_pad  , \T_ED[13]_pad  , \T_ED[14]_pad  , \T_ED[15]_pad  , \T_ED[1]_pad  , \T_ED[2]_pad  , \T_ED[3]_pad  , \T_ED[4]_pad  , \T_ED[5]_pad  , \T_ED[6]_pad  , \T_ED[7]_pad  , \T_ED[8]_pad  , \T_ED[9]_pad  , T_ICE_RSTn_pad , T_ID_pad , T_IMS_pad , T_IRDn_pad , \T_IRQ0n_pad  , \T_IRQ1n_pad  , \T_IRQ2n_pad  , \T_IRQE0n_pad  , \T_IRQE1n_pad  , \T_IRQL1n_pad  , T_ISn_pad , T_IWRn_pad , T_MMAP_pad , \T_PIOin[0]_pad  , \T_PIOin[10]_pad  , \T_PIOin[11]_pad  , \T_PIOin[1]_pad  , \T_PIOin[2]_pad  , \T_PIOin[3]_pad  , \T_PIOin[4]_pad  , \T_PIOin[5]_pad  , \T_PIOin[6]_pad  , \T_PIOin[7]_pad  , \T_PIOin[8]_pad  , \T_PIOin[9]_pad  , T_PWDn_pad , \T_RD0_pad  , \T_RD1_pad  , \T_RFS0_pad  , \T_RFS1_pad  , T_RSTn_pad , \T_SCLK0_pad  , \T_SCLK1_pad  , T_Sel_PLL_pad , \T_TFS0_pad  , \T_TFS1_pad  , \T_TMODE[0]_pad  , \T_TMODE[1]_pad  , \auctl_BSack_reg/NET0131  , \auctl_DSack_reg/NET0131  , \auctl_R0Sack_reg/NET0131  , \auctl_R1Sack_reg/NET0131  , \auctl_RST_reg/P0001  , \auctl_STEAL_reg/NET0131  , \auctl_T0Sack_reg/NET0131  , \auctl_T1Sack_reg/NET0131  , \bdma_BCTL_reg[0]/NET0131  , \bdma_BCTL_reg[10]/NET0131  , \bdma_BCTL_reg[11]/NET0131  , \bdma_BCTL_reg[12]/NET0131  , \bdma_BCTL_reg[13]/NET0131  , \bdma_BCTL_reg[14]/NET0131  , \bdma_BCTL_reg[15]/NET0131  , \bdma_BCTL_reg[1]/NET0131  , \bdma_BCTL_reg[2]/NET0131  , \bdma_BCTL_reg[3]/NET0131  , \bdma_BCTL_reg[4]/NET0131  , \bdma_BCTL_reg[5]/NET0131  , \bdma_BCTL_reg[6]/NET0131  , \bdma_BCTL_reg[7]/NET0131  , \bdma_BCTL_reg[8]/NET0131  , \bdma_BCTL_reg[9]/NET0131  , \bdma_BDMA_boot_reg/NET0131_reg_syn_10  , \bdma_BDMA_boot_reg/NET0131_reg_syn_2  , \bdma_BDMA_boot_reg/NET0131_reg_syn_8  , \bdma_BDMAmode_reg/NET0131  , \bdma_BEAD_reg[0]/NET0131  , \bdma_BEAD_reg[10]/NET0131  , \bdma_BEAD_reg[11]/NET0131  , \bdma_BEAD_reg[12]/NET0131  , \bdma_BEAD_reg[13]/NET0131  , \bdma_BEAD_reg[1]/NET0131  , \bdma_BEAD_reg[2]/NET0131  , \bdma_BEAD_reg[3]/NET0131  , \bdma_BEAD_reg[4]/NET0131  , \bdma_BEAD_reg[5]/NET0131  , \bdma_BEAD_reg[6]/NET0131  , \bdma_BEAD_reg[7]/NET0131  , \bdma_BEAD_reg[8]/NET0131  , \bdma_BEAD_reg[9]/NET0131  , \bdma_BIAD_reg[0]/NET0131  , \bdma_BIAD_reg[10]/NET0131  , \bdma_BIAD_reg[11]/NET0131  , \bdma_BIAD_reg[12]/NET0131  , \bdma_BIAD_reg[13]/NET0131  , \bdma_BIAD_reg[1]/NET0131  , \bdma_BIAD_reg[2]/NET0131  , \bdma_BIAD_reg[3]/NET0131  , \bdma_BIAD_reg[4]/NET0131  , \bdma_BIAD_reg[5]/NET0131  , \bdma_BIAD_reg[6]/NET0131  , \bdma_BIAD_reg[7]/NET0131  , \bdma_BIAD_reg[8]/NET0131  , \bdma_BIAD_reg[9]/NET0131  , \bdma_BM_cyc_reg/P0001  , \bdma_BMcyc_del_reg/P0001  , \bdma_BOVL_reg[0]/NET0131  , \bdma_BOVL_reg[10]/NET0131  , \bdma_BOVL_reg[11]/NET0131  , \bdma_BOVL_reg[1]/NET0131  , \bdma_BOVL_reg[2]/NET0131  , \bdma_BOVL_reg[3]/NET0131  , \bdma_BOVL_reg[4]/NET0131  , \bdma_BOVL_reg[5]/NET0131  , \bdma_BOVL_reg[6]/NET0131  , \bdma_BOVL_reg[7]/NET0131  , \bdma_BOVL_reg[8]/NET0131  , \bdma_BOVL_reg[9]/NET0131  , \bdma_BRST_s2_reg/NET0131  , \bdma_BRdataBUF_reg[0]/P0001  , \bdma_BRdataBUF_reg[10]/P0001  , \bdma_BRdataBUF_reg[11]/P0001  , \bdma_BRdataBUF_reg[12]/P0001  , \bdma_BRdataBUF_reg[13]/P0001  , \bdma_BRdataBUF_reg[14]/P0001  , \bdma_BRdataBUF_reg[15]/P0001  , \bdma_BRdataBUF_reg[16]/P0001  , \bdma_BRdataBUF_reg[17]/P0001  , \bdma_BRdataBUF_reg[18]/P0001  , \bdma_BRdataBUF_reg[19]/P0001  , \bdma_BRdataBUF_reg[1]/P0001  , \bdma_BRdataBUF_reg[20]/P0001  , \bdma_BRdataBUF_reg[21]/P0001  , \bdma_BRdataBUF_reg[22]/P0001  , \bdma_BRdataBUF_reg[23]/P0001  , \bdma_BRdataBUF_reg[2]/P0001  , \bdma_BRdataBUF_reg[3]/P0001  , \bdma_BRdataBUF_reg[4]/P0001  , \bdma_BRdataBUF_reg[5]/P0001  , \bdma_BRdataBUF_reg[6]/P0001  , \bdma_BRdataBUF_reg[7]/P0001  , \bdma_BRdataBUF_reg[8]/P0001  , \bdma_BRdataBUF_reg[9]/P0001  , \bdma_BSreq_reg/NET0131  , \bdma_BWCOUNT_reg[0]/NET0131  , \bdma_BWCOUNT_reg[10]/NET0131  , \bdma_BWCOUNT_reg[11]/NET0131  , \bdma_BWCOUNT_reg[12]/NET0131  , \bdma_BWCOUNT_reg[13]/NET0131  , \bdma_BWCOUNT_reg[1]/NET0131  , \bdma_BWCOUNT_reg[2]/NET0131  , \bdma_BWCOUNT_reg[3]/NET0131  , \bdma_BWCOUNT_reg[4]/NET0131  , \bdma_BWCOUNT_reg[5]/NET0131_reg_syn_2  , \bdma_BWCOUNT_reg[5]/NET0131_reg_syn_8  , \bdma_BWCOUNT_reg[6]/NET0131  , \bdma_BWCOUNT_reg[7]/NET0131  , \bdma_BWCOUNT_reg[8]/NET0131  , \bdma_BWCOUNT_reg[9]/NET0131  , \bdma_BWRn_reg/NET0131  , \bdma_BWcnt_reg[0]/NET0131  , \bdma_BWcnt_reg[1]/NET0131  , \bdma_BWcnt_reg[2]/NET0131  , \bdma_BWcnt_reg[3]/NET0131  , \bdma_BWcnt_reg[4]/NET0131  , \bdma_BWdataBUF_h_reg[0]/P0001  , \bdma_BWdataBUF_h_reg[10]/P0001  , \bdma_BWdataBUF_h_reg[11]/P0001  , \bdma_BWdataBUF_h_reg[12]/P0001  , \bdma_BWdataBUF_h_reg[13]/P0001  , \bdma_BWdataBUF_h_reg[14]/P0001  , \bdma_BWdataBUF_h_reg[15]/P0001  , \bdma_BWdataBUF_h_reg[16]/P0001  , \bdma_BWdataBUF_h_reg[17]/P0001  , \bdma_BWdataBUF_h_reg[18]/P0001  , \bdma_BWdataBUF_h_reg[19]/P0001  , \bdma_BWdataBUF_h_reg[1]/P0001  , \bdma_BWdataBUF_h_reg[20]/P0001  , \bdma_BWdataBUF_h_reg[21]/P0001  , \bdma_BWdataBUF_h_reg[22]/P0001  , \bdma_BWdataBUF_h_reg[23]/P0001  , \bdma_BWdataBUF_h_reg[2]/P0001  , \bdma_BWdataBUF_h_reg[3]/P0001  , \bdma_BWdataBUF_h_reg[4]/P0001  , \bdma_BWdataBUF_h_reg[5]/P0001  , \bdma_BWdataBUF_h_reg[6]/P0001  , \bdma_BWdataBUF_h_reg[7]/P0001  , \bdma_BWdataBUF_h_reg[8]/P0001  , \bdma_BWdataBUF_h_reg[9]/P0001  , \bdma_BWdataBUF_reg[0]/P0001  , \bdma_BWdataBUF_reg[1]/P0001  , \bdma_BWdataBUF_reg[2]/P0001  , \bdma_BWdataBUF_reg[3]/P0001  , \bdma_BWdataBUF_reg[4]/P0001  , \bdma_BWdataBUF_reg[5]/P0001  , \bdma_BWdataBUF_reg[6]/P0001  , \bdma_BWdataBUF_reg[7]/P0001  , \bdma_CMcnt_reg[0]/NET0131  , \bdma_CMcnt_reg[1]/NET0131  , \bdma_DM_2nd_reg/NET0131  , \bdma_RST_pin_reg/P0001  , \bdma_WRlat_reg/P0001  , \clkc_Awake_reg/NET0131  , \clkc_CLKOUT_reg/NET0131  , \clkc_CTR_cnt_reg[0]/NET0131  , \clkc_CTR_cnt_reg[1]/NET0131  , \clkc_Cnt128_reg/NET0131  , \clkc_Cnt4096_reg/NET0131  , \clkc_Cnt4096_s1_reg/NET0131  , \clkc_Cnt4096_s2_reg/NET0131  , \clkc_DSPoff_reg/NET0131  , \clkc_OSCoff_reg/NET0131  , \clkc_OSCoff_set_reg/P0001  , \clkc_OUTcnt_reg[0]/NET0131  , \clkc_OUTcnt_reg[1]/NET0131  , \clkc_OUTcnt_reg[2]/NET0131  , \clkc_OUTcnt_reg[3]/NET0131  , \clkc_OUTcnt_reg[4]/NET0131  , \clkc_OUTcnt_reg[5]/NET0131  , \clkc_OUTcnt_reg[6]/NET0131  , \clkc_RSTtext_reg/P0001  , \clkc_SIDLE_s1_reg/NET0131  , \clkc_SIDLE_s2_reg/NET0131  , \clkc_SLEEP_reg/NET0131  , \clkc_STBY_reg/NET0131  , \clkc_STDcnt_reg[0]/NET0131  , \clkc_STDcnt_reg[10]/NET0131  , \clkc_STDcnt_reg[1]/NET0131  , \clkc_STDcnt_reg[2]/NET0131  , \clkc_STDcnt_reg[3]/NET0131  , \clkc_STDcnt_reg[4]/NET0131  , \clkc_STDcnt_reg[5]/NET0131  , \clkc_STDcnt_reg[6]/NET0131  , \clkc_STDcnt_reg[7]/NET0131  , \clkc_STDcnt_reg[8]/NET0131  , \clkc_STDcnt_reg[9]/NET0131  , \clkc_SlowDn_reg/NET0131  , \clkc_SlowDn_s1_reg/P0001  , \clkc_SlowDn_s2_reg/P0001  , \clkc_ckSTDCLK_STDCLK_reg_Q_reg/NET0131  , \clkc_ckr_reg_DO_reg[0]/NET0131  , \clkc_ckr_reg_DO_reg[10]/NET0131  , \clkc_ckr_reg_DO_reg[11]/NET0131  , \clkc_ckr_reg_DO_reg[12]/NET0131  , \clkc_ckr_reg_DO_reg[13]/NET0131  , \clkc_ckr_reg_DO_reg[14]/NET0131  , \clkc_ckr_reg_DO_reg[15]/NET0131  , \clkc_ckr_reg_DO_reg[1]/NET0131  , \clkc_ckr_reg_DO_reg[2]/NET0131  , \clkc_ckr_reg_DO_reg[3]/NET0131  , \clkc_ckr_reg_DO_reg[4]/NET0131  , \clkc_ckr_reg_DO_reg[5]/NET0131  , \clkc_ckr_reg_DO_reg[6]/NET0131  , \clkc_ckr_reg_DO_reg[7]/NET0131  , \clkc_ckr_reg_DO_reg[8]/NET0131  , \clkc_ckr_reg_DO_reg[9]/NET0131  , \clkc_oscntr_reg_DO_reg[0]/NET0131  , \clkc_oscntr_reg_DO_reg[10]/NET0131  , \clkc_oscntr_reg_DO_reg[11]/NET0131  , \clkc_oscntr_reg_DO_reg[1]/NET0131  , \clkc_oscntr_reg_DO_reg[2]/NET0131  , \clkc_oscntr_reg_DO_reg[3]/NET0131  , \clkc_oscntr_reg_DO_reg[4]/NET0131  , \clkc_oscntr_reg_DO_reg[5]/NET0131  , \clkc_oscntr_reg_DO_reg[6]/NET0131  , \clkc_oscntr_reg_DO_reg[7]/NET0131  , \clkc_oscntr_reg_DO_reg[8]/NET0131  , \clkc_oscntr_reg_DO_reg[9]/NET0131  , \core_c_dec_ALUop_E_reg/P0001  , \core_c_dec_BR_Ed_reg/P0001  , \core_c_dec_Call_Ed_reg/P0001  , \core_c_dec_DIVQ_E_reg/P0001  , \core_c_dec_DIVS_E_reg/P0001  , \core_c_dec_DU_Eg_reg/P0001  , \core_c_dec_Double_E_reg/P0001  , \core_c_dec_Dummy_E_reg/NET0131  , \core_c_dec_EXIT_E_reg/P0001  , \core_c_dec_IDLE_Eg_reg/P0001  , \core_c_dec_IRE_reg[0]/NET0131  , \core_c_dec_IRE_reg[10]/NET0131  , \core_c_dec_IRE_reg[11]/NET0131  , \core_c_dec_IRE_reg[12]/NET0131  , \core_c_dec_IRE_reg[13]/NET0131  , \core_c_dec_IRE_reg[14]/NET0131  , \core_c_dec_IRE_reg[15]/NET0131  , \core_c_dec_IRE_reg[16]/NET0131  , \core_c_dec_IRE_reg[17]/NET0131  , \core_c_dec_IRE_reg[18]/NET0131  , \core_c_dec_IRE_reg[19]/NET0131  , \core_c_dec_IRE_reg[1]/NET0131  , \core_c_dec_IRE_reg[2]/NET0131  , \core_c_dec_IRE_reg[3]/NET0131  , \core_c_dec_IRE_reg[4]/NET0131  , \core_c_dec_IRE_reg[5]/NET0131  , \core_c_dec_IRE_reg[6]/NET0131  , \core_c_dec_IRE_reg[7]/NET0131  , \core_c_dec_IRE_reg[8]/NET0131  , \core_c_dec_IRE_reg[9]/NET0131  , \core_c_dec_IR_reg[0]/NET0131  , \core_c_dec_IR_reg[10]/NET0131  , \core_c_dec_IR_reg[11]/NET0131  , \core_c_dec_IR_reg[12]/NET0131  , \core_c_dec_IR_reg[13]/NET0131  , \core_c_dec_IR_reg[14]/NET0131  , \core_c_dec_IR_reg[15]/NET0131  , \core_c_dec_IR_reg[16]/NET0131  , \core_c_dec_IR_reg[17]/NET0131  , \core_c_dec_IR_reg[18]/NET0131  , \core_c_dec_IR_reg[19]/NET0131  , \core_c_dec_IR_reg[1]/NET0131  , \core_c_dec_IR_reg[20]/NET0131  , \core_c_dec_IR_reg[21]/NET0131  , \core_c_dec_IR_reg[22]/NET0131  , \core_c_dec_IR_reg[23]/NET0131  , \core_c_dec_IR_reg[2]/NET0131  , \core_c_dec_IR_reg[3]/NET0131  , \core_c_dec_IR_reg[4]/NET0131  , \core_c_dec_IR_reg[5]/NET0131  , \core_c_dec_IR_reg[6]/NET0131  , \core_c_dec_IR_reg[7]/NET0131  , \core_c_dec_IR_reg[8]/NET0131  , \core_c_dec_IR_reg[9]/NET0131  , \core_c_dec_Long_Cg_reg/P0001  , \core_c_dec_Long_Eg_reg/P0001  , \core_c_dec_MACdep_Eg_reg/P0001  , \core_c_dec_MACop_E_reg/P0001  , \core_c_dec_MFALU_Ei_reg/NET0131  , \core_c_dec_MFAR_E_reg/P0001  , \core_c_dec_MFASTAT_E_reg/P0001  , \core_c_dec_MFAX0_E_reg/P0001  , \core_c_dec_MFAX1_E_reg/P0001  , \core_c_dec_MFAY0_E_reg/P0001  , \core_c_dec_MFAY1_E_reg/P0001  , \core_c_dec_MFCNTR_E_reg/P0001  , \core_c_dec_MFDAG1_Ei_reg/NET0131  , \core_c_dec_MFDAG2_Ei_reg/NET0131  , \core_c_dec_MFDMOVL_E_reg/P0001  , \core_c_dec_MFICNTL_E_reg/P0001  , \core_c_dec_MFIDR_E_reg/P0001  , \core_c_dec_MFIMASK_E_reg/P0001  , \core_c_dec_MFIreg_E_reg[0]/P0001  , \core_c_dec_MFIreg_E_reg[1]/P0001  , \core_c_dec_MFIreg_E_reg[2]/P0001  , \core_c_dec_MFIreg_E_reg[3]/P0001  , \core_c_dec_MFIreg_E_reg[4]/P0001  , \core_c_dec_MFIreg_E_reg[5]/P0001  , \core_c_dec_MFIreg_E_reg[6]/P0001  , \core_c_dec_MFIreg_E_reg[7]/P0001  , \core_c_dec_MFLreg_E_reg[0]/P0001  , \core_c_dec_MFLreg_E_reg[1]/P0001  , \core_c_dec_MFLreg_E_reg[2]/P0001  , \core_c_dec_MFLreg_E_reg[3]/P0001  , \core_c_dec_MFLreg_E_reg[4]/P0001  , \core_c_dec_MFLreg_E_reg[5]/P0001  , \core_c_dec_MFLreg_E_reg[6]/P0001  , \core_c_dec_MFLreg_E_reg[7]/P0001  , \core_c_dec_MFMAC_Ei_reg/NET0131  , \core_c_dec_MFMR0_E_reg/P0001  , \core_c_dec_MFMR1_E_reg/P0001  , \core_c_dec_MFMR2_E_reg/P0001  , \core_c_dec_MFMSTAT_E_reg/P0001  , \core_c_dec_MFMX0_E_reg/P0001  , \core_c_dec_MFMX1_E_reg/P0001  , \core_c_dec_MFMY0_E_reg/P0001  , \core_c_dec_MFMY1_E_reg/P0001  , \core_c_dec_MFMreg_E_reg[0]/P0001  , \core_c_dec_MFMreg_E_reg[1]/P0001  , \core_c_dec_MFMreg_E_reg[2]/P0001  , \core_c_dec_MFMreg_E_reg[3]/P0001  , \core_c_dec_MFMreg_E_reg[4]/P0001  , \core_c_dec_MFMreg_E_reg[5]/P0001  , \core_c_dec_MFMreg_E_reg[6]/P0001  , \core_c_dec_MFMreg_E_reg[7]/P0001  , \core_c_dec_MFPMOVL_E_reg/P0001  , \core_c_dec_MFPSQ_Ei_reg/NET0131  , \core_c_dec_MFRX0_E_reg/P0001  , \core_c_dec_MFRX1_E_reg/P0001  , \core_c_dec_MFSB_E_reg/P0001  , \core_c_dec_MFSE_E_reg/P0001  , \core_c_dec_MFSHT_Ei_reg/NET0131  , \core_c_dec_MFSI_E_reg/P0001  , \core_c_dec_MFSPT_Ei_reg/NET0131  , \core_c_dec_MFSR0_E_reg/P0001  , \core_c_dec_MFSR1_E_reg/P0001  , \core_c_dec_MFSSTAT_E_reg/P0001  , \core_c_dec_MFTX0_E_reg/P0001  , \core_c_dec_MFTX1_E_reg/P0001  , \core_c_dec_MFtoppcs_Eg_reg/P0001  , \core_c_dec_MTAR_E_reg/P0001  , \core_c_dec_MTASTAT_E_reg/P0001  , \core_c_dec_MTAX0_E_reg/P0001  , \core_c_dec_MTAX1_E_reg/P0001  , \core_c_dec_MTAY0_E_reg/P0001  , \core_c_dec_MTAY1_E_reg/P0001  , \core_c_dec_MTCNTR_Eg_reg/P0001  , \core_c_dec_MTDMOVL_E_reg/P0001  , \core_c_dec_MTICNTL_Eg_reg/P0001  , \core_c_dec_MTIDR_E_reg/P0001  , \core_c_dec_MTIFC_Eg_reg/P0001  , \core_c_dec_MTIMASK_Eg_reg/P0001  , \core_c_dec_MTIreg_E_reg[0]/P0001  , \core_c_dec_MTIreg_E_reg[1]/P0001  , \core_c_dec_MTIreg_E_reg[2]/P0001  , \core_c_dec_MTIreg_E_reg[3]/P0001  , \core_c_dec_MTIreg_E_reg[4]/P0001  , \core_c_dec_MTIreg_E_reg[5]/P0001  , \core_c_dec_MTIreg_E_reg[6]/P0001  , \core_c_dec_MTIreg_E_reg[7]/P0001  , \core_c_dec_MTLreg_E_reg[0]/P0001  , \core_c_dec_MTLreg_E_reg[1]/P0001  , \core_c_dec_MTLreg_E_reg[2]/P0001  , \core_c_dec_MTLreg_E_reg[3]/P0001  , \core_c_dec_MTLreg_E_reg[4]/P0001  , \core_c_dec_MTLreg_E_reg[5]/P0001  , \core_c_dec_MTLreg_E_reg[6]/P0001  , \core_c_dec_MTLreg_E_reg[7]/P0001  , \core_c_dec_MTMR0_E_reg/P0001  , \core_c_dec_MTMR1_E_reg/P0001  , \core_c_dec_MTMR2_E_reg/P0001  , \core_c_dec_MTMSTAT_Eg_reg/P0001  , \core_c_dec_MTMX0_E_reg/P0001  , \core_c_dec_MTMX1_E_reg/P0001  , \core_c_dec_MTMY0_E_reg/P0001  , \core_c_dec_MTMY1_E_reg/P0001  , \core_c_dec_MTMreg_E_reg[0]/P0001  , \core_c_dec_MTMreg_E_reg[1]/P0001  , \core_c_dec_MTMreg_E_reg[2]/P0001  , \core_c_dec_MTMreg_E_reg[3]/P0001  , \core_c_dec_MTMreg_E_reg[4]/P0001  , \core_c_dec_MTMreg_E_reg[5]/P0001  , \core_c_dec_MTMreg_E_reg[6]/P0001  , \core_c_dec_MTMreg_E_reg[7]/P0001  , \core_c_dec_MTOWRCNTR_Eg_reg/P0001  , \core_c_dec_MTPMOVL_E_reg/P0001  , \core_c_dec_MTRX0_E_reg/P0001  , \core_c_dec_MTRX1_E_reg/P0001  , \core_c_dec_MTSB_E_reg/P0001  , \core_c_dec_MTSE_E_reg/P0001  , \core_c_dec_MTSI_E_reg/P0001  , \core_c_dec_MTSR0_E_reg/P0001  , \core_c_dec_MTSR1_E_reg/P0001  , \core_c_dec_MTTX0_E_reg/P0001  , \core_c_dec_MTTX1_E_reg/P0001  , \core_c_dec_MTtoppcs_Eg_reg/P0001  , \core_c_dec_Modctl_Eg_reg/P0001  , \core_c_dec_MpopLP_Eg_reg/P0001  , \core_c_dec_NOP_E_reg/P0001  , \core_c_dec_Nrti_Ed_reg/P0001  , \core_c_dec_Nseq_Ed_reg/P0001  , \core_c_dec_PPclr_reg/P0001  , \core_c_dec_Post1_E_reg/P0001  , \core_c_dec_Post2_E_reg/P0001  , \core_c_dec_Prderr_Cg_reg/NET0131  , \core_c_dec_RET_Ed_reg/P0001  , \core_c_dec_RTI_Ed_reg/P0001  , \core_c_dec_SHTop_E_reg/P0001  , \core_c_dec_Stkctl_Eg_reg/P0001  , \core_c_dec_Usecond_E_reg/P0001  , \core_c_dec_accCM_E_reg/NET0131  , \core_c_dec_accPM_E_reg/P0001  , \core_c_dec_cdAM_E_reg/P0001  , \core_c_dec_imSHT_E_reg/P0001  , \core_c_dec_imm14_E_reg/P0001  , \core_c_dec_imm16_E_reg/P0001  , \core_c_dec_pMFALU_Ei_reg/NET0131  , \core_c_dec_pMFMAC_Ei_reg/NET0131  , \core_c_dec_pMFSHT_Ei_reg/NET0131  , \core_c_dec_rdCM_E_reg/NET0131  , \core_c_dec_satMR_E_reg/P0001  , \core_c_dec_updAF_E_reg/P0001  , \core_c_dec_updAR_E_reg/P0001  , \core_c_dec_updMF_E_reg/P0001  , \core_c_dec_updMR_E_reg/P0001  , \core_c_dec_updSR_E_reg/P0001  , \core_c_psq_CE_reg/NET0131  , \core_c_psq_CNTR_reg_DO_reg[0]/NET0131  , \core_c_psq_CNTR_reg_DO_reg[10]/NET0131  , \core_c_psq_CNTR_reg_DO_reg[11]/NET0131  , \core_c_psq_CNTR_reg_DO_reg[12]/NET0131  , \core_c_psq_CNTR_reg_DO_reg[13]/NET0131  , \core_c_psq_CNTR_reg_DO_reg[1]/NET0131  , \core_c_psq_CNTR_reg_DO_reg[2]/NET0131  , \core_c_psq_CNTR_reg_DO_reg[3]/NET0131  , \core_c_psq_CNTR_reg_DO_reg[4]/NET0131  , \core_c_psq_CNTR_reg_DO_reg[5]/NET0131  , \core_c_psq_CNTR_reg_DO_reg[6]/NET0131  , \core_c_psq_CNTR_reg_DO_reg[7]/NET0131  , \core_c_psq_CNTR_reg_DO_reg[8]/NET0131  , \core_c_psq_CNTR_reg_DO_reg[9]/NET0131  , \core_c_psq_CNTRval_reg/NET0131  , \core_c_psq_DMOVL_reg_DO_reg[0]/NET0131  , \core_c_psq_DMOVL_reg_DO_reg[1]/NET0131  , \core_c_psq_DMOVL_reg_DO_reg[2]/NET0131  , \core_c_psq_DMOVL_reg_DO_reg[3]/NET0131  , \core_c_psq_DRA_reg[0]/P0001  , \core_c_psq_DRA_reg[10]/P0001  , \core_c_psq_DRA_reg[11]/P0001  , \core_c_psq_DRA_reg[12]/P0001  , \core_c_psq_DRA_reg[13]/P0001  , \core_c_psq_DRA_reg[1]/P0001  , \core_c_psq_DRA_reg[2]/P0001  , \core_c_psq_DRA_reg[3]/P0001  , \core_c_psq_DRA_reg[4]/P0001  , \core_c_psq_DRA_reg[5]/P0001  , \core_c_psq_DRA_reg[6]/P0001  , \core_c_psq_DRA_reg[7]/P0001  , \core_c_psq_DRA_reg[8]/P0001  , \core_c_psq_DRA_reg[9]/P0001  , \core_c_psq_ECYC_reg/P0001  , \core_c_psq_EXA_reg[0]/P0001  , \core_c_psq_EXA_reg[10]/P0001  , \core_c_psq_EXA_reg[11]/P0001  , \core_c_psq_EXA_reg[12]/P0001  , \core_c_psq_EXA_reg[13]/P0001  , \core_c_psq_EXA_reg[1]/P0001  , \core_c_psq_EXA_reg[2]/P0001  , \core_c_psq_EXA_reg[3]/P0001  , \core_c_psq_EXA_reg[4]/P0001  , \core_c_psq_EXA_reg[5]/P0001  , \core_c_psq_EXA_reg[6]/P0001  , \core_c_psq_EXA_reg[7]/P0001  , \core_c_psq_EXA_reg[8]/P0001  , \core_c_psq_EXA_reg[9]/P0001  , \core_c_psq_Eqend_D_reg/P0001  , \core_c_psq_Eqend_Ed_reg/P0001  , \core_c_psq_ICNTL_reg_DO_reg[0]/NET0131  , \core_c_psq_ICNTL_reg_DO_reg[1]/NET0131  , \core_c_psq_ICNTL_reg_DO_reg[2]/NET0131  , \core_c_psq_ICNTL_reg_DO_reg[4]/NET0131  , \core_c_psq_IFA_reg[0]/P0001  , \core_c_psq_IFA_reg[10]/P0001  , \core_c_psq_IFA_reg[11]/P0001  , \core_c_psq_IFA_reg[12]/P0001  , \core_c_psq_IFA_reg[13]/P0001  , \core_c_psq_IFA_reg[1]/P0001  , \core_c_psq_IFA_reg[2]/P0001  , \core_c_psq_IFA_reg[3]/P0001  , \core_c_psq_IFA_reg[4]/P0001  , \core_c_psq_IFA_reg[5]/P0001  , \core_c_psq_IFA_reg[6]/P0001  , \core_c_psq_IFA_reg[7]/P0001  , \core_c_psq_IFA_reg[8]/P0001  , \core_c_psq_IFA_reg[9]/P0001  , \core_c_psq_IFC_reg[0]/NET0131  , \core_c_psq_IFC_reg[10]/NET0131  , \core_c_psq_IFC_reg[11]/NET0131  , \core_c_psq_IFC_reg[12]/NET0131  , \core_c_psq_IFC_reg[13]/NET0131  , \core_c_psq_IFC_reg[14]/NET0131  , \core_c_psq_IFC_reg[15]/NET0131  , \core_c_psq_IFC_reg[1]/NET0131  , \core_c_psq_IFC_reg[2]/NET0131  , \core_c_psq_IFC_reg[3]/NET0131  , \core_c_psq_IFC_reg[4]/NET0131  , \core_c_psq_IFC_reg[5]/NET0131  , \core_c_psq_IFC_reg[6]/NET0131  , \core_c_psq_IFC_reg[7]/NET0131  , \core_c_psq_IFC_reg[8]/NET0131  , \core_c_psq_IFC_reg[9]/NET0131  , \core_c_psq_IMASK_reg[0]/NET0131  , \core_c_psq_IMASK_reg[1]/NET0131  , \core_c_psq_IMASK_reg[2]/NET0131  , \core_c_psq_IMASK_reg[3]/NET0131  , \core_c_psq_IMASK_reg[4]/NET0131  , \core_c_psq_IMASK_reg[5]/NET0131  , \core_c_psq_IMASK_reg[6]/NET0131  , \core_c_psq_IMASK_reg[7]/NET0131  , \core_c_psq_IMASK_reg[8]/NET0131  , \core_c_psq_IMASK_reg[9]/NET0131  , \core_c_psq_INT_en_reg/NET0131  , \core_c_psq_Iact_E_reg[0]/NET0131  , \core_c_psq_Iact_E_reg[10]/NET0131  , \core_c_psq_Iact_E_reg[1]/NET0131  , \core_c_psq_Iact_E_reg[2]/NET0131  , \core_c_psq_Iact_E_reg[3]/NET0131  , \core_c_psq_Iact_E_reg[4]/NET0131  , \core_c_psq_Iact_E_reg[5]/NET0131  , \core_c_psq_Iact_E_reg[6]/NET0131  , \core_c_psq_Iact_E_reg[7]/NET0131  , \core_c_psq_Iact_E_reg[8]/NET0131  , \core_c_psq_Iact_E_reg[9]/NET0131  , \core_c_psq_Iflag_reg[0]/NET0131  , \core_c_psq_Iflag_reg[10]/NET0131  , \core_c_psq_Iflag_reg[11]/NET0131  , \core_c_psq_Iflag_reg[12]/NET0131  , \core_c_psq_Iflag_reg[1]/NET0131  , \core_c_psq_Iflag_reg[2]/NET0131  , \core_c_psq_Iflag_reg[3]/NET0131  , \core_c_psq_Iflag_reg[4]/NET0131  , \core_c_psq_Iflag_reg[5]/NET0131  , \core_c_psq_Iflag_reg[6]/NET0131  , \core_c_psq_Iflag_reg[7]/NET0131  , \core_c_psq_Iflag_reg[8]/NET0131  , \core_c_psq_Iflag_reg[9]/NET0131  , \core_c_psq_MGNT_reg/NET0131  , \core_c_psq_MREQ_reg/NET0131  , \core_c_psq_MSTAT_reg_DO_reg[0]/P0002  , \core_c_psq_MSTAT_reg_DO_reg[1]/NET0131  , \core_c_psq_MSTAT_reg_DO_reg[2]/NET0131  , \core_c_psq_MSTAT_reg_DO_reg[3]/NET0131  , \core_c_psq_MSTAT_reg_DO_reg[4]/NET0131  , \core_c_psq_MSTAT_reg_DO_reg[5]/NET0131  , \core_c_psq_MSTAT_reg_DO_reg[6]/NET0131  , \core_c_psq_PCS2or3_reg/NET0131  , \core_c_psq_PCS_reg[0]/NET0131  , \core_c_psq_PCS_reg[10]/NET0131  , \core_c_psq_PCS_reg[11]/NET0131  , \core_c_psq_PCS_reg[12]/NET0131  , \core_c_psq_PCS_reg[13]/NET0131  , \core_c_psq_PCS_reg[14]/NET0131  , \core_c_psq_PCS_reg[15]/NET0131  , \core_c_psq_PCS_reg[1]/NET0131  , \core_c_psq_PCS_reg[2]/NET0131  , \core_c_psq_PCS_reg[3]/NET0131  , \core_c_psq_PCS_reg[4]/NET0131  , \core_c_psq_PCS_reg[5]/NET0131  , \core_c_psq_PCS_reg[6]/NET0131  , \core_c_psq_PCS_reg[7]/NET0131  , \core_c_psq_PCS_reg[8]/NET0131  , \core_c_psq_PMOVL_regh_DO_reg[0]/NET0131  , \core_c_psq_PMOVL_regh_DO_reg[1]/NET0131  , \core_c_psq_PMOVL_regh_DO_reg[2]/NET0131  , \core_c_psq_PMOVL_regh_DO_reg[3]/NET0131  , \core_c_psq_PMOVL_regl_DO_reg[0]/NET0131  , \core_c_psq_PMOVL_regl_DO_reg[1]/NET0131  , \core_c_psq_PMOVL_regl_DO_reg[2]/NET0131  , \core_c_psq_PMOVL_regl_DO_reg[3]/NET0131  , \core_c_psq_SRST_reg/P0001  , \core_c_psq_SSTAT_reg[0]/NET0131  , \core_c_psq_SSTAT_reg[1]/NET0131  , \core_c_psq_SSTAT_reg[2]/NET0131  , \core_c_psq_SSTAT_reg[3]/NET0131  , \core_c_psq_SSTAT_reg[4]/NET0131  , \core_c_psq_SSTAT_reg[5]/NET0131  , \core_c_psq_SSTAT_reg[6]/NET0131  , \core_c_psq_SSTAT_reg[7]/NET0131  , \core_c_psq_TRAP_Eg_reg/NET0131  , \core_c_psq_TRAP_R_L_reg/NET0131  , \core_c_psq_T_IRQ0_s1_reg/P0001  , \core_c_psq_T_IRQ0p_reg/P0001  , \core_c_psq_T_IRQ1_s1_reg/P0001  , \core_c_psq_T_IRQ1p_reg/P0001  , \core_c_psq_T_IRQ2_s1_reg/P0001  , \core_c_psq_T_IRQ2p_reg/P0001  , \core_c_psq_T_IRQE0_reg/P0001  , \core_c_psq_T_IRQE0_s1_reg/P0001  , \core_c_psq_T_IRQE1_reg/P0001  , \core_c_psq_T_IRQE1_s1_reg/P0001  , \core_c_psq_T_IRQL0p_reg/P0001  , \core_c_psq_T_IRQL1p_reg/P0001  , \core_c_psq_T_PWRDN_reg/P0001  , \core_c_psq_T_PWRDN_s1_reg/P0001  , \core_c_psq_Taddr_Eb_reg[0]/P0001  , \core_c_psq_Taddr_Eb_reg[10]/P0001  , \core_c_psq_Taddr_Eb_reg[11]/P0001  , \core_c_psq_Taddr_Eb_reg[12]/P0001  , \core_c_psq_Taddr_Eb_reg[13]/P0001  , \core_c_psq_Taddr_Eb_reg[1]/P0001  , \core_c_psq_Taddr_Eb_reg[2]/P0001  , \core_c_psq_Taddr_Eb_reg[3]/P0001  , \core_c_psq_Taddr_Eb_reg[4]/P0001  , \core_c_psq_Taddr_Eb_reg[5]/P0001  , \core_c_psq_Taddr_Eb_reg[6]/P0001  , \core_c_psq_Taddr_Eb_reg[7]/P0001  , \core_c_psq_Taddr_Eb_reg[8]/P0001  , \core_c_psq_Taddr_Eb_reg[9]/P0001  , \core_c_psq_cntstk_cnts4x14_CNTcell_reg[0][0]/P0001  , \core_c_psq_cntstk_cnts4x14_CNTcell_reg[0][10]/P0001  , \core_c_psq_cntstk_cnts4x14_CNTcell_reg[0][11]/P0001  , \core_c_psq_cntstk_cnts4x14_CNTcell_reg[0][12]/P0001  , \core_c_psq_cntstk_cnts4x14_CNTcell_reg[0][13]/P0001  , \core_c_psq_cntstk_cnts4x14_CNTcell_reg[0][1]/P0001  , \core_c_psq_cntstk_cnts4x14_CNTcell_reg[0][2]/P0001  , \core_c_psq_cntstk_cnts4x14_CNTcell_reg[0][3]/P0001  , \core_c_psq_cntstk_cnts4x14_CNTcell_reg[0][4]/P0001  , \core_c_psq_cntstk_cnts4x14_CNTcell_reg[0][5]/P0001  , \core_c_psq_cntstk_cnts4x14_CNTcell_reg[0][6]/P0001  , \core_c_psq_cntstk_cnts4x14_CNTcell_reg[0][7]/P0001  , \core_c_psq_cntstk_cnts4x14_CNTcell_reg[0][8]/P0001  , \core_c_psq_cntstk_cnts4x14_CNTcell_reg[0][9]/P0001  , \core_c_psq_cntstk_cnts4x14_CNTcell_reg[1][0]/P0001  , \core_c_psq_cntstk_cnts4x14_CNTcell_reg[1][10]/P0001  , \core_c_psq_cntstk_cnts4x14_CNTcell_reg[1][11]/P0001  , \core_c_psq_cntstk_cnts4x14_CNTcell_reg[1][12]/P0001  , \core_c_psq_cntstk_cnts4x14_CNTcell_reg[1][13]/P0001  , \core_c_psq_cntstk_cnts4x14_CNTcell_reg[1][1]/P0001  , \core_c_psq_cntstk_cnts4x14_CNTcell_reg[1][2]/P0001  , \core_c_psq_cntstk_cnts4x14_CNTcell_reg[1][3]/P0001  , \core_c_psq_cntstk_cnts4x14_CNTcell_reg[1][4]/P0001  , \core_c_psq_cntstk_cnts4x14_CNTcell_reg[1][5]/P0001  , \core_c_psq_cntstk_cnts4x14_CNTcell_reg[1][6]/P0001  , \core_c_psq_cntstk_cnts4x14_CNTcell_reg[1][7]/P0001  , \core_c_psq_cntstk_cnts4x14_CNTcell_reg[1][8]/P0001  , \core_c_psq_cntstk_cnts4x14_CNTcell_reg[1][9]/P0001  , \core_c_psq_cntstk_cnts4x14_CNTcell_reg[2][0]/P0001  , \core_c_psq_cntstk_cnts4x14_CNTcell_reg[2][10]/P0001  , \core_c_psq_cntstk_cnts4x14_CNTcell_reg[2][11]/P0001  , \core_c_psq_cntstk_cnts4x14_CNTcell_reg[2][12]/P0001  , \core_c_psq_cntstk_cnts4x14_CNTcell_reg[2][13]/P0001  , \core_c_psq_cntstk_cnts4x14_CNTcell_reg[2][1]/P0001  , \core_c_psq_cntstk_cnts4x14_CNTcell_reg[2][2]/P0001  , \core_c_psq_cntstk_cnts4x14_CNTcell_reg[2][3]/P0001  , \core_c_psq_cntstk_cnts4x14_CNTcell_reg[2][4]/P0001  , \core_c_psq_cntstk_cnts4x14_CNTcell_reg[2][5]/P0001  , \core_c_psq_cntstk_cnts4x14_CNTcell_reg[2][6]/P0001  , \core_c_psq_cntstk_cnts4x14_CNTcell_reg[2][7]/P0001  , \core_c_psq_cntstk_cnts4x14_CNTcell_reg[2][8]/P0001  , \core_c_psq_cntstk_cnts4x14_CNTcell_reg[2][9]/P0001  , \core_c_psq_cntstk_cnts4x14_CNTcell_reg[3][0]/P0001  , \core_c_psq_cntstk_cnts4x14_CNTcell_reg[3][10]/P0001  , \core_c_psq_cntstk_cnts4x14_CNTcell_reg[3][11]/P0001  , \core_c_psq_cntstk_cnts4x14_CNTcell_reg[3][12]/P0001  , \core_c_psq_cntstk_cnts4x14_CNTcell_reg[3][13]/P0001  , \core_c_psq_cntstk_cnts4x14_CNTcell_reg[3][1]/P0001  , \core_c_psq_cntstk_cnts4x14_CNTcell_reg[3][2]/P0001  , \core_c_psq_cntstk_cnts4x14_CNTcell_reg[3][3]/P0001  , \core_c_psq_cntstk_cnts4x14_CNTcell_reg[3][4]/P0001  , \core_c_psq_cntstk_cnts4x14_CNTcell_reg[3][5]/P0001  , \core_c_psq_cntstk_cnts4x14_CNTcell_reg[3][6]/P0001  , \core_c_psq_cntstk_cnts4x14_CNTcell_reg[3][7]/P0001  , \core_c_psq_cntstk_cnts4x14_CNTcell_reg[3][8]/P0001  , \core_c_psq_cntstk_cnts4x14_CNTcell_reg[3][9]/P0001  , \core_c_psq_cntstk_ptr_reg[0]/NET0131  , \core_c_psq_cntstk_ptr_reg[1]/NET0131  , \core_c_psq_cntstk_ptr_reg[2]/NET0131  , \core_c_psq_irq0_de_IN_syn_reg/P0001  , \core_c_psq_irq0_de_OUT_reg/P0001  , \core_c_psq_irq1_de_IN_syn_reg/P0001  , \core_c_psq_irq1_de_OUT_reg/P0001  , \core_c_psq_irq2_de_IN_syn_reg/P0001  , \core_c_psq_irq2_de_OUT_reg/P0001  , \core_c_psq_irql0_de_IN_syn_reg/P0001  , \core_c_psq_irql0_de_OUT_reg/P0001  , \core_c_psq_irql1_de_IN_syn_reg/P0001  , \core_c_psq_irql1_de_OUT_reg/P0001  , \core_c_psq_lpstk_lps4x22_LPcell_reg[0][0]/P0001  , \core_c_psq_lpstk_lps4x22_LPcell_reg[0][10]/P0001  , \core_c_psq_lpstk_lps4x22_LPcell_reg[0][11]/P0001  , \core_c_psq_lpstk_lps4x22_LPcell_reg[0][12]/P0001  , \core_c_psq_lpstk_lps4x22_LPcell_reg[0][13]/P0001  , \core_c_psq_lpstk_lps4x22_LPcell_reg[0][14]/P0001  , \core_c_psq_lpstk_lps4x22_LPcell_reg[0][15]/P0001  , \core_c_psq_lpstk_lps4x22_LPcell_reg[0][16]/P0001  , \core_c_psq_lpstk_lps4x22_LPcell_reg[0][17]/P0001  , \core_c_psq_lpstk_lps4x22_LPcell_reg[0][18]/P0001  , \core_c_psq_lpstk_lps4x22_LPcell_reg[0][19]/P0001  , \core_c_psq_lpstk_lps4x22_LPcell_reg[0][1]/P0001  , \core_c_psq_lpstk_lps4x22_LPcell_reg[0][20]/P0001  , \core_c_psq_lpstk_lps4x22_LPcell_reg[0][21]/P0001  , \core_c_psq_lpstk_lps4x22_LPcell_reg[0][2]/P0001  , \core_c_psq_lpstk_lps4x22_LPcell_reg[0][3]/P0001  , \core_c_psq_lpstk_lps4x22_LPcell_reg[0][4]/P0001  , \core_c_psq_lpstk_lps4x22_LPcell_reg[0][5]/P0001  , \core_c_psq_lpstk_lps4x22_LPcell_reg[0][6]/P0001  , \core_c_psq_lpstk_lps4x22_LPcell_reg[0][7]/P0001  , \core_c_psq_lpstk_lps4x22_LPcell_reg[0][8]/P0001  , \core_c_psq_lpstk_lps4x22_LPcell_reg[0][9]/P0001  , \core_c_psq_lpstk_lps4x22_LPcell_reg[1][0]/P0001  , \core_c_psq_lpstk_lps4x22_LPcell_reg[1][10]/P0001  , \core_c_psq_lpstk_lps4x22_LPcell_reg[1][11]/P0001  , \core_c_psq_lpstk_lps4x22_LPcell_reg[1][12]/P0001  , \core_c_psq_lpstk_lps4x22_LPcell_reg[1][13]/P0001  , \core_c_psq_lpstk_lps4x22_LPcell_reg[1][14]/P0001  , \core_c_psq_lpstk_lps4x22_LPcell_reg[1][15]/P0001  , \core_c_psq_lpstk_lps4x22_LPcell_reg[1][16]/P0001  , \core_c_psq_lpstk_lps4x22_LPcell_reg[1][17]/P0001  , \core_c_psq_lpstk_lps4x22_LPcell_reg[1][18]/P0001  , \core_c_psq_lpstk_lps4x22_LPcell_reg[1][19]/P0001  , \core_c_psq_lpstk_lps4x22_LPcell_reg[1][1]/P0001  , \core_c_psq_lpstk_lps4x22_LPcell_reg[1][20]/P0001  , \core_c_psq_lpstk_lps4x22_LPcell_reg[1][21]/P0001  , \core_c_psq_lpstk_lps4x22_LPcell_reg[1][2]/P0001  , \core_c_psq_lpstk_lps4x22_LPcell_reg[1][3]/P0001  , \core_c_psq_lpstk_lps4x22_LPcell_reg[1][4]/P0001  , \core_c_psq_lpstk_lps4x22_LPcell_reg[1][5]/P0001  , \core_c_psq_lpstk_lps4x22_LPcell_reg[1][6]/P0001  , \core_c_psq_lpstk_lps4x22_LPcell_reg[1][7]/P0001  , \core_c_psq_lpstk_lps4x22_LPcell_reg[1][8]/P0001  , \core_c_psq_lpstk_lps4x22_LPcell_reg[1][9]/P0001  , \core_c_psq_lpstk_lps4x22_LPcell_reg[2][0]/P0001  , \core_c_psq_lpstk_lps4x22_LPcell_reg[2][10]/P0001  , \core_c_psq_lpstk_lps4x22_LPcell_reg[2][11]/P0001  , \core_c_psq_lpstk_lps4x22_LPcell_reg[2][12]/P0001  , \core_c_psq_lpstk_lps4x22_LPcell_reg[2][13]/P0001  , \core_c_psq_lpstk_lps4x22_LPcell_reg[2][14]/P0001  , \core_c_psq_lpstk_lps4x22_LPcell_reg[2][15]/P0001  , \core_c_psq_lpstk_lps4x22_LPcell_reg[2][16]/P0001  , \core_c_psq_lpstk_lps4x22_LPcell_reg[2][17]/P0001  , \core_c_psq_lpstk_lps4x22_LPcell_reg[2][18]/P0001  , \core_c_psq_lpstk_lps4x22_LPcell_reg[2][19]/P0001  , \core_c_psq_lpstk_lps4x22_LPcell_reg[2][1]/P0001  , \core_c_psq_lpstk_lps4x22_LPcell_reg[2][20]/P0001  , \core_c_psq_lpstk_lps4x22_LPcell_reg[2][21]/P0001  , \core_c_psq_lpstk_lps4x22_LPcell_reg[2][2]/P0001  , \core_c_psq_lpstk_lps4x22_LPcell_reg[2][3]/P0001  , \core_c_psq_lpstk_lps4x22_LPcell_reg[2][4]/P0001  , \core_c_psq_lpstk_lps4x22_LPcell_reg[2][5]/P0001  , \core_c_psq_lpstk_lps4x22_LPcell_reg[2][6]/P0001  , \core_c_psq_lpstk_lps4x22_LPcell_reg[2][7]/P0001  , \core_c_psq_lpstk_lps4x22_LPcell_reg[2][8]/P0001  , \core_c_psq_lpstk_lps4x22_LPcell_reg[2][9]/P0001  , \core_c_psq_lpstk_lps4x22_LPcell_reg[3][0]/P0001  , \core_c_psq_lpstk_lps4x22_LPcell_reg[3][10]/P0001  , \core_c_psq_lpstk_lps4x22_LPcell_reg[3][11]/P0001  , \core_c_psq_lpstk_lps4x22_LPcell_reg[3][12]/P0001  , \core_c_psq_lpstk_lps4x22_LPcell_reg[3][13]/P0001  , \core_c_psq_lpstk_lps4x22_LPcell_reg[3][14]/P0001  , \core_c_psq_lpstk_lps4x22_LPcell_reg[3][15]/P0001  , \core_c_psq_lpstk_lps4x22_LPcell_reg[3][16]/P0001  , \core_c_psq_lpstk_lps4x22_LPcell_reg[3][17]/P0001  , \core_c_psq_lpstk_lps4x22_LPcell_reg[3][18]/P0001  , \core_c_psq_lpstk_lps4x22_LPcell_reg[3][19]/P0001  , \core_c_psq_lpstk_lps4x22_LPcell_reg[3][1]/P0001  , \core_c_psq_lpstk_lps4x22_LPcell_reg[3][20]/P0001  , \core_c_psq_lpstk_lps4x22_LPcell_reg[3][21]/P0001  , \core_c_psq_lpstk_lps4x22_LPcell_reg[3][2]/P0001  , \core_c_psq_lpstk_lps4x22_LPcell_reg[3][3]/P0001  , \core_c_psq_lpstk_lps4x22_LPcell_reg[3][4]/P0001  , \core_c_psq_lpstk_lps4x22_LPcell_reg[3][5]/P0001  , \core_c_psq_lpstk_lps4x22_LPcell_reg[3][6]/P0001  , \core_c_psq_lpstk_lps4x22_LPcell_reg[3][7]/P0001  , \core_c_psq_lpstk_lps4x22_LPcell_reg[3][8]/P0001  , \core_c_psq_lpstk_lps4x22_LPcell_reg[3][9]/P0001  , \core_c_psq_lpstk_ptr_reg[0]/NET0131  , \core_c_psq_lpstk_ptr_reg[1]/NET0131  , \core_c_psq_lpstk_ptr_reg[2]/NET0131  , \core_c_psq_pcstk_cnts16x14_PCcell_reg[0][0]/P0001  , \core_c_psq_pcstk_cnts16x14_PCcell_reg[0][10]/P0001  , \core_c_psq_pcstk_cnts16x14_PCcell_reg[0][11]/P0001  , \core_c_psq_pcstk_cnts16x14_PCcell_reg[0][12]/P0001  , \core_c_psq_pcstk_cnts16x14_PCcell_reg[0][13]/P0001  , \core_c_psq_pcstk_cnts16x14_PCcell_reg[0][1]/P0001  , \core_c_psq_pcstk_cnts16x14_PCcell_reg[0][2]/P0001  , \core_c_psq_pcstk_cnts16x14_PCcell_reg[0][3]/P0001  , \core_c_psq_pcstk_cnts16x14_PCcell_reg[0][4]/P0001  , \core_c_psq_pcstk_cnts16x14_PCcell_reg[0][5]/P0001  , \core_c_psq_pcstk_cnts16x14_PCcell_reg[0][6]/P0001  , \core_c_psq_pcstk_cnts16x14_PCcell_reg[0][7]/P0001  , \core_c_psq_pcstk_cnts16x14_PCcell_reg[0][8]/P0001  , \core_c_psq_pcstk_cnts16x14_PCcell_reg[0][9]/P0001  , \core_c_psq_pcstk_cnts16x14_PCcell_reg[10][0]/P0001  , \core_c_psq_pcstk_cnts16x14_PCcell_reg[10][10]/P0001  , \core_c_psq_pcstk_cnts16x14_PCcell_reg[10][11]/P0001  , \core_c_psq_pcstk_cnts16x14_PCcell_reg[10][12]/P0001  , \core_c_psq_pcstk_cnts16x14_PCcell_reg[10][13]/P0001  , \core_c_psq_pcstk_cnts16x14_PCcell_reg[10][1]/P0001  , \core_c_psq_pcstk_cnts16x14_PCcell_reg[10][2]/P0001  , \core_c_psq_pcstk_cnts16x14_PCcell_reg[10][3]/P0001  , \core_c_psq_pcstk_cnts16x14_PCcell_reg[10][4]/P0001  , \core_c_psq_pcstk_cnts16x14_PCcell_reg[10][5]/P0001  , \core_c_psq_pcstk_cnts16x14_PCcell_reg[10][6]/P0001  , \core_c_psq_pcstk_cnts16x14_PCcell_reg[10][7]/P0001  , \core_c_psq_pcstk_cnts16x14_PCcell_reg[10][8]/P0001  , \core_c_psq_pcstk_cnts16x14_PCcell_reg[10][9]/P0001  , \core_c_psq_pcstk_cnts16x14_PCcell_reg[11][0]/P0001  , \core_c_psq_pcstk_cnts16x14_PCcell_reg[11][10]/P0001  , \core_c_psq_pcstk_cnts16x14_PCcell_reg[11][11]/P0001  , \core_c_psq_pcstk_cnts16x14_PCcell_reg[11][12]/P0001  , \core_c_psq_pcstk_cnts16x14_PCcell_reg[11][13]/P0001  , \core_c_psq_pcstk_cnts16x14_PCcell_reg[11][1]/P0001  , \core_c_psq_pcstk_cnts16x14_PCcell_reg[11][2]/P0001  , \core_c_psq_pcstk_cnts16x14_PCcell_reg[11][3]/P0001  , \core_c_psq_pcstk_cnts16x14_PCcell_reg[11][4]/P0001  , \core_c_psq_pcstk_cnts16x14_PCcell_reg[11][5]/P0001  , \core_c_psq_pcstk_cnts16x14_PCcell_reg[11][6]/P0001  , \core_c_psq_pcstk_cnts16x14_PCcell_reg[11][7]/P0001  , \core_c_psq_pcstk_cnts16x14_PCcell_reg[11][8]/P0001  , \core_c_psq_pcstk_cnts16x14_PCcell_reg[11][9]/P0001  , \core_c_psq_pcstk_cnts16x14_PCcell_reg[12][0]/P0001  , \core_c_psq_pcstk_cnts16x14_PCcell_reg[12][10]/P0001  , \core_c_psq_pcstk_cnts16x14_PCcell_reg[12][11]/P0001  , \core_c_psq_pcstk_cnts16x14_PCcell_reg[12][12]/P0001  , \core_c_psq_pcstk_cnts16x14_PCcell_reg[12][13]/P0001  , \core_c_psq_pcstk_cnts16x14_PCcell_reg[12][1]/P0001  , \core_c_psq_pcstk_cnts16x14_PCcell_reg[12][2]/P0001  , \core_c_psq_pcstk_cnts16x14_PCcell_reg[12][3]/P0001  , \core_c_psq_pcstk_cnts16x14_PCcell_reg[12][4]/P0001  , \core_c_psq_pcstk_cnts16x14_PCcell_reg[12][5]/P0001  , \core_c_psq_pcstk_cnts16x14_PCcell_reg[12][6]/P0001  , \core_c_psq_pcstk_cnts16x14_PCcell_reg[12][7]/P0001  , \core_c_psq_pcstk_cnts16x14_PCcell_reg[12][8]/P0001  , \core_c_psq_pcstk_cnts16x14_PCcell_reg[12][9]/P0001  , \core_c_psq_pcstk_cnts16x14_PCcell_reg[13][0]/P0001  , \core_c_psq_pcstk_cnts16x14_PCcell_reg[13][10]/P0001  , \core_c_psq_pcstk_cnts16x14_PCcell_reg[13][11]/P0001  , \core_c_psq_pcstk_cnts16x14_PCcell_reg[13][12]/P0001  , \core_c_psq_pcstk_cnts16x14_PCcell_reg[13][13]/P0001  , \core_c_psq_pcstk_cnts16x14_PCcell_reg[13][1]/P0001  , \core_c_psq_pcstk_cnts16x14_PCcell_reg[13][2]/P0001  , \core_c_psq_pcstk_cnts16x14_PCcell_reg[13][3]/P0001  , \core_c_psq_pcstk_cnts16x14_PCcell_reg[13][4]/P0001  , \core_c_psq_pcstk_cnts16x14_PCcell_reg[13][5]/P0001  , \core_c_psq_pcstk_cnts16x14_PCcell_reg[13][6]/P0001  , \core_c_psq_pcstk_cnts16x14_PCcell_reg[13][7]/P0001  , \core_c_psq_pcstk_cnts16x14_PCcell_reg[13][8]/P0001  , \core_c_psq_pcstk_cnts16x14_PCcell_reg[13][9]/P0001  , \core_c_psq_pcstk_cnts16x14_PCcell_reg[14][0]/P0001  , \core_c_psq_pcstk_cnts16x14_PCcell_reg[14][10]/P0001  , \core_c_psq_pcstk_cnts16x14_PCcell_reg[14][11]/P0001  , \core_c_psq_pcstk_cnts16x14_PCcell_reg[14][12]/P0001  , \core_c_psq_pcstk_cnts16x14_PCcell_reg[14][13]/P0001  , \core_c_psq_pcstk_cnts16x14_PCcell_reg[14][1]/P0001  , \core_c_psq_pcstk_cnts16x14_PCcell_reg[14][2]/P0001  , \core_c_psq_pcstk_cnts16x14_PCcell_reg[14][3]/P0001  , \core_c_psq_pcstk_cnts16x14_PCcell_reg[14][4]/P0001  , \core_c_psq_pcstk_cnts16x14_PCcell_reg[14][5]/P0001  , \core_c_psq_pcstk_cnts16x14_PCcell_reg[14][6]/P0001  , \core_c_psq_pcstk_cnts16x14_PCcell_reg[14][7]/P0001  , \core_c_psq_pcstk_cnts16x14_PCcell_reg[14][8]/P0001  , \core_c_psq_pcstk_cnts16x14_PCcell_reg[14][9]/P0001  , \core_c_psq_pcstk_cnts16x14_PCcell_reg[15][0]/P0001  , \core_c_psq_pcstk_cnts16x14_PCcell_reg[15][10]/P0001  , \core_c_psq_pcstk_cnts16x14_PCcell_reg[15][11]/P0001  , \core_c_psq_pcstk_cnts16x14_PCcell_reg[15][12]/P0001  , \core_c_psq_pcstk_cnts16x14_PCcell_reg[15][13]/P0001  , \core_c_psq_pcstk_cnts16x14_PCcell_reg[15][1]/P0001  , \core_c_psq_pcstk_cnts16x14_PCcell_reg[15][2]/P0001  , \core_c_psq_pcstk_cnts16x14_PCcell_reg[15][3]/P0001  , \core_c_psq_pcstk_cnts16x14_PCcell_reg[15][4]/P0001  , \core_c_psq_pcstk_cnts16x14_PCcell_reg[15][5]/P0001  , \core_c_psq_pcstk_cnts16x14_PCcell_reg[15][6]/P0001  , \core_c_psq_pcstk_cnts16x14_PCcell_reg[15][7]/P0001  , \core_c_psq_pcstk_cnts16x14_PCcell_reg[15][8]/P0001  , \core_c_psq_pcstk_cnts16x14_PCcell_reg[15][9]/P0001  , \core_c_psq_pcstk_cnts16x14_PCcell_reg[1][0]/P0001  , \core_c_psq_pcstk_cnts16x14_PCcell_reg[1][10]/P0001  , \core_c_psq_pcstk_cnts16x14_PCcell_reg[1][11]/P0001  , \core_c_psq_pcstk_cnts16x14_PCcell_reg[1][12]/P0001  , \core_c_psq_pcstk_cnts16x14_PCcell_reg[1][13]/P0001  , \core_c_psq_pcstk_cnts16x14_PCcell_reg[1][1]/P0001  , \core_c_psq_pcstk_cnts16x14_PCcell_reg[1][2]/P0001  , \core_c_psq_pcstk_cnts16x14_PCcell_reg[1][3]/P0001  , \core_c_psq_pcstk_cnts16x14_PCcell_reg[1][4]/P0001  , \core_c_psq_pcstk_cnts16x14_PCcell_reg[1][5]/P0001  , \core_c_psq_pcstk_cnts16x14_PCcell_reg[1][6]/P0001  , \core_c_psq_pcstk_cnts16x14_PCcell_reg[1][7]/P0001  , \core_c_psq_pcstk_cnts16x14_PCcell_reg[1][8]/P0001  , \core_c_psq_pcstk_cnts16x14_PCcell_reg[1][9]/P0001  , \core_c_psq_pcstk_cnts16x14_PCcell_reg[2][0]/P0001  , \core_c_psq_pcstk_cnts16x14_PCcell_reg[2][10]/P0001  , \core_c_psq_pcstk_cnts16x14_PCcell_reg[2][11]/P0001  , \core_c_psq_pcstk_cnts16x14_PCcell_reg[2][12]/P0001  , \core_c_psq_pcstk_cnts16x14_PCcell_reg[2][13]/P0001  , \core_c_psq_pcstk_cnts16x14_PCcell_reg[2][1]/P0001  , \core_c_psq_pcstk_cnts16x14_PCcell_reg[2][2]/P0001  , \core_c_psq_pcstk_cnts16x14_PCcell_reg[2][3]/P0001  , \core_c_psq_pcstk_cnts16x14_PCcell_reg[2][4]/P0001  , \core_c_psq_pcstk_cnts16x14_PCcell_reg[2][5]/P0001  , \core_c_psq_pcstk_cnts16x14_PCcell_reg[2][6]/P0001  , \core_c_psq_pcstk_cnts16x14_PCcell_reg[2][7]/P0001  , \core_c_psq_pcstk_cnts16x14_PCcell_reg[2][8]/P0001  , \core_c_psq_pcstk_cnts16x14_PCcell_reg[2][9]/P0001  , \core_c_psq_pcstk_cnts16x14_PCcell_reg[3][0]/P0001  , \core_c_psq_pcstk_cnts16x14_PCcell_reg[3][10]/P0001  , \core_c_psq_pcstk_cnts16x14_PCcell_reg[3][11]/P0001  , \core_c_psq_pcstk_cnts16x14_PCcell_reg[3][12]/P0001  , \core_c_psq_pcstk_cnts16x14_PCcell_reg[3][13]/P0001  , \core_c_psq_pcstk_cnts16x14_PCcell_reg[3][1]/P0001  , \core_c_psq_pcstk_cnts16x14_PCcell_reg[3][2]/P0001  , \core_c_psq_pcstk_cnts16x14_PCcell_reg[3][3]/P0001  , \core_c_psq_pcstk_cnts16x14_PCcell_reg[3][4]/P0001  , \core_c_psq_pcstk_cnts16x14_PCcell_reg[3][5]/P0001  , \core_c_psq_pcstk_cnts16x14_PCcell_reg[3][6]/P0001  , \core_c_psq_pcstk_cnts16x14_PCcell_reg[3][7]/P0001  , \core_c_psq_pcstk_cnts16x14_PCcell_reg[3][8]/P0001  , \core_c_psq_pcstk_cnts16x14_PCcell_reg[3][9]/P0001  , \core_c_psq_pcstk_cnts16x14_PCcell_reg[4][0]/P0001  , \core_c_psq_pcstk_cnts16x14_PCcell_reg[4][10]/P0001  , \core_c_psq_pcstk_cnts16x14_PCcell_reg[4][11]/P0001  , \core_c_psq_pcstk_cnts16x14_PCcell_reg[4][12]/P0001  , \core_c_psq_pcstk_cnts16x14_PCcell_reg[4][13]/P0001  , \core_c_psq_pcstk_cnts16x14_PCcell_reg[4][1]/P0001  , \core_c_psq_pcstk_cnts16x14_PCcell_reg[4][2]/P0001  , \core_c_psq_pcstk_cnts16x14_PCcell_reg[4][3]/P0001  , \core_c_psq_pcstk_cnts16x14_PCcell_reg[4][4]/P0001  , \core_c_psq_pcstk_cnts16x14_PCcell_reg[4][5]/P0001  , \core_c_psq_pcstk_cnts16x14_PCcell_reg[4][6]/P0001  , \core_c_psq_pcstk_cnts16x14_PCcell_reg[4][7]/P0001  , \core_c_psq_pcstk_cnts16x14_PCcell_reg[4][8]/P0001  , \core_c_psq_pcstk_cnts16x14_PCcell_reg[4][9]/P0001  , \core_c_psq_pcstk_cnts16x14_PCcell_reg[5][0]/P0001  , \core_c_psq_pcstk_cnts16x14_PCcell_reg[5][10]/P0001  , \core_c_psq_pcstk_cnts16x14_PCcell_reg[5][11]/P0001  , \core_c_psq_pcstk_cnts16x14_PCcell_reg[5][12]/P0001  , \core_c_psq_pcstk_cnts16x14_PCcell_reg[5][13]/P0001  , \core_c_psq_pcstk_cnts16x14_PCcell_reg[5][1]/P0001  , \core_c_psq_pcstk_cnts16x14_PCcell_reg[5][2]/P0001  , \core_c_psq_pcstk_cnts16x14_PCcell_reg[5][3]/P0001  , \core_c_psq_pcstk_cnts16x14_PCcell_reg[5][4]/P0001  , \core_c_psq_pcstk_cnts16x14_PCcell_reg[5][5]/P0001  , \core_c_psq_pcstk_cnts16x14_PCcell_reg[5][6]/P0001  , \core_c_psq_pcstk_cnts16x14_PCcell_reg[5][7]/P0001  , \core_c_psq_pcstk_cnts16x14_PCcell_reg[5][8]/P0001  , \core_c_psq_pcstk_cnts16x14_PCcell_reg[5][9]/P0001  , \core_c_psq_pcstk_cnts16x14_PCcell_reg[6][0]/P0001  , \core_c_psq_pcstk_cnts16x14_PCcell_reg[6][10]/P0001  , \core_c_psq_pcstk_cnts16x14_PCcell_reg[6][11]/P0001  , \core_c_psq_pcstk_cnts16x14_PCcell_reg[6][12]/P0001  , \core_c_psq_pcstk_cnts16x14_PCcell_reg[6][13]/P0001  , \core_c_psq_pcstk_cnts16x14_PCcell_reg[6][1]/P0001  , \core_c_psq_pcstk_cnts16x14_PCcell_reg[6][2]/P0001  , \core_c_psq_pcstk_cnts16x14_PCcell_reg[6][3]/P0001  , \core_c_psq_pcstk_cnts16x14_PCcell_reg[6][4]/P0001  , \core_c_psq_pcstk_cnts16x14_PCcell_reg[6][5]/P0001  , \core_c_psq_pcstk_cnts16x14_PCcell_reg[6][6]/P0001  , \core_c_psq_pcstk_cnts16x14_PCcell_reg[6][7]/P0001  , \core_c_psq_pcstk_cnts16x14_PCcell_reg[6][8]/P0001  , \core_c_psq_pcstk_cnts16x14_PCcell_reg[6][9]/P0001  , \core_c_psq_pcstk_cnts16x14_PCcell_reg[7][0]/P0001  , \core_c_psq_pcstk_cnts16x14_PCcell_reg[7][10]/P0001  , \core_c_psq_pcstk_cnts16x14_PCcell_reg[7][11]/P0001  , \core_c_psq_pcstk_cnts16x14_PCcell_reg[7][12]/P0001  , \core_c_psq_pcstk_cnts16x14_PCcell_reg[7][13]/P0001  , \core_c_psq_pcstk_cnts16x14_PCcell_reg[7][1]/P0001  , \core_c_psq_pcstk_cnts16x14_PCcell_reg[7][2]/P0001  , \core_c_psq_pcstk_cnts16x14_PCcell_reg[7][3]/P0001  , \core_c_psq_pcstk_cnts16x14_PCcell_reg[7][4]/P0001  , \core_c_psq_pcstk_cnts16x14_PCcell_reg[7][5]/P0001  , \core_c_psq_pcstk_cnts16x14_PCcell_reg[7][6]/P0001  , \core_c_psq_pcstk_cnts16x14_PCcell_reg[7][7]/P0001  , \core_c_psq_pcstk_cnts16x14_PCcell_reg[7][8]/P0001  , \core_c_psq_pcstk_cnts16x14_PCcell_reg[7][9]/P0001  , \core_c_psq_pcstk_cnts16x14_PCcell_reg[8][0]/P0001  , \core_c_psq_pcstk_cnts16x14_PCcell_reg[8][10]/P0001  , \core_c_psq_pcstk_cnts16x14_PCcell_reg[8][11]/P0001  , \core_c_psq_pcstk_cnts16x14_PCcell_reg[8][12]/P0001  , \core_c_psq_pcstk_cnts16x14_PCcell_reg[8][13]/P0001  , \core_c_psq_pcstk_cnts16x14_PCcell_reg[8][1]/P0001  , \core_c_psq_pcstk_cnts16x14_PCcell_reg[8][2]/P0001  , \core_c_psq_pcstk_cnts16x14_PCcell_reg[8][3]/P0001  , \core_c_psq_pcstk_cnts16x14_PCcell_reg[8][4]/P0001  , \core_c_psq_pcstk_cnts16x14_PCcell_reg[8][5]/P0001  , \core_c_psq_pcstk_cnts16x14_PCcell_reg[8][6]/P0001  , \core_c_psq_pcstk_cnts16x14_PCcell_reg[8][7]/P0001  , \core_c_psq_pcstk_cnts16x14_PCcell_reg[8][8]/P0001  , \core_c_psq_pcstk_cnts16x14_PCcell_reg[8][9]/P0001  , \core_c_psq_pcstk_cnts16x14_PCcell_reg[9][0]/P0001  , \core_c_psq_pcstk_cnts16x14_PCcell_reg[9][10]/P0001  , \core_c_psq_pcstk_cnts16x14_PCcell_reg[9][11]/P0001  , \core_c_psq_pcstk_cnts16x14_PCcell_reg[9][12]/P0001  , \core_c_psq_pcstk_cnts16x14_PCcell_reg[9][13]/P0001  , \core_c_psq_pcstk_cnts16x14_PCcell_reg[9][1]/P0001  , \core_c_psq_pcstk_cnts16x14_PCcell_reg[9][2]/P0001  , \core_c_psq_pcstk_cnts16x14_PCcell_reg[9][3]/P0001  , \core_c_psq_pcstk_cnts16x14_PCcell_reg[9][4]/P0001  , \core_c_psq_pcstk_cnts16x14_PCcell_reg[9][5]/P0001  , \core_c_psq_pcstk_cnts16x14_PCcell_reg[9][6]/P0001  , \core_c_psq_pcstk_cnts16x14_PCcell_reg[9][7]/P0001  , \core_c_psq_pcstk_cnts16x14_PCcell_reg[9][8]/P0001  , \core_c_psq_pcstk_cnts16x14_PCcell_reg[9][9]/P0001  , \core_c_psq_pcstk_ptr_reg[0]/NET0131  , \core_c_psq_pcstk_ptr_reg[1]/NET0131  , \core_c_psq_pcstk_ptr_reg[2]/NET0131  , \core_c_psq_pcstk_ptr_reg[3]/NET0131  , \core_c_psq_pcstk_ptr_reg[4]/NET0131  , \core_c_psq_ststk_ptr_reg[0]/NET0131  , \core_c_psq_ststk_ptr_reg[1]/NET0131  , \core_c_psq_ststk_ptr_reg[2]/NET0131  , \core_c_psq_ststk_sts7x23_STcell_reg[0][0]/P0001  , \core_c_psq_ststk_sts7x23_STcell_reg[0][10]/P0001  , \core_c_psq_ststk_sts7x23_STcell_reg[0][11]/P0001  , \core_c_psq_ststk_sts7x23_STcell_reg[0][12]/P0001  , \core_c_psq_ststk_sts7x23_STcell_reg[0][13]/P0001  , \core_c_psq_ststk_sts7x23_STcell_reg[0][14]/P0001  , \core_c_psq_ststk_sts7x23_STcell_reg[0][15]/P0001  , \core_c_psq_ststk_sts7x23_STcell_reg[0][16]/P0001  , \core_c_psq_ststk_sts7x23_STcell_reg[0][17]/P0001  , \core_c_psq_ststk_sts7x23_STcell_reg[0][18]/P0001  , \core_c_psq_ststk_sts7x23_STcell_reg[0][19]/P0001  , \core_c_psq_ststk_sts7x23_STcell_reg[0][1]/P0001  , \core_c_psq_ststk_sts7x23_STcell_reg[0][20]/P0001  , \core_c_psq_ststk_sts7x23_STcell_reg[0][21]/P0001  , \core_c_psq_ststk_sts7x23_STcell_reg[0][22]/P0001  , \core_c_psq_ststk_sts7x23_STcell_reg[0][23]/P0001  , \core_c_psq_ststk_sts7x23_STcell_reg[0][24]/P0001  , \core_c_psq_ststk_sts7x23_STcell_reg[0][2]/P0001  , \core_c_psq_ststk_sts7x23_STcell_reg[0][3]/P0001  , \core_c_psq_ststk_sts7x23_STcell_reg[0][4]/P0001  , \core_c_psq_ststk_sts7x23_STcell_reg[0][5]/P0001  , \core_c_psq_ststk_sts7x23_STcell_reg[0][6]/P0001  , \core_c_psq_ststk_sts7x23_STcell_reg[0][7]/P0001  , \core_c_psq_ststk_sts7x23_STcell_reg[0][8]/P0001  , \core_c_psq_ststk_sts7x23_STcell_reg[0][9]/P0001  , \core_c_psq_ststk_sts7x23_STcell_reg[1][0]/P0001  , \core_c_psq_ststk_sts7x23_STcell_reg[1][10]/P0001  , \core_c_psq_ststk_sts7x23_STcell_reg[1][11]/P0001  , \core_c_psq_ststk_sts7x23_STcell_reg[1][12]/P0001  , \core_c_psq_ststk_sts7x23_STcell_reg[1][13]/P0001  , \core_c_psq_ststk_sts7x23_STcell_reg[1][14]/P0001  , \core_c_psq_ststk_sts7x23_STcell_reg[1][15]/P0001  , \core_c_psq_ststk_sts7x23_STcell_reg[1][16]/P0001  , \core_c_psq_ststk_sts7x23_STcell_reg[1][17]/P0001  , \core_c_psq_ststk_sts7x23_STcell_reg[1][18]/P0001  , \core_c_psq_ststk_sts7x23_STcell_reg[1][19]/P0001  , \core_c_psq_ststk_sts7x23_STcell_reg[1][1]/P0001  , \core_c_psq_ststk_sts7x23_STcell_reg[1][20]/P0001  , \core_c_psq_ststk_sts7x23_STcell_reg[1][21]/P0001  , \core_c_psq_ststk_sts7x23_STcell_reg[1][22]/P0001  , \core_c_psq_ststk_sts7x23_STcell_reg[1][23]/P0001  , \core_c_psq_ststk_sts7x23_STcell_reg[1][24]/P0001  , \core_c_psq_ststk_sts7x23_STcell_reg[1][2]/P0001  , \core_c_psq_ststk_sts7x23_STcell_reg[1][3]/P0001  , \core_c_psq_ststk_sts7x23_STcell_reg[1][4]/P0001  , \core_c_psq_ststk_sts7x23_STcell_reg[1][5]/P0001  , \core_c_psq_ststk_sts7x23_STcell_reg[1][6]/P0001  , \core_c_psq_ststk_sts7x23_STcell_reg[1][7]/P0001  , \core_c_psq_ststk_sts7x23_STcell_reg[1][8]/P0001  , \core_c_psq_ststk_sts7x23_STcell_reg[1][9]/P0001  , \core_c_psq_ststk_sts7x23_STcell_reg[2][0]/P0001  , \core_c_psq_ststk_sts7x23_STcell_reg[2][10]/P0001  , \core_c_psq_ststk_sts7x23_STcell_reg[2][11]/P0001  , \core_c_psq_ststk_sts7x23_STcell_reg[2][12]/P0001  , \core_c_psq_ststk_sts7x23_STcell_reg[2][13]/P0001  , \core_c_psq_ststk_sts7x23_STcell_reg[2][14]/P0001  , \core_c_psq_ststk_sts7x23_STcell_reg[2][15]/P0001  , \core_c_psq_ststk_sts7x23_STcell_reg[2][16]/P0001  , \core_c_psq_ststk_sts7x23_STcell_reg[2][17]/P0001  , \core_c_psq_ststk_sts7x23_STcell_reg[2][18]/P0001  , \core_c_psq_ststk_sts7x23_STcell_reg[2][19]/P0001  , \core_c_psq_ststk_sts7x23_STcell_reg[2][1]/P0001  , \core_c_psq_ststk_sts7x23_STcell_reg[2][20]/P0001  , \core_c_psq_ststk_sts7x23_STcell_reg[2][21]/P0001  , \core_c_psq_ststk_sts7x23_STcell_reg[2][22]/P0001  , \core_c_psq_ststk_sts7x23_STcell_reg[2][23]/P0001  , \core_c_psq_ststk_sts7x23_STcell_reg[2][24]/P0001  , \core_c_psq_ststk_sts7x23_STcell_reg[2][2]/P0001  , \core_c_psq_ststk_sts7x23_STcell_reg[2][3]/P0001  , \core_c_psq_ststk_sts7x23_STcell_reg[2][4]/P0001  , \core_c_psq_ststk_sts7x23_STcell_reg[2][5]/P0001  , \core_c_psq_ststk_sts7x23_STcell_reg[2][6]/P0001  , \core_c_psq_ststk_sts7x23_STcell_reg[2][7]/P0001  , \core_c_psq_ststk_sts7x23_STcell_reg[2][8]/P0001  , \core_c_psq_ststk_sts7x23_STcell_reg[2][9]/P0001  , \core_c_psq_ststk_sts7x23_STcell_reg[3][0]/P0001  , \core_c_psq_ststk_sts7x23_STcell_reg[3][10]/P0001  , \core_c_psq_ststk_sts7x23_STcell_reg[3][11]/P0001  , \core_c_psq_ststk_sts7x23_STcell_reg[3][12]/P0001  , \core_c_psq_ststk_sts7x23_STcell_reg[3][13]/P0001  , \core_c_psq_ststk_sts7x23_STcell_reg[3][14]/P0001  , \core_c_psq_ststk_sts7x23_STcell_reg[3][15]/P0001  , \core_c_psq_ststk_sts7x23_STcell_reg[3][16]/P0001  , \core_c_psq_ststk_sts7x23_STcell_reg[3][17]/P0001  , \core_c_psq_ststk_sts7x23_STcell_reg[3][18]/P0001  , \core_c_psq_ststk_sts7x23_STcell_reg[3][19]/P0001  , \core_c_psq_ststk_sts7x23_STcell_reg[3][1]/P0001  , \core_c_psq_ststk_sts7x23_STcell_reg[3][20]/P0001  , \core_c_psq_ststk_sts7x23_STcell_reg[3][21]/P0001  , \core_c_psq_ststk_sts7x23_STcell_reg[3][22]/P0001  , \core_c_psq_ststk_sts7x23_STcell_reg[3][23]/P0001  , \core_c_psq_ststk_sts7x23_STcell_reg[3][24]/P0001  , \core_c_psq_ststk_sts7x23_STcell_reg[3][2]/P0001  , \core_c_psq_ststk_sts7x23_STcell_reg[3][3]/P0001  , \core_c_psq_ststk_sts7x23_STcell_reg[3][4]/P0001  , \core_c_psq_ststk_sts7x23_STcell_reg[3][5]/P0001  , \core_c_psq_ststk_sts7x23_STcell_reg[3][6]/P0001  , \core_c_psq_ststk_sts7x23_STcell_reg[3][7]/P0001  , \core_c_psq_ststk_sts7x23_STcell_reg[3][8]/P0001  , \core_c_psq_ststk_sts7x23_STcell_reg[3][9]/P0001  , \core_c_psq_ststk_sts7x23_STcell_reg[4][0]/P0001  , \core_c_psq_ststk_sts7x23_STcell_reg[4][10]/P0001  , \core_c_psq_ststk_sts7x23_STcell_reg[4][11]/P0001  , \core_c_psq_ststk_sts7x23_STcell_reg[4][12]/P0001  , \core_c_psq_ststk_sts7x23_STcell_reg[4][13]/P0001  , \core_c_psq_ststk_sts7x23_STcell_reg[4][14]/P0001  , \core_c_psq_ststk_sts7x23_STcell_reg[4][15]/P0001  , \core_c_psq_ststk_sts7x23_STcell_reg[4][16]/P0001  , \core_c_psq_ststk_sts7x23_STcell_reg[4][17]/P0001  , \core_c_psq_ststk_sts7x23_STcell_reg[4][18]/P0001  , \core_c_psq_ststk_sts7x23_STcell_reg[4][19]/P0001  , \core_c_psq_ststk_sts7x23_STcell_reg[4][1]/P0001  , \core_c_psq_ststk_sts7x23_STcell_reg[4][20]/P0001  , \core_c_psq_ststk_sts7x23_STcell_reg[4][21]/P0001  , \core_c_psq_ststk_sts7x23_STcell_reg[4][22]/P0001  , \core_c_psq_ststk_sts7x23_STcell_reg[4][23]/P0001  , \core_c_psq_ststk_sts7x23_STcell_reg[4][24]/P0001  , \core_c_psq_ststk_sts7x23_STcell_reg[4][2]/P0001  , \core_c_psq_ststk_sts7x23_STcell_reg[4][3]/P0001  , \core_c_psq_ststk_sts7x23_STcell_reg[4][4]/P0001  , \core_c_psq_ststk_sts7x23_STcell_reg[4][5]/P0001  , \core_c_psq_ststk_sts7x23_STcell_reg[4][6]/P0001  , \core_c_psq_ststk_sts7x23_STcell_reg[4][7]/P0001  , \core_c_psq_ststk_sts7x23_STcell_reg[4][8]/P0001  , \core_c_psq_ststk_sts7x23_STcell_reg[4][9]/P0001  , \core_c_psq_ststk_sts7x23_STcell_reg[5][0]/P0001  , \core_c_psq_ststk_sts7x23_STcell_reg[5][10]/P0001  , \core_c_psq_ststk_sts7x23_STcell_reg[5][11]/P0001  , \core_c_psq_ststk_sts7x23_STcell_reg[5][12]/P0001  , \core_c_psq_ststk_sts7x23_STcell_reg[5][13]/P0001  , \core_c_psq_ststk_sts7x23_STcell_reg[5][14]/P0001  , \core_c_psq_ststk_sts7x23_STcell_reg[5][15]/P0001  , \core_c_psq_ststk_sts7x23_STcell_reg[5][16]/P0001  , \core_c_psq_ststk_sts7x23_STcell_reg[5][17]/P0001  , \core_c_psq_ststk_sts7x23_STcell_reg[5][18]/P0001  , \core_c_psq_ststk_sts7x23_STcell_reg[5][19]/P0001  , \core_c_psq_ststk_sts7x23_STcell_reg[5][1]/P0001  , \core_c_psq_ststk_sts7x23_STcell_reg[5][20]/P0001  , \core_c_psq_ststk_sts7x23_STcell_reg[5][21]/P0001  , \core_c_psq_ststk_sts7x23_STcell_reg[5][22]/P0001  , \core_c_psq_ststk_sts7x23_STcell_reg[5][23]/P0001  , \core_c_psq_ststk_sts7x23_STcell_reg[5][24]/P0001  , \core_c_psq_ststk_sts7x23_STcell_reg[5][2]/P0001  , \core_c_psq_ststk_sts7x23_STcell_reg[5][3]/P0001  , \core_c_psq_ststk_sts7x23_STcell_reg[5][4]/P0001  , \core_c_psq_ststk_sts7x23_STcell_reg[5][5]/P0001  , \core_c_psq_ststk_sts7x23_STcell_reg[5][6]/P0001  , \core_c_psq_ststk_sts7x23_STcell_reg[5][7]/P0001  , \core_c_psq_ststk_sts7x23_STcell_reg[5][8]/P0001  , \core_c_psq_ststk_sts7x23_STcell_reg[5][9]/P0001  , \core_c_psq_ststk_sts7x23_STcell_reg[6][0]/P0001  , \core_c_psq_ststk_sts7x23_STcell_reg[6][10]/P0001  , \core_c_psq_ststk_sts7x23_STcell_reg[6][11]/P0001  , \core_c_psq_ststk_sts7x23_STcell_reg[6][12]/P0001  , \core_c_psq_ststk_sts7x23_STcell_reg[6][13]/P0001  , \core_c_psq_ststk_sts7x23_STcell_reg[6][14]/P0001  , \core_c_psq_ststk_sts7x23_STcell_reg[6][15]/P0001  , \core_c_psq_ststk_sts7x23_STcell_reg[6][16]/P0001  , \core_c_psq_ststk_sts7x23_STcell_reg[6][17]/P0001  , \core_c_psq_ststk_sts7x23_STcell_reg[6][18]/P0001  , \core_c_psq_ststk_sts7x23_STcell_reg[6][19]/P0001  , \core_c_psq_ststk_sts7x23_STcell_reg[6][1]/P0001  , \core_c_psq_ststk_sts7x23_STcell_reg[6][20]/P0001  , \core_c_psq_ststk_sts7x23_STcell_reg[6][21]/P0001  , \core_c_psq_ststk_sts7x23_STcell_reg[6][22]/P0001  , \core_c_psq_ststk_sts7x23_STcell_reg[6][23]/P0001  , \core_c_psq_ststk_sts7x23_STcell_reg[6][24]/P0001  , \core_c_psq_ststk_sts7x23_STcell_reg[6][2]/P0001  , \core_c_psq_ststk_sts7x23_STcell_reg[6][3]/P0001  , \core_c_psq_ststk_sts7x23_STcell_reg[6][4]/P0001  , \core_c_psq_ststk_sts7x23_STcell_reg[6][5]/P0001  , \core_c_psq_ststk_sts7x23_STcell_reg[6][6]/P0001  , \core_c_psq_ststk_sts7x23_STcell_reg[6][7]/P0001  , \core_c_psq_ststk_sts7x23_STcell_reg[6][8]/P0001  , \core_c_psq_ststk_sts7x23_STcell_reg[6][9]/P0001  , \core_dag_ilm1reg_DMA_pi_DO_reg[0]/NET0131  , \core_dag_ilm1reg_DMA_pi_DO_reg[10]/NET0131  , \core_dag_ilm1reg_DMA_pi_DO_reg[11]/NET0131  , \core_dag_ilm1reg_DMA_pi_DO_reg[12]/NET0131  , \core_dag_ilm1reg_DMA_pi_DO_reg[13]/NET0131  , \core_dag_ilm1reg_DMA_pi_DO_reg[1]/NET0131  , \core_dag_ilm1reg_DMA_pi_DO_reg[2]/NET0131  , \core_dag_ilm1reg_DMA_pi_DO_reg[3]/NET0131  , \core_dag_ilm1reg_DMA_pi_DO_reg[4]/NET0131  , \core_dag_ilm1reg_DMA_pi_DO_reg[5]/NET0131  , \core_dag_ilm1reg_DMA_pi_DO_reg[6]/NET0131  , \core_dag_ilm1reg_DMA_pi_DO_reg[7]/NET0131  , \core_dag_ilm1reg_DMA_pi_DO_reg[8]/NET0131  , \core_dag_ilm1reg_DMA_pi_DO_reg[9]/NET0131  , \core_dag_ilm1reg_I0_we_DO_reg[0]/NET0131  , \core_dag_ilm1reg_I0_we_DO_reg[10]/NET0131  , \core_dag_ilm1reg_I0_we_DO_reg[11]/NET0131  , \core_dag_ilm1reg_I0_we_DO_reg[12]/NET0131  , \core_dag_ilm1reg_I0_we_DO_reg[13]/NET0131  , \core_dag_ilm1reg_I0_we_DO_reg[1]/NET0131  , \core_dag_ilm1reg_I0_we_DO_reg[2]/NET0131  , \core_dag_ilm1reg_I0_we_DO_reg[3]/NET0131  , \core_dag_ilm1reg_I0_we_DO_reg[4]/NET0131  , \core_dag_ilm1reg_I0_we_DO_reg[5]/NET0131  , \core_dag_ilm1reg_I0_we_DO_reg[6]/NET0131  , \core_dag_ilm1reg_I0_we_DO_reg[7]/NET0131  , \core_dag_ilm1reg_I0_we_DO_reg[8]/NET0131  , \core_dag_ilm1reg_I0_we_DO_reg[9]/NET0131  , \core_dag_ilm1reg_I1_we_DO_reg[0]/NET0131  , \core_dag_ilm1reg_I1_we_DO_reg[10]/NET0131  , \core_dag_ilm1reg_I1_we_DO_reg[11]/NET0131  , \core_dag_ilm1reg_I1_we_DO_reg[12]/NET0131  , \core_dag_ilm1reg_I1_we_DO_reg[13]/NET0131  , \core_dag_ilm1reg_I1_we_DO_reg[1]/NET0131  , \core_dag_ilm1reg_I1_we_DO_reg[2]/NET0131  , \core_dag_ilm1reg_I1_we_DO_reg[3]/NET0131  , \core_dag_ilm1reg_I1_we_DO_reg[4]/NET0131  , \core_dag_ilm1reg_I1_we_DO_reg[5]/NET0131  , \core_dag_ilm1reg_I1_we_DO_reg[6]/NET0131  , \core_dag_ilm1reg_I1_we_DO_reg[7]/NET0131  , \core_dag_ilm1reg_I1_we_DO_reg[8]/NET0131  , \core_dag_ilm1reg_I1_we_DO_reg[9]/NET0131  , \core_dag_ilm1reg_I2_we_DO_reg[0]/NET0131  , \core_dag_ilm1reg_I2_we_DO_reg[10]/NET0131  , \core_dag_ilm1reg_I2_we_DO_reg[11]/NET0131  , \core_dag_ilm1reg_I2_we_DO_reg[12]/NET0131  , \core_dag_ilm1reg_I2_we_DO_reg[13]/NET0131  , \core_dag_ilm1reg_I2_we_DO_reg[1]/NET0131  , \core_dag_ilm1reg_I2_we_DO_reg[2]/NET0131  , \core_dag_ilm1reg_I2_we_DO_reg[3]/NET0131  , \core_dag_ilm1reg_I2_we_DO_reg[4]/NET0131  , \core_dag_ilm1reg_I2_we_DO_reg[5]/NET0131  , \core_dag_ilm1reg_I2_we_DO_reg[6]/NET0131  , \core_dag_ilm1reg_I2_we_DO_reg[7]/NET0131  , \core_dag_ilm1reg_I2_we_DO_reg[8]/NET0131  , \core_dag_ilm1reg_I2_we_DO_reg[9]/NET0131  , \core_dag_ilm1reg_I3_we_DO_reg[0]/NET0131  , \core_dag_ilm1reg_I3_we_DO_reg[10]/NET0131  , \core_dag_ilm1reg_I3_we_DO_reg[11]/NET0131  , \core_dag_ilm1reg_I3_we_DO_reg[12]/NET0131  , \core_dag_ilm1reg_I3_we_DO_reg[13]/NET0131  , \core_dag_ilm1reg_I3_we_DO_reg[1]/NET0131  , \core_dag_ilm1reg_I3_we_DO_reg[2]/NET0131  , \core_dag_ilm1reg_I3_we_DO_reg[3]/NET0131  , \core_dag_ilm1reg_I3_we_DO_reg[4]/NET0131  , \core_dag_ilm1reg_I3_we_DO_reg[5]/NET0131  , \core_dag_ilm1reg_I3_we_DO_reg[6]/NET0131  , \core_dag_ilm1reg_I3_we_DO_reg[7]/NET0131  , \core_dag_ilm1reg_I3_we_DO_reg[8]/NET0131  , \core_dag_ilm1reg_I3_we_DO_reg[9]/NET0131  , \core_dag_ilm1reg_I_reg[0]/NET0131  , \core_dag_ilm1reg_I_reg[10]/NET0131  , \core_dag_ilm1reg_I_reg[11]/NET0131  , \core_dag_ilm1reg_I_reg[12]/NET0131  , \core_dag_ilm1reg_I_reg[13]/NET0131  , \core_dag_ilm1reg_I_reg[1]/NET0131  , \core_dag_ilm1reg_I_reg[2]/NET0131  , \core_dag_ilm1reg_I_reg[3]/NET0131  , \core_dag_ilm1reg_I_reg[4]/NET0131  , \core_dag_ilm1reg_I_reg[5]/NET0131  , \core_dag_ilm1reg_I_reg[6]/NET0131  , \core_dag_ilm1reg_I_reg[7]/NET0131  , \core_dag_ilm1reg_I_reg[8]/NET0131  , \core_dag_ilm1reg_I_reg[9]/NET0131  , \core_dag_ilm1reg_L0_we_DO_reg[0]/NET0131  , \core_dag_ilm1reg_L0_we_DO_reg[10]/NET0131  , \core_dag_ilm1reg_L0_we_DO_reg[11]/NET0131  , \core_dag_ilm1reg_L0_we_DO_reg[12]/NET0131  , \core_dag_ilm1reg_L0_we_DO_reg[13]/NET0131  , \core_dag_ilm1reg_L0_we_DO_reg[1]/NET0131  , \core_dag_ilm1reg_L0_we_DO_reg[2]/NET0131  , \core_dag_ilm1reg_L0_we_DO_reg[3]/NET0131  , \core_dag_ilm1reg_L0_we_DO_reg[4]/NET0131  , \core_dag_ilm1reg_L0_we_DO_reg[5]/NET0131  , \core_dag_ilm1reg_L0_we_DO_reg[6]/NET0131  , \core_dag_ilm1reg_L0_we_DO_reg[7]/NET0131  , \core_dag_ilm1reg_L0_we_DO_reg[8]/NET0131  , \core_dag_ilm1reg_L0_we_DO_reg[9]/NET0131  , \core_dag_ilm1reg_L1_we_DO_reg[0]/NET0131  , \core_dag_ilm1reg_L1_we_DO_reg[10]/NET0131  , \core_dag_ilm1reg_L1_we_DO_reg[11]/NET0131  , \core_dag_ilm1reg_L1_we_DO_reg[12]/NET0131  , \core_dag_ilm1reg_L1_we_DO_reg[13]/NET0131  , \core_dag_ilm1reg_L1_we_DO_reg[1]/NET0131  , \core_dag_ilm1reg_L1_we_DO_reg[2]/NET0131  , \core_dag_ilm1reg_L1_we_DO_reg[3]/NET0131  , \core_dag_ilm1reg_L1_we_DO_reg[4]/NET0131  , \core_dag_ilm1reg_L1_we_DO_reg[5]/NET0131  , \core_dag_ilm1reg_L1_we_DO_reg[6]/NET0131  , \core_dag_ilm1reg_L1_we_DO_reg[7]/NET0131  , \core_dag_ilm1reg_L1_we_DO_reg[8]/NET0131  , \core_dag_ilm1reg_L1_we_DO_reg[9]/NET0131  , \core_dag_ilm1reg_L2_we_DO_reg[0]/NET0131  , \core_dag_ilm1reg_L2_we_DO_reg[10]/NET0131  , \core_dag_ilm1reg_L2_we_DO_reg[11]/NET0131  , \core_dag_ilm1reg_L2_we_DO_reg[12]/NET0131  , \core_dag_ilm1reg_L2_we_DO_reg[13]/NET0131  , \core_dag_ilm1reg_L2_we_DO_reg[1]/NET0131  , \core_dag_ilm1reg_L2_we_DO_reg[2]/NET0131  , \core_dag_ilm1reg_L2_we_DO_reg[3]/NET0131  , \core_dag_ilm1reg_L2_we_DO_reg[4]/NET0131  , \core_dag_ilm1reg_L2_we_DO_reg[5]/NET0131  , \core_dag_ilm1reg_L2_we_DO_reg[6]/NET0131  , \core_dag_ilm1reg_L2_we_DO_reg[7]/NET0131  , \core_dag_ilm1reg_L2_we_DO_reg[8]/NET0131  , \core_dag_ilm1reg_L2_we_DO_reg[9]/NET0131  , \core_dag_ilm1reg_L3_we_DO_reg[0]/NET0131  , \core_dag_ilm1reg_L3_we_DO_reg[10]/NET0131  , \core_dag_ilm1reg_L3_we_DO_reg[11]/NET0131  , \core_dag_ilm1reg_L3_we_DO_reg[12]/NET0131  , \core_dag_ilm1reg_L3_we_DO_reg[13]/NET0131  , \core_dag_ilm1reg_L3_we_DO_reg[1]/NET0131  , \core_dag_ilm1reg_L3_we_DO_reg[2]/NET0131  , \core_dag_ilm1reg_L3_we_DO_reg[3]/NET0131  , \core_dag_ilm1reg_L3_we_DO_reg[4]/NET0131  , \core_dag_ilm1reg_L3_we_DO_reg[5]/NET0131  , \core_dag_ilm1reg_L3_we_DO_reg[6]/NET0131  , \core_dag_ilm1reg_L3_we_DO_reg[7]/NET0131  , \core_dag_ilm1reg_L3_we_DO_reg[8]/NET0131  , \core_dag_ilm1reg_L3_we_DO_reg[9]/NET0131  , \core_dag_ilm1reg_L_reg[0]/NET0131  , \core_dag_ilm1reg_L_reg[10]/NET0131  , \core_dag_ilm1reg_L_reg[11]/NET0131  , \core_dag_ilm1reg_L_reg[12]/NET0131  , \core_dag_ilm1reg_L_reg[13]/NET0131  , \core_dag_ilm1reg_L_reg[1]/NET0131  , \core_dag_ilm1reg_L_reg[2]/NET0131  , \core_dag_ilm1reg_L_reg[3]/NET0131  , \core_dag_ilm1reg_L_reg[4]/NET0131  , \core_dag_ilm1reg_L_reg[5]/NET0131  , \core_dag_ilm1reg_L_reg[6]/NET0131  , \core_dag_ilm1reg_L_reg[7]/NET0131  , \core_dag_ilm1reg_L_reg[8]/NET0131  , \core_dag_ilm1reg_L_reg[9]/NET0131  , \core_dag_ilm1reg_M0_we_DO_reg[0]/NET0131  , \core_dag_ilm1reg_M0_we_DO_reg[10]/NET0131  , \core_dag_ilm1reg_M0_we_DO_reg[11]/NET0131  , \core_dag_ilm1reg_M0_we_DO_reg[12]/NET0131  , \core_dag_ilm1reg_M0_we_DO_reg[13]/NET0131  , \core_dag_ilm1reg_M0_we_DO_reg[1]/NET0131  , \core_dag_ilm1reg_M0_we_DO_reg[2]/NET0131  , \core_dag_ilm1reg_M0_we_DO_reg[3]/NET0131  , \core_dag_ilm1reg_M0_we_DO_reg[4]/NET0131  , \core_dag_ilm1reg_M0_we_DO_reg[5]/NET0131  , \core_dag_ilm1reg_M0_we_DO_reg[6]/NET0131  , \core_dag_ilm1reg_M0_we_DO_reg[7]/NET0131  , \core_dag_ilm1reg_M0_we_DO_reg[8]/NET0131  , \core_dag_ilm1reg_M0_we_DO_reg[9]/NET0131  , \core_dag_ilm1reg_M1_we_DO_reg[0]/NET0131  , \core_dag_ilm1reg_M1_we_DO_reg[10]/NET0131  , \core_dag_ilm1reg_M1_we_DO_reg[11]/NET0131  , \core_dag_ilm1reg_M1_we_DO_reg[12]/NET0131  , \core_dag_ilm1reg_M1_we_DO_reg[13]/NET0131  , \core_dag_ilm1reg_M1_we_DO_reg[1]/NET0131  , \core_dag_ilm1reg_M1_we_DO_reg[2]/NET0131  , \core_dag_ilm1reg_M1_we_DO_reg[3]/NET0131  , \core_dag_ilm1reg_M1_we_DO_reg[4]/NET0131  , \core_dag_ilm1reg_M1_we_DO_reg[5]/NET0131  , \core_dag_ilm1reg_M1_we_DO_reg[6]/NET0131  , \core_dag_ilm1reg_M1_we_DO_reg[7]/NET0131  , \core_dag_ilm1reg_M1_we_DO_reg[8]/NET0131  , \core_dag_ilm1reg_M1_we_DO_reg[9]/NET0131  , \core_dag_ilm1reg_M2_we_DO_reg[0]/NET0131  , \core_dag_ilm1reg_M2_we_DO_reg[10]/NET0131  , \core_dag_ilm1reg_M2_we_DO_reg[11]/NET0131  , \core_dag_ilm1reg_M2_we_DO_reg[12]/NET0131  , \core_dag_ilm1reg_M2_we_DO_reg[13]/NET0131  , \core_dag_ilm1reg_M2_we_DO_reg[1]/NET0131  , \core_dag_ilm1reg_M2_we_DO_reg[2]/NET0131  , \core_dag_ilm1reg_M2_we_DO_reg[3]/NET0131  , \core_dag_ilm1reg_M2_we_DO_reg[4]/NET0131  , \core_dag_ilm1reg_M2_we_DO_reg[5]/NET0131  , \core_dag_ilm1reg_M2_we_DO_reg[6]/NET0131  , \core_dag_ilm1reg_M2_we_DO_reg[7]/NET0131  , \core_dag_ilm1reg_M2_we_DO_reg[8]/NET0131  , \core_dag_ilm1reg_M2_we_DO_reg[9]/NET0131  , \core_dag_ilm1reg_M3_we_DO_reg[0]/NET0131  , \core_dag_ilm1reg_M3_we_DO_reg[10]/NET0131  , \core_dag_ilm1reg_M3_we_DO_reg[11]/NET0131  , \core_dag_ilm1reg_M3_we_DO_reg[12]/NET0131  , \core_dag_ilm1reg_M3_we_DO_reg[13]/NET0131  , \core_dag_ilm1reg_M3_we_DO_reg[1]/NET0131  , \core_dag_ilm1reg_M3_we_DO_reg[2]/NET0131  , \core_dag_ilm1reg_M3_we_DO_reg[3]/NET0131  , \core_dag_ilm1reg_M3_we_DO_reg[4]/NET0131  , \core_dag_ilm1reg_M3_we_DO_reg[5]/NET0131  , \core_dag_ilm1reg_M3_we_DO_reg[6]/NET0131  , \core_dag_ilm1reg_M3_we_DO_reg[7]/NET0131  , \core_dag_ilm1reg_M3_we_DO_reg[8]/NET0131  , \core_dag_ilm1reg_M3_we_DO_reg[9]/NET0131  , \core_dag_ilm1reg_M_reg[0]/NET0131  , \core_dag_ilm1reg_M_reg[10]/NET0131  , \core_dag_ilm1reg_M_reg[11]/NET0131  , \core_dag_ilm1reg_M_reg[12]/NET0131  , \core_dag_ilm1reg_M_reg[13]/NET0131  , \core_dag_ilm1reg_M_reg[1]/NET0131  , \core_dag_ilm1reg_M_reg[2]/NET0131  , \core_dag_ilm1reg_M_reg[3]/NET0131  , \core_dag_ilm1reg_M_reg[4]/NET0131  , \core_dag_ilm1reg_M_reg[5]/NET0131  , \core_dag_ilm1reg_M_reg[6]/NET0131  , \core_dag_ilm1reg_M_reg[7]/NET0131  , \core_dag_ilm1reg_M_reg[8]/NET0131  , \core_dag_ilm1reg_M_reg[9]/NET0131  , \core_dag_ilm1reg_STAC_pi_DO_reg[0]/NET0131  , \core_dag_ilm1reg_STAC_pi_DO_reg[10]/NET0131  , \core_dag_ilm1reg_STAC_pi_DO_reg[11]/NET0131  , \core_dag_ilm1reg_STAC_pi_DO_reg[12]/NET0131  , \core_dag_ilm1reg_STAC_pi_DO_reg[13]/NET0131  , \core_dag_ilm1reg_STAC_pi_DO_reg[1]/NET0131  , \core_dag_ilm1reg_STAC_pi_DO_reg[2]/NET0131  , \core_dag_ilm1reg_STAC_pi_DO_reg[3]/NET0131  , \core_dag_ilm1reg_STAC_pi_DO_reg[4]/NET0131  , \core_dag_ilm1reg_STAC_pi_DO_reg[5]/NET0131  , \core_dag_ilm1reg_STAC_pi_DO_reg[6]/NET0131  , \core_dag_ilm1reg_STAC_pi_DO_reg[7]/NET0131  , \core_dag_ilm1reg_STAC_pi_DO_reg[8]/NET0131  , \core_dag_ilm1reg_STAC_pi_DO_reg[9]/NET0131  , \core_dag_ilm1reg_STEALI_E_reg[0]/P0001  , \core_dag_ilm1reg_STEALI_E_reg[1]/P0001  , \core_dag_ilm1reg_STEALI_E_reg[2]/P0001  , \core_dag_ilm2reg_I4_we_DO_reg[0]/NET0131  , \core_dag_ilm2reg_I4_we_DO_reg[10]/NET0131  , \core_dag_ilm2reg_I4_we_DO_reg[11]/NET0131  , \core_dag_ilm2reg_I4_we_DO_reg[12]/NET0131  , \core_dag_ilm2reg_I4_we_DO_reg[13]/NET0131  , \core_dag_ilm2reg_I4_we_DO_reg[1]/NET0131  , \core_dag_ilm2reg_I4_we_DO_reg[2]/NET0131  , \core_dag_ilm2reg_I4_we_DO_reg[3]/NET0131  , \core_dag_ilm2reg_I4_we_DO_reg[4]/NET0131  , \core_dag_ilm2reg_I4_we_DO_reg[5]/NET0131  , \core_dag_ilm2reg_I4_we_DO_reg[6]/NET0131  , \core_dag_ilm2reg_I4_we_DO_reg[7]/NET0131  , \core_dag_ilm2reg_I4_we_DO_reg[8]/NET0131  , \core_dag_ilm2reg_I4_we_DO_reg[9]/NET0131  , \core_dag_ilm2reg_I5_we_DO_reg[0]/NET0131  , \core_dag_ilm2reg_I5_we_DO_reg[10]/NET0131  , \core_dag_ilm2reg_I5_we_DO_reg[11]/NET0131  , \core_dag_ilm2reg_I5_we_DO_reg[12]/NET0131  , \core_dag_ilm2reg_I5_we_DO_reg[13]/NET0131  , \core_dag_ilm2reg_I5_we_DO_reg[1]/NET0131  , \core_dag_ilm2reg_I5_we_DO_reg[2]/NET0131  , \core_dag_ilm2reg_I5_we_DO_reg[3]/NET0131  , \core_dag_ilm2reg_I5_we_DO_reg[4]/NET0131  , \core_dag_ilm2reg_I5_we_DO_reg[5]/NET0131  , \core_dag_ilm2reg_I5_we_DO_reg[6]/NET0131  , \core_dag_ilm2reg_I5_we_DO_reg[7]/NET0131  , \core_dag_ilm2reg_I5_we_DO_reg[8]/NET0131  , \core_dag_ilm2reg_I5_we_DO_reg[9]/NET0131  , \core_dag_ilm2reg_I6_we_DO_reg[0]/NET0131  , \core_dag_ilm2reg_I6_we_DO_reg[10]/NET0131  , \core_dag_ilm2reg_I6_we_DO_reg[11]/NET0131  , \core_dag_ilm2reg_I6_we_DO_reg[12]/NET0131  , \core_dag_ilm2reg_I6_we_DO_reg[13]/NET0131  , \core_dag_ilm2reg_I6_we_DO_reg[1]/NET0131  , \core_dag_ilm2reg_I6_we_DO_reg[2]/NET0131  , \core_dag_ilm2reg_I6_we_DO_reg[3]/NET0131  , \core_dag_ilm2reg_I6_we_DO_reg[4]/NET0131  , \core_dag_ilm2reg_I6_we_DO_reg[5]/NET0131  , \core_dag_ilm2reg_I6_we_DO_reg[6]/NET0131  , \core_dag_ilm2reg_I6_we_DO_reg[7]/NET0131  , \core_dag_ilm2reg_I6_we_DO_reg[8]/NET0131  , \core_dag_ilm2reg_I6_we_DO_reg[9]/NET0131  , \core_dag_ilm2reg_I7_we_DO_reg[0]/NET0131  , \core_dag_ilm2reg_I7_we_DO_reg[10]/NET0131  , \core_dag_ilm2reg_I7_we_DO_reg[11]/NET0131  , \core_dag_ilm2reg_I7_we_DO_reg[12]/NET0131  , \core_dag_ilm2reg_I7_we_DO_reg[13]/NET0131  , \core_dag_ilm2reg_I7_we_DO_reg[1]/NET0131  , \core_dag_ilm2reg_I7_we_DO_reg[2]/NET0131  , \core_dag_ilm2reg_I7_we_DO_reg[3]/NET0131  , \core_dag_ilm2reg_I7_we_DO_reg[4]/NET0131  , \core_dag_ilm2reg_I7_we_DO_reg[5]/NET0131  , \core_dag_ilm2reg_I7_we_DO_reg[6]/NET0131  , \core_dag_ilm2reg_I7_we_DO_reg[7]/NET0131  , \core_dag_ilm2reg_I7_we_DO_reg[8]/NET0131  , \core_dag_ilm2reg_I7_we_DO_reg[9]/NET0131  , \core_dag_ilm2reg_IL_E_reg[0]/P0001  , \core_dag_ilm2reg_IL_E_reg[1]/P0001  , \core_dag_ilm2reg_I_reg[0]/NET0131  , \core_dag_ilm2reg_I_reg[10]/NET0131  , \core_dag_ilm2reg_I_reg[11]/NET0131  , \core_dag_ilm2reg_I_reg[12]/NET0131  , \core_dag_ilm2reg_I_reg[13]/NET0131  , \core_dag_ilm2reg_I_reg[1]/NET0131  , \core_dag_ilm2reg_I_reg[2]/NET0131  , \core_dag_ilm2reg_I_reg[3]/NET0131  , \core_dag_ilm2reg_I_reg[4]/NET0131  , \core_dag_ilm2reg_I_reg[5]/NET0131  , \core_dag_ilm2reg_I_reg[6]/NET0131  , \core_dag_ilm2reg_I_reg[7]/NET0131  , \core_dag_ilm2reg_I_reg[8]/NET0131  , \core_dag_ilm2reg_I_reg[9]/NET0131  , \core_dag_ilm2reg_L4_we_DO_reg[0]/NET0131  , \core_dag_ilm2reg_L4_we_DO_reg[10]/NET0131  , \core_dag_ilm2reg_L4_we_DO_reg[11]/NET0131  , \core_dag_ilm2reg_L4_we_DO_reg[12]/NET0131  , \core_dag_ilm2reg_L4_we_DO_reg[13]/NET0131  , \core_dag_ilm2reg_L4_we_DO_reg[1]/NET0131  , \core_dag_ilm2reg_L4_we_DO_reg[2]/NET0131  , \core_dag_ilm2reg_L4_we_DO_reg[3]/NET0131  , \core_dag_ilm2reg_L4_we_DO_reg[4]/NET0131  , \core_dag_ilm2reg_L4_we_DO_reg[5]/NET0131  , \core_dag_ilm2reg_L4_we_DO_reg[6]/NET0131  , \core_dag_ilm2reg_L4_we_DO_reg[7]/NET0131  , \core_dag_ilm2reg_L4_we_DO_reg[8]/NET0131  , \core_dag_ilm2reg_L4_we_DO_reg[9]/NET0131  , \core_dag_ilm2reg_L5_we_DO_reg[0]/NET0131  , \core_dag_ilm2reg_L5_we_DO_reg[10]/NET0131  , \core_dag_ilm2reg_L5_we_DO_reg[11]/NET0131  , \core_dag_ilm2reg_L5_we_DO_reg[12]/NET0131  , \core_dag_ilm2reg_L5_we_DO_reg[13]/NET0131  , \core_dag_ilm2reg_L5_we_DO_reg[1]/NET0131  , \core_dag_ilm2reg_L5_we_DO_reg[2]/NET0131  , \core_dag_ilm2reg_L5_we_DO_reg[3]/NET0131  , \core_dag_ilm2reg_L5_we_DO_reg[4]/NET0131  , \core_dag_ilm2reg_L5_we_DO_reg[5]/NET0131  , \core_dag_ilm2reg_L5_we_DO_reg[6]/NET0131  , \core_dag_ilm2reg_L5_we_DO_reg[7]/NET0131  , \core_dag_ilm2reg_L5_we_DO_reg[8]/NET0131  , \core_dag_ilm2reg_L5_we_DO_reg[9]/NET0131  , \core_dag_ilm2reg_L6_we_DO_reg[0]/NET0131  , \core_dag_ilm2reg_L6_we_DO_reg[10]/NET0131  , \core_dag_ilm2reg_L6_we_DO_reg[11]/NET0131  , \core_dag_ilm2reg_L6_we_DO_reg[12]/NET0131  , \core_dag_ilm2reg_L6_we_DO_reg[13]/NET0131  , \core_dag_ilm2reg_L6_we_DO_reg[1]/NET0131  , \core_dag_ilm2reg_L6_we_DO_reg[2]/NET0131  , \core_dag_ilm2reg_L6_we_DO_reg[3]/NET0131  , \core_dag_ilm2reg_L6_we_DO_reg[4]/NET0131  , \core_dag_ilm2reg_L6_we_DO_reg[5]/NET0131  , \core_dag_ilm2reg_L6_we_DO_reg[6]/NET0131  , \core_dag_ilm2reg_L6_we_DO_reg[7]/NET0131  , \core_dag_ilm2reg_L6_we_DO_reg[8]/NET0131  , \core_dag_ilm2reg_L6_we_DO_reg[9]/NET0131  , \core_dag_ilm2reg_L7_we_DO_reg[0]/NET0131  , \core_dag_ilm2reg_L7_we_DO_reg[10]/NET0131  , \core_dag_ilm2reg_L7_we_DO_reg[11]/NET0131  , \core_dag_ilm2reg_L7_we_DO_reg[12]/NET0131  , \core_dag_ilm2reg_L7_we_DO_reg[13]/NET0131  , \core_dag_ilm2reg_L7_we_DO_reg[1]/NET0131  , \core_dag_ilm2reg_L7_we_DO_reg[2]/NET0131  , \core_dag_ilm2reg_L7_we_DO_reg[3]/NET0131  , \core_dag_ilm2reg_L7_we_DO_reg[4]/NET0131  , \core_dag_ilm2reg_L7_we_DO_reg[5]/NET0131  , \core_dag_ilm2reg_L7_we_DO_reg[6]/NET0131  , \core_dag_ilm2reg_L7_we_DO_reg[7]/NET0131  , \core_dag_ilm2reg_L7_we_DO_reg[8]/NET0131  , \core_dag_ilm2reg_L7_we_DO_reg[9]/NET0131  , \core_dag_ilm2reg_L_reg[0]/NET0131  , \core_dag_ilm2reg_L_reg[10]/NET0131  , \core_dag_ilm2reg_L_reg[11]/NET0131  , \core_dag_ilm2reg_L_reg[12]/NET0131  , \core_dag_ilm2reg_L_reg[13]/NET0131  , \core_dag_ilm2reg_L_reg[1]/NET0131  , \core_dag_ilm2reg_L_reg[2]/NET0131  , \core_dag_ilm2reg_L_reg[3]/NET0131  , \core_dag_ilm2reg_L_reg[4]/NET0131  , \core_dag_ilm2reg_L_reg[5]/NET0131  , \core_dag_ilm2reg_L_reg[6]/NET0131  , \core_dag_ilm2reg_L_reg[7]/NET0131  , \core_dag_ilm2reg_L_reg[8]/NET0131  , \core_dag_ilm2reg_L_reg[9]/NET0131  , \core_dag_ilm2reg_M4_we_DO_reg[0]/NET0131  , \core_dag_ilm2reg_M4_we_DO_reg[10]/NET0131  , \core_dag_ilm2reg_M4_we_DO_reg[11]/NET0131  , \core_dag_ilm2reg_M4_we_DO_reg[12]/NET0131  , \core_dag_ilm2reg_M4_we_DO_reg[13]/NET0131  , \core_dag_ilm2reg_M4_we_DO_reg[1]/NET0131  , \core_dag_ilm2reg_M4_we_DO_reg[2]/NET0131  , \core_dag_ilm2reg_M4_we_DO_reg[3]/NET0131  , \core_dag_ilm2reg_M4_we_DO_reg[4]/NET0131  , \core_dag_ilm2reg_M4_we_DO_reg[5]/NET0131  , \core_dag_ilm2reg_M4_we_DO_reg[6]/NET0131  , \core_dag_ilm2reg_M4_we_DO_reg[7]/NET0131  , \core_dag_ilm2reg_M4_we_DO_reg[8]/NET0131  , \core_dag_ilm2reg_M4_we_DO_reg[9]/NET0131  , \core_dag_ilm2reg_M5_we_DO_reg[0]/NET0131  , \core_dag_ilm2reg_M5_we_DO_reg[10]/NET0131  , \core_dag_ilm2reg_M5_we_DO_reg[11]/NET0131  , \core_dag_ilm2reg_M5_we_DO_reg[12]/NET0131  , \core_dag_ilm2reg_M5_we_DO_reg[13]/NET0131  , \core_dag_ilm2reg_M5_we_DO_reg[1]/NET0131  , \core_dag_ilm2reg_M5_we_DO_reg[2]/NET0131  , \core_dag_ilm2reg_M5_we_DO_reg[3]/NET0131  , \core_dag_ilm2reg_M5_we_DO_reg[4]/NET0131  , \core_dag_ilm2reg_M5_we_DO_reg[5]/NET0131  , \core_dag_ilm2reg_M5_we_DO_reg[6]/NET0131  , \core_dag_ilm2reg_M5_we_DO_reg[7]/NET0131  , \core_dag_ilm2reg_M5_we_DO_reg[8]/NET0131  , \core_dag_ilm2reg_M5_we_DO_reg[9]/NET0131  , \core_dag_ilm2reg_M6_we_DO_reg[0]/NET0131  , \core_dag_ilm2reg_M6_we_DO_reg[10]/NET0131  , \core_dag_ilm2reg_M6_we_DO_reg[11]/NET0131  , \core_dag_ilm2reg_M6_we_DO_reg[12]/NET0131  , \core_dag_ilm2reg_M6_we_DO_reg[13]/NET0131  , \core_dag_ilm2reg_M6_we_DO_reg[1]/NET0131  , \core_dag_ilm2reg_M6_we_DO_reg[2]/NET0131  , \core_dag_ilm2reg_M6_we_DO_reg[3]/NET0131  , \core_dag_ilm2reg_M6_we_DO_reg[4]/NET0131  , \core_dag_ilm2reg_M6_we_DO_reg[5]/NET0131  , \core_dag_ilm2reg_M6_we_DO_reg[6]/NET0131  , \core_dag_ilm2reg_M6_we_DO_reg[7]/NET0131  , \core_dag_ilm2reg_M6_we_DO_reg[8]/NET0131  , \core_dag_ilm2reg_M6_we_DO_reg[9]/NET0131  , \core_dag_ilm2reg_M7_we_DO_reg[0]/NET0131  , \core_dag_ilm2reg_M7_we_DO_reg[10]/NET0131  , \core_dag_ilm2reg_M7_we_DO_reg[11]/NET0131  , \core_dag_ilm2reg_M7_we_DO_reg[12]/NET0131  , \core_dag_ilm2reg_M7_we_DO_reg[13]/NET0131  , \core_dag_ilm2reg_M7_we_DO_reg[1]/NET0131  , \core_dag_ilm2reg_M7_we_DO_reg[2]/NET0131  , \core_dag_ilm2reg_M7_we_DO_reg[3]/NET0131  , \core_dag_ilm2reg_M7_we_DO_reg[4]/NET0131  , \core_dag_ilm2reg_M7_we_DO_reg[5]/NET0131  , \core_dag_ilm2reg_M7_we_DO_reg[6]/NET0131  , \core_dag_ilm2reg_M7_we_DO_reg[7]/NET0131  , \core_dag_ilm2reg_M7_we_DO_reg[8]/NET0131  , \core_dag_ilm2reg_M7_we_DO_reg[9]/NET0131  , \core_dag_ilm2reg_M_E_reg[0]/NET0131  , \core_dag_ilm2reg_M_E_reg[1]/NET0131  , \core_dag_ilm2reg_M_reg[0]/NET0131  , \core_dag_ilm2reg_M_reg[10]/NET0131  , \core_dag_ilm2reg_M_reg[11]/NET0131  , \core_dag_ilm2reg_M_reg[12]/NET0131  , \core_dag_ilm2reg_M_reg[13]/NET0131  , \core_dag_ilm2reg_M_reg[1]/NET0131  , \core_dag_ilm2reg_M_reg[2]/NET0131  , \core_dag_ilm2reg_M_reg[3]/NET0131  , \core_dag_ilm2reg_M_reg[4]/NET0131  , \core_dag_ilm2reg_M_reg[5]/NET0131  , \core_dag_ilm2reg_M_reg[6]/NET0131  , \core_dag_ilm2reg_M_reg[7]/NET0131  , \core_dag_ilm2reg_M_reg[8]/NET0131  , \core_dag_ilm2reg_M_reg[9]/NET0131  , \core_dag_ilm2reg_PMA_pi_DO_reg[0]/NET0131  , \core_dag_ilm2reg_PMA_pi_DO_reg[10]/NET0131  , \core_dag_ilm2reg_PMA_pi_DO_reg[11]/NET0131  , \core_dag_ilm2reg_PMA_pi_DO_reg[12]/NET0131  , \core_dag_ilm2reg_PMA_pi_DO_reg[13]/NET0131  , \core_dag_ilm2reg_PMA_pi_DO_reg[1]/NET0131  , \core_dag_ilm2reg_PMA_pi_DO_reg[2]/NET0131  , \core_dag_ilm2reg_PMA_pi_DO_reg[3]/NET0131  , \core_dag_ilm2reg_PMA_pi_DO_reg[4]/NET0131  , \core_dag_ilm2reg_PMA_pi_DO_reg[5]/NET0131  , \core_dag_ilm2reg_PMA_pi_DO_reg[6]/NET0131  , \core_dag_ilm2reg_PMA_pi_DO_reg[7]/NET0131  , \core_dag_ilm2reg_PMA_pi_DO_reg[8]/NET0131  , \core_dag_ilm2reg_PMA_pi_DO_reg[9]/NET0131  , \core_dag_modulo1_R0wrap_reg/P0001  , \core_dag_modulo1_R1wrap_reg/P0001  , \core_dag_modulo1_T0wrap_reg/P0001  , \core_dag_modulo1_T1wrap_reg/P0001  , \core_eu_ea_alu_ea_dec_AMF_E_reg[0]/NET0131  , \core_eu_ea_alu_ea_dec_AMF_E_reg[1]/NET0131  , \core_eu_ea_alu_ea_dec_AMF_E_reg[2]/NET0131  , \core_eu_ea_alu_ea_dec_AMF_E_reg[3]/NET0131  , \core_eu_ea_alu_ea_dec_AMF_E_reg[4]/NET0131  , \core_eu_ea_alu_ea_dec_piconst_DO_reg[0]/P0001  , \core_eu_ea_alu_ea_dec_piconst_DO_reg[10]/P0001  , \core_eu_ea_alu_ea_dec_piconst_DO_reg[11]/P0001  , \core_eu_ea_alu_ea_dec_piconst_DO_reg[12]/P0001  , \core_eu_ea_alu_ea_dec_piconst_DO_reg[13]/P0001  , \core_eu_ea_alu_ea_dec_piconst_DO_reg[14]/P0001  , \core_eu_ea_alu_ea_dec_piconst_DO_reg[15]/P0001  , \core_eu_ea_alu_ea_dec_piconst_DO_reg[1]/P0001  , \core_eu_ea_alu_ea_dec_piconst_DO_reg[2]/P0001  , \core_eu_ea_alu_ea_dec_piconst_DO_reg[3]/P0001  , \core_eu_ea_alu_ea_dec_piconst_DO_reg[4]/P0001  , \core_eu_ea_alu_ea_dec_piconst_DO_reg[5]/P0001  , \core_eu_ea_alu_ea_dec_piconst_DO_reg[6]/P0001  , \core_eu_ea_alu_ea_dec_piconst_DO_reg[7]/P0001  , \core_eu_ea_alu_ea_dec_piconst_DO_reg[8]/P0001  , \core_eu_ea_alu_ea_dec_piconst_DO_reg[9]/P0001  , \core_eu_ea_alu_ea_reg_afrwe_DO_reg[0]/P0001  , \core_eu_ea_alu_ea_reg_afrwe_DO_reg[10]/P0001  , \core_eu_ea_alu_ea_reg_afrwe_DO_reg[11]/P0001  , \core_eu_ea_alu_ea_reg_afrwe_DO_reg[12]/P0001  , \core_eu_ea_alu_ea_reg_afrwe_DO_reg[13]/P0001  , \core_eu_ea_alu_ea_reg_afrwe_DO_reg[14]/P0001  , \core_eu_ea_alu_ea_reg_afrwe_DO_reg[15]/P0001  , \core_eu_ea_alu_ea_reg_afrwe_DO_reg[1]/P0001  , \core_eu_ea_alu_ea_reg_afrwe_DO_reg[2]/P0001  , \core_eu_ea_alu_ea_reg_afrwe_DO_reg[3]/P0001  , \core_eu_ea_alu_ea_reg_afrwe_DO_reg[4]/P0001  , \core_eu_ea_alu_ea_reg_afrwe_DO_reg[5]/P0001  , \core_eu_ea_alu_ea_reg_afrwe_DO_reg[6]/P0001  , \core_eu_ea_alu_ea_reg_afrwe_DO_reg[7]/P0001  , \core_eu_ea_alu_ea_reg_afrwe_DO_reg[8]/P0001  , \core_eu_ea_alu_ea_reg_afrwe_DO_reg[9]/P0001  , \core_eu_ea_alu_ea_reg_afswe_DO_reg[0]/P0001  , \core_eu_ea_alu_ea_reg_afswe_DO_reg[10]/P0001  , \core_eu_ea_alu_ea_reg_afswe_DO_reg[11]/P0001  , \core_eu_ea_alu_ea_reg_afswe_DO_reg[12]/P0001  , \core_eu_ea_alu_ea_reg_afswe_DO_reg[13]/P0001  , \core_eu_ea_alu_ea_reg_afswe_DO_reg[14]/P0001  , \core_eu_ea_alu_ea_reg_afswe_DO_reg[15]/P0001  , \core_eu_ea_alu_ea_reg_afswe_DO_reg[1]/P0001  , \core_eu_ea_alu_ea_reg_afswe_DO_reg[2]/P0001  , \core_eu_ea_alu_ea_reg_afswe_DO_reg[3]/P0001  , \core_eu_ea_alu_ea_reg_afswe_DO_reg[4]/P0001  , \core_eu_ea_alu_ea_reg_afswe_DO_reg[5]/P0001  , \core_eu_ea_alu_ea_reg_afswe_DO_reg[6]/P0001  , \core_eu_ea_alu_ea_reg_afswe_DO_reg[7]/P0001  , \core_eu_ea_alu_ea_reg_afswe_DO_reg[8]/P0001  , \core_eu_ea_alu_ea_reg_afswe_DO_reg[9]/P0001  , \core_eu_ea_alu_ea_reg_arrwe_DO_reg[0]/P0001  , \core_eu_ea_alu_ea_reg_arrwe_DO_reg[10]/P0001  , \core_eu_ea_alu_ea_reg_arrwe_DO_reg[11]/P0001  , \core_eu_ea_alu_ea_reg_arrwe_DO_reg[12]/P0001  , \core_eu_ea_alu_ea_reg_arrwe_DO_reg[13]/P0001  , \core_eu_ea_alu_ea_reg_arrwe_DO_reg[14]/P0001  , \core_eu_ea_alu_ea_reg_arrwe_DO_reg[15]/P0001  , \core_eu_ea_alu_ea_reg_arrwe_DO_reg[1]/P0001  , \core_eu_ea_alu_ea_reg_arrwe_DO_reg[2]/P0001  , \core_eu_ea_alu_ea_reg_arrwe_DO_reg[3]/P0001  , \core_eu_ea_alu_ea_reg_arrwe_DO_reg[4]/P0001  , \core_eu_ea_alu_ea_reg_arrwe_DO_reg[5]/P0001  , \core_eu_ea_alu_ea_reg_arrwe_DO_reg[6]/P0001  , \core_eu_ea_alu_ea_reg_arrwe_DO_reg[7]/P0001  , \core_eu_ea_alu_ea_reg_arrwe_DO_reg[8]/P0001  , \core_eu_ea_alu_ea_reg_arrwe_DO_reg[9]/P0001  , \core_eu_ea_alu_ea_reg_arswe_DO_reg[0]/P0001  , \core_eu_ea_alu_ea_reg_arswe_DO_reg[10]/P0001  , \core_eu_ea_alu_ea_reg_arswe_DO_reg[11]/P0001  , \core_eu_ea_alu_ea_reg_arswe_DO_reg[12]/P0001  , \core_eu_ea_alu_ea_reg_arswe_DO_reg[13]/P0001  , \core_eu_ea_alu_ea_reg_arswe_DO_reg[14]/P0001  , \core_eu_ea_alu_ea_reg_arswe_DO_reg[15]/P0001  , \core_eu_ea_alu_ea_reg_arswe_DO_reg[1]/P0001  , \core_eu_ea_alu_ea_reg_arswe_DO_reg[2]/P0001  , \core_eu_ea_alu_ea_reg_arswe_DO_reg[3]/P0001  , \core_eu_ea_alu_ea_reg_arswe_DO_reg[4]/P0001  , \core_eu_ea_alu_ea_reg_arswe_DO_reg[5]/P0001  , \core_eu_ea_alu_ea_reg_arswe_DO_reg[6]/P0001  , \core_eu_ea_alu_ea_reg_arswe_DO_reg[7]/P0001  , \core_eu_ea_alu_ea_reg_arswe_DO_reg[8]/P0001  , \core_eu_ea_alu_ea_reg_arswe_DO_reg[9]/P0001  , \core_eu_ea_alu_ea_reg_ax0rwe_DO_reg[0]/P0001  , \core_eu_ea_alu_ea_reg_ax0rwe_DO_reg[10]/P0001  , \core_eu_ea_alu_ea_reg_ax0rwe_DO_reg[11]/P0001  , \core_eu_ea_alu_ea_reg_ax0rwe_DO_reg[12]/P0001  , \core_eu_ea_alu_ea_reg_ax0rwe_DO_reg[13]/P0001  , \core_eu_ea_alu_ea_reg_ax0rwe_DO_reg[14]/P0001  , \core_eu_ea_alu_ea_reg_ax0rwe_DO_reg[15]/P0001  , \core_eu_ea_alu_ea_reg_ax0rwe_DO_reg[1]/P0001  , \core_eu_ea_alu_ea_reg_ax0rwe_DO_reg[2]/P0001  , \core_eu_ea_alu_ea_reg_ax0rwe_DO_reg[3]/P0001  , \core_eu_ea_alu_ea_reg_ax0rwe_DO_reg[4]/P0001  , \core_eu_ea_alu_ea_reg_ax0rwe_DO_reg[5]/P0001  , \core_eu_ea_alu_ea_reg_ax0rwe_DO_reg[6]/P0001  , \core_eu_ea_alu_ea_reg_ax0rwe_DO_reg[7]/P0001  , \core_eu_ea_alu_ea_reg_ax0rwe_DO_reg[8]/P0001  , \core_eu_ea_alu_ea_reg_ax0rwe_DO_reg[9]/P0001  , \core_eu_ea_alu_ea_reg_ax0swe_DO_reg[0]/P0001  , \core_eu_ea_alu_ea_reg_ax0swe_DO_reg[10]/P0001  , \core_eu_ea_alu_ea_reg_ax0swe_DO_reg[11]/P0001  , \core_eu_ea_alu_ea_reg_ax0swe_DO_reg[12]/P0001  , \core_eu_ea_alu_ea_reg_ax0swe_DO_reg[13]/P0001  , \core_eu_ea_alu_ea_reg_ax0swe_DO_reg[14]/P0001  , \core_eu_ea_alu_ea_reg_ax0swe_DO_reg[15]/P0001  , \core_eu_ea_alu_ea_reg_ax0swe_DO_reg[1]/P0001  , \core_eu_ea_alu_ea_reg_ax0swe_DO_reg[2]/P0001  , \core_eu_ea_alu_ea_reg_ax0swe_DO_reg[3]/P0001  , \core_eu_ea_alu_ea_reg_ax0swe_DO_reg[4]/P0001  , \core_eu_ea_alu_ea_reg_ax0swe_DO_reg[5]/P0001  , \core_eu_ea_alu_ea_reg_ax0swe_DO_reg[6]/P0001  , \core_eu_ea_alu_ea_reg_ax0swe_DO_reg[7]/P0001  , \core_eu_ea_alu_ea_reg_ax0swe_DO_reg[8]/P0001  , \core_eu_ea_alu_ea_reg_ax0swe_DO_reg[9]/P0001  , \core_eu_ea_alu_ea_reg_ax1rwe_DO_reg[0]/P0001  , \core_eu_ea_alu_ea_reg_ax1rwe_DO_reg[10]/P0001  , \core_eu_ea_alu_ea_reg_ax1rwe_DO_reg[11]/P0001  , \core_eu_ea_alu_ea_reg_ax1rwe_DO_reg[12]/P0001  , \core_eu_ea_alu_ea_reg_ax1rwe_DO_reg[13]/P0001  , \core_eu_ea_alu_ea_reg_ax1rwe_DO_reg[14]/P0001  , \core_eu_ea_alu_ea_reg_ax1rwe_DO_reg[15]/P0001  , \core_eu_ea_alu_ea_reg_ax1rwe_DO_reg[1]/P0001  , \core_eu_ea_alu_ea_reg_ax1rwe_DO_reg[2]/P0001  , \core_eu_ea_alu_ea_reg_ax1rwe_DO_reg[3]/P0001  , \core_eu_ea_alu_ea_reg_ax1rwe_DO_reg[4]/P0001  , \core_eu_ea_alu_ea_reg_ax1rwe_DO_reg[5]/P0001  , \core_eu_ea_alu_ea_reg_ax1rwe_DO_reg[6]/P0001  , \core_eu_ea_alu_ea_reg_ax1rwe_DO_reg[7]/P0001  , \core_eu_ea_alu_ea_reg_ax1rwe_DO_reg[8]/P0001  , \core_eu_ea_alu_ea_reg_ax1rwe_DO_reg[9]/P0001  , \core_eu_ea_alu_ea_reg_ax1swe_DO_reg[0]/P0001  , \core_eu_ea_alu_ea_reg_ax1swe_DO_reg[10]/P0001  , \core_eu_ea_alu_ea_reg_ax1swe_DO_reg[11]/P0001  , \core_eu_ea_alu_ea_reg_ax1swe_DO_reg[12]/P0001  , \core_eu_ea_alu_ea_reg_ax1swe_DO_reg[13]/P0001  , \core_eu_ea_alu_ea_reg_ax1swe_DO_reg[14]/P0001  , \core_eu_ea_alu_ea_reg_ax1swe_DO_reg[15]/P0001  , \core_eu_ea_alu_ea_reg_ax1swe_DO_reg[1]/P0001  , \core_eu_ea_alu_ea_reg_ax1swe_DO_reg[2]/P0001  , \core_eu_ea_alu_ea_reg_ax1swe_DO_reg[3]/P0001  , \core_eu_ea_alu_ea_reg_ax1swe_DO_reg[4]/P0001  , \core_eu_ea_alu_ea_reg_ax1swe_DO_reg[5]/P0001  , \core_eu_ea_alu_ea_reg_ax1swe_DO_reg[6]/P0001  , \core_eu_ea_alu_ea_reg_ax1swe_DO_reg[7]/P0001  , \core_eu_ea_alu_ea_reg_ax1swe_DO_reg[8]/P0001  , \core_eu_ea_alu_ea_reg_ax1swe_DO_reg[9]/P0001  , \core_eu_ea_alu_ea_reg_ay0rwe_DO_reg[0]/P0001  , \core_eu_ea_alu_ea_reg_ay0rwe_DO_reg[10]/P0001  , \core_eu_ea_alu_ea_reg_ay0rwe_DO_reg[11]/P0001  , \core_eu_ea_alu_ea_reg_ay0rwe_DO_reg[12]/P0001  , \core_eu_ea_alu_ea_reg_ay0rwe_DO_reg[13]/P0001  , \core_eu_ea_alu_ea_reg_ay0rwe_DO_reg[14]/P0001  , \core_eu_ea_alu_ea_reg_ay0rwe_DO_reg[15]/P0001  , \core_eu_ea_alu_ea_reg_ay0rwe_DO_reg[1]/P0001  , \core_eu_ea_alu_ea_reg_ay0rwe_DO_reg[2]/P0001  , \core_eu_ea_alu_ea_reg_ay0rwe_DO_reg[3]/P0001  , \core_eu_ea_alu_ea_reg_ay0rwe_DO_reg[4]/P0001  , \core_eu_ea_alu_ea_reg_ay0rwe_DO_reg[5]/P0001  , \core_eu_ea_alu_ea_reg_ay0rwe_DO_reg[6]/P0001  , \core_eu_ea_alu_ea_reg_ay0rwe_DO_reg[7]/P0001  , \core_eu_ea_alu_ea_reg_ay0rwe_DO_reg[8]/P0001  , \core_eu_ea_alu_ea_reg_ay0rwe_DO_reg[9]/P0001  , \core_eu_ea_alu_ea_reg_ay0swe_DO_reg[0]/P0001  , \core_eu_ea_alu_ea_reg_ay0swe_DO_reg[10]/P0001  , \core_eu_ea_alu_ea_reg_ay0swe_DO_reg[11]/P0001  , \core_eu_ea_alu_ea_reg_ay0swe_DO_reg[12]/P0001  , \core_eu_ea_alu_ea_reg_ay0swe_DO_reg[13]/P0001  , \core_eu_ea_alu_ea_reg_ay0swe_DO_reg[14]/P0001  , \core_eu_ea_alu_ea_reg_ay0swe_DO_reg[15]/P0001  , \core_eu_ea_alu_ea_reg_ay0swe_DO_reg[1]/P0001  , \core_eu_ea_alu_ea_reg_ay0swe_DO_reg[2]/P0001  , \core_eu_ea_alu_ea_reg_ay0swe_DO_reg[3]/P0001  , \core_eu_ea_alu_ea_reg_ay0swe_DO_reg[4]/P0001  , \core_eu_ea_alu_ea_reg_ay0swe_DO_reg[5]/P0001  , \core_eu_ea_alu_ea_reg_ay0swe_DO_reg[6]/P0001  , \core_eu_ea_alu_ea_reg_ay0swe_DO_reg[7]/P0001  , \core_eu_ea_alu_ea_reg_ay0swe_DO_reg[8]/P0001  , \core_eu_ea_alu_ea_reg_ay0swe_DO_reg[9]/P0001  , \core_eu_ea_alu_ea_reg_ay1rwe_DO_reg[0]/P0001  , \core_eu_ea_alu_ea_reg_ay1rwe_DO_reg[10]/P0001  , \core_eu_ea_alu_ea_reg_ay1rwe_DO_reg[11]/P0001  , \core_eu_ea_alu_ea_reg_ay1rwe_DO_reg[12]/P0001  , \core_eu_ea_alu_ea_reg_ay1rwe_DO_reg[13]/P0001  , \core_eu_ea_alu_ea_reg_ay1rwe_DO_reg[14]/P0001  , \core_eu_ea_alu_ea_reg_ay1rwe_DO_reg[15]/P0001  , \core_eu_ea_alu_ea_reg_ay1rwe_DO_reg[1]/P0001  , \core_eu_ea_alu_ea_reg_ay1rwe_DO_reg[2]/P0001  , \core_eu_ea_alu_ea_reg_ay1rwe_DO_reg[3]/P0001  , \core_eu_ea_alu_ea_reg_ay1rwe_DO_reg[4]/P0001  , \core_eu_ea_alu_ea_reg_ay1rwe_DO_reg[5]/P0001  , \core_eu_ea_alu_ea_reg_ay1rwe_DO_reg[6]/P0001  , \core_eu_ea_alu_ea_reg_ay1rwe_DO_reg[7]/P0001  , \core_eu_ea_alu_ea_reg_ay1rwe_DO_reg[8]/P0001  , \core_eu_ea_alu_ea_reg_ay1rwe_DO_reg[9]/P0001  , \core_eu_ea_alu_ea_reg_ay1swe_DO_reg[0]/P0001  , \core_eu_ea_alu_ea_reg_ay1swe_DO_reg[10]/P0001  , \core_eu_ea_alu_ea_reg_ay1swe_DO_reg[11]/P0001  , \core_eu_ea_alu_ea_reg_ay1swe_DO_reg[12]/P0001  , \core_eu_ea_alu_ea_reg_ay1swe_DO_reg[13]/P0001  , \core_eu_ea_alu_ea_reg_ay1swe_DO_reg[14]/P0001  , \core_eu_ea_alu_ea_reg_ay1swe_DO_reg[15]/P0001  , \core_eu_ea_alu_ea_reg_ay1swe_DO_reg[1]/P0001  , \core_eu_ea_alu_ea_reg_ay1swe_DO_reg[2]/P0001  , \core_eu_ea_alu_ea_reg_ay1swe_DO_reg[3]/P0001  , \core_eu_ea_alu_ea_reg_ay1swe_DO_reg[4]/P0001  , \core_eu_ea_alu_ea_reg_ay1swe_DO_reg[5]/P0001  , \core_eu_ea_alu_ea_reg_ay1swe_DO_reg[6]/P0001  , \core_eu_ea_alu_ea_reg_ay1swe_DO_reg[7]/P0001  , \core_eu_ea_alu_ea_reg_ay1swe_DO_reg[8]/P0001  , \core_eu_ea_alu_ea_reg_ay1swe_DO_reg[9]/P0001  , \core_eu_ec_cun_AC_reg/P0001  , \core_eu_ec_cun_AN_reg/P0001  , \core_eu_ec_cun_AQ_reg/P0001  , \core_eu_ec_cun_AS_reg/P0001  , \core_eu_ec_cun_AV_reg/P0001  , \core_eu_ec_cun_AZ_reg/P0001  , \core_eu_ec_cun_COND_E_reg[0]/P0001  , \core_eu_ec_cun_COND_E_reg[1]/P0001  , \core_eu_ec_cun_COND_E_reg[2]/P0001  , \core_eu_ec_cun_COND_E_reg[3]/P0001  , \core_eu_ec_cun_MV_reg/P0000_reg_syn_2  , \core_eu_ec_cun_MVi_pre_C_reg/P0001  , \core_eu_ec_cun_SS_reg/P0001  , \core_eu_ec_cun_TERM_E_reg[0]/P0001  , \core_eu_ec_cun_TERM_E_reg[1]/P0001  , \core_eu_ec_cun_TERM_E_reg[2]/P0001  , \core_eu_ec_cun_TERM_E_reg[3]/P0001  , \core_eu_ec_cun_condOK_CE_reg/P0001  , \core_eu_ec_cun_mven_FFout_reg/NET0131  , \core_eu_ec_cun_termOK_CE_reg/P0001  , \core_eu_ec_cun_updateMV_C_reg/P0001  , \core_eu_em_mac_em_dec_emcorepi_DO_reg[0]/P0001  , \core_eu_em_mac_em_dec_emcorepi_DO_reg[10]/P0001  , \core_eu_em_mac_em_dec_emcorepi_DO_reg[1]/P0001  , \core_eu_em_mac_em_dec_emcorepi_DO_reg[2]/P0001  , \core_eu_em_mac_em_dec_emcorepi_DO_reg[3]/P0001  , \core_eu_em_mac_em_reg_Sq_E_reg/P0001  , \core_eu_em_mac_em_reg_mfrwe_DO_reg[0]/P0001  , \core_eu_em_mac_em_reg_mfrwe_DO_reg[10]/P0001  , \core_eu_em_mac_em_reg_mfrwe_DO_reg[11]/P0001  , \core_eu_em_mac_em_reg_mfrwe_DO_reg[12]/P0001  , \core_eu_em_mac_em_reg_mfrwe_DO_reg[13]/P0001  , \core_eu_em_mac_em_reg_mfrwe_DO_reg[14]/P0001  , \core_eu_em_mac_em_reg_mfrwe_DO_reg[15]/P0001  , \core_eu_em_mac_em_reg_mfrwe_DO_reg[1]/P0001  , \core_eu_em_mac_em_reg_mfrwe_DO_reg[2]/P0001  , \core_eu_em_mac_em_reg_mfrwe_DO_reg[3]/P0001  , \core_eu_em_mac_em_reg_mfrwe_DO_reg[4]/P0001  , \core_eu_em_mac_em_reg_mfrwe_DO_reg[5]/P0001  , \core_eu_em_mac_em_reg_mfrwe_DO_reg[6]/P0001  , \core_eu_em_mac_em_reg_mfrwe_DO_reg[7]/P0001  , \core_eu_em_mac_em_reg_mfrwe_DO_reg[8]/P0001  , \core_eu_em_mac_em_reg_mfrwe_DO_reg[9]/P0001  , \core_eu_em_mac_em_reg_mfswe_DO_reg[0]/P0001  , \core_eu_em_mac_em_reg_mfswe_DO_reg[10]/P0001  , \core_eu_em_mac_em_reg_mfswe_DO_reg[11]/P0001  , \core_eu_em_mac_em_reg_mfswe_DO_reg[12]/P0001  , \core_eu_em_mac_em_reg_mfswe_DO_reg[13]/P0001  , \core_eu_em_mac_em_reg_mfswe_DO_reg[14]/P0001  , \core_eu_em_mac_em_reg_mfswe_DO_reg[15]/P0001  , \core_eu_em_mac_em_reg_mfswe_DO_reg[1]/P0001  , \core_eu_em_mac_em_reg_mfswe_DO_reg[2]/P0001  , \core_eu_em_mac_em_reg_mfswe_DO_reg[3]/P0001  , \core_eu_em_mac_em_reg_mfswe_DO_reg[4]/P0001  , \core_eu_em_mac_em_reg_mfswe_DO_reg[5]/P0001  , \core_eu_em_mac_em_reg_mfswe_DO_reg[6]/P0001  , \core_eu_em_mac_em_reg_mfswe_DO_reg[7]/P0001  , \core_eu_em_mac_em_reg_mfswe_DO_reg[8]/P0001  , \core_eu_em_mac_em_reg_mfswe_DO_reg[9]/P0001  , \core_eu_em_mac_em_reg_mr0rwe_DO_reg[0]/P0001  , \core_eu_em_mac_em_reg_mr0rwe_DO_reg[10]/P0001  , \core_eu_em_mac_em_reg_mr0rwe_DO_reg[11]/P0001  , \core_eu_em_mac_em_reg_mr0rwe_DO_reg[12]/P0001  , \core_eu_em_mac_em_reg_mr0rwe_DO_reg[13]/P0001  , \core_eu_em_mac_em_reg_mr0rwe_DO_reg[14]/P0001  , \core_eu_em_mac_em_reg_mr0rwe_DO_reg[15]/P0001  , \core_eu_em_mac_em_reg_mr0rwe_DO_reg[1]/P0001  , \core_eu_em_mac_em_reg_mr0rwe_DO_reg[2]/P0001  , \core_eu_em_mac_em_reg_mr0rwe_DO_reg[3]/P0001  , \core_eu_em_mac_em_reg_mr0rwe_DO_reg[4]/P0001  , \core_eu_em_mac_em_reg_mr0rwe_DO_reg[5]/P0001  , \core_eu_em_mac_em_reg_mr0rwe_DO_reg[6]/P0001  , \core_eu_em_mac_em_reg_mr0rwe_DO_reg[7]/P0001  , \core_eu_em_mac_em_reg_mr0rwe_DO_reg[8]/P0001  , \core_eu_em_mac_em_reg_mr0rwe_DO_reg[9]/P0001  , \core_eu_em_mac_em_reg_mr0swe_DO_reg[0]/P0001  , \core_eu_em_mac_em_reg_mr0swe_DO_reg[10]/P0001  , \core_eu_em_mac_em_reg_mr0swe_DO_reg[11]/P0001  , \core_eu_em_mac_em_reg_mr0swe_DO_reg[12]/P0001  , \core_eu_em_mac_em_reg_mr0swe_DO_reg[13]/P0001  , \core_eu_em_mac_em_reg_mr0swe_DO_reg[14]/P0001  , \core_eu_em_mac_em_reg_mr0swe_DO_reg[15]/P0001  , \core_eu_em_mac_em_reg_mr0swe_DO_reg[1]/P0001  , \core_eu_em_mac_em_reg_mr0swe_DO_reg[2]/P0001  , \core_eu_em_mac_em_reg_mr0swe_DO_reg[3]/P0001  , \core_eu_em_mac_em_reg_mr0swe_DO_reg[4]/P0001  , \core_eu_em_mac_em_reg_mr0swe_DO_reg[5]/P0001  , \core_eu_em_mac_em_reg_mr0swe_DO_reg[6]/P0001  , \core_eu_em_mac_em_reg_mr0swe_DO_reg[7]/P0001  , \core_eu_em_mac_em_reg_mr0swe_DO_reg[8]/P0001  , \core_eu_em_mac_em_reg_mr0swe_DO_reg[9]/P0001  , \core_eu_em_mac_em_reg_mr1rwe_DO_reg[0]/P0001  , \core_eu_em_mac_em_reg_mr1rwe_DO_reg[10]/P0001  , \core_eu_em_mac_em_reg_mr1rwe_DO_reg[11]/P0001  , \core_eu_em_mac_em_reg_mr1rwe_DO_reg[12]/P0001  , \core_eu_em_mac_em_reg_mr1rwe_DO_reg[13]/P0001  , \core_eu_em_mac_em_reg_mr1rwe_DO_reg[14]/P0001  , \core_eu_em_mac_em_reg_mr1rwe_DO_reg[15]/P0001  , \core_eu_em_mac_em_reg_mr1rwe_DO_reg[1]/P0001  , \core_eu_em_mac_em_reg_mr1rwe_DO_reg[2]/P0001  , \core_eu_em_mac_em_reg_mr1rwe_DO_reg[3]/P0001  , \core_eu_em_mac_em_reg_mr1rwe_DO_reg[4]/P0001  , \core_eu_em_mac_em_reg_mr1rwe_DO_reg[5]/P0001  , \core_eu_em_mac_em_reg_mr1rwe_DO_reg[6]/P0001  , \core_eu_em_mac_em_reg_mr1rwe_DO_reg[7]/P0001  , \core_eu_em_mac_em_reg_mr1rwe_DO_reg[8]/P0001  , \core_eu_em_mac_em_reg_mr1rwe_DO_reg[9]/P0001  , \core_eu_em_mac_em_reg_mr1swe_DO_reg[0]/P0001  , \core_eu_em_mac_em_reg_mr1swe_DO_reg[10]/P0001  , \core_eu_em_mac_em_reg_mr1swe_DO_reg[11]/P0001  , \core_eu_em_mac_em_reg_mr1swe_DO_reg[12]/P0001  , \core_eu_em_mac_em_reg_mr1swe_DO_reg[13]/P0001  , \core_eu_em_mac_em_reg_mr1swe_DO_reg[14]/P0001  , \core_eu_em_mac_em_reg_mr1swe_DO_reg[15]/P0001  , \core_eu_em_mac_em_reg_mr1swe_DO_reg[1]/P0001  , \core_eu_em_mac_em_reg_mr1swe_DO_reg[2]/P0001  , \core_eu_em_mac_em_reg_mr1swe_DO_reg[3]/P0001  , \core_eu_em_mac_em_reg_mr1swe_DO_reg[4]/P0001  , \core_eu_em_mac_em_reg_mr1swe_DO_reg[5]/P0001  , \core_eu_em_mac_em_reg_mr1swe_DO_reg[6]/P0001  , \core_eu_em_mac_em_reg_mr1swe_DO_reg[7]/P0001  , \core_eu_em_mac_em_reg_mr1swe_DO_reg[8]/P0001  , \core_eu_em_mac_em_reg_mr1swe_DO_reg[9]/P0001  , \core_eu_em_mac_em_reg_mr2rwe_DO_reg[0]/P0001  , \core_eu_em_mac_em_reg_mr2rwe_DO_reg[1]/P0001  , \core_eu_em_mac_em_reg_mr2rwe_DO_reg[2]/P0001  , \core_eu_em_mac_em_reg_mr2rwe_DO_reg[3]/P0001  , \core_eu_em_mac_em_reg_mr2rwe_DO_reg[4]/P0001  , \core_eu_em_mac_em_reg_mr2rwe_DO_reg[5]/P0001  , \core_eu_em_mac_em_reg_mr2rwe_DO_reg[6]/P0001  , \core_eu_em_mac_em_reg_mr2rwe_DO_reg[7]/P0001  , \core_eu_em_mac_em_reg_mr2swe_DO_reg[0]/P0001  , \core_eu_em_mac_em_reg_mr2swe_DO_reg[1]/P0001  , \core_eu_em_mac_em_reg_mr2swe_DO_reg[2]/P0001  , \core_eu_em_mac_em_reg_mr2swe_DO_reg[3]/P0001  , \core_eu_em_mac_em_reg_mr2swe_DO_reg[4]/P0001  , \core_eu_em_mac_em_reg_mr2swe_DO_reg[5]/P0001  , \core_eu_em_mac_em_reg_mr2swe_DO_reg[6]/P0001  , \core_eu_em_mac_em_reg_mr2swe_DO_reg[7]/P0001  , \core_eu_em_mac_em_reg_mrovfwe_DO_reg[0]/P0001  , \core_eu_em_mac_em_reg_mrovfwe_DO_reg[1]/P0001  , \core_eu_em_mac_em_reg_mrovfwe_DO_reg[2]/P0001  , \core_eu_em_mac_em_reg_mrovfwe_DO_reg[3]/P0001  , \core_eu_em_mac_em_reg_mrovfwe_DO_reg[4]/P0001  , \core_eu_em_mac_em_reg_mrovfwe_DO_reg[5]/P0001  , \core_eu_em_mac_em_reg_mrovfwe_DO_reg[6]/P0001  , \core_eu_em_mac_em_reg_mrovfwe_DO_reg[7]/P0001  , \core_eu_em_mac_em_reg_mrovfwe_DO_reg[8]/P0001  , \core_eu_em_mac_em_reg_mx0rwe_DO_reg[0]/P0001  , \core_eu_em_mac_em_reg_mx0rwe_DO_reg[10]/P0001  , \core_eu_em_mac_em_reg_mx0rwe_DO_reg[11]/P0001  , \core_eu_em_mac_em_reg_mx0rwe_DO_reg[12]/P0001  , \core_eu_em_mac_em_reg_mx0rwe_DO_reg[13]/P0001  , \core_eu_em_mac_em_reg_mx0rwe_DO_reg[14]/P0001  , \core_eu_em_mac_em_reg_mx0rwe_DO_reg[15]/P0001  , \core_eu_em_mac_em_reg_mx0rwe_DO_reg[1]/P0001  , \core_eu_em_mac_em_reg_mx0rwe_DO_reg[2]/P0001  , \core_eu_em_mac_em_reg_mx0rwe_DO_reg[3]/P0001  , \core_eu_em_mac_em_reg_mx0rwe_DO_reg[4]/P0001  , \core_eu_em_mac_em_reg_mx0rwe_DO_reg[5]/P0001  , \core_eu_em_mac_em_reg_mx0rwe_DO_reg[6]/P0001  , \core_eu_em_mac_em_reg_mx0rwe_DO_reg[7]/P0001  , \core_eu_em_mac_em_reg_mx0rwe_DO_reg[8]/P0001  , \core_eu_em_mac_em_reg_mx0rwe_DO_reg[9]/P0001  , \core_eu_em_mac_em_reg_mx0swe_DO_reg[0]/P0001  , \core_eu_em_mac_em_reg_mx0swe_DO_reg[10]/P0001  , \core_eu_em_mac_em_reg_mx0swe_DO_reg[11]/P0001  , \core_eu_em_mac_em_reg_mx0swe_DO_reg[12]/P0001  , \core_eu_em_mac_em_reg_mx0swe_DO_reg[13]/P0001  , \core_eu_em_mac_em_reg_mx0swe_DO_reg[14]/P0001  , \core_eu_em_mac_em_reg_mx0swe_DO_reg[15]/P0001  , \core_eu_em_mac_em_reg_mx0swe_DO_reg[1]/P0001  , \core_eu_em_mac_em_reg_mx0swe_DO_reg[2]/P0001  , \core_eu_em_mac_em_reg_mx0swe_DO_reg[3]/P0001  , \core_eu_em_mac_em_reg_mx0swe_DO_reg[4]/P0001  , \core_eu_em_mac_em_reg_mx0swe_DO_reg[5]/P0001  , \core_eu_em_mac_em_reg_mx0swe_DO_reg[6]/P0001  , \core_eu_em_mac_em_reg_mx0swe_DO_reg[7]/P0001  , \core_eu_em_mac_em_reg_mx0swe_DO_reg[8]/P0001  , \core_eu_em_mac_em_reg_mx0swe_DO_reg[9]/P0001  , \core_eu_em_mac_em_reg_mx1rwe_DO_reg[0]/P0001  , \core_eu_em_mac_em_reg_mx1rwe_DO_reg[10]/P0001  , \core_eu_em_mac_em_reg_mx1rwe_DO_reg[11]/P0001  , \core_eu_em_mac_em_reg_mx1rwe_DO_reg[12]/P0001  , \core_eu_em_mac_em_reg_mx1rwe_DO_reg[13]/P0001  , \core_eu_em_mac_em_reg_mx1rwe_DO_reg[14]/P0001  , \core_eu_em_mac_em_reg_mx1rwe_DO_reg[15]/P0001  , \core_eu_em_mac_em_reg_mx1rwe_DO_reg[1]/P0001  , \core_eu_em_mac_em_reg_mx1rwe_DO_reg[2]/P0001  , \core_eu_em_mac_em_reg_mx1rwe_DO_reg[3]/P0001  , \core_eu_em_mac_em_reg_mx1rwe_DO_reg[4]/P0001  , \core_eu_em_mac_em_reg_mx1rwe_DO_reg[5]/P0001  , \core_eu_em_mac_em_reg_mx1rwe_DO_reg[6]/P0001  , \core_eu_em_mac_em_reg_mx1rwe_DO_reg[7]/P0001  , \core_eu_em_mac_em_reg_mx1rwe_DO_reg[8]/P0001  , \core_eu_em_mac_em_reg_mx1rwe_DO_reg[9]/P0001  , \core_eu_em_mac_em_reg_mx1swe_DO_reg[0]/P0001  , \core_eu_em_mac_em_reg_mx1swe_DO_reg[10]/P0001  , \core_eu_em_mac_em_reg_mx1swe_DO_reg[11]/P0001  , \core_eu_em_mac_em_reg_mx1swe_DO_reg[12]/P0001  , \core_eu_em_mac_em_reg_mx1swe_DO_reg[13]/P0001  , \core_eu_em_mac_em_reg_mx1swe_DO_reg[14]/P0001  , \core_eu_em_mac_em_reg_mx1swe_DO_reg[15]/P0001  , \core_eu_em_mac_em_reg_mx1swe_DO_reg[1]/P0001  , \core_eu_em_mac_em_reg_mx1swe_DO_reg[2]/P0001  , \core_eu_em_mac_em_reg_mx1swe_DO_reg[3]/P0001  , \core_eu_em_mac_em_reg_mx1swe_DO_reg[4]/P0001  , \core_eu_em_mac_em_reg_mx1swe_DO_reg[5]/P0001  , \core_eu_em_mac_em_reg_mx1swe_DO_reg[6]/P0001  , \core_eu_em_mac_em_reg_mx1swe_DO_reg[7]/P0001  , \core_eu_em_mac_em_reg_mx1swe_DO_reg[8]/P0001  , \core_eu_em_mac_em_reg_mx1swe_DO_reg[9]/P0001  , \core_eu_em_mac_em_reg_mxopwe_DO_reg[0]/P0001  , \core_eu_em_mac_em_reg_mxopwe_DO_reg[10]/P0001  , \core_eu_em_mac_em_reg_mxopwe_DO_reg[11]/P0001  , \core_eu_em_mac_em_reg_mxopwe_DO_reg[12]/P0001  , \core_eu_em_mac_em_reg_mxopwe_DO_reg[13]/P0001  , \core_eu_em_mac_em_reg_mxopwe_DO_reg[14]/P0001  , \core_eu_em_mac_em_reg_mxopwe_DO_reg[15]/P0001  , \core_eu_em_mac_em_reg_mxopwe_DO_reg[1]/P0001  , \core_eu_em_mac_em_reg_mxopwe_DO_reg[2]/P0001  , \core_eu_em_mac_em_reg_mxopwe_DO_reg[3]/P0001  , \core_eu_em_mac_em_reg_mxopwe_DO_reg[4]/P0001  , \core_eu_em_mac_em_reg_mxopwe_DO_reg[5]/P0001  , \core_eu_em_mac_em_reg_mxopwe_DO_reg[6]/P0001  , \core_eu_em_mac_em_reg_mxopwe_DO_reg[7]/P0001  , \core_eu_em_mac_em_reg_mxopwe_DO_reg[8]/P0001  , \core_eu_em_mac_em_reg_mxopwe_DO_reg[9]/P0001  , \core_eu_em_mac_em_reg_my0rwe_DO_reg[0]/P0001  , \core_eu_em_mac_em_reg_my0rwe_DO_reg[10]/P0001  , \core_eu_em_mac_em_reg_my0rwe_DO_reg[11]/P0001  , \core_eu_em_mac_em_reg_my0rwe_DO_reg[12]/P0001  , \core_eu_em_mac_em_reg_my0rwe_DO_reg[13]/P0001  , \core_eu_em_mac_em_reg_my0rwe_DO_reg[14]/P0001  , \core_eu_em_mac_em_reg_my0rwe_DO_reg[15]/P0001  , \core_eu_em_mac_em_reg_my0rwe_DO_reg[1]/P0001  , \core_eu_em_mac_em_reg_my0rwe_DO_reg[2]/P0001  , \core_eu_em_mac_em_reg_my0rwe_DO_reg[3]/P0001  , \core_eu_em_mac_em_reg_my0rwe_DO_reg[4]/P0001  , \core_eu_em_mac_em_reg_my0rwe_DO_reg[5]/P0001  , \core_eu_em_mac_em_reg_my0rwe_DO_reg[6]/P0001  , \core_eu_em_mac_em_reg_my0rwe_DO_reg[7]/P0001  , \core_eu_em_mac_em_reg_my0rwe_DO_reg[8]/P0001  , \core_eu_em_mac_em_reg_my0rwe_DO_reg[9]/P0001  , \core_eu_em_mac_em_reg_my0swe_DO_reg[0]/P0001  , \core_eu_em_mac_em_reg_my0swe_DO_reg[10]/P0001  , \core_eu_em_mac_em_reg_my0swe_DO_reg[11]/P0001  , \core_eu_em_mac_em_reg_my0swe_DO_reg[12]/P0001  , \core_eu_em_mac_em_reg_my0swe_DO_reg[13]/P0001  , \core_eu_em_mac_em_reg_my0swe_DO_reg[14]/P0001  , \core_eu_em_mac_em_reg_my0swe_DO_reg[15]/P0001  , \core_eu_em_mac_em_reg_my0swe_DO_reg[1]/P0001  , \core_eu_em_mac_em_reg_my0swe_DO_reg[2]/P0001  , \core_eu_em_mac_em_reg_my0swe_DO_reg[3]/P0001  , \core_eu_em_mac_em_reg_my0swe_DO_reg[4]/P0001  , \core_eu_em_mac_em_reg_my0swe_DO_reg[5]/P0001  , \core_eu_em_mac_em_reg_my0swe_DO_reg[6]/P0001  , \core_eu_em_mac_em_reg_my0swe_DO_reg[7]/P0001  , \core_eu_em_mac_em_reg_my0swe_DO_reg[8]/P0001  , \core_eu_em_mac_em_reg_my0swe_DO_reg[9]/P0001  , \core_eu_em_mac_em_reg_my1rwe_DO_reg[0]/P0001  , \core_eu_em_mac_em_reg_my1rwe_DO_reg[10]/P0001  , \core_eu_em_mac_em_reg_my1rwe_DO_reg[11]/P0001  , \core_eu_em_mac_em_reg_my1rwe_DO_reg[12]/P0001  , \core_eu_em_mac_em_reg_my1rwe_DO_reg[13]/P0001  , \core_eu_em_mac_em_reg_my1rwe_DO_reg[14]/P0001  , \core_eu_em_mac_em_reg_my1rwe_DO_reg[15]/P0001  , \core_eu_em_mac_em_reg_my1rwe_DO_reg[1]/P0001  , \core_eu_em_mac_em_reg_my1rwe_DO_reg[2]/P0001  , \core_eu_em_mac_em_reg_my1rwe_DO_reg[3]/P0001  , \core_eu_em_mac_em_reg_my1rwe_DO_reg[4]/P0001  , \core_eu_em_mac_em_reg_my1rwe_DO_reg[5]/P0001  , \core_eu_em_mac_em_reg_my1rwe_DO_reg[6]/P0001  , \core_eu_em_mac_em_reg_my1rwe_DO_reg[7]/P0001  , \core_eu_em_mac_em_reg_my1rwe_DO_reg[8]/P0001  , \core_eu_em_mac_em_reg_my1rwe_DO_reg[9]/P0001  , \core_eu_em_mac_em_reg_my1swe_DO_reg[0]/P0001  , \core_eu_em_mac_em_reg_my1swe_DO_reg[10]/P0001  , \core_eu_em_mac_em_reg_my1swe_DO_reg[11]/P0001  , \core_eu_em_mac_em_reg_my1swe_DO_reg[12]/P0001  , \core_eu_em_mac_em_reg_my1swe_DO_reg[13]/P0001  , \core_eu_em_mac_em_reg_my1swe_DO_reg[14]/P0001  , \core_eu_em_mac_em_reg_my1swe_DO_reg[15]/P0001  , \core_eu_em_mac_em_reg_my1swe_DO_reg[1]/P0001  , \core_eu_em_mac_em_reg_my1swe_DO_reg[2]/P0001  , \core_eu_em_mac_em_reg_my1swe_DO_reg[3]/P0001  , \core_eu_em_mac_em_reg_my1swe_DO_reg[4]/P0001  , \core_eu_em_mac_em_reg_my1swe_DO_reg[5]/P0001  , \core_eu_em_mac_em_reg_my1swe_DO_reg[6]/P0001  , \core_eu_em_mac_em_reg_my1swe_DO_reg[7]/P0001  , \core_eu_em_mac_em_reg_my1swe_DO_reg[8]/P0001  , \core_eu_em_mac_em_reg_my1swe_DO_reg[9]/P0001  , \core_eu_em_mac_em_reg_myopwe_DO_reg[0]/P0001  , \core_eu_em_mac_em_reg_myopwe_DO_reg[10]/P0001  , \core_eu_em_mac_em_reg_myopwe_DO_reg[11]/P0001  , \core_eu_em_mac_em_reg_myopwe_DO_reg[12]/P0001  , \core_eu_em_mac_em_reg_myopwe_DO_reg[13]/P0001  , \core_eu_em_mac_em_reg_myopwe_DO_reg[14]/P0001  , \core_eu_em_mac_em_reg_myopwe_DO_reg[15]/P0001  , \core_eu_em_mac_em_reg_myopwe_DO_reg[1]/P0001  , \core_eu_em_mac_em_reg_myopwe_DO_reg[2]/P0001  , \core_eu_em_mac_em_reg_myopwe_DO_reg[3]/P0001  , \core_eu_em_mac_em_reg_myopwe_DO_reg[4]/P0001  , \core_eu_em_mac_em_reg_myopwe_DO_reg[5]/P0001  , \core_eu_em_mac_em_reg_myopwe_DO_reg[6]/P0001  , \core_eu_em_mac_em_reg_myopwe_DO_reg[7]/P0001  , \core_eu_em_mac_em_reg_myopwe_DO_reg[8]/P0001  , \core_eu_em_mac_em_reg_myopwe_DO_reg[9]/P0001  , \core_eu_em_mac_em_reg_s0_reg/P0000_reg_syn_2  , \core_eu_em_mac_em_reg_s1_reg/P0000_reg_syn_2  , \core_eu_em_mac_em_reg_s2_reg/P0000_reg_syn_2  , \core_eu_es_sht_es_reg_SBr_reg[0]/P0001  , \core_eu_es_sht_es_reg_SBr_reg[1]/P0001  , \core_eu_es_sht_es_reg_SBr_reg[2]/P0001  , \core_eu_es_sht_es_reg_SBr_reg[3]/P0001  , \core_eu_es_sht_es_reg_SBr_reg[4]/P0001  , \core_eu_es_sht_es_reg_SBs_reg[0]/P0001  , \core_eu_es_sht_es_reg_SBs_reg[1]/P0001  , \core_eu_es_sht_es_reg_SBs_reg[2]/P0001  , \core_eu_es_sht_es_reg_SBs_reg[3]/P0001  , \core_eu_es_sht_es_reg_SBs_reg[4]/P0001  , \core_eu_es_sht_es_reg_serwe_DO_reg[0]/P0001  , \core_eu_es_sht_es_reg_serwe_DO_reg[1]/P0001  , \core_eu_es_sht_es_reg_serwe_DO_reg[2]/P0001  , \core_eu_es_sht_es_reg_serwe_DO_reg[3]/P0001  , \core_eu_es_sht_es_reg_serwe_DO_reg[4]/P0001  , \core_eu_es_sht_es_reg_serwe_DO_reg[5]/P0001  , \core_eu_es_sht_es_reg_serwe_DO_reg[6]/P0001  , \core_eu_es_sht_es_reg_serwe_DO_reg[7]/P0001  , \core_eu_es_sht_es_reg_seswe_DO_reg[0]/P0001  , \core_eu_es_sht_es_reg_seswe_DO_reg[1]/P0001  , \core_eu_es_sht_es_reg_seswe_DO_reg[2]/P0001  , \core_eu_es_sht_es_reg_seswe_DO_reg[3]/P0001  , \core_eu_es_sht_es_reg_seswe_DO_reg[4]/P0001  , \core_eu_es_sht_es_reg_seswe_DO_reg[5]/P0001  , \core_eu_es_sht_es_reg_seswe_DO_reg[6]/P0001  , \core_eu_es_sht_es_reg_seswe_DO_reg[7]/P0001  , \core_eu_es_sht_es_reg_sirwe_DO_reg[0]/P0001  , \core_eu_es_sht_es_reg_sirwe_DO_reg[10]/P0001  , \core_eu_es_sht_es_reg_sirwe_DO_reg[11]/P0001  , \core_eu_es_sht_es_reg_sirwe_DO_reg[12]/P0001  , \core_eu_es_sht_es_reg_sirwe_DO_reg[13]/P0001  , \core_eu_es_sht_es_reg_sirwe_DO_reg[14]/P0001  , \core_eu_es_sht_es_reg_sirwe_DO_reg[15]/P0001  , \core_eu_es_sht_es_reg_sirwe_DO_reg[1]/P0001  , \core_eu_es_sht_es_reg_sirwe_DO_reg[2]/P0001  , \core_eu_es_sht_es_reg_sirwe_DO_reg[3]/P0001  , \core_eu_es_sht_es_reg_sirwe_DO_reg[4]/P0001  , \core_eu_es_sht_es_reg_sirwe_DO_reg[5]/P0001  , \core_eu_es_sht_es_reg_sirwe_DO_reg[6]/P0001  , \core_eu_es_sht_es_reg_sirwe_DO_reg[7]/P0001  , \core_eu_es_sht_es_reg_sirwe_DO_reg[8]/P0001  , \core_eu_es_sht_es_reg_sirwe_DO_reg[9]/P0001  , \core_eu_es_sht_es_reg_siswe_DO_reg[0]/P0001  , \core_eu_es_sht_es_reg_siswe_DO_reg[10]/P0001  , \core_eu_es_sht_es_reg_siswe_DO_reg[11]/P0001  , \core_eu_es_sht_es_reg_siswe_DO_reg[12]/P0001  , \core_eu_es_sht_es_reg_siswe_DO_reg[13]/P0001  , \core_eu_es_sht_es_reg_siswe_DO_reg[14]/P0001  , \core_eu_es_sht_es_reg_siswe_DO_reg[15]/P0001  , \core_eu_es_sht_es_reg_siswe_DO_reg[1]/P0001  , \core_eu_es_sht_es_reg_siswe_DO_reg[2]/P0001  , \core_eu_es_sht_es_reg_siswe_DO_reg[3]/P0001  , \core_eu_es_sht_es_reg_siswe_DO_reg[4]/P0001  , \core_eu_es_sht_es_reg_siswe_DO_reg[5]/P0001  , \core_eu_es_sht_es_reg_siswe_DO_reg[6]/P0001  , \core_eu_es_sht_es_reg_siswe_DO_reg[7]/P0001  , \core_eu_es_sht_es_reg_siswe_DO_reg[8]/P0001  , \core_eu_es_sht_es_reg_siswe_DO_reg[9]/P0001  , \core_eu_es_sht_es_reg_sr0rwe_DO_reg[0]/P0001  , \core_eu_es_sht_es_reg_sr0rwe_DO_reg[10]/P0001  , \core_eu_es_sht_es_reg_sr0rwe_DO_reg[11]/P0001  , \core_eu_es_sht_es_reg_sr0rwe_DO_reg[12]/P0001  , \core_eu_es_sht_es_reg_sr0rwe_DO_reg[13]/P0001  , \core_eu_es_sht_es_reg_sr0rwe_DO_reg[14]/P0001  , \core_eu_es_sht_es_reg_sr0rwe_DO_reg[15]/P0001  , \core_eu_es_sht_es_reg_sr0rwe_DO_reg[1]/P0001  , \core_eu_es_sht_es_reg_sr0rwe_DO_reg[2]/P0001  , \core_eu_es_sht_es_reg_sr0rwe_DO_reg[3]/P0001  , \core_eu_es_sht_es_reg_sr0rwe_DO_reg[4]/P0001  , \core_eu_es_sht_es_reg_sr0rwe_DO_reg[5]/P0001  , \core_eu_es_sht_es_reg_sr0rwe_DO_reg[6]/P0001  , \core_eu_es_sht_es_reg_sr0rwe_DO_reg[7]/P0001  , \core_eu_es_sht_es_reg_sr0rwe_DO_reg[8]/P0001  , \core_eu_es_sht_es_reg_sr0rwe_DO_reg[9]/P0001  , \core_eu_es_sht_es_reg_sr0swe_DO_reg[0]/P0001  , \core_eu_es_sht_es_reg_sr0swe_DO_reg[10]/P0001  , \core_eu_es_sht_es_reg_sr0swe_DO_reg[11]/P0001  , \core_eu_es_sht_es_reg_sr0swe_DO_reg[12]/P0001  , \core_eu_es_sht_es_reg_sr0swe_DO_reg[13]/P0001  , \core_eu_es_sht_es_reg_sr0swe_DO_reg[14]/P0001  , \core_eu_es_sht_es_reg_sr0swe_DO_reg[15]/P0001  , \core_eu_es_sht_es_reg_sr0swe_DO_reg[1]/P0001  , \core_eu_es_sht_es_reg_sr0swe_DO_reg[2]/P0001  , \core_eu_es_sht_es_reg_sr0swe_DO_reg[3]/P0001  , \core_eu_es_sht_es_reg_sr0swe_DO_reg[4]/P0001  , \core_eu_es_sht_es_reg_sr0swe_DO_reg[5]/P0001  , \core_eu_es_sht_es_reg_sr0swe_DO_reg[6]/P0001  , \core_eu_es_sht_es_reg_sr0swe_DO_reg[7]/P0001  , \core_eu_es_sht_es_reg_sr0swe_DO_reg[8]/P0001  , \core_eu_es_sht_es_reg_sr0swe_DO_reg[9]/P0001  , \core_eu_es_sht_es_reg_sr1rwe_DO_reg[0]/P0001  , \core_eu_es_sht_es_reg_sr1rwe_DO_reg[10]/P0001  , \core_eu_es_sht_es_reg_sr1rwe_DO_reg[11]/P0001  , \core_eu_es_sht_es_reg_sr1rwe_DO_reg[12]/P0001  , \core_eu_es_sht_es_reg_sr1rwe_DO_reg[13]/P0001  , \core_eu_es_sht_es_reg_sr1rwe_DO_reg[14]/P0001  , \core_eu_es_sht_es_reg_sr1rwe_DO_reg[15]/P0001  , \core_eu_es_sht_es_reg_sr1rwe_DO_reg[1]/P0001  , \core_eu_es_sht_es_reg_sr1rwe_DO_reg[2]/P0001  , \core_eu_es_sht_es_reg_sr1rwe_DO_reg[3]/P0001  , \core_eu_es_sht_es_reg_sr1rwe_DO_reg[4]/P0001  , \core_eu_es_sht_es_reg_sr1rwe_DO_reg[5]/P0001  , \core_eu_es_sht_es_reg_sr1rwe_DO_reg[6]/P0001  , \core_eu_es_sht_es_reg_sr1rwe_DO_reg[7]/P0001  , \core_eu_es_sht_es_reg_sr1rwe_DO_reg[8]/P0001  , \core_eu_es_sht_es_reg_sr1rwe_DO_reg[9]/P0001  , \core_eu_es_sht_es_reg_sr1swe_DO_reg[0]/P0001  , \core_eu_es_sht_es_reg_sr1swe_DO_reg[10]/P0001  , \core_eu_es_sht_es_reg_sr1swe_DO_reg[11]/P0001  , \core_eu_es_sht_es_reg_sr1swe_DO_reg[12]/P0001  , \core_eu_es_sht_es_reg_sr1swe_DO_reg[13]/P0001  , \core_eu_es_sht_es_reg_sr1swe_DO_reg[14]/P0001  , \core_eu_es_sht_es_reg_sr1swe_DO_reg[15]/P0001  , \core_eu_es_sht_es_reg_sr1swe_DO_reg[1]/P0001  , \core_eu_es_sht_es_reg_sr1swe_DO_reg[2]/P0001  , \core_eu_es_sht_es_reg_sr1swe_DO_reg[3]/P0001  , \core_eu_es_sht_es_reg_sr1swe_DO_reg[4]/P0001  , \core_eu_es_sht_es_reg_sr1swe_DO_reg[5]/P0001  , \core_eu_es_sht_es_reg_sr1swe_DO_reg[6]/P0001  , \core_eu_es_sht_es_reg_sr1swe_DO_reg[7]/P0001  , \core_eu_es_sht_es_reg_sr1swe_DO_reg[8]/P0001  , \core_eu_es_sht_es_reg_sr1swe_DO_reg[9]/P0001  , \emc_DMDoe_reg/NET0131  , \emc_DMDreg_reg[0]/P0001  , \emc_DMDreg_reg[10]/P0001  , \emc_DMDreg_reg[11]/P0001  , \emc_DMDreg_reg[12]/P0001  , \emc_DMDreg_reg[13]/P0001  , \emc_DMDreg_reg[14]/P0001  , \emc_DMDreg_reg[15]/P0001  , \emc_DMDreg_reg[1]/P0001  , \emc_DMDreg_reg[2]/P0001  , \emc_DMDreg_reg[3]/P0001  , \emc_DMDreg_reg[4]/P0001  , \emc_DMDreg_reg[5]/P0001  , \emc_DMDreg_reg[6]/P0001  , \emc_DMDreg_reg[7]/P0001  , \emc_DMDreg_reg[8]/P0001  , \emc_DMDreg_reg[9]/P0001  , \emc_DMcst_reg/NET0131  , \emc_ECMA_reg[0]/P0001  , \emc_ECMA_reg[10]/P0001  , \emc_ECMA_reg[11]/P0001  , \emc_ECMA_reg[12]/P0001  , \emc_ECMA_reg[1]/P0001  , \emc_ECMA_reg[2]/P0001  , \emc_ECMA_reg[3]/P0001  , \emc_ECMA_reg[4]/P0001  , \emc_ECMA_reg[5]/P0001  , \emc_ECMA_reg[6]/P0001  , \emc_ECMA_reg[7]/P0001  , \emc_ECMA_reg[8]/P0001  , \emc_ECMA_reg[9]/P0001  , \emc_ECMDreg_reg[0]/P0001  , \emc_ECMDreg_reg[10]/P0001  , \emc_ECMDreg_reg[11]/P0001  , \emc_ECMDreg_reg[12]/P0001  , \emc_ECMDreg_reg[13]/P0001  , \emc_ECMDreg_reg[14]/P0001  , \emc_ECMDreg_reg[15]/P0001  , \emc_ECMDreg_reg[16]/P0001  , \emc_ECMDreg_reg[17]/P0001  , \emc_ECMDreg_reg[18]/P0001  , \emc_ECMDreg_reg[19]/P0001  , \emc_ECMDreg_reg[1]/P0001  , \emc_ECMDreg_reg[20]/P0001  , \emc_ECMDreg_reg[21]/P0001  , \emc_ECMDreg_reg[22]/P0001  , \emc_ECMDreg_reg[23]/P0001  , \emc_ECMDreg_reg[2]/P0001  , \emc_ECMDreg_reg[3]/P0001  , \emc_ECMDreg_reg[4]/P0001  , \emc_ECMDreg_reg[5]/P0001  , \emc_ECMDreg_reg[6]/P0001  , \emc_ECMDreg_reg[7]/P0001  , \emc_ECMDreg_reg[8]/P0001  , \emc_ECMDreg_reg[9]/P0001  , \emc_ECMcs_reg/NET0131  , \emc_ECS_reg[0]/NET0131  , \emc_ECS_reg[1]/NET0131  , \emc_ECS_reg[2]/NET0131  , \emc_ECS_reg[3]/NET0131  , \emc_ED_oei_reg/P0001  , \emc_EXTC_Eg_syn_reg/P0001  , \emc_IOcst_reg/NET0131  , \emc_PMDoe_reg/NET0131  , \emc_PMDreg_reg[0]/P0001  , \emc_PMDreg_reg[10]/P0001  , \emc_PMDreg_reg[11]/P0001  , \emc_PMDreg_reg[12]/P0001  , \emc_PMDreg_reg[13]/P0001  , \emc_PMDreg_reg[14]/P0001  , \emc_PMDreg_reg[15]/P0001  , \emc_PMDreg_reg[1]/P0001  , \emc_PMDreg_reg[2]/P0001  , \emc_PMDreg_reg[3]/P0001  , \emc_PMDreg_reg[4]/P0001  , \emc_PMDreg_reg[5]/P0001  , \emc_PMDreg_reg[6]/P0001  , \emc_PMDreg_reg[7]/P0001  , \emc_PMDreg_reg[8]/P0001  , \emc_PMDreg_reg[9]/P0001  , \emc_PMcst_reg/NET0131  , \emc_RWcnt_reg[0]/P0001  , \emc_RWcnt_reg[1]/P0001  , \emc_RWcnt_reg[2]/P0001  , \emc_RWcnt_reg[3]/P0001  , \emc_RWcnt_reg[4]/P0001  , \emc_RWcnt_reg[5]/P0001  , \emc_WRn_h_reg/P0001  , \emc_WSCRext_reg_DO_reg[0]/NET0131  , \emc_WSCRext_reg_DO_reg[1]/NET0131  , \emc_WSCRext_reg_DO_reg[2]/NET0131  , \emc_WSCRext_reg_DO_reg[3]/NET0131  , \emc_WSCRext_reg_DO_reg[4]/NET0131  , \emc_WSCRext_reg_DO_reg[5]/NET0131  , \emc_WSCRext_reg_DO_reg[6]/NET0131  , \emc_WSCRext_reg_DO_reg[7]/NET0131  , \emc_WSCRreg_DO_reg[0]/NET0131  , \emc_WSCRreg_DO_reg[10]/NET0131  , \emc_WSCRreg_DO_reg[11]/NET0131  , \emc_WSCRreg_DO_reg[12]/NET0131  , \emc_WSCRreg_DO_reg[13]/NET0131  , \emc_WSCRreg_DO_reg[14]/NET0131  , \emc_WSCRreg_DO_reg[1]/NET0131  , \emc_WSCRreg_DO_reg[2]/NET0131  , \emc_WSCRreg_DO_reg[3]/NET0131  , \emc_WSCRreg_DO_reg[4]/NET0131  , \emc_WSCRreg_DO_reg[5]/NET0131  , \emc_WSCRreg_DO_reg[6]/NET0131  , \emc_WSCRreg_DO_reg[7]/NET0131  , \emc_WSCRreg_DO_reg[8]/NET0131  , \emc_WSCRreg_DO_reg[9]/NET0131  , \emc_eRDY_reg/NET0131  , \emc_selDMDi_reg/P0001  , \emc_selPMDi_reg/P0001  , \idma_CM_oe_reg/P0001  , \idma_CMo_oe0_reg/P0001  , \idma_CMo_oe1_reg/P0001  , \idma_CMo_oe2_reg/P0001  , \idma_CMo_oe3_reg/P0001  , \idma_CMo_oe4_reg/P0001  , \idma_CMo_oe5_reg/P0001  , \idma_CMo_oe6_reg/P0001  , \idma_CMo_oe7_reg/P0001  , \idma_DCTL_reg[0]/NET0131  , \idma_DCTL_reg[10]/NET0131  , \idma_DCTL_reg[11]/NET0131  , \idma_DCTL_reg[12]/NET0131  , \idma_DCTL_reg[13]/NET0131  , \idma_DCTL_reg[14]/NET0131  , \idma_DCTL_reg[1]/NET0131  , \idma_DCTL_reg[2]/NET0131  , \idma_DCTL_reg[3]/NET0131  , \idma_DCTL_reg[4]/NET0131  , \idma_DCTL_reg[5]/NET0131  , \idma_DCTL_reg[6]/NET0131  , \idma_DCTL_reg[7]/NET0131  , \idma_DCTL_reg[8]/NET0131  , \idma_DCTL_reg[9]/NET0131  , \idma_DOVL_reg[0]/NET0131  , \idma_DOVL_reg[10]/NET0131  , \idma_DOVL_reg[11]/NET0131  , \idma_DOVL_reg[1]/NET0131  , \idma_DOVL_reg[2]/NET0131  , \idma_DOVL_reg[3]/NET0131  , \idma_DOVL_reg[4]/NET0131  , \idma_DOVL_reg[5]/NET0131  , \idma_DOVL_reg[6]/NET0131  , \idma_DOVL_reg[7]/NET0131  , \idma_DOVL_reg[8]/NET0131  , \idma_DOVL_reg[9]/NET0131  , \idma_DSreq_reg/NET0131  , \idma_DTMP_H_reg[0]/P0001  , \idma_DTMP_H_reg[10]/P0001  , \idma_DTMP_H_reg[11]/P0001  , \idma_DTMP_H_reg[12]/P0001  , \idma_DTMP_H_reg[13]/P0001  , \idma_DTMP_H_reg[14]/P0001  , \idma_DTMP_H_reg[15]/P0001  , \idma_DTMP_H_reg[1]/P0001  , \idma_DTMP_H_reg[2]/P0001  , \idma_DTMP_H_reg[3]/P0001  , \idma_DTMP_H_reg[4]/P0001  , \idma_DTMP_H_reg[5]/P0001  , \idma_DTMP_H_reg[6]/P0001  , \idma_DTMP_H_reg[7]/P0001  , \idma_DTMP_H_reg[8]/P0001  , \idma_DTMP_H_reg[9]/P0001  , \idma_DTMP_L_reg[0]/P0001  , \idma_DTMP_L_reg[1]/P0001  , \idma_DTMP_L_reg[2]/P0001  , \idma_DTMP_L_reg[3]/P0001  , \idma_DTMP_L_reg[4]/P0001  , \idma_DTMP_L_reg[5]/P0001  , \idma_DTMP_L_reg[6]/P0001  , \idma_DTMP_L_reg[7]/P0001  , \idma_IADi_reg[0]/P0001  , \idma_IADi_reg[10]/P0001  , \idma_IADi_reg[11]/P0001  , \idma_IADi_reg[12]/P0001  , \idma_IADi_reg[13]/P0001  , \idma_IADi_reg[14]/P0001  , \idma_IADi_reg[15]/P0001  , \idma_IADi_reg[1]/P0001  , \idma_IADi_reg[2]/P0001  , \idma_IADi_reg[3]/P0001  , \idma_IADi_reg[4]/P0001  , \idma_IADi_reg[5]/P0001  , \idma_IADi_reg[6]/P0001  , \idma_IADi_reg[7]/P0001  , \idma_IADi_reg[8]/P0001  , \idma_IADi_reg[9]/P0001  , \idma_IAL_reg/P0001  , \idma_IDMA_boot_reg/NET0131_reg_syn_10  , \idma_IDMA_boot_reg/NET0131_reg_syn_2  , \idma_IDMA_boot_reg/NET0131_reg_syn_8  , \idma_IRDn_reg/P0001  , \idma_ISn_reg/P0001  , \idma_IWRn_reg/P0001  , \idma_PCrd_1st_reg/NET0131  , \idma_PM_1st_reg/NET0131  , \idma_RDCMD_d1_reg/P0001  , \idma_RDCMD_reg/P0001  , \idma_RDcnt_reg[0]/NET0131  , \idma_RDcnt_reg[1]/NET0131  , \idma_RDcnt_reg[2]/NET0131  , \idma_RDcyc_reg/NET0131  , \idma_WRCMD_d1_reg/P0001  , \idma_WRCMD_reg/P0001  , \idma_WRcnt_reg[0]/NET0131  , \idma_WRcnt_reg[1]/NET0131  , \idma_WRcnt_reg[2]/NET0131  , \idma_WRcyc_reg/NET0131  , \idma_WRtrue_reg/NET0131  , \memc_DM_oe_reg/P0001  , \memc_DMo_oe0_reg/P0001  , \memc_DMo_oe1_reg/P0001  , \memc_DMo_oe2_reg/P0001  , \memc_DMo_oe3_reg/P0001  , \memc_DMo_oe4_reg/P0001  , \memc_DMo_oe5_reg/P0001  , \memc_DMo_oe6_reg/P0001  , \memc_DMo_oe7_reg/P0001  , \memc_Dread_E_reg/NET0131  , \memc_Dwrite_C_reg/NET0131  , \memc_Dwrite_E_reg/NET0131  , \memc_EXTC_E_reg/NET0131  , \memc_EXTC_Eg_reg/NET0131_reg_syn_10  , \memc_EXTC_Eg_reg/NET0131_reg_syn_2  , \memc_EXTC_Eg_reg/NET0131_reg_syn_8  , \memc_IOcmd_E_reg/NET0131  , \memc_LDaST_Eg_reg/NET0131  , \memc_MMR_web_reg/NET0131  , \memc_PMo_oe0_reg/P0001  , \memc_PMo_oe1_reg/P0001  , \memc_PMo_oe2_reg/P0001  , \memc_PMo_oe3_reg/P0001  , \memc_PMo_oe4_reg/P0001  , \memc_PMo_oe5_reg/P0001  , \memc_PMo_oe6_reg/P0001  , \memc_PMo_oe7_reg/P0001  , \memc_Pread_E_reg/NET0131  , \memc_Pwrite_C_reg/NET0131  , \memc_Pwrite_E_reg/NET0131  , \memc_STI_Cg_reg/NET0131  , \memc_accDM_E_reg/NET0131  , \memc_accPM_E_reg/NET0131  , \memc_ldSREG_E_reg/NET0131  , \memc_selMIO_E_reg/P0001  , \memc_usysr_DO_reg[0]/NET0131  , \memc_usysr_DO_reg[10]/NET0131  , \memc_usysr_DO_reg[11]/NET0131  , \memc_usysr_DO_reg[12]/NET0131  , \memc_usysr_DO_reg[13]/NET0131  , \memc_usysr_DO_reg[14]/NET0131  , \memc_usysr_DO_reg[15]/NET0131  , \memc_usysr_DO_reg[1]/NET0131  , \memc_usysr_DO_reg[2]/NET0131  , \memc_usysr_DO_reg[3]/NET0131  , \memc_usysr_DO_reg[4]/NET0131  , \memc_usysr_DO_reg[5]/NET0131  , \memc_usysr_DO_reg[6]/NET0131  , \memc_usysr_DO_reg[7]/NET0131  , \memc_usysr_DO_reg[8]/NET0131  , \memc_usysr_DO_reg[9]/NET0131  , \pio_PINT_reg[0]/NET0131  , \pio_PINT_reg[10]/NET0131  , \pio_PINT_reg[11]/NET0131  , \pio_PINT_reg[1]/NET0131  , \pio_PINT_reg[2]/NET0131  , \pio_PINT_reg[3]/NET0131  , \pio_PINT_reg[4]/NET0131  , \pio_PINT_reg[5]/NET0131  , \pio_PINT_reg[6]/NET0131  , \pio_PINT_reg[7]/NET0131  , \pio_PINT_reg[8]/NET0131  , \pio_PINT_reg[9]/NET0131  , \pio_PIO_IN_P_reg[0]/P0001  , \pio_PIO_IN_P_reg[10]/P0001  , \pio_PIO_IN_P_reg[11]/P0001  , \pio_PIO_IN_P_reg[1]/P0001  , \pio_PIO_IN_P_reg[2]/P0001  , \pio_PIO_IN_P_reg[3]/P0001  , \pio_PIO_IN_P_reg[4]/P0001  , \pio_PIO_IN_P_reg[5]/P0001  , \pio_PIO_IN_P_reg[6]/P0001  , \pio_PIO_IN_P_reg[7]/P0001  , \pio_PIO_IN_P_reg[8]/P0001  , \pio_PIO_IN_P_reg[9]/P0001  , \pio_PIO_RES_OUT_reg[0]/P0001  , \pio_PIO_RES_OUT_reg[10]/P0001  , \pio_PIO_RES_OUT_reg[11]/P0001  , \pio_PIO_RES_OUT_reg[1]/P0001  , \pio_PIO_RES_OUT_reg[2]/P0001  , \pio_PIO_RES_OUT_reg[3]/P0001  , \pio_PIO_RES_OUT_reg[4]/P0001  , \pio_PIO_RES_OUT_reg[5]/P0001  , \pio_PIO_RES_OUT_reg[6]/P0001  , \pio_PIO_RES_OUT_reg[7]/P0001  , \pio_PIO_RES_OUT_reg[8]/P0001  , \pio_PIO_RES_OUT_reg[9]/P0001  , \pio_PIO_RES_reg[0]/NET0131  , \pio_PIO_RES_reg[10]/NET0131  , \pio_PIO_RES_reg[11]/NET0131  , \pio_PIO_RES_reg[1]/NET0131  , \pio_PIO_RES_reg[2]/NET0131  , \pio_PIO_RES_reg[3]/NET0131  , \pio_PIO_RES_reg[4]/NET0131  , \pio_PIO_RES_reg[5]/NET0131  , \pio_PIO_RES_reg[6]/NET0131  , \pio_PIO_RES_reg[7]/NET0131  , \pio_PIO_RES_reg[8]/NET0131  , \pio_PIO_RES_reg[9]/NET0131  , \pio_pmask_reg_DO_reg[0]/NET0131  , \pio_pmask_reg_DO_reg[10]/NET0131  , \pio_pmask_reg_DO_reg[11]/NET0131  , \pio_pmask_reg_DO_reg[1]/NET0131  , \pio_pmask_reg_DO_reg[2]/NET0131  , \pio_pmask_reg_DO_reg[3]/NET0131  , \pio_pmask_reg_DO_reg[4]/NET0131  , \pio_pmask_reg_DO_reg[5]/NET0131  , \pio_pmask_reg_DO_reg[6]/NET0131  , \pio_pmask_reg_DO_reg[7]/NET0131  , \pio_pmask_reg_DO_reg[8]/NET0131  , \pio_pmask_reg_DO_reg[9]/NET0131  , \regout_STD_C_reg[0]/P0001  , \regout_STD_C_reg[10]/P0001  , \regout_STD_C_reg[11]/P0001  , \regout_STD_C_reg[12]/P0001  , \regout_STD_C_reg[13]/P0001  , \regout_STD_C_reg[14]/P0001  , \regout_STD_C_reg[15]/P0001  , \regout_STD_C_reg[1]/P0001  , \regout_STD_C_reg[2]/P0001  , \regout_STD_C_reg[3]/P0001  , \regout_STD_C_reg[4]/P0001  , \regout_STD_C_reg[5]/P0001  , \regout_STD_C_reg[6]/P0001  , \regout_STD_C_reg[7]/P0001  , \regout_STD_C_reg[8]/P0001  , \regout_STD_C_reg[9]/P0001  , \sice_CLR_I_reg/NET0131  , \sice_CLR_M_reg/NET0131  , \sice_CMRW_reg/NET0131  , \sice_DBR1_reg[0]/P0001  , \sice_DBR1_reg[10]/P0001  , \sice_DBR1_reg[11]/P0001  , \sice_DBR1_reg[12]/P0001  , \sice_DBR1_reg[13]/P0001  , \sice_DBR1_reg[14]/P0001  , \sice_DBR1_reg[15]/P0001  , \sice_DBR1_reg[16]/P0001  , \sice_DBR1_reg[17]/P0001  , \sice_DBR1_reg[18]/P0001  , \sice_DBR1_reg[1]/P0001  , \sice_DBR1_reg[2]/P0001  , \sice_DBR1_reg[3]/P0001  , \sice_DBR1_reg[4]/P0001  , \sice_DBR1_reg[5]/P0001  , \sice_DBR1_reg[6]/P0001  , \sice_DBR1_reg[7]/P0001  , \sice_DBR1_reg[8]/P0001  , \sice_DBR1_reg[9]/P0001  , \sice_DBR2_reg[0]/P0001  , \sice_DBR2_reg[10]/P0001  , \sice_DBR2_reg[11]/P0001  , \sice_DBR2_reg[12]/P0001  , \sice_DBR2_reg[13]/P0001  , \sice_DBR2_reg[14]/P0001  , \sice_DBR2_reg[15]/P0001  , \sice_DBR2_reg[16]/P0001  , \sice_DBR2_reg[17]/P0001  , \sice_DBR2_reg[18]/P0001  , \sice_DBR2_reg[1]/P0001  , \sice_DBR2_reg[2]/P0001  , \sice_DBR2_reg[3]/P0001  , \sice_DBR2_reg[4]/P0001  , \sice_DBR2_reg[5]/P0001  , \sice_DBR2_reg[6]/P0001  , \sice_DBR2_reg[7]/P0001  , \sice_DBR2_reg[8]/P0001  , \sice_DBR2_reg[9]/P0001  , \sice_DMR1_reg[0]/NET0131  , \sice_DMR1_reg[10]/NET0131  , \sice_DMR1_reg[11]/NET0131  , \sice_DMR1_reg[12]/NET0131  , \sice_DMR1_reg[13]/NET0131  , \sice_DMR1_reg[14]/NET0131  , \sice_DMR1_reg[15]/NET0131  , \sice_DMR1_reg[16]/NET0131  , \sice_DMR1_reg[17]/NET0131  , \sice_DMR1_reg[1]/NET0131  , \sice_DMR1_reg[2]/NET0131  , \sice_DMR1_reg[3]/NET0131  , \sice_DMR1_reg[4]/NET0131  , \sice_DMR1_reg[5]/NET0131  , \sice_DMR1_reg[6]/NET0131  , \sice_DMR1_reg[7]/NET0131  , \sice_DMR1_reg[8]/NET0131  , \sice_DMR1_reg[9]/NET0131  , \sice_DMR2_reg[0]/NET0131  , \sice_DMR2_reg[10]/NET0131  , \sice_DMR2_reg[11]/NET0131  , \sice_DMR2_reg[12]/NET0131  , \sice_DMR2_reg[13]/NET0131  , \sice_DMR2_reg[14]/NET0131  , \sice_DMR2_reg[15]/NET0131  , \sice_DMR2_reg[16]/NET0131  , \sice_DMR2_reg[17]/NET0131  , \sice_DMR2_reg[1]/NET0131  , \sice_DMR2_reg[2]/NET0131  , \sice_DMR2_reg[3]/NET0131  , \sice_DMR2_reg[4]/NET0131  , \sice_DMR2_reg[5]/NET0131  , \sice_DMR2_reg[6]/NET0131  , \sice_DMR2_reg[7]/NET0131  , \sice_DMR2_reg[8]/NET0131  , \sice_DMR2_reg[9]/NET0131  , \sice_GOICE_1_reg/NET0131  , \sice_GOICE_2_reg/NET0131  , \sice_GOICE_s1_reg/NET0131  , \sice_GOICE_syn_reg/P0001  , \sice_GO_NX_reg/NET0131  , \sice_GO_NXi_reg/NET0131  , \sice_HALT_E_reg/P0001  , \sice_IAR_reg[0]/NET0131  , \sice_IAR_reg[1]/NET0131  , \sice_IAR_reg[2]/NET0131  , \sice_IAR_reg[3]/NET0131  , \sice_IBR1_reg[0]/P0001  , \sice_IBR1_reg[10]/P0001  , \sice_IBR1_reg[11]/P0001  , \sice_IBR1_reg[12]/P0001  , \sice_IBR1_reg[13]/P0001  , \sice_IBR1_reg[14]/P0001  , \sice_IBR1_reg[15]/P0001  , \sice_IBR1_reg[16]/P0001  , \sice_IBR1_reg[17]/P0001  , \sice_IBR1_reg[1]/P0001  , \sice_IBR1_reg[2]/P0001  , \sice_IBR1_reg[3]/P0001  , \sice_IBR1_reg[4]/P0001  , \sice_IBR1_reg[5]/P0001  , \sice_IBR1_reg[6]/P0001  , \sice_IBR1_reg[7]/P0001  , \sice_IBR1_reg[8]/P0001  , \sice_IBR1_reg[9]/P0001  , \sice_IBR2_reg[0]/P0001  , \sice_IBR2_reg[10]/P0001  , \sice_IBR2_reg[11]/P0001  , \sice_IBR2_reg[12]/P0001  , \sice_IBR2_reg[13]/P0001  , \sice_IBR2_reg[14]/P0001  , \sice_IBR2_reg[15]/P0001  , \sice_IBR2_reg[16]/P0001  , \sice_IBR2_reg[17]/P0001  , \sice_IBR2_reg[1]/P0001  , \sice_IBR2_reg[2]/P0001  , \sice_IBR2_reg[3]/P0001  , \sice_IBR2_reg[4]/P0001  , \sice_IBR2_reg[5]/P0001  , \sice_IBR2_reg[6]/P0001  , \sice_IBR2_reg[7]/P0001  , \sice_IBR2_reg[8]/P0001  , \sice_IBR2_reg[9]/P0001  , \sice_ICS_reg[0]/NET0131  , \sice_ICS_reg[1]/NET0131  , \sice_ICS_reg[2]/NET0131  , \sice_ICYC_clr_reg/NET0131  , \sice_ICYC_en_reg/NET0131  , \sice_ICYC_en_syn_reg/P0001  , \sice_ICYC_reg[0]/NET0131  , \sice_ICYC_reg[10]/NET0131  , \sice_ICYC_reg[11]/NET0131  , \sice_ICYC_reg[12]/NET0131  , \sice_ICYC_reg[13]/NET0131  , \sice_ICYC_reg[14]/NET0131  , \sice_ICYC_reg[15]/NET0131  , \sice_ICYC_reg[16]/NET0131  , \sice_ICYC_reg[17]/NET0131  , \sice_ICYC_reg[18]/NET0131  , \sice_ICYC_reg[19]/NET0131  , \sice_ICYC_reg[1]/NET0131  , \sice_ICYC_reg[20]/NET0131  , \sice_ICYC_reg[21]/NET0131  , \sice_ICYC_reg[22]/NET0131  , \sice_ICYC_reg[23]/NET0131  , \sice_ICYC_reg[2]/NET0131  , \sice_ICYC_reg[3]/NET0131  , \sice_ICYC_reg[4]/NET0131  , \sice_ICYC_reg[5]/NET0131  , \sice_ICYC_reg[6]/NET0131  , \sice_ICYC_reg[7]/NET0131  , \sice_ICYC_reg[8]/NET0131  , \sice_ICYC_reg[9]/NET0131  , \sice_IDONE_reg/NET0131  , \sice_IIRC_reg[0]/NET0131  , \sice_IIRC_reg[10]/NET0131  , \sice_IIRC_reg[11]/NET0131  , \sice_IIRC_reg[12]/NET0131  , \sice_IIRC_reg[13]/NET0131  , \sice_IIRC_reg[14]/NET0131  , \sice_IIRC_reg[15]/NET0131  , \sice_IIRC_reg[16]/NET0131  , \sice_IIRC_reg[17]/NET0131  , \sice_IIRC_reg[18]/NET0131  , \sice_IIRC_reg[19]/NET0131  , \sice_IIRC_reg[1]/NET0131  , \sice_IIRC_reg[20]/NET0131  , \sice_IIRC_reg[21]/NET0131  , \sice_IIRC_reg[22]/NET0131  , \sice_IIRC_reg[23]/NET0131  , \sice_IIRC_reg[2]/NET0131  , \sice_IIRC_reg[3]/NET0131  , \sice_IIRC_reg[4]/NET0131  , \sice_IIRC_reg[5]/NET0131  , \sice_IIRC_reg[6]/NET0131  , \sice_IIRC_reg[7]/NET0131  , \sice_IIRC_reg[8]/NET0131  , \sice_IIRC_reg[9]/NET0131  , \sice_IMR1_reg[0]/NET0131  , \sice_IMR1_reg[10]/NET0131  , \sice_IMR1_reg[11]/NET0131  , \sice_IMR1_reg[12]/NET0131  , \sice_IMR1_reg[13]/NET0131  , \sice_IMR1_reg[14]/NET0131  , \sice_IMR1_reg[15]/NET0131  , \sice_IMR1_reg[16]/NET0131  , \sice_IMR1_reg[17]/NET0131  , \sice_IMR1_reg[1]/NET0131  , \sice_IMR1_reg[2]/NET0131  , \sice_IMR1_reg[3]/NET0131  , \sice_IMR1_reg[4]/NET0131  , \sice_IMR1_reg[5]/NET0131  , \sice_IMR1_reg[6]/NET0131  , \sice_IMR1_reg[7]/NET0131  , \sice_IMR1_reg[8]/NET0131  , \sice_IMR1_reg[9]/NET0131  , \sice_IMR2_reg[0]/NET0131  , \sice_IMR2_reg[10]/NET0131  , \sice_IMR2_reg[11]/NET0131  , \sice_IMR2_reg[12]/NET0131  , \sice_IMR2_reg[13]/NET0131  , \sice_IMR2_reg[14]/NET0131  , \sice_IMR2_reg[15]/NET0131  , \sice_IMR2_reg[16]/NET0131  , \sice_IMR2_reg[17]/NET0131  , \sice_IMR2_reg[1]/NET0131  , \sice_IMR2_reg[2]/NET0131  , \sice_IMR2_reg[3]/NET0131  , \sice_IMR2_reg[4]/NET0131  , \sice_IMR2_reg[5]/NET0131  , \sice_IMR2_reg[6]/NET0131  , \sice_IMR2_reg[7]/NET0131  , \sice_IMR2_reg[8]/NET0131  , \sice_IMR2_reg[9]/NET0131  , \sice_IRR_reg[0]/P0001  , \sice_IRR_reg[10]/P0001  , \sice_IRR_reg[11]/P0001  , \sice_IRR_reg[12]/P0001  , \sice_IRR_reg[13]/P0001  , \sice_IRR_reg[1]/P0001  , \sice_IRR_reg[2]/P0001  , \sice_IRR_reg[3]/P0001  , \sice_IRR_reg[4]/P0001  , \sice_IRR_reg[5]/P0001  , \sice_IRR_reg[6]/P0001  , \sice_IRR_reg[7]/P0001  , \sice_IRR_reg[8]/P0001  , \sice_IRR_reg[9]/P0001  , \sice_IRST_reg/NET0131  , \sice_IRST_syn_reg/P0001  , \sice_ITR_reg[0]/NET0131  , \sice_ITR_reg[1]/NET0131  , \sice_ITR_reg[2]/NET0131  , \sice_OE_reg/P0001  , \sice_RCS_reg[0]/NET0131  , \sice_RCS_reg[1]/NET0131  , \sice_RST_req_reg/NET0131  , \sice_SPC_reg[0]/P0001  , \sice_SPC_reg[10]/P0001  , \sice_SPC_reg[11]/P0001  , \sice_SPC_reg[12]/P0001  , \sice_SPC_reg[13]/P0001  , \sice_SPC_reg[14]/P0001  , \sice_SPC_reg[15]/P0001  , \sice_SPC_reg[16]/P0001  , \sice_SPC_reg[17]/P0001  , \sice_SPC_reg[18]/P0001  , \sice_SPC_reg[19]/P0001  , \sice_SPC_reg[1]/P0001  , \sice_SPC_reg[20]/P0001  , \sice_SPC_reg[21]/P0001  , \sice_SPC_reg[22]/P0001  , \sice_SPC_reg[23]/P0001  , \sice_SPC_reg[2]/P0001  , \sice_SPC_reg[3]/P0001  , \sice_SPC_reg[4]/P0001  , \sice_SPC_reg[5]/P0001  , \sice_SPC_reg[6]/P0001  , \sice_SPC_reg[7]/P0001  , \sice_SPC_reg[8]/P0001  , \sice_SPC_reg[9]/P0001  , \sice_UpdDR_sd1_reg/P0001  , \sice_UpdDR_sd2_reg/P0001  , \sice_idr0_reg_DO_reg[0]/P0001  , \sice_idr0_reg_DO_reg[10]/P0001  , \sice_idr0_reg_DO_reg[11]/P0001  , \sice_idr0_reg_DO_reg[1]/P0001  , \sice_idr0_reg_DO_reg[2]/P0001  , \sice_idr0_reg_DO_reg[3]/P0001  , \sice_idr0_reg_DO_reg[4]/P0001  , \sice_idr0_reg_DO_reg[5]/P0001  , \sice_idr0_reg_DO_reg[6]/P0001  , \sice_idr0_reg_DO_reg[7]/P0001  , \sice_idr0_reg_DO_reg[8]/P0001  , \sice_idr0_reg_DO_reg[9]/P0001  , \sice_idr1_reg_DO_reg[0]/P0001  , \sice_idr1_reg_DO_reg[10]/P0001  , \sice_idr1_reg_DO_reg[11]/P0001  , \sice_idr1_reg_DO_reg[1]/P0001  , \sice_idr1_reg_DO_reg[2]/P0001  , \sice_idr1_reg_DO_reg[3]/P0001  , \sice_idr1_reg_DO_reg[4]/P0001  , \sice_idr1_reg_DO_reg[5]/P0001  , \sice_idr1_reg_DO_reg[6]/P0001  , \sice_idr1_reg_DO_reg[7]/P0001  , \sice_idr1_reg_DO_reg[8]/P0001  , \sice_idr1_reg_DO_reg[9]/P0001  , \sport0_cfg_FSi_cnt_reg[0]/NET0131  , \sport0_cfg_FSi_cnt_reg[10]/NET0131  , \sport0_cfg_FSi_cnt_reg[11]/NET0131  , \sport0_cfg_FSi_cnt_reg[12]/NET0131  , \sport0_cfg_FSi_cnt_reg[13]/NET0131  , \sport0_cfg_FSi_cnt_reg[14]/NET0131  , \sport0_cfg_FSi_cnt_reg[15]/NET0131  , \sport0_cfg_FSi_cnt_reg[1]/NET0131  , \sport0_cfg_FSi_cnt_reg[2]/NET0131  , \sport0_cfg_FSi_cnt_reg[3]/NET0131  , \sport0_cfg_FSi_cnt_reg[4]/NET0131  , \sport0_cfg_FSi_cnt_reg[5]/NET0131  , \sport0_cfg_FSi_cnt_reg[6]/NET0131  , \sport0_cfg_FSi_cnt_reg[7]/NET0131  , \sport0_cfg_FSi_cnt_reg[8]/NET0131  , \sport0_cfg_FSi_cnt_reg[9]/NET0131  , \sport0_cfg_FSi_reg/NET0131  , \sport0_cfg_RFSg_d1_reg/NET0131  , \sport0_cfg_RFSg_d2_reg/NET0131  , \sport0_cfg_RFSg_d3_reg/NET0131  , \sport0_cfg_RFSgi_d_reg/NET0131  , \sport0_cfg_SCLKi_cnt_reg[0]/NET0131  , \sport0_cfg_SCLKi_cnt_reg[10]/NET0131  , \sport0_cfg_SCLKi_cnt_reg[11]/NET0131  , \sport0_cfg_SCLKi_cnt_reg[12]/NET0131  , \sport0_cfg_SCLKi_cnt_reg[13]/NET0131  , \sport0_cfg_SCLKi_cnt_reg[14]/NET0131  , \sport0_cfg_SCLKi_cnt_reg[15]/NET0131  , \sport0_cfg_SCLKi_cnt_reg[1]/NET0131  , \sport0_cfg_SCLKi_cnt_reg[2]/NET0131  , \sport0_cfg_SCLKi_cnt_reg[3]/NET0131  , \sport0_cfg_SCLKi_cnt_reg[4]/NET0131  , \sport0_cfg_SCLKi_cnt_reg[5]/NET0131  , \sport0_cfg_SCLKi_cnt_reg[6]/NET0131  , \sport0_cfg_SCLKi_cnt_reg[7]/NET0131  , \sport0_cfg_SCLKi_cnt_reg[8]/NET0131  , \sport0_cfg_SCLKi_cnt_reg[9]/NET0131  , \sport0_cfg_SCLKi_h_reg/NET0131  , \sport0_cfg_SP_ENg_D1_reg/P0001  , \sport0_cfg_SP_ENg_reg/NET0131  , \sport0_cfg_TFSg_d1_reg/NET0131  , \sport0_cfg_TFSg_d2_reg/NET0131  , \sport0_cfg_TFSg_d3_reg/NET0131  , \sport0_cfg_TFSgi_d_reg/NET0131  , \sport0_regs_AUTO_a_reg[12]/NET0131  , \sport0_regs_AUTO_a_reg[13]/NET0131  , \sport0_regs_AUTO_a_reg[14]/NET0131  , \sport0_regs_AUTO_a_reg[15]/NET0131  , \sport0_regs_AUTOreg_DO_reg[0]/NET0131  , \sport0_regs_AUTOreg_DO_reg[10]/NET0131  , \sport0_regs_AUTOreg_DO_reg[11]/NET0131  , \sport0_regs_AUTOreg_DO_reg[1]/NET0131  , \sport0_regs_AUTOreg_DO_reg[2]/NET0131  , \sport0_regs_AUTOreg_DO_reg[3]/NET0131  , \sport0_regs_AUTOreg_DO_reg[4]/NET0131  , \sport0_regs_AUTOreg_DO_reg[5]/NET0131  , \sport0_regs_AUTOreg_DO_reg[6]/NET0131  , \sport0_regs_AUTOreg_DO_reg[7]/NET0131  , \sport0_regs_AUTOreg_DO_reg[8]/NET0131  , \sport0_regs_AUTOreg_DO_reg[9]/NET0131  , \sport0_regs_FSDIVreg_DO_reg[0]/NET0131  , \sport0_regs_FSDIVreg_DO_reg[10]/NET0131  , \sport0_regs_FSDIVreg_DO_reg[11]/NET0131  , \sport0_regs_FSDIVreg_DO_reg[12]/NET0131  , \sport0_regs_FSDIVreg_DO_reg[13]/NET0131  , \sport0_regs_FSDIVreg_DO_reg[14]/NET0131  , \sport0_regs_FSDIVreg_DO_reg[15]/NET0131  , \sport0_regs_FSDIVreg_DO_reg[1]/NET0131  , \sport0_regs_FSDIVreg_DO_reg[2]/NET0131  , \sport0_regs_FSDIVreg_DO_reg[3]/NET0131  , \sport0_regs_FSDIVreg_DO_reg[4]/NET0131  , \sport0_regs_FSDIVreg_DO_reg[5]/NET0131  , \sport0_regs_FSDIVreg_DO_reg[6]/NET0131  , \sport0_regs_FSDIVreg_DO_reg[7]/NET0131  , \sport0_regs_FSDIVreg_DO_reg[8]/NET0131  , \sport0_regs_FSDIVreg_DO_reg[9]/NET0131  , \sport0_regs_MWORDreg_DO_reg[0]/NET0131  , \sport0_regs_MWORDreg_DO_reg[10]/NET0131  , \sport0_regs_MWORDreg_DO_reg[1]/NET0131  , \sport0_regs_MWORDreg_DO_reg[2]/NET0131  , \sport0_regs_MWORDreg_DO_reg[3]/NET0131  , \sport0_regs_MWORDreg_DO_reg[4]/NET0131  , \sport0_regs_MWORDreg_DO_reg[5]/NET0131  , \sport0_regs_MWORDreg_DO_reg[6]/NET0131  , \sport0_regs_MWORDreg_DO_reg[7]/NET0131  , \sport0_regs_MWORDreg_DO_reg[8]/NET0131  , \sport0_regs_MWORDreg_DO_reg[9]/NET0131  , \sport0_regs_SCLKDIVreg_DO_reg[0]/NET0131  , \sport0_regs_SCLKDIVreg_DO_reg[10]/NET0131  , \sport0_regs_SCLKDIVreg_DO_reg[11]/NET0131  , \sport0_regs_SCLKDIVreg_DO_reg[12]/NET0131  , \sport0_regs_SCLKDIVreg_DO_reg[13]/NET0131  , \sport0_regs_SCLKDIVreg_DO_reg[14]/NET0131  , \sport0_regs_SCLKDIVreg_DO_reg[15]/NET0131  , \sport0_regs_SCLKDIVreg_DO_reg[1]/NET0131  , \sport0_regs_SCLKDIVreg_DO_reg[2]/NET0131  , \sport0_regs_SCLKDIVreg_DO_reg[3]/NET0131  , \sport0_regs_SCLKDIVreg_DO_reg[4]/NET0131  , \sport0_regs_SCLKDIVreg_DO_reg[5]/NET0131  , \sport0_regs_SCLKDIVreg_DO_reg[6]/NET0131  , \sport0_regs_SCLKDIVreg_DO_reg[7]/NET0131  , \sport0_regs_SCLKDIVreg_DO_reg[8]/NET0131  , \sport0_regs_SCLKDIVreg_DO_reg[9]/NET0131  , \sport0_regs_SCTLreg_DO_reg[0]/NET0131  , \sport0_regs_SCTLreg_DO_reg[10]/NET0131  , \sport0_regs_SCTLreg_DO_reg[11]/NET0131  , \sport0_regs_SCTLreg_DO_reg[12]/NET0131  , \sport0_regs_SCTLreg_DO_reg[13]/NET0131  , \sport0_regs_SCTLreg_DO_reg[15]/NET0131  , \sport0_regs_SCTLreg_DO_reg[1]/NET0131  , \sport0_regs_SCTLreg_DO_reg[2]/NET0131  , \sport0_regs_SCTLreg_DO_reg[3]/NET0131  , \sport0_regs_SCTLreg_DO_reg[4]/NET0131  , \sport0_regs_SCTLreg_DO_reg[5]/NET0131  , \sport0_regs_SCTLreg_DO_reg[6]/NET0131  , \sport0_regs_SCTLreg_DO_reg[7]/NET0131  , \sport0_rxctl_Bcnt_reg[0]/NET0131  , \sport0_rxctl_Bcnt_reg[1]/NET0131  , \sport0_rxctl_Bcnt_reg[2]/NET0131  , \sport0_rxctl_Bcnt_reg[3]/NET0131  , \sport0_rxctl_Bcnt_reg[4]/NET0131  , \sport0_rxctl_ISRa_reg/P0001  , \sport0_rxctl_LMcnt_reg[0]/NET0131  , \sport0_rxctl_LMcnt_reg[1]/NET0131  , \sport0_rxctl_LMcnt_reg[2]/NET0131  , \sport0_rxctl_LMcnt_reg[3]/NET0131  , \sport0_rxctl_LMcnt_reg[4]/NET0131  , \sport0_rxctl_RCS_reg[0]/NET0131  , \sport0_rxctl_RCS_reg[1]/NET0131  , \sport0_rxctl_RCS_reg[2]/NET0131  , \sport0_rxctl_RSreq_reg/NET0131  , \sport0_rxctl_RXSHT_reg[0]/P0001  , \sport0_rxctl_RXSHT_reg[10]/P0001  , \sport0_rxctl_RXSHT_reg[11]/P0001  , \sport0_rxctl_RXSHT_reg[12]/P0001  , \sport0_rxctl_RXSHT_reg[13]/P0001  , \sport0_rxctl_RXSHT_reg[14]/P0001  , \sport0_rxctl_RXSHT_reg[15]/P0001  , \sport0_rxctl_RXSHT_reg[1]/P0001  , \sport0_rxctl_RXSHT_reg[2]/P0001  , \sport0_rxctl_RXSHT_reg[3]/P0001  , \sport0_rxctl_RXSHT_reg[4]/P0001  , \sport0_rxctl_RXSHT_reg[5]/P0001  , \sport0_rxctl_RXSHT_reg[6]/P0001  , \sport0_rxctl_RXSHT_reg[7]/P0001  , \sport0_rxctl_RXSHT_reg[8]/P0001  , \sport0_rxctl_RXSHT_reg[9]/P0001  , \sport0_rxctl_RX_reg[0]/P0001  , \sport0_rxctl_RX_reg[10]/P0001  , \sport0_rxctl_RX_reg[11]/P0001  , \sport0_rxctl_RX_reg[12]/P0001  , \sport0_rxctl_RX_reg[13]/P0001  , \sport0_rxctl_RX_reg[14]/P0001  , \sport0_rxctl_RX_reg[15]/P0001  , \sport0_rxctl_RX_reg[1]/P0001  , \sport0_rxctl_RX_reg[2]/P0001  , \sport0_rxctl_RX_reg[3]/P0001  , \sport0_rxctl_RX_reg[4]/P0001  , \sport0_rxctl_RX_reg[5]/P0001  , \sport0_rxctl_RX_reg[6]/P0001  , \sport0_rxctl_RX_reg[7]/P0001  , \sport0_rxctl_RX_reg[8]/P0001  , \sport0_rxctl_RX_reg[9]/P0001  , \sport0_rxctl_SLOT1_EXT_reg[2]/NET0131  , \sport0_rxctl_SLOT1_EXT_reg[3]/NET0131  , \sport0_rxctl_TAG_SLOT_reg/P0001  , \sport0_rxctl_Wcnt_reg[0]/NET0131  , \sport0_rxctl_Wcnt_reg[1]/NET0131  , \sport0_rxctl_Wcnt_reg[2]/NET0131  , \sport0_rxctl_Wcnt_reg[3]/NET0131  , \sport0_rxctl_Wcnt_reg[4]/NET0131  , \sport0_rxctl_Wcnt_reg[5]/NET0131  , \sport0_rxctl_Wcnt_reg[6]/NET0131  , \sport0_rxctl_Wcnt_reg[7]/NET0131  , \sport0_rxctl_a_sync1_reg/P0001  , \sport0_rxctl_a_sync2_reg/P0001  , \sport0_rxctl_ldRX_cmp_reg/P0001  , \sport0_rxctl_sht2nd_reg/P0001  , \sport0_txctl_Bcnt_reg[0]/NET0131  , \sport0_txctl_Bcnt_reg[1]/NET0131  , \sport0_txctl_Bcnt_reg[2]/NET0131  , \sport0_txctl_Bcnt_reg[3]/NET0131  , \sport0_txctl_Bcnt_reg[4]/NET0131  , \sport0_txctl_SP_EN_D1_reg/P0001  , \sport0_txctl_TCS_reg[0]/NET0131  , \sport0_txctl_TCS_reg[1]/NET0131  , \sport0_txctl_TCS_reg[2]/NET0131  , \sport0_txctl_TSreq_reg/NET0131  , \sport0_txctl_TSreqi_reg/NET0131  , \sport0_txctl_TXSHT_reg[0]/P0001  , \sport0_txctl_TXSHT_reg[10]/P0001  , \sport0_txctl_TXSHT_reg[11]/P0001  , \sport0_txctl_TXSHT_reg[12]/P0001  , \sport0_txctl_TXSHT_reg[13]/P0001  , \sport0_txctl_TXSHT_reg[14]/P0001  , \sport0_txctl_TXSHT_reg[15]/P0001  , \sport0_txctl_TXSHT_reg[1]/P0001  , \sport0_txctl_TXSHT_reg[2]/P0001  , \sport0_txctl_TXSHT_reg[3]/P0001  , \sport0_txctl_TXSHT_reg[4]/P0001  , \sport0_txctl_TXSHT_reg[5]/P0001  , \sport0_txctl_TXSHT_reg[6]/P0001  , \sport0_txctl_TXSHT_reg[7]/P0001  , \sport0_txctl_TXSHT_reg[8]/P0001  , \sport0_txctl_TXSHT_reg[9]/P0001  , \sport0_txctl_TX_reg[0]/P0001  , \sport0_txctl_TX_reg[10]/P0001  , \sport0_txctl_TX_reg[11]/P0001  , \sport0_txctl_TX_reg[12]/P0001  , \sport0_txctl_TX_reg[13]/P0001  , \sport0_txctl_TX_reg[14]/P0001  , \sport0_txctl_TX_reg[15]/P0001  , \sport0_txctl_TX_reg[1]/P0001  , \sport0_txctl_TX_reg[2]/P0001  , \sport0_txctl_TX_reg[3]/P0001  , \sport0_txctl_TX_reg[4]/P0001  , \sport0_txctl_TX_reg[5]/P0001  , \sport0_txctl_TX_reg[6]/P0001  , \sport0_txctl_TX_reg[7]/P0001  , \sport0_txctl_TX_reg[8]/P0001  , \sport0_txctl_TX_reg[9]/P0001  , \sport0_txctl_Wcnt_reg[0]/NET0131  , \sport0_txctl_Wcnt_reg[1]/NET0131  , \sport0_txctl_Wcnt_reg[2]/NET0131  , \sport0_txctl_Wcnt_reg[3]/NET0131  , \sport0_txctl_Wcnt_reg[4]/NET0131  , \sport0_txctl_Wcnt_reg[5]/NET0131  , \sport0_txctl_Wcnt_reg[6]/NET0131  , \sport0_txctl_Wcnt_reg[7]/NET0131  , \sport0_txctl_b_sync1_reg/P0001  , \sport0_txctl_c_sync1_reg/P0001  , \sport0_txctl_c_sync2_reg/P0001  , \sport0_txctl_ldTX_cmp_reg/P0001  , \sport1_cfg_FSi_cnt_reg[0]/NET0131  , \sport1_cfg_FSi_cnt_reg[10]/NET0131  , \sport1_cfg_FSi_cnt_reg[11]/NET0131  , \sport1_cfg_FSi_cnt_reg[12]/NET0131  , \sport1_cfg_FSi_cnt_reg[13]/NET0131  , \sport1_cfg_FSi_cnt_reg[14]/NET0131  , \sport1_cfg_FSi_cnt_reg[15]/NET0131  , \sport1_cfg_FSi_cnt_reg[1]/NET0131  , \sport1_cfg_FSi_cnt_reg[2]/NET0131  , \sport1_cfg_FSi_cnt_reg[3]/NET0131  , \sport1_cfg_FSi_cnt_reg[4]/NET0131  , \sport1_cfg_FSi_cnt_reg[5]/NET0131  , \sport1_cfg_FSi_cnt_reg[6]/NET0131  , \sport1_cfg_FSi_cnt_reg[7]/NET0131  , \sport1_cfg_FSi_cnt_reg[8]/NET0131  , \sport1_cfg_FSi_cnt_reg[9]/NET0131  , \sport1_cfg_FSi_reg/NET0131  , \sport1_cfg_RFSg_d1_reg/NET0131  , \sport1_cfg_RFSg_d2_reg/NET0131  , \sport1_cfg_RFSg_d3_reg/NET0131  , \sport1_cfg_RFSgi_d_reg/NET0131  , \sport1_cfg_SCLKi_cnt_reg[0]/NET0131  , \sport1_cfg_SCLKi_cnt_reg[10]/NET0131  , \sport1_cfg_SCLKi_cnt_reg[11]/NET0131  , \sport1_cfg_SCLKi_cnt_reg[12]/NET0131  , \sport1_cfg_SCLKi_cnt_reg[13]/NET0131  , \sport1_cfg_SCLKi_cnt_reg[14]/NET0131  , \sport1_cfg_SCLKi_cnt_reg[15]/NET0131  , \sport1_cfg_SCLKi_cnt_reg[1]/NET0131  , \sport1_cfg_SCLKi_cnt_reg[2]/NET0131  , \sport1_cfg_SCLKi_cnt_reg[3]/NET0131  , \sport1_cfg_SCLKi_cnt_reg[4]/NET0131  , \sport1_cfg_SCLKi_cnt_reg[5]/NET0131  , \sport1_cfg_SCLKi_cnt_reg[6]/NET0131  , \sport1_cfg_SCLKi_cnt_reg[7]/NET0131  , \sport1_cfg_SCLKi_cnt_reg[8]/NET0131  , \sport1_cfg_SCLKi_cnt_reg[9]/NET0131  , \sport1_cfg_SCLKi_h_reg/NET0131  , \sport1_cfg_SP_ENg_D1_reg/P0001  , \sport1_cfg_SP_ENg_reg/NET0131  , \sport1_cfg_TFSg_d1_reg/NET0131  , \sport1_cfg_TFSg_d2_reg/NET0131  , \sport1_cfg_TFSg_d3_reg/NET0131  , \sport1_cfg_TFSgi_d_reg/NET0131  , \sport1_regs_AUTOreg_DO_reg[0]/NET0131  , \sport1_regs_AUTOreg_DO_reg[10]/NET0131  , \sport1_regs_AUTOreg_DO_reg[11]/NET0131  , \sport1_regs_AUTOreg_DO_reg[1]/NET0131  , \sport1_regs_AUTOreg_DO_reg[2]/NET0131  , \sport1_regs_AUTOreg_DO_reg[3]/NET0131  , \sport1_regs_AUTOreg_DO_reg[4]/NET0131  , \sport1_regs_AUTOreg_DO_reg[5]/NET0131  , \sport1_regs_AUTOreg_DO_reg[6]/NET0131  , \sport1_regs_AUTOreg_DO_reg[7]/NET0131  , \sport1_regs_AUTOreg_DO_reg[8]/NET0131  , \sport1_regs_AUTOreg_DO_reg[9]/NET0131  , \sport1_regs_FSDIVreg_DO_reg[0]/NET0131  , \sport1_regs_FSDIVreg_DO_reg[10]/NET0131  , \sport1_regs_FSDIVreg_DO_reg[11]/NET0131  , \sport1_regs_FSDIVreg_DO_reg[12]/NET0131  , \sport1_regs_FSDIVreg_DO_reg[13]/NET0131  , \sport1_regs_FSDIVreg_DO_reg[14]/NET0131  , \sport1_regs_FSDIVreg_DO_reg[15]/NET0131  , \sport1_regs_FSDIVreg_DO_reg[1]/NET0131  , \sport1_regs_FSDIVreg_DO_reg[2]/NET0131  , \sport1_regs_FSDIVreg_DO_reg[3]/NET0131  , \sport1_regs_FSDIVreg_DO_reg[4]/NET0131  , \sport1_regs_FSDIVreg_DO_reg[5]/NET0131  , \sport1_regs_FSDIVreg_DO_reg[6]/NET0131  , \sport1_regs_FSDIVreg_DO_reg[7]/NET0131  , \sport1_regs_FSDIVreg_DO_reg[8]/NET0131  , \sport1_regs_FSDIVreg_DO_reg[9]/NET0131  , \sport1_regs_MWORDreg_DO_reg[0]/NET0131  , \sport1_regs_MWORDreg_DO_reg[10]/NET0131  , \sport1_regs_MWORDreg_DO_reg[1]/NET0131  , \sport1_regs_MWORDreg_DO_reg[2]/NET0131  , \sport1_regs_MWORDreg_DO_reg[3]/NET0131  , \sport1_regs_MWORDreg_DO_reg[4]/NET0131  , \sport1_regs_MWORDreg_DO_reg[5]/NET0131  , \sport1_regs_MWORDreg_DO_reg[6]/NET0131  , \sport1_regs_MWORDreg_DO_reg[7]/NET0131  , \sport1_regs_MWORDreg_DO_reg[8]/NET0131  , \sport1_regs_MWORDreg_DO_reg[9]/NET0131  , \sport1_regs_SCLKDIVreg_DO_reg[0]/NET0131  , \sport1_regs_SCLKDIVreg_DO_reg[10]/NET0131  , \sport1_regs_SCLKDIVreg_DO_reg[11]/NET0131  , \sport1_regs_SCLKDIVreg_DO_reg[12]/NET0131  , \sport1_regs_SCLKDIVreg_DO_reg[13]/NET0131  , \sport1_regs_SCLKDIVreg_DO_reg[14]/NET0131  , \sport1_regs_SCLKDIVreg_DO_reg[15]/NET0131  , \sport1_regs_SCLKDIVreg_DO_reg[1]/NET0131  , \sport1_regs_SCLKDIVreg_DO_reg[2]/NET0131  , \sport1_regs_SCLKDIVreg_DO_reg[3]/NET0131  , \sport1_regs_SCLKDIVreg_DO_reg[4]/NET0131  , \sport1_regs_SCLKDIVreg_DO_reg[5]/NET0131  , \sport1_regs_SCLKDIVreg_DO_reg[6]/NET0131  , \sport1_regs_SCLKDIVreg_DO_reg[7]/NET0131  , \sport1_regs_SCLKDIVreg_DO_reg[8]/NET0131  , \sport1_regs_SCLKDIVreg_DO_reg[9]/NET0131  , \sport1_regs_SCTLreg_DO_reg[0]/NET0131  , \sport1_regs_SCTLreg_DO_reg[10]/NET0131  , \sport1_regs_SCTLreg_DO_reg[11]/NET0131  , \sport1_regs_SCTLreg_DO_reg[12]/NET0131  , \sport1_regs_SCTLreg_DO_reg[13]/NET0131  , \sport1_regs_SCTLreg_DO_reg[15]/NET0131  , \sport1_regs_SCTLreg_DO_reg[1]/NET0131  , \sport1_regs_SCTLreg_DO_reg[2]/NET0131  , \sport1_regs_SCTLreg_DO_reg[3]/NET0131  , \sport1_regs_SCTLreg_DO_reg[4]/NET0131  , \sport1_regs_SCTLreg_DO_reg[5]/NET0131  , \sport1_regs_SCTLreg_DO_reg[6]/NET0131  , \sport1_regs_SCTLreg_DO_reg[7]/NET0131  , \sport1_rxctl_Bcnt_reg[0]/NET0131  , \sport1_rxctl_Bcnt_reg[1]/NET0131  , \sport1_rxctl_Bcnt_reg[2]/NET0131  , \sport1_rxctl_Bcnt_reg[3]/NET0131  , \sport1_rxctl_Bcnt_reg[4]/NET0131  , \sport1_rxctl_ISRa_reg/P0001  , \sport1_rxctl_LMcnt_reg[0]/NET0131  , \sport1_rxctl_LMcnt_reg[1]/NET0131  , \sport1_rxctl_LMcnt_reg[2]/NET0131  , \sport1_rxctl_LMcnt_reg[3]/NET0131  , \sport1_rxctl_LMcnt_reg[4]/NET0131  , \sport1_rxctl_RCS_reg[0]/NET0131  , \sport1_rxctl_RCS_reg[1]/NET0131  , \sport1_rxctl_RCS_reg[2]/NET0131  , \sport1_rxctl_RSreq_reg/NET0131  , \sport1_rxctl_RXSHT_reg[0]/P0001  , \sport1_rxctl_RXSHT_reg[10]/P0001  , \sport1_rxctl_RXSHT_reg[11]/P0001  , \sport1_rxctl_RXSHT_reg[12]/P0001  , \sport1_rxctl_RXSHT_reg[13]/P0001  , \sport1_rxctl_RXSHT_reg[14]/P0001  , \sport1_rxctl_RXSHT_reg[15]/P0001  , \sport1_rxctl_RXSHT_reg[1]/P0001  , \sport1_rxctl_RXSHT_reg[2]/P0001  , \sport1_rxctl_RXSHT_reg[3]/P0001  , \sport1_rxctl_RXSHT_reg[4]/P0001  , \sport1_rxctl_RXSHT_reg[5]/P0001  , \sport1_rxctl_RXSHT_reg[6]/P0001  , \sport1_rxctl_RXSHT_reg[7]/P0001  , \sport1_rxctl_RXSHT_reg[8]/P0001  , \sport1_rxctl_RXSHT_reg[9]/P0001  , \sport1_rxctl_RX_reg[0]/P0001  , \sport1_rxctl_RX_reg[10]/P0001  , \sport1_rxctl_RX_reg[11]/P0001  , \sport1_rxctl_RX_reg[12]/P0001  , \sport1_rxctl_RX_reg[13]/P0001  , \sport1_rxctl_RX_reg[14]/P0001  , \sport1_rxctl_RX_reg[15]/P0001  , \sport1_rxctl_RX_reg[1]/P0001  , \sport1_rxctl_RX_reg[2]/P0001  , \sport1_rxctl_RX_reg[3]/P0001  , \sport1_rxctl_RX_reg[4]/P0001  , \sport1_rxctl_RX_reg[5]/P0001  , \sport1_rxctl_RX_reg[6]/P0001  , \sport1_rxctl_RX_reg[7]/P0001  , \sport1_rxctl_RX_reg[8]/P0001  , \sport1_rxctl_RX_reg[9]/P0001  , \sport1_rxctl_SLOT1_EXT_reg[2]/NET0131  , \sport1_rxctl_SLOT1_EXT_reg[3]/NET0131  , \sport1_rxctl_TAG_SLOT_reg/P0001  , \sport1_rxctl_Wcnt_reg[0]/NET0131  , \sport1_rxctl_Wcnt_reg[1]/NET0131  , \sport1_rxctl_Wcnt_reg[2]/NET0131  , \sport1_rxctl_Wcnt_reg[3]/NET0131  , \sport1_rxctl_Wcnt_reg[4]/NET0131  , \sport1_rxctl_Wcnt_reg[5]/NET0131  , \sport1_rxctl_Wcnt_reg[6]/NET0131  , \sport1_rxctl_Wcnt_reg[7]/NET0131  , \sport1_rxctl_a_sync1_reg/P0001  , \sport1_rxctl_a_sync2_reg/P0001  , \sport1_rxctl_sht2nd_reg/P0001  , \sport1_txctl_Bcnt_reg[0]/NET0131  , \sport1_txctl_Bcnt_reg[1]/NET0131  , \sport1_txctl_Bcnt_reg[2]/NET0131  , \sport1_txctl_Bcnt_reg[3]/NET0131  , \sport1_txctl_Bcnt_reg[4]/NET0131  , \sport1_txctl_SP_EN_D1_reg/P0001  , \sport1_txctl_TCS_reg[0]/NET0131  , \sport1_txctl_TCS_reg[1]/NET0131  , \sport1_txctl_TCS_reg[2]/NET0131  , \sport1_txctl_TSreq_reg/NET0131  , \sport1_txctl_TSreqi_reg/NET0131  , \sport1_txctl_TXSHT_reg[0]/P0001  , \sport1_txctl_TXSHT_reg[10]/P0001  , \sport1_txctl_TXSHT_reg[11]/P0001  , \sport1_txctl_TXSHT_reg[12]/P0001  , \sport1_txctl_TXSHT_reg[13]/P0001  , \sport1_txctl_TXSHT_reg[14]/P0001  , \sport1_txctl_TXSHT_reg[15]/P0001  , \sport1_txctl_TXSHT_reg[1]/P0001  , \sport1_txctl_TXSHT_reg[2]/P0001  , \sport1_txctl_TXSHT_reg[3]/P0001  , \sport1_txctl_TXSHT_reg[4]/P0001  , \sport1_txctl_TXSHT_reg[5]/P0001  , \sport1_txctl_TXSHT_reg[6]/P0001  , \sport1_txctl_TXSHT_reg[7]/P0001  , \sport1_txctl_TXSHT_reg[8]/P0001  , \sport1_txctl_TXSHT_reg[9]/P0001  , \sport1_txctl_TX_reg[0]/P0001  , \sport1_txctl_TX_reg[10]/P0001  , \sport1_txctl_TX_reg[11]/P0001  , \sport1_txctl_TX_reg[12]/P0001  , \sport1_txctl_TX_reg[13]/P0001  , \sport1_txctl_TX_reg[14]/P0001  , \sport1_txctl_TX_reg[15]/P0001  , \sport1_txctl_TX_reg[1]/P0001  , \sport1_txctl_TX_reg[2]/P0001  , \sport1_txctl_TX_reg[3]/P0001  , \sport1_txctl_TX_reg[4]/P0001  , \sport1_txctl_TX_reg[5]/P0001  , \sport1_txctl_TX_reg[6]/P0001  , \sport1_txctl_TX_reg[7]/P0001  , \sport1_txctl_TX_reg[8]/P0001  , \sport1_txctl_TX_reg[9]/P0001  , \sport1_txctl_Wcnt_reg[0]/NET0131  , \sport1_txctl_Wcnt_reg[1]/NET0131  , \sport1_txctl_Wcnt_reg[2]/NET0131  , \sport1_txctl_Wcnt_reg[3]/NET0131  , \sport1_txctl_Wcnt_reg[4]/NET0131  , \sport1_txctl_Wcnt_reg[5]/NET0131  , \sport1_txctl_Wcnt_reg[6]/NET0131  , \sport1_txctl_Wcnt_reg[7]/NET0131  , \sport1_txctl_c_sync1_reg/P0001  , \sport1_txctl_c_sync2_reg/P0001  , \tm_MSTAT5_syn_reg/NET0131  , \tm_TCR_TMP_reg[0]/NET0131  , \tm_TCR_TMP_reg[10]/NET0131  , \tm_TCR_TMP_reg[11]/NET0131  , \tm_TCR_TMP_reg[12]/NET0131  , \tm_TCR_TMP_reg[13]/NET0131  , \tm_TCR_TMP_reg[14]/NET0131  , \tm_TCR_TMP_reg[15]/NET0131  , \tm_TCR_TMP_reg[1]/NET0131  , \tm_TCR_TMP_reg[2]/NET0131  , \tm_TCR_TMP_reg[3]/NET0131  , \tm_TCR_TMP_reg[4]/NET0131  , \tm_TCR_TMP_reg[5]/NET0131  , \tm_TCR_TMP_reg[6]/NET0131  , \tm_TCR_TMP_reg[7]/NET0131  , \tm_TCR_TMP_reg[8]/NET0131  , \tm_TCR_TMP_reg[9]/NET0131  , \tm_TINT_GEN1_reg/NET0131  , \tm_TINT_GEN2_reg/NET0131  , \tm_TSR_TMP_reg[0]/NET0131  , \tm_TSR_TMP_reg[1]/NET0131  , \tm_TSR_TMP_reg[2]/NET0131  , \tm_TSR_TMP_reg[3]/NET0131  , \tm_TSR_TMP_reg[4]/NET0131  , \tm_TSR_TMP_reg[5]/NET0131  , \tm_TSR_TMP_reg[6]/NET0131  , \tm_TSR_TMP_reg[7]/NET0131  , \tm_WR_TCR_KEEP_TO_TMCLK_p_reg/NET0131  , \tm_WR_TCR_TMP_GEN1_reg/P0001  , \tm_WR_TCR_TMP_GEN2_reg/P0001  , \tm_WR_TCR_p_reg/P0001  , \tm_WR_TSR_KEEP_TO_TMCLK_p_reg/NET0131  , \tm_WR_TSR_TMP_GEN1_reg/P0001  , \tm_WR_TSR_TMP_GEN2_reg/P0001  , \tm_WR_TSR_p_reg/P0001  , \tm_tcr_reg_DO_reg[0]/NET0131  , \tm_tcr_reg_DO_reg[10]/NET0131  , \tm_tcr_reg_DO_reg[11]/NET0131  , \tm_tcr_reg_DO_reg[12]/NET0131  , \tm_tcr_reg_DO_reg[13]/NET0131  , \tm_tcr_reg_DO_reg[14]/NET0131  , \tm_tcr_reg_DO_reg[15]/NET0131  , \tm_tcr_reg_DO_reg[1]/NET0131  , \tm_tcr_reg_DO_reg[2]/NET0131  , \tm_tcr_reg_DO_reg[3]/NET0131  , \tm_tcr_reg_DO_reg[4]/NET0131  , \tm_tcr_reg_DO_reg[5]/NET0131  , \tm_tcr_reg_DO_reg[6]/NET0131  , \tm_tcr_reg_DO_reg[7]/NET0131  , \tm_tcr_reg_DO_reg[8]/NET0131  , \tm_tcr_reg_DO_reg[9]/NET0131  , \tm_tpr_reg_DO_reg[0]/NET0131  , \tm_tpr_reg_DO_reg[10]/NET0131  , \tm_tpr_reg_DO_reg[11]/NET0131  , \tm_tpr_reg_DO_reg[12]/NET0131  , \tm_tpr_reg_DO_reg[13]/NET0131  , \tm_tpr_reg_DO_reg[14]/NET0131  , \tm_tpr_reg_DO_reg[15]/NET0131  , \tm_tpr_reg_DO_reg[1]/NET0131  , \tm_tpr_reg_DO_reg[2]/NET0131  , \tm_tpr_reg_DO_reg[3]/NET0131  , \tm_tpr_reg_DO_reg[4]/NET0131  , \tm_tpr_reg_DO_reg[5]/NET0131  , \tm_tpr_reg_DO_reg[6]/NET0131  , \tm_tpr_reg_DO_reg[7]/NET0131  , \tm_tpr_reg_DO_reg[8]/NET0131  , \tm_tpr_reg_DO_reg[9]/NET0131  , \tm_tsr_reg_DO_reg[0]/NET0131  , \tm_tsr_reg_DO_reg[1]/NET0131  , \tm_tsr_reg_DO_reg[2]/NET0131  , \tm_tsr_reg_DO_reg[3]/NET0131  , \tm_tsr_reg_DO_reg[4]/NET0131  , \tm_tsr_reg_DO_reg[5]/NET0131  , \tm_tsr_reg_DO_reg[6]/NET0131  , \tm_tsr_reg_DO_reg[7]/NET0131  , \tm_tsr_reg_DO_reg[8]/NET0131  , CLKO_pad , \CMAinx[0]_pad  , \CMAinx[10]_pad  , \CMAinx[11]_pad  , \CMAinx[1]_pad  , \CMAinx[2]_pad  , \CMAinx[3]_pad  , \CMAinx[4]_pad  , \CMAinx[5]_pad  , \CMAinx[6]_pad  , \CMAinx[7]_pad  , \CMAinx[8]_pad  , \CMAinx[9]_pad  , CMSn_pad , CM_cs_pad , \CM_wd[0]_pad  , \CM_wd[10]_pad  , \CM_wd[11]_pad  , \CM_wd[12]_pad  , \CM_wd[13]_pad  , \CM_wd[14]_pad  , \CM_wd[15]_pad  , \CM_wd[16]_pad  , \CM_wd[17]_pad  , \CM_wd[18]_pad  , \CM_wd[19]_pad  , \CM_wd[1]_pad  , \CM_wd[20]_pad  , \CM_wd[21]_pad  , \CM_wd[22]_pad  , \CM_wd[23]_pad  , \CM_wd[2]_pad  , \CM_wd[3]_pad  , \CM_wd[4]_pad  , \CM_wd[5]_pad  , \CM_wd[6]_pad  , \CM_wd[7]_pad  , \CM_wd[8]_pad  , \CM_wd[9]_pad  , CM_web_pad , \CMo_cs0_pad  , \CMo_cs1_pad  , \CMo_cs2_pad  , \CMo_cs3_pad  , \CMo_cs4_pad  , \CMo_cs5_pad  , \CMo_cs6_pad  , \CMo_cs7_pad  , \DMAinx[0]_pad  , \DMAinx[10]_pad  , \DMAinx[11]_pad  , \DMAinx[12]_pad  , \DMAinx[13]_pad  , \DMAinx[1]_pad  , \DMAinx[2]_pad  , \DMAinx[3]_pad  , \DMAinx[4]_pad  , \DMAinx[5]_pad  , \DMAinx[6]_pad  , \DMAinx[7]_pad  , \DMAinx[8]_pad  , \DMAinx[9]_pad  , DMSn_pad , DM_cs_pad , \DM_wd[0]_pad  , \DM_wd[10]_pad  , \DM_wd[11]_pad  , \DM_wd[12]_pad  , \DM_wd[13]_pad  , \DM_wd[14]_pad  , \DM_wd[15]_pad  , \DM_wd[1]_pad  , \DM_wd[2]_pad  , \DM_wd[3]_pad  , \DM_wd[4]_pad  , \DM_wd[5]_pad  , \DM_wd[6]_pad  , \DM_wd[7]_pad  , \DM_wd[8]_pad  , \DM_wd[9]_pad  , \DMo_cs0_pad  , \DMo_cs1_pad  , \DMo_cs2_pad  , \DMo_cs3_pad  , \DMo_cs4_pad  , \DMo_cs5_pad  , \DMo_cs6_pad  , \DMo_cs7_pad  , \DSPCLK_cm1_pad  , \EA_do[0]_pad  , \EA_do[10]_pad  , \EA_do[12]_pad  , \EA_do[13]_pad  , \EA_do[14]_pad  , \EA_do[1]_pad  , \EA_do[2]_pad  , \EA_do[3]_pad  , \EA_do[4]_pad  , \EA_do[5]_pad  , \EA_do[6]_pad  , \EA_do[7]_pad  , \EA_do[8]_pad  , \EA_do[9]_pad  , EA_oe_pad , \ED_do[0]_pad  , \ED_do[10]_pad  , \ED_do[11]_pad  , \ED_do[12]_pad  , \ED_do[13]_pad  , \ED_do[14]_pad  , \ED_do[15]_pad  , \ED_do[1]_pad  , \ED_do[2]_pad  , \ED_do[3]_pad  , \ED_do[4]_pad  , \ED_do[5]_pad  , \ED_do[6]_pad  , \ED_do[7]_pad  , \ED_do[8]_pad  , \ED_do[9]_pad  , \ED_oe_14_8_pad  , \ED_oe_7_0_pad  , \IAD_do[0]_pad  , \IAD_do[10]_pad  , \IAD_do[11]_pad  , \IAD_do[12]_pad  , \IAD_do[13]_pad  , \IAD_do[14]_pad  , \IAD_do[15]_pad  , \IAD_do[1]_pad  , \IAD_do[2]_pad  , \IAD_do[3]_pad  , \IAD_do[4]_pad  , \IAD_do[5]_pad  , \IAD_do[6]_pad  , \IAD_do[7]_pad  , \IAD_do[8]_pad  , \IAD_do[9]_pad  , IAD_oe_pad , IDoe_pad , IOSn_pad , \PMAinx[0]_pad  , \PMAinx[10]_pad  , \PMAinx[11]_pad  , \PMAinx[1]_pad  , \PMAinx[2]_pad  , \PMAinx[3]_pad  , \PMAinx[4]_pad  , \PMAinx[5]_pad  , \PMAinx[6]_pad  , \PMAinx[7]_pad  , \PMAinx[8]_pad  , \PMAinx[9]_pad  , \PM_wd[0]_pad  , \PM_wd[10]_pad  , \PM_wd[11]_pad  , \PM_wd[12]_pad  , \PM_wd[13]_pad  , \PM_wd[14]_pad  , \PM_wd[15]_pad  , \PM_wd[1]_pad  , \PM_wd[2]_pad  , \PM_wd[3]_pad  , \PM_wd[4]_pad  , \PM_wd[5]_pad  , \PM_wd[6]_pad  , \PM_wd[7]_pad  , \PM_wd[8]_pad  , \PM_wd[9]_pad  , \PMo_cs0_pad  , \PMo_cs1_pad  , \PMo_cs2_pad  , \PMo_cs3_pad  , \PMo_cs4_pad  , \PMo_cs5_pad  , \PMo_cs6_pad  , \PMo_cs7_pad  , \PMo_oe0_pad  , \RFS0_pad  , \RFS1_pad  , \SCLK0_pad  , \SCLK1_pad  , \TD0_pad  , \TD1_pad  , \TFS0_pad  , \TFS1_pad  , \T_ISn_syn_2  , WRn_pad , XTALoffn_pad , \_al_n0  , \bdma_BDMA_boot_reg/NET0131_reg_syn_3  , \bdma_BDMA_boot_reg/n0  , \bdma_BM_cyc_reg/P0000  , \bdma_BWCOUNT_reg[5]/NET0131_reg_syn_3  , \core_c_psq_MGNT_reg/P0001  , \core_c_psq_cntstk_cnts4x14_CNTcell_reg[0][5]/P0001_reg_syn_3  , \core_c_psq_cntstk_cnts4x14_CNTcell_reg[1][5]/P0001_reg_syn_3  , \core_c_psq_cntstk_cnts4x14_CNTcell_reg[2][5]/P0001_reg_syn_3  , \core_c_psq_cntstk_cnts4x14_CNTcell_reg[3][5]/P0001_reg_syn_3  , \core_eu_ea_alu_ea_reg_afrwe_DO_reg[12]/P0001_reg_syn_3  , \core_eu_ea_alu_ea_reg_afrwe_DO_reg[14]/P0001_reg_syn_3  , \core_eu_ea_alu_ea_reg_afrwe_DO_reg[1]/P0001_reg_syn_3  , \core_eu_ea_alu_ea_reg_afrwe_DO_reg[2]/P0001_reg_syn_3  , \core_eu_ea_alu_ea_reg_afrwe_DO_reg[4]/P0001_reg_syn_3  , \core_eu_ea_alu_ea_reg_afrwe_DO_reg[6]/P0001_reg_syn_3  , \core_eu_ea_alu_ea_reg_afrwe_DO_reg[9]/P0001_reg_syn_3  , \core_eu_ea_alu_ea_reg_afswe_DO_reg[12]/P0001_reg_syn_3  , \core_eu_ea_alu_ea_reg_afswe_DO_reg[14]/P0001_reg_syn_3  , \core_eu_ea_alu_ea_reg_afswe_DO_reg[1]/P0001_reg_syn_3  , \core_eu_ea_alu_ea_reg_afswe_DO_reg[2]/P0001_reg_syn_3  , \core_eu_ea_alu_ea_reg_afswe_DO_reg[4]/P0001_reg_syn_3  , \core_eu_ea_alu_ea_reg_afswe_DO_reg[6]/P0001_reg_syn_3  , \core_eu_ea_alu_ea_reg_afswe_DO_reg[9]/P0001_reg_syn_3  , \core_eu_ec_cun_MVi_pre_C_reg/P0001_reg_syn_3  , \core_eu_em_mac_em_reg_Sq_E_reg/P0001_reg_syn_3  , \emc_DMDreg_reg[8]/P0001_reg_syn_3  , \emc_DMDreg_reg[9]/P0001_reg_syn_3  , \emc_ECMcs_reg/P0001  , \emc_PMDreg_reg[8]/P0001_reg_syn_3  , \emc_PMDreg_reg[9]/P0001_reg_syn_3  , \g10/_0_  , \g1000/_0_  , \g10000/_0_  , \g10001/_0_  , \g10002/_0_  , \g10003/_0_  , \g10004/_0_  , \g10005/_0_  , \g10007/_0_  , \g10008/_0_  , \g10009/_0_  , \g1001/_3_  , \g10010/_0_  , \g10011/_0_  , \g10012/_0_  , \g10013/_0_  , \g10014/_0_  , \g10015/_0_  , \g10016/_0_  , \g10017/_0_  , \g10018/_0_  , \g10019/_0_  , \g1002/_3_  , \g10020/_0_  , \g10021/_0_  , \g10022/_0_  , \g10023/_0_  , \g10024/_0_  , \g10025/_0_  , \g10026/_0_  , \g10027/_0_  , \g10028/_0_  , \g10029/_0_  , \g1003/_0_  , \g10030/_0_  , \g10031/_0_  , \g10032/_0_  , \g10033/_0_  , \g10034/_0_  , \g10035/_0_  , \g10036/_0_  , \g10037/_0_  , \g10038/_0_  , \g10039/_0_  , \g10040/_0_  , \g10041/_0_  , \g10042/_0_  , \g10043/_0_  , \g10044/_0_  , \g10045/_0_  , \g10046/_0_  , \g10047/_0_  , \g10048/_0_  , \g10049/_0_  , \g10050/_0_  , \g10051/_0_  , \g10052/_0_  , \g10053/_0_  , \g10054/_0_  , \g10055/_0_  , \g10056/_0_  , \g10057/_0_  , \g10058/_0_  , \g10059/_0_  , \g10060/_0_  , \g10061/_0_  , \g10062/_0_  , \g10063/_0_  , \g10064/_0_  , \g10065/_0_  , \g10066/_0_  , \g10067/_0_  , \g10068/_0_  , \g10069/_0_  , \g10070/_0_  , \g10071/_0_  , \g10072/_0_  , \g10073/_0_  , \g10074/_0_  , \g10075/_0_  , \g10076/_0_  , \g10077/_0_  , \g10078/_0_  , \g10080/_0_  , \g10081/_0_  , \g10083/_0_  , \g10089/_0_  , \g1009/_0_  , \g10090/_0_  , \g10091/_0_  , \g10092/_0_  , \g10093/_0_  , \g10094/_0_  , \g1010/_0_  , \g10108/_3_  , \g1011/_0_  , \g10110/_0_  , \g10111/_0_  , \g10113/_3_  , \g10115/_3_  , \g1013/_0_  , \g1014/_0_  , \g10152/_0_  , \g10153/_0_  , \g10154/_0_  , \g10155/_0_  , \g10156/_0_  , \g10157/_0_  , \g10158/_0_  , \g10159/_0_  , \g1016/_0_  , \g10160/_0_  , \g10161/_0_  , \g10162/_0_  , \g10163/_0_  , \g10164/_0_  , \g10165/_0_  , \g1017/_0_  , \g10170/_3_  , \g1018/_0_  , \g10190/_3_  , \g10194/_3_  , \g10198/_0_  , \g10199/_0_  , \g102/_0_  , \g103/_0_  , \g104/_0_  , \g105/_0_  , \g10598/_0_  , \g106/_0_  , \g10667/_0_  , \g10683/_0_  , \g10685/_0_  , \g107/_0_  , \g10721/_0_  , \g10758/_0_  , \g10765/_0_  , \g10778/_0_  , \g10791/_0_  , \g108/_0_  , \g10887/_0_  , \g1089/_0_  , \g109/_0_  , \g1090/_0_  , \g1091/_0_  , \g1092/_0_  , \g10923/_0_  , \g1093/_0_  , \g10930/_0_  , \g10931/_0_  , \g10936/_0_  , \g1097/_0_  , \g11/_0_  , \g110/_0_  , \g1101/_0_  , \g11013/_0_  , \g1102/_0_  , \g1103/_0_  , \g11032/_0_  , \g1104/_0_  , \g1105/_0_  , \g1107/_0_  , \g11074/_0_  , \g11077/_0_  , \g1108/_0_  , \g1109/_0_  , \g11112/_0_  , \g11115/_0_  , \g11116/_0_  , \g11119/_0_  , \g11120/_0_  , \g1113/_0_  , \g1115/_0_  , \g1116/_0_  , \g1117/_0_  , \g11267/_0_  , \g11281/_0_  , \g11287/_0_  , \g11300/_0_  , \g11323/_0_  , \g11325/_2__syn_2  , \g11345/_2_  , \g11470/_0_  , \g11471/_0_  , \g11472/_0_  , \g11473/_0_  , \g11474/_0_  , \g11476/_0_  , \g11477/_0_  , \g11496/_0_  , \g11497/_0_  , \g11498/_0_  , \g11499/_0_  , \g11500/_0_  , \g11501/_0_  , \g11502/_0_  , \g11503/_0_  , \g11504/_0_  , \g11505/_0_  , \g11506/_0_  , \g11507/_0_  , \g11509/_0_  , \g11510/_0_  , \g11515/_0_  , \g11516/_0_  , \g11520/_0_  , \g11521/_0_  , \g11576/_0_  , \g11577/_0_  , \g11578/_0_  , \g11579/_0_  , \g11580/_0_  , \g11581/_0_  , \g11582/_0_  , \g11583/_0_  , \g11584/_0_  , \g11585/_0_  , \g11586/_0_  , \g11587/_0_  , \g11588/_0_  , \g11589/_0_  , \g11591/_0_  , \g11593/_0_  , \g11595/_0_  , \g11596/_0_  , \g11597/_0_  , \g11605/_0_  , \g11606/_0_  , \g11607/_0_  , \g11608/_0_  , \g11609/_0_  , \g11610/_0_  , \g11611/_0_  , \g11612/_0_  , \g11613/_0_  , \g11615/_0_  , \g11616/_0_  , \g11617/_0_  , \g11651/_3_  , \g11704/_0_  , \g11705/_0_  , \g11709/_0_  , \g11722/_0_  , \g11723/_0_  , \g119/_0_  , \g1192/_0_  , \g11994/_0_  , \g120/_0_  , \g1200/_0_  , \g12003/_0_  , \g1201/_0_  , \g12019/_0_  , \g1203/_3_  , \g1204/_3_  , \g1207/_0_  , \g1208/_0_  , \g12092/_0_  , \g1210/_0_  , \g1211/_0_  , \g1212/_0_  , \g1213/_0_  , \g12145/_0_  , \g12155/_0_  , \g12186/_0_  , \g12187/_0_  , \g12192/_0_  , \g12201/_0_  , \g12202/_0_  , \g12203/_0_  , \g12204/_0_  , \g12207/_0_  , \g12229/_3_  , \g12267/_0_  , \g12276/_0_  , \g12278/_0_  , \g12279/_0_  , \g12280/_0_  , \g12302/_0_  , \g12316/_0_  , \g12317/_0_  , \g12319/_0_  , \g12328/_3_  , \g1233/_0_  , \g12348/_0_  , \g12351/_0_  , \g12352/_0_  , \g12353/_0_  , \g12354/_0_  , \g12355/_0_  , \g1237/_0_  , \g124/_0_  , \g12444/_0_  , \g125/_0_  , \g12637/_0_  , \g12639/_0_  , \g12658/_0_  , \g12659/_0_  , \g12660/_0_  , \g12663/_0_  , \g12664/_0_  , \g12665/_0_  , \g12672/_3_  , \g12673/_3_  , \g12674/_3_  , \g12675/_3_  , \g12676/_3_  , \g12677/_3_  , \g12678/_0_  , \g12679/_3_  , \g12697/_3_  , \g12701/_3_  , \g12711/_2_  , \g12713/_2_  , \g12715/_2_  , \g12717/_2_  , \g12718/_2__syn_2  , \g1272/_0_  , \g12728/_1__syn_2  , \g12730/_3_  , \g12741/_1__syn_2  , \g12746/_0__syn_2  , \g12748/_0_  , \g12749/_0_  , \g12759/_1__syn_2  , \g12760/_0_  , \g12762/_0_  , \g12763/_0_  , \g12764/_0_  , \g12765/_0_  , \g12766/_0_  , \g12767/_0_  , \g12768/_0_  , \g12769/_0_  , \g12770/_0_  , \g12771/_0_  , \g12772/_0_  , \g12773/_0_  , \g12774/_0_  , \g12775/_0_  , \g12776/_0_  , \g12777/_0_  , \g12778/_0_  , \g12779/_0_  , \g1278/_0_  , \g12780/_0_  , \g12781/_0_  , \g12782/_0_  , \g12783/_0_  , \g12784/_0_  , \g12785/_0_  , \g12786/_0_  , \g12787/_0_  , \g12788/_0_  , \g12789/_0_  , \g12790/_0_  , \g12791/_0_  , \g12792/_0_  , \g12793/_0_  , \g12794/_0_  , \g12795/_0_  , \g12796/_0_  , \g12797/_0_  , \g12798/_0_  , \g12799/_0_  , \g12800/_0_  , \g12801/_0_  , \g12802/_0_  , \g12803/_0_  , \g12804/_0_  , \g12805/_0_  , \g12806/_0_  , \g12807/_0_  , \g12808/_0_  , \g12809/_0_  , \g1281/_0_  , \g12810/_0_  , \g12811/_0_  , \g12812/_0_  , \g12813/_0_  , \g12814/_0_  , \g12815/_0_  , \g12816/_0_  , \g12817/_0_  , \g12818/_0_  , \g12819/_0_  , \g1282/_0_  , \g12820/_0_  , \g12821/_0_  , \g12822/_0_  , \g12823/_0_  , \g12824/_0_  , \g12825/_0_  , \g12826/_0_  , \g12827/_0_  , \g12828/_0_  , \g12829/_0_  , \g12830/_0_  , \g12831/_0_  , \g12832/_0_  , \g12833/_0_  , \g12835/_0_  , \g12836/_0_  , \g12838/_0_  , \g12848/_0_  , \g12849/_0_  , \g1285/_0_  , \g12850/_0_  , \g12857/_0_  , \g12858/_0_  , \g12859/_0_  , \g12861/_0_  , \g12862/_0_  , \g12868/_0_  , \g12869/_0_  , \g1287/_0_  , \g12870/_0_  , \g12871/_0_  , \g12872/_0_  , \g12873/_0_  , \g12874/_0_  , \g12875/_0_  , \g12876/_0_  , \g12877/_0_  , \g12878/_0_  , \g12879/_0_  , \g12880/_0_  , \g12881/_0_  , \g12882/_0_  , \g12883/_0_  , \g12884/_0_  , \g12885/_0_  , \g12886/_0_  , \g12887/_0_  , \g12888/_0_  , \g12889/_0_  , \g1289/_0_  , \g12890/_0_  , \g12891/_0_  , \g12894/_0_  , \g12898/_0_  , \g12899/_0_  , \g12900/_0_  , \g12901/_0_  , \g12902/_0_  , \g12903/_0_  , \g12906/_0_  , \g12907/_0_  , \g12908/_0_  , \g12912/_0_  , \g12913/_0_  , \g12914/_0_  , \g12915/_0_  , \g12916/_0_  , \g12917/_0_  , \g12918/_0_  , \g12919/_0_  , \g12920/_0_  , \g12921/_0_  , \g12922/_0_  , \g12923/_0_  , \g12924/_0_  , \g12925/_0_  , \g12926/_0_  , \g12932/_0_  , \g12933/_0_  , \g12936/_0_  , \g12955/_0_  , \g13015/_0_  , \g13016/_0_  , \g13017/_0_  , \g13018/_0_  , \g13019/_0_  , \g13020/_0_  , \g13021/_0_  , \g13024/_0_  , \g13025/_0_  , \g13027/_0_  , \g13028/_0_  , \g13030/_0_  , \g13031/_0_  , \g13033/_0_  , \g13047/_0_  , \g13060/_0_  , \g13062/_0_  , \g13063/_0_  , \g13064/_0_  , \g13067/_0_  , \g13068/_0_  , \g13069/_0_  , \g13070/_0_  , \g13072/_0_  , \g13094/_0_  , \g13104/_0_  , \g13110/_0_  , \g13114/_0_  , \g13115/_0_  , \g13116/_0_  , \g13117/_0_  , \g13118/_0_  , \g13119/_0_  , \g13120/_0_  , \g13121/_0_  , \g13124/_0_  , \g13125/_0_  , \g13127/_0_  , \g13128/_0_  , \g13129/_0_  , \g13130/_0_  , \g13131/_0_  , \g13132/_0_  , \g13133/_0_  , \g13134/_0_  , \g13138/_0_  , \g13139/_0_  , \g13140/_0_  , \g13141/_0_  , \g13142/_0_  , \g13143/_0_  , \g13144/_0_  , \g13146/_0_  , \g13150/_0_  , \g13152/_0_  , \g13154/_0_  , \g13155/_0_  , \g13156/_0_  , \g13157/_0_  , \g13158/_0_  , \g1320/_3_  , \g13266/_0_  , \g13269/_0_  , \g13274/_0_  , \g13277/_0_  , \g13280/_0_  , \g13283/_0_  , \g13294/_0_  , \g13330/_0_  , \g13333/_0_  , \g13334/_0_  , \g13335/_0_  , \g13336/_0_  , \g13337/_0_  , \g13338/_0_  , \g13345/_0_  , \g13346/_0_  , \g13347/_0_  , \g13348/_0_  , \g13349/_0_  , \g13350/_0_  , \g13351/_0_  , \g13352/_0_  , \g13486/_0_  , \g13488/_0_  , \g13508/_0_  , \g13509/_0_  , \g13510/_0_  , \g13511/_0_  , \g13512/_0_  , \g13513/_0_  , \g13514/_0_  , \g13515/_0_  , \g13516/_0_  , \g13517/_0_  , \g13518/_0_  , \g13519/_0_  , \g13520/_0_  , \g13521/_0_  , \g13540/_0_  , \g13541/_0_  , \g13542/_0_  , \g13543/_0_  , \g13544/_0_  , \g13545/_0_  , \g13546/_0_  , \g13547/_0_  , \g13548/_0_  , \g13549/_0_  , \g13550/_0_  , \g13551/_0_  , \g13552/_0_  , \g13553/_0_  , \g13554/_0_  , \g13555/_0_  , \g13556/_0_  , \g13557/_0_  , \g13558/_0_  , \g13559/_0_  , \g13560/_0_  , \g13561/_0_  , \g13562/_0_  , \g13563/_0_  , \g13564/_0_  , \g13565/_0_  , \g13566/_0_  , \g13567/_0_  , \g13568/_0_  , \g13569/_0_  , \g13570/_0_  , \g13571/_0_  , \g13572/_0_  , \g137/_3_  , \g1387/_3_  , \g1388/_3_  , \g1389/_0_  , \g139/_0_  , \g1390/_0_  , \g1393/_0_  , \g140/_0_  , \g141/_0_  , \g14173/_0_  , \g14176/_0_  , \g142/_3_  , \g14273/_1__syn_2  , \g14274/_0_  , \g14280/_0_  , \g14281/_0_  , \g143/_3_  , \g14354/_3__syn_2  , \g14370/_0_  , \g14385/_0_  , \g14386/_0_  , \g144/_3_  , \g14407/_0_  , \g14412/_0_  , \g14435/_0_  , \g14439/_0_  , \g145/_0_  , \g14522/_0_  , \g14528/_0_  , \g14533/_0_  , \g14581/_1_  , \g14582/_0_  , \g146/_3_  , \g14671/_0_  , \g14672/_0_  , \g147/_0_  , \g1473/_0_  , \g148/_0_  , \g14826/_0_  , \g149/_0_  , \g14908/_0_  , \g14911/_0_  , \g14936/_2_  , \g1494/_0_  , \g1495/_0_  , \g14950/_2_  , \g14953/_2_  , \g15003/_0_  , \g15004/_0_  , \g15006/_0_  , \g15007/_0_  , \g15008/_0_  , \g15009/_0_  , \g15010/_0_  , \g15011/_0_  , \g15012/_0_  , \g15013/_0_  , \g15014/_0_  , \g15015/_0_  , \g15016/_0_  , \g15017/_0_  , \g15018/_0_  , \g15019/_0_  , \g15035/_0_  , \g15036/_0_  , \g15038/_0_  , \g15039/_0_  , \g15040/_0_  , \g15041/_0_  , \g15042/_0_  , \g15043/_0_  , \g15044/_0_  , \g15045/_0_  , \g15046/_0_  , \g15056/_00_  , \g151/_0_  , \g15193/_0_  , \g152/_0_  , \g15256/_0_  , \g153/_0_  , \g15393/_0_  , \g15394/_0_  , \g15395/_0_  , \g15396/_0_  , \g15397/_0_  , \g15398/_0_  , \g15399/_0_  , \g154/_0_  , \g15400/_0_  , \g15401/_0_  , \g15402/_0_  , \g15403/_0_  , \g15404/_0_  , \g15405/_0_  , \g15406/_0_  , \g15407/_0_  , \g15408/_0_  , \g15473/_0_  , \g15650/_0_  , \g15651/_0_  , \g15652/_0_  , \g15653/_0_  , \g15662/_0_  , \g15663/_0_  , \g15664/_0_  , \g15665/_0_  , \g15666/_0_  , \g15667/_0_  , \g15668/_0_  , \g15669/_0_  , \g15670/_0_  , \g15671/_0_  , \g15672/_0_  , \g15673/_0_  , \g15674/_0_  , \g15675/_0_  , \g1569/_0_  , \g1570/_0_  , \g1575/_0_  , \g1576/_0_  , \g15922/_1_  , \g15970/_0_  , \g16059/_0_  , \g1606/_3_  , \g16124/_0_  , \g16144/_0_  , \g16202/_0_  , \g16214/_0_  , \g16247/_0_  , \g16257/_0_  , \g16274/_1_  , \g16324/_0_  , \g16343/_1__syn_2  , \g16381/_0_  , \g16383/_0_  , \g16386/_0_  , \g16414/_1__syn_2  , \g16416/_0__syn_2  , \g16448/_0_  , \g16460/_1_  , \g16625/_3_  , \g16662/_0_  , \g16668/_1__syn_2  , \g16692/_0_  , \g16721/_0_  , \g16723/_0_  , \g16725/_0_  , \g16726/_0_  , \g16727/_0_  , \g16728/_0_  , \g16729/_0_  , \g16730/_0_  , \g16731/_0_  , \g16732/_0_  , \g16733/_0_  , \g16734/_0_  , \g16735/_0_  , \g16736/_0_  , \g16737/_0_  , \g16738/_0_  , \g16739/_0_  , \g16740/_0_  , \g16741/_0_  , \g16742/_0_  , \g16743/_0_  , \g16747/_0_  , \g16748/_0_  , \g16749/_0_  , \g16750/_0_  , \g16753/_0_  , \g16754/_0_  , \g16755/_0_  , \g16756/_0_  , \g16757/_0_  , \g16758/_0_  , \g16761/_0_  , \g16765/_0_  , \g16766/_0_  , \g16767/_0_  , \g16768/_0_  , \g16769/_0_  , \g16772/_0_  , \g16785/_0_  , \g16786/_0_  , \g16787/_0_  , \g16788/_0_  , \g16789/_0_  , \g16790/_0_  , \g16791/_0_  , \g16804/_0_  , \g16805/_0_  , \g16806/_0_  , \g16807/_0_  , \g16808/_0_  , \g16809/_0_  , \g16810/_0_  , \g16811/_0_  , \g16812/_0_  , \g16813/_0_  , \g16814/_0_  , \g16815/_0_  , \g16816/_0_  , \g16817/_0_  , \g16819/_0_  , \g16822/_0_  , \g16823/_0_  , \g16824/_0_  , \g16825/_0_  , \g16828/_0_  , \g16829/_0_  , \g16830/_0_  , \g16831/_0_  , \g16832/_0_  , \g16833/_0_  , \g16834/_0_  , \g16835/_0_  , \g16836/_0_  , \g16837/_0_  , \g16840/_0_  , \g16841/_0_  , \g16842/_0_  , \g16843/_0_  , \g16846/_0_  , \g16847/_0_  , \g16848/_0_  , \g16849/_0_  , \g16850/_0_  , \g16851/_0_  , \g16852/_0_  , \g16853/_0_  , \g16854/_0_  , \g16855/_0_  , \g16856/_0_  , \g16857/_0_  , \g16859/_0_  , \g16862/_0_  , \g16865/_0_  , \g16866/_0_  , \g16867/_0_  , \g16868/_0_  , \g16869/_0_  , \g16870/_0_  , \g16871/_0_  , \g16872/_0_  , \g16873/_0_  , \g16874/_0_  , \g16875/_0_  , \g16876/_0_  , \g16877/_0_  , \g16878/_0_  , \g16879/_0_  , \g16880/_0_  , \g16881/_0_  , \g16882/_0_  , \g16884/_0_  , \g16887/_0_  , \g16891/_0_  , \g16892/_0_  , \g16893/_0_  , \g16894/_0_  , \g16895/_0_  , \g16897/_0_  , \g16898/_0_  , \g16899/_0_  , \g16900/_0_  , \g16901/_0_  , \g16902/_0_  , \g16903/_0_  , \g16904/_0_  , \g16905/_0_  , \g16906/_0_  , \g16907/_0_  , \g16908/_0_  , \g16909/_0_  , \g16910/_0_  , \g16912/_0_  , \g16914/_0_  , \g16915/_0_  , \g16950/_0_  , \g16951/_0_  , \g16952/_0_  , \g16953/_0_  , \g16954/_0_  , \g16955/_0_  , \g16956/_0_  , \g16957/_0_  , \g16958/_0_  , \g16959/_0_  , \g16960/_0_  , \g16961/_0_  , \g16962/_0_  , \g16963/_0_  , \g16964/_0_  , \g16965/_0_  , \g16966/_0_  , \g16967/_0_  , \g16968/_0_  , \g16970/_0_  , \g17102/_3_  , \g17106/_0_  , \g17107/_0_  , \g17109/_0_  , \g17110/_0_  , \g17111/_0_  , \g17112/_0_  , \g17115/_0_  , \g17116/_0_  , \g17119/_0_  , \g17120/_0_  , \g17122/_0_  , \g17123/_0_  , \g17124/_0_  , \g17125/_0_  , \g17126/_0_  , \g17127/_0_  , \g17128/_0_  , \g17130/_0_  , \g17131/_0_  , \g17132/_0_  , \g17133/_0_  , \g17134/_0_  , \g17135/_0_  , \g17136/_0_  , \g17137/_0_  , \g17138/_0_  , \g17140/_0_  , \g17141/_0_  , \g17142/_0_  , \g17143/_0_  , \g17144/_0_  , \g17145/_0_  , \g17146/_0_  , \g17147/_0_  , \g17148/_0_  , \g17149/_0_  , \g17150/_0_  , \g17151/_0_  , \g17152/_0_  , \g17153/_0_  , \g17154/_0_  , \g17155/_0_  , \g17157/_0_  , \g17159/_0_  , \g17160/_0_  , \g17161/_0_  , \g17162/_0_  , \g17163/_0_  , \g17164/_0_  , \g17165/_0_  , \g17166/_0_  , \g17168/_0_  , \g17171/_0_  , \g17173/_0_  , \g17177/_0_  , \g17178/_0_  , \g17179/_0_  , \g17180/_0_  , \g17182/_0_  , \g17183/_0_  , \g17184/_0_  , \g17185/_0_  , \g17186/_0_  , \g17188/_0_  , \g17189/_0_  , \g17190/_0_  , \g17191/_0_  , \g17193/_0_  , \g17194/_0_  , \g17195/_0_  , \g17196/_0_  , \g17197/_0_  , \g17198/_0_  , \g17199/_0_  , \g17200/_0_  , \g17201/_0_  , \g17202/_0_  , \g17203/_0_  , \g17204/_0_  , \g17205/_0_  , \g17206/_0_  , \g17207/_0_  , \g17208/_0_  , \g17209/_0_  , \g17210/_0_  , \g17211/_0_  , \g17212/_0_  , \g17213/_0_  , \g17214/_0_  , \g17215/_0_  , \g17216/_0_  , \g17217/_0_  , \g17218/_0_  , \g17219/_0_  , \g17223/_0_  , \g17224/_0_  , \g17225/_0_  , \g17226/_0_  , \g17227/_0_  , \g17228/_0_  , \g17229/_0_  , \g17231/_0_  , \g17232/_0_  , \g17233/_0_  , \g17234/_0_  , \g17237/_0_  , \g17239/_0_  , \g17240/_0_  , \g17243/_0_  , \g17246/_0_  , \g17247/_0_  , \g17248/_0_  , \g17249/_0_  , \g17250/_0_  , \g17251/_0_  , \g17252/_0_  , \g17253/_0_  , \g17254/_0_  , \g17258/_0_  , \g17261/_0_  , \g17262/_0_  , \g17269/_0_  , \g17271/_0_  , \g17274/_0_  , \g17275/_0_  , \g17276/_0_  , \g17277/_0_  , \g17278/_0_  , \g17279/_0_  , \g17280/_0_  , \g17281/_0_  , \g17282/_0_  , \g17283/_0_  , \g17285/_0_  , \g17290/_0_  , \g17292/_0_  , \g17293/_0_  , \g17296/_0_  , \g17297/_0_  , \g17298/_0_  , \g173/_0_  , \g17303/_0_  , \g17304/_0_  , \g17305/_0_  , \g17306/_0_  , \g17307/_0_  , \g17308/_0_  , \g17309/_0_  , \g17310/_0_  , \g17311/_0_  , \g17312/_0_  , \g17314/_0_  , \g17315/_0_  , \g17316/_0_  , \g17317/_0_  , \g17318/_0_  , \g17319/_0_  , \g17320/_0_  , \g17321/_0_  , \g17322/_0_  , \g17323/_0_  , \g17324/_0_  , \g17325/_0_  , \g17326/_0_  , \g17327/_0_  , \g17328/_0_  , \g17329/_0_  , \g17330/_0_  , \g17331/_0_  , \g17332/_0_  , \g17333/_0_  , \g17335/_0_  , \g17336/_0_  , \g17337/_0_  , \g17338/_0_  , \g17339/_0_  , \g17340/_0_  , \g17342/_0_  , \g17343/_0_  , \g17347/_0_  , \g17350/_0_  , \g17354/_0_  , \g17356/_0_  , \g17357/_0_  , \g17358/_0_  , \g17359/_0_  , \g17360/_0_  , \g17415/_0_  , \g17441/_0_  , \g17442/_0_  , \g17451/_0_  , \g17457/_0_  , \g17458/_0_  , \g17459/_0_  , \g17460/_0_  , \g17461/_0_  , \g17462/_0_  , \g17463/_0_  , \g17464/_0_  , \g17465/_0_  , \g17466/_0_  , \g17467/_0_  , \g17468/_0_  , \g17469/_0_  , \g17470/_0_  , \g17471/_0_  , \g17472/_0_  , \g175/_3_  , \g1750/_0_  , \g176/_3_  , \g17619/_0_  , \g17620/_0_  , \g1763/_3_  , \g1764/_3_  , \g1768/_0_  , \g1769/_0_  , \g177/_3_  , \g17737/_0_  , \g17747/_0_  , \g178/_3_  , \g17814/_1_  , \g17815/_0_  , \g17821/_1_  , \g17821/_1__syn_2  , \g17872/_0_  , \g179/_3_  , \g17902/_0_  , \g180/_3_  , \g18020/_1_  , \g18057/_0_  , \g18096/_0_  , \g18099/_0_  , \g18107/_0_  , \g18133/_0_  , \g18140/_1_  , \g18153/_0_  , \g182/_0_  , \g18218/_0_  , \g18244/_0_  , \g18262/_0_  , \g18267/_0_  , \g18387/_1__syn_2  , \g184/_0_  , \g18478/_1_  , \g18585/_3_  , \g18608/_0_  , \g18609/_0_  , \g18613/_0_  , \g18618/_0_  , \g18647/_0_  , \g18687/_2_  , \g18707/_0_  , \g18748/_0_  , \g18753/_0_  , \g18758/_0_  , \g18759/_0_  , \g18760/_0_  , \g18761/_0_  , \g18762/_0_  , \g18763/_0_  , \g18764/_0_  , \g18765/_0_  , \g18766/_0_  , \g18767/_0_  , \g18768/_0_  , \g18770/_0_  , \g18771/_0_  , \g18788/_0_  , \g18796/_0_  , \g18800/_0_  , \g18801/_0_  , \g18802/_0_  , \g18803/_0_  , \g18804/_0_  , \g18805/_0_  , \g18807/_0_  , \g18840/_0_  , \g18843/_0_  , \g18844/_0_  , \g18846/_0_  , \g18847/_0_  , \g18848/_0_  , \g18849/_0_  , \g18850/_0_  , \g18851/_0_  , \g18852/_0_  , \g18853/_0_  , \g18854/_0_  , \g18855/_0_  , \g18856/_0_  , \g18858/_0_  , \g18860/_0_  , \g18861/_0_  , \g18863/_0_  , \g18864/_0_  , \g18866/_0_  , \g18867/_0_  , \g18868/_0_  , \g18869/_0_  , \g18870/_0_  , \g18871/_0_  , \g18872/_0_  , \g18873/_0_  , \g18874/_0_  , \g18875/_0_  , \g18876/_0_  , \g18877/_0_  , \g18878/_0_  , \g18879/_0_  , \g18880/_0_  , \g18881/_0_  , \g18882/_0_  , \g18883/_0_  , \g18888/_0_  , \g18892/_0_  , \g18895/_0_  , \g18896/_0_  , \g18897/_0_  , \g18905/_0_  , \g18908/_0_  , \g18909/_0_  , \g18912/_0_  , \g18918/_0_  , \g18919/_0_  , \g18920/_0_  , \g18921/_0_  , \g18922/_0_  , \g18924/_0_  , \g18925/_0_  , \g18927/_0_  , \g18930/_0_  , \g18966/_0_  , \g18968/_0_  , \g18970/_0_  , \g18974/_0_  , \g18975/_0_  , \g18977/_0_  , \g18981/_0_  , \g18983/_0_  , \g18985/_0_  , \g18987/_0_  , \g18989/_0_  , \g18991/_0_  , \g18992/_0_  , \g18993/_0_  , \g18994/_0_  , \g18995/_0_  , \g18996/_0_  , \g18997/_0_  , \g18998/_0_  , \g18999/_0_  , \g19001/_0_  , \g19003/_0_  , \g19005/_0_  , \g19006/_0_  , \g19014/_0_  , \g19016/_0_  , \g19018/_0_  , \g19020/_0_  , \g19022/_0_  , \g19056/_3_  , \g19058/_3_  , \g19060/_3_  , \g19062/_3_  , \g1910/_0_  , \g19186/_0_  , \g19188/_0_  , \g19235/_0_  , \g19239/_0_  , \g19244/_0_  , \g19253/_0_  , \g19254/_0_  , \g19259/_0_  , \g19261/_0_  , \g19267/_0_  , \g19277/_0_  , \g19278/_0_  , \g19280/_0_  , \g19281/_0_  , \g19282/_0_  , \g19283/_0_  , \g19284/_0_  , \g19285/_0_  , \g19286/_0_  , \g19287/_0_  , \g19288/_0_  , \g19289/_0_  , \g19290/_0_  , \g19291/_0_  , \g19292/_0_  , \g19293/_0_  , \g19294/_0_  , \g19295/_0_  , \g19296/_0_  , \g19297/_0_  , \g19298/_0_  , \g19299/_0_  , \g19300/_0_  , \g19301/_0_  , \g19302/_0_  , \g19303/_0_  , \g19304/_0_  , \g19305/_0_  , \g19306/_0_  , \g19307/_0_  , \g19308/_0_  , \g19315/_0_  , \g19316/_0_  , \g19317/_0_  , \g19318/_0_  , \g19319/_0_  , \g19320/_0_  , \g19321/_0_  , \g19322/_0_  , \g19323/_0_  , \g19325/_3_  , \g19326/_3_  , \g19333/_3_  , \g19341/_3_  , \g19347/_3_  , \g19377/_3_  , \g19381/_3_  , \g19393/_0_  , \g19401/_0_  , \g19402/_0_  , \g195/_2_  , \g19513/_0_  , \g19514/_0_  , \g19515/_0_  , \g19516/_0_  , \g1952/_3_  , \g19529/_0_  , \g19530/_0_  , \g19531/_0_  , \g19532/_0_  , \g19533/_0_  , \g19534/_0_  , \g19535/_0_  , \g19536/_0_  , \g19537/_0_  , \g19539/_0_  , \g19546/_0_  , \g19552/_0_  , \g19553/_0_  , \g19562/_0_  , \g19563/_0_  , \g19564/_0_  , \g19572/_0_  , \g19575/_0_  , \g19615/_0_  , \g19686/_0_  , \g19688/_0_  , \g197/_0_  , \g19729/_0_  , \g19774/_0_  , \g19777/_0_  , \g19791/_0_  , \g19818/_0_  , \g19819/_0_  , \g19828/_0_  , \g19852/_1_  , \g19860/_0_  , \g19861/_0_  , \g19864/_0_  , \g19886/_0_  , \g19887/_0_  , \g199/_0_  , \g19908/_0_  , \g19918/_0_  , \g19927/_0_  , \g19933/_0_  , \g200/_0_  , \g20019/_0_  , \g20046/_0_  , \g20068/_1_  , \g20080/_1_  , \g201/_0_  , \g20137/_0_  , \g20139/_0_  , \g20141/_0_  , \g20152/_1_  , \g20154/_00_  , \g202/_0_  , \g20206/_0_  , \g20211/_2_  , \g20217/_2_  , \g20239/_0_  , \g20265/_2_  , \g20266/_0_  , \g20272/_2_  , \g20278/_2_  , \g20283/_0_  , \g20285/_2_  , \g20288/_2__syn_2  , \g20293/_0_  , \g20295/_2_  , \g203/_0_  , \g20302/_2_  , \g20303/_2_  , \g20304/_2_  , \g20311/_2_  , \g20326/_0_  , \g20330/_0_  , \g2034/_0_  , \g20345/_0_  , \g20346/_0_  , \g2035/_0_  , \g20363/_0_  , \g20364/_0_  , \g204/_0_  , \g2047/_0_  , \g20483/_0_  , \g20493/_00_  , \g205/_0_  , \g20569/_0_  , \g20570/_0_  , \g20571/_0_  , \g206/_0_  , \g20613/_0_  , \g20615/_0_  , \g20657/_1__syn_2  , \g20660/_0_  , \g20685/_0_  , \g207/_0_  , \g20713/_1_  , \g20747/_1_  , \g20784/_0_  , \g20820/_1_  , \g20859/_0_  , \g20873/_2_  , \g20886/_0_  , \g20887/_0_  , \g20891/_2__syn_2  , \g20907/_2_  , \g20936/_2__syn_2  , \g20937/_1_  , \g20955/_0_  , \g20959/_2__syn_2  , \g20967/_0_  , \g20971/_2__syn_2  , \g20974/_1__syn_2  , \g21015/_1_  , \g21051/_2_  , \g21079/_1_  , \g21081/_1_  , \g21087/_2__syn_2  , \g21114/_1_  , \g21116/_1_  , \g21120/_2__syn_2  , \g21147/_0_  , \g21179/_1_  , \g21185/_1_  , \g21223/_0_  , \g21242/_0_  , \g21253/_0_  , \g21257/_0_  , \g21323/_1_  , \g21324/_1_  , \g21366/_0_  , \g21385/_2_  , \g21464/_0_  , \g21475/_3_  , \g21481/_0_  , \g21482/_0_  , \g21494/_3_  , \g21500/_3_  , \g21507/_3_  , \g21511/_3_  , \g21537/_1_  , \g21568/_0_  , \g21591/_0_  , \g21604/_0_  , \g21605/_3_  , \g21606/_0_  , \g21607/_0_  , \g21608/_0_  , \g21609/_0_  , \g21610/_0_  , \g21611/_0_  , \g21612/_0_  , \g21613/_0_  , \g21614/_0_  , \g21615/_0_  , \g21616/_0_  , \g21617/_0_  , \g21618/_0_  , \g21621/_0_  , \g21640/_0_  , \g21678/_0_  , \g21679/_0_  , \g21686/_0_  , \g21692/_3_  , \g21696/_0_  , \g21698/_0_  , \g21702/_3_  , \g21707/_0_  , \g21709/_0_  , \g21728/_0_  , \g21729/_0_  , \g21731/_0_  , \g21732/_0_  , \g21733/_0_  , \g21736/_0_  , \g21744/_3_  , \g21753/_0_  , \g21754/_0_  , \g21755/_0_  , \g21756/_0_  , \g21757/_0_  , \g21759/_0_  , \g21761/_0_  , \g21763/_0_  , \g21764/_0_  , \g21766/_0_  , \g2180/_0_  , \g21853/_3_  , \g21861/_3_  , \g21863/_3_  , \g21869/_3_  , \g2187/_0_  , \g21875/_3_  , \g21877/_3_  , \g21879/_3_  , \g2188/_0_  , \g21900/_0_  , \g22080/_0_  , \g22082/_0_  , \g22135/_0_  , \g22145/_1_  , \g22225/_0_  , \g223/_0_  , \g22354/_0_  , \g224/_0_  , \g22412/_0_  , \g22415/_1__syn_2  , \g225/_0_  , \g2257/_0_  , \g226/_3_  , \g22624/_0_  , \g227/_3_  , \g22702/_0_  , \g22919/_1__syn_2  , \g22933/_0_  , \g22954/_0_  , \g22989/_1_  , \g23529/_0_  , \g23539/_0_  , \g2362/_2_  , \g23766/_0_  , \g24/_3_  , \g24018/_0_  , \g2416/_0_  , \g2420/_0_  , \g24213/_0_  , \g24301/_0_  , \g2479/_0_  , \g248/_3_  , \g2480/_0_  , \g2481/_0_  , \g2482/_0_  , \g2483/_0_  , \g2484/_0_  , \g2485/_0_  , \g2486/_0_  , \g2487/_0_  , \g2488/_0_  , \g249/_3_  , \g2490/_0_  , \g2491/_0_  , \g2492/_0_  , \g2493/_0_  , \g2494/_0_  , \g2495/_0_  , \g2496/_0_  , \g2497/_0_  , \g2507/_0_  , \g2508/_0_  , \g2509/_0_  , \g2510/_0_  , \g2511/_0_  , \g2512/_0_  , \g2513/_0_  , \g2514/_0_  , \g2515/_0_  , \g2516/_0_  , \g25237/_0_  , \g2558/_0_  , \g2562/_0_  , \g2563/_0_  , \g2564/_0_  , \g2565/_0_  , \g2566/_0_  , \g2567/_0_  , \g2699/_0_  , \g27/_2_  , \g271/_0_  , \g272/_3_  , \g273/_3_  , \g274/_3_  , \g275/_3_  , \g276/_3_  , \g277/_3_  , \g2787/_3_  , \g2788/_3_  , \g279/_0_  , \g2795/_0_  , \g2796/_0_  , \g280/_0_  , \g2842/_3_  , \g29/_1_  , \g2927/_0_  , \g2978/_0_  , \g2979/_0_  , \g2980/_0_  , \g2981/_0_  , \g2982/_0_  , \g2983/_0_  , \g2984/_0_  , \g2985/_0_  , \g3021/_3_  , \g3022/_3_  , \g3023/_3_  , \g3024/_3_  , \g3025/_3_  , \g3026/_3_  , \g3027/_3_  , \g3028/_3_  , \g3029/_3_  , \g3030/_3_  , \g3031/_3_  , \g3032/_3_  , \g3033/_3_  , \g3034/_3_  , \g3035/_3_  , \g3036/_3_  , \g3037/_3_  , \g3038/_3_  , \g3039/_3_  , \g3040/_3_  , \g3041/_3_  , \g3042/_3_  , \g3049/_0_  , \g3050/_0_  , \g3051/_0_  , \g3052/_0_  , \g3053/_0_  , \g3054/_0_  , \g3058/_0_  , \g3059/_0_  , \g3088/_0_  , \g3089/_0_  , \g3090/_0_  , \g3091/_0_  , \g3092/_0_  , \g3093/_0_  , \g3094/_0_  , \g3095/_0_  , \g314/_0_  , \g3147/_3_  , \g3148/_3_  , \g3189/_0_  , \g3190/_0_  , \g3191/_0_  , \g3192/_0_  , \g3193/_0_  , \g3194/_0_  , \g3195/_0_  , \g3196/_0_  , \g3197/_0_  , \g3198/_0_  , \g3199/_0_  , \g32/_0_  , \g320/_3_  , \g3200/_0_  , \g3201/_0_  , \g3202/_0_  , \g3203/_0_  , \g3204/_0_  , \g321/_3_  , \g325/_3_  , \g3271/_2_  , \g33/_0_  , \g3363/_0_  , \g3413/_0_  , \g3414/_0_  , \g352/_0_  , \g355/_0_  , \g356/_3_  , \g357/_3_  , \g35_dup/_1_  , \g36/_3_  , \g365/_3_  , \g366/_3_  , \g367/_3_  , \g368/_3_  , \g3687/_0_  , \g369/_3_  , \g37/_3_  , \g370/_3_  , \g372/_3_  , \g374/_3_  , \g3740/_0_  , \g375/_3_  , \g376/_3_  , \g3878/_0_  , \g3879/_0_  , \g388/_3_  , \g3880/_0_  , \g3881/_0_  , \g3882/_0_  , \g389/_3_  , \g3894/_0_  , \g3895/_0_  , \g3896/_0_  , \g3897/_0_  , \g3898/_0_  , \g392/_3_  , \g393/_3_  , \g394/_3_  , \g395/_3_  , \g396/_3_  , \g397/_3_  , \g398/_3_  , \g399/_3_  , \g401/_3_  , \g402/_3_  , \g404/_3_  , \g4048/_0_  , \g405/_3_  , \g4050/_0_  , \g406/_3_  , \g407/_3_  , \g410/_3_  , \g411/_3_  , \g412/_3_  , \g413/_3_  , \g415/_3_  , \g416/_3_  , \g42/_0_  , \g4216/_3_  , \g4217/_3_  , \g4218/_3_  , \g4219/_3_  , \g4296/_0_  , \g4297/_0_  , \g4298/_0_  , \g4299/_0_  , \g43/_0_  , \g4300/_0_  , \g4301/_0_  , \g4302/_0_  , \g4303/_0_  , \g4304/_0_  , \g4305/_0_  , \g4306/_0_  , \g4307/_0_  , \g4308/_0_  , \g4309/_0_  , \g4310/_0_  , \g4311/_0_  , \g4312/_0_  , \g4313/_0_  , \g4314/_0_  , \g4315/_0_  , \g4316/_0_  , \g4317/_0_  , \g4318/_0_  , \g4319/_0_  , \g4320/_0_  , \g4321/_0_  , \g4322/_0_  , \g4323/_0_  , \g436/_0_  , \g44/_0_  , \g448/_3_  , \g45/_0_  , \g4587/_0_  , \g4588/_0_  , \g46/_0_  , \g4601/_0_  , \g4602/_0_  , \g4613/_3_  , \g4614/_3_  , \g4615/_3_  , \g463/_0_  , \g465/_0_  , \g4653/_0_  , \g4654/_0_  , \g4655/_0_  , \g4656/_0_  , \g4659/_0_  , \g466/_0_  , \g468/_3_  , \g469/_3_  , \g4697/_0_  , \g47/_3_  , \g470/_0_  , \g471/_0_  , \g4755/_0_  , \g476/_0_  , \g48/_3_  , \g480/_00_  , \g4839/_0_  , \g4840/_0_  , \g485/_3_  , \g4854/_0_  , \g4855/_0_  , \g4859/_0_  , \g486/_3_  , \g4860/_0_  , \g4880/_0_  , \g4881/_0_  , \g4882/_0_  , \g4883/_0_  , \g4884/_0_  , \g4885/_0_  , \g4886/_0_  , \g4887/_0_  , \g4888/_0_  , \g49/_0_  , \g494/_0_  , \g499/_1_  , \g50/_0_  , \g5002/_0_  , \g5003/_0_  , \g5009/_0_  , \g5010/_0_  , \g5011/_0_  , \g5014/_0_  , \g51/_0_  , \g5105/_0_  , \g5129/_2_  , \g5132/_0_  , \g5135/_0_  , \g5168/_0_  , \g5169/_0_  , \g5173/_0_  , \g5224/_0_  , \g5225/_0_  , \g5226/_0_  , \g5227/_0_  , \g5334/_0_  , \g5335/_0_  , \g5336/_0_  , \g5337/_0_  , \g5338/_0_  , \g5339/_0_  , \g5340/_0_  , \g5341/_0_  , \g5342/_0_  , \g5343/_0_  , \g5344/_0_  , \g5345/_0_  , \g5346/_0_  , \g5347/_0_  , \g5348/_0_  , \g5349/_0_  , \g5395/_0_  , \g54/_0_  , \g5434/_0_  , \g5447/_0_  , \g5450/_0_  , \g5451/_0_  , \g5452/_0_  , \g5453/_0_  , \g5454/_0_  , \g5461/_0_  , \g5483/_0_  , \g5484/_0_  , \g5492/_0_  , \g5493/_0_  , \g5496/_3_  , \g5497/_3_  , \g55/_0_  , \g5500/_0_  , \g5502/_0_  , \g5503/_0_  , \g5506/_0_  , \g5511/_0_  , \g5518/_0_  , \g5519/_0_  , \g5520/_0_  , \g5522/_0_  , \g5523/_0_  , \g5524/_0_  , \g5525/_0_  , \g5532/_0_  , \g5533/_0_  , \g5534/_0_  , \g5535/_0_  , \g5536/_0_  , \g5537/_0_  , \g5538/_0_  , \g5546/_0_  , \g5555/_00_  , \g5593/_0_  , \g5614/_2_  , \g567/_0_  , \g5677/_0_  , \g5678/_0_  , \g5682/_0_  , \g5683/_0_  , \g5684/_0_  , \g5686/_0_  , \g5687/_0_  , \g5689/_0_  , \g5690/_0_  , \g5691/_0_  , \g5692/_0_  , \g5698/_0_  , \g5699/_0_  , \g5700/_0_  , \g5701/_0_  , \g5702/_0_  , \g5703/_0_  , \g5704/_0_  , \g5709/_0_  , \g5711/_0_  , \g5714/_0_  , \g572/_0_  , \g5723/_0_  , \g5724/_0_  , \g5725/_0_  , \g573/_0_  , \g5739/_0_  , \g5740/_0_  , \g575/_0_  , \g5756/_0_  , \g5757/_0_  , \g5758/_0_  , \g5759/_0_  , \g576/_0_  , \g5760/_0_  , \g5761/_0_  , \g5762/_0_  , \g5763/_0_  , \g577/_0_  , \g5772/_0_  , \g5773/_0_  , \g5774/_0_  , \g5775/_0_  , \g5776/_0_  , \g5777/_0_  , \g578/_0_  , \g5781/_0_  , \g5783/_0_  , \g5784/_0_  , \g5785/_0_  , \g5786/_0_  , \g5787/_0_  , \g5788/_0_  , \g5789/_0_  , \g579/_0_  , \g5790/_0_  , \g5791/_0_  , \g5792/_0_  , \g5794/_0_  , \g5795/_0_  , \g5796/_0_  , \g580/_0_  , \g5801/_0_  , \g5802/_0_  , \g5803/_0_  , \g5804/_0_  , \g5805/_0_  , \g581/_0_  , \g5814/_0_  , \g582/_0_  , \g583/_0_  , \g5849/_3_  , \g585/_0_  , \g586/_0_  , \g587/_0_  , \g588/_0_  , \g589/_0_  , \g590/_0_  , \g591/_0_  , \g592/_0_  , \g593/_0_  , \g594/_0_  , \g595/_0_  , \g596/_0_  , \g597/_0_  , \g5971/_0_  , \g5972/_0_  , \g5976/_0_  , \g598/_0_  , \g5989/_0_  , \g599/_0_  , \g600/_0_  , \g601/_0_  , \g602/_0_  , \g603/_0_  , \g604/_0_  , \g605/_0_  , \g6092/_0_  , \g6093/_2_  , \g6094/_0_  , \g6114/_0_  , \g614/_3_  , \g6148/_0_  , \g6149/_0_  , \g6171/_0_  , \g6172/_0_  , \g6173/_0_  , \g6174/_0_  , \g6175/_0_  , \g6176/_0_  , \g6177/_0_  , \g6178/_0_  , \g6179/_0_  , \g6180/_0_  , \g6181/_0_  , \g6182/_0_  , \g6183/_0_  , \g6184/_0_  , \g6185/_0_  , \g6186/_0_  , \g6187/_0_  , \g6193/_0_  , \g6196/_0_  , \g6197/_0_  , \g6198/_3_  , \g6200/_2_  , \g6202/_2_  , \g6203/_3_  , \g6204/_3_  , \g6209/_0_  , \g6211/_0_  , \g6215/_0_  , \g6217/_0_  , \g6219/_0_  , \g6220/_0_  , \g6222/_0_  , \g6224/_0_  , \g6228/_0_  , \g6238/_0_  , \g6239/_0_  , \g6240/_0_  , \g6242/_0_  , \g6243/_0_  , \g6244/_0_  , \g6245/_0_  , \g6246/_0_  , \g6248/_0_  , \g6249/_0_  , \g6259/_0_  , \g6260/_0_  , \g6261/_0_  , \g6262/_0_  , \g6263/_0_  , \g6264/_0_  , \g6265/_0_  , \g6266/_0_  , \g6267/_0_  , \g6268/_0_  , \g6269/_0_  , \g6270/_0_  , \g6271/_0_  , \g6272/_0_  , \g6277/_0_  , \g6318/_0_  , \g6326/_0_  , \g6329/_0_  , \g6330/_0_  , \g6331/_0_  , \g6332/_0_  , \g6333/_0_  , \g6334/_0_  , \g6335/_0_  , \g6336/_0_  , \g6337/_0_  , \g6338/_0_  , \g6339/_0_  , \g6340/_0_  , \g6341/_0_  , \g6342/_0_  , \g6343/_0_  , \g6344/_0_  , \g6345/_0_  , \g6346/_0_  , \g6347/_0_  , \g6348/_0_  , \g6349/_0_  , \g6350/_0_  , \g6351/_0_  , \g6352/_0_  , \g6353/_0_  , \g6354/_0_  , \g6355/_0_  , \g6361/_0_  , \g637/_0_  , \g638/_0_  , \g639/_3_  , \g64/_3_  , \g640/_3_  , \g6419/_0_  , \g6442/_0_  , \g6442/_1_  , \g6489/_0_  , \g6490/_0_  , \g65/_3_  , \g6513/_0_  , \g6515/_0_  , \g6571/_0_  , \g6588/_0_  , \g6589/_0_  , \g6638/_0_  , \g6639/_0_  , \g6653/_0_  , \g6654/_3_  , \g6655/_0_  , \g6656/_0_  , \g6657/_0_  , \g6687/_0_  , \g6688/_0_  , \g6689/_0_  , \g6690/_0_  , \g6691/_0_  , \g6692/_0_  , \g6693/_0_  , \g6694/_0_  , \g6701/_0_  , \g6706/_0_  , \g6711/_0_  , \g6727/_0_  , \g6728/_0_  , \g6736/_0_  , \g6739/_0_  , \g6742/_0_  , \g6746/_0_  , \g6752/_0_  , \g6771/_0_  , \g684/_0_  , \g685/_0_  , \g686/_0_  , \g687/_0_  , \g688/_0_  , \g689/_0_  , \g690/_0_  , \g691/_0_  , \g692/_0_  , \g693/_0_  , \g696/_3_  , \g697/_3_  , \g699/_0_  , \g7/_0_  , \g700/_0_  , \g7005/_0_  , \g7056/_0_  , \g7057/_0_  , \g7058/_0_  , \g7060/_0_  , \g7075/_0_  , \g7086/_0_  , \g7087/_0_  , \g7089/_0_  , \g7108/_0_  , \g7109/_0_  , \g7112/_0_  , \g7172/_2_  , \g7210/_2_  , \g7211/_0_  , \g7212/_0_  , \g7213/_0_  , \g7214/_0_  , \g7215/_0_  , \g7216/_0_  , \g7217/_3_  , \g7218/_0_  , \g7219/_0_  , \g7220/_0_  , \g7222/_0_  , \g7227/_2_  , \g723/_3_  , \g7234/_0_  , \g7237/_3_  , \g7238/_3_  , \g7239/_3_  , \g724/_3_  , \g7240/_3_  , \g7241/_3_  , \g7242/_3_  , \g7243/_3_  , \g7244/_0_  , \g7245/_0_  , \g7246/_0_  , \g7247/_0_  , \g7248/_0_  , \g7249/_0_  , \g7250/_0_  , \g7251/_0_  , \g7253/_0_  , \g7254/_0_  , \g7255/_0_  , \g7256/_0_  , \g7257/_0_  , \g7258/_0_  , \g7261/_0_  , \g7264/_0_  , \g7265/_0_  , \g7266/_0_  , \g7267/_0_  , \g7268/_0_  , \g7269/_0_  , \g7278/_0_  , \g7279/_0_  , \g7280/_0_  , \g7281/_0_  , \g7282/_0_  , \g7283/_0_  , \g7284/_0_  , \g7285/_0_  , \g7286/_3_  , \g7288/_3_  , \g7291/_0_  , \g7296/_3_  , \g73/_0_  , \g7302/_3_  , \g7306/_3_  , \g7310/_3_  , \g7311/_3_  , \g7312/_3_  , \g7313/_3_  , \g7314/_3_  , \g7315/_3_  , \g7316/_3_  , \g7317/_3_  , \g7323/_3_  , \g7324/_3_  , \g7325/_3_  , \g7327/_0_  , \g7362/_0_  , \g74/_0_  , \g75/_0_  , \g7512/_0_  , \g7513/_0_  , \g7514/_0_  , \g7515/_0_  , \g7516/_0_  , \g7518/_0_  , \g7528/_0_  , \g7529/_0_  , \g7548/_0_  , \g7549/_0_  , \g7550/_0_  , \g7575/_0_  , \g7576/_0_  , \g7577/_0_  , \g7578/_0_  , \g7579/_0_  , \g7580/_0_  , \g7581/_0_  , \g7582/_0_  , \g7583/_0_  , \g7584/_0_  , \g7585/_0_  , \g7586/_0_  , \g7587/_0_  , \g7588/_0_  , \g7589/_0_  , \g7590/_0_  , \g7591/_0_  , \g7592/_0_  , \g7593/_0_  , \g7594/_0_  , \g7595/_0_  , \g7596/_0_  , \g7597/_0_  , \g7598/_0_  , \g7599/_0_  , \g76/_0_  , \g7600/_0_  , \g7601/_0_  , \g7602/_0_  , \g7603/_0_  , \g7604/_0_  , \g7614/_0_  , \g7618/_0_  , \g762/_0_  , \g7634/_0_  , \g766/_0_  , \g767/_0_  , \g768/_0_  , \g769/_0_  , \g77/_0_  , \g770/_3_  , \g771/_3_  , \g7715/_0_  , \g774/_0_  , \g7746/_0_  , \g7753/_0_  , \g7754/_0_  , \g7755/_0_  , \g7756/_0_  , \g7757/_0_  , \g7758/_0_  , \g7759/_0_  , \g7760/_0_  , \g7761/_0_  , \g7762/_0_  , \g7763/_0_  , \g7764/_0_  , \g7765/_0_  , \g7766/_0_  , \g7778/_0_  , \g7779/_0_  , \g7780/_0_  , \g7781/_0_  , \g7782/_0_  , \g7784/_0_  , \g78/_0_  , \g7800/_0_  , \g7823/_3_  , \g7837/_0_  , \g7841/_0_  , \g7842/_0_  , \g7843/_0_  , \g7844/_0_  , \g7845/_0_  , \g7846/_0_  , \g7847/_0_  , \g7849/_0_  , \g7850/_0_  , \g7852/_0_  , \g7854/_0_  , \g7855/_0_  , \g7857/_0_  , \g7858/_0_  , \g7859/_0_  , \g7860/_0_  , \g7861/_0_  , \g7862/_0_  , \g7863/_0_  , \g7864/_0_  , \g7865/_0_  , \g7866/_0_  , \g7867/_0_  , \g7868/_0_  , \g7869/_0_  , \g7870/_0_  , \g7871/_0_  , \g79211/_3_  , \g79258/_3_  , \g79299/_3_  , \g79316/_2_  , \g79342/_3_  , \g79401/_3_  , \g79452/_3_  , \g79457/_3_  , \g7951/_0_  , \g79541/_3_  , \g7958/_0_  , \g79598/_3_  , \g79654/_3_  , \g79675/_3_  , \g7971/_0_  , \g7972/_0_  , \g7973/_3_  , \g79753/_3_  , \g7976/_3_  , \g79855/_3_  , \g79858/_3_  , \g79997/_3_  , \g8/_0_  , \g80008/_3_  , \g80011/_0_  , \g80104/_0_  , \g80172/_1_  , \g80195/_3_  , \g80238/_3_  , \g80290/_2_  , \g80294/_0_  , \g80302/_0_  , \g80327/_0_  , \g80360/_3_  , \g80373/_0_  , \g80401/_0_  , \g80410/_0_  , \g80475/_0_  , \g80476/_0_  , \g80516/_3_  , \g80536/_0_  , \g80537/_0_  , \g80572/_0_  , \g80573/_0_  , \g80609/_2_  , \g80610/_2_  , \g80676/_0_  , \g80798/_0_  , \g80807/_0_  , \g80890/_2_  , \g80904/_0_  , \g81719/_2_  , \g81746/_0_  , \g81775/_0_  , \g81872/_0_  , \g81961/_0_  , \g81968/_0_  , \g82096/_0_  , \g82123/_0_  , \g82147/_0_  , \g82147/_1_  , \g82335/_0_  , \g82338/_2_  , \g82368/_0_  , \g82460/_2_  , \g82469/_0_  , \g82481/_0_  , \g82625/_1_  , \g82711/_0_  , \g82772/_0_  , \g82946/_0_  , \g82947/_0_  , \g82956/_0_  , \g83003/_0_  , \g83006/_1_  , \g83415/_0_  , \g83498/_0_  , \g837/_0_  , \g838/_0_  , \g83863/_0_  , \g839/_0_  , \g84049/_3_  , \g84050/_3_  , \g84077/_2_  , \g842/_0_  , \g84245/_0_  , \g843/_0_  , \g844/_0_  , \g84448/_0_  , \g84478/_3_  , \g845/_0_  , \g846/_0_  , \g847/_0_  , \g848/_0_  , \g8487/_0_  , \g8488/_0_  , \g8489/_0_  , \g849/_0_  , \g8490/_0_  , \g84904/_0_  , \g8491/_0_  , \g8492/_0_  , \g8493/_0_  , \g8494/_0_  , \g8496/_0_  , \g8517/_0_  , \g8534/_0_  , \g8538/_0_  , \g8540/_0_  , \g8576/_2_  , \g8597/_0_  , \g8598/_0_  , \g8599/_0_  , \g8600/_0_  , \g8601/_0_  , \g8602/_0_  , \g8603/_0_  , \g8605/_0_  , \g8606/_0_  , \g8607/_0_  , \g8608/_0_  , \g8609/_0_  , \g8610/_0_  , \g8611/_0_  , \g8612/_0_  , \g8613/_0_  , \g8614/_0_  , \g8615/_0_  , \g8617/_0_  , \g8643/_0_  , \g8644/_0_  , \g8645/_0_  , \g8646/_0_  , \g8647/_0_  , \g8648/_0_  , \g8650/_0_  , \g8651/_0_  , \g8652/_0_  , \g8653/_0_  , \g8654/_0_  , \g8655/_0_  , \g8656/_0_  , \g8657/_0_  , \g8658/_0_  , \g8659/_0_  , \g8660/_0_  , \g8665/_00_  , \g8666/_00_  , \g8667/_00_  , \g8668/_00_  , \g8669/_00_  , \g86715/_0_  , \g86745/_3_  , \g8691/_0_  , \g8700/_0_  , \g8701/_0_  , \g8702/_0_  , \g8703/_0_  , \g8704/_0_  , \g8705/_0_  , \g87063/_0_  , \g87114/_0_  , \g8712/_0_  , \g8713/_0_  , \g8714/_0_  , \g87171/_1_  , \g87252/_1_  , \g87298/_0_  , \g8730/_0_  , \g8741/_0_  , \g8747/_0_  , \g87480/_0_  , \g87484/_2_  , \g87488/_1__syn_2  , \g8761/_0_  , \g8762/_0_  , \g8763/_0_  , \g8764/_0_  , \g8765/_0_  , \g8775/_0_  , \g8776/_0_  , \g8777/_0_  , \g8778/_0_  , \g8784/_0_  , \g8804/_0_  , \g8807/_0_  , \g8808/_0_  , \g8809/_0_  , \g8810/_0_  , \g8811/_0_  , \g8812/_0_  , \g8813/_0_  , \g8814/_0_  , \g8815/_0_  , \g8816/_0_  , \g8817/_0_  , \g8818/_0_  , \g8819/_0_  , \g8820/_0_  , \g8821/_0_  , \g8822/_0_  , \g8823/_0_  , \g8824/_0_  , \g8825/_0_  , \g8826/_0_  , \g8827/_0_  , \g8828/_0_  , \g8829/_0_  , \g8830/_0_  , \g8831/_0_  , \g8832/_0_  , \g8833/_0_  , \g8834/_0_  , \g8835/_0_  , \g8836/_0_  , \g8837/_0_  , \g8838/_0_  , \g8839/_0_  , \g8840/_0_  , \g8842/_0_  , \g8843/_0_  , \g8846/_0_  , \g8848/_0_  , \g8857/_0_  , \g8895/_0_  , \g8902/_3_  , \g8903/_3_  , \g8904/_3_  , \g8905/_3_  , \g8906/_3_  , \g8909/_0_  , \g8910/_0_  , \g8911/_0_  , \g8924/_3_  , \g8926/_3_  , \g8927/_3_  , \g8943/_0_  , \g8944/_0_  , \g8958/_3_  , \g8960/_00_  , \g8961/_3_  , \g8965/_0_  , \g8966/_0_  , \g8967/_0_  , \g8968/_0_  , \g9/_0_  , \g9123/_0_  , \g9125/_0_  , \g9126/_0_  , \g913/_0_  , \g915/_0_  , \g916/_0_  , \g917/_0_  , \g918/_0_  , \g919/_0_  , \g920/_3_  , \g921/_3_  , \g925/_0_  , \g926/_0_  , \g927/_0_  , \g928/_0_  , \g929/_0_  , \g930/_0_  , \g9336/_0_  , \g9337/_0_  , \g939/_3_  , \g9396/_0_  , \g9397/_0_  , \g9399/_0_  , \g9400/_0_  , \g9401/_0_  , \g9402/_0_  , \g9403/_0_  , \g9404/_0_  , \g9415/_0_  , \g9418/_0_  , \g9419/_0_  , \g9420/_0_  , \g9446/_0_  , \g9465/_0_  , \g9493/_0_  , \g9536/_0_  , \g9537/_0_  , \g9538/_0_  , \g9539/_0_  , \g9540/_0_  , \g9541/_0_  , \g9542/_0_  , \g955/_2_  , \g9561/_0_  , \g9562/_0_  , \g9563/_0_  , \g9564/_0_  , \g9565/_0_  , \g9566/_0_  , \g9567/_0_  , \g9568/_0_  , \g9569/_0_  , \g9570/_0_  , \g9571/_0_  , \g9572/_0_  , \g9573/_0_  , \g9574/_0_  , \g9575/_0_  , \g9576/_0_  , \g9577/_0_  , \g9578/_0_  , \g9579/_0_  , \g9580/_0_  , \g9581/_0_  , \g9582/_0_  , \g9583/_0_  , \g9584/_0_  , \g9585/_0_  , \g9586/_0_  , \g9587/_0_  , \g9588/_0_  , \g9589/_0_  , \g9590/_0_  , \g9591/_0_  , \g9592/_0_  , \g9593/_0_  , \g9594/_0_  , \g9595/_0_  , \g9596/_0_  , \g9597/_0_  , \g9598/_0_  , \g9599/_0_  , \g9600/_0_  , \g9601/_0_  , \g9602/_0_  , \g9603/_0_  , \g9604/_0_  , \g9605/_0_  , \g9606/_0_  , \g9607/_0_  , \g9608/_0_  , \g9609/_0_  , \g9610/_0_  , \g9611/_0_  , \g9612/_0_  , \g9613/_0_  , \g9614/_0_  , \g9615/_0_  , \g9616/_0_  , \g9617/_0_  , \g9618/_0_  , \g9619/_0_  , \g9620/_0_  , \g9621/_0_  , \g9622/_0_  , \g9623/_0_  , \g9624/_0_  , \g9625/_0_  , \g9626/_0_  , \g9627/_0_  , \g9628/_0_  , \g9629/_0_  , \g9630/_0_  , \g9631/_0_  , \g9632/_0_  , \g9633/_0_  , \g9634/_0_  , \g9635/_0_  , \g9636/_0_  , \g9637/_0_  , \g9638/_0_  , \g9639/_0_  , \g9640/_0_  , \g9641/_0_  , \g9642/_0_  , \g9643/_0_  , \g9644/_0_  , \g9645/_0_  , \g9646/_0_  , \g9647/_0_  , \g9648/_0_  , \g9649/_0_  , \g9650/_0_  , \g9651/_0_  , \g9652/_0_  , \g9653/_0_  , \g9654/_0_  , \g9655/_0_  , \g9656/_0_  , \g9657/_0_  , \g9658/_0_  , \g9659/_0_  , \g9660/_0_  , \g9661/_0_  , \g9662/_0_  , \g9663/_0_  , \g9664/_0_  , \g9665/_0_  , \g9666/_0_  , \g9667/_0_  , \g9668/_0_  , \g9669/_0_  , \g9670/_0_  , \g9671/_0_  , \g9672/_0_  , \g9673/_0_  , \g9674/_0_  , \g9675/_0_  , \g9676/_0_  , \g9677/_0_  , \g9678/_0_  , \g9681/_0_  , \g9683/_0_  , \g9689/_0_  , \g9692/_0_  , \g9694/_0_  , \g9695/_0_  , \g9701/_0_  , \g9702/_0_  , \g9703/_0_  , \g9704/_0_  , \g9709/_0_  , \g9710/_0_  , \g9711/_0_  , \g9712/_0_  , \g9720/_0_  , \g9721/_0_  , \g9722/_0_  , \g9726/_0_  , \g9733/_0_  , \g9734/_0_  , \g9735/_0_  , \g9736/_0_  , \g9737/_0_  , \g9738/_0_  , \g9739/_0_  , \g9740/_0_  , \g9741/_0_  , \g9742/_0_  , \g9743/_0_  , \g9744/_0_  , \g9745/_0_  , \g9746/_0_  , \g9747/_0_  , \g9748/_0_  , \g9749/_0_  , \g9750/_0_  , \g9751/_0_  , \g9752/_0_  , \g9753/_0_  , \g9754/_0_  , \g9755/_0_  , \g9756/_0_  , \g9757/_0_  , \g9758/_0_  , \g9759/_0_  , \g9760/_0_  , \g9761/_0_  , \g9762/_0_  , \g9763/_0_  , \g9764/_0_  , \g9765/_0_  , \g9766/_0_  , \g9767/_0_  , \g9768/_0_  , \g9769/_0_  , \g9770/_0_  , \g9771/_0_  , \g9772/_0_  , \g9773/_0_  , \g9774/_0_  , \g9775/_0_  , \g9776/_0_  , \g9777/_0_  , \g9778/_0_  , \g9779/_0_  , \g9780/_0_  , \g9781/_0_  , \g9782/_0_  , \g9783/_0_  , \g9784/_0_  , \g9785/_0_  , \g9786/_0_  , \g9787/_0_  , \g9788/_0_  , \g9789/_0_  , \g9790/_0_  , \g9791/_0_  , \g9792/_0_  , \g9793/_0_  , \g9794/_0_  , \g9795/_0_  , \g9796/_0_  , \g9797/_0_  , \g9798/_0_  , \g9799/_0_  , \g9800/_0_  , \g9801/_0_  , \g9802/_0_  , \g9803/_0_  , \g9804/_0_  , \g9805/_0_  , \g9806/_0_  , \g9807/_0_  , \g9808/_0_  , \g9809/_0_  , \g9810/_0_  , \g9811/_0_  , \g9812/_0_  , \g9813/_0_  , \g9814/_0_  , \g9815/_0_  , \g9816/_0_  , \g9817/_0_  , \g9818/_0_  , \g9819/_0_  , \g9820/_0_  , \g9821/_0_  , \g9822/_0_  , \g9823/_0_  , \g9824/_0_  , \g9825/_0_  , \g9826/_0_  , \g9827/_0_  , \g9828/_0_  , \g9829/_0_  , \g9830/_0_  , \g9831/_0_  , \g9832/_0_  , \g9833/_0_  , \g9835/_0_  , \g9836/_0_  , \g9837/_0_  , \g9838/_0_  , \g9839/_0_  , \g9840/_0_  , \g9841/_0_  , \g9842/_0_  , \g9844/_0_  , \g9845/_0_  , \g9846/_0_  , \g9848/_0_  , \g9849/_0_  , \g9850/_0_  , \g9851/_0_  , \g9853/_0_  , \g9854/_0_  , \g9855/_0_  , \g9856/_0_  , \g9857/_0_  , \g9858/_0_  , \g9859/_0_  , \g9860/_0_  , \g9862/_0_  , \g9863/_0_  , \g9864/_0_  , \g9865/_0_  , \g9867/_0_  , \g9868/_0_  , \g9876/_0_  , \g9877/_0_  , \g9878/_0_  , \g9879/_0_  , \g9880/_0_  , \g9881/_0_  , \g9898/_0_  , \g9900/_0_  , \g9901/_0_  , \g9902/_0_  , \g9903/_0_  , \g9904/_0_  , \g9905/_0_  , \g9906/_0_  , \g9907/_0_  , \g9908/_0_  , \g9909/_0_  , \g9910/_0_  , \g9911/_0_  , \g9912/_0_  , \g9913/_0_  , \g9914/_0_  , \g9915/_0_  , \g9916/_0_  , \g9917/_0_  , \g9918/_0_  , \g9919/_0_  , \g992/_0_  , \g9920/_0_  , \g9921/_0_  , \g9922/_0_  , \g9923/_0_  , \g9924/_0_  , \g9925/_0_  , \g9926/_0_  , \g9927/_0_  , \g9928/_0_  , \g9929/_0_  , \g9930/_0_  , \g9931/_0_  , \g9932/_0_  , \g9933/_0_  , \g9934/_0_  , \g9935/_0_  , \g9936/_0_  , \g9937/_0_  , \g9938/_0_  , \g9939/_0_  , \g9940/_0_  , \g9941/_0_  , \g9942/_0_  , \g9943/_0_  , \g9944/_0_  , \g9945/_0_  , \g9946/_0_  , \g9947/_0_  , \g9948/_0_  , \g9949/_0_  , \g9950/_0_  , \g9951/_0_  , \g9952/_0_  , \g9953/_0_  , \g9954/_0_  , \g9955/_0_  , \g9956/_0_  , \g9957/_0_  , \g9958/_0_  , \g9959/_0_  , \g9960/_0_  , \g9961/_0_  , \g9962/_0_  , \g9963/_0_  , \g9964/_0_  , \g9965/_0_  , \g9966/_0_  , \g9967/_0_  , \g9968/_0_  , \g9969/_0_  , \g9970/_0_  , \g9971/_0_  , \g9972/_0_  , \g9973/_0_  , \g9974/_0_  , \g9975/_0_  , \g9976/_0_  , \g9977/_0_  , \g9978/_0_  , \g9979/_0_  , \g9980/_0_  , \g9981/_0_  , \g9982/_0_  , \g9983/_0_  , \g9984/_0_  , \g9985/_0_  , \g9987/_0_  , \g9988/_0_  , \g9989/_0_  , \g999/_0_  , \g9990/_0_  , \g9991/_0_  , \g9992/_0_  , \g9993/_0_  , \g9994/_0_  , \g9995/_0_  , \g9996/_0_  , \g9997/_0_  , \g9998/_0_  , \g9999/_0_  , \idma_IDMA_boot_reg/NET0131_reg_syn_3  , \memc_EXTC_Eg_reg/NET0131  , \memc_EXTC_Eg_reg/NET0131_reg_syn_3  , \memc_EXTC_Eg_reg/n0  , \pio_PIO_IN_P_reg[0]/P0001_reg_syn_3  , \pio_PIO_IN_P_reg[10]/P0001_reg_syn_3  , \pio_PIO_IN_P_reg[11]/P0001_reg_syn_3  , \pio_PIO_IN_P_reg[1]/P0001_reg_syn_3  , \pio_PIO_IN_P_reg[2]/P0001_reg_syn_3  , \pio_PIO_IN_P_reg[3]/P0001_reg_syn_3  , \pio_PIO_IN_P_reg[4]/P0001_reg_syn_3  , \pio_PIO_IN_P_reg[5]/P0001_reg_syn_3  , \pio_PIO_IN_P_reg[6]/P0001_reg_syn_3  , \pio_PIO_IN_P_reg[7]/P0001_reg_syn_3  , \pio_PIO_IN_P_reg[8]/P0001_reg_syn_3  , \pio_PIO_IN_P_reg[9]/P0001_reg_syn_3  , \pio_PIO_RES_OUT_reg[0]/P0001_reg_syn_3  , \pio_PIO_RES_OUT_reg[10]/P0001_reg_syn_3  , \pio_PIO_RES_OUT_reg[2]/P0001_reg_syn_3  , \pio_PIO_RES_OUT_reg[4]/P0001_reg_syn_3  , \pio_PIO_RES_OUT_reg[6]/P0001_reg_syn_3  , \sice_GO_NXi_reg/NET0131_reg_syn_3  , \sport0_rxctl_RXSHT_reg[0]/P0001_reg_syn_3  , \sport0_rxctl_RXSHT_reg[1]/P0001_reg_syn_3  , \sport1_rxctl_RXSHT_reg[0]/P0001_reg_syn_3  , \sport1_rxctl_RXSHT_reg[1]/P0001_reg_syn_3  );
  input \CM_rd0[0]_pad  ;
  input \CM_rd0[10]_pad  ;
  input \CM_rd0[11]_pad  ;
  input \CM_rd0[12]_pad  ;
  input \CM_rd0[13]_pad  ;
  input \CM_rd0[14]_pad  ;
  input \CM_rd0[15]_pad  ;
  input \CM_rd0[16]_pad  ;
  input \CM_rd0[17]_pad  ;
  input \CM_rd0[18]_pad  ;
  input \CM_rd0[19]_pad  ;
  input \CM_rd0[1]_pad  ;
  input \CM_rd0[20]_pad  ;
  input \CM_rd0[21]_pad  ;
  input \CM_rd0[22]_pad  ;
  input \CM_rd0[23]_pad  ;
  input \CM_rd0[2]_pad  ;
  input \CM_rd0[3]_pad  ;
  input \CM_rd0[4]_pad  ;
  input \CM_rd0[5]_pad  ;
  input \CM_rd0[6]_pad  ;
  input \CM_rd0[7]_pad  ;
  input \CM_rd0[8]_pad  ;
  input \CM_rd0[9]_pad  ;
  input \CM_rd1[0]_pad  ;
  input \CM_rd1[10]_pad  ;
  input \CM_rd1[11]_pad  ;
  input \CM_rd1[12]_pad  ;
  input \CM_rd1[13]_pad  ;
  input \CM_rd1[14]_pad  ;
  input \CM_rd1[15]_pad  ;
  input \CM_rd1[16]_pad  ;
  input \CM_rd1[17]_pad  ;
  input \CM_rd1[18]_pad  ;
  input \CM_rd1[19]_pad  ;
  input \CM_rd1[1]_pad  ;
  input \CM_rd1[20]_pad  ;
  input \CM_rd1[21]_pad  ;
  input \CM_rd1[22]_pad  ;
  input \CM_rd1[23]_pad  ;
  input \CM_rd1[2]_pad  ;
  input \CM_rd1[3]_pad  ;
  input \CM_rd1[4]_pad  ;
  input \CM_rd1[5]_pad  ;
  input \CM_rd1[6]_pad  ;
  input \CM_rd1[7]_pad  ;
  input \CM_rd1[8]_pad  ;
  input \CM_rd1[9]_pad  ;
  input \CM_rd2[0]_pad  ;
  input \CM_rd2[10]_pad  ;
  input \CM_rd2[11]_pad  ;
  input \CM_rd2[12]_pad  ;
  input \CM_rd2[13]_pad  ;
  input \CM_rd2[14]_pad  ;
  input \CM_rd2[15]_pad  ;
  input \CM_rd2[16]_pad  ;
  input \CM_rd2[17]_pad  ;
  input \CM_rd2[18]_pad  ;
  input \CM_rd2[19]_pad  ;
  input \CM_rd2[1]_pad  ;
  input \CM_rd2[20]_pad  ;
  input \CM_rd2[21]_pad  ;
  input \CM_rd2[22]_pad  ;
  input \CM_rd2[23]_pad  ;
  input \CM_rd2[2]_pad  ;
  input \CM_rd2[3]_pad  ;
  input \CM_rd2[4]_pad  ;
  input \CM_rd2[5]_pad  ;
  input \CM_rd2[6]_pad  ;
  input \CM_rd2[7]_pad  ;
  input \CM_rd2[8]_pad  ;
  input \CM_rd2[9]_pad  ;
  input \CM_rd3[0]_pad  ;
  input \CM_rd3[10]_pad  ;
  input \CM_rd3[11]_pad  ;
  input \CM_rd3[12]_pad  ;
  input \CM_rd3[13]_pad  ;
  input \CM_rd3[14]_pad  ;
  input \CM_rd3[15]_pad  ;
  input \CM_rd3[16]_pad  ;
  input \CM_rd3[17]_pad  ;
  input \CM_rd3[18]_pad  ;
  input \CM_rd3[19]_pad  ;
  input \CM_rd3[1]_pad  ;
  input \CM_rd3[20]_pad  ;
  input \CM_rd3[21]_pad  ;
  input \CM_rd3[22]_pad  ;
  input \CM_rd3[23]_pad  ;
  input \CM_rd3[2]_pad  ;
  input \CM_rd3[3]_pad  ;
  input \CM_rd3[4]_pad  ;
  input \CM_rd3[5]_pad  ;
  input \CM_rd3[6]_pad  ;
  input \CM_rd3[7]_pad  ;
  input \CM_rd3[8]_pad  ;
  input \CM_rd3[9]_pad  ;
  input \CM_rd4[0]_pad  ;
  input \CM_rd4[10]_pad  ;
  input \CM_rd4[11]_pad  ;
  input \CM_rd4[12]_pad  ;
  input \CM_rd4[13]_pad  ;
  input \CM_rd4[14]_pad  ;
  input \CM_rd4[15]_pad  ;
  input \CM_rd4[16]_pad  ;
  input \CM_rd4[17]_pad  ;
  input \CM_rd4[18]_pad  ;
  input \CM_rd4[19]_pad  ;
  input \CM_rd4[1]_pad  ;
  input \CM_rd4[20]_pad  ;
  input \CM_rd4[21]_pad  ;
  input \CM_rd4[22]_pad  ;
  input \CM_rd4[23]_pad  ;
  input \CM_rd4[2]_pad  ;
  input \CM_rd4[3]_pad  ;
  input \CM_rd4[4]_pad  ;
  input \CM_rd4[5]_pad  ;
  input \CM_rd4[6]_pad  ;
  input \CM_rd4[7]_pad  ;
  input \CM_rd4[8]_pad  ;
  input \CM_rd4[9]_pad  ;
  input \CM_rd5[0]_pad  ;
  input \CM_rd5[10]_pad  ;
  input \CM_rd5[11]_pad  ;
  input \CM_rd5[12]_pad  ;
  input \CM_rd5[13]_pad  ;
  input \CM_rd5[14]_pad  ;
  input \CM_rd5[15]_pad  ;
  input \CM_rd5[16]_pad  ;
  input \CM_rd5[17]_pad  ;
  input \CM_rd5[18]_pad  ;
  input \CM_rd5[19]_pad  ;
  input \CM_rd5[1]_pad  ;
  input \CM_rd5[20]_pad  ;
  input \CM_rd5[21]_pad  ;
  input \CM_rd5[22]_pad  ;
  input \CM_rd5[23]_pad  ;
  input \CM_rd5[2]_pad  ;
  input \CM_rd5[3]_pad  ;
  input \CM_rd5[4]_pad  ;
  input \CM_rd5[5]_pad  ;
  input \CM_rd5[6]_pad  ;
  input \CM_rd5[7]_pad  ;
  input \CM_rd5[8]_pad  ;
  input \CM_rd5[9]_pad  ;
  input \CM_rd6[0]_pad  ;
  input \CM_rd6[10]_pad  ;
  input \CM_rd6[11]_pad  ;
  input \CM_rd6[12]_pad  ;
  input \CM_rd6[13]_pad  ;
  input \CM_rd6[14]_pad  ;
  input \CM_rd6[15]_pad  ;
  input \CM_rd6[16]_pad  ;
  input \CM_rd6[17]_pad  ;
  input \CM_rd6[18]_pad  ;
  input \CM_rd6[19]_pad  ;
  input \CM_rd6[1]_pad  ;
  input \CM_rd6[20]_pad  ;
  input \CM_rd6[21]_pad  ;
  input \CM_rd6[22]_pad  ;
  input \CM_rd6[23]_pad  ;
  input \CM_rd6[2]_pad  ;
  input \CM_rd6[3]_pad  ;
  input \CM_rd6[4]_pad  ;
  input \CM_rd6[5]_pad  ;
  input \CM_rd6[6]_pad  ;
  input \CM_rd6[7]_pad  ;
  input \CM_rd6[8]_pad  ;
  input \CM_rd6[9]_pad  ;
  input \CM_rd7[0]_pad  ;
  input \CM_rd7[10]_pad  ;
  input \CM_rd7[11]_pad  ;
  input \CM_rd7[12]_pad  ;
  input \CM_rd7[13]_pad  ;
  input \CM_rd7[14]_pad  ;
  input \CM_rd7[15]_pad  ;
  input \CM_rd7[16]_pad  ;
  input \CM_rd7[17]_pad  ;
  input \CM_rd7[18]_pad  ;
  input \CM_rd7[19]_pad  ;
  input \CM_rd7[1]_pad  ;
  input \CM_rd7[20]_pad  ;
  input \CM_rd7[21]_pad  ;
  input \CM_rd7[22]_pad  ;
  input \CM_rd7[23]_pad  ;
  input \CM_rd7[2]_pad  ;
  input \CM_rd7[3]_pad  ;
  input \CM_rd7[4]_pad  ;
  input \CM_rd7[5]_pad  ;
  input \CM_rd7[6]_pad  ;
  input \CM_rd7[7]_pad  ;
  input \CM_rd7[8]_pad  ;
  input \CM_rd7[9]_pad  ;
  input \CM_rdm[0]_pad  ;
  input \CM_rdm[10]_pad  ;
  input \CM_rdm[11]_pad  ;
  input \CM_rdm[12]_pad  ;
  input \CM_rdm[13]_pad  ;
  input \CM_rdm[14]_pad  ;
  input \CM_rdm[15]_pad  ;
  input \CM_rdm[16]_pad  ;
  input \CM_rdm[17]_pad  ;
  input \CM_rdm[18]_pad  ;
  input \CM_rdm[19]_pad  ;
  input \CM_rdm[1]_pad  ;
  input \CM_rdm[20]_pad  ;
  input \CM_rdm[21]_pad  ;
  input \CM_rdm[22]_pad  ;
  input \CM_rdm[23]_pad  ;
  input \CM_rdm[2]_pad  ;
  input \CM_rdm[3]_pad  ;
  input \CM_rdm[4]_pad  ;
  input \CM_rdm[5]_pad  ;
  input \CM_rdm[6]_pad  ;
  input \CM_rdm[7]_pad  ;
  input \CM_rdm[8]_pad  ;
  input \CM_rdm[9]_pad  ;
  input \DM_rd0[0]_pad  ;
  input \DM_rd0[10]_pad  ;
  input \DM_rd0[11]_pad  ;
  input \DM_rd0[12]_pad  ;
  input \DM_rd0[13]_pad  ;
  input \DM_rd0[14]_pad  ;
  input \DM_rd0[15]_pad  ;
  input \DM_rd0[1]_pad  ;
  input \DM_rd0[2]_pad  ;
  input \DM_rd0[3]_pad  ;
  input \DM_rd0[4]_pad  ;
  input \DM_rd0[5]_pad  ;
  input \DM_rd0[6]_pad  ;
  input \DM_rd0[7]_pad  ;
  input \DM_rd0[8]_pad  ;
  input \DM_rd0[9]_pad  ;
  input \DM_rd1[0]_pad  ;
  input \DM_rd1[10]_pad  ;
  input \DM_rd1[11]_pad  ;
  input \DM_rd1[12]_pad  ;
  input \DM_rd1[13]_pad  ;
  input \DM_rd1[14]_pad  ;
  input \DM_rd1[15]_pad  ;
  input \DM_rd1[1]_pad  ;
  input \DM_rd1[2]_pad  ;
  input \DM_rd1[3]_pad  ;
  input \DM_rd1[4]_pad  ;
  input \DM_rd1[5]_pad  ;
  input \DM_rd1[6]_pad  ;
  input \DM_rd1[7]_pad  ;
  input \DM_rd1[8]_pad  ;
  input \DM_rd1[9]_pad  ;
  input \DM_rd2[0]_pad  ;
  input \DM_rd2[10]_pad  ;
  input \DM_rd2[11]_pad  ;
  input \DM_rd2[12]_pad  ;
  input \DM_rd2[13]_pad  ;
  input \DM_rd2[14]_pad  ;
  input \DM_rd2[15]_pad  ;
  input \DM_rd2[1]_pad  ;
  input \DM_rd2[2]_pad  ;
  input \DM_rd2[3]_pad  ;
  input \DM_rd2[4]_pad  ;
  input \DM_rd2[5]_pad  ;
  input \DM_rd2[6]_pad  ;
  input \DM_rd2[7]_pad  ;
  input \DM_rd2[8]_pad  ;
  input \DM_rd2[9]_pad  ;
  input \DM_rd3[0]_pad  ;
  input \DM_rd3[10]_pad  ;
  input \DM_rd3[11]_pad  ;
  input \DM_rd3[12]_pad  ;
  input \DM_rd3[13]_pad  ;
  input \DM_rd3[14]_pad  ;
  input \DM_rd3[15]_pad  ;
  input \DM_rd3[1]_pad  ;
  input \DM_rd3[2]_pad  ;
  input \DM_rd3[3]_pad  ;
  input \DM_rd3[4]_pad  ;
  input \DM_rd3[5]_pad  ;
  input \DM_rd3[6]_pad  ;
  input \DM_rd3[7]_pad  ;
  input \DM_rd3[8]_pad  ;
  input \DM_rd3[9]_pad  ;
  input \DM_rd4[0]_pad  ;
  input \DM_rd4[10]_pad  ;
  input \DM_rd4[11]_pad  ;
  input \DM_rd4[12]_pad  ;
  input \DM_rd4[13]_pad  ;
  input \DM_rd4[14]_pad  ;
  input \DM_rd4[15]_pad  ;
  input \DM_rd4[1]_pad  ;
  input \DM_rd4[2]_pad  ;
  input \DM_rd4[3]_pad  ;
  input \DM_rd4[4]_pad  ;
  input \DM_rd4[5]_pad  ;
  input \DM_rd4[6]_pad  ;
  input \DM_rd4[7]_pad  ;
  input \DM_rd4[8]_pad  ;
  input \DM_rd4[9]_pad  ;
  input \DM_rd5[0]_pad  ;
  input \DM_rd5[10]_pad  ;
  input \DM_rd5[11]_pad  ;
  input \DM_rd5[12]_pad  ;
  input \DM_rd5[13]_pad  ;
  input \DM_rd5[14]_pad  ;
  input \DM_rd5[15]_pad  ;
  input \DM_rd5[1]_pad  ;
  input \DM_rd5[2]_pad  ;
  input \DM_rd5[3]_pad  ;
  input \DM_rd5[4]_pad  ;
  input \DM_rd5[5]_pad  ;
  input \DM_rd5[6]_pad  ;
  input \DM_rd5[7]_pad  ;
  input \DM_rd5[8]_pad  ;
  input \DM_rd5[9]_pad  ;
  input \DM_rd6[0]_pad  ;
  input \DM_rd6[10]_pad  ;
  input \DM_rd6[11]_pad  ;
  input \DM_rd6[12]_pad  ;
  input \DM_rd6[13]_pad  ;
  input \DM_rd6[14]_pad  ;
  input \DM_rd6[15]_pad  ;
  input \DM_rd6[1]_pad  ;
  input \DM_rd6[2]_pad  ;
  input \DM_rd6[3]_pad  ;
  input \DM_rd6[4]_pad  ;
  input \DM_rd6[5]_pad  ;
  input \DM_rd6[6]_pad  ;
  input \DM_rd6[7]_pad  ;
  input \DM_rd6[8]_pad  ;
  input \DM_rd6[9]_pad  ;
  input \DM_rd7[0]_pad  ;
  input \DM_rd7[10]_pad  ;
  input \DM_rd7[11]_pad  ;
  input \DM_rd7[12]_pad  ;
  input \DM_rd7[13]_pad  ;
  input \DM_rd7[14]_pad  ;
  input \DM_rd7[15]_pad  ;
  input \DM_rd7[1]_pad  ;
  input \DM_rd7[2]_pad  ;
  input \DM_rd7[3]_pad  ;
  input \DM_rd7[4]_pad  ;
  input \DM_rd7[5]_pad  ;
  input \DM_rd7[6]_pad  ;
  input \DM_rd7[7]_pad  ;
  input \DM_rd7[8]_pad  ;
  input \DM_rd7[9]_pad  ;
  input \DM_rdm[0]_pad  ;
  input \DM_rdm[10]_pad  ;
  input \DM_rdm[11]_pad  ;
  input \DM_rdm[12]_pad  ;
  input \DM_rdm[13]_pad  ;
  input \DM_rdm[14]_pad  ;
  input \DM_rdm[15]_pad  ;
  input \DM_rdm[1]_pad  ;
  input \DM_rdm[2]_pad  ;
  input \DM_rdm[3]_pad  ;
  input \DM_rdm[4]_pad  ;
  input \DM_rdm[5]_pad  ;
  input \DM_rdm[6]_pad  ;
  input \DM_rdm[7]_pad  ;
  input \DM_rdm[8]_pad  ;
  input \DM_rdm[9]_pad  ;
  input IACKn_pad ;
  input \IRFS0_pad  ;
  input \IRFS1_pad  ;
  input \ISCLK0_pad  ;
  input \ISCLK1_pad  ;
  input \ITFS0_pad  ;
  input \ITFS1_pad  ;
  input \PIO_oe[0]_pad  ;
  input \PIO_oe[10]_pad  ;
  input \PIO_oe[11]_pad  ;
  input \PIO_oe[1]_pad  ;
  input \PIO_oe[2]_pad  ;
  input \PIO_oe[3]_pad  ;
  input \PIO_oe[4]_pad  ;
  input \PIO_oe[5]_pad  ;
  input \PIO_oe[6]_pad  ;
  input \PIO_oe[7]_pad  ;
  input \PIO_oe[8]_pad  ;
  input \PIO_oe[9]_pad  ;
  input \PIO_out[0]_pad  ;
  input \PIO_out[10]_pad  ;
  input \PIO_out[11]_pad  ;
  input \PIO_out[1]_pad  ;
  input \PIO_out[2]_pad  ;
  input \PIO_out[3]_pad  ;
  input \PIO_out[4]_pad  ;
  input \PIO_out[5]_pad  ;
  input \PIO_out[6]_pad  ;
  input \PIO_out[7]_pad  ;
  input \PIO_out[8]_pad  ;
  input \PIO_out[9]_pad  ;
  input PM_bdry_sel_pad ;
  input \PM_rd0[0]_pad  ;
  input \PM_rd0[10]_pad  ;
  input \PM_rd0[11]_pad  ;
  input \PM_rd0[12]_pad  ;
  input \PM_rd0[13]_pad  ;
  input \PM_rd0[14]_pad  ;
  input \PM_rd0[15]_pad  ;
  input \PM_rd0[1]_pad  ;
  input \PM_rd0[2]_pad  ;
  input \PM_rd0[3]_pad  ;
  input \PM_rd0[4]_pad  ;
  input \PM_rd0[5]_pad  ;
  input \PM_rd0[6]_pad  ;
  input \PM_rd0[7]_pad  ;
  input \PM_rd0[8]_pad  ;
  input \PM_rd0[9]_pad  ;
  input \PM_rd1[0]_pad  ;
  input \PM_rd1[10]_pad  ;
  input \PM_rd1[11]_pad  ;
  input \PM_rd1[12]_pad  ;
  input \PM_rd1[13]_pad  ;
  input \PM_rd1[14]_pad  ;
  input \PM_rd1[15]_pad  ;
  input \PM_rd1[1]_pad  ;
  input \PM_rd1[2]_pad  ;
  input \PM_rd1[3]_pad  ;
  input \PM_rd1[4]_pad  ;
  input \PM_rd1[5]_pad  ;
  input \PM_rd1[6]_pad  ;
  input \PM_rd1[7]_pad  ;
  input \PM_rd1[8]_pad  ;
  input \PM_rd1[9]_pad  ;
  input \PM_rd2[0]_pad  ;
  input \PM_rd2[10]_pad  ;
  input \PM_rd2[11]_pad  ;
  input \PM_rd2[12]_pad  ;
  input \PM_rd2[13]_pad  ;
  input \PM_rd2[14]_pad  ;
  input \PM_rd2[15]_pad  ;
  input \PM_rd2[1]_pad  ;
  input \PM_rd2[2]_pad  ;
  input \PM_rd2[3]_pad  ;
  input \PM_rd2[4]_pad  ;
  input \PM_rd2[5]_pad  ;
  input \PM_rd2[6]_pad  ;
  input \PM_rd2[7]_pad  ;
  input \PM_rd2[8]_pad  ;
  input \PM_rd2[9]_pad  ;
  input \PM_rd3[0]_pad  ;
  input \PM_rd3[10]_pad  ;
  input \PM_rd3[11]_pad  ;
  input \PM_rd3[12]_pad  ;
  input \PM_rd3[13]_pad  ;
  input \PM_rd3[14]_pad  ;
  input \PM_rd3[15]_pad  ;
  input \PM_rd3[1]_pad  ;
  input \PM_rd3[2]_pad  ;
  input \PM_rd3[3]_pad  ;
  input \PM_rd3[4]_pad  ;
  input \PM_rd3[5]_pad  ;
  input \PM_rd3[6]_pad  ;
  input \PM_rd3[7]_pad  ;
  input \PM_rd3[8]_pad  ;
  input \PM_rd3[9]_pad  ;
  input \PM_rd4[0]_pad  ;
  input \PM_rd4[10]_pad  ;
  input \PM_rd4[11]_pad  ;
  input \PM_rd4[12]_pad  ;
  input \PM_rd4[13]_pad  ;
  input \PM_rd4[14]_pad  ;
  input \PM_rd4[15]_pad  ;
  input \PM_rd4[1]_pad  ;
  input \PM_rd4[2]_pad  ;
  input \PM_rd4[3]_pad  ;
  input \PM_rd4[4]_pad  ;
  input \PM_rd4[5]_pad  ;
  input \PM_rd4[6]_pad  ;
  input \PM_rd4[7]_pad  ;
  input \PM_rd4[8]_pad  ;
  input \PM_rd4[9]_pad  ;
  input \PM_rd5[0]_pad  ;
  input \PM_rd5[10]_pad  ;
  input \PM_rd5[11]_pad  ;
  input \PM_rd5[12]_pad  ;
  input \PM_rd5[13]_pad  ;
  input \PM_rd5[14]_pad  ;
  input \PM_rd5[15]_pad  ;
  input \PM_rd5[1]_pad  ;
  input \PM_rd5[2]_pad  ;
  input \PM_rd5[3]_pad  ;
  input \PM_rd5[4]_pad  ;
  input \PM_rd5[5]_pad  ;
  input \PM_rd5[6]_pad  ;
  input \PM_rd5[7]_pad  ;
  input \PM_rd5[8]_pad  ;
  input \PM_rd5[9]_pad  ;
  input \PM_rd6[0]_pad  ;
  input \PM_rd6[10]_pad  ;
  input \PM_rd6[11]_pad  ;
  input \PM_rd6[12]_pad  ;
  input \PM_rd6[13]_pad  ;
  input \PM_rd6[14]_pad  ;
  input \PM_rd6[15]_pad  ;
  input \PM_rd6[1]_pad  ;
  input \PM_rd6[2]_pad  ;
  input \PM_rd6[3]_pad  ;
  input \PM_rd6[4]_pad  ;
  input \PM_rd6[5]_pad  ;
  input \PM_rd6[6]_pad  ;
  input \PM_rd6[7]_pad  ;
  input \PM_rd6[8]_pad  ;
  input \PM_rd6[9]_pad  ;
  input \PM_rd7[0]_pad  ;
  input \PM_rd7[10]_pad  ;
  input \PM_rd7[11]_pad  ;
  input \PM_rd7[12]_pad  ;
  input \PM_rd7[13]_pad  ;
  input \PM_rd7[14]_pad  ;
  input \PM_rd7[15]_pad  ;
  input \PM_rd7[1]_pad  ;
  input \PM_rd7[2]_pad  ;
  input \PM_rd7[3]_pad  ;
  input \PM_rd7[4]_pad  ;
  input \PM_rd7[5]_pad  ;
  input \PM_rd7[6]_pad  ;
  input \PM_rd7[7]_pad  ;
  input \PM_rd7[8]_pad  ;
  input \PM_rd7[9]_pad  ;
  input PWDACK_pad ;
  input T_BMODE_pad ;
  input T_BRn_pad ;
  input T_CLKI_OSC_pad ;
  input T_CLKI_PLL_pad ;
  input \T_ED[0]_pad  ;
  input \T_ED[10]_pad  ;
  input \T_ED[11]_pad  ;
  input \T_ED[12]_pad  ;
  input \T_ED[13]_pad  ;
  input \T_ED[14]_pad  ;
  input \T_ED[15]_pad  ;
  input \T_ED[1]_pad  ;
  input \T_ED[2]_pad  ;
  input \T_ED[3]_pad  ;
  input \T_ED[4]_pad  ;
  input \T_ED[5]_pad  ;
  input \T_ED[6]_pad  ;
  input \T_ED[7]_pad  ;
  input \T_ED[8]_pad  ;
  input \T_ED[9]_pad  ;
  input T_ICE_RSTn_pad ;
  input T_ID_pad ;
  input T_IMS_pad ;
  input T_IRDn_pad ;
  input \T_IRQ0n_pad  ;
  input \T_IRQ1n_pad  ;
  input \T_IRQ2n_pad  ;
  input \T_IRQE0n_pad  ;
  input \T_IRQE1n_pad  ;
  input \T_IRQL1n_pad  ;
  input T_ISn_pad ;
  input T_IWRn_pad ;
  input T_MMAP_pad ;
  input \T_PIOin[0]_pad  ;
  input \T_PIOin[10]_pad  ;
  input \T_PIOin[11]_pad  ;
  input \T_PIOin[1]_pad  ;
  input \T_PIOin[2]_pad  ;
  input \T_PIOin[3]_pad  ;
  input \T_PIOin[4]_pad  ;
  input \T_PIOin[5]_pad  ;
  input \T_PIOin[6]_pad  ;
  input \T_PIOin[7]_pad  ;
  input \T_PIOin[8]_pad  ;
  input \T_PIOin[9]_pad  ;
  input T_PWDn_pad ;
  input \T_RD0_pad  ;
  input \T_RD1_pad  ;
  input \T_RFS0_pad  ;
  input \T_RFS1_pad  ;
  input T_RSTn_pad ;
  input \T_SCLK0_pad  ;
  input \T_SCLK1_pad  ;
  input T_Sel_PLL_pad ;
  input \T_TFS0_pad  ;
  input \T_TFS1_pad  ;
  input \T_TMODE[0]_pad  ;
  input \T_TMODE[1]_pad  ;
  input \auctl_BSack_reg/NET0131  ;
  input \auctl_DSack_reg/NET0131  ;
  input \auctl_R0Sack_reg/NET0131  ;
  input \auctl_R1Sack_reg/NET0131  ;
  input \auctl_RST_reg/P0001  ;
  input \auctl_STEAL_reg/NET0131  ;
  input \auctl_T0Sack_reg/NET0131  ;
  input \auctl_T1Sack_reg/NET0131  ;
  input \bdma_BCTL_reg[0]/NET0131  ;
  input \bdma_BCTL_reg[10]/NET0131  ;
  input \bdma_BCTL_reg[11]/NET0131  ;
  input \bdma_BCTL_reg[12]/NET0131  ;
  input \bdma_BCTL_reg[13]/NET0131  ;
  input \bdma_BCTL_reg[14]/NET0131  ;
  input \bdma_BCTL_reg[15]/NET0131  ;
  input \bdma_BCTL_reg[1]/NET0131  ;
  input \bdma_BCTL_reg[2]/NET0131  ;
  input \bdma_BCTL_reg[3]/NET0131  ;
  input \bdma_BCTL_reg[4]/NET0131  ;
  input \bdma_BCTL_reg[5]/NET0131  ;
  input \bdma_BCTL_reg[6]/NET0131  ;
  input \bdma_BCTL_reg[7]/NET0131  ;
  input \bdma_BCTL_reg[8]/NET0131  ;
  input \bdma_BCTL_reg[9]/NET0131  ;
  input \bdma_BDMA_boot_reg/NET0131_reg_syn_10  ;
  input \bdma_BDMA_boot_reg/NET0131_reg_syn_2  ;
  input \bdma_BDMA_boot_reg/NET0131_reg_syn_8  ;
  input \bdma_BDMAmode_reg/NET0131  ;
  input \bdma_BEAD_reg[0]/NET0131  ;
  input \bdma_BEAD_reg[10]/NET0131  ;
  input \bdma_BEAD_reg[11]/NET0131  ;
  input \bdma_BEAD_reg[12]/NET0131  ;
  input \bdma_BEAD_reg[13]/NET0131  ;
  input \bdma_BEAD_reg[1]/NET0131  ;
  input \bdma_BEAD_reg[2]/NET0131  ;
  input \bdma_BEAD_reg[3]/NET0131  ;
  input \bdma_BEAD_reg[4]/NET0131  ;
  input \bdma_BEAD_reg[5]/NET0131  ;
  input \bdma_BEAD_reg[6]/NET0131  ;
  input \bdma_BEAD_reg[7]/NET0131  ;
  input \bdma_BEAD_reg[8]/NET0131  ;
  input \bdma_BEAD_reg[9]/NET0131  ;
  input \bdma_BIAD_reg[0]/NET0131  ;
  input \bdma_BIAD_reg[10]/NET0131  ;
  input \bdma_BIAD_reg[11]/NET0131  ;
  input \bdma_BIAD_reg[12]/NET0131  ;
  input \bdma_BIAD_reg[13]/NET0131  ;
  input \bdma_BIAD_reg[1]/NET0131  ;
  input \bdma_BIAD_reg[2]/NET0131  ;
  input \bdma_BIAD_reg[3]/NET0131  ;
  input \bdma_BIAD_reg[4]/NET0131  ;
  input \bdma_BIAD_reg[5]/NET0131  ;
  input \bdma_BIAD_reg[6]/NET0131  ;
  input \bdma_BIAD_reg[7]/NET0131  ;
  input \bdma_BIAD_reg[8]/NET0131  ;
  input \bdma_BIAD_reg[9]/NET0131  ;
  input \bdma_BM_cyc_reg/P0001  ;
  input \bdma_BMcyc_del_reg/P0001  ;
  input \bdma_BOVL_reg[0]/NET0131  ;
  input \bdma_BOVL_reg[10]/NET0131  ;
  input \bdma_BOVL_reg[11]/NET0131  ;
  input \bdma_BOVL_reg[1]/NET0131  ;
  input \bdma_BOVL_reg[2]/NET0131  ;
  input \bdma_BOVL_reg[3]/NET0131  ;
  input \bdma_BOVL_reg[4]/NET0131  ;
  input \bdma_BOVL_reg[5]/NET0131  ;
  input \bdma_BOVL_reg[6]/NET0131  ;
  input \bdma_BOVL_reg[7]/NET0131  ;
  input \bdma_BOVL_reg[8]/NET0131  ;
  input \bdma_BOVL_reg[9]/NET0131  ;
  input \bdma_BRST_s2_reg/NET0131  ;
  input \bdma_BRdataBUF_reg[0]/P0001  ;
  input \bdma_BRdataBUF_reg[10]/P0001  ;
  input \bdma_BRdataBUF_reg[11]/P0001  ;
  input \bdma_BRdataBUF_reg[12]/P0001  ;
  input \bdma_BRdataBUF_reg[13]/P0001  ;
  input \bdma_BRdataBUF_reg[14]/P0001  ;
  input \bdma_BRdataBUF_reg[15]/P0001  ;
  input \bdma_BRdataBUF_reg[16]/P0001  ;
  input \bdma_BRdataBUF_reg[17]/P0001  ;
  input \bdma_BRdataBUF_reg[18]/P0001  ;
  input \bdma_BRdataBUF_reg[19]/P0001  ;
  input \bdma_BRdataBUF_reg[1]/P0001  ;
  input \bdma_BRdataBUF_reg[20]/P0001  ;
  input \bdma_BRdataBUF_reg[21]/P0001  ;
  input \bdma_BRdataBUF_reg[22]/P0001  ;
  input \bdma_BRdataBUF_reg[23]/P0001  ;
  input \bdma_BRdataBUF_reg[2]/P0001  ;
  input \bdma_BRdataBUF_reg[3]/P0001  ;
  input \bdma_BRdataBUF_reg[4]/P0001  ;
  input \bdma_BRdataBUF_reg[5]/P0001  ;
  input \bdma_BRdataBUF_reg[6]/P0001  ;
  input \bdma_BRdataBUF_reg[7]/P0001  ;
  input \bdma_BRdataBUF_reg[8]/P0001  ;
  input \bdma_BRdataBUF_reg[9]/P0001  ;
  input \bdma_BSreq_reg/NET0131  ;
  input \bdma_BWCOUNT_reg[0]/NET0131  ;
  input \bdma_BWCOUNT_reg[10]/NET0131  ;
  input \bdma_BWCOUNT_reg[11]/NET0131  ;
  input \bdma_BWCOUNT_reg[12]/NET0131  ;
  input \bdma_BWCOUNT_reg[13]/NET0131  ;
  input \bdma_BWCOUNT_reg[1]/NET0131  ;
  input \bdma_BWCOUNT_reg[2]/NET0131  ;
  input \bdma_BWCOUNT_reg[3]/NET0131  ;
  input \bdma_BWCOUNT_reg[4]/NET0131  ;
  input \bdma_BWCOUNT_reg[5]/NET0131_reg_syn_2  ;
  input \bdma_BWCOUNT_reg[5]/NET0131_reg_syn_8  ;
  input \bdma_BWCOUNT_reg[6]/NET0131  ;
  input \bdma_BWCOUNT_reg[7]/NET0131  ;
  input \bdma_BWCOUNT_reg[8]/NET0131  ;
  input \bdma_BWCOUNT_reg[9]/NET0131  ;
  input \bdma_BWRn_reg/NET0131  ;
  input \bdma_BWcnt_reg[0]/NET0131  ;
  input \bdma_BWcnt_reg[1]/NET0131  ;
  input \bdma_BWcnt_reg[2]/NET0131  ;
  input \bdma_BWcnt_reg[3]/NET0131  ;
  input \bdma_BWcnt_reg[4]/NET0131  ;
  input \bdma_BWdataBUF_h_reg[0]/P0001  ;
  input \bdma_BWdataBUF_h_reg[10]/P0001  ;
  input \bdma_BWdataBUF_h_reg[11]/P0001  ;
  input \bdma_BWdataBUF_h_reg[12]/P0001  ;
  input \bdma_BWdataBUF_h_reg[13]/P0001  ;
  input \bdma_BWdataBUF_h_reg[14]/P0001  ;
  input \bdma_BWdataBUF_h_reg[15]/P0001  ;
  input \bdma_BWdataBUF_h_reg[16]/P0001  ;
  input \bdma_BWdataBUF_h_reg[17]/P0001  ;
  input \bdma_BWdataBUF_h_reg[18]/P0001  ;
  input \bdma_BWdataBUF_h_reg[19]/P0001  ;
  input \bdma_BWdataBUF_h_reg[1]/P0001  ;
  input \bdma_BWdataBUF_h_reg[20]/P0001  ;
  input \bdma_BWdataBUF_h_reg[21]/P0001  ;
  input \bdma_BWdataBUF_h_reg[22]/P0001  ;
  input \bdma_BWdataBUF_h_reg[23]/P0001  ;
  input \bdma_BWdataBUF_h_reg[2]/P0001  ;
  input \bdma_BWdataBUF_h_reg[3]/P0001  ;
  input \bdma_BWdataBUF_h_reg[4]/P0001  ;
  input \bdma_BWdataBUF_h_reg[5]/P0001  ;
  input \bdma_BWdataBUF_h_reg[6]/P0001  ;
  input \bdma_BWdataBUF_h_reg[7]/P0001  ;
  input \bdma_BWdataBUF_h_reg[8]/P0001  ;
  input \bdma_BWdataBUF_h_reg[9]/P0001  ;
  input \bdma_BWdataBUF_reg[0]/P0001  ;
  input \bdma_BWdataBUF_reg[1]/P0001  ;
  input \bdma_BWdataBUF_reg[2]/P0001  ;
  input \bdma_BWdataBUF_reg[3]/P0001  ;
  input \bdma_BWdataBUF_reg[4]/P0001  ;
  input \bdma_BWdataBUF_reg[5]/P0001  ;
  input \bdma_BWdataBUF_reg[6]/P0001  ;
  input \bdma_BWdataBUF_reg[7]/P0001  ;
  input \bdma_CMcnt_reg[0]/NET0131  ;
  input \bdma_CMcnt_reg[1]/NET0131  ;
  input \bdma_DM_2nd_reg/NET0131  ;
  input \bdma_RST_pin_reg/P0001  ;
  input \bdma_WRlat_reg/P0001  ;
  input \clkc_Awake_reg/NET0131  ;
  input \clkc_CLKOUT_reg/NET0131  ;
  input \clkc_CTR_cnt_reg[0]/NET0131  ;
  input \clkc_CTR_cnt_reg[1]/NET0131  ;
  input \clkc_Cnt128_reg/NET0131  ;
  input \clkc_Cnt4096_reg/NET0131  ;
  input \clkc_Cnt4096_s1_reg/NET0131  ;
  input \clkc_Cnt4096_s2_reg/NET0131  ;
  input \clkc_DSPoff_reg/NET0131  ;
  input \clkc_OSCoff_reg/NET0131  ;
  input \clkc_OSCoff_set_reg/P0001  ;
  input \clkc_OUTcnt_reg[0]/NET0131  ;
  input \clkc_OUTcnt_reg[1]/NET0131  ;
  input \clkc_OUTcnt_reg[2]/NET0131  ;
  input \clkc_OUTcnt_reg[3]/NET0131  ;
  input \clkc_OUTcnt_reg[4]/NET0131  ;
  input \clkc_OUTcnt_reg[5]/NET0131  ;
  input \clkc_OUTcnt_reg[6]/NET0131  ;
  input \clkc_RSTtext_reg/P0001  ;
  input \clkc_SIDLE_s1_reg/NET0131  ;
  input \clkc_SIDLE_s2_reg/NET0131  ;
  input \clkc_SLEEP_reg/NET0131  ;
  input \clkc_STBY_reg/NET0131  ;
  input \clkc_STDcnt_reg[0]/NET0131  ;
  input \clkc_STDcnt_reg[10]/NET0131  ;
  input \clkc_STDcnt_reg[1]/NET0131  ;
  input \clkc_STDcnt_reg[2]/NET0131  ;
  input \clkc_STDcnt_reg[3]/NET0131  ;
  input \clkc_STDcnt_reg[4]/NET0131  ;
  input \clkc_STDcnt_reg[5]/NET0131  ;
  input \clkc_STDcnt_reg[6]/NET0131  ;
  input \clkc_STDcnt_reg[7]/NET0131  ;
  input \clkc_STDcnt_reg[8]/NET0131  ;
  input \clkc_STDcnt_reg[9]/NET0131  ;
  input \clkc_SlowDn_reg/NET0131  ;
  input \clkc_SlowDn_s1_reg/P0001  ;
  input \clkc_SlowDn_s2_reg/P0001  ;
  input \clkc_ckSTDCLK_STDCLK_reg_Q_reg/NET0131  ;
  input \clkc_ckr_reg_DO_reg[0]/NET0131  ;
  input \clkc_ckr_reg_DO_reg[10]/NET0131  ;
  input \clkc_ckr_reg_DO_reg[11]/NET0131  ;
  input \clkc_ckr_reg_DO_reg[12]/NET0131  ;
  input \clkc_ckr_reg_DO_reg[13]/NET0131  ;
  input \clkc_ckr_reg_DO_reg[14]/NET0131  ;
  input \clkc_ckr_reg_DO_reg[15]/NET0131  ;
  input \clkc_ckr_reg_DO_reg[1]/NET0131  ;
  input \clkc_ckr_reg_DO_reg[2]/NET0131  ;
  input \clkc_ckr_reg_DO_reg[3]/NET0131  ;
  input \clkc_ckr_reg_DO_reg[4]/NET0131  ;
  input \clkc_ckr_reg_DO_reg[5]/NET0131  ;
  input \clkc_ckr_reg_DO_reg[6]/NET0131  ;
  input \clkc_ckr_reg_DO_reg[7]/NET0131  ;
  input \clkc_ckr_reg_DO_reg[8]/NET0131  ;
  input \clkc_ckr_reg_DO_reg[9]/NET0131  ;
  input \clkc_oscntr_reg_DO_reg[0]/NET0131  ;
  input \clkc_oscntr_reg_DO_reg[10]/NET0131  ;
  input \clkc_oscntr_reg_DO_reg[11]/NET0131  ;
  input \clkc_oscntr_reg_DO_reg[1]/NET0131  ;
  input \clkc_oscntr_reg_DO_reg[2]/NET0131  ;
  input \clkc_oscntr_reg_DO_reg[3]/NET0131  ;
  input \clkc_oscntr_reg_DO_reg[4]/NET0131  ;
  input \clkc_oscntr_reg_DO_reg[5]/NET0131  ;
  input \clkc_oscntr_reg_DO_reg[6]/NET0131  ;
  input \clkc_oscntr_reg_DO_reg[7]/NET0131  ;
  input \clkc_oscntr_reg_DO_reg[8]/NET0131  ;
  input \clkc_oscntr_reg_DO_reg[9]/NET0131  ;
  input \core_c_dec_ALUop_E_reg/P0001  ;
  input \core_c_dec_BR_Ed_reg/P0001  ;
  input \core_c_dec_Call_Ed_reg/P0001  ;
  input \core_c_dec_DIVQ_E_reg/P0001  ;
  input \core_c_dec_DIVS_E_reg/P0001  ;
  input \core_c_dec_DU_Eg_reg/P0001  ;
  input \core_c_dec_Double_E_reg/P0001  ;
  input \core_c_dec_Dummy_E_reg/NET0131  ;
  input \core_c_dec_EXIT_E_reg/P0001  ;
  input \core_c_dec_IDLE_Eg_reg/P0001  ;
  input \core_c_dec_IRE_reg[0]/NET0131  ;
  input \core_c_dec_IRE_reg[10]/NET0131  ;
  input \core_c_dec_IRE_reg[11]/NET0131  ;
  input \core_c_dec_IRE_reg[12]/NET0131  ;
  input \core_c_dec_IRE_reg[13]/NET0131  ;
  input \core_c_dec_IRE_reg[14]/NET0131  ;
  input \core_c_dec_IRE_reg[15]/NET0131  ;
  input \core_c_dec_IRE_reg[16]/NET0131  ;
  input \core_c_dec_IRE_reg[17]/NET0131  ;
  input \core_c_dec_IRE_reg[18]/NET0131  ;
  input \core_c_dec_IRE_reg[19]/NET0131  ;
  input \core_c_dec_IRE_reg[1]/NET0131  ;
  input \core_c_dec_IRE_reg[2]/NET0131  ;
  input \core_c_dec_IRE_reg[3]/NET0131  ;
  input \core_c_dec_IRE_reg[4]/NET0131  ;
  input \core_c_dec_IRE_reg[5]/NET0131  ;
  input \core_c_dec_IRE_reg[6]/NET0131  ;
  input \core_c_dec_IRE_reg[7]/NET0131  ;
  input \core_c_dec_IRE_reg[8]/NET0131  ;
  input \core_c_dec_IRE_reg[9]/NET0131  ;
  input \core_c_dec_IR_reg[0]/NET0131  ;
  input \core_c_dec_IR_reg[10]/NET0131  ;
  input \core_c_dec_IR_reg[11]/NET0131  ;
  input \core_c_dec_IR_reg[12]/NET0131  ;
  input \core_c_dec_IR_reg[13]/NET0131  ;
  input \core_c_dec_IR_reg[14]/NET0131  ;
  input \core_c_dec_IR_reg[15]/NET0131  ;
  input \core_c_dec_IR_reg[16]/NET0131  ;
  input \core_c_dec_IR_reg[17]/NET0131  ;
  input \core_c_dec_IR_reg[18]/NET0131  ;
  input \core_c_dec_IR_reg[19]/NET0131  ;
  input \core_c_dec_IR_reg[1]/NET0131  ;
  input \core_c_dec_IR_reg[20]/NET0131  ;
  input \core_c_dec_IR_reg[21]/NET0131  ;
  input \core_c_dec_IR_reg[22]/NET0131  ;
  input \core_c_dec_IR_reg[23]/NET0131  ;
  input \core_c_dec_IR_reg[2]/NET0131  ;
  input \core_c_dec_IR_reg[3]/NET0131  ;
  input \core_c_dec_IR_reg[4]/NET0131  ;
  input \core_c_dec_IR_reg[5]/NET0131  ;
  input \core_c_dec_IR_reg[6]/NET0131  ;
  input \core_c_dec_IR_reg[7]/NET0131  ;
  input \core_c_dec_IR_reg[8]/NET0131  ;
  input \core_c_dec_IR_reg[9]/NET0131  ;
  input \core_c_dec_Long_Cg_reg/P0001  ;
  input \core_c_dec_Long_Eg_reg/P0001  ;
  input \core_c_dec_MACdep_Eg_reg/P0001  ;
  input \core_c_dec_MACop_E_reg/P0001  ;
  input \core_c_dec_MFALU_Ei_reg/NET0131  ;
  input \core_c_dec_MFAR_E_reg/P0001  ;
  input \core_c_dec_MFASTAT_E_reg/P0001  ;
  input \core_c_dec_MFAX0_E_reg/P0001  ;
  input \core_c_dec_MFAX1_E_reg/P0001  ;
  input \core_c_dec_MFAY0_E_reg/P0001  ;
  input \core_c_dec_MFAY1_E_reg/P0001  ;
  input \core_c_dec_MFCNTR_E_reg/P0001  ;
  input \core_c_dec_MFDAG1_Ei_reg/NET0131  ;
  input \core_c_dec_MFDAG2_Ei_reg/NET0131  ;
  input \core_c_dec_MFDMOVL_E_reg/P0001  ;
  input \core_c_dec_MFICNTL_E_reg/P0001  ;
  input \core_c_dec_MFIDR_E_reg/P0001  ;
  input \core_c_dec_MFIMASK_E_reg/P0001  ;
  input \core_c_dec_MFIreg_E_reg[0]/P0001  ;
  input \core_c_dec_MFIreg_E_reg[1]/P0001  ;
  input \core_c_dec_MFIreg_E_reg[2]/P0001  ;
  input \core_c_dec_MFIreg_E_reg[3]/P0001  ;
  input \core_c_dec_MFIreg_E_reg[4]/P0001  ;
  input \core_c_dec_MFIreg_E_reg[5]/P0001  ;
  input \core_c_dec_MFIreg_E_reg[6]/P0001  ;
  input \core_c_dec_MFIreg_E_reg[7]/P0001  ;
  input \core_c_dec_MFLreg_E_reg[0]/P0001  ;
  input \core_c_dec_MFLreg_E_reg[1]/P0001  ;
  input \core_c_dec_MFLreg_E_reg[2]/P0001  ;
  input \core_c_dec_MFLreg_E_reg[3]/P0001  ;
  input \core_c_dec_MFLreg_E_reg[4]/P0001  ;
  input \core_c_dec_MFLreg_E_reg[5]/P0001  ;
  input \core_c_dec_MFLreg_E_reg[6]/P0001  ;
  input \core_c_dec_MFLreg_E_reg[7]/P0001  ;
  input \core_c_dec_MFMAC_Ei_reg/NET0131  ;
  input \core_c_dec_MFMR0_E_reg/P0001  ;
  input \core_c_dec_MFMR1_E_reg/P0001  ;
  input \core_c_dec_MFMR2_E_reg/P0001  ;
  input \core_c_dec_MFMSTAT_E_reg/P0001  ;
  input \core_c_dec_MFMX0_E_reg/P0001  ;
  input \core_c_dec_MFMX1_E_reg/P0001  ;
  input \core_c_dec_MFMY0_E_reg/P0001  ;
  input \core_c_dec_MFMY1_E_reg/P0001  ;
  input \core_c_dec_MFMreg_E_reg[0]/P0001  ;
  input \core_c_dec_MFMreg_E_reg[1]/P0001  ;
  input \core_c_dec_MFMreg_E_reg[2]/P0001  ;
  input \core_c_dec_MFMreg_E_reg[3]/P0001  ;
  input \core_c_dec_MFMreg_E_reg[4]/P0001  ;
  input \core_c_dec_MFMreg_E_reg[5]/P0001  ;
  input \core_c_dec_MFMreg_E_reg[6]/P0001  ;
  input \core_c_dec_MFMreg_E_reg[7]/P0001  ;
  input \core_c_dec_MFPMOVL_E_reg/P0001  ;
  input \core_c_dec_MFPSQ_Ei_reg/NET0131  ;
  input \core_c_dec_MFRX0_E_reg/P0001  ;
  input \core_c_dec_MFRX1_E_reg/P0001  ;
  input \core_c_dec_MFSB_E_reg/P0001  ;
  input \core_c_dec_MFSE_E_reg/P0001  ;
  input \core_c_dec_MFSHT_Ei_reg/NET0131  ;
  input \core_c_dec_MFSI_E_reg/P0001  ;
  input \core_c_dec_MFSPT_Ei_reg/NET0131  ;
  input \core_c_dec_MFSR0_E_reg/P0001  ;
  input \core_c_dec_MFSR1_E_reg/P0001  ;
  input \core_c_dec_MFSSTAT_E_reg/P0001  ;
  input \core_c_dec_MFTX0_E_reg/P0001  ;
  input \core_c_dec_MFTX1_E_reg/P0001  ;
  input \core_c_dec_MFtoppcs_Eg_reg/P0001  ;
  input \core_c_dec_MTAR_E_reg/P0001  ;
  input \core_c_dec_MTASTAT_E_reg/P0001  ;
  input \core_c_dec_MTAX0_E_reg/P0001  ;
  input \core_c_dec_MTAX1_E_reg/P0001  ;
  input \core_c_dec_MTAY0_E_reg/P0001  ;
  input \core_c_dec_MTAY1_E_reg/P0001  ;
  input \core_c_dec_MTCNTR_Eg_reg/P0001  ;
  input \core_c_dec_MTDMOVL_E_reg/P0001  ;
  input \core_c_dec_MTICNTL_Eg_reg/P0001  ;
  input \core_c_dec_MTIDR_E_reg/P0001  ;
  input \core_c_dec_MTIFC_Eg_reg/P0001  ;
  input \core_c_dec_MTIMASK_Eg_reg/P0001  ;
  input \core_c_dec_MTIreg_E_reg[0]/P0001  ;
  input \core_c_dec_MTIreg_E_reg[1]/P0001  ;
  input \core_c_dec_MTIreg_E_reg[2]/P0001  ;
  input \core_c_dec_MTIreg_E_reg[3]/P0001  ;
  input \core_c_dec_MTIreg_E_reg[4]/P0001  ;
  input \core_c_dec_MTIreg_E_reg[5]/P0001  ;
  input \core_c_dec_MTIreg_E_reg[6]/P0001  ;
  input \core_c_dec_MTIreg_E_reg[7]/P0001  ;
  input \core_c_dec_MTLreg_E_reg[0]/P0001  ;
  input \core_c_dec_MTLreg_E_reg[1]/P0001  ;
  input \core_c_dec_MTLreg_E_reg[2]/P0001  ;
  input \core_c_dec_MTLreg_E_reg[3]/P0001  ;
  input \core_c_dec_MTLreg_E_reg[4]/P0001  ;
  input \core_c_dec_MTLreg_E_reg[5]/P0001  ;
  input \core_c_dec_MTLreg_E_reg[6]/P0001  ;
  input \core_c_dec_MTLreg_E_reg[7]/P0001  ;
  input \core_c_dec_MTMR0_E_reg/P0001  ;
  input \core_c_dec_MTMR1_E_reg/P0001  ;
  input \core_c_dec_MTMR2_E_reg/P0001  ;
  input \core_c_dec_MTMSTAT_Eg_reg/P0001  ;
  input \core_c_dec_MTMX0_E_reg/P0001  ;
  input \core_c_dec_MTMX1_E_reg/P0001  ;
  input \core_c_dec_MTMY0_E_reg/P0001  ;
  input \core_c_dec_MTMY1_E_reg/P0001  ;
  input \core_c_dec_MTMreg_E_reg[0]/P0001  ;
  input \core_c_dec_MTMreg_E_reg[1]/P0001  ;
  input \core_c_dec_MTMreg_E_reg[2]/P0001  ;
  input \core_c_dec_MTMreg_E_reg[3]/P0001  ;
  input \core_c_dec_MTMreg_E_reg[4]/P0001  ;
  input \core_c_dec_MTMreg_E_reg[5]/P0001  ;
  input \core_c_dec_MTMreg_E_reg[6]/P0001  ;
  input \core_c_dec_MTMreg_E_reg[7]/P0001  ;
  input \core_c_dec_MTOWRCNTR_Eg_reg/P0001  ;
  input \core_c_dec_MTPMOVL_E_reg/P0001  ;
  input \core_c_dec_MTRX0_E_reg/P0001  ;
  input \core_c_dec_MTRX1_E_reg/P0001  ;
  input \core_c_dec_MTSB_E_reg/P0001  ;
  input \core_c_dec_MTSE_E_reg/P0001  ;
  input \core_c_dec_MTSI_E_reg/P0001  ;
  input \core_c_dec_MTSR0_E_reg/P0001  ;
  input \core_c_dec_MTSR1_E_reg/P0001  ;
  input \core_c_dec_MTTX0_E_reg/P0001  ;
  input \core_c_dec_MTTX1_E_reg/P0001  ;
  input \core_c_dec_MTtoppcs_Eg_reg/P0001  ;
  input \core_c_dec_Modctl_Eg_reg/P0001  ;
  input \core_c_dec_MpopLP_Eg_reg/P0001  ;
  input \core_c_dec_NOP_E_reg/P0001  ;
  input \core_c_dec_Nrti_Ed_reg/P0001  ;
  input \core_c_dec_Nseq_Ed_reg/P0001  ;
  input \core_c_dec_PPclr_reg/P0001  ;
  input \core_c_dec_Post1_E_reg/P0001  ;
  input \core_c_dec_Post2_E_reg/P0001  ;
  input \core_c_dec_Prderr_Cg_reg/NET0131  ;
  input \core_c_dec_RET_Ed_reg/P0001  ;
  input \core_c_dec_RTI_Ed_reg/P0001  ;
  input \core_c_dec_SHTop_E_reg/P0001  ;
  input \core_c_dec_Stkctl_Eg_reg/P0001  ;
  input \core_c_dec_Usecond_E_reg/P0001  ;
  input \core_c_dec_accCM_E_reg/NET0131  ;
  input \core_c_dec_accPM_E_reg/P0001  ;
  input \core_c_dec_cdAM_E_reg/P0001  ;
  input \core_c_dec_imSHT_E_reg/P0001  ;
  input \core_c_dec_imm14_E_reg/P0001  ;
  input \core_c_dec_imm16_E_reg/P0001  ;
  input \core_c_dec_pMFALU_Ei_reg/NET0131  ;
  input \core_c_dec_pMFMAC_Ei_reg/NET0131  ;
  input \core_c_dec_pMFSHT_Ei_reg/NET0131  ;
  input \core_c_dec_rdCM_E_reg/NET0131  ;
  input \core_c_dec_satMR_E_reg/P0001  ;
  input \core_c_dec_updAF_E_reg/P0001  ;
  input \core_c_dec_updAR_E_reg/P0001  ;
  input \core_c_dec_updMF_E_reg/P0001  ;
  input \core_c_dec_updMR_E_reg/P0001  ;
  input \core_c_dec_updSR_E_reg/P0001  ;
  input \core_c_psq_CE_reg/NET0131  ;
  input \core_c_psq_CNTR_reg_DO_reg[0]/NET0131  ;
  input \core_c_psq_CNTR_reg_DO_reg[10]/NET0131  ;
  input \core_c_psq_CNTR_reg_DO_reg[11]/NET0131  ;
  input \core_c_psq_CNTR_reg_DO_reg[12]/NET0131  ;
  input \core_c_psq_CNTR_reg_DO_reg[13]/NET0131  ;
  input \core_c_psq_CNTR_reg_DO_reg[1]/NET0131  ;
  input \core_c_psq_CNTR_reg_DO_reg[2]/NET0131  ;
  input \core_c_psq_CNTR_reg_DO_reg[3]/NET0131  ;
  input \core_c_psq_CNTR_reg_DO_reg[4]/NET0131  ;
  input \core_c_psq_CNTR_reg_DO_reg[5]/NET0131  ;
  input \core_c_psq_CNTR_reg_DO_reg[6]/NET0131  ;
  input \core_c_psq_CNTR_reg_DO_reg[7]/NET0131  ;
  input \core_c_psq_CNTR_reg_DO_reg[8]/NET0131  ;
  input \core_c_psq_CNTR_reg_DO_reg[9]/NET0131  ;
  input \core_c_psq_CNTRval_reg/NET0131  ;
  input \core_c_psq_DMOVL_reg_DO_reg[0]/NET0131  ;
  input \core_c_psq_DMOVL_reg_DO_reg[1]/NET0131  ;
  input \core_c_psq_DMOVL_reg_DO_reg[2]/NET0131  ;
  input \core_c_psq_DMOVL_reg_DO_reg[3]/NET0131  ;
  input \core_c_psq_DRA_reg[0]/P0001  ;
  input \core_c_psq_DRA_reg[10]/P0001  ;
  input \core_c_psq_DRA_reg[11]/P0001  ;
  input \core_c_psq_DRA_reg[12]/P0001  ;
  input \core_c_psq_DRA_reg[13]/P0001  ;
  input \core_c_psq_DRA_reg[1]/P0001  ;
  input \core_c_psq_DRA_reg[2]/P0001  ;
  input \core_c_psq_DRA_reg[3]/P0001  ;
  input \core_c_psq_DRA_reg[4]/P0001  ;
  input \core_c_psq_DRA_reg[5]/P0001  ;
  input \core_c_psq_DRA_reg[6]/P0001  ;
  input \core_c_psq_DRA_reg[7]/P0001  ;
  input \core_c_psq_DRA_reg[8]/P0001  ;
  input \core_c_psq_DRA_reg[9]/P0001  ;
  input \core_c_psq_ECYC_reg/P0001  ;
  input \core_c_psq_EXA_reg[0]/P0001  ;
  input \core_c_psq_EXA_reg[10]/P0001  ;
  input \core_c_psq_EXA_reg[11]/P0001  ;
  input \core_c_psq_EXA_reg[12]/P0001  ;
  input \core_c_psq_EXA_reg[13]/P0001  ;
  input \core_c_psq_EXA_reg[1]/P0001  ;
  input \core_c_psq_EXA_reg[2]/P0001  ;
  input \core_c_psq_EXA_reg[3]/P0001  ;
  input \core_c_psq_EXA_reg[4]/P0001  ;
  input \core_c_psq_EXA_reg[5]/P0001  ;
  input \core_c_psq_EXA_reg[6]/P0001  ;
  input \core_c_psq_EXA_reg[7]/P0001  ;
  input \core_c_psq_EXA_reg[8]/P0001  ;
  input \core_c_psq_EXA_reg[9]/P0001  ;
  input \core_c_psq_Eqend_D_reg/P0001  ;
  input \core_c_psq_Eqend_Ed_reg/P0001  ;
  input \core_c_psq_ICNTL_reg_DO_reg[0]/NET0131  ;
  input \core_c_psq_ICNTL_reg_DO_reg[1]/NET0131  ;
  input \core_c_psq_ICNTL_reg_DO_reg[2]/NET0131  ;
  input \core_c_psq_ICNTL_reg_DO_reg[4]/NET0131  ;
  input \core_c_psq_IFA_reg[0]/P0001  ;
  input \core_c_psq_IFA_reg[10]/P0001  ;
  input \core_c_psq_IFA_reg[11]/P0001  ;
  input \core_c_psq_IFA_reg[12]/P0001  ;
  input \core_c_psq_IFA_reg[13]/P0001  ;
  input \core_c_psq_IFA_reg[1]/P0001  ;
  input \core_c_psq_IFA_reg[2]/P0001  ;
  input \core_c_psq_IFA_reg[3]/P0001  ;
  input \core_c_psq_IFA_reg[4]/P0001  ;
  input \core_c_psq_IFA_reg[5]/P0001  ;
  input \core_c_psq_IFA_reg[6]/P0001  ;
  input \core_c_psq_IFA_reg[7]/P0001  ;
  input \core_c_psq_IFA_reg[8]/P0001  ;
  input \core_c_psq_IFA_reg[9]/P0001  ;
  input \core_c_psq_IFC_reg[0]/NET0131  ;
  input \core_c_psq_IFC_reg[10]/NET0131  ;
  input \core_c_psq_IFC_reg[11]/NET0131  ;
  input \core_c_psq_IFC_reg[12]/NET0131  ;
  input \core_c_psq_IFC_reg[13]/NET0131  ;
  input \core_c_psq_IFC_reg[14]/NET0131  ;
  input \core_c_psq_IFC_reg[15]/NET0131  ;
  input \core_c_psq_IFC_reg[1]/NET0131  ;
  input \core_c_psq_IFC_reg[2]/NET0131  ;
  input \core_c_psq_IFC_reg[3]/NET0131  ;
  input \core_c_psq_IFC_reg[4]/NET0131  ;
  input \core_c_psq_IFC_reg[5]/NET0131  ;
  input \core_c_psq_IFC_reg[6]/NET0131  ;
  input \core_c_psq_IFC_reg[7]/NET0131  ;
  input \core_c_psq_IFC_reg[8]/NET0131  ;
  input \core_c_psq_IFC_reg[9]/NET0131  ;
  input \core_c_psq_IMASK_reg[0]/NET0131  ;
  input \core_c_psq_IMASK_reg[1]/NET0131  ;
  input \core_c_psq_IMASK_reg[2]/NET0131  ;
  input \core_c_psq_IMASK_reg[3]/NET0131  ;
  input \core_c_psq_IMASK_reg[4]/NET0131  ;
  input \core_c_psq_IMASK_reg[5]/NET0131  ;
  input \core_c_psq_IMASK_reg[6]/NET0131  ;
  input \core_c_psq_IMASK_reg[7]/NET0131  ;
  input \core_c_psq_IMASK_reg[8]/NET0131  ;
  input \core_c_psq_IMASK_reg[9]/NET0131  ;
  input \core_c_psq_INT_en_reg/NET0131  ;
  input \core_c_psq_Iact_E_reg[0]/NET0131  ;
  input \core_c_psq_Iact_E_reg[10]/NET0131  ;
  input \core_c_psq_Iact_E_reg[1]/NET0131  ;
  input \core_c_psq_Iact_E_reg[2]/NET0131  ;
  input \core_c_psq_Iact_E_reg[3]/NET0131  ;
  input \core_c_psq_Iact_E_reg[4]/NET0131  ;
  input \core_c_psq_Iact_E_reg[5]/NET0131  ;
  input \core_c_psq_Iact_E_reg[6]/NET0131  ;
  input \core_c_psq_Iact_E_reg[7]/NET0131  ;
  input \core_c_psq_Iact_E_reg[8]/NET0131  ;
  input \core_c_psq_Iact_E_reg[9]/NET0131  ;
  input \core_c_psq_Iflag_reg[0]/NET0131  ;
  input \core_c_psq_Iflag_reg[10]/NET0131  ;
  input \core_c_psq_Iflag_reg[11]/NET0131  ;
  input \core_c_psq_Iflag_reg[12]/NET0131  ;
  input \core_c_psq_Iflag_reg[1]/NET0131  ;
  input \core_c_psq_Iflag_reg[2]/NET0131  ;
  input \core_c_psq_Iflag_reg[3]/NET0131  ;
  input \core_c_psq_Iflag_reg[4]/NET0131  ;
  input \core_c_psq_Iflag_reg[5]/NET0131  ;
  input \core_c_psq_Iflag_reg[6]/NET0131  ;
  input \core_c_psq_Iflag_reg[7]/NET0131  ;
  input \core_c_psq_Iflag_reg[8]/NET0131  ;
  input \core_c_psq_Iflag_reg[9]/NET0131  ;
  input \core_c_psq_MGNT_reg/NET0131  ;
  input \core_c_psq_MREQ_reg/NET0131  ;
  input \core_c_psq_MSTAT_reg_DO_reg[0]/P0002  ;
  input \core_c_psq_MSTAT_reg_DO_reg[1]/NET0131  ;
  input \core_c_psq_MSTAT_reg_DO_reg[2]/NET0131  ;
  input \core_c_psq_MSTAT_reg_DO_reg[3]/NET0131  ;
  input \core_c_psq_MSTAT_reg_DO_reg[4]/NET0131  ;
  input \core_c_psq_MSTAT_reg_DO_reg[5]/NET0131  ;
  input \core_c_psq_MSTAT_reg_DO_reg[6]/NET0131  ;
  input \core_c_psq_PCS2or3_reg/NET0131  ;
  input \core_c_psq_PCS_reg[0]/NET0131  ;
  input \core_c_psq_PCS_reg[10]/NET0131  ;
  input \core_c_psq_PCS_reg[11]/NET0131  ;
  input \core_c_psq_PCS_reg[12]/NET0131  ;
  input \core_c_psq_PCS_reg[13]/NET0131  ;
  input \core_c_psq_PCS_reg[14]/NET0131  ;
  input \core_c_psq_PCS_reg[15]/NET0131  ;
  input \core_c_psq_PCS_reg[1]/NET0131  ;
  input \core_c_psq_PCS_reg[2]/NET0131  ;
  input \core_c_psq_PCS_reg[3]/NET0131  ;
  input \core_c_psq_PCS_reg[4]/NET0131  ;
  input \core_c_psq_PCS_reg[5]/NET0131  ;
  input \core_c_psq_PCS_reg[6]/NET0131  ;
  input \core_c_psq_PCS_reg[7]/NET0131  ;
  input \core_c_psq_PCS_reg[8]/NET0131  ;
  input \core_c_psq_PMOVL_regh_DO_reg[0]/NET0131  ;
  input \core_c_psq_PMOVL_regh_DO_reg[1]/NET0131  ;
  input \core_c_psq_PMOVL_regh_DO_reg[2]/NET0131  ;
  input \core_c_psq_PMOVL_regh_DO_reg[3]/NET0131  ;
  input \core_c_psq_PMOVL_regl_DO_reg[0]/NET0131  ;
  input \core_c_psq_PMOVL_regl_DO_reg[1]/NET0131  ;
  input \core_c_psq_PMOVL_regl_DO_reg[2]/NET0131  ;
  input \core_c_psq_PMOVL_regl_DO_reg[3]/NET0131  ;
  input \core_c_psq_SRST_reg/P0001  ;
  input \core_c_psq_SSTAT_reg[0]/NET0131  ;
  input \core_c_psq_SSTAT_reg[1]/NET0131  ;
  input \core_c_psq_SSTAT_reg[2]/NET0131  ;
  input \core_c_psq_SSTAT_reg[3]/NET0131  ;
  input \core_c_psq_SSTAT_reg[4]/NET0131  ;
  input \core_c_psq_SSTAT_reg[5]/NET0131  ;
  input \core_c_psq_SSTAT_reg[6]/NET0131  ;
  input \core_c_psq_SSTAT_reg[7]/NET0131  ;
  input \core_c_psq_TRAP_Eg_reg/NET0131  ;
  input \core_c_psq_TRAP_R_L_reg/NET0131  ;
  input \core_c_psq_T_IRQ0_s1_reg/P0001  ;
  input \core_c_psq_T_IRQ0p_reg/P0001  ;
  input \core_c_psq_T_IRQ1_s1_reg/P0001  ;
  input \core_c_psq_T_IRQ1p_reg/P0001  ;
  input \core_c_psq_T_IRQ2_s1_reg/P0001  ;
  input \core_c_psq_T_IRQ2p_reg/P0001  ;
  input \core_c_psq_T_IRQE0_reg/P0001  ;
  input \core_c_psq_T_IRQE0_s1_reg/P0001  ;
  input \core_c_psq_T_IRQE1_reg/P0001  ;
  input \core_c_psq_T_IRQE1_s1_reg/P0001  ;
  input \core_c_psq_T_IRQL0p_reg/P0001  ;
  input \core_c_psq_T_IRQL1p_reg/P0001  ;
  input \core_c_psq_T_PWRDN_reg/P0001  ;
  input \core_c_psq_T_PWRDN_s1_reg/P0001  ;
  input \core_c_psq_Taddr_Eb_reg[0]/P0001  ;
  input \core_c_psq_Taddr_Eb_reg[10]/P0001  ;
  input \core_c_psq_Taddr_Eb_reg[11]/P0001  ;
  input \core_c_psq_Taddr_Eb_reg[12]/P0001  ;
  input \core_c_psq_Taddr_Eb_reg[13]/P0001  ;
  input \core_c_psq_Taddr_Eb_reg[1]/P0001  ;
  input \core_c_psq_Taddr_Eb_reg[2]/P0001  ;
  input \core_c_psq_Taddr_Eb_reg[3]/P0001  ;
  input \core_c_psq_Taddr_Eb_reg[4]/P0001  ;
  input \core_c_psq_Taddr_Eb_reg[5]/P0001  ;
  input \core_c_psq_Taddr_Eb_reg[6]/P0001  ;
  input \core_c_psq_Taddr_Eb_reg[7]/P0001  ;
  input \core_c_psq_Taddr_Eb_reg[8]/P0001  ;
  input \core_c_psq_Taddr_Eb_reg[9]/P0001  ;
  input \core_c_psq_cntstk_cnts4x14_CNTcell_reg[0][0]/P0001  ;
  input \core_c_psq_cntstk_cnts4x14_CNTcell_reg[0][10]/P0001  ;
  input \core_c_psq_cntstk_cnts4x14_CNTcell_reg[0][11]/P0001  ;
  input \core_c_psq_cntstk_cnts4x14_CNTcell_reg[0][12]/P0001  ;
  input \core_c_psq_cntstk_cnts4x14_CNTcell_reg[0][13]/P0001  ;
  input \core_c_psq_cntstk_cnts4x14_CNTcell_reg[0][1]/P0001  ;
  input \core_c_psq_cntstk_cnts4x14_CNTcell_reg[0][2]/P0001  ;
  input \core_c_psq_cntstk_cnts4x14_CNTcell_reg[0][3]/P0001  ;
  input \core_c_psq_cntstk_cnts4x14_CNTcell_reg[0][4]/P0001  ;
  input \core_c_psq_cntstk_cnts4x14_CNTcell_reg[0][5]/P0001  ;
  input \core_c_psq_cntstk_cnts4x14_CNTcell_reg[0][6]/P0001  ;
  input \core_c_psq_cntstk_cnts4x14_CNTcell_reg[0][7]/P0001  ;
  input \core_c_psq_cntstk_cnts4x14_CNTcell_reg[0][8]/P0001  ;
  input \core_c_psq_cntstk_cnts4x14_CNTcell_reg[0][9]/P0001  ;
  input \core_c_psq_cntstk_cnts4x14_CNTcell_reg[1][0]/P0001  ;
  input \core_c_psq_cntstk_cnts4x14_CNTcell_reg[1][10]/P0001  ;
  input \core_c_psq_cntstk_cnts4x14_CNTcell_reg[1][11]/P0001  ;
  input \core_c_psq_cntstk_cnts4x14_CNTcell_reg[1][12]/P0001  ;
  input \core_c_psq_cntstk_cnts4x14_CNTcell_reg[1][13]/P0001  ;
  input \core_c_psq_cntstk_cnts4x14_CNTcell_reg[1][1]/P0001  ;
  input \core_c_psq_cntstk_cnts4x14_CNTcell_reg[1][2]/P0001  ;
  input \core_c_psq_cntstk_cnts4x14_CNTcell_reg[1][3]/P0001  ;
  input \core_c_psq_cntstk_cnts4x14_CNTcell_reg[1][4]/P0001  ;
  input \core_c_psq_cntstk_cnts4x14_CNTcell_reg[1][5]/P0001  ;
  input \core_c_psq_cntstk_cnts4x14_CNTcell_reg[1][6]/P0001  ;
  input \core_c_psq_cntstk_cnts4x14_CNTcell_reg[1][7]/P0001  ;
  input \core_c_psq_cntstk_cnts4x14_CNTcell_reg[1][8]/P0001  ;
  input \core_c_psq_cntstk_cnts4x14_CNTcell_reg[1][9]/P0001  ;
  input \core_c_psq_cntstk_cnts4x14_CNTcell_reg[2][0]/P0001  ;
  input \core_c_psq_cntstk_cnts4x14_CNTcell_reg[2][10]/P0001  ;
  input \core_c_psq_cntstk_cnts4x14_CNTcell_reg[2][11]/P0001  ;
  input \core_c_psq_cntstk_cnts4x14_CNTcell_reg[2][12]/P0001  ;
  input \core_c_psq_cntstk_cnts4x14_CNTcell_reg[2][13]/P0001  ;
  input \core_c_psq_cntstk_cnts4x14_CNTcell_reg[2][1]/P0001  ;
  input \core_c_psq_cntstk_cnts4x14_CNTcell_reg[2][2]/P0001  ;
  input \core_c_psq_cntstk_cnts4x14_CNTcell_reg[2][3]/P0001  ;
  input \core_c_psq_cntstk_cnts4x14_CNTcell_reg[2][4]/P0001  ;
  input \core_c_psq_cntstk_cnts4x14_CNTcell_reg[2][5]/P0001  ;
  input \core_c_psq_cntstk_cnts4x14_CNTcell_reg[2][6]/P0001  ;
  input \core_c_psq_cntstk_cnts4x14_CNTcell_reg[2][7]/P0001  ;
  input \core_c_psq_cntstk_cnts4x14_CNTcell_reg[2][8]/P0001  ;
  input \core_c_psq_cntstk_cnts4x14_CNTcell_reg[2][9]/P0001  ;
  input \core_c_psq_cntstk_cnts4x14_CNTcell_reg[3][0]/P0001  ;
  input \core_c_psq_cntstk_cnts4x14_CNTcell_reg[3][10]/P0001  ;
  input \core_c_psq_cntstk_cnts4x14_CNTcell_reg[3][11]/P0001  ;
  input \core_c_psq_cntstk_cnts4x14_CNTcell_reg[3][12]/P0001  ;
  input \core_c_psq_cntstk_cnts4x14_CNTcell_reg[3][13]/P0001  ;
  input \core_c_psq_cntstk_cnts4x14_CNTcell_reg[3][1]/P0001  ;
  input \core_c_psq_cntstk_cnts4x14_CNTcell_reg[3][2]/P0001  ;
  input \core_c_psq_cntstk_cnts4x14_CNTcell_reg[3][3]/P0001  ;
  input \core_c_psq_cntstk_cnts4x14_CNTcell_reg[3][4]/P0001  ;
  input \core_c_psq_cntstk_cnts4x14_CNTcell_reg[3][5]/P0001  ;
  input \core_c_psq_cntstk_cnts4x14_CNTcell_reg[3][6]/P0001  ;
  input \core_c_psq_cntstk_cnts4x14_CNTcell_reg[3][7]/P0001  ;
  input \core_c_psq_cntstk_cnts4x14_CNTcell_reg[3][8]/P0001  ;
  input \core_c_psq_cntstk_cnts4x14_CNTcell_reg[3][9]/P0001  ;
  input \core_c_psq_cntstk_ptr_reg[0]/NET0131  ;
  input \core_c_psq_cntstk_ptr_reg[1]/NET0131  ;
  input \core_c_psq_cntstk_ptr_reg[2]/NET0131  ;
  input \core_c_psq_irq0_de_IN_syn_reg/P0001  ;
  input \core_c_psq_irq0_de_OUT_reg/P0001  ;
  input \core_c_psq_irq1_de_IN_syn_reg/P0001  ;
  input \core_c_psq_irq1_de_OUT_reg/P0001  ;
  input \core_c_psq_irq2_de_IN_syn_reg/P0001  ;
  input \core_c_psq_irq2_de_OUT_reg/P0001  ;
  input \core_c_psq_irql0_de_IN_syn_reg/P0001  ;
  input \core_c_psq_irql0_de_OUT_reg/P0001  ;
  input \core_c_psq_irql1_de_IN_syn_reg/P0001  ;
  input \core_c_psq_irql1_de_OUT_reg/P0001  ;
  input \core_c_psq_lpstk_lps4x22_LPcell_reg[0][0]/P0001  ;
  input \core_c_psq_lpstk_lps4x22_LPcell_reg[0][10]/P0001  ;
  input \core_c_psq_lpstk_lps4x22_LPcell_reg[0][11]/P0001  ;
  input \core_c_psq_lpstk_lps4x22_LPcell_reg[0][12]/P0001  ;
  input \core_c_psq_lpstk_lps4x22_LPcell_reg[0][13]/P0001  ;
  input \core_c_psq_lpstk_lps4x22_LPcell_reg[0][14]/P0001  ;
  input \core_c_psq_lpstk_lps4x22_LPcell_reg[0][15]/P0001  ;
  input \core_c_psq_lpstk_lps4x22_LPcell_reg[0][16]/P0001  ;
  input \core_c_psq_lpstk_lps4x22_LPcell_reg[0][17]/P0001  ;
  input \core_c_psq_lpstk_lps4x22_LPcell_reg[0][18]/P0001  ;
  input \core_c_psq_lpstk_lps4x22_LPcell_reg[0][19]/P0001  ;
  input \core_c_psq_lpstk_lps4x22_LPcell_reg[0][1]/P0001  ;
  input \core_c_psq_lpstk_lps4x22_LPcell_reg[0][20]/P0001  ;
  input \core_c_psq_lpstk_lps4x22_LPcell_reg[0][21]/P0001  ;
  input \core_c_psq_lpstk_lps4x22_LPcell_reg[0][2]/P0001  ;
  input \core_c_psq_lpstk_lps4x22_LPcell_reg[0][3]/P0001  ;
  input \core_c_psq_lpstk_lps4x22_LPcell_reg[0][4]/P0001  ;
  input \core_c_psq_lpstk_lps4x22_LPcell_reg[0][5]/P0001  ;
  input \core_c_psq_lpstk_lps4x22_LPcell_reg[0][6]/P0001  ;
  input \core_c_psq_lpstk_lps4x22_LPcell_reg[0][7]/P0001  ;
  input \core_c_psq_lpstk_lps4x22_LPcell_reg[0][8]/P0001  ;
  input \core_c_psq_lpstk_lps4x22_LPcell_reg[0][9]/P0001  ;
  input \core_c_psq_lpstk_lps4x22_LPcell_reg[1][0]/P0001  ;
  input \core_c_psq_lpstk_lps4x22_LPcell_reg[1][10]/P0001  ;
  input \core_c_psq_lpstk_lps4x22_LPcell_reg[1][11]/P0001  ;
  input \core_c_psq_lpstk_lps4x22_LPcell_reg[1][12]/P0001  ;
  input \core_c_psq_lpstk_lps4x22_LPcell_reg[1][13]/P0001  ;
  input \core_c_psq_lpstk_lps4x22_LPcell_reg[1][14]/P0001  ;
  input \core_c_psq_lpstk_lps4x22_LPcell_reg[1][15]/P0001  ;
  input \core_c_psq_lpstk_lps4x22_LPcell_reg[1][16]/P0001  ;
  input \core_c_psq_lpstk_lps4x22_LPcell_reg[1][17]/P0001  ;
  input \core_c_psq_lpstk_lps4x22_LPcell_reg[1][18]/P0001  ;
  input \core_c_psq_lpstk_lps4x22_LPcell_reg[1][19]/P0001  ;
  input \core_c_psq_lpstk_lps4x22_LPcell_reg[1][1]/P0001  ;
  input \core_c_psq_lpstk_lps4x22_LPcell_reg[1][20]/P0001  ;
  input \core_c_psq_lpstk_lps4x22_LPcell_reg[1][21]/P0001  ;
  input \core_c_psq_lpstk_lps4x22_LPcell_reg[1][2]/P0001  ;
  input \core_c_psq_lpstk_lps4x22_LPcell_reg[1][3]/P0001  ;
  input \core_c_psq_lpstk_lps4x22_LPcell_reg[1][4]/P0001  ;
  input \core_c_psq_lpstk_lps4x22_LPcell_reg[1][5]/P0001  ;
  input \core_c_psq_lpstk_lps4x22_LPcell_reg[1][6]/P0001  ;
  input \core_c_psq_lpstk_lps4x22_LPcell_reg[1][7]/P0001  ;
  input \core_c_psq_lpstk_lps4x22_LPcell_reg[1][8]/P0001  ;
  input \core_c_psq_lpstk_lps4x22_LPcell_reg[1][9]/P0001  ;
  input \core_c_psq_lpstk_lps4x22_LPcell_reg[2][0]/P0001  ;
  input \core_c_psq_lpstk_lps4x22_LPcell_reg[2][10]/P0001  ;
  input \core_c_psq_lpstk_lps4x22_LPcell_reg[2][11]/P0001  ;
  input \core_c_psq_lpstk_lps4x22_LPcell_reg[2][12]/P0001  ;
  input \core_c_psq_lpstk_lps4x22_LPcell_reg[2][13]/P0001  ;
  input \core_c_psq_lpstk_lps4x22_LPcell_reg[2][14]/P0001  ;
  input \core_c_psq_lpstk_lps4x22_LPcell_reg[2][15]/P0001  ;
  input \core_c_psq_lpstk_lps4x22_LPcell_reg[2][16]/P0001  ;
  input \core_c_psq_lpstk_lps4x22_LPcell_reg[2][17]/P0001  ;
  input \core_c_psq_lpstk_lps4x22_LPcell_reg[2][18]/P0001  ;
  input \core_c_psq_lpstk_lps4x22_LPcell_reg[2][19]/P0001  ;
  input \core_c_psq_lpstk_lps4x22_LPcell_reg[2][1]/P0001  ;
  input \core_c_psq_lpstk_lps4x22_LPcell_reg[2][20]/P0001  ;
  input \core_c_psq_lpstk_lps4x22_LPcell_reg[2][21]/P0001  ;
  input \core_c_psq_lpstk_lps4x22_LPcell_reg[2][2]/P0001  ;
  input \core_c_psq_lpstk_lps4x22_LPcell_reg[2][3]/P0001  ;
  input \core_c_psq_lpstk_lps4x22_LPcell_reg[2][4]/P0001  ;
  input \core_c_psq_lpstk_lps4x22_LPcell_reg[2][5]/P0001  ;
  input \core_c_psq_lpstk_lps4x22_LPcell_reg[2][6]/P0001  ;
  input \core_c_psq_lpstk_lps4x22_LPcell_reg[2][7]/P0001  ;
  input \core_c_psq_lpstk_lps4x22_LPcell_reg[2][8]/P0001  ;
  input \core_c_psq_lpstk_lps4x22_LPcell_reg[2][9]/P0001  ;
  input \core_c_psq_lpstk_lps4x22_LPcell_reg[3][0]/P0001  ;
  input \core_c_psq_lpstk_lps4x22_LPcell_reg[3][10]/P0001  ;
  input \core_c_psq_lpstk_lps4x22_LPcell_reg[3][11]/P0001  ;
  input \core_c_psq_lpstk_lps4x22_LPcell_reg[3][12]/P0001  ;
  input \core_c_psq_lpstk_lps4x22_LPcell_reg[3][13]/P0001  ;
  input \core_c_psq_lpstk_lps4x22_LPcell_reg[3][14]/P0001  ;
  input \core_c_psq_lpstk_lps4x22_LPcell_reg[3][15]/P0001  ;
  input \core_c_psq_lpstk_lps4x22_LPcell_reg[3][16]/P0001  ;
  input \core_c_psq_lpstk_lps4x22_LPcell_reg[3][17]/P0001  ;
  input \core_c_psq_lpstk_lps4x22_LPcell_reg[3][18]/P0001  ;
  input \core_c_psq_lpstk_lps4x22_LPcell_reg[3][19]/P0001  ;
  input \core_c_psq_lpstk_lps4x22_LPcell_reg[3][1]/P0001  ;
  input \core_c_psq_lpstk_lps4x22_LPcell_reg[3][20]/P0001  ;
  input \core_c_psq_lpstk_lps4x22_LPcell_reg[3][21]/P0001  ;
  input \core_c_psq_lpstk_lps4x22_LPcell_reg[3][2]/P0001  ;
  input \core_c_psq_lpstk_lps4x22_LPcell_reg[3][3]/P0001  ;
  input \core_c_psq_lpstk_lps4x22_LPcell_reg[3][4]/P0001  ;
  input \core_c_psq_lpstk_lps4x22_LPcell_reg[3][5]/P0001  ;
  input \core_c_psq_lpstk_lps4x22_LPcell_reg[3][6]/P0001  ;
  input \core_c_psq_lpstk_lps4x22_LPcell_reg[3][7]/P0001  ;
  input \core_c_psq_lpstk_lps4x22_LPcell_reg[3][8]/P0001  ;
  input \core_c_psq_lpstk_lps4x22_LPcell_reg[3][9]/P0001  ;
  input \core_c_psq_lpstk_ptr_reg[0]/NET0131  ;
  input \core_c_psq_lpstk_ptr_reg[1]/NET0131  ;
  input \core_c_psq_lpstk_ptr_reg[2]/NET0131  ;
  input \core_c_psq_pcstk_cnts16x14_PCcell_reg[0][0]/P0001  ;
  input \core_c_psq_pcstk_cnts16x14_PCcell_reg[0][10]/P0001  ;
  input \core_c_psq_pcstk_cnts16x14_PCcell_reg[0][11]/P0001  ;
  input \core_c_psq_pcstk_cnts16x14_PCcell_reg[0][12]/P0001  ;
  input \core_c_psq_pcstk_cnts16x14_PCcell_reg[0][13]/P0001  ;
  input \core_c_psq_pcstk_cnts16x14_PCcell_reg[0][1]/P0001  ;
  input \core_c_psq_pcstk_cnts16x14_PCcell_reg[0][2]/P0001  ;
  input \core_c_psq_pcstk_cnts16x14_PCcell_reg[0][3]/P0001  ;
  input \core_c_psq_pcstk_cnts16x14_PCcell_reg[0][4]/P0001  ;
  input \core_c_psq_pcstk_cnts16x14_PCcell_reg[0][5]/P0001  ;
  input \core_c_psq_pcstk_cnts16x14_PCcell_reg[0][6]/P0001  ;
  input \core_c_psq_pcstk_cnts16x14_PCcell_reg[0][7]/P0001  ;
  input \core_c_psq_pcstk_cnts16x14_PCcell_reg[0][8]/P0001  ;
  input \core_c_psq_pcstk_cnts16x14_PCcell_reg[0][9]/P0001  ;
  input \core_c_psq_pcstk_cnts16x14_PCcell_reg[10][0]/P0001  ;
  input \core_c_psq_pcstk_cnts16x14_PCcell_reg[10][10]/P0001  ;
  input \core_c_psq_pcstk_cnts16x14_PCcell_reg[10][11]/P0001  ;
  input \core_c_psq_pcstk_cnts16x14_PCcell_reg[10][12]/P0001  ;
  input \core_c_psq_pcstk_cnts16x14_PCcell_reg[10][13]/P0001  ;
  input \core_c_psq_pcstk_cnts16x14_PCcell_reg[10][1]/P0001  ;
  input \core_c_psq_pcstk_cnts16x14_PCcell_reg[10][2]/P0001  ;
  input \core_c_psq_pcstk_cnts16x14_PCcell_reg[10][3]/P0001  ;
  input \core_c_psq_pcstk_cnts16x14_PCcell_reg[10][4]/P0001  ;
  input \core_c_psq_pcstk_cnts16x14_PCcell_reg[10][5]/P0001  ;
  input \core_c_psq_pcstk_cnts16x14_PCcell_reg[10][6]/P0001  ;
  input \core_c_psq_pcstk_cnts16x14_PCcell_reg[10][7]/P0001  ;
  input \core_c_psq_pcstk_cnts16x14_PCcell_reg[10][8]/P0001  ;
  input \core_c_psq_pcstk_cnts16x14_PCcell_reg[10][9]/P0001  ;
  input \core_c_psq_pcstk_cnts16x14_PCcell_reg[11][0]/P0001  ;
  input \core_c_psq_pcstk_cnts16x14_PCcell_reg[11][10]/P0001  ;
  input \core_c_psq_pcstk_cnts16x14_PCcell_reg[11][11]/P0001  ;
  input \core_c_psq_pcstk_cnts16x14_PCcell_reg[11][12]/P0001  ;
  input \core_c_psq_pcstk_cnts16x14_PCcell_reg[11][13]/P0001  ;
  input \core_c_psq_pcstk_cnts16x14_PCcell_reg[11][1]/P0001  ;
  input \core_c_psq_pcstk_cnts16x14_PCcell_reg[11][2]/P0001  ;
  input \core_c_psq_pcstk_cnts16x14_PCcell_reg[11][3]/P0001  ;
  input \core_c_psq_pcstk_cnts16x14_PCcell_reg[11][4]/P0001  ;
  input \core_c_psq_pcstk_cnts16x14_PCcell_reg[11][5]/P0001  ;
  input \core_c_psq_pcstk_cnts16x14_PCcell_reg[11][6]/P0001  ;
  input \core_c_psq_pcstk_cnts16x14_PCcell_reg[11][7]/P0001  ;
  input \core_c_psq_pcstk_cnts16x14_PCcell_reg[11][8]/P0001  ;
  input \core_c_psq_pcstk_cnts16x14_PCcell_reg[11][9]/P0001  ;
  input \core_c_psq_pcstk_cnts16x14_PCcell_reg[12][0]/P0001  ;
  input \core_c_psq_pcstk_cnts16x14_PCcell_reg[12][10]/P0001  ;
  input \core_c_psq_pcstk_cnts16x14_PCcell_reg[12][11]/P0001  ;
  input \core_c_psq_pcstk_cnts16x14_PCcell_reg[12][12]/P0001  ;
  input \core_c_psq_pcstk_cnts16x14_PCcell_reg[12][13]/P0001  ;
  input \core_c_psq_pcstk_cnts16x14_PCcell_reg[12][1]/P0001  ;
  input \core_c_psq_pcstk_cnts16x14_PCcell_reg[12][2]/P0001  ;
  input \core_c_psq_pcstk_cnts16x14_PCcell_reg[12][3]/P0001  ;
  input \core_c_psq_pcstk_cnts16x14_PCcell_reg[12][4]/P0001  ;
  input \core_c_psq_pcstk_cnts16x14_PCcell_reg[12][5]/P0001  ;
  input \core_c_psq_pcstk_cnts16x14_PCcell_reg[12][6]/P0001  ;
  input \core_c_psq_pcstk_cnts16x14_PCcell_reg[12][7]/P0001  ;
  input \core_c_psq_pcstk_cnts16x14_PCcell_reg[12][8]/P0001  ;
  input \core_c_psq_pcstk_cnts16x14_PCcell_reg[12][9]/P0001  ;
  input \core_c_psq_pcstk_cnts16x14_PCcell_reg[13][0]/P0001  ;
  input \core_c_psq_pcstk_cnts16x14_PCcell_reg[13][10]/P0001  ;
  input \core_c_psq_pcstk_cnts16x14_PCcell_reg[13][11]/P0001  ;
  input \core_c_psq_pcstk_cnts16x14_PCcell_reg[13][12]/P0001  ;
  input \core_c_psq_pcstk_cnts16x14_PCcell_reg[13][13]/P0001  ;
  input \core_c_psq_pcstk_cnts16x14_PCcell_reg[13][1]/P0001  ;
  input \core_c_psq_pcstk_cnts16x14_PCcell_reg[13][2]/P0001  ;
  input \core_c_psq_pcstk_cnts16x14_PCcell_reg[13][3]/P0001  ;
  input \core_c_psq_pcstk_cnts16x14_PCcell_reg[13][4]/P0001  ;
  input \core_c_psq_pcstk_cnts16x14_PCcell_reg[13][5]/P0001  ;
  input \core_c_psq_pcstk_cnts16x14_PCcell_reg[13][6]/P0001  ;
  input \core_c_psq_pcstk_cnts16x14_PCcell_reg[13][7]/P0001  ;
  input \core_c_psq_pcstk_cnts16x14_PCcell_reg[13][8]/P0001  ;
  input \core_c_psq_pcstk_cnts16x14_PCcell_reg[13][9]/P0001  ;
  input \core_c_psq_pcstk_cnts16x14_PCcell_reg[14][0]/P0001  ;
  input \core_c_psq_pcstk_cnts16x14_PCcell_reg[14][10]/P0001  ;
  input \core_c_psq_pcstk_cnts16x14_PCcell_reg[14][11]/P0001  ;
  input \core_c_psq_pcstk_cnts16x14_PCcell_reg[14][12]/P0001  ;
  input \core_c_psq_pcstk_cnts16x14_PCcell_reg[14][13]/P0001  ;
  input \core_c_psq_pcstk_cnts16x14_PCcell_reg[14][1]/P0001  ;
  input \core_c_psq_pcstk_cnts16x14_PCcell_reg[14][2]/P0001  ;
  input \core_c_psq_pcstk_cnts16x14_PCcell_reg[14][3]/P0001  ;
  input \core_c_psq_pcstk_cnts16x14_PCcell_reg[14][4]/P0001  ;
  input \core_c_psq_pcstk_cnts16x14_PCcell_reg[14][5]/P0001  ;
  input \core_c_psq_pcstk_cnts16x14_PCcell_reg[14][6]/P0001  ;
  input \core_c_psq_pcstk_cnts16x14_PCcell_reg[14][7]/P0001  ;
  input \core_c_psq_pcstk_cnts16x14_PCcell_reg[14][8]/P0001  ;
  input \core_c_psq_pcstk_cnts16x14_PCcell_reg[14][9]/P0001  ;
  input \core_c_psq_pcstk_cnts16x14_PCcell_reg[15][0]/P0001  ;
  input \core_c_psq_pcstk_cnts16x14_PCcell_reg[15][10]/P0001  ;
  input \core_c_psq_pcstk_cnts16x14_PCcell_reg[15][11]/P0001  ;
  input \core_c_psq_pcstk_cnts16x14_PCcell_reg[15][12]/P0001  ;
  input \core_c_psq_pcstk_cnts16x14_PCcell_reg[15][13]/P0001  ;
  input \core_c_psq_pcstk_cnts16x14_PCcell_reg[15][1]/P0001  ;
  input \core_c_psq_pcstk_cnts16x14_PCcell_reg[15][2]/P0001  ;
  input \core_c_psq_pcstk_cnts16x14_PCcell_reg[15][3]/P0001  ;
  input \core_c_psq_pcstk_cnts16x14_PCcell_reg[15][4]/P0001  ;
  input \core_c_psq_pcstk_cnts16x14_PCcell_reg[15][5]/P0001  ;
  input \core_c_psq_pcstk_cnts16x14_PCcell_reg[15][6]/P0001  ;
  input \core_c_psq_pcstk_cnts16x14_PCcell_reg[15][7]/P0001  ;
  input \core_c_psq_pcstk_cnts16x14_PCcell_reg[15][8]/P0001  ;
  input \core_c_psq_pcstk_cnts16x14_PCcell_reg[15][9]/P0001  ;
  input \core_c_psq_pcstk_cnts16x14_PCcell_reg[1][0]/P0001  ;
  input \core_c_psq_pcstk_cnts16x14_PCcell_reg[1][10]/P0001  ;
  input \core_c_psq_pcstk_cnts16x14_PCcell_reg[1][11]/P0001  ;
  input \core_c_psq_pcstk_cnts16x14_PCcell_reg[1][12]/P0001  ;
  input \core_c_psq_pcstk_cnts16x14_PCcell_reg[1][13]/P0001  ;
  input \core_c_psq_pcstk_cnts16x14_PCcell_reg[1][1]/P0001  ;
  input \core_c_psq_pcstk_cnts16x14_PCcell_reg[1][2]/P0001  ;
  input \core_c_psq_pcstk_cnts16x14_PCcell_reg[1][3]/P0001  ;
  input \core_c_psq_pcstk_cnts16x14_PCcell_reg[1][4]/P0001  ;
  input \core_c_psq_pcstk_cnts16x14_PCcell_reg[1][5]/P0001  ;
  input \core_c_psq_pcstk_cnts16x14_PCcell_reg[1][6]/P0001  ;
  input \core_c_psq_pcstk_cnts16x14_PCcell_reg[1][7]/P0001  ;
  input \core_c_psq_pcstk_cnts16x14_PCcell_reg[1][8]/P0001  ;
  input \core_c_psq_pcstk_cnts16x14_PCcell_reg[1][9]/P0001  ;
  input \core_c_psq_pcstk_cnts16x14_PCcell_reg[2][0]/P0001  ;
  input \core_c_psq_pcstk_cnts16x14_PCcell_reg[2][10]/P0001  ;
  input \core_c_psq_pcstk_cnts16x14_PCcell_reg[2][11]/P0001  ;
  input \core_c_psq_pcstk_cnts16x14_PCcell_reg[2][12]/P0001  ;
  input \core_c_psq_pcstk_cnts16x14_PCcell_reg[2][13]/P0001  ;
  input \core_c_psq_pcstk_cnts16x14_PCcell_reg[2][1]/P0001  ;
  input \core_c_psq_pcstk_cnts16x14_PCcell_reg[2][2]/P0001  ;
  input \core_c_psq_pcstk_cnts16x14_PCcell_reg[2][3]/P0001  ;
  input \core_c_psq_pcstk_cnts16x14_PCcell_reg[2][4]/P0001  ;
  input \core_c_psq_pcstk_cnts16x14_PCcell_reg[2][5]/P0001  ;
  input \core_c_psq_pcstk_cnts16x14_PCcell_reg[2][6]/P0001  ;
  input \core_c_psq_pcstk_cnts16x14_PCcell_reg[2][7]/P0001  ;
  input \core_c_psq_pcstk_cnts16x14_PCcell_reg[2][8]/P0001  ;
  input \core_c_psq_pcstk_cnts16x14_PCcell_reg[2][9]/P0001  ;
  input \core_c_psq_pcstk_cnts16x14_PCcell_reg[3][0]/P0001  ;
  input \core_c_psq_pcstk_cnts16x14_PCcell_reg[3][10]/P0001  ;
  input \core_c_psq_pcstk_cnts16x14_PCcell_reg[3][11]/P0001  ;
  input \core_c_psq_pcstk_cnts16x14_PCcell_reg[3][12]/P0001  ;
  input \core_c_psq_pcstk_cnts16x14_PCcell_reg[3][13]/P0001  ;
  input \core_c_psq_pcstk_cnts16x14_PCcell_reg[3][1]/P0001  ;
  input \core_c_psq_pcstk_cnts16x14_PCcell_reg[3][2]/P0001  ;
  input \core_c_psq_pcstk_cnts16x14_PCcell_reg[3][3]/P0001  ;
  input \core_c_psq_pcstk_cnts16x14_PCcell_reg[3][4]/P0001  ;
  input \core_c_psq_pcstk_cnts16x14_PCcell_reg[3][5]/P0001  ;
  input \core_c_psq_pcstk_cnts16x14_PCcell_reg[3][6]/P0001  ;
  input \core_c_psq_pcstk_cnts16x14_PCcell_reg[3][7]/P0001  ;
  input \core_c_psq_pcstk_cnts16x14_PCcell_reg[3][8]/P0001  ;
  input \core_c_psq_pcstk_cnts16x14_PCcell_reg[3][9]/P0001  ;
  input \core_c_psq_pcstk_cnts16x14_PCcell_reg[4][0]/P0001  ;
  input \core_c_psq_pcstk_cnts16x14_PCcell_reg[4][10]/P0001  ;
  input \core_c_psq_pcstk_cnts16x14_PCcell_reg[4][11]/P0001  ;
  input \core_c_psq_pcstk_cnts16x14_PCcell_reg[4][12]/P0001  ;
  input \core_c_psq_pcstk_cnts16x14_PCcell_reg[4][13]/P0001  ;
  input \core_c_psq_pcstk_cnts16x14_PCcell_reg[4][1]/P0001  ;
  input \core_c_psq_pcstk_cnts16x14_PCcell_reg[4][2]/P0001  ;
  input \core_c_psq_pcstk_cnts16x14_PCcell_reg[4][3]/P0001  ;
  input \core_c_psq_pcstk_cnts16x14_PCcell_reg[4][4]/P0001  ;
  input \core_c_psq_pcstk_cnts16x14_PCcell_reg[4][5]/P0001  ;
  input \core_c_psq_pcstk_cnts16x14_PCcell_reg[4][6]/P0001  ;
  input \core_c_psq_pcstk_cnts16x14_PCcell_reg[4][7]/P0001  ;
  input \core_c_psq_pcstk_cnts16x14_PCcell_reg[4][8]/P0001  ;
  input \core_c_psq_pcstk_cnts16x14_PCcell_reg[4][9]/P0001  ;
  input \core_c_psq_pcstk_cnts16x14_PCcell_reg[5][0]/P0001  ;
  input \core_c_psq_pcstk_cnts16x14_PCcell_reg[5][10]/P0001  ;
  input \core_c_psq_pcstk_cnts16x14_PCcell_reg[5][11]/P0001  ;
  input \core_c_psq_pcstk_cnts16x14_PCcell_reg[5][12]/P0001  ;
  input \core_c_psq_pcstk_cnts16x14_PCcell_reg[5][13]/P0001  ;
  input \core_c_psq_pcstk_cnts16x14_PCcell_reg[5][1]/P0001  ;
  input \core_c_psq_pcstk_cnts16x14_PCcell_reg[5][2]/P0001  ;
  input \core_c_psq_pcstk_cnts16x14_PCcell_reg[5][3]/P0001  ;
  input \core_c_psq_pcstk_cnts16x14_PCcell_reg[5][4]/P0001  ;
  input \core_c_psq_pcstk_cnts16x14_PCcell_reg[5][5]/P0001  ;
  input \core_c_psq_pcstk_cnts16x14_PCcell_reg[5][6]/P0001  ;
  input \core_c_psq_pcstk_cnts16x14_PCcell_reg[5][7]/P0001  ;
  input \core_c_psq_pcstk_cnts16x14_PCcell_reg[5][8]/P0001  ;
  input \core_c_psq_pcstk_cnts16x14_PCcell_reg[5][9]/P0001  ;
  input \core_c_psq_pcstk_cnts16x14_PCcell_reg[6][0]/P0001  ;
  input \core_c_psq_pcstk_cnts16x14_PCcell_reg[6][10]/P0001  ;
  input \core_c_psq_pcstk_cnts16x14_PCcell_reg[6][11]/P0001  ;
  input \core_c_psq_pcstk_cnts16x14_PCcell_reg[6][12]/P0001  ;
  input \core_c_psq_pcstk_cnts16x14_PCcell_reg[6][13]/P0001  ;
  input \core_c_psq_pcstk_cnts16x14_PCcell_reg[6][1]/P0001  ;
  input \core_c_psq_pcstk_cnts16x14_PCcell_reg[6][2]/P0001  ;
  input \core_c_psq_pcstk_cnts16x14_PCcell_reg[6][3]/P0001  ;
  input \core_c_psq_pcstk_cnts16x14_PCcell_reg[6][4]/P0001  ;
  input \core_c_psq_pcstk_cnts16x14_PCcell_reg[6][5]/P0001  ;
  input \core_c_psq_pcstk_cnts16x14_PCcell_reg[6][6]/P0001  ;
  input \core_c_psq_pcstk_cnts16x14_PCcell_reg[6][7]/P0001  ;
  input \core_c_psq_pcstk_cnts16x14_PCcell_reg[6][8]/P0001  ;
  input \core_c_psq_pcstk_cnts16x14_PCcell_reg[6][9]/P0001  ;
  input \core_c_psq_pcstk_cnts16x14_PCcell_reg[7][0]/P0001  ;
  input \core_c_psq_pcstk_cnts16x14_PCcell_reg[7][10]/P0001  ;
  input \core_c_psq_pcstk_cnts16x14_PCcell_reg[7][11]/P0001  ;
  input \core_c_psq_pcstk_cnts16x14_PCcell_reg[7][12]/P0001  ;
  input \core_c_psq_pcstk_cnts16x14_PCcell_reg[7][13]/P0001  ;
  input \core_c_psq_pcstk_cnts16x14_PCcell_reg[7][1]/P0001  ;
  input \core_c_psq_pcstk_cnts16x14_PCcell_reg[7][2]/P0001  ;
  input \core_c_psq_pcstk_cnts16x14_PCcell_reg[7][3]/P0001  ;
  input \core_c_psq_pcstk_cnts16x14_PCcell_reg[7][4]/P0001  ;
  input \core_c_psq_pcstk_cnts16x14_PCcell_reg[7][5]/P0001  ;
  input \core_c_psq_pcstk_cnts16x14_PCcell_reg[7][6]/P0001  ;
  input \core_c_psq_pcstk_cnts16x14_PCcell_reg[7][7]/P0001  ;
  input \core_c_psq_pcstk_cnts16x14_PCcell_reg[7][8]/P0001  ;
  input \core_c_psq_pcstk_cnts16x14_PCcell_reg[7][9]/P0001  ;
  input \core_c_psq_pcstk_cnts16x14_PCcell_reg[8][0]/P0001  ;
  input \core_c_psq_pcstk_cnts16x14_PCcell_reg[8][10]/P0001  ;
  input \core_c_psq_pcstk_cnts16x14_PCcell_reg[8][11]/P0001  ;
  input \core_c_psq_pcstk_cnts16x14_PCcell_reg[8][12]/P0001  ;
  input \core_c_psq_pcstk_cnts16x14_PCcell_reg[8][13]/P0001  ;
  input \core_c_psq_pcstk_cnts16x14_PCcell_reg[8][1]/P0001  ;
  input \core_c_psq_pcstk_cnts16x14_PCcell_reg[8][2]/P0001  ;
  input \core_c_psq_pcstk_cnts16x14_PCcell_reg[8][3]/P0001  ;
  input \core_c_psq_pcstk_cnts16x14_PCcell_reg[8][4]/P0001  ;
  input \core_c_psq_pcstk_cnts16x14_PCcell_reg[8][5]/P0001  ;
  input \core_c_psq_pcstk_cnts16x14_PCcell_reg[8][6]/P0001  ;
  input \core_c_psq_pcstk_cnts16x14_PCcell_reg[8][7]/P0001  ;
  input \core_c_psq_pcstk_cnts16x14_PCcell_reg[8][8]/P0001  ;
  input \core_c_psq_pcstk_cnts16x14_PCcell_reg[8][9]/P0001  ;
  input \core_c_psq_pcstk_cnts16x14_PCcell_reg[9][0]/P0001  ;
  input \core_c_psq_pcstk_cnts16x14_PCcell_reg[9][10]/P0001  ;
  input \core_c_psq_pcstk_cnts16x14_PCcell_reg[9][11]/P0001  ;
  input \core_c_psq_pcstk_cnts16x14_PCcell_reg[9][12]/P0001  ;
  input \core_c_psq_pcstk_cnts16x14_PCcell_reg[9][13]/P0001  ;
  input \core_c_psq_pcstk_cnts16x14_PCcell_reg[9][1]/P0001  ;
  input \core_c_psq_pcstk_cnts16x14_PCcell_reg[9][2]/P0001  ;
  input \core_c_psq_pcstk_cnts16x14_PCcell_reg[9][3]/P0001  ;
  input \core_c_psq_pcstk_cnts16x14_PCcell_reg[9][4]/P0001  ;
  input \core_c_psq_pcstk_cnts16x14_PCcell_reg[9][5]/P0001  ;
  input \core_c_psq_pcstk_cnts16x14_PCcell_reg[9][6]/P0001  ;
  input \core_c_psq_pcstk_cnts16x14_PCcell_reg[9][7]/P0001  ;
  input \core_c_psq_pcstk_cnts16x14_PCcell_reg[9][8]/P0001  ;
  input \core_c_psq_pcstk_cnts16x14_PCcell_reg[9][9]/P0001  ;
  input \core_c_psq_pcstk_ptr_reg[0]/NET0131  ;
  input \core_c_psq_pcstk_ptr_reg[1]/NET0131  ;
  input \core_c_psq_pcstk_ptr_reg[2]/NET0131  ;
  input \core_c_psq_pcstk_ptr_reg[3]/NET0131  ;
  input \core_c_psq_pcstk_ptr_reg[4]/NET0131  ;
  input \core_c_psq_ststk_ptr_reg[0]/NET0131  ;
  input \core_c_psq_ststk_ptr_reg[1]/NET0131  ;
  input \core_c_psq_ststk_ptr_reg[2]/NET0131  ;
  input \core_c_psq_ststk_sts7x23_STcell_reg[0][0]/P0001  ;
  input \core_c_psq_ststk_sts7x23_STcell_reg[0][10]/P0001  ;
  input \core_c_psq_ststk_sts7x23_STcell_reg[0][11]/P0001  ;
  input \core_c_psq_ststk_sts7x23_STcell_reg[0][12]/P0001  ;
  input \core_c_psq_ststk_sts7x23_STcell_reg[0][13]/P0001  ;
  input \core_c_psq_ststk_sts7x23_STcell_reg[0][14]/P0001  ;
  input \core_c_psq_ststk_sts7x23_STcell_reg[0][15]/P0001  ;
  input \core_c_psq_ststk_sts7x23_STcell_reg[0][16]/P0001  ;
  input \core_c_psq_ststk_sts7x23_STcell_reg[0][17]/P0001  ;
  input \core_c_psq_ststk_sts7x23_STcell_reg[0][18]/P0001  ;
  input \core_c_psq_ststk_sts7x23_STcell_reg[0][19]/P0001  ;
  input \core_c_psq_ststk_sts7x23_STcell_reg[0][1]/P0001  ;
  input \core_c_psq_ststk_sts7x23_STcell_reg[0][20]/P0001  ;
  input \core_c_psq_ststk_sts7x23_STcell_reg[0][21]/P0001  ;
  input \core_c_psq_ststk_sts7x23_STcell_reg[0][22]/P0001  ;
  input \core_c_psq_ststk_sts7x23_STcell_reg[0][23]/P0001  ;
  input \core_c_psq_ststk_sts7x23_STcell_reg[0][24]/P0001  ;
  input \core_c_psq_ststk_sts7x23_STcell_reg[0][2]/P0001  ;
  input \core_c_psq_ststk_sts7x23_STcell_reg[0][3]/P0001  ;
  input \core_c_psq_ststk_sts7x23_STcell_reg[0][4]/P0001  ;
  input \core_c_psq_ststk_sts7x23_STcell_reg[0][5]/P0001  ;
  input \core_c_psq_ststk_sts7x23_STcell_reg[0][6]/P0001  ;
  input \core_c_psq_ststk_sts7x23_STcell_reg[0][7]/P0001  ;
  input \core_c_psq_ststk_sts7x23_STcell_reg[0][8]/P0001  ;
  input \core_c_psq_ststk_sts7x23_STcell_reg[0][9]/P0001  ;
  input \core_c_psq_ststk_sts7x23_STcell_reg[1][0]/P0001  ;
  input \core_c_psq_ststk_sts7x23_STcell_reg[1][10]/P0001  ;
  input \core_c_psq_ststk_sts7x23_STcell_reg[1][11]/P0001  ;
  input \core_c_psq_ststk_sts7x23_STcell_reg[1][12]/P0001  ;
  input \core_c_psq_ststk_sts7x23_STcell_reg[1][13]/P0001  ;
  input \core_c_psq_ststk_sts7x23_STcell_reg[1][14]/P0001  ;
  input \core_c_psq_ststk_sts7x23_STcell_reg[1][15]/P0001  ;
  input \core_c_psq_ststk_sts7x23_STcell_reg[1][16]/P0001  ;
  input \core_c_psq_ststk_sts7x23_STcell_reg[1][17]/P0001  ;
  input \core_c_psq_ststk_sts7x23_STcell_reg[1][18]/P0001  ;
  input \core_c_psq_ststk_sts7x23_STcell_reg[1][19]/P0001  ;
  input \core_c_psq_ststk_sts7x23_STcell_reg[1][1]/P0001  ;
  input \core_c_psq_ststk_sts7x23_STcell_reg[1][20]/P0001  ;
  input \core_c_psq_ststk_sts7x23_STcell_reg[1][21]/P0001  ;
  input \core_c_psq_ststk_sts7x23_STcell_reg[1][22]/P0001  ;
  input \core_c_psq_ststk_sts7x23_STcell_reg[1][23]/P0001  ;
  input \core_c_psq_ststk_sts7x23_STcell_reg[1][24]/P0001  ;
  input \core_c_psq_ststk_sts7x23_STcell_reg[1][2]/P0001  ;
  input \core_c_psq_ststk_sts7x23_STcell_reg[1][3]/P0001  ;
  input \core_c_psq_ststk_sts7x23_STcell_reg[1][4]/P0001  ;
  input \core_c_psq_ststk_sts7x23_STcell_reg[1][5]/P0001  ;
  input \core_c_psq_ststk_sts7x23_STcell_reg[1][6]/P0001  ;
  input \core_c_psq_ststk_sts7x23_STcell_reg[1][7]/P0001  ;
  input \core_c_psq_ststk_sts7x23_STcell_reg[1][8]/P0001  ;
  input \core_c_psq_ststk_sts7x23_STcell_reg[1][9]/P0001  ;
  input \core_c_psq_ststk_sts7x23_STcell_reg[2][0]/P0001  ;
  input \core_c_psq_ststk_sts7x23_STcell_reg[2][10]/P0001  ;
  input \core_c_psq_ststk_sts7x23_STcell_reg[2][11]/P0001  ;
  input \core_c_psq_ststk_sts7x23_STcell_reg[2][12]/P0001  ;
  input \core_c_psq_ststk_sts7x23_STcell_reg[2][13]/P0001  ;
  input \core_c_psq_ststk_sts7x23_STcell_reg[2][14]/P0001  ;
  input \core_c_psq_ststk_sts7x23_STcell_reg[2][15]/P0001  ;
  input \core_c_psq_ststk_sts7x23_STcell_reg[2][16]/P0001  ;
  input \core_c_psq_ststk_sts7x23_STcell_reg[2][17]/P0001  ;
  input \core_c_psq_ststk_sts7x23_STcell_reg[2][18]/P0001  ;
  input \core_c_psq_ststk_sts7x23_STcell_reg[2][19]/P0001  ;
  input \core_c_psq_ststk_sts7x23_STcell_reg[2][1]/P0001  ;
  input \core_c_psq_ststk_sts7x23_STcell_reg[2][20]/P0001  ;
  input \core_c_psq_ststk_sts7x23_STcell_reg[2][21]/P0001  ;
  input \core_c_psq_ststk_sts7x23_STcell_reg[2][22]/P0001  ;
  input \core_c_psq_ststk_sts7x23_STcell_reg[2][23]/P0001  ;
  input \core_c_psq_ststk_sts7x23_STcell_reg[2][24]/P0001  ;
  input \core_c_psq_ststk_sts7x23_STcell_reg[2][2]/P0001  ;
  input \core_c_psq_ststk_sts7x23_STcell_reg[2][3]/P0001  ;
  input \core_c_psq_ststk_sts7x23_STcell_reg[2][4]/P0001  ;
  input \core_c_psq_ststk_sts7x23_STcell_reg[2][5]/P0001  ;
  input \core_c_psq_ststk_sts7x23_STcell_reg[2][6]/P0001  ;
  input \core_c_psq_ststk_sts7x23_STcell_reg[2][7]/P0001  ;
  input \core_c_psq_ststk_sts7x23_STcell_reg[2][8]/P0001  ;
  input \core_c_psq_ststk_sts7x23_STcell_reg[2][9]/P0001  ;
  input \core_c_psq_ststk_sts7x23_STcell_reg[3][0]/P0001  ;
  input \core_c_psq_ststk_sts7x23_STcell_reg[3][10]/P0001  ;
  input \core_c_psq_ststk_sts7x23_STcell_reg[3][11]/P0001  ;
  input \core_c_psq_ststk_sts7x23_STcell_reg[3][12]/P0001  ;
  input \core_c_psq_ststk_sts7x23_STcell_reg[3][13]/P0001  ;
  input \core_c_psq_ststk_sts7x23_STcell_reg[3][14]/P0001  ;
  input \core_c_psq_ststk_sts7x23_STcell_reg[3][15]/P0001  ;
  input \core_c_psq_ststk_sts7x23_STcell_reg[3][16]/P0001  ;
  input \core_c_psq_ststk_sts7x23_STcell_reg[3][17]/P0001  ;
  input \core_c_psq_ststk_sts7x23_STcell_reg[3][18]/P0001  ;
  input \core_c_psq_ststk_sts7x23_STcell_reg[3][19]/P0001  ;
  input \core_c_psq_ststk_sts7x23_STcell_reg[3][1]/P0001  ;
  input \core_c_psq_ststk_sts7x23_STcell_reg[3][20]/P0001  ;
  input \core_c_psq_ststk_sts7x23_STcell_reg[3][21]/P0001  ;
  input \core_c_psq_ststk_sts7x23_STcell_reg[3][22]/P0001  ;
  input \core_c_psq_ststk_sts7x23_STcell_reg[3][23]/P0001  ;
  input \core_c_psq_ststk_sts7x23_STcell_reg[3][24]/P0001  ;
  input \core_c_psq_ststk_sts7x23_STcell_reg[3][2]/P0001  ;
  input \core_c_psq_ststk_sts7x23_STcell_reg[3][3]/P0001  ;
  input \core_c_psq_ststk_sts7x23_STcell_reg[3][4]/P0001  ;
  input \core_c_psq_ststk_sts7x23_STcell_reg[3][5]/P0001  ;
  input \core_c_psq_ststk_sts7x23_STcell_reg[3][6]/P0001  ;
  input \core_c_psq_ststk_sts7x23_STcell_reg[3][7]/P0001  ;
  input \core_c_psq_ststk_sts7x23_STcell_reg[3][8]/P0001  ;
  input \core_c_psq_ststk_sts7x23_STcell_reg[3][9]/P0001  ;
  input \core_c_psq_ststk_sts7x23_STcell_reg[4][0]/P0001  ;
  input \core_c_psq_ststk_sts7x23_STcell_reg[4][10]/P0001  ;
  input \core_c_psq_ststk_sts7x23_STcell_reg[4][11]/P0001  ;
  input \core_c_psq_ststk_sts7x23_STcell_reg[4][12]/P0001  ;
  input \core_c_psq_ststk_sts7x23_STcell_reg[4][13]/P0001  ;
  input \core_c_psq_ststk_sts7x23_STcell_reg[4][14]/P0001  ;
  input \core_c_psq_ststk_sts7x23_STcell_reg[4][15]/P0001  ;
  input \core_c_psq_ststk_sts7x23_STcell_reg[4][16]/P0001  ;
  input \core_c_psq_ststk_sts7x23_STcell_reg[4][17]/P0001  ;
  input \core_c_psq_ststk_sts7x23_STcell_reg[4][18]/P0001  ;
  input \core_c_psq_ststk_sts7x23_STcell_reg[4][19]/P0001  ;
  input \core_c_psq_ststk_sts7x23_STcell_reg[4][1]/P0001  ;
  input \core_c_psq_ststk_sts7x23_STcell_reg[4][20]/P0001  ;
  input \core_c_psq_ststk_sts7x23_STcell_reg[4][21]/P0001  ;
  input \core_c_psq_ststk_sts7x23_STcell_reg[4][22]/P0001  ;
  input \core_c_psq_ststk_sts7x23_STcell_reg[4][23]/P0001  ;
  input \core_c_psq_ststk_sts7x23_STcell_reg[4][24]/P0001  ;
  input \core_c_psq_ststk_sts7x23_STcell_reg[4][2]/P0001  ;
  input \core_c_psq_ststk_sts7x23_STcell_reg[4][3]/P0001  ;
  input \core_c_psq_ststk_sts7x23_STcell_reg[4][4]/P0001  ;
  input \core_c_psq_ststk_sts7x23_STcell_reg[4][5]/P0001  ;
  input \core_c_psq_ststk_sts7x23_STcell_reg[4][6]/P0001  ;
  input \core_c_psq_ststk_sts7x23_STcell_reg[4][7]/P0001  ;
  input \core_c_psq_ststk_sts7x23_STcell_reg[4][8]/P0001  ;
  input \core_c_psq_ststk_sts7x23_STcell_reg[4][9]/P0001  ;
  input \core_c_psq_ststk_sts7x23_STcell_reg[5][0]/P0001  ;
  input \core_c_psq_ststk_sts7x23_STcell_reg[5][10]/P0001  ;
  input \core_c_psq_ststk_sts7x23_STcell_reg[5][11]/P0001  ;
  input \core_c_psq_ststk_sts7x23_STcell_reg[5][12]/P0001  ;
  input \core_c_psq_ststk_sts7x23_STcell_reg[5][13]/P0001  ;
  input \core_c_psq_ststk_sts7x23_STcell_reg[5][14]/P0001  ;
  input \core_c_psq_ststk_sts7x23_STcell_reg[5][15]/P0001  ;
  input \core_c_psq_ststk_sts7x23_STcell_reg[5][16]/P0001  ;
  input \core_c_psq_ststk_sts7x23_STcell_reg[5][17]/P0001  ;
  input \core_c_psq_ststk_sts7x23_STcell_reg[5][18]/P0001  ;
  input \core_c_psq_ststk_sts7x23_STcell_reg[5][19]/P0001  ;
  input \core_c_psq_ststk_sts7x23_STcell_reg[5][1]/P0001  ;
  input \core_c_psq_ststk_sts7x23_STcell_reg[5][20]/P0001  ;
  input \core_c_psq_ststk_sts7x23_STcell_reg[5][21]/P0001  ;
  input \core_c_psq_ststk_sts7x23_STcell_reg[5][22]/P0001  ;
  input \core_c_psq_ststk_sts7x23_STcell_reg[5][23]/P0001  ;
  input \core_c_psq_ststk_sts7x23_STcell_reg[5][24]/P0001  ;
  input \core_c_psq_ststk_sts7x23_STcell_reg[5][2]/P0001  ;
  input \core_c_psq_ststk_sts7x23_STcell_reg[5][3]/P0001  ;
  input \core_c_psq_ststk_sts7x23_STcell_reg[5][4]/P0001  ;
  input \core_c_psq_ststk_sts7x23_STcell_reg[5][5]/P0001  ;
  input \core_c_psq_ststk_sts7x23_STcell_reg[5][6]/P0001  ;
  input \core_c_psq_ststk_sts7x23_STcell_reg[5][7]/P0001  ;
  input \core_c_psq_ststk_sts7x23_STcell_reg[5][8]/P0001  ;
  input \core_c_psq_ststk_sts7x23_STcell_reg[5][9]/P0001  ;
  input \core_c_psq_ststk_sts7x23_STcell_reg[6][0]/P0001  ;
  input \core_c_psq_ststk_sts7x23_STcell_reg[6][10]/P0001  ;
  input \core_c_psq_ststk_sts7x23_STcell_reg[6][11]/P0001  ;
  input \core_c_psq_ststk_sts7x23_STcell_reg[6][12]/P0001  ;
  input \core_c_psq_ststk_sts7x23_STcell_reg[6][13]/P0001  ;
  input \core_c_psq_ststk_sts7x23_STcell_reg[6][14]/P0001  ;
  input \core_c_psq_ststk_sts7x23_STcell_reg[6][15]/P0001  ;
  input \core_c_psq_ststk_sts7x23_STcell_reg[6][16]/P0001  ;
  input \core_c_psq_ststk_sts7x23_STcell_reg[6][17]/P0001  ;
  input \core_c_psq_ststk_sts7x23_STcell_reg[6][18]/P0001  ;
  input \core_c_psq_ststk_sts7x23_STcell_reg[6][19]/P0001  ;
  input \core_c_psq_ststk_sts7x23_STcell_reg[6][1]/P0001  ;
  input \core_c_psq_ststk_sts7x23_STcell_reg[6][20]/P0001  ;
  input \core_c_psq_ststk_sts7x23_STcell_reg[6][21]/P0001  ;
  input \core_c_psq_ststk_sts7x23_STcell_reg[6][22]/P0001  ;
  input \core_c_psq_ststk_sts7x23_STcell_reg[6][23]/P0001  ;
  input \core_c_psq_ststk_sts7x23_STcell_reg[6][24]/P0001  ;
  input \core_c_psq_ststk_sts7x23_STcell_reg[6][2]/P0001  ;
  input \core_c_psq_ststk_sts7x23_STcell_reg[6][3]/P0001  ;
  input \core_c_psq_ststk_sts7x23_STcell_reg[6][4]/P0001  ;
  input \core_c_psq_ststk_sts7x23_STcell_reg[6][5]/P0001  ;
  input \core_c_psq_ststk_sts7x23_STcell_reg[6][6]/P0001  ;
  input \core_c_psq_ststk_sts7x23_STcell_reg[6][7]/P0001  ;
  input \core_c_psq_ststk_sts7x23_STcell_reg[6][8]/P0001  ;
  input \core_c_psq_ststk_sts7x23_STcell_reg[6][9]/P0001  ;
  input \core_dag_ilm1reg_DMA_pi_DO_reg[0]/NET0131  ;
  input \core_dag_ilm1reg_DMA_pi_DO_reg[10]/NET0131  ;
  input \core_dag_ilm1reg_DMA_pi_DO_reg[11]/NET0131  ;
  input \core_dag_ilm1reg_DMA_pi_DO_reg[12]/NET0131  ;
  input \core_dag_ilm1reg_DMA_pi_DO_reg[13]/NET0131  ;
  input \core_dag_ilm1reg_DMA_pi_DO_reg[1]/NET0131  ;
  input \core_dag_ilm1reg_DMA_pi_DO_reg[2]/NET0131  ;
  input \core_dag_ilm1reg_DMA_pi_DO_reg[3]/NET0131  ;
  input \core_dag_ilm1reg_DMA_pi_DO_reg[4]/NET0131  ;
  input \core_dag_ilm1reg_DMA_pi_DO_reg[5]/NET0131  ;
  input \core_dag_ilm1reg_DMA_pi_DO_reg[6]/NET0131  ;
  input \core_dag_ilm1reg_DMA_pi_DO_reg[7]/NET0131  ;
  input \core_dag_ilm1reg_DMA_pi_DO_reg[8]/NET0131  ;
  input \core_dag_ilm1reg_DMA_pi_DO_reg[9]/NET0131  ;
  input \core_dag_ilm1reg_I0_we_DO_reg[0]/NET0131  ;
  input \core_dag_ilm1reg_I0_we_DO_reg[10]/NET0131  ;
  input \core_dag_ilm1reg_I0_we_DO_reg[11]/NET0131  ;
  input \core_dag_ilm1reg_I0_we_DO_reg[12]/NET0131  ;
  input \core_dag_ilm1reg_I0_we_DO_reg[13]/NET0131  ;
  input \core_dag_ilm1reg_I0_we_DO_reg[1]/NET0131  ;
  input \core_dag_ilm1reg_I0_we_DO_reg[2]/NET0131  ;
  input \core_dag_ilm1reg_I0_we_DO_reg[3]/NET0131  ;
  input \core_dag_ilm1reg_I0_we_DO_reg[4]/NET0131  ;
  input \core_dag_ilm1reg_I0_we_DO_reg[5]/NET0131  ;
  input \core_dag_ilm1reg_I0_we_DO_reg[6]/NET0131  ;
  input \core_dag_ilm1reg_I0_we_DO_reg[7]/NET0131  ;
  input \core_dag_ilm1reg_I0_we_DO_reg[8]/NET0131  ;
  input \core_dag_ilm1reg_I0_we_DO_reg[9]/NET0131  ;
  input \core_dag_ilm1reg_I1_we_DO_reg[0]/NET0131  ;
  input \core_dag_ilm1reg_I1_we_DO_reg[10]/NET0131  ;
  input \core_dag_ilm1reg_I1_we_DO_reg[11]/NET0131  ;
  input \core_dag_ilm1reg_I1_we_DO_reg[12]/NET0131  ;
  input \core_dag_ilm1reg_I1_we_DO_reg[13]/NET0131  ;
  input \core_dag_ilm1reg_I1_we_DO_reg[1]/NET0131  ;
  input \core_dag_ilm1reg_I1_we_DO_reg[2]/NET0131  ;
  input \core_dag_ilm1reg_I1_we_DO_reg[3]/NET0131  ;
  input \core_dag_ilm1reg_I1_we_DO_reg[4]/NET0131  ;
  input \core_dag_ilm1reg_I1_we_DO_reg[5]/NET0131  ;
  input \core_dag_ilm1reg_I1_we_DO_reg[6]/NET0131  ;
  input \core_dag_ilm1reg_I1_we_DO_reg[7]/NET0131  ;
  input \core_dag_ilm1reg_I1_we_DO_reg[8]/NET0131  ;
  input \core_dag_ilm1reg_I1_we_DO_reg[9]/NET0131  ;
  input \core_dag_ilm1reg_I2_we_DO_reg[0]/NET0131  ;
  input \core_dag_ilm1reg_I2_we_DO_reg[10]/NET0131  ;
  input \core_dag_ilm1reg_I2_we_DO_reg[11]/NET0131  ;
  input \core_dag_ilm1reg_I2_we_DO_reg[12]/NET0131  ;
  input \core_dag_ilm1reg_I2_we_DO_reg[13]/NET0131  ;
  input \core_dag_ilm1reg_I2_we_DO_reg[1]/NET0131  ;
  input \core_dag_ilm1reg_I2_we_DO_reg[2]/NET0131  ;
  input \core_dag_ilm1reg_I2_we_DO_reg[3]/NET0131  ;
  input \core_dag_ilm1reg_I2_we_DO_reg[4]/NET0131  ;
  input \core_dag_ilm1reg_I2_we_DO_reg[5]/NET0131  ;
  input \core_dag_ilm1reg_I2_we_DO_reg[6]/NET0131  ;
  input \core_dag_ilm1reg_I2_we_DO_reg[7]/NET0131  ;
  input \core_dag_ilm1reg_I2_we_DO_reg[8]/NET0131  ;
  input \core_dag_ilm1reg_I2_we_DO_reg[9]/NET0131  ;
  input \core_dag_ilm1reg_I3_we_DO_reg[0]/NET0131  ;
  input \core_dag_ilm1reg_I3_we_DO_reg[10]/NET0131  ;
  input \core_dag_ilm1reg_I3_we_DO_reg[11]/NET0131  ;
  input \core_dag_ilm1reg_I3_we_DO_reg[12]/NET0131  ;
  input \core_dag_ilm1reg_I3_we_DO_reg[13]/NET0131  ;
  input \core_dag_ilm1reg_I3_we_DO_reg[1]/NET0131  ;
  input \core_dag_ilm1reg_I3_we_DO_reg[2]/NET0131  ;
  input \core_dag_ilm1reg_I3_we_DO_reg[3]/NET0131  ;
  input \core_dag_ilm1reg_I3_we_DO_reg[4]/NET0131  ;
  input \core_dag_ilm1reg_I3_we_DO_reg[5]/NET0131  ;
  input \core_dag_ilm1reg_I3_we_DO_reg[6]/NET0131  ;
  input \core_dag_ilm1reg_I3_we_DO_reg[7]/NET0131  ;
  input \core_dag_ilm1reg_I3_we_DO_reg[8]/NET0131  ;
  input \core_dag_ilm1reg_I3_we_DO_reg[9]/NET0131  ;
  input \core_dag_ilm1reg_I_reg[0]/NET0131  ;
  input \core_dag_ilm1reg_I_reg[10]/NET0131  ;
  input \core_dag_ilm1reg_I_reg[11]/NET0131  ;
  input \core_dag_ilm1reg_I_reg[12]/NET0131  ;
  input \core_dag_ilm1reg_I_reg[13]/NET0131  ;
  input \core_dag_ilm1reg_I_reg[1]/NET0131  ;
  input \core_dag_ilm1reg_I_reg[2]/NET0131  ;
  input \core_dag_ilm1reg_I_reg[3]/NET0131  ;
  input \core_dag_ilm1reg_I_reg[4]/NET0131  ;
  input \core_dag_ilm1reg_I_reg[5]/NET0131  ;
  input \core_dag_ilm1reg_I_reg[6]/NET0131  ;
  input \core_dag_ilm1reg_I_reg[7]/NET0131  ;
  input \core_dag_ilm1reg_I_reg[8]/NET0131  ;
  input \core_dag_ilm1reg_I_reg[9]/NET0131  ;
  input \core_dag_ilm1reg_L0_we_DO_reg[0]/NET0131  ;
  input \core_dag_ilm1reg_L0_we_DO_reg[10]/NET0131  ;
  input \core_dag_ilm1reg_L0_we_DO_reg[11]/NET0131  ;
  input \core_dag_ilm1reg_L0_we_DO_reg[12]/NET0131  ;
  input \core_dag_ilm1reg_L0_we_DO_reg[13]/NET0131  ;
  input \core_dag_ilm1reg_L0_we_DO_reg[1]/NET0131  ;
  input \core_dag_ilm1reg_L0_we_DO_reg[2]/NET0131  ;
  input \core_dag_ilm1reg_L0_we_DO_reg[3]/NET0131  ;
  input \core_dag_ilm1reg_L0_we_DO_reg[4]/NET0131  ;
  input \core_dag_ilm1reg_L0_we_DO_reg[5]/NET0131  ;
  input \core_dag_ilm1reg_L0_we_DO_reg[6]/NET0131  ;
  input \core_dag_ilm1reg_L0_we_DO_reg[7]/NET0131  ;
  input \core_dag_ilm1reg_L0_we_DO_reg[8]/NET0131  ;
  input \core_dag_ilm1reg_L0_we_DO_reg[9]/NET0131  ;
  input \core_dag_ilm1reg_L1_we_DO_reg[0]/NET0131  ;
  input \core_dag_ilm1reg_L1_we_DO_reg[10]/NET0131  ;
  input \core_dag_ilm1reg_L1_we_DO_reg[11]/NET0131  ;
  input \core_dag_ilm1reg_L1_we_DO_reg[12]/NET0131  ;
  input \core_dag_ilm1reg_L1_we_DO_reg[13]/NET0131  ;
  input \core_dag_ilm1reg_L1_we_DO_reg[1]/NET0131  ;
  input \core_dag_ilm1reg_L1_we_DO_reg[2]/NET0131  ;
  input \core_dag_ilm1reg_L1_we_DO_reg[3]/NET0131  ;
  input \core_dag_ilm1reg_L1_we_DO_reg[4]/NET0131  ;
  input \core_dag_ilm1reg_L1_we_DO_reg[5]/NET0131  ;
  input \core_dag_ilm1reg_L1_we_DO_reg[6]/NET0131  ;
  input \core_dag_ilm1reg_L1_we_DO_reg[7]/NET0131  ;
  input \core_dag_ilm1reg_L1_we_DO_reg[8]/NET0131  ;
  input \core_dag_ilm1reg_L1_we_DO_reg[9]/NET0131  ;
  input \core_dag_ilm1reg_L2_we_DO_reg[0]/NET0131  ;
  input \core_dag_ilm1reg_L2_we_DO_reg[10]/NET0131  ;
  input \core_dag_ilm1reg_L2_we_DO_reg[11]/NET0131  ;
  input \core_dag_ilm1reg_L2_we_DO_reg[12]/NET0131  ;
  input \core_dag_ilm1reg_L2_we_DO_reg[13]/NET0131  ;
  input \core_dag_ilm1reg_L2_we_DO_reg[1]/NET0131  ;
  input \core_dag_ilm1reg_L2_we_DO_reg[2]/NET0131  ;
  input \core_dag_ilm1reg_L2_we_DO_reg[3]/NET0131  ;
  input \core_dag_ilm1reg_L2_we_DO_reg[4]/NET0131  ;
  input \core_dag_ilm1reg_L2_we_DO_reg[5]/NET0131  ;
  input \core_dag_ilm1reg_L2_we_DO_reg[6]/NET0131  ;
  input \core_dag_ilm1reg_L2_we_DO_reg[7]/NET0131  ;
  input \core_dag_ilm1reg_L2_we_DO_reg[8]/NET0131  ;
  input \core_dag_ilm1reg_L2_we_DO_reg[9]/NET0131  ;
  input \core_dag_ilm1reg_L3_we_DO_reg[0]/NET0131  ;
  input \core_dag_ilm1reg_L3_we_DO_reg[10]/NET0131  ;
  input \core_dag_ilm1reg_L3_we_DO_reg[11]/NET0131  ;
  input \core_dag_ilm1reg_L3_we_DO_reg[12]/NET0131  ;
  input \core_dag_ilm1reg_L3_we_DO_reg[13]/NET0131  ;
  input \core_dag_ilm1reg_L3_we_DO_reg[1]/NET0131  ;
  input \core_dag_ilm1reg_L3_we_DO_reg[2]/NET0131  ;
  input \core_dag_ilm1reg_L3_we_DO_reg[3]/NET0131  ;
  input \core_dag_ilm1reg_L3_we_DO_reg[4]/NET0131  ;
  input \core_dag_ilm1reg_L3_we_DO_reg[5]/NET0131  ;
  input \core_dag_ilm1reg_L3_we_DO_reg[6]/NET0131  ;
  input \core_dag_ilm1reg_L3_we_DO_reg[7]/NET0131  ;
  input \core_dag_ilm1reg_L3_we_DO_reg[8]/NET0131  ;
  input \core_dag_ilm1reg_L3_we_DO_reg[9]/NET0131  ;
  input \core_dag_ilm1reg_L_reg[0]/NET0131  ;
  input \core_dag_ilm1reg_L_reg[10]/NET0131  ;
  input \core_dag_ilm1reg_L_reg[11]/NET0131  ;
  input \core_dag_ilm1reg_L_reg[12]/NET0131  ;
  input \core_dag_ilm1reg_L_reg[13]/NET0131  ;
  input \core_dag_ilm1reg_L_reg[1]/NET0131  ;
  input \core_dag_ilm1reg_L_reg[2]/NET0131  ;
  input \core_dag_ilm1reg_L_reg[3]/NET0131  ;
  input \core_dag_ilm1reg_L_reg[4]/NET0131  ;
  input \core_dag_ilm1reg_L_reg[5]/NET0131  ;
  input \core_dag_ilm1reg_L_reg[6]/NET0131  ;
  input \core_dag_ilm1reg_L_reg[7]/NET0131  ;
  input \core_dag_ilm1reg_L_reg[8]/NET0131  ;
  input \core_dag_ilm1reg_L_reg[9]/NET0131  ;
  input \core_dag_ilm1reg_M0_we_DO_reg[0]/NET0131  ;
  input \core_dag_ilm1reg_M0_we_DO_reg[10]/NET0131  ;
  input \core_dag_ilm1reg_M0_we_DO_reg[11]/NET0131  ;
  input \core_dag_ilm1reg_M0_we_DO_reg[12]/NET0131  ;
  input \core_dag_ilm1reg_M0_we_DO_reg[13]/NET0131  ;
  input \core_dag_ilm1reg_M0_we_DO_reg[1]/NET0131  ;
  input \core_dag_ilm1reg_M0_we_DO_reg[2]/NET0131  ;
  input \core_dag_ilm1reg_M0_we_DO_reg[3]/NET0131  ;
  input \core_dag_ilm1reg_M0_we_DO_reg[4]/NET0131  ;
  input \core_dag_ilm1reg_M0_we_DO_reg[5]/NET0131  ;
  input \core_dag_ilm1reg_M0_we_DO_reg[6]/NET0131  ;
  input \core_dag_ilm1reg_M0_we_DO_reg[7]/NET0131  ;
  input \core_dag_ilm1reg_M0_we_DO_reg[8]/NET0131  ;
  input \core_dag_ilm1reg_M0_we_DO_reg[9]/NET0131  ;
  input \core_dag_ilm1reg_M1_we_DO_reg[0]/NET0131  ;
  input \core_dag_ilm1reg_M1_we_DO_reg[10]/NET0131  ;
  input \core_dag_ilm1reg_M1_we_DO_reg[11]/NET0131  ;
  input \core_dag_ilm1reg_M1_we_DO_reg[12]/NET0131  ;
  input \core_dag_ilm1reg_M1_we_DO_reg[13]/NET0131  ;
  input \core_dag_ilm1reg_M1_we_DO_reg[1]/NET0131  ;
  input \core_dag_ilm1reg_M1_we_DO_reg[2]/NET0131  ;
  input \core_dag_ilm1reg_M1_we_DO_reg[3]/NET0131  ;
  input \core_dag_ilm1reg_M1_we_DO_reg[4]/NET0131  ;
  input \core_dag_ilm1reg_M1_we_DO_reg[5]/NET0131  ;
  input \core_dag_ilm1reg_M1_we_DO_reg[6]/NET0131  ;
  input \core_dag_ilm1reg_M1_we_DO_reg[7]/NET0131  ;
  input \core_dag_ilm1reg_M1_we_DO_reg[8]/NET0131  ;
  input \core_dag_ilm1reg_M1_we_DO_reg[9]/NET0131  ;
  input \core_dag_ilm1reg_M2_we_DO_reg[0]/NET0131  ;
  input \core_dag_ilm1reg_M2_we_DO_reg[10]/NET0131  ;
  input \core_dag_ilm1reg_M2_we_DO_reg[11]/NET0131  ;
  input \core_dag_ilm1reg_M2_we_DO_reg[12]/NET0131  ;
  input \core_dag_ilm1reg_M2_we_DO_reg[13]/NET0131  ;
  input \core_dag_ilm1reg_M2_we_DO_reg[1]/NET0131  ;
  input \core_dag_ilm1reg_M2_we_DO_reg[2]/NET0131  ;
  input \core_dag_ilm1reg_M2_we_DO_reg[3]/NET0131  ;
  input \core_dag_ilm1reg_M2_we_DO_reg[4]/NET0131  ;
  input \core_dag_ilm1reg_M2_we_DO_reg[5]/NET0131  ;
  input \core_dag_ilm1reg_M2_we_DO_reg[6]/NET0131  ;
  input \core_dag_ilm1reg_M2_we_DO_reg[7]/NET0131  ;
  input \core_dag_ilm1reg_M2_we_DO_reg[8]/NET0131  ;
  input \core_dag_ilm1reg_M2_we_DO_reg[9]/NET0131  ;
  input \core_dag_ilm1reg_M3_we_DO_reg[0]/NET0131  ;
  input \core_dag_ilm1reg_M3_we_DO_reg[10]/NET0131  ;
  input \core_dag_ilm1reg_M3_we_DO_reg[11]/NET0131  ;
  input \core_dag_ilm1reg_M3_we_DO_reg[12]/NET0131  ;
  input \core_dag_ilm1reg_M3_we_DO_reg[13]/NET0131  ;
  input \core_dag_ilm1reg_M3_we_DO_reg[1]/NET0131  ;
  input \core_dag_ilm1reg_M3_we_DO_reg[2]/NET0131  ;
  input \core_dag_ilm1reg_M3_we_DO_reg[3]/NET0131  ;
  input \core_dag_ilm1reg_M3_we_DO_reg[4]/NET0131  ;
  input \core_dag_ilm1reg_M3_we_DO_reg[5]/NET0131  ;
  input \core_dag_ilm1reg_M3_we_DO_reg[6]/NET0131  ;
  input \core_dag_ilm1reg_M3_we_DO_reg[7]/NET0131  ;
  input \core_dag_ilm1reg_M3_we_DO_reg[8]/NET0131  ;
  input \core_dag_ilm1reg_M3_we_DO_reg[9]/NET0131  ;
  input \core_dag_ilm1reg_M_reg[0]/NET0131  ;
  input \core_dag_ilm1reg_M_reg[10]/NET0131  ;
  input \core_dag_ilm1reg_M_reg[11]/NET0131  ;
  input \core_dag_ilm1reg_M_reg[12]/NET0131  ;
  input \core_dag_ilm1reg_M_reg[13]/NET0131  ;
  input \core_dag_ilm1reg_M_reg[1]/NET0131  ;
  input \core_dag_ilm1reg_M_reg[2]/NET0131  ;
  input \core_dag_ilm1reg_M_reg[3]/NET0131  ;
  input \core_dag_ilm1reg_M_reg[4]/NET0131  ;
  input \core_dag_ilm1reg_M_reg[5]/NET0131  ;
  input \core_dag_ilm1reg_M_reg[6]/NET0131  ;
  input \core_dag_ilm1reg_M_reg[7]/NET0131  ;
  input \core_dag_ilm1reg_M_reg[8]/NET0131  ;
  input \core_dag_ilm1reg_M_reg[9]/NET0131  ;
  input \core_dag_ilm1reg_STAC_pi_DO_reg[0]/NET0131  ;
  input \core_dag_ilm1reg_STAC_pi_DO_reg[10]/NET0131  ;
  input \core_dag_ilm1reg_STAC_pi_DO_reg[11]/NET0131  ;
  input \core_dag_ilm1reg_STAC_pi_DO_reg[12]/NET0131  ;
  input \core_dag_ilm1reg_STAC_pi_DO_reg[13]/NET0131  ;
  input \core_dag_ilm1reg_STAC_pi_DO_reg[1]/NET0131  ;
  input \core_dag_ilm1reg_STAC_pi_DO_reg[2]/NET0131  ;
  input \core_dag_ilm1reg_STAC_pi_DO_reg[3]/NET0131  ;
  input \core_dag_ilm1reg_STAC_pi_DO_reg[4]/NET0131  ;
  input \core_dag_ilm1reg_STAC_pi_DO_reg[5]/NET0131  ;
  input \core_dag_ilm1reg_STAC_pi_DO_reg[6]/NET0131  ;
  input \core_dag_ilm1reg_STAC_pi_DO_reg[7]/NET0131  ;
  input \core_dag_ilm1reg_STAC_pi_DO_reg[8]/NET0131  ;
  input \core_dag_ilm1reg_STAC_pi_DO_reg[9]/NET0131  ;
  input \core_dag_ilm1reg_STEALI_E_reg[0]/P0001  ;
  input \core_dag_ilm1reg_STEALI_E_reg[1]/P0001  ;
  input \core_dag_ilm1reg_STEALI_E_reg[2]/P0001  ;
  input \core_dag_ilm2reg_I4_we_DO_reg[0]/NET0131  ;
  input \core_dag_ilm2reg_I4_we_DO_reg[10]/NET0131  ;
  input \core_dag_ilm2reg_I4_we_DO_reg[11]/NET0131  ;
  input \core_dag_ilm2reg_I4_we_DO_reg[12]/NET0131  ;
  input \core_dag_ilm2reg_I4_we_DO_reg[13]/NET0131  ;
  input \core_dag_ilm2reg_I4_we_DO_reg[1]/NET0131  ;
  input \core_dag_ilm2reg_I4_we_DO_reg[2]/NET0131  ;
  input \core_dag_ilm2reg_I4_we_DO_reg[3]/NET0131  ;
  input \core_dag_ilm2reg_I4_we_DO_reg[4]/NET0131  ;
  input \core_dag_ilm2reg_I4_we_DO_reg[5]/NET0131  ;
  input \core_dag_ilm2reg_I4_we_DO_reg[6]/NET0131  ;
  input \core_dag_ilm2reg_I4_we_DO_reg[7]/NET0131  ;
  input \core_dag_ilm2reg_I4_we_DO_reg[8]/NET0131  ;
  input \core_dag_ilm2reg_I4_we_DO_reg[9]/NET0131  ;
  input \core_dag_ilm2reg_I5_we_DO_reg[0]/NET0131  ;
  input \core_dag_ilm2reg_I5_we_DO_reg[10]/NET0131  ;
  input \core_dag_ilm2reg_I5_we_DO_reg[11]/NET0131  ;
  input \core_dag_ilm2reg_I5_we_DO_reg[12]/NET0131  ;
  input \core_dag_ilm2reg_I5_we_DO_reg[13]/NET0131  ;
  input \core_dag_ilm2reg_I5_we_DO_reg[1]/NET0131  ;
  input \core_dag_ilm2reg_I5_we_DO_reg[2]/NET0131  ;
  input \core_dag_ilm2reg_I5_we_DO_reg[3]/NET0131  ;
  input \core_dag_ilm2reg_I5_we_DO_reg[4]/NET0131  ;
  input \core_dag_ilm2reg_I5_we_DO_reg[5]/NET0131  ;
  input \core_dag_ilm2reg_I5_we_DO_reg[6]/NET0131  ;
  input \core_dag_ilm2reg_I5_we_DO_reg[7]/NET0131  ;
  input \core_dag_ilm2reg_I5_we_DO_reg[8]/NET0131  ;
  input \core_dag_ilm2reg_I5_we_DO_reg[9]/NET0131  ;
  input \core_dag_ilm2reg_I6_we_DO_reg[0]/NET0131  ;
  input \core_dag_ilm2reg_I6_we_DO_reg[10]/NET0131  ;
  input \core_dag_ilm2reg_I6_we_DO_reg[11]/NET0131  ;
  input \core_dag_ilm2reg_I6_we_DO_reg[12]/NET0131  ;
  input \core_dag_ilm2reg_I6_we_DO_reg[13]/NET0131  ;
  input \core_dag_ilm2reg_I6_we_DO_reg[1]/NET0131  ;
  input \core_dag_ilm2reg_I6_we_DO_reg[2]/NET0131  ;
  input \core_dag_ilm2reg_I6_we_DO_reg[3]/NET0131  ;
  input \core_dag_ilm2reg_I6_we_DO_reg[4]/NET0131  ;
  input \core_dag_ilm2reg_I6_we_DO_reg[5]/NET0131  ;
  input \core_dag_ilm2reg_I6_we_DO_reg[6]/NET0131  ;
  input \core_dag_ilm2reg_I6_we_DO_reg[7]/NET0131  ;
  input \core_dag_ilm2reg_I6_we_DO_reg[8]/NET0131  ;
  input \core_dag_ilm2reg_I6_we_DO_reg[9]/NET0131  ;
  input \core_dag_ilm2reg_I7_we_DO_reg[0]/NET0131  ;
  input \core_dag_ilm2reg_I7_we_DO_reg[10]/NET0131  ;
  input \core_dag_ilm2reg_I7_we_DO_reg[11]/NET0131  ;
  input \core_dag_ilm2reg_I7_we_DO_reg[12]/NET0131  ;
  input \core_dag_ilm2reg_I7_we_DO_reg[13]/NET0131  ;
  input \core_dag_ilm2reg_I7_we_DO_reg[1]/NET0131  ;
  input \core_dag_ilm2reg_I7_we_DO_reg[2]/NET0131  ;
  input \core_dag_ilm2reg_I7_we_DO_reg[3]/NET0131  ;
  input \core_dag_ilm2reg_I7_we_DO_reg[4]/NET0131  ;
  input \core_dag_ilm2reg_I7_we_DO_reg[5]/NET0131  ;
  input \core_dag_ilm2reg_I7_we_DO_reg[6]/NET0131  ;
  input \core_dag_ilm2reg_I7_we_DO_reg[7]/NET0131  ;
  input \core_dag_ilm2reg_I7_we_DO_reg[8]/NET0131  ;
  input \core_dag_ilm2reg_I7_we_DO_reg[9]/NET0131  ;
  input \core_dag_ilm2reg_IL_E_reg[0]/P0001  ;
  input \core_dag_ilm2reg_IL_E_reg[1]/P0001  ;
  input \core_dag_ilm2reg_I_reg[0]/NET0131  ;
  input \core_dag_ilm2reg_I_reg[10]/NET0131  ;
  input \core_dag_ilm2reg_I_reg[11]/NET0131  ;
  input \core_dag_ilm2reg_I_reg[12]/NET0131  ;
  input \core_dag_ilm2reg_I_reg[13]/NET0131  ;
  input \core_dag_ilm2reg_I_reg[1]/NET0131  ;
  input \core_dag_ilm2reg_I_reg[2]/NET0131  ;
  input \core_dag_ilm2reg_I_reg[3]/NET0131  ;
  input \core_dag_ilm2reg_I_reg[4]/NET0131  ;
  input \core_dag_ilm2reg_I_reg[5]/NET0131  ;
  input \core_dag_ilm2reg_I_reg[6]/NET0131  ;
  input \core_dag_ilm2reg_I_reg[7]/NET0131  ;
  input \core_dag_ilm2reg_I_reg[8]/NET0131  ;
  input \core_dag_ilm2reg_I_reg[9]/NET0131  ;
  input \core_dag_ilm2reg_L4_we_DO_reg[0]/NET0131  ;
  input \core_dag_ilm2reg_L4_we_DO_reg[10]/NET0131  ;
  input \core_dag_ilm2reg_L4_we_DO_reg[11]/NET0131  ;
  input \core_dag_ilm2reg_L4_we_DO_reg[12]/NET0131  ;
  input \core_dag_ilm2reg_L4_we_DO_reg[13]/NET0131  ;
  input \core_dag_ilm2reg_L4_we_DO_reg[1]/NET0131  ;
  input \core_dag_ilm2reg_L4_we_DO_reg[2]/NET0131  ;
  input \core_dag_ilm2reg_L4_we_DO_reg[3]/NET0131  ;
  input \core_dag_ilm2reg_L4_we_DO_reg[4]/NET0131  ;
  input \core_dag_ilm2reg_L4_we_DO_reg[5]/NET0131  ;
  input \core_dag_ilm2reg_L4_we_DO_reg[6]/NET0131  ;
  input \core_dag_ilm2reg_L4_we_DO_reg[7]/NET0131  ;
  input \core_dag_ilm2reg_L4_we_DO_reg[8]/NET0131  ;
  input \core_dag_ilm2reg_L4_we_DO_reg[9]/NET0131  ;
  input \core_dag_ilm2reg_L5_we_DO_reg[0]/NET0131  ;
  input \core_dag_ilm2reg_L5_we_DO_reg[10]/NET0131  ;
  input \core_dag_ilm2reg_L5_we_DO_reg[11]/NET0131  ;
  input \core_dag_ilm2reg_L5_we_DO_reg[12]/NET0131  ;
  input \core_dag_ilm2reg_L5_we_DO_reg[13]/NET0131  ;
  input \core_dag_ilm2reg_L5_we_DO_reg[1]/NET0131  ;
  input \core_dag_ilm2reg_L5_we_DO_reg[2]/NET0131  ;
  input \core_dag_ilm2reg_L5_we_DO_reg[3]/NET0131  ;
  input \core_dag_ilm2reg_L5_we_DO_reg[4]/NET0131  ;
  input \core_dag_ilm2reg_L5_we_DO_reg[5]/NET0131  ;
  input \core_dag_ilm2reg_L5_we_DO_reg[6]/NET0131  ;
  input \core_dag_ilm2reg_L5_we_DO_reg[7]/NET0131  ;
  input \core_dag_ilm2reg_L5_we_DO_reg[8]/NET0131  ;
  input \core_dag_ilm2reg_L5_we_DO_reg[9]/NET0131  ;
  input \core_dag_ilm2reg_L6_we_DO_reg[0]/NET0131  ;
  input \core_dag_ilm2reg_L6_we_DO_reg[10]/NET0131  ;
  input \core_dag_ilm2reg_L6_we_DO_reg[11]/NET0131  ;
  input \core_dag_ilm2reg_L6_we_DO_reg[12]/NET0131  ;
  input \core_dag_ilm2reg_L6_we_DO_reg[13]/NET0131  ;
  input \core_dag_ilm2reg_L6_we_DO_reg[1]/NET0131  ;
  input \core_dag_ilm2reg_L6_we_DO_reg[2]/NET0131  ;
  input \core_dag_ilm2reg_L6_we_DO_reg[3]/NET0131  ;
  input \core_dag_ilm2reg_L6_we_DO_reg[4]/NET0131  ;
  input \core_dag_ilm2reg_L6_we_DO_reg[5]/NET0131  ;
  input \core_dag_ilm2reg_L6_we_DO_reg[6]/NET0131  ;
  input \core_dag_ilm2reg_L6_we_DO_reg[7]/NET0131  ;
  input \core_dag_ilm2reg_L6_we_DO_reg[8]/NET0131  ;
  input \core_dag_ilm2reg_L6_we_DO_reg[9]/NET0131  ;
  input \core_dag_ilm2reg_L7_we_DO_reg[0]/NET0131  ;
  input \core_dag_ilm2reg_L7_we_DO_reg[10]/NET0131  ;
  input \core_dag_ilm2reg_L7_we_DO_reg[11]/NET0131  ;
  input \core_dag_ilm2reg_L7_we_DO_reg[12]/NET0131  ;
  input \core_dag_ilm2reg_L7_we_DO_reg[13]/NET0131  ;
  input \core_dag_ilm2reg_L7_we_DO_reg[1]/NET0131  ;
  input \core_dag_ilm2reg_L7_we_DO_reg[2]/NET0131  ;
  input \core_dag_ilm2reg_L7_we_DO_reg[3]/NET0131  ;
  input \core_dag_ilm2reg_L7_we_DO_reg[4]/NET0131  ;
  input \core_dag_ilm2reg_L7_we_DO_reg[5]/NET0131  ;
  input \core_dag_ilm2reg_L7_we_DO_reg[6]/NET0131  ;
  input \core_dag_ilm2reg_L7_we_DO_reg[7]/NET0131  ;
  input \core_dag_ilm2reg_L7_we_DO_reg[8]/NET0131  ;
  input \core_dag_ilm2reg_L7_we_DO_reg[9]/NET0131  ;
  input \core_dag_ilm2reg_L_reg[0]/NET0131  ;
  input \core_dag_ilm2reg_L_reg[10]/NET0131  ;
  input \core_dag_ilm2reg_L_reg[11]/NET0131  ;
  input \core_dag_ilm2reg_L_reg[12]/NET0131  ;
  input \core_dag_ilm2reg_L_reg[13]/NET0131  ;
  input \core_dag_ilm2reg_L_reg[1]/NET0131  ;
  input \core_dag_ilm2reg_L_reg[2]/NET0131  ;
  input \core_dag_ilm2reg_L_reg[3]/NET0131  ;
  input \core_dag_ilm2reg_L_reg[4]/NET0131  ;
  input \core_dag_ilm2reg_L_reg[5]/NET0131  ;
  input \core_dag_ilm2reg_L_reg[6]/NET0131  ;
  input \core_dag_ilm2reg_L_reg[7]/NET0131  ;
  input \core_dag_ilm2reg_L_reg[8]/NET0131  ;
  input \core_dag_ilm2reg_L_reg[9]/NET0131  ;
  input \core_dag_ilm2reg_M4_we_DO_reg[0]/NET0131  ;
  input \core_dag_ilm2reg_M4_we_DO_reg[10]/NET0131  ;
  input \core_dag_ilm2reg_M4_we_DO_reg[11]/NET0131  ;
  input \core_dag_ilm2reg_M4_we_DO_reg[12]/NET0131  ;
  input \core_dag_ilm2reg_M4_we_DO_reg[13]/NET0131  ;
  input \core_dag_ilm2reg_M4_we_DO_reg[1]/NET0131  ;
  input \core_dag_ilm2reg_M4_we_DO_reg[2]/NET0131  ;
  input \core_dag_ilm2reg_M4_we_DO_reg[3]/NET0131  ;
  input \core_dag_ilm2reg_M4_we_DO_reg[4]/NET0131  ;
  input \core_dag_ilm2reg_M4_we_DO_reg[5]/NET0131  ;
  input \core_dag_ilm2reg_M4_we_DO_reg[6]/NET0131  ;
  input \core_dag_ilm2reg_M4_we_DO_reg[7]/NET0131  ;
  input \core_dag_ilm2reg_M4_we_DO_reg[8]/NET0131  ;
  input \core_dag_ilm2reg_M4_we_DO_reg[9]/NET0131  ;
  input \core_dag_ilm2reg_M5_we_DO_reg[0]/NET0131  ;
  input \core_dag_ilm2reg_M5_we_DO_reg[10]/NET0131  ;
  input \core_dag_ilm2reg_M5_we_DO_reg[11]/NET0131  ;
  input \core_dag_ilm2reg_M5_we_DO_reg[12]/NET0131  ;
  input \core_dag_ilm2reg_M5_we_DO_reg[13]/NET0131  ;
  input \core_dag_ilm2reg_M5_we_DO_reg[1]/NET0131  ;
  input \core_dag_ilm2reg_M5_we_DO_reg[2]/NET0131  ;
  input \core_dag_ilm2reg_M5_we_DO_reg[3]/NET0131  ;
  input \core_dag_ilm2reg_M5_we_DO_reg[4]/NET0131  ;
  input \core_dag_ilm2reg_M5_we_DO_reg[5]/NET0131  ;
  input \core_dag_ilm2reg_M5_we_DO_reg[6]/NET0131  ;
  input \core_dag_ilm2reg_M5_we_DO_reg[7]/NET0131  ;
  input \core_dag_ilm2reg_M5_we_DO_reg[8]/NET0131  ;
  input \core_dag_ilm2reg_M5_we_DO_reg[9]/NET0131  ;
  input \core_dag_ilm2reg_M6_we_DO_reg[0]/NET0131  ;
  input \core_dag_ilm2reg_M6_we_DO_reg[10]/NET0131  ;
  input \core_dag_ilm2reg_M6_we_DO_reg[11]/NET0131  ;
  input \core_dag_ilm2reg_M6_we_DO_reg[12]/NET0131  ;
  input \core_dag_ilm2reg_M6_we_DO_reg[13]/NET0131  ;
  input \core_dag_ilm2reg_M6_we_DO_reg[1]/NET0131  ;
  input \core_dag_ilm2reg_M6_we_DO_reg[2]/NET0131  ;
  input \core_dag_ilm2reg_M6_we_DO_reg[3]/NET0131  ;
  input \core_dag_ilm2reg_M6_we_DO_reg[4]/NET0131  ;
  input \core_dag_ilm2reg_M6_we_DO_reg[5]/NET0131  ;
  input \core_dag_ilm2reg_M6_we_DO_reg[6]/NET0131  ;
  input \core_dag_ilm2reg_M6_we_DO_reg[7]/NET0131  ;
  input \core_dag_ilm2reg_M6_we_DO_reg[8]/NET0131  ;
  input \core_dag_ilm2reg_M6_we_DO_reg[9]/NET0131  ;
  input \core_dag_ilm2reg_M7_we_DO_reg[0]/NET0131  ;
  input \core_dag_ilm2reg_M7_we_DO_reg[10]/NET0131  ;
  input \core_dag_ilm2reg_M7_we_DO_reg[11]/NET0131  ;
  input \core_dag_ilm2reg_M7_we_DO_reg[12]/NET0131  ;
  input \core_dag_ilm2reg_M7_we_DO_reg[13]/NET0131  ;
  input \core_dag_ilm2reg_M7_we_DO_reg[1]/NET0131  ;
  input \core_dag_ilm2reg_M7_we_DO_reg[2]/NET0131  ;
  input \core_dag_ilm2reg_M7_we_DO_reg[3]/NET0131  ;
  input \core_dag_ilm2reg_M7_we_DO_reg[4]/NET0131  ;
  input \core_dag_ilm2reg_M7_we_DO_reg[5]/NET0131  ;
  input \core_dag_ilm2reg_M7_we_DO_reg[6]/NET0131  ;
  input \core_dag_ilm2reg_M7_we_DO_reg[7]/NET0131  ;
  input \core_dag_ilm2reg_M7_we_DO_reg[8]/NET0131  ;
  input \core_dag_ilm2reg_M7_we_DO_reg[9]/NET0131  ;
  input \core_dag_ilm2reg_M_E_reg[0]/NET0131  ;
  input \core_dag_ilm2reg_M_E_reg[1]/NET0131  ;
  input \core_dag_ilm2reg_M_reg[0]/NET0131  ;
  input \core_dag_ilm2reg_M_reg[10]/NET0131  ;
  input \core_dag_ilm2reg_M_reg[11]/NET0131  ;
  input \core_dag_ilm2reg_M_reg[12]/NET0131  ;
  input \core_dag_ilm2reg_M_reg[13]/NET0131  ;
  input \core_dag_ilm2reg_M_reg[1]/NET0131  ;
  input \core_dag_ilm2reg_M_reg[2]/NET0131  ;
  input \core_dag_ilm2reg_M_reg[3]/NET0131  ;
  input \core_dag_ilm2reg_M_reg[4]/NET0131  ;
  input \core_dag_ilm2reg_M_reg[5]/NET0131  ;
  input \core_dag_ilm2reg_M_reg[6]/NET0131  ;
  input \core_dag_ilm2reg_M_reg[7]/NET0131  ;
  input \core_dag_ilm2reg_M_reg[8]/NET0131  ;
  input \core_dag_ilm2reg_M_reg[9]/NET0131  ;
  input \core_dag_ilm2reg_PMA_pi_DO_reg[0]/NET0131  ;
  input \core_dag_ilm2reg_PMA_pi_DO_reg[10]/NET0131  ;
  input \core_dag_ilm2reg_PMA_pi_DO_reg[11]/NET0131  ;
  input \core_dag_ilm2reg_PMA_pi_DO_reg[12]/NET0131  ;
  input \core_dag_ilm2reg_PMA_pi_DO_reg[13]/NET0131  ;
  input \core_dag_ilm2reg_PMA_pi_DO_reg[1]/NET0131  ;
  input \core_dag_ilm2reg_PMA_pi_DO_reg[2]/NET0131  ;
  input \core_dag_ilm2reg_PMA_pi_DO_reg[3]/NET0131  ;
  input \core_dag_ilm2reg_PMA_pi_DO_reg[4]/NET0131  ;
  input \core_dag_ilm2reg_PMA_pi_DO_reg[5]/NET0131  ;
  input \core_dag_ilm2reg_PMA_pi_DO_reg[6]/NET0131  ;
  input \core_dag_ilm2reg_PMA_pi_DO_reg[7]/NET0131  ;
  input \core_dag_ilm2reg_PMA_pi_DO_reg[8]/NET0131  ;
  input \core_dag_ilm2reg_PMA_pi_DO_reg[9]/NET0131  ;
  input \core_dag_modulo1_R0wrap_reg/P0001  ;
  input \core_dag_modulo1_R1wrap_reg/P0001  ;
  input \core_dag_modulo1_T0wrap_reg/P0001  ;
  input \core_dag_modulo1_T1wrap_reg/P0001  ;
  input \core_eu_ea_alu_ea_dec_AMF_E_reg[0]/NET0131  ;
  input \core_eu_ea_alu_ea_dec_AMF_E_reg[1]/NET0131  ;
  input \core_eu_ea_alu_ea_dec_AMF_E_reg[2]/NET0131  ;
  input \core_eu_ea_alu_ea_dec_AMF_E_reg[3]/NET0131  ;
  input \core_eu_ea_alu_ea_dec_AMF_E_reg[4]/NET0131  ;
  input \core_eu_ea_alu_ea_dec_piconst_DO_reg[0]/P0001  ;
  input \core_eu_ea_alu_ea_dec_piconst_DO_reg[10]/P0001  ;
  input \core_eu_ea_alu_ea_dec_piconst_DO_reg[11]/P0001  ;
  input \core_eu_ea_alu_ea_dec_piconst_DO_reg[12]/P0001  ;
  input \core_eu_ea_alu_ea_dec_piconst_DO_reg[13]/P0001  ;
  input \core_eu_ea_alu_ea_dec_piconst_DO_reg[14]/P0001  ;
  input \core_eu_ea_alu_ea_dec_piconst_DO_reg[15]/P0001  ;
  input \core_eu_ea_alu_ea_dec_piconst_DO_reg[1]/P0001  ;
  input \core_eu_ea_alu_ea_dec_piconst_DO_reg[2]/P0001  ;
  input \core_eu_ea_alu_ea_dec_piconst_DO_reg[3]/P0001  ;
  input \core_eu_ea_alu_ea_dec_piconst_DO_reg[4]/P0001  ;
  input \core_eu_ea_alu_ea_dec_piconst_DO_reg[5]/P0001  ;
  input \core_eu_ea_alu_ea_dec_piconst_DO_reg[6]/P0001  ;
  input \core_eu_ea_alu_ea_dec_piconst_DO_reg[7]/P0001  ;
  input \core_eu_ea_alu_ea_dec_piconst_DO_reg[8]/P0001  ;
  input \core_eu_ea_alu_ea_dec_piconst_DO_reg[9]/P0001  ;
  input \core_eu_ea_alu_ea_reg_afrwe_DO_reg[0]/P0001  ;
  input \core_eu_ea_alu_ea_reg_afrwe_DO_reg[10]/P0001  ;
  input \core_eu_ea_alu_ea_reg_afrwe_DO_reg[11]/P0001  ;
  input \core_eu_ea_alu_ea_reg_afrwe_DO_reg[12]/P0001  ;
  input \core_eu_ea_alu_ea_reg_afrwe_DO_reg[13]/P0001  ;
  input \core_eu_ea_alu_ea_reg_afrwe_DO_reg[14]/P0001  ;
  input \core_eu_ea_alu_ea_reg_afrwe_DO_reg[15]/P0001  ;
  input \core_eu_ea_alu_ea_reg_afrwe_DO_reg[1]/P0001  ;
  input \core_eu_ea_alu_ea_reg_afrwe_DO_reg[2]/P0001  ;
  input \core_eu_ea_alu_ea_reg_afrwe_DO_reg[3]/P0001  ;
  input \core_eu_ea_alu_ea_reg_afrwe_DO_reg[4]/P0001  ;
  input \core_eu_ea_alu_ea_reg_afrwe_DO_reg[5]/P0001  ;
  input \core_eu_ea_alu_ea_reg_afrwe_DO_reg[6]/P0001  ;
  input \core_eu_ea_alu_ea_reg_afrwe_DO_reg[7]/P0001  ;
  input \core_eu_ea_alu_ea_reg_afrwe_DO_reg[8]/P0001  ;
  input \core_eu_ea_alu_ea_reg_afrwe_DO_reg[9]/P0001  ;
  input \core_eu_ea_alu_ea_reg_afswe_DO_reg[0]/P0001  ;
  input \core_eu_ea_alu_ea_reg_afswe_DO_reg[10]/P0001  ;
  input \core_eu_ea_alu_ea_reg_afswe_DO_reg[11]/P0001  ;
  input \core_eu_ea_alu_ea_reg_afswe_DO_reg[12]/P0001  ;
  input \core_eu_ea_alu_ea_reg_afswe_DO_reg[13]/P0001  ;
  input \core_eu_ea_alu_ea_reg_afswe_DO_reg[14]/P0001  ;
  input \core_eu_ea_alu_ea_reg_afswe_DO_reg[15]/P0001  ;
  input \core_eu_ea_alu_ea_reg_afswe_DO_reg[1]/P0001  ;
  input \core_eu_ea_alu_ea_reg_afswe_DO_reg[2]/P0001  ;
  input \core_eu_ea_alu_ea_reg_afswe_DO_reg[3]/P0001  ;
  input \core_eu_ea_alu_ea_reg_afswe_DO_reg[4]/P0001  ;
  input \core_eu_ea_alu_ea_reg_afswe_DO_reg[5]/P0001  ;
  input \core_eu_ea_alu_ea_reg_afswe_DO_reg[6]/P0001  ;
  input \core_eu_ea_alu_ea_reg_afswe_DO_reg[7]/P0001  ;
  input \core_eu_ea_alu_ea_reg_afswe_DO_reg[8]/P0001  ;
  input \core_eu_ea_alu_ea_reg_afswe_DO_reg[9]/P0001  ;
  input \core_eu_ea_alu_ea_reg_arrwe_DO_reg[0]/P0001  ;
  input \core_eu_ea_alu_ea_reg_arrwe_DO_reg[10]/P0001  ;
  input \core_eu_ea_alu_ea_reg_arrwe_DO_reg[11]/P0001  ;
  input \core_eu_ea_alu_ea_reg_arrwe_DO_reg[12]/P0001  ;
  input \core_eu_ea_alu_ea_reg_arrwe_DO_reg[13]/P0001  ;
  input \core_eu_ea_alu_ea_reg_arrwe_DO_reg[14]/P0001  ;
  input \core_eu_ea_alu_ea_reg_arrwe_DO_reg[15]/P0001  ;
  input \core_eu_ea_alu_ea_reg_arrwe_DO_reg[1]/P0001  ;
  input \core_eu_ea_alu_ea_reg_arrwe_DO_reg[2]/P0001  ;
  input \core_eu_ea_alu_ea_reg_arrwe_DO_reg[3]/P0001  ;
  input \core_eu_ea_alu_ea_reg_arrwe_DO_reg[4]/P0001  ;
  input \core_eu_ea_alu_ea_reg_arrwe_DO_reg[5]/P0001  ;
  input \core_eu_ea_alu_ea_reg_arrwe_DO_reg[6]/P0001  ;
  input \core_eu_ea_alu_ea_reg_arrwe_DO_reg[7]/P0001  ;
  input \core_eu_ea_alu_ea_reg_arrwe_DO_reg[8]/P0001  ;
  input \core_eu_ea_alu_ea_reg_arrwe_DO_reg[9]/P0001  ;
  input \core_eu_ea_alu_ea_reg_arswe_DO_reg[0]/P0001  ;
  input \core_eu_ea_alu_ea_reg_arswe_DO_reg[10]/P0001  ;
  input \core_eu_ea_alu_ea_reg_arswe_DO_reg[11]/P0001  ;
  input \core_eu_ea_alu_ea_reg_arswe_DO_reg[12]/P0001  ;
  input \core_eu_ea_alu_ea_reg_arswe_DO_reg[13]/P0001  ;
  input \core_eu_ea_alu_ea_reg_arswe_DO_reg[14]/P0001  ;
  input \core_eu_ea_alu_ea_reg_arswe_DO_reg[15]/P0001  ;
  input \core_eu_ea_alu_ea_reg_arswe_DO_reg[1]/P0001  ;
  input \core_eu_ea_alu_ea_reg_arswe_DO_reg[2]/P0001  ;
  input \core_eu_ea_alu_ea_reg_arswe_DO_reg[3]/P0001  ;
  input \core_eu_ea_alu_ea_reg_arswe_DO_reg[4]/P0001  ;
  input \core_eu_ea_alu_ea_reg_arswe_DO_reg[5]/P0001  ;
  input \core_eu_ea_alu_ea_reg_arswe_DO_reg[6]/P0001  ;
  input \core_eu_ea_alu_ea_reg_arswe_DO_reg[7]/P0001  ;
  input \core_eu_ea_alu_ea_reg_arswe_DO_reg[8]/P0001  ;
  input \core_eu_ea_alu_ea_reg_arswe_DO_reg[9]/P0001  ;
  input \core_eu_ea_alu_ea_reg_ax0rwe_DO_reg[0]/P0001  ;
  input \core_eu_ea_alu_ea_reg_ax0rwe_DO_reg[10]/P0001  ;
  input \core_eu_ea_alu_ea_reg_ax0rwe_DO_reg[11]/P0001  ;
  input \core_eu_ea_alu_ea_reg_ax0rwe_DO_reg[12]/P0001  ;
  input \core_eu_ea_alu_ea_reg_ax0rwe_DO_reg[13]/P0001  ;
  input \core_eu_ea_alu_ea_reg_ax0rwe_DO_reg[14]/P0001  ;
  input \core_eu_ea_alu_ea_reg_ax0rwe_DO_reg[15]/P0001  ;
  input \core_eu_ea_alu_ea_reg_ax0rwe_DO_reg[1]/P0001  ;
  input \core_eu_ea_alu_ea_reg_ax0rwe_DO_reg[2]/P0001  ;
  input \core_eu_ea_alu_ea_reg_ax0rwe_DO_reg[3]/P0001  ;
  input \core_eu_ea_alu_ea_reg_ax0rwe_DO_reg[4]/P0001  ;
  input \core_eu_ea_alu_ea_reg_ax0rwe_DO_reg[5]/P0001  ;
  input \core_eu_ea_alu_ea_reg_ax0rwe_DO_reg[6]/P0001  ;
  input \core_eu_ea_alu_ea_reg_ax0rwe_DO_reg[7]/P0001  ;
  input \core_eu_ea_alu_ea_reg_ax0rwe_DO_reg[8]/P0001  ;
  input \core_eu_ea_alu_ea_reg_ax0rwe_DO_reg[9]/P0001  ;
  input \core_eu_ea_alu_ea_reg_ax0swe_DO_reg[0]/P0001  ;
  input \core_eu_ea_alu_ea_reg_ax0swe_DO_reg[10]/P0001  ;
  input \core_eu_ea_alu_ea_reg_ax0swe_DO_reg[11]/P0001  ;
  input \core_eu_ea_alu_ea_reg_ax0swe_DO_reg[12]/P0001  ;
  input \core_eu_ea_alu_ea_reg_ax0swe_DO_reg[13]/P0001  ;
  input \core_eu_ea_alu_ea_reg_ax0swe_DO_reg[14]/P0001  ;
  input \core_eu_ea_alu_ea_reg_ax0swe_DO_reg[15]/P0001  ;
  input \core_eu_ea_alu_ea_reg_ax0swe_DO_reg[1]/P0001  ;
  input \core_eu_ea_alu_ea_reg_ax0swe_DO_reg[2]/P0001  ;
  input \core_eu_ea_alu_ea_reg_ax0swe_DO_reg[3]/P0001  ;
  input \core_eu_ea_alu_ea_reg_ax0swe_DO_reg[4]/P0001  ;
  input \core_eu_ea_alu_ea_reg_ax0swe_DO_reg[5]/P0001  ;
  input \core_eu_ea_alu_ea_reg_ax0swe_DO_reg[6]/P0001  ;
  input \core_eu_ea_alu_ea_reg_ax0swe_DO_reg[7]/P0001  ;
  input \core_eu_ea_alu_ea_reg_ax0swe_DO_reg[8]/P0001  ;
  input \core_eu_ea_alu_ea_reg_ax0swe_DO_reg[9]/P0001  ;
  input \core_eu_ea_alu_ea_reg_ax1rwe_DO_reg[0]/P0001  ;
  input \core_eu_ea_alu_ea_reg_ax1rwe_DO_reg[10]/P0001  ;
  input \core_eu_ea_alu_ea_reg_ax1rwe_DO_reg[11]/P0001  ;
  input \core_eu_ea_alu_ea_reg_ax1rwe_DO_reg[12]/P0001  ;
  input \core_eu_ea_alu_ea_reg_ax1rwe_DO_reg[13]/P0001  ;
  input \core_eu_ea_alu_ea_reg_ax1rwe_DO_reg[14]/P0001  ;
  input \core_eu_ea_alu_ea_reg_ax1rwe_DO_reg[15]/P0001  ;
  input \core_eu_ea_alu_ea_reg_ax1rwe_DO_reg[1]/P0001  ;
  input \core_eu_ea_alu_ea_reg_ax1rwe_DO_reg[2]/P0001  ;
  input \core_eu_ea_alu_ea_reg_ax1rwe_DO_reg[3]/P0001  ;
  input \core_eu_ea_alu_ea_reg_ax1rwe_DO_reg[4]/P0001  ;
  input \core_eu_ea_alu_ea_reg_ax1rwe_DO_reg[5]/P0001  ;
  input \core_eu_ea_alu_ea_reg_ax1rwe_DO_reg[6]/P0001  ;
  input \core_eu_ea_alu_ea_reg_ax1rwe_DO_reg[7]/P0001  ;
  input \core_eu_ea_alu_ea_reg_ax1rwe_DO_reg[8]/P0001  ;
  input \core_eu_ea_alu_ea_reg_ax1rwe_DO_reg[9]/P0001  ;
  input \core_eu_ea_alu_ea_reg_ax1swe_DO_reg[0]/P0001  ;
  input \core_eu_ea_alu_ea_reg_ax1swe_DO_reg[10]/P0001  ;
  input \core_eu_ea_alu_ea_reg_ax1swe_DO_reg[11]/P0001  ;
  input \core_eu_ea_alu_ea_reg_ax1swe_DO_reg[12]/P0001  ;
  input \core_eu_ea_alu_ea_reg_ax1swe_DO_reg[13]/P0001  ;
  input \core_eu_ea_alu_ea_reg_ax1swe_DO_reg[14]/P0001  ;
  input \core_eu_ea_alu_ea_reg_ax1swe_DO_reg[15]/P0001  ;
  input \core_eu_ea_alu_ea_reg_ax1swe_DO_reg[1]/P0001  ;
  input \core_eu_ea_alu_ea_reg_ax1swe_DO_reg[2]/P0001  ;
  input \core_eu_ea_alu_ea_reg_ax1swe_DO_reg[3]/P0001  ;
  input \core_eu_ea_alu_ea_reg_ax1swe_DO_reg[4]/P0001  ;
  input \core_eu_ea_alu_ea_reg_ax1swe_DO_reg[5]/P0001  ;
  input \core_eu_ea_alu_ea_reg_ax1swe_DO_reg[6]/P0001  ;
  input \core_eu_ea_alu_ea_reg_ax1swe_DO_reg[7]/P0001  ;
  input \core_eu_ea_alu_ea_reg_ax1swe_DO_reg[8]/P0001  ;
  input \core_eu_ea_alu_ea_reg_ax1swe_DO_reg[9]/P0001  ;
  input \core_eu_ea_alu_ea_reg_ay0rwe_DO_reg[0]/P0001  ;
  input \core_eu_ea_alu_ea_reg_ay0rwe_DO_reg[10]/P0001  ;
  input \core_eu_ea_alu_ea_reg_ay0rwe_DO_reg[11]/P0001  ;
  input \core_eu_ea_alu_ea_reg_ay0rwe_DO_reg[12]/P0001  ;
  input \core_eu_ea_alu_ea_reg_ay0rwe_DO_reg[13]/P0001  ;
  input \core_eu_ea_alu_ea_reg_ay0rwe_DO_reg[14]/P0001  ;
  input \core_eu_ea_alu_ea_reg_ay0rwe_DO_reg[15]/P0001  ;
  input \core_eu_ea_alu_ea_reg_ay0rwe_DO_reg[1]/P0001  ;
  input \core_eu_ea_alu_ea_reg_ay0rwe_DO_reg[2]/P0001  ;
  input \core_eu_ea_alu_ea_reg_ay0rwe_DO_reg[3]/P0001  ;
  input \core_eu_ea_alu_ea_reg_ay0rwe_DO_reg[4]/P0001  ;
  input \core_eu_ea_alu_ea_reg_ay0rwe_DO_reg[5]/P0001  ;
  input \core_eu_ea_alu_ea_reg_ay0rwe_DO_reg[6]/P0001  ;
  input \core_eu_ea_alu_ea_reg_ay0rwe_DO_reg[7]/P0001  ;
  input \core_eu_ea_alu_ea_reg_ay0rwe_DO_reg[8]/P0001  ;
  input \core_eu_ea_alu_ea_reg_ay0rwe_DO_reg[9]/P0001  ;
  input \core_eu_ea_alu_ea_reg_ay0swe_DO_reg[0]/P0001  ;
  input \core_eu_ea_alu_ea_reg_ay0swe_DO_reg[10]/P0001  ;
  input \core_eu_ea_alu_ea_reg_ay0swe_DO_reg[11]/P0001  ;
  input \core_eu_ea_alu_ea_reg_ay0swe_DO_reg[12]/P0001  ;
  input \core_eu_ea_alu_ea_reg_ay0swe_DO_reg[13]/P0001  ;
  input \core_eu_ea_alu_ea_reg_ay0swe_DO_reg[14]/P0001  ;
  input \core_eu_ea_alu_ea_reg_ay0swe_DO_reg[15]/P0001  ;
  input \core_eu_ea_alu_ea_reg_ay0swe_DO_reg[1]/P0001  ;
  input \core_eu_ea_alu_ea_reg_ay0swe_DO_reg[2]/P0001  ;
  input \core_eu_ea_alu_ea_reg_ay0swe_DO_reg[3]/P0001  ;
  input \core_eu_ea_alu_ea_reg_ay0swe_DO_reg[4]/P0001  ;
  input \core_eu_ea_alu_ea_reg_ay0swe_DO_reg[5]/P0001  ;
  input \core_eu_ea_alu_ea_reg_ay0swe_DO_reg[6]/P0001  ;
  input \core_eu_ea_alu_ea_reg_ay0swe_DO_reg[7]/P0001  ;
  input \core_eu_ea_alu_ea_reg_ay0swe_DO_reg[8]/P0001  ;
  input \core_eu_ea_alu_ea_reg_ay0swe_DO_reg[9]/P0001  ;
  input \core_eu_ea_alu_ea_reg_ay1rwe_DO_reg[0]/P0001  ;
  input \core_eu_ea_alu_ea_reg_ay1rwe_DO_reg[10]/P0001  ;
  input \core_eu_ea_alu_ea_reg_ay1rwe_DO_reg[11]/P0001  ;
  input \core_eu_ea_alu_ea_reg_ay1rwe_DO_reg[12]/P0001  ;
  input \core_eu_ea_alu_ea_reg_ay1rwe_DO_reg[13]/P0001  ;
  input \core_eu_ea_alu_ea_reg_ay1rwe_DO_reg[14]/P0001  ;
  input \core_eu_ea_alu_ea_reg_ay1rwe_DO_reg[15]/P0001  ;
  input \core_eu_ea_alu_ea_reg_ay1rwe_DO_reg[1]/P0001  ;
  input \core_eu_ea_alu_ea_reg_ay1rwe_DO_reg[2]/P0001  ;
  input \core_eu_ea_alu_ea_reg_ay1rwe_DO_reg[3]/P0001  ;
  input \core_eu_ea_alu_ea_reg_ay1rwe_DO_reg[4]/P0001  ;
  input \core_eu_ea_alu_ea_reg_ay1rwe_DO_reg[5]/P0001  ;
  input \core_eu_ea_alu_ea_reg_ay1rwe_DO_reg[6]/P0001  ;
  input \core_eu_ea_alu_ea_reg_ay1rwe_DO_reg[7]/P0001  ;
  input \core_eu_ea_alu_ea_reg_ay1rwe_DO_reg[8]/P0001  ;
  input \core_eu_ea_alu_ea_reg_ay1rwe_DO_reg[9]/P0001  ;
  input \core_eu_ea_alu_ea_reg_ay1swe_DO_reg[0]/P0001  ;
  input \core_eu_ea_alu_ea_reg_ay1swe_DO_reg[10]/P0001  ;
  input \core_eu_ea_alu_ea_reg_ay1swe_DO_reg[11]/P0001  ;
  input \core_eu_ea_alu_ea_reg_ay1swe_DO_reg[12]/P0001  ;
  input \core_eu_ea_alu_ea_reg_ay1swe_DO_reg[13]/P0001  ;
  input \core_eu_ea_alu_ea_reg_ay1swe_DO_reg[14]/P0001  ;
  input \core_eu_ea_alu_ea_reg_ay1swe_DO_reg[15]/P0001  ;
  input \core_eu_ea_alu_ea_reg_ay1swe_DO_reg[1]/P0001  ;
  input \core_eu_ea_alu_ea_reg_ay1swe_DO_reg[2]/P0001  ;
  input \core_eu_ea_alu_ea_reg_ay1swe_DO_reg[3]/P0001  ;
  input \core_eu_ea_alu_ea_reg_ay1swe_DO_reg[4]/P0001  ;
  input \core_eu_ea_alu_ea_reg_ay1swe_DO_reg[5]/P0001  ;
  input \core_eu_ea_alu_ea_reg_ay1swe_DO_reg[6]/P0001  ;
  input \core_eu_ea_alu_ea_reg_ay1swe_DO_reg[7]/P0001  ;
  input \core_eu_ea_alu_ea_reg_ay1swe_DO_reg[8]/P0001  ;
  input \core_eu_ea_alu_ea_reg_ay1swe_DO_reg[9]/P0001  ;
  input \core_eu_ec_cun_AC_reg/P0001  ;
  input \core_eu_ec_cun_AN_reg/P0001  ;
  input \core_eu_ec_cun_AQ_reg/P0001  ;
  input \core_eu_ec_cun_AS_reg/P0001  ;
  input \core_eu_ec_cun_AV_reg/P0001  ;
  input \core_eu_ec_cun_AZ_reg/P0001  ;
  input \core_eu_ec_cun_COND_E_reg[0]/P0001  ;
  input \core_eu_ec_cun_COND_E_reg[1]/P0001  ;
  input \core_eu_ec_cun_COND_E_reg[2]/P0001  ;
  input \core_eu_ec_cun_COND_E_reg[3]/P0001  ;
  input \core_eu_ec_cun_MV_reg/P0000_reg_syn_2  ;
  input \core_eu_ec_cun_MVi_pre_C_reg/P0001  ;
  input \core_eu_ec_cun_SS_reg/P0001  ;
  input \core_eu_ec_cun_TERM_E_reg[0]/P0001  ;
  input \core_eu_ec_cun_TERM_E_reg[1]/P0001  ;
  input \core_eu_ec_cun_TERM_E_reg[2]/P0001  ;
  input \core_eu_ec_cun_TERM_E_reg[3]/P0001  ;
  input \core_eu_ec_cun_condOK_CE_reg/P0001  ;
  input \core_eu_ec_cun_mven_FFout_reg/NET0131  ;
  input \core_eu_ec_cun_termOK_CE_reg/P0001  ;
  input \core_eu_ec_cun_updateMV_C_reg/P0001  ;
  input \core_eu_em_mac_em_dec_emcorepi_DO_reg[0]/P0001  ;
  input \core_eu_em_mac_em_dec_emcorepi_DO_reg[10]/P0001  ;
  input \core_eu_em_mac_em_dec_emcorepi_DO_reg[1]/P0001  ;
  input \core_eu_em_mac_em_dec_emcorepi_DO_reg[2]/P0001  ;
  input \core_eu_em_mac_em_dec_emcorepi_DO_reg[3]/P0001  ;
  input \core_eu_em_mac_em_reg_Sq_E_reg/P0001  ;
  input \core_eu_em_mac_em_reg_mfrwe_DO_reg[0]/P0001  ;
  input \core_eu_em_mac_em_reg_mfrwe_DO_reg[10]/P0001  ;
  input \core_eu_em_mac_em_reg_mfrwe_DO_reg[11]/P0001  ;
  input \core_eu_em_mac_em_reg_mfrwe_DO_reg[12]/P0001  ;
  input \core_eu_em_mac_em_reg_mfrwe_DO_reg[13]/P0001  ;
  input \core_eu_em_mac_em_reg_mfrwe_DO_reg[14]/P0001  ;
  input \core_eu_em_mac_em_reg_mfrwe_DO_reg[15]/P0001  ;
  input \core_eu_em_mac_em_reg_mfrwe_DO_reg[1]/P0001  ;
  input \core_eu_em_mac_em_reg_mfrwe_DO_reg[2]/P0001  ;
  input \core_eu_em_mac_em_reg_mfrwe_DO_reg[3]/P0001  ;
  input \core_eu_em_mac_em_reg_mfrwe_DO_reg[4]/P0001  ;
  input \core_eu_em_mac_em_reg_mfrwe_DO_reg[5]/P0001  ;
  input \core_eu_em_mac_em_reg_mfrwe_DO_reg[6]/P0001  ;
  input \core_eu_em_mac_em_reg_mfrwe_DO_reg[7]/P0001  ;
  input \core_eu_em_mac_em_reg_mfrwe_DO_reg[8]/P0001  ;
  input \core_eu_em_mac_em_reg_mfrwe_DO_reg[9]/P0001  ;
  input \core_eu_em_mac_em_reg_mfswe_DO_reg[0]/P0001  ;
  input \core_eu_em_mac_em_reg_mfswe_DO_reg[10]/P0001  ;
  input \core_eu_em_mac_em_reg_mfswe_DO_reg[11]/P0001  ;
  input \core_eu_em_mac_em_reg_mfswe_DO_reg[12]/P0001  ;
  input \core_eu_em_mac_em_reg_mfswe_DO_reg[13]/P0001  ;
  input \core_eu_em_mac_em_reg_mfswe_DO_reg[14]/P0001  ;
  input \core_eu_em_mac_em_reg_mfswe_DO_reg[15]/P0001  ;
  input \core_eu_em_mac_em_reg_mfswe_DO_reg[1]/P0001  ;
  input \core_eu_em_mac_em_reg_mfswe_DO_reg[2]/P0001  ;
  input \core_eu_em_mac_em_reg_mfswe_DO_reg[3]/P0001  ;
  input \core_eu_em_mac_em_reg_mfswe_DO_reg[4]/P0001  ;
  input \core_eu_em_mac_em_reg_mfswe_DO_reg[5]/P0001  ;
  input \core_eu_em_mac_em_reg_mfswe_DO_reg[6]/P0001  ;
  input \core_eu_em_mac_em_reg_mfswe_DO_reg[7]/P0001  ;
  input \core_eu_em_mac_em_reg_mfswe_DO_reg[8]/P0001  ;
  input \core_eu_em_mac_em_reg_mfswe_DO_reg[9]/P0001  ;
  input \core_eu_em_mac_em_reg_mr0rwe_DO_reg[0]/P0001  ;
  input \core_eu_em_mac_em_reg_mr0rwe_DO_reg[10]/P0001  ;
  input \core_eu_em_mac_em_reg_mr0rwe_DO_reg[11]/P0001  ;
  input \core_eu_em_mac_em_reg_mr0rwe_DO_reg[12]/P0001  ;
  input \core_eu_em_mac_em_reg_mr0rwe_DO_reg[13]/P0001  ;
  input \core_eu_em_mac_em_reg_mr0rwe_DO_reg[14]/P0001  ;
  input \core_eu_em_mac_em_reg_mr0rwe_DO_reg[15]/P0001  ;
  input \core_eu_em_mac_em_reg_mr0rwe_DO_reg[1]/P0001  ;
  input \core_eu_em_mac_em_reg_mr0rwe_DO_reg[2]/P0001  ;
  input \core_eu_em_mac_em_reg_mr0rwe_DO_reg[3]/P0001  ;
  input \core_eu_em_mac_em_reg_mr0rwe_DO_reg[4]/P0001  ;
  input \core_eu_em_mac_em_reg_mr0rwe_DO_reg[5]/P0001  ;
  input \core_eu_em_mac_em_reg_mr0rwe_DO_reg[6]/P0001  ;
  input \core_eu_em_mac_em_reg_mr0rwe_DO_reg[7]/P0001  ;
  input \core_eu_em_mac_em_reg_mr0rwe_DO_reg[8]/P0001  ;
  input \core_eu_em_mac_em_reg_mr0rwe_DO_reg[9]/P0001  ;
  input \core_eu_em_mac_em_reg_mr0swe_DO_reg[0]/P0001  ;
  input \core_eu_em_mac_em_reg_mr0swe_DO_reg[10]/P0001  ;
  input \core_eu_em_mac_em_reg_mr0swe_DO_reg[11]/P0001  ;
  input \core_eu_em_mac_em_reg_mr0swe_DO_reg[12]/P0001  ;
  input \core_eu_em_mac_em_reg_mr0swe_DO_reg[13]/P0001  ;
  input \core_eu_em_mac_em_reg_mr0swe_DO_reg[14]/P0001  ;
  input \core_eu_em_mac_em_reg_mr0swe_DO_reg[15]/P0001  ;
  input \core_eu_em_mac_em_reg_mr0swe_DO_reg[1]/P0001  ;
  input \core_eu_em_mac_em_reg_mr0swe_DO_reg[2]/P0001  ;
  input \core_eu_em_mac_em_reg_mr0swe_DO_reg[3]/P0001  ;
  input \core_eu_em_mac_em_reg_mr0swe_DO_reg[4]/P0001  ;
  input \core_eu_em_mac_em_reg_mr0swe_DO_reg[5]/P0001  ;
  input \core_eu_em_mac_em_reg_mr0swe_DO_reg[6]/P0001  ;
  input \core_eu_em_mac_em_reg_mr0swe_DO_reg[7]/P0001  ;
  input \core_eu_em_mac_em_reg_mr0swe_DO_reg[8]/P0001  ;
  input \core_eu_em_mac_em_reg_mr0swe_DO_reg[9]/P0001  ;
  input \core_eu_em_mac_em_reg_mr1rwe_DO_reg[0]/P0001  ;
  input \core_eu_em_mac_em_reg_mr1rwe_DO_reg[10]/P0001  ;
  input \core_eu_em_mac_em_reg_mr1rwe_DO_reg[11]/P0001  ;
  input \core_eu_em_mac_em_reg_mr1rwe_DO_reg[12]/P0001  ;
  input \core_eu_em_mac_em_reg_mr1rwe_DO_reg[13]/P0001  ;
  input \core_eu_em_mac_em_reg_mr1rwe_DO_reg[14]/P0001  ;
  input \core_eu_em_mac_em_reg_mr1rwe_DO_reg[15]/P0001  ;
  input \core_eu_em_mac_em_reg_mr1rwe_DO_reg[1]/P0001  ;
  input \core_eu_em_mac_em_reg_mr1rwe_DO_reg[2]/P0001  ;
  input \core_eu_em_mac_em_reg_mr1rwe_DO_reg[3]/P0001  ;
  input \core_eu_em_mac_em_reg_mr1rwe_DO_reg[4]/P0001  ;
  input \core_eu_em_mac_em_reg_mr1rwe_DO_reg[5]/P0001  ;
  input \core_eu_em_mac_em_reg_mr1rwe_DO_reg[6]/P0001  ;
  input \core_eu_em_mac_em_reg_mr1rwe_DO_reg[7]/P0001  ;
  input \core_eu_em_mac_em_reg_mr1rwe_DO_reg[8]/P0001  ;
  input \core_eu_em_mac_em_reg_mr1rwe_DO_reg[9]/P0001  ;
  input \core_eu_em_mac_em_reg_mr1swe_DO_reg[0]/P0001  ;
  input \core_eu_em_mac_em_reg_mr1swe_DO_reg[10]/P0001  ;
  input \core_eu_em_mac_em_reg_mr1swe_DO_reg[11]/P0001  ;
  input \core_eu_em_mac_em_reg_mr1swe_DO_reg[12]/P0001  ;
  input \core_eu_em_mac_em_reg_mr1swe_DO_reg[13]/P0001  ;
  input \core_eu_em_mac_em_reg_mr1swe_DO_reg[14]/P0001  ;
  input \core_eu_em_mac_em_reg_mr1swe_DO_reg[15]/P0001  ;
  input \core_eu_em_mac_em_reg_mr1swe_DO_reg[1]/P0001  ;
  input \core_eu_em_mac_em_reg_mr1swe_DO_reg[2]/P0001  ;
  input \core_eu_em_mac_em_reg_mr1swe_DO_reg[3]/P0001  ;
  input \core_eu_em_mac_em_reg_mr1swe_DO_reg[4]/P0001  ;
  input \core_eu_em_mac_em_reg_mr1swe_DO_reg[5]/P0001  ;
  input \core_eu_em_mac_em_reg_mr1swe_DO_reg[6]/P0001  ;
  input \core_eu_em_mac_em_reg_mr1swe_DO_reg[7]/P0001  ;
  input \core_eu_em_mac_em_reg_mr1swe_DO_reg[8]/P0001  ;
  input \core_eu_em_mac_em_reg_mr1swe_DO_reg[9]/P0001  ;
  input \core_eu_em_mac_em_reg_mr2rwe_DO_reg[0]/P0001  ;
  input \core_eu_em_mac_em_reg_mr2rwe_DO_reg[1]/P0001  ;
  input \core_eu_em_mac_em_reg_mr2rwe_DO_reg[2]/P0001  ;
  input \core_eu_em_mac_em_reg_mr2rwe_DO_reg[3]/P0001  ;
  input \core_eu_em_mac_em_reg_mr2rwe_DO_reg[4]/P0001  ;
  input \core_eu_em_mac_em_reg_mr2rwe_DO_reg[5]/P0001  ;
  input \core_eu_em_mac_em_reg_mr2rwe_DO_reg[6]/P0001  ;
  input \core_eu_em_mac_em_reg_mr2rwe_DO_reg[7]/P0001  ;
  input \core_eu_em_mac_em_reg_mr2swe_DO_reg[0]/P0001  ;
  input \core_eu_em_mac_em_reg_mr2swe_DO_reg[1]/P0001  ;
  input \core_eu_em_mac_em_reg_mr2swe_DO_reg[2]/P0001  ;
  input \core_eu_em_mac_em_reg_mr2swe_DO_reg[3]/P0001  ;
  input \core_eu_em_mac_em_reg_mr2swe_DO_reg[4]/P0001  ;
  input \core_eu_em_mac_em_reg_mr2swe_DO_reg[5]/P0001  ;
  input \core_eu_em_mac_em_reg_mr2swe_DO_reg[6]/P0001  ;
  input \core_eu_em_mac_em_reg_mr2swe_DO_reg[7]/P0001  ;
  input \core_eu_em_mac_em_reg_mrovfwe_DO_reg[0]/P0001  ;
  input \core_eu_em_mac_em_reg_mrovfwe_DO_reg[1]/P0001  ;
  input \core_eu_em_mac_em_reg_mrovfwe_DO_reg[2]/P0001  ;
  input \core_eu_em_mac_em_reg_mrovfwe_DO_reg[3]/P0001  ;
  input \core_eu_em_mac_em_reg_mrovfwe_DO_reg[4]/P0001  ;
  input \core_eu_em_mac_em_reg_mrovfwe_DO_reg[5]/P0001  ;
  input \core_eu_em_mac_em_reg_mrovfwe_DO_reg[6]/P0001  ;
  input \core_eu_em_mac_em_reg_mrovfwe_DO_reg[7]/P0001  ;
  input \core_eu_em_mac_em_reg_mrovfwe_DO_reg[8]/P0001  ;
  input \core_eu_em_mac_em_reg_mx0rwe_DO_reg[0]/P0001  ;
  input \core_eu_em_mac_em_reg_mx0rwe_DO_reg[10]/P0001  ;
  input \core_eu_em_mac_em_reg_mx0rwe_DO_reg[11]/P0001  ;
  input \core_eu_em_mac_em_reg_mx0rwe_DO_reg[12]/P0001  ;
  input \core_eu_em_mac_em_reg_mx0rwe_DO_reg[13]/P0001  ;
  input \core_eu_em_mac_em_reg_mx0rwe_DO_reg[14]/P0001  ;
  input \core_eu_em_mac_em_reg_mx0rwe_DO_reg[15]/P0001  ;
  input \core_eu_em_mac_em_reg_mx0rwe_DO_reg[1]/P0001  ;
  input \core_eu_em_mac_em_reg_mx0rwe_DO_reg[2]/P0001  ;
  input \core_eu_em_mac_em_reg_mx0rwe_DO_reg[3]/P0001  ;
  input \core_eu_em_mac_em_reg_mx0rwe_DO_reg[4]/P0001  ;
  input \core_eu_em_mac_em_reg_mx0rwe_DO_reg[5]/P0001  ;
  input \core_eu_em_mac_em_reg_mx0rwe_DO_reg[6]/P0001  ;
  input \core_eu_em_mac_em_reg_mx0rwe_DO_reg[7]/P0001  ;
  input \core_eu_em_mac_em_reg_mx0rwe_DO_reg[8]/P0001  ;
  input \core_eu_em_mac_em_reg_mx0rwe_DO_reg[9]/P0001  ;
  input \core_eu_em_mac_em_reg_mx0swe_DO_reg[0]/P0001  ;
  input \core_eu_em_mac_em_reg_mx0swe_DO_reg[10]/P0001  ;
  input \core_eu_em_mac_em_reg_mx0swe_DO_reg[11]/P0001  ;
  input \core_eu_em_mac_em_reg_mx0swe_DO_reg[12]/P0001  ;
  input \core_eu_em_mac_em_reg_mx0swe_DO_reg[13]/P0001  ;
  input \core_eu_em_mac_em_reg_mx0swe_DO_reg[14]/P0001  ;
  input \core_eu_em_mac_em_reg_mx0swe_DO_reg[15]/P0001  ;
  input \core_eu_em_mac_em_reg_mx0swe_DO_reg[1]/P0001  ;
  input \core_eu_em_mac_em_reg_mx0swe_DO_reg[2]/P0001  ;
  input \core_eu_em_mac_em_reg_mx0swe_DO_reg[3]/P0001  ;
  input \core_eu_em_mac_em_reg_mx0swe_DO_reg[4]/P0001  ;
  input \core_eu_em_mac_em_reg_mx0swe_DO_reg[5]/P0001  ;
  input \core_eu_em_mac_em_reg_mx0swe_DO_reg[6]/P0001  ;
  input \core_eu_em_mac_em_reg_mx0swe_DO_reg[7]/P0001  ;
  input \core_eu_em_mac_em_reg_mx0swe_DO_reg[8]/P0001  ;
  input \core_eu_em_mac_em_reg_mx0swe_DO_reg[9]/P0001  ;
  input \core_eu_em_mac_em_reg_mx1rwe_DO_reg[0]/P0001  ;
  input \core_eu_em_mac_em_reg_mx1rwe_DO_reg[10]/P0001  ;
  input \core_eu_em_mac_em_reg_mx1rwe_DO_reg[11]/P0001  ;
  input \core_eu_em_mac_em_reg_mx1rwe_DO_reg[12]/P0001  ;
  input \core_eu_em_mac_em_reg_mx1rwe_DO_reg[13]/P0001  ;
  input \core_eu_em_mac_em_reg_mx1rwe_DO_reg[14]/P0001  ;
  input \core_eu_em_mac_em_reg_mx1rwe_DO_reg[15]/P0001  ;
  input \core_eu_em_mac_em_reg_mx1rwe_DO_reg[1]/P0001  ;
  input \core_eu_em_mac_em_reg_mx1rwe_DO_reg[2]/P0001  ;
  input \core_eu_em_mac_em_reg_mx1rwe_DO_reg[3]/P0001  ;
  input \core_eu_em_mac_em_reg_mx1rwe_DO_reg[4]/P0001  ;
  input \core_eu_em_mac_em_reg_mx1rwe_DO_reg[5]/P0001  ;
  input \core_eu_em_mac_em_reg_mx1rwe_DO_reg[6]/P0001  ;
  input \core_eu_em_mac_em_reg_mx1rwe_DO_reg[7]/P0001  ;
  input \core_eu_em_mac_em_reg_mx1rwe_DO_reg[8]/P0001  ;
  input \core_eu_em_mac_em_reg_mx1rwe_DO_reg[9]/P0001  ;
  input \core_eu_em_mac_em_reg_mx1swe_DO_reg[0]/P0001  ;
  input \core_eu_em_mac_em_reg_mx1swe_DO_reg[10]/P0001  ;
  input \core_eu_em_mac_em_reg_mx1swe_DO_reg[11]/P0001  ;
  input \core_eu_em_mac_em_reg_mx1swe_DO_reg[12]/P0001  ;
  input \core_eu_em_mac_em_reg_mx1swe_DO_reg[13]/P0001  ;
  input \core_eu_em_mac_em_reg_mx1swe_DO_reg[14]/P0001  ;
  input \core_eu_em_mac_em_reg_mx1swe_DO_reg[15]/P0001  ;
  input \core_eu_em_mac_em_reg_mx1swe_DO_reg[1]/P0001  ;
  input \core_eu_em_mac_em_reg_mx1swe_DO_reg[2]/P0001  ;
  input \core_eu_em_mac_em_reg_mx1swe_DO_reg[3]/P0001  ;
  input \core_eu_em_mac_em_reg_mx1swe_DO_reg[4]/P0001  ;
  input \core_eu_em_mac_em_reg_mx1swe_DO_reg[5]/P0001  ;
  input \core_eu_em_mac_em_reg_mx1swe_DO_reg[6]/P0001  ;
  input \core_eu_em_mac_em_reg_mx1swe_DO_reg[7]/P0001  ;
  input \core_eu_em_mac_em_reg_mx1swe_DO_reg[8]/P0001  ;
  input \core_eu_em_mac_em_reg_mx1swe_DO_reg[9]/P0001  ;
  input \core_eu_em_mac_em_reg_mxopwe_DO_reg[0]/P0001  ;
  input \core_eu_em_mac_em_reg_mxopwe_DO_reg[10]/P0001  ;
  input \core_eu_em_mac_em_reg_mxopwe_DO_reg[11]/P0001  ;
  input \core_eu_em_mac_em_reg_mxopwe_DO_reg[12]/P0001  ;
  input \core_eu_em_mac_em_reg_mxopwe_DO_reg[13]/P0001  ;
  input \core_eu_em_mac_em_reg_mxopwe_DO_reg[14]/P0001  ;
  input \core_eu_em_mac_em_reg_mxopwe_DO_reg[15]/P0001  ;
  input \core_eu_em_mac_em_reg_mxopwe_DO_reg[1]/P0001  ;
  input \core_eu_em_mac_em_reg_mxopwe_DO_reg[2]/P0001  ;
  input \core_eu_em_mac_em_reg_mxopwe_DO_reg[3]/P0001  ;
  input \core_eu_em_mac_em_reg_mxopwe_DO_reg[4]/P0001  ;
  input \core_eu_em_mac_em_reg_mxopwe_DO_reg[5]/P0001  ;
  input \core_eu_em_mac_em_reg_mxopwe_DO_reg[6]/P0001  ;
  input \core_eu_em_mac_em_reg_mxopwe_DO_reg[7]/P0001  ;
  input \core_eu_em_mac_em_reg_mxopwe_DO_reg[8]/P0001  ;
  input \core_eu_em_mac_em_reg_mxopwe_DO_reg[9]/P0001  ;
  input \core_eu_em_mac_em_reg_my0rwe_DO_reg[0]/P0001  ;
  input \core_eu_em_mac_em_reg_my0rwe_DO_reg[10]/P0001  ;
  input \core_eu_em_mac_em_reg_my0rwe_DO_reg[11]/P0001  ;
  input \core_eu_em_mac_em_reg_my0rwe_DO_reg[12]/P0001  ;
  input \core_eu_em_mac_em_reg_my0rwe_DO_reg[13]/P0001  ;
  input \core_eu_em_mac_em_reg_my0rwe_DO_reg[14]/P0001  ;
  input \core_eu_em_mac_em_reg_my0rwe_DO_reg[15]/P0001  ;
  input \core_eu_em_mac_em_reg_my0rwe_DO_reg[1]/P0001  ;
  input \core_eu_em_mac_em_reg_my0rwe_DO_reg[2]/P0001  ;
  input \core_eu_em_mac_em_reg_my0rwe_DO_reg[3]/P0001  ;
  input \core_eu_em_mac_em_reg_my0rwe_DO_reg[4]/P0001  ;
  input \core_eu_em_mac_em_reg_my0rwe_DO_reg[5]/P0001  ;
  input \core_eu_em_mac_em_reg_my0rwe_DO_reg[6]/P0001  ;
  input \core_eu_em_mac_em_reg_my0rwe_DO_reg[7]/P0001  ;
  input \core_eu_em_mac_em_reg_my0rwe_DO_reg[8]/P0001  ;
  input \core_eu_em_mac_em_reg_my0rwe_DO_reg[9]/P0001  ;
  input \core_eu_em_mac_em_reg_my0swe_DO_reg[0]/P0001  ;
  input \core_eu_em_mac_em_reg_my0swe_DO_reg[10]/P0001  ;
  input \core_eu_em_mac_em_reg_my0swe_DO_reg[11]/P0001  ;
  input \core_eu_em_mac_em_reg_my0swe_DO_reg[12]/P0001  ;
  input \core_eu_em_mac_em_reg_my0swe_DO_reg[13]/P0001  ;
  input \core_eu_em_mac_em_reg_my0swe_DO_reg[14]/P0001  ;
  input \core_eu_em_mac_em_reg_my0swe_DO_reg[15]/P0001  ;
  input \core_eu_em_mac_em_reg_my0swe_DO_reg[1]/P0001  ;
  input \core_eu_em_mac_em_reg_my0swe_DO_reg[2]/P0001  ;
  input \core_eu_em_mac_em_reg_my0swe_DO_reg[3]/P0001  ;
  input \core_eu_em_mac_em_reg_my0swe_DO_reg[4]/P0001  ;
  input \core_eu_em_mac_em_reg_my0swe_DO_reg[5]/P0001  ;
  input \core_eu_em_mac_em_reg_my0swe_DO_reg[6]/P0001  ;
  input \core_eu_em_mac_em_reg_my0swe_DO_reg[7]/P0001  ;
  input \core_eu_em_mac_em_reg_my0swe_DO_reg[8]/P0001  ;
  input \core_eu_em_mac_em_reg_my0swe_DO_reg[9]/P0001  ;
  input \core_eu_em_mac_em_reg_my1rwe_DO_reg[0]/P0001  ;
  input \core_eu_em_mac_em_reg_my1rwe_DO_reg[10]/P0001  ;
  input \core_eu_em_mac_em_reg_my1rwe_DO_reg[11]/P0001  ;
  input \core_eu_em_mac_em_reg_my1rwe_DO_reg[12]/P0001  ;
  input \core_eu_em_mac_em_reg_my1rwe_DO_reg[13]/P0001  ;
  input \core_eu_em_mac_em_reg_my1rwe_DO_reg[14]/P0001  ;
  input \core_eu_em_mac_em_reg_my1rwe_DO_reg[15]/P0001  ;
  input \core_eu_em_mac_em_reg_my1rwe_DO_reg[1]/P0001  ;
  input \core_eu_em_mac_em_reg_my1rwe_DO_reg[2]/P0001  ;
  input \core_eu_em_mac_em_reg_my1rwe_DO_reg[3]/P0001  ;
  input \core_eu_em_mac_em_reg_my1rwe_DO_reg[4]/P0001  ;
  input \core_eu_em_mac_em_reg_my1rwe_DO_reg[5]/P0001  ;
  input \core_eu_em_mac_em_reg_my1rwe_DO_reg[6]/P0001  ;
  input \core_eu_em_mac_em_reg_my1rwe_DO_reg[7]/P0001  ;
  input \core_eu_em_mac_em_reg_my1rwe_DO_reg[8]/P0001  ;
  input \core_eu_em_mac_em_reg_my1rwe_DO_reg[9]/P0001  ;
  input \core_eu_em_mac_em_reg_my1swe_DO_reg[0]/P0001  ;
  input \core_eu_em_mac_em_reg_my1swe_DO_reg[10]/P0001  ;
  input \core_eu_em_mac_em_reg_my1swe_DO_reg[11]/P0001  ;
  input \core_eu_em_mac_em_reg_my1swe_DO_reg[12]/P0001  ;
  input \core_eu_em_mac_em_reg_my1swe_DO_reg[13]/P0001  ;
  input \core_eu_em_mac_em_reg_my1swe_DO_reg[14]/P0001  ;
  input \core_eu_em_mac_em_reg_my1swe_DO_reg[15]/P0001  ;
  input \core_eu_em_mac_em_reg_my1swe_DO_reg[1]/P0001  ;
  input \core_eu_em_mac_em_reg_my1swe_DO_reg[2]/P0001  ;
  input \core_eu_em_mac_em_reg_my1swe_DO_reg[3]/P0001  ;
  input \core_eu_em_mac_em_reg_my1swe_DO_reg[4]/P0001  ;
  input \core_eu_em_mac_em_reg_my1swe_DO_reg[5]/P0001  ;
  input \core_eu_em_mac_em_reg_my1swe_DO_reg[6]/P0001  ;
  input \core_eu_em_mac_em_reg_my1swe_DO_reg[7]/P0001  ;
  input \core_eu_em_mac_em_reg_my1swe_DO_reg[8]/P0001  ;
  input \core_eu_em_mac_em_reg_my1swe_DO_reg[9]/P0001  ;
  input \core_eu_em_mac_em_reg_myopwe_DO_reg[0]/P0001  ;
  input \core_eu_em_mac_em_reg_myopwe_DO_reg[10]/P0001  ;
  input \core_eu_em_mac_em_reg_myopwe_DO_reg[11]/P0001  ;
  input \core_eu_em_mac_em_reg_myopwe_DO_reg[12]/P0001  ;
  input \core_eu_em_mac_em_reg_myopwe_DO_reg[13]/P0001  ;
  input \core_eu_em_mac_em_reg_myopwe_DO_reg[14]/P0001  ;
  input \core_eu_em_mac_em_reg_myopwe_DO_reg[15]/P0001  ;
  input \core_eu_em_mac_em_reg_myopwe_DO_reg[1]/P0001  ;
  input \core_eu_em_mac_em_reg_myopwe_DO_reg[2]/P0001  ;
  input \core_eu_em_mac_em_reg_myopwe_DO_reg[3]/P0001  ;
  input \core_eu_em_mac_em_reg_myopwe_DO_reg[4]/P0001  ;
  input \core_eu_em_mac_em_reg_myopwe_DO_reg[5]/P0001  ;
  input \core_eu_em_mac_em_reg_myopwe_DO_reg[6]/P0001  ;
  input \core_eu_em_mac_em_reg_myopwe_DO_reg[7]/P0001  ;
  input \core_eu_em_mac_em_reg_myopwe_DO_reg[8]/P0001  ;
  input \core_eu_em_mac_em_reg_myopwe_DO_reg[9]/P0001  ;
  input \core_eu_em_mac_em_reg_s0_reg/P0000_reg_syn_2  ;
  input \core_eu_em_mac_em_reg_s1_reg/P0000_reg_syn_2  ;
  input \core_eu_em_mac_em_reg_s2_reg/P0000_reg_syn_2  ;
  input \core_eu_es_sht_es_reg_SBr_reg[0]/P0001  ;
  input \core_eu_es_sht_es_reg_SBr_reg[1]/P0001  ;
  input \core_eu_es_sht_es_reg_SBr_reg[2]/P0001  ;
  input \core_eu_es_sht_es_reg_SBr_reg[3]/P0001  ;
  input \core_eu_es_sht_es_reg_SBr_reg[4]/P0001  ;
  input \core_eu_es_sht_es_reg_SBs_reg[0]/P0001  ;
  input \core_eu_es_sht_es_reg_SBs_reg[1]/P0001  ;
  input \core_eu_es_sht_es_reg_SBs_reg[2]/P0001  ;
  input \core_eu_es_sht_es_reg_SBs_reg[3]/P0001  ;
  input \core_eu_es_sht_es_reg_SBs_reg[4]/P0001  ;
  input \core_eu_es_sht_es_reg_serwe_DO_reg[0]/P0001  ;
  input \core_eu_es_sht_es_reg_serwe_DO_reg[1]/P0001  ;
  input \core_eu_es_sht_es_reg_serwe_DO_reg[2]/P0001  ;
  input \core_eu_es_sht_es_reg_serwe_DO_reg[3]/P0001  ;
  input \core_eu_es_sht_es_reg_serwe_DO_reg[4]/P0001  ;
  input \core_eu_es_sht_es_reg_serwe_DO_reg[5]/P0001  ;
  input \core_eu_es_sht_es_reg_serwe_DO_reg[6]/P0001  ;
  input \core_eu_es_sht_es_reg_serwe_DO_reg[7]/P0001  ;
  input \core_eu_es_sht_es_reg_seswe_DO_reg[0]/P0001  ;
  input \core_eu_es_sht_es_reg_seswe_DO_reg[1]/P0001  ;
  input \core_eu_es_sht_es_reg_seswe_DO_reg[2]/P0001  ;
  input \core_eu_es_sht_es_reg_seswe_DO_reg[3]/P0001  ;
  input \core_eu_es_sht_es_reg_seswe_DO_reg[4]/P0001  ;
  input \core_eu_es_sht_es_reg_seswe_DO_reg[5]/P0001  ;
  input \core_eu_es_sht_es_reg_seswe_DO_reg[6]/P0001  ;
  input \core_eu_es_sht_es_reg_seswe_DO_reg[7]/P0001  ;
  input \core_eu_es_sht_es_reg_sirwe_DO_reg[0]/P0001  ;
  input \core_eu_es_sht_es_reg_sirwe_DO_reg[10]/P0001  ;
  input \core_eu_es_sht_es_reg_sirwe_DO_reg[11]/P0001  ;
  input \core_eu_es_sht_es_reg_sirwe_DO_reg[12]/P0001  ;
  input \core_eu_es_sht_es_reg_sirwe_DO_reg[13]/P0001  ;
  input \core_eu_es_sht_es_reg_sirwe_DO_reg[14]/P0001  ;
  input \core_eu_es_sht_es_reg_sirwe_DO_reg[15]/P0001  ;
  input \core_eu_es_sht_es_reg_sirwe_DO_reg[1]/P0001  ;
  input \core_eu_es_sht_es_reg_sirwe_DO_reg[2]/P0001  ;
  input \core_eu_es_sht_es_reg_sirwe_DO_reg[3]/P0001  ;
  input \core_eu_es_sht_es_reg_sirwe_DO_reg[4]/P0001  ;
  input \core_eu_es_sht_es_reg_sirwe_DO_reg[5]/P0001  ;
  input \core_eu_es_sht_es_reg_sirwe_DO_reg[6]/P0001  ;
  input \core_eu_es_sht_es_reg_sirwe_DO_reg[7]/P0001  ;
  input \core_eu_es_sht_es_reg_sirwe_DO_reg[8]/P0001  ;
  input \core_eu_es_sht_es_reg_sirwe_DO_reg[9]/P0001  ;
  input \core_eu_es_sht_es_reg_siswe_DO_reg[0]/P0001  ;
  input \core_eu_es_sht_es_reg_siswe_DO_reg[10]/P0001  ;
  input \core_eu_es_sht_es_reg_siswe_DO_reg[11]/P0001  ;
  input \core_eu_es_sht_es_reg_siswe_DO_reg[12]/P0001  ;
  input \core_eu_es_sht_es_reg_siswe_DO_reg[13]/P0001  ;
  input \core_eu_es_sht_es_reg_siswe_DO_reg[14]/P0001  ;
  input \core_eu_es_sht_es_reg_siswe_DO_reg[15]/P0001  ;
  input \core_eu_es_sht_es_reg_siswe_DO_reg[1]/P0001  ;
  input \core_eu_es_sht_es_reg_siswe_DO_reg[2]/P0001  ;
  input \core_eu_es_sht_es_reg_siswe_DO_reg[3]/P0001  ;
  input \core_eu_es_sht_es_reg_siswe_DO_reg[4]/P0001  ;
  input \core_eu_es_sht_es_reg_siswe_DO_reg[5]/P0001  ;
  input \core_eu_es_sht_es_reg_siswe_DO_reg[6]/P0001  ;
  input \core_eu_es_sht_es_reg_siswe_DO_reg[7]/P0001  ;
  input \core_eu_es_sht_es_reg_siswe_DO_reg[8]/P0001  ;
  input \core_eu_es_sht_es_reg_siswe_DO_reg[9]/P0001  ;
  input \core_eu_es_sht_es_reg_sr0rwe_DO_reg[0]/P0001  ;
  input \core_eu_es_sht_es_reg_sr0rwe_DO_reg[10]/P0001  ;
  input \core_eu_es_sht_es_reg_sr0rwe_DO_reg[11]/P0001  ;
  input \core_eu_es_sht_es_reg_sr0rwe_DO_reg[12]/P0001  ;
  input \core_eu_es_sht_es_reg_sr0rwe_DO_reg[13]/P0001  ;
  input \core_eu_es_sht_es_reg_sr0rwe_DO_reg[14]/P0001  ;
  input \core_eu_es_sht_es_reg_sr0rwe_DO_reg[15]/P0001  ;
  input \core_eu_es_sht_es_reg_sr0rwe_DO_reg[1]/P0001  ;
  input \core_eu_es_sht_es_reg_sr0rwe_DO_reg[2]/P0001  ;
  input \core_eu_es_sht_es_reg_sr0rwe_DO_reg[3]/P0001  ;
  input \core_eu_es_sht_es_reg_sr0rwe_DO_reg[4]/P0001  ;
  input \core_eu_es_sht_es_reg_sr0rwe_DO_reg[5]/P0001  ;
  input \core_eu_es_sht_es_reg_sr0rwe_DO_reg[6]/P0001  ;
  input \core_eu_es_sht_es_reg_sr0rwe_DO_reg[7]/P0001  ;
  input \core_eu_es_sht_es_reg_sr0rwe_DO_reg[8]/P0001  ;
  input \core_eu_es_sht_es_reg_sr0rwe_DO_reg[9]/P0001  ;
  input \core_eu_es_sht_es_reg_sr0swe_DO_reg[0]/P0001  ;
  input \core_eu_es_sht_es_reg_sr0swe_DO_reg[10]/P0001  ;
  input \core_eu_es_sht_es_reg_sr0swe_DO_reg[11]/P0001  ;
  input \core_eu_es_sht_es_reg_sr0swe_DO_reg[12]/P0001  ;
  input \core_eu_es_sht_es_reg_sr0swe_DO_reg[13]/P0001  ;
  input \core_eu_es_sht_es_reg_sr0swe_DO_reg[14]/P0001  ;
  input \core_eu_es_sht_es_reg_sr0swe_DO_reg[15]/P0001  ;
  input \core_eu_es_sht_es_reg_sr0swe_DO_reg[1]/P0001  ;
  input \core_eu_es_sht_es_reg_sr0swe_DO_reg[2]/P0001  ;
  input \core_eu_es_sht_es_reg_sr0swe_DO_reg[3]/P0001  ;
  input \core_eu_es_sht_es_reg_sr0swe_DO_reg[4]/P0001  ;
  input \core_eu_es_sht_es_reg_sr0swe_DO_reg[5]/P0001  ;
  input \core_eu_es_sht_es_reg_sr0swe_DO_reg[6]/P0001  ;
  input \core_eu_es_sht_es_reg_sr0swe_DO_reg[7]/P0001  ;
  input \core_eu_es_sht_es_reg_sr0swe_DO_reg[8]/P0001  ;
  input \core_eu_es_sht_es_reg_sr0swe_DO_reg[9]/P0001  ;
  input \core_eu_es_sht_es_reg_sr1rwe_DO_reg[0]/P0001  ;
  input \core_eu_es_sht_es_reg_sr1rwe_DO_reg[10]/P0001  ;
  input \core_eu_es_sht_es_reg_sr1rwe_DO_reg[11]/P0001  ;
  input \core_eu_es_sht_es_reg_sr1rwe_DO_reg[12]/P0001  ;
  input \core_eu_es_sht_es_reg_sr1rwe_DO_reg[13]/P0001  ;
  input \core_eu_es_sht_es_reg_sr1rwe_DO_reg[14]/P0001  ;
  input \core_eu_es_sht_es_reg_sr1rwe_DO_reg[15]/P0001  ;
  input \core_eu_es_sht_es_reg_sr1rwe_DO_reg[1]/P0001  ;
  input \core_eu_es_sht_es_reg_sr1rwe_DO_reg[2]/P0001  ;
  input \core_eu_es_sht_es_reg_sr1rwe_DO_reg[3]/P0001  ;
  input \core_eu_es_sht_es_reg_sr1rwe_DO_reg[4]/P0001  ;
  input \core_eu_es_sht_es_reg_sr1rwe_DO_reg[5]/P0001  ;
  input \core_eu_es_sht_es_reg_sr1rwe_DO_reg[6]/P0001  ;
  input \core_eu_es_sht_es_reg_sr1rwe_DO_reg[7]/P0001  ;
  input \core_eu_es_sht_es_reg_sr1rwe_DO_reg[8]/P0001  ;
  input \core_eu_es_sht_es_reg_sr1rwe_DO_reg[9]/P0001  ;
  input \core_eu_es_sht_es_reg_sr1swe_DO_reg[0]/P0001  ;
  input \core_eu_es_sht_es_reg_sr1swe_DO_reg[10]/P0001  ;
  input \core_eu_es_sht_es_reg_sr1swe_DO_reg[11]/P0001  ;
  input \core_eu_es_sht_es_reg_sr1swe_DO_reg[12]/P0001  ;
  input \core_eu_es_sht_es_reg_sr1swe_DO_reg[13]/P0001  ;
  input \core_eu_es_sht_es_reg_sr1swe_DO_reg[14]/P0001  ;
  input \core_eu_es_sht_es_reg_sr1swe_DO_reg[15]/P0001  ;
  input \core_eu_es_sht_es_reg_sr1swe_DO_reg[1]/P0001  ;
  input \core_eu_es_sht_es_reg_sr1swe_DO_reg[2]/P0001  ;
  input \core_eu_es_sht_es_reg_sr1swe_DO_reg[3]/P0001  ;
  input \core_eu_es_sht_es_reg_sr1swe_DO_reg[4]/P0001  ;
  input \core_eu_es_sht_es_reg_sr1swe_DO_reg[5]/P0001  ;
  input \core_eu_es_sht_es_reg_sr1swe_DO_reg[6]/P0001  ;
  input \core_eu_es_sht_es_reg_sr1swe_DO_reg[7]/P0001  ;
  input \core_eu_es_sht_es_reg_sr1swe_DO_reg[8]/P0001  ;
  input \core_eu_es_sht_es_reg_sr1swe_DO_reg[9]/P0001  ;
  input \emc_DMDoe_reg/NET0131  ;
  input \emc_DMDreg_reg[0]/P0001  ;
  input \emc_DMDreg_reg[10]/P0001  ;
  input \emc_DMDreg_reg[11]/P0001  ;
  input \emc_DMDreg_reg[12]/P0001  ;
  input \emc_DMDreg_reg[13]/P0001  ;
  input \emc_DMDreg_reg[14]/P0001  ;
  input \emc_DMDreg_reg[15]/P0001  ;
  input \emc_DMDreg_reg[1]/P0001  ;
  input \emc_DMDreg_reg[2]/P0001  ;
  input \emc_DMDreg_reg[3]/P0001  ;
  input \emc_DMDreg_reg[4]/P0001  ;
  input \emc_DMDreg_reg[5]/P0001  ;
  input \emc_DMDreg_reg[6]/P0001  ;
  input \emc_DMDreg_reg[7]/P0001  ;
  input \emc_DMDreg_reg[8]/P0001  ;
  input \emc_DMDreg_reg[9]/P0001  ;
  input \emc_DMcst_reg/NET0131  ;
  input \emc_ECMA_reg[0]/P0001  ;
  input \emc_ECMA_reg[10]/P0001  ;
  input \emc_ECMA_reg[11]/P0001  ;
  input \emc_ECMA_reg[12]/P0001  ;
  input \emc_ECMA_reg[1]/P0001  ;
  input \emc_ECMA_reg[2]/P0001  ;
  input \emc_ECMA_reg[3]/P0001  ;
  input \emc_ECMA_reg[4]/P0001  ;
  input \emc_ECMA_reg[5]/P0001  ;
  input \emc_ECMA_reg[6]/P0001  ;
  input \emc_ECMA_reg[7]/P0001  ;
  input \emc_ECMA_reg[8]/P0001  ;
  input \emc_ECMA_reg[9]/P0001  ;
  input \emc_ECMDreg_reg[0]/P0001  ;
  input \emc_ECMDreg_reg[10]/P0001  ;
  input \emc_ECMDreg_reg[11]/P0001  ;
  input \emc_ECMDreg_reg[12]/P0001  ;
  input \emc_ECMDreg_reg[13]/P0001  ;
  input \emc_ECMDreg_reg[14]/P0001  ;
  input \emc_ECMDreg_reg[15]/P0001  ;
  input \emc_ECMDreg_reg[16]/P0001  ;
  input \emc_ECMDreg_reg[17]/P0001  ;
  input \emc_ECMDreg_reg[18]/P0001  ;
  input \emc_ECMDreg_reg[19]/P0001  ;
  input \emc_ECMDreg_reg[1]/P0001  ;
  input \emc_ECMDreg_reg[20]/P0001  ;
  input \emc_ECMDreg_reg[21]/P0001  ;
  input \emc_ECMDreg_reg[22]/P0001  ;
  input \emc_ECMDreg_reg[23]/P0001  ;
  input \emc_ECMDreg_reg[2]/P0001  ;
  input \emc_ECMDreg_reg[3]/P0001  ;
  input \emc_ECMDreg_reg[4]/P0001  ;
  input \emc_ECMDreg_reg[5]/P0001  ;
  input \emc_ECMDreg_reg[6]/P0001  ;
  input \emc_ECMDreg_reg[7]/P0001  ;
  input \emc_ECMDreg_reg[8]/P0001  ;
  input \emc_ECMDreg_reg[9]/P0001  ;
  input \emc_ECMcs_reg/NET0131  ;
  input \emc_ECS_reg[0]/NET0131  ;
  input \emc_ECS_reg[1]/NET0131  ;
  input \emc_ECS_reg[2]/NET0131  ;
  input \emc_ECS_reg[3]/NET0131  ;
  input \emc_ED_oei_reg/P0001  ;
  input \emc_EXTC_Eg_syn_reg/P0001  ;
  input \emc_IOcst_reg/NET0131  ;
  input \emc_PMDoe_reg/NET0131  ;
  input \emc_PMDreg_reg[0]/P0001  ;
  input \emc_PMDreg_reg[10]/P0001  ;
  input \emc_PMDreg_reg[11]/P0001  ;
  input \emc_PMDreg_reg[12]/P0001  ;
  input \emc_PMDreg_reg[13]/P0001  ;
  input \emc_PMDreg_reg[14]/P0001  ;
  input \emc_PMDreg_reg[15]/P0001  ;
  input \emc_PMDreg_reg[1]/P0001  ;
  input \emc_PMDreg_reg[2]/P0001  ;
  input \emc_PMDreg_reg[3]/P0001  ;
  input \emc_PMDreg_reg[4]/P0001  ;
  input \emc_PMDreg_reg[5]/P0001  ;
  input \emc_PMDreg_reg[6]/P0001  ;
  input \emc_PMDreg_reg[7]/P0001  ;
  input \emc_PMDreg_reg[8]/P0001  ;
  input \emc_PMDreg_reg[9]/P0001  ;
  input \emc_PMcst_reg/NET0131  ;
  input \emc_RWcnt_reg[0]/P0001  ;
  input \emc_RWcnt_reg[1]/P0001  ;
  input \emc_RWcnt_reg[2]/P0001  ;
  input \emc_RWcnt_reg[3]/P0001  ;
  input \emc_RWcnt_reg[4]/P0001  ;
  input \emc_RWcnt_reg[5]/P0001  ;
  input \emc_WRn_h_reg/P0001  ;
  input \emc_WSCRext_reg_DO_reg[0]/NET0131  ;
  input \emc_WSCRext_reg_DO_reg[1]/NET0131  ;
  input \emc_WSCRext_reg_DO_reg[2]/NET0131  ;
  input \emc_WSCRext_reg_DO_reg[3]/NET0131  ;
  input \emc_WSCRext_reg_DO_reg[4]/NET0131  ;
  input \emc_WSCRext_reg_DO_reg[5]/NET0131  ;
  input \emc_WSCRext_reg_DO_reg[6]/NET0131  ;
  input \emc_WSCRext_reg_DO_reg[7]/NET0131  ;
  input \emc_WSCRreg_DO_reg[0]/NET0131  ;
  input \emc_WSCRreg_DO_reg[10]/NET0131  ;
  input \emc_WSCRreg_DO_reg[11]/NET0131  ;
  input \emc_WSCRreg_DO_reg[12]/NET0131  ;
  input \emc_WSCRreg_DO_reg[13]/NET0131  ;
  input \emc_WSCRreg_DO_reg[14]/NET0131  ;
  input \emc_WSCRreg_DO_reg[1]/NET0131  ;
  input \emc_WSCRreg_DO_reg[2]/NET0131  ;
  input \emc_WSCRreg_DO_reg[3]/NET0131  ;
  input \emc_WSCRreg_DO_reg[4]/NET0131  ;
  input \emc_WSCRreg_DO_reg[5]/NET0131  ;
  input \emc_WSCRreg_DO_reg[6]/NET0131  ;
  input \emc_WSCRreg_DO_reg[7]/NET0131  ;
  input \emc_WSCRreg_DO_reg[8]/NET0131  ;
  input \emc_WSCRreg_DO_reg[9]/NET0131  ;
  input \emc_eRDY_reg/NET0131  ;
  input \emc_selDMDi_reg/P0001  ;
  input \emc_selPMDi_reg/P0001  ;
  input \idma_CM_oe_reg/P0001  ;
  input \idma_CMo_oe0_reg/P0001  ;
  input \idma_CMo_oe1_reg/P0001  ;
  input \idma_CMo_oe2_reg/P0001  ;
  input \idma_CMo_oe3_reg/P0001  ;
  input \idma_CMo_oe4_reg/P0001  ;
  input \idma_CMo_oe5_reg/P0001  ;
  input \idma_CMo_oe6_reg/P0001  ;
  input \idma_CMo_oe7_reg/P0001  ;
  input \idma_DCTL_reg[0]/NET0131  ;
  input \idma_DCTL_reg[10]/NET0131  ;
  input \idma_DCTL_reg[11]/NET0131  ;
  input \idma_DCTL_reg[12]/NET0131  ;
  input \idma_DCTL_reg[13]/NET0131  ;
  input \idma_DCTL_reg[14]/NET0131  ;
  input \idma_DCTL_reg[1]/NET0131  ;
  input \idma_DCTL_reg[2]/NET0131  ;
  input \idma_DCTL_reg[3]/NET0131  ;
  input \idma_DCTL_reg[4]/NET0131  ;
  input \idma_DCTL_reg[5]/NET0131  ;
  input \idma_DCTL_reg[6]/NET0131  ;
  input \idma_DCTL_reg[7]/NET0131  ;
  input \idma_DCTL_reg[8]/NET0131  ;
  input \idma_DCTL_reg[9]/NET0131  ;
  input \idma_DOVL_reg[0]/NET0131  ;
  input \idma_DOVL_reg[10]/NET0131  ;
  input \idma_DOVL_reg[11]/NET0131  ;
  input \idma_DOVL_reg[1]/NET0131  ;
  input \idma_DOVL_reg[2]/NET0131  ;
  input \idma_DOVL_reg[3]/NET0131  ;
  input \idma_DOVL_reg[4]/NET0131  ;
  input \idma_DOVL_reg[5]/NET0131  ;
  input \idma_DOVL_reg[6]/NET0131  ;
  input \idma_DOVL_reg[7]/NET0131  ;
  input \idma_DOVL_reg[8]/NET0131  ;
  input \idma_DOVL_reg[9]/NET0131  ;
  input \idma_DSreq_reg/NET0131  ;
  input \idma_DTMP_H_reg[0]/P0001  ;
  input \idma_DTMP_H_reg[10]/P0001  ;
  input \idma_DTMP_H_reg[11]/P0001  ;
  input \idma_DTMP_H_reg[12]/P0001  ;
  input \idma_DTMP_H_reg[13]/P0001  ;
  input \idma_DTMP_H_reg[14]/P0001  ;
  input \idma_DTMP_H_reg[15]/P0001  ;
  input \idma_DTMP_H_reg[1]/P0001  ;
  input \idma_DTMP_H_reg[2]/P0001  ;
  input \idma_DTMP_H_reg[3]/P0001  ;
  input \idma_DTMP_H_reg[4]/P0001  ;
  input \idma_DTMP_H_reg[5]/P0001  ;
  input \idma_DTMP_H_reg[6]/P0001  ;
  input \idma_DTMP_H_reg[7]/P0001  ;
  input \idma_DTMP_H_reg[8]/P0001  ;
  input \idma_DTMP_H_reg[9]/P0001  ;
  input \idma_DTMP_L_reg[0]/P0001  ;
  input \idma_DTMP_L_reg[1]/P0001  ;
  input \idma_DTMP_L_reg[2]/P0001  ;
  input \idma_DTMP_L_reg[3]/P0001  ;
  input \idma_DTMP_L_reg[4]/P0001  ;
  input \idma_DTMP_L_reg[5]/P0001  ;
  input \idma_DTMP_L_reg[6]/P0001  ;
  input \idma_DTMP_L_reg[7]/P0001  ;
  input \idma_IADi_reg[0]/P0001  ;
  input \idma_IADi_reg[10]/P0001  ;
  input \idma_IADi_reg[11]/P0001  ;
  input \idma_IADi_reg[12]/P0001  ;
  input \idma_IADi_reg[13]/P0001  ;
  input \idma_IADi_reg[14]/P0001  ;
  input \idma_IADi_reg[15]/P0001  ;
  input \idma_IADi_reg[1]/P0001  ;
  input \idma_IADi_reg[2]/P0001  ;
  input \idma_IADi_reg[3]/P0001  ;
  input \idma_IADi_reg[4]/P0001  ;
  input \idma_IADi_reg[5]/P0001  ;
  input \idma_IADi_reg[6]/P0001  ;
  input \idma_IADi_reg[7]/P0001  ;
  input \idma_IADi_reg[8]/P0001  ;
  input \idma_IADi_reg[9]/P0001  ;
  input \idma_IAL_reg/P0001  ;
  input \idma_IDMA_boot_reg/NET0131_reg_syn_10  ;
  input \idma_IDMA_boot_reg/NET0131_reg_syn_2  ;
  input \idma_IDMA_boot_reg/NET0131_reg_syn_8  ;
  input \idma_IRDn_reg/P0001  ;
  input \idma_ISn_reg/P0001  ;
  input \idma_IWRn_reg/P0001  ;
  input \idma_PCrd_1st_reg/NET0131  ;
  input \idma_PM_1st_reg/NET0131  ;
  input \idma_RDCMD_d1_reg/P0001  ;
  input \idma_RDCMD_reg/P0001  ;
  input \idma_RDcnt_reg[0]/NET0131  ;
  input \idma_RDcnt_reg[1]/NET0131  ;
  input \idma_RDcnt_reg[2]/NET0131  ;
  input \idma_RDcyc_reg/NET0131  ;
  input \idma_WRCMD_d1_reg/P0001  ;
  input \idma_WRCMD_reg/P0001  ;
  input \idma_WRcnt_reg[0]/NET0131  ;
  input \idma_WRcnt_reg[1]/NET0131  ;
  input \idma_WRcnt_reg[2]/NET0131  ;
  input \idma_WRcyc_reg/NET0131  ;
  input \idma_WRtrue_reg/NET0131  ;
  input \memc_DM_oe_reg/P0001  ;
  input \memc_DMo_oe0_reg/P0001  ;
  input \memc_DMo_oe1_reg/P0001  ;
  input \memc_DMo_oe2_reg/P0001  ;
  input \memc_DMo_oe3_reg/P0001  ;
  input \memc_DMo_oe4_reg/P0001  ;
  input \memc_DMo_oe5_reg/P0001  ;
  input \memc_DMo_oe6_reg/P0001  ;
  input \memc_DMo_oe7_reg/P0001  ;
  input \memc_Dread_E_reg/NET0131  ;
  input \memc_Dwrite_C_reg/NET0131  ;
  input \memc_Dwrite_E_reg/NET0131  ;
  input \memc_EXTC_E_reg/NET0131  ;
  input \memc_EXTC_Eg_reg/NET0131_reg_syn_10  ;
  input \memc_EXTC_Eg_reg/NET0131_reg_syn_2  ;
  input \memc_EXTC_Eg_reg/NET0131_reg_syn_8  ;
  input \memc_IOcmd_E_reg/NET0131  ;
  input \memc_LDaST_Eg_reg/NET0131  ;
  input \memc_MMR_web_reg/NET0131  ;
  input \memc_PMo_oe0_reg/P0001  ;
  input \memc_PMo_oe1_reg/P0001  ;
  input \memc_PMo_oe2_reg/P0001  ;
  input \memc_PMo_oe3_reg/P0001  ;
  input \memc_PMo_oe4_reg/P0001  ;
  input \memc_PMo_oe5_reg/P0001  ;
  input \memc_PMo_oe6_reg/P0001  ;
  input \memc_PMo_oe7_reg/P0001  ;
  input \memc_Pread_E_reg/NET0131  ;
  input \memc_Pwrite_C_reg/NET0131  ;
  input \memc_Pwrite_E_reg/NET0131  ;
  input \memc_STI_Cg_reg/NET0131  ;
  input \memc_accDM_E_reg/NET0131  ;
  input \memc_accPM_E_reg/NET0131  ;
  input \memc_ldSREG_E_reg/NET0131  ;
  input \memc_selMIO_E_reg/P0001  ;
  input \memc_usysr_DO_reg[0]/NET0131  ;
  input \memc_usysr_DO_reg[10]/NET0131  ;
  input \memc_usysr_DO_reg[11]/NET0131  ;
  input \memc_usysr_DO_reg[12]/NET0131  ;
  input \memc_usysr_DO_reg[13]/NET0131  ;
  input \memc_usysr_DO_reg[14]/NET0131  ;
  input \memc_usysr_DO_reg[15]/NET0131  ;
  input \memc_usysr_DO_reg[1]/NET0131  ;
  input \memc_usysr_DO_reg[2]/NET0131  ;
  input \memc_usysr_DO_reg[3]/NET0131  ;
  input \memc_usysr_DO_reg[4]/NET0131  ;
  input \memc_usysr_DO_reg[5]/NET0131  ;
  input \memc_usysr_DO_reg[6]/NET0131  ;
  input \memc_usysr_DO_reg[7]/NET0131  ;
  input \memc_usysr_DO_reg[8]/NET0131  ;
  input \memc_usysr_DO_reg[9]/NET0131  ;
  input \pio_PINT_reg[0]/NET0131  ;
  input \pio_PINT_reg[10]/NET0131  ;
  input \pio_PINT_reg[11]/NET0131  ;
  input \pio_PINT_reg[1]/NET0131  ;
  input \pio_PINT_reg[2]/NET0131  ;
  input \pio_PINT_reg[3]/NET0131  ;
  input \pio_PINT_reg[4]/NET0131  ;
  input \pio_PINT_reg[5]/NET0131  ;
  input \pio_PINT_reg[6]/NET0131  ;
  input \pio_PINT_reg[7]/NET0131  ;
  input \pio_PINT_reg[8]/NET0131  ;
  input \pio_PINT_reg[9]/NET0131  ;
  input \pio_PIO_IN_P_reg[0]/P0001  ;
  input \pio_PIO_IN_P_reg[10]/P0001  ;
  input \pio_PIO_IN_P_reg[11]/P0001  ;
  input \pio_PIO_IN_P_reg[1]/P0001  ;
  input \pio_PIO_IN_P_reg[2]/P0001  ;
  input \pio_PIO_IN_P_reg[3]/P0001  ;
  input \pio_PIO_IN_P_reg[4]/P0001  ;
  input \pio_PIO_IN_P_reg[5]/P0001  ;
  input \pio_PIO_IN_P_reg[6]/P0001  ;
  input \pio_PIO_IN_P_reg[7]/P0001  ;
  input \pio_PIO_IN_P_reg[8]/P0001  ;
  input \pio_PIO_IN_P_reg[9]/P0001  ;
  input \pio_PIO_RES_OUT_reg[0]/P0001  ;
  input \pio_PIO_RES_OUT_reg[10]/P0001  ;
  input \pio_PIO_RES_OUT_reg[11]/P0001  ;
  input \pio_PIO_RES_OUT_reg[1]/P0001  ;
  input \pio_PIO_RES_OUT_reg[2]/P0001  ;
  input \pio_PIO_RES_OUT_reg[3]/P0001  ;
  input \pio_PIO_RES_OUT_reg[4]/P0001  ;
  input \pio_PIO_RES_OUT_reg[5]/P0001  ;
  input \pio_PIO_RES_OUT_reg[6]/P0001  ;
  input \pio_PIO_RES_OUT_reg[7]/P0001  ;
  input \pio_PIO_RES_OUT_reg[8]/P0001  ;
  input \pio_PIO_RES_OUT_reg[9]/P0001  ;
  input \pio_PIO_RES_reg[0]/NET0131  ;
  input \pio_PIO_RES_reg[10]/NET0131  ;
  input \pio_PIO_RES_reg[11]/NET0131  ;
  input \pio_PIO_RES_reg[1]/NET0131  ;
  input \pio_PIO_RES_reg[2]/NET0131  ;
  input \pio_PIO_RES_reg[3]/NET0131  ;
  input \pio_PIO_RES_reg[4]/NET0131  ;
  input \pio_PIO_RES_reg[5]/NET0131  ;
  input \pio_PIO_RES_reg[6]/NET0131  ;
  input \pio_PIO_RES_reg[7]/NET0131  ;
  input \pio_PIO_RES_reg[8]/NET0131  ;
  input \pio_PIO_RES_reg[9]/NET0131  ;
  input \pio_pmask_reg_DO_reg[0]/NET0131  ;
  input \pio_pmask_reg_DO_reg[10]/NET0131  ;
  input \pio_pmask_reg_DO_reg[11]/NET0131  ;
  input \pio_pmask_reg_DO_reg[1]/NET0131  ;
  input \pio_pmask_reg_DO_reg[2]/NET0131  ;
  input \pio_pmask_reg_DO_reg[3]/NET0131  ;
  input \pio_pmask_reg_DO_reg[4]/NET0131  ;
  input \pio_pmask_reg_DO_reg[5]/NET0131  ;
  input \pio_pmask_reg_DO_reg[6]/NET0131  ;
  input \pio_pmask_reg_DO_reg[7]/NET0131  ;
  input \pio_pmask_reg_DO_reg[8]/NET0131  ;
  input \pio_pmask_reg_DO_reg[9]/NET0131  ;
  input \regout_STD_C_reg[0]/P0001  ;
  input \regout_STD_C_reg[10]/P0001  ;
  input \regout_STD_C_reg[11]/P0001  ;
  input \regout_STD_C_reg[12]/P0001  ;
  input \regout_STD_C_reg[13]/P0001  ;
  input \regout_STD_C_reg[14]/P0001  ;
  input \regout_STD_C_reg[15]/P0001  ;
  input \regout_STD_C_reg[1]/P0001  ;
  input \regout_STD_C_reg[2]/P0001  ;
  input \regout_STD_C_reg[3]/P0001  ;
  input \regout_STD_C_reg[4]/P0001  ;
  input \regout_STD_C_reg[5]/P0001  ;
  input \regout_STD_C_reg[6]/P0001  ;
  input \regout_STD_C_reg[7]/P0001  ;
  input \regout_STD_C_reg[8]/P0001  ;
  input \regout_STD_C_reg[9]/P0001  ;
  input \sice_CLR_I_reg/NET0131  ;
  input \sice_CLR_M_reg/NET0131  ;
  input \sice_CMRW_reg/NET0131  ;
  input \sice_DBR1_reg[0]/P0001  ;
  input \sice_DBR1_reg[10]/P0001  ;
  input \sice_DBR1_reg[11]/P0001  ;
  input \sice_DBR1_reg[12]/P0001  ;
  input \sice_DBR1_reg[13]/P0001  ;
  input \sice_DBR1_reg[14]/P0001  ;
  input \sice_DBR1_reg[15]/P0001  ;
  input \sice_DBR1_reg[16]/P0001  ;
  input \sice_DBR1_reg[17]/P0001  ;
  input \sice_DBR1_reg[18]/P0001  ;
  input \sice_DBR1_reg[1]/P0001  ;
  input \sice_DBR1_reg[2]/P0001  ;
  input \sice_DBR1_reg[3]/P0001  ;
  input \sice_DBR1_reg[4]/P0001  ;
  input \sice_DBR1_reg[5]/P0001  ;
  input \sice_DBR1_reg[6]/P0001  ;
  input \sice_DBR1_reg[7]/P0001  ;
  input \sice_DBR1_reg[8]/P0001  ;
  input \sice_DBR1_reg[9]/P0001  ;
  input \sice_DBR2_reg[0]/P0001  ;
  input \sice_DBR2_reg[10]/P0001  ;
  input \sice_DBR2_reg[11]/P0001  ;
  input \sice_DBR2_reg[12]/P0001  ;
  input \sice_DBR2_reg[13]/P0001  ;
  input \sice_DBR2_reg[14]/P0001  ;
  input \sice_DBR2_reg[15]/P0001  ;
  input \sice_DBR2_reg[16]/P0001  ;
  input \sice_DBR2_reg[17]/P0001  ;
  input \sice_DBR2_reg[18]/P0001  ;
  input \sice_DBR2_reg[1]/P0001  ;
  input \sice_DBR2_reg[2]/P0001  ;
  input \sice_DBR2_reg[3]/P0001  ;
  input \sice_DBR2_reg[4]/P0001  ;
  input \sice_DBR2_reg[5]/P0001  ;
  input \sice_DBR2_reg[6]/P0001  ;
  input \sice_DBR2_reg[7]/P0001  ;
  input \sice_DBR2_reg[8]/P0001  ;
  input \sice_DBR2_reg[9]/P0001  ;
  input \sice_DMR1_reg[0]/NET0131  ;
  input \sice_DMR1_reg[10]/NET0131  ;
  input \sice_DMR1_reg[11]/NET0131  ;
  input \sice_DMR1_reg[12]/NET0131  ;
  input \sice_DMR1_reg[13]/NET0131  ;
  input \sice_DMR1_reg[14]/NET0131  ;
  input \sice_DMR1_reg[15]/NET0131  ;
  input \sice_DMR1_reg[16]/NET0131  ;
  input \sice_DMR1_reg[17]/NET0131  ;
  input \sice_DMR1_reg[1]/NET0131  ;
  input \sice_DMR1_reg[2]/NET0131  ;
  input \sice_DMR1_reg[3]/NET0131  ;
  input \sice_DMR1_reg[4]/NET0131  ;
  input \sice_DMR1_reg[5]/NET0131  ;
  input \sice_DMR1_reg[6]/NET0131  ;
  input \sice_DMR1_reg[7]/NET0131  ;
  input \sice_DMR1_reg[8]/NET0131  ;
  input \sice_DMR1_reg[9]/NET0131  ;
  input \sice_DMR2_reg[0]/NET0131  ;
  input \sice_DMR2_reg[10]/NET0131  ;
  input \sice_DMR2_reg[11]/NET0131  ;
  input \sice_DMR2_reg[12]/NET0131  ;
  input \sice_DMR2_reg[13]/NET0131  ;
  input \sice_DMR2_reg[14]/NET0131  ;
  input \sice_DMR2_reg[15]/NET0131  ;
  input \sice_DMR2_reg[16]/NET0131  ;
  input \sice_DMR2_reg[17]/NET0131  ;
  input \sice_DMR2_reg[1]/NET0131  ;
  input \sice_DMR2_reg[2]/NET0131  ;
  input \sice_DMR2_reg[3]/NET0131  ;
  input \sice_DMR2_reg[4]/NET0131  ;
  input \sice_DMR2_reg[5]/NET0131  ;
  input \sice_DMR2_reg[6]/NET0131  ;
  input \sice_DMR2_reg[7]/NET0131  ;
  input \sice_DMR2_reg[8]/NET0131  ;
  input \sice_DMR2_reg[9]/NET0131  ;
  input \sice_GOICE_1_reg/NET0131  ;
  input \sice_GOICE_2_reg/NET0131  ;
  input \sice_GOICE_s1_reg/NET0131  ;
  input \sice_GOICE_syn_reg/P0001  ;
  input \sice_GO_NX_reg/NET0131  ;
  input \sice_GO_NXi_reg/NET0131  ;
  input \sice_HALT_E_reg/P0001  ;
  input \sice_IAR_reg[0]/NET0131  ;
  input \sice_IAR_reg[1]/NET0131  ;
  input \sice_IAR_reg[2]/NET0131  ;
  input \sice_IAR_reg[3]/NET0131  ;
  input \sice_IBR1_reg[0]/P0001  ;
  input \sice_IBR1_reg[10]/P0001  ;
  input \sice_IBR1_reg[11]/P0001  ;
  input \sice_IBR1_reg[12]/P0001  ;
  input \sice_IBR1_reg[13]/P0001  ;
  input \sice_IBR1_reg[14]/P0001  ;
  input \sice_IBR1_reg[15]/P0001  ;
  input \sice_IBR1_reg[16]/P0001  ;
  input \sice_IBR1_reg[17]/P0001  ;
  input \sice_IBR1_reg[1]/P0001  ;
  input \sice_IBR1_reg[2]/P0001  ;
  input \sice_IBR1_reg[3]/P0001  ;
  input \sice_IBR1_reg[4]/P0001  ;
  input \sice_IBR1_reg[5]/P0001  ;
  input \sice_IBR1_reg[6]/P0001  ;
  input \sice_IBR1_reg[7]/P0001  ;
  input \sice_IBR1_reg[8]/P0001  ;
  input \sice_IBR1_reg[9]/P0001  ;
  input \sice_IBR2_reg[0]/P0001  ;
  input \sice_IBR2_reg[10]/P0001  ;
  input \sice_IBR2_reg[11]/P0001  ;
  input \sice_IBR2_reg[12]/P0001  ;
  input \sice_IBR2_reg[13]/P0001  ;
  input \sice_IBR2_reg[14]/P0001  ;
  input \sice_IBR2_reg[15]/P0001  ;
  input \sice_IBR2_reg[16]/P0001  ;
  input \sice_IBR2_reg[17]/P0001  ;
  input \sice_IBR2_reg[1]/P0001  ;
  input \sice_IBR2_reg[2]/P0001  ;
  input \sice_IBR2_reg[3]/P0001  ;
  input \sice_IBR2_reg[4]/P0001  ;
  input \sice_IBR2_reg[5]/P0001  ;
  input \sice_IBR2_reg[6]/P0001  ;
  input \sice_IBR2_reg[7]/P0001  ;
  input \sice_IBR2_reg[8]/P0001  ;
  input \sice_IBR2_reg[9]/P0001  ;
  input \sice_ICS_reg[0]/NET0131  ;
  input \sice_ICS_reg[1]/NET0131  ;
  input \sice_ICS_reg[2]/NET0131  ;
  input \sice_ICYC_clr_reg/NET0131  ;
  input \sice_ICYC_en_reg/NET0131  ;
  input \sice_ICYC_en_syn_reg/P0001  ;
  input \sice_ICYC_reg[0]/NET0131  ;
  input \sice_ICYC_reg[10]/NET0131  ;
  input \sice_ICYC_reg[11]/NET0131  ;
  input \sice_ICYC_reg[12]/NET0131  ;
  input \sice_ICYC_reg[13]/NET0131  ;
  input \sice_ICYC_reg[14]/NET0131  ;
  input \sice_ICYC_reg[15]/NET0131  ;
  input \sice_ICYC_reg[16]/NET0131  ;
  input \sice_ICYC_reg[17]/NET0131  ;
  input \sice_ICYC_reg[18]/NET0131  ;
  input \sice_ICYC_reg[19]/NET0131  ;
  input \sice_ICYC_reg[1]/NET0131  ;
  input \sice_ICYC_reg[20]/NET0131  ;
  input \sice_ICYC_reg[21]/NET0131  ;
  input \sice_ICYC_reg[22]/NET0131  ;
  input \sice_ICYC_reg[23]/NET0131  ;
  input \sice_ICYC_reg[2]/NET0131  ;
  input \sice_ICYC_reg[3]/NET0131  ;
  input \sice_ICYC_reg[4]/NET0131  ;
  input \sice_ICYC_reg[5]/NET0131  ;
  input \sice_ICYC_reg[6]/NET0131  ;
  input \sice_ICYC_reg[7]/NET0131  ;
  input \sice_ICYC_reg[8]/NET0131  ;
  input \sice_ICYC_reg[9]/NET0131  ;
  input \sice_IDONE_reg/NET0131  ;
  input \sice_IIRC_reg[0]/NET0131  ;
  input \sice_IIRC_reg[10]/NET0131  ;
  input \sice_IIRC_reg[11]/NET0131  ;
  input \sice_IIRC_reg[12]/NET0131  ;
  input \sice_IIRC_reg[13]/NET0131  ;
  input \sice_IIRC_reg[14]/NET0131  ;
  input \sice_IIRC_reg[15]/NET0131  ;
  input \sice_IIRC_reg[16]/NET0131  ;
  input \sice_IIRC_reg[17]/NET0131  ;
  input \sice_IIRC_reg[18]/NET0131  ;
  input \sice_IIRC_reg[19]/NET0131  ;
  input \sice_IIRC_reg[1]/NET0131  ;
  input \sice_IIRC_reg[20]/NET0131  ;
  input \sice_IIRC_reg[21]/NET0131  ;
  input \sice_IIRC_reg[22]/NET0131  ;
  input \sice_IIRC_reg[23]/NET0131  ;
  input \sice_IIRC_reg[2]/NET0131  ;
  input \sice_IIRC_reg[3]/NET0131  ;
  input \sice_IIRC_reg[4]/NET0131  ;
  input \sice_IIRC_reg[5]/NET0131  ;
  input \sice_IIRC_reg[6]/NET0131  ;
  input \sice_IIRC_reg[7]/NET0131  ;
  input \sice_IIRC_reg[8]/NET0131  ;
  input \sice_IIRC_reg[9]/NET0131  ;
  input \sice_IMR1_reg[0]/NET0131  ;
  input \sice_IMR1_reg[10]/NET0131  ;
  input \sice_IMR1_reg[11]/NET0131  ;
  input \sice_IMR1_reg[12]/NET0131  ;
  input \sice_IMR1_reg[13]/NET0131  ;
  input \sice_IMR1_reg[14]/NET0131  ;
  input \sice_IMR1_reg[15]/NET0131  ;
  input \sice_IMR1_reg[16]/NET0131  ;
  input \sice_IMR1_reg[17]/NET0131  ;
  input \sice_IMR1_reg[1]/NET0131  ;
  input \sice_IMR1_reg[2]/NET0131  ;
  input \sice_IMR1_reg[3]/NET0131  ;
  input \sice_IMR1_reg[4]/NET0131  ;
  input \sice_IMR1_reg[5]/NET0131  ;
  input \sice_IMR1_reg[6]/NET0131  ;
  input \sice_IMR1_reg[7]/NET0131  ;
  input \sice_IMR1_reg[8]/NET0131  ;
  input \sice_IMR1_reg[9]/NET0131  ;
  input \sice_IMR2_reg[0]/NET0131  ;
  input \sice_IMR2_reg[10]/NET0131  ;
  input \sice_IMR2_reg[11]/NET0131  ;
  input \sice_IMR2_reg[12]/NET0131  ;
  input \sice_IMR2_reg[13]/NET0131  ;
  input \sice_IMR2_reg[14]/NET0131  ;
  input \sice_IMR2_reg[15]/NET0131  ;
  input \sice_IMR2_reg[16]/NET0131  ;
  input \sice_IMR2_reg[17]/NET0131  ;
  input \sice_IMR2_reg[1]/NET0131  ;
  input \sice_IMR2_reg[2]/NET0131  ;
  input \sice_IMR2_reg[3]/NET0131  ;
  input \sice_IMR2_reg[4]/NET0131  ;
  input \sice_IMR2_reg[5]/NET0131  ;
  input \sice_IMR2_reg[6]/NET0131  ;
  input \sice_IMR2_reg[7]/NET0131  ;
  input \sice_IMR2_reg[8]/NET0131  ;
  input \sice_IMR2_reg[9]/NET0131  ;
  input \sice_IRR_reg[0]/P0001  ;
  input \sice_IRR_reg[10]/P0001  ;
  input \sice_IRR_reg[11]/P0001  ;
  input \sice_IRR_reg[12]/P0001  ;
  input \sice_IRR_reg[13]/P0001  ;
  input \sice_IRR_reg[1]/P0001  ;
  input \sice_IRR_reg[2]/P0001  ;
  input \sice_IRR_reg[3]/P0001  ;
  input \sice_IRR_reg[4]/P0001  ;
  input \sice_IRR_reg[5]/P0001  ;
  input \sice_IRR_reg[6]/P0001  ;
  input \sice_IRR_reg[7]/P0001  ;
  input \sice_IRR_reg[8]/P0001  ;
  input \sice_IRR_reg[9]/P0001  ;
  input \sice_IRST_reg/NET0131  ;
  input \sice_IRST_syn_reg/P0001  ;
  input \sice_ITR_reg[0]/NET0131  ;
  input \sice_ITR_reg[1]/NET0131  ;
  input \sice_ITR_reg[2]/NET0131  ;
  input \sice_OE_reg/P0001  ;
  input \sice_RCS_reg[0]/NET0131  ;
  input \sice_RCS_reg[1]/NET0131  ;
  input \sice_RST_req_reg/NET0131  ;
  input \sice_SPC_reg[0]/P0001  ;
  input \sice_SPC_reg[10]/P0001  ;
  input \sice_SPC_reg[11]/P0001  ;
  input \sice_SPC_reg[12]/P0001  ;
  input \sice_SPC_reg[13]/P0001  ;
  input \sice_SPC_reg[14]/P0001  ;
  input \sice_SPC_reg[15]/P0001  ;
  input \sice_SPC_reg[16]/P0001  ;
  input \sice_SPC_reg[17]/P0001  ;
  input \sice_SPC_reg[18]/P0001  ;
  input \sice_SPC_reg[19]/P0001  ;
  input \sice_SPC_reg[1]/P0001  ;
  input \sice_SPC_reg[20]/P0001  ;
  input \sice_SPC_reg[21]/P0001  ;
  input \sice_SPC_reg[22]/P0001  ;
  input \sice_SPC_reg[23]/P0001  ;
  input \sice_SPC_reg[2]/P0001  ;
  input \sice_SPC_reg[3]/P0001  ;
  input \sice_SPC_reg[4]/P0001  ;
  input \sice_SPC_reg[5]/P0001  ;
  input \sice_SPC_reg[6]/P0001  ;
  input \sice_SPC_reg[7]/P0001  ;
  input \sice_SPC_reg[8]/P0001  ;
  input \sice_SPC_reg[9]/P0001  ;
  input \sice_UpdDR_sd1_reg/P0001  ;
  input \sice_UpdDR_sd2_reg/P0001  ;
  input \sice_idr0_reg_DO_reg[0]/P0001  ;
  input \sice_idr0_reg_DO_reg[10]/P0001  ;
  input \sice_idr0_reg_DO_reg[11]/P0001  ;
  input \sice_idr0_reg_DO_reg[1]/P0001  ;
  input \sice_idr0_reg_DO_reg[2]/P0001  ;
  input \sice_idr0_reg_DO_reg[3]/P0001  ;
  input \sice_idr0_reg_DO_reg[4]/P0001  ;
  input \sice_idr0_reg_DO_reg[5]/P0001  ;
  input \sice_idr0_reg_DO_reg[6]/P0001  ;
  input \sice_idr0_reg_DO_reg[7]/P0001  ;
  input \sice_idr0_reg_DO_reg[8]/P0001  ;
  input \sice_idr0_reg_DO_reg[9]/P0001  ;
  input \sice_idr1_reg_DO_reg[0]/P0001  ;
  input \sice_idr1_reg_DO_reg[10]/P0001  ;
  input \sice_idr1_reg_DO_reg[11]/P0001  ;
  input \sice_idr1_reg_DO_reg[1]/P0001  ;
  input \sice_idr1_reg_DO_reg[2]/P0001  ;
  input \sice_idr1_reg_DO_reg[3]/P0001  ;
  input \sice_idr1_reg_DO_reg[4]/P0001  ;
  input \sice_idr1_reg_DO_reg[5]/P0001  ;
  input \sice_idr1_reg_DO_reg[6]/P0001  ;
  input \sice_idr1_reg_DO_reg[7]/P0001  ;
  input \sice_idr1_reg_DO_reg[8]/P0001  ;
  input \sice_idr1_reg_DO_reg[9]/P0001  ;
  input \sport0_cfg_FSi_cnt_reg[0]/NET0131  ;
  input \sport0_cfg_FSi_cnt_reg[10]/NET0131  ;
  input \sport0_cfg_FSi_cnt_reg[11]/NET0131  ;
  input \sport0_cfg_FSi_cnt_reg[12]/NET0131  ;
  input \sport0_cfg_FSi_cnt_reg[13]/NET0131  ;
  input \sport0_cfg_FSi_cnt_reg[14]/NET0131  ;
  input \sport0_cfg_FSi_cnt_reg[15]/NET0131  ;
  input \sport0_cfg_FSi_cnt_reg[1]/NET0131  ;
  input \sport0_cfg_FSi_cnt_reg[2]/NET0131  ;
  input \sport0_cfg_FSi_cnt_reg[3]/NET0131  ;
  input \sport0_cfg_FSi_cnt_reg[4]/NET0131  ;
  input \sport0_cfg_FSi_cnt_reg[5]/NET0131  ;
  input \sport0_cfg_FSi_cnt_reg[6]/NET0131  ;
  input \sport0_cfg_FSi_cnt_reg[7]/NET0131  ;
  input \sport0_cfg_FSi_cnt_reg[8]/NET0131  ;
  input \sport0_cfg_FSi_cnt_reg[9]/NET0131  ;
  input \sport0_cfg_FSi_reg/NET0131  ;
  input \sport0_cfg_RFSg_d1_reg/NET0131  ;
  input \sport0_cfg_RFSg_d2_reg/NET0131  ;
  input \sport0_cfg_RFSg_d3_reg/NET0131  ;
  input \sport0_cfg_RFSgi_d_reg/NET0131  ;
  input \sport0_cfg_SCLKi_cnt_reg[0]/NET0131  ;
  input \sport0_cfg_SCLKi_cnt_reg[10]/NET0131  ;
  input \sport0_cfg_SCLKi_cnt_reg[11]/NET0131  ;
  input \sport0_cfg_SCLKi_cnt_reg[12]/NET0131  ;
  input \sport0_cfg_SCLKi_cnt_reg[13]/NET0131  ;
  input \sport0_cfg_SCLKi_cnt_reg[14]/NET0131  ;
  input \sport0_cfg_SCLKi_cnt_reg[15]/NET0131  ;
  input \sport0_cfg_SCLKi_cnt_reg[1]/NET0131  ;
  input \sport0_cfg_SCLKi_cnt_reg[2]/NET0131  ;
  input \sport0_cfg_SCLKi_cnt_reg[3]/NET0131  ;
  input \sport0_cfg_SCLKi_cnt_reg[4]/NET0131  ;
  input \sport0_cfg_SCLKi_cnt_reg[5]/NET0131  ;
  input \sport0_cfg_SCLKi_cnt_reg[6]/NET0131  ;
  input \sport0_cfg_SCLKi_cnt_reg[7]/NET0131  ;
  input \sport0_cfg_SCLKi_cnt_reg[8]/NET0131  ;
  input \sport0_cfg_SCLKi_cnt_reg[9]/NET0131  ;
  input \sport0_cfg_SCLKi_h_reg/NET0131  ;
  input \sport0_cfg_SP_ENg_D1_reg/P0001  ;
  input \sport0_cfg_SP_ENg_reg/NET0131  ;
  input \sport0_cfg_TFSg_d1_reg/NET0131  ;
  input \sport0_cfg_TFSg_d2_reg/NET0131  ;
  input \sport0_cfg_TFSg_d3_reg/NET0131  ;
  input \sport0_cfg_TFSgi_d_reg/NET0131  ;
  input \sport0_regs_AUTO_a_reg[12]/NET0131  ;
  input \sport0_regs_AUTO_a_reg[13]/NET0131  ;
  input \sport0_regs_AUTO_a_reg[14]/NET0131  ;
  input \sport0_regs_AUTO_a_reg[15]/NET0131  ;
  input \sport0_regs_AUTOreg_DO_reg[0]/NET0131  ;
  input \sport0_regs_AUTOreg_DO_reg[10]/NET0131  ;
  input \sport0_regs_AUTOreg_DO_reg[11]/NET0131  ;
  input \sport0_regs_AUTOreg_DO_reg[1]/NET0131  ;
  input \sport0_regs_AUTOreg_DO_reg[2]/NET0131  ;
  input \sport0_regs_AUTOreg_DO_reg[3]/NET0131  ;
  input \sport0_regs_AUTOreg_DO_reg[4]/NET0131  ;
  input \sport0_regs_AUTOreg_DO_reg[5]/NET0131  ;
  input \sport0_regs_AUTOreg_DO_reg[6]/NET0131  ;
  input \sport0_regs_AUTOreg_DO_reg[7]/NET0131  ;
  input \sport0_regs_AUTOreg_DO_reg[8]/NET0131  ;
  input \sport0_regs_AUTOreg_DO_reg[9]/NET0131  ;
  input \sport0_regs_FSDIVreg_DO_reg[0]/NET0131  ;
  input \sport0_regs_FSDIVreg_DO_reg[10]/NET0131  ;
  input \sport0_regs_FSDIVreg_DO_reg[11]/NET0131  ;
  input \sport0_regs_FSDIVreg_DO_reg[12]/NET0131  ;
  input \sport0_regs_FSDIVreg_DO_reg[13]/NET0131  ;
  input \sport0_regs_FSDIVreg_DO_reg[14]/NET0131  ;
  input \sport0_regs_FSDIVreg_DO_reg[15]/NET0131  ;
  input \sport0_regs_FSDIVreg_DO_reg[1]/NET0131  ;
  input \sport0_regs_FSDIVreg_DO_reg[2]/NET0131  ;
  input \sport0_regs_FSDIVreg_DO_reg[3]/NET0131  ;
  input \sport0_regs_FSDIVreg_DO_reg[4]/NET0131  ;
  input \sport0_regs_FSDIVreg_DO_reg[5]/NET0131  ;
  input \sport0_regs_FSDIVreg_DO_reg[6]/NET0131  ;
  input \sport0_regs_FSDIVreg_DO_reg[7]/NET0131  ;
  input \sport0_regs_FSDIVreg_DO_reg[8]/NET0131  ;
  input \sport0_regs_FSDIVreg_DO_reg[9]/NET0131  ;
  input \sport0_regs_MWORDreg_DO_reg[0]/NET0131  ;
  input \sport0_regs_MWORDreg_DO_reg[10]/NET0131  ;
  input \sport0_regs_MWORDreg_DO_reg[1]/NET0131  ;
  input \sport0_regs_MWORDreg_DO_reg[2]/NET0131  ;
  input \sport0_regs_MWORDreg_DO_reg[3]/NET0131  ;
  input \sport0_regs_MWORDreg_DO_reg[4]/NET0131  ;
  input \sport0_regs_MWORDreg_DO_reg[5]/NET0131  ;
  input \sport0_regs_MWORDreg_DO_reg[6]/NET0131  ;
  input \sport0_regs_MWORDreg_DO_reg[7]/NET0131  ;
  input \sport0_regs_MWORDreg_DO_reg[8]/NET0131  ;
  input \sport0_regs_MWORDreg_DO_reg[9]/NET0131  ;
  input \sport0_regs_SCLKDIVreg_DO_reg[0]/NET0131  ;
  input \sport0_regs_SCLKDIVreg_DO_reg[10]/NET0131  ;
  input \sport0_regs_SCLKDIVreg_DO_reg[11]/NET0131  ;
  input \sport0_regs_SCLKDIVreg_DO_reg[12]/NET0131  ;
  input \sport0_regs_SCLKDIVreg_DO_reg[13]/NET0131  ;
  input \sport0_regs_SCLKDIVreg_DO_reg[14]/NET0131  ;
  input \sport0_regs_SCLKDIVreg_DO_reg[15]/NET0131  ;
  input \sport0_regs_SCLKDIVreg_DO_reg[1]/NET0131  ;
  input \sport0_regs_SCLKDIVreg_DO_reg[2]/NET0131  ;
  input \sport0_regs_SCLKDIVreg_DO_reg[3]/NET0131  ;
  input \sport0_regs_SCLKDIVreg_DO_reg[4]/NET0131  ;
  input \sport0_regs_SCLKDIVreg_DO_reg[5]/NET0131  ;
  input \sport0_regs_SCLKDIVreg_DO_reg[6]/NET0131  ;
  input \sport0_regs_SCLKDIVreg_DO_reg[7]/NET0131  ;
  input \sport0_regs_SCLKDIVreg_DO_reg[8]/NET0131  ;
  input \sport0_regs_SCLKDIVreg_DO_reg[9]/NET0131  ;
  input \sport0_regs_SCTLreg_DO_reg[0]/NET0131  ;
  input \sport0_regs_SCTLreg_DO_reg[10]/NET0131  ;
  input \sport0_regs_SCTLreg_DO_reg[11]/NET0131  ;
  input \sport0_regs_SCTLreg_DO_reg[12]/NET0131  ;
  input \sport0_regs_SCTLreg_DO_reg[13]/NET0131  ;
  input \sport0_regs_SCTLreg_DO_reg[15]/NET0131  ;
  input \sport0_regs_SCTLreg_DO_reg[1]/NET0131  ;
  input \sport0_regs_SCTLreg_DO_reg[2]/NET0131  ;
  input \sport0_regs_SCTLreg_DO_reg[3]/NET0131  ;
  input \sport0_regs_SCTLreg_DO_reg[4]/NET0131  ;
  input \sport0_regs_SCTLreg_DO_reg[5]/NET0131  ;
  input \sport0_regs_SCTLreg_DO_reg[6]/NET0131  ;
  input \sport0_regs_SCTLreg_DO_reg[7]/NET0131  ;
  input \sport0_rxctl_Bcnt_reg[0]/NET0131  ;
  input \sport0_rxctl_Bcnt_reg[1]/NET0131  ;
  input \sport0_rxctl_Bcnt_reg[2]/NET0131  ;
  input \sport0_rxctl_Bcnt_reg[3]/NET0131  ;
  input \sport0_rxctl_Bcnt_reg[4]/NET0131  ;
  input \sport0_rxctl_ISRa_reg/P0001  ;
  input \sport0_rxctl_LMcnt_reg[0]/NET0131  ;
  input \sport0_rxctl_LMcnt_reg[1]/NET0131  ;
  input \sport0_rxctl_LMcnt_reg[2]/NET0131  ;
  input \sport0_rxctl_LMcnt_reg[3]/NET0131  ;
  input \sport0_rxctl_LMcnt_reg[4]/NET0131  ;
  input \sport0_rxctl_RCS_reg[0]/NET0131  ;
  input \sport0_rxctl_RCS_reg[1]/NET0131  ;
  input \sport0_rxctl_RCS_reg[2]/NET0131  ;
  input \sport0_rxctl_RSreq_reg/NET0131  ;
  input \sport0_rxctl_RXSHT_reg[0]/P0001  ;
  input \sport0_rxctl_RXSHT_reg[10]/P0001  ;
  input \sport0_rxctl_RXSHT_reg[11]/P0001  ;
  input \sport0_rxctl_RXSHT_reg[12]/P0001  ;
  input \sport0_rxctl_RXSHT_reg[13]/P0001  ;
  input \sport0_rxctl_RXSHT_reg[14]/P0001  ;
  input \sport0_rxctl_RXSHT_reg[15]/P0001  ;
  input \sport0_rxctl_RXSHT_reg[1]/P0001  ;
  input \sport0_rxctl_RXSHT_reg[2]/P0001  ;
  input \sport0_rxctl_RXSHT_reg[3]/P0001  ;
  input \sport0_rxctl_RXSHT_reg[4]/P0001  ;
  input \sport0_rxctl_RXSHT_reg[5]/P0001  ;
  input \sport0_rxctl_RXSHT_reg[6]/P0001  ;
  input \sport0_rxctl_RXSHT_reg[7]/P0001  ;
  input \sport0_rxctl_RXSHT_reg[8]/P0001  ;
  input \sport0_rxctl_RXSHT_reg[9]/P0001  ;
  input \sport0_rxctl_RX_reg[0]/P0001  ;
  input \sport0_rxctl_RX_reg[10]/P0001  ;
  input \sport0_rxctl_RX_reg[11]/P0001  ;
  input \sport0_rxctl_RX_reg[12]/P0001  ;
  input \sport0_rxctl_RX_reg[13]/P0001  ;
  input \sport0_rxctl_RX_reg[14]/P0001  ;
  input \sport0_rxctl_RX_reg[15]/P0001  ;
  input \sport0_rxctl_RX_reg[1]/P0001  ;
  input \sport0_rxctl_RX_reg[2]/P0001  ;
  input \sport0_rxctl_RX_reg[3]/P0001  ;
  input \sport0_rxctl_RX_reg[4]/P0001  ;
  input \sport0_rxctl_RX_reg[5]/P0001  ;
  input \sport0_rxctl_RX_reg[6]/P0001  ;
  input \sport0_rxctl_RX_reg[7]/P0001  ;
  input \sport0_rxctl_RX_reg[8]/P0001  ;
  input \sport0_rxctl_RX_reg[9]/P0001  ;
  input \sport0_rxctl_SLOT1_EXT_reg[2]/NET0131  ;
  input \sport0_rxctl_SLOT1_EXT_reg[3]/NET0131  ;
  input \sport0_rxctl_TAG_SLOT_reg/P0001  ;
  input \sport0_rxctl_Wcnt_reg[0]/NET0131  ;
  input \sport0_rxctl_Wcnt_reg[1]/NET0131  ;
  input \sport0_rxctl_Wcnt_reg[2]/NET0131  ;
  input \sport0_rxctl_Wcnt_reg[3]/NET0131  ;
  input \sport0_rxctl_Wcnt_reg[4]/NET0131  ;
  input \sport0_rxctl_Wcnt_reg[5]/NET0131  ;
  input \sport0_rxctl_Wcnt_reg[6]/NET0131  ;
  input \sport0_rxctl_Wcnt_reg[7]/NET0131  ;
  input \sport0_rxctl_a_sync1_reg/P0001  ;
  input \sport0_rxctl_a_sync2_reg/P0001  ;
  input \sport0_rxctl_ldRX_cmp_reg/P0001  ;
  input \sport0_rxctl_sht2nd_reg/P0001  ;
  input \sport0_txctl_Bcnt_reg[0]/NET0131  ;
  input \sport0_txctl_Bcnt_reg[1]/NET0131  ;
  input \sport0_txctl_Bcnt_reg[2]/NET0131  ;
  input \sport0_txctl_Bcnt_reg[3]/NET0131  ;
  input \sport0_txctl_Bcnt_reg[4]/NET0131  ;
  input \sport0_txctl_SP_EN_D1_reg/P0001  ;
  input \sport0_txctl_TCS_reg[0]/NET0131  ;
  input \sport0_txctl_TCS_reg[1]/NET0131  ;
  input \sport0_txctl_TCS_reg[2]/NET0131  ;
  input \sport0_txctl_TSreq_reg/NET0131  ;
  input \sport0_txctl_TSreqi_reg/NET0131  ;
  input \sport0_txctl_TXSHT_reg[0]/P0001  ;
  input \sport0_txctl_TXSHT_reg[10]/P0001  ;
  input \sport0_txctl_TXSHT_reg[11]/P0001  ;
  input \sport0_txctl_TXSHT_reg[12]/P0001  ;
  input \sport0_txctl_TXSHT_reg[13]/P0001  ;
  input \sport0_txctl_TXSHT_reg[14]/P0001  ;
  input \sport0_txctl_TXSHT_reg[15]/P0001  ;
  input \sport0_txctl_TXSHT_reg[1]/P0001  ;
  input \sport0_txctl_TXSHT_reg[2]/P0001  ;
  input \sport0_txctl_TXSHT_reg[3]/P0001  ;
  input \sport0_txctl_TXSHT_reg[4]/P0001  ;
  input \sport0_txctl_TXSHT_reg[5]/P0001  ;
  input \sport0_txctl_TXSHT_reg[6]/P0001  ;
  input \sport0_txctl_TXSHT_reg[7]/P0001  ;
  input \sport0_txctl_TXSHT_reg[8]/P0001  ;
  input \sport0_txctl_TXSHT_reg[9]/P0001  ;
  input \sport0_txctl_TX_reg[0]/P0001  ;
  input \sport0_txctl_TX_reg[10]/P0001  ;
  input \sport0_txctl_TX_reg[11]/P0001  ;
  input \sport0_txctl_TX_reg[12]/P0001  ;
  input \sport0_txctl_TX_reg[13]/P0001  ;
  input \sport0_txctl_TX_reg[14]/P0001  ;
  input \sport0_txctl_TX_reg[15]/P0001  ;
  input \sport0_txctl_TX_reg[1]/P0001  ;
  input \sport0_txctl_TX_reg[2]/P0001  ;
  input \sport0_txctl_TX_reg[3]/P0001  ;
  input \sport0_txctl_TX_reg[4]/P0001  ;
  input \sport0_txctl_TX_reg[5]/P0001  ;
  input \sport0_txctl_TX_reg[6]/P0001  ;
  input \sport0_txctl_TX_reg[7]/P0001  ;
  input \sport0_txctl_TX_reg[8]/P0001  ;
  input \sport0_txctl_TX_reg[9]/P0001  ;
  input \sport0_txctl_Wcnt_reg[0]/NET0131  ;
  input \sport0_txctl_Wcnt_reg[1]/NET0131  ;
  input \sport0_txctl_Wcnt_reg[2]/NET0131  ;
  input \sport0_txctl_Wcnt_reg[3]/NET0131  ;
  input \sport0_txctl_Wcnt_reg[4]/NET0131  ;
  input \sport0_txctl_Wcnt_reg[5]/NET0131  ;
  input \sport0_txctl_Wcnt_reg[6]/NET0131  ;
  input \sport0_txctl_Wcnt_reg[7]/NET0131  ;
  input \sport0_txctl_b_sync1_reg/P0001  ;
  input \sport0_txctl_c_sync1_reg/P0001  ;
  input \sport0_txctl_c_sync2_reg/P0001  ;
  input \sport0_txctl_ldTX_cmp_reg/P0001  ;
  input \sport1_cfg_FSi_cnt_reg[0]/NET0131  ;
  input \sport1_cfg_FSi_cnt_reg[10]/NET0131  ;
  input \sport1_cfg_FSi_cnt_reg[11]/NET0131  ;
  input \sport1_cfg_FSi_cnt_reg[12]/NET0131  ;
  input \sport1_cfg_FSi_cnt_reg[13]/NET0131  ;
  input \sport1_cfg_FSi_cnt_reg[14]/NET0131  ;
  input \sport1_cfg_FSi_cnt_reg[15]/NET0131  ;
  input \sport1_cfg_FSi_cnt_reg[1]/NET0131  ;
  input \sport1_cfg_FSi_cnt_reg[2]/NET0131  ;
  input \sport1_cfg_FSi_cnt_reg[3]/NET0131  ;
  input \sport1_cfg_FSi_cnt_reg[4]/NET0131  ;
  input \sport1_cfg_FSi_cnt_reg[5]/NET0131  ;
  input \sport1_cfg_FSi_cnt_reg[6]/NET0131  ;
  input \sport1_cfg_FSi_cnt_reg[7]/NET0131  ;
  input \sport1_cfg_FSi_cnt_reg[8]/NET0131  ;
  input \sport1_cfg_FSi_cnt_reg[9]/NET0131  ;
  input \sport1_cfg_FSi_reg/NET0131  ;
  input \sport1_cfg_RFSg_d1_reg/NET0131  ;
  input \sport1_cfg_RFSg_d2_reg/NET0131  ;
  input \sport1_cfg_RFSg_d3_reg/NET0131  ;
  input \sport1_cfg_RFSgi_d_reg/NET0131  ;
  input \sport1_cfg_SCLKi_cnt_reg[0]/NET0131  ;
  input \sport1_cfg_SCLKi_cnt_reg[10]/NET0131  ;
  input \sport1_cfg_SCLKi_cnt_reg[11]/NET0131  ;
  input \sport1_cfg_SCLKi_cnt_reg[12]/NET0131  ;
  input \sport1_cfg_SCLKi_cnt_reg[13]/NET0131  ;
  input \sport1_cfg_SCLKi_cnt_reg[14]/NET0131  ;
  input \sport1_cfg_SCLKi_cnt_reg[15]/NET0131  ;
  input \sport1_cfg_SCLKi_cnt_reg[1]/NET0131  ;
  input \sport1_cfg_SCLKi_cnt_reg[2]/NET0131  ;
  input \sport1_cfg_SCLKi_cnt_reg[3]/NET0131  ;
  input \sport1_cfg_SCLKi_cnt_reg[4]/NET0131  ;
  input \sport1_cfg_SCLKi_cnt_reg[5]/NET0131  ;
  input \sport1_cfg_SCLKi_cnt_reg[6]/NET0131  ;
  input \sport1_cfg_SCLKi_cnt_reg[7]/NET0131  ;
  input \sport1_cfg_SCLKi_cnt_reg[8]/NET0131  ;
  input \sport1_cfg_SCLKi_cnt_reg[9]/NET0131  ;
  input \sport1_cfg_SCLKi_h_reg/NET0131  ;
  input \sport1_cfg_SP_ENg_D1_reg/P0001  ;
  input \sport1_cfg_SP_ENg_reg/NET0131  ;
  input \sport1_cfg_TFSg_d1_reg/NET0131  ;
  input \sport1_cfg_TFSg_d2_reg/NET0131  ;
  input \sport1_cfg_TFSg_d3_reg/NET0131  ;
  input \sport1_cfg_TFSgi_d_reg/NET0131  ;
  input \sport1_regs_AUTOreg_DO_reg[0]/NET0131  ;
  input \sport1_regs_AUTOreg_DO_reg[10]/NET0131  ;
  input \sport1_regs_AUTOreg_DO_reg[11]/NET0131  ;
  input \sport1_regs_AUTOreg_DO_reg[1]/NET0131  ;
  input \sport1_regs_AUTOreg_DO_reg[2]/NET0131  ;
  input \sport1_regs_AUTOreg_DO_reg[3]/NET0131  ;
  input \sport1_regs_AUTOreg_DO_reg[4]/NET0131  ;
  input \sport1_regs_AUTOreg_DO_reg[5]/NET0131  ;
  input \sport1_regs_AUTOreg_DO_reg[6]/NET0131  ;
  input \sport1_regs_AUTOreg_DO_reg[7]/NET0131  ;
  input \sport1_regs_AUTOreg_DO_reg[8]/NET0131  ;
  input \sport1_regs_AUTOreg_DO_reg[9]/NET0131  ;
  input \sport1_regs_FSDIVreg_DO_reg[0]/NET0131  ;
  input \sport1_regs_FSDIVreg_DO_reg[10]/NET0131  ;
  input \sport1_regs_FSDIVreg_DO_reg[11]/NET0131  ;
  input \sport1_regs_FSDIVreg_DO_reg[12]/NET0131  ;
  input \sport1_regs_FSDIVreg_DO_reg[13]/NET0131  ;
  input \sport1_regs_FSDIVreg_DO_reg[14]/NET0131  ;
  input \sport1_regs_FSDIVreg_DO_reg[15]/NET0131  ;
  input \sport1_regs_FSDIVreg_DO_reg[1]/NET0131  ;
  input \sport1_regs_FSDIVreg_DO_reg[2]/NET0131  ;
  input \sport1_regs_FSDIVreg_DO_reg[3]/NET0131  ;
  input \sport1_regs_FSDIVreg_DO_reg[4]/NET0131  ;
  input \sport1_regs_FSDIVreg_DO_reg[5]/NET0131  ;
  input \sport1_regs_FSDIVreg_DO_reg[6]/NET0131  ;
  input \sport1_regs_FSDIVreg_DO_reg[7]/NET0131  ;
  input \sport1_regs_FSDIVreg_DO_reg[8]/NET0131  ;
  input \sport1_regs_FSDIVreg_DO_reg[9]/NET0131  ;
  input \sport1_regs_MWORDreg_DO_reg[0]/NET0131  ;
  input \sport1_regs_MWORDreg_DO_reg[10]/NET0131  ;
  input \sport1_regs_MWORDreg_DO_reg[1]/NET0131  ;
  input \sport1_regs_MWORDreg_DO_reg[2]/NET0131  ;
  input \sport1_regs_MWORDreg_DO_reg[3]/NET0131  ;
  input \sport1_regs_MWORDreg_DO_reg[4]/NET0131  ;
  input \sport1_regs_MWORDreg_DO_reg[5]/NET0131  ;
  input \sport1_regs_MWORDreg_DO_reg[6]/NET0131  ;
  input \sport1_regs_MWORDreg_DO_reg[7]/NET0131  ;
  input \sport1_regs_MWORDreg_DO_reg[8]/NET0131  ;
  input \sport1_regs_MWORDreg_DO_reg[9]/NET0131  ;
  input \sport1_regs_SCLKDIVreg_DO_reg[0]/NET0131  ;
  input \sport1_regs_SCLKDIVreg_DO_reg[10]/NET0131  ;
  input \sport1_regs_SCLKDIVreg_DO_reg[11]/NET0131  ;
  input \sport1_regs_SCLKDIVreg_DO_reg[12]/NET0131  ;
  input \sport1_regs_SCLKDIVreg_DO_reg[13]/NET0131  ;
  input \sport1_regs_SCLKDIVreg_DO_reg[14]/NET0131  ;
  input \sport1_regs_SCLKDIVreg_DO_reg[15]/NET0131  ;
  input \sport1_regs_SCLKDIVreg_DO_reg[1]/NET0131  ;
  input \sport1_regs_SCLKDIVreg_DO_reg[2]/NET0131  ;
  input \sport1_regs_SCLKDIVreg_DO_reg[3]/NET0131  ;
  input \sport1_regs_SCLKDIVreg_DO_reg[4]/NET0131  ;
  input \sport1_regs_SCLKDIVreg_DO_reg[5]/NET0131  ;
  input \sport1_regs_SCLKDIVreg_DO_reg[6]/NET0131  ;
  input \sport1_regs_SCLKDIVreg_DO_reg[7]/NET0131  ;
  input \sport1_regs_SCLKDIVreg_DO_reg[8]/NET0131  ;
  input \sport1_regs_SCLKDIVreg_DO_reg[9]/NET0131  ;
  input \sport1_regs_SCTLreg_DO_reg[0]/NET0131  ;
  input \sport1_regs_SCTLreg_DO_reg[10]/NET0131  ;
  input \sport1_regs_SCTLreg_DO_reg[11]/NET0131  ;
  input \sport1_regs_SCTLreg_DO_reg[12]/NET0131  ;
  input \sport1_regs_SCTLreg_DO_reg[13]/NET0131  ;
  input \sport1_regs_SCTLreg_DO_reg[15]/NET0131  ;
  input \sport1_regs_SCTLreg_DO_reg[1]/NET0131  ;
  input \sport1_regs_SCTLreg_DO_reg[2]/NET0131  ;
  input \sport1_regs_SCTLreg_DO_reg[3]/NET0131  ;
  input \sport1_regs_SCTLreg_DO_reg[4]/NET0131  ;
  input \sport1_regs_SCTLreg_DO_reg[5]/NET0131  ;
  input \sport1_regs_SCTLreg_DO_reg[6]/NET0131  ;
  input \sport1_regs_SCTLreg_DO_reg[7]/NET0131  ;
  input \sport1_rxctl_Bcnt_reg[0]/NET0131  ;
  input \sport1_rxctl_Bcnt_reg[1]/NET0131  ;
  input \sport1_rxctl_Bcnt_reg[2]/NET0131  ;
  input \sport1_rxctl_Bcnt_reg[3]/NET0131  ;
  input \sport1_rxctl_Bcnt_reg[4]/NET0131  ;
  input \sport1_rxctl_ISRa_reg/P0001  ;
  input \sport1_rxctl_LMcnt_reg[0]/NET0131  ;
  input \sport1_rxctl_LMcnt_reg[1]/NET0131  ;
  input \sport1_rxctl_LMcnt_reg[2]/NET0131  ;
  input \sport1_rxctl_LMcnt_reg[3]/NET0131  ;
  input \sport1_rxctl_LMcnt_reg[4]/NET0131  ;
  input \sport1_rxctl_RCS_reg[0]/NET0131  ;
  input \sport1_rxctl_RCS_reg[1]/NET0131  ;
  input \sport1_rxctl_RCS_reg[2]/NET0131  ;
  input \sport1_rxctl_RSreq_reg/NET0131  ;
  input \sport1_rxctl_RXSHT_reg[0]/P0001  ;
  input \sport1_rxctl_RXSHT_reg[10]/P0001  ;
  input \sport1_rxctl_RXSHT_reg[11]/P0001  ;
  input \sport1_rxctl_RXSHT_reg[12]/P0001  ;
  input \sport1_rxctl_RXSHT_reg[13]/P0001  ;
  input \sport1_rxctl_RXSHT_reg[14]/P0001  ;
  input \sport1_rxctl_RXSHT_reg[15]/P0001  ;
  input \sport1_rxctl_RXSHT_reg[1]/P0001  ;
  input \sport1_rxctl_RXSHT_reg[2]/P0001  ;
  input \sport1_rxctl_RXSHT_reg[3]/P0001  ;
  input \sport1_rxctl_RXSHT_reg[4]/P0001  ;
  input \sport1_rxctl_RXSHT_reg[5]/P0001  ;
  input \sport1_rxctl_RXSHT_reg[6]/P0001  ;
  input \sport1_rxctl_RXSHT_reg[7]/P0001  ;
  input \sport1_rxctl_RXSHT_reg[8]/P0001  ;
  input \sport1_rxctl_RXSHT_reg[9]/P0001  ;
  input \sport1_rxctl_RX_reg[0]/P0001  ;
  input \sport1_rxctl_RX_reg[10]/P0001  ;
  input \sport1_rxctl_RX_reg[11]/P0001  ;
  input \sport1_rxctl_RX_reg[12]/P0001  ;
  input \sport1_rxctl_RX_reg[13]/P0001  ;
  input \sport1_rxctl_RX_reg[14]/P0001  ;
  input \sport1_rxctl_RX_reg[15]/P0001  ;
  input \sport1_rxctl_RX_reg[1]/P0001  ;
  input \sport1_rxctl_RX_reg[2]/P0001  ;
  input \sport1_rxctl_RX_reg[3]/P0001  ;
  input \sport1_rxctl_RX_reg[4]/P0001  ;
  input \sport1_rxctl_RX_reg[5]/P0001  ;
  input \sport1_rxctl_RX_reg[6]/P0001  ;
  input \sport1_rxctl_RX_reg[7]/P0001  ;
  input \sport1_rxctl_RX_reg[8]/P0001  ;
  input \sport1_rxctl_RX_reg[9]/P0001  ;
  input \sport1_rxctl_SLOT1_EXT_reg[2]/NET0131  ;
  input \sport1_rxctl_SLOT1_EXT_reg[3]/NET0131  ;
  input \sport1_rxctl_TAG_SLOT_reg/P0001  ;
  input \sport1_rxctl_Wcnt_reg[0]/NET0131  ;
  input \sport1_rxctl_Wcnt_reg[1]/NET0131  ;
  input \sport1_rxctl_Wcnt_reg[2]/NET0131  ;
  input \sport1_rxctl_Wcnt_reg[3]/NET0131  ;
  input \sport1_rxctl_Wcnt_reg[4]/NET0131  ;
  input \sport1_rxctl_Wcnt_reg[5]/NET0131  ;
  input \sport1_rxctl_Wcnt_reg[6]/NET0131  ;
  input \sport1_rxctl_Wcnt_reg[7]/NET0131  ;
  input \sport1_rxctl_a_sync1_reg/P0001  ;
  input \sport1_rxctl_a_sync2_reg/P0001  ;
  input \sport1_rxctl_sht2nd_reg/P0001  ;
  input \sport1_txctl_Bcnt_reg[0]/NET0131  ;
  input \sport1_txctl_Bcnt_reg[1]/NET0131  ;
  input \sport1_txctl_Bcnt_reg[2]/NET0131  ;
  input \sport1_txctl_Bcnt_reg[3]/NET0131  ;
  input \sport1_txctl_Bcnt_reg[4]/NET0131  ;
  input \sport1_txctl_SP_EN_D1_reg/P0001  ;
  input \sport1_txctl_TCS_reg[0]/NET0131  ;
  input \sport1_txctl_TCS_reg[1]/NET0131  ;
  input \sport1_txctl_TCS_reg[2]/NET0131  ;
  input \sport1_txctl_TSreq_reg/NET0131  ;
  input \sport1_txctl_TSreqi_reg/NET0131  ;
  input \sport1_txctl_TXSHT_reg[0]/P0001  ;
  input \sport1_txctl_TXSHT_reg[10]/P0001  ;
  input \sport1_txctl_TXSHT_reg[11]/P0001  ;
  input \sport1_txctl_TXSHT_reg[12]/P0001  ;
  input \sport1_txctl_TXSHT_reg[13]/P0001  ;
  input \sport1_txctl_TXSHT_reg[14]/P0001  ;
  input \sport1_txctl_TXSHT_reg[15]/P0001  ;
  input \sport1_txctl_TXSHT_reg[1]/P0001  ;
  input \sport1_txctl_TXSHT_reg[2]/P0001  ;
  input \sport1_txctl_TXSHT_reg[3]/P0001  ;
  input \sport1_txctl_TXSHT_reg[4]/P0001  ;
  input \sport1_txctl_TXSHT_reg[5]/P0001  ;
  input \sport1_txctl_TXSHT_reg[6]/P0001  ;
  input \sport1_txctl_TXSHT_reg[7]/P0001  ;
  input \sport1_txctl_TXSHT_reg[8]/P0001  ;
  input \sport1_txctl_TXSHT_reg[9]/P0001  ;
  input \sport1_txctl_TX_reg[0]/P0001  ;
  input \sport1_txctl_TX_reg[10]/P0001  ;
  input \sport1_txctl_TX_reg[11]/P0001  ;
  input \sport1_txctl_TX_reg[12]/P0001  ;
  input \sport1_txctl_TX_reg[13]/P0001  ;
  input \sport1_txctl_TX_reg[14]/P0001  ;
  input \sport1_txctl_TX_reg[15]/P0001  ;
  input \sport1_txctl_TX_reg[1]/P0001  ;
  input \sport1_txctl_TX_reg[2]/P0001  ;
  input \sport1_txctl_TX_reg[3]/P0001  ;
  input \sport1_txctl_TX_reg[4]/P0001  ;
  input \sport1_txctl_TX_reg[5]/P0001  ;
  input \sport1_txctl_TX_reg[6]/P0001  ;
  input \sport1_txctl_TX_reg[7]/P0001  ;
  input \sport1_txctl_TX_reg[8]/P0001  ;
  input \sport1_txctl_TX_reg[9]/P0001  ;
  input \sport1_txctl_Wcnt_reg[0]/NET0131  ;
  input \sport1_txctl_Wcnt_reg[1]/NET0131  ;
  input \sport1_txctl_Wcnt_reg[2]/NET0131  ;
  input \sport1_txctl_Wcnt_reg[3]/NET0131  ;
  input \sport1_txctl_Wcnt_reg[4]/NET0131  ;
  input \sport1_txctl_Wcnt_reg[5]/NET0131  ;
  input \sport1_txctl_Wcnt_reg[6]/NET0131  ;
  input \sport1_txctl_Wcnt_reg[7]/NET0131  ;
  input \sport1_txctl_c_sync1_reg/P0001  ;
  input \sport1_txctl_c_sync2_reg/P0001  ;
  input \tm_MSTAT5_syn_reg/NET0131  ;
  input \tm_TCR_TMP_reg[0]/NET0131  ;
  input \tm_TCR_TMP_reg[10]/NET0131  ;
  input \tm_TCR_TMP_reg[11]/NET0131  ;
  input \tm_TCR_TMP_reg[12]/NET0131  ;
  input \tm_TCR_TMP_reg[13]/NET0131  ;
  input \tm_TCR_TMP_reg[14]/NET0131  ;
  input \tm_TCR_TMP_reg[15]/NET0131  ;
  input \tm_TCR_TMP_reg[1]/NET0131  ;
  input \tm_TCR_TMP_reg[2]/NET0131  ;
  input \tm_TCR_TMP_reg[3]/NET0131  ;
  input \tm_TCR_TMP_reg[4]/NET0131  ;
  input \tm_TCR_TMP_reg[5]/NET0131  ;
  input \tm_TCR_TMP_reg[6]/NET0131  ;
  input \tm_TCR_TMP_reg[7]/NET0131  ;
  input \tm_TCR_TMP_reg[8]/NET0131  ;
  input \tm_TCR_TMP_reg[9]/NET0131  ;
  input \tm_TINT_GEN1_reg/NET0131  ;
  input \tm_TINT_GEN2_reg/NET0131  ;
  input \tm_TSR_TMP_reg[0]/NET0131  ;
  input \tm_TSR_TMP_reg[1]/NET0131  ;
  input \tm_TSR_TMP_reg[2]/NET0131  ;
  input \tm_TSR_TMP_reg[3]/NET0131  ;
  input \tm_TSR_TMP_reg[4]/NET0131  ;
  input \tm_TSR_TMP_reg[5]/NET0131  ;
  input \tm_TSR_TMP_reg[6]/NET0131  ;
  input \tm_TSR_TMP_reg[7]/NET0131  ;
  input \tm_WR_TCR_KEEP_TO_TMCLK_p_reg/NET0131  ;
  input \tm_WR_TCR_TMP_GEN1_reg/P0001  ;
  input \tm_WR_TCR_TMP_GEN2_reg/P0001  ;
  input \tm_WR_TCR_p_reg/P0001  ;
  input \tm_WR_TSR_KEEP_TO_TMCLK_p_reg/NET0131  ;
  input \tm_WR_TSR_TMP_GEN1_reg/P0001  ;
  input \tm_WR_TSR_TMP_GEN2_reg/P0001  ;
  input \tm_WR_TSR_p_reg/P0001  ;
  input \tm_tcr_reg_DO_reg[0]/NET0131  ;
  input \tm_tcr_reg_DO_reg[10]/NET0131  ;
  input \tm_tcr_reg_DO_reg[11]/NET0131  ;
  input \tm_tcr_reg_DO_reg[12]/NET0131  ;
  input \tm_tcr_reg_DO_reg[13]/NET0131  ;
  input \tm_tcr_reg_DO_reg[14]/NET0131  ;
  input \tm_tcr_reg_DO_reg[15]/NET0131  ;
  input \tm_tcr_reg_DO_reg[1]/NET0131  ;
  input \tm_tcr_reg_DO_reg[2]/NET0131  ;
  input \tm_tcr_reg_DO_reg[3]/NET0131  ;
  input \tm_tcr_reg_DO_reg[4]/NET0131  ;
  input \tm_tcr_reg_DO_reg[5]/NET0131  ;
  input \tm_tcr_reg_DO_reg[6]/NET0131  ;
  input \tm_tcr_reg_DO_reg[7]/NET0131  ;
  input \tm_tcr_reg_DO_reg[8]/NET0131  ;
  input \tm_tcr_reg_DO_reg[9]/NET0131  ;
  input \tm_tpr_reg_DO_reg[0]/NET0131  ;
  input \tm_tpr_reg_DO_reg[10]/NET0131  ;
  input \tm_tpr_reg_DO_reg[11]/NET0131  ;
  input \tm_tpr_reg_DO_reg[12]/NET0131  ;
  input \tm_tpr_reg_DO_reg[13]/NET0131  ;
  input \tm_tpr_reg_DO_reg[14]/NET0131  ;
  input \tm_tpr_reg_DO_reg[15]/NET0131  ;
  input \tm_tpr_reg_DO_reg[1]/NET0131  ;
  input \tm_tpr_reg_DO_reg[2]/NET0131  ;
  input \tm_tpr_reg_DO_reg[3]/NET0131  ;
  input \tm_tpr_reg_DO_reg[4]/NET0131  ;
  input \tm_tpr_reg_DO_reg[5]/NET0131  ;
  input \tm_tpr_reg_DO_reg[6]/NET0131  ;
  input \tm_tpr_reg_DO_reg[7]/NET0131  ;
  input \tm_tpr_reg_DO_reg[8]/NET0131  ;
  input \tm_tpr_reg_DO_reg[9]/NET0131  ;
  input \tm_tsr_reg_DO_reg[0]/NET0131  ;
  input \tm_tsr_reg_DO_reg[1]/NET0131  ;
  input \tm_tsr_reg_DO_reg[2]/NET0131  ;
  input \tm_tsr_reg_DO_reg[3]/NET0131  ;
  input \tm_tsr_reg_DO_reg[4]/NET0131  ;
  input \tm_tsr_reg_DO_reg[5]/NET0131  ;
  input \tm_tsr_reg_DO_reg[6]/NET0131  ;
  input \tm_tsr_reg_DO_reg[7]/NET0131  ;
  input \tm_tsr_reg_DO_reg[8]/NET0131  ;
  output CLKO_pad ;
  output \CMAinx[0]_pad  ;
  output \CMAinx[10]_pad  ;
  output \CMAinx[11]_pad  ;
  output \CMAinx[1]_pad  ;
  output \CMAinx[2]_pad  ;
  output \CMAinx[3]_pad  ;
  output \CMAinx[4]_pad  ;
  output \CMAinx[5]_pad  ;
  output \CMAinx[6]_pad  ;
  output \CMAinx[7]_pad  ;
  output \CMAinx[8]_pad  ;
  output \CMAinx[9]_pad  ;
  output CMSn_pad ;
  output CM_cs_pad ;
  output \CM_wd[0]_pad  ;
  output \CM_wd[10]_pad  ;
  output \CM_wd[11]_pad  ;
  output \CM_wd[12]_pad  ;
  output \CM_wd[13]_pad  ;
  output \CM_wd[14]_pad  ;
  output \CM_wd[15]_pad  ;
  output \CM_wd[16]_pad  ;
  output \CM_wd[17]_pad  ;
  output \CM_wd[18]_pad  ;
  output \CM_wd[19]_pad  ;
  output \CM_wd[1]_pad  ;
  output \CM_wd[20]_pad  ;
  output \CM_wd[21]_pad  ;
  output \CM_wd[22]_pad  ;
  output \CM_wd[23]_pad  ;
  output \CM_wd[2]_pad  ;
  output \CM_wd[3]_pad  ;
  output \CM_wd[4]_pad  ;
  output \CM_wd[5]_pad  ;
  output \CM_wd[6]_pad  ;
  output \CM_wd[7]_pad  ;
  output \CM_wd[8]_pad  ;
  output \CM_wd[9]_pad  ;
  output CM_web_pad ;
  output \CMo_cs0_pad  ;
  output \CMo_cs1_pad  ;
  output \CMo_cs2_pad  ;
  output \CMo_cs3_pad  ;
  output \CMo_cs4_pad  ;
  output \CMo_cs5_pad  ;
  output \CMo_cs6_pad  ;
  output \CMo_cs7_pad  ;
  output \DMAinx[0]_pad  ;
  output \DMAinx[10]_pad  ;
  output \DMAinx[11]_pad  ;
  output \DMAinx[12]_pad  ;
  output \DMAinx[13]_pad  ;
  output \DMAinx[1]_pad  ;
  output \DMAinx[2]_pad  ;
  output \DMAinx[3]_pad  ;
  output \DMAinx[4]_pad  ;
  output \DMAinx[5]_pad  ;
  output \DMAinx[6]_pad  ;
  output \DMAinx[7]_pad  ;
  output \DMAinx[8]_pad  ;
  output \DMAinx[9]_pad  ;
  output DMSn_pad ;
  output DM_cs_pad ;
  output \DM_wd[0]_pad  ;
  output \DM_wd[10]_pad  ;
  output \DM_wd[11]_pad  ;
  output \DM_wd[12]_pad  ;
  output \DM_wd[13]_pad  ;
  output \DM_wd[14]_pad  ;
  output \DM_wd[15]_pad  ;
  output \DM_wd[1]_pad  ;
  output \DM_wd[2]_pad  ;
  output \DM_wd[3]_pad  ;
  output \DM_wd[4]_pad  ;
  output \DM_wd[5]_pad  ;
  output \DM_wd[6]_pad  ;
  output \DM_wd[7]_pad  ;
  output \DM_wd[8]_pad  ;
  output \DM_wd[9]_pad  ;
  output \DMo_cs0_pad  ;
  output \DMo_cs1_pad  ;
  output \DMo_cs2_pad  ;
  output \DMo_cs3_pad  ;
  output \DMo_cs4_pad  ;
  output \DMo_cs5_pad  ;
  output \DMo_cs6_pad  ;
  output \DMo_cs7_pad  ;
  output \DSPCLK_cm1_pad  ;
  output \EA_do[0]_pad  ;
  output \EA_do[10]_pad  ;
  output \EA_do[12]_pad  ;
  output \EA_do[13]_pad  ;
  output \EA_do[14]_pad  ;
  output \EA_do[1]_pad  ;
  output \EA_do[2]_pad  ;
  output \EA_do[3]_pad  ;
  output \EA_do[4]_pad  ;
  output \EA_do[5]_pad  ;
  output \EA_do[6]_pad  ;
  output \EA_do[7]_pad  ;
  output \EA_do[8]_pad  ;
  output \EA_do[9]_pad  ;
  output EA_oe_pad ;
  output \ED_do[0]_pad  ;
  output \ED_do[10]_pad  ;
  output \ED_do[11]_pad  ;
  output \ED_do[12]_pad  ;
  output \ED_do[13]_pad  ;
  output \ED_do[14]_pad  ;
  output \ED_do[15]_pad  ;
  output \ED_do[1]_pad  ;
  output \ED_do[2]_pad  ;
  output \ED_do[3]_pad  ;
  output \ED_do[4]_pad  ;
  output \ED_do[5]_pad  ;
  output \ED_do[6]_pad  ;
  output \ED_do[7]_pad  ;
  output \ED_do[8]_pad  ;
  output \ED_do[9]_pad  ;
  output \ED_oe_14_8_pad  ;
  output \ED_oe_7_0_pad  ;
  output \IAD_do[0]_pad  ;
  output \IAD_do[10]_pad  ;
  output \IAD_do[11]_pad  ;
  output \IAD_do[12]_pad  ;
  output \IAD_do[13]_pad  ;
  output \IAD_do[14]_pad  ;
  output \IAD_do[15]_pad  ;
  output \IAD_do[1]_pad  ;
  output \IAD_do[2]_pad  ;
  output \IAD_do[3]_pad  ;
  output \IAD_do[4]_pad  ;
  output \IAD_do[5]_pad  ;
  output \IAD_do[6]_pad  ;
  output \IAD_do[7]_pad  ;
  output \IAD_do[8]_pad  ;
  output \IAD_do[9]_pad  ;
  output IAD_oe_pad ;
  output IDoe_pad ;
  output IOSn_pad ;
  output \PMAinx[0]_pad  ;
  output \PMAinx[10]_pad  ;
  output \PMAinx[11]_pad  ;
  output \PMAinx[1]_pad  ;
  output \PMAinx[2]_pad  ;
  output \PMAinx[3]_pad  ;
  output \PMAinx[4]_pad  ;
  output \PMAinx[5]_pad  ;
  output \PMAinx[6]_pad  ;
  output \PMAinx[7]_pad  ;
  output \PMAinx[8]_pad  ;
  output \PMAinx[9]_pad  ;
  output \PM_wd[0]_pad  ;
  output \PM_wd[10]_pad  ;
  output \PM_wd[11]_pad  ;
  output \PM_wd[12]_pad  ;
  output \PM_wd[13]_pad  ;
  output \PM_wd[14]_pad  ;
  output \PM_wd[15]_pad  ;
  output \PM_wd[1]_pad  ;
  output \PM_wd[2]_pad  ;
  output \PM_wd[3]_pad  ;
  output \PM_wd[4]_pad  ;
  output \PM_wd[5]_pad  ;
  output \PM_wd[6]_pad  ;
  output \PM_wd[7]_pad  ;
  output \PM_wd[8]_pad  ;
  output \PM_wd[9]_pad  ;
  output \PMo_cs0_pad  ;
  output \PMo_cs1_pad  ;
  output \PMo_cs2_pad  ;
  output \PMo_cs3_pad  ;
  output \PMo_cs4_pad  ;
  output \PMo_cs5_pad  ;
  output \PMo_cs6_pad  ;
  output \PMo_cs7_pad  ;
  output \PMo_oe0_pad  ;
  output \RFS0_pad  ;
  output \RFS1_pad  ;
  output \SCLK0_pad  ;
  output \SCLK1_pad  ;
  output \TD0_pad  ;
  output \TD1_pad  ;
  output \TFS0_pad  ;
  output \TFS1_pad  ;
  output \T_ISn_syn_2  ;
  output WRn_pad ;
  output XTALoffn_pad ;
  output \_al_n0  ;
  output \bdma_BDMA_boot_reg/NET0131_reg_syn_3  ;
  output \bdma_BDMA_boot_reg/n0  ;
  output \bdma_BM_cyc_reg/P0000  ;
  output \bdma_BWCOUNT_reg[5]/NET0131_reg_syn_3  ;
  output \core_c_psq_MGNT_reg/P0001  ;
  output \core_c_psq_cntstk_cnts4x14_CNTcell_reg[0][5]/P0001_reg_syn_3  ;
  output \core_c_psq_cntstk_cnts4x14_CNTcell_reg[1][5]/P0001_reg_syn_3  ;
  output \core_c_psq_cntstk_cnts4x14_CNTcell_reg[2][5]/P0001_reg_syn_3  ;
  output \core_c_psq_cntstk_cnts4x14_CNTcell_reg[3][5]/P0001_reg_syn_3  ;
  output \core_eu_ea_alu_ea_reg_afrwe_DO_reg[12]/P0001_reg_syn_3  ;
  output \core_eu_ea_alu_ea_reg_afrwe_DO_reg[14]/P0001_reg_syn_3  ;
  output \core_eu_ea_alu_ea_reg_afrwe_DO_reg[1]/P0001_reg_syn_3  ;
  output \core_eu_ea_alu_ea_reg_afrwe_DO_reg[2]/P0001_reg_syn_3  ;
  output \core_eu_ea_alu_ea_reg_afrwe_DO_reg[4]/P0001_reg_syn_3  ;
  output \core_eu_ea_alu_ea_reg_afrwe_DO_reg[6]/P0001_reg_syn_3  ;
  output \core_eu_ea_alu_ea_reg_afrwe_DO_reg[9]/P0001_reg_syn_3  ;
  output \core_eu_ea_alu_ea_reg_afswe_DO_reg[12]/P0001_reg_syn_3  ;
  output \core_eu_ea_alu_ea_reg_afswe_DO_reg[14]/P0001_reg_syn_3  ;
  output \core_eu_ea_alu_ea_reg_afswe_DO_reg[1]/P0001_reg_syn_3  ;
  output \core_eu_ea_alu_ea_reg_afswe_DO_reg[2]/P0001_reg_syn_3  ;
  output \core_eu_ea_alu_ea_reg_afswe_DO_reg[4]/P0001_reg_syn_3  ;
  output \core_eu_ea_alu_ea_reg_afswe_DO_reg[6]/P0001_reg_syn_3  ;
  output \core_eu_ea_alu_ea_reg_afswe_DO_reg[9]/P0001_reg_syn_3  ;
  output \core_eu_ec_cun_MVi_pre_C_reg/P0001_reg_syn_3  ;
  output \core_eu_em_mac_em_reg_Sq_E_reg/P0001_reg_syn_3  ;
  output \emc_DMDreg_reg[8]/P0001_reg_syn_3  ;
  output \emc_DMDreg_reg[9]/P0001_reg_syn_3  ;
  output \emc_ECMcs_reg/P0001  ;
  output \emc_PMDreg_reg[8]/P0001_reg_syn_3  ;
  output \emc_PMDreg_reg[9]/P0001_reg_syn_3  ;
  output \g10/_0_  ;
  output \g1000/_0_  ;
  output \g10000/_0_  ;
  output \g10001/_0_  ;
  output \g10002/_0_  ;
  output \g10003/_0_  ;
  output \g10004/_0_  ;
  output \g10005/_0_  ;
  output \g10007/_0_  ;
  output \g10008/_0_  ;
  output \g10009/_0_  ;
  output \g1001/_3_  ;
  output \g10010/_0_  ;
  output \g10011/_0_  ;
  output \g10012/_0_  ;
  output \g10013/_0_  ;
  output \g10014/_0_  ;
  output \g10015/_0_  ;
  output \g10016/_0_  ;
  output \g10017/_0_  ;
  output \g10018/_0_  ;
  output \g10019/_0_  ;
  output \g1002/_3_  ;
  output \g10020/_0_  ;
  output \g10021/_0_  ;
  output \g10022/_0_  ;
  output \g10023/_0_  ;
  output \g10024/_0_  ;
  output \g10025/_0_  ;
  output \g10026/_0_  ;
  output \g10027/_0_  ;
  output \g10028/_0_  ;
  output \g10029/_0_  ;
  output \g1003/_0_  ;
  output \g10030/_0_  ;
  output \g10031/_0_  ;
  output \g10032/_0_  ;
  output \g10033/_0_  ;
  output \g10034/_0_  ;
  output \g10035/_0_  ;
  output \g10036/_0_  ;
  output \g10037/_0_  ;
  output \g10038/_0_  ;
  output \g10039/_0_  ;
  output \g10040/_0_  ;
  output \g10041/_0_  ;
  output \g10042/_0_  ;
  output \g10043/_0_  ;
  output \g10044/_0_  ;
  output \g10045/_0_  ;
  output \g10046/_0_  ;
  output \g10047/_0_  ;
  output \g10048/_0_  ;
  output \g10049/_0_  ;
  output \g10050/_0_  ;
  output \g10051/_0_  ;
  output \g10052/_0_  ;
  output \g10053/_0_  ;
  output \g10054/_0_  ;
  output \g10055/_0_  ;
  output \g10056/_0_  ;
  output \g10057/_0_  ;
  output \g10058/_0_  ;
  output \g10059/_0_  ;
  output \g10060/_0_  ;
  output \g10061/_0_  ;
  output \g10062/_0_  ;
  output \g10063/_0_  ;
  output \g10064/_0_  ;
  output \g10065/_0_  ;
  output \g10066/_0_  ;
  output \g10067/_0_  ;
  output \g10068/_0_  ;
  output \g10069/_0_  ;
  output \g10070/_0_  ;
  output \g10071/_0_  ;
  output \g10072/_0_  ;
  output \g10073/_0_  ;
  output \g10074/_0_  ;
  output \g10075/_0_  ;
  output \g10076/_0_  ;
  output \g10077/_0_  ;
  output \g10078/_0_  ;
  output \g10080/_0_  ;
  output \g10081/_0_  ;
  output \g10083/_0_  ;
  output \g10089/_0_  ;
  output \g1009/_0_  ;
  output \g10090/_0_  ;
  output \g10091/_0_  ;
  output \g10092/_0_  ;
  output \g10093/_0_  ;
  output \g10094/_0_  ;
  output \g1010/_0_  ;
  output \g10108/_3_  ;
  output \g1011/_0_  ;
  output \g10110/_0_  ;
  output \g10111/_0_  ;
  output \g10113/_3_  ;
  output \g10115/_3_  ;
  output \g1013/_0_  ;
  output \g1014/_0_  ;
  output \g10152/_0_  ;
  output \g10153/_0_  ;
  output \g10154/_0_  ;
  output \g10155/_0_  ;
  output \g10156/_0_  ;
  output \g10157/_0_  ;
  output \g10158/_0_  ;
  output \g10159/_0_  ;
  output \g1016/_0_  ;
  output \g10160/_0_  ;
  output \g10161/_0_  ;
  output \g10162/_0_  ;
  output \g10163/_0_  ;
  output \g10164/_0_  ;
  output \g10165/_0_  ;
  output \g1017/_0_  ;
  output \g10170/_3_  ;
  output \g1018/_0_  ;
  output \g10190/_3_  ;
  output \g10194/_3_  ;
  output \g10198/_0_  ;
  output \g10199/_0_  ;
  output \g102/_0_  ;
  output \g103/_0_  ;
  output \g104/_0_  ;
  output \g105/_0_  ;
  output \g10598/_0_  ;
  output \g106/_0_  ;
  output \g10667/_0_  ;
  output \g10683/_0_  ;
  output \g10685/_0_  ;
  output \g107/_0_  ;
  output \g10721/_0_  ;
  output \g10758/_0_  ;
  output \g10765/_0_  ;
  output \g10778/_0_  ;
  output \g10791/_0_  ;
  output \g108/_0_  ;
  output \g10887/_0_  ;
  output \g1089/_0_  ;
  output \g109/_0_  ;
  output \g1090/_0_  ;
  output \g1091/_0_  ;
  output \g1092/_0_  ;
  output \g10923/_0_  ;
  output \g1093/_0_  ;
  output \g10930/_0_  ;
  output \g10931/_0_  ;
  output \g10936/_0_  ;
  output \g1097/_0_  ;
  output \g11/_0_  ;
  output \g110/_0_  ;
  output \g1101/_0_  ;
  output \g11013/_0_  ;
  output \g1102/_0_  ;
  output \g1103/_0_  ;
  output \g11032/_0_  ;
  output \g1104/_0_  ;
  output \g1105/_0_  ;
  output \g1107/_0_  ;
  output \g11074/_0_  ;
  output \g11077/_0_  ;
  output \g1108/_0_  ;
  output \g1109/_0_  ;
  output \g11112/_0_  ;
  output \g11115/_0_  ;
  output \g11116/_0_  ;
  output \g11119/_0_  ;
  output \g11120/_0_  ;
  output \g1113/_0_  ;
  output \g1115/_0_  ;
  output \g1116/_0_  ;
  output \g1117/_0_  ;
  output \g11267/_0_  ;
  output \g11281/_0_  ;
  output \g11287/_0_  ;
  output \g11300/_0_  ;
  output \g11323/_0_  ;
  output \g11325/_2__syn_2  ;
  output \g11345/_2_  ;
  output \g11470/_0_  ;
  output \g11471/_0_  ;
  output \g11472/_0_  ;
  output \g11473/_0_  ;
  output \g11474/_0_  ;
  output \g11476/_0_  ;
  output \g11477/_0_  ;
  output \g11496/_0_  ;
  output \g11497/_0_  ;
  output \g11498/_0_  ;
  output \g11499/_0_  ;
  output \g11500/_0_  ;
  output \g11501/_0_  ;
  output \g11502/_0_  ;
  output \g11503/_0_  ;
  output \g11504/_0_  ;
  output \g11505/_0_  ;
  output \g11506/_0_  ;
  output \g11507/_0_  ;
  output \g11509/_0_  ;
  output \g11510/_0_  ;
  output \g11515/_0_  ;
  output \g11516/_0_  ;
  output \g11520/_0_  ;
  output \g11521/_0_  ;
  output \g11576/_0_  ;
  output \g11577/_0_  ;
  output \g11578/_0_  ;
  output \g11579/_0_  ;
  output \g11580/_0_  ;
  output \g11581/_0_  ;
  output \g11582/_0_  ;
  output \g11583/_0_  ;
  output \g11584/_0_  ;
  output \g11585/_0_  ;
  output \g11586/_0_  ;
  output \g11587/_0_  ;
  output \g11588/_0_  ;
  output \g11589/_0_  ;
  output \g11591/_0_  ;
  output \g11593/_0_  ;
  output \g11595/_0_  ;
  output \g11596/_0_  ;
  output \g11597/_0_  ;
  output \g11605/_0_  ;
  output \g11606/_0_  ;
  output \g11607/_0_  ;
  output \g11608/_0_  ;
  output \g11609/_0_  ;
  output \g11610/_0_  ;
  output \g11611/_0_  ;
  output \g11612/_0_  ;
  output \g11613/_0_  ;
  output \g11615/_0_  ;
  output \g11616/_0_  ;
  output \g11617/_0_  ;
  output \g11651/_3_  ;
  output \g11704/_0_  ;
  output \g11705/_0_  ;
  output \g11709/_0_  ;
  output \g11722/_0_  ;
  output \g11723/_0_  ;
  output \g119/_0_  ;
  output \g1192/_0_  ;
  output \g11994/_0_  ;
  output \g120/_0_  ;
  output \g1200/_0_  ;
  output \g12003/_0_  ;
  output \g1201/_0_  ;
  output \g12019/_0_  ;
  output \g1203/_3_  ;
  output \g1204/_3_  ;
  output \g1207/_0_  ;
  output \g1208/_0_  ;
  output \g12092/_0_  ;
  output \g1210/_0_  ;
  output \g1211/_0_  ;
  output \g1212/_0_  ;
  output \g1213/_0_  ;
  output \g12145/_0_  ;
  output \g12155/_0_  ;
  output \g12186/_0_  ;
  output \g12187/_0_  ;
  output \g12192/_0_  ;
  output \g12201/_0_  ;
  output \g12202/_0_  ;
  output \g12203/_0_  ;
  output \g12204/_0_  ;
  output \g12207/_0_  ;
  output \g12229/_3_  ;
  output \g12267/_0_  ;
  output \g12276/_0_  ;
  output \g12278/_0_  ;
  output \g12279/_0_  ;
  output \g12280/_0_  ;
  output \g12302/_0_  ;
  output \g12316/_0_  ;
  output \g12317/_0_  ;
  output \g12319/_0_  ;
  output \g12328/_3_  ;
  output \g1233/_0_  ;
  output \g12348/_0_  ;
  output \g12351/_0_  ;
  output \g12352/_0_  ;
  output \g12353/_0_  ;
  output \g12354/_0_  ;
  output \g12355/_0_  ;
  output \g1237/_0_  ;
  output \g124/_0_  ;
  output \g12444/_0_  ;
  output \g125/_0_  ;
  output \g12637/_0_  ;
  output \g12639/_0_  ;
  output \g12658/_0_  ;
  output \g12659/_0_  ;
  output \g12660/_0_  ;
  output \g12663/_0_  ;
  output \g12664/_0_  ;
  output \g12665/_0_  ;
  output \g12672/_3_  ;
  output \g12673/_3_  ;
  output \g12674/_3_  ;
  output \g12675/_3_  ;
  output \g12676/_3_  ;
  output \g12677/_3_  ;
  output \g12678/_0_  ;
  output \g12679/_3_  ;
  output \g12697/_3_  ;
  output \g12701/_3_  ;
  output \g12711/_2_  ;
  output \g12713/_2_  ;
  output \g12715/_2_  ;
  output \g12717/_2_  ;
  output \g12718/_2__syn_2  ;
  output \g1272/_0_  ;
  output \g12728/_1__syn_2  ;
  output \g12730/_3_  ;
  output \g12741/_1__syn_2  ;
  output \g12746/_0__syn_2  ;
  output \g12748/_0_  ;
  output \g12749/_0_  ;
  output \g12759/_1__syn_2  ;
  output \g12760/_0_  ;
  output \g12762/_0_  ;
  output \g12763/_0_  ;
  output \g12764/_0_  ;
  output \g12765/_0_  ;
  output \g12766/_0_  ;
  output \g12767/_0_  ;
  output \g12768/_0_  ;
  output \g12769/_0_  ;
  output \g12770/_0_  ;
  output \g12771/_0_  ;
  output \g12772/_0_  ;
  output \g12773/_0_  ;
  output \g12774/_0_  ;
  output \g12775/_0_  ;
  output \g12776/_0_  ;
  output \g12777/_0_  ;
  output \g12778/_0_  ;
  output \g12779/_0_  ;
  output \g1278/_0_  ;
  output \g12780/_0_  ;
  output \g12781/_0_  ;
  output \g12782/_0_  ;
  output \g12783/_0_  ;
  output \g12784/_0_  ;
  output \g12785/_0_  ;
  output \g12786/_0_  ;
  output \g12787/_0_  ;
  output \g12788/_0_  ;
  output \g12789/_0_  ;
  output \g12790/_0_  ;
  output \g12791/_0_  ;
  output \g12792/_0_  ;
  output \g12793/_0_  ;
  output \g12794/_0_  ;
  output \g12795/_0_  ;
  output \g12796/_0_  ;
  output \g12797/_0_  ;
  output \g12798/_0_  ;
  output \g12799/_0_  ;
  output \g12800/_0_  ;
  output \g12801/_0_  ;
  output \g12802/_0_  ;
  output \g12803/_0_  ;
  output \g12804/_0_  ;
  output \g12805/_0_  ;
  output \g12806/_0_  ;
  output \g12807/_0_  ;
  output \g12808/_0_  ;
  output \g12809/_0_  ;
  output \g1281/_0_  ;
  output \g12810/_0_  ;
  output \g12811/_0_  ;
  output \g12812/_0_  ;
  output \g12813/_0_  ;
  output \g12814/_0_  ;
  output \g12815/_0_  ;
  output \g12816/_0_  ;
  output \g12817/_0_  ;
  output \g12818/_0_  ;
  output \g12819/_0_  ;
  output \g1282/_0_  ;
  output \g12820/_0_  ;
  output \g12821/_0_  ;
  output \g12822/_0_  ;
  output \g12823/_0_  ;
  output \g12824/_0_  ;
  output \g12825/_0_  ;
  output \g12826/_0_  ;
  output \g12827/_0_  ;
  output \g12828/_0_  ;
  output \g12829/_0_  ;
  output \g12830/_0_  ;
  output \g12831/_0_  ;
  output \g12832/_0_  ;
  output \g12833/_0_  ;
  output \g12835/_0_  ;
  output \g12836/_0_  ;
  output \g12838/_0_  ;
  output \g12848/_0_  ;
  output \g12849/_0_  ;
  output \g1285/_0_  ;
  output \g12850/_0_  ;
  output \g12857/_0_  ;
  output \g12858/_0_  ;
  output \g12859/_0_  ;
  output \g12861/_0_  ;
  output \g12862/_0_  ;
  output \g12868/_0_  ;
  output \g12869/_0_  ;
  output \g1287/_0_  ;
  output \g12870/_0_  ;
  output \g12871/_0_  ;
  output \g12872/_0_  ;
  output \g12873/_0_  ;
  output \g12874/_0_  ;
  output \g12875/_0_  ;
  output \g12876/_0_  ;
  output \g12877/_0_  ;
  output \g12878/_0_  ;
  output \g12879/_0_  ;
  output \g12880/_0_  ;
  output \g12881/_0_  ;
  output \g12882/_0_  ;
  output \g12883/_0_  ;
  output \g12884/_0_  ;
  output \g12885/_0_  ;
  output \g12886/_0_  ;
  output \g12887/_0_  ;
  output \g12888/_0_  ;
  output \g12889/_0_  ;
  output \g1289/_0_  ;
  output \g12890/_0_  ;
  output \g12891/_0_  ;
  output \g12894/_0_  ;
  output \g12898/_0_  ;
  output \g12899/_0_  ;
  output \g12900/_0_  ;
  output \g12901/_0_  ;
  output \g12902/_0_  ;
  output \g12903/_0_  ;
  output \g12906/_0_  ;
  output \g12907/_0_  ;
  output \g12908/_0_  ;
  output \g12912/_0_  ;
  output \g12913/_0_  ;
  output \g12914/_0_  ;
  output \g12915/_0_  ;
  output \g12916/_0_  ;
  output \g12917/_0_  ;
  output \g12918/_0_  ;
  output \g12919/_0_  ;
  output \g12920/_0_  ;
  output \g12921/_0_  ;
  output \g12922/_0_  ;
  output \g12923/_0_  ;
  output \g12924/_0_  ;
  output \g12925/_0_  ;
  output \g12926/_0_  ;
  output \g12932/_0_  ;
  output \g12933/_0_  ;
  output \g12936/_0_  ;
  output \g12955/_0_  ;
  output \g13015/_0_  ;
  output \g13016/_0_  ;
  output \g13017/_0_  ;
  output \g13018/_0_  ;
  output \g13019/_0_  ;
  output \g13020/_0_  ;
  output \g13021/_0_  ;
  output \g13024/_0_  ;
  output \g13025/_0_  ;
  output \g13027/_0_  ;
  output \g13028/_0_  ;
  output \g13030/_0_  ;
  output \g13031/_0_  ;
  output \g13033/_0_  ;
  output \g13047/_0_  ;
  output \g13060/_0_  ;
  output \g13062/_0_  ;
  output \g13063/_0_  ;
  output \g13064/_0_  ;
  output \g13067/_0_  ;
  output \g13068/_0_  ;
  output \g13069/_0_  ;
  output \g13070/_0_  ;
  output \g13072/_0_  ;
  output \g13094/_0_  ;
  output \g13104/_0_  ;
  output \g13110/_0_  ;
  output \g13114/_0_  ;
  output \g13115/_0_  ;
  output \g13116/_0_  ;
  output \g13117/_0_  ;
  output \g13118/_0_  ;
  output \g13119/_0_  ;
  output \g13120/_0_  ;
  output \g13121/_0_  ;
  output \g13124/_0_  ;
  output \g13125/_0_  ;
  output \g13127/_0_  ;
  output \g13128/_0_  ;
  output \g13129/_0_  ;
  output \g13130/_0_  ;
  output \g13131/_0_  ;
  output \g13132/_0_  ;
  output \g13133/_0_  ;
  output \g13134/_0_  ;
  output \g13138/_0_  ;
  output \g13139/_0_  ;
  output \g13140/_0_  ;
  output \g13141/_0_  ;
  output \g13142/_0_  ;
  output \g13143/_0_  ;
  output \g13144/_0_  ;
  output \g13146/_0_  ;
  output \g13150/_0_  ;
  output \g13152/_0_  ;
  output \g13154/_0_  ;
  output \g13155/_0_  ;
  output \g13156/_0_  ;
  output \g13157/_0_  ;
  output \g13158/_0_  ;
  output \g1320/_3_  ;
  output \g13266/_0_  ;
  output \g13269/_0_  ;
  output \g13274/_0_  ;
  output \g13277/_0_  ;
  output \g13280/_0_  ;
  output \g13283/_0_  ;
  output \g13294/_0_  ;
  output \g13330/_0_  ;
  output \g13333/_0_  ;
  output \g13334/_0_  ;
  output \g13335/_0_  ;
  output \g13336/_0_  ;
  output \g13337/_0_  ;
  output \g13338/_0_  ;
  output \g13345/_0_  ;
  output \g13346/_0_  ;
  output \g13347/_0_  ;
  output \g13348/_0_  ;
  output \g13349/_0_  ;
  output \g13350/_0_  ;
  output \g13351/_0_  ;
  output \g13352/_0_  ;
  output \g13486/_0_  ;
  output \g13488/_0_  ;
  output \g13508/_0_  ;
  output \g13509/_0_  ;
  output \g13510/_0_  ;
  output \g13511/_0_  ;
  output \g13512/_0_  ;
  output \g13513/_0_  ;
  output \g13514/_0_  ;
  output \g13515/_0_  ;
  output \g13516/_0_  ;
  output \g13517/_0_  ;
  output \g13518/_0_  ;
  output \g13519/_0_  ;
  output \g13520/_0_  ;
  output \g13521/_0_  ;
  output \g13540/_0_  ;
  output \g13541/_0_  ;
  output \g13542/_0_  ;
  output \g13543/_0_  ;
  output \g13544/_0_  ;
  output \g13545/_0_  ;
  output \g13546/_0_  ;
  output \g13547/_0_  ;
  output \g13548/_0_  ;
  output \g13549/_0_  ;
  output \g13550/_0_  ;
  output \g13551/_0_  ;
  output \g13552/_0_  ;
  output \g13553/_0_  ;
  output \g13554/_0_  ;
  output \g13555/_0_  ;
  output \g13556/_0_  ;
  output \g13557/_0_  ;
  output \g13558/_0_  ;
  output \g13559/_0_  ;
  output \g13560/_0_  ;
  output \g13561/_0_  ;
  output \g13562/_0_  ;
  output \g13563/_0_  ;
  output \g13564/_0_  ;
  output \g13565/_0_  ;
  output \g13566/_0_  ;
  output \g13567/_0_  ;
  output \g13568/_0_  ;
  output \g13569/_0_  ;
  output \g13570/_0_  ;
  output \g13571/_0_  ;
  output \g13572/_0_  ;
  output \g137/_3_  ;
  output \g1387/_3_  ;
  output \g1388/_3_  ;
  output \g1389/_0_  ;
  output \g139/_0_  ;
  output \g1390/_0_  ;
  output \g1393/_0_  ;
  output \g140/_0_  ;
  output \g141/_0_  ;
  output \g14173/_0_  ;
  output \g14176/_0_  ;
  output \g142/_3_  ;
  output \g14273/_1__syn_2  ;
  output \g14274/_0_  ;
  output \g14280/_0_  ;
  output \g14281/_0_  ;
  output \g143/_3_  ;
  output \g14354/_3__syn_2  ;
  output \g14370/_0_  ;
  output \g14385/_0_  ;
  output \g14386/_0_  ;
  output \g144/_3_  ;
  output \g14407/_0_  ;
  output \g14412/_0_  ;
  output \g14435/_0_  ;
  output \g14439/_0_  ;
  output \g145/_0_  ;
  output \g14522/_0_  ;
  output \g14528/_0_  ;
  output \g14533/_0_  ;
  output \g14581/_1_  ;
  output \g14582/_0_  ;
  output \g146/_3_  ;
  output \g14671/_0_  ;
  output \g14672/_0_  ;
  output \g147/_0_  ;
  output \g1473/_0_  ;
  output \g148/_0_  ;
  output \g14826/_0_  ;
  output \g149/_0_  ;
  output \g14908/_0_  ;
  output \g14911/_0_  ;
  output \g14936/_2_  ;
  output \g1494/_0_  ;
  output \g1495/_0_  ;
  output \g14950/_2_  ;
  output \g14953/_2_  ;
  output \g15003/_0_  ;
  output \g15004/_0_  ;
  output \g15006/_0_  ;
  output \g15007/_0_  ;
  output \g15008/_0_  ;
  output \g15009/_0_  ;
  output \g15010/_0_  ;
  output \g15011/_0_  ;
  output \g15012/_0_  ;
  output \g15013/_0_  ;
  output \g15014/_0_  ;
  output \g15015/_0_  ;
  output \g15016/_0_  ;
  output \g15017/_0_  ;
  output \g15018/_0_  ;
  output \g15019/_0_  ;
  output \g15035/_0_  ;
  output \g15036/_0_  ;
  output \g15038/_0_  ;
  output \g15039/_0_  ;
  output \g15040/_0_  ;
  output \g15041/_0_  ;
  output \g15042/_0_  ;
  output \g15043/_0_  ;
  output \g15044/_0_  ;
  output \g15045/_0_  ;
  output \g15046/_0_  ;
  output \g15056/_00_  ;
  output \g151/_0_  ;
  output \g15193/_0_  ;
  output \g152/_0_  ;
  output \g15256/_0_  ;
  output \g153/_0_  ;
  output \g15393/_0_  ;
  output \g15394/_0_  ;
  output \g15395/_0_  ;
  output \g15396/_0_  ;
  output \g15397/_0_  ;
  output \g15398/_0_  ;
  output \g15399/_0_  ;
  output \g154/_0_  ;
  output \g15400/_0_  ;
  output \g15401/_0_  ;
  output \g15402/_0_  ;
  output \g15403/_0_  ;
  output \g15404/_0_  ;
  output \g15405/_0_  ;
  output \g15406/_0_  ;
  output \g15407/_0_  ;
  output \g15408/_0_  ;
  output \g15473/_0_  ;
  output \g15650/_0_  ;
  output \g15651/_0_  ;
  output \g15652/_0_  ;
  output \g15653/_0_  ;
  output \g15662/_0_  ;
  output \g15663/_0_  ;
  output \g15664/_0_  ;
  output \g15665/_0_  ;
  output \g15666/_0_  ;
  output \g15667/_0_  ;
  output \g15668/_0_  ;
  output \g15669/_0_  ;
  output \g15670/_0_  ;
  output \g15671/_0_  ;
  output \g15672/_0_  ;
  output \g15673/_0_  ;
  output \g15674/_0_  ;
  output \g15675/_0_  ;
  output \g1569/_0_  ;
  output \g1570/_0_  ;
  output \g1575/_0_  ;
  output \g1576/_0_  ;
  output \g15922/_1_  ;
  output \g15970/_0_  ;
  output \g16059/_0_  ;
  output \g1606/_3_  ;
  output \g16124/_0_  ;
  output \g16144/_0_  ;
  output \g16202/_0_  ;
  output \g16214/_0_  ;
  output \g16247/_0_  ;
  output \g16257/_0_  ;
  output \g16274/_1_  ;
  output \g16324/_0_  ;
  output \g16343/_1__syn_2  ;
  output \g16381/_0_  ;
  output \g16383/_0_  ;
  output \g16386/_0_  ;
  output \g16414/_1__syn_2  ;
  output \g16416/_0__syn_2  ;
  output \g16448/_0_  ;
  output \g16460/_1_  ;
  output \g16625/_3_  ;
  output \g16662/_0_  ;
  output \g16668/_1__syn_2  ;
  output \g16692/_0_  ;
  output \g16721/_0_  ;
  output \g16723/_0_  ;
  output \g16725/_0_  ;
  output \g16726/_0_  ;
  output \g16727/_0_  ;
  output \g16728/_0_  ;
  output \g16729/_0_  ;
  output \g16730/_0_  ;
  output \g16731/_0_  ;
  output \g16732/_0_  ;
  output \g16733/_0_  ;
  output \g16734/_0_  ;
  output \g16735/_0_  ;
  output \g16736/_0_  ;
  output \g16737/_0_  ;
  output \g16738/_0_  ;
  output \g16739/_0_  ;
  output \g16740/_0_  ;
  output \g16741/_0_  ;
  output \g16742/_0_  ;
  output \g16743/_0_  ;
  output \g16747/_0_  ;
  output \g16748/_0_  ;
  output \g16749/_0_  ;
  output \g16750/_0_  ;
  output \g16753/_0_  ;
  output \g16754/_0_  ;
  output \g16755/_0_  ;
  output \g16756/_0_  ;
  output \g16757/_0_  ;
  output \g16758/_0_  ;
  output \g16761/_0_  ;
  output \g16765/_0_  ;
  output \g16766/_0_  ;
  output \g16767/_0_  ;
  output \g16768/_0_  ;
  output \g16769/_0_  ;
  output \g16772/_0_  ;
  output \g16785/_0_  ;
  output \g16786/_0_  ;
  output \g16787/_0_  ;
  output \g16788/_0_  ;
  output \g16789/_0_  ;
  output \g16790/_0_  ;
  output \g16791/_0_  ;
  output \g16804/_0_  ;
  output \g16805/_0_  ;
  output \g16806/_0_  ;
  output \g16807/_0_  ;
  output \g16808/_0_  ;
  output \g16809/_0_  ;
  output \g16810/_0_  ;
  output \g16811/_0_  ;
  output \g16812/_0_  ;
  output \g16813/_0_  ;
  output \g16814/_0_  ;
  output \g16815/_0_  ;
  output \g16816/_0_  ;
  output \g16817/_0_  ;
  output \g16819/_0_  ;
  output \g16822/_0_  ;
  output \g16823/_0_  ;
  output \g16824/_0_  ;
  output \g16825/_0_  ;
  output \g16828/_0_  ;
  output \g16829/_0_  ;
  output \g16830/_0_  ;
  output \g16831/_0_  ;
  output \g16832/_0_  ;
  output \g16833/_0_  ;
  output \g16834/_0_  ;
  output \g16835/_0_  ;
  output \g16836/_0_  ;
  output \g16837/_0_  ;
  output \g16840/_0_  ;
  output \g16841/_0_  ;
  output \g16842/_0_  ;
  output \g16843/_0_  ;
  output \g16846/_0_  ;
  output \g16847/_0_  ;
  output \g16848/_0_  ;
  output \g16849/_0_  ;
  output \g16850/_0_  ;
  output \g16851/_0_  ;
  output \g16852/_0_  ;
  output \g16853/_0_  ;
  output \g16854/_0_  ;
  output \g16855/_0_  ;
  output \g16856/_0_  ;
  output \g16857/_0_  ;
  output \g16859/_0_  ;
  output \g16862/_0_  ;
  output \g16865/_0_  ;
  output \g16866/_0_  ;
  output \g16867/_0_  ;
  output \g16868/_0_  ;
  output \g16869/_0_  ;
  output \g16870/_0_  ;
  output \g16871/_0_  ;
  output \g16872/_0_  ;
  output \g16873/_0_  ;
  output \g16874/_0_  ;
  output \g16875/_0_  ;
  output \g16876/_0_  ;
  output \g16877/_0_  ;
  output \g16878/_0_  ;
  output \g16879/_0_  ;
  output \g16880/_0_  ;
  output \g16881/_0_  ;
  output \g16882/_0_  ;
  output \g16884/_0_  ;
  output \g16887/_0_  ;
  output \g16891/_0_  ;
  output \g16892/_0_  ;
  output \g16893/_0_  ;
  output \g16894/_0_  ;
  output \g16895/_0_  ;
  output \g16897/_0_  ;
  output \g16898/_0_  ;
  output \g16899/_0_  ;
  output \g16900/_0_  ;
  output \g16901/_0_  ;
  output \g16902/_0_  ;
  output \g16903/_0_  ;
  output \g16904/_0_  ;
  output \g16905/_0_  ;
  output \g16906/_0_  ;
  output \g16907/_0_  ;
  output \g16908/_0_  ;
  output \g16909/_0_  ;
  output \g16910/_0_  ;
  output \g16912/_0_  ;
  output \g16914/_0_  ;
  output \g16915/_0_  ;
  output \g16950/_0_  ;
  output \g16951/_0_  ;
  output \g16952/_0_  ;
  output \g16953/_0_  ;
  output \g16954/_0_  ;
  output \g16955/_0_  ;
  output \g16956/_0_  ;
  output \g16957/_0_  ;
  output \g16958/_0_  ;
  output \g16959/_0_  ;
  output \g16960/_0_  ;
  output \g16961/_0_  ;
  output \g16962/_0_  ;
  output \g16963/_0_  ;
  output \g16964/_0_  ;
  output \g16965/_0_  ;
  output \g16966/_0_  ;
  output \g16967/_0_  ;
  output \g16968/_0_  ;
  output \g16970/_0_  ;
  output \g17102/_3_  ;
  output \g17106/_0_  ;
  output \g17107/_0_  ;
  output \g17109/_0_  ;
  output \g17110/_0_  ;
  output \g17111/_0_  ;
  output \g17112/_0_  ;
  output \g17115/_0_  ;
  output \g17116/_0_  ;
  output \g17119/_0_  ;
  output \g17120/_0_  ;
  output \g17122/_0_  ;
  output \g17123/_0_  ;
  output \g17124/_0_  ;
  output \g17125/_0_  ;
  output \g17126/_0_  ;
  output \g17127/_0_  ;
  output \g17128/_0_  ;
  output \g17130/_0_  ;
  output \g17131/_0_  ;
  output \g17132/_0_  ;
  output \g17133/_0_  ;
  output \g17134/_0_  ;
  output \g17135/_0_  ;
  output \g17136/_0_  ;
  output \g17137/_0_  ;
  output \g17138/_0_  ;
  output \g17140/_0_  ;
  output \g17141/_0_  ;
  output \g17142/_0_  ;
  output \g17143/_0_  ;
  output \g17144/_0_  ;
  output \g17145/_0_  ;
  output \g17146/_0_  ;
  output \g17147/_0_  ;
  output \g17148/_0_  ;
  output \g17149/_0_  ;
  output \g17150/_0_  ;
  output \g17151/_0_  ;
  output \g17152/_0_  ;
  output \g17153/_0_  ;
  output \g17154/_0_  ;
  output \g17155/_0_  ;
  output \g17157/_0_  ;
  output \g17159/_0_  ;
  output \g17160/_0_  ;
  output \g17161/_0_  ;
  output \g17162/_0_  ;
  output \g17163/_0_  ;
  output \g17164/_0_  ;
  output \g17165/_0_  ;
  output \g17166/_0_  ;
  output \g17168/_0_  ;
  output \g17171/_0_  ;
  output \g17173/_0_  ;
  output \g17177/_0_  ;
  output \g17178/_0_  ;
  output \g17179/_0_  ;
  output \g17180/_0_  ;
  output \g17182/_0_  ;
  output \g17183/_0_  ;
  output \g17184/_0_  ;
  output \g17185/_0_  ;
  output \g17186/_0_  ;
  output \g17188/_0_  ;
  output \g17189/_0_  ;
  output \g17190/_0_  ;
  output \g17191/_0_  ;
  output \g17193/_0_  ;
  output \g17194/_0_  ;
  output \g17195/_0_  ;
  output \g17196/_0_  ;
  output \g17197/_0_  ;
  output \g17198/_0_  ;
  output \g17199/_0_  ;
  output \g17200/_0_  ;
  output \g17201/_0_  ;
  output \g17202/_0_  ;
  output \g17203/_0_  ;
  output \g17204/_0_  ;
  output \g17205/_0_  ;
  output \g17206/_0_  ;
  output \g17207/_0_  ;
  output \g17208/_0_  ;
  output \g17209/_0_  ;
  output \g17210/_0_  ;
  output \g17211/_0_  ;
  output \g17212/_0_  ;
  output \g17213/_0_  ;
  output \g17214/_0_  ;
  output \g17215/_0_  ;
  output \g17216/_0_  ;
  output \g17217/_0_  ;
  output \g17218/_0_  ;
  output \g17219/_0_  ;
  output \g17223/_0_  ;
  output \g17224/_0_  ;
  output \g17225/_0_  ;
  output \g17226/_0_  ;
  output \g17227/_0_  ;
  output \g17228/_0_  ;
  output \g17229/_0_  ;
  output \g17231/_0_  ;
  output \g17232/_0_  ;
  output \g17233/_0_  ;
  output \g17234/_0_  ;
  output \g17237/_0_  ;
  output \g17239/_0_  ;
  output \g17240/_0_  ;
  output \g17243/_0_  ;
  output \g17246/_0_  ;
  output \g17247/_0_  ;
  output \g17248/_0_  ;
  output \g17249/_0_  ;
  output \g17250/_0_  ;
  output \g17251/_0_  ;
  output \g17252/_0_  ;
  output \g17253/_0_  ;
  output \g17254/_0_  ;
  output \g17258/_0_  ;
  output \g17261/_0_  ;
  output \g17262/_0_  ;
  output \g17269/_0_  ;
  output \g17271/_0_  ;
  output \g17274/_0_  ;
  output \g17275/_0_  ;
  output \g17276/_0_  ;
  output \g17277/_0_  ;
  output \g17278/_0_  ;
  output \g17279/_0_  ;
  output \g17280/_0_  ;
  output \g17281/_0_  ;
  output \g17282/_0_  ;
  output \g17283/_0_  ;
  output \g17285/_0_  ;
  output \g17290/_0_  ;
  output \g17292/_0_  ;
  output \g17293/_0_  ;
  output \g17296/_0_  ;
  output \g17297/_0_  ;
  output \g17298/_0_  ;
  output \g173/_0_  ;
  output \g17303/_0_  ;
  output \g17304/_0_  ;
  output \g17305/_0_  ;
  output \g17306/_0_  ;
  output \g17307/_0_  ;
  output \g17308/_0_  ;
  output \g17309/_0_  ;
  output \g17310/_0_  ;
  output \g17311/_0_  ;
  output \g17312/_0_  ;
  output \g17314/_0_  ;
  output \g17315/_0_  ;
  output \g17316/_0_  ;
  output \g17317/_0_  ;
  output \g17318/_0_  ;
  output \g17319/_0_  ;
  output \g17320/_0_  ;
  output \g17321/_0_  ;
  output \g17322/_0_  ;
  output \g17323/_0_  ;
  output \g17324/_0_  ;
  output \g17325/_0_  ;
  output \g17326/_0_  ;
  output \g17327/_0_  ;
  output \g17328/_0_  ;
  output \g17329/_0_  ;
  output \g17330/_0_  ;
  output \g17331/_0_  ;
  output \g17332/_0_  ;
  output \g17333/_0_  ;
  output \g17335/_0_  ;
  output \g17336/_0_  ;
  output \g17337/_0_  ;
  output \g17338/_0_  ;
  output \g17339/_0_  ;
  output \g17340/_0_  ;
  output \g17342/_0_  ;
  output \g17343/_0_  ;
  output \g17347/_0_  ;
  output \g17350/_0_  ;
  output \g17354/_0_  ;
  output \g17356/_0_  ;
  output \g17357/_0_  ;
  output \g17358/_0_  ;
  output \g17359/_0_  ;
  output \g17360/_0_  ;
  output \g17415/_0_  ;
  output \g17441/_0_  ;
  output \g17442/_0_  ;
  output \g17451/_0_  ;
  output \g17457/_0_  ;
  output \g17458/_0_  ;
  output \g17459/_0_  ;
  output \g17460/_0_  ;
  output \g17461/_0_  ;
  output \g17462/_0_  ;
  output \g17463/_0_  ;
  output \g17464/_0_  ;
  output \g17465/_0_  ;
  output \g17466/_0_  ;
  output \g17467/_0_  ;
  output \g17468/_0_  ;
  output \g17469/_0_  ;
  output \g17470/_0_  ;
  output \g17471/_0_  ;
  output \g17472/_0_  ;
  output \g175/_3_  ;
  output \g1750/_0_  ;
  output \g176/_3_  ;
  output \g17619/_0_  ;
  output \g17620/_0_  ;
  output \g1763/_3_  ;
  output \g1764/_3_  ;
  output \g1768/_0_  ;
  output \g1769/_0_  ;
  output \g177/_3_  ;
  output \g17737/_0_  ;
  output \g17747/_0_  ;
  output \g178/_3_  ;
  output \g17814/_1_  ;
  output \g17815/_0_  ;
  output \g17821/_1_  ;
  output \g17821/_1__syn_2  ;
  output \g17872/_0_  ;
  output \g179/_3_  ;
  output \g17902/_0_  ;
  output \g180/_3_  ;
  output \g18020/_1_  ;
  output \g18057/_0_  ;
  output \g18096/_0_  ;
  output \g18099/_0_  ;
  output \g18107/_0_  ;
  output \g18133/_0_  ;
  output \g18140/_1_  ;
  output \g18153/_0_  ;
  output \g182/_0_  ;
  output \g18218/_0_  ;
  output \g18244/_0_  ;
  output \g18262/_0_  ;
  output \g18267/_0_  ;
  output \g18387/_1__syn_2  ;
  output \g184/_0_  ;
  output \g18478/_1_  ;
  output \g18585/_3_  ;
  output \g18608/_0_  ;
  output \g18609/_0_  ;
  output \g18613/_0_  ;
  output \g18618/_0_  ;
  output \g18647/_0_  ;
  output \g18687/_2_  ;
  output \g18707/_0_  ;
  output \g18748/_0_  ;
  output \g18753/_0_  ;
  output \g18758/_0_  ;
  output \g18759/_0_  ;
  output \g18760/_0_  ;
  output \g18761/_0_  ;
  output \g18762/_0_  ;
  output \g18763/_0_  ;
  output \g18764/_0_  ;
  output \g18765/_0_  ;
  output \g18766/_0_  ;
  output \g18767/_0_  ;
  output \g18768/_0_  ;
  output \g18770/_0_  ;
  output \g18771/_0_  ;
  output \g18788/_0_  ;
  output \g18796/_0_  ;
  output \g18800/_0_  ;
  output \g18801/_0_  ;
  output \g18802/_0_  ;
  output \g18803/_0_  ;
  output \g18804/_0_  ;
  output \g18805/_0_  ;
  output \g18807/_0_  ;
  output \g18840/_0_  ;
  output \g18843/_0_  ;
  output \g18844/_0_  ;
  output \g18846/_0_  ;
  output \g18847/_0_  ;
  output \g18848/_0_  ;
  output \g18849/_0_  ;
  output \g18850/_0_  ;
  output \g18851/_0_  ;
  output \g18852/_0_  ;
  output \g18853/_0_  ;
  output \g18854/_0_  ;
  output \g18855/_0_  ;
  output \g18856/_0_  ;
  output \g18858/_0_  ;
  output \g18860/_0_  ;
  output \g18861/_0_  ;
  output \g18863/_0_  ;
  output \g18864/_0_  ;
  output \g18866/_0_  ;
  output \g18867/_0_  ;
  output \g18868/_0_  ;
  output \g18869/_0_  ;
  output \g18870/_0_  ;
  output \g18871/_0_  ;
  output \g18872/_0_  ;
  output \g18873/_0_  ;
  output \g18874/_0_  ;
  output \g18875/_0_  ;
  output \g18876/_0_  ;
  output \g18877/_0_  ;
  output \g18878/_0_  ;
  output \g18879/_0_  ;
  output \g18880/_0_  ;
  output \g18881/_0_  ;
  output \g18882/_0_  ;
  output \g18883/_0_  ;
  output \g18888/_0_  ;
  output \g18892/_0_  ;
  output \g18895/_0_  ;
  output \g18896/_0_  ;
  output \g18897/_0_  ;
  output \g18905/_0_  ;
  output \g18908/_0_  ;
  output \g18909/_0_  ;
  output \g18912/_0_  ;
  output \g18918/_0_  ;
  output \g18919/_0_  ;
  output \g18920/_0_  ;
  output \g18921/_0_  ;
  output \g18922/_0_  ;
  output \g18924/_0_  ;
  output \g18925/_0_  ;
  output \g18927/_0_  ;
  output \g18930/_0_  ;
  output \g18966/_0_  ;
  output \g18968/_0_  ;
  output \g18970/_0_  ;
  output \g18974/_0_  ;
  output \g18975/_0_  ;
  output \g18977/_0_  ;
  output \g18981/_0_  ;
  output \g18983/_0_  ;
  output \g18985/_0_  ;
  output \g18987/_0_  ;
  output \g18989/_0_  ;
  output \g18991/_0_  ;
  output \g18992/_0_  ;
  output \g18993/_0_  ;
  output \g18994/_0_  ;
  output \g18995/_0_  ;
  output \g18996/_0_  ;
  output \g18997/_0_  ;
  output \g18998/_0_  ;
  output \g18999/_0_  ;
  output \g19001/_0_  ;
  output \g19003/_0_  ;
  output \g19005/_0_  ;
  output \g19006/_0_  ;
  output \g19014/_0_  ;
  output \g19016/_0_  ;
  output \g19018/_0_  ;
  output \g19020/_0_  ;
  output \g19022/_0_  ;
  output \g19056/_3_  ;
  output \g19058/_3_  ;
  output \g19060/_3_  ;
  output \g19062/_3_  ;
  output \g1910/_0_  ;
  output \g19186/_0_  ;
  output \g19188/_0_  ;
  output \g19235/_0_  ;
  output \g19239/_0_  ;
  output \g19244/_0_  ;
  output \g19253/_0_  ;
  output \g19254/_0_  ;
  output \g19259/_0_  ;
  output \g19261/_0_  ;
  output \g19267/_0_  ;
  output \g19277/_0_  ;
  output \g19278/_0_  ;
  output \g19280/_0_  ;
  output \g19281/_0_  ;
  output \g19282/_0_  ;
  output \g19283/_0_  ;
  output \g19284/_0_  ;
  output \g19285/_0_  ;
  output \g19286/_0_  ;
  output \g19287/_0_  ;
  output \g19288/_0_  ;
  output \g19289/_0_  ;
  output \g19290/_0_  ;
  output \g19291/_0_  ;
  output \g19292/_0_  ;
  output \g19293/_0_  ;
  output \g19294/_0_  ;
  output \g19295/_0_  ;
  output \g19296/_0_  ;
  output \g19297/_0_  ;
  output \g19298/_0_  ;
  output \g19299/_0_  ;
  output \g19300/_0_  ;
  output \g19301/_0_  ;
  output \g19302/_0_  ;
  output \g19303/_0_  ;
  output \g19304/_0_  ;
  output \g19305/_0_  ;
  output \g19306/_0_  ;
  output \g19307/_0_  ;
  output \g19308/_0_  ;
  output \g19315/_0_  ;
  output \g19316/_0_  ;
  output \g19317/_0_  ;
  output \g19318/_0_  ;
  output \g19319/_0_  ;
  output \g19320/_0_  ;
  output \g19321/_0_  ;
  output \g19322/_0_  ;
  output \g19323/_0_  ;
  output \g19325/_3_  ;
  output \g19326/_3_  ;
  output \g19333/_3_  ;
  output \g19341/_3_  ;
  output \g19347/_3_  ;
  output \g19377/_3_  ;
  output \g19381/_3_  ;
  output \g19393/_0_  ;
  output \g19401/_0_  ;
  output \g19402/_0_  ;
  output \g195/_2_  ;
  output \g19513/_0_  ;
  output \g19514/_0_  ;
  output \g19515/_0_  ;
  output \g19516/_0_  ;
  output \g1952/_3_  ;
  output \g19529/_0_  ;
  output \g19530/_0_  ;
  output \g19531/_0_  ;
  output \g19532/_0_  ;
  output \g19533/_0_  ;
  output \g19534/_0_  ;
  output \g19535/_0_  ;
  output \g19536/_0_  ;
  output \g19537/_0_  ;
  output \g19539/_0_  ;
  output \g19546/_0_  ;
  output \g19552/_0_  ;
  output \g19553/_0_  ;
  output \g19562/_0_  ;
  output \g19563/_0_  ;
  output \g19564/_0_  ;
  output \g19572/_0_  ;
  output \g19575/_0_  ;
  output \g19615/_0_  ;
  output \g19686/_0_  ;
  output \g19688/_0_  ;
  output \g197/_0_  ;
  output \g19729/_0_  ;
  output \g19774/_0_  ;
  output \g19777/_0_  ;
  output \g19791/_0_  ;
  output \g19818/_0_  ;
  output \g19819/_0_  ;
  output \g19828/_0_  ;
  output \g19852/_1_  ;
  output \g19860/_0_  ;
  output \g19861/_0_  ;
  output \g19864/_0_  ;
  output \g19886/_0_  ;
  output \g19887/_0_  ;
  output \g199/_0_  ;
  output \g19908/_0_  ;
  output \g19918/_0_  ;
  output \g19927/_0_  ;
  output \g19933/_0_  ;
  output \g200/_0_  ;
  output \g20019/_0_  ;
  output \g20046/_0_  ;
  output \g20068/_1_  ;
  output \g20080/_1_  ;
  output \g201/_0_  ;
  output \g20137/_0_  ;
  output \g20139/_0_  ;
  output \g20141/_0_  ;
  output \g20152/_1_  ;
  output \g20154/_00_  ;
  output \g202/_0_  ;
  output \g20206/_0_  ;
  output \g20211/_2_  ;
  output \g20217/_2_  ;
  output \g20239/_0_  ;
  output \g20265/_2_  ;
  output \g20266/_0_  ;
  output \g20272/_2_  ;
  output \g20278/_2_  ;
  output \g20283/_0_  ;
  output \g20285/_2_  ;
  output \g20288/_2__syn_2  ;
  output \g20293/_0_  ;
  output \g20295/_2_  ;
  output \g203/_0_  ;
  output \g20302/_2_  ;
  output \g20303/_2_  ;
  output \g20304/_2_  ;
  output \g20311/_2_  ;
  output \g20326/_0_  ;
  output \g20330/_0_  ;
  output \g2034/_0_  ;
  output \g20345/_0_  ;
  output \g20346/_0_  ;
  output \g2035/_0_  ;
  output \g20363/_0_  ;
  output \g20364/_0_  ;
  output \g204/_0_  ;
  output \g2047/_0_  ;
  output \g20483/_0_  ;
  output \g20493/_00_  ;
  output \g205/_0_  ;
  output \g20569/_0_  ;
  output \g20570/_0_  ;
  output \g20571/_0_  ;
  output \g206/_0_  ;
  output \g20613/_0_  ;
  output \g20615/_0_  ;
  output \g20657/_1__syn_2  ;
  output \g20660/_0_  ;
  output \g20685/_0_  ;
  output \g207/_0_  ;
  output \g20713/_1_  ;
  output \g20747/_1_  ;
  output \g20784/_0_  ;
  output \g20820/_1_  ;
  output \g20859/_0_  ;
  output \g20873/_2_  ;
  output \g20886/_0_  ;
  output \g20887/_0_  ;
  output \g20891/_2__syn_2  ;
  output \g20907/_2_  ;
  output \g20936/_2__syn_2  ;
  output \g20937/_1_  ;
  output \g20955/_0_  ;
  output \g20959/_2__syn_2  ;
  output \g20967/_0_  ;
  output \g20971/_2__syn_2  ;
  output \g20974/_1__syn_2  ;
  output \g21015/_1_  ;
  output \g21051/_2_  ;
  output \g21079/_1_  ;
  output \g21081/_1_  ;
  output \g21087/_2__syn_2  ;
  output \g21114/_1_  ;
  output \g21116/_1_  ;
  output \g21120/_2__syn_2  ;
  output \g21147/_0_  ;
  output \g21179/_1_  ;
  output \g21185/_1_  ;
  output \g21223/_0_  ;
  output \g21242/_0_  ;
  output \g21253/_0_  ;
  output \g21257/_0_  ;
  output \g21323/_1_  ;
  output \g21324/_1_  ;
  output \g21366/_0_  ;
  output \g21385/_2_  ;
  output \g21464/_0_  ;
  output \g21475/_3_  ;
  output \g21481/_0_  ;
  output \g21482/_0_  ;
  output \g21494/_3_  ;
  output \g21500/_3_  ;
  output \g21507/_3_  ;
  output \g21511/_3_  ;
  output \g21537/_1_  ;
  output \g21568/_0_  ;
  output \g21591/_0_  ;
  output \g21604/_0_  ;
  output \g21605/_3_  ;
  output \g21606/_0_  ;
  output \g21607/_0_  ;
  output \g21608/_0_  ;
  output \g21609/_0_  ;
  output \g21610/_0_  ;
  output \g21611/_0_  ;
  output \g21612/_0_  ;
  output \g21613/_0_  ;
  output \g21614/_0_  ;
  output \g21615/_0_  ;
  output \g21616/_0_  ;
  output \g21617/_0_  ;
  output \g21618/_0_  ;
  output \g21621/_0_  ;
  output \g21640/_0_  ;
  output \g21678/_0_  ;
  output \g21679/_0_  ;
  output \g21686/_0_  ;
  output \g21692/_3_  ;
  output \g21696/_0_  ;
  output \g21698/_0_  ;
  output \g21702/_3_  ;
  output \g21707/_0_  ;
  output \g21709/_0_  ;
  output \g21728/_0_  ;
  output \g21729/_0_  ;
  output \g21731/_0_  ;
  output \g21732/_0_  ;
  output \g21733/_0_  ;
  output \g21736/_0_  ;
  output \g21744/_3_  ;
  output \g21753/_0_  ;
  output \g21754/_0_  ;
  output \g21755/_0_  ;
  output \g21756/_0_  ;
  output \g21757/_0_  ;
  output \g21759/_0_  ;
  output \g21761/_0_  ;
  output \g21763/_0_  ;
  output \g21764/_0_  ;
  output \g21766/_0_  ;
  output \g2180/_0_  ;
  output \g21853/_3_  ;
  output \g21861/_3_  ;
  output \g21863/_3_  ;
  output \g21869/_3_  ;
  output \g2187/_0_  ;
  output \g21875/_3_  ;
  output \g21877/_3_  ;
  output \g21879/_3_  ;
  output \g2188/_0_  ;
  output \g21900/_0_  ;
  output \g22080/_0_  ;
  output \g22082/_0_  ;
  output \g22135/_0_  ;
  output \g22145/_1_  ;
  output \g22225/_0_  ;
  output \g223/_0_  ;
  output \g22354/_0_  ;
  output \g224/_0_  ;
  output \g22412/_0_  ;
  output \g22415/_1__syn_2  ;
  output \g225/_0_  ;
  output \g2257/_0_  ;
  output \g226/_3_  ;
  output \g22624/_0_  ;
  output \g227/_3_  ;
  output \g22702/_0_  ;
  output \g22919/_1__syn_2  ;
  output \g22933/_0_  ;
  output \g22954/_0_  ;
  output \g22989/_1_  ;
  output \g23529/_0_  ;
  output \g23539/_0_  ;
  output \g2362/_2_  ;
  output \g23766/_0_  ;
  output \g24/_3_  ;
  output \g24018/_0_  ;
  output \g2416/_0_  ;
  output \g2420/_0_  ;
  output \g24213/_0_  ;
  output \g24301/_0_  ;
  output \g2479/_0_  ;
  output \g248/_3_  ;
  output \g2480/_0_  ;
  output \g2481/_0_  ;
  output \g2482/_0_  ;
  output \g2483/_0_  ;
  output \g2484/_0_  ;
  output \g2485/_0_  ;
  output \g2486/_0_  ;
  output \g2487/_0_  ;
  output \g2488/_0_  ;
  output \g249/_3_  ;
  output \g2490/_0_  ;
  output \g2491/_0_  ;
  output \g2492/_0_  ;
  output \g2493/_0_  ;
  output \g2494/_0_  ;
  output \g2495/_0_  ;
  output \g2496/_0_  ;
  output \g2497/_0_  ;
  output \g2507/_0_  ;
  output \g2508/_0_  ;
  output \g2509/_0_  ;
  output \g2510/_0_  ;
  output \g2511/_0_  ;
  output \g2512/_0_  ;
  output \g2513/_0_  ;
  output \g2514/_0_  ;
  output \g2515/_0_  ;
  output \g2516/_0_  ;
  output \g25237/_0_  ;
  output \g2558/_0_  ;
  output \g2562/_0_  ;
  output \g2563/_0_  ;
  output \g2564/_0_  ;
  output \g2565/_0_  ;
  output \g2566/_0_  ;
  output \g2567/_0_  ;
  output \g2699/_0_  ;
  output \g27/_2_  ;
  output \g271/_0_  ;
  output \g272/_3_  ;
  output \g273/_3_  ;
  output \g274/_3_  ;
  output \g275/_3_  ;
  output \g276/_3_  ;
  output \g277/_3_  ;
  output \g2787/_3_  ;
  output \g2788/_3_  ;
  output \g279/_0_  ;
  output \g2795/_0_  ;
  output \g2796/_0_  ;
  output \g280/_0_  ;
  output \g2842/_3_  ;
  output \g29/_1_  ;
  output \g2927/_0_  ;
  output \g2978/_0_  ;
  output \g2979/_0_  ;
  output \g2980/_0_  ;
  output \g2981/_0_  ;
  output \g2982/_0_  ;
  output \g2983/_0_  ;
  output \g2984/_0_  ;
  output \g2985/_0_  ;
  output \g3021/_3_  ;
  output \g3022/_3_  ;
  output \g3023/_3_  ;
  output \g3024/_3_  ;
  output \g3025/_3_  ;
  output \g3026/_3_  ;
  output \g3027/_3_  ;
  output \g3028/_3_  ;
  output \g3029/_3_  ;
  output \g3030/_3_  ;
  output \g3031/_3_  ;
  output \g3032/_3_  ;
  output \g3033/_3_  ;
  output \g3034/_3_  ;
  output \g3035/_3_  ;
  output \g3036/_3_  ;
  output \g3037/_3_  ;
  output \g3038/_3_  ;
  output \g3039/_3_  ;
  output \g3040/_3_  ;
  output \g3041/_3_  ;
  output \g3042/_3_  ;
  output \g3049/_0_  ;
  output \g3050/_0_  ;
  output \g3051/_0_  ;
  output \g3052/_0_  ;
  output \g3053/_0_  ;
  output \g3054/_0_  ;
  output \g3058/_0_  ;
  output \g3059/_0_  ;
  output \g3088/_0_  ;
  output \g3089/_0_  ;
  output \g3090/_0_  ;
  output \g3091/_0_  ;
  output \g3092/_0_  ;
  output \g3093/_0_  ;
  output \g3094/_0_  ;
  output \g3095/_0_  ;
  output \g314/_0_  ;
  output \g3147/_3_  ;
  output \g3148/_3_  ;
  output \g3189/_0_  ;
  output \g3190/_0_  ;
  output \g3191/_0_  ;
  output \g3192/_0_  ;
  output \g3193/_0_  ;
  output \g3194/_0_  ;
  output \g3195/_0_  ;
  output \g3196/_0_  ;
  output \g3197/_0_  ;
  output \g3198/_0_  ;
  output \g3199/_0_  ;
  output \g32/_0_  ;
  output \g320/_3_  ;
  output \g3200/_0_  ;
  output \g3201/_0_  ;
  output \g3202/_0_  ;
  output \g3203/_0_  ;
  output \g3204/_0_  ;
  output \g321/_3_  ;
  output \g325/_3_  ;
  output \g3271/_2_  ;
  output \g33/_0_  ;
  output \g3363/_0_  ;
  output \g3413/_0_  ;
  output \g3414/_0_  ;
  output \g352/_0_  ;
  output \g355/_0_  ;
  output \g356/_3_  ;
  output \g357/_3_  ;
  output \g35_dup/_1_  ;
  output \g36/_3_  ;
  output \g365/_3_  ;
  output \g366/_3_  ;
  output \g367/_3_  ;
  output \g368/_3_  ;
  output \g3687/_0_  ;
  output \g369/_3_  ;
  output \g37/_3_  ;
  output \g370/_3_  ;
  output \g372/_3_  ;
  output \g374/_3_  ;
  output \g3740/_0_  ;
  output \g375/_3_  ;
  output \g376/_3_  ;
  output \g3878/_0_  ;
  output \g3879/_0_  ;
  output \g388/_3_  ;
  output \g3880/_0_  ;
  output \g3881/_0_  ;
  output \g3882/_0_  ;
  output \g389/_3_  ;
  output \g3894/_0_  ;
  output \g3895/_0_  ;
  output \g3896/_0_  ;
  output \g3897/_0_  ;
  output \g3898/_0_  ;
  output \g392/_3_  ;
  output \g393/_3_  ;
  output \g394/_3_  ;
  output \g395/_3_  ;
  output \g396/_3_  ;
  output \g397/_3_  ;
  output \g398/_3_  ;
  output \g399/_3_  ;
  output \g401/_3_  ;
  output \g402/_3_  ;
  output \g404/_3_  ;
  output \g4048/_0_  ;
  output \g405/_3_  ;
  output \g4050/_0_  ;
  output \g406/_3_  ;
  output \g407/_3_  ;
  output \g410/_3_  ;
  output \g411/_3_  ;
  output \g412/_3_  ;
  output \g413/_3_  ;
  output \g415/_3_  ;
  output \g416/_3_  ;
  output \g42/_0_  ;
  output \g4216/_3_  ;
  output \g4217/_3_  ;
  output \g4218/_3_  ;
  output \g4219/_3_  ;
  output \g4296/_0_  ;
  output \g4297/_0_  ;
  output \g4298/_0_  ;
  output \g4299/_0_  ;
  output \g43/_0_  ;
  output \g4300/_0_  ;
  output \g4301/_0_  ;
  output \g4302/_0_  ;
  output \g4303/_0_  ;
  output \g4304/_0_  ;
  output \g4305/_0_  ;
  output \g4306/_0_  ;
  output \g4307/_0_  ;
  output \g4308/_0_  ;
  output \g4309/_0_  ;
  output \g4310/_0_  ;
  output \g4311/_0_  ;
  output \g4312/_0_  ;
  output \g4313/_0_  ;
  output \g4314/_0_  ;
  output \g4315/_0_  ;
  output \g4316/_0_  ;
  output \g4317/_0_  ;
  output \g4318/_0_  ;
  output \g4319/_0_  ;
  output \g4320/_0_  ;
  output \g4321/_0_  ;
  output \g4322/_0_  ;
  output \g4323/_0_  ;
  output \g436/_0_  ;
  output \g44/_0_  ;
  output \g448/_3_  ;
  output \g45/_0_  ;
  output \g4587/_0_  ;
  output \g4588/_0_  ;
  output \g46/_0_  ;
  output \g4601/_0_  ;
  output \g4602/_0_  ;
  output \g4613/_3_  ;
  output \g4614/_3_  ;
  output \g4615/_3_  ;
  output \g463/_0_  ;
  output \g465/_0_  ;
  output \g4653/_0_  ;
  output \g4654/_0_  ;
  output \g4655/_0_  ;
  output \g4656/_0_  ;
  output \g4659/_0_  ;
  output \g466/_0_  ;
  output \g468/_3_  ;
  output \g469/_3_  ;
  output \g4697/_0_  ;
  output \g47/_3_  ;
  output \g470/_0_  ;
  output \g471/_0_  ;
  output \g4755/_0_  ;
  output \g476/_0_  ;
  output \g48/_3_  ;
  output \g480/_00_  ;
  output \g4839/_0_  ;
  output \g4840/_0_  ;
  output \g485/_3_  ;
  output \g4854/_0_  ;
  output \g4855/_0_  ;
  output \g4859/_0_  ;
  output \g486/_3_  ;
  output \g4860/_0_  ;
  output \g4880/_0_  ;
  output \g4881/_0_  ;
  output \g4882/_0_  ;
  output \g4883/_0_  ;
  output \g4884/_0_  ;
  output \g4885/_0_  ;
  output \g4886/_0_  ;
  output \g4887/_0_  ;
  output \g4888/_0_  ;
  output \g49/_0_  ;
  output \g494/_0_  ;
  output \g499/_1_  ;
  output \g50/_0_  ;
  output \g5002/_0_  ;
  output \g5003/_0_  ;
  output \g5009/_0_  ;
  output \g5010/_0_  ;
  output \g5011/_0_  ;
  output \g5014/_0_  ;
  output \g51/_0_  ;
  output \g5105/_0_  ;
  output \g5129/_2_  ;
  output \g5132/_0_  ;
  output \g5135/_0_  ;
  output \g5168/_0_  ;
  output \g5169/_0_  ;
  output \g5173/_0_  ;
  output \g5224/_0_  ;
  output \g5225/_0_  ;
  output \g5226/_0_  ;
  output \g5227/_0_  ;
  output \g5334/_0_  ;
  output \g5335/_0_  ;
  output \g5336/_0_  ;
  output \g5337/_0_  ;
  output \g5338/_0_  ;
  output \g5339/_0_  ;
  output \g5340/_0_  ;
  output \g5341/_0_  ;
  output \g5342/_0_  ;
  output \g5343/_0_  ;
  output \g5344/_0_  ;
  output \g5345/_0_  ;
  output \g5346/_0_  ;
  output \g5347/_0_  ;
  output \g5348/_0_  ;
  output \g5349/_0_  ;
  output \g5395/_0_  ;
  output \g54/_0_  ;
  output \g5434/_0_  ;
  output \g5447/_0_  ;
  output \g5450/_0_  ;
  output \g5451/_0_  ;
  output \g5452/_0_  ;
  output \g5453/_0_  ;
  output \g5454/_0_  ;
  output \g5461/_0_  ;
  output \g5483/_0_  ;
  output \g5484/_0_  ;
  output \g5492/_0_  ;
  output \g5493/_0_  ;
  output \g5496/_3_  ;
  output \g5497/_3_  ;
  output \g55/_0_  ;
  output \g5500/_0_  ;
  output \g5502/_0_  ;
  output \g5503/_0_  ;
  output \g5506/_0_  ;
  output \g5511/_0_  ;
  output \g5518/_0_  ;
  output \g5519/_0_  ;
  output \g5520/_0_  ;
  output \g5522/_0_  ;
  output \g5523/_0_  ;
  output \g5524/_0_  ;
  output \g5525/_0_  ;
  output \g5532/_0_  ;
  output \g5533/_0_  ;
  output \g5534/_0_  ;
  output \g5535/_0_  ;
  output \g5536/_0_  ;
  output \g5537/_0_  ;
  output \g5538/_0_  ;
  output \g5546/_0_  ;
  output \g5555/_00_  ;
  output \g5593/_0_  ;
  output \g5614/_2_  ;
  output \g567/_0_  ;
  output \g5677/_0_  ;
  output \g5678/_0_  ;
  output \g5682/_0_  ;
  output \g5683/_0_  ;
  output \g5684/_0_  ;
  output \g5686/_0_  ;
  output \g5687/_0_  ;
  output \g5689/_0_  ;
  output \g5690/_0_  ;
  output \g5691/_0_  ;
  output \g5692/_0_  ;
  output \g5698/_0_  ;
  output \g5699/_0_  ;
  output \g5700/_0_  ;
  output \g5701/_0_  ;
  output \g5702/_0_  ;
  output \g5703/_0_  ;
  output \g5704/_0_  ;
  output \g5709/_0_  ;
  output \g5711/_0_  ;
  output \g5714/_0_  ;
  output \g572/_0_  ;
  output \g5723/_0_  ;
  output \g5724/_0_  ;
  output \g5725/_0_  ;
  output \g573/_0_  ;
  output \g5739/_0_  ;
  output \g5740/_0_  ;
  output \g575/_0_  ;
  output \g5756/_0_  ;
  output \g5757/_0_  ;
  output \g5758/_0_  ;
  output \g5759/_0_  ;
  output \g576/_0_  ;
  output \g5760/_0_  ;
  output \g5761/_0_  ;
  output \g5762/_0_  ;
  output \g5763/_0_  ;
  output \g577/_0_  ;
  output \g5772/_0_  ;
  output \g5773/_0_  ;
  output \g5774/_0_  ;
  output \g5775/_0_  ;
  output \g5776/_0_  ;
  output \g5777/_0_  ;
  output \g578/_0_  ;
  output \g5781/_0_  ;
  output \g5783/_0_  ;
  output \g5784/_0_  ;
  output \g5785/_0_  ;
  output \g5786/_0_  ;
  output \g5787/_0_  ;
  output \g5788/_0_  ;
  output \g5789/_0_  ;
  output \g579/_0_  ;
  output \g5790/_0_  ;
  output \g5791/_0_  ;
  output \g5792/_0_  ;
  output \g5794/_0_  ;
  output \g5795/_0_  ;
  output \g5796/_0_  ;
  output \g580/_0_  ;
  output \g5801/_0_  ;
  output \g5802/_0_  ;
  output \g5803/_0_  ;
  output \g5804/_0_  ;
  output \g5805/_0_  ;
  output \g581/_0_  ;
  output \g5814/_0_  ;
  output \g582/_0_  ;
  output \g583/_0_  ;
  output \g5849/_3_  ;
  output \g585/_0_  ;
  output \g586/_0_  ;
  output \g587/_0_  ;
  output \g588/_0_  ;
  output \g589/_0_  ;
  output \g590/_0_  ;
  output \g591/_0_  ;
  output \g592/_0_  ;
  output \g593/_0_  ;
  output \g594/_0_  ;
  output \g595/_0_  ;
  output \g596/_0_  ;
  output \g597/_0_  ;
  output \g5971/_0_  ;
  output \g5972/_0_  ;
  output \g5976/_0_  ;
  output \g598/_0_  ;
  output \g5989/_0_  ;
  output \g599/_0_  ;
  output \g600/_0_  ;
  output \g601/_0_  ;
  output \g602/_0_  ;
  output \g603/_0_  ;
  output \g604/_0_  ;
  output \g605/_0_  ;
  output \g6092/_0_  ;
  output \g6093/_2_  ;
  output \g6094/_0_  ;
  output \g6114/_0_  ;
  output \g614/_3_  ;
  output \g6148/_0_  ;
  output \g6149/_0_  ;
  output \g6171/_0_  ;
  output \g6172/_0_  ;
  output \g6173/_0_  ;
  output \g6174/_0_  ;
  output \g6175/_0_  ;
  output \g6176/_0_  ;
  output \g6177/_0_  ;
  output \g6178/_0_  ;
  output \g6179/_0_  ;
  output \g6180/_0_  ;
  output \g6181/_0_  ;
  output \g6182/_0_  ;
  output \g6183/_0_  ;
  output \g6184/_0_  ;
  output \g6185/_0_  ;
  output \g6186/_0_  ;
  output \g6187/_0_  ;
  output \g6193/_0_  ;
  output \g6196/_0_  ;
  output \g6197/_0_  ;
  output \g6198/_3_  ;
  output \g6200/_2_  ;
  output \g6202/_2_  ;
  output \g6203/_3_  ;
  output \g6204/_3_  ;
  output \g6209/_0_  ;
  output \g6211/_0_  ;
  output \g6215/_0_  ;
  output \g6217/_0_  ;
  output \g6219/_0_  ;
  output \g6220/_0_  ;
  output \g6222/_0_  ;
  output \g6224/_0_  ;
  output \g6228/_0_  ;
  output \g6238/_0_  ;
  output \g6239/_0_  ;
  output \g6240/_0_  ;
  output \g6242/_0_  ;
  output \g6243/_0_  ;
  output \g6244/_0_  ;
  output \g6245/_0_  ;
  output \g6246/_0_  ;
  output \g6248/_0_  ;
  output \g6249/_0_  ;
  output \g6259/_0_  ;
  output \g6260/_0_  ;
  output \g6261/_0_  ;
  output \g6262/_0_  ;
  output \g6263/_0_  ;
  output \g6264/_0_  ;
  output \g6265/_0_  ;
  output \g6266/_0_  ;
  output \g6267/_0_  ;
  output \g6268/_0_  ;
  output \g6269/_0_  ;
  output \g6270/_0_  ;
  output \g6271/_0_  ;
  output \g6272/_0_  ;
  output \g6277/_0_  ;
  output \g6318/_0_  ;
  output \g6326/_0_  ;
  output \g6329/_0_  ;
  output \g6330/_0_  ;
  output \g6331/_0_  ;
  output \g6332/_0_  ;
  output \g6333/_0_  ;
  output \g6334/_0_  ;
  output \g6335/_0_  ;
  output \g6336/_0_  ;
  output \g6337/_0_  ;
  output \g6338/_0_  ;
  output \g6339/_0_  ;
  output \g6340/_0_  ;
  output \g6341/_0_  ;
  output \g6342/_0_  ;
  output \g6343/_0_  ;
  output \g6344/_0_  ;
  output \g6345/_0_  ;
  output \g6346/_0_  ;
  output \g6347/_0_  ;
  output \g6348/_0_  ;
  output \g6349/_0_  ;
  output \g6350/_0_  ;
  output \g6351/_0_  ;
  output \g6352/_0_  ;
  output \g6353/_0_  ;
  output \g6354/_0_  ;
  output \g6355/_0_  ;
  output \g6361/_0_  ;
  output \g637/_0_  ;
  output \g638/_0_  ;
  output \g639/_3_  ;
  output \g64/_3_  ;
  output \g640/_3_  ;
  output \g6419/_0_  ;
  output \g6442/_0_  ;
  output \g6442/_1_  ;
  output \g6489/_0_  ;
  output \g6490/_0_  ;
  output \g65/_3_  ;
  output \g6513/_0_  ;
  output \g6515/_0_  ;
  output \g6571/_0_  ;
  output \g6588/_0_  ;
  output \g6589/_0_  ;
  output \g6638/_0_  ;
  output \g6639/_0_  ;
  output \g6653/_0_  ;
  output \g6654/_3_  ;
  output \g6655/_0_  ;
  output \g6656/_0_  ;
  output \g6657/_0_  ;
  output \g6687/_0_  ;
  output \g6688/_0_  ;
  output \g6689/_0_  ;
  output \g6690/_0_  ;
  output \g6691/_0_  ;
  output \g6692/_0_  ;
  output \g6693/_0_  ;
  output \g6694/_0_  ;
  output \g6701/_0_  ;
  output \g6706/_0_  ;
  output \g6711/_0_  ;
  output \g6727/_0_  ;
  output \g6728/_0_  ;
  output \g6736/_0_  ;
  output \g6739/_0_  ;
  output \g6742/_0_  ;
  output \g6746/_0_  ;
  output \g6752/_0_  ;
  output \g6771/_0_  ;
  output \g684/_0_  ;
  output \g685/_0_  ;
  output \g686/_0_  ;
  output \g687/_0_  ;
  output \g688/_0_  ;
  output \g689/_0_  ;
  output \g690/_0_  ;
  output \g691/_0_  ;
  output \g692/_0_  ;
  output \g693/_0_  ;
  output \g696/_3_  ;
  output \g697/_3_  ;
  output \g699/_0_  ;
  output \g7/_0_  ;
  output \g700/_0_  ;
  output \g7005/_0_  ;
  output \g7056/_0_  ;
  output \g7057/_0_  ;
  output \g7058/_0_  ;
  output \g7060/_0_  ;
  output \g7075/_0_  ;
  output \g7086/_0_  ;
  output \g7087/_0_  ;
  output \g7089/_0_  ;
  output \g7108/_0_  ;
  output \g7109/_0_  ;
  output \g7112/_0_  ;
  output \g7172/_2_  ;
  output \g7210/_2_  ;
  output \g7211/_0_  ;
  output \g7212/_0_  ;
  output \g7213/_0_  ;
  output \g7214/_0_  ;
  output \g7215/_0_  ;
  output \g7216/_0_  ;
  output \g7217/_3_  ;
  output \g7218/_0_  ;
  output \g7219/_0_  ;
  output \g7220/_0_  ;
  output \g7222/_0_  ;
  output \g7227/_2_  ;
  output \g723/_3_  ;
  output \g7234/_0_  ;
  output \g7237/_3_  ;
  output \g7238/_3_  ;
  output \g7239/_3_  ;
  output \g724/_3_  ;
  output \g7240/_3_  ;
  output \g7241/_3_  ;
  output \g7242/_3_  ;
  output \g7243/_3_  ;
  output \g7244/_0_  ;
  output \g7245/_0_  ;
  output \g7246/_0_  ;
  output \g7247/_0_  ;
  output \g7248/_0_  ;
  output \g7249/_0_  ;
  output \g7250/_0_  ;
  output \g7251/_0_  ;
  output \g7253/_0_  ;
  output \g7254/_0_  ;
  output \g7255/_0_  ;
  output \g7256/_0_  ;
  output \g7257/_0_  ;
  output \g7258/_0_  ;
  output \g7261/_0_  ;
  output \g7264/_0_  ;
  output \g7265/_0_  ;
  output \g7266/_0_  ;
  output \g7267/_0_  ;
  output \g7268/_0_  ;
  output \g7269/_0_  ;
  output \g7278/_0_  ;
  output \g7279/_0_  ;
  output \g7280/_0_  ;
  output \g7281/_0_  ;
  output \g7282/_0_  ;
  output \g7283/_0_  ;
  output \g7284/_0_  ;
  output \g7285/_0_  ;
  output \g7286/_3_  ;
  output \g7288/_3_  ;
  output \g7291/_0_  ;
  output \g7296/_3_  ;
  output \g73/_0_  ;
  output \g7302/_3_  ;
  output \g7306/_3_  ;
  output \g7310/_3_  ;
  output \g7311/_3_  ;
  output \g7312/_3_  ;
  output \g7313/_3_  ;
  output \g7314/_3_  ;
  output \g7315/_3_  ;
  output \g7316/_3_  ;
  output \g7317/_3_  ;
  output \g7323/_3_  ;
  output \g7324/_3_  ;
  output \g7325/_3_  ;
  output \g7327/_0_  ;
  output \g7362/_0_  ;
  output \g74/_0_  ;
  output \g75/_0_  ;
  output \g7512/_0_  ;
  output \g7513/_0_  ;
  output \g7514/_0_  ;
  output \g7515/_0_  ;
  output \g7516/_0_  ;
  output \g7518/_0_  ;
  output \g7528/_0_  ;
  output \g7529/_0_  ;
  output \g7548/_0_  ;
  output \g7549/_0_  ;
  output \g7550/_0_  ;
  output \g7575/_0_  ;
  output \g7576/_0_  ;
  output \g7577/_0_  ;
  output \g7578/_0_  ;
  output \g7579/_0_  ;
  output \g7580/_0_  ;
  output \g7581/_0_  ;
  output \g7582/_0_  ;
  output \g7583/_0_  ;
  output \g7584/_0_  ;
  output \g7585/_0_  ;
  output \g7586/_0_  ;
  output \g7587/_0_  ;
  output \g7588/_0_  ;
  output \g7589/_0_  ;
  output \g7590/_0_  ;
  output \g7591/_0_  ;
  output \g7592/_0_  ;
  output \g7593/_0_  ;
  output \g7594/_0_  ;
  output \g7595/_0_  ;
  output \g7596/_0_  ;
  output \g7597/_0_  ;
  output \g7598/_0_  ;
  output \g7599/_0_  ;
  output \g76/_0_  ;
  output \g7600/_0_  ;
  output \g7601/_0_  ;
  output \g7602/_0_  ;
  output \g7603/_0_  ;
  output \g7604/_0_  ;
  output \g7614/_0_  ;
  output \g7618/_0_  ;
  output \g762/_0_  ;
  output \g7634/_0_  ;
  output \g766/_0_  ;
  output \g767/_0_  ;
  output \g768/_0_  ;
  output \g769/_0_  ;
  output \g77/_0_  ;
  output \g770/_3_  ;
  output \g771/_3_  ;
  output \g7715/_0_  ;
  output \g774/_0_  ;
  output \g7746/_0_  ;
  output \g7753/_0_  ;
  output \g7754/_0_  ;
  output \g7755/_0_  ;
  output \g7756/_0_  ;
  output \g7757/_0_  ;
  output \g7758/_0_  ;
  output \g7759/_0_  ;
  output \g7760/_0_  ;
  output \g7761/_0_  ;
  output \g7762/_0_  ;
  output \g7763/_0_  ;
  output \g7764/_0_  ;
  output \g7765/_0_  ;
  output \g7766/_0_  ;
  output \g7778/_0_  ;
  output \g7779/_0_  ;
  output \g7780/_0_  ;
  output \g7781/_0_  ;
  output \g7782/_0_  ;
  output \g7784/_0_  ;
  output \g78/_0_  ;
  output \g7800/_0_  ;
  output \g7823/_3_  ;
  output \g7837/_0_  ;
  output \g7841/_0_  ;
  output \g7842/_0_  ;
  output \g7843/_0_  ;
  output \g7844/_0_  ;
  output \g7845/_0_  ;
  output \g7846/_0_  ;
  output \g7847/_0_  ;
  output \g7849/_0_  ;
  output \g7850/_0_  ;
  output \g7852/_0_  ;
  output \g7854/_0_  ;
  output \g7855/_0_  ;
  output \g7857/_0_  ;
  output \g7858/_0_  ;
  output \g7859/_0_  ;
  output \g7860/_0_  ;
  output \g7861/_0_  ;
  output \g7862/_0_  ;
  output \g7863/_0_  ;
  output \g7864/_0_  ;
  output \g7865/_0_  ;
  output \g7866/_0_  ;
  output \g7867/_0_  ;
  output \g7868/_0_  ;
  output \g7869/_0_  ;
  output \g7870/_0_  ;
  output \g7871/_0_  ;
  output \g79211/_3_  ;
  output \g79258/_3_  ;
  output \g79299/_3_  ;
  output \g79316/_2_  ;
  output \g79342/_3_  ;
  output \g79401/_3_  ;
  output \g79452/_3_  ;
  output \g79457/_3_  ;
  output \g7951/_0_  ;
  output \g79541/_3_  ;
  output \g7958/_0_  ;
  output \g79598/_3_  ;
  output \g79654/_3_  ;
  output \g79675/_3_  ;
  output \g7971/_0_  ;
  output \g7972/_0_  ;
  output \g7973/_3_  ;
  output \g79753/_3_  ;
  output \g7976/_3_  ;
  output \g79855/_3_  ;
  output \g79858/_3_  ;
  output \g79997/_3_  ;
  output \g8/_0_  ;
  output \g80008/_3_  ;
  output \g80011/_0_  ;
  output \g80104/_0_  ;
  output \g80172/_1_  ;
  output \g80195/_3_  ;
  output \g80238/_3_  ;
  output \g80290/_2_  ;
  output \g80294/_0_  ;
  output \g80302/_0_  ;
  output \g80327/_0_  ;
  output \g80360/_3_  ;
  output \g80373/_0_  ;
  output \g80401/_0_  ;
  output \g80410/_0_  ;
  output \g80475/_0_  ;
  output \g80476/_0_  ;
  output \g80516/_3_  ;
  output \g80536/_0_  ;
  output \g80537/_0_  ;
  output \g80572/_0_  ;
  output \g80573/_0_  ;
  output \g80609/_2_  ;
  output \g80610/_2_  ;
  output \g80676/_0_  ;
  output \g80798/_0_  ;
  output \g80807/_0_  ;
  output \g80890/_2_  ;
  output \g80904/_0_  ;
  output \g81719/_2_  ;
  output \g81746/_0_  ;
  output \g81775/_0_  ;
  output \g81872/_0_  ;
  output \g81961/_0_  ;
  output \g81968/_0_  ;
  output \g82096/_0_  ;
  output \g82123/_0_  ;
  output \g82147/_0_  ;
  output \g82147/_1_  ;
  output \g82335/_0_  ;
  output \g82338/_2_  ;
  output \g82368/_0_  ;
  output \g82460/_2_  ;
  output \g82469/_0_  ;
  output \g82481/_0_  ;
  output \g82625/_1_  ;
  output \g82711/_0_  ;
  output \g82772/_0_  ;
  output \g82946/_0_  ;
  output \g82947/_0_  ;
  output \g82956/_0_  ;
  output \g83003/_0_  ;
  output \g83006/_1_  ;
  output \g83415/_0_  ;
  output \g83498/_0_  ;
  output \g837/_0_  ;
  output \g838/_0_  ;
  output \g83863/_0_  ;
  output \g839/_0_  ;
  output \g84049/_3_  ;
  output \g84050/_3_  ;
  output \g84077/_2_  ;
  output \g842/_0_  ;
  output \g84245/_0_  ;
  output \g843/_0_  ;
  output \g844/_0_  ;
  output \g84448/_0_  ;
  output \g84478/_3_  ;
  output \g845/_0_  ;
  output \g846/_0_  ;
  output \g847/_0_  ;
  output \g848/_0_  ;
  output \g8487/_0_  ;
  output \g8488/_0_  ;
  output \g8489/_0_  ;
  output \g849/_0_  ;
  output \g8490/_0_  ;
  output \g84904/_0_  ;
  output \g8491/_0_  ;
  output \g8492/_0_  ;
  output \g8493/_0_  ;
  output \g8494/_0_  ;
  output \g8496/_0_  ;
  output \g8517/_0_  ;
  output \g8534/_0_  ;
  output \g8538/_0_  ;
  output \g8540/_0_  ;
  output \g8576/_2_  ;
  output \g8597/_0_  ;
  output \g8598/_0_  ;
  output \g8599/_0_  ;
  output \g8600/_0_  ;
  output \g8601/_0_  ;
  output \g8602/_0_  ;
  output \g8603/_0_  ;
  output \g8605/_0_  ;
  output \g8606/_0_  ;
  output \g8607/_0_  ;
  output \g8608/_0_  ;
  output \g8609/_0_  ;
  output \g8610/_0_  ;
  output \g8611/_0_  ;
  output \g8612/_0_  ;
  output \g8613/_0_  ;
  output \g8614/_0_  ;
  output \g8615/_0_  ;
  output \g8617/_0_  ;
  output \g8643/_0_  ;
  output \g8644/_0_  ;
  output \g8645/_0_  ;
  output \g8646/_0_  ;
  output \g8647/_0_  ;
  output \g8648/_0_  ;
  output \g8650/_0_  ;
  output \g8651/_0_  ;
  output \g8652/_0_  ;
  output \g8653/_0_  ;
  output \g8654/_0_  ;
  output \g8655/_0_  ;
  output \g8656/_0_  ;
  output \g8657/_0_  ;
  output \g8658/_0_  ;
  output \g8659/_0_  ;
  output \g8660/_0_  ;
  output \g8665/_00_  ;
  output \g8666/_00_  ;
  output \g8667/_00_  ;
  output \g8668/_00_  ;
  output \g8669/_00_  ;
  output \g86715/_0_  ;
  output \g86745/_3_  ;
  output \g8691/_0_  ;
  output \g8700/_0_  ;
  output \g8701/_0_  ;
  output \g8702/_0_  ;
  output \g8703/_0_  ;
  output \g8704/_0_  ;
  output \g8705/_0_  ;
  output \g87063/_0_  ;
  output \g87114/_0_  ;
  output \g8712/_0_  ;
  output \g8713/_0_  ;
  output \g8714/_0_  ;
  output \g87171/_1_  ;
  output \g87252/_1_  ;
  output \g87298/_0_  ;
  output \g8730/_0_  ;
  output \g8741/_0_  ;
  output \g8747/_0_  ;
  output \g87480/_0_  ;
  output \g87484/_2_  ;
  output \g87488/_1__syn_2  ;
  output \g8761/_0_  ;
  output \g8762/_0_  ;
  output \g8763/_0_  ;
  output \g8764/_0_  ;
  output \g8765/_0_  ;
  output \g8775/_0_  ;
  output \g8776/_0_  ;
  output \g8777/_0_  ;
  output \g8778/_0_  ;
  output \g8784/_0_  ;
  output \g8804/_0_  ;
  output \g8807/_0_  ;
  output \g8808/_0_  ;
  output \g8809/_0_  ;
  output \g8810/_0_  ;
  output \g8811/_0_  ;
  output \g8812/_0_  ;
  output \g8813/_0_  ;
  output \g8814/_0_  ;
  output \g8815/_0_  ;
  output \g8816/_0_  ;
  output \g8817/_0_  ;
  output \g8818/_0_  ;
  output \g8819/_0_  ;
  output \g8820/_0_  ;
  output \g8821/_0_  ;
  output \g8822/_0_  ;
  output \g8823/_0_  ;
  output \g8824/_0_  ;
  output \g8825/_0_  ;
  output \g8826/_0_  ;
  output \g8827/_0_  ;
  output \g8828/_0_  ;
  output \g8829/_0_  ;
  output \g8830/_0_  ;
  output \g8831/_0_  ;
  output \g8832/_0_  ;
  output \g8833/_0_  ;
  output \g8834/_0_  ;
  output \g8835/_0_  ;
  output \g8836/_0_  ;
  output \g8837/_0_  ;
  output \g8838/_0_  ;
  output \g8839/_0_  ;
  output \g8840/_0_  ;
  output \g8842/_0_  ;
  output \g8843/_0_  ;
  output \g8846/_0_  ;
  output \g8848/_0_  ;
  output \g8857/_0_  ;
  output \g8895/_0_  ;
  output \g8902/_3_  ;
  output \g8903/_3_  ;
  output \g8904/_3_  ;
  output \g8905/_3_  ;
  output \g8906/_3_  ;
  output \g8909/_0_  ;
  output \g8910/_0_  ;
  output \g8911/_0_  ;
  output \g8924/_3_  ;
  output \g8926/_3_  ;
  output \g8927/_3_  ;
  output \g8943/_0_  ;
  output \g8944/_0_  ;
  output \g8958/_3_  ;
  output \g8960/_00_  ;
  output \g8961/_3_  ;
  output \g8965/_0_  ;
  output \g8966/_0_  ;
  output \g8967/_0_  ;
  output \g8968/_0_  ;
  output \g9/_0_  ;
  output \g9123/_0_  ;
  output \g9125/_0_  ;
  output \g9126/_0_  ;
  output \g913/_0_  ;
  output \g915/_0_  ;
  output \g916/_0_  ;
  output \g917/_0_  ;
  output \g918/_0_  ;
  output \g919/_0_  ;
  output \g920/_3_  ;
  output \g921/_3_  ;
  output \g925/_0_  ;
  output \g926/_0_  ;
  output \g927/_0_  ;
  output \g928/_0_  ;
  output \g929/_0_  ;
  output \g930/_0_  ;
  output \g9336/_0_  ;
  output \g9337/_0_  ;
  output \g939/_3_  ;
  output \g9396/_0_  ;
  output \g9397/_0_  ;
  output \g9399/_0_  ;
  output \g9400/_0_  ;
  output \g9401/_0_  ;
  output \g9402/_0_  ;
  output \g9403/_0_  ;
  output \g9404/_0_  ;
  output \g9415/_0_  ;
  output \g9418/_0_  ;
  output \g9419/_0_  ;
  output \g9420/_0_  ;
  output \g9446/_0_  ;
  output \g9465/_0_  ;
  output \g9493/_0_  ;
  output \g9536/_0_  ;
  output \g9537/_0_  ;
  output \g9538/_0_  ;
  output \g9539/_0_  ;
  output \g9540/_0_  ;
  output \g9541/_0_  ;
  output \g9542/_0_  ;
  output \g955/_2_  ;
  output \g9561/_0_  ;
  output \g9562/_0_  ;
  output \g9563/_0_  ;
  output \g9564/_0_  ;
  output \g9565/_0_  ;
  output \g9566/_0_  ;
  output \g9567/_0_  ;
  output \g9568/_0_  ;
  output \g9569/_0_  ;
  output \g9570/_0_  ;
  output \g9571/_0_  ;
  output \g9572/_0_  ;
  output \g9573/_0_  ;
  output \g9574/_0_  ;
  output \g9575/_0_  ;
  output \g9576/_0_  ;
  output \g9577/_0_  ;
  output \g9578/_0_  ;
  output \g9579/_0_  ;
  output \g9580/_0_  ;
  output \g9581/_0_  ;
  output \g9582/_0_  ;
  output \g9583/_0_  ;
  output \g9584/_0_  ;
  output \g9585/_0_  ;
  output \g9586/_0_  ;
  output \g9587/_0_  ;
  output \g9588/_0_  ;
  output \g9589/_0_  ;
  output \g9590/_0_  ;
  output \g9591/_0_  ;
  output \g9592/_0_  ;
  output \g9593/_0_  ;
  output \g9594/_0_  ;
  output \g9595/_0_  ;
  output \g9596/_0_  ;
  output \g9597/_0_  ;
  output \g9598/_0_  ;
  output \g9599/_0_  ;
  output \g9600/_0_  ;
  output \g9601/_0_  ;
  output \g9602/_0_  ;
  output \g9603/_0_  ;
  output \g9604/_0_  ;
  output \g9605/_0_  ;
  output \g9606/_0_  ;
  output \g9607/_0_  ;
  output \g9608/_0_  ;
  output \g9609/_0_  ;
  output \g9610/_0_  ;
  output \g9611/_0_  ;
  output \g9612/_0_  ;
  output \g9613/_0_  ;
  output \g9614/_0_  ;
  output \g9615/_0_  ;
  output \g9616/_0_  ;
  output \g9617/_0_  ;
  output \g9618/_0_  ;
  output \g9619/_0_  ;
  output \g9620/_0_  ;
  output \g9621/_0_  ;
  output \g9622/_0_  ;
  output \g9623/_0_  ;
  output \g9624/_0_  ;
  output \g9625/_0_  ;
  output \g9626/_0_  ;
  output \g9627/_0_  ;
  output \g9628/_0_  ;
  output \g9629/_0_  ;
  output \g9630/_0_  ;
  output \g9631/_0_  ;
  output \g9632/_0_  ;
  output \g9633/_0_  ;
  output \g9634/_0_  ;
  output \g9635/_0_  ;
  output \g9636/_0_  ;
  output \g9637/_0_  ;
  output \g9638/_0_  ;
  output \g9639/_0_  ;
  output \g9640/_0_  ;
  output \g9641/_0_  ;
  output \g9642/_0_  ;
  output \g9643/_0_  ;
  output \g9644/_0_  ;
  output \g9645/_0_  ;
  output \g9646/_0_  ;
  output \g9647/_0_  ;
  output \g9648/_0_  ;
  output \g9649/_0_  ;
  output \g9650/_0_  ;
  output \g9651/_0_  ;
  output \g9652/_0_  ;
  output \g9653/_0_  ;
  output \g9654/_0_  ;
  output \g9655/_0_  ;
  output \g9656/_0_  ;
  output \g9657/_0_  ;
  output \g9658/_0_  ;
  output \g9659/_0_  ;
  output \g9660/_0_  ;
  output \g9661/_0_  ;
  output \g9662/_0_  ;
  output \g9663/_0_  ;
  output \g9664/_0_  ;
  output \g9665/_0_  ;
  output \g9666/_0_  ;
  output \g9667/_0_  ;
  output \g9668/_0_  ;
  output \g9669/_0_  ;
  output \g9670/_0_  ;
  output \g9671/_0_  ;
  output \g9672/_0_  ;
  output \g9673/_0_  ;
  output \g9674/_0_  ;
  output \g9675/_0_  ;
  output \g9676/_0_  ;
  output \g9677/_0_  ;
  output \g9678/_0_  ;
  output \g9681/_0_  ;
  output \g9683/_0_  ;
  output \g9689/_0_  ;
  output \g9692/_0_  ;
  output \g9694/_0_  ;
  output \g9695/_0_  ;
  output \g9701/_0_  ;
  output \g9702/_0_  ;
  output \g9703/_0_  ;
  output \g9704/_0_  ;
  output \g9709/_0_  ;
  output \g9710/_0_  ;
  output \g9711/_0_  ;
  output \g9712/_0_  ;
  output \g9720/_0_  ;
  output \g9721/_0_  ;
  output \g9722/_0_  ;
  output \g9726/_0_  ;
  output \g9733/_0_  ;
  output \g9734/_0_  ;
  output \g9735/_0_  ;
  output \g9736/_0_  ;
  output \g9737/_0_  ;
  output \g9738/_0_  ;
  output \g9739/_0_  ;
  output \g9740/_0_  ;
  output \g9741/_0_  ;
  output \g9742/_0_  ;
  output \g9743/_0_  ;
  output \g9744/_0_  ;
  output \g9745/_0_  ;
  output \g9746/_0_  ;
  output \g9747/_0_  ;
  output \g9748/_0_  ;
  output \g9749/_0_  ;
  output \g9750/_0_  ;
  output \g9751/_0_  ;
  output \g9752/_0_  ;
  output \g9753/_0_  ;
  output \g9754/_0_  ;
  output \g9755/_0_  ;
  output \g9756/_0_  ;
  output \g9757/_0_  ;
  output \g9758/_0_  ;
  output \g9759/_0_  ;
  output \g9760/_0_  ;
  output \g9761/_0_  ;
  output \g9762/_0_  ;
  output \g9763/_0_  ;
  output \g9764/_0_  ;
  output \g9765/_0_  ;
  output \g9766/_0_  ;
  output \g9767/_0_  ;
  output \g9768/_0_  ;
  output \g9769/_0_  ;
  output \g9770/_0_  ;
  output \g9771/_0_  ;
  output \g9772/_0_  ;
  output \g9773/_0_  ;
  output \g9774/_0_  ;
  output \g9775/_0_  ;
  output \g9776/_0_  ;
  output \g9777/_0_  ;
  output \g9778/_0_  ;
  output \g9779/_0_  ;
  output \g9780/_0_  ;
  output \g9781/_0_  ;
  output \g9782/_0_  ;
  output \g9783/_0_  ;
  output \g9784/_0_  ;
  output \g9785/_0_  ;
  output \g9786/_0_  ;
  output \g9787/_0_  ;
  output \g9788/_0_  ;
  output \g9789/_0_  ;
  output \g9790/_0_  ;
  output \g9791/_0_  ;
  output \g9792/_0_  ;
  output \g9793/_0_  ;
  output \g9794/_0_  ;
  output \g9795/_0_  ;
  output \g9796/_0_  ;
  output \g9797/_0_  ;
  output \g9798/_0_  ;
  output \g9799/_0_  ;
  output \g9800/_0_  ;
  output \g9801/_0_  ;
  output \g9802/_0_  ;
  output \g9803/_0_  ;
  output \g9804/_0_  ;
  output \g9805/_0_  ;
  output \g9806/_0_  ;
  output \g9807/_0_  ;
  output \g9808/_0_  ;
  output \g9809/_0_  ;
  output \g9810/_0_  ;
  output \g9811/_0_  ;
  output \g9812/_0_  ;
  output \g9813/_0_  ;
  output \g9814/_0_  ;
  output \g9815/_0_  ;
  output \g9816/_0_  ;
  output \g9817/_0_  ;
  output \g9818/_0_  ;
  output \g9819/_0_  ;
  output \g9820/_0_  ;
  output \g9821/_0_  ;
  output \g9822/_0_  ;
  output \g9823/_0_  ;
  output \g9824/_0_  ;
  output \g9825/_0_  ;
  output \g9826/_0_  ;
  output \g9827/_0_  ;
  output \g9828/_0_  ;
  output \g9829/_0_  ;
  output \g9830/_0_  ;
  output \g9831/_0_  ;
  output \g9832/_0_  ;
  output \g9833/_0_  ;
  output \g9835/_0_  ;
  output \g9836/_0_  ;
  output \g9837/_0_  ;
  output \g9838/_0_  ;
  output \g9839/_0_  ;
  output \g9840/_0_  ;
  output \g9841/_0_  ;
  output \g9842/_0_  ;
  output \g9844/_0_  ;
  output \g9845/_0_  ;
  output \g9846/_0_  ;
  output \g9848/_0_  ;
  output \g9849/_0_  ;
  output \g9850/_0_  ;
  output \g9851/_0_  ;
  output \g9853/_0_  ;
  output \g9854/_0_  ;
  output \g9855/_0_  ;
  output \g9856/_0_  ;
  output \g9857/_0_  ;
  output \g9858/_0_  ;
  output \g9859/_0_  ;
  output \g9860/_0_  ;
  output \g9862/_0_  ;
  output \g9863/_0_  ;
  output \g9864/_0_  ;
  output \g9865/_0_  ;
  output \g9867/_0_  ;
  output \g9868/_0_  ;
  output \g9876/_0_  ;
  output \g9877/_0_  ;
  output \g9878/_0_  ;
  output \g9879/_0_  ;
  output \g9880/_0_  ;
  output \g9881/_0_  ;
  output \g9898/_0_  ;
  output \g9900/_0_  ;
  output \g9901/_0_  ;
  output \g9902/_0_  ;
  output \g9903/_0_  ;
  output \g9904/_0_  ;
  output \g9905/_0_  ;
  output \g9906/_0_  ;
  output \g9907/_0_  ;
  output \g9908/_0_  ;
  output \g9909/_0_  ;
  output \g9910/_0_  ;
  output \g9911/_0_  ;
  output \g9912/_0_  ;
  output \g9913/_0_  ;
  output \g9914/_0_  ;
  output \g9915/_0_  ;
  output \g9916/_0_  ;
  output \g9917/_0_  ;
  output \g9918/_0_  ;
  output \g9919/_0_  ;
  output \g992/_0_  ;
  output \g9920/_0_  ;
  output \g9921/_0_  ;
  output \g9922/_0_  ;
  output \g9923/_0_  ;
  output \g9924/_0_  ;
  output \g9925/_0_  ;
  output \g9926/_0_  ;
  output \g9927/_0_  ;
  output \g9928/_0_  ;
  output \g9929/_0_  ;
  output \g9930/_0_  ;
  output \g9931/_0_  ;
  output \g9932/_0_  ;
  output \g9933/_0_  ;
  output \g9934/_0_  ;
  output \g9935/_0_  ;
  output \g9936/_0_  ;
  output \g9937/_0_  ;
  output \g9938/_0_  ;
  output \g9939/_0_  ;
  output \g9940/_0_  ;
  output \g9941/_0_  ;
  output \g9942/_0_  ;
  output \g9943/_0_  ;
  output \g9944/_0_  ;
  output \g9945/_0_  ;
  output \g9946/_0_  ;
  output \g9947/_0_  ;
  output \g9948/_0_  ;
  output \g9949/_0_  ;
  output \g9950/_0_  ;
  output \g9951/_0_  ;
  output \g9952/_0_  ;
  output \g9953/_0_  ;
  output \g9954/_0_  ;
  output \g9955/_0_  ;
  output \g9956/_0_  ;
  output \g9957/_0_  ;
  output \g9958/_0_  ;
  output \g9959/_0_  ;
  output \g9960/_0_  ;
  output \g9961/_0_  ;
  output \g9962/_0_  ;
  output \g9963/_0_  ;
  output \g9964/_0_  ;
  output \g9965/_0_  ;
  output \g9966/_0_  ;
  output \g9967/_0_  ;
  output \g9968/_0_  ;
  output \g9969/_0_  ;
  output \g9970/_0_  ;
  output \g9971/_0_  ;
  output \g9972/_0_  ;
  output \g9973/_0_  ;
  output \g9974/_0_  ;
  output \g9975/_0_  ;
  output \g9976/_0_  ;
  output \g9977/_0_  ;
  output \g9978/_0_  ;
  output \g9979/_0_  ;
  output \g9980/_0_  ;
  output \g9981/_0_  ;
  output \g9982/_0_  ;
  output \g9983/_0_  ;
  output \g9984/_0_  ;
  output \g9985/_0_  ;
  output \g9987/_0_  ;
  output \g9988/_0_  ;
  output \g9989/_0_  ;
  output \g999/_0_  ;
  output \g9990/_0_  ;
  output \g9991/_0_  ;
  output \g9992/_0_  ;
  output \g9993/_0_  ;
  output \g9994/_0_  ;
  output \g9995/_0_  ;
  output \g9996/_0_  ;
  output \g9997/_0_  ;
  output \g9998/_0_  ;
  output \g9999/_0_  ;
  output \idma_IDMA_boot_reg/NET0131_reg_syn_3  ;
  output \memc_EXTC_Eg_reg/NET0131  ;
  output \memc_EXTC_Eg_reg/NET0131_reg_syn_3  ;
  output \memc_EXTC_Eg_reg/n0  ;
  output \pio_PIO_IN_P_reg[0]/P0001_reg_syn_3  ;
  output \pio_PIO_IN_P_reg[10]/P0001_reg_syn_3  ;
  output \pio_PIO_IN_P_reg[11]/P0001_reg_syn_3  ;
  output \pio_PIO_IN_P_reg[1]/P0001_reg_syn_3  ;
  output \pio_PIO_IN_P_reg[2]/P0001_reg_syn_3  ;
  output \pio_PIO_IN_P_reg[3]/P0001_reg_syn_3  ;
  output \pio_PIO_IN_P_reg[4]/P0001_reg_syn_3  ;
  output \pio_PIO_IN_P_reg[5]/P0001_reg_syn_3  ;
  output \pio_PIO_IN_P_reg[6]/P0001_reg_syn_3  ;
  output \pio_PIO_IN_P_reg[7]/P0001_reg_syn_3  ;
  output \pio_PIO_IN_P_reg[8]/P0001_reg_syn_3  ;
  output \pio_PIO_IN_P_reg[9]/P0001_reg_syn_3  ;
  output \pio_PIO_RES_OUT_reg[0]/P0001_reg_syn_3  ;
  output \pio_PIO_RES_OUT_reg[10]/P0001_reg_syn_3  ;
  output \pio_PIO_RES_OUT_reg[2]/P0001_reg_syn_3  ;
  output \pio_PIO_RES_OUT_reg[4]/P0001_reg_syn_3  ;
  output \pio_PIO_RES_OUT_reg[6]/P0001_reg_syn_3  ;
  output \sice_GO_NXi_reg/NET0131_reg_syn_3  ;
  output \sport0_rxctl_RXSHT_reg[0]/P0001_reg_syn_3  ;
  output \sport0_rxctl_RXSHT_reg[1]/P0001_reg_syn_3  ;
  output \sport1_rxctl_RXSHT_reg[0]/P0001_reg_syn_3  ;
  output \sport1_rxctl_RXSHT_reg[1]/P0001_reg_syn_3  ;
  wire n4047 , n4048 , n4049 , n4050 , n4051 , n4052 , n4053 , n4054 , n4055 , n4056 , n4057 , n4058 , n4059 , n4060 , n4061 , n4062 , n4063 , n4064 , n4065 , n4066 , n4067 , n4068 , n4069 , n4070 , n4071 , n4072 , n4073 , n4074 , n4075 , n4076 , n4077 , n4078 , n4079 , n4080 , n4081 , n4082 , n4083 , n4084 , n4085 , n4086 , n4087 , n4088 , n4089 , n4090 , n4091 , n4092 , n4093 , n4094 , n4095 , n4096 , n4097 , n4098 , n4099 , n4100 , n4101 , n4102 , n4103 , n4104 , n4105 , n4106 , n4107 , n4108 , n4109 , n4110 , n4111 , n4112 , n4113 , n4114 , n4115 , n4116 , n4117 , n4118 , n4119 , n4120 , n4121 , n4122 , n4123 , n4124 , n4125 , n4126 , n4127 , n4128 , n4129 , n4130 , n4131 , n4132 , n4133 , n4134 , n4135 , n4136 , n4137 , n4138 , n4139 , n4140 , n4141 , n4142 , n4143 , n4144 , n4145 , n4146 , n4147 , n4148 , n4149 , n4150 , n4151 , n4152 , n4153 , n4154 , n4155 , n4156 , n4157 , n4158 , n4159 , n4160 , n4161 , n4162 , n4163 , n4164 , n4165 , n4166 , n4167 , n4168 , n4169 , n4170 , n4171 , n4172 , n4173 , n4174 , n4175 , n4176 , n4177 , n4178 , n4179 , n4180 , n4181 , n4182 , n4183 , n4184 , n4185 , n4186 , n4187 , n4188 , n4189 , n4190 , n4191 , n4192 , n4193 , n4194 , n4195 , n4196 , n4197 , n4198 , n4199 , n4200 , n4201 , n4202 , n4203 , n4204 , n4205 , n4206 , n4207 , n4208 , n4209 , n4210 , n4211 , n4212 , n4213 , n4214 , n4215 , n4216 , n4217 , n4218 , n4219 , n4220 , n4221 , n4222 , n4223 , n4224 , n4225 , n4226 , n4227 , n4228 , n4229 , n4230 , n4231 , n4232 , n4233 , n4234 , n4235 , n4236 , n4237 , n4238 , n4239 , n4240 , n4241 , n4242 , n4243 , n4244 , n4245 , n4246 , n4247 , n4248 , n4249 , n4250 , n4251 , n4252 , n4253 , n4254 , n4255 , n4256 , n4257 , n4258 , n4259 , n4260 , n4261 , n4262 , n4263 , n4264 , n4265 , n4266 , n4267 , n4268 , n4269 , n4270 , n4271 , n4272 , n4273 , n4274 , n4275 , n4276 , n4277 , n4278 , n4279 , n4280 , n4281 , n4282 , n4283 , n4284 , n4285 , n4286 , n4287 , n4288 , n4289 , n4290 , n4291 , n4292 , n4293 , n4294 , n4295 , n4296 , n4297 , n4298 , n4299 , n4300 , n4301 , n4302 , n4303 , n4304 , n4305 , n4306 , n4307 , n4308 , n4309 , n4310 , n4311 , n4312 , n4313 , n4314 , n4315 , n4316 , n4317 , n4318 , n4319 , n4320 , n4321 , n4322 , n4323 , n4324 , n4325 , n4326 , n4327 , n4328 , n4329 , n4330 , n4331 , n4332 , n4333 , n4334 , n4335 , n4336 , n4337 , n4338 , n4339 , n4340 , n4341 , n4342 , n4343 , n4344 , n4345 , n4346 , n4347 , n4348 , n4349 , n4350 , n4351 , n4352 , n4353 , n4354 , n4355 , n4356 , n4357 , n4358 , n4359 , n4360 , n4361 , n4362 , n4363 , n4364 , n4365 , n4366 , n4367 , n4368 , n4369 , n4370 , n4371 , n4372 , n4373 , n4374 , n4375 , n4376 , n4377 , n4378 , n4379 , n4380 , n4381 , n4382 , n4383 , n4384 , n4385 , n4386 , n4387 , n4388 , n4389 , n4390 , n4391 , n4392 , n4393 , n4394 , n4395 , n4396 , n4397 , n4398 , n4399 , n4400 , n4401 , n4402 , n4403 , n4404 , n4405 , n4406 , n4407 , n4408 , n4409 , n4410 , n4411 , n4412 , n4413 , n4414 , n4415 , n4416 , n4417 , n4418 , n4419 , n4420 , n4421 , n4422 , n4423 , n4424 , n4425 , n4426 , n4427 , n4428 , n4429 , n4430 , n4431 , n4432 , n4433 , n4434 , n4435 , n4436 , n4437 , n4438 , n4439 , n4440 , n4441 , n4442 , n4443 , n4444 , n4445 , n4446 , n4447 , n4448 , n4449 , n4450 , n4451 , n4452 , n4453 , n4454 , n4455 , n4456 , n4457 , n4458 , n4459 , n4460 , n4461 , n4462 , n4463 , n4464 , n4465 , n4466 , n4467 , n4468 , n4469 , n4470 , n4471 , n4472 , n4473 , n4474 , n4475 , n4476 , n4477 , n4478 , n4479 , n4480 , n4481 , n4482 , n4483 , n4484 , n4485 , n4486 , n4487 , n4488 , n4489 , n4490 , n4491 , n4492 , n4493 , n4494 , n4495 , n4496 , n4497 , n4498 , n4499 , n4500 , n4501 , n4502 , n4503 , n4504 , n4505 , n4506 , n4507 , n4508 , n4509 , n4510 , n4511 , n4512 , n4513 , n4514 , n4515 , n4516 , n4517 , n4518 , n4519 , n4520 , n4521 , n4522 , n4523 , n4524 , n4525 , n4526 , n4527 , n4528 , n4529 , n4530 , n4531 , n4532 , n4533 , n4534 , n4535 , n4536 , n4537 , n4538 , n4539 , n4540 , n4541 , n4542 , n4543 , n4544 , n4545 , n4546 , n4547 , n4548 , n4549 , n4550 , n4551 , n4552 , n4553 , n4554 , n4555 , n4556 , n4557 , n4558 , n4559 , n4560 , n4561 , n4562 , n4563 , n4564 , n4565 , n4566 , n4567 , n4568 , n4569 , n4570 , n4571 , n4572 , n4573 , n4574 , n4575 , n4576 , n4577 , n4578 , n4579 , n4580 , n4581 , n4582 , n4583 , n4584 , n4585 , n4586 , n4587 , n4588 , n4589 , n4590 , n4591 , n4592 , n4593 , n4594 , n4595 , n4596 , n4597 , n4598 , n4599 , n4600 , n4601 , n4602 , n4603 , n4604 , n4605 , n4606 , n4607 , n4608 , n4609 , n4610 , n4611 , n4612 , n4613 , n4614 , n4615 , n4616 , n4617 , n4618 , n4619 , n4620 , n4621 , n4622 , n4623 , n4624 , n4625 , n4626 , n4627 , n4628 , n4629 , n4630 , n4631 , n4632 , n4633 , n4634 , n4635 , n4636 , n4637 , n4638 , n4639 , n4640 , n4641 , n4642 , n4643 , n4644 , n4645 , n4646 , n4647 , n4648 , n4649 , n4650 , n4651 , n4652 , n4653 , n4654 , n4655 , n4656 , n4657 , n4658 , n4659 , n4660 , n4661 , n4662 , n4663 , n4664 , n4665 , n4666 , n4667 , n4668 , n4669 , n4670 , n4671 , n4672 , n4673 , n4674 , n4675 , n4676 , n4677 , n4678 , n4679 , n4680 , n4681 , n4682 , n4683 , n4684 , n4685 , n4686 , n4687 , n4688 , n4689 , n4690 , n4691 , n4692 , n4693 , n4694 , n4695 , n4696 , n4697 , n4698 , n4699 , n4700 , n4701 , n4702 , n4703 , n4704 , n4705 , n4706 , n4707 , n4708 , n4709 , n4710 , n4711 , n4712 , n4713 , n4714 , n4715 , n4716 , n4717 , n4718 , n4719 , n4720 , n4721 , n4722 , n4723 , n4724 , n4725 , n4726 , n4727 , n4728 , n4729 , n4730 , n4731 , n4732 , n4733 , n4734 , n4735 , n4736 , n4737 , n4738 , n4739 , n4740 , n4741 , n4742 , n4743 , n4744 , n4745 , n4746 , n4747 , n4748 , n4749 , n4750 , n4751 , n4752 , n4753 , n4754 , n4755 , n4756 , n4757 , n4758 , n4759 , n4760 , n4761 , n4762 , n4763 , n4764 , n4765 , n4766 , n4767 , n4768 , n4769 , n4770 , n4771 , n4772 , n4773 , n4774 , n4775 , n4776 , n4777 , n4778 , n4779 , n4780 , n4781 , n4782 , n4783 , n4784 , n4785 , n4786 , n4787 , n4788 , n4789 , n4790 , n4791 , n4792 , n4793 , n4794 , n4795 , n4796 , n4797 , n4798 , n4799 , n4800 , n4801 , n4802 , n4803 , n4804 , n4805 , n4806 , n4807 , n4808 , n4809 , n4810 , n4811 , n4812 , n4813 , n4814 , n4815 , n4816 , n4817 , n4818 , n4819 , n4820 , n4821 , n4822 , n4823 , n4824 , n4825 , n4826 , n4827 , n4828 , n4829 , n4830 , n4831 , n4832 , n4833 , n4834 , n4835 , n4836 , n4837 , n4838 , n4839 , n4840 , n4841 , n4842 , n4843 , n4844 , n4845 , n4846 , n4847 , n4848 , n4849 , n4850 , n4851 , n4852 , n4853 , n4854 , n4855 , n4856 , n4857 , n4858 , n4859 , n4860 , n4861 , n4862 , n4863 , n4864 , n4865 , n4866 , n4867 , n4868 , n4869 , n4870 , n4871 , n4872 , n4873 , n4874 , n4875 , n4876 , n4877 , n4878 , n4879 , n4880 , n4881 , n4882 , n4883 , n4884 , n4885 , n4886 , n4887 , n4888 , n4889 , n4890 , n4891 , n4892 , n4893 , n4894 , n4895 , n4896 , n4897 , n4898 , n4899 , n4900 , n4901 , n4902 , n4903 , n4904 , n4905 , n4906 , n4907 , n4908 , n4909 , n4910 , n4911 , n4912 , n4913 , n4914 , n4915 , n4916 , n4917 , n4918 , n4919 , n4920 , n4921 , n4922 , n4923 , n4924 , n4925 , n4926 , n4927 , n4928 , n4929 , n4930 , n4931 , n4932 , n4933 , n4934 , n4935 , n4936 , n4937 , n4938 , n4939 , n4940 , n4941 , n4942 , n4943 , n4944 , n4945 , n4946 , n4947 , n4948 , n4949 , n4950 , n4951 , n4952 , n4953 , n4954 , n4955 , n4956 , n4957 , n4958 , n4959 , n4960 , n4961 , n4962 , n4963 , n4964 , n4965 , n4966 , n4967 , n4968 , n4969 , n4970 , n4971 , n4972 , n4973 , n4974 , n4975 , n4976 , n4977 , n4978 , n4979 , n4980 , n4981 , n4982 , n4983 , n4984 , n4985 , n4986 , n4987 , n4988 , n4989 , n4990 , n4991 , n4992 , n4993 , n4994 , n4995 , n4996 , n4997 , n4998 , n4999 , n5000 , n5001 , n5002 , n5003 , n5004 , n5005 , n5006 , n5007 , n5008 , n5009 , n5010 , n5011 , n5012 , n5013 , n5014 , n5015 , n5016 , n5017 , n5018 , n5019 , n5020 , n5021 , n5022 , n5023 , n5024 , n5025 , n5026 , n5027 , n5028 , n5029 , n5030 , n5031 , n5032 , n5033 , n5034 , n5035 , n5036 , n5037 , n5038 , n5039 , n5040 , n5041 , n5042 , n5043 , n5044 , n5045 , n5046 , n5047 , n5048 , n5049 , n5050 , n5051 , n5052 , n5053 , n5054 , n5055 , n5056 , n5057 , n5058 , n5059 , n5060 , n5061 , n5062 , n5063 , n5064 , n5065 , n5066 , n5067 , n5068 , n5069 , n5070 , n5071 , n5072 , n5073 , n5074 , n5075 , n5076 , n5077 , n5078 , n5079 , n5080 , n5081 , n5082 , n5083 , n5084 , n5085 , n5086 , n5087 , n5088 , n5089 , n5090 , n5091 , n5092 , n5093 , n5094 , n5095 , n5096 , n5097 , n5098 , n5099 , n5100 , n5101 , n5102 , n5103 , n5104 , n5105 , n5106 , n5107 , n5108 , n5109 , n5110 , n5111 , n5112 , n5113 , n5114 , n5115 , n5116 , n5117 , n5118 , n5119 , n5120 , n5121 , n5122 , n5123 , n5124 , n5125 , n5126 , n5127 , n5128 , n5129 , n5130 , n5131 , n5132 , n5133 , n5134 , n5135 , n5136 , n5137 , n5138 , n5139 , n5140 , n5141 , n5142 , n5143 , n5144 , n5145 , n5146 , n5147 , n5148 , n5149 , n5150 , n5151 , n5152 , n5153 , n5154 , n5155 , n5156 , n5157 , n5158 , n5159 , n5160 , n5161 , n5162 , n5163 , n5164 , n5165 , n5166 , n5167 , n5168 , n5169 , n5170 , n5171 , n5172 , n5173 , n5174 , n5175 , n5176 , n5177 , n5178 , n5179 , n5180 , n5181 , n5182 , n5183 , n5184 , n5185 , n5186 , n5187 , n5188 , n5189 , n5190 , n5191 , n5192 , n5193 , n5194 , n5195 , n5196 , n5197 , n5198 , n5199 , n5200 , n5201 , n5202 , n5203 , n5204 , n5205 , n5206 , n5207 , n5208 , n5209 , n5210 , n5211 , n5212 , n5213 , n5214 , n5215 , n5216 , n5217 , n5218 , n5219 , n5220 , n5221 , n5222 , n5223 , n5224 , n5225 , n5226 , n5227 , n5228 , n5229 , n5230 , n5231 , n5232 , n5233 , n5234 , n5235 , n5236 , n5237 , n5238 , n5239 , n5240 , n5241 , n5242 , n5243 , n5244 , n5245 , n5246 , n5247 , n5248 , n5249 , n5250 , n5251 , n5252 , n5253 , n5254 , n5255 , n5256 , n5257 , n5258 , n5259 , n5260 , n5261 , n5262 , n5263 , n5264 , n5265 , n5266 , n5267 , n5268 , n5269 , n5270 , n5271 , n5272 , n5273 , n5274 , n5275 , n5276 , n5277 , n5278 , n5279 , n5280 , n5281 , n5282 , n5283 , n5284 , n5285 , n5286 , n5287 , n5288 , n5289 , n5290 , n5291 , n5292 , n5293 , n5294 , n5295 , n5296 , n5297 , n5298 , n5299 , n5300 , n5301 , n5302 , n5303 , n5304 , n5305 , n5306 , n5307 , n5308 , n5309 , n5310 , n5311 , n5312 , n5313 , n5314 , n5315 , n5316 , n5317 , n5318 , n5319 , n5320 , n5321 , n5322 , n5323 , n5324 , n5325 , n5326 , n5327 , n5328 , n5329 , n5330 , n5331 , n5332 , n5333 , n5334 , n5335 , n5336 , n5337 , n5338 , n5339 , n5340 , n5341 , n5342 , n5343 , n5344 , n5345 , n5346 , n5347 , n5348 , n5349 , n5350 , n5351 , n5352 , n5353 , n5354 , n5355 , n5356 , n5357 , n5358 , n5359 , n5360 , n5361 , n5362 , n5363 , n5364 , n5365 , n5366 , n5367 , n5368 , n5369 , n5370 , n5371 , n5372 , n5373 , n5374 , n5375 , n5376 , n5377 , n5378 , n5379 , n5380 , n5381 , n5382 , n5383 , n5384 , n5385 , n5386 , n5387 , n5388 , n5389 , n5390 , n5391 , n5392 , n5393 , n5394 , n5395 , n5396 , n5397 , n5398 , n5399 , n5400 , n5401 , n5402 , n5403 , n5404 , n5405 , n5406 , n5407 , n5408 , n5409 , n5410 , n5411 , n5412 , n5413 , n5414 , n5415 , n5416 , n5417 , n5418 , n5419 , n5420 , n5421 , n5422 , n5423 , n5424 , n5425 , n5426 , n5427 , n5428 , n5429 , n5430 , n5431 , n5432 , n5433 , n5434 , n5435 , n5436 , n5437 , n5438 , n5439 , n5440 , n5441 , n5442 , n5443 , n5444 , n5445 , n5446 , n5447 , n5448 , n5449 , n5450 , n5451 , n5452 , n5453 , n5454 , n5455 , n5456 , n5457 , n5458 , n5459 , n5460 , n5461 , n5462 , n5463 , n5464 , n5465 , n5466 , n5467 , n5468 , n5469 , n5470 , n5471 , n5472 , n5473 , n5474 , n5475 , n5476 , n5477 , n5478 , n5479 , n5480 , n5481 , n5482 , n5483 , n5484 , n5485 , n5486 , n5487 , n5488 , n5489 , n5490 , n5491 , n5492 , n5493 , n5494 , n5495 , n5496 , n5497 , n5498 , n5499 , n5500 , n5501 , n5502 , n5503 , n5504 , n5505 , n5506 , n5507 , n5508 , n5509 , n5510 , n5511 , n5512 , n5513 , n5514 , n5515 , n5516 , n5517 , n5518 , n5519 , n5520 , n5521 , n5522 , n5523 , n5524 , n5525 , n5526 , n5527 , n5528 , n5529 , n5530 , n5531 , n5532 , n5533 , n5534 , n5535 , n5536 , n5537 , n5538 , n5539 , n5540 , n5541 , n5542 , n5543 , n5544 , n5545 , n5546 , n5547 , n5548 , n5549 , n5550 , n5551 , n5552 , n5553 , n5554 , n5555 , n5556 , n5557 , n5558 , n5559 , n5560 , n5561 , n5562 , n5563 , n5564 , n5565 , n5566 , n5567 , n5568 , n5569 , n5570 , n5571 , n5572 , n5573 , n5574 , n5575 , n5576 , n5577 , n5578 , n5579 , n5580 , n5581 , n5582 , n5583 , n5584 , n5585 , n5586 , n5587 , n5588 , n5589 , n5590 , n5591 , n5592 , n5593 , n5594 , n5595 , n5596 , n5597 , n5598 , n5599 , n5600 , n5601 , n5602 , n5603 , n5604 , n5605 , n5606 , n5607 , n5608 , n5609 , n5610 , n5611 , n5612 , n5613 , n5614 , n5615 , n5616 , n5617 , n5618 , n5619 , n5620 , n5621 , n5622 , n5623 , n5624 , n5625 , n5626 , n5627 , n5628 , n5629 , n5630 , n5631 , n5632 , n5633 , n5634 , n5635 , n5636 , n5637 , n5638 , n5639 , n5640 , n5641 , n5642 , n5643 , n5644 , n5645 , n5646 , n5647 , n5648 , n5649 , n5650 , n5651 , n5652 , n5653 , n5654 , n5655 , n5656 , n5657 , n5658 , n5659 , n5660 , n5661 , n5662 , n5663 , n5664 , n5665 , n5666 , n5667 , n5668 , n5669 , n5670 , n5671 , n5672 , n5673 , n5674 , n5675 , n5676 , n5677 , n5678 , n5679 , n5680 , n5681 , n5682 , n5683 , n5684 , n5685 , n5686 , n5687 , n5688 , n5689 , n5690 , n5691 , n5692 , n5693 , n5694 , n5695 , n5696 , n5697 , n5698 , n5699 , n5700 , n5701 , n5702 , n5703 , n5704 , n5705 , n5706 , n5707 , n5708 , n5709 , n5710 , n5711 , n5712 , n5713 , n5714 , n5715 , n5716 , n5717 , n5718 , n5719 , n5720 , n5721 , n5722 , n5723 , n5724 , n5725 , n5726 , n5727 , n5728 , n5729 , n5730 , n5731 , n5732 , n5733 , n5734 , n5735 , n5736 , n5737 , n5738 , n5739 , n5740 , n5741 , n5742 , n5743 , n5744 , n5745 , n5746 , n5747 , n5748 , n5749 , n5750 , n5751 , n5752 , n5753 , n5754 , n5755 , n5756 , n5757 , n5758 , n5759 , n5760 , n5761 , n5762 , n5763 , n5764 , n5765 , n5766 , n5767 , n5768 , n5769 , n5770 , n5771 , n5772 , n5773 , n5774 , n5775 , n5776 , n5777 , n5778 , n5779 , n5780 , n5781 , n5782 , n5783 , n5784 , n5785 , n5786 , n5787 , n5788 , n5789 , n5790 , n5791 , n5792 , n5793 , n5794 , n5795 , n5796 , n5797 , n5798 , n5799 , n5800 , n5801 , n5802 , n5803 , n5804 , n5805 , n5806 , n5807 , n5808 , n5809 , n5810 , n5811 , n5812 , n5813 , n5814 , n5815 , n5816 , n5817 , n5818 , n5819 , n5820 , n5821 , n5822 , n5823 , n5824 , n5825 , n5826 , n5827 , n5828 , n5829 , n5830 , n5831 , n5832 , n5833 , n5834 , n5835 , n5836 , n5837 , n5838 , n5839 , n5840 , n5841 , n5842 , n5843 , n5844 , n5845 , n5846 , n5847 , n5848 , n5849 , n5850 , n5851 , n5852 , n5853 , n5854 , n5855 , n5856 , n5857 , n5858 , n5859 , n5860 , n5861 , n5862 , n5863 , n5864 , n5865 , n5866 , n5867 , n5868 , n5869 , n5870 , n5871 , n5872 , n5873 , n5874 , n5875 , n5876 , n5877 , n5878 , n5879 , n5880 , n5881 , n5882 , n5883 , n5884 , n5885 , n5886 , n5887 , n5888 , n5889 , n5890 , n5891 , n5892 , n5893 , n5894 , n5895 , n5896 , n5897 , n5898 , n5899 , n5900 , n5901 , n5902 , n5903 , n5904 , n5905 , n5906 , n5907 , n5908 , n5909 , n5910 , n5911 , n5912 , n5913 , n5914 , n5915 , n5916 , n5917 , n5918 , n5919 , n5920 , n5921 , n5922 , n5923 , n5924 , n5925 , n5926 , n5927 , n5928 , n5929 , n5930 , n5931 , n5932 , n5933 , n5934 , n5935 , n5936 , n5937 , n5938 , n5939 , n5940 , n5941 , n5942 , n5943 , n5944 , n5945 , n5946 , n5947 , n5948 , n5949 , n5950 , n5951 , n5952 , n5953 , n5954 , n5955 , n5956 , n5957 , n5958 , n5959 , n5960 , n5961 , n5962 , n5963 , n5964 , n5965 , n5966 , n5967 , n5968 , n5969 , n5970 , n5971 , n5972 , n5973 , n5974 , n5975 , n5976 , n5977 , n5978 , n5979 , n5980 , n5981 , n5982 , n5983 , n5984 , n5985 , n5986 , n5987 , n5988 , n5989 , n5990 , n5991 , n5992 , n5993 , n5994 , n5995 , n5996 , n5997 , n5998 , n5999 , n6000 , n6001 , n6002 , n6003 , n6004 , n6005 , n6006 , n6007 , n6008 , n6009 , n6010 , n6011 , n6012 , n6013 , n6014 , n6015 , n6016 , n6017 , n6018 , n6019 , n6020 , n6021 , n6022 , n6023 , n6024 , n6025 , n6026 , n6027 , n6028 , n6029 , n6030 , n6031 , n6032 , n6033 , n6034 , n6035 , n6036 , n6037 , n6038 , n6039 , n6040 , n6041 , n6042 , n6043 , n6044 , n6045 , n6046 , n6047 , n6048 , n6049 , n6050 , n6051 , n6052 , n6053 , n6054 , n6055 , n6056 , n6057 , n6058 , n6059 , n6060 , n6061 , n6062 , n6063 , n6064 , n6065 , n6066 , n6067 , n6068 , n6069 , n6070 , n6071 , n6072 , n6073 , n6074 , n6075 , n6076 , n6077 , n6078 , n6079 , n6080 , n6081 , n6082 , n6083 , n6084 , n6085 , n6086 , n6087 , n6088 , n6089 , n6090 , n6091 , n6092 , n6093 , n6094 , n6095 , n6096 , n6097 , n6098 , n6099 , n6100 , n6101 , n6102 , n6103 , n6104 , n6105 , n6106 , n6107 , n6108 , n6109 , n6110 , n6111 , n6112 , n6113 , n6114 , n6115 , n6116 , n6117 , n6118 , n6119 , n6120 , n6121 , n6122 , n6123 , n6124 , n6125 , n6126 , n6127 , n6128 , n6129 , n6130 , n6131 , n6132 , n6133 , n6134 , n6135 , n6136 , n6137 , n6138 , n6139 , n6140 , n6141 , n6142 , n6143 , n6144 , n6145 , n6146 , n6147 , n6148 , n6149 , n6150 , n6151 , n6152 , n6153 , n6154 , n6155 , n6156 , n6157 , n6158 , n6159 , n6160 , n6161 , n6162 , n6163 , n6164 , n6165 , n6166 , n6167 , n6168 , n6169 , n6170 , n6171 , n6172 , n6173 , n6174 , n6175 , n6176 , n6177 , n6178 , n6179 , n6180 , n6181 , n6182 , n6183 , n6184 , n6185 , n6186 , n6187 , n6188 , n6189 , n6190 , n6191 , n6192 , n6193 , n6194 , n6195 , n6196 , n6197 , n6198 , n6199 , n6200 , n6201 , n6202 , n6203 , n6204 , n6205 , n6206 , n6207 , n6208 , n6209 , n6210 , n6211 , n6212 , n6213 , n6214 , n6215 , n6216 , n6217 , n6218 , n6219 , n6220 , n6221 , n6222 , n6223 , n6224 , n6225 , n6226 , n6227 , n6228 , n6229 , n6230 , n6231 , n6232 , n6233 , n6234 , n6235 , n6236 , n6237 , n6238 , n6239 , n6240 , n6241 , n6242 , n6243 , n6244 , n6245 , n6246 , n6247 , n6248 , n6249 , n6250 , n6251 , n6252 , n6253 , n6254 , n6255 , n6256 , n6257 , n6258 , n6259 , n6260 , n6261 , n6262 , n6263 , n6264 , n6265 , n6266 , n6267 , n6268 , n6269 , n6270 , n6271 , n6272 , n6273 , n6274 , n6275 , n6276 , n6277 , n6278 , n6279 , n6280 , n6281 , n6282 , n6283 , n6284 , n6285 , n6286 , n6287 , n6288 , n6289 , n6290 , n6291 , n6292 , n6293 , n6294 , n6295 , n6296 , n6297 , n6298 , n6299 , n6300 , n6301 , n6302 , n6303 , n6304 , n6305 , n6306 , n6307 , n6308 , n6309 , n6310 , n6311 , n6312 , n6313 , n6314 , n6315 , n6316 , n6317 , n6318 , n6319 , n6320 , n6321 , n6322 , n6323 , n6324 , n6325 , n6326 , n6327 , n6328 , n6329 , n6330 , n6331 , n6332 , n6333 , n6334 , n6335 , n6336 , n6337 , n6338 , n6339 , n6340 , n6341 , n6342 , n6343 , n6344 , n6345 , n6346 , n6347 , n6348 , n6349 , n6350 , n6351 , n6352 , n6353 , n6354 , n6355 , n6356 , n6357 , n6358 , n6359 , n6360 , n6361 , n6362 , n6363 , n6364 , n6365 , n6366 , n6367 , n6368 , n6369 , n6370 , n6371 , n6372 , n6373 , n6374 , n6375 , n6376 , n6377 , n6378 , n6379 , n6380 , n6381 , n6382 , n6383 , n6384 , n6385 , n6386 , n6387 , n6388 , n6389 , n6390 , n6391 , n6392 , n6393 , n6394 , n6395 , n6396 , n6397 , n6398 , n6399 , n6400 , n6401 , n6402 , n6403 , n6404 , n6405 , n6406 , n6407 , n6408 , n6409 , n6410 , n6411 , n6412 , n6413 , n6414 , n6415 , n6416 , n6417 , n6418 , n6419 , n6420 , n6421 , n6422 , n6423 , n6424 , n6425 , n6426 , n6427 , n6428 , n6429 , n6430 , n6431 , n6432 , n6433 , n6434 , n6435 , n6436 , n6437 , n6438 , n6439 , n6440 , n6441 , n6442 , n6443 , n6444 , n6445 , n6446 , n6447 , n6448 , n6449 , n6450 , n6451 , n6452 , n6453 , n6454 , n6455 , n6456 , n6457 , n6458 , n6459 , n6460 , n6461 , n6462 , n6463 , n6464 , n6465 , n6466 , n6467 , n6468 , n6469 , n6470 , n6471 , n6472 , n6473 , n6474 , n6475 , n6476 , n6477 , n6478 , n6479 , n6480 , n6481 , n6482 , n6483 , n6484 , n6485 , n6486 , n6487 , n6488 , n6489 , n6490 , n6491 , n6492 , n6493 , n6494 , n6495 , n6496 , n6497 , n6498 , n6499 , n6500 , n6501 , n6502 , n6503 , n6504 , n6505 , n6506 , n6507 , n6508 , n6509 , n6510 , n6511 , n6512 , n6513 , n6514 , n6515 , n6516 , n6517 , n6518 , n6519 , n6520 , n6521 , n6522 , n6523 , n6524 , n6525 , n6526 , n6527 , n6528 , n6529 , n6530 , n6531 , n6532 , n6533 , n6534 , n6535 , n6536 , n6537 , n6538 , n6539 , n6540 , n6541 , n6542 , n6543 , n6544 , n6545 , n6546 , n6547 , n6548 , n6549 , n6550 , n6551 , n6552 , n6553 , n6554 , n6555 , n6556 , n6557 , n6558 , n6559 , n6560 , n6561 , n6562 , n6563 , n6564 , n6565 , n6566 , n6567 , n6568 , n6569 , n6570 , n6571 , n6572 , n6573 , n6574 , n6575 , n6576 , n6577 , n6578 , n6579 , n6580 , n6581 , n6582 , n6583 , n6584 , n6585 , n6586 , n6587 , n6588 , n6589 , n6590 , n6591 , n6592 , n6593 , n6594 , n6595 , n6596 , n6597 , n6598 , n6599 , n6600 , n6601 , n6602 , n6603 , n6604 , n6605 , n6606 , n6607 , n6608 , n6609 , n6610 , n6611 , n6612 , n6613 , n6614 , n6615 , n6616 , n6617 , n6618 , n6619 , n6620 , n6621 , n6622 , n6623 , n6624 , n6625 , n6626 , n6627 , n6628 , n6629 , n6630 , n6631 , n6632 , n6633 , n6634 , n6635 , n6636 , n6637 , n6638 , n6639 , n6640 , n6641 , n6642 , n6643 , n6644 , n6645 , n6646 , n6647 , n6648 , n6649 , n6650 , n6651 , n6652 , n6653 , n6654 , n6655 , n6656 , n6657 , n6658 , n6659 , n6660 , n6661 , n6662 , n6663 , n6664 , n6665 , n6666 , n6667 , n6668 , n6669 , n6670 , n6671 , n6672 , n6673 , n6674 , n6675 , n6676 , n6677 , n6678 , n6679 , n6680 , n6681 , n6682 , n6683 , n6684 , n6685 , n6686 , n6687 , n6688 , n6689 , n6690 , n6691 , n6692 , n6693 , n6694 , n6695 , n6696 , n6697 , n6698 , n6699 , n6700 , n6701 , n6702 , n6703 , n6704 , n6705 , n6706 , n6707 , n6708 , n6709 , n6710 , n6711 , n6712 , n6713 , n6714 , n6715 , n6716 , n6717 , n6718 , n6719 , n6720 , n6721 , n6722 , n6723 , n6724 , n6725 , n6726 , n6727 , n6728 , n6729 , n6730 , n6731 , n6732 , n6733 , n6734 , n6735 , n6736 , n6737 , n6738 , n6739 , n6740 , n6741 , n6742 , n6743 , n6744 , n6745 , n6746 , n6747 , n6748 , n6749 , n6750 , n6751 , n6752 , n6753 , n6754 , n6755 , n6756 , n6757 , n6758 , n6759 , n6760 , n6761 , n6762 , n6763 , n6764 , n6765 , n6766 , n6767 , n6768 , n6769 , n6770 , n6771 , n6772 , n6773 , n6774 , n6775 , n6776 , n6777 , n6778 , n6779 , n6780 , n6781 , n6782 , n6783 , n6784 , n6785 , n6786 , n6787 , n6788 , n6789 , n6790 , n6791 , n6792 , n6793 , n6794 , n6795 , n6796 , n6797 , n6798 , n6799 , n6800 , n6801 , n6802 , n6803 , n6804 , n6805 , n6806 , n6807 , n6808 , n6809 , n6810 , n6811 , n6812 , n6813 , n6814 , n6815 , n6816 , n6817 , n6818 , n6819 , n6820 , n6821 , n6822 , n6823 , n6824 , n6825 , n6826 , n6827 , n6828 , n6829 , n6830 , n6831 , n6832 , n6833 , n6834 , n6835 , n6836 , n6837 , n6838 , n6839 , n6840 , n6841 , n6842 , n6843 , n6844 , n6845 , n6846 , n6847 , n6848 , n6849 , n6850 , n6851 , n6852 , n6853 , n6854 , n6855 , n6856 , n6857 , n6858 , n6859 , n6860 , n6861 , n6862 , n6863 , n6864 , n6865 , n6866 , n6867 , n6868 , n6869 , n6870 , n6871 , n6872 , n6873 , n6874 , n6875 , n6876 , n6877 , n6878 , n6879 , n6880 , n6881 , n6882 , n6883 , n6884 , n6885 , n6886 , n6887 , n6888 , n6889 , n6890 , n6891 , n6892 , n6893 , n6894 , n6895 , n6896 , n6897 , n6898 , n6899 , n6900 , n6901 , n6902 , n6903 , n6904 , n6905 , n6906 , n6907 , n6908 , n6909 , n6910 , n6911 , n6912 , n6913 , n6914 , n6915 , n6916 , n6917 , n6918 , n6919 , n6920 , n6921 , n6922 , n6923 , n6924 , n6925 , n6926 , n6927 , n6928 , n6929 , n6930 , n6931 , n6932 , n6933 , n6934 , n6935 , n6936 , n6937 , n6938 , n6939 , n6940 , n6941 , n6942 , n6943 , n6944 , n6945 , n6946 , n6947 , n6948 , n6949 , n6950 , n6951 , n6952 , n6953 , n6954 , n6955 , n6956 , n6957 , n6958 , n6959 , n6960 , n6961 , n6962 , n6963 , n6964 , n6965 , n6966 , n6967 , n6968 , n6969 , n6970 , n6971 , n6972 , n6973 , n6974 , n6975 , n6976 , n6977 , n6978 , n6979 , n6980 , n6981 , n6982 , n6983 , n6984 , n6985 , n6986 , n6987 , n6988 , n6989 , n6990 , n6991 , n6992 , n6993 , n6994 , n6995 , n6996 , n6997 , n6998 , n6999 , n7000 , n7001 , n7002 , n7003 , n7004 , n7005 , n7006 , n7007 , n7008 , n7009 , n7010 , n7011 , n7012 , n7013 , n7014 , n7015 , n7016 , n7017 , n7018 , n7019 , n7020 , n7021 , n7022 , n7023 , n7024 , n7025 , n7026 , n7027 , n7028 , n7029 , n7030 , n7031 , n7032 , n7033 , n7034 , n7035 , n7036 , n7037 , n7038 , n7039 , n7040 , n7041 , n7042 , n7043 , n7044 , n7045 , n7046 , n7047 , n7048 , n7049 , n7050 , n7051 , n7052 , n7053 , n7054 , n7055 , n7056 , n7057 , n7058 , n7059 , n7060 , n7061 , n7062 , n7063 , n7064 , n7065 , n7066 , n7067 , n7068 , n7069 , n7070 , n7071 , n7072 , n7073 , n7074 , n7075 , n7076 , n7077 , n7078 , n7079 , n7080 , n7081 , n7082 , n7083 , n7084 , n7085 , n7086 , n7087 , n7088 , n7089 , n7090 , n7091 , n7092 , n7093 , n7094 , n7095 , n7096 , n7097 , n7098 , n7099 , n7100 , n7101 , n7102 , n7103 , n7104 , n7105 , n7106 , n7107 , n7108 , n7109 , n7110 , n7111 , n7112 , n7113 , n7114 , n7115 , n7116 , n7117 , n7118 , n7119 , n7120 , n7121 , n7122 , n7123 , n7124 , n7125 , n7126 , n7127 , n7128 , n7129 , n7130 , n7131 , n7132 , n7133 , n7134 , n7135 , n7136 , n7137 , n7138 , n7139 , n7140 , n7141 , n7142 , n7143 , n7144 , n7145 , n7146 , n7147 , n7148 , n7149 , n7150 , n7151 , n7152 , n7153 , n7154 , n7155 , n7156 , n7157 , n7158 , n7159 , n7160 , n7161 , n7162 , n7163 , n7164 , n7165 , n7166 , n7167 , n7168 , n7169 , n7170 , n7171 , n7172 , n7173 , n7174 , n7175 , n7176 , n7177 , n7178 , n7179 , n7180 , n7181 , n7182 , n7183 , n7184 , n7185 , n7186 , n7187 , n7188 , n7189 , n7190 , n7191 , n7192 , n7193 , n7194 , n7195 , n7196 , n7197 , n7198 , n7199 , n7200 , n7201 , n7202 , n7203 , n7204 , n7205 , n7206 , n7207 , n7208 , n7209 , n7210 , n7211 , n7212 , n7213 , n7214 , n7215 , n7216 , n7217 , n7218 , n7219 , n7220 , n7221 , n7222 , n7223 , n7224 , n7225 , n7226 , n7227 , n7228 , n7229 , n7230 , n7231 , n7232 , n7233 , n7234 , n7235 , n7236 , n7237 , n7238 , n7239 , n7240 , n7241 , n7242 , n7243 , n7244 , n7245 , n7246 , n7247 , n7248 , n7249 , n7250 , n7251 , n7252 , n7253 , n7254 , n7255 , n7256 , n7257 , n7258 , n7259 , n7260 , n7261 , n7262 , n7263 , n7264 , n7265 , n7266 , n7267 , n7268 , n7269 , n7270 , n7271 , n7272 , n7273 , n7274 , n7275 , n7276 , n7277 , n7278 , n7279 , n7280 , n7281 , n7282 , n7283 , n7284 , n7285 , n7286 , n7287 , n7288 , n7289 , n7290 , n7291 , n7292 , n7293 , n7294 , n7295 , n7296 , n7297 , n7298 , n7299 , n7300 , n7301 , n7302 , n7303 , n7304 , n7305 , n7306 , n7307 , n7308 , n7309 , n7310 , n7311 , n7312 , n7313 , n7314 , n7315 , n7316 , n7317 , n7318 , n7319 , n7320 , n7321 , n7322 , n7323 , n7324 , n7325 , n7326 , n7327 , n7328 , n7329 , n7330 , n7331 , n7332 , n7333 , n7334 , n7335 , n7336 , n7337 , n7338 , n7339 , n7340 , n7341 , n7342 , n7343 , n7344 , n7345 , n7346 , n7347 , n7348 , n7349 , n7350 , n7351 , n7352 , n7353 , n7354 , n7355 , n7356 , n7357 , n7358 , n7359 , n7360 , n7361 , n7362 , n7363 , n7364 , n7365 , n7366 , n7367 , n7368 , n7369 , n7370 , n7371 , n7372 , n7373 , n7374 , n7375 , n7376 , n7377 , n7378 , n7379 , n7380 , n7381 , n7382 , n7383 , n7384 , n7385 , n7386 , n7387 , n7388 , n7389 , n7390 , n7391 , n7392 , n7393 , n7394 , n7395 , n7396 , n7397 , n7398 , n7399 , n7400 , n7401 , n7402 , n7403 , n7404 , n7405 , n7406 , n7407 , n7408 , n7409 , n7410 , n7411 , n7412 , n7413 , n7414 , n7415 , n7416 , n7417 , n7418 , n7419 , n7420 , n7421 , n7422 , n7423 , n7424 , n7425 , n7426 , n7427 , n7428 , n7429 , n7430 , n7431 , n7432 , n7433 , n7434 , n7435 , n7436 , n7437 , n7438 , n7439 , n7440 , n7441 , n7442 , n7443 , n7444 , n7445 , n7446 , n7447 , n7448 , n7449 , n7450 , n7451 , n7452 , n7453 , n7454 , n7455 , n7456 , n7457 , n7458 , n7459 , n7460 , n7461 , n7462 , n7463 , n7464 , n7465 , n7466 , n7467 , n7468 , n7469 , n7470 , n7471 , n7472 , n7473 , n7474 , n7475 , n7476 , n7477 , n7478 , n7479 , n7480 , n7481 , n7482 , n7483 , n7484 , n7485 , n7486 , n7487 , n7488 , n7489 , n7490 , n7491 , n7492 , n7493 , n7494 , n7495 , n7496 , n7497 , n7498 , n7499 , n7500 , n7501 , n7502 , n7503 , n7504 , n7505 , n7506 , n7507 , n7508 , n7509 , n7510 , n7511 , n7512 , n7513 , n7514 , n7515 , n7516 , n7517 , n7518 , n7519 , n7520 , n7521 , n7522 , n7523 , n7524 , n7525 , n7526 , n7527 , n7528 , n7529 , n7530 , n7531 , n7532 , n7533 , n7534 , n7535 , n7536 , n7537 , n7538 , n7539 , n7540 , n7541 , n7542 , n7543 , n7544 , n7545 , n7546 , n7547 , n7548 , n7549 , n7550 , n7551 , n7552 , n7553 , n7554 , n7555 , n7556 , n7557 , n7558 , n7559 , n7560 , n7561 , n7562 , n7563 , n7564 , n7565 , n7566 , n7567 , n7568 , n7569 , n7570 , n7571 , n7572 , n7573 , n7574 , n7575 , n7576 , n7577 , n7578 , n7579 , n7580 , n7581 , n7582 , n7583 , n7584 , n7585 , n7586 , n7587 , n7588 , n7589 , n7590 , n7591 , n7592 , n7593 , n7594 , n7595 , n7596 , n7597 , n7598 , n7599 , n7600 , n7601 , n7602 , n7603 , n7604 , n7605 , n7606 , n7607 , n7608 , n7609 , n7610 , n7611 , n7612 , n7613 , n7614 , n7615 , n7616 , n7617 , n7618 , n7619 , n7620 , n7621 , n7622 , n7623 , n7624 , n7625 , n7626 , n7627 , n7628 , n7629 , n7630 , n7631 , n7632 , n7633 , n7634 , n7635 , n7636 , n7637 , n7638 , n7639 , n7640 , n7641 , n7642 , n7643 , n7644 , n7645 , n7646 , n7647 , n7648 , n7649 , n7650 , n7651 , n7652 , n7653 , n7654 , n7655 , n7656 , n7657 , n7658 , n7659 , n7660 , n7661 , n7662 , n7663 , n7664 , n7665 , n7666 , n7667 , n7668 , n7669 , n7670 , n7671 , n7672 , n7673 , n7674 , n7675 , n7676 , n7677 , n7678 , n7679 , n7680 , n7681 , n7682 , n7683 , n7684 , n7685 , n7686 , n7687 , n7688 , n7689 , n7690 , n7691 , n7692 , n7693 , n7694 , n7695 , n7696 , n7697 , n7698 , n7699 , n7700 , n7701 , n7702 , n7703 , n7704 , n7705 , n7706 , n7707 , n7708 , n7709 , n7710 , n7711 , n7712 , n7713 , n7714 , n7715 , n7716 , n7717 , n7718 , n7719 , n7720 , n7721 , n7722 , n7723 , n7724 , n7725 , n7726 , n7727 , n7728 , n7729 , n7730 , n7731 , n7732 , n7733 , n7734 , n7735 , n7736 , n7737 , n7738 , n7739 , n7740 , n7741 , n7742 , n7743 , n7744 , n7745 , n7746 , n7747 , n7748 , n7749 , n7750 , n7751 , n7752 , n7753 , n7754 , n7755 , n7756 , n7757 , n7758 , n7759 , n7760 , n7761 , n7762 , n7763 , n7764 , n7765 , n7766 , n7767 , n7768 , n7769 , n7770 , n7771 , n7772 , n7773 , n7774 , n7775 , n7776 , n7777 , n7778 , n7779 , n7780 , n7781 , n7782 , n7783 , n7784 , n7785 , n7786 , n7787 , n7788 , n7789 , n7790 , n7791 , n7792 , n7793 , n7794 , n7795 , n7796 , n7797 , n7798 , n7799 , n7800 , n7801 , n7802 , n7803 , n7804 , n7805 , n7806 , n7807 , n7808 , n7809 , n7810 , n7811 , n7812 , n7813 , n7814 , n7815 , n7816 , n7817 , n7818 , n7819 , n7820 , n7821 , n7822 , n7823 , n7824 , n7825 , n7826 , n7827 , n7828 , n7829 , n7830 , n7831 , n7832 , n7833 , n7834 , n7835 , n7836 , n7837 , n7838 , n7839 , n7840 , n7841 , n7842 , n7843 , n7844 , n7845 , n7846 , n7847 , n7848 , n7849 , n7850 , n7851 , n7852 , n7853 , n7854 , n7855 , n7856 , n7857 , n7858 , n7859 , n7860 , n7861 , n7862 , n7863 , n7864 , n7865 , n7866 , n7867 , n7868 , n7869 , n7870 , n7871 , n7872 , n7873 , n7874 , n7875 , n7876 , n7877 , n7878 , n7879 , n7880 , n7881 , n7882 , n7883 , n7884 , n7885 , n7886 , n7887 , n7888 , n7889 , n7890 , n7891 , n7892 , n7893 , n7894 , n7895 , n7896 , n7897 , n7898 , n7899 , n7900 , n7901 , n7902 , n7903 , n7904 , n7905 , n7906 , n7907 , n7908 , n7909 , n7910 , n7911 , n7912 , n7913 , n7914 , n7915 , n7916 , n7917 , n7918 , n7919 , n7920 , n7921 , n7922 , n7923 , n7924 , n7925 , n7926 , n7927 , n7928 , n7929 , n7930 , n7931 , n7932 , n7933 , n7934 , n7935 , n7936 , n7937 , n7938 , n7939 , n7940 , n7941 , n7942 , n7943 , n7944 , n7945 , n7946 , n7947 , n7948 , n7949 , n7950 , n7951 , n7952 , n7953 , n7954 , n7955 , n7956 , n7957 , n7958 , n7959 , n7960 , n7961 , n7962 , n7963 , n7964 , n7965 , n7966 , n7967 , n7968 , n7969 , n7970 , n7971 , n7972 , n7973 , n7974 , n7975 , n7976 , n7977 , n7978 , n7979 , n7980 , n7981 , n7982 , n7983 , n7984 , n7985 , n7986 , n7987 , n7988 , n7989 , n7990 , n7991 , n7992 , n7993 , n7994 , n7995 , n7996 , n7997 , n7998 , n7999 , n8000 , n8001 , n8002 , n8003 , n8004 , n8005 , n8006 , n8007 , n8008 , n8009 , n8010 , n8011 , n8012 , n8013 , n8014 , n8015 , n8016 , n8017 , n8018 , n8019 , n8020 , n8021 , n8022 , n8023 , n8024 , n8025 , n8026 , n8027 , n8028 , n8029 , n8030 , n8031 , n8032 , n8033 , n8034 , n8035 , n8036 , n8037 , n8038 , n8039 , n8040 , n8041 , n8042 , n8043 , n8044 , n8045 , n8046 , n8047 , n8048 , n8049 , n8050 , n8051 , n8052 , n8053 , n8054 , n8055 , n8056 , n8057 , n8058 , n8059 , n8060 , n8061 , n8062 , n8063 , n8064 , n8065 , n8066 , n8067 , n8068 , n8069 , n8070 , n8071 , n8072 , n8073 , n8074 , n8075 , n8076 , n8077 , n8078 , n8079 , n8080 , n8081 , n8082 , n8083 , n8084 , n8085 , n8086 , n8087 , n8088 , n8089 , n8090 , n8091 , n8092 , n8093 , n8094 , n8095 , n8096 , n8097 , n8098 , n8099 , n8100 , n8101 , n8102 , n8103 , n8104 , n8105 , n8106 , n8107 , n8108 , n8109 , n8110 , n8111 , n8112 , n8113 , n8114 , n8115 , n8116 , n8117 , n8118 , n8119 , n8120 , n8121 , n8122 , n8123 , n8124 , n8125 , n8126 , n8127 , n8128 , n8129 , n8130 , n8131 , n8132 , n8133 , n8134 , n8135 , n8136 , n8137 , n8138 , n8139 , n8140 , n8141 , n8142 , n8143 , n8144 , n8145 , n8146 , n8147 , n8148 , n8149 , n8150 , n8151 , n8152 , n8153 , n8154 , n8155 , n8156 , n8157 , n8158 , n8159 , n8160 , n8161 , n8162 , n8163 , n8164 , n8165 , n8166 , n8167 , n8168 , n8169 , n8170 , n8171 , n8172 , n8173 , n8174 , n8175 , n8176 , n8177 , n8178 , n8179 , n8180 , n8181 , n8182 , n8183 , n8184 , n8185 , n8186 , n8187 , n8188 , n8189 , n8190 , n8191 , n8192 , n8193 , n8194 , n8195 , n8196 , n8197 , n8198 , n8199 , n8200 , n8201 , n8202 , n8203 , n8204 , n8205 , n8206 , n8207 , n8208 , n8209 , n8210 , n8211 , n8212 , n8213 , n8214 , n8215 , n8216 , n8217 , n8218 , n8219 , n8220 , n8221 , n8222 , n8223 , n8224 , n8225 , n8226 , n8227 , n8228 , n8229 , n8230 , n8231 , n8232 , n8233 , n8234 , n8235 , n8236 , n8237 , n8238 , n8239 , n8240 , n8241 , n8242 , n8243 , n8244 , n8245 , n8246 , n8247 , n8248 , n8249 , n8250 , n8251 , n8252 , n8253 , n8254 , n8255 , n8256 , n8257 , n8258 , n8259 , n8260 , n8261 , n8262 , n8263 , n8264 , n8265 , n8266 , n8267 , n8268 , n8269 , n8270 , n8271 , n8272 , n8273 , n8274 , n8275 , n8276 , n8277 , n8278 , n8279 , n8280 , n8281 , n8282 , n8283 , n8284 , n8285 , n8286 , n8287 , n8288 , n8289 , n8290 , n8291 , n8292 , n8293 , n8294 , n8295 , n8296 , n8297 , n8298 , n8299 , n8300 , n8301 , n8302 , n8303 , n8304 , n8305 , n8306 , n8307 , n8308 , n8309 , n8310 , n8311 , n8312 , n8313 , n8314 , n8315 , n8316 , n8317 , n8318 , n8319 , n8320 , n8321 , n8322 , n8323 , n8324 , n8325 , n8326 , n8327 , n8328 , n8329 , n8330 , n8331 , n8332 , n8333 , n8334 , n8335 , n8336 , n8337 , n8338 , n8339 , n8340 , n8341 , n8342 , n8343 , n8344 , n8345 , n8346 , n8347 , n8348 , n8349 , n8350 , n8351 , n8352 , n8353 , n8354 , n8355 , n8356 , n8357 , n8358 , n8359 , n8360 , n8361 , n8362 , n8363 , n8364 , n8365 , n8366 , n8367 , n8368 , n8369 , n8370 , n8371 , n8372 , n8373 , n8374 , n8375 , n8376 , n8377 , n8378 , n8379 , n8380 , n8381 , n8382 , n8383 , n8384 , n8385 , n8386 , n8387 , n8388 , n8389 , n8390 , n8391 , n8392 , n8393 , n8394 , n8395 , n8396 , n8397 , n8398 , n8399 , n8400 , n8401 , n8402 , n8403 , n8404 , n8405 , n8406 , n8407 , n8408 , n8409 , n8410 , n8411 , n8412 , n8413 , n8414 , n8415 , n8416 , n8417 , n8418 , n8419 , n8420 , n8421 , n8422 , n8423 , n8424 , n8425 , n8426 , n8427 , n8428 , n8429 , n8430 , n8431 , n8432 , n8433 , n8434 , n8435 , n8436 , n8437 , n8438 , n8439 , n8440 , n8441 , n8442 , n8443 , n8444 , n8445 , n8446 , n8447 , n8448 , n8449 , n8450 , n8451 , n8452 , n8453 , n8454 , n8455 , n8456 , n8457 , n8458 , n8459 , n8460 , n8461 , n8462 , n8463 , n8464 , n8465 , n8466 , n8467 , n8468 , n8469 , n8470 , n8471 , n8472 , n8473 , n8474 , n8475 , n8476 , n8477 , n8478 , n8479 , n8480 , n8481 , n8482 , n8483 , n8484 , n8485 , n8486 , n8487 , n8488 , n8489 , n8490 , n8491 , n8492 , n8493 , n8494 , n8495 , n8496 , n8497 , n8498 , n8499 , n8500 , n8501 , n8502 , n8503 , n8504 , n8505 , n8506 , n8507 , n8508 , n8509 , n8510 , n8511 , n8512 , n8513 , n8514 , n8515 , n8516 , n8517 , n8518 , n8519 , n8520 , n8521 , n8522 , n8523 , n8524 , n8525 , n8526 , n8527 , n8528 , n8529 , n8530 , n8531 , n8532 , n8533 , n8534 , n8535 , n8536 , n8537 , n8538 , n8539 , n8540 , n8541 , n8542 , n8543 , n8544 , n8545 , n8546 , n8547 , n8548 , n8549 , n8550 , n8551 , n8552 , n8553 , n8554 , n8555 , n8556 , n8557 , n8558 , n8559 , n8560 , n8561 , n8562 , n8563 , n8564 , n8565 , n8566 , n8567 , n8568 , n8569 , n8570 , n8571 , n8572 , n8573 , n8574 , n8575 , n8576 , n8577 , n8578 , n8579 , n8580 , n8581 , n8582 , n8583 , n8584 , n8585 , n8586 , n8587 , n8588 , n8589 , n8590 , n8591 , n8592 , n8593 , n8594 , n8595 , n8596 , n8597 , n8598 , n8599 , n8600 , n8601 , n8602 , n8603 , n8604 , n8605 , n8606 , n8607 , n8608 , n8609 , n8610 , n8611 , n8612 , n8613 , n8614 , n8615 , n8616 , n8617 , n8618 , n8619 , n8620 , n8621 , n8622 , n8623 , n8624 , n8625 , n8626 , n8627 , n8628 , n8629 , n8630 , n8631 , n8632 , n8633 , n8634 , n8635 , n8636 , n8637 , n8638 , n8639 , n8640 , n8641 , n8642 , n8643 , n8644 , n8645 , n8646 , n8647 , n8648 , n8649 , n8650 , n8651 , n8652 , n8653 , n8654 , n8655 , n8656 , n8657 , n8658 , n8659 , n8660 , n8661 , n8662 , n8663 , n8664 , n8665 , n8666 , n8667 , n8668 , n8669 , n8670 , n8671 , n8672 , n8673 , n8674 , n8675 , n8676 , n8677 , n8678 , n8679 , n8680 , n8681 , n8682 , n8683 , n8684 , n8685 , n8686 , n8687 , n8688 , n8689 , n8690 , n8691 , n8692 , n8693 , n8694 , n8695 , n8696 , n8697 , n8698 , n8699 , n8700 , n8701 , n8702 , n8703 , n8704 , n8705 , n8706 , n8707 , n8708 , n8709 , n8710 , n8711 , n8712 , n8713 , n8714 , n8715 , n8716 , n8717 , n8718 , n8719 , n8720 , n8721 , n8722 , n8723 , n8724 , n8725 , n8726 , n8727 , n8728 , n8729 , n8730 , n8731 , n8732 , n8733 , n8734 , n8735 , n8736 , n8737 , n8738 , n8739 , n8740 , n8741 , n8742 , n8743 , n8744 , n8745 , n8746 , n8747 , n8748 , n8749 , n8750 , n8751 , n8752 , n8753 , n8754 , n8755 , n8756 , n8757 , n8758 , n8759 , n8760 , n8761 , n8762 , n8763 , n8764 , n8765 , n8766 , n8767 , n8768 , n8769 , n8770 , n8771 , n8772 , n8773 , n8774 , n8775 , n8776 , n8777 , n8778 , n8779 , n8780 , n8781 , n8782 , n8783 , n8784 , n8785 , n8786 , n8787 , n8788 , n8789 , n8790 , n8791 , n8792 , n8793 , n8794 , n8795 , n8796 , n8797 , n8798 , n8799 , n8800 , n8801 , n8802 , n8803 , n8804 , n8805 , n8806 , n8807 , n8808 , n8809 , n8810 , n8811 , n8812 , n8813 , n8814 , n8815 , n8816 , n8817 , n8818 , n8819 , n8820 , n8821 , n8822 , n8823 , n8824 , n8825 , n8826 , n8827 , n8828 , n8829 , n8830 , n8831 , n8832 , n8833 , n8834 , n8835 , n8836 , n8837 , n8838 , n8839 , n8840 , n8841 , n8842 , n8843 , n8844 , n8845 , n8846 , n8847 , n8848 , n8849 , n8850 , n8851 , n8852 , n8853 , n8854 , n8855 , n8856 , n8857 , n8858 , n8859 , n8860 , n8861 , n8862 , n8863 , n8864 , n8865 , n8866 , n8867 , n8868 , n8869 , n8870 , n8871 , n8872 , n8873 , n8874 , n8875 , n8876 , n8877 , n8878 , n8879 , n8880 , n8881 , n8882 , n8883 , n8884 , n8885 , n8886 , n8887 , n8888 , n8889 , n8890 , n8891 , n8892 , n8893 , n8894 , n8895 , n8896 , n8897 , n8898 , n8899 , n8900 , n8901 , n8902 , n8903 , n8904 , n8905 , n8906 , n8907 , n8908 , n8909 , n8910 , n8911 , n8912 , n8913 , n8914 , n8915 , n8916 , n8917 , n8918 , n8919 , n8920 , n8921 , n8922 , n8923 , n8924 , n8925 , n8926 , n8927 , n8928 , n8929 , n8930 , n8931 , n8932 , n8933 , n8934 , n8935 , n8936 , n8937 , n8938 , n8939 , n8940 , n8941 , n8942 , n8943 , n8944 , n8945 , n8946 , n8947 , n8948 , n8949 , n8950 , n8951 , n8952 , n8953 , n8954 , n8955 , n8956 , n8957 , n8958 , n8959 , n8960 , n8961 , n8962 , n8963 , n8964 , n8965 , n8966 , n8967 , n8968 , n8969 , n8970 , n8971 , n8972 , n8973 , n8974 , n8975 , n8976 , n8977 , n8978 , n8979 , n8980 , n8981 , n8982 , n8983 , n8984 , n8985 , n8986 , n8987 , n8988 , n8989 , n8990 , n8991 , n8992 , n8993 , n8994 , n8995 , n8996 , n8997 , n8998 , n8999 , n9000 , n9001 , n9002 , n9003 , n9004 , n9005 , n9006 , n9007 , n9008 , n9009 , n9010 , n9011 , n9012 , n9013 , n9014 , n9015 , n9016 , n9017 , n9018 , n9019 , n9020 , n9021 , n9022 , n9023 , n9024 , n9025 , n9026 , n9027 , n9028 , n9029 , n9030 , n9031 , n9032 , n9033 , n9034 , n9035 , n9036 , n9037 , n9038 , n9039 , n9040 , n9041 , n9042 , n9043 , n9044 , n9045 , n9046 , n9047 , n9048 , n9049 , n9050 , n9051 , n9052 , n9053 , n9054 , n9055 , n9056 , n9057 , n9058 , n9059 , n9060 , n9061 , n9062 , n9063 , n9064 , n9065 , n9066 , n9067 , n9068 , n9069 , n9070 , n9071 , n9072 , n9073 , n9074 , n9075 , n9076 , n9077 , n9078 , n9079 , n9080 , n9081 , n9082 , n9083 , n9084 , n9085 , n9086 , n9087 , n9088 , n9089 , n9090 , n9091 , n9092 , n9093 , n9094 , n9095 , n9096 , n9097 , n9098 , n9099 , n9100 , n9101 , n9102 , n9103 , n9104 , n9105 , n9106 , n9107 , n9108 , n9109 , n9110 , n9111 , n9112 , n9113 , n9114 , n9115 , n9116 , n9117 , n9118 , n9119 , n9120 , n9121 , n9122 , n9123 , n9124 , n9125 , n9126 , n9127 , n9128 , n9129 , n9130 , n9131 , n9132 , n9133 , n9134 , n9135 , n9136 , n9137 , n9138 , n9139 , n9140 , n9141 , n9142 , n9143 , n9144 , n9145 , n9146 , n9147 , n9148 , n9149 , n9150 , n9151 , n9152 , n9153 , n9154 , n9155 , n9156 , n9157 , n9158 , n9159 , n9160 , n9161 , n9162 , n9163 , n9164 , n9165 , n9166 , n9167 , n9168 , n9169 , n9170 , n9171 , n9172 , n9173 , n9174 , n9175 , n9176 , n9177 , n9178 , n9179 , n9180 , n9181 , n9182 , n9183 , n9184 , n9185 , n9186 , n9187 , n9188 , n9189 , n9190 , n9191 , n9192 , n9193 , n9194 , n9195 , n9196 , n9197 , n9198 , n9199 , n9200 , n9201 , n9202 , n9203 , n9204 , n9205 , n9206 , n9207 , n9208 , n9209 , n9210 , n9211 , n9212 , n9213 , n9214 , n9215 , n9216 , n9217 , n9218 , n9219 , n9220 , n9221 , n9222 , n9223 , n9224 , n9225 , n9226 , n9227 , n9228 , n9229 , n9230 , n9231 , n9232 , n9233 , n9234 , n9235 , n9236 , n9237 , n9238 , n9239 , n9240 , n9241 , n9242 , n9243 , n9244 , n9245 , n9246 , n9247 , n9248 , n9249 , n9250 , n9251 , n9252 , n9253 , n9254 , n9255 , n9256 , n9257 , n9258 , n9259 , n9260 , n9261 , n9262 , n9263 , n9264 , n9265 , n9266 , n9267 , n9268 , n9269 , n9270 , n9271 , n9272 , n9273 , n9274 , n9275 , n9276 , n9277 , n9278 , n9279 , n9280 , n9281 , n9282 , n9283 , n9284 , n9285 , n9286 , n9287 , n9288 , n9289 , n9290 , n9291 , n9292 , n9293 , n9294 , n9295 , n9296 , n9297 , n9298 , n9299 , n9300 , n9301 , n9302 , n9303 , n9304 , n9305 , n9306 , n9307 , n9308 , n9309 , n9310 , n9311 , n9312 , n9313 , n9314 , n9315 , n9316 , n9317 , n9318 , n9319 , n9320 , n9321 , n9322 , n9323 , n9324 , n9325 , n9326 , n9327 , n9328 , n9329 , n9330 , n9331 , n9332 , n9333 , n9334 , n9335 , n9336 , n9337 , n9338 , n9339 , n9340 , n9341 , n9342 , n9343 , n9344 , n9345 , n9346 , n9347 , n9348 , n9349 , n9350 , n9351 , n9352 , n9353 , n9354 , n9355 , n9356 , n9357 , n9358 , n9359 , n9360 , n9361 , n9362 , n9363 , n9364 , n9365 , n9366 , n9367 , n9368 , n9369 , n9370 , n9371 , n9372 , n9373 , n9374 , n9375 , n9376 , n9377 , n9378 , n9379 , n9380 , n9381 , n9382 , n9383 , n9384 , n9385 , n9386 , n9387 , n9388 , n9389 , n9390 , n9391 , n9392 , n9393 , n9394 , n9395 , n9396 , n9397 , n9398 , n9399 , n9400 , n9401 , n9402 , n9403 , n9404 , n9405 , n9406 , n9407 , n9408 , n9409 , n9410 , n9411 , n9412 , n9413 , n9414 , n9415 , n9416 , n9417 , n9418 , n9419 , n9420 , n9421 , n9422 , n9423 , n9424 , n9425 , n9426 , n9427 , n9428 , n9429 , n9430 , n9431 , n9432 , n9433 , n9434 , n9435 , n9436 , n9437 , n9438 , n9439 , n9440 , n9441 , n9442 , n9443 , n9444 , n9445 , n9446 , n9447 , n9448 , n9449 , n9450 , n9451 , n9452 , n9453 , n9454 , n9455 , n9456 , n9457 , n9458 , n9459 , n9460 , n9461 , n9462 , n9463 , n9464 , n9465 , n9466 , n9467 , n9468 , n9469 , n9470 , n9471 , n9472 , n9473 , n9474 , n9475 , n9476 , n9477 , n9478 , n9479 , n9480 , n9481 , n9482 , n9483 , n9484 , n9485 , n9486 , n9487 , n9488 , n9489 , n9490 , n9491 , n9492 , n9493 , n9494 , n9495 , n9496 , n9497 , n9498 , n9499 , n9500 , n9501 , n9502 , n9503 , n9504 , n9505 , n9506 , n9507 , n9508 , n9509 , n9510 , n9511 , n9512 , n9513 , n9514 , n9515 , n9516 , n9517 , n9518 , n9519 , n9520 , n9521 , n9522 , n9523 , n9524 , n9525 , n9526 , n9527 , n9528 , n9529 , n9530 , n9531 , n9532 , n9533 , n9534 , n9535 , n9536 , n9537 , n9538 , n9539 , n9540 , n9541 , n9542 , n9543 , n9544 , n9545 , n9546 , n9547 , n9548 , n9549 , n9550 , n9551 , n9552 , n9553 , n9554 , n9555 , n9556 , n9557 , n9558 , n9559 , n9560 , n9561 , n9562 , n9563 , n9564 , n9565 , n9566 , n9567 , n9568 , n9569 , n9570 , n9571 , n9572 , n9573 , n9574 , n9575 , n9576 , n9577 , n9578 , n9579 , n9580 , n9581 , n9582 , n9583 , n9584 , n9585 , n9586 , n9587 , n9588 , n9589 , n9590 , n9591 , n9592 , n9593 , n9594 , n9595 , n9596 , n9597 , n9598 , n9599 , n9600 , n9601 , n9602 , n9603 , n9604 , n9605 , n9606 , n9607 , n9608 , n9609 , n9610 , n9611 , n9612 , n9613 , n9614 , n9615 , n9616 , n9617 , n9618 , n9619 , n9620 , n9621 , n9622 , n9623 , n9624 , n9625 , n9626 , n9627 , n9628 , n9629 , n9630 , n9631 , n9632 , n9633 , n9634 , n9635 , n9636 , n9637 , n9638 , n9639 , n9640 , n9641 , n9642 , n9643 , n9644 , n9645 , n9646 , n9647 , n9648 , n9649 , n9650 , n9651 , n9652 , n9653 , n9654 , n9655 , n9656 , n9657 , n9658 , n9659 , n9660 , n9661 , n9662 , n9663 , n9664 , n9665 , n9666 , n9667 , n9668 , n9669 , n9670 , n9671 , n9672 , n9673 , n9674 , n9675 , n9676 , n9677 , n9678 , n9679 , n9680 , n9681 , n9682 , n9683 , n9684 , n9685 , n9686 , n9687 , n9688 , n9689 , n9690 , n9691 , n9692 , n9693 , n9694 , n9695 , n9696 , n9697 , n9698 , n9699 , n9700 , n9701 , n9702 , n9703 , n9704 , n9705 , n9706 , n9707 , n9708 , n9709 , n9710 , n9711 , n9712 , n9713 , n9714 , n9715 , n9716 , n9717 , n9718 , n9719 , n9720 , n9721 , n9722 , n9723 , n9724 , n9725 , n9726 , n9727 , n9728 , n9729 , n9730 , n9731 , n9732 , n9733 , n9734 , n9735 , n9736 , n9737 , n9738 , n9739 , n9740 , n9741 , n9742 , n9743 , n9744 , n9745 , n9746 , n9747 , n9748 , n9749 , n9750 , n9751 , n9752 , n9753 , n9754 , n9755 , n9756 , n9757 , n9758 , n9759 , n9760 , n9761 , n9762 , n9763 , n9764 , n9765 , n9766 , n9767 , n9768 , n9769 , n9770 , n9771 , n9772 , n9773 , n9774 , n9775 , n9776 , n9777 , n9778 , n9779 , n9780 , n9781 , n9782 , n9783 , n9784 , n9785 , n9786 , n9787 , n9788 , n9789 , n9790 , n9791 , n9792 , n9793 , n9794 , n9795 , n9796 , n9797 , n9798 , n9799 , n9800 , n9801 , n9802 , n9803 , n9804 , n9805 , n9806 , n9807 , n9808 , n9809 , n9810 , n9811 , n9812 , n9813 , n9814 , n9815 , n9816 , n9817 , n9818 , n9819 , n9820 , n9821 , n9822 , n9823 , n9824 , n9825 , n9826 , n9827 , n9828 , n9829 , n9830 , n9831 , n9832 , n9833 , n9834 , n9835 , n9836 , n9837 , n9838 , n9839 , n9840 , n9841 , n9842 , n9843 , n9844 , n9845 , n9846 , n9847 , n9848 , n9849 , n9850 , n9851 , n9852 , n9853 , n9854 , n9855 , n9856 , n9857 , n9858 , n9859 , n9860 , n9861 , n9862 , n9863 , n9864 , n9865 , n9866 , n9867 , n9868 , n9869 , n9870 , n9871 , n9872 , n9873 , n9874 , n9875 , n9876 , n9877 , n9878 , n9879 , n9880 , n9881 , n9882 , n9883 , n9884 , n9885 , n9886 , n9887 , n9888 , n9889 , n9890 , n9891 , n9892 , n9893 , n9894 , n9895 , n9896 , n9897 , n9898 , n9899 , n9900 , n9901 , n9902 , n9903 , n9904 , n9905 , n9906 , n9907 , n9908 , n9909 , n9910 , n9911 , n9912 , n9913 , n9914 , n9915 , n9916 , n9917 , n9918 , n9919 , n9920 , n9921 , n9922 , n9923 , n9924 , n9925 , n9926 , n9927 , n9928 , n9929 , n9930 , n9931 , n9932 , n9933 , n9934 , n9935 , n9936 , n9937 , n9938 , n9939 , n9940 , n9941 , n9942 , n9943 , n9944 , n9945 , n9946 , n9947 , n9948 , n9949 , n9950 , n9951 , n9952 , n9953 , n9954 , n9955 , n9956 , n9957 , n9958 , n9959 , n9960 , n9961 , n9962 , n9963 , n9964 , n9965 , n9966 , n9967 , n9968 , n9969 , n9970 , n9971 , n9972 , n9973 , n9974 , n9975 , n9976 , n9977 , n9978 , n9979 , n9980 , n9981 , n9982 , n9983 , n9984 , n9985 , n9986 , n9987 , n9988 , n9989 , n9990 , n9991 , n9992 , n9993 , n9994 , n9995 , n9996 , n9997 , n9998 , n9999 , n10000 , n10001 , n10002 , n10003 , n10004 , n10005 , n10006 , n10007 , n10008 , n10009 , n10010 , n10011 , n10012 , n10013 , n10014 , n10015 , n10016 , n10017 , n10018 , n10019 , n10020 , n10021 , n10022 , n10023 , n10024 , n10025 , n10026 , n10027 , n10028 , n10029 , n10030 , n10031 , n10032 , n10033 , n10034 , n10035 , n10036 , n10037 , n10038 , n10039 , n10040 , n10041 , n10042 , n10043 , n10044 , n10045 , n10046 , n10047 , n10048 , n10049 , n10050 , n10051 , n10052 , n10053 , n10054 , n10055 , n10056 , n10057 , n10058 , n10059 , n10060 , n10061 , n10062 , n10063 , n10064 , n10065 , n10066 , n10067 , n10068 , n10069 , n10070 , n10071 , n10072 , n10073 , n10074 , n10075 , n10076 , n10077 , n10078 , n10079 , n10080 , n10081 , n10082 , n10083 , n10084 , n10085 , n10086 , n10087 , n10088 , n10089 , n10090 , n10091 , n10092 , n10093 , n10094 , n10095 , n10096 , n10097 , n10098 , n10099 , n10100 , n10101 , n10102 , n10103 , n10104 , n10105 , n10106 , n10107 , n10108 , n10109 , n10110 , n10111 , n10112 , n10113 , n10114 , n10115 , n10116 , n10117 , n10118 , n10119 , n10120 , n10121 , n10122 , n10123 , n10124 , n10125 , n10126 , n10127 , n10128 , n10129 , n10130 , n10131 , n10132 , n10133 , n10134 , n10135 , n10136 , n10137 , n10138 , n10139 , n10140 , n10141 , n10142 , n10143 , n10144 , n10145 , n10146 , n10147 , n10148 , n10149 , n10150 , n10151 , n10152 , n10153 , n10154 , n10155 , n10156 , n10157 , n10158 , n10159 , n10160 , n10161 , n10162 , n10163 , n10164 , n10165 , n10166 , n10167 , n10168 , n10169 , n10170 , n10171 , n10172 , n10173 , n10174 , n10175 , n10176 , n10177 , n10178 , n10179 , n10180 , n10181 , n10182 , n10183 , n10184 , n10185 , n10186 , n10187 , n10188 , n10189 , n10190 , n10191 , n10192 , n10193 , n10194 , n10195 , n10196 , n10197 , n10198 , n10199 , n10200 , n10201 , n10202 , n10203 , n10204 , n10205 , n10206 , n10207 , n10208 , n10209 , n10210 , n10211 , n10212 , n10213 , n10214 , n10215 , n10216 , n10217 , n10218 , n10219 , n10220 , n10221 , n10222 , n10223 , n10224 , n10225 , n10226 , n10227 , n10228 , n10229 , n10230 , n10231 , n10232 , n10233 , n10234 , n10235 , n10236 , n10237 , n10238 , n10239 , n10240 , n10241 , n10242 , n10243 , n10244 , n10245 , n10246 , n10247 , n10248 , n10249 , n10250 , n10251 , n10252 , n10253 , n10254 , n10255 , n10256 , n10257 , n10258 , n10259 , n10260 , n10261 , n10262 , n10263 , n10264 , n10265 , n10266 , n10267 , n10268 , n10269 , n10270 , n10271 , n10272 , n10273 , n10274 , n10275 , n10276 , n10277 , n10278 , n10279 , n10280 , n10281 , n10282 , n10283 , n10284 , n10285 , n10286 , n10287 , n10288 , n10289 , n10290 , n10291 , n10292 , n10293 , n10294 , n10295 , n10296 , n10297 , n10298 , n10299 , n10300 , n10301 , n10302 , n10303 , n10304 , n10305 , n10306 , n10307 , n10308 , n10309 , n10310 , n10311 , n10312 , n10313 , n10314 , n10315 , n10316 , n10317 , n10318 , n10319 , n10320 , n10321 , n10322 , n10323 , n10324 , n10325 , n10326 , n10327 , n10328 , n10329 , n10330 , n10331 , n10332 , n10333 , n10334 , n10335 , n10336 , n10337 , n10338 , n10339 , n10340 , n10341 , n10342 , n10343 , n10344 , n10345 , n10346 , n10347 , n10348 , n10349 , n10350 , n10351 , n10352 , n10353 , n10354 , n10355 , n10356 , n10357 , n10358 , n10359 , n10360 , n10361 , n10362 , n10363 , n10364 , n10365 , n10366 , n10367 , n10368 , n10369 , n10370 , n10371 , n10372 , n10373 , n10374 , n10375 , n10376 , n10377 , n10378 , n10379 , n10380 , n10381 , n10382 , n10383 , n10384 , n10385 , n10386 , n10387 , n10388 , n10389 , n10390 , n10391 , n10392 , n10393 , n10394 , n10395 , n10396 , n10397 , n10398 , n10399 , n10400 , n10401 , n10402 , n10403 , n10404 , n10405 , n10406 , n10407 , n10408 , n10409 , n10410 , n10411 , n10412 , n10413 , n10414 , n10415 , n10416 , n10417 , n10418 , n10419 , n10420 , n10421 , n10422 , n10423 , n10424 , n10425 , n10426 , n10427 , n10428 , n10429 , n10430 , n10431 , n10432 , n10433 , n10434 , n10435 , n10436 , n10437 , n10438 , n10439 , n10440 , n10441 , n10442 , n10443 , n10444 , n10445 , n10446 , n10447 , n10448 , n10449 , n10450 , n10451 , n10452 , n10453 , n10454 , n10455 , n10456 , n10457 , n10458 , n10459 , n10460 , n10461 , n10462 , n10463 , n10464 , n10465 , n10466 , n10467 , n10468 , n10469 , n10470 , n10471 , n10472 , n10473 , n10474 , n10475 , n10476 , n10477 , n10478 , n10479 , n10480 , n10481 , n10482 , n10483 , n10484 , n10485 , n10486 , n10487 , n10488 , n10489 , n10490 , n10491 , n10492 , n10493 , n10494 , n10495 , n10496 , n10497 , n10498 , n10499 , n10500 , n10501 , n10502 , n10503 , n10504 , n10505 , n10506 , n10507 , n10508 , n10509 , n10510 , n10511 , n10512 , n10513 , n10514 , n10515 , n10516 , n10517 , n10518 , n10519 , n10520 , n10521 , n10522 , n10523 , n10524 , n10525 , n10526 , n10527 , n10528 , n10529 , n10530 , n10531 , n10532 , n10533 , n10534 , n10535 , n10536 , n10537 , n10538 , n10539 , n10540 , n10541 , n10542 , n10543 , n10544 , n10545 , n10546 , n10547 , n10548 , n10549 , n10550 , n10551 , n10552 , n10553 , n10554 , n10555 , n10556 , n10557 , n10558 , n10559 , n10560 , n10561 , n10562 , n10563 , n10564 , n10565 , n10566 , n10567 , n10568 , n10569 , n10570 , n10571 , n10572 , n10573 , n10574 , n10575 , n10576 , n10577 , n10578 , n10579 , n10580 , n10581 , n10582 , n10583 , n10584 , n10585 , n10586 , n10587 , n10588 , n10589 , n10590 , n10591 , n10592 , n10593 , n10594 , n10595 , n10596 , n10597 , n10598 , n10599 , n10600 , n10601 , n10602 , n10603 , n10604 , n10605 , n10606 , n10607 , n10608 , n10609 , n10610 , n10611 , n10612 , n10613 , n10614 , n10615 , n10616 , n10617 , n10618 , n10619 , n10620 , n10621 , n10622 , n10623 , n10624 , n10625 , n10626 , n10627 , n10628 , n10629 , n10630 , n10631 , n10632 , n10633 , n10634 , n10635 , n10636 , n10637 , n10638 , n10639 , n10640 , n10641 , n10642 , n10643 , n10644 , n10645 , n10646 , n10647 , n10648 , n10649 , n10650 , n10651 , n10652 , n10653 , n10654 , n10655 , n10656 , n10657 , n10658 , n10659 , n10660 , n10661 , n10662 , n10663 , n10664 , n10665 , n10666 , n10667 , n10668 , n10669 , n10670 , n10671 , n10672 , n10673 , n10674 , n10675 , n10676 , n10677 , n10678 , n10679 , n10680 , n10681 , n10682 , n10683 , n10684 , n10685 , n10686 , n10687 , n10688 , n10689 , n10690 , n10691 , n10692 , n10693 , n10694 , n10695 , n10696 , n10697 , n10698 , n10699 , n10700 , n10701 , n10702 , n10703 , n10704 , n10705 , n10706 , n10707 , n10708 , n10709 , n10710 , n10711 , n10712 , n10713 , n10714 , n10715 , n10716 , n10717 , n10718 , n10719 , n10720 , n10721 , n10722 , n10723 , n10724 , n10725 , n10726 , n10727 , n10728 , n10729 , n10730 , n10731 , n10732 , n10733 , n10734 , n10735 , n10736 , n10737 , n10738 , n10739 , n10740 , n10741 , n10742 , n10743 , n10744 , n10745 , n10746 , n10747 , n10748 , n10749 , n10750 , n10751 , n10752 , n10753 , n10754 , n10755 , n10756 , n10757 , n10758 , n10759 , n10760 , n10761 , n10762 , n10763 , n10764 , n10765 , n10766 , n10767 , n10768 , n10769 , n10770 , n10771 , n10772 , n10773 , n10774 , n10775 , n10776 , n10777 , n10778 , n10779 , n10780 , n10781 , n10782 , n10783 , n10784 , n10785 , n10786 , n10787 , n10788 , n10789 , n10790 , n10791 , n10792 , n10793 , n10794 , n10795 , n10796 , n10797 , n10798 , n10799 , n10800 , n10801 , n10802 , n10803 , n10804 , n10805 , n10806 , n10807 , n10808 , n10809 , n10810 , n10811 , n10812 , n10813 , n10814 , n10815 , n10816 , n10817 , n10818 , n10819 , n10820 , n10821 , n10822 , n10823 , n10824 , n10825 , n10826 , n10827 , n10828 , n10829 , n10830 , n10831 , n10832 , n10833 , n10834 , n10835 , n10836 , n10837 , n10838 , n10839 , n10840 , n10841 , n10842 , n10843 , n10844 , n10845 , n10846 , n10847 , n10848 , n10849 , n10850 , n10851 , n10852 , n10853 , n10854 , n10855 , n10856 , n10857 , n10858 , n10859 , n10860 , n10861 , n10862 , n10863 , n10864 , n10865 , n10866 , n10867 , n10868 , n10869 , n10870 , n10871 , n10872 , n10873 , n10874 , n10875 , n10876 , n10877 , n10878 , n10879 , n10880 , n10881 , n10882 , n10883 , n10884 , n10885 , n10886 , n10887 , n10888 , n10889 , n10890 , n10891 , n10892 , n10893 , n10894 , n10895 , n10896 , n10897 , n10898 , n10899 , n10900 , n10901 , n10902 , n10903 , n10904 , n10905 , n10906 , n10907 , n10908 , n10909 , n10910 , n10911 , n10912 , n10913 , n10914 , n10915 , n10916 , n10917 , n10918 , n10919 , n10920 , n10921 , n10922 , n10923 , n10924 , n10925 , n10926 , n10927 , n10928 , n10929 , n10930 , n10931 , n10932 , n10933 , n10934 , n10935 , n10936 , n10937 , n10938 , n10939 , n10940 , n10941 , n10942 , n10943 , n10944 , n10945 , n10946 , n10947 , n10948 , n10949 , n10950 , n10951 , n10952 , n10953 , n10954 , n10955 , n10956 , n10957 , n10958 , n10959 , n10960 , n10961 , n10962 , n10963 , n10964 , n10965 , n10966 , n10967 , n10968 , n10969 , n10970 , n10971 , n10972 , n10973 , n10974 , n10975 , n10976 , n10977 , n10978 , n10979 , n10980 , n10981 , n10982 , n10983 , n10984 , n10985 , n10986 , n10987 , n10988 , n10989 , n10990 , n10991 , n10992 , n10993 , n10994 , n10995 , n10996 , n10997 , n10998 , n10999 , n11000 , n11001 , n11002 , n11003 , n11004 , n11005 , n11006 , n11007 , n11008 , n11009 , n11010 , n11011 , n11012 , n11013 , n11014 , n11015 , n11016 , n11017 , n11018 , n11019 , n11020 , n11021 , n11022 , n11023 , n11024 , n11025 , n11026 , n11027 , n11028 , n11029 , n11030 , n11031 , n11032 , n11033 , n11034 , n11035 , n11036 , n11037 , n11038 , n11039 , n11040 , n11041 , n11042 , n11043 , n11044 , n11045 , n11046 , n11047 , n11048 , n11049 , n11050 , n11051 , n11052 , n11053 , n11054 , n11055 , n11056 , n11057 , n11058 , n11059 , n11060 , n11061 , n11062 , n11063 , n11064 , n11065 , n11066 , n11067 , n11068 , n11069 , n11070 , n11071 , n11072 , n11073 , n11074 , n11075 , n11076 , n11077 , n11078 , n11079 , n11080 , n11081 , n11082 , n11083 , n11084 , n11085 , n11086 , n11087 , n11088 , n11089 , n11090 , n11091 , n11092 , n11093 , n11094 , n11095 , n11096 , n11097 , n11098 , n11099 , n11100 , n11101 , n11102 , n11103 , n11104 , n11105 , n11106 , n11107 , n11108 , n11109 , n11110 , n11111 , n11112 , n11113 , n11114 , n11115 , n11116 , n11117 , n11118 , n11119 , n11120 , n11121 , n11122 , n11123 , n11124 , n11125 , n11126 , n11127 , n11128 , n11129 , n11130 , n11131 , n11132 , n11133 , n11134 , n11135 , n11136 , n11137 , n11138 , n11139 , n11140 , n11141 , n11142 , n11143 , n11144 , n11145 , n11146 , n11147 , n11148 , n11149 , n11150 , n11151 , n11152 , n11153 , n11154 , n11155 , n11156 , n11157 , n11158 , n11159 , n11160 , n11161 , n11162 , n11163 , n11164 , n11165 , n11166 , n11167 , n11168 , n11169 , n11170 , n11171 , n11172 , n11173 , n11174 , n11175 , n11176 , n11177 , n11178 , n11179 , n11180 , n11181 , n11182 , n11183 , n11184 , n11185 , n11186 , n11187 , n11188 , n11189 , n11190 , n11191 , n11192 , n11193 , n11194 , n11195 , n11196 , n11197 , n11198 , n11199 , n11200 , n11201 , n11202 , n11203 , n11204 , n11205 , n11206 , n11207 , n11208 , n11209 , n11210 , n11211 , n11212 , n11213 , n11214 , n11215 , n11216 , n11217 , n11218 , n11219 , n11220 , n11221 , n11222 , n11223 , n11224 , n11225 , n11226 , n11227 , n11228 , n11229 , n11230 , n11231 , n11232 , n11233 , n11234 , n11235 , n11236 , n11237 , n11238 , n11239 , n11240 , n11241 , n11242 , n11243 , n11244 , n11245 , n11246 , n11247 , n11248 , n11249 , n11250 , n11251 , n11252 , n11253 , n11254 , n11255 , n11256 , n11257 , n11258 , n11259 , n11260 , n11261 , n11262 , n11263 , n11264 , n11265 , n11266 , n11267 , n11268 , n11269 , n11270 , n11271 , n11272 , n11273 , n11274 , n11275 , n11276 , n11277 , n11278 , n11279 , n11280 , n11281 , n11282 , n11283 , n11284 , n11285 , n11286 , n11287 , n11288 , n11289 , n11290 , n11291 , n11292 , n11293 , n11294 , n11295 , n11296 , n11297 , n11298 , n11299 , n11300 , n11301 , n11302 , n11303 , n11304 , n11305 , n11306 , n11307 , n11308 , n11309 , n11310 , n11311 , n11312 , n11313 , n11314 , n11315 , n11316 , n11317 , n11318 , n11319 , n11320 , n11321 , n11322 , n11323 , n11324 , n11325 , n11326 , n11327 , n11328 , n11329 , n11330 , n11331 , n11332 , n11333 , n11334 , n11335 , n11336 , n11337 , n11338 , n11339 , n11340 , n11341 , n11342 , n11343 , n11344 , n11345 , n11346 , n11347 , n11348 , n11349 , n11350 , n11351 , n11352 , n11353 , n11354 , n11355 , n11356 , n11357 , n11358 , n11359 , n11360 , n11361 , n11362 , n11363 , n11364 , n11365 , n11366 , n11367 , n11368 , n11369 , n11370 , n11371 , n11372 , n11373 , n11374 , n11375 , n11376 , n11377 , n11378 , n11379 , n11380 , n11381 , n11382 , n11383 , n11384 , n11385 , n11386 , n11387 , n11388 , n11389 , n11390 , n11391 , n11392 , n11393 , n11394 , n11395 , n11396 , n11397 , n11398 , n11399 , n11400 , n11401 , n11402 , n11403 , n11404 , n11405 , n11406 , n11407 , n11408 , n11409 , n11410 , n11411 , n11412 , n11413 , n11414 , n11415 , n11416 , n11417 , n11418 , n11419 , n11420 , n11421 , n11422 , n11423 , n11424 , n11425 , n11426 , n11427 , n11428 , n11429 , n11430 , n11431 , n11432 , n11433 , n11434 , n11435 , n11436 , n11437 , n11438 , n11439 , n11440 , n11441 , n11442 , n11443 , n11444 , n11445 , n11446 , n11447 , n11448 , n11449 , n11450 , n11451 , n11452 , n11453 , n11454 , n11455 , n11456 , n11457 , n11458 , n11459 , n11460 , n11461 , n11462 , n11463 , n11464 , n11465 , n11466 , n11467 , n11468 , n11469 , n11470 , n11471 , n11472 , n11473 , n11474 , n11475 , n11476 , n11477 , n11478 , n11479 , n11480 , n11481 , n11482 , n11483 , n11484 , n11485 , n11486 , n11487 , n11488 , n11489 , n11490 , n11491 , n11492 , n11493 , n11494 , n11495 , n11496 , n11497 , n11498 , n11499 , n11500 , n11501 , n11502 , n11503 , n11504 , n11505 , n11506 , n11507 , n11508 , n11509 , n11510 , n11511 , n11512 , n11513 , n11514 , n11515 , n11516 , n11517 , n11518 , n11519 , n11520 , n11521 , n11522 , n11523 , n11524 , n11525 , n11526 , n11527 , n11528 , n11529 , n11530 , n11531 , n11532 , n11533 , n11534 , n11535 , n11536 , n11537 , n11538 , n11539 , n11540 , n11541 , n11542 , n11543 , n11544 , n11545 , n11546 , n11547 , n11548 , n11549 , n11550 , n11551 , n11552 , n11553 , n11554 , n11555 , n11556 , n11557 , n11558 , n11559 , n11560 , n11561 , n11562 , n11563 , n11564 , n11565 , n11566 , n11567 , n11568 , n11569 , n11570 , n11571 , n11572 , n11573 , n11574 , n11575 , n11576 , n11577 , n11578 , n11579 , n11580 , n11581 , n11582 , n11583 , n11584 , n11585 , n11586 , n11587 , n11588 , n11589 , n11590 , n11591 , n11592 , n11593 , n11594 , n11595 , n11596 , n11597 , n11598 , n11599 , n11600 , n11601 , n11602 , n11603 , n11604 , n11605 , n11606 , n11607 , n11608 , n11609 , n11610 , n11611 , n11612 , n11613 , n11614 , n11615 , n11616 , n11617 , n11618 , n11619 , n11620 , n11621 , n11622 , n11623 , n11624 , n11625 , n11626 , n11627 , n11628 , n11629 , n11630 , n11631 , n11632 , n11633 , n11634 , n11635 , n11636 , n11637 , n11638 , n11639 , n11640 , n11641 , n11642 , n11643 , n11644 , n11645 , n11646 , n11647 , n11648 , n11649 , n11650 , n11651 , n11652 , n11653 , n11654 , n11655 , n11656 , n11657 , n11658 , n11659 , n11660 , n11661 , n11662 , n11663 , n11664 , n11665 , n11666 , n11667 , n11668 , n11669 , n11670 , n11671 , n11672 , n11673 , n11674 , n11675 , n11676 , n11677 , n11678 , n11679 , n11680 , n11681 , n11682 , n11683 , n11684 , n11685 , n11686 , n11687 , n11688 , n11689 , n11690 , n11691 , n11692 , n11693 , n11694 , n11695 , n11696 , n11697 , n11698 , n11699 , n11700 , n11701 , n11702 , n11703 , n11704 , n11705 , n11706 , n11707 , n11708 , n11709 , n11710 , n11711 , n11712 , n11713 , n11714 , n11715 , n11716 , n11717 , n11718 , n11719 , n11720 , n11721 , n11722 , n11723 , n11724 , n11725 , n11726 , n11727 , n11728 , n11729 , n11730 , n11731 , n11732 , n11733 , n11734 , n11735 , n11736 , n11737 , n11738 , n11739 , n11740 , n11741 , n11742 , n11743 , n11744 , n11745 , n11746 , n11747 , n11748 , n11749 , n11750 , n11751 , n11752 , n11753 , n11754 , n11755 , n11756 , n11757 , n11758 , n11759 , n11760 , n11761 , n11762 , n11763 , n11764 , n11765 , n11766 , n11767 , n11768 , n11769 , n11770 , n11771 , n11772 , n11773 , n11774 , n11775 , n11776 , n11777 , n11778 , n11779 , n11780 , n11781 , n11782 , n11783 , n11784 , n11785 , n11786 , n11787 , n11788 , n11789 , n11790 , n11791 , n11792 , n11793 , n11794 , n11795 , n11796 , n11797 , n11798 , n11799 , n11800 , n11801 , n11802 , n11803 , n11804 , n11805 , n11806 , n11807 , n11808 , n11809 , n11810 , n11811 , n11812 , n11813 , n11814 , n11815 , n11816 , n11817 , n11818 , n11819 , n11820 , n11821 , n11822 , n11823 , n11824 , n11825 , n11826 , n11827 , n11828 , n11829 , n11830 , n11831 , n11832 , n11833 , n11834 , n11835 , n11836 , n11837 , n11838 , n11839 , n11840 , n11841 , n11842 , n11843 , n11844 , n11845 , n11846 , n11847 , n11848 , n11849 , n11850 , n11851 , n11852 , n11853 , n11854 , n11855 , n11856 , n11857 , n11858 , n11859 , n11860 , n11861 , n11862 , n11863 , n11864 , n11865 , n11866 , n11867 , n11868 , n11869 , n11870 , n11871 , n11872 , n11873 , n11874 , n11875 , n11876 , n11877 , n11878 , n11879 , n11880 , n11881 , n11882 , n11883 , n11884 , n11885 , n11886 , n11887 , n11888 , n11889 , n11890 , n11891 , n11892 , n11893 , n11894 , n11895 , n11896 , n11897 , n11898 , n11899 , n11900 , n11901 , n11902 , n11903 , n11904 , n11905 , n11906 , n11907 , n11908 , n11909 , n11910 , n11911 , n11912 , n11913 , n11914 , n11915 , n11916 , n11917 , n11918 , n11919 , n11920 , n11921 , n11922 , n11923 , n11924 , n11925 , n11926 , n11927 , n11928 , n11929 , n11930 , n11931 , n11932 , n11933 , n11934 , n11935 , n11936 , n11937 , n11938 , n11939 , n11940 , n11941 , n11942 , n11943 , n11944 , n11945 , n11946 , n11947 , n11948 , n11949 , n11950 , n11951 , n11952 , n11953 , n11954 , n11955 , n11956 , n11957 , n11958 , n11959 , n11960 , n11961 , n11962 , n11963 , n11964 , n11965 , n11966 , n11967 , n11968 , n11969 , n11970 , n11971 , n11972 , n11973 , n11974 , n11975 , n11976 , n11977 , n11978 , n11979 , n11980 , n11981 , n11982 , n11983 , n11984 , n11985 , n11986 , n11987 , n11988 , n11989 , n11990 , n11991 , n11992 , n11993 , n11994 , n11995 , n11996 , n11997 , n11998 , n11999 , n12000 , n12001 , n12002 , n12003 , n12004 , n12005 , n12006 , n12007 , n12008 , n12009 , n12010 , n12011 , n12012 , n12013 , n12014 , n12015 , n12016 , n12017 , n12018 , n12019 , n12020 , n12021 , n12022 , n12023 , n12024 , n12025 , n12026 , n12027 , n12028 , n12029 , n12030 , n12031 , n12032 , n12033 , n12034 , n12035 , n12036 , n12037 , n12038 , n12039 , n12040 , n12041 , n12042 , n12043 , n12044 , n12045 , n12046 , n12047 , n12048 , n12049 , n12050 , n12051 , n12052 , n12053 , n12054 , n12055 , n12056 , n12057 , n12058 , n12059 , n12060 , n12061 , n12062 , n12063 , n12064 , n12065 , n12066 , n12067 , n12068 , n12069 , n12070 , n12071 , n12072 , n12073 , n12074 , n12075 , n12076 , n12077 , n12078 , n12079 , n12080 , n12081 , n12082 , n12083 , n12084 , n12085 , n12086 , n12087 , n12088 , n12089 , n12090 , n12091 , n12092 , n12093 , n12094 , n12095 , n12096 , n12097 , n12098 , n12099 , n12100 , n12101 , n12102 , n12103 , n12104 , n12105 , n12106 , n12107 , n12108 , n12109 , n12110 , n12111 , n12112 , n12113 , n12114 , n12115 , n12116 , n12117 , n12118 , n12119 , n12120 , n12121 , n12122 , n12123 , n12124 , n12125 , n12126 , n12127 , n12128 , n12129 , n12130 , n12131 , n12132 , n12133 , n12134 , n12135 , n12136 , n12137 , n12138 , n12139 , n12140 , n12141 , n12142 , n12143 , n12144 , n12145 , n12146 , n12147 , n12148 , n12149 , n12150 , n12151 , n12152 , n12153 , n12154 , n12155 , n12156 , n12157 , n12158 , n12159 , n12160 , n12161 , n12162 , n12163 , n12164 , n12165 , n12166 , n12167 , n12168 , n12169 , n12170 , n12171 , n12172 , n12173 , n12174 , n12175 , n12176 , n12177 , n12178 , n12179 , n12180 , n12181 , n12182 , n12183 , n12184 , n12185 , n12186 , n12187 , n12188 , n12189 , n12190 , n12191 , n12192 , n12193 , n12194 , n12195 , n12196 , n12197 , n12198 , n12199 , n12200 , n12201 , n12202 , n12203 , n12204 , n12205 , n12206 , n12207 , n12208 , n12209 , n12210 , n12211 , n12212 , n12213 , n12214 , n12215 , n12216 , n12217 , n12218 , n12219 , n12220 , n12221 , n12222 , n12223 , n12224 , n12225 , n12226 , n12227 , n12228 , n12229 , n12230 , n12231 , n12232 , n12233 , n12234 , n12235 , n12236 , n12237 , n12238 , n12239 , n12240 , n12241 , n12242 , n12243 , n12244 , n12245 , n12246 , n12247 , n12248 , n12249 , n12250 , n12251 , n12252 , n12253 , n12254 , n12255 , n12256 , n12257 , n12258 , n12259 , n12260 , n12261 , n12262 , n12263 , n12264 , n12265 , n12266 , n12267 , n12268 , n12269 , n12270 , n12271 , n12272 , n12273 , n12274 , n12275 , n12276 , n12277 , n12278 , n12279 , n12280 , n12281 , n12282 , n12283 , n12284 , n12285 , n12286 , n12287 , n12288 , n12289 , n12290 , n12291 , n12292 , n12293 , n12294 , n12295 , n12296 , n12297 , n12298 , n12299 , n12300 , n12301 , n12302 , n12303 , n12304 , n12305 , n12306 , n12307 , n12308 , n12309 , n12310 , n12311 , n12312 , n12313 , n12314 , n12315 , n12316 , n12317 , n12318 , n12319 , n12320 , n12321 , n12322 , n12323 , n12324 , n12325 , n12326 , n12327 , n12328 , n12329 , n12330 , n12331 , n12332 , n12333 , n12334 , n12335 , n12336 , n12337 , n12338 , n12339 , n12340 , n12341 , n12342 , n12343 , n12344 , n12345 , n12346 , n12347 , n12348 , n12349 , n12350 , n12351 , n12352 , n12353 , n12354 , n12355 , n12356 , n12357 , n12358 , n12359 , n12360 , n12361 , n12362 , n12363 , n12364 , n12365 , n12366 , n12367 , n12368 , n12369 , n12370 , n12371 , n12372 , n12373 , n12374 , n12375 , n12376 , n12377 , n12378 , n12379 , n12380 , n12381 , n12382 , n12383 , n12384 , n12385 , n12386 , n12387 , n12388 , n12389 , n12390 , n12391 , n12392 , n12393 , n12394 , n12395 , n12396 , n12397 , n12398 , n12399 , n12400 , n12401 , n12402 , n12403 , n12404 , n12405 , n12406 , n12407 , n12408 , n12409 , n12410 , n12411 , n12412 , n12413 , n12414 , n12415 , n12416 , n12417 , n12418 , n12419 , n12420 , n12421 , n12422 , n12423 , n12424 , n12425 , n12426 , n12427 , n12428 , n12429 , n12430 , n12431 , n12432 , n12433 , n12434 , n12435 , n12436 , n12437 , n12438 , n12439 , n12440 , n12441 , n12442 , n12443 , n12444 , n12445 , n12446 , n12447 , n12448 , n12449 , n12450 , n12451 , n12452 , n12453 , n12454 , n12455 , n12456 , n12457 , n12458 , n12459 , n12460 , n12461 , n12462 , n12463 , n12464 , n12465 , n12466 , n12467 , n12468 , n12469 , n12470 , n12471 , n12472 , n12473 , n12474 , n12475 , n12476 , n12477 , n12478 , n12479 , n12480 , n12481 , n12482 , n12483 , n12484 , n12485 , n12486 , n12487 , n12488 , n12489 , n12490 , n12491 , n12492 , n12493 , n12494 , n12495 , n12496 , n12497 , n12498 , n12499 , n12500 , n12501 , n12502 , n12503 , n12504 , n12505 , n12506 , n12507 , n12508 , n12509 , n12510 , n12511 , n12512 , n12513 , n12514 , n12515 , n12516 , n12517 , n12518 , n12519 , n12520 , n12521 , n12522 , n12523 , n12524 , n12525 , n12526 , n12527 , n12528 , n12529 , n12530 , n12531 , n12532 , n12533 , n12534 , n12535 , n12536 , n12537 , n12538 , n12539 , n12540 , n12541 , n12542 , n12543 , n12544 , n12545 , n12546 , n12547 , n12548 , n12549 , n12550 , n12551 , n12552 , n12553 , n12554 , n12555 , n12556 , n12557 , n12558 , n12559 , n12560 , n12561 , n12562 , n12563 , n12564 , n12565 , n12566 , n12567 , n12568 , n12569 , n12570 , n12571 , n12572 , n12573 , n12574 , n12575 , n12576 , n12577 , n12578 , n12579 , n12580 , n12581 , n12582 , n12583 , n12584 , n12585 , n12586 , n12587 , n12588 , n12589 , n12590 , n12591 , n12592 , n12593 , n12594 , n12595 , n12596 , n12597 , n12598 , n12599 , n12600 , n12601 , n12602 , n12603 , n12604 , n12605 , n12606 , n12607 , n12608 , n12609 , n12610 , n12611 , n12612 , n12613 , n12614 , n12615 , n12616 , n12617 , n12618 , n12619 , n12620 , n12621 , n12622 , n12623 , n12624 , n12625 , n12626 , n12627 , n12628 , n12629 , n12630 , n12631 , n12632 , n12633 , n12634 , n12635 , n12636 , n12637 , n12638 , n12639 , n12640 , n12641 , n12642 , n12643 , n12644 , n12645 , n12646 , n12647 , n12648 , n12649 , n12650 , n12651 , n12652 , n12653 , n12654 , n12655 , n12656 , n12657 , n12658 , n12659 , n12660 , n12661 , n12662 , n12663 , n12664 , n12665 , n12666 , n12667 , n12668 , n12669 , n12670 , n12671 , n12672 , n12673 , n12674 , n12675 , n12676 , n12677 , n12678 , n12679 , n12680 , n12681 , n12682 , n12683 , n12684 , n12685 , n12686 , n12687 , n12688 , n12689 , n12690 , n12691 , n12692 , n12693 , n12694 , n12695 , n12696 , n12697 , n12698 , n12699 , n12700 , n12701 , n12702 , n12703 , n12704 , n12705 , n12706 , n12707 , n12708 , n12709 , n12710 , n12711 , n12712 , n12713 , n12714 , n12715 , n12716 , n12717 , n12718 , n12719 , n12720 , n12721 , n12722 , n12723 , n12724 , n12725 , n12726 , n12727 , n12728 , n12729 , n12730 , n12731 , n12732 , n12733 , n12734 , n12735 , n12736 , n12737 , n12738 , n12739 , n12740 , n12741 , n12742 , n12743 , n12744 , n12745 , n12746 , n12747 , n12748 , n12749 , n12750 , n12751 , n12752 , n12753 , n12754 , n12755 , n12756 , n12757 , n12758 , n12759 , n12760 , n12761 , n12762 , n12763 , n12764 , n12765 , n12766 , n12767 , n12768 , n12769 , n12770 , n12771 , n12772 , n12773 , n12774 , n12775 , n12776 , n12777 , n12778 , n12779 , n12780 , n12781 , n12782 , n12783 , n12784 , n12785 , n12786 , n12787 , n12788 , n12789 , n12790 , n12791 , n12792 , n12793 , n12794 , n12795 , n12796 , n12797 , n12798 , n12799 , n12800 , n12801 , n12802 , n12803 , n12804 , n12805 , n12806 , n12807 , n12808 , n12809 , n12810 , n12811 , n12812 , n12813 , n12814 , n12815 , n12816 , n12817 , n12818 , n12819 , n12820 , n12821 , n12822 , n12823 , n12824 , n12825 , n12826 , n12827 , n12828 , n12829 , n12830 , n12831 , n12832 , n12833 , n12834 , n12835 , n12836 , n12837 , n12838 , n12839 , n12840 , n12841 , n12842 , n12843 , n12844 , n12845 , n12846 , n12847 , n12848 , n12849 , n12850 , n12851 , n12852 , n12853 , n12854 , n12855 , n12856 , n12857 , n12858 , n12859 , n12860 , n12861 , n12862 , n12863 , n12864 , n12865 , n12866 , n12867 , n12868 , n12869 , n12870 , n12871 , n12872 , n12873 , n12874 , n12875 , n12876 , n12877 , n12878 , n12879 , n12880 , n12881 , n12882 , n12883 , n12884 , n12885 , n12886 , n12887 , n12888 , n12889 , n12890 , n12891 , n12892 , n12893 , n12894 , n12895 , n12896 , n12897 , n12898 , n12899 , n12900 , n12901 , n12902 , n12903 , n12904 , n12905 , n12906 , n12907 , n12908 , n12909 , n12910 , n12911 , n12912 , n12913 , n12914 , n12915 , n12916 , n12917 , n12918 , n12919 , n12920 , n12921 , n12922 , n12923 , n12924 , n12925 , n12926 , n12927 , n12928 , n12929 , n12930 , n12931 , n12932 , n12933 , n12934 , n12935 , n12936 , n12937 , n12938 , n12939 , n12940 , n12941 , n12942 , n12943 , n12944 , n12945 , n12946 , n12947 , n12948 , n12949 , n12950 , n12951 , n12952 , n12953 , n12954 , n12955 , n12956 , n12957 , n12958 , n12959 , n12960 , n12961 , n12962 , n12963 , n12964 , n12965 , n12966 , n12967 , n12968 , n12969 , n12970 , n12971 , n12972 , n12973 , n12974 , n12975 , n12976 , n12977 , n12978 , n12979 , n12980 , n12981 , n12982 , n12983 , n12984 , n12985 , n12986 , n12987 , n12988 , n12989 , n12990 , n12991 , n12992 , n12993 , n12994 , n12995 , n12996 , n12997 , n12998 , n12999 , n13000 , n13001 , n13002 , n13003 , n13004 , n13005 , n13006 , n13007 , n13008 , n13009 , n13010 , n13011 , n13012 , n13013 , n13014 , n13015 , n13016 , n13017 , n13018 , n13019 , n13020 , n13021 , n13022 , n13023 , n13024 , n13025 , n13026 , n13027 , n13028 , n13029 , n13030 , n13031 , n13032 , n13033 , n13034 , n13035 , n13036 , n13037 , n13038 , n13039 , n13040 , n13041 , n13042 , n13043 , n13044 , n13045 , n13046 , n13047 , n13048 , n13049 , n13050 , n13051 , n13052 , n13053 , n13054 , n13055 , n13056 , n13057 , n13058 , n13059 , n13060 , n13061 , n13062 , n13063 , n13064 , n13065 , n13066 , n13067 , n13068 , n13069 , n13070 , n13071 , n13072 , n13073 , n13074 , n13075 , n13076 , n13077 , n13078 , n13079 , n13080 , n13081 , n13082 , n13083 , n13084 , n13085 , n13086 , n13087 , n13088 , n13089 , n13090 , n13091 , n13092 , n13093 , n13094 , n13095 , n13096 , n13097 , n13098 , n13099 , n13100 , n13101 , n13102 , n13103 , n13104 , n13105 , n13106 , n13107 , n13108 , n13109 , n13110 , n13111 , n13112 , n13113 , n13114 , n13115 , n13116 , n13117 , n13118 , n13119 , n13120 , n13121 , n13122 , n13123 , n13124 , n13125 , n13126 , n13127 , n13128 , n13129 , n13130 , n13131 , n13132 , n13133 , n13134 , n13135 , n13136 , n13137 , n13138 , n13139 , n13140 , n13141 , n13142 , n13143 , n13144 , n13145 , n13146 , n13147 , n13148 , n13149 , n13150 , n13151 , n13152 , n13153 , n13154 , n13155 , n13156 , n13157 , n13158 , n13159 , n13160 , n13161 , n13162 , n13163 , n13164 , n13165 , n13166 , n13167 , n13168 , n13169 , n13170 , n13171 , n13172 , n13173 , n13174 , n13175 , n13176 , n13177 , n13178 , n13179 , n13180 , n13181 , n13182 , n13183 , n13184 , n13185 , n13186 , n13187 , n13188 , n13189 , n13190 , n13191 , n13192 , n13193 , n13194 , n13195 , n13196 , n13197 , n13198 , n13199 , n13200 , n13201 , n13202 , n13203 , n13204 , n13205 , n13206 , n13207 , n13208 , n13209 , n13210 , n13211 , n13212 , n13213 , n13214 , n13215 , n13216 , n13217 , n13218 , n13219 , n13220 , n13221 , n13222 , n13223 , n13224 , n13225 , n13226 , n13227 , n13228 , n13229 , n13230 , n13231 , n13232 , n13233 , n13234 , n13235 , n13236 , n13237 , n13238 , n13239 , n13240 , n13241 , n13242 , n13243 , n13244 , n13245 , n13246 , n13247 , n13248 , n13249 , n13250 , n13251 , n13252 , n13253 , n13254 , n13255 , n13256 , n13257 , n13258 , n13259 , n13260 , n13261 , n13262 , n13263 , n13264 , n13265 , n13266 , n13267 , n13268 , n13269 , n13270 , n13271 , n13272 , n13273 , n13274 , n13275 , n13276 , n13277 , n13278 , n13279 , n13280 , n13281 , n13282 , n13283 , n13284 , n13285 , n13286 , n13287 , n13288 , n13289 , n13290 , n13291 , n13292 , n13293 , n13294 , n13295 , n13296 , n13297 , n13298 , n13299 , n13300 , n13301 , n13302 , n13303 , n13304 , n13305 , n13306 , n13307 , n13308 , n13309 , n13310 , n13311 , n13312 , n13313 , n13314 , n13315 , n13316 , n13317 , n13318 , n13319 , n13320 , n13321 , n13322 , n13323 , n13324 , n13325 , n13326 , n13327 , n13328 , n13329 , n13330 , n13331 , n13332 , n13333 , n13334 , n13335 , n13336 , n13337 , n13338 , n13339 , n13340 , n13341 , n13342 , n13343 , n13344 , n13345 , n13346 , n13347 , n13348 , n13349 , n13350 , n13351 , n13352 , n13353 , n13354 , n13355 , n13356 , n13357 , n13358 , n13359 , n13360 , n13361 , n13362 , n13363 , n13364 , n13365 , n13366 , n13367 , n13368 , n13369 , n13370 , n13371 , n13372 , n13373 , n13374 , n13375 , n13376 , n13377 , n13378 , n13379 , n13380 , n13381 , n13382 , n13383 , n13384 , n13385 , n13386 , n13387 , n13388 , n13389 , n13390 , n13391 , n13392 , n13393 , n13394 , n13395 , n13396 , n13397 , n13398 , n13399 , n13400 , n13401 , n13402 , n13403 , n13404 , n13405 , n13406 , n13407 , n13408 , n13409 , n13410 , n13411 , n13412 , n13413 , n13414 , n13415 , n13416 , n13417 , n13418 , n13419 , n13420 , n13421 , n13422 , n13423 , n13424 , n13425 , n13426 , n13427 , n13428 , n13429 , n13430 , n13431 , n13432 , n13433 , n13434 , n13435 , n13436 , n13437 , n13438 , n13439 , n13440 , n13441 , n13442 , n13443 , n13444 , n13445 , n13446 , n13447 , n13448 , n13449 , n13450 , n13451 , n13452 , n13453 , n13454 , n13455 , n13456 , n13457 , n13458 , n13459 , n13460 , n13461 , n13462 , n13463 , n13464 , n13465 , n13466 , n13467 , n13468 , n13469 , n13470 , n13471 , n13472 , n13473 , n13474 , n13475 , n13476 , n13477 , n13478 , n13479 , n13480 , n13481 , n13482 , n13483 , n13484 , n13485 , n13486 , n13487 , n13488 , n13489 , n13490 , n13491 , n13492 , n13493 , n13494 , n13495 , n13496 , n13497 , n13498 , n13499 , n13500 , n13501 , n13502 , n13503 , n13504 , n13505 , n13506 , n13507 , n13508 , n13509 , n13510 , n13511 , n13512 , n13513 , n13514 , n13515 , n13516 , n13517 , n13518 , n13519 , n13520 , n13521 , n13522 , n13523 , n13524 , n13525 , n13526 , n13527 , n13528 , n13529 , n13530 , n13531 , n13532 , n13533 , n13534 , n13535 , n13536 , n13537 , n13538 , n13539 , n13540 , n13541 , n13542 , n13543 , n13544 , n13545 , n13546 , n13547 , n13548 , n13549 , n13550 , n13551 , n13552 , n13553 , n13554 , n13555 , n13556 , n13557 , n13558 , n13559 , n13560 , n13561 , n13562 , n13563 , n13564 , n13565 , n13566 , n13567 , n13568 , n13569 , n13570 , n13571 , n13572 , n13573 , n13574 , n13575 , n13576 , n13577 , n13578 , n13579 , n13580 , n13581 , n13582 , n13583 , n13584 , n13585 , n13586 , n13587 , n13588 , n13589 , n13590 , n13591 , n13592 , n13593 , n13594 , n13595 , n13596 , n13597 , n13598 , n13599 , n13600 , n13601 , n13602 , n13603 , n13604 , n13605 , n13606 , n13607 , n13608 , n13609 , n13610 , n13611 , n13612 , n13613 , n13614 , n13615 , n13616 , n13617 , n13618 , n13619 , n13620 , n13621 , n13622 , n13623 , n13624 , n13625 , n13626 , n13627 , n13628 , n13629 , n13630 , n13631 , n13632 , n13633 , n13634 , n13635 , n13636 , n13637 , n13638 , n13639 , n13640 , n13641 , n13642 , n13643 , n13644 , n13645 , n13646 , n13647 , n13648 , n13649 , n13650 , n13651 , n13652 , n13653 , n13654 , n13655 , n13656 , n13657 , n13658 , n13659 , n13660 , n13661 , n13662 , n13663 , n13664 , n13665 , n13666 , n13667 , n13668 , n13669 , n13670 , n13671 , n13672 , n13673 , n13674 , n13675 , n13676 , n13677 , n13678 , n13679 , n13680 , n13681 , n13682 , n13683 , n13684 , n13685 , n13686 , n13687 , n13688 , n13689 , n13690 , n13691 , n13692 , n13693 , n13694 , n13695 , n13696 , n13697 , n13698 , n13699 , n13700 , n13701 , n13702 , n13703 , n13704 , n13705 , n13706 , n13707 , n13708 , n13709 , n13710 , n13711 , n13712 , n13713 , n13714 , n13715 , n13716 , n13717 , n13718 , n13719 , n13720 , n13721 , n13722 , n13723 , n13724 , n13725 , n13726 , n13727 , n13728 , n13729 , n13730 , n13731 , n13732 , n13733 , n13734 , n13735 , n13736 , n13737 , n13738 , n13739 , n13740 , n13741 , n13742 , n13743 , n13744 , n13745 , n13746 , n13747 , n13748 , n13749 , n13750 , n13751 , n13752 , n13753 , n13754 , n13755 , n13756 , n13757 , n13758 , n13759 , n13760 , n13761 , n13762 , n13763 , n13764 , n13765 , n13766 , n13767 , n13768 , n13769 , n13770 , n13771 , n13772 , n13773 , n13774 , n13775 , n13776 , n13777 , n13778 , n13779 , n13780 , n13781 , n13782 , n13783 , n13784 , n13785 , n13786 , n13787 , n13788 , n13789 , n13790 , n13791 , n13792 , n13793 , n13794 , n13795 , n13796 , n13797 , n13798 , n13799 , n13800 , n13801 , n13802 , n13803 , n13804 , n13805 , n13806 , n13807 , n13808 , n13809 , n13810 , n13811 , n13812 , n13813 , n13814 , n13815 , n13816 , n13817 , n13818 , n13819 , n13820 , n13821 , n13822 , n13823 , n13824 , n13825 , n13826 , n13827 , n13828 , n13829 , n13830 , n13831 , n13832 , n13833 , n13834 , n13835 , n13836 , n13837 , n13838 , n13839 , n13840 , n13841 , n13842 , n13843 , n13844 , n13845 , n13846 , n13847 , n13848 , n13849 , n13850 , n13851 , n13852 , n13853 , n13854 , n13855 , n13856 , n13857 , n13858 , n13859 , n13860 , n13861 , n13862 , n13863 , n13864 , n13865 , n13866 , n13867 , n13868 , n13869 , n13870 , n13871 , n13872 , n13873 , n13874 , n13875 , n13876 , n13877 , n13878 , n13879 , n13880 , n13881 , n13882 , n13883 , n13884 , n13885 , n13886 , n13887 , n13888 , n13889 , n13890 , n13891 , n13892 , n13893 , n13894 , n13895 , n13896 , n13897 , n13898 , n13899 , n13900 , n13901 , n13902 , n13903 , n13904 , n13905 , n13906 , n13907 , n13908 , n13909 , n13910 , n13911 , n13912 , n13913 , n13914 , n13915 , n13916 , n13917 , n13918 , n13919 , n13920 , n13921 , n13922 , n13923 , n13924 , n13925 , n13926 , n13927 , n13928 , n13929 , n13930 , n13931 , n13932 , n13933 , n13934 , n13935 , n13936 , n13937 , n13938 , n13939 , n13940 , n13941 , n13942 , n13943 , n13944 , n13945 , n13946 , n13947 , n13948 , n13949 , n13950 , n13951 , n13952 , n13953 , n13954 , n13955 , n13956 , n13957 , n13958 , n13959 , n13960 , n13961 , n13962 , n13963 , n13964 , n13965 , n13966 , n13967 , n13968 , n13969 , n13970 , n13971 , n13972 , n13973 , n13974 , n13975 , n13976 , n13977 , n13978 , n13979 , n13980 , n13981 , n13982 , n13983 , n13984 , n13985 , n13986 , n13987 , n13988 , n13989 , n13990 , n13991 , n13992 , n13993 , n13994 , n13995 , n13996 , n13997 , n13998 , n13999 , n14000 , n14001 , n14002 , n14003 , n14004 , n14005 , n14006 , n14007 , n14008 , n14009 , n14010 , n14011 , n14012 , n14013 , n14014 , n14015 , n14016 , n14017 , n14018 , n14019 , n14020 , n14021 , n14022 , n14023 , n14024 , n14025 , n14026 , n14027 , n14028 , n14029 , n14030 , n14031 , n14032 , n14033 , n14034 , n14035 , n14036 , n14037 , n14038 , n14039 , n14040 , n14041 , n14042 , n14043 , n14044 , n14045 , n14046 , n14047 , n14048 , n14049 , n14050 , n14051 , n14052 , n14053 , n14054 , n14055 , n14056 , n14057 , n14058 , n14059 , n14060 , n14061 , n14062 , n14063 , n14064 , n14065 , n14066 , n14067 , n14068 , n14069 , n14070 , n14071 , n14072 , n14073 , n14074 , n14075 , n14076 , n14077 , n14078 , n14079 , n14080 , n14081 , n14082 , n14083 , n14084 , n14085 , n14086 , n14087 , n14088 , n14089 , n14090 , n14091 , n14092 , n14093 , n14094 , n14095 , n14096 , n14097 , n14098 , n14099 , n14100 , n14101 , n14102 , n14103 , n14104 , n14105 , n14106 , n14107 , n14108 , n14109 , n14110 , n14111 , n14112 , n14113 , n14114 , n14115 , n14116 , n14117 , n14118 , n14119 , n14120 , n14121 , n14122 , n14123 , n14124 , n14125 , n14126 , n14127 , n14128 , n14129 , n14130 , n14131 , n14132 , n14133 , n14134 , n14135 , n14136 , n14137 , n14138 , n14139 , n14140 , n14141 , n14142 , n14143 , n14144 , n14145 , n14146 , n14147 , n14148 , n14149 , n14150 , n14151 , n14152 , n14153 , n14154 , n14155 , n14156 , n14157 , n14158 , n14159 , n14160 , n14161 , n14162 , n14163 , n14164 , n14165 , n14166 , n14167 , n14168 , n14169 , n14170 , n14171 , n14172 , n14173 , n14174 , n14175 , n14176 , n14177 , n14178 , n14179 , n14180 , n14181 , n14182 , n14183 , n14184 , n14185 , n14186 , n14187 , n14188 , n14189 , n14190 , n14191 , n14192 , n14193 , n14194 , n14195 , n14196 , n14197 , n14198 , n14199 , n14200 , n14201 , n14202 , n14203 , n14204 , n14205 , n14206 , n14207 , n14208 , n14209 , n14210 , n14211 , n14212 , n14213 , n14214 , n14215 , n14216 , n14217 , n14218 , n14219 , n14220 , n14221 , n14222 , n14223 , n14224 , n14225 , n14226 , n14227 , n14228 , n14229 , n14230 , n14231 , n14232 , n14233 , n14234 , n14235 , n14236 , n14237 , n14238 , n14239 , n14240 , n14241 , n14242 , n14243 , n14244 , n14245 , n14246 , n14247 , n14248 , n14249 , n14250 , n14251 , n14252 , n14253 , n14254 , n14255 , n14256 , n14257 , n14258 , n14259 , n14260 , n14261 , n14262 , n14263 , n14264 , n14265 , n14266 , n14267 , n14268 , n14269 , n14270 , n14271 , n14272 , n14273 , n14274 , n14275 , n14276 , n14277 , n14278 , n14279 , n14280 , n14281 , n14282 , n14283 , n14284 , n14285 , n14286 , n14287 , n14288 , n14289 , n14290 , n14291 , n14292 , n14293 , n14294 , n14295 , n14296 , n14297 , n14298 , n14299 , n14300 , n14301 , n14302 , n14303 , n14304 , n14305 , n14306 , n14307 , n14308 , n14309 , n14310 , n14311 , n14312 , n14313 , n14314 , n14315 , n14316 , n14317 , n14318 , n14319 , n14320 , n14321 , n14322 , n14323 , n14324 , n14325 , n14326 , n14327 , n14328 , n14329 , n14330 , n14331 , n14332 , n14333 , n14334 , n14335 , n14336 , n14337 , n14338 , n14339 , n14340 , n14341 , n14342 , n14343 , n14344 , n14345 , n14346 , n14347 , n14348 , n14349 , n14350 , n14351 , n14352 , n14353 , n14354 , n14355 , n14356 , n14357 , n14358 , n14359 , n14360 , n14361 , n14362 , n14363 , n14364 , n14365 , n14366 , n14367 , n14368 , n14369 , n14370 , n14371 , n14372 , n14373 , n14374 , n14375 , n14376 , n14377 , n14378 , n14379 , n14380 , n14381 , n14382 , n14383 , n14384 , n14385 , n14386 , n14387 , n14388 , n14389 , n14390 , n14391 , n14392 , n14393 , n14394 , n14395 , n14396 , n14397 , n14398 , n14399 , n14400 , n14401 , n14402 , n14403 , n14404 , n14405 , n14406 , n14407 , n14408 , n14409 , n14410 , n14411 , n14412 , n14413 , n14414 , n14415 , n14416 , n14417 , n14418 , n14419 , n14420 , n14421 , n14422 , n14423 , n14424 , n14425 , n14426 , n14427 , n14428 , n14429 , n14430 , n14431 , n14432 , n14433 , n14434 , n14435 , n14436 , n14437 , n14438 , n14439 , n14440 , n14441 , n14442 , n14443 , n14444 , n14445 , n14446 , n14447 , n14448 , n14449 , n14450 , n14451 , n14452 , n14453 , n14454 , n14455 , n14456 , n14457 , n14458 , n14459 , n14460 , n14461 , n14462 , n14463 , n14464 , n14465 , n14466 , n14467 , n14468 , n14469 , n14470 , n14471 , n14472 , n14473 , n14474 , n14475 , n14476 , n14477 , n14478 , n14479 , n14480 , n14481 , n14482 , n14483 , n14484 , n14485 , n14486 , n14487 , n14488 , n14489 , n14490 , n14491 , n14492 , n14493 , n14494 , n14495 , n14496 , n14497 , n14498 , n14499 , n14500 , n14501 , n14502 , n14503 , n14504 , n14505 , n14506 , n14507 , n14508 , n14509 , n14510 , n14511 , n14512 , n14513 , n14514 , n14515 , n14516 , n14517 , n14518 , n14519 , n14520 , n14521 , n14522 , n14523 , n14524 , n14525 , n14526 , n14527 , n14528 , n14529 , n14530 , n14531 , n14532 , n14533 , n14534 , n14535 , n14536 , n14537 , n14538 , n14539 , n14540 , n14541 , n14542 , n14543 , n14544 , n14545 , n14546 , n14547 , n14548 , n14549 , n14550 , n14551 , n14552 , n14553 , n14554 , n14555 , n14556 , n14557 , n14558 , n14559 , n14560 , n14561 , n14562 , n14563 , n14564 , n14565 , n14566 , n14567 , n14568 , n14569 , n14570 , n14571 , n14572 , n14573 , n14574 , n14575 , n14576 , n14577 , n14578 , n14579 , n14580 , n14581 , n14582 , n14583 , n14584 , n14585 , n14586 , n14587 , n14588 , n14589 , n14590 , n14591 , n14592 , n14593 , n14594 , n14595 , n14596 , n14597 , n14598 , n14599 , n14600 , n14601 , n14602 , n14603 , n14604 , n14605 , n14606 , n14607 , n14608 , n14609 , n14610 , n14611 , n14612 , n14613 , n14614 , n14615 , n14616 , n14617 , n14618 , n14619 , n14620 , n14621 , n14622 , n14623 , n14624 , n14625 , n14626 , n14627 , n14628 , n14629 , n14630 , n14631 , n14632 , n14633 , n14634 , n14635 , n14636 , n14637 , n14638 , n14639 , n14640 , n14641 , n14642 , n14643 , n14644 , n14645 , n14646 , n14647 , n14648 , n14649 , n14650 , n14651 , n14652 , n14653 , n14654 , n14655 , n14656 , n14657 , n14658 , n14659 , n14660 , n14661 , n14662 , n14663 , n14664 , n14665 , n14666 , n14667 , n14668 , n14669 , n14670 , n14671 , n14672 , n14673 , n14674 , n14675 , n14676 , n14677 , n14678 , n14679 , n14680 , n14681 , n14682 , n14683 , n14684 , n14685 , n14686 , n14687 , n14688 , n14689 , n14690 , n14691 , n14692 , n14693 , n14694 , n14695 , n14696 , n14697 , n14698 , n14699 , n14700 , n14701 , n14702 , n14703 , n14704 , n14705 , n14706 , n14707 , n14708 , n14709 , n14710 , n14711 , n14712 , n14713 , n14714 , n14715 , n14716 , n14717 , n14718 , n14719 , n14720 , n14721 , n14722 , n14723 , n14724 , n14725 , n14726 , n14727 , n14728 , n14729 , n14730 , n14731 , n14732 , n14733 , n14734 , n14735 , n14736 , n14737 , n14738 , n14739 , n14740 , n14741 , n14742 , n14743 , n14744 , n14745 , n14746 , n14747 , n14748 , n14749 , n14750 , n14751 , n14752 , n14753 , n14754 , n14755 , n14756 , n14757 , n14758 , n14759 , n14760 , n14761 , n14762 , n14763 , n14764 , n14765 , n14766 , n14767 , n14768 , n14769 , n14770 , n14771 , n14772 , n14773 , n14774 , n14775 , n14776 , n14777 , n14778 , n14779 , n14780 , n14781 , n14782 , n14783 , n14784 , n14785 , n14786 , n14787 , n14788 , n14789 , n14790 , n14791 , n14792 , n14793 , n14794 , n14795 , n14796 , n14797 , n14798 , n14799 , n14800 , n14801 , n14802 , n14803 , n14804 , n14805 , n14806 , n14807 , n14808 , n14809 , n14810 , n14811 , n14812 , n14813 , n14814 , n14815 , n14816 , n14817 , n14818 , n14819 , n14820 , n14821 , n14822 , n14823 , n14824 , n14825 , n14826 , n14827 , n14828 , n14829 , n14830 , n14831 , n14832 , n14833 , n14834 , n14835 , n14836 , n14837 , n14838 , n14839 , n14840 , n14841 , n14842 , n14843 , n14844 , n14845 , n14846 , n14847 , n14848 , n14849 , n14850 , n14851 , n14852 , n14853 , n14854 , n14855 , n14856 , n14857 , n14858 , n14859 , n14860 , n14861 , n14862 , n14863 , n14864 , n14865 , n14866 , n14867 , n14868 , n14869 , n14870 , n14871 , n14872 , n14873 , n14874 , n14875 , n14876 , n14877 , n14878 , n14879 , n14880 , n14881 , n14882 , n14883 , n14884 , n14885 , n14886 , n14887 , n14888 , n14889 , n14890 , n14891 , n14892 , n14893 , n14894 , n14895 , n14896 , n14897 , n14898 , n14899 , n14900 , n14901 , n14902 , n14903 , n14904 , n14905 , n14906 , n14907 , n14908 , n14909 , n14910 , n14911 , n14912 , n14913 , n14914 , n14915 , n14916 , n14917 , n14918 , n14919 , n14920 , n14921 , n14922 , n14923 , n14924 , n14925 , n14926 , n14927 , n14928 , n14929 , n14930 , n14931 , n14932 , n14933 , n14934 , n14935 , n14936 , n14937 , n14938 , n14939 , n14940 , n14941 , n14942 , n14943 , n14944 , n14945 , n14946 , n14947 , n14948 , n14949 , n14950 , n14951 , n14952 , n14953 , n14954 , n14955 , n14956 , n14957 , n14958 , n14959 , n14960 , n14961 , n14962 , n14963 , n14964 , n14965 , n14966 , n14967 , n14968 , n14969 , n14970 , n14971 , n14972 , n14973 , n14974 , n14975 , n14976 , n14977 , n14978 , n14979 , n14980 , n14981 , n14982 , n14983 , n14984 , n14985 , n14986 , n14987 , n14988 , n14989 , n14990 , n14991 , n14992 , n14993 , n14994 , n14995 , n14996 , n14997 , n14998 , n14999 , n15000 , n15001 , n15002 , n15003 , n15004 , n15005 , n15006 , n15007 , n15008 , n15009 , n15010 , n15011 , n15012 , n15013 , n15014 , n15015 , n15016 , n15017 , n15018 , n15019 , n15020 , n15021 , n15022 , n15023 , n15024 , n15025 , n15026 , n15027 , n15028 , n15029 , n15030 , n15031 , n15032 , n15033 , n15034 , n15035 , n15036 , n15037 , n15038 , n15039 , n15040 , n15041 , n15042 , n15043 , n15044 , n15045 , n15046 , n15047 , n15048 , n15049 , n15050 , n15051 , n15052 , n15053 , n15054 , n15055 , n15056 , n15057 , n15058 , n15059 , n15060 , n15061 , n15062 , n15063 , n15064 , n15065 , n15066 , n15067 , n15068 , n15069 , n15070 , n15071 , n15072 , n15073 , n15074 , n15075 , n15076 , n15077 , n15078 , n15079 , n15080 , n15081 , n15082 , n15083 , n15084 , n15085 , n15086 , n15087 , n15088 , n15089 , n15090 , n15091 , n15092 , n15093 , n15094 , n15095 , n15096 , n15097 , n15098 , n15099 , n15100 , n15101 , n15102 , n15103 , n15104 , n15105 , n15106 , n15107 , n15108 , n15109 , n15110 , n15111 , n15112 , n15113 , n15114 , n15115 , n15116 , n15117 , n15118 , n15119 , n15120 , n15121 , n15122 , n15123 , n15124 , n15125 , n15126 , n15127 , n15128 , n15129 , n15130 , n15131 , n15132 , n15133 , n15134 , n15135 , n15136 , n15137 , n15138 , n15139 , n15140 , n15141 , n15142 , n15143 , n15144 , n15145 , n15146 , n15147 , n15148 , n15149 , n15150 , n15151 , n15152 , n15153 , n15154 , n15155 , n15156 , n15157 , n15158 , n15159 , n15160 , n15161 , n15162 , n15163 , n15164 , n15165 , n15166 , n15167 , n15168 , n15169 , n15170 , n15171 , n15172 , n15173 , n15174 , n15175 , n15176 , n15177 , n15178 , n15179 , n15180 , n15181 , n15182 , n15183 , n15184 , n15185 , n15186 , n15187 , n15188 , n15189 , n15190 , n15191 , n15192 , n15193 , n15194 , n15195 , n15196 , n15197 , n15198 , n15199 , n15200 , n15201 , n15202 , n15203 , n15204 , n15205 , n15206 , n15207 , n15208 , n15209 , n15210 , n15211 , n15212 , n15213 , n15214 , n15215 , n15216 , n15217 , n15218 , n15219 , n15220 , n15221 , n15222 , n15223 , n15224 , n15225 , n15226 , n15227 , n15228 , n15229 , n15230 , n15231 , n15232 , n15233 , n15234 , n15235 , n15236 , n15237 , n15238 , n15239 , n15240 , n15241 , n15242 , n15243 , n15244 , n15245 , n15246 , n15247 , n15248 , n15249 , n15250 , n15251 , n15252 , n15253 , n15254 , n15255 , n15256 , n15257 , n15258 , n15259 , n15260 , n15261 , n15262 , n15263 , n15264 , n15265 , n15266 , n15267 , n15268 , n15269 , n15270 , n15271 , n15272 , n15273 , n15274 , n15275 , n15276 , n15277 , n15278 , n15279 , n15280 , n15281 , n15282 , n15283 , n15284 , n15285 , n15286 , n15287 , n15288 , n15289 , n15290 , n15291 , n15292 , n15293 , n15294 , n15295 , n15296 , n15297 , n15298 , n15299 , n15300 , n15301 , n15302 , n15303 , n15304 , n15305 , n15306 , n15307 , n15308 , n15309 , n15310 , n15311 , n15312 , n15313 , n15314 , n15315 , n15316 , n15317 , n15318 , n15319 , n15320 , n15321 , n15322 , n15323 , n15324 , n15325 , n15326 , n15327 , n15328 , n15329 , n15330 , n15331 , n15332 , n15333 , n15334 , n15335 , n15336 , n15337 , n15338 , n15339 , n15340 , n15341 , n15342 , n15343 , n15344 , n15345 , n15346 , n15347 , n15348 , n15349 , n15350 , n15351 , n15352 , n15353 , n15354 , n15355 , n15356 , n15357 , n15358 , n15359 , n15360 , n15361 , n15362 , n15363 , n15364 , n15365 , n15366 , n15367 , n15368 , n15369 , n15370 , n15371 , n15372 , n15373 , n15374 , n15375 , n15376 , n15377 , n15378 , n15379 , n15380 , n15381 , n15382 , n15383 , n15384 , n15385 , n15386 , n15387 , n15388 , n15389 , n15390 , n15391 , n15392 , n15393 , n15394 , n15395 , n15396 , n15397 , n15398 , n15399 , n15400 , n15401 , n15402 , n15403 , n15404 , n15405 , n15406 , n15407 , n15408 , n15409 , n15410 , n15411 , n15412 , n15413 , n15414 , n15415 , n15416 , n15417 , n15418 , n15419 , n15420 , n15421 , n15422 , n15423 , n15424 , n15425 , n15426 , n15427 , n15428 , n15429 , n15430 , n15431 , n15432 , n15433 , n15434 , n15435 , n15436 , n15437 , n15438 , n15439 , n15440 , n15441 , n15442 , n15443 , n15444 , n15445 , n15446 , n15447 , n15448 , n15449 , n15450 , n15451 , n15452 , n15453 , n15454 , n15455 , n15456 , n15457 , n15458 , n15459 , n15460 , n15461 , n15462 , n15463 , n15464 , n15465 , n15466 , n15467 , n15468 , n15469 , n15470 , n15471 , n15472 , n15473 , n15474 , n15475 , n15476 , n15477 , n15478 , n15479 , n15480 , n15481 , n15482 , n15483 , n15484 , n15485 , n15486 , n15487 , n15488 , n15489 , n15490 , n15491 , n15492 , n15493 , n15494 , n15495 , n15496 , n15497 , n15498 , n15499 , n15500 , n15501 , n15502 , n15503 , n15504 , n15505 , n15506 , n15507 , n15508 , n15509 , n15510 , n15511 , n15512 , n15513 , n15514 , n15515 , n15516 , n15517 , n15518 , n15519 , n15520 , n15521 , n15522 , n15523 , n15524 , n15525 , n15526 , n15527 , n15528 , n15529 , n15530 , n15531 , n15532 , n15533 , n15534 , n15535 , n15536 , n15537 , n15538 , n15539 , n15540 , n15541 , n15542 , n15543 , n15544 , n15545 , n15546 , n15547 , n15548 , n15549 , n15550 , n15551 , n15552 , n15553 , n15554 , n15555 , n15556 , n15557 , n15558 , n15559 , n15560 , n15561 , n15562 , n15563 , n15564 , n15565 , n15566 , n15567 , n15568 , n15569 , n15570 , n15571 , n15572 , n15573 , n15574 , n15575 , n15576 , n15577 , n15578 , n15579 , n15580 , n15581 , n15582 , n15583 , n15584 , n15585 , n15586 , n15587 , n15588 , n15589 , n15590 , n15591 , n15592 , n15593 , n15594 , n15595 , n15596 , n15597 , n15598 , n15599 , n15600 , n15601 , n15602 , n15603 , n15604 , n15605 , n15606 , n15607 , n15608 , n15609 , n15610 , n15611 , n15612 , n15613 , n15614 , n15615 , n15616 , n15617 , n15618 , n15619 , n15620 , n15621 , n15622 , n15623 , n15624 , n15625 , n15626 , n15627 , n15628 , n15629 , n15630 , n15631 , n15632 , n15633 , n15634 , n15635 , n15636 , n15637 , n15638 , n15639 , n15640 , n15641 , n15642 , n15643 , n15644 , n15645 , n15646 , n15647 , n15648 , n15649 , n15650 , n15651 , n15652 , n15653 , n15654 , n15655 , n15656 , n15657 , n15658 , n15659 , n15660 , n15661 , n15662 , n15663 , n15664 , n15665 , n15666 , n15667 , n15668 , n15669 , n15670 , n15671 , n15672 , n15673 , n15674 , n15675 , n15676 , n15677 , n15678 , n15679 , n15680 , n15681 , n15682 , n15683 , n15684 , n15685 , n15686 , n15687 , n15688 , n15689 , n15690 , n15691 , n15692 , n15693 , n15694 , n15695 , n15696 , n15697 , n15698 , n15699 , n15700 , n15701 , n15702 , n15703 , n15704 , n15705 , n15706 , n15707 , n15708 , n15709 , n15710 , n15711 , n15712 , n15713 , n15714 , n15715 , n15716 , n15717 , n15718 , n15719 , n15720 , n15721 , n15722 , n15723 , n15724 , n15725 , n15726 , n15727 , n15728 , n15729 , n15730 , n15731 , n15732 , n15733 , n15734 , n15735 , n15736 , n15737 , n15738 , n15739 , n15740 , n15741 , n15742 , n15743 , n15744 , n15745 , n15746 , n15747 , n15748 , n15749 , n15750 , n15751 , n15752 , n15753 , n15754 , n15755 , n15756 , n15757 , n15758 , n15759 , n15760 , n15761 , n15762 , n15763 , n15764 , n15765 , n15766 , n15767 , n15768 , n15769 , n15770 , n15771 , n15772 , n15773 , n15774 , n15775 , n15776 , n15777 , n15778 , n15779 , n15780 , n15781 , n15782 , n15783 , n15784 , n15785 , n15786 , n15787 , n15788 , n15789 , n15790 , n15791 , n15792 , n15793 , n15794 , n15795 , n15796 , n15797 , n15798 , n15799 , n15800 , n15801 , n15802 , n15803 , n15804 , n15805 , n15806 , n15807 , n15808 , n15809 , n15810 , n15811 , n15812 , n15813 , n15814 , n15815 , n15816 , n15817 , n15818 , n15819 , n15820 , n15821 , n15822 , n15823 , n15824 , n15825 , n15826 , n15827 , n15828 , n15829 , n15830 , n15831 , n15832 , n15833 , n15834 , n15835 , n15836 , n15837 , n15838 , n15839 , n15840 , n15841 , n15842 , n15843 , n15844 , n15845 , n15846 , n15847 , n15848 , n15849 , n15850 , n15851 , n15852 , n15853 , n15854 , n15855 , n15856 , n15857 , n15858 , n15859 , n15860 , n15861 , n15862 , n15863 , n15864 , n15865 , n15866 , n15867 , n15868 , n15869 , n15870 , n15871 , n15872 , n15873 , n15874 , n15875 , n15876 , n15877 , n15878 , n15879 , n15880 , n15881 , n15882 , n15883 , n15884 , n15885 , n15886 , n15887 , n15888 , n15889 , n15890 , n15891 , n15892 , n15893 , n15894 , n15895 , n15896 , n15897 , n15898 , n15899 , n15900 , n15901 , n15902 , n15903 , n15904 , n15905 , n15906 , n15907 , n15908 , n15909 , n15910 , n15911 , n15912 , n15913 , n15914 , n15915 , n15916 , n15917 , n15918 , n15919 , n15920 , n15921 , n15922 , n15923 , n15924 , n15925 , n15926 , n15927 , n15928 , n15929 , n15930 , n15931 , n15932 , n15933 , n15934 , n15935 , n15936 , n15937 , n15938 , n15939 , n15940 , n15941 , n15942 , n15943 , n15944 , n15945 , n15946 , n15947 , n15948 , n15949 , n15950 , n15951 , n15952 , n15953 , n15954 , n15955 , n15956 , n15957 , n15958 , n15959 , n15960 , n15961 , n15962 , n15963 , n15964 , n15965 , n15966 , n15967 , n15968 , n15969 , n15970 , n15971 , n15972 , n15973 , n15974 , n15975 , n15976 , n15977 , n15978 , n15979 , n15980 , n15981 , n15982 , n15983 , n15984 , n15985 , n15986 , n15987 , n15988 , n15989 , n15990 , n15991 , n15992 , n15993 , n15994 , n15995 , n15996 , n15997 , n15998 , n15999 , n16000 , n16001 , n16002 , n16003 , n16004 , n16005 , n16006 , n16007 , n16008 , n16009 , n16010 , n16011 , n16012 , n16013 , n16014 , n16015 , n16016 , n16017 , n16018 , n16019 , n16020 , n16021 , n16022 , n16023 , n16024 , n16025 , n16026 , n16027 , n16028 , n16029 , n16030 , n16031 , n16032 , n16033 , n16034 , n16035 , n16036 , n16037 , n16038 , n16039 , n16040 , n16041 , n16042 , n16043 , n16044 , n16045 , n16046 , n16047 , n16048 , n16049 , n16050 , n16051 , n16052 , n16053 , n16054 , n16055 , n16056 , n16057 , n16058 , n16059 , n16060 , n16061 , n16062 , n16063 , n16064 , n16065 , n16066 , n16067 , n16068 , n16069 , n16070 , n16071 , n16072 , n16073 , n16074 , n16075 , n16076 , n16077 , n16078 , n16079 , n16080 , n16081 , n16082 , n16083 , n16084 , n16085 , n16086 , n16087 , n16088 , n16089 , n16090 , n16091 , n16092 , n16093 , n16094 , n16095 , n16096 , n16097 , n16098 , n16099 , n16100 , n16101 , n16102 , n16103 , n16104 , n16105 , n16106 , n16107 , n16108 , n16109 , n16110 , n16111 , n16112 , n16113 , n16114 , n16115 , n16116 , n16117 , n16118 , n16119 , n16120 , n16121 , n16122 , n16123 , n16124 , n16125 , n16126 , n16127 , n16128 , n16129 , n16130 , n16131 , n16132 , n16133 , n16134 , n16135 , n16136 , n16137 , n16138 , n16139 , n16140 , n16141 , n16142 , n16143 , n16144 , n16145 , n16146 , n16147 , n16148 , n16149 , n16150 , n16151 , n16152 , n16153 , n16154 , n16155 , n16156 , n16157 , n16158 , n16159 , n16160 , n16161 , n16162 , n16163 , n16164 , n16165 , n16166 , n16167 , n16168 , n16169 , n16170 , n16171 , n16172 , n16173 , n16174 , n16175 , n16176 , n16177 , n16178 , n16179 , n16180 , n16181 , n16182 , n16183 , n16184 , n16185 , n16186 , n16187 , n16188 , n16189 , n16190 , n16191 , n16192 , n16193 , n16194 , n16195 , n16196 , n16197 , n16198 , n16199 , n16200 , n16201 , n16202 , n16203 , n16204 , n16205 , n16206 , n16207 , n16208 , n16209 , n16210 , n16211 , n16212 , n16213 , n16214 , n16215 , n16216 , n16217 , n16218 , n16219 , n16220 , n16221 , n16222 , n16223 , n16224 , n16225 , n16226 , n16227 , n16228 , n16229 , n16230 , n16231 , n16232 , n16233 , n16234 , n16235 , n16236 , n16237 , n16238 , n16239 , n16240 , n16241 , n16242 , n16243 , n16244 , n16245 , n16246 , n16247 , n16248 , n16249 , n16250 , n16251 , n16252 , n16253 , n16254 , n16255 , n16256 , n16257 , n16258 , n16259 , n16260 , n16261 , n16262 , n16263 , n16264 , n16265 , n16266 , n16267 , n16268 , n16269 , n16270 , n16271 , n16272 , n16273 , n16274 , n16275 , n16276 , n16277 , n16278 , n16279 , n16280 , n16281 , n16282 , n16283 , n16284 , n16285 , n16286 , n16287 , n16288 , n16289 , n16290 , n16291 , n16292 , n16293 , n16294 , n16295 , n16296 , n16297 , n16298 , n16299 , n16300 , n16301 , n16302 , n16303 , n16304 , n16305 , n16306 , n16307 , n16308 , n16309 , n16310 , n16311 , n16312 , n16313 , n16314 , n16315 , n16316 , n16317 , n16318 , n16319 , n16320 , n16321 , n16322 , n16323 , n16324 , n16325 , n16326 , n16327 , n16328 , n16329 , n16330 , n16331 , n16332 , n16333 , n16334 , n16335 , n16336 , n16337 , n16338 , n16339 , n16340 , n16341 , n16342 , n16343 , n16344 , n16345 , n16346 , n16347 , n16348 , n16349 , n16350 , n16351 , n16352 , n16353 , n16354 , n16355 , n16356 , n16357 , n16358 , n16359 , n16360 , n16361 , n16362 , n16363 , n16364 , n16365 , n16366 , n16367 , n16368 , n16369 , n16370 , n16371 , n16372 , n16373 , n16374 , n16375 , n16376 , n16377 , n16378 , n16379 , n16380 , n16381 , n16382 , n16383 , n16384 , n16385 , n16386 , n16387 , n16388 , n16389 , n16390 , n16391 , n16392 , n16393 , n16394 , n16395 , n16396 , n16397 , n16398 , n16399 , n16400 , n16401 , n16402 , n16403 , n16404 , n16405 , n16406 , n16407 , n16408 , n16409 , n16410 , n16411 , n16412 , n16413 , n16414 , n16415 , n16416 , n16417 , n16418 , n16419 , n16420 , n16421 , n16422 , n16423 , n16424 , n16425 , n16426 , n16427 , n16428 , n16429 , n16430 , n16431 , n16432 , n16433 , n16434 , n16435 , n16436 , n16437 , n16438 , n16439 , n16440 , n16441 , n16442 , n16443 , n16444 , n16445 , n16446 , n16447 , n16448 , n16449 , n16450 , n16451 , n16452 , n16453 , n16454 , n16455 , n16456 , n16457 , n16458 , n16459 , n16460 , n16461 , n16462 , n16463 , n16464 , n16465 , n16466 , n16467 , n16468 , n16469 , n16470 , n16471 , n16472 , n16473 , n16474 , n16475 , n16476 , n16477 , n16478 , n16479 , n16480 , n16481 , n16482 , n16483 , n16484 , n16485 , n16486 , n16487 , n16488 , n16489 , n16490 , n16491 , n16492 , n16493 , n16494 , n16495 , n16496 , n16497 , n16498 , n16499 , n16500 , n16501 , n16502 , n16503 , n16504 , n16505 , n16506 , n16507 , n16508 , n16509 , n16510 , n16511 , n16512 , n16513 , n16514 , n16515 , n16516 , n16517 , n16518 , n16519 , n16520 , n16521 , n16522 , n16523 , n16524 , n16525 , n16526 , n16527 , n16528 , n16529 , n16530 , n16531 , n16532 , n16533 , n16534 , n16535 , n16536 , n16537 , n16538 , n16539 , n16540 , n16541 , n16542 , n16543 , n16544 , n16545 , n16546 , n16547 , n16548 , n16549 , n16550 , n16551 , n16552 , n16553 , n16554 , n16555 , n16556 , n16557 , n16558 , n16559 , n16560 , n16561 , n16562 , n16563 , n16564 , n16565 , n16566 , n16567 , n16568 , n16569 , n16570 , n16571 , n16572 , n16573 , n16574 , n16575 , n16576 , n16577 , n16578 , n16579 , n16580 , n16581 , n16582 , n16583 , n16584 , n16585 , n16586 , n16587 , n16588 , n16589 , n16590 , n16591 , n16592 , n16593 , n16594 , n16595 , n16596 , n16597 , n16598 , n16599 , n16600 , n16601 , n16602 , n16603 , n16604 , n16605 , n16606 , n16607 , n16608 , n16609 , n16610 , n16611 , n16612 , n16613 , n16614 , n16615 , n16616 , n16617 , n16618 , n16619 , n16620 , n16621 , n16622 , n16623 , n16624 , n16625 , n16626 , n16627 , n16628 , n16629 , n16630 , n16631 , n16632 , n16633 , n16634 , n16635 , n16636 , n16637 , n16638 , n16639 , n16640 , n16641 , n16642 , n16643 , n16644 , n16645 , n16646 , n16647 , n16648 , n16649 , n16650 , n16651 , n16652 , n16653 , n16654 , n16655 , n16656 , n16657 , n16658 , n16659 , n16660 , n16661 , n16662 , n16663 , n16664 , n16665 , n16666 , n16667 , n16668 , n16669 , n16670 , n16671 , n16672 , n16673 , n16674 , n16675 , n16676 , n16677 , n16678 , n16679 , n16680 , n16681 , n16682 , n16683 , n16684 , n16685 , n16686 , n16687 , n16688 , n16689 , n16690 , n16691 , n16692 , n16693 , n16694 , n16695 , n16696 , n16697 , n16698 , n16699 , n16700 , n16701 , n16702 , n16703 , n16704 , n16705 , n16706 , n16707 , n16708 , n16709 , n16710 , n16711 , n16712 , n16713 , n16714 , n16715 , n16716 , n16717 , n16718 , n16719 , n16720 , n16721 , n16722 , n16723 , n16724 , n16725 , n16726 , n16727 , n16728 , n16729 , n16730 , n16731 , n16732 , n16733 , n16734 , n16735 , n16736 , n16737 , n16738 , n16739 , n16740 , n16741 , n16742 , n16743 , n16744 , n16745 , n16746 , n16747 , n16748 , n16749 , n16750 , n16751 , n16752 , n16753 , n16754 , n16755 , n16756 , n16757 , n16758 , n16759 , n16760 , n16761 , n16762 , n16763 , n16764 , n16765 , n16766 , n16767 , n16768 , n16769 , n16770 , n16771 , n16772 , n16773 , n16774 , n16775 , n16776 , n16777 , n16778 , n16779 , n16780 , n16781 , n16782 , n16783 , n16784 , n16785 , n16786 , n16787 , n16788 , n16789 , n16790 , n16791 , n16792 , n16793 , n16794 , n16795 , n16796 , n16797 , n16798 , n16799 , n16800 , n16801 , n16802 , n16803 , n16804 , n16805 , n16806 , n16807 , n16808 , n16809 , n16810 , n16811 , n16812 , n16813 , n16814 , n16815 , n16816 , n16817 , n16818 , n16819 , n16820 , n16821 , n16822 , n16823 , n16824 , n16825 , n16826 , n16827 , n16828 , n16829 , n16830 , n16831 , n16832 , n16833 , n16834 , n16835 , n16836 , n16837 , n16838 , n16839 , n16840 , n16841 , n16842 , n16843 , n16844 , n16845 , n16846 , n16847 , n16848 , n16849 , n16850 , n16851 , n16852 , n16853 , n16854 , n16855 , n16856 , n16857 , n16858 , n16859 , n16860 , n16861 , n16862 , n16863 , n16864 , n16865 , n16866 , n16867 , n16868 , n16869 , n16870 , n16871 , n16872 , n16873 , n16874 , n16875 , n16876 , n16877 , n16878 , n16879 , n16880 , n16881 , n16882 , n16883 , n16884 , n16885 , n16886 , n16887 , n16888 , n16889 , n16890 , n16891 , n16892 , n16893 , n16894 , n16895 , n16896 , n16897 , n16898 , n16899 , n16900 , n16901 , n16902 , n16903 , n16904 , n16905 , n16906 , n16907 , n16908 , n16909 , n16910 , n16911 , n16912 , n16913 , n16914 , n16915 , n16916 , n16917 , n16918 , n16919 , n16920 , n16921 , n16922 , n16923 , n16924 , n16925 , n16926 , n16927 , n16928 , n16929 , n16930 , n16931 , n16932 , n16933 , n16934 , n16935 , n16936 , n16937 , n16938 , n16939 , n16940 , n16941 , n16942 , n16943 , n16944 , n16945 , n16946 , n16947 , n16948 , n16949 , n16950 , n16951 , n16952 , n16953 , n16954 , n16955 , n16956 , n16957 , n16958 , n16959 , n16960 , n16961 , n16962 , n16963 , n16964 , n16965 , n16966 , n16967 , n16968 , n16969 , n16970 , n16971 , n16972 , n16973 , n16974 , n16975 , n16976 , n16977 , n16978 , n16979 , n16980 , n16981 , n16982 , n16983 , n16984 , n16985 , n16986 , n16987 , n16988 , n16989 , n16990 , n16991 , n16992 , n16993 , n16994 , n16995 , n16996 , n16997 , n16998 , n16999 , n17000 , n17001 , n17002 , n17003 , n17004 , n17005 , n17006 , n17007 , n17008 , n17009 , n17010 , n17011 , n17012 , n17013 , n17014 , n17015 , n17016 , n17017 , n17018 , n17019 , n17020 , n17021 , n17022 , n17023 , n17024 , n17025 , n17026 , n17027 , n17028 , n17029 , n17030 , n17031 , n17032 , n17033 , n17034 , n17035 , n17036 , n17037 , n17038 , n17039 , n17040 , n17041 , n17042 , n17043 , n17044 , n17045 , n17046 , n17047 , n17048 , n17049 , n17050 , n17051 , n17052 , n17053 , n17054 , n17055 , n17056 , n17057 , n17058 , n17059 , n17060 , n17061 , n17062 , n17063 , n17064 , n17065 , n17066 , n17067 , n17068 , n17069 , n17070 , n17071 , n17072 , n17073 , n17074 , n17075 , n17076 , n17077 , n17078 , n17079 , n17080 , n17081 , n17082 , n17083 , n17084 , n17085 , n17086 , n17087 , n17088 , n17089 , n17090 , n17091 , n17092 , n17093 , n17094 , n17095 , n17096 , n17097 , n17098 , n17099 , n17100 , n17101 , n17102 , n17103 , n17104 , n17105 , n17106 , n17107 , n17108 , n17109 , n17110 , n17111 , n17112 , n17113 , n17114 , n17115 , n17116 , n17117 , n17118 , n17119 , n17120 , n17121 , n17122 , n17123 , n17124 , n17125 , n17126 , n17127 , n17128 , n17129 , n17130 , n17131 , n17132 , n17133 , n17134 , n17135 , n17136 , n17137 , n17138 , n17139 , n17140 , n17141 , n17142 , n17143 , n17144 , n17145 , n17146 , n17147 , n17148 , n17149 , n17150 , n17151 , n17152 , n17153 , n17154 , n17155 , n17156 , n17157 , n17158 , n17159 , n17160 , n17161 , n17162 , n17163 , n17164 , n17165 , n17166 , n17167 , n17168 , n17169 , n17170 , n17171 , n17172 , n17173 , n17174 , n17175 , n17176 , n17177 , n17178 , n17179 , n17180 , n17181 , n17182 , n17183 , n17184 , n17185 , n17186 , n17187 , n17188 , n17189 , n17190 , n17191 , n17192 , n17193 , n17194 , n17195 , n17196 , n17197 , n17198 , n17199 , n17200 , n17201 , n17202 , n17203 , n17204 , n17205 , n17206 , n17207 , n17208 , n17209 , n17210 , n17211 , n17212 , n17213 , n17214 , n17215 , n17216 , n17217 , n17218 , n17219 , n17220 , n17221 , n17222 , n17223 , n17224 , n17225 , n17226 , n17227 , n17228 , n17229 , n17230 , n17231 , n17232 , n17233 , n17234 , n17235 , n17236 , n17237 , n17238 , n17239 , n17240 , n17241 , n17242 , n17243 , n17244 , n17245 , n17246 , n17247 , n17248 , n17249 , n17250 , n17251 , n17252 , n17253 , n17254 , n17255 , n17256 , n17257 , n17258 , n17259 , n17260 , n17261 , n17262 , n17263 , n17264 , n17265 , n17266 , n17267 , n17268 , n17269 , n17270 , n17271 , n17272 , n17273 , n17274 , n17275 , n17276 , n17277 , n17278 , n17279 , n17280 , n17281 , n17282 , n17283 , n17284 , n17285 , n17286 , n17287 , n17288 , n17289 , n17290 , n17291 , n17292 , n17293 , n17294 , n17295 , n17296 , n17297 , n17298 , n17299 , n17300 , n17301 , n17302 , n17303 , n17304 , n17305 , n17306 , n17307 , n17308 , n17309 , n17310 , n17311 , n17312 , n17313 , n17314 , n17315 , n17316 , n17317 , n17318 , n17319 , n17320 , n17321 , n17322 , n17323 , n17324 , n17325 , n17326 , n17327 , n17328 , n17329 , n17330 , n17331 , n17332 , n17333 , n17334 , n17335 , n17336 , n17337 , n17338 , n17339 , n17340 , n17341 , n17342 , n17343 , n17344 , n17345 , n17346 , n17347 , n17348 , n17349 , n17350 , n17351 , n17352 , n17353 , n17354 , n17355 , n17356 , n17357 , n17358 , n17359 , n17360 , n17361 , n17362 , n17363 , n17364 , n17365 , n17366 , n17367 , n17368 , n17369 , n17370 , n17371 , n17372 , n17373 , n17374 , n17375 , n17376 , n17377 , n17378 , n17379 , n17380 , n17381 , n17382 , n17383 , n17384 , n17385 , n17386 , n17387 , n17388 , n17389 , n17390 , n17391 , n17392 , n17393 , n17394 , n17395 , n17396 , n17397 , n17398 , n17399 , n17400 , n17401 , n17402 , n17403 , n17404 , n17405 , n17406 , n17407 , n17408 , n17409 , n17410 , n17411 , n17412 , n17413 , n17414 , n17415 , n17416 , n17417 , n17418 , n17419 , n17420 , n17421 , n17422 , n17423 , n17424 , n17425 , n17426 , n17427 , n17428 , n17429 , n17430 , n17431 , n17432 , n17433 , n17434 , n17435 , n17436 , n17437 , n17438 , n17439 , n17440 , n17441 , n17442 , n17443 , n17444 , n17445 , n17446 , n17447 , n17448 , n17449 , n17450 , n17451 , n17452 , n17453 , n17454 , n17455 , n17456 , n17457 , n17458 , n17459 , n17460 , n17461 , n17462 , n17463 , n17464 , n17465 , n17466 , n17467 , n17468 , n17469 , n17470 , n17471 , n17472 , n17473 , n17474 , n17475 , n17476 , n17477 , n17478 , n17479 , n17480 , n17481 , n17482 , n17483 , n17484 , n17485 , n17486 , n17487 , n17488 , n17489 , n17490 , n17491 , n17492 , n17493 , n17494 , n17495 , n17496 , n17497 , n17498 , n17499 , n17500 , n17501 , n17502 , n17503 , n17504 , n17505 , n17506 , n17507 , n17508 , n17509 , n17510 , n17511 , n17512 , n17513 , n17514 , n17515 , n17516 , n17517 , n17518 , n17519 , n17520 , n17521 , n17522 , n17523 , n17524 , n17525 , n17526 , n17527 , n17528 , n17529 , n17530 , n17531 , n17532 , n17533 , n17534 , n17535 , n17536 , n17537 , n17538 , n17539 , n17540 , n17541 , n17542 , n17543 , n17544 , n17545 , n17546 , n17547 , n17548 , n17549 , n17550 , n17551 , n17552 , n17553 , n17554 , n17555 , n17556 , n17557 , n17558 , n17559 , n17560 , n17561 , n17562 , n17563 , n17564 , n17565 , n17566 , n17567 , n17568 , n17569 , n17570 , n17571 , n17572 , n17573 , n17574 , n17575 , n17576 , n17577 , n17578 , n17579 , n17580 , n17581 , n17582 , n17583 , n17584 , n17585 , n17586 , n17587 , n17588 , n17589 , n17590 , n17591 , n17592 , n17593 , n17594 , n17595 , n17596 , n17597 , n17598 , n17599 , n17600 , n17601 , n17602 , n17603 , n17604 , n17605 , n17606 , n17607 , n17608 , n17609 , n17610 , n17611 , n17612 , n17613 , n17614 , n17615 , n17616 , n17617 , n17618 , n17619 , n17620 , n17621 , n17622 , n17623 , n17624 , n17625 , n17626 , n17627 , n17628 , n17629 , n17630 , n17631 , n17632 , n17633 , n17634 , n17635 , n17636 , n17637 , n17638 , n17639 , n17640 , n17641 , n17642 , n17643 , n17644 , n17645 , n17646 , n17647 , n17648 , n17649 , n17650 , n17651 , n17652 , n17653 , n17654 , n17655 , n17656 , n17657 , n17658 , n17659 , n17660 , n17661 , n17662 , n17663 , n17664 , n17665 , n17666 , n17667 , n17668 , n17669 , n17670 , n17671 , n17672 , n17673 , n17674 , n17675 , n17676 , n17677 , n17678 , n17679 , n17680 , n17681 , n17682 , n17683 , n17684 , n17685 , n17686 , n17687 , n17688 , n17689 , n17690 , n17691 , n17692 , n17693 , n17694 , n17695 , n17696 , n17697 , n17698 , n17699 , n17700 , n17701 , n17702 , n17703 , n17704 , n17705 , n17706 , n17707 , n17708 , n17709 , n17710 , n17711 , n17712 , n17713 , n17714 , n17715 , n17716 , n17717 , n17718 , n17719 , n17720 , n17721 , n17722 , n17723 , n17724 , n17725 , n17726 , n17727 , n17728 , n17729 , n17730 , n17731 , n17732 , n17733 , n17734 , n17735 , n17736 , n17737 , n17738 , n17739 , n17740 , n17741 , n17742 , n17743 , n17744 , n17745 , n17746 , n17747 , n17748 , n17749 , n17750 , n17751 , n17752 , n17753 , n17754 , n17755 , n17756 , n17757 , n17758 , n17759 , n17760 , n17761 , n17762 , n17763 , n17764 , n17765 , n17766 , n17767 , n17768 , n17769 , n17770 , n17771 , n17772 , n17773 , n17774 , n17775 , n17776 , n17777 , n17778 , n17779 , n17780 , n17781 , n17782 , n17783 , n17784 , n17785 , n17786 , n17787 , n17788 , n17789 , n17790 , n17791 , n17792 , n17793 , n17794 , n17795 , n17796 , n17797 , n17798 , n17799 , n17800 , n17801 , n17802 , n17803 , n17804 , n17805 , n17806 , n17807 , n17808 , n17809 , n17810 , n17811 , n17812 , n17813 , n17814 , n17815 , n17816 , n17817 , n17818 , n17819 , n17820 , n17821 , n17822 , n17823 , n17824 , n17825 , n17826 , n17827 , n17828 , n17829 , n17830 , n17831 , n17832 , n17833 , n17834 , n17835 , n17836 , n17837 , n17838 , n17839 , n17840 , n17841 , n17842 , n17843 , n17844 , n17845 , n17846 , n17847 , n17848 , n17849 , n17850 , n17851 , n17852 , n17853 , n17854 , n17855 , n17856 , n17857 , n17858 , n17859 , n17860 , n17861 , n17862 , n17863 , n17864 , n17865 , n17866 , n17867 , n17868 , n17869 , n17870 , n17871 , n17872 , n17873 , n17874 , n17875 , n17876 , n17877 , n17878 , n17879 , n17880 , n17881 , n17882 , n17883 , n17884 , n17885 , n17886 , n17887 , n17888 , n17889 , n17890 , n17891 , n17892 , n17893 , n17894 , n17895 , n17896 , n17897 , n17898 , n17899 , n17900 , n17901 , n17902 , n17903 , n17904 , n17905 , n17906 , n17907 , n17908 , n17909 , n17910 , n17911 , n17912 , n17913 , n17914 , n17915 , n17916 , n17917 , n17918 , n17919 , n17920 , n17921 , n17922 , n17923 , n17924 , n17925 , n17926 , n17927 , n17928 , n17929 , n17930 , n17931 , n17932 , n17933 , n17934 , n17935 , n17936 , n17937 , n17938 , n17939 , n17940 , n17941 , n17942 , n17943 , n17944 , n17945 , n17946 , n17947 , n17948 , n17949 , n17950 , n17951 , n17952 , n17953 , n17954 , n17955 , n17956 , n17957 , n17958 , n17959 , n17960 , n17961 , n17962 , n17963 , n17964 , n17965 , n17966 , n17967 , n17968 , n17969 , n17970 , n17971 , n17972 , n17973 , n17974 , n17975 , n17976 , n17977 , n17978 , n17979 , n17980 , n17981 , n17982 , n17983 , n17984 , n17985 , n17986 , n17987 , n17988 , n17989 , n17990 , n17991 , n17992 , n17993 , n17994 , n17995 , n17996 , n17997 , n17998 , n17999 , n18000 , n18001 , n18002 , n18003 , n18004 , n18005 , n18006 , n18007 , n18008 , n18009 , n18010 , n18011 , n18012 , n18013 , n18014 , n18015 , n18016 , n18017 , n18018 , n18019 , n18020 , n18021 , n18022 , n18023 , n18024 , n18025 , n18026 , n18027 , n18028 , n18029 , n18030 , n18031 , n18032 , n18033 , n18034 , n18035 , n18036 , n18037 , n18038 , n18039 , n18040 , n18041 , n18042 , n18043 , n18044 , n18045 , n18046 , n18047 , n18048 , n18049 , n18050 , n18051 , n18052 , n18053 , n18054 , n18055 , n18056 , n18057 , n18058 , n18059 , n18060 , n18061 , n18062 , n18063 , n18064 , n18065 , n18066 , n18067 , n18068 , n18069 , n18070 , n18071 , n18072 , n18073 , n18074 , n18075 , n18076 , n18077 , n18078 , n18079 , n18080 , n18081 , n18082 , n18083 , n18084 , n18085 , n18086 , n18087 , n18088 , n18089 , n18090 , n18091 , n18092 , n18093 , n18094 , n18095 , n18096 , n18097 , n18098 , n18099 , n18100 , n18101 , n18102 , n18103 , n18104 , n18105 , n18106 , n18107 , n18108 , n18109 , n18110 , n18111 , n18112 , n18113 , n18114 , n18115 , n18116 , n18117 , n18118 , n18119 , n18120 , n18121 , n18122 , n18123 , n18124 , n18125 , n18126 , n18127 , n18128 , n18129 , n18130 , n18131 , n18132 , n18133 , n18134 , n18135 , n18136 , n18137 , n18138 , n18139 , n18140 , n18141 , n18142 , n18143 , n18144 , n18145 , n18146 , n18147 , n18148 , n18149 , n18150 , n18151 , n18152 , n18153 , n18154 , n18155 , n18156 , n18157 , n18158 , n18159 , n18160 , n18161 , n18162 , n18163 , n18164 , n18165 , n18166 , n18167 , n18168 , n18169 , n18170 , n18171 , n18172 , n18173 , n18174 , n18175 , n18176 , n18177 , n18178 , n18179 , n18180 , n18181 , n18182 , n18183 , n18184 , n18185 , n18186 , n18187 , n18188 , n18189 , n18190 , n18191 , n18192 , n18193 , n18194 , n18195 , n18196 , n18197 , n18198 , n18199 , n18200 , n18201 , n18202 , n18203 , n18204 , n18205 , n18206 , n18207 , n18208 , n18209 , n18210 , n18211 , n18212 , n18213 , n18214 , n18215 , n18216 , n18217 , n18218 , n18219 , n18220 , n18221 , n18222 , n18223 , n18224 , n18225 , n18226 , n18227 , n18228 , n18229 , n18230 , n18231 , n18232 , n18233 , n18234 , n18235 , n18236 , n18237 , n18238 , n18239 , n18240 , n18241 , n18242 , n18243 , n18244 , n18245 , n18246 , n18247 , n18248 , n18249 , n18250 , n18251 , n18252 , n18253 , n18254 , n18255 , n18256 , n18257 , n18258 , n18259 , n18260 , n18261 , n18262 , n18263 , n18264 , n18265 , n18266 , n18267 , n18268 , n18269 , n18270 , n18271 , n18272 , n18273 , n18274 , n18275 , n18276 , n18277 , n18278 , n18279 , n18280 , n18281 , n18282 , n18283 , n18284 , n18285 , n18286 , n18287 , n18288 , n18289 , n18290 , n18291 , n18292 , n18293 , n18294 , n18295 , n18296 , n18297 , n18298 , n18299 , n18300 , n18301 , n18302 , n18303 , n18304 , n18305 , n18306 , n18307 , n18308 , n18309 , n18310 , n18311 , n18312 , n18313 , n18314 , n18315 , n18316 , n18317 , n18318 , n18319 , n18320 , n18321 , n18322 , n18323 , n18324 , n18325 , n18326 , n18327 , n18328 , n18329 , n18330 , n18331 , n18332 , n18333 , n18334 , n18335 , n18336 , n18337 , n18338 , n18339 , n18340 , n18341 , n18342 , n18343 , n18344 , n18345 , n18346 , n18347 , n18348 , n18349 , n18350 , n18351 , n18352 , n18353 , n18354 , n18355 , n18356 , n18357 , n18358 , n18359 , n18360 , n18361 , n18362 , n18363 , n18364 , n18365 , n18366 , n18367 , n18368 , n18369 , n18370 , n18371 , n18372 , n18373 , n18374 , n18375 , n18376 , n18377 , n18378 , n18379 , n18380 , n18381 , n18382 , n18383 , n18384 , n18385 , n18386 , n18387 , n18388 , n18389 , n18390 , n18391 , n18392 , n18393 , n18394 , n18395 , n18396 , n18397 , n18398 , n18399 , n18400 , n18401 , n18402 , n18403 , n18404 , n18405 , n18406 , n18407 , n18408 , n18409 , n18410 , n18411 , n18412 , n18413 , n18414 , n18415 , n18416 , n18417 , n18418 , n18419 , n18420 , n18421 , n18422 , n18423 , n18424 , n18425 , n18426 , n18427 , n18428 , n18429 , n18430 , n18431 , n18432 , n18433 , n18434 , n18435 , n18436 , n18437 , n18438 , n18439 , n18440 , n18441 , n18442 , n18443 , n18444 , n18445 , n18446 , n18447 , n18448 , n18449 , n18450 , n18451 , n18452 , n18453 , n18454 , n18455 , n18456 , n18457 , n18458 , n18459 , n18460 , n18461 , n18462 , n18463 , n18464 , n18465 , n18466 , n18467 , n18468 , n18469 , n18470 , n18471 , n18472 , n18473 , n18474 , n18475 , n18476 , n18477 , n18478 , n18479 , n18480 , n18481 , n18482 , n18483 , n18484 , n18485 , n18486 , n18487 , n18488 , n18489 , n18490 , n18491 , n18492 , n18493 , n18494 , n18495 , n18496 , n18497 , n18498 , n18499 , n18500 , n18501 , n18502 , n18503 , n18504 , n18505 , n18506 , n18507 , n18508 , n18509 , n18510 , n18511 , n18512 , n18513 , n18514 , n18515 , n18516 , n18517 , n18518 , n18519 , n18520 , n18521 , n18522 , n18523 , n18524 , n18525 , n18526 , n18527 , n18528 , n18529 , n18530 , n18531 , n18532 , n18533 , n18534 , n18535 , n18536 , n18537 , n18538 , n18539 , n18540 , n18541 , n18542 , n18543 , n18544 , n18545 , n18546 , n18547 , n18548 , n18549 , n18550 , n18551 , n18552 , n18553 , n18554 , n18555 , n18556 , n18557 , n18558 , n18559 , n18560 , n18561 , n18562 , n18563 , n18564 , n18565 , n18566 , n18567 , n18568 , n18569 , n18570 , n18571 , n18572 , n18573 , n18574 , n18575 , n18576 , n18577 , n18578 , n18579 , n18580 , n18581 , n18582 , n18583 , n18584 , n18585 , n18586 , n18587 , n18588 , n18589 , n18590 , n18591 , n18592 , n18593 , n18594 , n18595 , n18596 , n18597 , n18598 , n18599 , n18600 , n18601 , n18602 , n18603 , n18604 , n18605 , n18606 , n18607 , n18608 , n18609 , n18610 , n18611 , n18612 , n18613 , n18614 , n18615 , n18616 , n18617 , n18618 , n18619 , n18620 , n18621 , n18622 , n18623 , n18624 , n18625 , n18626 , n18627 , n18628 , n18629 , n18630 , n18631 , n18632 , n18633 , n18634 , n18635 , n18636 , n18637 , n18638 , n18639 , n18640 , n18641 , n18642 , n18643 , n18644 , n18645 , n18646 , n18647 , n18648 , n18649 , n18650 , n18651 , n18652 , n18653 , n18654 , n18655 , n18656 , n18657 , n18658 , n18659 , n18660 , n18661 , n18662 , n18663 , n18664 , n18665 , n18666 , n18667 , n18668 , n18669 , n18670 , n18671 , n18672 , n18673 , n18674 , n18675 , n18676 , n18677 , n18678 , n18679 , n18680 , n18681 , n18682 , n18683 , n18684 , n18685 , n18686 , n18687 , n18688 , n18689 , n18690 , n18691 , n18692 , n18693 , n18694 , n18695 , n18696 , n18697 , n18698 , n18699 , n18700 , n18701 , n18702 , n18703 , n18704 , n18705 , n18706 , n18707 , n18708 , n18709 , n18710 , n18711 , n18712 , n18713 , n18714 , n18715 , n18716 , n18717 , n18718 , n18719 , n18720 , n18721 , n18722 , n18723 , n18724 , n18725 , n18726 , n18727 , n18728 , n18729 , n18730 , n18731 , n18732 , n18733 , n18734 , n18735 , n18736 , n18737 , n18738 , n18739 , n18740 , n18741 , n18742 , n18743 , n18744 , n18745 , n18746 , n18747 , n18748 , n18749 , n18750 , n18751 , n18752 , n18753 , n18754 , n18755 , n18756 , n18757 , n18758 , n18759 , n18760 , n18761 , n18762 , n18763 , n18764 , n18765 , n18766 , n18767 , n18768 , n18769 , n18770 , n18771 , n18772 , n18773 , n18774 , n18775 , n18776 , n18777 , n18778 , n18779 , n18780 , n18781 , n18782 , n18783 , n18784 , n18785 , n18786 , n18787 , n18788 , n18789 , n18790 , n18791 , n18792 , n18793 , n18794 , n18795 , n18796 , n18797 , n18798 , n18799 , n18800 , n18801 , n18802 , n18803 , n18804 , n18805 , n18806 , n18807 , n18808 , n18809 , n18810 , n18811 , n18812 , n18813 , n18814 , n18815 , n18816 , n18817 , n18818 , n18819 , n18820 , n18821 , n18822 , n18823 , n18824 , n18825 , n18826 , n18827 , n18828 , n18829 , n18830 , n18831 , n18832 , n18833 , n18834 , n18835 , n18836 , n18837 , n18838 , n18839 , n18840 , n18841 , n18842 , n18843 , n18844 , n18845 , n18846 , n18847 , n18848 , n18849 , n18850 , n18851 , n18852 , n18853 , n18854 , n18855 , n18856 , n18857 , n18858 , n18859 , n18860 , n18861 , n18862 , n18863 , n18864 , n18865 , n18866 , n18867 , n18868 , n18869 , n18870 , n18871 , n18872 , n18873 , n18874 , n18875 , n18876 , n18877 , n18878 , n18879 , n18880 , n18881 , n18882 , n18883 , n18884 , n18885 , n18886 , n18887 , n18888 , n18889 , n18890 , n18891 , n18892 , n18893 , n18894 , n18895 , n18896 , n18897 , n18898 , n18899 , n18900 , n18901 , n18902 , n18903 , n18904 , n18905 , n18906 , n18907 , n18908 , n18909 , n18910 , n18911 , n18912 , n18913 , n18914 , n18915 , n18916 , n18917 , n18918 , n18919 , n18920 , n18921 , n18922 , n18923 , n18924 , n18925 , n18926 , n18927 , n18928 , n18929 , n18930 , n18931 , n18932 , n18933 , n18934 , n18935 , n18936 , n18937 , n18938 , n18939 , n18940 , n18941 , n18942 , n18943 , n18944 , n18945 , n18946 , n18947 , n18948 , n18949 , n18950 , n18951 , n18952 , n18953 , n18954 , n18955 , n18956 , n18957 , n18958 , n18959 , n18960 , n18961 , n18962 , n18963 , n18964 , n18965 , n18966 , n18967 , n18968 , n18969 , n18970 , n18971 , n18972 , n18973 , n18974 , n18975 , n18976 , n18977 , n18978 , n18979 , n18980 , n18981 , n18982 , n18983 , n18984 , n18985 , n18986 , n18987 , n18988 , n18989 , n18990 , n18991 , n18992 , n18993 , n18994 , n18995 , n18996 , n18997 , n18998 , n18999 , n19000 , n19001 , n19002 , n19003 , n19004 , n19005 , n19006 , n19007 , n19008 , n19009 , n19010 , n19011 , n19012 , n19013 , n19014 , n19015 , n19016 , n19017 , n19018 , n19019 , n19020 , n19021 , n19022 , n19023 , n19024 , n19025 , n19026 , n19027 , n19028 , n19029 , n19030 , n19031 , n19032 , n19033 , n19034 , n19035 , n19036 , n19037 , n19038 , n19039 , n19040 , n19041 , n19042 , n19043 , n19044 , n19045 , n19046 , n19047 , n19048 , n19049 , n19050 , n19051 , n19052 , n19053 , n19054 , n19055 , n19056 , n19057 , n19058 , n19059 , n19060 , n19061 , n19062 , n19063 , n19064 , n19065 , n19066 , n19067 , n19068 , n19069 , n19070 , n19071 , n19072 , n19073 , n19074 , n19075 , n19076 , n19077 , n19078 , n19079 , n19080 , n19081 , n19082 , n19083 , n19084 , n19085 , n19086 , n19087 , n19088 , n19089 , n19090 , n19091 , n19092 , n19093 , n19094 , n19095 , n19096 , n19097 , n19098 , n19099 , n19100 , n19101 , n19102 , n19103 , n19104 , n19105 , n19106 , n19107 , n19108 , n19109 , n19110 , n19111 , n19112 , n19113 , n19114 , n19115 , n19116 , n19117 , n19118 , n19119 , n19120 , n19121 , n19122 , n19123 , n19124 , n19125 , n19126 , n19127 , n19128 , n19129 , n19130 , n19131 , n19132 , n19133 , n19134 , n19135 , n19136 , n19137 , n19138 , n19139 , n19140 , n19141 , n19142 , n19143 , n19144 , n19145 , n19146 , n19147 , n19148 , n19149 , n19150 , n19151 , n19152 , n19153 , n19154 , n19155 , n19156 , n19157 , n19158 , n19159 , n19160 , n19161 , n19162 , n19163 , n19164 , n19165 , n19166 , n19167 , n19168 , n19169 , n19170 , n19171 , n19172 , n19173 , n19174 , n19175 , n19176 , n19177 , n19178 , n19179 , n19180 , n19181 , n19182 , n19183 , n19184 , n19185 , n19186 , n19187 , n19188 , n19189 , n19190 , n19191 , n19192 , n19193 , n19194 , n19195 , n19196 , n19197 , n19198 , n19199 , n19200 , n19201 , n19202 , n19203 , n19204 , n19205 , n19206 , n19207 , n19208 , n19209 , n19210 , n19211 , n19212 , n19213 , n19214 , n19215 , n19216 , n19217 , n19218 , n19219 , n19220 , n19221 , n19222 , n19223 , n19224 , n19225 , n19226 , n19227 , n19228 , n19229 , n19230 , n19231 , n19232 , n19233 , n19234 , n19235 , n19236 , n19237 , n19238 , n19239 , n19240 , n19241 , n19242 , n19243 , n19244 , n19245 , n19246 , n19247 , n19248 , n19249 , n19250 , n19251 , n19252 , n19253 , n19254 , n19255 , n19256 , n19257 , n19258 , n19259 , n19260 , n19261 , n19262 , n19263 , n19264 , n19265 , n19266 , n19267 , n19268 , n19269 , n19270 , n19271 , n19272 , n19273 , n19274 , n19275 , n19276 , n19277 , n19278 , n19279 , n19280 , n19281 , n19282 , n19283 , n19284 , n19285 , n19286 , n19287 , n19288 , n19289 , n19290 , n19291 , n19292 , n19293 , n19294 , n19295 , n19296 , n19297 , n19298 , n19299 , n19300 , n19301 , n19302 , n19303 , n19304 , n19305 , n19306 , n19307 , n19308 , n19309 , n19310 , n19311 , n19312 , n19313 , n19314 , n19315 , n19316 , n19317 , n19318 , n19319 , n19320 , n19321 , n19322 , n19323 , n19324 , n19325 , n19326 , n19327 , n19328 , n19329 , n19330 , n19331 , n19332 , n19333 , n19334 , n19335 , n19336 , n19337 , n19338 , n19339 , n19340 , n19341 , n19342 , n19343 , n19344 , n19345 , n19346 , n19347 , n19348 , n19349 , n19350 , n19351 , n19352 , n19353 , n19354 , n19355 , n19356 , n19357 , n19358 , n19359 , n19360 , n19361 , n19362 , n19363 , n19364 , n19365 , n19366 , n19367 , n19368 , n19369 , n19370 , n19371 , n19372 , n19373 , n19374 , n19375 , n19376 , n19377 , n19378 , n19379 , n19380 , n19381 , n19382 , n19383 , n19384 , n19385 , n19386 , n19387 , n19388 , n19389 , n19390 , n19391 , n19392 , n19393 , n19394 , n19395 , n19396 , n19397 , n19398 , n19399 , n19400 , n19401 , n19402 , n19403 , n19404 , n19405 , n19406 , n19407 , n19408 , n19409 , n19410 , n19411 , n19412 , n19413 , n19414 , n19415 , n19416 , n19417 , n19418 , n19419 , n19420 , n19421 , n19422 , n19423 , n19424 , n19425 , n19426 , n19427 , n19428 , n19429 , n19430 , n19431 , n19432 , n19433 , n19434 , n19435 , n19436 , n19437 , n19438 , n19439 , n19440 , n19441 , n19442 , n19443 , n19444 , n19445 , n19446 , n19447 , n19448 , n19449 , n19450 , n19451 , n19452 , n19453 , n19454 , n19455 , n19456 , n19457 , n19458 , n19459 , n19460 , n19461 , n19462 , n19463 , n19464 , n19465 , n19466 , n19467 , n19468 , n19469 , n19470 , n19471 , n19472 , n19473 , n19474 , n19475 , n19476 , n19477 , n19478 , n19479 , n19480 , n19481 , n19482 , n19483 , n19484 , n19485 , n19486 , n19487 , n19488 , n19489 , n19490 , n19491 , n19492 , n19493 , n19494 , n19495 , n19496 , n19497 , n19498 , n19499 , n19500 , n19501 , n19502 , n19503 , n19504 , n19505 , n19506 , n19507 , n19508 , n19509 , n19510 , n19511 , n19512 , n19513 , n19514 , n19515 , n19516 , n19517 , n19518 , n19519 , n19520 , n19521 , n19522 , n19523 , n19524 , n19525 , n19526 , n19527 , n19528 , n19529 , n19530 , n19531 , n19532 , n19533 , n19534 , n19535 , n19536 , n19537 , n19538 , n19539 , n19540 , n19541 , n19542 , n19543 , n19544 , n19545 , n19546 , n19547 , n19548 , n19549 , n19550 , n19551 , n19552 , n19553 , n19554 , n19555 , n19556 , n19557 , n19558 , n19559 , n19560 , n19561 , n19562 , n19563 , n19564 , n19565 , n19566 , n19567 , n19568 , n19569 , n19570 , n19571 , n19572 , n19573 , n19574 , n19575 , n19576 , n19577 , n19578 , n19579 , n19580 , n19581 , n19582 , n19583 , n19584 , n19585 , n19586 , n19587 , n19588 , n19589 , n19590 , n19591 , n19592 , n19593 , n19594 , n19595 , n19596 , n19597 , n19598 , n19599 , n19600 , n19601 , n19602 , n19603 , n19604 , n19605 , n19606 , n19607 , n19608 , n19609 , n19610 , n19611 , n19612 , n19613 , n19614 , n19615 , n19616 , n19617 , n19618 , n19619 , n19620 , n19621 , n19622 , n19623 , n19624 , n19625 , n19626 , n19627 , n19628 , n19629 , n19630 , n19631 , n19632 , n19633 , n19634 , n19635 , n19636 , n19637 , n19638 , n19639 , n19640 , n19641 , n19642 , n19643 , n19644 , n19645 , n19646 , n19647 , n19648 , n19649 , n19650 , n19651 , n19652 , n19653 , n19654 , n19655 , n19656 , n19657 , n19658 , n19659 , n19660 , n19661 , n19662 , n19663 , n19664 , n19665 , n19666 , n19667 , n19668 , n19669 , n19670 , n19671 , n19672 , n19673 , n19674 , n19675 , n19676 , n19677 , n19678 , n19679 , n19680 , n19681 , n19682 , n19683 , n19684 , n19685 , n19686 , n19687 , n19688 , n19689 , n19690 , n19691 , n19692 , n19693 , n19694 , n19695 , n19696 , n19697 , n19698 , n19699 , n19700 , n19701 , n19702 , n19703 , n19704 , n19705 , n19706 , n19707 , n19708 , n19709 , n19710 , n19711 , n19712 , n19713 , n19714 , n19715 , n19716 , n19717 , n19718 , n19719 , n19720 , n19721 , n19722 , n19723 , n19724 , n19725 , n19726 , n19727 , n19728 , n19729 , n19730 , n19731 , n19732 , n19733 , n19734 , n19735 , n19736 , n19737 , n19738 , n19739 , n19740 , n19741 , n19742 , n19743 , n19744 , n19745 , n19746 , n19747 , n19748 , n19749 , n19750 , n19751 , n19752 , n19753 , n19754 , n19755 , n19756 , n19757 , n19758 , n19759 , n19760 , n19761 , n19762 , n19763 , n19764 , n19765 , n19766 , n19767 , n19768 , n19769 , n19770 , n19771 , n19772 , n19773 , n19774 , n19775 , n19776 , n19777 , n19778 , n19779 , n19780 , n19781 , n19782 , n19783 , n19784 , n19785 , n19786 , n19787 , n19788 , n19789 , n19790 , n19791 , n19792 , n19793 , n19794 , n19795 , n19796 , n19797 , n19798 , n19799 , n19800 , n19801 , n19802 , n19803 , n19804 , n19805 , n19806 , n19807 , n19808 , n19809 , n19810 , n19811 , n19812 , n19813 , n19814 , n19815 , n19816 , n19817 , n19818 , n19819 , n19820 , n19821 , n19822 , n19823 , n19824 , n19825 , n19826 , n19827 , n19828 , n19829 , n19830 , n19831 , n19832 , n19833 , n19834 , n19835 , n19836 , n19837 , n19838 , n19839 , n19840 , n19841 , n19842 , n19843 , n19844 , n19845 , n19846 , n19847 , n19848 , n19849 , n19850 , n19851 , n19852 , n19853 , n19854 , n19855 , n19856 , n19857 , n19858 , n19859 , n19860 , n19861 , n19862 , n19863 , n19864 , n19865 , n19866 , n19867 , n19868 , n19869 , n19870 , n19871 , n19872 , n19873 , n19874 , n19875 , n19876 , n19877 , n19878 , n19879 , n19880 , n19881 , n19882 , n19883 , n19884 , n19885 , n19886 , n19887 , n19888 , n19889 , n19890 , n19891 , n19892 , n19893 , n19894 , n19895 , n19896 , n19897 , n19898 , n19899 , n19900 , n19901 , n19902 , n19903 , n19904 , n19905 , n19906 , n19907 , n19908 , n19909 , n19910 , n19911 , n19912 , n19913 , n19914 , n19915 , n19916 , n19917 , n19918 , n19919 , n19920 , n19921 , n19922 , n19923 , n19924 , n19925 , n19926 , n19927 , n19928 , n19929 , n19930 , n19931 , n19932 , n19933 , n19934 , n19935 , n19936 , n19937 , n19938 , n19939 , n19940 , n19941 , n19942 , n19943 , n19944 , n19945 , n19946 , n19947 , n19948 , n19949 , n19950 , n19951 , n19952 , n19953 , n19954 , n19955 , n19956 , n19957 , n19958 , n19959 , n19960 , n19961 , n19962 , n19963 , n19964 , n19965 , n19966 , n19967 , n19968 , n19969 , n19970 , n19971 , n19972 , n19973 , n19974 , n19975 , n19976 , n19977 , n19978 , n19979 , n19980 , n19981 , n19982 , n19983 , n19984 , n19985 , n19986 , n19987 , n19988 , n19989 , n19990 , n19991 , n19992 , n19993 , n19994 , n19995 , n19996 , n19997 , n19998 , n19999 , n20000 , n20001 , n20002 , n20003 , n20004 , n20005 , n20006 , n20007 , n20008 , n20009 , n20010 , n20011 , n20012 , n20013 , n20014 , n20015 , n20016 , n20017 , n20018 , n20019 , n20020 , n20021 , n20022 , n20023 , n20024 , n20025 , n20026 , n20027 , n20028 , n20029 , n20030 , n20031 , n20032 , n20033 , n20034 , n20035 , n20036 , n20037 , n20038 , n20039 , n20040 , n20041 , n20042 , n20043 , n20044 , n20045 , n20046 , n20047 , n20048 , n20049 , n20050 , n20051 , n20052 , n20053 , n20054 , n20055 , n20056 , n20057 , n20058 , n20059 , n20060 , n20061 , n20062 , n20063 , n20064 , n20065 , n20066 , n20067 , n20068 , n20069 , n20070 , n20071 , n20072 , n20073 , n20074 , n20075 , n20076 , n20077 , n20078 , n20079 , n20080 , n20081 , n20082 , n20083 , n20084 , n20085 , n20086 , n20087 , n20088 , n20089 , n20090 , n20091 , n20092 , n20093 , n20094 , n20095 , n20096 , n20097 , n20098 , n20099 , n20100 , n20101 , n20102 , n20103 , n20104 , n20105 , n20106 , n20107 , n20108 , n20109 , n20110 , n20111 , n20112 , n20113 , n20114 , n20115 , n20116 , n20117 , n20118 , n20119 , n20120 , n20121 , n20122 , n20123 , n20124 , n20125 , n20126 , n20127 , n20128 , n20129 , n20130 , n20131 , n20132 , n20133 , n20134 , n20135 , n20136 , n20137 , n20138 , n20139 , n20140 , n20141 , n20142 , n20143 , n20144 , n20145 , n20146 , n20147 , n20148 , n20149 , n20150 , n20151 , n20152 , n20153 , n20154 , n20155 , n20156 , n20157 , n20158 , n20159 , n20160 , n20161 , n20162 , n20163 , n20164 , n20165 , n20166 , n20167 , n20168 , n20169 , n20170 , n20171 , n20172 , n20173 , n20174 , n20175 , n20176 , n20177 , n20178 , n20179 , n20180 , n20181 , n20182 , n20183 , n20184 , n20185 , n20186 , n20187 , n20188 , n20189 , n20190 , n20191 , n20192 , n20193 , n20194 , n20195 , n20196 , n20197 , n20198 , n20199 , n20200 , n20201 , n20202 , n20203 , n20204 , n20205 , n20206 , n20207 , n20208 , n20209 , n20210 , n20211 , n20212 , n20213 , n20214 , n20215 , n20216 , n20217 , n20218 , n20219 , n20220 , n20221 , n20222 , n20223 , n20224 , n20225 , n20226 , n20227 , n20228 , n20229 , n20230 , n20231 , n20232 , n20233 , n20234 , n20235 , n20236 , n20237 , n20238 , n20239 , n20240 , n20241 , n20242 , n20243 , n20244 , n20245 , n20246 , n20247 , n20248 , n20249 , n20250 , n20251 , n20252 , n20253 , n20254 , n20255 , n20256 , n20257 , n20258 , n20259 , n20260 , n20261 , n20262 , n20263 , n20264 , n20265 , n20266 , n20267 , n20268 , n20269 , n20270 , n20271 , n20272 , n20273 , n20274 , n20275 , n20276 , n20277 , n20278 , n20279 , n20280 , n20281 , n20282 , n20283 , n20284 , n20285 , n20286 , n20287 , n20288 , n20289 , n20290 , n20291 , n20292 , n20293 , n20294 , n20295 , n20296 , n20297 , n20298 , n20299 , n20300 , n20301 , n20302 , n20303 , n20304 , n20305 , n20306 , n20307 , n20308 , n20309 , n20310 , n20311 , n20312 , n20313 , n20314 , n20315 , n20316 , n20317 , n20318 , n20319 , n20320 , n20321 , n20322 , n20323 , n20324 , n20325 , n20326 , n20327 , n20328 , n20329 , n20330 , n20331 , n20332 , n20333 , n20334 , n20335 , n20336 , n20337 , n20338 , n20339 , n20340 , n20341 , n20342 , n20343 , n20344 , n20345 , n20346 , n20347 , n20348 , n20349 , n20350 , n20351 , n20352 , n20353 , n20354 , n20355 , n20356 , n20357 , n20358 , n20359 , n20360 , n20361 , n20362 , n20363 , n20364 , n20365 , n20366 , n20367 , n20368 , n20369 , n20370 , n20371 , n20372 , n20373 , n20374 , n20375 , n20376 , n20377 , n20378 , n20379 , n20380 , n20381 , n20382 , n20383 , n20384 , n20385 , n20386 , n20387 , n20388 , n20389 , n20390 , n20391 , n20392 , n20393 , n20394 , n20395 , n20396 , n20397 , n20398 , n20399 , n20400 , n20401 , n20402 , n20403 , n20404 , n20405 , n20406 , n20407 , n20408 , n20409 , n20410 , n20411 , n20412 , n20413 , n20414 , n20415 , n20416 , n20417 , n20418 , n20419 , n20420 , n20421 , n20422 , n20423 , n20424 , n20425 , n20426 , n20427 , n20428 , n20429 , n20430 , n20431 , n20432 , n20433 , n20434 , n20435 , n20436 , n20437 , n20438 , n20439 , n20440 , n20441 , n20442 , n20443 , n20444 , n20445 , n20446 , n20447 , n20448 , n20449 , n20450 , n20451 , n20452 , n20453 , n20454 , n20455 , n20456 , n20457 , n20458 , n20459 , n20460 , n20461 , n20462 , n20463 , n20464 , n20465 , n20466 , n20467 , n20468 , n20469 , n20470 , n20471 , n20472 , n20473 , n20474 , n20475 , n20476 , n20477 , n20478 , n20479 , n20480 , n20481 , n20482 , n20483 , n20484 , n20485 , n20486 , n20487 , n20488 , n20489 , n20490 , n20491 , n20492 , n20493 , n20494 , n20495 , n20496 , n20497 , n20498 , n20499 , n20500 , n20501 , n20502 , n20503 , n20504 , n20505 , n20506 , n20507 , n20508 , n20509 , n20510 , n20511 , n20512 , n20513 , n20514 , n20515 , n20516 , n20517 , n20518 , n20519 , n20520 , n20521 , n20522 , n20523 , n20524 , n20525 , n20526 , n20527 , n20528 , n20529 , n20530 , n20531 , n20532 , n20533 , n20534 , n20535 , n20536 , n20537 , n20538 , n20539 , n20540 , n20541 , n20542 , n20543 , n20544 , n20545 , n20546 , n20547 , n20548 , n20549 , n20550 , n20551 , n20552 , n20553 , n20554 , n20555 , n20556 , n20557 , n20558 , n20559 , n20560 , n20561 , n20562 , n20563 , n20564 , n20565 , n20566 , n20567 , n20568 , n20569 , n20570 , n20571 , n20572 , n20573 , n20574 , n20575 , n20576 , n20577 , n20578 , n20579 , n20580 , n20581 , n20582 , n20583 , n20584 , n20585 , n20586 , n20587 , n20588 , n20589 , n20590 , n20591 , n20592 , n20593 , n20594 , n20595 , n20596 , n20597 , n20598 , n20599 , n20600 , n20601 , n20602 , n20603 , n20604 , n20605 , n20606 , n20607 , n20608 , n20609 , n20610 , n20611 , n20612 , n20613 , n20614 , n20615 , n20616 , n20617 , n20618 , n20619 , n20620 , n20621 , n20622 , n20623 , n20624 , n20625 , n20626 , n20627 , n20628 , n20629 , n20630 , n20631 , n20632 , n20633 , n20634 , n20635 , n20636 , n20637 , n20638 , n20639 , n20640 , n20641 , n20642 , n20643 , n20644 , n20645 , n20646 , n20647 , n20648 , n20649 , n20650 , n20651 , n20652 , n20653 , n20654 , n20655 , n20656 , n20657 , n20658 , n20659 , n20660 , n20661 , n20662 , n20663 , n20664 , n20665 , n20666 , n20667 , n20668 , n20669 , n20670 , n20671 , n20672 , n20673 , n20674 , n20675 , n20676 , n20677 , n20678 , n20679 , n20680 , n20681 , n20682 , n20683 , n20684 , n20685 , n20686 , n20687 , n20688 , n20689 , n20690 , n20691 , n20692 , n20693 , n20694 , n20695 , n20696 , n20697 , n20698 , n20699 , n20700 , n20701 , n20702 , n20703 , n20704 , n20705 , n20706 , n20707 , n20708 , n20709 , n20710 , n20711 , n20712 , n20713 , n20714 , n20715 , n20716 , n20717 , n20718 , n20719 , n20720 , n20721 , n20722 , n20723 , n20724 , n20725 , n20726 , n20727 , n20728 , n20729 , n20730 , n20731 , n20732 , n20733 , n20734 , n20735 , n20736 , n20737 , n20738 , n20739 , n20740 , n20741 , n20742 , n20743 , n20744 , n20745 , n20746 , n20747 , n20748 , n20749 , n20750 , n20751 , n20752 , n20753 , n20754 , n20755 , n20756 , n20757 , n20758 , n20759 , n20760 , n20761 , n20762 , n20763 , n20764 , n20765 , n20766 , n20767 , n20768 , n20769 , n20770 , n20771 , n20772 , n20773 , n20774 , n20775 , n20776 , n20777 , n20778 , n20779 , n20780 , n20781 , n20782 , n20783 , n20784 , n20785 , n20786 , n20787 , n20788 , n20789 , n20790 , n20791 , n20792 , n20793 , n20794 , n20795 , n20796 , n20797 , n20798 , n20799 , n20800 , n20801 , n20802 , n20803 , n20804 , n20805 , n20806 , n20807 , n20808 , n20809 , n20810 , n20811 , n20812 , n20813 , n20814 , n20815 , n20816 , n20817 , n20818 , n20819 , n20820 , n20821 , n20822 , n20823 , n20824 , n20825 , n20826 , n20827 , n20828 , n20829 , n20830 , n20831 , n20832 , n20833 , n20834 , n20835 , n20836 , n20837 , n20838 , n20839 , n20840 , n20841 , n20842 , n20843 , n20844 , n20845 , n20846 , n20847 , n20848 , n20849 , n20850 , n20851 , n20852 , n20853 , n20854 , n20855 , n20856 , n20857 , n20858 , n20859 , n20860 , n20861 , n20862 , n20863 , n20864 , n20865 , n20866 , n20867 , n20868 , n20869 , n20870 , n20871 , n20872 , n20873 , n20874 , n20875 , n20876 , n20877 , n20878 , n20879 , n20880 , n20881 , n20882 , n20883 , n20884 , n20885 , n20886 , n20887 , n20888 , n20889 , n20890 , n20891 , n20892 , n20893 , n20894 , n20895 , n20896 , n20897 , n20898 , n20899 , n20900 , n20901 , n20902 , n20903 , n20904 , n20905 , n20906 , n20907 , n20908 , n20909 , n20910 , n20911 , n20912 , n20913 , n20914 , n20915 , n20916 , n20917 , n20918 , n20919 , n20920 , n20921 , n20922 , n20923 , n20924 , n20925 , n20926 , n20927 , n20928 , n20929 , n20930 , n20931 , n20932 , n20933 , n20934 , n20935 , n20936 , n20937 , n20938 , n20939 , n20940 , n20941 , n20942 , n20943 , n20944 , n20945 , n20946 , n20947 , n20948 , n20949 , n20950 , n20951 , n20952 , n20953 , n20954 , n20955 , n20956 , n20957 , n20958 , n20959 , n20960 , n20961 , n20962 , n20963 , n20964 , n20965 , n20966 , n20967 , n20968 , n20969 , n20970 , n20971 , n20972 , n20973 , n20974 , n20975 , n20976 , n20977 , n20978 , n20979 , n20980 , n20981 , n20982 , n20983 , n20984 , n20985 , n20986 , n20987 , n20988 , n20989 , n20990 , n20991 , n20992 , n20993 , n20994 , n20995 , n20996 , n20997 , n20998 , n20999 , n21000 , n21001 , n21002 , n21003 , n21004 , n21005 , n21006 , n21007 , n21008 , n21009 , n21010 , n21011 , n21012 , n21013 , n21014 , n21015 , n21016 , n21017 , n21018 , n21019 , n21020 , n21021 , n21022 , n21023 , n21024 , n21025 , n21026 , n21027 , n21028 , n21029 , n21030 , n21031 , n21032 , n21033 , n21034 , n21035 , n21036 , n21037 , n21038 , n21039 , n21040 , n21041 , n21042 , n21043 , n21044 , n21045 , n21046 , n21047 , n21048 , n21049 , n21050 , n21051 , n21052 , n21053 , n21054 , n21055 , n21056 , n21057 , n21058 , n21059 , n21060 , n21061 , n21062 , n21063 , n21064 , n21065 , n21066 , n21067 , n21068 , n21069 , n21070 , n21071 , n21072 , n21073 , n21074 , n21075 , n21076 , n21077 , n21078 , n21079 , n21080 , n21081 , n21082 , n21083 , n21084 , n21085 , n21086 , n21087 , n21088 , n21089 , n21090 , n21091 , n21092 , n21093 , n21094 , n21095 , n21096 , n21097 , n21098 , n21099 , n21100 , n21101 , n21102 , n21103 , n21104 , n21105 , n21106 , n21107 , n21108 , n21109 , n21110 , n21111 , n21112 , n21113 , n21114 , n21115 , n21116 , n21117 , n21118 , n21119 , n21120 , n21121 , n21122 , n21123 , n21124 , n21125 , n21126 , n21127 , n21128 , n21129 , n21130 , n21131 , n21132 , n21133 , n21134 , n21135 , n21136 , n21137 , n21138 , n21139 , n21140 , n21141 , n21142 , n21143 , n21144 , n21145 , n21146 , n21147 , n21148 , n21149 , n21150 , n21151 , n21152 , n21153 , n21154 , n21155 , n21156 , n21157 , n21158 , n21159 , n21160 , n21161 , n21162 , n21163 , n21164 , n21165 , n21166 , n21167 , n21168 , n21169 , n21170 , n21171 , n21172 , n21173 , n21174 , n21175 , n21176 , n21177 , n21178 , n21179 , n21180 , n21181 , n21182 , n21183 , n21184 , n21185 , n21186 , n21187 , n21188 , n21189 , n21190 , n21191 , n21192 , n21193 , n21194 , n21195 , n21196 , n21197 , n21198 , n21199 , n21200 , n21201 , n21202 , n21203 , n21204 , n21205 , n21206 , n21207 , n21208 , n21209 , n21210 , n21211 , n21212 , n21213 , n21214 , n21215 , n21216 , n21217 , n21218 , n21219 , n21220 , n21221 , n21222 , n21223 , n21224 , n21225 , n21226 , n21227 , n21228 , n21229 , n21230 , n21231 , n21232 , n21233 , n21234 , n21235 , n21236 , n21237 , n21238 , n21239 , n21240 , n21241 , n21242 , n21243 , n21244 , n21245 , n21246 , n21247 , n21248 , n21249 , n21250 , n21251 , n21252 , n21253 , n21254 , n21255 , n21256 , n21257 , n21258 , n21259 , n21260 , n21261 , n21262 , n21263 , n21264 , n21265 , n21266 , n21267 , n21268 , n21269 , n21270 , n21271 , n21272 , n21273 , n21274 , n21275 , n21276 , n21277 , n21278 , n21279 , n21280 , n21281 , n21282 , n21283 , n21284 , n21285 , n21286 , n21287 , n21288 , n21289 , n21290 , n21291 , n21292 , n21293 , n21294 , n21295 , n21296 , n21297 , n21298 , n21299 , n21300 , n21301 , n21302 , n21303 , n21304 , n21305 , n21306 , n21307 , n21308 , n21309 , n21310 , n21311 , n21312 , n21313 , n21314 , n21315 , n21316 , n21317 , n21318 , n21319 , n21320 , n21321 , n21322 , n21323 , n21324 , n21325 , n21326 , n21327 , n21328 , n21329 , n21330 , n21331 , n21332 , n21333 , n21334 , n21335 , n21336 , n21337 , n21338 , n21339 , n21340 , n21341 , n21342 , n21343 , n21344 , n21345 , n21346 , n21347 , n21348 , n21349 , n21350 , n21351 , n21352 , n21353 , n21354 , n21355 , n21356 , n21357 , n21358 , n21359 , n21360 , n21361 , n21362 , n21363 , n21364 , n21365 , n21366 , n21367 , n21368 , n21369 , n21370 , n21371 , n21372 , n21373 , n21374 , n21375 , n21376 , n21377 , n21378 , n21379 , n21380 , n21381 , n21382 , n21383 , n21384 , n21385 , n21386 , n21387 , n21388 , n21389 , n21390 , n21391 , n21392 , n21393 , n21394 , n21395 , n21396 , n21397 , n21398 , n21399 , n21400 , n21401 , n21402 , n21403 , n21404 , n21405 , n21406 , n21407 , n21408 , n21409 , n21410 , n21411 , n21412 , n21413 , n21414 , n21415 , n21416 , n21417 , n21418 , n21419 , n21420 , n21421 , n21422 , n21423 , n21424 , n21425 , n21426 , n21427 , n21428 , n21429 , n21430 , n21431 , n21432 , n21433 , n21434 , n21435 , n21436 , n21437 , n21438 , n21439 , n21440 , n21441 , n21442 , n21443 , n21444 , n21445 , n21446 , n21447 , n21448 , n21449 , n21450 , n21451 , n21452 , n21453 , n21454 , n21455 , n21456 , n21457 , n21458 , n21459 , n21460 , n21461 , n21462 , n21463 , n21464 , n21465 , n21466 , n21467 , n21468 , n21469 , n21470 , n21471 , n21472 , n21473 , n21474 , n21475 , n21476 , n21477 , n21478 , n21479 , n21480 , n21481 , n21482 , n21483 , n21484 , n21485 , n21486 , n21487 , n21488 , n21489 , n21490 , n21491 , n21492 , n21493 , n21494 , n21495 , n21496 , n21497 , n21498 , n21499 , n21500 , n21501 , n21502 , n21503 , n21504 , n21505 , n21506 , n21507 , n21508 , n21509 , n21510 , n21511 , n21512 , n21513 , n21514 , n21515 , n21516 , n21517 , n21518 , n21519 , n21520 , n21521 , n21522 , n21523 , n21524 , n21525 , n21526 , n21527 , n21528 , n21529 , n21530 , n21531 , n21532 , n21533 , n21534 , n21535 , n21536 , n21537 , n21538 , n21539 , n21540 , n21541 , n21542 , n21543 , n21544 , n21545 , n21546 , n21547 , n21548 , n21549 , n21550 , n21551 , n21552 , n21553 , n21554 , n21555 , n21556 , n21557 , n21558 , n21559 , n21560 , n21561 , n21562 , n21563 , n21564 , n21565 , n21566 , n21567 , n21568 , n21569 , n21570 , n21571 , n21572 , n21573 , n21574 , n21575 , n21576 , n21577 , n21578 , n21579 , n21580 , n21581 , n21582 , n21583 , n21584 , n21585 , n21586 , n21587 , n21588 , n21589 , n21590 , n21591 , n21592 , n21593 , n21594 , n21595 , n21596 , n21597 , n21598 , n21599 , n21600 , n21601 , n21602 , n21603 , n21604 , n21605 , n21606 , n21607 , n21608 , n21609 , n21610 , n21611 , n21612 , n21613 , n21614 , n21615 , n21616 , n21617 , n21618 , n21619 , n21620 , n21621 , n21622 , n21623 , n21624 , n21625 , n21626 , n21627 , n21628 , n21629 , n21630 , n21631 , n21632 , n21633 , n21634 , n21635 , n21636 , n21637 , n21638 , n21639 , n21640 , n21641 , n21642 , n21643 , n21644 , n21645 , n21646 , n21647 , n21648 , n21649 , n21650 , n21651 , n21652 , n21653 , n21654 , n21655 , n21656 , n21657 , n21658 , n21659 , n21660 , n21661 , n21662 , n21663 , n21664 , n21665 , n21666 , n21667 , n21668 , n21669 , n21670 , n21671 , n21672 , n21673 , n21674 , n21675 , n21676 , n21677 , n21678 , n21679 , n21680 , n21681 , n21682 , n21683 , n21684 , n21685 , n21686 , n21687 , n21688 , n21689 , n21690 , n21691 , n21692 , n21693 , n21694 , n21695 , n21696 , n21697 , n21698 , n21699 , n21700 , n21701 , n21702 , n21703 , n21704 , n21705 , n21706 , n21707 , n21708 , n21709 , n21710 , n21711 , n21712 , n21713 , n21714 , n21715 , n21716 , n21717 , n21718 , n21719 , n21720 , n21721 , n21722 , n21723 , n21724 , n21725 , n21726 , n21727 , n21728 , n21729 , n21730 , n21731 , n21732 , n21733 , n21734 , n21735 , n21736 , n21737 , n21738 , n21739 , n21740 , n21741 , n21742 , n21743 , n21744 , n21745 , n21746 , n21747 , n21748 , n21749 , n21750 , n21751 , n21752 , n21753 , n21754 , n21755 , n21756 , n21757 , n21758 , n21759 , n21760 , n21761 , n21762 , n21763 , n21764 , n21765 , n21766 , n21767 , n21768 , n21769 , n21770 , n21771 , n21772 , n21773 , n21774 , n21775 , n21776 , n21777 , n21778 , n21779 , n21780 , n21781 , n21782 , n21783 , n21784 , n21785 , n21786 , n21787 , n21788 , n21789 , n21790 , n21791 , n21792 , n21793 , n21794 , n21795 , n21796 , n21797 , n21798 , n21799 , n21800 , n21801 , n21802 , n21803 , n21804 , n21805 , n21806 , n21807 , n21808 , n21809 , n21810 , n21811 , n21812 , n21813 , n21814 , n21815 , n21816 , n21817 , n21818 , n21819 , n21820 , n21821 , n21822 , n21823 , n21824 , n21825 , n21826 , n21827 , n21828 , n21829 , n21830 , n21831 , n21832 , n21833 , n21834 , n21835 , n21836 , n21837 , n21838 , n21839 , n21840 , n21841 , n21842 , n21843 , n21844 , n21845 , n21846 , n21847 , n21848 , n21849 , n21850 , n21851 , n21852 , n21853 , n21854 , n21855 , n21856 , n21857 , n21858 , n21859 , n21860 , n21861 , n21862 , n21863 , n21864 , n21865 , n21866 , n21867 , n21868 , n21869 , n21870 , n21871 , n21872 , n21873 , n21874 , n21875 , n21876 , n21877 , n21878 , n21879 , n21880 , n21881 , n21882 , n21883 , n21884 , n21885 , n21886 , n21887 , n21888 , n21889 , n21890 , n21891 , n21892 , n21893 , n21894 , n21895 , n21896 , n21897 , n21898 , n21899 , n21900 , n21901 , n21902 , n21903 , n21904 , n21905 , n21906 , n21907 , n21908 , n21909 , n21910 , n21911 , n21912 , n21913 , n21914 , n21915 , n21916 , n21917 , n21918 , n21919 , n21920 , n21921 , n21922 , n21923 , n21924 , n21925 , n21926 , n21927 , n21928 , n21929 , n21930 , n21931 , n21932 , n21933 , n21934 , n21935 , n21936 , n21937 , n21938 , n21939 , n21940 , n21941 , n21942 , n21943 , n21944 , n21945 , n21946 , n21947 , n21948 , n21949 , n21950 , n21951 , n21952 , n21953 , n21954 , n21955 , n21956 , n21957 , n21958 , n21959 , n21960 , n21961 , n21962 , n21963 , n21964 , n21965 , n21966 , n21967 , n21968 , n21969 , n21970 , n21971 , n21972 , n21973 , n21974 , n21975 , n21976 , n21977 , n21978 , n21979 , n21980 , n21981 , n21982 , n21983 , n21984 , n21985 , n21986 , n21987 , n21988 , n21989 , n21990 , n21991 , n21992 , n21993 , n21994 , n21995 , n21996 , n21997 , n21998 , n21999 , n22000 , n22001 , n22002 , n22003 , n22004 , n22005 , n22006 , n22007 , n22008 , n22009 , n22010 , n22011 , n22012 , n22013 , n22014 , n22015 , n22016 , n22017 , n22018 , n22019 , n22020 , n22021 , n22022 , n22023 , n22024 , n22025 , n22026 , n22027 , n22028 , n22029 , n22030 , n22031 , n22032 , n22033 , n22034 , n22035 , n22036 , n22037 , n22038 , n22039 , n22040 , n22041 , n22042 , n22043 , n22044 , n22045 , n22046 , n22047 , n22048 , n22049 , n22050 , n22051 , n22052 , n22053 , n22054 , n22055 , n22056 , n22057 , n22058 , n22059 , n22060 , n22061 , n22062 , n22063 , n22064 , n22065 , n22066 , n22067 , n22068 , n22069 , n22070 , n22071 , n22072 , n22073 , n22074 , n22075 , n22076 , n22077 , n22078 , n22079 , n22080 , n22081 , n22082 , n22083 , n22084 , n22085 , n22086 , n22087 , n22088 , n22089 , n22090 , n22091 , n22092 , n22093 , n22094 , n22095 , n22096 , n22097 , n22098 , n22099 , n22100 , n22101 , n22102 , n22103 , n22104 , n22105 , n22106 , n22107 , n22108 , n22109 , n22110 , n22111 , n22112 , n22113 , n22114 , n22115 , n22116 , n22117 , n22118 , n22119 , n22120 , n22121 , n22122 , n22123 , n22124 , n22125 , n22126 , n22127 , n22128 , n22129 , n22130 , n22131 , n22132 , n22133 , n22134 , n22135 , n22136 , n22137 , n22138 , n22139 , n22140 , n22141 , n22142 , n22143 , n22144 , n22145 , n22146 , n22147 , n22148 , n22149 , n22150 , n22151 , n22152 , n22153 , n22154 , n22155 , n22156 , n22157 , n22158 , n22159 , n22160 , n22161 , n22162 , n22163 , n22164 , n22165 , n22166 , n22167 , n22168 , n22169 , n22170 , n22171 , n22172 , n22173 , n22174 , n22175 , n22176 , n22177 , n22178 , n22179 , n22180 , n22181 , n22182 , n22183 , n22184 , n22185 , n22186 , n22187 , n22188 , n22189 , n22190 , n22191 , n22192 , n22193 , n22194 , n22195 , n22196 , n22197 , n22198 , n22199 , n22200 , n22201 , n22202 , n22203 , n22204 , n22205 , n22206 , n22207 , n22208 , n22209 , n22210 , n22211 , n22212 , n22213 , n22214 , n22215 , n22216 , n22217 , n22218 , n22219 , n22220 , n22221 , n22222 , n22223 , n22224 , n22225 , n22226 , n22227 , n22228 , n22229 , n22230 , n22231 , n22232 , n22233 , n22234 , n22235 , n22236 , n22237 , n22238 , n22239 , n22240 , n22241 , n22242 , n22243 , n22244 , n22245 , n22246 , n22247 , n22248 , n22249 , n22250 , n22251 , n22252 , n22253 , n22254 , n22255 , n22256 , n22257 , n22258 , n22259 , n22260 , n22261 , n22262 , n22263 , n22264 , n22265 , n22266 , n22267 , n22268 , n22269 , n22270 , n22271 , n22272 , n22273 , n22274 , n22275 , n22276 , n22277 , n22278 , n22279 , n22280 , n22281 , n22282 , n22283 , n22284 , n22285 , n22286 , n22287 , n22288 , n22289 , n22290 , n22291 , n22292 , n22293 , n22294 , n22295 , n22296 , n22297 , n22298 , n22299 , n22300 , n22301 , n22302 , n22303 , n22304 , n22305 , n22306 , n22307 , n22308 , n22309 , n22310 , n22311 , n22312 , n22313 , n22314 , n22315 , n22316 , n22317 , n22318 , n22319 , n22320 , n22321 , n22322 , n22323 , n22324 , n22325 , n22326 , n22327 , n22328 , n22329 , n22330 , n22331 , n22332 , n22333 , n22334 , n22335 , n22336 , n22337 , n22338 , n22339 , n22340 , n22341 , n22342 , n22343 , n22344 , n22345 , n22346 , n22347 , n22348 , n22349 , n22350 , n22351 , n22352 , n22353 , n22354 , n22355 , n22356 , n22357 , n22358 , n22359 , n22360 , n22361 , n22362 , n22363 , n22364 , n22365 , n22366 , n22367 , n22368 , n22369 , n22370 , n22371 , n22372 , n22373 , n22374 , n22375 , n22376 , n22377 , n22378 , n22379 , n22380 , n22381 , n22382 , n22383 , n22384 , n22385 , n22386 , n22387 , n22388 , n22389 , n22390 , n22391 , n22392 , n22393 , n22394 , n22395 , n22396 , n22397 , n22398 , n22399 , n22400 , n22401 , n22402 , n22403 , n22404 , n22405 , n22406 , n22407 , n22408 , n22409 , n22410 , n22411 , n22412 , n22413 , n22414 , n22415 , n22416 , n22417 , n22418 , n22419 , n22420 , n22421 , n22422 , n22423 , n22424 , n22425 , n22426 , n22427 , n22428 , n22429 , n22430 , n22431 , n22432 , n22433 , n22434 , n22435 , n22436 , n22437 , n22438 , n22439 , n22440 , n22441 , n22442 , n22443 , n22444 , n22445 , n22446 , n22447 , n22448 , n22449 , n22450 , n22451 , n22452 , n22453 , n22454 , n22455 , n22456 , n22457 , n22458 , n22459 , n22460 , n22461 , n22462 , n22463 , n22464 , n22465 , n22466 , n22467 , n22468 , n22469 , n22470 , n22471 , n22472 , n22473 , n22474 , n22475 , n22476 , n22477 , n22478 , n22479 , n22480 , n22481 , n22482 , n22483 , n22484 , n22485 , n22486 , n22487 , n22488 , n22489 , n22490 , n22491 , n22492 , n22493 , n22494 , n22495 , n22496 , n22497 , n22498 , n22499 , n22500 , n22501 , n22502 , n22503 , n22504 , n22505 , n22506 , n22507 , n22508 , n22509 , n22510 , n22511 , n22512 , n22513 , n22514 , n22515 , n22516 , n22517 , n22518 , n22519 , n22520 , n22521 , n22522 , n22523 , n22524 , n22525 , n22526 , n22527 , n22528 , n22529 , n22530 , n22531 , n22532 , n22533 , n22534 , n22535 , n22536 , n22537 , n22538 , n22539 , n22540 , n22541 , n22542 , n22543 , n22544 , n22545 , n22546 , n22547 , n22548 , n22549 , n22550 , n22551 , n22552 , n22553 , n22554 , n22555 , n22556 , n22557 , n22558 , n22559 , n22560 , n22561 , n22562 , n22563 , n22564 , n22565 , n22566 , n22567 , n22568 , n22569 , n22570 , n22571 , n22572 , n22573 , n22574 , n22575 , n22576 , n22577 , n22578 , n22579 , n22580 , n22581 , n22582 , n22583 , n22584 , n22585 , n22586 , n22587 , n22588 , n22589 , n22590 , n22591 , n22592 , n22593 , n22594 , n22595 , n22596 , n22597 , n22598 , n22599 , n22600 , n22601 , n22602 , n22603 , n22604 , n22605 , n22606 , n22607 , n22608 , n22609 , n22610 , n22611 , n22612 , n22613 , n22614 , n22615 , n22616 , n22617 , n22618 , n22619 , n22620 , n22621 , n22622 , n22623 , n22624 , n22625 , n22626 , n22627 , n22628 , n22629 , n22630 , n22631 , n22632 , n22633 , n22634 , n22635 , n22636 , n22637 , n22638 , n22639 , n22640 , n22641 , n22642 , n22643 , n22644 , n22645 , n22646 , n22647 , n22648 , n22649 , n22650 , n22651 , n22652 , n22653 , n22654 , n22655 , n22656 , n22657 , n22658 , n22659 , n22660 , n22661 , n22662 , n22663 , n22664 , n22665 , n22666 , n22667 , n22668 , n22669 , n22670 , n22671 , n22672 , n22673 , n22674 , n22675 , n22676 , n22677 , n22678 , n22679 , n22680 , n22681 , n22682 , n22683 , n22684 , n22685 , n22686 , n22687 , n22688 , n22689 , n22690 , n22691 , n22692 , n22693 , n22694 , n22695 , n22696 , n22697 , n22698 , n22699 , n22700 , n22701 , n22702 , n22703 , n22704 , n22705 , n22706 , n22707 , n22708 , n22709 , n22710 , n22711 , n22712 , n22713 , n22714 , n22715 , n22716 , n22717 , n22718 , n22719 , n22720 , n22721 , n22722 , n22723 , n22724 , n22725 , n22726 , n22727 , n22728 , n22729 , n22730 , n22731 , n22732 , n22733 , n22734 , n22735 , n22736 , n22737 , n22738 , n22739 , n22740 , n22741 , n22742 , n22743 , n22744 , n22745 , n22746 , n22747 , n22748 , n22749 , n22750 , n22751 , n22752 , n22753 , n22754 , n22755 , n22756 , n22757 , n22758 , n22759 , n22760 , n22761 , n22762 , n22763 , n22764 , n22765 , n22766 , n22767 , n22768 , n22769 , n22770 , n22771 , n22772 , n22773 , n22774 , n22775 , n22776 , n22777 , n22778 , n22779 , n22780 , n22781 , n22782 , n22783 , n22784 , n22785 , n22786 , n22787 , n22788 , n22789 , n22790 , n22791 , n22792 , n22793 , n22794 , n22795 , n22796 , n22797 , n22798 , n22799 , n22800 , n22801 , n22802 , n22803 , n22804 , n22805 , n22806 , n22807 , n22808 , n22809 , n22810 , n22811 , n22812 , n22813 , n22814 , n22815 , n22816 , n22817 , n22818 , n22819 , n22820 , n22821 , n22822 , n22823 , n22824 , n22825 , n22826 , n22827 , n22828 , n22829 , n22830 , n22831 , n22832 , n22833 , n22834 , n22835 , n22836 , n22837 , n22838 , n22839 , n22840 , n22841 , n22842 , n22843 , n22844 , n22845 , n22846 , n22847 , n22848 , n22849 , n22850 , n22851 , n22852 , n22853 , n22854 , n22855 , n22856 , n22857 , n22858 , n22859 , n22860 , n22861 , n22862 , n22863 , n22864 , n22865 , n22866 , n22867 , n22868 , n22869 , n22870 , n22871 , n22872 , n22873 , n22874 , n22875 , n22876 , n22877 , n22878 , n22879 , n22880 , n22881 , n22882 , n22883 , n22884 , n22885 , n22886 , n22887 , n22888 , n22889 , n22890 , n22891 , n22892 , n22893 , n22894 , n22895 , n22896 , n22897 , n22898 , n22899 , n22900 , n22901 , n22902 , n22903 , n22904 , n22905 , n22906 , n22907 , n22908 , n22909 , n22910 , n22911 , n22912 , n22913 , n22914 , n22915 , n22916 , n22917 , n22918 , n22919 , n22920 , n22921 , n22922 , n22923 , n22924 , n22925 , n22926 , n22927 , n22928 , n22929 , n22930 , n22931 , n22932 , n22933 , n22934 , n22935 , n22936 , n22937 , n22938 , n22939 , n22940 , n22941 , n22942 , n22943 , n22944 , n22945 , n22946 , n22947 , n22948 , n22949 , n22950 , n22951 , n22952 , n22953 , n22954 , n22955 , n22956 , n22957 , n22958 , n22959 , n22960 , n22961 , n22962 , n22963 , n22964 , n22965 , n22966 , n22967 , n22968 , n22969 , n22970 , n22971 , n22972 , n22973 , n22974 , n22975 , n22976 , n22977 , n22978 , n22979 , n22980 , n22981 , n22982 , n22983 , n22984 , n22985 , n22986 , n22987 , n22988 , n22989 , n22990 , n22991 , n22992 , n22993 , n22994 , n22995 , n22996 , n22997 , n22998 , n22999 , n23000 , n23001 , n23002 , n23003 , n23004 , n23005 , n23006 , n23007 , n23008 , n23009 , n23010 , n23011 , n23012 , n23013 , n23014 , n23015 , n23016 , n23017 , n23018 , n23019 , n23020 , n23021 , n23022 , n23023 , n23024 , n23025 , n23026 , n23027 , n23028 , n23029 , n23030 , n23031 , n23032 , n23033 , n23034 , n23035 , n23036 , n23037 , n23038 , n23039 , n23040 , n23041 , n23042 , n23043 , n23044 , n23045 , n23046 , n23047 , n23048 , n23049 , n23050 , n23051 , n23052 , n23053 , n23054 , n23055 , n23056 , n23057 , n23058 , n23059 , n23060 , n23061 , n23062 , n23063 , n23064 , n23065 , n23066 , n23067 , n23068 , n23069 , n23070 , n23071 , n23072 , n23073 , n23074 , n23075 , n23076 , n23077 , n23078 , n23079 , n23080 , n23081 , n23082 , n23083 , n23084 , n23085 , n23086 , n23087 , n23088 , n23089 , n23090 , n23091 , n23092 , n23093 , n23094 , n23095 , n23096 , n23097 , n23098 , n23099 , n23100 , n23101 , n23102 , n23103 , n23104 , n23105 , n23106 , n23107 , n23108 , n23109 , n23110 , n23111 , n23112 , n23113 , n23114 , n23115 , n23116 , n23117 , n23118 , n23119 , n23120 , n23121 , n23122 , n23123 , n23124 , n23125 , n23126 , n23127 , n23128 , n23129 , n23130 , n23131 , n23132 , n23133 , n23134 , n23135 , n23136 , n23137 , n23138 , n23139 , n23140 , n23141 , n23142 , n23143 , n23144 , n23145 , n23146 , n23147 , n23148 , n23149 , n23150 , n23151 , n23152 , n23153 , n23154 , n23155 , n23156 , n23157 , n23158 , n23159 , n23160 , n23161 , n23162 , n23163 , n23164 , n23165 , n23166 , n23167 , n23168 , n23169 , n23170 , n23171 , n23172 , n23173 , n23174 , n23175 , n23176 , n23177 , n23178 , n23179 , n23180 , n23181 , n23182 , n23183 , n23184 , n23185 , n23186 , n23187 , n23188 , n23189 , n23190 , n23191 , n23192 , n23193 , n23194 , n23195 , n23196 , n23197 , n23198 , n23199 , n23200 , n23201 , n23202 , n23203 , n23204 , n23205 , n23206 , n23207 , n23208 , n23209 , n23210 , n23211 , n23212 , n23213 , n23214 , n23215 , n23216 , n23217 , n23218 , n23219 , n23220 , n23221 , n23222 , n23223 , n23224 , n23225 , n23226 , n23227 , n23228 , n23229 , n23230 , n23231 , n23232 , n23233 , n23234 , n23235 , n23236 , n23237 , n23238 , n23239 , n23240 , n23241 , n23242 , n23243 , n23244 , n23245 , n23246 , n23247 , n23248 , n23249 , n23250 , n23251 , n23252 , n23253 , n23254 , n23255 , n23256 , n23257 , n23258 , n23259 , n23260 , n23261 , n23262 , n23263 , n23264 , n23265 , n23266 , n23267 , n23268 , n23269 , n23270 , n23271 , n23272 , n23273 , n23274 , n23275 , n23276 , n23277 , n23278 , n23279 , n23280 , n23281 , n23282 , n23283 , n23284 , n23285 , n23286 , n23287 , n23288 , n23289 , n23290 , n23291 , n23292 , n23293 , n23294 , n23295 , n23296 , n23297 , n23298 , n23299 , n23300 , n23301 , n23302 , n23303 , n23304 , n23305 , n23306 , n23307 , n23308 , n23309 , n23310 , n23311 , n23312 , n23313 , n23314 , n23315 , n23316 , n23317 , n23318 , n23319 , n23320 , n23321 , n23322 , n23323 , n23324 , n23325 , n23326 , n23327 , n23328 , n23329 , n23330 , n23331 , n23332 , n23333 , n23334 , n23335 , n23336 , n23337 , n23338 , n23339 , n23340 , n23341 , n23342 , n23343 , n23344 , n23345 , n23346 , n23347 , n23348 , n23349 , n23350 , n23351 , n23352 , n23353 , n23354 , n23355 , n23356 , n23357 , n23358 , n23359 , n23360 , n23361 , n23362 , n23363 , n23364 , n23365 , n23366 , n23367 , n23368 , n23369 , n23370 , n23371 , n23372 , n23373 , n23374 , n23375 , n23376 , n23377 , n23378 , n23379 , n23380 , n23381 , n23382 , n23383 , n23384 , n23385 , n23386 , n23387 , n23388 , n23389 , n23390 , n23391 , n23392 , n23393 , n23394 , n23395 , n23396 , n23397 , n23398 , n23399 , n23400 , n23401 , n23402 , n23403 , n23404 , n23405 , n23406 , n23407 , n23408 , n23409 , n23410 , n23411 , n23412 , n23413 , n23414 , n23415 , n23416 , n23417 , n23418 , n23419 , n23420 , n23421 , n23422 , n23423 , n23424 , n23425 , n23426 , n23427 , n23428 , n23429 , n23430 , n23431 , n23432 , n23433 , n23434 , n23435 , n23436 , n23437 , n23438 , n23439 , n23440 , n23441 , n23442 , n23443 , n23444 , n23445 , n23446 , n23447 , n23448 , n23449 , n23450 , n23451 , n23452 , n23453 , n23454 , n23455 , n23456 , n23457 , n23458 , n23459 , n23460 , n23461 , n23462 , n23463 , n23464 , n23465 , n23466 , n23467 , n23468 , n23469 , n23470 , n23471 , n23472 , n23473 , n23474 , n23475 , n23476 , n23477 , n23478 , n23479 , n23480 , n23481 , n23482 , n23483 , n23484 , n23485 , n23486 , n23487 , n23488 , n23489 , n23490 , n23491 , n23492 , n23493 , n23494 , n23495 , n23496 , n23497 , n23498 , n23499 , n23500 , n23501 , n23502 , n23503 , n23504 , n23505 , n23506 , n23507 , n23508 , n23509 , n23510 , n23511 , n23512 , n23513 , n23514 , n23515 , n23516 , n23517 , n23518 , n23519 , n23520 , n23521 , n23522 , n23523 , n23524 , n23525 , n23526 , n23527 , n23528 , n23529 , n23530 , n23531 , n23532 , n23533 , n23534 , n23535 , n23536 , n23537 , n23538 , n23539 , n23540 , n23541 , n23542 , n23543 , n23544 , n23545 , n23546 , n23547 , n23548 , n23549 , n23550 , n23551 , n23552 , n23553 , n23554 , n23555 , n23556 , n23557 , n23558 , n23559 , n23560 , n23561 , n23562 , n23563 , n23564 , n23565 , n23566 , n23567 , n23568 , n23569 , n23570 , n23571 , n23572 , n23573 , n23574 , n23575 , n23576 , n23577 , n23578 , n23579 , n23580 , n23581 , n23582 , n23583 , n23584 , n23585 , n23586 , n23587 , n23588 , n23589 , n23590 , n23591 , n23592 , n23593 , n23594 , n23595 , n23596 , n23597 , n23598 , n23599 , n23600 , n23601 , n23602 , n23603 , n23604 , n23605 , n23606 , n23607 , n23608 , n23609 , n23610 , n23611 , n23612 , n23613 , n23614 , n23615 , n23616 , n23617 , n23618 , n23619 , n23620 , n23621 , n23622 , n23623 , n23624 , n23625 , n23626 , n23627 , n23628 , n23629 , n23630 , n23631 , n23632 , n23633 , n23634 , n23635 , n23636 , n23637 , n23638 , n23639 , n23640 , n23641 , n23642 , n23643 , n23644 , n23645 , n23646 , n23647 , n23648 , n23649 , n23650 , n23651 , n23652 , n23653 , n23654 , n23655 , n23656 , n23657 , n23658 , n23659 , n23660 , n23661 , n23662 , n23663 , n23664 , n23665 , n23666 , n23667 , n23668 , n23669 , n23670 , n23671 , n23672 , n23673 , n23674 , n23675 , n23676 , n23677 , n23678 , n23679 , n23680 , n23681 , n23682 , n23683 , n23684 , n23685 , n23686 , n23687 , n23688 , n23689 , n23690 , n23691 , n23692 , n23693 , n23694 , n23695 , n23696 , n23697 , n23698 , n23699 , n23700 , n23701 , n23702 , n23703 , n23704 , n23705 , n23706 , n23707 , n23708 , n23709 , n23710 , n23711 , n23712 , n23713 , n23714 , n23715 , n23716 , n23717 , n23718 , n23719 , n23720 , n23721 , n23722 , n23723 , n23724 , n23725 , n23726 , n23727 , n23728 , n23729 , n23730 , n23731 , n23732 , n23733 , n23734 , n23735 , n23736 , n23737 , n23738 , n23739 , n23740 , n23741 , n23742 , n23743 , n23744 , n23745 , n23746 , n23747 , n23748 , n23749 , n23750 , n23751 , n23752 , n23753 , n23754 , n23755 , n23756 , n23757 , n23758 , n23759 , n23760 , n23761 , n23762 , n23763 , n23764 , n23765 , n23766 , n23767 , n23768 , n23769 , n23770 , n23771 , n23772 , n23773 , n23774 , n23775 , n23776 , n23777 , n23778 , n23779 , n23780 , n23781 , n23782 , n23783 , n23784 , n23785 , n23786 , n23787 , n23788 , n23789 , n23790 , n23791 , n23792 , n23793 , n23794 , n23795 , n23796 , n23797 , n23798 , n23799 , n23800 , n23801 , n23802 , n23803 , n23804 , n23805 , n23806 , n23807 , n23808 , n23809 , n23810 , n23811 , n23812 , n23813 , n23814 , n23815 , n23816 , n23817 , n23818 , n23819 , n23820 , n23821 , n23822 , n23823 , n23824 , n23825 , n23826 , n23827 , n23828 , n23829 , n23830 , n23831 , n23832 , n23833 , n23834 , n23835 , n23836 , n23837 , n23838 , n23839 , n23840 , n23841 , n23842 , n23843 , n23844 , n23845 , n23846 , n23847 , n23848 , n23849 , n23850 , n23851 , n23852 , n23853 , n23854 , n23855 , n23856 , n23857 , n23858 , n23859 , n23860 , n23861 , n23862 , n23863 , n23864 , n23865 , n23866 , n23867 , n23868 , n23869 , n23870 , n23871 , n23872 , n23873 , n23874 , n23875 , n23876 , n23877 , n23878 , n23879 , n23880 , n23881 , n23882 , n23883 , n23884 , n23885 , n23886 , n23887 , n23888 , n23889 , n23890 , n23891 , n23892 , n23893 , n23894 , n23895 , n23896 , n23897 , n23898 , n23899 , n23900 , n23901 , n23902 , n23903 , n23904 , n23905 , n23906 , n23907 , n23908 , n23909 , n23910 , n23911 , n23912 , n23913 , n23914 , n23915 , n23916 , n23917 , n23918 , n23919 , n23920 , n23921 , n23922 , n23923 , n23924 , n23925 , n23926 , n23927 , n23928 , n23929 , n23930 , n23931 , n23932 , n23933 , n23934 , n23935 , n23936 , n23937 , n23938 , n23939 , n23940 , n23941 , n23942 , n23943 , n23944 , n23945 , n23946 , n23947 , n23948 , n23949 , n23950 , n23951 , n23952 , n23953 , n23954 , n23955 , n23956 , n23957 , n23958 , n23959 , n23960 , n23961 , n23962 , n23963 , n23964 , n23965 , n23966 , n23967 , n23968 , n23969 , n23970 , n23971 , n23972 , n23973 , n23974 , n23975 , n23976 , n23977 , n23978 , n23979 , n23980 , n23981 , n23982 , n23983 , n23984 , n23985 , n23986 , n23987 , n23988 , n23989 , n23990 , n23991 , n23992 , n23993 , n23994 , n23995 , n23996 , n23997 , n23998 , n23999 , n24000 , n24001 , n24002 , n24003 , n24004 , n24005 , n24006 , n24007 , n24008 , n24009 , n24010 , n24011 , n24012 , n24013 , n24014 , n24015 , n24016 , n24017 , n24018 , n24019 , n24020 , n24021 , n24022 , n24023 , n24024 , n24025 , n24026 , n24027 , n24028 , n24029 , n24030 , n24031 , n24032 , n24033 , n24034 , n24035 , n24036 , n24037 , n24038 , n24039 , n24040 , n24041 , n24042 , n24043 , n24044 , n24045 , n24046 , n24047 , n24048 , n24049 , n24050 , n24051 , n24052 , n24053 , n24054 , n24055 , n24056 , n24057 , n24058 , n24059 , n24060 , n24061 , n24062 , n24063 , n24064 , n24065 , n24066 , n24067 , n24068 , n24069 , n24070 , n24071 , n24072 , n24073 , n24074 , n24075 , n24076 , n24077 , n24078 , n24079 , n24080 , n24081 , n24082 , n24083 , n24084 , n24085 , n24086 , n24087 , n24088 , n24089 , n24090 , n24091 , n24092 , n24093 , n24094 , n24095 , n24096 , n24097 , n24098 , n24099 , n24100 , n24101 , n24102 , n24103 , n24104 , n24105 , n24106 , n24107 , n24108 , n24109 , n24110 , n24111 , n24112 , n24113 , n24114 , n24115 , n24116 , n24117 , n24118 , n24119 , n24120 , n24121 , n24122 , n24123 , n24124 , n24125 , n24126 , n24127 , n24128 , n24129 , n24130 , n24131 , n24132 , n24133 , n24134 , n24135 , n24136 , n24137 , n24138 , n24139 , n24140 , n24141 , n24142 , n24143 , n24144 , n24145 , n24146 , n24147 , n24148 , n24149 , n24150 , n24151 , n24152 , n24153 , n24154 , n24155 , n24156 , n24157 , n24158 , n24159 , n24160 , n24161 , n24162 , n24163 , n24164 , n24165 , n24166 , n24167 , n24168 , n24169 , n24170 , n24171 , n24172 , n24173 , n24174 , n24175 , n24176 , n24177 , n24178 , n24179 , n24180 , n24181 , n24182 , n24183 , n24184 , n24185 , n24186 , n24187 , n24188 , n24189 , n24190 , n24191 , n24192 , n24193 , n24194 , n24195 , n24196 , n24197 , n24198 , n24199 , n24200 , n24201 , n24202 , n24203 , n24204 , n24205 , n24206 , n24207 , n24208 , n24209 , n24210 , n24211 , n24212 , n24213 , n24214 , n24215 , n24216 , n24217 , n24218 , n24219 , n24220 , n24221 , n24222 , n24223 , n24224 , n24225 , n24226 , n24227 , n24228 , n24229 , n24230 , n24231 , n24232 , n24233 , n24234 , n24235 , n24236 , n24237 , n24238 , n24239 , n24240 , n24241 , n24242 , n24243 , n24244 , n24245 , n24246 , n24247 , n24248 , n24249 , n24250 , n24251 , n24252 , n24253 , n24254 , n24255 , n24256 , n24257 , n24258 , n24259 , n24260 , n24261 , n24262 , n24263 , n24264 , n24265 , n24266 , n24267 , n24268 , n24269 , n24270 , n24271 , n24272 , n24273 , n24274 , n24275 , n24276 , n24277 , n24278 , n24279 , n24280 , n24281 , n24282 , n24283 , n24284 , n24285 , n24286 , n24287 , n24288 , n24289 , n24290 , n24291 , n24292 , n24293 , n24294 , n24295 , n24296 , n24297 , n24298 , n24299 , n24300 , n24301 , n24302 , n24303 , n24304 , n24305 , n24306 , n24307 , n24308 , n24309 , n24310 , n24311 , n24312 , n24313 , n24314 , n24315 , n24316 , n24317 , n24318 , n24319 , n24320 , n24321 , n24322 , n24323 , n24324 , n24325 , n24326 , n24327 , n24328 , n24329 , n24330 , n24331 , n24332 , n24333 , n24334 , n24335 , n24336 , n24337 , n24338 , n24339 , n24340 , n24341 , n24342 , n24343 , n24344 , n24345 , n24346 , n24347 , n24348 , n24349 , n24350 , n24351 , n24352 , n24353 , n24354 , n24355 , n24356 , n24357 , n24358 , n24359 , n24360 , n24361 , n24362 , n24363 , n24364 , n24365 , n24366 , n24367 , n24368 , n24369 , n24370 , n24371 , n24372 , n24373 , n24374 , n24375 , n24376 , n24377 , n24378 , n24379 , n24380 , n24381 , n24382 , n24383 , n24384 , n24385 , n24386 , n24387 , n24388 , n24389 , n24390 , n24391 , n24392 , n24393 , n24394 , n24395 , n24396 , n24397 , n24398 , n24399 , n24400 , n24401 , n24402 , n24403 , n24404 , n24405 , n24406 , n24407 , n24408 , n24409 , n24410 , n24411 , n24412 , n24413 , n24414 , n24415 , n24416 , n24417 , n24418 , n24419 , n24420 , n24421 , n24422 , n24423 , n24424 , n24425 , n24426 , n24427 , n24428 , n24429 , n24430 , n24431 , n24432 , n24433 , n24434 , n24435 , n24436 , n24437 , n24438 , n24439 , n24440 , n24441 , n24442 , n24443 , n24444 , n24445 , n24446 , n24447 , n24448 , n24449 , n24450 , n24451 , n24452 , n24453 , n24454 , n24455 , n24456 , n24457 , n24458 , n24459 , n24460 , n24461 , n24462 , n24463 , n24464 , n24465 , n24466 , n24467 , n24468 , n24469 , n24470 , n24471 , n24472 , n24473 , n24474 , n24475 , n24476 , n24477 , n24478 , n24479 , n24480 , n24481 , n24482 , n24483 , n24484 , n24485 , n24486 , n24487 , n24488 , n24489 , n24490 , n24491 , n24492 , n24493 , n24494 , n24495 , n24496 , n24497 , n24498 , n24499 , n24500 , n24501 , n24502 , n24503 , n24504 , n24505 , n24506 , n24507 , n24508 , n24509 , n24510 , n24511 , n24512 , n24513 , n24514 , n24515 , n24516 , n24517 , n24518 , n24519 , n24520 , n24521 , n24522 , n24523 , n24524 , n24525 , n24526 , n24527 , n24528 , n24529 , n24530 , n24531 , n24532 , n24533 , n24534 , n24535 , n24536 , n24537 , n24538 , n24539 , n24540 , n24541 , n24542 , n24543 , n24544 , n24545 , n24546 , n24547 , n24548 , n24549 , n24550 , n24551 , n24552 , n24553 , n24554 , n24555 , n24556 , n24557 , n24558 , n24559 , n24560 , n24561 , n24562 , n24563 , n24564 , n24565 , n24566 , n24567 , n24568 , n24569 , n24570 , n24571 , n24572 , n24573 , n24574 , n24575 , n24576 , n24577 , n24578 , n24579 , n24580 , n24581 , n24582 , n24583 , n24584 , n24585 , n24586 , n24587 , n24588 , n24589 , n24590 , n24591 , n24592 , n24593 , n24594 , n24595 , n24596 , n24597 , n24598 , n24599 , n24600 , n24601 , n24602 , n24603 , n24604 , n24605 , n24606 , n24607 , n24608 , n24609 , n24610 , n24611 , n24612 , n24613 , n24614 , n24615 , n24616 , n24617 , n24618 , n24619 , n24620 , n24621 , n24622 , n24623 , n24624 , n24625 , n24626 , n24627 , n24628 , n24629 , n24630 , n24631 , n24632 , n24633 , n24634 , n24635 , n24636 , n24637 , n24638 , n24639 , n24640 , n24641 , n24642 , n24643 , n24644 , n24645 , n24646 , n24647 , n24648 , n24649 , n24650 , n24651 , n24652 , n24653 , n24654 , n24655 , n24656 , n24657 , n24658 , n24659 , n24660 , n24661 , n24662 , n24663 , n24664 , n24665 , n24666 , n24667 , n24668 , n24669 , n24670 , n24671 , n24672 , n24673 , n24674 , n24675 , n24676 , n24677 , n24678 , n24679 , n24680 , n24681 , n24682 , n24683 , n24684 , n24685 , n24686 , n24687 , n24688 , n24689 , n24690 , n24691 , n24692 , n24693 , n24694 , n24695 , n24696 , n24697 , n24698 , n24699 , n24700 , n24701 , n24702 , n24703 , n24704 , n24705 , n24706 , n24707 , n24708 , n24709 , n24710 , n24711 , n24712 , n24713 , n24714 , n24715 , n24716 , n24717 , n24718 , n24719 , n24720 , n24721 , n24722 , n24723 , n24724 , n24725 , n24726 , n24727 , n24728 , n24729 , n24730 , n24731 , n24732 , n24733 , n24734 , n24735 , n24736 , n24737 , n24738 , n24739 , n24740 , n24741 , n24742 , n24743 , n24744 , n24745 , n24746 , n24747 , n24748 , n24749 , n24750 , n24751 , n24752 , n24753 , n24754 , n24755 , n24756 , n24757 , n24758 , n24759 , n24760 , n24761 , n24762 , n24763 , n24764 , n24765 , n24766 , n24767 , n24768 , n24769 , n24770 , n24771 , n24772 , n24773 , n24774 , n24775 , n24776 , n24777 , n24778 , n24779 , n24780 , n24781 , n24782 , n24783 , n24784 , n24785 , n24786 , n24787 , n24788 , n24789 , n24790 , n24791 , n24792 , n24793 , n24794 , n24795 , n24796 , n24797 , n24798 , n24799 , n24800 , n24801 , n24802 , n24803 , n24804 , n24805 , n24806 , n24807 , n24808 , n24809 , n24810 , n24811 , n24812 , n24813 , n24814 , n24815 , n24816 , n24817 , n24818 , n24819 , n24820 , n24821 , n24822 , n24823 , n24824 , n24825 , n24826 , n24827 , n24828 , n24829 , n24830 , n24831 , n24832 , n24833 , n24834 , n24835 , n24836 , n24837 , n24838 , n24839 , n24840 , n24841 , n24842 , n24843 , n24844 , n24845 , n24846 , n24847 , n24848 , n24849 , n24850 , n24851 , n24852 , n24853 , n24854 , n24855 , n24856 , n24857 , n24858 , n24859 , n24860 , n24861 , n24862 , n24863 , n24864 , n24865 , n24866 , n24867 , n24868 , n24869 , n24870 , n24871 , n24872 , n24873 , n24874 , n24875 , n24876 , n24877 , n24878 , n24879 , n24880 , n24881 , n24882 , n24883 , n24884 , n24885 , n24886 , n24887 , n24888 , n24889 , n24890 , n24891 , n24892 , n24893 , n24894 , n24895 , n24896 , n24897 , n24898 , n24899 , n24900 , n24901 , n24902 , n24903 , n24904 , n24905 , n24906 , n24907 , n24908 , n24909 , n24910 , n24911 , n24912 , n24913 , n24914 , n24915 , n24916 , n24917 , n24918 , n24919 , n24920 , n24921 , n24922 , n24923 , n24924 , n24925 , n24926 , n24927 , n24928 , n24929 , n24930 , n24931 , n24932 , n24933 , n24934 , n24935 , n24936 , n24937 , n24938 , n24939 , n24940 , n24941 , n24942 , n24943 , n24944 , n24945 , n24946 , n24947 , n24948 , n24949 , n24950 , n24951 , n24952 , n24953 , n24954 , n24955 , n24956 , n24957 , n24958 , n24959 , n24960 , n24961 , n24962 , n24963 , n24964 , n24965 , n24966 , n24967 , n24968 , n24969 , n24970 , n24971 , n24972 , n24973 , n24974 , n24975 , n24976 , n24977 , n24978 , n24979 , n24980 , n24981 , n24982 , n24983 , n24984 , n24985 , n24986 , n24987 , n24988 , n24989 , n24990 , n24991 , n24992 , n24993 , n24994 , n24995 , n24996 , n24997 , n24998 , n24999 , n25000 , n25001 , n25002 , n25003 , n25004 , n25005 , n25006 , n25007 , n25008 , n25009 , n25010 , n25011 , n25012 , n25013 , n25014 , n25015 , n25016 , n25017 , n25018 , n25019 , n25020 , n25021 , n25022 , n25023 , n25024 , n25025 , n25026 , n25027 , n25028 , n25029 , n25030 , n25031 , n25032 , n25033 , n25034 , n25035 , n25036 , n25037 , n25038 , n25039 , n25040 , n25041 , n25042 , n25043 , n25044 , n25045 , n25046 , n25047 , n25048 , n25049 , n25050 , n25051 , n25052 , n25053 , n25054 , n25055 , n25056 , n25057 , n25058 , n25059 , n25060 , n25061 , n25062 , n25063 , n25064 , n25065 , n25066 , n25067 , n25068 , n25069 , n25070 , n25071 , n25072 , n25073 , n25074 , n25075 , n25076 , n25077 , n25078 , n25079 , n25080 , n25081 , n25082 , n25083 , n25084 , n25085 , n25086 , n25087 , n25088 , n25089 , n25090 , n25091 , n25092 , n25093 , n25094 , n25095 , n25096 , n25097 , n25098 , n25099 , n25100 , n25101 , n25102 , n25103 , n25104 , n25105 , n25106 , n25107 , n25108 , n25109 , n25110 , n25111 , n25112 , n25113 , n25114 , n25115 , n25116 , n25117 , n25118 , n25119 , n25120 , n25121 , n25122 , n25123 , n25124 , n25125 , n25126 , n25127 , n25128 , n25129 , n25130 , n25131 , n25132 , n25133 , n25134 , n25135 , n25136 , n25137 , n25138 , n25139 , n25140 , n25141 , n25142 , n25143 , n25144 , n25145 , n25146 , n25147 , n25148 , n25149 , n25150 , n25151 , n25152 , n25153 , n25154 , n25155 , n25156 , n25157 , n25158 , n25159 , n25160 , n25161 , n25162 , n25163 , n25164 , n25165 , n25166 , n25167 , n25168 , n25169 , n25170 , n25171 , n25172 , n25173 , n25174 , n25175 , n25176 , n25177 , n25178 , n25179 , n25180 , n25181 , n25182 , n25183 , n25184 , n25185 , n25186 , n25187 , n25188 , n25189 , n25190 , n25191 , n25192 , n25193 , n25194 , n25195 , n25196 , n25197 , n25198 , n25199 , n25200 , n25201 , n25202 , n25203 , n25204 , n25205 , n25206 , n25207 , n25208 , n25209 , n25210 , n25211 , n25212 , n25213 , n25214 , n25215 , n25216 , n25217 , n25218 , n25219 , n25220 , n25221 , n25222 , n25223 , n25224 , n25225 , n25226 , n25227 , n25228 , n25229 , n25230 , n25231 , n25232 , n25233 , n25234 , n25235 , n25236 , n25237 , n25238 , n25239 , n25240 , n25241 , n25242 , n25243 , n25244 , n25245 , n25246 , n25247 , n25248 , n25249 , n25250 , n25251 , n25252 , n25253 , n25254 , n25255 , n25256 , n25257 , n25258 , n25259 , n25260 , n25261 , n25262 , n25263 , n25264 , n25265 , n25266 , n25267 , n25268 , n25269 , n25270 , n25271 , n25272 , n25273 , n25274 , n25275 , n25276 , n25277 , n25278 , n25279 , n25280 , n25281 , n25282 , n25283 , n25284 , n25285 , n25286 , n25287 , n25288 , n25289 , n25290 , n25291 , n25292 , n25293 , n25294 , n25295 , n25296 , n25297 , n25298 , n25299 , n25300 , n25301 , n25302 , n25303 , n25304 , n25305 , n25306 , n25307 , n25308 , n25309 , n25310 , n25311 , n25312 , n25313 , n25314 , n25315 , n25316 , n25317 , n25318 , n25319 , n25320 , n25321 , n25322 , n25323 , n25324 , n25325 , n25326 , n25327 , n25328 , n25329 , n25330 , n25331 , n25332 , n25333 , n25334 , n25335 , n25336 , n25337 , n25338 , n25339 , n25340 , n25341 , n25342 , n25343 , n25344 , n25345 , n25346 , n25347 , n25348 , n25349 , n25350 , n25351 , n25352 , n25353 , n25354 , n25355 , n25356 , n25357 , n25358 , n25359 , n25360 , n25361 , n25362 , n25363 , n25364 , n25365 , n25366 , n25367 , n25368 , n25369 , n25370 , n25371 , n25372 , n25373 , n25374 , n25375 , n25376 , n25377 , n25378 , n25379 , n25380 , n25381 , n25382 , n25383 , n25384 , n25385 , n25386 , n25387 , n25388 , n25389 , n25390 , n25391 , n25392 , n25393 , n25394 , n25395 , n25396 , n25397 , n25398 , n25399 , n25400 , n25401 , n25402 , n25403 , n25404 , n25405 , n25406 , n25407 , n25408 , n25409 , n25410 , n25411 , n25412 , n25413 , n25414 , n25415 , n25416 , n25417 , n25418 , n25419 , n25420 , n25421 , n25422 , n25423 , n25424 , n25425 , n25426 , n25427 , n25428 , n25429 , n25430 , n25431 , n25432 , n25433 , n25434 , n25435 , n25436 , n25437 , n25438 , n25439 , n25440 , n25441 , n25442 , n25443 , n25444 , n25445 , n25446 , n25447 , n25448 , n25449 , n25450 , n25451 , n25452 , n25453 , n25454 , n25455 , n25456 , n25457 , n25458 , n25459 , n25460 , n25461 , n25462 , n25463 , n25464 , n25465 , n25466 , n25467 , n25468 , n25469 , n25470 , n25471 , n25472 , n25473 , n25474 , n25475 , n25476 , n25477 , n25478 , n25479 , n25480 , n25481 , n25482 , n25483 , n25484 , n25485 , n25486 , n25487 , n25488 , n25489 , n25490 , n25491 , n25492 , n25493 , n25494 , n25495 , n25496 , n25497 , n25498 , n25499 , n25500 , n25501 , n25502 , n25503 , n25504 , n25505 , n25506 , n25507 , n25508 , n25509 , n25510 , n25511 , n25512 , n25513 , n25514 , n25515 , n25516 , n25517 , n25518 , n25519 , n25520 , n25521 , n25522 , n25523 , n25524 , n25525 , n25526 , n25527 , n25528 , n25529 , n25530 , n25531 , n25532 , n25533 , n25534 , n25535 , n25536 , n25537 , n25538 , n25539 , n25540 , n25541 , n25542 , n25543 , n25544 , n25545 , n25546 , n25547 , n25548 , n25549 , n25550 , n25551 , n25552 , n25553 , n25554 , n25555 , n25556 , n25557 , n25558 , n25559 , n25560 , n25561 , n25562 , n25563 , n25564 , n25565 , n25566 , n25567 , n25568 , n25569 , n25570 , n25571 , n25572 , n25573 , n25574 , n25575 , n25576 , n25577 , n25578 , n25579 , n25580 , n25581 , n25582 , n25583 , n25584 , n25585 , n25586 , n25587 , n25588 , n25589 , n25590 , n25591 , n25592 , n25593 , n25594 , n25595 , n25596 , n25597 , n25598 , n25599 , n25600 , n25601 , n25602 , n25603 , n25604 , n25605 , n25606 , n25607 , n25608 , n25609 , n25610 , n25611 , n25612 , n25613 , n25614 , n25615 , n25616 , n25617 , n25618 , n25619 , n25620 , n25621 , n25622 , n25623 , n25624 , n25625 , n25626 , n25627 , n25628 , n25629 , n25630 , n25631 , n25632 , n25633 , n25634 , n25635 , n25636 , n25637 , n25638 , n25639 , n25640 , n25641 , n25642 , n25643 , n25644 , n25645 , n25646 , n25647 , n25648 , n25649 , n25650 , n25651 , n25652 , n25653 , n25654 , n25655 , n25656 , n25657 , n25658 , n25659 , n25660 , n25661 , n25662 , n25663 , n25664 , n25665 , n25666 , n25667 , n25668 , n25669 , n25670 , n25671 , n25672 , n25673 , n25674 , n25675 , n25676 , n25677 , n25678 , n25679 , n25680 , n25681 , n25682 , n25683 , n25684 , n25685 , n25686 , n25687 , n25688 , n25689 , n25690 , n25691 , n25692 , n25693 , n25694 , n25695 , n25696 , n25697 , n25698 , n25699 , n25700 , n25701 , n25702 , n25703 , n25704 , n25705 , n25706 , n25707 , n25708 , n25709 , n25710 , n25711 , n25712 , n25713 , n25714 , n25715 , n25716 , n25717 , n25718 , n25719 , n25720 , n25721 , n25722 , n25723 , n25724 , n25725 , n25726 , n25727 , n25728 , n25729 , n25730 , n25731 , n25732 , n25733 , n25734 , n25735 , n25736 , n25737 , n25738 , n25739 , n25740 , n25741 , n25742 , n25743 , n25744 , n25745 , n25746 , n25747 , n25748 , n25749 , n25750 , n25751 , n25752 , n25753 , n25754 , n25755 , n25756 , n25757 , n25758 , n25759 , n25760 , n25761 , n25762 , n25763 , n25764 , n25765 , n25766 , n25767 , n25768 , n25769 , n25770 , n25771 , n25772 , n25773 , n25774 , n25775 , n25776 , n25777 , n25778 , n25779 , n25780 , n25781 , n25782 , n25783 , n25784 , n25785 , n25786 , n25787 , n25788 , n25789 , n25790 , n25791 , n25792 , n25793 , n25794 , n25795 , n25796 , n25797 , n25798 , n25799 , n25800 , n25801 , n25802 , n25803 , n25804 , n25805 , n25806 , n25807 , n25808 , n25809 , n25810 , n25811 , n25812 , n25813 , n25814 , n25815 , n25816 , n25817 , n25818 , n25819 , n25820 , n25821 , n25822 , n25823 , n25824 , n25825 , n25826 , n25827 , n25828 , n25829 , n25830 , n25831 , n25832 , n25833 , n25834 , n25835 , n25836 , n25837 , n25838 , n25839 , n25840 , n25841 , n25842 , n25843 , n25844 , n25845 , n25846 , n25847 , n25848 , n25849 , n25850 , n25851 , n25852 , n25853 , n25854 , n25855 , n25856 , n25857 , n25858 , n25859 , n25860 , n25861 , n25862 , n25863 , n25864 , n25865 , n25866 , n25867 , n25868 , n25869 , n25870 , n25871 , n25872 , n25873 , n25874 , n25875 , n25876 , n25877 , n25878 , n25879 , n25880 , n25881 , n25882 , n25883 , n25884 , n25885 , n25886 , n25887 , n25888 , n25889 , n25890 , n25891 , n25892 , n25893 , n25894 , n25895 , n25896 , n25897 , n25898 , n25899 , n25900 , n25901 , n25902 , n25903 , n25904 , n25905 , n25906 , n25907 , n25908 , n25909 , n25910 , n25911 , n25912 , n25913 , n25914 , n25915 , n25916 , n25917 , n25918 , n25919 , n25920 , n25921 , n25922 , n25923 , n25924 , n25925 , n25926 , n25927 , n25928 , n25929 , n25930 , n25931 , n25932 , n25933 , n25934 , n25935 , n25936 , n25937 , n25938 , n25939 , n25940 , n25941 , n25942 , n25943 , n25944 , n25945 , n25946 , n25947 , n25948 , n25949 , n25950 , n25951 , n25952 , n25953 , n25954 , n25955 , n25956 , n25957 , n25958 , n25959 , n25960 , n25961 , n25962 , n25963 , n25964 , n25965 , n25966 , n25967 , n25968 , n25969 , n25970 , n25971 , n25972 , n25973 , n25974 , n25975 , n25976 , n25977 , n25978 , n25979 , n25980 , n25981 , n25982 , n25983 , n25984 , n25985 , n25986 , n25987 , n25988 , n25989 , n25990 , n25991 , n25992 , n25993 , n25994 , n25995 , n25996 , n25997 , n25998 , n25999 , n26000 , n26001 , n26002 , n26003 , n26004 , n26005 , n26006 , n26007 , n26008 , n26009 , n26010 , n26011 , n26012 , n26013 , n26014 , n26015 , n26016 , n26017 , n26018 , n26019 , n26020 , n26021 , n26022 , n26023 , n26024 , n26025 , n26026 , n26027 , n26028 , n26029 , n26030 , n26031 , n26032 , n26033 , n26034 , n26035 , n26036 , n26037 , n26038 , n26039 , n26040 , n26041 , n26042 , n26043 , n26044 , n26045 , n26046 , n26047 , n26048 , n26049 , n26050 , n26051 , n26052 , n26053 , n26054 , n26055 , n26056 , n26057 , n26058 , n26059 , n26060 , n26061 , n26062 , n26063 , n26064 , n26065 , n26066 , n26067 , n26068 , n26069 , n26070 , n26071 , n26072 , n26073 , n26074 , n26075 , n26076 , n26077 , n26078 , n26079 , n26080 , n26081 , n26082 , n26083 , n26084 , n26085 , n26086 , n26087 , n26088 , n26089 , n26090 , n26091 , n26092 , n26093 , n26094 , n26095 , n26096 , n26097 , n26098 , n26099 , n26100 , n26101 , n26102 , n26103 , n26104 , n26105 , n26106 , n26107 , n26108 , n26109 , n26110 , n26111 , n26112 , n26113 , n26114 , n26115 , n26116 , n26117 , n26118 , n26119 , n26120 , n26121 , n26122 , n26123 , n26124 , n26125 , n26126 , n26127 , n26128 , n26129 , n26130 , n26131 , n26132 , n26133 , n26134 , n26135 , n26136 , n26137 , n26138 , n26139 , n26140 , n26141 , n26142 , n26143 , n26144 , n26145 , n26146 , n26147 , n26148 , n26149 , n26150 , n26151 , n26152 , n26153 , n26154 , n26155 , n26156 , n26157 , n26158 , n26159 , n26160 , n26161 , n26162 , n26163 , n26164 , n26165 , n26166 , n26167 , n26168 , n26169 , n26170 , n26171 , n26172 , n26173 , n26174 , n26175 , n26176 , n26177 , n26178 , n26179 , n26180 , n26181 , n26182 , n26183 , n26184 , n26185 , n26186 , n26187 , n26188 , n26189 , n26190 , n26191 , n26192 , n26193 , n26194 , n26195 , n26196 , n26197 , n26198 , n26199 , n26200 , n26201 , n26202 , n26203 , n26204 , n26205 , n26206 , n26207 , n26208 , n26209 , n26210 , n26211 , n26212 , n26213 , n26214 , n26215 , n26216 , n26217 , n26218 , n26219 , n26220 , n26221 , n26222 , n26223 , n26224 , n26225 , n26226 , n26227 , n26228 , n26229 , n26230 , n26231 , n26232 , n26233 , n26234 , n26235 , n26236 , n26237 , n26238 , n26239 , n26240 , n26241 , n26242 , n26243 , n26244 , n26245 , n26246 , n26247 , n26248 , n26249 , n26250 , n26251 , n26252 , n26253 , n26254 , n26255 , n26256 , n26257 , n26258 , n26259 , n26260 , n26261 , n26262 , n26263 , n26264 , n26265 , n26266 , n26267 , n26268 , n26269 , n26270 , n26271 , n26272 , n26273 , n26274 , n26275 , n26276 , n26277 , n26278 , n26279 , n26280 , n26281 , n26282 , n26283 , n26284 , n26285 , n26286 , n26287 , n26288 , n26289 , n26290 , n26291 , n26292 , n26293 , n26294 , n26295 , n26296 , n26297 , n26298 , n26299 , n26300 , n26301 , n26302 , n26303 , n26304 , n26305 , n26306 , n26307 , n26308 , n26309 , n26310 , n26311 , n26312 , n26313 , n26314 , n26315 , n26316 , n26317 , n26318 , n26319 , n26320 , n26321 , n26322 , n26323 , n26324 , n26325 , n26326 , n26327 , n26328 , n26329 , n26330 , n26331 , n26332 , n26333 , n26334 , n26335 , n26336 , n26337 , n26338 , n26339 , n26340 , n26341 , n26342 , n26343 , n26344 , n26345 , n26346 , n26347 , n26348 , n26349 , n26350 , n26351 , n26352 , n26353 , n26354 , n26355 , n26356 , n26357 , n26358 , n26359 , n26360 , n26361 , n26362 , n26363 , n26364 , n26365 , n26366 , n26367 , n26368 , n26369 , n26370 , n26371 , n26372 , n26373 , n26374 , n26375 , n26376 , n26377 , n26378 , n26379 , n26380 , n26381 , n26382 , n26383 , n26384 , n26385 , n26386 , n26387 , n26388 , n26389 , n26390 , n26391 , n26392 , n26393 , n26394 , n26395 , n26396 , n26397 , n26398 , n26399 , n26400 , n26401 , n26402 , n26403 , n26404 , n26405 , n26406 , n26407 , n26408 , n26409 , n26410 , n26411 , n26412 , n26413 , n26414 , n26415 , n26416 , n26417 , n26418 , n26419 , n26420 , n26421 , n26422 , n26423 , n26424 , n26425 , n26426 , n26427 , n26428 , n26429 , n26430 , n26431 , n26432 , n26433 , n26434 , n26435 , n26436 , n26437 , n26438 , n26439 , n26440 , n26441 , n26442 , n26443 , n26444 , n26445 , n26446 , n26447 , n26448 , n26449 , n26450 , n26451 , n26452 , n26453 , n26454 , n26455 , n26456 , n26457 , n26458 , n26459 , n26460 , n26461 , n26462 , n26463 , n26464 , n26465 , n26466 , n26467 , n26468 , n26469 , n26470 , n26471 , n26472 , n26473 , n26474 , n26475 , n26476 , n26477 , n26478 , n26479 , n26480 , n26481 , n26482 , n26483 , n26484 , n26485 , n26486 , n26487 , n26488 , n26489 , n26490 , n26491 , n26492 , n26493 , n26494 , n26495 , n26496 , n26497 , n26498 , n26499 , n26500 , n26501 , n26502 , n26503 , n26504 , n26505 , n26506 , n26507 , n26508 , n26509 , n26510 , n26511 , n26512 , n26513 , n26514 , n26515 , n26516 , n26517 , n26518 , n26519 , n26520 , n26521 , n26522 , n26523 , n26524 , n26525 , n26526 , n26527 , n26528 , n26529 , n26530 , n26531 , n26532 , n26533 , n26534 , n26535 , n26536 , n26537 , n26538 , n26539 , n26540 , n26541 , n26542 , n26543 , n26544 , n26545 , n26546 , n26547 , n26548 , n26549 , n26550 , n26551 , n26552 , n26553 , n26554 , n26555 , n26556 , n26557 , n26558 , n26559 , n26560 , n26561 , n26562 , n26563 , n26564 , n26565 , n26566 , n26567 , n26568 , n26569 , n26570 , n26571 , n26572 , n26573 , n26574 , n26575 , n26576 , n26577 , n26578 , n26579 , n26580 , n26581 , n26582 , n26583 , n26584 , n26585 , n26586 , n26587 , n26588 , n26589 , n26590 , n26591 , n26592 , n26593 , n26594 , n26595 , n26596 , n26597 , n26598 , n26599 , n26600 , n26601 , n26602 , n26603 , n26604 , n26605 , n26606 , n26607 , n26608 , n26609 , n26610 , n26611 , n26612 , n26613 , n26614 , n26615 , n26616 , n26617 , n26618 , n26619 , n26620 , n26621 , n26622 , n26623 , n26624 , n26625 , n26626 , n26627 , n26628 , n26629 , n26630 , n26631 , n26632 , n26633 , n26634 , n26635 , n26636 , n26637 , n26638 , n26639 , n26640 , n26641 , n26642 , n26643 , n26644 , n26645 , n26646 , n26647 , n26648 , n26649 , n26650 , n26651 , n26652 , n26653 , n26654 , n26655 , n26656 , n26657 , n26658 , n26659 , n26660 , n26661 , n26662 , n26663 , n26664 , n26665 , n26666 , n26667 , n26668 , n26669 , n26670 , n26671 , n26672 , n26673 , n26674 , n26675 , n26676 , n26677 , n26678 , n26679 , n26680 , n26681 , n26682 , n26683 , n26684 , n26685 , n26686 , n26687 , n26688 , n26689 , n26690 , n26691 , n26692 , n26693 , n26694 , n26695 , n26696 , n26697 , n26698 , n26699 , n26700 , n26701 , n26702 , n26703 , n26704 , n26705 , n26706 , n26707 , n26708 , n26709 , n26710 , n26711 , n26712 , n26713 , n26714 , n26715 , n26716 , n26717 , n26718 , n26719 , n26720 , n26721 , n26722 , n26723 , n26724 , n26725 , n26726 , n26727 , n26728 , n26729 , n26730 , n26731 , n26732 , n26733 , n26734 , n26735 , n26736 , n26737 , n26738 , n26739 , n26740 , n26741 , n26742 , n26743 , n26744 , n26745 , n26746 , n26747 , n26748 , n26749 , n26750 , n26751 , n26752 , n26753 , n26754 , n26755 , n26756 , n26757 , n26758 , n26759 , n26760 , n26761 , n26762 , n26763 , n26764 , n26765 , n26766 , n26767 , n26768 , n26769 , n26770 , n26771 , n26772 , n26773 , n26774 , n26775 , n26776 , n26777 , n26778 , n26779 , n26780 , n26781 , n26782 , n26783 , n26784 , n26785 , n26786 , n26787 , n26788 , n26789 , n26790 , n26791 , n26792 , n26793 , n26794 , n26795 , n26796 , n26797 , n26798 , n26799 , n26800 , n26801 , n26802 , n26803 , n26804 , n26805 , n26806 , n26807 , n26808 , n26809 , n26810 , n26811 , n26812 , n26813 , n26814 , n26815 , n26816 , n26817 , n26818 , n26819 , n26820 , n26821 , n26822 , n26823 , n26824 , n26825 , n26826 , n26827 , n26828 , n26829 , n26830 , n26831 , n26832 , n26833 , n26834 , n26835 , n26836 , n26837 , n26838 , n26839 , n26840 , n26841 , n26842 , n26843 , n26844 , n26845 , n26846 , n26847 , n26848 , n26849 , n26850 , n26851 , n26852 , n26853 , n26854 , n26855 , n26856 , n26857 , n26858 , n26859 , n26860 , n26861 , n26862 , n26863 , n26864 , n26865 , n26866 , n26867 , n26868 , n26869 , n26870 , n26871 , n26872 , n26873 , n26874 , n26875 , n26876 , n26877 , n26878 , n26879 , n26880 , n26881 , n26882 , n26883 , n26884 , n26885 , n26886 , n26887 , n26888 , n26889 , n26890 , n26891 , n26892 , n26893 , n26894 , n26895 , n26896 , n26897 , n26898 , n26899 , n26900 , n26901 , n26902 , n26903 , n26904 , n26905 , n26906 , n26907 , n26908 , n26909 , n26910 , n26911 , n26912 , n26913 , n26914 , n26915 , n26916 , n26917 , n26918 , n26919 , n26920 , n26921 , n26922 , n26923 , n26924 , n26925 , n26926 , n26927 , n26928 , n26929 , n26930 , n26931 , n26932 , n26933 , n26934 , n26935 , n26936 , n26937 , n26938 , n26939 , n26940 , n26941 , n26942 , n26943 , n26944 , n26945 , n26946 , n26947 , n26948 , n26949 , n26950 , n26951 , n26952 , n26953 , n26954 , n26955 , n26956 , n26957 , n26958 , n26959 , n26960 , n26961 , n26962 , n26963 , n26964 , n26965 , n26966 , n26967 , n26968 , n26969 , n26970 , n26971 , n26972 , n26973 , n26974 , n26975 , n26976 , n26977 , n26978 , n26979 , n26980 , n26981 , n26982 , n26983 , n26984 , n26985 , n26986 , n26987 , n26988 , n26989 , n26990 , n26991 , n26992 , n26993 , n26994 , n26995 , n26996 , n26997 , n26998 , n26999 , n27000 , n27001 , n27002 , n27003 , n27004 , n27005 , n27006 , n27007 , n27008 , n27009 , n27010 , n27011 , n27012 , n27013 , n27014 , n27015 , n27016 , n27017 , n27018 , n27019 , n27020 , n27021 , n27022 , n27023 , n27024 , n27025 , n27026 , n27027 , n27028 , n27029 , n27030 , n27031 , n27032 , n27033 , n27034 , n27035 , n27036 , n27037 , n27038 , n27039 , n27040 , n27041 , n27042 , n27043 , n27044 , n27045 , n27046 , n27047 , n27048 , n27049 , n27050 , n27051 , n27052 , n27053 , n27054 , n27055 , n27056 , n27057 , n27058 , n27059 , n27060 , n27061 , n27062 , n27063 , n27064 , n27065 , n27066 , n27067 , n27068 , n27069 , n27070 , n27071 , n27072 , n27073 , n27074 , n27075 , n27076 , n27077 , n27078 , n27079 , n27080 , n27081 , n27082 , n27083 , n27084 , n27085 , n27086 , n27087 , n27088 , n27089 , n27090 , n27091 , n27092 , n27093 , n27094 , n27095 , n27096 , n27097 , n27098 , n27099 , n27100 , n27101 , n27102 , n27103 , n27104 , n27105 , n27106 , n27107 , n27108 , n27109 , n27110 , n27111 , n27112 , n27113 , n27114 , n27115 , n27116 , n27117 , n27118 , n27119 , n27120 , n27121 , n27122 , n27123 , n27124 , n27125 , n27126 , n27127 , n27128 , n27129 , n27130 , n27131 , n27132 , n27133 , n27134 , n27135 , n27136 , n27137 , n27138 , n27139 , n27140 , n27141 , n27142 , n27143 , n27144 , n27145 , n27146 , n27147 , n27148 , n27149 , n27150 , n27151 , n27152 , n27153 , n27154 , n27155 , n27156 , n27157 , n27158 , n27159 , n27160 , n27161 , n27162 , n27163 , n27164 , n27165 , n27166 , n27167 , n27168 , n27169 , n27170 , n27171 , n27172 , n27173 , n27174 , n27175 , n27176 , n27177 , n27178 , n27179 , n27180 , n27181 , n27182 , n27183 , n27184 , n27185 , n27186 , n27187 , n27188 , n27189 , n27190 , n27191 , n27192 , n27193 , n27194 , n27195 , n27196 , n27197 , n27198 , n27199 , n27200 , n27201 , n27202 , n27203 , n27204 , n27205 , n27206 , n27207 , n27208 , n27209 , n27210 , n27211 , n27212 , n27213 , n27214 , n27215 , n27216 , n27217 , n27218 , n27219 , n27220 , n27221 , n27222 , n27223 , n27224 , n27225 , n27226 , n27227 , n27228 , n27229 , n27230 , n27231 , n27232 , n27233 , n27234 , n27235 , n27236 , n27237 , n27238 , n27239 , n27240 , n27241 , n27242 , n27243 , n27244 , n27245 , n27246 , n27247 , n27248 , n27249 , n27250 , n27251 , n27252 , n27253 , n27254 , n27255 , n27256 , n27257 , n27258 , n27259 , n27260 , n27261 , n27262 , n27263 , n27264 , n27265 , n27266 , n27267 , n27268 , n27269 , n27270 , n27271 , n27272 , n27273 , n27274 , n27275 , n27276 , n27277 , n27278 , n27279 , n27280 , n27281 , n27282 , n27283 , n27284 , n27285 , n27286 , n27287 , n27288 , n27289 , n27290 , n27291 , n27292 , n27293 , n27294 , n27295 , n27296 , n27297 , n27298 , n27299 , n27300 , n27301 , n27302 , n27303 , n27304 , n27305 , n27306 , n27307 , n27308 , n27309 , n27310 , n27311 , n27312 , n27313 , n27314 , n27315 , n27316 , n27317 , n27318 , n27319 , n27320 , n27321 , n27322 , n27323 , n27324 , n27325 , n27326 , n27327 , n27328 , n27329 , n27330 , n27331 , n27332 , n27333 , n27334 , n27335 , n27336 , n27337 , n27338 , n27339 , n27340 , n27341 , n27342 , n27343 , n27344 , n27345 , n27346 , n27347 , n27348 , n27349 , n27350 , n27351 , n27352 , n27353 , n27354 , n27355 , n27356 , n27357 , n27358 , n27359 , n27360 , n27361 , n27362 , n27363 , n27364 , n27365 , n27366 , n27367 , n27368 , n27369 , n27370 , n27371 , n27372 , n27373 , n27374 , n27375 , n27376 , n27377 , n27378 , n27379 , n27380 , n27381 , n27382 , n27383 , n27384 , n27385 , n27386 , n27387 , n27388 , n27389 , n27390 , n27391 , n27392 , n27393 , n27394 , n27395 , n27396 , n27397 , n27398 , n27399 , n27400 , n27401 , n27402 , n27403 , n27404 , n27405 , n27406 , n27407 , n27408 , n27409 , n27410 , n27411 , n27412 , n27413 , n27414 , n27415 , n27416 , n27417 , n27418 , n27419 , n27420 , n27421 , n27422 , n27423 , n27424 , n27425 , n27426 , n27427 , n27428 , n27429 , n27430 , n27431 , n27432 , n27433 , n27434 , n27435 , n27436 , n27437 , n27438 , n27439 , n27440 , n27441 , n27442 , n27443 , n27444 , n27445 , n27446 , n27447 , n27448 , n27449 , n27450 , n27451 , n27452 , n27453 , n27454 , n27455 , n27456 , n27457 , n27458 , n27459 , n27460 , n27461 , n27462 , n27463 , n27464 , n27465 , n27466 , n27467 , n27468 , n27469 , n27470 , n27471 , n27472 , n27473 , n27474 , n27475 , n27476 , n27477 , n27478 , n27479 , n27480 , n27481 , n27482 , n27483 , n27484 , n27485 , n27486 , n27487 , n27488 , n27489 , n27490 , n27491 , n27492 , n27493 , n27494 , n27495 , n27496 , n27497 , n27498 , n27499 , n27500 , n27501 , n27502 , n27503 , n27504 , n27505 , n27506 , n27507 , n27508 , n27509 , n27510 , n27511 , n27512 , n27513 , n27514 , n27515 , n27516 , n27517 , n27518 , n27519 , n27520 , n27521 , n27522 , n27523 , n27524 , n27525 , n27526 , n27527 , n27528 , n27529 , n27530 , n27531 , n27532 , n27533 , n27534 , n27535 , n27536 , n27537 , n27538 , n27539 , n27540 , n27541 , n27542 , n27543 , n27544 , n27545 , n27546 , n27547 , n27548 , n27549 , n27550 , n27551 , n27552 , n27553 , n27554 , n27555 , n27556 , n27557 , n27558 , n27559 , n27560 , n27561 , n27562 , n27563 , n27564 , n27565 , n27566 , n27567 , n27568 , n27569 , n27570 , n27571 , n27572 , n27573 , n27574 , n27575 , n27576 , n27577 , n27578 , n27579 , n27580 , n27581 , n27582 , n27583 , n27584 , n27585 , n27586 , n27587 , n27588 , n27589 , n27590 , n27591 , n27592 , n27593 , n27594 , n27595 , n27596 , n27597 , n27598 , n27599 , n27600 , n27601 , n27602 , n27603 , n27604 , n27605 , n27606 , n27607 , n27608 , n27609 , n27610 , n27611 , n27612 , n27613 , n27614 , n27615 , n27616 , n27617 , n27618 , n27619 , n27620 , n27621 , n27622 , n27623 , n27624 , n27625 , n27626 , n27627 , n27628 , n27629 , n27630 , n27631 , n27632 , n27633 , n27634 , n27635 , n27636 , n27637 , n27638 , n27639 , n27640 , n27641 , n27642 , n27643 , n27644 , n27645 , n27646 , n27647 , n27648 , n27649 , n27650 , n27651 , n27652 , n27653 , n27654 , n27655 , n27656 , n27657 , n27658 , n27659 , n27660 , n27661 , n27662 , n27663 , n27664 , n27665 , n27666 , n27667 , n27668 , n27669 , n27670 , n27671 , n27672 , n27673 , n27674 , n27675 , n27676 , n27677 , n27678 , n27679 , n27680 , n27681 , n27682 , n27683 , n27684 , n27685 , n27686 , n27687 , n27688 , n27689 , n27690 , n27691 , n27692 , n27693 , n27694 , n27695 , n27696 , n27697 , n27698 , n27699 , n27700 , n27701 , n27702 , n27703 , n27704 , n27705 , n27706 , n27707 , n27708 , n27709 , n27710 , n27711 , n27712 , n27713 , n27714 , n27715 , n27716 , n27717 , n27718 , n27719 , n27720 , n27721 , n27722 , n27723 , n27724 , n27725 , n27726 , n27727 , n27728 , n27729 , n27730 , n27731 , n27732 , n27733 , n27734 , n27735 , n27736 , n27737 , n27738 , n27739 , n27740 , n27741 , n27742 , n27743 , n27744 , n27745 , n27746 , n27747 , n27748 , n27749 , n27750 , n27751 , n27752 , n27753 , n27754 , n27755 , n27756 , n27757 , n27758 , n27759 , n27760 , n27761 , n27762 , n27763 , n27764 , n27765 , n27766 , n27767 , n27768 , n27769 , n27770 , n27771 , n27772 , n27773 , n27774 , n27775 , n27776 , n27777 , n27778 , n27779 , n27780 , n27781 , n27782 , n27783 , n27784 , n27785 , n27786 , n27787 , n27788 , n27789 , n27790 , n27791 , n27792 , n27793 , n27794 , n27795 , n27796 , n27797 , n27798 , n27799 , n27800 , n27801 , n27802 , n27803 , n27804 , n27805 , n27806 , n27807 , n27808 , n27809 , n27810 , n27811 , n27812 , n27813 , n27814 , n27815 , n27816 , n27817 , n27818 , n27819 , n27820 , n27821 , n27822 , n27823 , n27824 , n27825 , n27826 , n27827 , n27828 , n27829 , n27830 , n27831 , n27832 , n27833 , n27834 , n27835 , n27836 , n27837 , n27838 , n27839 , n27840 , n27841 , n27842 , n27843 , n27844 , n27845 , n27846 , n27847 , n27848 , n27849 , n27850 , n27851 , n27852 , n27853 , n27854 , n27855 , n27856 , n27857 , n27858 , n27859 , n27860 , n27861 , n27862 , n27863 , n27864 , n27865 , n27866 , n27867 , n27868 , n27869 , n27870 , n27871 , n27872 , n27873 , n27874 , n27875 , n27876 , n27877 , n27878 , n27879 , n27880 , n27881 , n27882 , n27883 , n27884 , n27885 , n27886 , n27887 , n27888 , n27889 , n27890 , n27891 , n27892 , n27893 , n27894 , n27895 , n27896 , n27897 , n27898 , n27899 , n27900 , n27901 , n27902 , n27903 , n27904 , n27905 , n27906 , n27907 , n27908 , n27909 , n27910 , n27911 , n27912 , n27913 , n27914 , n27915 , n27916 , n27917 , n27918 , n27919 , n27920 , n27921 , n27922 , n27923 , n27924 , n27925 , n27926 , n27927 , n27928 , n27929 , n27930 , n27931 , n27932 , n27933 , n27934 , n27935 , n27936 , n27937 , n27938 , n27939 , n27940 , n27941 , n27942 , n27943 , n27944 , n27945 , n27946 , n27947 , n27948 , n27949 , n27950 , n27951 , n27952 , n27953 , n27954 , n27955 , n27956 , n27957 , n27958 , n27959 , n27960 , n27961 , n27962 , n27963 , n27964 , n27965 , n27966 , n27967 , n27968 , n27969 , n27970 , n27971 , n27972 , n27973 , n27974 , n27975 , n27976 , n27977 , n27978 , n27979 , n27980 , n27981 , n27982 , n27983 , n27984 , n27985 , n27986 , n27987 , n27988 , n27989 , n27990 , n27991 , n27992 , n27993 , n27994 , n27995 , n27996 , n27997 , n27998 , n27999 , n28000 , n28001 , n28002 , n28003 , n28004 , n28005 , n28006 , n28007 , n28008 , n28009 , n28010 , n28011 , n28012 , n28013 , n28014 , n28015 , n28016 , n28017 , n28018 , n28019 , n28020 , n28021 , n28022 , n28023 , n28024 , n28025 , n28026 , n28027 , n28028 , n28029 , n28030 , n28031 , n28032 , n28033 , n28034 , n28035 , n28036 , n28037 , n28038 , n28039 , n28040 , n28041 , n28042 , n28043 , n28044 , n28045 , n28046 , n28047 , n28048 , n28049 , n28050 , n28051 , n28052 , n28053 , n28054 , n28055 , n28056 , n28057 , n28058 , n28059 , n28060 , n28061 , n28062 , n28063 , n28064 , n28065 , n28066 , n28067 , n28068 , n28069 , n28070 , n28071 , n28072 , n28073 , n28074 , n28075 , n28076 , n28077 , n28078 , n28079 , n28080 , n28081 , n28082 , n28083 , n28084 , n28085 , n28086 , n28087 , n28088 , n28089 , n28090 , n28091 , n28092 , n28093 , n28094 , n28095 , n28096 , n28097 , n28098 , n28099 , n28100 , n28101 , n28102 , n28103 , n28104 , n28105 , n28106 , n28107 , n28108 , n28109 , n28110 , n28111 , n28112 , n28113 , n28114 , n28115 , n28116 , n28117 , n28118 , n28119 , n28120 , n28121 , n28122 , n28123 , n28124 , n28125 , n28126 , n28127 , n28128 , n28129 , n28130 , n28131 , n28132 , n28133 , n28134 , n28135 , n28136 , n28137 , n28138 , n28139 , n28140 , n28141 , n28142 , n28143 , n28144 , n28145 , n28146 , n28147 , n28148 , n28149 , n28150 , n28151 , n28152 , n28153 , n28154 , n28155 , n28156 , n28157 , n28158 , n28159 , n28160 , n28161 , n28162 , n28163 , n28164 , n28165 , n28166 , n28167 , n28168 , n28169 , n28170 , n28171 , n28172 , n28173 , n28174 , n28175 , n28176 , n28177 , n28178 , n28179 , n28180 , n28181 , n28182 , n28183 , n28184 , n28185 , n28186 , n28187 , n28188 , n28189 , n28190 , n28191 , n28192 , n28193 , n28194 , n28195 , n28196 , n28197 , n28198 , n28199 , n28200 , n28201 , n28202 , n28203 , n28204 , n28205 , n28206 , n28207 , n28208 , n28209 , n28210 , n28211 , n28212 , n28213 , n28214 , n28215 , n28216 , n28217 , n28218 , n28219 , n28220 , n28221 , n28222 , n28223 , n28224 , n28225 , n28226 , n28227 , n28228 , n28229 , n28230 , n28231 , n28232 , n28233 , n28234 , n28235 , n28236 , n28237 , n28238 , n28239 , n28240 , n28241 , n28242 , n28243 , n28244 , n28245 , n28246 , n28247 , n28248 , n28249 , n28250 , n28251 , n28252 , n28253 , n28254 , n28255 , n28256 , n28257 , n28258 , n28259 , n28260 , n28261 , n28262 , n28263 , n28264 , n28265 , n28266 , n28267 , n28268 , n28269 , n28270 , n28271 , n28272 , n28273 , n28274 , n28275 , n28276 , n28277 , n28278 , n28279 , n28280 , n28281 , n28282 , n28283 , n28284 , n28285 , n28286 , n28287 , n28288 , n28289 , n28290 , n28291 , n28292 , n28293 , n28294 , n28295 , n28296 , n28297 , n28298 , n28299 , n28300 , n28301 , n28302 , n28303 , n28304 , n28305 , n28306 , n28307 , n28308 , n28309 , n28310 , n28311 , n28312 , n28313 , n28314 , n28315 , n28316 , n28317 , n28318 , n28319 , n28320 , n28321 , n28322 , n28323 , n28324 , n28325 , n28326 , n28327 , n28328 , n28329 , n28330 , n28331 , n28332 , n28333 , n28334 , n28335 , n28336 , n28337 , n28338 , n28339 , n28340 , n28341 , n28342 , n28343 , n28344 , n28345 , n28346 , n28347 , n28348 , n28349 , n28350 , n28351 , n28352 , n28353 , n28354 , n28355 , n28356 , n28357 , n28358 , n28359 , n28360 , n28361 , n28362 , n28363 , n28364 , n28365 , n28366 , n28367 , n28368 , n28369 , n28370 , n28371 , n28372 , n28373 , n28374 , n28375 , n28376 , n28377 , n28378 , n28379 , n28380 , n28381 , n28382 , n28383 , n28384 , n28385 , n28386 , n28387 , n28388 , n28389 , n28390 , n28391 , n28392 , n28393 , n28394 , n28395 , n28396 , n28397 , n28398 , n28399 , n28400 , n28401 , n28402 , n28403 , n28404 , n28405 , n28406 , n28407 , n28408 , n28409 , n28410 , n28411 , n28412 , n28413 , n28414 , n28415 , n28416 , n28417 , n28418 , n28419 , n28420 , n28421 , n28422 , n28423 , n28424 , n28425 , n28426 , n28427 , n28428 , n28429 , n28430 , n28431 , n28432 , n28433 , n28434 , n28435 , n28436 , n28437 , n28438 , n28439 , n28440 , n28441 , n28442 , n28443 , n28444 , n28445 , n28446 , n28447 , n28448 , n28449 , n28450 , n28451 , n28452 , n28453 , n28454 , n28455 , n28456 , n28457 , n28458 , n28459 , n28460 , n28461 , n28462 , n28463 , n28464 , n28465 , n28466 , n28467 , n28468 , n28469 , n28470 , n28471 , n28472 , n28473 , n28474 , n28475 , n28476 , n28477 , n28478 , n28479 , n28480 , n28481 , n28482 , n28483 , n28484 , n28485 , n28486 , n28487 , n28488 , n28489 , n28490 , n28491 , n28492 , n28493 , n28494 , n28495 , n28496 , n28497 , n28498 , n28499 , n28500 , n28501 , n28502 , n28503 , n28504 , n28505 , n28506 , n28507 , n28508 , n28509 , n28510 , n28511 , n28512 , n28513 , n28514 , n28515 , n28516 , n28517 , n28518 , n28519 , n28520 , n28521 , n28522 , n28523 , n28524 , n28525 , n28526 , n28527 , n28528 , n28529 , n28530 , n28531 , n28532 , n28533 , n28534 , n28535 , n28536 , n28537 , n28538 , n28539 , n28540 , n28541 , n28542 , n28543 , n28544 , n28545 , n28546 , n28547 , n28548 , n28549 , n28550 , n28551 , n28552 , n28553 , n28554 , n28555 , n28556 , n28557 , n28558 , n28559 , n28560 , n28561 , n28562 , n28563 , n28564 , n28565 , n28566 , n28567 , n28568 , n28569 , n28570 , n28571 , n28572 , n28573 , n28574 , n28575 , n28576 , n28577 , n28578 , n28579 , n28580 , n28581 , n28582 , n28583 , n28584 , n28585 , n28586 , n28587 , n28588 , n28589 , n28590 , n28591 , n28592 , n28593 , n28594 , n28595 , n28596 , n28597 , n28598 , n28599 , n28600 , n28601 , n28602 , n28603 , n28604 , n28605 , n28606 , n28607 , n28608 , n28609 , n28610 , n28611 , n28612 , n28613 , n28614 , n28615 , n28616 , n28617 , n28618 , n28619 , n28620 , n28621 , n28622 , n28623 , n28624 , n28625 , n28626 , n28627 , n28628 , n28629 , n28630 , n28631 , n28632 , n28633 , n28634 , n28635 , n28636 , n28637 , n28638 , n28639 , n28640 , n28641 , n28642 , n28643 , n28644 , n28645 , n28646 , n28647 , n28648 , n28649 , n28650 , n28651 , n28652 , n28653 , n28654 , n28655 , n28656 , n28657 , n28658 , n28659 , n28660 , n28661 , n28662 , n28663 , n28664 , n28665 , n28666 , n28667 , n28668 , n28669 , n28670 , n28671 , n28672 , n28673 , n28674 , n28675 , n28676 , n28677 , n28678 , n28679 , n28680 , n28681 , n28682 , n28683 , n28684 , n28685 , n28686 , n28687 , n28688 , n28689 , n28690 , n28691 , n28692 , n28693 , n28694 , n28695 , n28696 , n28697 , n28698 , n28699 , n28700 , n28701 , n28702 , n28703 , n28704 , n28705 , n28706 , n28707 , n28708 , n28709 , n28710 , n28711 , n28712 , n28713 , n28714 , n28715 , n28716 , n28717 , n28718 , n28719 , n28720 , n28721 , n28722 , n28723 , n28724 , n28725 , n28726 , n28727 , n28728 , n28729 , n28730 , n28731 , n28732 , n28733 , n28734 , n28735 , n28736 , n28737 , n28738 , n28739 , n28740 , n28741 , n28742 , n28743 , n28744 , n28745 , n28746 , n28747 , n28748 , n28749 , n28750 , n28751 , n28752 , n28753 , n28754 , n28755 , n28756 , n28757 , n28758 , n28759 , n28760 , n28761 , n28762 , n28763 , n28764 , n28765 , n28766 , n28767 , n28768 , n28769 , n28770 , n28771 , n28772 , n28773 , n28774 , n28775 , n28776 , n28777 , n28778 , n28779 , n28780 , n28781 , n28782 , n28783 , n28784 , n28785 , n28786 , n28787 , n28788 , n28789 , n28790 , n28791 , n28792 , n28793 , n28794 , n28795 , n28796 , n28797 , n28798 , n28799 , n28800 , n28801 , n28802 , n28803 , n28804 , n28805 , n28806 , n28807 , n28808 , n28809 , n28810 , n28811 , n28812 , n28813 , n28814 , n28815 , n28816 , n28817 , n28818 , n28819 , n28820 , n28821 , n28822 , n28823 , n28824 , n28825 , n28826 , n28827 , n28828 , n28829 , n28830 , n28831 , n28832 , n28833 , n28834 , n28835 , n28836 , n28837 , n28838 , n28839 , n28840 , n28841 , n28842 , n28843 , n28844 , n28845 , n28846 , n28847 , n28848 , n28849 , n28850 , n28851 , n28852 , n28853 , n28854 , n28855 , n28856 , n28857 , n28858 , n28859 , n28860 , n28861 , n28862 , n28863 , n28864 , n28865 , n28866 , n28867 , n28868 , n28869 , n28870 , n28871 , n28872 , n28873 , n28874 , n28875 , n28876 , n28877 , n28878 , n28879 , n28880 , n28881 , n28882 , n28883 , n28884 , n28885 , n28886 , n28887 , n28888 , n28889 , n28890 , n28891 , n28892 , n28893 , n28894 , n28895 , n28896 , n28897 , n28898 , n28899 , n28900 , n28901 , n28902 , n28903 , n28904 , n28905 , n28906 , n28907 , n28908 , n28909 , n28910 , n28911 , n28912 , n28913 , n28914 , n28915 , n28916 , n28917 , n28918 , n28919 , n28920 , n28921 , n28922 , n28923 , n28924 , n28925 , n28926 , n28927 , n28928 , n28929 , n28930 , n28931 , n28932 , n28933 , n28934 , n28935 , n28936 , n28937 , n28938 , n28939 , n28940 , n28941 , n28942 , n28943 , n28944 , n28945 , n28946 , n28947 , n28948 , n28949 , n28950 , n28951 , n28952 , n28953 , n28954 , n28955 , n28956 , n28957 , n28958 , n28959 , n28960 , n28961 , n28962 , n28963 , n28964 , n28965 , n28966 , n28967 , n28968 , n28969 , n28970 , n28971 , n28972 , n28973 , n28974 , n28975 , n28976 , n28977 , n28978 , n28979 , n28980 , n28981 , n28982 , n28983 , n28984 , n28985 , n28986 , n28987 , n28988 , n28989 , n28990 , n28991 , n28992 , n28993 , n28994 , n28995 , n28996 , n28997 , n28998 , n28999 , n29000 , n29001 , n29002 , n29003 , n29004 , n29005 , n29006 , n29007 , n29008 , n29009 , n29010 , n29011 , n29012 , n29013 , n29014 , n29015 , n29016 , n29017 , n29018 , n29019 , n29020 , n29021 , n29022 , n29023 , n29024 , n29025 , n29026 , n29027 , n29028 , n29029 , n29030 , n29031 , n29032 , n29033 , n29034 , n29035 , n29036 , n29037 , n29038 , n29039 , n29040 , n29041 , n29042 , n29043 , n29044 , n29045 , n29046 , n29047 , n29048 , n29049 , n29050 , n29051 , n29052 , n29053 , n29054 , n29055 , n29056 , n29057 , n29058 , n29059 , n29060 , n29061 , n29062 , n29063 , n29064 , n29065 , n29066 , n29067 , n29068 , n29069 , n29070 , n29071 , n29072 , n29073 , n29074 , n29075 , n29076 , n29077 , n29078 , n29079 , n29080 , n29081 , n29082 , n29083 , n29084 , n29085 , n29086 , n29087 , n29088 , n29089 , n29090 , n29091 , n29092 , n29093 , n29094 , n29095 , n29096 , n29097 , n29098 , n29099 , n29100 , n29101 , n29102 , n29103 , n29104 , n29105 , n29106 , n29107 , n29108 , n29109 , n29110 , n29111 , n29112 , n29113 , n29114 , n29115 , n29116 , n29117 , n29118 , n29119 , n29120 , n29121 , n29122 , n29123 , n29124 , n29125 , n29126 , n29127 , n29128 , n29129 , n29130 , n29131 , n29132 , n29133 , n29134 , n29135 , n29136 , n29137 , n29138 , n29139 , n29140 , n29141 , n29142 , n29143 , n29144 , n29145 , n29146 , n29147 , n29148 , n29149 , n29150 , n29151 , n29152 , n29153 , n29154 , n29155 , n29156 , n29157 , n29158 , n29159 , n29160 , n29161 , n29162 , n29163 , n29164 , n29165 , n29166 , n29167 , n29168 , n29169 , n29170 , n29171 , n29172 , n29173 , n29174 , n29175 , n29176 , n29177 , n29178 , n29179 , n29180 , n29181 , n29182 , n29183 , n29184 , n29185 , n29186 , n29187 , n29188 , n29189 , n29190 , n29191 , n29192 , n29193 , n29194 , n29195 , n29196 , n29197 , n29198 , n29199 , n29200 , n29201 , n29202 , n29203 , n29204 , n29205 , n29206 , n29207 , n29208 , n29209 , n29210 , n29211 , n29212 , n29213 , n29214 , n29215 , n29216 , n29217 , n29218 , n29219 , n29220 , n29221 , n29222 , n29223 , n29224 , n29225 , n29226 , n29227 , n29228 , n29229 , n29230 , n29231 , n29232 , n29233 , n29234 , n29235 , n29236 , n29237 , n29238 , n29239 , n29240 , n29241 , n29242 , n29243 , n29244 , n29245 , n29246 , n29247 , n29248 , n29249 , n29250 , n29251 , n29252 , n29253 , n29254 , n29255 , n29256 , n29257 , n29258 , n29259 , n29260 , n29261 , n29262 , n29263 , n29264 , n29265 , n29266 , n29267 , n29268 , n29269 , n29270 , n29271 , n29272 , n29273 , n29274 , n29275 , n29276 , n29277 , n29278 , n29279 , n29280 , n29281 , n29282 , n29283 , n29284 , n29285 , n29286 , n29287 , n29288 , n29289 , n29290 , n29291 , n29292 , n29293 , n29294 , n29295 , n29296 , n29297 , n29298 , n29299 , n29300 , n29301 , n29302 , n29303 , n29304 , n29305 , n29306 , n29307 , n29308 , n29309 , n29310 , n29311 , n29312 , n29313 , n29314 , n29315 , n29316 , n29317 , n29318 , n29319 , n29320 , n29321 , n29322 , n29323 , n29324 , n29325 , n29326 , n29327 , n29328 , n29329 , n29330 , n29331 , n29332 , n29333 , n29334 , n29335 , n29336 , n29337 , n29338 , n29339 , n29340 , n29341 , n29342 , n29343 , n29344 , n29345 , n29346 , n29347 , n29348 , n29349 , n29350 , n29351 , n29352 , n29353 , n29354 , n29355 , n29356 , n29357 , n29358 , n29359 , n29360 , n29361 , n29362 , n29363 , n29364 , n29365 , n29366 , n29367 , n29368 , n29369 , n29370 , n29371 , n29372 , n29373 , n29374 , n29375 , n29376 , n29377 , n29378 , n29379 , n29380 , n29381 , n29382 , n29383 , n29384 , n29385 , n29386 , n29387 , n29388 , n29389 , n29390 , n29391 , n29392 , n29393 , n29394 , n29395 , n29396 , n29397 , n29398 , n29399 , n29400 , n29401 , n29402 , n29403 , n29404 , n29405 , n29406 , n29407 , n29408 , n29409 , n29410 , n29411 , n29412 , n29413 , n29414 , n29415 , n29416 , n29417 , n29418 , n29419 , n29420 , n29421 , n29422 , n29423 , n29424 , n29425 , n29426 , n29427 , n29428 , n29429 , n29430 , n29431 , n29432 , n29433 , n29434 , n29435 , n29436 , n29437 , n29438 , n29439 , n29440 , n29441 , n29442 , n29443 , n29444 , n29445 , n29446 , n29447 , n29448 , n29449 , n29450 , n29451 , n29452 , n29453 , n29454 , n29455 , n29456 , n29457 , n29458 , n29459 , n29460 , n29461 , n29462 , n29463 , n29464 , n29465 , n29466 , n29467 , n29468 , n29469 , n29470 , n29471 , n29472 , n29473 , n29474 , n29475 , n29476 , n29477 , n29478 , n29479 , n29480 , n29481 , n29482 , n29483 , n29484 , n29485 , n29486 , n29487 , n29488 , n29489 , n29490 , n29491 , n29492 , n29493 , n29494 , n29495 , n29496 , n29497 , n29498 , n29499 , n29500 , n29501 , n29502 , n29503 , n29504 , n29505 , n29506 , n29507 , n29508 , n29509 , n29510 , n29511 , n29512 , n29513 , n29514 , n29515 , n29516 , n29517 , n29518 , n29519 , n29520 , n29521 , n29522 , n29523 , n29524 , n29525 , n29526 , n29527 , n29528 , n29529 , n29530 , n29531 , n29532 , n29533 , n29534 , n29535 , n29536 , n29537 , n29538 , n29539 , n29540 , n29541 , n29542 , n29543 , n29544 , n29545 , n29546 , n29547 , n29548 , n29549 , n29550 , n29551 , n29552 , n29553 , n29554 , n29555 , n29556 , n29557 , n29558 , n29559 , n29560 , n29561 , n29562 , n29563 , n29564 , n29565 , n29566 , n29567 , n29568 , n29569 , n29570 , n29571 , n29572 , n29573 , n29574 , n29575 , n29576 , n29577 , n29578 , n29579 , n29580 , n29581 , n29582 , n29583 , n29584 , n29585 , n29586 , n29587 , n29588 , n29589 , n29590 , n29591 , n29592 , n29593 , n29594 , n29595 , n29596 , n29597 , n29598 , n29599 , n29600 , n29601 , n29602 , n29603 , n29604 , n29605 , n29606 , n29607 , n29608 , n29609 , n29610 , n29611 , n29612 , n29613 , n29614 , n29615 , n29616 , n29617 , n29618 , n29619 , n29620 , n29621 , n29622 , n29623 , n29624 , n29625 , n29626 , n29627 , n29628 , n29629 , n29630 , n29631 , n29632 , n29633 , n29634 , n29635 , n29636 , n29637 , n29638 , n29639 , n29640 , n29641 , n29642 , n29643 , n29644 , n29645 , n29646 , n29647 , n29648 , n29649 , n29650 , n29651 , n29652 , n29653 , n29654 , n29655 , n29656 , n29657 , n29658 , n29659 , n29660 , n29661 , n29662 , n29663 , n29664 , n29665 , n29666 , n29667 , n29668 , n29669 , n29670 , n29671 , n29672 , n29673 , n29674 , n29675 , n29676 , n29677 , n29678 , n29679 , n29680 , n29681 , n29682 , n29683 , n29684 , n29685 , n29686 , n29687 , n29688 , n29689 , n29690 , n29691 , n29692 , n29693 , n29694 , n29695 , n29696 , n29697 , n29698 , n29699 , n29700 , n29701 , n29702 , n29703 , n29704 , n29705 , n29706 , n29707 , n29708 , n29709 , n29710 , n29711 , n29712 , n29713 , n29714 , n29715 , n29716 , n29717 , n29718 , n29719 , n29720 , n29721 , n29722 , n29723 , n29724 , n29725 , n29726 , n29727 , n29728 , n29729 , n29730 , n29731 , n29732 , n29733 , n29734 , n29735 , n29736 , n29737 , n29738 , n29739 , n29740 , n29741 , n29742 , n29743 , n29744 , n29745 , n29746 , n29747 , n29748 , n29749 , n29750 , n29751 , n29752 , n29753 , n29754 , n29755 , n29756 , n29757 , n29758 , n29759 , n29760 , n29761 , n29762 , n29763 , n29764 , n29765 , n29766 , n29767 , n29768 , n29769 , n29770 , n29771 , n29772 , n29773 , n29774 , n29775 , n29776 , n29777 , n29778 , n29779 , n29780 , n29781 , n29782 , n29783 , n29784 , n29785 , n29786 , n29787 , n29788 , n29789 , n29790 , n29791 , n29792 , n29793 , n29794 , n29795 , n29796 , n29797 , n29798 , n29799 , n29800 , n29801 , n29802 , n29803 , n29804 , n29805 , n29806 , n29807 , n29808 , n29809 , n29810 , n29811 , n29812 , n29813 , n29814 , n29815 , n29816 , n29817 , n29818 , n29819 , n29820 , n29821 , n29822 , n29823 , n29824 , n29825 , n29826 , n29827 , n29828 , n29829 , n29830 , n29831 , n29832 , n29833 , n29834 , n29835 , n29836 , n29837 , n29838 , n29839 , n29840 , n29841 , n29842 , n29843 , n29844 , n29845 , n29846 , n29847 , n29848 , n29849 , n29850 , n29851 , n29852 , n29853 , n29854 , n29855 , n29856 , n29857 , n29858 , n29859 , n29860 , n29861 , n29862 , n29863 , n29864 , n29865 , n29866 , n29867 , n29868 , n29869 , n29870 , n29871 , n29872 , n29873 , n29874 , n29875 , n29876 , n29877 , n29878 , n29879 , n29880 , n29881 , n29882 , n29883 , n29884 , n29885 , n29886 , n29887 , n29888 , n29889 , n29890 , n29891 , n29892 , n29893 , n29894 , n29895 , n29896 , n29897 , n29898 , n29899 , n29900 , n29901 , n29902 , n29903 , n29904 , n29905 , n29906 , n29907 , n29908 , n29909 , n29910 , n29911 , n29912 , n29913 , n29914 , n29915 , n29916 , n29917 , n29918 , n29919 , n29920 , n29921 , n29922 , n29923 , n29924 , n29925 , n29926 , n29927 , n29928 , n29929 , n29930 , n29931 , n29932 , n29933 , n29934 , n29935 , n29936 , n29937 , n29938 , n29939 , n29940 , n29941 , n29942 , n29943 , n29944 , n29945 , n29946 , n29947 , n29948 , n29949 , n29950 , n29951 , n29952 , n29953 , n29954 , n29955 , n29956 , n29957 , n29958 , n29959 , n29960 , n29961 , n29962 , n29963 , n29964 , n29965 , n29966 , n29967 , n29968 , n29969 , n29970 , n29971 , n29972 , n29973 , n29974 , n29975 , n29976 , n29977 , n29978 , n29979 , n29980 , n29981 , n29982 , n29983 , n29984 , n29985 , n29986 , n29987 , n29988 , n29989 , n29990 , n29991 , n29992 , n29993 , n29994 , n29995 , n29996 , n29997 , n29998 , n29999 , n30000 , n30001 , n30002 , n30003 , n30004 , n30005 , n30006 , n30007 , n30008 , n30009 , n30010 , n30011 , n30012 , n30013 , n30014 , n30015 , n30016 , n30017 , n30018 , n30019 , n30020 , n30021 , n30022 , n30023 , n30024 , n30025 , n30026 , n30027 , n30028 , n30029 , n30030 , n30031 , n30032 , n30033 , n30034 , n30035 , n30036 , n30037 , n30038 , n30039 , n30040 , n30041 , n30042 , n30043 , n30044 , n30045 , n30046 , n30047 , n30048 , n30049 , n30050 , n30051 , n30052 , n30053 , n30054 , n30055 , n30056 , n30057 , n30058 , n30059 , n30060 , n30061 , n30062 , n30063 , n30064 , n30065 , n30066 , n30067 , n30068 , n30069 , n30070 , n30071 , n30072 , n30073 , n30074 , n30075 , n30076 , n30077 , n30078 , n30079 , n30080 , n30081 , n30082 , n30083 , n30084 , n30085 , n30086 , n30087 , n30088 , n30089 , n30090 , n30091 , n30092 , n30093 , n30094 , n30095 , n30096 , n30097 , n30098 , n30099 , n30100 , n30101 , n30102 , n30103 , n30104 , n30105 , n30106 , n30107 , n30108 , n30109 , n30110 , n30111 , n30112 , n30113 , n30114 , n30115 , n30116 , n30117 , n30118 , n30119 , n30120 , n30121 , n30122 , n30123 , n30124 , n30125 , n30126 , n30127 , n30128 , n30129 , n30130 , n30131 , n30132 , n30133 , n30134 , n30135 , n30136 , n30137 , n30138 , n30139 , n30140 , n30141 , n30142 , n30143 , n30144 , n30145 , n30146 , n30147 , n30148 , n30149 , n30150 , n30151 , n30152 , n30153 , n30154 , n30155 , n30156 , n30157 , n30158 , n30159 , n30160 , n30161 , n30162 , n30163 , n30164 , n30165 , n30166 , n30167 , n30168 , n30169 , n30170 , n30171 , n30172 , n30173 , n30174 , n30175 , n30176 , n30177 , n30178 , n30179 , n30180 , n30181 , n30182 , n30183 , n30184 , n30185 , n30186 , n30187 , n30188 , n30189 , n30190 , n30191 , n30192 , n30193 , n30194 , n30195 , n30196 , n30197 , n30198 , n30199 , n30200 , n30201 , n30202 , n30203 , n30204 , n30205 , n30206 , n30207 , n30208 , n30209 , n30210 , n30211 , n30212 , n30213 , n30214 , n30215 , n30216 , n30217 , n30218 , n30219 , n30220 , n30221 , n30222 , n30223 , n30224 , n30225 , n30226 , n30227 , n30228 , n30229 , n30230 , n30231 , n30232 , n30233 , n30234 , n30235 , n30236 , n30237 , n30238 , n30239 , n30240 , n30241 , n30242 , n30243 , n30244 , n30245 , n30246 , n30247 , n30248 , n30249 , n30250 , n30251 , n30252 , n30253 , n30254 , n30255 , n30256 , n30257 , n30258 , n30259 , n30260 , n30261 , n30262 , n30263 , n30264 , n30265 , n30266 , n30267 , n30268 , n30269 , n30270 , n30271 , n30272 , n30273 , n30274 , n30275 , n30276 , n30277 , n30278 , n30279 , n30280 , n30281 , n30282 , n30283 , n30284 , n30285 , n30286 , n30287 , n30288 , n30289 , n30290 , n30291 , n30292 , n30293 , n30294 , n30295 , n30296 , n30297 , n30298 , n30299 , n30300 , n30301 , n30302 , n30303 , n30304 , n30305 , n30306 , n30307 , n30308 , n30309 , n30310 , n30311 , n30312 , n30313 , n30314 , n30315 , n30316 , n30317 , n30318 , n30319 , n30320 , n30321 , n30322 , n30323 , n30324 , n30325 , n30326 , n30327 , n30328 , n30329 , n30330 , n30331 , n30332 , n30333 , n30334 , n30335 , n30336 , n30337 , n30338 , n30339 , n30340 , n30341 , n30342 , n30343 , n30344 , n30345 , n30346 , n30347 , n30348 , n30349 , n30350 , n30351 , n30352 , n30353 , n30354 , n30355 , n30356 , n30357 , n30358 , n30359 , n30360 , n30361 , n30362 , n30363 , n30364 , n30365 , n30366 , n30367 , n30368 , n30369 , n30370 , n30371 , n30372 , n30373 , n30374 , n30375 , n30376 , n30377 , n30378 , n30379 , n30380 , n30381 , n30382 , n30383 , n30384 , n30385 , n30386 , n30387 , n30388 , n30389 , n30390 , n30391 , n30392 , n30393 , n30394 , n30395 , n30396 , n30397 , n30398 , n30399 , n30400 , n30401 , n30402 , n30403 , n30404 , n30405 , n30406 , n30407 , n30408 , n30409 , n30410 , n30411 , n30412 , n30413 , n30414 , n30415 , n30416 , n30417 , n30418 , n30419 , n30420 , n30421 , n30422 , n30423 , n30424 , n30425 , n30426 , n30427 , n30428 , n30429 , n30430 , n30431 , n30432 , n30433 , n30434 , n30435 , n30436 , n30437 , n30438 , n30439 , n30440 , n30441 , n30442 , n30443 , n30444 , n30445 , n30446 , n30447 , n30448 , n30449 , n30450 , n30451 , n30452 , n30453 , n30454 , n30455 , n30456 , n30457 , n30458 , n30459 , n30460 , n30461 , n30462 , n30463 , n30464 , n30465 , n30466 , n30467 , n30468 , n30469 , n30470 , n30471 , n30472 , n30473 , n30474 , n30475 , n30476 , n30477 , n30478 , n30479 , n30480 , n30481 , n30482 , n30483 , n30484 , n30485 , n30486 , n30487 , n30488 , n30489 , n30490 , n30491 , n30492 , n30493 , n30494 , n30495 , n30496 , n30497 , n30498 , n30499 , n30500 , n30501 , n30502 , n30503 , n30504 , n30505 , n30506 , n30507 , n30508 , n30509 , n30510 , n30511 , n30512 , n30513 , n30514 , n30515 , n30516 , n30517 , n30518 , n30519 , n30520 , n30521 , n30522 , n30523 , n30524 , n30525 , n30526 , n30527 , n30528 , n30529 , n30530 , n30531 , n30532 , n30533 , n30534 , n30535 , n30536 , n30537 , n30538 , n30539 , n30540 , n30541 , n30542 , n30543 , n30544 , n30545 , n30546 , n30547 , n30548 , n30549 , n30550 , n30551 , n30552 , n30553 , n30554 , n30555 , n30556 , n30557 , n30558 , n30559 , n30560 , n30561 , n30562 , n30563 , n30564 , n30565 , n30566 , n30567 , n30568 , n30569 , n30570 , n30571 , n30572 , n30573 , n30574 , n30575 , n30576 , n30577 , n30578 , n30579 , n30580 , n30581 , n30582 , n30583 , n30584 , n30585 , n30586 , n30587 , n30588 , n30589 , n30590 , n30591 , n30592 , n30593 , n30594 , n30595 , n30596 , n30597 , n30598 , n30599 , n30600 , n30601 , n30602 , n30603 , n30604 , n30605 , n30606 , n30607 , n30608 , n30609 , n30610 , n30611 , n30612 , n30613 , n30614 , n30615 , n30616 , n30617 , n30618 , n30619 , n30620 , n30621 , n30622 , n30623 , n30624 , n30625 , n30626 , n30627 , n30628 , n30629 , n30630 , n30631 , n30632 , n30633 , n30634 , n30635 , n30636 , n30637 , n30638 , n30639 , n30640 , n30641 , n30642 , n30643 , n30644 , n30645 , n30646 , n30647 , n30648 , n30649 , n30650 , n30651 , n30652 , n30653 , n30654 , n30655 , n30656 , n30657 , n30658 , n30659 , n30660 , n30661 , n30662 , n30663 , n30664 , n30665 , n30666 , n30667 , n30668 , n30669 , n30670 , n30671 , n30672 , n30673 , n30674 , n30675 , n30676 , n30677 , n30678 , n30679 , n30680 , n30681 , n30682 , n30683 , n30684 , n30685 , n30686 , n30687 , n30688 , n30689 , n30690 , n30691 , n30692 , n30693 , n30694 , n30695 , n30696 , n30697 , n30698 , n30699 , n30700 , n30701 , n30702 , n30703 , n30704 , n30705 , n30706 , n30707 , n30708 , n30709 , n30710 , n30711 , n30712 , n30713 , n30714 , n30715 , n30716 , n30717 , n30718 , n30719 , n30720 , n30721 , n30722 , n30723 , n30724 , n30725 , n30726 , n30727 , n30728 , n30729 , n30730 , n30731 , n30732 , n30733 , n30734 , n30735 , n30736 , n30737 , n30738 , n30739 , n30740 , n30741 , n30742 , n30743 , n30744 , n30745 , n30746 , n30747 , n30748 , n30749 , n30750 , n30751 , n30752 , n30753 , n30754 , n30755 , n30756 , n30757 , n30758 , n30759 , n30760 , n30761 , n30762 , n30763 , n30764 , n30765 , n30766 , n30767 , n30768 , n30769 , n30770 , n30771 , n30772 , n30773 , n30774 , n30775 , n30776 , n30777 , n30778 , n30779 , n30780 , n30781 , n30782 , n30783 , n30784 , n30785 , n30786 , n30787 , n30788 , n30789 , n30790 , n30791 , n30792 , n30793 , n30794 , n30795 , n30796 , n30797 , n30798 , n30799 , n30800 , n30801 , n30802 , n30803 , n30804 , n30805 , n30806 , n30807 , n30808 , n30809 , n30810 , n30811 , n30812 , n30813 , n30814 , n30815 , n30816 , n30817 , n30818 , n30819 , n30820 , n30821 , n30822 , n30823 , n30824 , n30825 , n30826 , n30827 , n30828 , n30829 , n30830 , n30831 , n30832 , n30833 , n30834 , n30835 , n30836 , n30837 , n30838 , n30839 , n30840 , n30841 , n30842 , n30843 , n30844 , n30845 , n30846 , n30847 , n30848 , n30849 , n30850 , n30851 , n30852 , n30853 , n30854 , n30855 , n30856 , n30857 , n30858 , n30859 , n30860 , n30861 , n30862 , n30863 , n30864 , n30865 , n30866 , n30867 , n30868 , n30869 , n30870 , n30871 , n30872 , n30873 , n30874 , n30875 , n30876 , n30877 , n30878 , n30879 , n30880 , n30881 , n30882 , n30883 , n30884 , n30885 , n30886 , n30887 , n30888 , n30889 , n30890 , n30891 , n30892 , n30893 , n30894 , n30895 , n30896 , n30897 , n30898 , n30899 , n30900 , n30901 , n30902 , n30903 , n30904 , n30905 , n30906 , n30907 , n30908 , n30909 , n30910 , n30911 , n30912 , n30913 , n30914 , n30915 , n30916 , n30917 , n30918 , n30919 , n30920 , n30921 , n30922 , n30923 , n30924 , n30925 , n30926 , n30927 , n30928 , n30929 , n30930 , n30931 , n30932 , n30933 , n30934 , n30935 , n30936 , n30937 , n30938 , n30939 , n30940 , n30941 , n30942 , n30943 , n30944 , n30945 , n30946 , n30947 , n30948 , n30949 , n30950 , n30951 , n30952 , n30953 , n30954 , n30955 , n30956 , n30957 , n30958 , n30959 , n30960 , n30961 , n30962 , n30963 , n30964 , n30965 , n30966 , n30967 , n30968 , n30969 , n30970 , n30971 , n30972 , n30973 , n30974 , n30975 , n30976 , n30977 , n30978 , n30979 , n30980 , n30981 , n30982 , n30983 , n30984 , n30985 , n30986 , n30987 , n30988 , n30989 , n30990 , n30991 , n30992 , n30993 , n30994 , n30995 , n30996 , n30997 , n30998 , n30999 , n31000 , n31001 , n31002 , n31003 , n31004 , n31005 , n31006 , n31007 , n31008 , n31009 , n31010 , n31011 , n31012 , n31013 , n31014 , n31015 , n31016 , n31017 , n31018 , n31019 , n31020 , n31021 , n31022 , n31023 , n31024 , n31025 , n31026 , n31027 , n31028 , n31029 , n31030 , n31031 , n31032 , n31033 , n31034 , n31035 , n31036 , n31037 , n31038 , n31039 , n31040 , n31041 , n31042 , n31043 , n31044 , n31045 , n31046 , n31047 , n31048 , n31049 , n31050 , n31051 , n31052 , n31053 , n31054 , n31055 , n31056 , n31057 , n31058 , n31059 , n31060 , n31061 , n31062 , n31063 , n31064 , n31065 , n31066 , n31067 , n31068 , n31069 , n31070 , n31071 , n31072 , n31073 , n31074 , n31075 , n31076 , n31077 , n31078 , n31079 , n31080 , n31081 , n31082 , n31083 , n31084 , n31085 , n31086 , n31087 , n31088 , n31089 , n31090 , n31091 , n31092 , n31093 , n31094 , n31095 , n31096 , n31097 , n31098 , n31099 , n31100 , n31101 , n31102 , n31103 , n31104 , n31105 , n31106 , n31107 , n31108 , n31109 , n31110 , n31111 , n31112 , n31113 , n31114 , n31115 , n31116 , n31117 , n31118 , n31119 , n31120 , n31121 , n31122 , n31123 , n31124 , n31125 , n31126 , n31127 , n31128 , n31129 , n31130 , n31131 , n31132 , n31133 , n31134 , n31135 , n31136 , n31137 , n31138 , n31139 , n31140 , n31141 , n31142 , n31143 , n31144 , n31145 , n31146 , n31147 , n31148 , n31149 , n31150 , n31151 , n31152 , n31153 , n31154 , n31155 , n31156 , n31157 , n31158 , n31159 , n31160 , n31161 , n31162 , n31163 , n31164 , n31165 , n31166 , n31167 , n31168 , n31169 , n31170 , n31171 , n31172 , n31173 , n31174 , n31175 , n31176 , n31177 , n31178 , n31179 , n31180 , n31181 , n31182 , n31183 , n31184 , n31185 , n31186 , n31187 , n31188 , n31189 , n31190 , n31191 , n31192 , n31193 , n31194 , n31195 , n31196 , n31197 , n31198 , n31199 , n31200 , n31201 , n31202 , n31203 , n31204 , n31205 , n31206 , n31207 , n31208 , n31209 , n31210 , n31211 , n31212 , n31213 , n31214 , n31215 , n31216 , n31217 , n31218 , n31219 , n31220 , n31221 , n31222 , n31223 , n31224 , n31225 , n31226 , n31227 , n31228 , n31229 , n31230 , n31231 , n31232 , n31233 , n31234 , n31235 , n31236 , n31237 , n31238 , n31239 , n31240 , n31241 , n31242 , n31243 , n31244 , n31245 , n31246 , n31247 , n31248 , n31249 , n31250 , n31251 , n31252 , n31253 , n31254 , n31255 , n31256 , n31257 , n31258 , n31259 , n31260 , n31261 , n31262 , n31263 , n31264 , n31265 , n31266 , n31267 , n31268 , n31269 , n31270 , n31271 , n31272 , n31273 , n31274 , n31275 , n31276 , n31277 , n31278 , n31279 , n31280 , n31281 , n31282 , n31283 , n31284 , n31285 , n31286 , n31287 , n31288 , n31289 , n31290 , n31291 , n31292 , n31293 , n31294 , n31295 , n31296 , n31297 , n31298 , n31299 , n31300 , n31301 , n31302 , n31303 , n31304 , n31305 , n31306 , n31307 , n31308 , n31309 , n31310 , n31311 , n31312 , n31313 , n31314 , n31315 , n31316 , n31317 , n31318 , n31319 , n31320 , n31321 , n31322 , n31323 , n31324 , n31325 , n31326 , n31327 , n31328 , n31329 , n31330 , n31331 , n31332 , n31333 , n31334 , n31335 , n31336 , n31337 , n31338 , n31339 , n31340 , n31341 , n31342 , n31343 , n31344 , n31345 , n31346 , n31347 , n31348 , n31349 , n31350 , n31351 , n31352 , n31353 , n31354 , n31355 , n31356 , n31357 , n31358 , n31359 , n31360 , n31361 , n31362 , n31363 , n31364 , n31365 , n31366 , n31367 , n31368 , n31369 , n31370 , n31371 , n31372 , n31373 , n31374 , n31375 , n31376 , n31377 , n31378 , n31379 , n31380 , n31381 , n31382 , n31383 , n31384 , n31385 , n31386 , n31387 , n31388 , n31389 , n31390 , n31391 , n31392 , n31393 , n31394 , n31395 , n31396 , n31397 , n31398 , n31399 , n31400 , n31401 , n31402 , n31403 , n31404 , n31405 , n31406 , n31407 , n31408 , n31409 , n31410 , n31411 , n31412 , n31413 , n31414 , n31415 , n31416 , n31417 , n31418 , n31419 , n31420 , n31421 , n31422 , n31423 , n31424 , n31425 , n31426 , n31427 , n31428 , n31429 , n31430 , n31431 , n31432 , n31433 , n31434 , n31435 , n31436 , n31437 , n31438 , n31439 , n31440 , n31441 , n31442 , n31443 , n31444 , n31445 , n31446 , n31447 , n31448 , n31449 , n31450 , n31451 , n31452 , n31453 , n31454 , n31455 , n31456 , n31457 , n31458 , n31459 , n31460 , n31461 , n31462 , n31463 , n31464 , n31465 , n31466 , n31467 , n31468 , n31469 , n31470 , n31471 , n31472 , n31473 , n31474 , n31475 , n31476 , n31477 , n31478 , n31479 , n31480 , n31481 , n31482 , n31483 , n31484 , n31485 , n31486 , n31487 , n31488 , n31489 , n31490 , n31491 , n31492 , n31493 , n31494 , n31495 , n31496 , n31497 , n31498 , n31499 , n31500 , n31501 , n31502 , n31503 , n31504 , n31505 , n31506 , n31507 , n31508 , n31509 , n31510 , n31511 , n31512 , n31513 , n31514 , n31515 , n31516 , n31517 , n31518 , n31519 , n31520 , n31521 , n31522 , n31523 , n31524 , n31525 , n31526 , n31527 , n31528 , n31529 , n31530 , n31531 , n31532 , n31533 , n31534 , n31535 , n31536 , n31537 , n31538 , n31539 , n31540 , n31541 , n31542 , n31543 , n31544 , n31545 , n31546 , n31547 , n31548 , n31549 , n31550 , n31551 , n31552 , n31553 , n31554 , n31555 , n31556 , n31557 , n31558 , n31559 , n31560 , n31561 , n31562 , n31563 , n31564 , n31565 , n31566 , n31567 , n31568 , n31569 , n31570 , n31571 , n31572 , n31573 , n31574 , n31575 , n31576 , n31577 , n31578 , n31579 , n31580 , n31581 , n31582 , n31583 , n31584 , n31585 , n31586 , n31587 , n31588 , n31589 , n31590 , n31591 , n31592 , n31593 , n31594 , n31595 , n31596 , n31597 , n31598 , n31599 , n31600 , n31601 , n31602 , n31603 , n31604 , n31605 , n31606 , n31607 , n31608 , n31609 , n31610 , n31611 , n31612 , n31613 , n31614 , n31615 , n31616 , n31617 , n31618 , n31619 , n31620 , n31621 , n31622 , n31623 , n31624 , n31625 , n31626 , n31627 , n31628 , n31629 , n31630 , n31631 , n31632 , n31633 , n31634 , n31635 , n31636 , n31637 , n31638 , n31639 , n31640 , n31641 , n31642 , n31643 , n31644 , n31645 , n31646 , n31647 , n31648 , n31649 , n31650 , n31651 , n31652 , n31653 , n31654 , n31655 , n31656 , n31657 , n31658 , n31659 , n31660 , n31661 , n31662 , n31663 , n31664 , n31665 , n31666 , n31667 , n31668 , n31669 , n31670 , n31671 , n31672 , n31673 , n31674 , n31675 , n31676 , n31677 , n31678 , n31679 , n31680 , n31681 , n31682 , n31683 , n31684 , n31685 , n31686 , n31687 , n31688 , n31689 , n31690 , n31691 , n31692 , n31693 , n31694 , n31695 , n31696 , n31697 , n31698 , n31699 , n31700 , n31701 , n31702 , n31703 , n31704 , n31705 , n31706 , n31707 , n31708 , n31709 , n31710 , n31711 , n31712 , n31713 , n31714 , n31715 , n31716 , n31717 , n31718 , n31719 , n31720 , n31721 , n31722 , n31723 , n31724 , n31725 , n31726 , n31727 , n31728 , n31729 , n31730 , n31731 , n31732 , n31733 , n31734 , n31735 , n31736 , n31737 , n31738 , n31739 , n31740 , n31741 , n31742 , n31743 , n31744 , n31745 , n31746 , n31747 , n31748 , n31749 , n31750 , n31751 , n31752 , n31753 , n31754 , n31755 , n31756 , n31757 , n31758 , n31759 , n31760 , n31761 , n31762 , n31763 , n31764 , n31765 , n31766 , n31767 , n31768 , n31769 , n31770 , n31771 , n31772 , n31773 , n31774 , n31775 , n31776 , n31777 , n31778 , n31779 , n31780 , n31781 , n31782 , n31783 , n31784 , n31785 , n31786 , n31787 , n31788 , n31789 , n31790 , n31791 , n31792 , n31793 , n31794 , n31795 , n31796 , n31797 , n31798 , n31799 , n31800 , n31801 , n31802 , n31803 , n31804 , n31805 , n31806 , n31807 , n31808 , n31809 , n31810 , n31811 , n31812 , n31813 , n31814 , n31815 , n31816 , n31817 , n31818 , n31819 , n31820 , n31821 , n31822 , n31823 , n31824 , n31825 , n31826 , n31827 , n31828 , n31829 , n31830 , n31831 , n31832 , n31833 , n31834 , n31835 , n31836 , n31837 , n31838 , n31839 , n31840 , n31841 , n31842 , n31843 , n31844 , n31845 , n31846 , n31847 , n31848 , n31849 , n31850 , n31851 , n31852 , n31853 , n31854 , n31855 , n31856 , n31857 , n31858 , n31859 , n31860 , n31861 , n31862 , n31863 , n31864 , n31865 , n31866 , n31867 , n31868 , n31869 , n31870 , n31871 , n31872 , n31873 , n31874 , n31875 , n31876 , n31877 , n31878 , n31879 , n31880 , n31881 , n31882 , n31883 , n31884 , n31885 , n31886 , n31887 , n31888 , n31889 , n31890 , n31891 , n31892 , n31893 , n31894 , n31895 , n31896 , n31897 , n31898 , n31899 , n31900 , n31901 , n31902 , n31903 , n31904 , n31905 , n31906 , n31907 , n31908 , n31909 , n31910 , n31911 , n31912 , n31913 , n31914 , n31915 , n31916 , n31917 , n31918 , n31919 , n31920 , n31921 , n31922 , n31923 , n31924 , n31925 , n31926 , n31927 , n31928 , n31929 , n31930 , n31931 , n31932 , n31933 , n31934 , n31935 , n31936 , n31937 , n31938 , n31939 , n31940 , n31941 , n31942 , n31943 , n31944 , n31945 , n31946 , n31947 , n31948 , n31949 , n31950 , n31951 , n31952 , n31953 , n31954 , n31955 , n31956 , n31957 , n31958 , n31959 , n31960 , n31961 , n31962 , n31963 , n31964 , n31965 , n31966 , n31967 , n31968 , n31969 , n31970 , n31971 , n31972 , n31973 , n31974 , n31975 , n31976 , n31977 , n31978 , n31979 , n31980 , n31981 , n31982 , n31983 , n31984 , n31985 , n31986 , n31987 , n31988 , n31989 , n31990 , n31991 , n31992 , n31993 , n31994 , n31995 , n31996 , n31997 , n31998 , n31999 , n32000 , n32001 , n32002 , n32003 , n32004 , n32005 , n32006 , n32007 , n32008 , n32009 , n32010 , n32011 , n32012 , n32013 , n32014 , n32015 , n32016 , n32017 , n32018 , n32019 , n32020 , n32021 , n32022 , n32023 , n32024 , n32025 , n32026 , n32027 , n32028 , n32029 , n32030 , n32031 , n32032 , n32033 , n32034 , n32035 , n32036 , n32037 , n32038 , n32039 , n32040 , n32041 , n32042 , n32043 , n32044 , n32045 , n32046 , n32047 , n32048 , n32049 , n32050 , n32051 , n32052 , n32053 , n32054 , n32055 , n32056 , n32057 , n32058 , n32059 , n32060 , n32061 , n32062 , n32063 , n32064 , n32065 , n32066 , n32067 , n32068 , n32069 , n32070 , n32071 , n32072 , n32073 , n32074 , n32075 , n32076 , n32077 , n32078 , n32079 , n32080 , n32081 , n32082 , n32083 , n32084 , n32085 , n32086 , n32087 , n32088 , n32089 , n32090 , n32091 , n32092 , n32093 , n32094 , n32095 , n32096 , n32097 , n32098 , n32099 , n32100 , n32101 , n32102 , n32103 , n32104 , n32105 , n32106 , n32107 , n32108 , n32109 , n32110 , n32111 , n32112 , n32113 , n32114 , n32115 , n32116 , n32117 , n32118 , n32119 , n32120 , n32121 , n32122 , n32123 , n32124 , n32125 , n32126 , n32127 , n32128 , n32129 , n32130 , n32131 , n32132 , n32133 , n32134 , n32135 , n32136 , n32137 , n32138 , n32139 , n32140 , n32141 , n32142 , n32143 , n32144 , n32145 , n32146 , n32147 , n32148 , n32149 , n32150 , n32151 , n32152 , n32153 , n32154 , n32155 , n32156 , n32157 , n32158 , n32159 , n32160 , n32161 , n32162 , n32163 , n32164 , n32165 , n32166 , n32167 , n32168 , n32169 , n32170 , n32171 , n32172 , n32173 , n32174 , n32175 , n32176 , n32177 , n32178 , n32179 , n32180 , n32181 , n32182 , n32183 , n32184 , n32185 , n32186 , n32187 , n32188 , n32189 , n32190 , n32191 , n32192 , n32193 , n32194 , n32195 , n32196 , n32197 , n32198 , n32199 , n32200 , n32201 , n32202 , n32203 , n32204 , n32205 , n32206 , n32207 , n32208 , n32209 , n32210 , n32211 , n32212 , n32213 , n32214 , n32215 , n32216 , n32217 , n32218 , n32219 , n32220 , n32221 , n32222 , n32223 , n32224 , n32225 , n32226 , n32227 , n32228 , n32229 , n32230 , n32231 , n32232 , n32233 , n32234 , n32235 , n32236 , n32237 , n32238 , n32239 , n32240 , n32241 , n32242 , n32243 , n32244 , n32245 , n32246 , n32247 , n32248 , n32249 , n32250 , n32251 , n32252 , n32253 , n32254 , n32255 , n32256 , n32257 , n32258 , n32259 , n32260 , n32261 , n32262 , n32263 , n32264 , n32265 , n32266 , n32267 , n32268 , n32269 , n32270 , n32271 , n32272 , n32273 , n32274 , n32275 , n32276 , n32277 , n32278 , n32279 , n32280 , n32281 , n32282 , n32283 , n32284 , n32285 , n32286 , n32287 , n32288 , n32289 , n32290 , n32291 , n32292 , n32293 , n32294 , n32295 , n32296 , n32297 , n32298 , n32299 , n32300 , n32301 , n32302 , n32303 , n32304 , n32305 , n32306 , n32307 , n32308 , n32309 , n32310 , n32311 , n32312 , n32313 , n32314 , n32315 , n32316 , n32317 , n32318 , n32319 , n32320 , n32321 , n32322 , n32323 , n32324 , n32325 , n32326 , n32327 , n32328 , n32329 , n32330 , n32331 , n32332 , n32333 , n32334 , n32335 , n32336 , n32337 , n32338 , n32339 , n32340 , n32341 , n32342 , n32343 , n32344 , n32345 , n32346 , n32347 , n32348 , n32349 , n32350 , n32351 , n32352 , n32353 , n32354 , n32355 , n32356 , n32357 , n32358 , n32359 , n32360 , n32361 , n32362 , n32363 , n32364 , n32365 , n32366 , n32367 , n32368 , n32369 , n32370 , n32371 , n32372 , n32373 , n32374 , n32375 , n32376 , n32377 , n32378 , n32379 , n32380 , n32381 , n32382 , n32383 , n32384 , n32385 , n32386 , n32387 , n32388 , n32389 , n32390 , n32391 , n32392 , n32393 , n32394 , n32395 , n32396 , n32397 , n32398 , n32399 , n32400 , n32401 , n32402 , n32403 , n32404 , n32405 , n32406 , n32407 , n32408 , n32409 , n32410 , n32411 , n32412 , n32413 , n32414 , n32415 , n32416 , n32417 , n32418 , n32419 , n32420 , n32421 , n32422 , n32423 , n32424 , n32425 , n32426 , n32427 , n32428 , n32429 , n32430 , n32431 , n32432 , n32433 , n32434 , n32435 , n32436 , n32437 , n32438 , n32439 , n32440 , n32441 , n32442 , n32443 , n32444 , n32445 , n32446 , n32447 , n32448 , n32449 , n32450 , n32451 , n32452 , n32453 , n32454 , n32455 , n32456 , n32457 , n32458 , n32459 , n32460 , n32461 , n32462 , n32463 , n32464 , n32465 , n32466 , n32467 , n32468 , n32469 , n32470 , n32471 , n32472 , n32473 , n32474 , n32475 , n32476 , n32477 , n32478 , n32479 , n32480 , n32481 , n32482 , n32483 , n32484 , n32485 , n32486 , n32487 , n32488 , n32489 , n32490 , n32491 , n32492 , n32493 , n32494 , n32495 , n32496 , n32497 , n32498 , n32499 , n32500 , n32501 , n32502 , n32503 , n32504 , n32505 , n32506 , n32507 , n32508 , n32509 , n32510 , n32511 , n32512 , n32513 , n32514 , n32515 , n32516 , n32517 , n32518 , n32519 , n32520 , n32521 , n32522 , n32523 , n32524 , n32525 , n32526 , n32527 , n32528 , n32529 , n32530 , n32531 , n32532 , n32533 , n32534 , n32535 , n32536 , n32537 , n32538 , n32539 , n32540 , n32541 , n32542 , n32543 , n32544 , n32545 , n32546 , n32547 , n32548 , n32549 , n32550 , n32551 , n32552 , n32553 , n32554 , n32555 , n32556 , n32557 , n32558 , n32559 , n32560 , n32561 , n32562 , n32563 , n32564 , n32565 , n32566 , n32567 , n32568 , n32569 , n32570 , n32571 , n32572 , n32573 , n32574 , n32575 , n32576 , n32577 , n32578 , n32579 , n32580 , n32581 , n32582 , n32583 , n32584 , n32585 , n32586 , n32587 , n32588 , n32589 , n32590 , n32591 , n32592 , n32593 , n32594 , n32595 , n32596 , n32597 , n32598 , n32599 , n32600 , n32601 , n32602 , n32603 , n32604 , n32605 , n32606 , n32607 , n32608 , n32609 , n32610 , n32611 , n32612 , n32613 , n32614 , n32615 , n32616 , n32617 , n32618 , n32619 , n32620 , n32621 , n32622 , n32623 , n32624 , n32625 , n32626 , n32627 , n32628 , n32629 , n32630 , n32631 , n32632 , n32633 , n32634 , n32635 , n32636 , n32637 , n32638 , n32639 , n32640 , n32641 , n32642 , n32643 , n32644 , n32645 , n32646 , n32647 , n32648 , n32649 , n32650 , n32651 , n32652 , n32653 , n32654 , n32655 , n32656 , n32657 , n32658 , n32659 , n32660 , n32661 , n32662 , n32663 , n32664 , n32665 , n32666 , n32667 , n32668 , n32669 , n32670 , n32671 , n32672 , n32673 , n32674 , n32675 , n32676 , n32677 , n32678 , n32679 , n32680 , n32681 , n32682 , n32683 , n32684 , n32685 , n32686 , n32687 , n32688 , n32689 , n32690 , n32691 , n32692 , n32693 , n32694 , n32695 , n32696 , n32697 , n32698 , n32699 , n32700 , n32701 , n32702 , n32703 , n32704 , n32705 , n32706 , n32707 , n32708 , n32709 , n32710 , n32711 , n32712 , n32713 , n32714 , n32715 , n32716 , n32717 , n32718 , n32719 , n32720 , n32721 , n32722 , n32723 , n32724 , n32725 , n32726 , n32727 , n32728 , n32729 , n32730 , n32731 , n32732 , n32733 , n32734 , n32735 , n32736 , n32737 , n32738 , n32739 , n32740 , n32741 , n32742 , n32743 , n32744 , n32745 , n32746 , n32747 , n32748 , n32749 , n32750 , n32751 , n32752 , n32753 , n32754 , n32755 , n32756 , n32757 , n32758 , n32759 , n32760 , n32761 , n32762 , n32763 , n32764 , n32765 , n32766 , n32767 , n32768 , n32769 , n32770 , n32771 , n32772 , n32773 , n32774 , n32775 , n32776 , n32777 , n32778 , n32779 , n32780 , n32781 , n32782 , n32783 , n32784 , n32785 , n32786 , n32787 , n32788 , n32789 , n32790 , n32791 , n32792 , n32793 , n32794 , n32795 , n32796 , n32797 , n32798 , n32799 , n32800 , n32801 , n32802 , n32803 , n32804 , n32805 , n32806 , n32807 , n32808 , n32809 , n32810 , n32811 , n32812 , n32813 , n32814 , n32815 , n32816 , n32817 , n32818 , n32819 , n32820 , n32821 , n32822 , n32823 , n32824 , n32825 , n32826 , n32827 , n32828 , n32829 , n32830 , n32831 , n32832 , n32833 , n32834 , n32835 , n32836 , n32837 , n32838 , n32839 , n32840 , n32841 , n32842 , n32843 , n32844 , n32845 , n32846 , n32847 , n32848 , n32849 , n32850 , n32851 , n32852 , n32853 , n32854 , n32855 , n32856 , n32857 , n32858 , n32859 , n32860 , n32861 , n32862 , n32863 , n32864 , n32865 , n32866 , n32867 , n32868 , n32869 , n32870 , n32871 , n32872 , n32873 , n32874 , n32875 , n32876 , n32877 , n32878 , n32879 , n32880 , n32881 , n32882 , n32883 , n32884 , n32885 , n32886 , n32887 , n32888 , n32889 , n32890 , n32891 , n32892 , n32893 , n32894 , n32895 , n32896 , n32897 , n32898 , n32899 , n32900 , n32901 , n32902 , n32903 , n32904 , n32905 , n32906 , n32907 , n32908 , n32909 , n32910 , n32911 , n32912 , n32913 , n32914 , n32915 , n32916 , n32917 , n32918 , n32919 , n32920 , n32921 , n32922 , n32923 , n32924 , n32925 , n32926 , n32927 , n32928 , n32929 , n32930 , n32931 , n32932 , n32933 , n32934 , n32935 , n32936 , n32937 , n32938 , n32939 , n32940 , n32941 , n32942 , n32943 , n32944 , n32945 , n32946 , n32947 , n32948 , n32949 , n32950 , n32951 , n32952 , n32953 , n32954 , n32955 , n32956 , n32957 , n32958 , n32959 , n32960 , n32961 , n32962 , n32963 , n32964 , n32965 , n32966 , n32967 , n32968 , n32969 , n32970 , n32971 , n32972 , n32973 , n32974 , n32975 , n32976 , n32977 , n32978 , n32979 , n32980 , n32981 , n32982 , n32983 , n32984 , n32985 , n32986 , n32987 , n32988 , n32989 , n32990 , n32991 , n32992 , n32993 , n32994 , n32995 , n32996 , n32997 , n32998 , n32999 , n33000 , n33001 , n33002 , n33003 , n33004 , n33005 , n33006 , n33007 , n33008 , n33009 , n33010 , n33011 , n33012 , n33013 , n33014 , n33015 , n33016 , n33017 , n33018 , n33019 , n33020 , n33021 , n33022 , n33023 , n33024 , n33025 , n33026 , n33027 , n33028 , n33029 , n33030 , n33031 , n33032 , n33033 , n33034 , n33035 , n33036 , n33037 , n33038 , n33039 , n33040 , n33041 , n33042 , n33043 , n33044 , n33045 , n33046 , n33047 , n33048 , n33049 , n33050 , n33051 , n33052 , n33053 , n33054 , n33055 , n33056 , n33057 , n33058 , n33059 , n33060 , n33061 , n33062 , n33063 , n33064 , n33065 , n33066 , n33067 , n33068 , n33069 , n33070 , n33071 , n33072 , n33073 , n33074 , n33075 , n33076 , n33077 , n33078 , n33079 , n33080 , n33081 , n33082 , n33083 , n33084 , n33085 , n33086 , n33087 , n33088 , n33089 , n33090 , n33091 , n33092 , n33093 , n33094 , n33095 , n33096 , n33097 , n33098 , n33099 , n33100 , n33101 , n33102 , n33103 , n33104 , n33105 , n33106 , n33107 , n33108 , n33109 , n33110 , n33111 , n33112 , n33113 , n33114 , n33115 , n33116 , n33117 , n33118 , n33119 , n33120 , n33121 , n33122 , n33123 , n33124 , n33125 , n33126 , n33127 , n33128 , n33129 , n33130 , n33131 , n33132 , n33133 , n33134 , n33135 , n33136 , n33137 , n33138 , n33139 , n33140 , n33141 , n33142 , n33143 , n33144 , n33145 , n33146 , n33147 , n33148 , n33149 , n33150 , n33151 , n33152 , n33153 , n33154 , n33155 , n33156 , n33157 , n33158 , n33159 , n33160 , n33161 , n33162 , n33163 , n33164 , n33165 , n33166 , n33167 , n33168 , n33169 , n33170 , n33171 , n33172 , n33173 , n33174 , n33175 , n33176 , n33177 , n33178 , n33179 , n33180 , n33181 , n33182 , n33183 , n33184 , n33185 , n33186 , n33187 , n33188 , n33189 , n33190 , n33191 , n33192 , n33193 , n33194 , n33195 , n33196 , n33197 , n33198 , n33199 , n33200 , n33201 , n33202 , n33203 , n33204 , n33205 , n33206 , n33207 , n33208 , n33209 , n33210 , n33211 , n33212 , n33213 , n33214 , n33215 , n33216 , n33217 , n33218 , n33219 , n33220 , n33221 , n33222 , n33223 , n33224 , n33225 , n33226 , n33227 , n33228 , n33229 , n33230 , n33231 , n33232 , n33233 , n33234 , n33235 , n33236 , n33237 , n33238 , n33239 , n33240 , n33241 , n33242 , n33243 , n33244 , n33245 , n33246 , n33247 , n33248 , n33249 , n33250 , n33251 , n33252 , n33253 , n33254 , n33255 , n33256 , n33257 , n33258 , n33259 , n33260 , n33261 , n33262 , n33263 , n33264 , n33265 , n33266 , n33267 , n33268 , n33269 , n33270 , n33271 , n33272 , n33273 , n33274 , n33275 , n33276 , n33277 , n33278 , n33279 , n33280 , n33281 , n33282 , n33283 , n33284 , n33285 , n33286 , n33287 , n33288 , n33289 , n33290 , n33291 , n33292 , n33293 , n33294 , n33295 , n33296 , n33297 , n33298 , n33299 , n33300 , n33301 , n33302 , n33303 , n33304 , n33305 , n33306 , n33307 , n33308 , n33309 , n33310 , n33311 , n33312 , n33313 , n33314 , n33315 , n33316 , n33317 , n33318 , n33319 , n33320 , n33321 , n33322 , n33323 , n33324 , n33325 , n33326 , n33327 , n33328 , n33329 , n33330 , n33331 , n33332 , n33333 , n33334 , n33335 , n33336 , n33337 , n33338 , n33339 , n33340 , n33341 , n33342 , n33343 , n33344 , n33345 , n33346 , n33347 , n33348 , n33349 , n33350 , n33351 , n33352 , n33353 , n33354 , n33355 , n33356 , n33357 , n33358 , n33359 , n33360 , n33361 , n33362 , n33363 , n33364 , n33365 , n33366 , n33367 , n33368 , n33369 , n33370 , n33371 , n33372 , n33373 , n33374 , n33375 , n33376 , n33377 , n33378 , n33379 , n33380 , n33381 , n33382 , n33383 , n33384 , n33385 , n33386 , n33387 , n33388 , n33389 , n33390 , n33391 , n33392 , n33393 , n33394 , n33395 , n33396 , n33397 , n33398 , n33399 , n33400 , n33401 , n33402 , n33403 , n33404 , n33405 , n33406 , n33407 , n33408 , n33409 , n33410 , n33411 , n33412 , n33413 , n33414 , n33415 , n33416 , n33417 , n33418 , n33419 , n33420 , n33421 , n33422 , n33423 , n33424 , n33425 , n33426 , n33427 , n33428 , n33429 , n33430 , n33431 , n33432 , n33433 , n33434 , n33435 , n33436 , n33437 , n33438 , n33439 , n33440 , n33441 , n33442 , n33443 , n33444 , n33445 , n33446 , n33447 , n33448 , n33449 , n33450 , n33451 , n33452 , n33453 , n33454 , n33455 , n33456 , n33457 , n33458 , n33459 , n33460 , n33461 , n33462 , n33463 , n33464 , n33465 , n33466 , n33467 , n33468 , n33469 , n33470 , n33471 , n33472 , n33473 , n33474 , n33475 , n33476 , n33477 , n33478 , n33479 , n33480 , n33481 , n33482 , n33483 , n33484 , n33485 , n33486 , n33487 , n33488 , n33489 , n33490 , n33491 , n33492 , n33493 , n33494 , n33495 , n33496 , n33497 , n33498 , n33499 , n33500 , n33501 , n33502 , n33503 , n33504 , n33505 , n33506 , n33507 , n33508 , n33509 , n33510 , n33511 , n33512 , n33513 , n33514 , n33515 , n33516 , n33517 , n33518 , n33519 , n33520 , n33521 , n33522 , n33523 , n33524 , n33525 , n33526 , n33527 , n33528 , n33529 , n33530 , n33531 , n33532 , n33533 , n33534 , n33535 , n33536 , n33537 , n33538 , n33539 , n33540 , n33541 , n33542 , n33543 , n33544 , n33545 , n33546 , n33547 , n33548 , n33549 , n33550 , n33551 , n33552 , n33553 , n33554 , n33555 , n33556 , n33557 , n33558 , n33559 , n33560 , n33561 , n33562 , n33563 , n33564 , n33565 , n33566 , n33567 , n33568 , n33569 , n33570 , n33571 , n33572 , n33573 , n33574 , n33575 , n33576 , n33577 , n33578 , n33579 , n33580 , n33581 , n33582 , n33583 , n33584 , n33585 , n33586 , n33587 , n33588 , n33589 , n33590 , n33591 , n33592 , n33593 , n33594 , n33595 , n33596 , n33597 , n33598 , n33599 , n33600 , n33601 , n33602 , n33603 , n33604 , n33605 , n33606 , n33607 , n33608 , n33609 , n33610 , n33611 , n33612 , n33613 , n33614 , n33615 , n33616 , n33617 , n33618 , n33619 , n33620 , n33621 , n33622 , n33623 , n33624 , n33625 , n33626 , n33627 , n33628 , n33629 , n33630 , n33631 , n33632 , n33633 , n33634 , n33635 , n33636 , n33637 , n33638 , n33639 , n33640 , n33641 , n33642 , n33643 , n33644 , n33645 , n33646 , n33647 , n33648 , n33649 , n33650 , n33651 , n33652 , n33653 , n33654 , n33655 , n33656 , n33657 , n33658 , n33659 , n33660 , n33661 , n33662 , n33663 , n33664 , n33665 , n33666 , n33667 , n33668 , n33669 , n33670 , n33671 , n33672 , n33673 , n33674 , n33675 , n33676 , n33677 , n33678 , n33679 , n33680 , n33681 , n33682 , n33683 , n33684 , n33685 , n33686 , n33687 , n33688 , n33689 , n33690 , n33691 , n33692 , n33693 , n33694 , n33695 , n33696 , n33697 , n33698 , n33699 , n33700 , n33701 , n33702 , n33703 , n33704 , n33705 , n33706 , n33707 , n33708 , n33709 , n33710 , n33711 , n33712 , n33713 , n33714 , n33715 , n33716 , n33717 , n33718 , n33719 , n33720 , n33721 , n33722 , n33723 , n33724 , n33725 , n33726 , n33727 , n33728 , n33729 , n33730 , n33731 , n33732 , n33733 , n33734 , n33735 , n33736 , n33737 , n33738 , n33739 , n33740 , n33741 , n33742 , n33743 , n33744 , n33745 , n33746 , n33747 , n33748 , n33749 , n33750 , n33751 , n33752 , n33753 , n33754 , n33755 , n33756 , n33757 , n33758 , n33759 , n33760 , n33761 , n33762 , n33763 , n33764 , n33765 , n33766 , n33767 , n33768 , n33769 , n33770 , n33771 , n33772 , n33773 , n33774 , n33775 , n33776 , n33777 , n33778 , n33779 , n33780 , n33781 , n33782 , n33783 , n33784 , n33785 , n33786 , n33787 , n33788 , n33789 , n33790 , n33791 , n33792 , n33793 , n33794 , n33795 , n33796 , n33797 , n33798 , n33799 , n33800 , n33801 , n33802 , n33803 , n33804 , n33805 , n33806 , n33807 , n33808 , n33809 , n33810 , n33811 , n33812 , n33813 , n33814 , n33815 , n33816 , n33817 , n33818 , n33819 , n33820 , n33821 , n33822 , n33823 , n33824 , n33825 , n33826 , n33827 , n33828 , n33829 , n33830 , n33831 , n33832 , n33833 , n33834 , n33835 , n33836 , n33837 , n33838 , n33839 , n33840 , n33841 , n33842 , n33843 , n33844 , n33845 , n33846 , n33847 , n33848 , n33849 , n33850 , n33851 , n33852 , n33853 , n33854 , n33855 , n33856 , n33857 , n33858 , n33859 , n33860 , n33861 , n33862 , n33863 , n33864 , n33865 , n33866 , n33867 , n33868 , n33869 , n33870 , n33871 , n33872 , n33873 , n33874 , n33875 , n33876 , n33877 , n33878 , n33879 , n33880 , n33881 , n33882 , n33883 , n33884 , n33885 , n33886 , n33887 , n33888 , n33889 , n33890 , n33891 , n33892 , n33893 , n33894 , n33895 , n33896 , n33897 , n33898 , n33899 , n33900 , n33901 , n33902 , n33903 , n33904 , n33905 , n33906 , n33907 , n33908 , n33909 , n33910 , n33911 , n33912 , n33913 , n33914 , n33915 , n33916 , n33917 , n33918 , n33919 , n33920 , n33921 , n33922 , n33923 , n33924 , n33925 , n33926 , n33927 , n33928 , n33929 , n33930 , n33931 , n33932 , n33933 , n33934 , n33935 , n33936 , n33937 , n33938 , n33939 , n33940 , n33941 , n33942 , n33943 , n33944 , n33945 , n33946 , n33947 , n33948 , n33949 , n33950 , n33951 , n33952 , n33953 , n33954 , n33955 , n33956 , n33957 , n33958 , n33959 , n33960 , n33961 , n33962 , n33963 , n33964 , n33965 , n33966 , n33967 , n33968 , n33969 , n33970 , n33971 , n33972 , n33973 , n33974 , n33975 , n33976 , n33977 , n33978 , n33979 , n33980 , n33981 , n33982 , n33983 , n33984 , n33985 , n33986 , n33987 , n33988 , n33989 , n33990 , n33991 , n33992 , n33993 , n33994 , n33995 , n33996 , n33997 , n33998 , n33999 , n34000 , n34001 , n34002 , n34003 , n34004 , n34005 , n34006 , n34007 , n34008 , n34009 , n34010 , n34011 , n34012 , n34013 , n34014 , n34015 , n34016 , n34017 , n34018 , n34019 , n34020 , n34021 , n34022 , n34023 , n34024 , n34025 , n34026 , n34027 , n34028 , n34029 , n34030 , n34031 , n34032 , n34033 , n34034 , n34035 , n34036 , n34037 , n34038 , n34039 , n34040 , n34041 , n34042 , n34043 , n34044 , n34045 , n34046 , n34047 , n34048 , n34049 , n34050 , n34051 , n34052 , n34053 , n34054 , n34055 , n34056 , n34057 , n34058 , n34059 , n34060 , n34061 , n34062 , n34063 , n34064 , n34065 , n34066 , n34067 , n34068 , n34069 , n34070 , n34071 , n34072 , n34073 , n34074 , n34075 , n34076 , n34077 , n34078 , n34079 , n34080 , n34081 , n34082 , n34083 , n34084 , n34085 , n34086 , n34087 , n34088 , n34089 , n34090 , n34091 , n34092 , n34093 , n34094 , n34095 , n34096 , n34097 , n34098 , n34099 , n34100 , n34101 , n34102 , n34103 , n34104 , n34105 , n34106 , n34107 , n34108 , n34109 , n34110 , n34111 , n34112 , n34113 , n34114 , n34115 , n34116 , n34117 , n34118 , n34119 , n34120 , n34121 , n34122 , n34123 , n34124 , n34125 , n34126 , n34127 , n34128 , n34129 , n34130 , n34131 , n34132 , n34133 , n34134 , n34135 , n34136 , n34137 , n34138 , n34139 , n34140 , n34141 , n34142 , n34143 , n34144 , n34145 , n34146 , n34147 , n34148 , n34149 , n34150 , n34151 , n34152 , n34153 , n34154 , n34155 , n34156 , n34157 , n34158 , n34159 , n34160 , n34161 , n34162 , n34163 , n34164 , n34165 , n34166 , n34167 , n34168 , n34169 , n34170 , n34171 , n34172 , n34173 , n34174 , n34175 , n34176 , n34177 , n34178 , n34179 , n34180 , n34181 , n34182 , n34183 , n34184 , n34185 , n34186 , n34187 , n34188 , n34189 , n34190 , n34191 , n34192 , n34193 , n34194 , n34195 , n34196 , n34197 , n34198 , n34199 , n34200 , n34201 , n34202 , n34203 , n34204 , n34205 , n34206 , n34207 , n34208 , n34209 , n34210 , n34211 , n34212 , n34213 , n34214 , n34215 , n34216 , n34217 , n34218 , n34219 , n34220 , n34221 , n34222 , n34223 , n34224 , n34225 , n34226 , n34227 , n34228 , n34229 , n34230 , n34231 , n34232 , n34233 , n34234 , n34235 , n34236 , n34237 , n34238 , n34239 , n34240 , n34241 , n34242 , n34243 , n34244 , n34245 , n34246 , n34247 , n34248 , n34249 , n34250 , n34251 , n34252 , n34253 , n34254 , n34255 , n34256 , n34257 , n34258 , n34259 , n34260 , n34261 , n34262 , n34263 , n34264 , n34265 , n34266 , n34267 , n34268 , n34269 , n34270 , n34271 , n34272 , n34273 , n34274 , n34275 , n34276 , n34277 , n34278 , n34279 , n34280 , n34281 , n34282 , n34283 , n34284 , n34285 , n34286 , n34287 , n34288 , n34289 , n34290 , n34291 , n34292 , n34293 , n34294 , n34295 , n34296 , n34297 , n34298 , n34299 , n34300 , n34301 , n34302 , n34303 , n34304 , n34305 , n34306 , n34307 , n34308 , n34309 , n34310 , n34311 , n34312 , n34313 , n34314 , n34315 , n34316 , n34317 , n34318 , n34319 , n34320 , n34321 , n34322 , n34323 , n34324 , n34325 , n34326 , n34327 , n34328 , n34329 , n34330 , n34331 , n34332 , n34333 , n34334 , n34335 , n34336 , n34337 , n34338 , n34339 , n34340 , n34341 , n34342 , n34343 , n34344 , n34345 , n34346 , n34347 , n34348 , n34349 , n34350 , n34351 , n34352 , n34353 , n34354 , n34355 , n34356 , n34357 , n34358 , n34359 , n34360 , n34361 , n34362 , n34363 , n34364 , n34365 , n34366 , n34367 , n34368 , n34369 , n34370 , n34371 , n34372 , n34373 , n34374 , n34375 , n34376 , n34377 , n34378 , n34379 , n34380 , n34381 , n34382 , n34383 , n34384 , n34385 , n34386 , n34387 , n34388 , n34389 , n34390 , n34391 , n34392 , n34393 , n34394 , n34395 , n34396 , n34397 , n34398 , n34399 , n34400 , n34401 , n34402 , n34403 , n34404 , n34405 , n34406 , n34407 , n34408 , n34409 , n34410 , n34411 , n34412 , n34413 , n34414 , n34415 , n34416 , n34417 , n34418 , n34419 , n34420 , n34421 , n34422 , n34423 , n34424 , n34425 , n34426 , n34427 , n34428 , n34429 , n34430 , n34431 , n34432 , n34433 , n34434 , n34435 , n34436 , n34437 , n34438 , n34439 , n34440 , n34441 , n34442 , n34443 , n34444 , n34445 , n34446 , n34447 , n34448 , n34449 , n34450 , n34451 , n34452 , n34453 , n34454 , n34455 , n34456 , n34457 , n34458 , n34459 , n34460 , n34461 , n34462 , n34463 , n34464 , n34465 , n34466 , n34467 , n34468 , n34469 , n34470 , n34471 , n34472 , n34473 , n34474 , n34475 , n34476 , n34477 , n34478 , n34479 , n34480 , n34481 , n34482 , n34483 , n34484 , n34485 , n34486 , n34487 , n34488 , n34489 , n34490 , n34491 , n34492 , n34493 , n34494 , n34495 , n34496 , n34497 , n34498 , n34499 , n34500 , n34501 , n34502 , n34503 , n34504 , n34505 , n34506 , n34507 , n34508 , n34509 , n34510 , n34511 , n34512 , n34513 , n34514 , n34515 , n34516 , n34517 , n34518 , n34519 , n34520 , n34521 , n34522 , n34523 , n34524 , n34525 , n34526 , n34527 , n34528 , n34529 , n34530 , n34531 , n34532 , n34533 , n34534 , n34535 , n34536 , n34537 , n34538 , n34539 , n34540 , n34541 , n34542 , n34543 , n34544 , n34545 , n34546 , n34547 , n34548 , n34549 , n34550 , n34551 , n34552 , n34553 , n34554 , n34555 , n34556 , n34557 , n34558 , n34559 , n34560 , n34561 , n34562 , n34563 , n34564 , n34565 , n34566 , n34567 , n34568 , n34569 , n34570 , n34571 , n34572 , n34573 , n34574 , n34575 , n34576 , n34577 , n34578 , n34579 , n34580 , n34581 , n34582 , n34583 , n34584 , n34585 , n34586 , n34587 , n34588 , n34589 , n34590 , n34591 , n34592 , n34593 , n34594 , n34595 , n34596 , n34597 , n34598 , n34599 , n34600 , n34601 , n34602 , n34603 , n34604 , n34605 , n34606 , n34607 , n34608 , n34609 , n34610 , n34611 , n34612 , n34613 , n34614 , n34615 , n34616 , n34617 , n34618 , n34619 , n34620 , n34621 , n34622 , n34623 , n34624 , n34625 , n34626 , n34627 , n34628 , n34629 , n34630 , n34631 , n34632 , n34633 , n34634 , n34635 , n34636 , n34637 , n34638 , n34639 , n34640 , n34641 , n34642 , n34643 , n34644 , n34645 , n34646 , n34647 , n34648 , n34649 , n34650 , n34651 , n34652 , n34653 , n34654 , n34655 , n34656 , n34657 , n34658 , n34659 , n34660 , n34661 , n34662 , n34663 , n34664 , n34665 , n34666 , n34667 , n34668 , n34669 , n34670 , n34671 , n34672 , n34673 , n34674 , n34675 , n34676 , n34677 , n34678 , n34679 , n34680 , n34681 , n34682 , n34683 , n34684 , n34685 , n34686 , n34687 , n34688 , n34689 , n34690 , n34691 , n34692 , n34693 , n34694 , n34695 , n34696 , n34697 , n34698 , n34699 , n34700 , n34701 , n34702 , n34703 , n34704 , n34705 , n34706 , n34707 , n34708 , n34709 , n34710 , n34711 , n34712 , n34713 , n34714 , n34715 , n34716 , n34717 , n34718 , n34719 , n34720 , n34721 , n34722 , n34723 , n34724 , n34725 , n34726 , n34727 , n34728 , n34729 , n34730 , n34731 , n34732 , n34733 , n34734 , n34735 , n34736 , n34737 , n34738 , n34739 , n34740 , n34741 , n34742 , n34743 , n34744 , n34745 , n34746 , n34747 , n34748 , n34749 , n34750 , n34751 , n34752 , n34753 , n34754 , n34755 , n34756 , n34757 , n34758 , n34759 , n34760 , n34761 , n34762 , n34763 , n34764 , n34765 , n34766 , n34767 , n34768 , n34769 , n34770 , n34771 , n34772 , n34773 , n34774 , n34775 , n34776 , n34777 , n34778 , n34779 , n34780 , n34781 , n34782 , n34783 , n34784 , n34785 , n34786 , n34787 , n34788 , n34789 , n34790 , n34791 , n34792 , n34793 , n34794 , n34795 , n34796 , n34797 , n34798 , n34799 , n34800 , n34801 , n34802 , n34803 , n34804 , n34805 , n34806 , n34807 , n34808 , n34809 , n34810 , n34811 , n34812 , n34813 , n34814 , n34815 , n34816 , n34817 , n34818 , n34819 , n34820 , n34821 , n34822 , n34823 , n34824 , n34825 , n34826 , n34827 , n34828 , n34829 , n34830 , n34831 , n34832 , n34833 , n34834 , n34835 , n34836 , n34837 , n34838 , n34839 , n34840 , n34841 , n34842 , n34843 , n34844 , n34845 , n34846 , n34847 , n34848 , n34849 , n34850 , n34851 , n34852 , n34853 , n34854 , n34855 , n34856 , n34857 , n34858 , n34859 , n34860 , n34861 , n34862 , n34863 , n34864 , n34865 , n34866 , n34867 , n34868 , n34869 , n34870 , n34871 , n34872 , n34873 , n34874 , n34875 , n34876 , n34877 , n34878 , n34879 , n34880 , n34881 , n34882 , n34883 , n34884 , n34885 , n34886 , n34887 , n34888 , n34889 , n34890 , n34891 , n34892 , n34893 , n34894 , n34895 , n34896 , n34897 , n34898 , n34899 , n34900 , n34901 , n34902 , n34903 , n34904 , n34905 , n34906 , n34907 , n34908 , n34909 , n34910 , n34911 , n34912 , n34913 , n34914 , n34915 , n34916 , n34917 , n34918 , n34919 , n34920 , n34921 , n34922 , n34923 , n34924 , n34925 , n34926 , n34927 , n34928 , n34929 , n34930 , n34931 , n34932 , n34933 , n34934 , n34935 , n34936 , n34937 , n34938 , n34939 , n34940 , n34941 , n34942 , n34943 , n34944 , n34945 , n34946 , n34947 , n34948 , n34949 , n34950 , n34951 , n34952 , n34953 , n34954 , n34955 , n34956 , n34957 , n34958 , n34959 , n34960 , n34961 , n34962 , n34963 , n34964 , n34965 , n34966 , n34967 , n34968 , n34969 , n34970 , n34971 , n34972 , n34973 , n34974 , n34975 , n34976 , n34977 , n34978 , n34979 , n34980 , n34981 , n34982 , n34983 , n34984 , n34985 , n34986 , n34987 , n34988 , n34989 , n34990 , n34991 , n34992 , n34993 , n34994 , n34995 , n34996 , n34997 , n34998 , n34999 , n35000 , n35001 , n35002 , n35003 , n35004 , n35005 , n35006 , n35007 , n35008 , n35009 , n35010 , n35011 , n35012 , n35013 , n35014 , n35015 , n35016 , n35017 , n35018 , n35019 , n35020 , n35021 , n35022 , n35023 , n35024 , n35025 , n35026 , n35027 , n35028 , n35029 , n35030 , n35031 , n35032 , n35033 , n35034 , n35035 , n35036 , n35037 , n35038 , n35039 , n35040 , n35041 , n35042 , n35043 , n35044 , n35045 , n35046 , n35047 , n35048 , n35049 , n35050 , n35051 , n35052 , n35053 , n35054 , n35055 , n35056 , n35057 , n35058 , n35059 , n35060 , n35061 , n35062 , n35063 , n35064 , n35065 , n35066 , n35067 , n35068 , n35069 , n35070 , n35071 , n35072 , n35073 , n35074 , n35075 , n35076 , n35077 , n35078 , n35079 , n35080 , n35081 , n35082 , n35083 , n35084 , n35085 , n35086 , n35087 , n35088 , n35089 , n35090 , n35091 , n35092 , n35093 , n35094 , n35095 , n35096 , n35097 , n35098 , n35099 , n35100 , n35101 , n35102 , n35103 , n35104 , n35105 , n35106 , n35107 , n35108 , n35109 , n35110 , n35111 , n35112 , n35113 , n35114 , n35115 , n35116 , n35117 , n35118 , n35119 , n35120 , n35121 , n35122 , n35123 , n35124 , n35125 , n35126 , n35127 , n35128 , n35129 , n35130 , n35131 , n35132 , n35133 , n35134 , n35135 , n35136 , n35137 , n35138 , n35139 , n35140 , n35141 , n35142 , n35143 , n35144 , n35145 , n35146 , n35147 , n35148 , n35149 , n35150 , n35151 , n35152 , n35153 , n35154 , n35155 , n35156 , n35157 , n35158 , n35159 , n35160 , n35161 , n35162 , n35163 , n35164 , n35165 , n35166 , n35167 , n35168 , n35169 , n35170 , n35171 , n35172 , n35173 , n35174 , n35175 , n35176 , n35177 , n35178 , n35179 , n35180 , n35181 , n35182 , n35183 , n35184 , n35185 , n35186 , n35187 , n35188 , n35189 , n35190 , n35191 , n35192 , n35193 , n35194 , n35195 , n35196 , n35197 , n35198 , n35199 , n35200 , n35201 , n35202 , n35203 , n35204 , n35205 , n35206 , n35207 , n35208 , n35209 , n35210 , n35211 , n35212 , n35213 , n35214 , n35215 , n35216 , n35217 , n35218 , n35219 , n35220 , n35221 , n35222 , n35223 , n35224 , n35225 , n35226 , n35227 , n35228 , n35229 , n35230 , n35231 , n35232 , n35233 , n35234 , n35235 , n35236 , n35237 , n35238 , n35239 , n35240 , n35241 , n35242 , n35243 , n35244 , n35245 , n35246 , n35247 , n35248 , n35249 , n35250 , n35251 , n35252 , n35253 , n35254 , n35255 , n35256 , n35257 , n35258 , n35259 , n35260 , n35261 , n35262 , n35263 , n35264 , n35265 , n35266 , n35267 , n35268 , n35269 , n35270 , n35271 , n35272 , n35273 , n35274 , n35275 , n35276 , n35277 , n35278 , n35279 , n35280 , n35281 , n35282 , n35283 , n35284 , n35285 , n35286 , n35287 , n35288 , n35289 , n35290 , n35291 , n35292 , n35293 , n35294 , n35295 , n35296 , n35297 , n35298 , n35299 , n35300 , n35301 , n35302 , n35303 , n35304 , n35305 , n35306 , n35307 , n35308 , n35309 , n35310 , n35311 , n35312 , n35313 , n35314 , n35315 , n35316 , n35317 , n35318 , n35319 , n35320 , n35321 , n35322 , n35323 , n35324 , n35325 , n35326 , n35327 , n35328 , n35329 , n35330 , n35331 , n35332 , n35333 , n35334 , n35335 , n35336 , n35337 , n35338 , n35339 , n35340 , n35341 , n35342 , n35343 , n35344 , n35345 , n35346 , n35347 , n35348 , n35349 , n35350 , n35351 , n35352 , n35353 , n35354 , n35355 , n35356 , n35357 , n35358 , n35359 , n35360 , n35361 , n35362 , n35363 , n35364 , n35365 , n35366 , n35367 , n35368 , n35369 , n35370 , n35371 , n35372 , n35373 , n35374 , n35375 , n35376 , n35377 , n35378 , n35379 , n35380 , n35381 , n35382 , n35383 , n35384 , n35385 , n35386 , n35387 , n35388 , n35389 , n35390 , n35391 , n35392 , n35393 , n35394 , n35395 , n35396 , n35397 , n35398 , n35399 , n35400 , n35401 , n35402 , n35403 , n35404 , n35405 , n35406 , n35407 , n35408 , n35409 , n35410 , n35411 , n35412 , n35413 , n35414 , n35415 , n35416 , n35417 , n35418 , n35419 , n35420 , n35421 , n35422 , n35423 , n35424 , n35425 , n35426 , n35427 , n35428 , n35429 , n35430 , n35431 , n35432 , n35433 , n35434 , n35435 , n35436 , n35437 , n35438 , n35439 , n35440 , n35441 , n35442 , n35443 , n35444 , n35445 , n35446 , n35447 , n35448 , n35449 , n35450 , n35451 , n35452 , n35453 , n35454 , n35455 , n35456 , n35457 , n35458 , n35459 , n35460 , n35461 , n35462 , n35463 , n35464 , n35465 , n35466 , n35467 , n35468 , n35469 , n35470 , n35471 , n35472 , n35473 , n35474 , n35475 , n35476 , n35477 , n35478 , n35479 , n35480 , n35481 , n35482 , n35483 , n35484 , n35485 , n35486 , n35487 , n35488 , n35489 , n35490 , n35491 , n35492 , n35493 , n35494 , n35495 , n35496 , n35497 , n35498 , n35499 , n35500 , n35501 , n35502 , n35503 , n35504 , n35505 , n35506 , n35507 , n35508 , n35509 , n35510 , n35511 , n35512 , n35513 , n35514 , n35515 , n35516 , n35517 , n35518 , n35519 , n35520 , n35521 , n35522 , n35523 , n35524 , n35525 , n35526 , n35527 , n35528 , n35529 , n35530 , n35531 , n35532 , n35533 , n35534 , n35535 , n35536 , n35537 , n35538 , n35539 , n35540 , n35541 , n35542 , n35543 , n35544 , n35545 , n35546 , n35547 , n35548 , n35549 , n35550 , n35551 , n35552 , n35553 , n35554 , n35555 , n35556 , n35557 , n35558 , n35559 , n35560 , n35561 , n35562 , n35563 , n35564 , n35565 , n35566 , n35567 , n35568 , n35569 , n35570 , n35571 , n35572 , n35573 , n35574 , n35575 , n35576 , n35577 , n35578 , n35579 , n35580 , n35581 , n35582 , n35583 , n35584 , n35585 , n35586 , n35587 , n35588 , n35589 , n35590 , n35591 , n35592 , n35593 , n35594 , n35595 , n35596 , n35597 , n35598 , n35599 , n35600 , n35601 , n35602 , n35603 , n35604 , n35605 , n35606 , n35607 , n35608 , n35609 , n35610 , n35611 , n35612 , n35613 , n35614 , n35615 , n35616 , n35617 , n35618 , n35619 , n35620 , n35621 , n35622 , n35623 , n35624 , n35625 , n35626 , n35627 , n35628 , n35629 , n35630 , n35631 , n35632 , n35633 , n35634 , n35635 , n35636 , n35637 , n35638 , n35639 , n35640 , n35641 , n35642 , n35643 , n35644 , n35645 , n35646 , n35647 , n35648 , n35649 , n35650 , n35651 , n35652 , n35653 , n35654 , n35655 , n35656 , n35657 , n35658 , n35659 , n35660 , n35661 , n35662 , n35663 , n35664 , n35665 , n35666 , n35667 , n35668 , n35669 , n35670 , n35671 , n35672 , n35673 , n35674 , n35675 , n35676 , n35677 , n35678 , n35679 , n35680 , n35681 , n35682 , n35683 , n35684 , n35685 , n35686 , n35687 , n35688 , n35689 , n35690 , n35691 , n35692 , n35693 , n35694 , n35695 , n35696 , n35697 , n35698 , n35699 , n35700 , n35701 , n35702 , n35703 , n35704 , n35705 , n35706 , n35707 , n35708 , n35709 , n35710 , n35711 , n35712 , n35713 , n35714 , n35715 , n35716 , n35717 , n35718 , n35719 , n35720 , n35721 , n35722 , n35723 , n35724 , n35725 , n35726 , n35727 , n35728 , n35729 , n35730 , n35731 , n35732 , n35733 , n35734 , n35735 , n35736 , n35737 , n35738 , n35739 , n35740 , n35741 , n35742 , n35743 , n35744 , n35745 , n35746 , n35747 , n35748 , n35749 , n35750 , n35751 , n35752 , n35753 , n35754 , n35755 , n35756 , n35757 , n35758 , n35759 , n35760 , n35761 , n35762 , n35763 , n35764 , n35765 , n35766 , n35767 , n35768 , n35769 , n35770 , n35771 , n35772 , n35773 , n35774 , n35775 , n35776 , n35777 , n35778 , n35779 , n35780 , n35781 , n35782 , n35783 , n35784 , n35785 , n35786 , n35787 , n35788 , n35789 , n35790 , n35791 , n35792 , n35793 , n35794 , n35795 , n35796 , n35797 , n35798 , n35799 , n35800 , n35801 , n35802 , n35803 , n35804 , n35805 , n35806 , n35807 , n35808 , n35809 , n35810 , n35811 , n35812 , n35813 , n35814 , n35815 , n35816 , n35817 , n35818 , n35819 , n35820 , n35821 , n35822 , n35823 , n35824 , n35825 , n35826 , n35827 , n35828 , n35829 , n35830 , n35831 , n35832 , n35833 , n35834 , n35835 , n35836 , n35837 , n35838 , n35839 , n35840 , n35841 , n35842 , n35843 , n35844 , n35845 , n35846 , n35847 , n35848 , n35849 , n35850 , n35851 , n35852 , n35853 , n35854 , n35855 , n35856 , n35857 , n35858 , n35859 , n35860 , n35861 , n35862 , n35863 , n35864 , n35865 , n35866 , n35867 , n35868 , n35869 , n35870 , n35871 , n35872 , n35873 , n35874 , n35875 , n35876 , n35877 , n35878 , n35879 , n35880 , n35881 , n35882 , n35883 , n35884 , n35885 , n35886 , n35887 , n35888 , n35889 , n35890 , n35891 , n35892 , n35893 , n35894 , n35895 , n35896 , n35897 , n35898 , n35899 , n35900 , n35901 , n35902 , n35903 , n35904 , n35905 , n35906 , n35907 , n35908 , n35909 , n35910 , n35911 , n35912 , n35913 , n35914 , n35915 , n35916 , n35917 , n35918 , n35919 , n35920 , n35921 , n35922 , n35923 , n35924 , n35925 , n35926 , n35927 , n35928 , n35929 , n35930 , n35931 , n35932 , n35933 , n35934 , n35935 , n35936 , n35937 , n35938 , n35939 , n35940 , n35941 , n35942 , n35943 , n35944 , n35945 , n35946 , n35947 , n35948 , n35949 , n35950 , n35951 , n35952 , n35953 , n35954 , n35955 , n35956 , n35957 , n35958 , n35959 , n35960 , n35961 , n35962 , n35963 , n35964 , n35965 , n35966 , n35967 , n35968 , n35969 , n35970 , n35971 , n35972 , n35973 , n35974 , n35975 , n35976 , n35977 , n35978 , n35979 , n35980 , n35981 , n35982 , n35983 , n35984 , n35985 , n35986 , n35987 , n35988 , n35989 , n35990 , n35991 , n35992 , n35993 , n35994 , n35995 , n35996 , n35997 , n35998 , n35999 , n36000 , n36001 , n36002 , n36003 , n36004 , n36005 , n36006 , n36007 , n36008 , n36009 , n36010 , n36011 , n36012 , n36013 , n36014 , n36015 , n36016 , n36017 , n36018 , n36019 , n36020 , n36021 , n36022 , n36023 , n36024 , n36025 , n36026 , n36027 , n36028 , n36029 , n36030 , n36031 , n36032 , n36033 , n36034 , n36035 , n36036 , n36037 , n36038 , n36039 , n36040 , n36041 , n36042 , n36043 , n36044 , n36045 , n36046 , n36047 , n36048 , n36049 , n36050 , n36051 , n36052 , n36053 , n36054 , n36055 , n36056 , n36057 , n36058 , n36059 , n36060 , n36061 , n36062 , n36063 , n36064 , n36065 , n36066 , n36067 , n36068 , n36069 , n36070 , n36071 , n36072 , n36073 , n36074 , n36075 , n36076 , n36077 , n36078 , n36079 , n36080 , n36081 , n36082 , n36083 , n36084 , n36085 , n36086 , n36087 , n36088 , n36089 , n36090 , n36091 , n36092 , n36093 , n36094 , n36095 , n36096 , n36097 , n36098 , n36099 , n36100 , n36101 , n36102 , n36103 , n36104 , n36105 , n36106 , n36107 , n36108 , n36109 , n36110 , n36111 , n36112 , n36113 , n36114 , n36115 , n36116 , n36117 , n36118 , n36119 , n36120 , n36121 , n36122 , n36123 , n36124 , n36125 , n36126 , n36127 , n36128 , n36129 , n36130 , n36131 , n36132 , n36133 , n36134 , n36135 , n36136 , n36137 , n36138 , n36139 , n36140 , n36141 , n36142 , n36143 , n36144 , n36145 , n36146 , n36147 , n36148 , n36149 , n36150 , n36151 , n36152 , n36153 , n36154 , n36155 , n36156 , n36157 , n36158 , n36159 , n36160 , n36161 , n36162 , n36163 , n36164 , n36165 , n36166 , n36167 , n36168 , n36169 , n36170 , n36171 , n36172 , n36173 , n36174 , n36175 , n36176 , n36177 , n36178 , n36179 , n36180 , n36181 , n36182 , n36183 , n36184 , n36185 , n36186 , n36187 , n36188 , n36189 , n36190 , n36191 , n36192 , n36193 , n36194 , n36195 , n36196 , n36197 , n36198 , n36199 , n36200 , n36201 , n36202 , n36203 , n36204 , n36205 , n36206 , n36207 , n36208 , n36209 , n36210 , n36211 , n36212 , n36213 , n36214 , n36215 , n36216 , n36217 , n36218 , n36219 , n36220 , n36221 , n36222 , n36223 , n36224 , n36225 , n36226 , n36227 , n36228 , n36229 , n36230 , n36231 , n36232 , n36233 , n36234 , n36235 , n36236 , n36237 , n36238 , n36239 , n36240 , n36241 , n36242 , n36243 , n36244 , n36245 , n36246 , n36247 , n36248 , n36249 , n36250 , n36251 , n36252 , n36253 , n36254 , n36255 , n36256 , n36257 , n36258 , n36259 , n36260 , n36261 , n36262 , n36263 , n36264 , n36265 , n36266 , n36267 , n36268 , n36269 , n36270 , n36271 , n36272 , n36273 , n36274 , n36275 , n36276 , n36277 , n36278 , n36279 , n36280 , n36281 , n36282 , n36283 , n36284 , n36285 , n36286 , n36287 , n36288 , n36289 , n36290 , n36291 , n36292 , n36293 , n36294 , n36295 , n36296 , n36297 , n36298 , n36299 , n36300 , n36301 , n36302 , n36303 , n36304 , n36305 , n36306 , n36307 , n36308 , n36309 , n36310 , n36311 , n36312 , n36313 , n36314 , n36315 , n36316 , n36317 , n36318 , n36319 , n36320 , n36321 , n36322 , n36323 , n36324 , n36325 , n36326 , n36327 , n36328 , n36329 , n36330 , n36331 , n36332 , n36333 , n36334 , n36335 , n36336 , n36337 , n36338 , n36339 , n36340 , n36341 , n36342 , n36343 , n36344 , n36345 , n36346 , n36347 , n36348 , n36349 , n36350 , n36351 , n36352 , n36353 , n36354 , n36355 , n36356 , n36357 , n36358 , n36359 , n36360 , n36361 , n36362 , n36363 , n36364 , n36365 , n36366 , n36367 , n36368 , n36369 , n36370 , n36371 , n36372 , n36373 , n36374 , n36375 , n36376 , n36377 , n36378 , n36379 , n36380 , n36381 , n36382 , n36383 , n36384 , n36385 , n36386 , n36387 , n36388 , n36389 , n36390 , n36391 , n36392 , n36393 , n36394 , n36395 , n36396 , n36397 , n36398 , n36399 , n36400 , n36401 , n36402 , n36403 , n36404 , n36405 , n36406 , n36407 , n36408 , n36409 , n36410 , n36411 , n36412 , n36413 , n36414 , n36415 , n36416 , n36417 , n36418 , n36419 , n36420 , n36421 , n36422 , n36423 , n36424 , n36425 , n36426 , n36427 , n36428 , n36429 , n36430 , n36431 , n36432 , n36433 , n36434 , n36435 , n36436 , n36437 , n36438 , n36439 , n36440 , n36441 , n36442 , n36443 , n36444 , n36445 , n36446 , n36447 , n36448 , n36449 , n36450 , n36451 , n36452 , n36453 , n36454 , n36455 , n36456 , n36457 , n36458 , n36459 , n36460 , n36461 , n36462 , n36463 , n36464 , n36465 , n36466 , n36467 , n36468 , n36469 , n36470 , n36471 , n36472 , n36473 , n36474 , n36475 , n36476 , n36477 , n36478 , n36479 , n36480 , n36481 , n36482 , n36483 , n36484 , n36485 , n36486 , n36487 , n36488 , n36489 , n36490 , n36491 , n36492 , n36493 , n36494 , n36495 , n36496 , n36497 , n36498 , n36499 , n36500 , n36501 , n36502 , n36503 , n36504 , n36505 , n36506 , n36507 , n36508 , n36509 , n36510 , n36511 , n36512 , n36513 , n36514 , n36515 , n36516 , n36517 , n36518 , n36519 , n36520 , n36521 , n36522 , n36523 , n36524 , n36525 , n36526 , n36527 , n36528 , n36529 , n36530 , n36531 , n36532 , n36533 , n36534 , n36535 , n36536 , n36537 , n36538 , n36539 , n36540 , n36541 , n36542 , n36543 , n36544 , n36545 , n36546 , n36547 , n36548 , n36549 , n36550 , n36551 , n36552 , n36553 , n36554 , n36555 , n36556 , n36557 , n36558 , n36559 , n36560 , n36561 , n36562 , n36563 , n36564 , n36565 , n36566 , n36567 , n36568 , n36569 , n36570 , n36571 , n36572 , n36573 , n36574 , n36575 , n36576 , n36577 , n36578 , n36579 , n36580 , n36581 , n36582 , n36583 , n36584 , n36585 , n36586 , n36587 , n36588 , n36589 , n36590 , n36591 , n36592 , n36593 , n36594 , n36595 , n36596 , n36597 , n36598 , n36599 , n36600 , n36601 , n36602 , n36603 , n36604 , n36605 , n36606 , n36607 , n36608 , n36609 , n36610 , n36611 , n36612 , n36613 , n36614 , n36615 , n36616 , n36617 , n36618 , n36619 , n36620 , n36621 , n36622 , n36623 , n36624 , n36625 , n36626 , n36627 , n36628 , n36629 , n36630 , n36631 , n36632 , n36633 , n36634 , n36635 , n36636 , n36637 , n36638 , n36639 , n36640 , n36641 , n36642 , n36643 , n36644 , n36645 , n36646 , n36647 , n36648 , n36649 , n36650 , n36651 , n36652 , n36653 , n36654 , n36655 , n36656 , n36657 , n36658 , n36659 , n36660 , n36661 , n36662 , n36663 , n36664 , n36665 , n36666 , n36667 , n36668 , n36669 , n36670 , n36671 , n36672 , n36673 , n36674 , n36675 , n36676 , n36677 , n36678 , n36679 , n36680 , n36681 , n36682 , n36683 , n36684 , n36685 , n36686 , n36687 , n36688 , n36689 , n36690 , n36691 , n36692 , n36693 , n36694 , n36695 , n36696 , n36697 , n36698 , n36699 , n36700 , n36701 , n36702 , n36703 , n36704 , n36705 , n36706 , n36707 , n36708 , n36709 , n36710 , n36711 , n36712 , n36713 , n36714 , n36715 , n36716 , n36717 , n36718 , n36719 , n36720 , n36721 , n36722 , n36723 , n36724 , n36725 , n36726 , n36727 , n36728 , n36729 , n36730 , n36731 , n36732 , n36733 , n36734 , n36735 , n36736 , n36737 , n36738 , n36739 , n36740 , n36741 , n36742 , n36743 , n36744 , n36745 , n36746 , n36747 , n36748 , n36749 , n36750 , n36751 , n36752 , n36753 , n36754 , n36755 , n36756 , n36757 , n36758 , n36759 , n36760 , n36761 , n36762 , n36763 , n36764 , n36765 , n36766 , n36767 , n36768 , n36769 , n36770 , n36771 , n36772 , n36773 , n36774 , n36775 , n36776 , n36777 , n36778 , n36779 , n36780 , n36781 , n36782 , n36783 , n36784 , n36785 , n36786 , n36787 , n36788 , n36789 , n36790 , n36791 , n36792 , n36793 , n36794 , n36795 , n36796 , n36797 , n36798 , n36799 , n36800 , n36801 , n36802 , n36803 , n36804 , n36805 , n36806 , n36807 , n36808 , n36809 , n36810 , n36811 , n36812 , n36813 , n36814 , n36815 , n36816 , n36817 , n36818 , n36819 , n36820 , n36821 , n36822 , n36823 , n36824 , n36825 , n36826 , n36827 , n36828 , n36829 , n36830 , n36831 , n36832 , n36833 , n36834 , n36835 , n36836 , n36837 , n36838 , n36839 , n36840 , n36841 , n36842 , n36843 , n36844 , n36845 , n36846 , n36847 , n36848 , n36849 , n36850 , n36851 , n36852 , n36853 , n36854 , n36855 , n36856 , n36857 , n36858 , n36859 , n36860 , n36861 , n36862 , n36863 , n36864 , n36865 , n36866 , n36867 , n36868 , n36869 , n36870 , n36871 , n36872 , n36873 , n36874 , n36875 , n36876 , n36877 , n36878 , n36879 , n36880 , n36881 , n36882 , n36883 , n36884 , n36885 , n36886 , n36887 , n36888 , n36889 , n36890 , n36891 , n36892 , n36893 , n36894 , n36895 , n36896 , n36897 , n36898 , n36899 , n36900 , n36901 , n36902 , n36903 , n36904 , n36905 , n36906 , n36907 , n36908 , n36909 , n36910 , n36911 , n36912 , n36913 , n36914 , n36915 , n36916 , n36917 , n36918 , n36919 , n36920 , n36921 , n36922 , n36923 , n36924 , n36925 , n36926 , n36927 , n36928 , n36929 , n36930 , n36931 , n36932 , n36933 , n36934 , n36935 , n36936 , n36937 , n36938 , n36939 , n36940 , n36941 , n36942 , n36943 , n36944 , n36945 , n36946 , n36947 , n36948 , n36949 , n36950 , n36951 , n36952 , n36953 , n36954 , n36955 , n36956 , n36957 , n36958 , n36959 , n36960 , n36961 , n36962 , n36963 , n36964 , n36965 , n36966 , n36967 , n36968 , n36969 , n36970 , n36971 , n36972 , n36973 , n36974 , n36975 , n36976 , n36977 , n36978 , n36979 , n36980 , n36981 , n36982 , n36983 , n36984 , n36985 , n36986 , n36987 , n36988 , n36989 , n36990 , n36991 , n36992 , n36993 , n36994 , n36995 , n36996 , n36997 , n36998 , n36999 , n37000 , n37001 , n37002 , n37003 , n37004 , n37005 , n37006 , n37007 , n37008 , n37009 , n37010 , n37011 , n37012 , n37013 , n37014 , n37015 , n37016 , n37017 , n37018 , n37019 , n37020 , n37021 , n37022 , n37023 , n37024 , n37025 , n37026 , n37027 , n37028 , n37029 , n37030 , n37031 , n37032 , n37033 , n37034 , n37035 , n37036 , n37037 , n37038 , n37039 , n37040 , n37041 , n37042 , n37043 , n37044 , n37045 , n37046 , n37047 , n37048 , n37049 , n37050 , n37051 , n37052 , n37053 , n37054 , n37055 , n37056 , n37057 , n37058 , n37059 , n37060 , n37061 , n37062 , n37063 , n37064 , n37065 , n37066 , n37067 , n37068 , n37069 , n37070 , n37071 , n37072 , n37073 , n37074 , n37075 , n37076 , n37077 , n37078 , n37079 , n37080 , n37081 , n37082 , n37083 , n37084 , n37085 , n37086 , n37087 , n37088 , n37089 , n37090 , n37091 , n37092 , n37093 , n37094 , n37095 , n37096 , n37097 , n37098 , n37099 , n37100 , n37101 , n37102 , n37103 , n37104 , n37105 , n37106 , n37107 , n37108 , n37109 , n37110 , n37111 , n37112 , n37113 , n37114 , n37115 , n37116 , n37117 , n37118 , n37119 , n37120 , n37121 , n37122 , n37123 , n37124 , n37125 , n37126 , n37127 , n37128 , n37129 , n37130 , n37131 , n37132 , n37133 , n37134 , n37135 , n37136 , n37137 , n37138 , n37139 , n37140 , n37141 , n37142 , n37143 , n37144 , n37145 , n37146 , n37147 , n37148 , n37149 , n37150 , n37151 , n37152 , n37153 , n37154 , n37155 , n37156 , n37157 , n37158 , n37159 , n37160 , n37161 , n37162 , n37163 , n37164 , n37165 , n37166 , n37167 , n37168 , n37169 , n37170 , n37171 , n37172 , n37173 , n37174 , n37175 , n37176 , n37177 , n37178 , n37179 , n37180 , n37181 , n37182 , n37183 , n37184 , n37185 , n37186 , n37187 , n37188 , n37189 , n37190 , n37191 , n37192 , n37193 , n37194 , n37195 , n37196 , n37197 , n37198 , n37199 , n37200 , n37201 , n37202 , n37203 , n37204 , n37205 , n37206 , n37207 , n37208 , n37209 , n37210 , n37211 , n37212 , n37213 , n37214 , n37215 , n37216 , n37217 , n37218 , n37219 , n37220 , n37221 , n37222 , n37223 , n37224 , n37225 , n37226 , n37227 , n37228 , n37229 , n37230 , n37231 , n37232 , n37233 , n37234 , n37235 , n37236 , n37237 , n37238 , n37239 , n37240 , n37241 , n37242 , n37243 , n37244 , n37245 , n37246 , n37247 , n37248 , n37249 , n37250 , n37251 , n37252 , n37253 , n37254 , n37255 , n37256 , n37257 , n37258 , n37259 , n37260 , n37261 , n37262 , n37263 , n37264 , n37265 , n37266 , n37267 , n37268 , n37269 , n37270 , n37271 , n37272 , n37273 , n37274 , n37275 , n37276 , n37277 , n37278 , n37279 , n37280 , n37281 , n37282 , n37283 , n37284 , n37285 , n37286 , n37287 , n37288 , n37289 , n37290 , n37291 , n37292 , n37293 , n37294 , n37295 , n37296 , n37297 , n37298 , n37299 , n37300 , n37301 , n37302 , n37303 , n37304 , n37305 , n37306 , n37307 , n37308 , n37309 , n37310 , n37311 , n37312 , n37313 , n37314 , n37315 , n37316 , n37317 , n37318 , n37319 , n37320 , n37321 , n37322 , n37323 , n37324 , n37325 , n37326 , n37327 , n37328 , n37329 , n37330 , n37331 , n37332 , n37333 , n37334 , n37335 , n37336 , n37337 , n37338 , n37339 , n37340 , n37341 , n37342 , n37343 , n37344 , n37345 , n37346 , n37347 , n37348 , n37349 , n37350 , n37351 , n37352 , n37353 , n37354 , n37355 , n37356 , n37357 , n37358 , n37359 , n37360 , n37361 , n37362 , n37363 , n37364 , n37365 , n37366 , n37367 , n37368 , n37369 , n37370 , n37371 , n37372 , n37373 , n37374 , n37375 , n37376 , n37377 , n37378 , n37379 , n37380 , n37381 , n37382 , n37383 , n37384 , n37385 , n37386 , n37387 , n37388 , n37389 , n37390 , n37391 , n37392 , n37393 , n37394 , n37395 , n37396 , n37397 , n37398 , n37399 , n37400 , n37401 , n37402 , n37403 , n37404 , n37405 , n37406 , n37407 , n37408 , n37409 , n37410 , n37411 , n37412 , n37413 , n37414 , n37415 , n37416 , n37417 , n37418 , n37419 , n37420 , n37421 , n37422 , n37423 , n37424 , n37425 , n37426 , n37427 , n37428 , n37429 , n37430 , n37431 , n37432 , n37433 , n37434 , n37435 , n37436 , n37437 , n37438 , n37439 , n37440 , n37441 , n37442 , n37443 , n37444 , n37445 , n37446 , n37447 , n37448 , n37449 , n37450 , n37451 , n37452 , n37453 , n37454 , n37455 , n37456 , n37457 , n37458 , n37459 , n37460 , n37461 , n37462 , n37463 , n37464 , n37465 , n37466 , n37467 , n37468 , n37469 , n37470 , n37471 , n37472 , n37473 , n37474 , n37475 , n37476 , n37477 , n37478 , n37479 , n37480 , n37481 , n37482 , n37483 , n37484 , n37485 , n37486 , n37487 , n37488 , n37489 , n37490 , n37491 , n37492 , n37493 , n37494 , n37495 , n37496 , n37497 , n37498 , n37499 , n37500 , n37501 , n37502 , n37503 , n37504 , n37505 , n37506 , n37507 , n37508 , n37509 , n37510 , n37511 , n37512 , n37513 , n37514 , n37515 , n37516 , n37517 , n37518 , n37519 , n37520 , n37521 , n37522 , n37523 , n37524 , n37525 , n37526 , n37527 , n37528 , n37529 , n37530 , n37531 , n37532 , n37533 , n37534 , n37535 , n37536 , n37537 , n37538 , n37539 , n37540 , n37541 , n37542 , n37543 , n37544 , n37545 , n37546 , n37547 , n37548 , n37549 , n37550 , n37551 , n37552 , n37553 , n37554 , n37555 , n37556 , n37557 , n37558 , n37559 , n37560 , n37561 , n37562 , n37563 , n37564 , n37565 , n37566 , n37567 , n37568 , n37569 , n37570 , n37571 , n37572 , n37573 , n37574 , n37575 , n37576 , n37577 , n37578 , n37579 , n37580 , n37581 , n37582 , n37583 , n37584 , n37585 , n37586 , n37587 , n37588 , n37589 , n37590 , n37591 , n37592 , n37593 , n37594 , n37595 , n37596 , n37597 , n37598 , n37599 , n37600 , n37601 , n37602 , n37603 , n37604 , n37605 , n37606 , n37607 , n37608 , n37609 , n37610 , n37611 , n37612 , n37613 , n37614 , n37615 , n37616 , n37617 , n37618 , n37619 , n37620 , n37621 , n37622 , n37623 , n37624 , n37625 , n37626 , n37627 , n37628 , n37629 , n37630 , n37631 , n37632 , n37633 , n37634 , n37635 , n37636 , n37637 , n37638 , n37639 , n37640 , n37641 , n37642 , n37643 , n37644 , n37645 , n37646 , n37647 , n37648 , n37649 , n37650 , n37651 , n37652 , n37653 , n37654 , n37655 , n37656 , n37657 , n37658 , n37659 , n37660 , n37661 , n37662 , n37663 , n37664 , n37665 , n37666 , n37667 , n37668 , n37669 , n37670 , n37671 , n37672 , n37673 , n37674 , n37675 , n37676 , n37677 , n37678 , n37679 , n37680 , n37681 , n37682 , n37683 , n37684 , n37685 , n37686 , n37687 , n37688 , n37689 , n37690 , n37691 , n37692 , n37693 , n37694 , n37695 , n37696 , n37697 , n37698 , n37699 , n37700 , n37701 , n37702 , n37703 , n37704 , n37705 , n37706 , n37707 , n37708 , n37709 , n37710 , n37711 , n37712 , n37713 , n37714 , n37715 , n37716 , n37717 , n37718 , n37719 , n37720 , n37721 , n37722 , n37723 , n37724 , n37725 , n37726 , n37727 , n37728 , n37729 , n37730 , n37731 , n37732 , n37733 , n37734 , n37735 , n37736 , n37737 , n37738 , n37739 , n37740 , n37741 , n37742 , n37743 , n37744 , n37745 , n37746 , n37747 , n37748 , n37749 , n37750 , n37751 , n37752 , n37753 , n37754 , n37755 , n37756 , n37757 , n37758 , n37759 , n37760 , n37761 , n37762 , n37763 , n37764 , n37765 , n37766 , n37767 , n37768 , n37769 , n37770 , n37771 , n37772 , n37773 , n37774 , n37775 , n37776 , n37777 , n37778 , n37779 , n37780 , n37781 , n37782 , n37783 , n37784 , n37785 , n37786 , n37787 , n37788 , n37789 , n37790 , n37791 , n37792 , n37793 , n37794 , n37795 , n37796 , n37797 , n37798 , n37799 , n37800 , n37801 , n37802 , n37803 , n37804 , n37805 , n37806 , n37807 , n37808 , n37809 , n37810 , n37811 , n37812 , n37813 , n37814 , n37815 , n37816 , n37817 , n37818 , n37819 , n37820 , n37821 , n37822 , n37823 , n37824 , n37825 , n37826 , n37827 , n37828 , n37829 , n37830 , n37831 , n37832 , n37833 , n37834 , n37835 , n37836 , n37837 , n37838 , n37839 , n37840 , n37841 , n37842 , n37843 , n37844 , n37845 , n37846 , n37847 , n37848 , n37849 , n37850 , n37851 , n37852 , n37853 , n37854 , n37855 , n37856 , n37857 , n37858 , n37859 , n37860 , n37861 , n37862 , n37863 , n37864 , n37865 , n37866 , n37867 , n37868 , n37869 , n37870 , n37871 , n37872 , n37873 , n37874 , n37875 , n37876 , n37877 , n37878 , n37879 , n37880 , n37881 , n37882 , n37883 , n37884 , n37885 , n37886 , n37887 , n37888 , n37889 , n37890 , n37891 , n37892 , n37893 , n37894 , n37895 , n37896 , n37897 , n37898 , n37899 , n37900 , n37901 , n37902 , n37903 , n37904 , n37905 , n37906 , n37907 , n37908 , n37909 , n37910 , n37911 , n37912 , n37913 , n37914 , n37915 , n37916 , n37917 , n37918 , n37919 , n37920 , n37921 , n37922 , n37923 , n37924 , n37925 , n37926 , n37927 , n37928 , n37929 , n37930 , n37931 , n37932 , n37933 , n37934 , n37935 , n37936 , n37937 , n37938 , n37939 , n37940 , n37941 , n37942 , n37943 , n37944 , n37945 , n37946 , n37947 , n37948 , n37949 , n37950 , n37951 , n37952 , n37953 , n37954 , n37955 , n37956 , n37957 , n37958 , n37959 , n37960 , n37961 , n37962 , n37963 , n37964 , n37965 , n37966 , n37967 , n37968 , n37969 , n37970 , n37971 , n37972 , n37973 , n37974 , n37975 , n37976 , n37977 , n37978 , n37979 , n37980 , n37981 , n37982 , n37983 , n37984 , n37985 , n37986 , n37987 , n37988 , n37989 , n37990 , n37991 , n37992 , n37993 , n37994 , n37995 , n37996 , n37997 , n37998 , n37999 , n38000 , n38001 , n38002 , n38003 , n38004 , n38005 , n38006 , n38007 , n38008 , n38009 , n38010 , n38011 , n38012 , n38013 , n38014 , n38015 , n38016 , n38017 , n38018 , n38019 , n38020 , n38021 , n38022 , n38023 , n38024 , n38025 , n38026 , n38027 , n38028 , n38029 , n38030 , n38031 , n38032 , n38033 , n38034 , n38035 , n38036 , n38037 , n38038 , n38039 , n38040 , n38041 , n38042 , n38043 , n38044 , n38045 , n38046 , n38047 , n38048 , n38049 , n38050 , n38051 , n38052 , n38053 , n38054 , n38055 , n38056 , n38057 , n38058 , n38059 , n38060 , n38061 , n38062 , n38063 , n38064 , n38065 , n38066 , n38067 , n38068 , n38069 , n38070 , n38071 , n38072 , n38073 , n38074 , n38075 , n38076 , n38077 , n38078 , n38079 , n38080 , n38081 , n38082 , n38083 , n38084 , n38085 , n38086 , n38087 , n38088 , n38089 , n38090 , n38091 , n38092 , n38093 , n38094 , n38095 , n38096 , n38097 , n38098 , n38099 , n38100 , n38101 , n38102 , n38103 , n38104 , n38105 , n38106 , n38107 , n38108 , n38109 , n38110 , n38111 , n38112 , n38113 , n38114 , n38115 , n38116 , n38117 , n38118 , n38119 , n38120 , n38121 , n38122 , n38123 , n38124 , n38125 , n38126 , n38127 , n38128 , n38129 , n38130 , n38131 , n38132 , n38133 , n38134 , n38135 , n38136 , n38137 , n38138 , n38139 , n38140 , n38141 , n38142 , n38143 , n38144 , n38145 , n38146 , n38147 , n38148 , n38149 , n38150 , n38151 , n38152 , n38153 , n38154 , n38155 , n38156 , n38157 , n38158 , n38159 , n38160 , n38161 , n38162 , n38163 , n38164 , n38165 , n38166 , n38167 , n38168 , n38169 , n38170 , n38171 , n38172 , n38173 , n38174 , n38175 , n38176 , n38177 , n38178 , n38179 , n38180 , n38181 , n38182 , n38183 , n38184 , n38185 , n38186 , n38187 , n38188 , n38189 , n38190 , n38191 , n38192 , n38193 , n38194 , n38195 , n38196 , n38197 , n38198 , n38199 , n38200 , n38201 , n38202 , n38203 , n38204 , n38205 , n38206 , n38207 , n38208 , n38209 , n38210 , n38211 , n38212 , n38213 , n38214 , n38215 , n38216 , n38217 , n38218 , n38219 , n38220 , n38221 , n38222 , n38223 , n38224 , n38225 , n38226 , n38227 , n38228 , n38229 , n38230 , n38231 , n38232 , n38233 , n38234 , n38235 , n38236 , n38237 , n38238 , n38239 , n38240 , n38241 , n38242 , n38243 , n38244 , n38245 , n38246 , n38247 , n38248 , n38249 , n38250 , n38251 , n38252 , n38253 , n38254 , n38255 , n38256 , n38257 , n38258 , n38259 , n38260 , n38261 , n38262 , n38263 , n38264 , n38265 , n38266 , n38267 , n38268 , n38269 , n38270 , n38271 , n38272 , n38273 , n38274 , n38275 , n38276 , n38277 , n38278 , n38279 , n38280 , n38281 , n38282 , n38283 , n38284 , n38285 , n38286 , n38287 , n38288 , n38289 , n38290 , n38291 , n38292 , n38293 , n38294 , n38295 , n38296 , n38297 , n38298 , n38299 , n38300 , n38301 , n38302 , n38303 , n38304 , n38305 , n38306 , n38307 , n38308 , n38309 , n38310 , n38311 , n38312 , n38313 , n38314 , n38315 , n38316 , n38317 , n38318 , n38319 , n38320 , n38321 , n38322 , n38323 , n38324 , n38325 , n38326 , n38327 , n38328 , n38329 , n38330 , n38331 , n38332 , n38333 , n38334 , n38335 , n38336 , n38337 , n38338 , n38339 , n38340 , n38341 , n38342 , n38343 , n38344 , n38345 , n38346 , n38347 , n38348 , n38349 , n38350 , n38351 , n38352 , n38353 , n38354 , n38355 , n38356 , n38357 , n38358 , n38359 , n38360 , n38361 , n38362 , n38363 , n38364 , n38365 , n38366 , n38367 , n38368 , n38369 , n38370 , n38371 , n38372 , n38373 , n38374 , n38375 , n38376 , n38377 , n38378 , n38379 , n38380 , n38381 , n38382 , n38383 , n38384 , n38385 , n38386 , n38387 , n38388 , n38389 , n38390 , n38391 , n38392 , n38393 , n38394 , n38395 , n38396 , n38397 , n38398 , n38399 , n38400 , n38401 , n38402 , n38403 , n38404 , n38405 , n38406 , n38407 , n38408 , n38409 , n38410 , n38411 , n38412 , n38413 , n38414 , n38415 , n38416 , n38417 , n38418 , n38419 , n38420 , n38421 , n38422 , n38423 , n38424 , n38425 , n38426 , n38427 , n38428 , n38429 , n38430 , n38431 , n38432 , n38433 , n38434 , n38435 , n38436 , n38437 , n38438 , n38439 , n38440 , n38441 , n38442 , n38443 , n38444 , n38445 , n38446 , n38447 , n38448 , n38449 , n38450 , n38451 , n38452 , n38453 , n38454 , n38455 , n38456 , n38457 , n38458 , n38459 , n38460 , n38461 , n38462 , n38463 , n38464 , n38465 , n38466 , n38467 , n38468 , n38469 , n38470 , n38471 , n38472 , n38473 , n38474 , n38475 , n38476 , n38477 , n38478 , n38479 , n38480 , n38481 , n38482 , n38483 , n38484 , n38485 , n38486 , n38487 , n38488 , n38489 , n38490 , n38491 , n38492 , n38493 , n38494 , n38495 , n38496 , n38497 , n38498 , n38499 , n38500 , n38501 , n38502 , n38503 , n38504 , n38505 , n38506 , n38507 , n38508 , n38509 , n38510 , n38511 , n38512 , n38513 , n38514 , n38515 , n38516 , n38517 , n38518 , n38519 , n38520 , n38521 , n38522 , n38523 , n38524 , n38525 , n38526 , n38527 , n38528 , n38529 , n38530 , n38531 , n38532 , n38533 , n38534 , n38535 , n38536 , n38537 , n38538 , n38539 , n38540 , n38541 , n38542 , n38543 , n38544 , n38545 , n38546 , n38547 , n38548 , n38549 , n38550 , n38551 , n38552 , n38553 , n38554 , n38555 , n38556 , n38557 , n38558 , n38559 , n38560 , n38561 , n38562 , n38563 , n38564 , n38565 , n38566 , n38567 , n38568 , n38569 , n38570 , n38571 , n38572 , n38573 , n38574 , n38575 , n38576 , n38577 , n38578 , n38579 , n38580 , n38581 , n38582 , n38583 , n38584 , n38585 , n38586 , n38587 , n38588 ;
  assign n4047 = \clkc_CLKOUT_reg/NET0131  & ~\clkc_ckr_reg_DO_reg[15]/NET0131  ;
  assign n4048 = \bdma_BSreq_reg/NET0131  & ~\core_c_psq_PCS_reg[3]/NET0131  ;
  assign n4049 = ~\core_c_psq_PCS_reg[3]/NET0131  & \sport1_rxctl_RSreq_reg/NET0131  ;
  assign n4050 = ~\core_c_psq_PCS_reg[3]/NET0131  & \sport0_txctl_TSreq_reg/NET0131  ;
  assign n4051 = ~\core_c_psq_PCS_reg[3]/NET0131  & \sport0_rxctl_RSreq_reg/NET0131  ;
  assign n4052 = ~n4050 & ~n4051 ;
  assign n4053 = ~\core_c_psq_PCS_reg[3]/NET0131  & \sport1_txctl_TSreq_reg/NET0131  ;
  assign n4054 = n4052 & ~n4053 ;
  assign n4055 = ~n4049 & n4054 ;
  assign n4056 = ~\idma_DSreq_reg/NET0131  & n4055 ;
  assign n4057 = ~n4048 & n4056 ;
  assign n4058 = ~\idma_IDMA_boot_reg/NET0131_reg_syn_10  & \idma_IDMA_boot_reg/NET0131_reg_syn_2  ;
  assign n4059 = \idma_IDMA_boot_reg/NET0131_reg_syn_10  & \idma_IDMA_boot_reg/NET0131_reg_syn_8  ;
  assign n4060 = ~n4058 & ~n4059 ;
  assign n4061 = ~\bdma_BDMA_boot_reg/NET0131_reg_syn_10  & \bdma_BDMA_boot_reg/NET0131_reg_syn_2  ;
  assign n4062 = \bdma_BDMA_boot_reg/NET0131_reg_syn_10  & \bdma_BDMA_boot_reg/NET0131_reg_syn_8  ;
  assign n4063 = ~n4061 & ~n4062 ;
  assign n4064 = n4060 & n4063 ;
  assign n4065 = \bdma_BM_cyc_reg/P0001  & \core_c_psq_ECYC_reg/P0001  ;
  assign n4066 = ~\memc_EXTC_Eg_reg/NET0131_reg_syn_10  & \memc_EXTC_Eg_reg/NET0131_reg_syn_2  ;
  assign n4067 = \memc_EXTC_Eg_reg/NET0131_reg_syn_10  & \memc_EXTC_Eg_reg/NET0131_reg_syn_8  ;
  assign n4068 = ~n4066 & ~n4067 ;
  assign n4069 = \core_c_psq_PCS_reg[2]/NET0131  & n4068 ;
  assign n4070 = \core_c_psq_PCS_reg[15]/NET0131  & \emc_eRDY_reg/NET0131  ;
  assign n4071 = ~n4069 & ~n4070 ;
  assign n4082 = ~\core_c_psq_TRAP_Eg_reg/NET0131  & ~\sice_HALT_E_reg/P0001  ;
  assign n4083 = ~\auctl_STEAL_reg/NET0131  & ~\core_c_dec_IDLE_Eg_reg/P0001  ;
  assign n4084 = n4082 & n4083 ;
  assign n4085 = ~\core_c_psq_MREQ_reg/NET0131  & n4084 ;
  assign n4080 = \core_c_psq_PCS2or3_reg/NET0131  & ~\memc_LDaST_Eg_reg/NET0131  ;
  assign n4081 = ~\core_c_psq_PCS_reg[12]/NET0131  & ~n4080 ;
  assign n4086 = ~\core_c_dec_MACdep_Eg_reg/P0001  & ~n4081 ;
  assign n4087 = n4085 & n4086 ;
  assign n4078 = ~\core_c_dec_MACdep_Eg_reg/P0001  & ~\core_c_psq_MGNT_reg/NET0131  ;
  assign n4079 = \core_c_psq_PCS_reg[11]/NET0131  & n4078 ;
  assign n4088 = ~\core_c_psq_PCS_reg[5]/NET0131  & ~\core_c_psq_PCS_reg[6]/NET0131  ;
  assign n4089 = ~n4079 & n4088 ;
  assign n4090 = ~n4087 & n4089 ;
  assign n4091 = n4068 & ~n4090 ;
  assign n4072 = ~\clkc_Awake_reg/NET0131  & ~\clkc_STBY_reg/NET0131  ;
  assign n4073 = \clkc_STBY_reg/NET0131  & ~\core_c_psq_TRAP_R_L_reg/NET0131  ;
  assign n4074 = ~\sice_GOICE_syn_reg/P0001  & n4073 ;
  assign n4075 = ~n4072 & ~n4074 ;
  assign n4076 = \core_c_psq_PCS_reg[4]/NET0131  & n4075 ;
  assign n4077 = \core_c_psq_PCS_reg[10]/NET0131  & \emc_eRDY_reg/NET0131  ;
  assign n4092 = ~n4076 & ~n4077 ;
  assign n4093 = ~n4091 & n4092 ;
  assign n4094 = n4071 & n4093 ;
  assign n4095 = ~\auctl_STEAL_reg/NET0131  & ~\clkc_STBY_reg/NET0131  ;
  assign n4096 = n4094 & n4095 ;
  assign n4097 = ~n4065 & n4096 ;
  assign n4098 = n4064 & n4097 ;
  assign n4099 = ~n4057 & ~n4098 ;
  assign n4100 = ~\core_c_dec_IR_reg[21]/NET0131  & ~\core_c_dec_IR_reg[22]/NET0131  ;
  assign n4101 = \core_c_dec_IR_reg[23]/NET0131  & n4100 ;
  assign n4102 = \core_c_psq_PCS_reg[3]/NET0131  & \sice_CMRW_reg/NET0131  ;
  assign n4103 = n4101 & n4102 ;
  assign n4104 = ~\core_c_dec_accCM_E_reg/NET0131  & ~n4103 ;
  assign n4105 = ~\core_c_psq_SRST_reg/P0001  & n4064 ;
  assign n4106 = \core_c_psq_PCS_reg[1]/NET0131  & ~n4105 ;
  assign n4107 = ~\auctl_STEAL_reg/NET0131  & \core_c_psq_PCS2or3_reg/NET0131  ;
  assign n4108 = ~\core_c_psq_PCS_reg[12]/NET0131  & ~n4107 ;
  assign n4109 = \core_c_psq_TRAP_Eg_reg/NET0131  & ~n4108 ;
  assign n4110 = \core_c_dec_EXIT_E_reg/P0001  & \core_c_psq_PCS_reg[2]/NET0131  ;
  assign n4111 = ~n4109 & ~n4110 ;
  assign n4112 = ~n4106 & n4111 ;
  assign n4113 = ~\core_c_psq_PCS_reg[11]/NET0131  & ~n4107 ;
  assign n4114 = ~\core_c_psq_TRAP_Eg_reg/NET0131  & \sice_HALT_E_reg/P0001  ;
  assign n4115 = ~n4113 & n4114 ;
  assign n4116 = n4112 & ~n4115 ;
  assign n4117 = ~\sice_GO_NX_reg/NET0131  & n4094 ;
  assign n4118 = n4116 & n4117 ;
  assign n4119 = n4104 & ~n4118 ;
  assign n4128 = ~n4099 & n4119 ;
  assign n4189 = ~\core_c_psq_pcstk_ptr_reg[1]/NET0131  & ~\core_c_psq_pcstk_ptr_reg[2]/NET0131  ;
  assign n4217 = ~\core_c_psq_pcstk_ptr_reg[0]/NET0131  & n4189 ;
  assign n4220 = \core_c_psq_pcstk_ptr_reg[3]/NET0131  & n4217 ;
  assign n4564 = \core_c_psq_pcstk_cnts16x14_PCcell_reg[8][0]/P0001  & n4220 ;
  assign n4207 = \core_c_psq_pcstk_ptr_reg[1]/NET0131  & \core_c_psq_pcstk_ptr_reg[2]/NET0131  ;
  assign n4208 = \core_c_psq_pcstk_ptr_reg[0]/NET0131  & n4207 ;
  assign n4209 = ~\core_c_psq_pcstk_ptr_reg[3]/NET0131  & n4208 ;
  assign n4567 = \core_c_psq_pcstk_cnts16x14_PCcell_reg[7][0]/P0001  & n4209 ;
  assign n4583 = ~n4564 & ~n4567 ;
  assign n4215 = \core_c_psq_pcstk_ptr_reg[3]/NET0131  & n4208 ;
  assign n4568 = \core_c_psq_pcstk_cnts16x14_PCcell_reg[15][0]/P0001  & n4215 ;
  assign n4218 = ~\core_c_psq_pcstk_ptr_reg[3]/NET0131  & n4217 ;
  assign n4569 = \core_c_psq_pcstk_cnts16x14_PCcell_reg[0][0]/P0001  & n4218 ;
  assign n4584 = ~n4568 & ~n4569 ;
  assign n4585 = n4583 & n4584 ;
  assign n4192 = ~\core_c_psq_pcstk_ptr_reg[1]/NET0131  & \core_c_psq_pcstk_ptr_reg[2]/NET0131  ;
  assign n4204 = \core_c_psq_pcstk_ptr_reg[0]/NET0131  & \core_c_psq_pcstk_ptr_reg[3]/NET0131  ;
  assign n4224 = n4192 & n4204 ;
  assign n4570 = \core_c_psq_pcstk_cnts16x14_PCcell_reg[13][0]/P0001  & n4224 ;
  assign n4193 = ~\core_c_psq_pcstk_ptr_reg[0]/NET0131  & \core_c_psq_pcstk_ptr_reg[3]/NET0131  ;
  assign n4199 = \core_c_psq_pcstk_ptr_reg[1]/NET0131  & ~\core_c_psq_pcstk_ptr_reg[2]/NET0131  ;
  assign n4202 = n4193 & n4199 ;
  assign n4571 = \core_c_psq_pcstk_cnts16x14_PCcell_reg[10][0]/P0001  & n4202 ;
  assign n4578 = ~n4570 & ~n4571 ;
  assign n4205 = n4199 & n4204 ;
  assign n4572 = \core_c_psq_pcstk_cnts16x14_PCcell_reg[11][0]/P0001  & n4205 ;
  assign n4196 = ~\core_c_psq_pcstk_ptr_reg[0]/NET0131  & ~\core_c_psq_pcstk_ptr_reg[3]/NET0131  ;
  assign n4211 = n4196 & n4199 ;
  assign n4573 = \core_c_psq_pcstk_cnts16x14_PCcell_reg[2][0]/P0001  & n4211 ;
  assign n4579 = ~n4572 & ~n4573 ;
  assign n4580 = n4578 & n4579 ;
  assign n4222 = n4193 & n4207 ;
  assign n4562 = \core_c_psq_pcstk_cnts16x14_PCcell_reg[14][0]/P0001  & n4222 ;
  assign n4197 = n4192 & n4196 ;
  assign n4563 = \core_c_psq_pcstk_cnts16x14_PCcell_reg[4][0]/P0001  & n4197 ;
  assign n4576 = ~n4562 & ~n4563 ;
  assign n4188 = \core_c_psq_pcstk_ptr_reg[0]/NET0131  & ~\core_c_psq_pcstk_ptr_reg[3]/NET0131  ;
  assign n4190 = n4188 & n4189 ;
  assign n4565 = \core_c_psq_pcstk_cnts16x14_PCcell_reg[1][0]/P0001  & n4190 ;
  assign n4226 = n4196 & n4207 ;
  assign n4566 = \core_c_psq_pcstk_cnts16x14_PCcell_reg[6][0]/P0001  & n4226 ;
  assign n4577 = ~n4565 & ~n4566 ;
  assign n4581 = n4576 & n4577 ;
  assign n4228 = n4189 & n4204 ;
  assign n4558 = \core_c_psq_pcstk_cnts16x14_PCcell_reg[9][0]/P0001  & n4228 ;
  assign n4213 = n4188 & n4192 ;
  assign n4559 = \core_c_psq_pcstk_cnts16x14_PCcell_reg[5][0]/P0001  & n4213 ;
  assign n4574 = ~n4558 & ~n4559 ;
  assign n4200 = n4188 & n4199 ;
  assign n4560 = \core_c_psq_pcstk_cnts16x14_PCcell_reg[3][0]/P0001  & n4200 ;
  assign n4194 = n4192 & n4193 ;
  assign n4561 = \core_c_psq_pcstk_cnts16x14_PCcell_reg[12][0]/P0001  & n4194 ;
  assign n4575 = ~n4560 & ~n4561 ;
  assign n4582 = n4574 & n4575 ;
  assign n4586 = n4581 & n4582 ;
  assign n4587 = n4580 & n4586 ;
  assign n4588 = n4585 & n4587 ;
  assign n4147 = \clkc_Cnt4096_reg/NET0131  & \clkc_Cnt4096_s2_reg/NET0131  ;
  assign n4148 = \sport0_regs_AUTO_a_reg[12]/NET0131  & n4147 ;
  assign n4149 = ~\bdma_RST_pin_reg/P0001  & ~\sice_RCS_reg[1]/NET0131  ;
  assign n4150 = ~n4148 & n4149 ;
  assign n4151 = ~\core_eu_ec_cun_mven_FFout_reg/NET0131  & n4150 ;
  assign n4152 = \core_eu_ec_cun_MV_reg/P0000_reg_syn_2  & n4151 ;
  assign n4164 = ~\core_eu_em_mac_em_reg_mrovfwe_DO_reg[6]/P0001  & ~\core_eu_em_mac_em_reg_mrovfwe_DO_reg[7]/P0001  ;
  assign n4165 = ~\core_eu_em_mac_em_reg_mrovfwe_DO_reg[8]/P0001  & n4164 ;
  assign n4161 = ~\core_eu_em_mac_em_reg_mrovfwe_DO_reg[0]/P0001  & ~\core_eu_em_mac_em_reg_mrovfwe_DO_reg[1]/P0001  ;
  assign n4162 = ~\core_eu_em_mac_em_reg_mrovfwe_DO_reg[2]/P0001  & ~\core_eu_em_mac_em_reg_mrovfwe_DO_reg[3]/P0001  ;
  assign n4163 = ~\core_eu_em_mac_em_reg_mrovfwe_DO_reg[4]/P0001  & ~\core_eu_em_mac_em_reg_mrovfwe_DO_reg[5]/P0001  ;
  assign n4166 = n4162 & n4163 ;
  assign n4167 = n4161 & n4166 ;
  assign n4168 = n4165 & n4167 ;
  assign n4156 = \core_eu_em_mac_em_reg_mrovfwe_DO_reg[6]/P0001  & \core_eu_em_mac_em_reg_mrovfwe_DO_reg[7]/P0001  ;
  assign n4157 = \core_eu_em_mac_em_reg_mrovfwe_DO_reg[8]/P0001  & n4156 ;
  assign n4153 = \core_eu_em_mac_em_reg_mrovfwe_DO_reg[0]/P0001  & \core_eu_em_mac_em_reg_mrovfwe_DO_reg[1]/P0001  ;
  assign n4154 = \core_eu_em_mac_em_reg_mrovfwe_DO_reg[2]/P0001  & \core_eu_em_mac_em_reg_mrovfwe_DO_reg[3]/P0001  ;
  assign n4155 = \core_eu_em_mac_em_reg_mrovfwe_DO_reg[4]/P0001  & \core_eu_em_mac_em_reg_mrovfwe_DO_reg[5]/P0001  ;
  assign n4158 = n4154 & n4155 ;
  assign n4159 = n4153 & n4158 ;
  assign n4160 = n4157 & n4159 ;
  assign n4169 = \core_eu_ec_cun_updateMV_C_reg/P0001  & ~n4160 ;
  assign n4170 = ~n4168 & n4169 ;
  assign n4171 = ~\core_eu_ec_cun_MVi_pre_C_reg/P0001  & ~n4170 ;
  assign n4172 = n4150 & ~n4171 ;
  assign n4173 = \core_eu_ec_cun_mven_FFout_reg/NET0131  & n4172 ;
  assign n4174 = ~n4152 & ~n4173 ;
  assign n4131 = ~\core_eu_ec_cun_COND_E_reg[0]/P0001  & \core_eu_ec_cun_COND_E_reg[3]/P0001  ;
  assign n4175 = ~\core_eu_ec_cun_COND_E_reg[1]/P0001  & \core_eu_ec_cun_COND_E_reg[2]/P0001  ;
  assign n4179 = n4131 & n4175 ;
  assign n4180 = ~n4174 & n4179 ;
  assign n4176 = \core_eu_ec_cun_COND_E_reg[0]/P0001  & \core_eu_ec_cun_COND_E_reg[3]/P0001  ;
  assign n4177 = n4175 & n4176 ;
  assign n4178 = n4174 & n4177 ;
  assign n4135 = ~\core_eu_ec_cun_AN_reg/P0001  & ~\core_eu_ec_cun_AV_reg/P0001  ;
  assign n4136 = \core_eu_ec_cun_AN_reg/P0001  & \core_eu_ec_cun_AV_reg/P0001  ;
  assign n4137 = ~n4135 & ~n4136 ;
  assign n4138 = ~\core_eu_ec_cun_AZ_reg/P0001  & ~n4137 ;
  assign n4139 = \core_eu_ec_cun_COND_E_reg[1]/P0001  & ~n4138 ;
  assign n4140 = ~\core_eu_ec_cun_AZ_reg/P0001  & ~\core_eu_ec_cun_COND_E_reg[1]/P0001  ;
  assign n4141 = ~n4139 & ~n4140 ;
  assign n4143 = ~\core_eu_ec_cun_COND_E_reg[0]/P0001  & ~n4141 ;
  assign n4142 = \core_eu_ec_cun_COND_E_reg[0]/P0001  & n4141 ;
  assign n4144 = ~\core_eu_ec_cun_COND_E_reg[2]/P0001  & ~\core_eu_ec_cun_COND_E_reg[3]/P0001  ;
  assign n4145 = ~n4142 & n4144 ;
  assign n4146 = ~n4143 & n4145 ;
  assign n4132 = ~\core_c_psq_CE_reg/NET0131  & \core_eu_ec_cun_COND_E_reg[1]/P0001  ;
  assign n4133 = \core_eu_ec_cun_COND_E_reg[2]/P0001  & n4132 ;
  assign n4134 = n4131 & n4133 ;
  assign n4181 = ~\core_eu_ec_cun_condOK_CE_reg/P0001  & ~n4134 ;
  assign n4182 = ~n4146 & n4181 ;
  assign n4183 = ~n4178 & n4182 ;
  assign n4184 = ~n4180 & n4183 ;
  assign n4130 = ~\core_c_dec_IDLE_Eg_reg/P0001  & \core_c_psq_Eqend_Ed_reg/P0001  ;
  assign n4280 = ~\core_eu_ec_cun_TERM_E_reg[0]/P0001  & ~n4174 ;
  assign n4278 = \core_eu_ec_cun_TERM_E_reg[0]/P0001  & n4174 ;
  assign n4279 = \core_eu_ec_cun_TERM_E_reg[2]/P0001  & \core_eu_ec_cun_TERM_E_reg[3]/P0001  ;
  assign n4281 = ~\core_eu_ec_cun_TERM_E_reg[1]/P0001  & n4279 ;
  assign n4282 = ~n4278 & n4281 ;
  assign n4283 = ~n4280 & n4282 ;
  assign n4287 = \core_eu_ec_cun_TERM_E_reg[1]/P0001  & ~n4138 ;
  assign n4288 = ~\core_eu_ec_cun_AZ_reg/P0001  & ~\core_eu_ec_cun_TERM_E_reg[1]/P0001  ;
  assign n4289 = ~n4287 & ~n4288 ;
  assign n4291 = \core_eu_ec_cun_TERM_E_reg[0]/P0001  & ~n4289 ;
  assign n4290 = ~\core_eu_ec_cun_TERM_E_reg[0]/P0001  & n4289 ;
  assign n4292 = ~\core_eu_ec_cun_TERM_E_reg[2]/P0001  & ~\core_eu_ec_cun_TERM_E_reg[3]/P0001  ;
  assign n4293 = ~n4290 & n4292 ;
  assign n4294 = ~n4291 & n4293 ;
  assign n4284 = \core_c_psq_CE_reg/NET0131  & ~\core_eu_ec_cun_TERM_E_reg[0]/P0001  ;
  assign n4285 = \core_eu_ec_cun_TERM_E_reg[1]/P0001  & n4284 ;
  assign n4286 = n4279 & n4285 ;
  assign n4295 = ~\core_eu_ec_cun_termOK_CE_reg/P0001  & ~n4286 ;
  assign n4296 = ~n4294 & n4295 ;
  assign n4297 = ~n4283 & n4296 ;
  assign n4401 = \core_c_psq_pcstk_cnts16x14_PCcell_reg[8][8]/P0001  & n4220 ;
  assign n4404 = \core_c_psq_pcstk_cnts16x14_PCcell_reg[7][8]/P0001  & n4209 ;
  assign n4420 = ~n4401 & ~n4404 ;
  assign n4405 = \core_c_psq_pcstk_cnts16x14_PCcell_reg[15][8]/P0001  & n4215 ;
  assign n4406 = \core_c_psq_pcstk_cnts16x14_PCcell_reg[0][8]/P0001  & n4218 ;
  assign n4421 = ~n4405 & ~n4406 ;
  assign n4422 = n4420 & n4421 ;
  assign n4407 = \core_c_psq_pcstk_cnts16x14_PCcell_reg[13][8]/P0001  & n4224 ;
  assign n4408 = \core_c_psq_pcstk_cnts16x14_PCcell_reg[10][8]/P0001  & n4202 ;
  assign n4415 = ~n4407 & ~n4408 ;
  assign n4409 = \core_c_psq_pcstk_cnts16x14_PCcell_reg[1][8]/P0001  & n4190 ;
  assign n4410 = \core_c_psq_pcstk_cnts16x14_PCcell_reg[3][8]/P0001  & n4200 ;
  assign n4416 = ~n4409 & ~n4410 ;
  assign n4417 = n4415 & n4416 ;
  assign n4399 = \core_c_psq_pcstk_cnts16x14_PCcell_reg[14][8]/P0001  & n4222 ;
  assign n4400 = \core_c_psq_pcstk_cnts16x14_PCcell_reg[4][8]/P0001  & n4197 ;
  assign n4413 = ~n4399 & ~n4400 ;
  assign n4402 = \core_c_psq_pcstk_cnts16x14_PCcell_reg[11][8]/P0001  & n4205 ;
  assign n4403 = \core_c_psq_pcstk_cnts16x14_PCcell_reg[6][8]/P0001  & n4226 ;
  assign n4414 = ~n4402 & ~n4403 ;
  assign n4418 = n4413 & n4414 ;
  assign n4395 = \core_c_psq_pcstk_cnts16x14_PCcell_reg[9][8]/P0001  & n4228 ;
  assign n4396 = \core_c_psq_pcstk_cnts16x14_PCcell_reg[5][8]/P0001  & n4213 ;
  assign n4411 = ~n4395 & ~n4396 ;
  assign n4397 = \core_c_psq_pcstk_cnts16x14_PCcell_reg[2][8]/P0001  & n4211 ;
  assign n4398 = \core_c_psq_pcstk_cnts16x14_PCcell_reg[12][8]/P0001  & n4194 ;
  assign n4412 = ~n4397 & ~n4398 ;
  assign n4419 = n4411 & n4412 ;
  assign n4423 = n4418 & n4419 ;
  assign n4424 = n4417 & n4423 ;
  assign n4425 = n4422 & n4424 ;
  assign n4662 = \core_c_psq_DRA_reg[8]/P0001  & n4425 ;
  assign n4336 = \core_c_psq_pcstk_cnts16x14_PCcell_reg[15][4]/P0001  & n4215 ;
  assign n4339 = \core_c_psq_pcstk_cnts16x14_PCcell_reg[0][4]/P0001  & n4218 ;
  assign n4355 = ~n4336 & ~n4339 ;
  assign n4340 = \core_c_psq_pcstk_cnts16x14_PCcell_reg[7][4]/P0001  & n4209 ;
  assign n4341 = \core_c_psq_pcstk_cnts16x14_PCcell_reg[8][4]/P0001  & n4220 ;
  assign n4356 = ~n4340 & ~n4341 ;
  assign n4357 = n4355 & n4356 ;
  assign n4342 = \core_c_psq_pcstk_cnts16x14_PCcell_reg[2][4]/P0001  & n4211 ;
  assign n4343 = \core_c_psq_pcstk_cnts16x14_PCcell_reg[9][4]/P0001  & n4228 ;
  assign n4350 = ~n4342 & ~n4343 ;
  assign n4344 = \core_c_psq_pcstk_cnts16x14_PCcell_reg[10][4]/P0001  & n4202 ;
  assign n4345 = \core_c_psq_pcstk_cnts16x14_PCcell_reg[13][4]/P0001  & n4224 ;
  assign n4351 = ~n4344 & ~n4345 ;
  assign n4352 = n4350 & n4351 ;
  assign n4334 = \core_c_psq_pcstk_cnts16x14_PCcell_reg[6][4]/P0001  & n4226 ;
  assign n4335 = \core_c_psq_pcstk_cnts16x14_PCcell_reg[5][4]/P0001  & n4213 ;
  assign n4348 = ~n4334 & ~n4335 ;
  assign n4337 = \core_c_psq_pcstk_cnts16x14_PCcell_reg[3][4]/P0001  & n4200 ;
  assign n4338 = \core_c_psq_pcstk_cnts16x14_PCcell_reg[1][4]/P0001  & n4190 ;
  assign n4349 = ~n4337 & ~n4338 ;
  assign n4353 = n4348 & n4349 ;
  assign n4330 = \core_c_psq_pcstk_cnts16x14_PCcell_reg[11][4]/P0001  & n4205 ;
  assign n4331 = \core_c_psq_pcstk_cnts16x14_PCcell_reg[12][4]/P0001  & n4194 ;
  assign n4346 = ~n4330 & ~n4331 ;
  assign n4332 = \core_c_psq_pcstk_cnts16x14_PCcell_reg[4][4]/P0001  & n4197 ;
  assign n4333 = \core_c_psq_pcstk_cnts16x14_PCcell_reg[14][4]/P0001  & n4222 ;
  assign n4347 = ~n4332 & ~n4333 ;
  assign n4354 = n4346 & n4347 ;
  assign n4358 = n4353 & n4354 ;
  assign n4359 = n4352 & n4358 ;
  assign n4360 = n4357 & n4359 ;
  assign n4663 = ~\core_c_psq_DRA_reg[4]/P0001  & ~n4360 ;
  assign n4708 = ~n4662 & ~n4663 ;
  assign n4670 = \core_c_psq_pcstk_cnts16x14_PCcell_reg[8][12]/P0001  & n4220 ;
  assign n4673 = \core_c_psq_pcstk_cnts16x14_PCcell_reg[7][12]/P0001  & n4209 ;
  assign n4689 = ~n4670 & ~n4673 ;
  assign n4674 = \core_c_psq_pcstk_cnts16x14_PCcell_reg[15][12]/P0001  & n4215 ;
  assign n4675 = \core_c_psq_pcstk_cnts16x14_PCcell_reg[0][12]/P0001  & n4218 ;
  assign n4690 = ~n4674 & ~n4675 ;
  assign n4691 = n4689 & n4690 ;
  assign n4676 = \core_c_psq_pcstk_cnts16x14_PCcell_reg[13][12]/P0001  & n4224 ;
  assign n4677 = \core_c_psq_pcstk_cnts16x14_PCcell_reg[10][12]/P0001  & n4202 ;
  assign n4684 = ~n4676 & ~n4677 ;
  assign n4678 = \core_c_psq_pcstk_cnts16x14_PCcell_reg[11][12]/P0001  & n4205 ;
  assign n4679 = \core_c_psq_pcstk_cnts16x14_PCcell_reg[2][12]/P0001  & n4211 ;
  assign n4685 = ~n4678 & ~n4679 ;
  assign n4686 = n4684 & n4685 ;
  assign n4668 = \core_c_psq_pcstk_cnts16x14_PCcell_reg[14][12]/P0001  & n4222 ;
  assign n4669 = \core_c_psq_pcstk_cnts16x14_PCcell_reg[4][12]/P0001  & n4197 ;
  assign n4682 = ~n4668 & ~n4669 ;
  assign n4671 = \core_c_psq_pcstk_cnts16x14_PCcell_reg[1][12]/P0001  & n4190 ;
  assign n4672 = \core_c_psq_pcstk_cnts16x14_PCcell_reg[6][12]/P0001  & n4226 ;
  assign n4683 = ~n4671 & ~n4672 ;
  assign n4687 = n4682 & n4683 ;
  assign n4664 = \core_c_psq_pcstk_cnts16x14_PCcell_reg[9][12]/P0001  & n4228 ;
  assign n4665 = \core_c_psq_pcstk_cnts16x14_PCcell_reg[5][12]/P0001  & n4213 ;
  assign n4680 = ~n4664 & ~n4665 ;
  assign n4666 = \core_c_psq_pcstk_cnts16x14_PCcell_reg[3][12]/P0001  & n4200 ;
  assign n4667 = \core_c_psq_pcstk_cnts16x14_PCcell_reg[12][12]/P0001  & n4194 ;
  assign n4681 = ~n4666 & ~n4667 ;
  assign n4688 = n4680 & n4681 ;
  assign n4692 = n4687 & n4688 ;
  assign n4693 = n4686 & n4692 ;
  assign n4694 = n4691 & n4693 ;
  assign n4695 = ~\core_c_psq_DRA_reg[12]/P0001  & ~n4694 ;
  assign n4696 = \core_c_psq_DRA_reg[12]/P0001  & n4694 ;
  assign n4709 = ~n4695 & ~n4696 ;
  assign n4710 = n4708 & n4709 ;
  assign n4530 = \core_c_psq_pcstk_cnts16x14_PCcell_reg[8][9]/P0001  & n4220 ;
  assign n4533 = \core_c_psq_pcstk_cnts16x14_PCcell_reg[15][9]/P0001  & n4215 ;
  assign n4549 = ~n4530 & ~n4533 ;
  assign n4534 = \core_c_psq_pcstk_cnts16x14_PCcell_reg[0][9]/P0001  & n4218 ;
  assign n4535 = \core_c_psq_pcstk_cnts16x14_PCcell_reg[7][9]/P0001  & n4209 ;
  assign n4550 = ~n4534 & ~n4535 ;
  assign n4551 = n4549 & n4550 ;
  assign n4536 = \core_c_psq_pcstk_cnts16x14_PCcell_reg[1][9]/P0001  & n4190 ;
  assign n4537 = \core_c_psq_pcstk_cnts16x14_PCcell_reg[14][9]/P0001  & n4222 ;
  assign n4544 = ~n4536 & ~n4537 ;
  assign n4538 = \core_c_psq_pcstk_cnts16x14_PCcell_reg[5][9]/P0001  & n4213 ;
  assign n4539 = \core_c_psq_pcstk_cnts16x14_PCcell_reg[3][9]/P0001  & n4200 ;
  assign n4545 = ~n4538 & ~n4539 ;
  assign n4546 = n4544 & n4545 ;
  assign n4528 = \core_c_psq_pcstk_cnts16x14_PCcell_reg[11][9]/P0001  & n4205 ;
  assign n4529 = \core_c_psq_pcstk_cnts16x14_PCcell_reg[6][9]/P0001  & n4226 ;
  assign n4542 = ~n4528 & ~n4529 ;
  assign n4531 = \core_c_psq_pcstk_cnts16x14_PCcell_reg[9][9]/P0001  & n4228 ;
  assign n4532 = \core_c_psq_pcstk_cnts16x14_PCcell_reg[4][9]/P0001  & n4197 ;
  assign n4543 = ~n4531 & ~n4532 ;
  assign n4547 = n4542 & n4543 ;
  assign n4524 = \core_c_psq_pcstk_cnts16x14_PCcell_reg[10][9]/P0001  & n4202 ;
  assign n4525 = \core_c_psq_pcstk_cnts16x14_PCcell_reg[2][9]/P0001  & n4211 ;
  assign n4540 = ~n4524 & ~n4525 ;
  assign n4526 = \core_c_psq_pcstk_cnts16x14_PCcell_reg[12][9]/P0001  & n4194 ;
  assign n4527 = \core_c_psq_pcstk_cnts16x14_PCcell_reg[13][9]/P0001  & n4224 ;
  assign n4541 = ~n4526 & ~n4527 ;
  assign n4548 = n4540 & n4541 ;
  assign n4552 = n4547 & n4548 ;
  assign n4553 = n4546 & n4552 ;
  assign n4554 = n4551 & n4553 ;
  assign n4658 = ~\core_c_psq_DRA_reg[9]/P0001  & ~n4554 ;
  assign n4465 = \core_c_psq_pcstk_cnts16x14_PCcell_reg[7][13]/P0001  & n4209 ;
  assign n4468 = \core_c_psq_pcstk_cnts16x14_PCcell_reg[15][13]/P0001  & n4215 ;
  assign n4484 = ~n4465 & ~n4468 ;
  assign n4469 = \core_c_psq_pcstk_cnts16x14_PCcell_reg[0][13]/P0001  & n4218 ;
  assign n4470 = \core_c_psq_pcstk_cnts16x14_PCcell_reg[8][13]/P0001  & n4220 ;
  assign n4485 = ~n4469 & ~n4470 ;
  assign n4486 = n4484 & n4485 ;
  assign n4471 = \core_c_psq_pcstk_cnts16x14_PCcell_reg[14][13]/P0001  & n4222 ;
  assign n4472 = \core_c_psq_pcstk_cnts16x14_PCcell_reg[13][13]/P0001  & n4224 ;
  assign n4479 = ~n4471 & ~n4472 ;
  assign n4473 = \core_c_psq_pcstk_cnts16x14_PCcell_reg[6][13]/P0001  & n4226 ;
  assign n4474 = \core_c_psq_pcstk_cnts16x14_PCcell_reg[9][13]/P0001  & n4228 ;
  assign n4480 = ~n4473 & ~n4474 ;
  assign n4481 = n4479 & n4480 ;
  assign n4463 = \core_c_psq_pcstk_cnts16x14_PCcell_reg[10][13]/P0001  & n4202 ;
  assign n4464 = \core_c_psq_pcstk_cnts16x14_PCcell_reg[11][13]/P0001  & n4205 ;
  assign n4477 = ~n4463 & ~n4464 ;
  assign n4466 = \core_c_psq_pcstk_cnts16x14_PCcell_reg[2][13]/P0001  & n4211 ;
  assign n4467 = \core_c_psq_pcstk_cnts16x14_PCcell_reg[5][13]/P0001  & n4213 ;
  assign n4478 = ~n4466 & ~n4467 ;
  assign n4482 = n4477 & n4478 ;
  assign n4459 = \core_c_psq_pcstk_cnts16x14_PCcell_reg[1][13]/P0001  & n4190 ;
  assign n4460 = \core_c_psq_pcstk_cnts16x14_PCcell_reg[12][13]/P0001  & n4194 ;
  assign n4475 = ~n4459 & ~n4460 ;
  assign n4461 = \core_c_psq_pcstk_cnts16x14_PCcell_reg[4][13]/P0001  & n4197 ;
  assign n4462 = \core_c_psq_pcstk_cnts16x14_PCcell_reg[3][13]/P0001  & n4200 ;
  assign n4476 = ~n4461 & ~n4462 ;
  assign n4483 = n4475 & n4476 ;
  assign n4487 = n4482 & n4483 ;
  assign n4488 = n4481 & n4487 ;
  assign n4489 = n4486 & n4488 ;
  assign n4659 = \core_c_psq_DRA_reg[13]/P0001  & n4489 ;
  assign n4706 = ~n4658 & ~n4659 ;
  assign n4252 = \core_c_psq_pcstk_cnts16x14_PCcell_reg[8][10]/P0001  & n4220 ;
  assign n4255 = \core_c_psq_pcstk_cnts16x14_PCcell_reg[7][10]/P0001  & n4209 ;
  assign n4271 = ~n4252 & ~n4255 ;
  assign n4256 = \core_c_psq_pcstk_cnts16x14_PCcell_reg[15][10]/P0001  & n4215 ;
  assign n4257 = \core_c_psq_pcstk_cnts16x14_PCcell_reg[0][10]/P0001  & n4218 ;
  assign n4272 = ~n4256 & ~n4257 ;
  assign n4273 = n4271 & n4272 ;
  assign n4258 = \core_c_psq_pcstk_cnts16x14_PCcell_reg[1][10]/P0001  & n4190 ;
  assign n4259 = \core_c_psq_pcstk_cnts16x14_PCcell_reg[14][10]/P0001  & n4222 ;
  assign n4266 = ~n4258 & ~n4259 ;
  assign n4260 = \core_c_psq_pcstk_cnts16x14_PCcell_reg[5][10]/P0001  & n4213 ;
  assign n4261 = \core_c_psq_pcstk_cnts16x14_PCcell_reg[3][10]/P0001  & n4200 ;
  assign n4267 = ~n4260 & ~n4261 ;
  assign n4268 = n4266 & n4267 ;
  assign n4250 = \core_c_psq_pcstk_cnts16x14_PCcell_reg[11][10]/P0001  & n4205 ;
  assign n4251 = \core_c_psq_pcstk_cnts16x14_PCcell_reg[6][10]/P0001  & n4226 ;
  assign n4264 = ~n4250 & ~n4251 ;
  assign n4253 = \core_c_psq_pcstk_cnts16x14_PCcell_reg[9][10]/P0001  & n4228 ;
  assign n4254 = \core_c_psq_pcstk_cnts16x14_PCcell_reg[4][10]/P0001  & n4197 ;
  assign n4265 = ~n4253 & ~n4254 ;
  assign n4269 = n4264 & n4265 ;
  assign n4246 = \core_c_psq_pcstk_cnts16x14_PCcell_reg[10][10]/P0001  & n4202 ;
  assign n4247 = \core_c_psq_pcstk_cnts16x14_PCcell_reg[2][10]/P0001  & n4211 ;
  assign n4262 = ~n4246 & ~n4247 ;
  assign n4248 = \core_c_psq_pcstk_cnts16x14_PCcell_reg[12][10]/P0001  & n4194 ;
  assign n4249 = \core_c_psq_pcstk_cnts16x14_PCcell_reg[13][10]/P0001  & n4224 ;
  assign n4263 = ~n4248 & ~n4249 ;
  assign n4270 = n4262 & n4263 ;
  assign n4274 = n4269 & n4270 ;
  assign n4275 = n4268 & n4274 ;
  assign n4276 = n4273 & n4275 ;
  assign n4660 = ~\core_c_psq_DRA_reg[10]/P0001  & ~n4276 ;
  assign n4632 = \core_c_psq_pcstk_cnts16x14_PCcell_reg[8][7]/P0001  & n4220 ;
  assign n4635 = \core_c_psq_pcstk_cnts16x14_PCcell_reg[7][7]/P0001  & n4209 ;
  assign n4651 = ~n4632 & ~n4635 ;
  assign n4636 = \core_c_psq_pcstk_cnts16x14_PCcell_reg[15][7]/P0001  & n4215 ;
  assign n4637 = \core_c_psq_pcstk_cnts16x14_PCcell_reg[0][7]/P0001  & n4218 ;
  assign n4652 = ~n4636 & ~n4637 ;
  assign n4653 = n4651 & n4652 ;
  assign n4638 = \core_c_psq_pcstk_cnts16x14_PCcell_reg[13][7]/P0001  & n4224 ;
  assign n4639 = \core_c_psq_pcstk_cnts16x14_PCcell_reg[10][7]/P0001  & n4202 ;
  assign n4646 = ~n4638 & ~n4639 ;
  assign n4640 = \core_c_psq_pcstk_cnts16x14_PCcell_reg[1][7]/P0001  & n4190 ;
  assign n4641 = \core_c_psq_pcstk_cnts16x14_PCcell_reg[14][7]/P0001  & n4222 ;
  assign n4647 = ~n4640 & ~n4641 ;
  assign n4648 = n4646 & n4647 ;
  assign n4630 = \core_c_psq_pcstk_cnts16x14_PCcell_reg[3][7]/P0001  & n4200 ;
  assign n4631 = \core_c_psq_pcstk_cnts16x14_PCcell_reg[4][7]/P0001  & n4197 ;
  assign n4644 = ~n4630 & ~n4631 ;
  assign n4633 = \core_c_psq_pcstk_cnts16x14_PCcell_reg[5][7]/P0001  & n4213 ;
  assign n4634 = \core_c_psq_pcstk_cnts16x14_PCcell_reg[6][7]/P0001  & n4226 ;
  assign n4645 = ~n4633 & ~n4634 ;
  assign n4649 = n4644 & n4645 ;
  assign n4626 = \core_c_psq_pcstk_cnts16x14_PCcell_reg[9][7]/P0001  & n4228 ;
  assign n4627 = \core_c_psq_pcstk_cnts16x14_PCcell_reg[11][7]/P0001  & n4205 ;
  assign n4642 = ~n4626 & ~n4627 ;
  assign n4628 = \core_c_psq_pcstk_cnts16x14_PCcell_reg[2][7]/P0001  & n4211 ;
  assign n4629 = \core_c_psq_pcstk_cnts16x14_PCcell_reg[12][7]/P0001  & n4194 ;
  assign n4643 = ~n4628 & ~n4629 ;
  assign n4650 = n4642 & n4643 ;
  assign n4654 = n4649 & n4650 ;
  assign n4655 = n4648 & n4654 ;
  assign n4656 = n4653 & n4655 ;
  assign n4661 = ~\core_c_psq_DRA_reg[7]/P0001  & ~n4656 ;
  assign n4707 = ~n4660 & ~n4661 ;
  assign n4711 = n4706 & n4707 ;
  assign n4589 = ~\core_c_psq_DRA_reg[0]/P0001  & ~n4588 ;
  assign n4304 = \core_c_psq_pcstk_cnts16x14_PCcell_reg[7][3]/P0001  & n4209 ;
  assign n4307 = \core_c_psq_pcstk_cnts16x14_PCcell_reg[15][3]/P0001  & n4215 ;
  assign n4323 = ~n4304 & ~n4307 ;
  assign n4308 = \core_c_psq_pcstk_cnts16x14_PCcell_reg[0][3]/P0001  & n4218 ;
  assign n4309 = \core_c_psq_pcstk_cnts16x14_PCcell_reg[8][3]/P0001  & n4220 ;
  assign n4324 = ~n4308 & ~n4309 ;
  assign n4325 = n4323 & n4324 ;
  assign n4310 = \core_c_psq_pcstk_cnts16x14_PCcell_reg[14][3]/P0001  & n4222 ;
  assign n4311 = \core_c_psq_pcstk_cnts16x14_PCcell_reg[13][3]/P0001  & n4224 ;
  assign n4318 = ~n4310 & ~n4311 ;
  assign n4312 = \core_c_psq_pcstk_cnts16x14_PCcell_reg[6][3]/P0001  & n4226 ;
  assign n4313 = \core_c_psq_pcstk_cnts16x14_PCcell_reg[9][3]/P0001  & n4228 ;
  assign n4319 = ~n4312 & ~n4313 ;
  assign n4320 = n4318 & n4319 ;
  assign n4302 = \core_c_psq_pcstk_cnts16x14_PCcell_reg[10][3]/P0001  & n4202 ;
  assign n4303 = \core_c_psq_pcstk_cnts16x14_PCcell_reg[11][3]/P0001  & n4205 ;
  assign n4316 = ~n4302 & ~n4303 ;
  assign n4305 = \core_c_psq_pcstk_cnts16x14_PCcell_reg[2][3]/P0001  & n4211 ;
  assign n4306 = \core_c_psq_pcstk_cnts16x14_PCcell_reg[5][3]/P0001  & n4213 ;
  assign n4317 = ~n4305 & ~n4306 ;
  assign n4321 = n4316 & n4317 ;
  assign n4298 = \core_c_psq_pcstk_cnts16x14_PCcell_reg[1][3]/P0001  & n4190 ;
  assign n4299 = \core_c_psq_pcstk_cnts16x14_PCcell_reg[12][3]/P0001  & n4194 ;
  assign n4314 = ~n4298 & ~n4299 ;
  assign n4300 = \core_c_psq_pcstk_cnts16x14_PCcell_reg[4][3]/P0001  & n4197 ;
  assign n4301 = \core_c_psq_pcstk_cnts16x14_PCcell_reg[3][3]/P0001  & n4200 ;
  assign n4315 = ~n4300 & ~n4301 ;
  assign n4322 = n4314 & n4315 ;
  assign n4326 = n4321 & n4322 ;
  assign n4327 = n4320 & n4326 ;
  assign n4328 = n4325 & n4327 ;
  assign n4590 = ~\core_c_psq_DRA_reg[3]/P0001  & ~n4328 ;
  assign n4704 = ~n4589 & ~n4590 ;
  assign n4591 = \core_c_psq_DRA_reg[0]/P0001  & n4588 ;
  assign n4657 = \core_c_psq_DRA_reg[7]/P0001  & n4656 ;
  assign n4705 = ~n4591 & ~n4657 ;
  assign n4712 = n4704 & n4705 ;
  assign n4719 = n4711 & n4712 ;
  assign n4720 = n4710 & n4719 ;
  assign n4329 = \core_c_psq_DRA_reg[3]/P0001  & n4328 ;
  assign n4361 = \core_c_psq_DRA_reg[4]/P0001  & n4360 ;
  assign n4698 = ~n4329 & ~n4361 ;
  assign n4368 = \core_c_psq_pcstk_cnts16x14_PCcell_reg[7][6]/P0001  & n4209 ;
  assign n4371 = \core_c_psq_pcstk_cnts16x14_PCcell_reg[15][6]/P0001  & n4215 ;
  assign n4387 = ~n4368 & ~n4371 ;
  assign n4372 = \core_c_psq_pcstk_cnts16x14_PCcell_reg[0][6]/P0001  & n4218 ;
  assign n4373 = \core_c_psq_pcstk_cnts16x14_PCcell_reg[8][6]/P0001  & n4220 ;
  assign n4388 = ~n4372 & ~n4373 ;
  assign n4389 = n4387 & n4388 ;
  assign n4374 = \core_c_psq_pcstk_cnts16x14_PCcell_reg[13][6]/P0001  & n4224 ;
  assign n4375 = \core_c_psq_pcstk_cnts16x14_PCcell_reg[1][6]/P0001  & n4190 ;
  assign n4382 = ~n4374 & ~n4375 ;
  assign n4376 = \core_c_psq_pcstk_cnts16x14_PCcell_reg[10][6]/P0001  & n4202 ;
  assign n4377 = \core_c_psq_pcstk_cnts16x14_PCcell_reg[11][6]/P0001  & n4205 ;
  assign n4383 = ~n4376 & ~n4377 ;
  assign n4384 = n4382 & n4383 ;
  assign n4366 = \core_c_psq_pcstk_cnts16x14_PCcell_reg[9][6]/P0001  & n4228 ;
  assign n4367 = \core_c_psq_pcstk_cnts16x14_PCcell_reg[4][6]/P0001  & n4197 ;
  assign n4380 = ~n4366 & ~n4367 ;
  assign n4369 = \core_c_psq_pcstk_cnts16x14_PCcell_reg[12][6]/P0001  & n4194 ;
  assign n4370 = \core_c_psq_pcstk_cnts16x14_PCcell_reg[3][6]/P0001  & n4200 ;
  assign n4381 = ~n4369 & ~n4370 ;
  assign n4385 = n4380 & n4381 ;
  assign n4362 = \core_c_psq_pcstk_cnts16x14_PCcell_reg[6][6]/P0001  & n4226 ;
  assign n4363 = \core_c_psq_pcstk_cnts16x14_PCcell_reg[14][6]/P0001  & n4222 ;
  assign n4378 = ~n4362 & ~n4363 ;
  assign n4364 = \core_c_psq_pcstk_cnts16x14_PCcell_reg[2][6]/P0001  & n4211 ;
  assign n4365 = \core_c_psq_pcstk_cnts16x14_PCcell_reg[5][6]/P0001  & n4213 ;
  assign n4379 = ~n4364 & ~n4365 ;
  assign n4386 = n4378 & n4379 ;
  assign n4390 = n4385 & n4386 ;
  assign n4391 = n4384 & n4390 ;
  assign n4392 = n4389 & n4391 ;
  assign n4393 = ~\core_c_psq_DRA_reg[6]/P0001  & ~n4392 ;
  assign n4394 = \core_c_psq_DRA_reg[6]/P0001  & n4392 ;
  assign n4699 = ~n4393 & ~n4394 ;
  assign n4715 = n4698 & n4699 ;
  assign n4598 = \core_c_psq_pcstk_cnts16x14_PCcell_reg[8][11]/P0001  & n4220 ;
  assign n4601 = \core_c_psq_pcstk_cnts16x14_PCcell_reg[15][11]/P0001  & n4215 ;
  assign n4617 = ~n4598 & ~n4601 ;
  assign n4602 = \core_c_psq_pcstk_cnts16x14_PCcell_reg[0][11]/P0001  & n4218 ;
  assign n4603 = \core_c_psq_pcstk_cnts16x14_PCcell_reg[7][11]/P0001  & n4209 ;
  assign n4618 = ~n4602 & ~n4603 ;
  assign n4619 = n4617 & n4618 ;
  assign n4604 = \core_c_psq_pcstk_cnts16x14_PCcell_reg[5][11]/P0001  & n4213 ;
  assign n4605 = \core_c_psq_pcstk_cnts16x14_PCcell_reg[10][11]/P0001  & n4202 ;
  assign n4612 = ~n4604 & ~n4605 ;
  assign n4606 = \core_c_psq_pcstk_cnts16x14_PCcell_reg[11][11]/P0001  & n4205 ;
  assign n4607 = \core_c_psq_pcstk_cnts16x14_PCcell_reg[6][11]/P0001  & n4226 ;
  assign n4613 = ~n4606 & ~n4607 ;
  assign n4614 = n4612 & n4613 ;
  assign n4596 = \core_c_psq_pcstk_cnts16x14_PCcell_reg[3][11]/P0001  & n4200 ;
  assign n4597 = \core_c_psq_pcstk_cnts16x14_PCcell_reg[12][11]/P0001  & n4194 ;
  assign n4610 = ~n4596 & ~n4597 ;
  assign n4599 = \core_c_psq_pcstk_cnts16x14_PCcell_reg[2][11]/P0001  & n4211 ;
  assign n4600 = \core_c_psq_pcstk_cnts16x14_PCcell_reg[13][11]/P0001  & n4224 ;
  assign n4611 = ~n4599 & ~n4600 ;
  assign n4615 = n4610 & n4611 ;
  assign n4592 = \core_c_psq_pcstk_cnts16x14_PCcell_reg[14][11]/P0001  & n4222 ;
  assign n4593 = \core_c_psq_pcstk_cnts16x14_PCcell_reg[1][11]/P0001  & n4190 ;
  assign n4608 = ~n4592 & ~n4593 ;
  assign n4594 = \core_c_psq_pcstk_cnts16x14_PCcell_reg[9][11]/P0001  & n4228 ;
  assign n4595 = \core_c_psq_pcstk_cnts16x14_PCcell_reg[4][11]/P0001  & n4197 ;
  assign n4609 = ~n4594 & ~n4595 ;
  assign n4616 = n4608 & n4609 ;
  assign n4620 = n4615 & n4616 ;
  assign n4621 = n4614 & n4620 ;
  assign n4622 = n4619 & n4621 ;
  assign n4623 = \core_c_psq_DRA_reg[11]/P0001  & ~n4622 ;
  assign n4624 = ~\core_c_psq_DRA_reg[11]/P0001  & n4622 ;
  assign n4625 = ~n4623 & ~n4624 ;
  assign n4210 = \core_c_psq_pcstk_cnts16x14_PCcell_reg[7][5]/P0001  & n4209 ;
  assign n4216 = \core_c_psq_pcstk_cnts16x14_PCcell_reg[15][5]/P0001  & n4215 ;
  assign n4239 = ~n4210 & ~n4216 ;
  assign n4219 = \core_c_psq_pcstk_cnts16x14_PCcell_reg[0][5]/P0001  & n4218 ;
  assign n4221 = \core_c_psq_pcstk_cnts16x14_PCcell_reg[8][5]/P0001  & n4220 ;
  assign n4240 = ~n4219 & ~n4221 ;
  assign n4241 = n4239 & n4240 ;
  assign n4223 = \core_c_psq_pcstk_cnts16x14_PCcell_reg[14][5]/P0001  & n4222 ;
  assign n4225 = \core_c_psq_pcstk_cnts16x14_PCcell_reg[13][5]/P0001  & n4224 ;
  assign n4234 = ~n4223 & ~n4225 ;
  assign n4227 = \core_c_psq_pcstk_cnts16x14_PCcell_reg[6][5]/P0001  & n4226 ;
  assign n4229 = \core_c_psq_pcstk_cnts16x14_PCcell_reg[9][5]/P0001  & n4228 ;
  assign n4235 = ~n4227 & ~n4229 ;
  assign n4236 = n4234 & n4235 ;
  assign n4203 = \core_c_psq_pcstk_cnts16x14_PCcell_reg[10][5]/P0001  & n4202 ;
  assign n4206 = \core_c_psq_pcstk_cnts16x14_PCcell_reg[11][5]/P0001  & n4205 ;
  assign n4232 = ~n4203 & ~n4206 ;
  assign n4212 = \core_c_psq_pcstk_cnts16x14_PCcell_reg[2][5]/P0001  & n4211 ;
  assign n4214 = \core_c_psq_pcstk_cnts16x14_PCcell_reg[5][5]/P0001  & n4213 ;
  assign n4233 = ~n4212 & ~n4214 ;
  assign n4237 = n4232 & n4233 ;
  assign n4191 = \core_c_psq_pcstk_cnts16x14_PCcell_reg[1][5]/P0001  & n4190 ;
  assign n4195 = \core_c_psq_pcstk_cnts16x14_PCcell_reg[12][5]/P0001  & n4194 ;
  assign n4230 = ~n4191 & ~n4195 ;
  assign n4198 = \core_c_psq_pcstk_cnts16x14_PCcell_reg[4][5]/P0001  & n4197 ;
  assign n4201 = \core_c_psq_pcstk_cnts16x14_PCcell_reg[3][5]/P0001  & n4200 ;
  assign n4231 = ~n4198 & ~n4201 ;
  assign n4238 = n4230 & n4231 ;
  assign n4242 = n4237 & n4238 ;
  assign n4243 = n4236 & n4242 ;
  assign n4244 = n4241 & n4243 ;
  assign n4245 = \core_c_psq_DRA_reg[5]/P0001  & n4244 ;
  assign n4277 = \core_c_psq_DRA_reg[10]/P0001  & n4276 ;
  assign n4697 = ~n4245 & ~n4277 ;
  assign n4716 = ~n4625 & n4697 ;
  assign n4717 = n4715 & n4716 ;
  assign n4523 = ~\core_c_psq_DRA_reg[5]/P0001  & ~n4244 ;
  assign n4555 = \core_c_psq_DRA_reg[9]/P0001  & n4554 ;
  assign n4702 = ~n4523 & ~n4555 ;
  assign n4497 = \core_c_psq_pcstk_cnts16x14_PCcell_reg[8][2]/P0001  & n4220 ;
  assign n4500 = \core_c_psq_pcstk_cnts16x14_PCcell_reg[7][2]/P0001  & n4209 ;
  assign n4516 = ~n4497 & ~n4500 ;
  assign n4501 = \core_c_psq_pcstk_cnts16x14_PCcell_reg[15][2]/P0001  & n4215 ;
  assign n4502 = \core_c_psq_pcstk_cnts16x14_PCcell_reg[0][2]/P0001  & n4218 ;
  assign n4517 = ~n4501 & ~n4502 ;
  assign n4518 = n4516 & n4517 ;
  assign n4503 = \core_c_psq_pcstk_cnts16x14_PCcell_reg[14][2]/P0001  & n4222 ;
  assign n4504 = \core_c_psq_pcstk_cnts16x14_PCcell_reg[10][2]/P0001  & n4202 ;
  assign n4511 = ~n4503 & ~n4504 ;
  assign n4505 = \core_c_psq_pcstk_cnts16x14_PCcell_reg[11][2]/P0001  & n4205 ;
  assign n4506 = \core_c_psq_pcstk_cnts16x14_PCcell_reg[6][2]/P0001  & n4226 ;
  assign n4512 = ~n4505 & ~n4506 ;
  assign n4513 = n4511 & n4512 ;
  assign n4495 = \core_c_psq_pcstk_cnts16x14_PCcell_reg[3][2]/P0001  & n4200 ;
  assign n4496 = \core_c_psq_pcstk_cnts16x14_PCcell_reg[12][2]/P0001  & n4194 ;
  assign n4509 = ~n4495 & ~n4496 ;
  assign n4498 = \core_c_psq_pcstk_cnts16x14_PCcell_reg[2][2]/P0001  & n4211 ;
  assign n4499 = \core_c_psq_pcstk_cnts16x14_PCcell_reg[13][2]/P0001  & n4224 ;
  assign n4510 = ~n4498 & ~n4499 ;
  assign n4514 = n4509 & n4510 ;
  assign n4491 = \core_c_psq_pcstk_cnts16x14_PCcell_reg[5][2]/P0001  & n4213 ;
  assign n4492 = \core_c_psq_pcstk_cnts16x14_PCcell_reg[1][2]/P0001  & n4190 ;
  assign n4507 = ~n4491 & ~n4492 ;
  assign n4493 = \core_c_psq_pcstk_cnts16x14_PCcell_reg[9][2]/P0001  & n4228 ;
  assign n4494 = \core_c_psq_pcstk_cnts16x14_PCcell_reg[4][2]/P0001  & n4197 ;
  assign n4508 = ~n4493 & ~n4494 ;
  assign n4515 = n4507 & n4508 ;
  assign n4519 = n4514 & n4515 ;
  assign n4520 = n4513 & n4519 ;
  assign n4521 = n4518 & n4520 ;
  assign n4556 = \core_c_psq_DRA_reg[2]/P0001  & n4521 ;
  assign n4433 = \core_c_psq_pcstk_cnts16x14_PCcell_reg[8][1]/P0001  & n4220 ;
  assign n4436 = \core_c_psq_pcstk_cnts16x14_PCcell_reg[7][1]/P0001  & n4209 ;
  assign n4452 = ~n4433 & ~n4436 ;
  assign n4437 = \core_c_psq_pcstk_cnts16x14_PCcell_reg[15][1]/P0001  & n4215 ;
  assign n4438 = \core_c_psq_pcstk_cnts16x14_PCcell_reg[0][1]/P0001  & n4218 ;
  assign n4453 = ~n4437 & ~n4438 ;
  assign n4454 = n4452 & n4453 ;
  assign n4439 = \core_c_psq_pcstk_cnts16x14_PCcell_reg[1][1]/P0001  & n4190 ;
  assign n4440 = \core_c_psq_pcstk_cnts16x14_PCcell_reg[14][1]/P0001  & n4222 ;
  assign n4447 = ~n4439 & ~n4440 ;
  assign n4441 = \core_c_psq_pcstk_cnts16x14_PCcell_reg[5][1]/P0001  & n4213 ;
  assign n4442 = \core_c_psq_pcstk_cnts16x14_PCcell_reg[3][1]/P0001  & n4200 ;
  assign n4448 = ~n4441 & ~n4442 ;
  assign n4449 = n4447 & n4448 ;
  assign n4431 = \core_c_psq_pcstk_cnts16x14_PCcell_reg[11][1]/P0001  & n4205 ;
  assign n4432 = \core_c_psq_pcstk_cnts16x14_PCcell_reg[6][1]/P0001  & n4226 ;
  assign n4445 = ~n4431 & ~n4432 ;
  assign n4434 = \core_c_psq_pcstk_cnts16x14_PCcell_reg[9][1]/P0001  & n4228 ;
  assign n4435 = \core_c_psq_pcstk_cnts16x14_PCcell_reg[4][1]/P0001  & n4197 ;
  assign n4446 = ~n4434 & ~n4435 ;
  assign n4450 = n4445 & n4446 ;
  assign n4427 = \core_c_psq_pcstk_cnts16x14_PCcell_reg[10][1]/P0001  & n4202 ;
  assign n4428 = \core_c_psq_pcstk_cnts16x14_PCcell_reg[2][1]/P0001  & n4211 ;
  assign n4443 = ~n4427 & ~n4428 ;
  assign n4429 = \core_c_psq_pcstk_cnts16x14_PCcell_reg[12][1]/P0001  & n4194 ;
  assign n4430 = \core_c_psq_pcstk_cnts16x14_PCcell_reg[13][1]/P0001  & n4224 ;
  assign n4444 = ~n4429 & ~n4430 ;
  assign n4451 = n4443 & n4444 ;
  assign n4455 = n4450 & n4451 ;
  assign n4456 = n4449 & n4455 ;
  assign n4457 = n4454 & n4456 ;
  assign n4557 = \core_c_psq_DRA_reg[1]/P0001  & n4457 ;
  assign n4703 = ~n4556 & ~n4557 ;
  assign n4713 = n4702 & n4703 ;
  assign n4426 = ~\core_c_psq_DRA_reg[8]/P0001  & ~n4425 ;
  assign n4458 = ~\core_c_psq_DRA_reg[1]/P0001  & ~n4457 ;
  assign n4700 = ~n4426 & ~n4458 ;
  assign n4490 = ~\core_c_psq_DRA_reg[13]/P0001  & ~n4489 ;
  assign n4522 = ~\core_c_psq_DRA_reg[2]/P0001  & ~n4521 ;
  assign n4701 = ~n4490 & ~n4522 ;
  assign n4714 = n4700 & n4701 ;
  assign n4718 = n4713 & n4714 ;
  assign n4721 = n4717 & n4718 ;
  assign n4722 = n4720 & n4721 ;
  assign n4723 = n4297 & n4722 ;
  assign n4724 = n4130 & ~n4723 ;
  assign n4725 = n4184 & ~n4724 ;
  assign n4786 = \core_c_dec_BR_Ed_reg/P0001  & \core_c_psq_Taddr_Eb_reg[13]/P0001  ;
  assign n4787 = ~\core_c_dec_BR_Ed_reg/P0001  & ~n4489 ;
  assign n4788 = ~n4786 & ~n4787 ;
  assign n4796 = ~\core_c_psq_DRA_reg[13]/P0001  & ~n4788 ;
  assign n4755 = \core_c_dec_BR_Ed_reg/P0001  & \core_c_psq_Taddr_Eb_reg[10]/P0001  ;
  assign n4756 = ~\core_c_dec_BR_Ed_reg/P0001  & ~n4276 ;
  assign n4757 = ~n4755 & ~n4756 ;
  assign n4797 = \core_c_psq_DRA_reg[10]/P0001  & n4757 ;
  assign n4808 = ~n4796 & ~n4797 ;
  assign n4782 = ~\core_c_dec_BR_Ed_reg/P0001  & ~n4656 ;
  assign n4783 = \core_c_dec_BR_Ed_reg/P0001  & \core_c_psq_Taddr_Eb_reg[7]/P0001  ;
  assign n4784 = ~n4782 & ~n4783 ;
  assign n4798 = ~\core_c_psq_DRA_reg[7]/P0001  & ~n4784 ;
  assign n4759 = ~\core_c_dec_BR_Ed_reg/P0001  & ~n4244 ;
  assign n4760 = \core_c_dec_BR_Ed_reg/P0001  & \core_c_psq_Taddr_Eb_reg[5]/P0001  ;
  assign n4761 = ~n4759 & ~n4760 ;
  assign n4799 = ~\core_c_psq_DRA_reg[5]/P0001  & ~n4761 ;
  assign n4809 = ~n4798 & ~n4799 ;
  assign n4810 = n4808 & n4809 ;
  assign n4776 = ~\core_c_dec_BR_Ed_reg/P0001  & ~n4328 ;
  assign n4777 = \core_c_dec_BR_Ed_reg/P0001  & \core_c_psq_Taddr_Eb_reg[3]/P0001  ;
  assign n4778 = ~n4776 & ~n4777 ;
  assign n4780 = ~\core_c_psq_DRA_reg[3]/P0001  & ~n4778 ;
  assign n4726 = \core_c_dec_BR_Ed_reg/P0001  & \core_c_psq_Taddr_Eb_reg[0]/P0001  ;
  assign n4727 = ~\core_c_dec_BR_Ed_reg/P0001  & ~n4588 ;
  assign n4728 = ~n4726 & ~n4727 ;
  assign n4781 = \core_c_psq_DRA_reg[0]/P0001  & n4728 ;
  assign n4806 = ~n4780 & ~n4781 ;
  assign n4785 = \core_c_psq_DRA_reg[7]/P0001  & n4784 ;
  assign n4789 = \core_c_psq_DRA_reg[13]/P0001  & n4788 ;
  assign n4807 = ~n4785 & ~n4789 ;
  assign n4811 = n4806 & n4807 ;
  assign n4764 = \core_c_dec_BR_Ed_reg/P0001  & \core_c_psq_Taddr_Eb_reg[6]/P0001  ;
  assign n4765 = ~\core_c_dec_BR_Ed_reg/P0001  & ~n4392 ;
  assign n4766 = ~n4764 & ~n4765 ;
  assign n4767 = \core_c_psq_DRA_reg[6]/P0001  & n4766 ;
  assign n4730 = ~\core_c_dec_BR_Ed_reg/P0001  & ~n4622 ;
  assign n4731 = \core_c_dec_BR_Ed_reg/P0001  & \core_c_psq_Taddr_Eb_reg[11]/P0001  ;
  assign n4732 = ~n4730 & ~n4731 ;
  assign n4774 = ~\core_c_psq_DRA_reg[11]/P0001  & ~n4732 ;
  assign n4804 = ~n4767 & ~n4774 ;
  assign n4775 = ~\core_c_psq_DRA_reg[6]/P0001  & ~n4766 ;
  assign n4779 = \core_c_psq_DRA_reg[3]/P0001  & n4778 ;
  assign n4805 = ~n4775 & ~n4779 ;
  assign n4812 = n4804 & n4805 ;
  assign n4819 = n4811 & n4812 ;
  assign n4820 = n4810 & n4819 ;
  assign n4743 = \core_c_dec_BR_Ed_reg/P0001  & ~\core_c_psq_Taddr_Eb_reg[4]/P0001  ;
  assign n4744 = ~\core_c_dec_BR_Ed_reg/P0001  & n4360 ;
  assign n4745 = ~n4743 & ~n4744 ;
  assign n4746 = ~\core_c_psq_DRA_reg[4]/P0001  & ~n4745 ;
  assign n4747 = \core_c_psq_DRA_reg[4]/P0001  & n4745 ;
  assign n4748 = ~n4746 & ~n4747 ;
  assign n4749 = \core_c_dec_BR_Ed_reg/P0001  & ~\core_c_psq_Taddr_Eb_reg[2]/P0001  ;
  assign n4750 = ~\core_c_dec_BR_Ed_reg/P0001  & n4521 ;
  assign n4751 = ~n4749 & ~n4750 ;
  assign n4752 = ~\core_c_psq_DRA_reg[2]/P0001  & ~n4751 ;
  assign n4753 = \core_c_psq_DRA_reg[2]/P0001  & n4751 ;
  assign n4754 = ~n4752 & ~n4753 ;
  assign n4815 = ~n4748 & ~n4754 ;
  assign n4768 = ~\core_c_dec_BR_Ed_reg/P0001  & ~n4457 ;
  assign n4769 = \core_c_dec_BR_Ed_reg/P0001  & \core_c_psq_Taddr_Eb_reg[1]/P0001  ;
  assign n4770 = ~n4768 & ~n4769 ;
  assign n4771 = \core_c_psq_DRA_reg[1]/P0001  & ~n4770 ;
  assign n4772 = ~\core_c_psq_DRA_reg[1]/P0001  & n4770 ;
  assign n4773 = ~n4771 & ~n4772 ;
  assign n4790 = \core_c_dec_BR_Ed_reg/P0001  & \core_c_psq_Taddr_Eb_reg[12]/P0001  ;
  assign n4791 = ~\core_c_dec_BR_Ed_reg/P0001  & ~n4694 ;
  assign n4792 = ~n4790 & ~n4791 ;
  assign n4793 = \core_c_psq_DRA_reg[12]/P0001  & ~n4792 ;
  assign n4794 = ~\core_c_psq_DRA_reg[12]/P0001  & n4792 ;
  assign n4795 = ~n4793 & ~n4794 ;
  assign n4816 = ~n4773 & ~n4795 ;
  assign n4817 = n4815 & n4816 ;
  assign n4739 = \core_c_dec_BR_Ed_reg/P0001  & \core_c_psq_Taddr_Eb_reg[9]/P0001  ;
  assign n4740 = ~\core_c_dec_BR_Ed_reg/P0001  & ~n4554 ;
  assign n4741 = ~n4739 & ~n4740 ;
  assign n4742 = ~\core_c_psq_DRA_reg[9]/P0001  & ~n4741 ;
  assign n4758 = ~\core_c_psq_DRA_reg[10]/P0001  & ~n4757 ;
  assign n4802 = ~n4742 & ~n4758 ;
  assign n4762 = \core_c_psq_DRA_reg[5]/P0001  & n4761 ;
  assign n4763 = \core_c_psq_DRA_reg[9]/P0001  & n4741 ;
  assign n4803 = ~n4762 & ~n4763 ;
  assign n4813 = n4802 & n4803 ;
  assign n4729 = ~\core_c_psq_DRA_reg[0]/P0001  & ~n4728 ;
  assign n4733 = \core_c_psq_DRA_reg[11]/P0001  & n4732 ;
  assign n4800 = ~n4729 & ~n4733 ;
  assign n4734 = ~\core_c_dec_BR_Ed_reg/P0001  & ~n4425 ;
  assign n4735 = \core_c_dec_BR_Ed_reg/P0001  & \core_c_psq_Taddr_Eb_reg[8]/P0001  ;
  assign n4736 = ~n4734 & ~n4735 ;
  assign n4737 = \core_c_psq_DRA_reg[8]/P0001  & n4736 ;
  assign n4738 = ~\core_c_psq_DRA_reg[8]/P0001  & ~n4736 ;
  assign n4801 = ~n4737 & ~n4738 ;
  assign n4814 = n4800 & n4801 ;
  assign n4818 = n4813 & n4814 ;
  assign n4821 = n4817 & n4818 ;
  assign n4822 = n4297 & n4821 ;
  assign n4823 = n4820 & n4822 ;
  assign n4824 = ~\core_c_dec_Nseq_Ed_reg/P0001  & ~n4823 ;
  assign n4825 = ~n4184 & ~n4824 ;
  assign n4826 = n4130 & ~n4825 ;
  assign n4827 = ~\core_c_dec_Nrti_Ed_reg/P0001  & ~\core_c_dec_RTI_Ed_reg/P0001  ;
  assign n4828 = ~n4826 & n4827 ;
  assign n4829 = ~n4725 & ~n4828 ;
  assign n4129 = ~\core_c_psq_TRAP_Eg_reg/NET0131  & n4105 ;
  assign n4185 = \core_c_dec_Nseq_Ed_reg/P0001  & ~n4184 ;
  assign n4839 = n4129 & n4185 ;
  assign n4840 = n4829 & n4839 ;
  assign n5052 = ~\core_c_dec_BR_Ed_reg/P0001  & n4840 ;
  assign n5053 = ~\core_c_dec_Long_Eg_reg/P0001  & ~n4829 ;
  assign n4844 = ~\core_c_dec_EXIT_E_reg/P0001  & ~\core_c_psq_PCS_reg[7]/NET0131  ;
  assign n4845 = ~\core_c_psq_lpstk_ptr_reg[0]/NET0131  & ~\core_c_psq_lpstk_ptr_reg[1]/NET0131  ;
  assign n4879 = \core_c_psq_lpstk_lps4x22_LPcell_reg[0][14]/P0001  & n4845 ;
  assign n4847 = \core_c_psq_lpstk_ptr_reg[0]/NET0131  & ~\core_c_psq_lpstk_ptr_reg[1]/NET0131  ;
  assign n4880 = \core_c_psq_lpstk_lps4x22_LPcell_reg[1][14]/P0001  & n4847 ;
  assign n4883 = ~n4879 & ~n4880 ;
  assign n4849 = \core_c_psq_lpstk_ptr_reg[0]/NET0131  & \core_c_psq_lpstk_ptr_reg[1]/NET0131  ;
  assign n4881 = \core_c_psq_lpstk_lps4x22_LPcell_reg[3][14]/P0001  & n4849 ;
  assign n4851 = ~\core_c_psq_lpstk_ptr_reg[0]/NET0131  & \core_c_psq_lpstk_ptr_reg[1]/NET0131  ;
  assign n4882 = \core_c_psq_lpstk_lps4x22_LPcell_reg[2][14]/P0001  & n4851 ;
  assign n4884 = ~n4881 & ~n4882 ;
  assign n4885 = n4883 & n4884 ;
  assign n4886 = \core_c_psq_IFA_reg[10]/P0001  & ~n4885 ;
  assign n4887 = ~\core_c_psq_IFA_reg[10]/P0001  & n4885 ;
  assign n4888 = ~n4886 & ~n4887 ;
  assign n4889 = \core_c_psq_lpstk_lps4x22_LPcell_reg[0][21]/P0001  & n4845 ;
  assign n4890 = \core_c_psq_lpstk_lps4x22_LPcell_reg[1][21]/P0001  & n4847 ;
  assign n4893 = ~n4889 & ~n4890 ;
  assign n4891 = \core_c_psq_lpstk_lps4x22_LPcell_reg[3][21]/P0001  & n4849 ;
  assign n4892 = \core_c_psq_lpstk_lps4x22_LPcell_reg[2][21]/P0001  & n4851 ;
  assign n4894 = ~n4891 & ~n4892 ;
  assign n4895 = n4893 & n4894 ;
  assign n4896 = \core_c_psq_PMOVL_regl_DO_reg[3]/NET0131  & ~n4895 ;
  assign n4897 = ~\core_c_psq_PMOVL_regl_DO_reg[3]/NET0131  & n4895 ;
  assign n4898 = ~n4896 & ~n4897 ;
  assign n5031 = ~n4888 & ~n4898 ;
  assign n4899 = \core_c_psq_lpstk_lps4x22_LPcell_reg[0][20]/P0001  & n4845 ;
  assign n4900 = \core_c_psq_lpstk_lps4x22_LPcell_reg[1][20]/P0001  & n4847 ;
  assign n4903 = ~n4899 & ~n4900 ;
  assign n4901 = \core_c_psq_lpstk_lps4x22_LPcell_reg[3][20]/P0001  & n4849 ;
  assign n4902 = \core_c_psq_lpstk_lps4x22_LPcell_reg[2][20]/P0001  & n4851 ;
  assign n4904 = ~n4901 & ~n4902 ;
  assign n4905 = n4903 & n4904 ;
  assign n4906 = \core_c_psq_PMOVL_regl_DO_reg[2]/NET0131  & ~n4905 ;
  assign n4907 = ~\core_c_psq_PMOVL_regl_DO_reg[2]/NET0131  & n4905 ;
  assign n4908 = ~n4906 & ~n4907 ;
  assign n4909 = \core_c_psq_lpstk_lps4x22_LPcell_reg[2][17]/P0001  & n4851 ;
  assign n4910 = \core_c_psq_lpstk_lps4x22_LPcell_reg[3][17]/P0001  & n4849 ;
  assign n4913 = ~n4909 & ~n4910 ;
  assign n4911 = \core_c_psq_lpstk_lps4x22_LPcell_reg[1][17]/P0001  & n4847 ;
  assign n4912 = \core_c_psq_lpstk_lps4x22_LPcell_reg[0][17]/P0001  & n4845 ;
  assign n4914 = ~n4911 & ~n4912 ;
  assign n4915 = n4913 & n4914 ;
  assign n4916 = \core_c_psq_IFA_reg[13]/P0001  & ~n4915 ;
  assign n4917 = ~\core_c_psq_IFA_reg[13]/P0001  & n4915 ;
  assign n4918 = ~n4916 & ~n4917 ;
  assign n5032 = ~n4908 & ~n4918 ;
  assign n5041 = n5031 & n5032 ;
  assign n4846 = \core_c_psq_lpstk_lps4x22_LPcell_reg[0][19]/P0001  & n4845 ;
  assign n4848 = \core_c_psq_lpstk_lps4x22_LPcell_reg[1][19]/P0001  & n4847 ;
  assign n4853 = ~n4846 & ~n4848 ;
  assign n4850 = \core_c_psq_lpstk_lps4x22_LPcell_reg[3][19]/P0001  & n4849 ;
  assign n4852 = \core_c_psq_lpstk_lps4x22_LPcell_reg[2][19]/P0001  & n4851 ;
  assign n4854 = ~n4850 & ~n4852 ;
  assign n4855 = n4853 & n4854 ;
  assign n4856 = \core_c_psq_PMOVL_regl_DO_reg[1]/NET0131  & ~n4855 ;
  assign n4857 = ~\core_c_psq_PMOVL_regl_DO_reg[1]/NET0131  & n4855 ;
  assign n4858 = ~n4856 & ~n4857 ;
  assign n5029 = ~\core_c_psq_lpstk_ptr_reg[2]/NET0131  & ~n4858 ;
  assign n4859 = \core_c_psq_lpstk_lps4x22_LPcell_reg[0][18]/P0001  & n4845 ;
  assign n4860 = \core_c_psq_lpstk_lps4x22_LPcell_reg[1][18]/P0001  & n4847 ;
  assign n4863 = ~n4859 & ~n4860 ;
  assign n4861 = \core_c_psq_lpstk_lps4x22_LPcell_reg[3][18]/P0001  & n4849 ;
  assign n4862 = \core_c_psq_lpstk_lps4x22_LPcell_reg[2][18]/P0001  & n4851 ;
  assign n4864 = ~n4861 & ~n4862 ;
  assign n4865 = n4863 & n4864 ;
  assign n4866 = \core_c_psq_PMOVL_regl_DO_reg[0]/NET0131  & ~n4865 ;
  assign n4867 = ~\core_c_psq_PMOVL_regl_DO_reg[0]/NET0131  & n4865 ;
  assign n4868 = ~n4866 & ~n4867 ;
  assign n4869 = \core_c_psq_lpstk_lps4x22_LPcell_reg[0][13]/P0001  & n4845 ;
  assign n4870 = \core_c_psq_lpstk_lps4x22_LPcell_reg[1][13]/P0001  & n4847 ;
  assign n4873 = ~n4869 & ~n4870 ;
  assign n4871 = \core_c_psq_lpstk_lps4x22_LPcell_reg[3][13]/P0001  & n4849 ;
  assign n4872 = \core_c_psq_lpstk_lps4x22_LPcell_reg[2][13]/P0001  & n4851 ;
  assign n4874 = ~n4871 & ~n4872 ;
  assign n4875 = n4873 & n4874 ;
  assign n4876 = \core_c_psq_IFA_reg[9]/P0001  & ~n4875 ;
  assign n4877 = ~\core_c_psq_IFA_reg[9]/P0001  & n4875 ;
  assign n4878 = ~n4876 & ~n4877 ;
  assign n5030 = ~n4868 & ~n4878 ;
  assign n5042 = n5029 & n5030 ;
  assign n5043 = n5041 & n5042 ;
  assign n5019 = \core_c_psq_lpstk_lps4x22_LPcell_reg[0][10]/P0001  & n4845 ;
  assign n5020 = \core_c_psq_lpstk_lps4x22_LPcell_reg[1][10]/P0001  & n4847 ;
  assign n5023 = ~n5019 & ~n5020 ;
  assign n5021 = \core_c_psq_lpstk_lps4x22_LPcell_reg[3][10]/P0001  & n4849 ;
  assign n5022 = \core_c_psq_lpstk_lps4x22_LPcell_reg[2][10]/P0001  & n4851 ;
  assign n5024 = ~n5021 & ~n5022 ;
  assign n5025 = n5023 & n5024 ;
  assign n5026 = \core_c_psq_IFA_reg[6]/P0001  & ~n5025 ;
  assign n5027 = ~\core_c_psq_IFA_reg[6]/P0001  & n5025 ;
  assign n5028 = ~n5026 & ~n5027 ;
  assign n4999 = \core_c_psq_lpstk_lps4x22_LPcell_reg[0][12]/P0001  & n4845 ;
  assign n5000 = \core_c_psq_lpstk_lps4x22_LPcell_reg[1][12]/P0001  & n4847 ;
  assign n5003 = ~n4999 & ~n5000 ;
  assign n5001 = \core_c_psq_lpstk_lps4x22_LPcell_reg[3][12]/P0001  & n4849 ;
  assign n5002 = \core_c_psq_lpstk_lps4x22_LPcell_reg[2][12]/P0001  & n4851 ;
  assign n5004 = ~n5001 & ~n5002 ;
  assign n5005 = n5003 & n5004 ;
  assign n5006 = \core_c_psq_IFA_reg[8]/P0001  & ~n5005 ;
  assign n5007 = ~\core_c_psq_IFA_reg[8]/P0001  & n5005 ;
  assign n5008 = ~n5006 & ~n5007 ;
  assign n5009 = \core_c_psq_lpstk_lps4x22_LPcell_reg[2][11]/P0001  & n4851 ;
  assign n5010 = \core_c_psq_lpstk_lps4x22_LPcell_reg[3][11]/P0001  & n4849 ;
  assign n5013 = ~n5009 & ~n5010 ;
  assign n5011 = \core_c_psq_lpstk_lps4x22_LPcell_reg[1][11]/P0001  & n4847 ;
  assign n5012 = \core_c_psq_lpstk_lps4x22_LPcell_reg[0][11]/P0001  & n4845 ;
  assign n5014 = ~n5011 & ~n5012 ;
  assign n5015 = n5013 & n5014 ;
  assign n5016 = \core_c_psq_IFA_reg[7]/P0001  & ~n5015 ;
  assign n5017 = ~\core_c_psq_IFA_reg[7]/P0001  & n5015 ;
  assign n5018 = ~n5016 & ~n5017 ;
  assign n5037 = ~n5008 & ~n5018 ;
  assign n5038 = ~n5028 & n5037 ;
  assign n4959 = \core_c_psq_lpstk_lps4x22_LPcell_reg[0][4]/P0001  & n4845 ;
  assign n4960 = \core_c_psq_lpstk_lps4x22_LPcell_reg[1][4]/P0001  & n4847 ;
  assign n4963 = ~n4959 & ~n4960 ;
  assign n4961 = \core_c_psq_lpstk_lps4x22_LPcell_reg[3][4]/P0001  & n4849 ;
  assign n4962 = \core_c_psq_lpstk_lps4x22_LPcell_reg[2][4]/P0001  & n4851 ;
  assign n4964 = ~n4961 & ~n4962 ;
  assign n4965 = n4963 & n4964 ;
  assign n4966 = \core_c_psq_IFA_reg[0]/P0001  & ~n4965 ;
  assign n4967 = ~\core_c_psq_IFA_reg[0]/P0001  & n4965 ;
  assign n4968 = ~n4966 & ~n4967 ;
  assign n4969 = \core_c_psq_lpstk_lps4x22_LPcell_reg[0][8]/P0001  & n4845 ;
  assign n4970 = \core_c_psq_lpstk_lps4x22_LPcell_reg[1][8]/P0001  & n4847 ;
  assign n4973 = ~n4969 & ~n4970 ;
  assign n4971 = \core_c_psq_lpstk_lps4x22_LPcell_reg[3][8]/P0001  & n4849 ;
  assign n4972 = \core_c_psq_lpstk_lps4x22_LPcell_reg[2][8]/P0001  & n4851 ;
  assign n4974 = ~n4971 & ~n4972 ;
  assign n4975 = n4973 & n4974 ;
  assign n4976 = \core_c_psq_IFA_reg[4]/P0001  & ~n4975 ;
  assign n4977 = ~\core_c_psq_IFA_reg[4]/P0001  & n4975 ;
  assign n4978 = ~n4976 & ~n4977 ;
  assign n5035 = ~n4968 & ~n4978 ;
  assign n4979 = \core_c_psq_lpstk_lps4x22_LPcell_reg[0][6]/P0001  & n4845 ;
  assign n4980 = \core_c_psq_lpstk_lps4x22_LPcell_reg[1][6]/P0001  & n4847 ;
  assign n4983 = ~n4979 & ~n4980 ;
  assign n4981 = \core_c_psq_lpstk_lps4x22_LPcell_reg[3][6]/P0001  & n4849 ;
  assign n4982 = \core_c_psq_lpstk_lps4x22_LPcell_reg[2][6]/P0001  & n4851 ;
  assign n4984 = ~n4981 & ~n4982 ;
  assign n4985 = n4983 & n4984 ;
  assign n4986 = \core_c_psq_IFA_reg[2]/P0001  & ~n4985 ;
  assign n4987 = ~\core_c_psq_IFA_reg[2]/P0001  & n4985 ;
  assign n4988 = ~n4986 & ~n4987 ;
  assign n4989 = \core_c_psq_lpstk_lps4x22_LPcell_reg[2][5]/P0001  & n4851 ;
  assign n4990 = \core_c_psq_lpstk_lps4x22_LPcell_reg[3][5]/P0001  & n4849 ;
  assign n4993 = ~n4989 & ~n4990 ;
  assign n4991 = \core_c_psq_lpstk_lps4x22_LPcell_reg[0][5]/P0001  & n4845 ;
  assign n4992 = \core_c_psq_lpstk_lps4x22_LPcell_reg[1][5]/P0001  & n4847 ;
  assign n4994 = ~n4991 & ~n4992 ;
  assign n4995 = n4993 & n4994 ;
  assign n4996 = \core_c_psq_IFA_reg[1]/P0001  & ~n4995 ;
  assign n4997 = ~\core_c_psq_IFA_reg[1]/P0001  & n4995 ;
  assign n4998 = ~n4996 & ~n4997 ;
  assign n5036 = ~n4988 & ~n4998 ;
  assign n5039 = n5035 & n5036 ;
  assign n4919 = \core_c_psq_lpstk_lps4x22_LPcell_reg[0][16]/P0001  & n4845 ;
  assign n4920 = \core_c_psq_lpstk_lps4x22_LPcell_reg[1][16]/P0001  & n4847 ;
  assign n4923 = ~n4919 & ~n4920 ;
  assign n4921 = \core_c_psq_lpstk_lps4x22_LPcell_reg[3][16]/P0001  & n4849 ;
  assign n4922 = \core_c_psq_lpstk_lps4x22_LPcell_reg[2][16]/P0001  & n4851 ;
  assign n4924 = ~n4921 & ~n4922 ;
  assign n4925 = n4923 & n4924 ;
  assign n4926 = \core_c_psq_IFA_reg[12]/P0001  & ~n4925 ;
  assign n4927 = ~\core_c_psq_IFA_reg[12]/P0001  & n4925 ;
  assign n4928 = ~n4926 & ~n4927 ;
  assign n4929 = \core_c_psq_lpstk_lps4x22_LPcell_reg[2][15]/P0001  & n4851 ;
  assign n4930 = \core_c_psq_lpstk_lps4x22_LPcell_reg[3][15]/P0001  & n4849 ;
  assign n4933 = ~n4929 & ~n4930 ;
  assign n4931 = \core_c_psq_lpstk_lps4x22_LPcell_reg[1][15]/P0001  & n4847 ;
  assign n4932 = \core_c_psq_lpstk_lps4x22_LPcell_reg[0][15]/P0001  & n4845 ;
  assign n4934 = ~n4931 & ~n4932 ;
  assign n4935 = n4933 & n4934 ;
  assign n4936 = \core_c_psq_IFA_reg[11]/P0001  & ~n4935 ;
  assign n4937 = ~\core_c_psq_IFA_reg[11]/P0001  & n4935 ;
  assign n4938 = ~n4936 & ~n4937 ;
  assign n5033 = ~n4928 & ~n4938 ;
  assign n4939 = \core_c_psq_lpstk_lps4x22_LPcell_reg[0][9]/P0001  & n4845 ;
  assign n4940 = \core_c_psq_lpstk_lps4x22_LPcell_reg[1][9]/P0001  & n4847 ;
  assign n4943 = ~n4939 & ~n4940 ;
  assign n4941 = \core_c_psq_lpstk_lps4x22_LPcell_reg[3][9]/P0001  & n4849 ;
  assign n4942 = \core_c_psq_lpstk_lps4x22_LPcell_reg[2][9]/P0001  & n4851 ;
  assign n4944 = ~n4941 & ~n4942 ;
  assign n4945 = n4943 & n4944 ;
  assign n4946 = \core_c_psq_IFA_reg[5]/P0001  & ~n4945 ;
  assign n4947 = ~\core_c_psq_IFA_reg[5]/P0001  & n4945 ;
  assign n4948 = ~n4946 & ~n4947 ;
  assign n4949 = \core_c_psq_lpstk_lps4x22_LPcell_reg[0][7]/P0001  & n4845 ;
  assign n4950 = \core_c_psq_lpstk_lps4x22_LPcell_reg[1][7]/P0001  & n4847 ;
  assign n4953 = ~n4949 & ~n4950 ;
  assign n4951 = \core_c_psq_lpstk_lps4x22_LPcell_reg[3][7]/P0001  & n4849 ;
  assign n4952 = \core_c_psq_lpstk_lps4x22_LPcell_reg[2][7]/P0001  & n4851 ;
  assign n4954 = ~n4951 & ~n4952 ;
  assign n4955 = n4953 & n4954 ;
  assign n4956 = \core_c_psq_IFA_reg[3]/P0001  & ~n4955 ;
  assign n4957 = ~\core_c_psq_IFA_reg[3]/P0001  & n4955 ;
  assign n4958 = ~n4956 & ~n4957 ;
  assign n5034 = ~n4948 & ~n4958 ;
  assign n5040 = n5033 & n5034 ;
  assign n5044 = n5039 & n5040 ;
  assign n5045 = n5038 & n5044 ;
  assign n5046 = n5043 & n5045 ;
  assign n5055 = n4844 & n5046 ;
  assign n5056 = n5053 & ~n5055 ;
  assign n4186 = n4130 & ~n4185 ;
  assign n4830 = n4186 & n4297 ;
  assign n5054 = ~n4830 & ~n5053 ;
  assign n5057 = n4129 & ~n5054 ;
  assign n5058 = ~n5056 & n5057 ;
  assign n5059 = ~n5052 & ~n5058 ;
  assign n5060 = ~n4588 & ~n5059 ;
  assign n4831 = ~n4185 & ~n4830 ;
  assign n4832 = n4829 & n4831 ;
  assign n4187 = \core_c_dec_Long_Eg_reg/P0001  & ~n4186 ;
  assign n4833 = ~\core_c_psq_PCS_reg[7]/NET0131  & ~n4187 ;
  assign n4834 = ~n4832 & n4833 ;
  assign n4835 = n4129 & ~n4834 ;
  assign n4836 = ~\core_c_psq_EXA_reg[0]/P0001  & n4835 ;
  assign n4842 = n4186 & ~n4297 ;
  assign n4843 = \core_c_dec_Long_Eg_reg/P0001  & ~n4842 ;
  assign n5047 = n4129 & n4844 ;
  assign n5048 = ~n5046 & n5047 ;
  assign n5049 = ~n4843 & n5048 ;
  assign n5050 = ~n4829 & n5049 ;
  assign n5051 = ~\core_c_psq_IFA_reg[0]/P0001  & n5050 ;
  assign n4837 = \core_c_dec_EXIT_E_reg/P0001  & n4129 ;
  assign n4838 = \sice_IRR_reg[0]/P0001  & n4837 ;
  assign n4841 = n4726 & n4840 ;
  assign n5061 = ~n4838 & ~n4841 ;
  assign n5062 = ~n5051 & n5061 ;
  assign n5063 = ~n4836 & n5062 ;
  assign n5064 = ~n5060 & n5063 ;
  assign n5065 = n4128 & ~n5064 ;
  assign n4120 = ~n4099 & ~n4119 ;
  assign n4121 = ~\core_c_dec_IR_reg[4]/NET0131  & ~n4117 ;
  assign n4122 = ~\core_c_dec_IRE_reg[4]/NET0131  & n4117 ;
  assign n4123 = ~n4121 & ~n4122 ;
  assign n4124 = ~n4104 & ~n4123 ;
  assign n4125 = ~\core_c_psq_IFA_reg[0]/P0001  & n4104 ;
  assign n4126 = ~n4124 & ~n4125 ;
  assign n4127 = n4120 & n4126 ;
  assign n5066 = n4048 & n4056 ;
  assign n5067 = \bdma_BIAD_reg[0]/NET0131  & n5066 ;
  assign n5068 = \idma_DSreq_reg/NET0131  & n4055 ;
  assign n5069 = \idma_DCTL_reg[0]/NET0131  & n5068 ;
  assign n5070 = ~n5067 & ~n5069 ;
  assign n5071 = n4099 & ~n5070 ;
  assign n5072 = ~n4127 & ~n5071 ;
  assign n5073 = ~n5065 & n5072 ;
  assign n5081 = ~n4276 & ~n5059 ;
  assign n5082 = \core_c_psq_EXA_reg[0]/P0001  & \core_c_psq_EXA_reg[1]/P0001  ;
  assign n5083 = \core_c_psq_EXA_reg[2]/P0001  & n5082 ;
  assign n5084 = \core_c_psq_EXA_reg[3]/P0001  & n5083 ;
  assign n5085 = \core_c_psq_EXA_reg[4]/P0001  & n5084 ;
  assign n5086 = \core_c_psq_EXA_reg[5]/P0001  & n5085 ;
  assign n5087 = \core_c_psq_EXA_reg[6]/P0001  & n5086 ;
  assign n5088 = \core_c_psq_EXA_reg[7]/P0001  & n5087 ;
  assign n5089 = \core_c_psq_EXA_reg[8]/P0001  & n5088 ;
  assign n5090 = \core_c_psq_EXA_reg[9]/P0001  & n5089 ;
  assign n5091 = ~\core_c_psq_EXA_reg[10]/P0001  & ~n5090 ;
  assign n5092 = \core_c_psq_EXA_reg[10]/P0001  & n5090 ;
  assign n5093 = ~n5091 & ~n5092 ;
  assign n5094 = n4835 & n5093 ;
  assign n5108 = n4755 & n4840 ;
  assign n5095 = \core_c_psq_IFA_reg[0]/P0001  & \core_c_psq_IFA_reg[1]/P0001  ;
  assign n5096 = \core_c_psq_IFA_reg[2]/P0001  & n5095 ;
  assign n5097 = \core_c_psq_IFA_reg[3]/P0001  & n5096 ;
  assign n5098 = \core_c_psq_IFA_reg[4]/P0001  & n5097 ;
  assign n5099 = \core_c_psq_IFA_reg[5]/P0001  & n5098 ;
  assign n5100 = \core_c_psq_IFA_reg[6]/P0001  & n5099 ;
  assign n5101 = \core_c_psq_IFA_reg[7]/P0001  & n5100 ;
  assign n5102 = \core_c_psq_IFA_reg[8]/P0001  & n5101 ;
  assign n5103 = \core_c_psq_IFA_reg[9]/P0001  & n5102 ;
  assign n5104 = ~\core_c_psq_IFA_reg[10]/P0001  & ~n5103 ;
  assign n5105 = \core_c_psq_IFA_reg[10]/P0001  & n5103 ;
  assign n5106 = ~n5104 & ~n5105 ;
  assign n5107 = n5050 & n5106 ;
  assign n5109 = \sice_IRR_reg[10]/P0001  & n4837 ;
  assign n5110 = ~n5107 & ~n5109 ;
  assign n5111 = ~n5108 & n5110 ;
  assign n5112 = ~n5094 & n5111 ;
  assign n5113 = ~n5081 & n5112 ;
  assign n5114 = n4128 & ~n5113 ;
  assign n5074 = ~\core_c_psq_IFA_reg[10]/P0001  & n4104 ;
  assign n5075 = ~\core_c_dec_IR_reg[14]/NET0131  & ~n4117 ;
  assign n5076 = ~\core_c_dec_IRE_reg[14]/NET0131  & n4117 ;
  assign n5077 = ~n5075 & ~n5076 ;
  assign n5078 = ~n4104 & ~n5077 ;
  assign n5079 = ~n5074 & ~n5078 ;
  assign n5080 = n4120 & n5079 ;
  assign n5115 = \bdma_BIAD_reg[10]/NET0131  & n5066 ;
  assign n5116 = \idma_DCTL_reg[10]/NET0131  & n5068 ;
  assign n5117 = ~n5115 & ~n5116 ;
  assign n5118 = n4099 & ~n5117 ;
  assign n5119 = ~n5080 & ~n5118 ;
  assign n5120 = ~n5114 & n5119 ;
  assign n5128 = ~n4622 & ~n5059 ;
  assign n5129 = ~\core_c_psq_EXA_reg[11]/P0001  & ~n5092 ;
  assign n5130 = \core_c_psq_EXA_reg[11]/P0001  & n5092 ;
  assign n5131 = ~n5129 & ~n5130 ;
  assign n5132 = n4835 & n5131 ;
  assign n5137 = n4731 & n4840 ;
  assign n5133 = ~\core_c_psq_IFA_reg[11]/P0001  & ~n5105 ;
  assign n5134 = \core_c_psq_IFA_reg[11]/P0001  & n5105 ;
  assign n5135 = ~n5133 & ~n5134 ;
  assign n5136 = n5050 & n5135 ;
  assign n5138 = \sice_IRR_reg[11]/P0001  & n4837 ;
  assign n5139 = ~n5136 & ~n5138 ;
  assign n5140 = ~n5137 & n5139 ;
  assign n5141 = ~n5132 & n5140 ;
  assign n5142 = ~n5128 & n5141 ;
  assign n5143 = n4128 & ~n5142 ;
  assign n5121 = ~\core_c_psq_IFA_reg[11]/P0001  & n4104 ;
  assign n5123 = \core_c_dec_IR_reg[15]/NET0131  & ~n4117 ;
  assign n5122 = \core_c_dec_IRE_reg[15]/NET0131  & n4117 ;
  assign n5124 = ~n4104 & ~n5122 ;
  assign n5125 = ~n5123 & n5124 ;
  assign n5126 = ~n5121 & ~n5125 ;
  assign n5127 = n4120 & n5126 ;
  assign n5144 = \bdma_BIAD_reg[11]/NET0131  & n5066 ;
  assign n5145 = \idma_DCTL_reg[11]/NET0131  & n5068 ;
  assign n5146 = ~n5144 & ~n5145 ;
  assign n5147 = n4099 & ~n5146 ;
  assign n5148 = ~n5127 & ~n5147 ;
  assign n5149 = ~n5143 & n5148 ;
  assign n5165 = ~n4457 & ~n5059 ;
  assign n5157 = ~\core_c_psq_EXA_reg[0]/P0001  & ~\core_c_psq_EXA_reg[1]/P0001  ;
  assign n5158 = ~n5082 & ~n5157 ;
  assign n5159 = n4835 & n5158 ;
  assign n5162 = ~\core_c_psq_IFA_reg[0]/P0001  & ~\core_c_psq_IFA_reg[1]/P0001  ;
  assign n5163 = ~n5095 & ~n5162 ;
  assign n5164 = n5050 & n5163 ;
  assign n5160 = \sice_IRR_reg[1]/P0001  & n4837 ;
  assign n5161 = n4769 & n4840 ;
  assign n5166 = ~n5160 & ~n5161 ;
  assign n5167 = ~n5164 & n5166 ;
  assign n5168 = ~n5159 & n5167 ;
  assign n5169 = ~n5165 & n5168 ;
  assign n5170 = n4128 & ~n5169 ;
  assign n5150 = ~\core_c_psq_IFA_reg[1]/P0001  & n4104 ;
  assign n5151 = ~\core_c_dec_IR_reg[5]/NET0131  & ~n4117 ;
  assign n5152 = ~\core_c_dec_IRE_reg[5]/NET0131  & n4117 ;
  assign n5153 = ~n5151 & ~n5152 ;
  assign n5154 = ~n4104 & ~n5153 ;
  assign n5155 = ~n5150 & ~n5154 ;
  assign n5156 = n4120 & n5155 ;
  assign n5171 = \bdma_BIAD_reg[1]/NET0131  & n5066 ;
  assign n5172 = \idma_DCTL_reg[1]/NET0131  & n5068 ;
  assign n5173 = ~n5171 & ~n5172 ;
  assign n5174 = n4099 & ~n5173 ;
  assign n5175 = ~n5156 & ~n5174 ;
  assign n5176 = ~n5170 & n5175 ;
  assign n5184 = ~n4521 & n5058 ;
  assign n5194 = ~\core_c_psq_EXA_reg[2]/P0001  & ~n5082 ;
  assign n5195 = ~n5083 & ~n5194 ;
  assign n5196 = n4835 & n5195 ;
  assign n5189 = \core_c_dec_BR_Ed_reg/P0001  & ~n4184 ;
  assign n5190 = ~\core_c_psq_Taddr_Eb_reg[2]/P0001  & n5189 ;
  assign n5191 = n4521 & ~n5189 ;
  assign n5192 = ~n5190 & ~n5191 ;
  assign n5193 = n4840 & n5192 ;
  assign n5186 = ~\core_c_psq_IFA_reg[2]/P0001  & ~n5095 ;
  assign n5187 = ~n5096 & ~n5186 ;
  assign n5188 = n5050 & n5187 ;
  assign n5185 = \sice_IRR_reg[2]/P0001  & n4837 ;
  assign n5197 = \core_c_psq_TRAP_Eg_reg/NET0131  & n4105 ;
  assign n5198 = ~\core_c_psq_Iact_E_reg[0]/NET0131  & ~\core_c_psq_Iact_E_reg[10]/NET0131  ;
  assign n5199 = ~\core_c_psq_Iact_E_reg[2]/NET0131  & ~\core_c_psq_Iact_E_reg[4]/NET0131  ;
  assign n5200 = ~\core_c_psq_Iact_E_reg[6]/NET0131  & ~\core_c_psq_Iact_E_reg[8]/NET0131  ;
  assign n5201 = n5199 & n5200 ;
  assign n5202 = n5198 & n5201 ;
  assign n5203 = n5197 & ~n5202 ;
  assign n5204 = ~n5185 & ~n5203 ;
  assign n5205 = ~n5188 & n5204 ;
  assign n5206 = ~n5193 & n5205 ;
  assign n5207 = ~n5196 & n5206 ;
  assign n5208 = ~n5184 & n5207 ;
  assign n5209 = n4128 & ~n5208 ;
  assign n5177 = ~\core_c_psq_IFA_reg[2]/P0001  & n4104 ;
  assign n5178 = ~\core_c_dec_IR_reg[6]/NET0131  & ~n4117 ;
  assign n5179 = ~\core_c_dec_IRE_reg[6]/NET0131  & n4117 ;
  assign n5180 = ~n5178 & ~n5179 ;
  assign n5181 = ~n4104 & ~n5180 ;
  assign n5182 = ~n5177 & ~n5181 ;
  assign n5183 = n4120 & n5182 ;
  assign n5210 = \bdma_BIAD_reg[2]/NET0131  & n5066 ;
  assign n5211 = \idma_DCTL_reg[2]/NET0131  & n5068 ;
  assign n5212 = ~n5210 & ~n5211 ;
  assign n5213 = n4099 & ~n5212 ;
  assign n5214 = ~n5183 & ~n5213 ;
  assign n5215 = ~n5209 & n5214 ;
  assign n5223 = ~n4328 & n5058 ;
  assign n5232 = ~\core_c_psq_EXA_reg[3]/P0001  & ~n5083 ;
  assign n5233 = ~n5084 & ~n5232 ;
  assign n5234 = n4835 & n5233 ;
  assign n5228 = ~\core_c_psq_Taddr_Eb_reg[3]/P0001  & n5189 ;
  assign n5229 = n4328 & ~n5189 ;
  assign n5230 = ~n5228 & ~n5229 ;
  assign n5231 = n4840 & n5230 ;
  assign n5225 = ~\core_c_psq_IFA_reg[3]/P0001  & ~n5096 ;
  assign n5226 = ~n5097 & ~n5225 ;
  assign n5227 = n5050 & n5226 ;
  assign n5224 = \sice_IRR_reg[3]/P0001  & n4837 ;
  assign n5235 = ~\core_c_psq_Iact_E_reg[2]/NET0131  & ~\core_c_psq_Iact_E_reg[5]/NET0131  ;
  assign n5236 = ~\core_c_psq_Iact_E_reg[10]/NET0131  & ~\core_c_psq_Iact_E_reg[1]/NET0131  ;
  assign n5237 = ~\core_c_psq_Iact_E_reg[6]/NET0131  & ~\core_c_psq_Iact_E_reg[9]/NET0131  ;
  assign n5238 = n5236 & n5237 ;
  assign n5239 = n5235 & n5238 ;
  assign n5240 = n5197 & ~n5239 ;
  assign n5241 = ~n5224 & ~n5240 ;
  assign n5242 = ~n5227 & n5241 ;
  assign n5243 = ~n5231 & n5242 ;
  assign n5244 = ~n5234 & n5243 ;
  assign n5245 = ~n5223 & n5244 ;
  assign n5246 = n4128 & ~n5245 ;
  assign n5216 = ~\core_c_psq_IFA_reg[3]/P0001  & n4104 ;
  assign n5217 = ~\core_c_dec_IR_reg[7]/NET0131  & ~n4117 ;
  assign n5218 = ~\core_c_dec_IRE_reg[7]/NET0131  & n4117 ;
  assign n5219 = ~n5217 & ~n5218 ;
  assign n5220 = ~n4104 & ~n5219 ;
  assign n5221 = ~n5216 & ~n5220 ;
  assign n5222 = n4120 & n5221 ;
  assign n5247 = \bdma_BIAD_reg[3]/NET0131  & n5066 ;
  assign n5248 = \idma_DCTL_reg[3]/NET0131  & n5068 ;
  assign n5249 = ~n5247 & ~n5248 ;
  assign n5250 = n4099 & ~n5249 ;
  assign n5251 = ~n5222 & ~n5250 ;
  assign n5252 = ~n5246 & n5251 ;
  assign n5260 = ~n4360 & n5058 ;
  assign n5269 = ~\core_c_psq_EXA_reg[4]/P0001  & ~n5084 ;
  assign n5270 = ~n5085 & ~n5269 ;
  assign n5271 = n4835 & n5270 ;
  assign n5265 = ~\core_c_psq_Taddr_Eb_reg[4]/P0001  & n5189 ;
  assign n5266 = n4360 & ~n5189 ;
  assign n5267 = ~n5265 & ~n5266 ;
  assign n5268 = n4840 & n5267 ;
  assign n5262 = ~\core_c_psq_IFA_reg[4]/P0001  & ~n5097 ;
  assign n5263 = ~n5098 & ~n5262 ;
  assign n5264 = n5050 & n5263 ;
  assign n5261 = \sice_IRR_reg[4]/P0001  & n4837 ;
  assign n5272 = ~\core_c_psq_Iact_E_reg[4]/NET0131  & ~\core_c_psq_Iact_E_reg[7]/NET0131  ;
  assign n5273 = n5235 & n5272 ;
  assign n5274 = n5197 & ~n5273 ;
  assign n5275 = ~n5261 & ~n5274 ;
  assign n5276 = ~n5264 & n5275 ;
  assign n5277 = ~n5268 & n5276 ;
  assign n5278 = ~n5271 & n5277 ;
  assign n5279 = ~n5260 & n5278 ;
  assign n5280 = n4128 & ~n5279 ;
  assign n5253 = ~\core_c_psq_IFA_reg[4]/P0001  & n4104 ;
  assign n5254 = ~\core_c_dec_IR_reg[8]/NET0131  & ~n4117 ;
  assign n5255 = ~\core_c_dec_IRE_reg[8]/NET0131  & n4117 ;
  assign n5256 = ~n5254 & ~n5255 ;
  assign n5257 = ~n4104 & ~n5256 ;
  assign n5258 = ~n5253 & ~n5257 ;
  assign n5259 = n4120 & n5258 ;
  assign n5281 = \bdma_BIAD_reg[4]/NET0131  & n5066 ;
  assign n5282 = \idma_DCTL_reg[4]/NET0131  & n5068 ;
  assign n5283 = ~n5281 & ~n5282 ;
  assign n5284 = n4099 & ~n5283 ;
  assign n5285 = ~n5259 & ~n5284 ;
  assign n5286 = ~n5280 & n5285 ;
  assign n5294 = ~n4244 & ~n5059 ;
  assign n5303 = ~\core_c_psq_EXA_reg[5]/P0001  & ~n5085 ;
  assign n5304 = ~n5086 & ~n5303 ;
  assign n5305 = n4835 & n5304 ;
  assign n5296 = ~\core_c_psq_IFA_reg[5]/P0001  & ~n5098 ;
  assign n5297 = ~n5099 & ~n5296 ;
  assign n5298 = n5050 & n5297 ;
  assign n5295 = n4760 & n4840 ;
  assign n5299 = ~\core_c_psq_Iact_E_reg[0]/NET0131  & ~\core_c_psq_Iact_E_reg[1]/NET0131  ;
  assign n5300 = ~\core_c_psq_Iact_E_reg[10]/NET0131  & ~\core_c_psq_Iact_E_reg[3]/NET0131  ;
  assign n5301 = n5299 & n5300 ;
  assign n5302 = n5197 & ~n5301 ;
  assign n5306 = \sice_IRR_reg[5]/P0001  & n4837 ;
  assign n5307 = ~n5302 & ~n5306 ;
  assign n5308 = ~n5295 & n5307 ;
  assign n5309 = ~n5298 & n5308 ;
  assign n5310 = ~n5305 & n5309 ;
  assign n5311 = ~n5294 & n5310 ;
  assign n5312 = n4128 & ~n5311 ;
  assign n5287 = ~\core_c_psq_IFA_reg[5]/P0001  & n4104 ;
  assign n5288 = ~\core_c_dec_IR_reg[9]/NET0131  & ~n4117 ;
  assign n5289 = ~\core_c_dec_IRE_reg[9]/NET0131  & n4117 ;
  assign n5290 = ~n5288 & ~n5289 ;
  assign n5291 = ~n4104 & ~n5290 ;
  assign n5292 = ~n5287 & ~n5291 ;
  assign n5293 = n4120 & n5292 ;
  assign n5313 = \bdma_BIAD_reg[5]/NET0131  & n5066 ;
  assign n5314 = \idma_DCTL_reg[5]/NET0131  & n5068 ;
  assign n5315 = ~n5313 & ~n5314 ;
  assign n5316 = n4099 & ~n5315 ;
  assign n5317 = ~n5293 & ~n5316 ;
  assign n5318 = ~n5312 & n5317 ;
  assign n5326 = ~n4392 & ~n5059 ;
  assign n5327 = ~\core_c_psq_EXA_reg[6]/P0001  & ~n5086 ;
  assign n5328 = ~n5087 & ~n5327 ;
  assign n5329 = n4835 & n5328 ;
  assign n5333 = n4764 & n4840 ;
  assign n5330 = ~\core_c_psq_IFA_reg[6]/P0001  & ~n5099 ;
  assign n5331 = ~n5100 & ~n5330 ;
  assign n5332 = n5050 & n5331 ;
  assign n5334 = \sice_IRR_reg[6]/P0001  & n4837 ;
  assign n5335 = ~n5332 & ~n5334 ;
  assign n5336 = ~n5333 & n5335 ;
  assign n5337 = ~n5329 & n5336 ;
  assign n5338 = ~n5326 & n5337 ;
  assign n5339 = n4128 & ~n5338 ;
  assign n5319 = ~\core_c_psq_IFA_reg[6]/P0001  & n4104 ;
  assign n5320 = ~\core_c_dec_IR_reg[10]/NET0131  & ~n4117 ;
  assign n5321 = ~\core_c_dec_IRE_reg[10]/NET0131  & n4117 ;
  assign n5322 = ~n5320 & ~n5321 ;
  assign n5323 = ~n4104 & ~n5322 ;
  assign n5324 = ~n5319 & ~n5323 ;
  assign n5325 = n4120 & n5324 ;
  assign n5340 = \bdma_BIAD_reg[6]/NET0131  & n5066 ;
  assign n5341 = \idma_DCTL_reg[6]/NET0131  & n5068 ;
  assign n5342 = ~n5340 & ~n5341 ;
  assign n5343 = n4099 & ~n5342 ;
  assign n5344 = ~n5325 & ~n5343 ;
  assign n5345 = ~n5339 & n5344 ;
  assign n5353 = ~n4656 & ~n5059 ;
  assign n5354 = ~\core_c_psq_EXA_reg[7]/P0001  & ~n5087 ;
  assign n5355 = ~n5088 & ~n5354 ;
  assign n5356 = n4835 & n5355 ;
  assign n5360 = n4783 & n4840 ;
  assign n5357 = ~\core_c_psq_IFA_reg[7]/P0001  & ~n5100 ;
  assign n5358 = ~n5101 & ~n5357 ;
  assign n5359 = n5050 & n5358 ;
  assign n5361 = \sice_IRR_reg[7]/P0001  & n4837 ;
  assign n5362 = ~n5359 & ~n5361 ;
  assign n5363 = ~n5360 & n5362 ;
  assign n5364 = ~n5356 & n5363 ;
  assign n5365 = ~n5353 & n5364 ;
  assign n5366 = n4128 & ~n5365 ;
  assign n5346 = ~\core_c_psq_IFA_reg[7]/P0001  & n4104 ;
  assign n5347 = ~\core_c_dec_IR_reg[11]/NET0131  & ~n4117 ;
  assign n5348 = ~\core_c_dec_IRE_reg[11]/NET0131  & n4117 ;
  assign n5349 = ~n5347 & ~n5348 ;
  assign n5350 = ~n4104 & ~n5349 ;
  assign n5351 = ~n5346 & ~n5350 ;
  assign n5352 = n4120 & n5351 ;
  assign n5367 = \bdma_BIAD_reg[7]/NET0131  & n5066 ;
  assign n5368 = \idma_DCTL_reg[7]/NET0131  & n5068 ;
  assign n5369 = ~n5367 & ~n5368 ;
  assign n5370 = n4099 & ~n5369 ;
  assign n5371 = ~n5352 & ~n5370 ;
  assign n5372 = ~n5366 & n5371 ;
  assign n5380 = ~n4425 & ~n5059 ;
  assign n5381 = ~\core_c_psq_EXA_reg[8]/P0001  & ~n5088 ;
  assign n5382 = ~n5089 & ~n5381 ;
  assign n5383 = n4835 & n5382 ;
  assign n5387 = n4735 & n4840 ;
  assign n5384 = ~\core_c_psq_IFA_reg[8]/P0001  & ~n5101 ;
  assign n5385 = ~n5102 & ~n5384 ;
  assign n5386 = n5050 & n5385 ;
  assign n5388 = \sice_IRR_reg[8]/P0001  & n4837 ;
  assign n5389 = ~n5386 & ~n5388 ;
  assign n5390 = ~n5387 & n5389 ;
  assign n5391 = ~n5383 & n5390 ;
  assign n5392 = ~n5380 & n5391 ;
  assign n5393 = n4128 & ~n5392 ;
  assign n5373 = ~\core_c_psq_IFA_reg[8]/P0001  & n4104 ;
  assign n5374 = ~\core_c_dec_IR_reg[12]/NET0131  & ~n4117 ;
  assign n5375 = ~\core_c_dec_IRE_reg[12]/NET0131  & n4117 ;
  assign n5376 = ~n5374 & ~n5375 ;
  assign n5377 = ~n4104 & ~n5376 ;
  assign n5378 = ~n5373 & ~n5377 ;
  assign n5379 = n4120 & n5378 ;
  assign n5394 = \bdma_BIAD_reg[8]/NET0131  & n5066 ;
  assign n5395 = \idma_DCTL_reg[8]/NET0131  & n5068 ;
  assign n5396 = ~n5394 & ~n5395 ;
  assign n5397 = n4099 & ~n5396 ;
  assign n5398 = ~n5379 & ~n5397 ;
  assign n5399 = ~n5393 & n5398 ;
  assign n5407 = ~n4554 & ~n5059 ;
  assign n5408 = ~\core_c_psq_EXA_reg[9]/P0001  & ~n5089 ;
  assign n5409 = ~n5090 & ~n5408 ;
  assign n5410 = n4835 & n5409 ;
  assign n5414 = n4739 & n4840 ;
  assign n5411 = ~\core_c_psq_IFA_reg[9]/P0001  & ~n5102 ;
  assign n5412 = ~n5103 & ~n5411 ;
  assign n5413 = n5050 & n5412 ;
  assign n5415 = \sice_IRR_reg[9]/P0001  & n4837 ;
  assign n5416 = ~n5413 & ~n5415 ;
  assign n5417 = ~n5414 & n5416 ;
  assign n5418 = ~n5410 & n5417 ;
  assign n5419 = ~n5407 & n5418 ;
  assign n5420 = n4128 & ~n5419 ;
  assign n5400 = ~\core_c_psq_IFA_reg[9]/P0001  & n4104 ;
  assign n5401 = ~\core_c_dec_IR_reg[13]/NET0131  & ~n4117 ;
  assign n5402 = ~\core_c_dec_IRE_reg[13]/NET0131  & n4117 ;
  assign n5403 = ~n5401 & ~n5402 ;
  assign n5404 = ~n4104 & ~n5403 ;
  assign n5405 = ~n5400 & ~n5404 ;
  assign n5406 = n4120 & n5405 ;
  assign n5421 = \bdma_BIAD_reg[9]/NET0131  & n5066 ;
  assign n5422 = \idma_DCTL_reg[9]/NET0131  & n5068 ;
  assign n5423 = ~n5421 & ~n5422 ;
  assign n5424 = n4099 & ~n5423 ;
  assign n5425 = ~n5406 & ~n5424 ;
  assign n5426 = ~n5420 & n5425 ;
  assign n5427 = ~\emc_ECS_reg[0]/NET0131  & ~\emc_ECS_reg[3]/NET0131  ;
  assign n5428 = \emc_ECS_reg[1]/NET0131  & \emc_ECS_reg[2]/NET0131  ;
  assign n5429 = n5427 & n5428 ;
  assign n5430 = \emc_ECS_reg[0]/NET0131  & ~\emc_ECS_reg[3]/NET0131  ;
  assign n5431 = ~\emc_ECS_reg[1]/NET0131  & \emc_ECS_reg[2]/NET0131  ;
  assign n5432 = n5430 & n5431 ;
  assign n5433 = ~\emc_ECS_reg[1]/NET0131  & ~\emc_ECS_reg[2]/NET0131  ;
  assign n5434 = n5430 & n5433 ;
  assign n5435 = \core_c_psq_DMOVL_reg_DO_reg[3]/NET0131  & ~\core_dag_ilm1reg_DMA_pi_DO_reg[13]/NET0131  ;
  assign n5436 = \core_c_dec_Double_E_reg/P0001  & n5435 ;
  assign n5437 = ~\emc_IOcst_reg/NET0131  & ~\emc_WSCRext_reg_DO_reg[1]/NET0131  ;
  assign n5438 = \emc_IOcst_reg/NET0131  & ~\emc_WSCRreg_DO_reg[3]/NET0131  ;
  assign n5439 = ~n5437 & ~n5438 ;
  assign n5440 = ~\emc_DMcst_reg/NET0131  & ~n5439 ;
  assign n5441 = \emc_DMcst_reg/NET0131  & ~\emc_WSCRreg_DO_reg[11]/NET0131  ;
  assign n5442 = ~n5440 & ~n5441 ;
  assign n5443 = ~\emc_PMcst_reg/NET0131  & ~n5442 ;
  assign n5444 = \emc_PMcst_reg/NET0131  & ~\emc_WSCRreg_DO_reg[7]/NET0131  ;
  assign n5445 = ~n5443 & ~n5444 ;
  assign n5498 = \emc_RWcnt_reg[3]/P0001  & ~n5445 ;
  assign n5486 = ~\emc_IOcst_reg/NET0131  & ~\memc_usysr_DO_reg[14]/NET0131  ;
  assign n5487 = \emc_IOcst_reg/NET0131  & ~\emc_WSCRreg_DO_reg[0]/NET0131  ;
  assign n5488 = ~n5486 & ~n5487 ;
  assign n5489 = ~\emc_DMcst_reg/NET0131  & ~n5488 ;
  assign n5490 = \emc_DMcst_reg/NET0131  & ~\emc_WSCRreg_DO_reg[8]/NET0131  ;
  assign n5491 = ~n5489 & ~n5490 ;
  assign n5492 = ~\emc_PMcst_reg/NET0131  & ~n5491 ;
  assign n5493 = \emc_PMcst_reg/NET0131  & ~\emc_WSCRreg_DO_reg[4]/NET0131  ;
  assign n5494 = ~n5492 & ~n5493 ;
  assign n5495 = ~\emc_RWcnt_reg[0]/P0001  & n5494 ;
  assign n5497 = \emc_RWcnt_reg[0]/P0001  & ~n5494 ;
  assign n5504 = ~n5495 & ~n5497 ;
  assign n5505 = ~n5498 & n5504 ;
  assign n5446 = ~\emc_RWcnt_reg[3]/P0001  & n5445 ;
  assign n5447 = \emc_PMcst_reg/NET0131  & ~\emc_WSCRext_reg_DO_reg[4]/NET0131  ;
  assign n5448 = ~\emc_DMcst_reg/NET0131  & \emc_IOcst_reg/NET0131  ;
  assign n5449 = \emc_WSCRext_reg_DO_reg[2]/NET0131  & n5448 ;
  assign n5450 = \emc_DMcst_reg/NET0131  & \emc_WSCRext_reg_DO_reg[6]/NET0131  ;
  assign n5451 = ~\emc_PMcst_reg/NET0131  & ~n5450 ;
  assign n5452 = ~n5449 & n5451 ;
  assign n5453 = ~n5447 & ~n5452 ;
  assign n5454 = ~\emc_RWcnt_reg[4]/P0001  & ~n5453 ;
  assign n5455 = \emc_RWcnt_reg[4]/P0001  & n5453 ;
  assign n5456 = ~n5454 & ~n5455 ;
  assign n5479 = \emc_PMcst_reg/NET0131  & ~\emc_WSCRext_reg_DO_reg[5]/NET0131  ;
  assign n5480 = \emc_WSCRext_reg_DO_reg[3]/NET0131  & n5448 ;
  assign n5481 = \emc_DMcst_reg/NET0131  & \emc_WSCRext_reg_DO_reg[7]/NET0131  ;
  assign n5482 = ~\emc_PMcst_reg/NET0131  & ~n5481 ;
  assign n5483 = ~n5480 & n5482 ;
  assign n5484 = ~n5479 & ~n5483 ;
  assign n5485 = ~\emc_RWcnt_reg[5]/P0001  & n5484 ;
  assign n5496 = \emc_RWcnt_reg[5]/P0001  & ~n5484 ;
  assign n5499 = ~n5485 & ~n5496 ;
  assign n5500 = ~n5456 & n5499 ;
  assign n5501 = ~n5446 & n5500 ;
  assign n5457 = ~\emc_IOcst_reg/NET0131  & ~\memc_usysr_DO_reg[15]/NET0131  ;
  assign n5458 = \emc_IOcst_reg/NET0131  & ~\emc_WSCRreg_DO_reg[1]/NET0131  ;
  assign n5459 = ~n5457 & ~n5458 ;
  assign n5460 = ~\emc_DMcst_reg/NET0131  & ~n5459 ;
  assign n5461 = \emc_DMcst_reg/NET0131  & ~\emc_WSCRreg_DO_reg[9]/NET0131  ;
  assign n5462 = ~n5460 & ~n5461 ;
  assign n5463 = ~\emc_PMcst_reg/NET0131  & ~n5462 ;
  assign n5464 = \emc_PMcst_reg/NET0131  & ~\emc_WSCRreg_DO_reg[5]/NET0131  ;
  assign n5465 = ~n5463 & ~n5464 ;
  assign n5466 = \emc_RWcnt_reg[1]/P0001  & ~n5465 ;
  assign n5467 = ~\emc_RWcnt_reg[1]/P0001  & n5465 ;
  assign n5502 = ~n5466 & ~n5467 ;
  assign n5468 = ~\emc_IOcst_reg/NET0131  & ~\emc_WSCRext_reg_DO_reg[0]/NET0131  ;
  assign n5469 = \emc_IOcst_reg/NET0131  & ~\emc_WSCRreg_DO_reg[2]/NET0131  ;
  assign n5470 = ~n5468 & ~n5469 ;
  assign n5471 = ~\emc_DMcst_reg/NET0131  & ~n5470 ;
  assign n5472 = \emc_DMcst_reg/NET0131  & ~\emc_WSCRreg_DO_reg[10]/NET0131  ;
  assign n5473 = ~n5471 & ~n5472 ;
  assign n5474 = ~\emc_PMcst_reg/NET0131  & ~n5473 ;
  assign n5475 = \emc_PMcst_reg/NET0131  & ~\emc_WSCRreg_DO_reg[6]/NET0131  ;
  assign n5476 = ~n5474 & ~n5475 ;
  assign n5477 = \emc_RWcnt_reg[2]/P0001  & ~n5476 ;
  assign n5478 = ~\emc_RWcnt_reg[2]/P0001  & n5476 ;
  assign n5503 = ~n5477 & ~n5478 ;
  assign n5506 = n5502 & n5503 ;
  assign n5507 = n5501 & n5506 ;
  assign n5508 = n5505 & n5507 ;
  assign n5509 = ~n5436 & n5508 ;
  assign n5510 = n5434 & ~n5509 ;
  assign n5522 = ~\emc_ECS_reg[0]/NET0131  & \emc_ECS_reg[3]/NET0131  ;
  assign n5523 = ~\emc_ECS_reg[2]/NET0131  & n5522 ;
  assign n5524 = n5508 & n5523 ;
  assign n5518 = \emc_ECS_reg[0]/NET0131  & \emc_ECS_reg[3]/NET0131  ;
  assign n5519 = n5433 & n5518 ;
  assign n5520 = ~n5432 & ~n5519 ;
  assign n5521 = ~n5508 & ~n5520 ;
  assign n5511 = ~\emc_DMcst_reg/NET0131  & ~\emc_IOcst_reg/NET0131  ;
  assign n5512 = ~\emc_PMcst_reg/NET0131  & n5511 ;
  assign n5513 = \core_c_psq_ECYC_reg/P0001  & ~\emc_eRDY_reg/NET0131  ;
  assign n5514 = ~n5512 & n5513 ;
  assign n5515 = ~\emc_ECS_reg[2]/NET0131  & ~n5514 ;
  assign n5516 = ~\emc_ECS_reg[1]/NET0131  & n5427 ;
  assign n5517 = ~n5515 & n5516 ;
  assign n5535 = \bdma_BCTL_reg[2]/NET0131  & ~\bdma_BCTL_reg[4]/NET0131  ;
  assign n5536 = ~\bdma_BCTL_reg[2]/NET0131  & ~\bdma_BCTL_reg[5]/NET0131  ;
  assign n5537 = ~n5535 & ~n5536 ;
  assign n5538 = ~\bdma_BWcnt_reg[1]/NET0131  & ~n5537 ;
  assign n5539 = \bdma_BWcnt_reg[1]/NET0131  & n5537 ;
  assign n5540 = ~n5538 & ~n5539 ;
  assign n5541 = \bdma_BCTL_reg[2]/NET0131  & ~\bdma_BCTL_reg[5]/NET0131  ;
  assign n5542 = ~\bdma_BCTL_reg[2]/NET0131  & ~\bdma_BCTL_reg[6]/NET0131  ;
  assign n5543 = ~n5541 & ~n5542 ;
  assign n5544 = \bdma_BWcnt_reg[2]/NET0131  & ~n5543 ;
  assign n5545 = ~\bdma_BWcnt_reg[2]/NET0131  & n5543 ;
  assign n5551 = ~n5544 & ~n5545 ;
  assign n5546 = \bdma_BCTL_reg[2]/NET0131  & ~\bdma_BCTL_reg[6]/NET0131  ;
  assign n5547 = ~\bdma_BCTL_reg[2]/NET0131  & ~\bdma_BCTL_reg[7]/NET0131  ;
  assign n5548 = ~n5546 & ~n5547 ;
  assign n5549 = \bdma_BWcnt_reg[3]/NET0131  & ~n5548 ;
  assign n5550 = ~\bdma_BWcnt_reg[3]/NET0131  & n5548 ;
  assign n5552 = ~n5549 & ~n5550 ;
  assign n5553 = n5551 & n5552 ;
  assign n5554 = ~n5540 & n5553 ;
  assign n5525 = ~\bdma_BCTL_reg[2]/NET0131  & ~\bdma_BCTL_reg[4]/NET0131  ;
  assign n5526 = \bdma_BWcnt_reg[0]/NET0131  & ~n5525 ;
  assign n5527 = ~\bdma_BWcnt_reg[0]/NET0131  & n5525 ;
  assign n5528 = ~n5526 & ~n5527 ;
  assign n5529 = \bdma_BCTL_reg[2]/NET0131  & ~\bdma_BCTL_reg[7]/NET0131  ;
  assign n5530 = \bdma_BWcnt_reg[4]/NET0131  & ~n5529 ;
  assign n5531 = ~\bdma_BWcnt_reg[4]/NET0131  & n5529 ;
  assign n5532 = ~n5530 & ~n5531 ;
  assign n5533 = ~n5528 & ~n5532 ;
  assign n5534 = n5431 & n5522 ;
  assign n5555 = n5533 & n5534 ;
  assign n5556 = n5554 & n5555 ;
  assign n5557 = ~n5517 & ~n5556 ;
  assign n5558 = ~n5521 & n5557 ;
  assign n5559 = ~n5524 & n5558 ;
  assign n5560 = ~n5510 & n5559 ;
  assign n5570 = ~\emc_PMcst_reg/NET0131  & ~\emc_eRDY_reg/NET0131  ;
  assign n5571 = n5427 & n5570 ;
  assign n5572 = n5433 & n5571 ;
  assign n5566 = ~\T_TMODE[1]_pad  & \bdma_BDMAmode_reg/NET0131  ;
  assign n5567 = ~\core_c_psq_ECYC_reg/P0001  & n5566 ;
  assign n5568 = \T_TMODE[1]_pad  & \core_c_psq_ECYC_reg/P0001  ;
  assign n5569 = ~n5567 & ~n5568 ;
  assign n5573 = n5511 & ~n5569 ;
  assign n5574 = n5572 & n5573 ;
  assign n5561 = n5431 & n5518 ;
  assign n5562 = \bdma_BSreq_reg/NET0131  & n5561 ;
  assign n5563 = n5428 & n5522 ;
  assign n5564 = ~\auctl_BSack_reg/NET0131  & n5563 ;
  assign n5565 = ~n5562 & ~n5564 ;
  assign n5577 = ~n5519 & ~n5523 ;
  assign n5575 = \T_TMODE[1]_pad  & \emc_ECS_reg[1]/NET0131  ;
  assign n5576 = n5427 & n5575 ;
  assign n5578 = ~n5534 & ~n5576 ;
  assign n5579 = n5577 & n5578 ;
  assign n5580 = n5565 & n5579 ;
  assign n5581 = ~n5574 & n5580 ;
  assign n5583 = ~n5434 & n5520 ;
  assign n5584 = n5508 & ~n5583 ;
  assign n5582 = \emc_ECS_reg[1]/NET0131  & n5523 ;
  assign n5585 = n5565 & ~n5582 ;
  assign n5586 = ~n5584 & n5585 ;
  assign n5587 = n5581 & n5586 ;
  assign n5589 = n5511 & ~n5567 ;
  assign n5588 = ~\core_c_psq_ECYC_reg/P0001  & ~n5511 ;
  assign n5590 = n5572 & ~n5588 ;
  assign n5591 = ~n5589 & n5590 ;
  assign n5592 = \emc_ECS_reg[1]/NET0131  & ~\emc_ECS_reg[2]/NET0131  ;
  assign n5593 = n5430 & n5592 ;
  assign n5594 = n5431 & ~n5518 ;
  assign n5595 = ~n5593 & ~n5594 ;
  assign n5596 = n5565 & n5595 ;
  assign n5597 = ~n5591 & n5596 ;
  assign n5598 = n5587 & ~n5597 ;
  assign n5599 = ~n5560 & n5598 ;
  assign n5600 = ~n5432 & ~n5599 ;
  assign n5601 = ~n5429 & n5600 ;
  assign n5610 = \emc_IOcst_reg/NET0131  & ~n5601 ;
  assign n5611 = \emc_WSCRreg_DO_reg[14]/NET0131  & n5610 ;
  assign n5602 = \emc_DMcst_reg/NET0131  & ~n5601 ;
  assign n5603 = \emc_WSCRreg_DO_reg[13]/NET0131  & n5602 ;
  assign n5604 = n5427 & n5592 ;
  assign n5605 = ~n5560 & n5597 ;
  assign n5606 = n5587 & n5605 ;
  assign n5607 = ~n5434 & ~n5606 ;
  assign n5608 = ~n5604 & n5607 ;
  assign n5609 = \emc_WSCRreg_DO_reg[12]/NET0131  & ~n5608 ;
  assign n5612 = ~n5603 & ~n5609 ;
  assign n5613 = ~n5611 & n5612 ;
  assign n5621 = ~n4694 & ~n5059 ;
  assign n5622 = \core_c_psq_EXA_reg[12]/P0001  & n5130 ;
  assign n5623 = ~\core_c_psq_EXA_reg[12]/P0001  & ~n5130 ;
  assign n5624 = ~n5622 & ~n5623 ;
  assign n5625 = n4835 & n5624 ;
  assign n5630 = n4790 & n4840 ;
  assign n5626 = \core_c_psq_IFA_reg[12]/P0001  & n5134 ;
  assign n5627 = ~\core_c_psq_IFA_reg[12]/P0001  & ~n5134 ;
  assign n5628 = ~n5626 & ~n5627 ;
  assign n5629 = n5050 & n5628 ;
  assign n5631 = \sice_IRR_reg[12]/P0001  & n4837 ;
  assign n5632 = ~n5629 & ~n5631 ;
  assign n5633 = ~n5630 & n5632 ;
  assign n5634 = ~n5625 & n5633 ;
  assign n5635 = ~n5621 & n5634 ;
  assign n5636 = n4128 & ~n5635 ;
  assign n5614 = ~\core_c_psq_IFA_reg[12]/P0001  & n4104 ;
  assign n5615 = ~\core_c_dec_IR_reg[16]/NET0131  & ~n4117 ;
  assign n5616 = ~\core_c_dec_IRE_reg[16]/NET0131  & n4117 ;
  assign n5617 = ~n5615 & ~n5616 ;
  assign n5618 = ~n4104 & ~n5617 ;
  assign n5619 = ~n5614 & ~n5618 ;
  assign n5620 = n4120 & n5619 ;
  assign n5637 = \bdma_BIAD_reg[12]/NET0131  & n5066 ;
  assign n5638 = \idma_DCTL_reg[12]/NET0131  & n5068 ;
  assign n5639 = ~n5637 & ~n5638 ;
  assign n5640 = n4099 & ~n5639 ;
  assign n5641 = ~n5620 & ~n5640 ;
  assign n5642 = ~n5636 & n5641 ;
  assign n5643 = PM_bdry_sel_pad & ~n5642 ;
  assign n5646 = ~n4489 & ~n5059 ;
  assign n5647 = ~\core_c_psq_EXA_reg[13]/P0001  & ~n5622 ;
  assign n5648 = \core_c_psq_EXA_reg[13]/P0001  & n5622 ;
  assign n5649 = ~n5647 & ~n5648 ;
  assign n5650 = n4835 & n5649 ;
  assign n5653 = ~\core_c_psq_IFA_reg[13]/P0001  & ~n5626 ;
  assign n5654 = \core_c_psq_IFA_reg[13]/P0001  & n5626 ;
  assign n5655 = ~n5653 & ~n5654 ;
  assign n5656 = n5050 & n5655 ;
  assign n5651 = n4786 & n4840 ;
  assign n5652 = \sice_IRR_reg[13]/P0001  & n4837 ;
  assign n5657 = ~n5651 & ~n5652 ;
  assign n5658 = ~n5656 & n5657 ;
  assign n5659 = ~n5650 & n5658 ;
  assign n5660 = ~n5646 & n5659 ;
  assign n5661 = n4128 & ~n5660 ;
  assign n5662 = ~\core_c_psq_IFA_reg[13]/P0001  & n4104 ;
  assign n5664 = \core_c_dec_IR_reg[17]/NET0131  & ~n4117 ;
  assign n5663 = \core_c_dec_IRE_reg[17]/NET0131  & n4117 ;
  assign n5665 = ~n4104 & ~n5663 ;
  assign n5666 = ~n5664 & n5665 ;
  assign n5667 = ~n5662 & ~n5666 ;
  assign n5668 = n4120 & n5667 ;
  assign n5644 = ~n4098 & n5066 ;
  assign n5645 = \bdma_BIAD_reg[13]/NET0131  & n5644 ;
  assign n5669 = \idma_DCTL_reg[13]/NET0131  & n5068 ;
  assign n5670 = n4099 & n5669 ;
  assign n5671 = ~n5645 & ~n5670 ;
  assign n5672 = ~n5668 & n5671 ;
  assign n5673 = ~n5661 & n5672 ;
  assign n5674 = ~n5643 & n5673 ;
  assign n5716 = ~\sice_GO_NX_reg/NET0131  & n4096 ;
  assign n5717 = n4064 & n5716 ;
  assign n5718 = ~n4065 & n5717 ;
  assign n5701 = \core_c_psq_MGNT_reg/NET0131  & \core_c_psq_PCS_reg[10]/NET0131  ;
  assign n5702 = \core_c_psq_PCS_reg[0]/NET0131  & n4105 ;
  assign n5703 = ~\core_c_psq_PCS2or3_reg/NET0131  & ~\core_c_psq_PCS_reg[13]/NET0131  ;
  assign n5704 = n4084 & ~n5703 ;
  assign n5705 = ~\core_c_psq_PCS_reg[1]/NET0131  & ~n5704 ;
  assign n5706 = ~n5702 & n5705 ;
  assign n5707 = \core_c_psq_MREQ_reg/NET0131  & ~n5706 ;
  assign n5708 = ~n5701 & ~n5707 ;
  assign n5685 = ~\core_c_psq_MGNT_reg/NET0131  & \core_c_psq_PCS_reg[10]/NET0131  ;
  assign n5686 = ~\core_c_psq_PCS2or3_reg/NET0131  & ~\core_c_psq_PCS_reg[11]/NET0131  ;
  assign n5687 = n4085 & ~n5686 ;
  assign n5688 = ~n5685 & ~n5687 ;
  assign n5689 = \core_c_dec_MACdep_Eg_reg/P0001  & ~n5688 ;
  assign n5690 = ~\auctl_STEAL_reg/NET0131  & \core_c_psq_PCS_reg[5]/NET0131  ;
  assign n5691 = ~\memc_STI_Cg_reg/NET0131  & n5690 ;
  assign n5692 = ~\core_c_psq_PCS_reg[11]/NET0131  & ~n5691 ;
  assign n5693 = \core_c_psq_PCS2or3_reg/NET0131  & \memc_LDaST_Eg_reg/NET0131  ;
  assign n5694 = n4085 & n5693 ;
  assign n5695 = n5692 & ~n5694 ;
  assign n5696 = ~n5689 & n5695 ;
  assign n5697 = \core_c_psq_PCS_reg[1]/NET0131  & ~\emc_eRDY_reg/NET0131  ;
  assign n5698 = \core_c_psq_PCS_reg[10]/NET0131  & ~n4068 ;
  assign n5699 = n4105 & n5698 ;
  assign n5700 = ~n5697 & ~n5699 ;
  assign n5709 = ~\core_c_psq_PCS_reg[7]/NET0131  & ~\core_c_psq_PCS_reg[8]/NET0131  ;
  assign n5710 = ~n4079 & n5709 ;
  assign n5711 = ~n4087 & n5710 ;
  assign n5712 = ~n4068 & ~n5711 ;
  assign n5713 = n5700 & ~n5712 ;
  assign n5714 = n5696 & n5713 ;
  assign n5715 = n5708 & n5714 ;
  assign n5675 = \core_c_psq_PCS_reg[6]/NET0131  & ~n4075 ;
  assign n5676 = ~\core_c_psq_PCS_reg[2]/NET0131  & ~n4107 ;
  assign n5677 = \core_c_dec_IDLE_Eg_reg/P0001  & n4082 ;
  assign n5678 = ~n5676 & n5677 ;
  assign n5679 = ~n5675 & ~n5678 ;
  assign n5719 = n4116 & n5679 ;
  assign n5720 = n5715 & n5719 ;
  assign n5721 = n5718 & n5720 ;
  assign n5681 = \clkc_Cnt4096_s1_reg/NET0131  & \clkc_Cnt4096_s2_reg/NET0131  ;
  assign n5682 = n4115 & ~n5681 ;
  assign n5683 = ~n5068 & n5682 ;
  assign n5684 = ~n5066 & n5683 ;
  assign n5680 = n4104 & ~n5679 ;
  assign n5722 = ~\T_TMODE[1]_pad  & ~n5680 ;
  assign n5723 = ~n5684 & n5722 ;
  assign n5724 = ~n5721 & n5723 ;
  assign n5725 = n5674 & n5724 ;
  assign n5728 = \bdma_BDMAmode_reg/NET0131  & \bdma_BM_cyc_reg/P0001  ;
  assign n5729 = ~\bdma_BCTL_reg[0]/NET0131  & ~\bdma_BCTL_reg[1]/NET0131  ;
  assign n5730 = n5728 & n5729 ;
  assign n5726 = ~PM_bdry_sel_pad & ~\bdma_BIAD_reg[12]/NET0131  ;
  assign n5727 = \bdma_BIAD_reg[13]/NET0131  & ~n5726 ;
  assign n5731 = ~\bdma_CMcnt_reg[0]/NET0131  & \bdma_CMcnt_reg[1]/NET0131  ;
  assign n5732 = ~n5727 & n5731 ;
  assign n5733 = n5730 & n5732 ;
  assign n5734 = ~\bdma_BCTL_reg[2]/NET0131  & n5733 ;
  assign n5735 = n5066 & n5734 ;
  assign n5736 = \sice_idr0_reg_DO_reg[0]/P0001  & ~n5735 ;
  assign n5737 = \bdma_BRdataBUF_reg[0]/P0001  & n5735 ;
  assign n5738 = ~n5736 & ~n5737 ;
  assign n5739 = ~n5068 & ~n5738 ;
  assign n5740 = \idma_DTMP_L_reg[0]/P0001  & n5068 ;
  assign n5741 = ~n5739 & ~n5740 ;
  assign n5742 = \sice_idr0_reg_DO_reg[10]/P0001  & ~n5735 ;
  assign n5743 = \bdma_BRdataBUF_reg[10]/P0001  & n5735 ;
  assign n5744 = ~n5742 & ~n5743 ;
  assign n5745 = ~n5068 & ~n5744 ;
  assign n5746 = \idma_DTMP_H_reg[2]/P0001  & n5068 ;
  assign n5747 = ~n5745 & ~n5746 ;
  assign n5748 = \sice_idr0_reg_DO_reg[11]/P0001  & ~n5735 ;
  assign n5749 = \bdma_BRdataBUF_reg[11]/P0001  & n5735 ;
  assign n5750 = ~n5748 & ~n5749 ;
  assign n5751 = ~n5068 & ~n5750 ;
  assign n5752 = \idma_DTMP_H_reg[3]/P0001  & n5068 ;
  assign n5753 = ~n5751 & ~n5752 ;
  assign n5754 = \sice_idr1_reg_DO_reg[0]/P0001  & ~n5735 ;
  assign n5755 = \bdma_BRdataBUF_reg[12]/P0001  & n5735 ;
  assign n5756 = ~n5754 & ~n5755 ;
  assign n5757 = ~n5068 & ~n5756 ;
  assign n5758 = \idma_DTMP_H_reg[4]/P0001  & n5068 ;
  assign n5759 = ~n5757 & ~n5758 ;
  assign n5760 = \sice_idr1_reg_DO_reg[1]/P0001  & ~n5735 ;
  assign n5761 = \bdma_BRdataBUF_reg[13]/P0001  & n5735 ;
  assign n5762 = ~n5760 & ~n5761 ;
  assign n5763 = ~n5068 & ~n5762 ;
  assign n5764 = \idma_DTMP_H_reg[5]/P0001  & n5068 ;
  assign n5765 = ~n5763 & ~n5764 ;
  assign n5766 = \sice_idr1_reg_DO_reg[2]/P0001  & ~n5735 ;
  assign n5767 = \bdma_BRdataBUF_reg[14]/P0001  & n5735 ;
  assign n5768 = ~n5766 & ~n5767 ;
  assign n5769 = ~n5068 & ~n5768 ;
  assign n5770 = \idma_DTMP_H_reg[6]/P0001  & n5068 ;
  assign n5771 = ~n5769 & ~n5770 ;
  assign n5772 = \sice_idr1_reg_DO_reg[3]/P0001  & ~n5735 ;
  assign n5773 = \bdma_BRdataBUF_reg[15]/P0001  & n5735 ;
  assign n5774 = ~n5772 & ~n5773 ;
  assign n5775 = ~n5068 & ~n5774 ;
  assign n5776 = \idma_DTMP_H_reg[7]/P0001  & n5068 ;
  assign n5777 = ~n5775 & ~n5776 ;
  assign n5778 = \sice_idr1_reg_DO_reg[4]/P0001  & ~n5735 ;
  assign n5779 = \bdma_BRdataBUF_reg[16]/P0001  & n5735 ;
  assign n5780 = ~n5778 & ~n5779 ;
  assign n5781 = ~n5068 & ~n5780 ;
  assign n5782 = \idma_DTMP_H_reg[8]/P0001  & n5068 ;
  assign n5783 = ~n5781 & ~n5782 ;
  assign n5784 = \sice_idr1_reg_DO_reg[5]/P0001  & ~n5735 ;
  assign n5785 = \bdma_BRdataBUF_reg[17]/P0001  & n5735 ;
  assign n5786 = ~n5784 & ~n5785 ;
  assign n5787 = ~n5068 & ~n5786 ;
  assign n5788 = \idma_DTMP_H_reg[9]/P0001  & n5068 ;
  assign n5789 = ~n5787 & ~n5788 ;
  assign n5790 = \sice_idr1_reg_DO_reg[6]/P0001  & ~n5735 ;
  assign n5791 = \bdma_BRdataBUF_reg[18]/P0001  & n5735 ;
  assign n5792 = ~n5790 & ~n5791 ;
  assign n5793 = ~n5068 & ~n5792 ;
  assign n5794 = \idma_DTMP_H_reg[10]/P0001  & n5068 ;
  assign n5795 = ~n5793 & ~n5794 ;
  assign n5796 = \sice_idr1_reg_DO_reg[7]/P0001  & ~n5735 ;
  assign n5797 = \bdma_BRdataBUF_reg[19]/P0001  & n5735 ;
  assign n5798 = ~n5796 & ~n5797 ;
  assign n5799 = ~n5068 & ~n5798 ;
  assign n5800 = \idma_DTMP_H_reg[11]/P0001  & n5068 ;
  assign n5801 = ~n5799 & ~n5800 ;
  assign n5802 = \sice_idr0_reg_DO_reg[1]/P0001  & ~n5735 ;
  assign n5803 = \bdma_BRdataBUF_reg[1]/P0001  & n5735 ;
  assign n5804 = ~n5802 & ~n5803 ;
  assign n5805 = ~n5068 & ~n5804 ;
  assign n5806 = \idma_DTMP_L_reg[1]/P0001  & n5068 ;
  assign n5807 = ~n5805 & ~n5806 ;
  assign n5808 = \sice_idr1_reg_DO_reg[8]/P0001  & ~n5735 ;
  assign n5809 = \bdma_BRdataBUF_reg[20]/P0001  & n5735 ;
  assign n5810 = ~n5808 & ~n5809 ;
  assign n5811 = ~n5068 & ~n5810 ;
  assign n5812 = \idma_DTMP_H_reg[12]/P0001  & n5068 ;
  assign n5813 = ~n5811 & ~n5812 ;
  assign n5814 = \sice_idr1_reg_DO_reg[9]/P0001  & ~n5735 ;
  assign n5815 = \bdma_BRdataBUF_reg[21]/P0001  & n5735 ;
  assign n5816 = ~n5814 & ~n5815 ;
  assign n5817 = ~n5068 & ~n5816 ;
  assign n5818 = \idma_DTMP_H_reg[13]/P0001  & n5068 ;
  assign n5819 = ~n5817 & ~n5818 ;
  assign n5820 = \sice_idr1_reg_DO_reg[10]/P0001  & ~n5735 ;
  assign n5821 = \bdma_BRdataBUF_reg[22]/P0001  & n5735 ;
  assign n5822 = ~n5820 & ~n5821 ;
  assign n5823 = ~n5068 & ~n5822 ;
  assign n5824 = \idma_DTMP_H_reg[14]/P0001  & n5068 ;
  assign n5825 = ~n5823 & ~n5824 ;
  assign n5826 = \sice_idr1_reg_DO_reg[11]/P0001  & ~n5735 ;
  assign n5827 = \bdma_BRdataBUF_reg[23]/P0001  & n5735 ;
  assign n5828 = ~n5826 & ~n5827 ;
  assign n5829 = ~n5068 & ~n5828 ;
  assign n5830 = \idma_DTMP_H_reg[15]/P0001  & n5068 ;
  assign n5831 = ~n5829 & ~n5830 ;
  assign n5832 = \sice_idr0_reg_DO_reg[2]/P0001  & ~n5735 ;
  assign n5833 = \bdma_BRdataBUF_reg[2]/P0001  & n5735 ;
  assign n5834 = ~n5832 & ~n5833 ;
  assign n5835 = ~n5068 & ~n5834 ;
  assign n5836 = \idma_DTMP_L_reg[2]/P0001  & n5068 ;
  assign n5837 = ~n5835 & ~n5836 ;
  assign n5838 = \sice_idr0_reg_DO_reg[3]/P0001  & ~n5735 ;
  assign n5839 = \bdma_BRdataBUF_reg[3]/P0001  & n5735 ;
  assign n5840 = ~n5838 & ~n5839 ;
  assign n5841 = ~n5068 & ~n5840 ;
  assign n5842 = \idma_DTMP_L_reg[3]/P0001  & n5068 ;
  assign n5843 = ~n5841 & ~n5842 ;
  assign n5844 = \sice_idr0_reg_DO_reg[4]/P0001  & ~n5735 ;
  assign n5845 = \bdma_BRdataBUF_reg[4]/P0001  & n5735 ;
  assign n5846 = ~n5844 & ~n5845 ;
  assign n5847 = ~n5068 & ~n5846 ;
  assign n5848 = \idma_DTMP_L_reg[4]/P0001  & n5068 ;
  assign n5849 = ~n5847 & ~n5848 ;
  assign n5850 = \sice_idr0_reg_DO_reg[5]/P0001  & ~n5735 ;
  assign n5851 = \bdma_BRdataBUF_reg[5]/P0001  & n5735 ;
  assign n5852 = ~n5850 & ~n5851 ;
  assign n5853 = ~n5068 & ~n5852 ;
  assign n5854 = \idma_DTMP_L_reg[5]/P0001  & n5068 ;
  assign n5855 = ~n5853 & ~n5854 ;
  assign n5856 = \sice_idr0_reg_DO_reg[6]/P0001  & ~n5735 ;
  assign n5857 = \bdma_BRdataBUF_reg[6]/P0001  & n5735 ;
  assign n5858 = ~n5856 & ~n5857 ;
  assign n5859 = ~n5068 & ~n5858 ;
  assign n5860 = \idma_DTMP_L_reg[6]/P0001  & n5068 ;
  assign n5861 = ~n5859 & ~n5860 ;
  assign n5862 = \sice_idr0_reg_DO_reg[7]/P0001  & ~n5735 ;
  assign n5863 = \bdma_BRdataBUF_reg[7]/P0001  & n5735 ;
  assign n5864 = ~n5862 & ~n5863 ;
  assign n5865 = ~n5068 & ~n5864 ;
  assign n5866 = \idma_DTMP_L_reg[7]/P0001  & n5068 ;
  assign n5867 = ~n5865 & ~n5866 ;
  assign n5868 = \sice_idr0_reg_DO_reg[8]/P0001  & ~n5735 ;
  assign n5869 = \bdma_BRdataBUF_reg[8]/P0001  & n5735 ;
  assign n5870 = ~n5868 & ~n5869 ;
  assign n5871 = ~n5068 & ~n5870 ;
  assign n5872 = \idma_DTMP_H_reg[0]/P0001  & n5068 ;
  assign n5873 = ~n5871 & ~n5872 ;
  assign n5874 = \sice_idr0_reg_DO_reg[9]/P0001  & ~n5735 ;
  assign n5875 = \bdma_BRdataBUF_reg[9]/P0001  & n5735 ;
  assign n5876 = ~n5874 & ~n5875 ;
  assign n5877 = ~n5068 & ~n5876 ;
  assign n5878 = \idma_DTMP_H_reg[1]/P0001  & n5068 ;
  assign n5879 = ~n5877 & ~n5878 ;
  assign n5880 = ~\idma_DCTL_reg[14]/NET0131  & n5068 ;
  assign n5881 = ~PM_bdry_sel_pad & ~\idma_DCTL_reg[12]/NET0131  ;
  assign n5882 = \idma_DCTL_reg[13]/NET0131  & ~n5881 ;
  assign n5883 = \idma_WRcyc_reg/NET0131  & ~n5882 ;
  assign n5884 = n5880 & n5883 ;
  assign n5885 = ~n5735 & ~n5884 ;
  assign n5886 = n5679 & ~n5885 ;
  assign n5887 = ~n5718 & n5886 ;
  assign n5888 = n4103 & ~n4117 ;
  assign n5889 = \core_c_dec_IR_reg[20]/NET0131  & ~n5679 ;
  assign n5890 = n5888 & n5889 ;
  assign n5891 = ~n5887 & ~n5890 ;
  assign n5892 = ~PM_bdry_sel_pad & n5642 ;
  assign n5893 = ~n5673 & ~n5892 ;
  assign n5895 = n5068 & ~n5718 ;
  assign n5899 = \idma_DOVL_reg[3]/NET0131  & n5895 ;
  assign n5894 = ~\core_c_psq_PMOVL_regl_DO_reg[3]/NET0131  & ~n5066 ;
  assign n5896 = ~\bdma_BOVL_reg[3]/NET0131  & n5066 ;
  assign n5897 = ~n5894 & ~n5896 ;
  assign n5898 = ~n5895 & n5897 ;
  assign n5900 = n5724 & ~n5898 ;
  assign n5901 = ~n5899 & n5900 ;
  assign n5902 = ~n5674 & n5901 ;
  assign n5903 = ~n5893 & n5902 ;
  assign n5904 = \core_c_psq_PMOVL_regl_DO_reg[2]/NET0131  & ~n5066 ;
  assign n5905 = \bdma_BOVL_reg[2]/NET0131  & n5066 ;
  assign n5906 = ~n5904 & ~n5905 ;
  assign n5907 = ~n5895 & ~n5906 ;
  assign n5908 = \idma_DOVL_reg[2]/NET0131  & n5895 ;
  assign n5909 = ~n5907 & ~n5908 ;
  assign n5910 = n5903 & n5909 ;
  assign n5911 = \core_c_psq_PMOVL_regl_DO_reg[1]/NET0131  & ~n5066 ;
  assign n5912 = \bdma_BOVL_reg[1]/NET0131  & n5066 ;
  assign n5913 = ~n5911 & ~n5912 ;
  assign n5914 = ~n5895 & ~n5913 ;
  assign n5915 = \idma_DOVL_reg[1]/NET0131  & n5895 ;
  assign n5916 = ~n5914 & ~n5915 ;
  assign n5917 = n5910 & n5916 ;
  assign n5918 = \core_c_psq_PMOVL_regl_DO_reg[0]/NET0131  & ~n5066 ;
  assign n5919 = \bdma_BOVL_reg[0]/NET0131  & n5066 ;
  assign n5920 = ~n5918 & ~n5919 ;
  assign n5921 = ~n5895 & ~n5920 ;
  assign n5922 = \idma_DOVL_reg[0]/NET0131  & n5895 ;
  assign n5923 = ~n5921 & ~n5922 ;
  assign n5924 = n5917 & n5923 ;
  assign n5925 = n5917 & ~n5923 ;
  assign n5926 = n5910 & ~n5916 ;
  assign n5927 = n5923 & n5926 ;
  assign n5928 = ~n5923 & n5926 ;
  assign n5929 = n5903 & ~n5909 ;
  assign n5930 = n5916 & n5929 ;
  assign n5931 = n5923 & n5930 ;
  assign n5932 = ~n5923 & n5930 ;
  assign n5933 = ~n5916 & n5929 ;
  assign n5934 = n5923 & n5933 ;
  assign n5935 = ~n5923 & n5933 ;
  assign n5936 = ~n4055 & ~n5716 ;
  assign n6022 = \core_c_dec_IR_reg[21]/NET0131  & ~\core_c_dec_IR_reg[22]/NET0131  ;
  assign n6023 = \core_c_dec_IR_reg[23]/NET0131  & n6022 ;
  assign n6107 = \core_c_dec_IR_reg[22]/NET0131  & \core_c_dec_IR_reg[23]/NET0131  ;
  assign n6108 = n4101 & ~n4102 ;
  assign n6109 = ~n6107 & ~n6108 ;
  assign n6110 = ~\core_c_dec_IR_reg[20]/NET0131  & ~n6109 ;
  assign n6111 = ~n6023 & ~n6110 ;
  assign n5950 = ~\sice_GO_NX_reg/NET0131  & n4093 ;
  assign n5951 = ~\core_c_dec_Dummy_E_reg/NET0131  & ~n5950 ;
  assign n5952 = ~\core_c_dec_Dummy_E_reg/NET0131  & ~\core_dag_ilm2reg_IL_E_reg[0]/P0001  ;
  assign n5953 = ~\auctl_R0Sack_reg/NET0131  & ~\auctl_R1Sack_reg/NET0131  ;
  assign n5954 = ~\auctl_T0Sack_reg/NET0131  & ~\auctl_T1Sack_reg/NET0131  ;
  assign n5955 = n5953 & n5954 ;
  assign n5956 = \core_c_dec_Post2_E_reg/P0001  & n5955 ;
  assign n5957 = ~\core_dag_ilm2reg_IL_E_reg[1]/P0001  & n5956 ;
  assign n5958 = n5952 & n5957 ;
  assign n5959 = ~\core_c_dec_MTIreg_E_reg[4]/P0001  & ~n5958 ;
  assign n5960 = n5951 & ~n5959 ;
  assign n5961 = ~\core_dag_ilm1reg_STEALI_E_reg[0]/P0001  & \core_dag_ilm1reg_STEALI_E_reg[2]/P0001  ;
  assign n5962 = ~\core_dag_ilm1reg_STEALI_E_reg[1]/P0001  & ~n5955 ;
  assign n5963 = n5961 & n5962 ;
  assign n5964 = ~n5960 & ~n5963 ;
  assign n5966 = n4049 & n4054 ;
  assign n5967 = \sport1_regs_AUTOreg_DO_reg[5]/NET0131  & n5966 ;
  assign n5968 = n4052 & n4053 ;
  assign n5969 = \sport1_regs_AUTOreg_DO_reg[10]/NET0131  & n5968 ;
  assign n5965 = \sport0_regs_AUTOreg_DO_reg[10]/NET0131  & n4050 ;
  assign n5970 = ~n4050 & n4051 ;
  assign n5971 = \sport0_regs_AUTOreg_DO_reg[5]/NET0131  & n5970 ;
  assign n5972 = ~n5965 & ~n5971 ;
  assign n5973 = ~n5969 & n5972 ;
  assign n5974 = ~n5967 & n5973 ;
  assign n5976 = \sport1_regs_AUTOreg_DO_reg[6]/NET0131  & n5966 ;
  assign n5977 = \sport1_regs_AUTOreg_DO_reg[11]/NET0131  & n5968 ;
  assign n5975 = \sport0_regs_AUTOreg_DO_reg[11]/NET0131  & n4050 ;
  assign n5978 = \sport0_regs_AUTOreg_DO_reg[6]/NET0131  & n5970 ;
  assign n5979 = ~n5975 & ~n5978 ;
  assign n5980 = ~n5977 & n5979 ;
  assign n5981 = ~n5976 & n5980 ;
  assign n5982 = n5974 & ~n5981 ;
  assign n5984 = \sport1_regs_AUTOreg_DO_reg[4]/NET0131  & n5966 ;
  assign n5985 = \sport1_regs_AUTOreg_DO_reg[9]/NET0131  & n5968 ;
  assign n5983 = \sport0_regs_AUTOreg_DO_reg[9]/NET0131  & n4050 ;
  assign n5986 = \sport0_regs_AUTOreg_DO_reg[4]/NET0131  & n5970 ;
  assign n5987 = ~n5983 & ~n5986 ;
  assign n5988 = ~n5985 & n5987 ;
  assign n5989 = ~n5984 & n5988 ;
  assign n5990 = n5982 & n5989 ;
  assign n5991 = ~n5964 & n5990 ;
  assign n5992 = \core_dag_ilm2reg_IL_E_reg[1]/P0001  & n5956 ;
  assign n5993 = ~\core_c_dec_Dummy_E_reg/NET0131  & \core_dag_ilm2reg_IL_E_reg[0]/P0001  ;
  assign n5994 = n5992 & n5993 ;
  assign n5995 = ~\core_c_dec_MTIreg_E_reg[7]/P0001  & ~n5994 ;
  assign n5996 = n5951 & ~n5995 ;
  assign n5997 = \core_dag_ilm1reg_STEALI_E_reg[1]/P0001  & ~n5955 ;
  assign n5998 = \core_dag_ilm1reg_STEALI_E_reg[0]/P0001  & \core_dag_ilm1reg_STEALI_E_reg[2]/P0001  ;
  assign n5999 = n5997 & n5998 ;
  assign n6000 = ~n5996 & ~n5999 ;
  assign n6001 = ~n5974 & ~n5981 ;
  assign n6002 = ~n5989 & n6001 ;
  assign n6003 = ~n6000 & n6002 ;
  assign n6018 = ~n5991 & ~n6003 ;
  assign n6004 = n5952 & n5992 ;
  assign n6005 = ~\core_c_dec_MTIreg_E_reg[6]/P0001  & ~n6004 ;
  assign n6006 = n5951 & ~n6005 ;
  assign n6007 = n5961 & n5997 ;
  assign n6008 = ~n6006 & ~n6007 ;
  assign n6009 = n5989 & n6001 ;
  assign n6010 = ~n6008 & n6009 ;
  assign n6011 = n5957 & n5993 ;
  assign n6012 = ~\core_c_dec_MTIreg_E_reg[5]/P0001  & ~n6011 ;
  assign n6013 = n5951 & ~n6012 ;
  assign n6014 = n5962 & n5998 ;
  assign n6015 = ~n6013 & ~n6014 ;
  assign n6016 = n5982 & ~n5989 ;
  assign n6017 = ~n6015 & n6016 ;
  assign n6019 = ~n6010 & ~n6017 ;
  assign n6020 = n6018 & n6019 ;
  assign n6021 = ~n4055 & n6020 ;
  assign n6024 = ~\core_c_dec_IR_reg[16]/NET0131  & ~\core_c_dec_IR_reg[17]/NET0131  ;
  assign n6025 = \core_c_dec_IR_reg[18]/NET0131  & \core_c_dec_IR_reg[19]/NET0131  ;
  assign n6026 = ~\core_c_dec_IR_reg[20]/NET0131  & ~\core_c_dec_IR_reg[23]/NET0131  ;
  assign n6027 = n4100 & n6026 ;
  assign n6028 = n6025 & n6027 ;
  assign n6029 = n6024 & n6028 ;
  assign n6030 = ~n6023 & ~n6029 ;
  assign n6031 = \core_c_dec_IR_reg[7]/NET0131  & ~n6030 ;
  assign n6032 = \core_c_dec_IR_reg[3]/NET0131  & n6030 ;
  assign n6033 = ~n6031 & ~n6032 ;
  assign n6034 = \core_c_dec_IR_reg[6]/NET0131  & ~n6030 ;
  assign n6035 = \core_c_dec_IR_reg[2]/NET0131  & n6030 ;
  assign n6036 = ~n6034 & ~n6035 ;
  assign n6037 = n6033 & n6036 ;
  assign n6038 = ~n5964 & n6037 ;
  assign n6039 = ~n6033 & ~n6036 ;
  assign n6040 = ~n6000 & n6039 ;
  assign n6045 = ~n6038 & ~n6040 ;
  assign n6041 = ~n6033 & n6036 ;
  assign n6042 = ~n6008 & n6041 ;
  assign n6043 = n6033 & ~n6036 ;
  assign n6044 = ~n6015 & n6043 ;
  assign n6046 = ~n6042 & ~n6044 ;
  assign n6047 = n6045 & n6046 ;
  assign n6048 = n4055 & n6047 ;
  assign n6049 = ~n6021 & ~n6048 ;
  assign n6114 = \core_c_dec_IR_reg[20]/NET0131  & ~n6109 ;
  assign n6115 = \core_c_dec_IR_reg[16]/NET0131  & ~\core_c_dec_IR_reg[17]/NET0131  ;
  assign n6116 = ~\core_c_dec_IR_reg[18]/NET0131  & ~\core_c_dec_IR_reg[19]/NET0131  ;
  assign n6117 = \core_c_dec_IR_reg[20]/NET0131  & ~\core_c_dec_IR_reg[23]/NET0131  ;
  assign n6118 = n4100 & n6117 ;
  assign n6119 = n6116 & n6118 ;
  assign n6120 = n6115 & n6119 ;
  assign n6121 = ~n6114 & ~n6120 ;
  assign n6122 = n6049 & ~n6121 ;
  assign n6123 = n6111 & ~n6122 ;
  assign n5940 = \core_dag_ilm1reg_DMA_pi_DO_reg[7]/NET0131  & \core_dag_ilm1reg_DMA_pi_DO_reg[8]/NET0131  ;
  assign n5941 = \core_dag_ilm1reg_DMA_pi_DO_reg[9]/NET0131  & n5940 ;
  assign n5937 = \core_dag_ilm1reg_DMA_pi_DO_reg[10]/NET0131  & \core_dag_ilm1reg_DMA_pi_DO_reg[11]/NET0131  ;
  assign n5938 = \core_dag_ilm1reg_DMA_pi_DO_reg[12]/NET0131  & \core_dag_ilm1reg_DMA_pi_DO_reg[13]/NET0131  ;
  assign n5939 = \core_dag_ilm1reg_DMA_pi_DO_reg[5]/NET0131  & \core_dag_ilm1reg_DMA_pi_DO_reg[6]/NET0131  ;
  assign n5942 = n5938 & n5939 ;
  assign n5943 = n5937 & n5942 ;
  assign n5944 = n5941 & n5943 ;
  assign n5945 = \memc_Dwrite_E_reg/NET0131  & ~\memc_EXTC_E_reg/NET0131  ;
  assign n5946 = ~n5944 & n5945 ;
  assign n5947 = ~\core_c_dec_Dummy_E_reg/NET0131  & n5946 ;
  assign n5948 = ~n4099 & ~n5947 ;
  assign n5949 = ~n4117 & n5948 ;
  assign n6050 = ~\core_dag_ilm1reg_STEALI_E_reg[0]/P0001  & ~\core_dag_ilm1reg_STEALI_E_reg[2]/P0001  ;
  assign n6051 = n5962 & n6050 ;
  assign n6052 = ~\core_c_dec_Dummy_E_reg/NET0131  & \core_c_dec_Post1_E_reg/P0001  ;
  assign n6053 = n5955 & n6052 ;
  assign n6054 = ~\core_c_dec_IRE_reg[3]/NET0131  & n6053 ;
  assign n6055 = ~\core_c_dec_IRE_reg[2]/NET0131  & n6054 ;
  assign n6056 = ~\core_c_dec_MTIreg_E_reg[0]/P0001  & ~n6055 ;
  assign n6057 = n5951 & ~n6056 ;
  assign n6058 = ~n6051 & ~n6057 ;
  assign n6059 = n5974 & n5981 ;
  assign n6060 = n5989 & n6059 ;
  assign n6061 = ~n6058 & n6060 ;
  assign n6087 = ~n4055 & ~n6061 ;
  assign n6079 = n5997 & n6050 ;
  assign n6080 = ~\core_c_dec_IRE_reg[2]/NET0131  & \core_c_dec_IRE_reg[3]/NET0131  ;
  assign n6081 = n6053 & n6080 ;
  assign n6082 = ~\core_c_dec_MTIreg_E_reg[2]/P0001  & ~n6081 ;
  assign n6083 = n5951 & ~n6082 ;
  assign n6084 = ~n6079 & ~n6083 ;
  assign n6076 = ~n5974 & n5981 ;
  assign n6085 = n5989 & n6076 ;
  assign n6086 = ~n6084 & n6085 ;
  assign n6062 = \core_dag_ilm1reg_STEALI_E_reg[0]/P0001  & ~\core_dag_ilm1reg_STEALI_E_reg[2]/P0001  ;
  assign n6063 = n5962 & n6062 ;
  assign n6064 = \core_c_dec_IRE_reg[2]/NET0131  & n6054 ;
  assign n6065 = ~\core_c_dec_MTIreg_E_reg[1]/P0001  & ~n6064 ;
  assign n6066 = n5951 & ~n6065 ;
  assign n6067 = ~n6063 & ~n6066 ;
  assign n6068 = ~n5989 & n6059 ;
  assign n6069 = ~n6067 & n6068 ;
  assign n6070 = n5997 & n6062 ;
  assign n6071 = \core_c_dec_IRE_reg[2]/NET0131  & \core_c_dec_IRE_reg[3]/NET0131  ;
  assign n6072 = n6053 & n6071 ;
  assign n6073 = ~\core_c_dec_MTIreg_E_reg[3]/P0001  & ~n6072 ;
  assign n6074 = n5951 & ~n6073 ;
  assign n6075 = ~n6070 & ~n6074 ;
  assign n6077 = ~n5989 & n6076 ;
  assign n6078 = ~n6075 & n6077 ;
  assign n6088 = ~n6069 & ~n6078 ;
  assign n6089 = ~n6086 & n6088 ;
  assign n6090 = n6087 & n6089 ;
  assign n6091 = \core_c_dec_IR_reg[2]/NET0131  & ~\core_c_dec_IR_reg[3]/NET0131  ;
  assign n6092 = ~n6067 & n6091 ;
  assign n6093 = ~\core_c_dec_IR_reg[2]/NET0131  & ~\core_c_dec_IR_reg[3]/NET0131  ;
  assign n6094 = ~n6058 & n6093 ;
  assign n6099 = ~n6092 & ~n6094 ;
  assign n6095 = ~\core_c_dec_IR_reg[2]/NET0131  & \core_c_dec_IR_reg[3]/NET0131  ;
  assign n6096 = ~n6084 & n6095 ;
  assign n6097 = \core_c_dec_IR_reg[2]/NET0131  & \core_c_dec_IR_reg[3]/NET0131  ;
  assign n6098 = ~n6075 & n6097 ;
  assign n6100 = ~n6096 & ~n6098 ;
  assign n6101 = n6099 & n6100 ;
  assign n6102 = n4055 & n6101 ;
  assign n6103 = ~n6090 & ~n6102 ;
  assign n6104 = ~n6049 & ~n6103 ;
  assign n6105 = n5949 & ~n6104 ;
  assign n6106 = ~\core_c_dec_Post1_E_reg/P0001  & n5955 ;
  assign n6112 = \core_c_psq_MSTAT_reg_DO_reg[1]/NET0131  & ~n6111 ;
  assign n6113 = n6106 & n6112 ;
  assign n6124 = n6105 & ~n6113 ;
  assign n6125 = ~n6123 & n6124 ;
  assign n6126 = ~n5936 & ~n6125 ;
  assign n6127 = ~\core_c_psq_MSTAT_reg_DO_reg[1]/NET0131  & ~n6111 ;
  assign n6128 = ~n5936 & ~n6127 ;
  assign n6129 = ~n6106 & ~n6128 ;
  assign n6130 = n6103 & n6129 ;
  assign n6131 = n5949 & ~n6111 ;
  assign n6132 = n6049 & n6131 ;
  assign n6133 = ~n6103 & n6132 ;
  assign n6134 = ~n6130 & ~n6133 ;
  assign n6135 = ~n6126 & n6134 ;
  assign n6177 = ~\core_dag_ilm1reg_L_reg[6]/NET0131  & ~\core_dag_ilm1reg_L_reg[7]/NET0131  ;
  assign n6178 = ~\core_dag_ilm1reg_L_reg[12]/NET0131  & ~\core_dag_ilm1reg_L_reg[13]/NET0131  ;
  assign n6179 = ~\core_dag_ilm1reg_L_reg[11]/NET0131  & n6178 ;
  assign n6180 = ~\core_dag_ilm1reg_L_reg[10]/NET0131  & ~\core_dag_ilm1reg_L_reg[9]/NET0131  ;
  assign n6181 = ~\core_dag_ilm1reg_L_reg[8]/NET0131  & n6180 ;
  assign n6182 = n6179 & n6181 ;
  assign n6183 = n6177 & n6182 ;
  assign n6184 = ~\core_dag_ilm1reg_L_reg[4]/NET0131  & ~\core_dag_ilm1reg_L_reg[5]/NET0131  ;
  assign n6185 = ~\core_dag_ilm1reg_L_reg[3]/NET0131  & n6184 ;
  assign n6186 = n6183 & n6185 ;
  assign n6187 = ~\core_dag_ilm1reg_L_reg[1]/NET0131  & ~\core_dag_ilm1reg_L_reg[2]/NET0131  ;
  assign n6188 = n6186 & n6187 ;
  assign n6189 = \core_dag_ilm1reg_L_reg[0]/NET0131  & ~n6188 ;
  assign n6190 = ~\core_dag_ilm1reg_L_reg[6]/NET0131  & n6184 ;
  assign n6191 = ~\core_dag_ilm1reg_L_reg[7]/NET0131  & ~\core_dag_ilm1reg_L_reg[8]/NET0131  ;
  assign n6192 = ~\core_dag_ilm1reg_L_reg[10]/NET0131  & n6179 ;
  assign n6193 = ~\core_dag_ilm1reg_L_reg[9]/NET0131  & n6192 ;
  assign n6194 = n6191 & n6193 ;
  assign n6195 = ~n6190 & ~n6194 ;
  assign n6196 = ~n6191 & ~n6193 ;
  assign n6204 = \core_dag_ilm1reg_L_reg[6]/NET0131  & ~n6184 ;
  assign n6201 = \core_dag_ilm1reg_L_reg[11]/NET0131  & ~n6178 ;
  assign n6198 = \core_dag_ilm1reg_L_reg[12]/NET0131  & \core_dag_ilm1reg_L_reg[13]/NET0131  ;
  assign n6199 = \core_dag_ilm1reg_L_reg[4]/NET0131  & \core_dag_ilm1reg_L_reg[5]/NET0131  ;
  assign n6208 = ~n6198 & ~n6199 ;
  assign n6211 = ~n6201 & n6208 ;
  assign n6212 = ~n6204 & n6211 ;
  assign n6197 = ~n6179 & ~n6180 ;
  assign n6203 = \core_dag_ilm1reg_L_reg[1]/NET0131  & \core_dag_ilm1reg_L_reg[2]/NET0131  ;
  assign n6200 = \core_dag_ilm1reg_L_reg[10]/NET0131  & \core_dag_ilm1reg_L_reg[9]/NET0131  ;
  assign n6202 = \core_dag_ilm1reg_L_reg[7]/NET0131  & \core_dag_ilm1reg_L_reg[8]/NET0131  ;
  assign n6209 = ~n6200 & ~n6202 ;
  assign n6210 = ~n6203 & n6209 ;
  assign n6213 = ~n6197 & n6210 ;
  assign n6214 = n6212 & n6213 ;
  assign n6215 = ~n6196 & n6214 ;
  assign n6216 = ~n6195 & n6215 ;
  assign n6205 = ~n6186 & ~n6187 ;
  assign n6206 = n6183 & n6184 ;
  assign n6207 = \core_dag_ilm1reg_L_reg[3]/NET0131  & ~n6206 ;
  assign n6217 = ~n6205 & ~n6207 ;
  assign n6218 = n6216 & n6217 ;
  assign n6219 = ~n6189 & n6218 ;
  assign n6220 = \core_dag_ilm1reg_L_reg[13]/NET0131  & ~n6219 ;
  assign n6221 = ~\core_dag_ilm1reg_L_reg[0]/NET0131  & ~\core_dag_ilm1reg_L_reg[1]/NET0131  ;
  assign n6222 = ~\core_dag_ilm1reg_L_reg[2]/NET0131  & n6221 ;
  assign n6223 = ~\core_dag_ilm1reg_L_reg[3]/NET0131  & n6222 ;
  assign n6224 = n6184 & n6223 ;
  assign n6225 = n6177 & n6224 ;
  assign n6226 = n6219 & n6225 ;
  assign n6227 = n6181 & n6226 ;
  assign n6228 = n6179 & n6227 ;
  assign n6229 = ~n6220 & ~n6228 ;
  assign n6230 = \core_dag_ilm1reg_I_reg[13]/NET0131  & ~n6229 ;
  assign n6231 = ~\core_dag_ilm1reg_L_reg[13]/NET0131  & ~n6230 ;
  assign n6232 = \core_dag_ilm1reg_L_reg[13]/NET0131  & ~\core_dag_ilm1reg_M_reg[13]/NET0131  ;
  assign n6233 = ~n6231 & ~n6232 ;
  assign n6299 = ~\core_dag_ilm1reg_L_reg[3]/NET0131  & ~\core_dag_ilm1reg_M_reg[13]/NET0131  ;
  assign n6300 = \core_dag_ilm1reg_L_reg[3]/NET0131  & \core_dag_ilm1reg_M_reg[13]/NET0131  ;
  assign n6301 = ~n6299 & ~n6300 ;
  assign n6235 = n6219 & ~n6223 ;
  assign n6294 = n6186 & ~n6219 ;
  assign n6295 = ~n6235 & ~n6294 ;
  assign n6296 = \core_dag_ilm1reg_I_reg[3]/NET0131  & n6295 ;
  assign n6297 = \core_dag_ilm1reg_M_reg[3]/NET0131  & n6296 ;
  assign n6298 = ~\core_dag_ilm1reg_M_reg[3]/NET0131  & ~n6296 ;
  assign n6310 = ~n6297 & ~n6298 ;
  assign n6311 = ~n6301 & n6310 ;
  assign n6312 = n6301 & ~n6310 ;
  assign n6313 = ~n6311 & ~n6312 ;
  assign n6314 = n6219 & ~n6222 ;
  assign n6315 = ~\core_dag_ilm1reg_L_reg[2]/NET0131  & n6186 ;
  assign n6316 = ~n6219 & n6315 ;
  assign n6317 = ~n6314 & ~n6316 ;
  assign n6318 = \core_dag_ilm1reg_I_reg[2]/NET0131  & n6317 ;
  assign n6319 = \core_dag_ilm1reg_M_reg[2]/NET0131  & n6318 ;
  assign n6320 = ~\core_dag_ilm1reg_M_reg[2]/NET0131  & ~n6318 ;
  assign n6321 = ~\core_dag_ilm1reg_L_reg[2]/NET0131  & ~\core_dag_ilm1reg_M_reg[13]/NET0131  ;
  assign n6322 = \core_dag_ilm1reg_L_reg[2]/NET0131  & \core_dag_ilm1reg_M_reg[13]/NET0131  ;
  assign n6323 = ~n6321 & ~n6322 ;
  assign n6324 = ~n6320 & ~n6323 ;
  assign n6325 = ~n6319 & ~n6324 ;
  assign n6326 = n6313 & ~n6325 ;
  assign n6327 = ~n6313 & n6325 ;
  assign n6329 = n6219 & ~n6221 ;
  assign n6328 = n6188 & ~n6218 ;
  assign n6330 = \core_dag_ilm1reg_I_reg[1]/NET0131  & ~n6328 ;
  assign n6331 = ~n6329 & n6330 ;
  assign n6332 = \core_dag_ilm1reg_M_reg[1]/NET0131  & n6331 ;
  assign n6333 = ~\core_dag_ilm1reg_M_reg[1]/NET0131  & ~n6331 ;
  assign n6334 = ~\core_dag_ilm1reg_L_reg[1]/NET0131  & ~\core_dag_ilm1reg_M_reg[13]/NET0131  ;
  assign n6335 = \core_dag_ilm1reg_L_reg[1]/NET0131  & \core_dag_ilm1reg_M_reg[13]/NET0131  ;
  assign n6336 = ~n6334 & ~n6335 ;
  assign n6337 = ~n6333 & ~n6336 ;
  assign n6338 = ~n6332 & ~n6337 ;
  assign n6339 = ~n6319 & ~n6320 ;
  assign n6340 = n6323 & ~n6339 ;
  assign n6341 = ~n6323 & n6339 ;
  assign n6342 = ~n6340 & ~n6341 ;
  assign n6343 = ~n6338 & n6342 ;
  assign n6344 = n6338 & ~n6342 ;
  assign n6346 = n6221 & n6316 ;
  assign n6345 = \core_dag_ilm1reg_L_reg[0]/NET0131  & n6219 ;
  assign n6347 = \core_dag_ilm1reg_I_reg[0]/NET0131  & ~n6345 ;
  assign n6348 = ~n6346 & n6347 ;
  assign n6349 = ~\core_dag_ilm1reg_M_reg[0]/NET0131  & ~n6348 ;
  assign n6350 = \core_dag_ilm1reg_M_reg[0]/NET0131  & n6348 ;
  assign n6351 = ~\core_dag_ilm1reg_L_reg[0]/NET0131  & ~\core_dag_ilm1reg_M_reg[13]/NET0131  ;
  assign n6352 = \core_dag_ilm1reg_L_reg[0]/NET0131  & \core_dag_ilm1reg_M_reg[13]/NET0131  ;
  assign n6353 = ~n6351 & ~n6352 ;
  assign n6354 = ~n6350 & n6353 ;
  assign n6355 = ~n6349 & ~n6354 ;
  assign n6356 = ~n6332 & ~n6333 ;
  assign n6357 = n6336 & ~n6356 ;
  assign n6358 = ~n6336 & n6356 ;
  assign n6359 = ~n6357 & ~n6358 ;
  assign n6360 = ~n6355 & ~n6359 ;
  assign n6361 = n6355 & n6359 ;
  assign n6362 = ~n6349 & ~n6350 ;
  assign n6363 = ~n6353 & n6362 ;
  assign n6364 = n6353 & ~n6362 ;
  assign n6365 = ~n6363 & ~n6364 ;
  assign n6366 = ~\core_dag_ilm1reg_M_reg[13]/NET0131  & n6365 ;
  assign n6367 = ~n6361 & ~n6366 ;
  assign n6368 = ~n6360 & ~n6367 ;
  assign n6369 = ~n6344 & n6368 ;
  assign n6370 = ~n6343 & ~n6369 ;
  assign n6371 = ~n6327 & ~n6370 ;
  assign n6372 = ~n6326 & ~n6371 ;
  assign n6236 = ~n6190 & n6219 ;
  assign n6234 = n6183 & ~n6219 ;
  assign n6237 = ~n6234 & ~n6235 ;
  assign n6238 = ~n6236 & n6237 ;
  assign n6239 = \core_dag_ilm1reg_I_reg[6]/NET0131  & n6238 ;
  assign n6240 = ~\core_dag_ilm1reg_M_reg[6]/NET0131  & ~n6239 ;
  assign n6241 = \core_dag_ilm1reg_M_reg[6]/NET0131  & n6239 ;
  assign n6242 = ~n6240 & ~n6241 ;
  assign n6243 = ~\core_dag_ilm1reg_L_reg[6]/NET0131  & ~\core_dag_ilm1reg_M_reg[13]/NET0131  ;
  assign n6244 = \core_dag_ilm1reg_L_reg[6]/NET0131  & \core_dag_ilm1reg_M_reg[13]/NET0131  ;
  assign n6245 = ~n6243 & ~n6244 ;
  assign n6246 = n6242 & ~n6245 ;
  assign n6247 = ~n6242 & n6245 ;
  assign n6248 = ~n6246 & ~n6247 ;
  assign n6249 = n6219 & ~n6224 ;
  assign n6250 = ~\core_dag_ilm1reg_L_reg[5]/NET0131  & n6234 ;
  assign n6251 = ~n6249 & ~n6250 ;
  assign n6252 = \core_dag_ilm1reg_I_reg[5]/NET0131  & n6251 ;
  assign n6253 = \core_dag_ilm1reg_M_reg[5]/NET0131  & n6252 ;
  assign n6254 = ~\core_dag_ilm1reg_M_reg[5]/NET0131  & ~n6252 ;
  assign n6255 = ~\core_dag_ilm1reg_L_reg[5]/NET0131  & ~\core_dag_ilm1reg_M_reg[13]/NET0131  ;
  assign n6256 = \core_dag_ilm1reg_L_reg[5]/NET0131  & \core_dag_ilm1reg_M_reg[13]/NET0131  ;
  assign n6257 = ~n6255 & ~n6256 ;
  assign n6258 = ~n6254 & ~n6257 ;
  assign n6259 = ~n6253 & ~n6258 ;
  assign n6260 = ~n6248 & n6259 ;
  assign n6261 = ~n6194 & ~n6219 ;
  assign n6262 = ~n6226 & ~n6261 ;
  assign n6263 = \core_dag_ilm1reg_I_reg[7]/NET0131  & ~n6262 ;
  assign n6264 = ~\core_dag_ilm1reg_M_reg[7]/NET0131  & ~n6263 ;
  assign n6265 = \core_dag_ilm1reg_M_reg[7]/NET0131  & n6263 ;
  assign n6266 = ~n6264 & ~n6265 ;
  assign n6267 = ~\core_dag_ilm1reg_L_reg[7]/NET0131  & ~\core_dag_ilm1reg_M_reg[13]/NET0131  ;
  assign n6268 = \core_dag_ilm1reg_L_reg[7]/NET0131  & \core_dag_ilm1reg_M_reg[13]/NET0131  ;
  assign n6269 = ~n6267 & ~n6268 ;
  assign n6270 = n6266 & ~n6269 ;
  assign n6271 = ~n6266 & n6269 ;
  assign n6272 = ~n6270 & ~n6271 ;
  assign n6273 = ~n6240 & ~n6245 ;
  assign n6274 = ~n6241 & ~n6273 ;
  assign n6275 = ~n6272 & n6274 ;
  assign n6276 = ~n6260 & ~n6275 ;
  assign n6277 = ~\core_dag_ilm1reg_L_reg[4]/NET0131  & n6223 ;
  assign n6278 = n6219 & ~n6277 ;
  assign n6279 = n6184 & n6234 ;
  assign n6280 = ~n6278 & ~n6279 ;
  assign n6281 = \core_dag_ilm1reg_I_reg[4]/NET0131  & n6280 ;
  assign n6282 = \core_dag_ilm1reg_M_reg[4]/NET0131  & n6281 ;
  assign n6283 = ~\core_dag_ilm1reg_M_reg[4]/NET0131  & ~n6281 ;
  assign n6284 = ~\core_dag_ilm1reg_L_reg[4]/NET0131  & ~\core_dag_ilm1reg_M_reg[13]/NET0131  ;
  assign n6285 = \core_dag_ilm1reg_L_reg[4]/NET0131  & \core_dag_ilm1reg_M_reg[13]/NET0131  ;
  assign n6286 = ~n6284 & ~n6285 ;
  assign n6287 = ~n6283 & ~n6286 ;
  assign n6288 = ~n6282 & ~n6287 ;
  assign n6289 = ~n6253 & ~n6254 ;
  assign n6290 = n6257 & ~n6289 ;
  assign n6291 = ~n6257 & n6289 ;
  assign n6292 = ~n6290 & ~n6291 ;
  assign n6293 = n6288 & ~n6292 ;
  assign n6302 = ~n6298 & ~n6301 ;
  assign n6303 = ~n6297 & ~n6302 ;
  assign n6304 = ~n6282 & ~n6283 ;
  assign n6305 = n6286 & ~n6304 ;
  assign n6306 = ~n6286 & n6304 ;
  assign n6307 = ~n6305 & ~n6306 ;
  assign n6308 = n6303 & ~n6307 ;
  assign n6309 = ~n6293 & ~n6308 ;
  assign n6373 = n6276 & n6309 ;
  assign n6374 = ~n6372 & n6373 ;
  assign n6377 = ~n6288 & n6292 ;
  assign n6378 = ~n6303 & n6307 ;
  assign n6379 = ~n6293 & n6378 ;
  assign n6380 = ~n6377 & ~n6379 ;
  assign n6381 = n6276 & ~n6380 ;
  assign n6375 = n6248 & ~n6259 ;
  assign n6376 = ~n6275 & n6375 ;
  assign n6382 = n6272 & ~n6274 ;
  assign n6383 = ~n6376 & ~n6382 ;
  assign n6384 = ~n6381 & n6383 ;
  assign n6385 = ~n6374 & n6384 ;
  assign n6386 = ~\core_dag_ilm1reg_L_reg[8]/NET0131  & n6226 ;
  assign n6387 = ~\core_dag_ilm1reg_L_reg[9]/NET0131  & n6386 ;
  assign n6388 = ~n6193 & ~n6219 ;
  assign n6389 = ~n6387 & ~n6388 ;
  assign n6390 = \core_dag_ilm1reg_I_reg[9]/NET0131  & ~n6389 ;
  assign n6391 = ~\core_dag_ilm1reg_M_reg[9]/NET0131  & ~n6390 ;
  assign n6392 = \core_dag_ilm1reg_M_reg[9]/NET0131  & n6390 ;
  assign n6393 = ~n6391 & ~n6392 ;
  assign n6394 = ~\core_dag_ilm1reg_L_reg[9]/NET0131  & ~\core_dag_ilm1reg_M_reg[13]/NET0131  ;
  assign n6395 = \core_dag_ilm1reg_L_reg[9]/NET0131  & \core_dag_ilm1reg_M_reg[13]/NET0131  ;
  assign n6396 = ~n6394 & ~n6395 ;
  assign n6397 = n6393 & ~n6396 ;
  assign n6398 = ~n6393 & n6396 ;
  assign n6399 = ~n6397 & ~n6398 ;
  assign n6400 = ~n6182 & ~n6219 ;
  assign n6401 = ~n6386 & ~n6400 ;
  assign n6402 = \core_dag_ilm1reg_I_reg[8]/NET0131  & ~n6401 ;
  assign n6403 = \core_dag_ilm1reg_M_reg[8]/NET0131  & n6402 ;
  assign n6404 = ~\core_dag_ilm1reg_M_reg[8]/NET0131  & ~n6402 ;
  assign n6405 = ~\core_dag_ilm1reg_L_reg[8]/NET0131  & ~\core_dag_ilm1reg_M_reg[13]/NET0131  ;
  assign n6406 = \core_dag_ilm1reg_L_reg[8]/NET0131  & \core_dag_ilm1reg_M_reg[13]/NET0131  ;
  assign n6407 = ~n6405 & ~n6406 ;
  assign n6408 = ~n6404 & ~n6407 ;
  assign n6409 = ~n6403 & ~n6408 ;
  assign n6410 = ~n6399 & n6409 ;
  assign n6411 = ~n6264 & ~n6269 ;
  assign n6412 = ~n6265 & ~n6411 ;
  assign n6413 = ~n6403 & ~n6404 ;
  assign n6414 = n6407 & ~n6413 ;
  assign n6415 = ~n6407 & n6413 ;
  assign n6416 = ~n6414 & ~n6415 ;
  assign n6417 = n6412 & ~n6416 ;
  assign n6418 = ~n6410 & ~n6417 ;
  assign n6419 = ~n6385 & n6418 ;
  assign n6420 = ~n6391 & ~n6396 ;
  assign n6421 = ~n6392 & ~n6420 ;
  assign n6422 = ~n6192 & ~n6219 ;
  assign n6423 = ~n6227 & ~n6422 ;
  assign n6424 = \core_dag_ilm1reg_I_reg[10]/NET0131  & ~n6423 ;
  assign n6425 = ~\core_dag_ilm1reg_M_reg[10]/NET0131  & ~n6424 ;
  assign n6426 = \core_dag_ilm1reg_M_reg[10]/NET0131  & n6424 ;
  assign n6427 = ~n6425 & ~n6426 ;
  assign n6428 = ~\core_dag_ilm1reg_L_reg[10]/NET0131  & ~\core_dag_ilm1reg_M_reg[13]/NET0131  ;
  assign n6429 = \core_dag_ilm1reg_L_reg[10]/NET0131  & \core_dag_ilm1reg_M_reg[13]/NET0131  ;
  assign n6430 = ~n6428 & ~n6429 ;
  assign n6431 = n6427 & ~n6430 ;
  assign n6432 = ~n6427 & n6430 ;
  assign n6433 = ~n6431 & ~n6432 ;
  assign n6434 = n6421 & ~n6433 ;
  assign n6435 = ~n6425 & ~n6430 ;
  assign n6436 = ~n6426 & ~n6435 ;
  assign n6437 = ~\core_dag_ilm1reg_L_reg[11]/NET0131  & n6181 ;
  assign n6438 = n6225 & n6437 ;
  assign n6439 = n6219 & ~n6438 ;
  assign n6440 = n6178 & ~n6219 ;
  assign n6441 = ~\core_dag_ilm1reg_L_reg[11]/NET0131  & n6440 ;
  assign n6442 = ~n6439 & ~n6441 ;
  assign n6443 = \core_dag_ilm1reg_I_reg[11]/NET0131  & n6442 ;
  assign n6444 = \core_dag_ilm1reg_M_reg[11]/NET0131  & n6443 ;
  assign n6445 = ~\core_dag_ilm1reg_M_reg[11]/NET0131  & ~n6443 ;
  assign n6446 = ~n6444 & ~n6445 ;
  assign n6447 = ~\core_dag_ilm1reg_L_reg[11]/NET0131  & ~\core_dag_ilm1reg_M_reg[13]/NET0131  ;
  assign n6448 = \core_dag_ilm1reg_L_reg[11]/NET0131  & \core_dag_ilm1reg_M_reg[13]/NET0131  ;
  assign n6449 = ~n6447 & ~n6448 ;
  assign n6450 = n6446 & ~n6449 ;
  assign n6451 = ~n6446 & n6449 ;
  assign n6452 = ~n6450 & ~n6451 ;
  assign n6453 = n6436 & ~n6452 ;
  assign n6454 = ~n6434 & ~n6453 ;
  assign n6455 = n6419 & n6454 ;
  assign n6456 = ~n6436 & n6452 ;
  assign n6457 = ~n6421 & n6433 ;
  assign n6458 = n6399 & ~n6409 ;
  assign n6459 = ~n6412 & n6416 ;
  assign n6460 = ~n6410 & n6459 ;
  assign n6461 = ~n6458 & ~n6460 ;
  assign n6462 = ~n6457 & n6461 ;
  assign n6463 = n6454 & ~n6462 ;
  assign n6464 = ~n6456 & ~n6463 ;
  assign n6465 = ~n6455 & n6464 ;
  assign n6466 = \core_dag_ilm1reg_L_reg[13]/NET0131  & n6230 ;
  assign n6467 = ~n6231 & ~n6466 ;
  assign n6468 = \core_dag_ilm1reg_L_reg[12]/NET0131  & n6219 ;
  assign n6469 = ~n6439 & ~n6440 ;
  assign n6470 = ~n6468 & n6469 ;
  assign n6471 = \core_dag_ilm1reg_I_reg[12]/NET0131  & n6470 ;
  assign n6472 = ~\core_dag_ilm1reg_M_reg[12]/NET0131  & ~n6471 ;
  assign n6473 = \core_dag_ilm1reg_M_reg[12]/NET0131  & n6471 ;
  assign n6474 = ~\core_dag_ilm1reg_L_reg[12]/NET0131  & ~\core_dag_ilm1reg_M_reg[13]/NET0131  ;
  assign n6475 = \core_dag_ilm1reg_L_reg[12]/NET0131  & \core_dag_ilm1reg_M_reg[13]/NET0131  ;
  assign n6476 = ~n6474 & ~n6475 ;
  assign n6477 = ~n6473 & n6476 ;
  assign n6478 = ~n6472 & ~n6477 ;
  assign n6479 = n6467 & ~n6478 ;
  assign n6480 = ~n6445 & ~n6449 ;
  assign n6481 = ~n6444 & ~n6480 ;
  assign n6482 = ~n6472 & ~n6473 ;
  assign n6483 = ~n6476 & n6482 ;
  assign n6484 = n6476 & ~n6482 ;
  assign n6485 = ~n6483 & ~n6484 ;
  assign n6486 = n6481 & ~n6485 ;
  assign n6487 = ~n6479 & ~n6486 ;
  assign n6488 = ~n6465 & n6487 ;
  assign n6489 = ~n6467 & n6478 ;
  assign n6490 = ~n6481 & n6485 ;
  assign n6491 = ~n6479 & n6490 ;
  assign n6492 = ~n6489 & ~n6491 ;
  assign n6493 = ~n6488 & n6492 ;
  assign n6494 = ~n6233 & n6493 ;
  assign n6495 = n6233 & ~n6493 ;
  assign n6496 = ~n6494 & ~n6495 ;
  assign n6532 = ~n6479 & ~n6489 ;
  assign n6533 = ~n6465 & ~n6486 ;
  assign n6534 = ~n6490 & ~n6533 ;
  assign n6535 = n6532 & ~n6534 ;
  assign n6536 = ~n6532 & n6534 ;
  assign n6537 = ~n6535 & ~n6536 ;
  assign n6538 = n6496 & ~n6537 ;
  assign n6497 = \core_dag_ilm1reg_M_reg[13]/NET0131  & ~n6230 ;
  assign n6498 = ~\core_dag_ilm1reg_M_reg[13]/NET0131  & n6230 ;
  assign n6499 = ~n6497 & ~n6498 ;
  assign n6500 = ~n6332 & ~n6350 ;
  assign n6501 = ~n6333 & ~n6500 ;
  assign n6502 = ~n6319 & ~n6501 ;
  assign n6503 = ~n6320 & ~n6502 ;
  assign n6504 = ~n6297 & ~n6503 ;
  assign n6505 = ~n6298 & ~n6504 ;
  assign n6506 = ~n6254 & ~n6283 ;
  assign n6507 = n6505 & n6506 ;
  assign n6508 = ~n6254 & n6282 ;
  assign n6509 = ~n6253 & ~n6508 ;
  assign n6510 = ~n6507 & n6509 ;
  assign n6511 = ~n6240 & ~n6510 ;
  assign n6512 = ~n6241 & ~n6265 ;
  assign n6513 = ~n6511 & n6512 ;
  assign n6514 = ~n6264 & ~n6513 ;
  assign n6515 = ~n6391 & ~n6404 ;
  assign n6516 = n6514 & n6515 ;
  assign n6517 = ~n6425 & ~n6445 ;
  assign n6518 = n6516 & n6517 ;
  assign n6520 = ~n6392 & ~n6403 ;
  assign n6521 = ~n6391 & ~n6520 ;
  assign n6522 = n6517 & n6521 ;
  assign n6519 = n6426 & ~n6445 ;
  assign n6523 = ~n6444 & ~n6519 ;
  assign n6524 = ~n6522 & n6523 ;
  assign n6525 = ~n6518 & n6524 ;
  assign n6526 = ~n6472 & ~n6525 ;
  assign n6527 = ~n6473 & ~n6526 ;
  assign n6528 = n6499 & n6527 ;
  assign n6529 = ~n6499 & ~n6527 ;
  assign n6530 = ~n6528 & ~n6529 ;
  assign n6531 = ~n6496 & ~n6530 ;
  assign n6539 = ~\core_dag_ilm1reg_M_reg[13]/NET0131  & ~n6531 ;
  assign n6540 = ~n6538 & n6539 ;
  assign n6541 = ~\core_dag_ilm1reg_I_reg[13]/NET0131  & ~n6537 ;
  assign n6542 = \core_dag_ilm1reg_M_reg[13]/NET0131  & n6530 ;
  assign n6543 = ~n6541 & n6542 ;
  assign n6544 = \core_dag_ilm1reg_I_reg[13]/NET0131  & n6229 ;
  assign n6545 = ~n6543 & ~n6544 ;
  assign n6546 = ~n6540 & n6545 ;
  assign n6547 = n6135 & ~n6546 ;
  assign n6136 = \core_dag_ilm1reg_I0_we_DO_reg[13]/NET0131  & n6058 ;
  assign n6137 = n6060 & n6136 ;
  assign n6144 = ~n4055 & ~n6137 ;
  assign n6142 = n6067 & n6068 ;
  assign n6143 = \core_dag_ilm1reg_I1_we_DO_reg[13]/NET0131  & n6142 ;
  assign n6138 = n6084 & n6085 ;
  assign n6139 = \core_dag_ilm1reg_I2_we_DO_reg[13]/NET0131  & n6138 ;
  assign n6140 = n6075 & n6077 ;
  assign n6141 = \core_dag_ilm1reg_I3_we_DO_reg[13]/NET0131  & n6140 ;
  assign n6145 = ~n6139 & ~n6141 ;
  assign n6146 = ~n6143 & n6145 ;
  assign n6147 = n6144 & n6146 ;
  assign n6148 = n6058 & n6093 ;
  assign n6149 = \core_dag_ilm1reg_I0_we_DO_reg[13]/NET0131  & n6148 ;
  assign n6150 = n6075 & n6097 ;
  assign n6151 = \core_dag_ilm1reg_I3_we_DO_reg[13]/NET0131  & n6150 ;
  assign n6156 = ~n6149 & ~n6151 ;
  assign n6152 = n6084 & n6095 ;
  assign n6153 = \core_dag_ilm1reg_I2_we_DO_reg[13]/NET0131  & n6152 ;
  assign n6154 = n6067 & n6091 ;
  assign n6155 = \core_dag_ilm1reg_I1_we_DO_reg[13]/NET0131  & n6154 ;
  assign n6157 = ~n6153 & ~n6155 ;
  assign n6158 = n6156 & n6157 ;
  assign n6159 = n4055 & n6158 ;
  assign n6160 = ~n6147 & ~n6159 ;
  assign n6161 = ~n6135 & n6160 ;
  assign n6164 = ~\core_c_dec_Post2_E_reg/P0001  & n5955 ;
  assign n6165 = ~n6121 & n6164 ;
  assign n6166 = n6049 & n6165 ;
  assign n6167 = n6111 & ~n6166 ;
  assign n6163 = n6103 & n6113 ;
  assign n6168 = n5949 & ~n6163 ;
  assign n6169 = ~n6167 & n6168 ;
  assign n6170 = ~n5936 & ~n6169 ;
  assign n6162 = n5936 & n6104 ;
  assign n6171 = ~n6131 & n6164 ;
  assign n6172 = ~n6103 & ~n6171 ;
  assign n6173 = \core_c_psq_MSTAT_reg_DO_reg[1]/NET0131  & n6131 ;
  assign n6174 = n6172 & ~n6173 ;
  assign n6175 = ~n6162 & ~n6174 ;
  assign n6176 = ~n6170 & n6175 ;
  assign n6548 = ~n6161 & n6176 ;
  assign n6549 = ~n6547 & n6548 ;
  assign n6550 = ~\core_dag_ilm2reg_L_reg[0]/NET0131  & ~\core_dag_ilm2reg_L_reg[1]/NET0131  ;
  assign n6551 = ~\core_dag_ilm2reg_L_reg[2]/NET0131  & n6550 ;
  assign n6552 = ~\core_dag_ilm2reg_L_reg[12]/NET0131  & ~\core_dag_ilm2reg_L_reg[13]/NET0131  ;
  assign n6553 = ~\core_dag_ilm2reg_L_reg[10]/NET0131  & ~\core_dag_ilm2reg_L_reg[11]/NET0131  ;
  assign n6554 = n6552 & n6553 ;
  assign n6555 = ~\core_dag_ilm2reg_L_reg[7]/NET0131  & ~\core_dag_ilm2reg_L_reg[8]/NET0131  ;
  assign n6556 = ~\core_dag_ilm2reg_L_reg[9]/NET0131  & n6555 ;
  assign n6557 = n6554 & n6556 ;
  assign n6558 = ~\core_dag_ilm2reg_L_reg[5]/NET0131  & ~\core_dag_ilm2reg_L_reg[6]/NET0131  ;
  assign n6559 = ~\core_dag_ilm2reg_L_reg[4]/NET0131  & n6558 ;
  assign n6560 = n6557 & n6559 ;
  assign n6561 = ~\core_dag_ilm2reg_L_reg[3]/NET0131  & n6560 ;
  assign n6562 = ~n6551 & ~n6561 ;
  assign n6563 = ~n6556 & ~n6558 ;
  assign n6564 = n6554 & ~n6563 ;
  assign n6565 = ~\core_dag_ilm2reg_L_reg[11]/NET0131  & n6552 ;
  assign n6566 = \core_dag_ilm2reg_L_reg[10]/NET0131  & ~n6565 ;
  assign n6567 = ~\core_dag_ilm2reg_L_reg[9]/NET0131  & n6558 ;
  assign n6568 = ~n6566 & n6567 ;
  assign n6569 = ~n6564 & ~n6568 ;
  assign n6570 = ~\core_dag_ilm2reg_L_reg[9]/NET0131  & n6554 ;
  assign n6571 = ~n6555 & ~n6570 ;
  assign n6577 = \core_dag_ilm2reg_L_reg[5]/NET0131  & \core_dag_ilm2reg_L_reg[6]/NET0131  ;
  assign n6575 = \core_dag_ilm2reg_L_reg[12]/NET0131  & \core_dag_ilm2reg_L_reg[13]/NET0131  ;
  assign n6576 = \core_dag_ilm2reg_L_reg[7]/NET0131  & \core_dag_ilm2reg_L_reg[8]/NET0131  ;
  assign n6581 = ~n6575 & ~n6576 ;
  assign n6582 = ~n6577 & n6581 ;
  assign n6572 = \core_dag_ilm2reg_L_reg[11]/NET0131  & ~n6552 ;
  assign n6573 = ~\core_dag_ilm2reg_L_reg[1]/NET0131  & ~\core_dag_ilm2reg_L_reg[2]/NET0131  ;
  assign n6574 = \core_dag_ilm2reg_L_reg[0]/NET0131  & ~n6573 ;
  assign n6583 = ~n6572 & ~n6574 ;
  assign n6584 = n6582 & n6583 ;
  assign n6585 = ~n6571 & n6584 ;
  assign n6586 = ~n6569 & n6585 ;
  assign n6578 = n6557 & n6558 ;
  assign n6579 = \core_dag_ilm2reg_L_reg[4]/NET0131  & ~n6578 ;
  assign n6580 = \core_dag_ilm2reg_L_reg[3]/NET0131  & ~n6560 ;
  assign n6587 = ~n6579 & ~n6580 ;
  assign n6588 = n6586 & n6587 ;
  assign n6589 = \core_dag_ilm2reg_L_reg[1]/NET0131  & \core_dag_ilm2reg_L_reg[2]/NET0131  ;
  assign n6590 = n6588 & ~n6589 ;
  assign n6591 = ~n6562 & n6590 ;
  assign n6592 = \core_dag_ilm2reg_L_reg[0]/NET0131  & n6591 ;
  assign n6594 = \core_dag_ilm2reg_I_reg[0]/NET0131  & ~n6592 ;
  assign n6595 = ~\core_dag_ilm2reg_M_reg[0]/NET0131  & ~n6594 ;
  assign n6596 = \core_dag_ilm2reg_M_reg[0]/NET0131  & n6594 ;
  assign n6597 = ~n6595 & ~n6596 ;
  assign n6598 = \core_dag_ilm2reg_L_reg[13]/NET0131  & ~n6591 ;
  assign n6599 = ~\core_dag_ilm2reg_L_reg[3]/NET0131  & n6551 ;
  assign n6600 = n6559 & n6599 ;
  assign n6601 = n6555 & n6600 ;
  assign n6602 = n6570 & n6601 ;
  assign n6603 = n6591 & n6602 ;
  assign n6604 = ~n6598 & ~n6603 ;
  assign n6605 = \core_dag_ilm2reg_I_reg[13]/NET0131  & ~n6604 ;
  assign n6606 = \core_dag_ilm2reg_M_reg[13]/NET0131  & n6605 ;
  assign n6611 = n6552 & ~n6591 ;
  assign n6607 = ~\core_dag_ilm2reg_L_reg[9]/NET0131  & n6601 ;
  assign n6608 = n6553 & n6607 ;
  assign n6609 = n6591 & ~n6608 ;
  assign n6610 = \core_dag_ilm2reg_L_reg[12]/NET0131  & n6591 ;
  assign n6612 = ~n6609 & ~n6610 ;
  assign n6613 = ~n6611 & n6612 ;
  assign n6614 = \core_dag_ilm2reg_I_reg[12]/NET0131  & n6613 ;
  assign n6615 = \core_dag_ilm2reg_M_reg[12]/NET0131  & n6614 ;
  assign n6616 = ~\core_dag_ilm2reg_M_reg[12]/NET0131  & ~n6614 ;
  assign n6617 = ~\core_dag_ilm2reg_L_reg[10]/NET0131  & n6607 ;
  assign n6618 = n6591 & ~n6617 ;
  assign n6619 = n6553 & n6611 ;
  assign n6620 = ~n6618 & ~n6619 ;
  assign n6621 = \core_dag_ilm2reg_I_reg[10]/NET0131  & n6620 ;
  assign n6622 = ~\core_dag_ilm2reg_M_reg[10]/NET0131  & ~n6621 ;
  assign n6623 = n6565 & ~n6591 ;
  assign n6624 = ~n6609 & ~n6623 ;
  assign n6625 = \core_dag_ilm2reg_I_reg[11]/NET0131  & n6624 ;
  assign n6626 = ~\core_dag_ilm2reg_M_reg[11]/NET0131  & ~n6625 ;
  assign n6627 = ~n6622 & ~n6626 ;
  assign n6628 = n6591 & ~n6607 ;
  assign n6629 = ~\core_dag_ilm2reg_L_reg[9]/NET0131  & n6619 ;
  assign n6630 = ~n6628 & ~n6629 ;
  assign n6631 = \core_dag_ilm2reg_I_reg[9]/NET0131  & n6630 ;
  assign n6632 = ~\core_dag_ilm2reg_M_reg[9]/NET0131  & ~n6631 ;
  assign n6633 = ~\core_dag_ilm2reg_L_reg[8]/NET0131  & n6629 ;
  assign n6634 = n6591 & ~n6601 ;
  assign n6635 = ~n6633 & ~n6634 ;
  assign n6636 = \core_dag_ilm2reg_I_reg[8]/NET0131  & n6635 ;
  assign n6637 = ~\core_dag_ilm2reg_M_reg[8]/NET0131  & ~n6636 ;
  assign n6638 = n6556 & n6619 ;
  assign n6639 = \core_dag_ilm2reg_L_reg[7]/NET0131  & n6591 ;
  assign n6640 = n6591 & ~n6600 ;
  assign n6641 = ~n6639 & ~n6640 ;
  assign n6642 = ~n6638 & n6641 ;
  assign n6643 = \core_dag_ilm2reg_I_reg[7]/NET0131  & n6642 ;
  assign n6644 = ~\core_dag_ilm2reg_M_reg[7]/NET0131  & ~n6643 ;
  assign n6645 = \core_dag_ilm2reg_M_reg[7]/NET0131  & n6643 ;
  assign n6646 = ~\core_dag_ilm2reg_L_reg[6]/NET0131  & n6638 ;
  assign n6647 = ~n6640 & ~n6646 ;
  assign n6648 = \core_dag_ilm2reg_I_reg[6]/NET0131  & n6647 ;
  assign n6649 = ~\core_dag_ilm2reg_M_reg[6]/NET0131  & ~n6648 ;
  assign n6650 = \core_dag_ilm2reg_M_reg[6]/NET0131  & n6648 ;
  assign n6651 = n6591 & ~n6599 ;
  assign n6652 = n6561 & ~n6590 ;
  assign n6653 = ~n6651 & ~n6652 ;
  assign n6654 = \core_dag_ilm2reg_I_reg[3]/NET0131  & n6653 ;
  assign n6655 = ~\core_dag_ilm2reg_M_reg[3]/NET0131  & ~n6654 ;
  assign n6656 = \core_dag_ilm2reg_M_reg[3]/NET0131  & n6654 ;
  assign n6657 = ~n6551 & n6591 ;
  assign n6658 = ~\core_dag_ilm2reg_L_reg[2]/NET0131  & n6561 ;
  assign n6659 = ~n6588 & n6658 ;
  assign n6660 = ~n6657 & ~n6659 ;
  assign n6661 = \core_dag_ilm2reg_I_reg[2]/NET0131  & n6660 ;
  assign n6662 = ~\core_dag_ilm2reg_M_reg[2]/NET0131  & ~n6661 ;
  assign n6663 = \core_dag_ilm2reg_M_reg[2]/NET0131  & n6661 ;
  assign n6664 = ~n6550 & n6591 ;
  assign n6665 = ~\core_dag_ilm2reg_L_reg[1]/NET0131  & n6659 ;
  assign n6666 = \core_dag_ilm2reg_I_reg[1]/NET0131  & ~n6665 ;
  assign n6667 = ~n6664 & n6666 ;
  assign n6668 = ~\core_dag_ilm2reg_M_reg[1]/NET0131  & ~n6667 ;
  assign n6669 = \core_dag_ilm2reg_M_reg[1]/NET0131  & n6667 ;
  assign n6670 = ~n6596 & ~n6669 ;
  assign n6671 = ~n6668 & ~n6670 ;
  assign n6672 = ~n6663 & ~n6671 ;
  assign n6673 = ~n6662 & ~n6672 ;
  assign n6674 = ~n6656 & ~n6673 ;
  assign n6675 = ~n6655 & ~n6674 ;
  assign n6676 = ~n6578 & ~n6591 ;
  assign n6677 = ~\core_dag_ilm2reg_L_reg[4]/NET0131  & n6599 ;
  assign n6678 = n6591 & n6677 ;
  assign n6679 = ~\core_dag_ilm2reg_L_reg[5]/NET0131  & n6678 ;
  assign n6680 = ~n6676 & ~n6679 ;
  assign n6681 = \core_dag_ilm2reg_I_reg[5]/NET0131  & ~n6680 ;
  assign n6682 = ~\core_dag_ilm2reg_M_reg[5]/NET0131  & ~n6681 ;
  assign n6683 = ~n6560 & ~n6591 ;
  assign n6684 = ~n6678 & ~n6683 ;
  assign n6685 = \core_dag_ilm2reg_I_reg[4]/NET0131  & ~n6684 ;
  assign n6686 = ~\core_dag_ilm2reg_M_reg[4]/NET0131  & ~n6685 ;
  assign n6687 = ~n6682 & ~n6686 ;
  assign n6688 = n6675 & n6687 ;
  assign n6689 = \core_dag_ilm2reg_M_reg[5]/NET0131  & n6681 ;
  assign n6690 = \core_dag_ilm2reg_M_reg[4]/NET0131  & n6685 ;
  assign n6691 = ~n6682 & n6690 ;
  assign n6692 = ~n6689 & ~n6691 ;
  assign n6693 = ~n6688 & n6692 ;
  assign n6694 = ~n6650 & n6693 ;
  assign n6695 = ~n6649 & ~n6694 ;
  assign n6696 = ~n6645 & ~n6695 ;
  assign n6697 = ~n6644 & ~n6696 ;
  assign n6698 = ~n6637 & n6697 ;
  assign n6699 = ~n6632 & n6698 ;
  assign n6700 = n6627 & n6699 ;
  assign n6701 = \core_dag_ilm2reg_M_reg[11]/NET0131  & n6625 ;
  assign n6702 = \core_dag_ilm2reg_M_reg[10]/NET0131  & n6621 ;
  assign n6703 = \core_dag_ilm2reg_M_reg[8]/NET0131  & n6636 ;
  assign n6704 = \core_dag_ilm2reg_M_reg[9]/NET0131  & n6631 ;
  assign n6705 = ~n6703 & ~n6704 ;
  assign n6706 = ~n6632 & ~n6705 ;
  assign n6707 = ~n6702 & ~n6706 ;
  assign n6708 = n6627 & ~n6707 ;
  assign n6709 = ~n6701 & ~n6708 ;
  assign n6710 = ~n6700 & n6709 ;
  assign n6711 = ~n6616 & ~n6710 ;
  assign n6712 = ~n6615 & ~n6711 ;
  assign n6713 = ~n6606 & n6712 ;
  assign n6714 = \core_dag_ilm2reg_M_reg[13]/NET0131  & ~n6713 ;
  assign n6715 = n6605 & ~n6712 ;
  assign n6716 = ~\core_dag_ilm2reg_M_reg[13]/NET0131  & ~n6715 ;
  assign n6717 = ~n6714 & ~n6716 ;
  assign n6718 = n6597 & ~n6717 ;
  assign n6719 = ~\core_dag_ilm2reg_L_reg[0]/NET0131  & ~\core_dag_ilm2reg_M_reg[13]/NET0131  ;
  assign n6720 = \core_dag_ilm2reg_L_reg[0]/NET0131  & \core_dag_ilm2reg_M_reg[13]/NET0131  ;
  assign n6721 = ~n6719 & ~n6720 ;
  assign n6722 = ~n6597 & n6721 ;
  assign n6723 = n6597 & ~n6721 ;
  assign n6724 = ~n6722 & ~n6723 ;
  assign n6725 = n6713 & n6724 ;
  assign n6726 = ~n6718 & ~n6725 ;
  assign n6727 = \core_dag_ilm2reg_M_reg[13]/NET0131  & ~n6726 ;
  assign n6593 = \core_dag_ilm2reg_I_reg[0]/NET0131  & n6592 ;
  assign n6728 = ~\core_dag_ilm2reg_L_reg[13]/NET0131  & ~n6605 ;
  assign n6729 = \core_dag_ilm2reg_L_reg[13]/NET0131  & ~\core_dag_ilm2reg_M_reg[13]/NET0131  ;
  assign n6730 = ~n6728 & ~n6729 ;
  assign n6731 = ~n6644 & ~n6645 ;
  assign n6732 = ~\core_dag_ilm2reg_L_reg[7]/NET0131  & ~\core_dag_ilm2reg_M_reg[13]/NET0131  ;
  assign n6733 = \core_dag_ilm2reg_L_reg[7]/NET0131  & \core_dag_ilm2reg_M_reg[13]/NET0131  ;
  assign n6734 = ~n6732 & ~n6733 ;
  assign n6735 = n6731 & ~n6734 ;
  assign n6736 = ~n6731 & n6734 ;
  assign n6737 = ~n6735 & ~n6736 ;
  assign n6738 = ~\core_dag_ilm2reg_L_reg[6]/NET0131  & ~\core_dag_ilm2reg_M_reg[13]/NET0131  ;
  assign n6739 = \core_dag_ilm2reg_L_reg[6]/NET0131  & \core_dag_ilm2reg_M_reg[13]/NET0131  ;
  assign n6740 = ~n6738 & ~n6739 ;
  assign n6741 = ~n6649 & ~n6740 ;
  assign n6742 = ~n6650 & ~n6741 ;
  assign n6743 = ~n6737 & n6742 ;
  assign n6744 = ~\core_dag_ilm2reg_L_reg[5]/NET0131  & ~\core_dag_ilm2reg_M_reg[13]/NET0131  ;
  assign n6745 = \core_dag_ilm2reg_L_reg[5]/NET0131  & \core_dag_ilm2reg_M_reg[13]/NET0131  ;
  assign n6746 = ~n6744 & ~n6745 ;
  assign n6747 = ~n6682 & ~n6746 ;
  assign n6748 = ~n6689 & ~n6747 ;
  assign n6749 = ~n6649 & ~n6650 ;
  assign n6750 = n6740 & ~n6749 ;
  assign n6751 = ~n6740 & n6749 ;
  assign n6752 = ~n6750 & ~n6751 ;
  assign n6753 = n6748 & ~n6752 ;
  assign n6754 = ~\core_dag_ilm2reg_L_reg[4]/NET0131  & ~\core_dag_ilm2reg_M_reg[13]/NET0131  ;
  assign n6755 = \core_dag_ilm2reg_L_reg[4]/NET0131  & \core_dag_ilm2reg_M_reg[13]/NET0131  ;
  assign n6756 = ~n6754 & ~n6755 ;
  assign n6757 = ~n6686 & ~n6756 ;
  assign n6758 = ~n6690 & ~n6757 ;
  assign n6759 = ~n6682 & ~n6689 ;
  assign n6760 = n6746 & ~n6759 ;
  assign n6761 = ~n6746 & n6759 ;
  assign n6762 = ~n6760 & ~n6761 ;
  assign n6763 = ~n6758 & n6762 ;
  assign n6764 = n6758 & ~n6762 ;
  assign n6765 = ~\core_dag_ilm2reg_L_reg[3]/NET0131  & ~\core_dag_ilm2reg_M_reg[13]/NET0131  ;
  assign n6766 = \core_dag_ilm2reg_L_reg[3]/NET0131  & \core_dag_ilm2reg_M_reg[13]/NET0131  ;
  assign n6767 = ~n6765 & ~n6766 ;
  assign n6768 = ~n6655 & ~n6767 ;
  assign n6769 = ~n6656 & ~n6768 ;
  assign n6770 = ~n6686 & ~n6690 ;
  assign n6771 = n6756 & ~n6770 ;
  assign n6772 = ~n6756 & n6770 ;
  assign n6773 = ~n6771 & ~n6772 ;
  assign n6774 = ~n6769 & n6773 ;
  assign n6775 = ~n6764 & n6774 ;
  assign n6776 = ~n6763 & ~n6775 ;
  assign n6777 = ~n6753 & ~n6776 ;
  assign n6778 = ~n6748 & n6752 ;
  assign n6779 = n6737 & ~n6742 ;
  assign n6780 = ~n6778 & ~n6779 ;
  assign n6781 = ~n6777 & n6780 ;
  assign n6782 = ~n6743 & ~n6781 ;
  assign n6783 = ~\core_dag_ilm2reg_L_reg[2]/NET0131  & ~\core_dag_ilm2reg_M_reg[13]/NET0131  ;
  assign n6784 = \core_dag_ilm2reg_L_reg[2]/NET0131  & \core_dag_ilm2reg_M_reg[13]/NET0131  ;
  assign n6785 = ~n6783 & ~n6784 ;
  assign n6786 = ~n6662 & ~n6785 ;
  assign n6787 = ~n6663 & ~n6786 ;
  assign n6788 = ~n6655 & ~n6656 ;
  assign n6789 = n6767 & ~n6788 ;
  assign n6790 = ~n6767 & n6788 ;
  assign n6791 = ~n6789 & ~n6790 ;
  assign n6792 = n6787 & ~n6791 ;
  assign n6793 = ~n6787 & n6791 ;
  assign n6794 = ~\core_dag_ilm2reg_L_reg[1]/NET0131  & ~\core_dag_ilm2reg_M_reg[13]/NET0131  ;
  assign n6795 = \core_dag_ilm2reg_L_reg[1]/NET0131  & \core_dag_ilm2reg_M_reg[13]/NET0131  ;
  assign n6796 = ~n6794 & ~n6795 ;
  assign n6797 = ~n6668 & ~n6796 ;
  assign n6798 = ~n6669 & ~n6797 ;
  assign n6799 = ~n6662 & ~n6663 ;
  assign n6800 = n6785 & ~n6799 ;
  assign n6801 = ~n6785 & n6799 ;
  assign n6802 = ~n6800 & ~n6801 ;
  assign n6803 = n6798 & ~n6802 ;
  assign n6804 = ~n6798 & n6802 ;
  assign n6805 = ~n6596 & n6721 ;
  assign n6806 = ~n6595 & ~n6805 ;
  assign n6807 = ~n6668 & ~n6669 ;
  assign n6808 = n6796 & ~n6807 ;
  assign n6809 = ~n6796 & n6807 ;
  assign n6810 = ~n6808 & ~n6809 ;
  assign n6811 = ~n6806 & ~n6810 ;
  assign n6812 = n6806 & n6810 ;
  assign n6813 = ~\core_dag_ilm2reg_M_reg[13]/NET0131  & n6724 ;
  assign n6814 = ~n6812 & ~n6813 ;
  assign n6815 = ~n6811 & ~n6814 ;
  assign n6816 = ~n6804 & ~n6815 ;
  assign n6817 = ~n6803 & ~n6816 ;
  assign n6818 = ~n6793 & ~n6817 ;
  assign n6819 = ~n6792 & ~n6818 ;
  assign n6820 = n6769 & ~n6773 ;
  assign n6821 = ~n6764 & ~n6820 ;
  assign n6822 = ~n6743 & n6821 ;
  assign n6823 = ~n6753 & n6822 ;
  assign n6824 = n6819 & n6823 ;
  assign n6825 = ~n6782 & ~n6824 ;
  assign n6826 = ~n6632 & ~n6704 ;
  assign n6827 = ~\core_dag_ilm2reg_L_reg[9]/NET0131  & ~\core_dag_ilm2reg_M_reg[13]/NET0131  ;
  assign n6828 = \core_dag_ilm2reg_L_reg[9]/NET0131  & \core_dag_ilm2reg_M_reg[13]/NET0131  ;
  assign n6829 = ~n6827 & ~n6828 ;
  assign n6830 = n6826 & ~n6829 ;
  assign n6831 = ~n6826 & n6829 ;
  assign n6832 = ~n6830 & ~n6831 ;
  assign n6833 = ~\core_dag_ilm2reg_L_reg[8]/NET0131  & ~\core_dag_ilm2reg_M_reg[13]/NET0131  ;
  assign n6834 = \core_dag_ilm2reg_L_reg[8]/NET0131  & \core_dag_ilm2reg_M_reg[13]/NET0131  ;
  assign n6835 = ~n6833 & ~n6834 ;
  assign n6836 = ~n6637 & ~n6835 ;
  assign n6837 = ~n6703 & ~n6836 ;
  assign n6838 = ~n6832 & n6837 ;
  assign n6839 = ~n6644 & ~n6734 ;
  assign n6840 = ~n6645 & ~n6839 ;
  assign n6841 = ~n6637 & ~n6703 ;
  assign n6842 = n6835 & ~n6841 ;
  assign n6843 = ~n6835 & n6841 ;
  assign n6844 = ~n6842 & ~n6843 ;
  assign n6845 = n6840 & ~n6844 ;
  assign n6846 = ~n6838 & ~n6845 ;
  assign n6847 = ~n6825 & n6846 ;
  assign n6848 = ~n6632 & ~n6829 ;
  assign n6849 = ~n6704 & ~n6848 ;
  assign n6850 = ~n6622 & ~n6702 ;
  assign n6851 = ~\core_dag_ilm2reg_L_reg[10]/NET0131  & ~\core_dag_ilm2reg_M_reg[13]/NET0131  ;
  assign n6852 = \core_dag_ilm2reg_L_reg[10]/NET0131  & \core_dag_ilm2reg_M_reg[13]/NET0131  ;
  assign n6853 = ~n6851 & ~n6852 ;
  assign n6854 = n6850 & ~n6853 ;
  assign n6855 = ~n6850 & n6853 ;
  assign n6856 = ~n6854 & ~n6855 ;
  assign n6857 = n6849 & ~n6856 ;
  assign n6858 = ~n6622 & ~n6853 ;
  assign n6859 = ~n6702 & ~n6858 ;
  assign n6860 = ~n6626 & ~n6701 ;
  assign n6861 = ~\core_dag_ilm2reg_L_reg[11]/NET0131  & ~\core_dag_ilm2reg_M_reg[13]/NET0131  ;
  assign n6862 = \core_dag_ilm2reg_L_reg[11]/NET0131  & \core_dag_ilm2reg_M_reg[13]/NET0131  ;
  assign n6863 = ~n6861 & ~n6862 ;
  assign n6864 = n6860 & ~n6863 ;
  assign n6865 = ~n6860 & n6863 ;
  assign n6866 = ~n6864 & ~n6865 ;
  assign n6867 = n6859 & ~n6866 ;
  assign n6868 = ~n6857 & ~n6867 ;
  assign n6869 = n6847 & n6868 ;
  assign n6872 = n6832 & ~n6837 ;
  assign n6873 = ~n6840 & n6844 ;
  assign n6874 = ~n6838 & n6873 ;
  assign n6875 = ~n6872 & ~n6874 ;
  assign n6876 = n6868 & ~n6875 ;
  assign n6870 = ~n6849 & n6856 ;
  assign n6871 = ~n6867 & n6870 ;
  assign n6877 = ~n6859 & n6866 ;
  assign n6878 = ~n6871 & ~n6877 ;
  assign n6879 = ~n6876 & n6878 ;
  assign n6880 = ~n6869 & n6879 ;
  assign n6881 = \core_dag_ilm2reg_L_reg[13]/NET0131  & n6605 ;
  assign n6882 = ~n6728 & ~n6881 ;
  assign n6883 = ~\core_dag_ilm2reg_L_reg[12]/NET0131  & ~\core_dag_ilm2reg_M_reg[13]/NET0131  ;
  assign n6884 = \core_dag_ilm2reg_L_reg[12]/NET0131  & \core_dag_ilm2reg_M_reg[13]/NET0131  ;
  assign n6885 = ~n6883 & ~n6884 ;
  assign n6886 = ~n6615 & n6885 ;
  assign n6887 = ~n6616 & ~n6886 ;
  assign n6888 = n6882 & ~n6887 ;
  assign n6889 = ~n6626 & ~n6863 ;
  assign n6890 = ~n6701 & ~n6889 ;
  assign n6891 = ~n6615 & ~n6616 ;
  assign n6892 = ~n6885 & n6891 ;
  assign n6893 = n6885 & ~n6891 ;
  assign n6894 = ~n6892 & ~n6893 ;
  assign n6895 = n6890 & ~n6894 ;
  assign n6896 = ~n6888 & ~n6895 ;
  assign n6897 = ~n6880 & n6896 ;
  assign n6898 = ~n6882 & n6887 ;
  assign n6899 = ~n6890 & n6894 ;
  assign n6900 = ~n6888 & n6899 ;
  assign n6901 = ~n6898 & ~n6900 ;
  assign n6902 = ~n6897 & n6901 ;
  assign n6903 = ~n6730 & n6902 ;
  assign n6904 = n6730 & ~n6902 ;
  assign n6905 = ~n6903 & ~n6904 ;
  assign n6907 = ~n6597 & ~n6905 ;
  assign n6906 = n6724 & n6905 ;
  assign n6908 = ~\core_dag_ilm2reg_M_reg[13]/NET0131  & ~n6906 ;
  assign n6909 = ~n6907 & n6908 ;
  assign n6910 = ~n6593 & ~n6909 ;
  assign n6911 = ~n6727 & n6910 ;
  assign n6912 = n6135 & ~n6911 ;
  assign n6913 = n5066 & ~n5718 ;
  assign n6915 = n5728 & ~n5729 ;
  assign n6914 = ~\bdma_BCTL_reg[1]/NET0131  & ~\bdma_DM_2nd_reg/NET0131  ;
  assign n6916 = ~\bdma_BCTL_reg[2]/NET0131  & ~n6914 ;
  assign n6917 = n6915 & n6916 ;
  assign n6918 = n6913 & n6917 ;
  assign n6919 = ~\bdma_BCTL_reg[1]/NET0131  & \bdma_DM_2nd_reg/NET0131  ;
  assign n6920 = \bdma_BCTL_reg[2]/NET0131  & ~n6919 ;
  assign n6921 = n6915 & n6920 ;
  assign n6922 = n5066 & n6921 ;
  assign n6923 = ~n5718 & n6922 ;
  assign n6924 = ~n6918 & ~n6923 ;
  assign n6958 = n5964 & n5990 ;
  assign n6959 = \core_dag_ilm2reg_I4_we_DO_reg[0]/NET0131  & n6958 ;
  assign n6960 = n6000 & n6002 ;
  assign n6961 = \core_dag_ilm2reg_I7_we_DO_reg[0]/NET0131  & n6960 ;
  assign n6966 = ~n6959 & ~n6961 ;
  assign n6962 = n6008 & n6009 ;
  assign n6963 = \core_dag_ilm2reg_I6_we_DO_reg[0]/NET0131  & n6962 ;
  assign n6964 = n6015 & n6016 ;
  assign n6965 = \core_dag_ilm2reg_I5_we_DO_reg[0]/NET0131  & n6964 ;
  assign n6967 = ~n6963 & ~n6965 ;
  assign n6968 = n6966 & n6967 ;
  assign n6969 = ~n4055 & n6968 ;
  assign n6970 = n6015 & n6043 ;
  assign n6971 = \core_dag_ilm2reg_I5_we_DO_reg[0]/NET0131  & n6970 ;
  assign n6972 = n6000 & n6039 ;
  assign n6973 = \core_dag_ilm2reg_I7_we_DO_reg[0]/NET0131  & n6972 ;
  assign n6978 = ~n6971 & ~n6973 ;
  assign n6974 = n6008 & n6041 ;
  assign n6975 = \core_dag_ilm2reg_I6_we_DO_reg[0]/NET0131  & n6974 ;
  assign n6976 = n5964 & n6037 ;
  assign n6977 = \core_dag_ilm2reg_I4_we_DO_reg[0]/NET0131  & n6976 ;
  assign n6979 = ~n6975 & ~n6977 ;
  assign n6980 = n6978 & n6979 ;
  assign n6981 = n4055 & n6980 ;
  assign n6982 = ~n6969 & ~n6981 ;
  assign n6983 = ~n6121 & n6982 ;
  assign n6936 = \core_dag_ilm1reg_I0_we_DO_reg[0]/NET0131  & n6058 ;
  assign n6937 = n6060 & n6936 ;
  assign n6941 = ~n4055 & ~n6937 ;
  assign n6940 = \core_dag_ilm1reg_I1_we_DO_reg[0]/NET0131  & n6142 ;
  assign n6938 = \core_dag_ilm1reg_I2_we_DO_reg[0]/NET0131  & n6138 ;
  assign n6939 = \core_dag_ilm1reg_I3_we_DO_reg[0]/NET0131  & n6140 ;
  assign n6942 = ~n6938 & ~n6939 ;
  assign n6943 = ~n6940 & n6942 ;
  assign n6944 = n6941 & n6943 ;
  assign n6945 = n6093 & n6936 ;
  assign n6946 = \core_dag_ilm1reg_I2_we_DO_reg[0]/NET0131  & n6152 ;
  assign n6949 = ~n6945 & ~n6946 ;
  assign n6947 = \core_dag_ilm1reg_I3_we_DO_reg[0]/NET0131  & n6150 ;
  assign n6948 = \core_dag_ilm1reg_I1_we_DO_reg[0]/NET0131  & n6154 ;
  assign n6950 = ~n6947 & ~n6948 ;
  assign n6951 = n6949 & n6950 ;
  assign n6952 = n4055 & n6951 ;
  assign n6953 = ~n6944 & ~n6952 ;
  assign n6954 = ~n6111 & n6953 ;
  assign n6955 = \core_c_dec_IR_reg[21]/NET0131  & \core_c_dec_IR_reg[22]/NET0131  ;
  assign n6956 = ~\core_c_dec_IR_reg[23]/NET0131  & n6955 ;
  assign n6957 = \core_c_dec_IR_reg[4]/NET0131  & n6956 ;
  assign n6984 = ~n6954 & ~n6957 ;
  assign n6985 = ~n6983 & n6984 ;
  assign n6986 = n5949 & ~n6985 ;
  assign n6928 = ~\core_c_dec_EXIT_E_reg/P0001  & \core_c_psq_PCS_reg[6]/NET0131  ;
  assign n6929 = ~\core_c_psq_PCS_reg[5]/NET0131  & ~n6928 ;
  assign n6930 = n5715 & n6929 ;
  assign n6931 = ~\core_c_dec_Dummy_E_reg/NET0131  & ~n4117 ;
  assign n6932 = ~n4099 & n5946 ;
  assign n6933 = n6931 & n6932 ;
  assign n6934 = n6930 & ~n6933 ;
  assign n6935 = \core_dag_ilm1reg_DMA_pi_DO_reg[0]/NET0131  & ~n6934 ;
  assign n6925 = \idma_DCTL_reg[14]/NET0131  & n5068 ;
  assign n6926 = ~n5717 & n6925 ;
  assign n6927 = \idma_DCTL_reg[0]/NET0131  & n6926 ;
  assign n6987 = ~\auctl_STEAL_reg/NET0131  & \core_c_psq_PCS_reg[7]/NET0131  ;
  assign n6988 = \memc_STI_Cg_reg/NET0131  & n6987 ;
  assign n6989 = \core_dag_ilm1reg_STAC_pi_DO_reg[0]/NET0131  & n6988 ;
  assign n6990 = ~n6927 & ~n6989 ;
  assign n6991 = ~n6935 & n6990 ;
  assign n6992 = ~n6986 & n6991 ;
  assign n6993 = n6924 & ~n6992 ;
  assign n6994 = \bdma_BIAD_reg[0]/NET0131  & ~n6924 ;
  assign n6995 = ~n6993 & ~n6994 ;
  assign n6996 = ~n6135 & ~n6995 ;
  assign n6997 = ~n6176 & ~n6996 ;
  assign n6998 = ~n6912 & n6997 ;
  assign n6999 = ~n6549 & ~n6998 ;
  assign n7000 = ~n6106 & n6112 ;
  assign n7001 = n6105 & ~n7000 ;
  assign n7002 = ~n6167 & n7001 ;
  assign n7003 = ~n5936 & ~n7002 ;
  assign n7004 = n6049 & n6172 ;
  assign n7005 = ~n7003 & ~n7004 ;
  assign n7006 = ~n6999 & ~n7005 ;
  assign n7009 = ~\memc_DMo_oe1_reg/P0001  & ~\memc_DMo_oe2_reg/P0001  ;
  assign n7010 = ~\memc_DMo_oe4_reg/P0001  & ~\memc_DMo_oe5_reg/P0001  ;
  assign n7011 = ~\memc_DMo_oe3_reg/P0001  & ~\memc_DMo_oe6_reg/P0001  ;
  assign n7012 = n7010 & n7011 ;
  assign n7013 = n7009 & n7012 ;
  assign n7014 = ~\memc_DMo_oe0_reg/P0001  & n7013 ;
  assign n7033 = ~\memc_DM_oe_reg/P0001  & \memc_DMo_oe7_reg/P0001  ;
  assign n7034 = n7014 & n7033 ;
  assign n7015 = \memc_DM_oe_reg/P0001  & ~\memc_DMo_oe7_reg/P0001  ;
  assign n7016 = n7014 & n7015 ;
  assign n7018 = ~\memc_DM_oe_reg/P0001  & ~\memc_DMo_oe7_reg/P0001  ;
  assign n7019 = ~\memc_DMo_oe0_reg/P0001  & n7018 ;
  assign n7024 = n7009 & n7019 ;
  assign n7025 = ~\memc_DMo_oe3_reg/P0001  & n7024 ;
  assign n7030 = \memc_DMo_oe6_reg/P0001  & n7010 ;
  assign n7031 = n7025 & n7030 ;
  assign n7046 = ~n7016 & ~n7031 ;
  assign n7047 = ~n7034 & n7046 ;
  assign n7026 = ~\memc_DMo_oe6_reg/P0001  & n7025 ;
  assign n7042 = ~\memc_DMo_oe4_reg/P0001  & \memc_DMo_oe5_reg/P0001  ;
  assign n7043 = n7026 & n7042 ;
  assign n7027 = \memc_DMo_oe4_reg/P0001  & ~\memc_DMo_oe5_reg/P0001  ;
  assign n7028 = n7026 & n7027 ;
  assign n7020 = n7012 & n7019 ;
  assign n7040 = ~\memc_DMo_oe1_reg/P0001  & \memc_DMo_oe2_reg/P0001  ;
  assign n7041 = n7020 & n7040 ;
  assign n7021 = \memc_DMo_oe1_reg/P0001  & ~\memc_DMo_oe2_reg/P0001  ;
  assign n7022 = n7020 & n7021 ;
  assign n7036 = \memc_DMo_oe3_reg/P0001  & ~\memc_DMo_oe6_reg/P0001  ;
  assign n7037 = n7010 & n7036 ;
  assign n7038 = n7024 & n7037 ;
  assign n7044 = ~n7022 & ~n7038 ;
  assign n7045 = ~n7041 & n7044 ;
  assign n7048 = ~n7028 & n7045 ;
  assign n7049 = ~n7043 & n7048 ;
  assign n7050 = n7047 & n7049 ;
  assign n7051 = \memc_DMo_oe0_reg/P0001  & n7018 ;
  assign n7052 = n7013 & n7051 ;
  assign n7053 = ~n7050 & ~n7052 ;
  assign n7054 = \DM_rd0[13]_pad  & ~n7053 ;
  assign n7017 = \DM_rdm[13]_pad  & n7016 ;
  assign n7032 = \DM_rd6[13]_pad  & n7031 ;
  assign n7060 = ~n7017 & ~n7032 ;
  assign n7035 = \DM_rd7[13]_pad  & n7034 ;
  assign n7057 = n7010 & n7026 ;
  assign n7061 = ~n7035 & ~n7057 ;
  assign n7062 = n7060 & n7061 ;
  assign n7055 = \DM_rd5[13]_pad  & n7043 ;
  assign n7029 = \DM_rd4[13]_pad  & n7028 ;
  assign n7056 = \DM_rd2[13]_pad  & n7041 ;
  assign n7023 = \DM_rd1[13]_pad  & n7022 ;
  assign n7039 = \DM_rd3[13]_pad  & n7038 ;
  assign n7058 = ~n7023 & ~n7039 ;
  assign n7059 = ~n7056 & n7058 ;
  assign n7063 = ~n7029 & n7059 ;
  assign n7064 = ~n7055 & n7063 ;
  assign n7065 = n7062 & n7064 ;
  assign n7066 = ~n7054 & n7065 ;
  assign n7067 = \regout_STD_C_reg[13]/P0001  & n6988 ;
  assign n7225 = ~\core_dag_ilm1reg_DMA_pi_DO_reg[2]/NET0131  & \memc_selMIO_E_reg/P0001  ;
  assign n7226 = \core_dag_ilm1reg_DMA_pi_DO_reg[0]/NET0131  & \core_dag_ilm1reg_DMA_pi_DO_reg[1]/NET0131  ;
  assign n7227 = n7225 & n7226 ;
  assign n7228 = ~\core_dag_ilm1reg_DMA_pi_DO_reg[3]/NET0131  & ~\core_dag_ilm1reg_DMA_pi_DO_reg[4]/NET0131  ;
  assign n7229 = n5944 & n7228 ;
  assign n7230 = n7227 & n7229 ;
  assign n7231 = \bdma_BCTL_reg[13]/NET0131  & n7230 ;
  assign n7236 = \core_dag_ilm1reg_DMA_pi_DO_reg[3]/NET0131  & \core_dag_ilm1reg_DMA_pi_DO_reg[4]/NET0131  ;
  assign n7241 = \core_dag_ilm1reg_DMA_pi_DO_reg[1]/NET0131  & \core_dag_ilm1reg_DMA_pi_DO_reg[2]/NET0131  ;
  assign n7242 = ~\core_dag_ilm1reg_DMA_pi_DO_reg[0]/NET0131  & \memc_selMIO_E_reg/P0001  ;
  assign n7243 = n7241 & n7242 ;
  assign n7251 = n7236 & n7243 ;
  assign n7252 = \emc_WSCRreg_DO_reg[13]/NET0131  & n7251 ;
  assign n7246 = ~\core_dag_ilm1reg_DMA_pi_DO_reg[3]/NET0131  & \core_dag_ilm1reg_DMA_pi_DO_reg[4]/NET0131  ;
  assign n7253 = \core_dag_ilm1reg_DMA_pi_DO_reg[0]/NET0131  & \memc_selMIO_E_reg/P0001  ;
  assign n7254 = ~\core_dag_ilm1reg_DMA_pi_DO_reg[1]/NET0131  & \core_dag_ilm1reg_DMA_pi_DO_reg[2]/NET0131  ;
  assign n7255 = n7253 & n7254 ;
  assign n7256 = n7246 & n7255 ;
  assign n7257 = \sport0_regs_SCLKDIVreg_DO_reg[13]/NET0131  & n7256 ;
  assign n7307 = ~n7252 & ~n7257 ;
  assign n7258 = n7242 & n7254 ;
  assign n7259 = n7246 & n7258 ;
  assign n7260 = \sport0_regs_FSDIVreg_DO_reg[13]/NET0131  & n7259 ;
  assign n7261 = ~\core_dag_ilm1reg_DMA_pi_DO_reg[0]/NET0131  & ~\core_dag_ilm1reg_DMA_pi_DO_reg[1]/NET0131  ;
  assign n7262 = n7225 & n7261 ;
  assign n7263 = n7236 & n7262 ;
  assign n7264 = ~\sport1_regs_MWORDreg_DO_reg[8]/NET0131  & ~\sport1_regs_MWORDreg_DO_reg[9]/NET0131  ;
  assign n7265 = \sport1_regs_MWORDreg_DO_reg[9]/NET0131  & ~\sport1_rxctl_SLOT1_EXT_reg[3]/NET0131  ;
  assign n7266 = ~n7264 & ~n7265 ;
  assign n7267 = n7263 & n7266 ;
  assign n7308 = ~n7260 & ~n7267 ;
  assign n7317 = n7307 & n7308 ;
  assign n7237 = ~\core_dag_ilm1reg_DMA_pi_DO_reg[0]/NET0131  & \core_dag_ilm1reg_DMA_pi_DO_reg[1]/NET0131  ;
  assign n7238 = n7225 & n7237 ;
  assign n7239 = n7236 & n7238 ;
  assign n7240 = \clkc_ckr_reg_DO_reg[13]/NET0131  & n7239 ;
  assign n7244 = n7228 & n7243 ;
  assign n7245 = \PIO_oe[9]_pad  & n7244 ;
  assign n7305 = ~n7240 & ~n7245 ;
  assign n7232 = \core_dag_ilm1reg_DMA_pi_DO_reg[0]/NET0131  & ~\core_dag_ilm1reg_DMA_pi_DO_reg[1]/NET0131  ;
  assign n7233 = n7225 & n7232 ;
  assign n7247 = n7233 & n7246 ;
  assign n7248 = \sport1_regs_SCLKDIVreg_DO_reg[13]/NET0131  & n7247 ;
  assign n7249 = n7243 & n7246 ;
  assign n7250 = \sport0_regs_SCTLreg_DO_reg[13]/NET0131  & n7249 ;
  assign n7306 = ~n7248 & ~n7250 ;
  assign n7318 = n7305 & n7306 ;
  assign n7319 = n7317 & n7318 ;
  assign n7322 = ~n7231 & n7319 ;
  assign n7234 = n7229 & n7233 ;
  assign n7235 = \bdma_BIAD_reg[13]/NET0131  & n7234 ;
  assign n7303 = n7229 & n7238 ;
  assign n7304 = \bdma_BEAD_reg[13]/NET0131  & n7303 ;
  assign n7323 = ~n7235 & ~n7304 ;
  assign n7324 = n7322 & n7323 ;
  assign n7283 = \core_dag_ilm1reg_DMA_pi_DO_reg[2]/NET0131  & ~\core_dag_ilm1reg_DMA_pi_DO_reg[3]/NET0131  ;
  assign n7284 = n7261 & n7283 ;
  assign n7285 = ~\core_dag_ilm1reg_DMA_pi_DO_reg[4]/NET0131  & n5944 ;
  assign n7286 = \memc_selMIO_E_reg/P0001  & n7285 ;
  assign n7287 = n7284 & n7286 ;
  assign n7288 = \bdma_BWCOUNT_reg[13]/NET0131  & n7287 ;
  assign n7275 = n7241 & n7253 ;
  assign n7301 = n7236 & n7275 ;
  assign n7302 = \memc_usysr_DO_reg[13]/NET0131  & n7301 ;
  assign n7297 = n7228 & n7275 ;
  assign n7298 = \pio_pmask_reg_DO_reg[9]/NET0131  & n7297 ;
  assign n7299 = n7228 & n7262 ;
  assign n7300 = \idma_DCTL_reg[13]/NET0131  & n7299 ;
  assign n7313 = ~n7298 & ~n7300 ;
  assign n7314 = ~n7302 & n7313 ;
  assign n7289 = n7236 & n7258 ;
  assign n7290 = \tm_TCR_TMP_reg[13]/NET0131  & n7289 ;
  assign n7291 = n7228 & n7255 ;
  assign n7292 = \PIO_out[9]_pad  & n7291 ;
  assign n7311 = ~n7290 & ~n7292 ;
  assign n7293 = n7236 & n7255 ;
  assign n7294 = \tm_tpr_reg_DO_reg[13]/NET0131  & n7293 ;
  assign n7295 = n7227 & n7246 ;
  assign n7296 = \sport0_regs_AUTO_a_reg[13]/NET0131  & n7295 ;
  assign n7312 = ~n7294 & ~n7296 ;
  assign n7315 = n7311 & n7312 ;
  assign n7268 = ~\core_dag_ilm1reg_DMA_pi_DO_reg[4]/NET0131  & \memc_selMIO_E_reg/P0001  ;
  assign n7269 = ~\core_dag_ilm1reg_DMA_pi_DO_reg[2]/NET0131  & \core_dag_ilm1reg_DMA_pi_DO_reg[3]/NET0131  ;
  assign n7270 = n7261 & n7269 ;
  assign n7271 = n7268 & n7270 ;
  assign n7272 = \pio_PINT_reg[9]/NET0131  & n7271 ;
  assign n7273 = n7246 & n7262 ;
  assign n7274 = \sport1_regs_FSDIVreg_DO_reg[13]/NET0131  & n7273 ;
  assign n7309 = ~n7272 & ~n7274 ;
  assign n7276 = n7246 & n7275 ;
  assign n7277 = ~\sport0_regs_MWORDreg_DO_reg[8]/NET0131  & ~\sport0_regs_MWORDreg_DO_reg[9]/NET0131  ;
  assign n7278 = \sport0_regs_MWORDreg_DO_reg[9]/NET0131  & ~\sport0_rxctl_SLOT1_EXT_reg[3]/NET0131  ;
  assign n7279 = ~n7277 & ~n7278 ;
  assign n7280 = n7276 & n7279 ;
  assign n7281 = n7238 & n7246 ;
  assign n7282 = \sport1_regs_SCTLreg_DO_reg[13]/NET0131  & n7281 ;
  assign n7310 = ~n7280 & ~n7282 ;
  assign n7316 = n7309 & n7310 ;
  assign n7320 = n7315 & n7316 ;
  assign n7321 = n7314 & n7320 ;
  assign n7325 = ~n7288 & n7321 ;
  assign n7326 = n7324 & n7325 ;
  assign n7327 = \memc_ldSREG_E_reg/NET0131  & ~n7326 ;
  assign n7215 = \core_c_dec_MFPSQ_Ei_reg/NET0131  & ~n6988 ;
  assign n7220 = \core_c_dec_MFtoppcs_Eg_reg/P0001  & ~n4489 ;
  assign n7216 = ~\core_c_dec_imm14_E_reg/P0001  & ~\core_c_dec_imm16_E_reg/P0001  ;
  assign n7217 = \core_c_dec_IRE_reg[17]/NET0131  & ~n7216 ;
  assign n7218 = \core_c_dec_MFCNTR_E_reg/P0001  & \core_c_psq_CNTR_reg_DO_reg[13]/NET0131  ;
  assign n7219 = \core_c_dec_MFIDR_E_reg/P0001  & \sice_idr1_reg_DO_reg[1]/P0001  ;
  assign n7221 = ~n7218 & ~n7219 ;
  assign n7222 = ~n7217 & n7221 ;
  assign n7223 = ~n7220 & n7222 ;
  assign n7224 = n7215 & ~n7223 ;
  assign n7128 = \core_c_dec_MFDAG2_Ei_reg/NET0131  & ~n6988 ;
  assign n7131 = \core_c_dec_MFMreg_E_reg[4]/P0001  & \core_dag_ilm2reg_M4_we_DO_reg[13]/NET0131  ;
  assign n7132 = \core_c_dec_MFMreg_E_reg[5]/P0001  & \core_dag_ilm2reg_M5_we_DO_reg[13]/NET0131  ;
  assign n7135 = ~n7131 & ~n7132 ;
  assign n7133 = \core_c_dec_MFMreg_E_reg[6]/P0001  & \core_dag_ilm2reg_M6_we_DO_reg[13]/NET0131  ;
  assign n7134 = \core_c_dec_MFMreg_E_reg[7]/P0001  & \core_dag_ilm2reg_M7_we_DO_reg[13]/NET0131  ;
  assign n7136 = ~n7133 & ~n7134 ;
  assign n7137 = n7135 & n7136 ;
  assign n7140 = \core_c_dec_MFIreg_E_reg[5]/P0001  & \core_dag_ilm2reg_I5_we_DO_reg[13]/NET0131  ;
  assign n7141 = \core_c_dec_MFLreg_E_reg[6]/P0001  & \core_dag_ilm2reg_L6_we_DO_reg[13]/NET0131  ;
  assign n7146 = ~n7140 & ~n7141 ;
  assign n7142 = \core_c_dec_MFIreg_E_reg[7]/P0001  & \core_dag_ilm2reg_I7_we_DO_reg[13]/NET0131  ;
  assign n7143 = \core_c_dec_MFLreg_E_reg[4]/P0001  & \core_dag_ilm2reg_L4_we_DO_reg[13]/NET0131  ;
  assign n7147 = ~n7142 & ~n7143 ;
  assign n7148 = n7146 & n7147 ;
  assign n7129 = \core_c_dec_MFLreg_E_reg[7]/P0001  & \core_dag_ilm2reg_L7_we_DO_reg[13]/NET0131  ;
  assign n7130 = \core_c_dec_MFIreg_E_reg[4]/P0001  & \core_dag_ilm2reg_I4_we_DO_reg[13]/NET0131  ;
  assign n7144 = ~n7129 & ~n7130 ;
  assign n7138 = \core_c_dec_MFLreg_E_reg[5]/P0001  & \core_dag_ilm2reg_L5_we_DO_reg[13]/NET0131  ;
  assign n7139 = \core_c_dec_MFIreg_E_reg[6]/P0001  & \core_dag_ilm2reg_I6_we_DO_reg[13]/NET0131  ;
  assign n7145 = ~n7138 & ~n7139 ;
  assign n7149 = n7144 & n7145 ;
  assign n7150 = n7148 & n7149 ;
  assign n7151 = n7137 & n7150 ;
  assign n7152 = n7128 & ~n7151 ;
  assign n7068 = \core_c_dec_MFDAG1_Ei_reg/NET0131  & ~n6988 ;
  assign n7072 = \core_c_dec_MFMreg_E_reg[0]/P0001  & \core_dag_ilm1reg_M0_we_DO_reg[13]/NET0131  ;
  assign n7073 = \core_c_dec_MFMreg_E_reg[1]/P0001  & \core_dag_ilm1reg_M1_we_DO_reg[13]/NET0131  ;
  assign n7076 = ~n7072 & ~n7073 ;
  assign n7074 = \core_c_dec_MFMreg_E_reg[2]/P0001  & \core_dag_ilm1reg_M2_we_DO_reg[13]/NET0131  ;
  assign n7075 = \core_c_dec_MFMreg_E_reg[3]/P0001  & \core_dag_ilm1reg_M3_we_DO_reg[13]/NET0131  ;
  assign n7077 = ~n7074 & ~n7075 ;
  assign n7078 = n7076 & n7077 ;
  assign n7080 = \core_c_dec_MFLreg_E_reg[1]/P0001  & \core_dag_ilm1reg_L1_we_DO_reg[13]/NET0131  ;
  assign n7081 = \core_c_dec_MFIreg_E_reg[2]/P0001  & \core_dag_ilm1reg_I2_we_DO_reg[13]/NET0131  ;
  assign n7086 = ~n7080 & ~n7081 ;
  assign n7082 = \core_c_dec_MFIreg_E_reg[3]/P0001  & \core_dag_ilm1reg_I3_we_DO_reg[13]/NET0131  ;
  assign n7083 = \core_c_dec_MFLreg_E_reg[0]/P0001  & \core_dag_ilm1reg_L0_we_DO_reg[13]/NET0131  ;
  assign n7087 = ~n7082 & ~n7083 ;
  assign n7088 = n7086 & n7087 ;
  assign n7069 = \core_c_dec_MFLreg_E_reg[3]/P0001  & \core_dag_ilm1reg_L3_we_DO_reg[13]/NET0131  ;
  assign n7070 = \core_c_dec_MFIreg_E_reg[0]/P0001  & \core_dag_ilm1reg_I0_we_DO_reg[13]/NET0131  ;
  assign n7084 = ~n7069 & ~n7070 ;
  assign n7071 = \core_c_dec_MFIreg_E_reg[1]/P0001  & \core_dag_ilm1reg_I1_we_DO_reg[13]/NET0131  ;
  assign n7079 = \core_c_dec_MFLreg_E_reg[2]/P0001  & \core_dag_ilm1reg_L2_we_DO_reg[13]/NET0131  ;
  assign n7085 = ~n7071 & ~n7079 ;
  assign n7089 = n7084 & n7085 ;
  assign n7090 = n7088 & n7089 ;
  assign n7091 = n7078 & n7090 ;
  assign n7092 = n7068 & ~n7091 ;
  assign n7119 = \core_c_dec_MFSPT_Ei_reg/NET0131  & ~n6988 ;
  assign n7120 = \core_c_dec_MFTX1_E_reg/P0001  & \sport1_txctl_TX_reg[13]/P0001  ;
  assign n7121 = \core_c_dec_MFTX0_E_reg/P0001  & \sport0_txctl_TX_reg[13]/P0001  ;
  assign n7124 = ~n7120 & ~n7121 ;
  assign n7122 = \core_c_dec_MFRX1_E_reg/P0001  & \sport1_rxctl_RX_reg[13]/P0001  ;
  assign n7123 = \core_c_dec_MFRX0_E_reg/P0001  & \sport0_rxctl_RX_reg[13]/P0001  ;
  assign n7125 = ~n7122 & ~n7123 ;
  assign n7126 = n7124 & n7125 ;
  assign n7127 = n7119 & ~n7126 ;
  assign n7328 = ~n7092 & ~n7127 ;
  assign n7329 = ~n7152 & n7328 ;
  assign n7179 = \core_c_dec_MFMAC_Ei_reg/NET0131  & ~n6988 ;
  assign n7204 = ~\core_c_psq_MSTAT_reg_DO_reg[0]/P0002  & \core_eu_em_mac_em_reg_mr2rwe_DO_reg[7]/P0001  ;
  assign n7205 = \core_c_psq_MSTAT_reg_DO_reg[0]/P0002  & \core_eu_em_mac_em_reg_mr2swe_DO_reg[7]/P0001  ;
  assign n7206 = ~n7204 & ~n7205 ;
  assign n7207 = \core_c_dec_MFMR2_E_reg/P0001  & ~n7206 ;
  assign n7196 = ~\core_c_psq_MSTAT_reg_DO_reg[0]/P0002  & \core_eu_em_mac_em_reg_my0rwe_DO_reg[13]/P0001  ;
  assign n7197 = \core_c_psq_MSTAT_reg_DO_reg[0]/P0002  & \core_eu_em_mac_em_reg_my0swe_DO_reg[13]/P0001  ;
  assign n7198 = ~n7196 & ~n7197 ;
  assign n7199 = \core_c_dec_MFMY0_E_reg/P0001  & ~n7198 ;
  assign n7200 = ~\core_c_psq_MSTAT_reg_DO_reg[0]/P0002  & \core_eu_em_mac_em_reg_mr1rwe_DO_reg[13]/P0001  ;
  assign n7201 = \core_c_psq_MSTAT_reg_DO_reg[0]/P0002  & \core_eu_em_mac_em_reg_mr1swe_DO_reg[13]/P0001  ;
  assign n7202 = ~n7200 & ~n7201 ;
  assign n7203 = \core_c_dec_MFMR1_E_reg/P0001  & ~n7202 ;
  assign n7210 = ~n7199 & ~n7203 ;
  assign n7211 = ~n7207 & n7210 ;
  assign n7180 = ~\core_c_psq_MSTAT_reg_DO_reg[0]/P0002  & \core_eu_em_mac_em_reg_mr0rwe_DO_reg[13]/P0001  ;
  assign n7181 = \core_c_psq_MSTAT_reg_DO_reg[0]/P0002  & \core_eu_em_mac_em_reg_mr0swe_DO_reg[13]/P0001  ;
  assign n7182 = ~n7180 & ~n7181 ;
  assign n7183 = \core_c_dec_MFMR0_E_reg/P0001  & ~n7182 ;
  assign n7184 = ~\core_c_psq_MSTAT_reg_DO_reg[0]/P0002  & \core_eu_em_mac_em_reg_mx1rwe_DO_reg[13]/P0001  ;
  assign n7185 = \core_c_psq_MSTAT_reg_DO_reg[0]/P0002  & \core_eu_em_mac_em_reg_mx1swe_DO_reg[13]/P0001  ;
  assign n7186 = ~n7184 & ~n7185 ;
  assign n7187 = \core_c_dec_MFMX1_E_reg/P0001  & ~n7186 ;
  assign n7208 = ~n7183 & ~n7187 ;
  assign n7188 = ~\core_c_psq_MSTAT_reg_DO_reg[0]/P0002  & \core_eu_em_mac_em_reg_my1rwe_DO_reg[13]/P0001  ;
  assign n7189 = \core_c_psq_MSTAT_reg_DO_reg[0]/P0002  & \core_eu_em_mac_em_reg_my1swe_DO_reg[13]/P0001  ;
  assign n7190 = ~n7188 & ~n7189 ;
  assign n7191 = \core_c_dec_MFMY1_E_reg/P0001  & ~n7190 ;
  assign n7192 = ~\core_c_psq_MSTAT_reg_DO_reg[0]/P0002  & \core_eu_em_mac_em_reg_mx0rwe_DO_reg[13]/P0001  ;
  assign n7193 = \core_c_psq_MSTAT_reg_DO_reg[0]/P0002  & \core_eu_em_mac_em_reg_mx0swe_DO_reg[13]/P0001  ;
  assign n7194 = ~n7192 & ~n7193 ;
  assign n7195 = \core_c_dec_MFMX0_E_reg/P0001  & ~n7194 ;
  assign n7209 = ~n7191 & ~n7195 ;
  assign n7212 = n7208 & n7209 ;
  assign n7213 = n7211 & n7212 ;
  assign n7214 = n7179 & ~n7213 ;
  assign n7093 = \core_c_dec_MFALU_Ei_reg/NET0131  & ~n6988 ;
  assign n7094 = ~\core_c_psq_MSTAT_reg_DO_reg[0]/P0002  & \core_eu_ea_alu_ea_reg_ax0rwe_DO_reg[13]/P0001  ;
  assign n7095 = \core_c_psq_MSTAT_reg_DO_reg[0]/P0002  & \core_eu_ea_alu_ea_reg_ax0swe_DO_reg[13]/P0001  ;
  assign n7096 = ~n7094 & ~n7095 ;
  assign n7097 = \core_c_dec_MFAX0_E_reg/P0001  & ~n7096 ;
  assign n7098 = ~\core_c_psq_MSTAT_reg_DO_reg[0]/P0002  & \core_eu_ea_alu_ea_reg_ax1rwe_DO_reg[13]/P0001  ;
  assign n7099 = \core_c_psq_MSTAT_reg_DO_reg[0]/P0002  & \core_eu_ea_alu_ea_reg_ax1swe_DO_reg[13]/P0001  ;
  assign n7100 = ~n7098 & ~n7099 ;
  assign n7101 = \core_c_dec_MFAX1_E_reg/P0001  & ~n7100 ;
  assign n7114 = ~n7097 & ~n7101 ;
  assign n7110 = ~\core_c_psq_MSTAT_reg_DO_reg[0]/P0002  & \core_eu_ea_alu_ea_reg_arrwe_DO_reg[13]/P0001  ;
  assign n7111 = \core_c_psq_MSTAT_reg_DO_reg[0]/P0002  & \core_eu_ea_alu_ea_reg_arswe_DO_reg[13]/P0001  ;
  assign n7112 = ~n7110 & ~n7111 ;
  assign n7113 = \core_c_dec_MFAR_E_reg/P0001  & ~n7112 ;
  assign n7102 = ~\core_c_psq_MSTAT_reg_DO_reg[0]/P0002  & \core_eu_ea_alu_ea_reg_ay0rwe_DO_reg[13]/P0001  ;
  assign n7103 = \core_c_psq_MSTAT_reg_DO_reg[0]/P0002  & \core_eu_ea_alu_ea_reg_ay0swe_DO_reg[13]/P0001  ;
  assign n7104 = ~n7102 & ~n7103 ;
  assign n7105 = \core_c_dec_MFAY0_E_reg/P0001  & ~n7104 ;
  assign n7106 = ~\core_c_psq_MSTAT_reg_DO_reg[0]/P0002  & \core_eu_ea_alu_ea_reg_ay1rwe_DO_reg[13]/P0001  ;
  assign n7107 = \core_c_psq_MSTAT_reg_DO_reg[0]/P0002  & \core_eu_ea_alu_ea_reg_ay1swe_DO_reg[13]/P0001  ;
  assign n7108 = ~n7106 & ~n7107 ;
  assign n7109 = \core_c_dec_MFAY1_E_reg/P0001  & ~n7108 ;
  assign n7115 = ~n7105 & ~n7109 ;
  assign n7116 = ~n7113 & n7115 ;
  assign n7117 = n7114 & n7116 ;
  assign n7118 = n7093 & ~n7117 ;
  assign n7153 = \core_c_dec_MFSHT_Ei_reg/NET0131  & ~n6988 ;
  assign n7166 = ~\core_c_psq_MSTAT_reg_DO_reg[0]/P0002  & \core_eu_es_sht_es_reg_SBr_reg[4]/P0001  ;
  assign n7167 = \core_c_psq_MSTAT_reg_DO_reg[0]/P0002  & \core_eu_es_sht_es_reg_SBs_reg[4]/P0001  ;
  assign n7168 = ~n7166 & ~n7167 ;
  assign n7169 = \core_c_dec_MFSB_E_reg/P0001  & ~n7168 ;
  assign n7170 = ~\core_c_psq_MSTAT_reg_DO_reg[0]/P0002  & \core_eu_es_sht_es_reg_serwe_DO_reg[7]/P0001  ;
  assign n7171 = \core_c_psq_MSTAT_reg_DO_reg[0]/P0002  & \core_eu_es_sht_es_reg_seswe_DO_reg[7]/P0001  ;
  assign n7172 = ~n7170 & ~n7171 ;
  assign n7173 = \core_c_dec_MFSE_E_reg/P0001  & ~n7172 ;
  assign n7174 = ~n7169 & ~n7173 ;
  assign n7162 = ~\core_c_psq_MSTAT_reg_DO_reg[0]/P0002  & \core_eu_es_sht_es_reg_sr0rwe_DO_reg[13]/P0001  ;
  assign n7163 = \core_c_psq_MSTAT_reg_DO_reg[0]/P0002  & \core_eu_es_sht_es_reg_sr0swe_DO_reg[13]/P0001  ;
  assign n7164 = ~n7162 & ~n7163 ;
  assign n7165 = \core_c_dec_MFSR0_E_reg/P0001  & ~n7164 ;
  assign n7154 = ~\core_c_psq_MSTAT_reg_DO_reg[0]/P0002  & \core_eu_es_sht_es_reg_sr1rwe_DO_reg[13]/P0001  ;
  assign n7155 = \core_c_psq_MSTAT_reg_DO_reg[0]/P0002  & \core_eu_es_sht_es_reg_sr1swe_DO_reg[13]/P0001  ;
  assign n7156 = ~n7154 & ~n7155 ;
  assign n7157 = \core_c_dec_MFSR1_E_reg/P0001  & ~n7156 ;
  assign n7158 = ~\core_c_psq_MSTAT_reg_DO_reg[0]/P0002  & \core_eu_es_sht_es_reg_sirwe_DO_reg[13]/P0001  ;
  assign n7159 = \core_c_psq_MSTAT_reg_DO_reg[0]/P0002  & \core_eu_es_sht_es_reg_siswe_DO_reg[13]/P0001  ;
  assign n7160 = ~n7158 & ~n7159 ;
  assign n7161 = \core_c_dec_MFSI_E_reg/P0001  & ~n7160 ;
  assign n7175 = ~n7157 & ~n7161 ;
  assign n7176 = ~n7165 & n7175 ;
  assign n7177 = n7174 & n7176 ;
  assign n7178 = n7153 & ~n7177 ;
  assign n7330 = ~n7118 & ~n7178 ;
  assign n7331 = ~n7214 & n7330 ;
  assign n7332 = n7329 & n7331 ;
  assign n7333 = ~n7224 & n7332 ;
  assign n7334 = ~n7327 & n7333 ;
  assign n7335 = ~n7067 & n7334 ;
  assign n7336 = ~\emc_DMDoe_reg/NET0131  & ~n7335 ;
  assign n7337 = \emc_DMDoe_reg/NET0131  & \emc_DMDreg_reg[13]/P0001  ;
  assign n7338 = n7057 & ~n7337 ;
  assign n7339 = ~n7336 & n7338 ;
  assign n7340 = ~n7066 & ~n7339 ;
  assign n7341 = ~n6135 & n7340 ;
  assign n7007 = ~n6953 & ~n6982 ;
  assign n7008 = n6135 & ~n7007 ;
  assign n7342 = ~n6176 & ~n7008 ;
  assign n7343 = ~n7341 & n7342 ;
  assign n7618 = n6365 & n6496 ;
  assign n7617 = ~n6362 & ~n6496 ;
  assign n7619 = ~\core_dag_ilm1reg_M_reg[13]/NET0131  & ~n7617 ;
  assign n7620 = ~n7618 & n7619 ;
  assign n7609 = \core_dag_ilm1reg_I_reg[0]/NET0131  & n6345 ;
  assign n7610 = n6497 & n6527 ;
  assign n7611 = n6498 & ~n6527 ;
  assign n7612 = ~n7610 & ~n7611 ;
  assign n7614 = ~n6365 & ~n7612 ;
  assign n7613 = ~n6362 & n7612 ;
  assign n7615 = \core_dag_ilm1reg_M_reg[13]/NET0131  & ~n7613 ;
  assign n7616 = ~n7614 & n7615 ;
  assign n7621 = ~n7609 & ~n7616 ;
  assign n7622 = ~n7620 & n7621 ;
  assign n7623 = ~n6135 & ~n7622 ;
  assign n7350 = \DM_rd0[0]_pad  & ~n7053 ;
  assign n7344 = \DM_rdm[0]_pad  & n7016 ;
  assign n7355 = ~n7057 & ~n7344 ;
  assign n7347 = \DM_rd6[0]_pad  & n7031 ;
  assign n7348 = \DM_rd7[0]_pad  & n7034 ;
  assign n7356 = ~n7347 & ~n7348 ;
  assign n7357 = n7355 & n7356 ;
  assign n7351 = \DM_rd4[0]_pad  & n7028 ;
  assign n7346 = \DM_rd5[0]_pad  & n7043 ;
  assign n7352 = \DM_rd2[0]_pad  & n7041 ;
  assign n7345 = \DM_rd1[0]_pad  & n7022 ;
  assign n7349 = \DM_rd3[0]_pad  & n7038 ;
  assign n7353 = ~n7345 & ~n7349 ;
  assign n7354 = ~n7352 & n7353 ;
  assign n7358 = ~n7346 & n7354 ;
  assign n7359 = ~n7351 & n7358 ;
  assign n7360 = n7357 & n7359 ;
  assign n7361 = ~n7350 & n7360 ;
  assign n7362 = \regout_STD_C_reg[0]/P0001  & n6988 ;
  assign n7523 = \bdma_BIAD_reg[0]/NET0131  & n7234 ;
  assign n7510 = \sport0_regs_SCTLreg_DO_reg[0]/NET0131  & n7249 ;
  assign n7511 = \PIO_oe[0]_pad  & n7244 ;
  assign n7548 = ~n7510 & ~n7511 ;
  assign n7512 = \sport0_regs_SCLKDIVreg_DO_reg[0]/NET0131  & n7256 ;
  assign n7513 = n7226 & n7269 ;
  assign n7514 = n7268 & n7513 ;
  assign n7515 = \emc_WSCRext_reg_DO_reg[0]/NET0131  & n7514 ;
  assign n7549 = ~n7512 & ~n7515 ;
  assign n7562 = n7548 & n7549 ;
  assign n7506 = \emc_WSCRreg_DO_reg[0]/NET0131  & n7251 ;
  assign n7521 = n7237 & n7268 ;
  assign n7522 = n7269 & n7521 ;
  assign n7546 = ~n7506 & ~n7522 ;
  assign n7507 = \sport0_regs_FSDIVreg_DO_reg[0]/NET0131  & n7259 ;
  assign n7508 = \sport1_regs_MWORDreg_DO_reg[0]/NET0131  & n7263 ;
  assign n7547 = ~n7507 & ~n7508 ;
  assign n7563 = n7546 & n7547 ;
  assign n7564 = n7562 & n7563 ;
  assign n7568 = ~n7523 & n7564 ;
  assign n7538 = \bdma_BEAD_reg[0]/NET0131  & n7303 ;
  assign n7539 = \bdma_BCTL_reg[0]/NET0131  & n7230 ;
  assign n7569 = ~n7538 & ~n7539 ;
  assign n7570 = n7568 & n7569 ;
  assign n7530 = n7232 & n7269 ;
  assign n7534 = n7286 & n7530 ;
  assign n7535 = \bdma_BOVL_reg[0]/NET0131  & n7534 ;
  assign n7509 = \bdma_BWCOUNT_reg[0]/NET0131  & n7287 ;
  assign n7520 = \tm_TCR_TMP_reg[0]/NET0131  & n7289 ;
  assign n7524 = \pio_pmask_reg_DO_reg[0]/NET0131  & n7297 ;
  assign n7552 = ~n7520 & ~n7524 ;
  assign n7525 = \core_dag_ilm1reg_DMA_pi_DO_reg[2]/NET0131  & \core_dag_ilm1reg_DMA_pi_DO_reg[3]/NET0131  ;
  assign n7526 = n7226 & n7525 ;
  assign n7527 = n7268 & n7526 ;
  assign n7528 = \sport1_regs_AUTOreg_DO_reg[0]/NET0131  & n7527 ;
  assign n7529 = \sport1_regs_SCLKDIVreg_DO_reg[0]/NET0131  & n7247 ;
  assign n7553 = ~n7528 & ~n7529 ;
  assign n7560 = n7552 & n7553 ;
  assign n7516 = \memc_usysr_DO_reg[0]/NET0131  & n7301 ;
  assign n7517 = \sport0_regs_AUTOreg_DO_reg[0]/NET0131  & n7295 ;
  assign n7550 = ~n7516 & ~n7517 ;
  assign n7518 = \idma_DCTL_reg[0]/NET0131  & n7299 ;
  assign n7519 = \pio_PINT_reg[0]/NET0131  & n7271 ;
  assign n7551 = ~n7518 & ~n7519 ;
  assign n7561 = n7550 & n7551 ;
  assign n7565 = n7560 & n7561 ;
  assign n7542 = \sport1_regs_SCTLreg_DO_reg[0]/NET0131  & n7281 ;
  assign n7543 = \clkc_ckr_reg_DO_reg[0]/NET0131  & n7239 ;
  assign n7556 = ~n7542 & ~n7543 ;
  assign n7544 = \sport0_regs_MWORDreg_DO_reg[0]/NET0131  & n7276 ;
  assign n7545 = \PIO_out[0]_pad  & n7291 ;
  assign n7557 = ~n7544 & ~n7545 ;
  assign n7558 = n7556 & n7557 ;
  assign n7531 = \core_dag_ilm1reg_DMA_pi_DO_reg[4]/NET0131  & \memc_selMIO_E_reg/P0001  ;
  assign n7532 = n7530 & n7531 ;
  assign n7533 = \idma_DOVL_reg[0]/NET0131  & n7532 ;
  assign n7536 = \tm_tpr_reg_DO_reg[0]/NET0131  & n7293 ;
  assign n7554 = ~n7533 & ~n7536 ;
  assign n7537 = \sport1_regs_FSDIVreg_DO_reg[0]/NET0131  & n7273 ;
  assign n7540 = n7227 & n7236 ;
  assign n7541 = \tm_tsr_reg_DO_reg[0]/NET0131  & n7540 ;
  assign n7555 = ~n7537 & ~n7541 ;
  assign n7559 = n7554 & n7555 ;
  assign n7566 = n7558 & n7559 ;
  assign n7567 = n7565 & n7566 ;
  assign n7571 = ~n7509 & n7567 ;
  assign n7572 = ~n7535 & n7571 ;
  assign n7573 = n7570 & n7572 ;
  assign n7574 = \memc_ldSREG_E_reg/NET0131  & ~n7573 ;
  assign n7578 = \core_c_dec_MFtoppcs_Eg_reg/P0001  & ~n4588 ;
  assign n7581 = \core_c_dec_MFDMOVL_E_reg/P0001  & \core_c_psq_DMOVL_reg_DO_reg[0]/NET0131  ;
  assign n7582 = \core_c_dec_MFIDR_E_reg/P0001  & \sice_idr0_reg_DO_reg[0]/P0001  ;
  assign n7587 = ~n7581 & ~n7582 ;
  assign n7583 = \core_c_dec_MFICNTL_E_reg/P0001  & \core_c_psq_ICNTL_reg_DO_reg[0]/NET0131  ;
  assign n7584 = \core_c_dec_MFCNTR_E_reg/P0001  & \core_c_psq_CNTR_reg_DO_reg[0]/NET0131  ;
  assign n7588 = ~n7583 & ~n7584 ;
  assign n7589 = n7587 & n7588 ;
  assign n7579 = \core_c_dec_IRE_reg[4]/NET0131  & ~n7216 ;
  assign n7575 = \core_c_dec_MFMSTAT_E_reg/P0001  & \core_c_psq_MSTAT_reg_DO_reg[0]/P0002  ;
  assign n7576 = \core_c_dec_MFIMASK_E_reg/P0001  & \core_c_psq_IMASK_reg[0]/NET0131  ;
  assign n7585 = ~n7575 & ~n7576 ;
  assign n7577 = \core_c_dec_MFSSTAT_E_reg/P0001  & \core_c_psq_SSTAT_reg[0]/NET0131  ;
  assign n7580 = \core_c_dec_MFPMOVL_E_reg/P0001  & \core_c_psq_PMOVL_regl_DO_reg[0]/NET0131  ;
  assign n7586 = ~n7577 & ~n7580 ;
  assign n7590 = n7585 & n7586 ;
  assign n7591 = ~n7579 & n7590 ;
  assign n7592 = n7589 & n7591 ;
  assign n7593 = ~n7578 & n7592 ;
  assign n7594 = n7215 & ~n7593 ;
  assign n7490 = \core_c_dec_MFLreg_E_reg[2]/P0001  & \core_dag_ilm1reg_L2_we_DO_reg[0]/NET0131  ;
  assign n7491 = \core_c_dec_MFMreg_E_reg[1]/P0001  & \core_dag_ilm1reg_M1_we_DO_reg[0]/NET0131  ;
  assign n7498 = ~n7490 & ~n7491 ;
  assign n7492 = \core_c_dec_MFMreg_E_reg[2]/P0001  & \core_dag_ilm1reg_M2_we_DO_reg[0]/NET0131  ;
  assign n7493 = \core_c_dec_MFMreg_E_reg[3]/P0001  & \core_dag_ilm1reg_M3_we_DO_reg[0]/NET0131  ;
  assign n7499 = ~n7492 & ~n7493 ;
  assign n7500 = n7498 & n7499 ;
  assign n7486 = \core_c_dec_MFLreg_E_reg[3]/P0001  & \core_dag_ilm1reg_L3_we_DO_reg[0]/NET0131  ;
  assign n7487 = \core_c_dec_MFMreg_E_reg[0]/P0001  & \core_dag_ilm1reg_M0_we_DO_reg[0]/NET0131  ;
  assign n7496 = ~n7486 & ~n7487 ;
  assign n7488 = \core_c_dec_MFIreg_E_reg[1]/P0001  & \core_dag_ilm1reg_I1_we_DO_reg[0]/NET0131  ;
  assign n7489 = \core_c_dec_MFIreg_E_reg[2]/P0001  & \core_dag_ilm1reg_I2_we_DO_reg[0]/NET0131  ;
  assign n7497 = ~n7488 & ~n7489 ;
  assign n7501 = n7496 & n7497 ;
  assign n7482 = \core_c_dec_MFIreg_E_reg[0]/P0001  & \core_dag_ilm1reg_I0_we_DO_reg[0]/NET0131  ;
  assign n7483 = \core_c_dec_MFIreg_E_reg[3]/P0001  & \core_dag_ilm1reg_I3_we_DO_reg[0]/NET0131  ;
  assign n7494 = ~n7482 & ~n7483 ;
  assign n7484 = \core_c_dec_MFLreg_E_reg[0]/P0001  & \core_dag_ilm1reg_L0_we_DO_reg[0]/NET0131  ;
  assign n7485 = \core_c_dec_MFLreg_E_reg[1]/P0001  & \core_dag_ilm1reg_L1_we_DO_reg[0]/NET0131  ;
  assign n7495 = ~n7484 & ~n7485 ;
  assign n7502 = n7494 & n7495 ;
  assign n7503 = n7501 & n7502 ;
  assign n7504 = n7500 & n7503 ;
  assign n7505 = n7068 & ~n7504 ;
  assign n7396 = \core_c_dec_MFIreg_E_reg[4]/P0001  & \core_dag_ilm2reg_I4_we_DO_reg[0]/NET0131  ;
  assign n7397 = \core_c_dec_MFIreg_E_reg[7]/P0001  & \core_dag_ilm2reg_I7_we_DO_reg[0]/NET0131  ;
  assign n7404 = ~n7396 & ~n7397 ;
  assign n7398 = \core_c_dec_MFLreg_E_reg[4]/P0001  & \core_dag_ilm2reg_L4_we_DO_reg[0]/NET0131  ;
  assign n7399 = \core_c_dec_MFLreg_E_reg[5]/P0001  & \core_dag_ilm2reg_L5_we_DO_reg[0]/NET0131  ;
  assign n7405 = ~n7398 & ~n7399 ;
  assign n7406 = n7404 & n7405 ;
  assign n7392 = \core_c_dec_MFIreg_E_reg[5]/P0001  & \core_dag_ilm2reg_I5_we_DO_reg[0]/NET0131  ;
  assign n7393 = \core_c_dec_MFIreg_E_reg[6]/P0001  & \core_dag_ilm2reg_I6_we_DO_reg[0]/NET0131  ;
  assign n7402 = ~n7392 & ~n7393 ;
  assign n7394 = \core_c_dec_MFMreg_E_reg[6]/P0001  & \core_dag_ilm2reg_M6_we_DO_reg[0]/NET0131  ;
  assign n7395 = \core_c_dec_MFMreg_E_reg[7]/P0001  & \core_dag_ilm2reg_M7_we_DO_reg[0]/NET0131  ;
  assign n7403 = ~n7394 & ~n7395 ;
  assign n7407 = n7402 & n7403 ;
  assign n7388 = \core_c_dec_MFMreg_E_reg[5]/P0001  & \core_dag_ilm2reg_M5_we_DO_reg[0]/NET0131  ;
  assign n7389 = \core_c_dec_MFLreg_E_reg[6]/P0001  & \core_dag_ilm2reg_L6_we_DO_reg[0]/NET0131  ;
  assign n7400 = ~n7388 & ~n7389 ;
  assign n7390 = \core_c_dec_MFLreg_E_reg[7]/P0001  & \core_dag_ilm2reg_L7_we_DO_reg[0]/NET0131  ;
  assign n7391 = \core_c_dec_MFMreg_E_reg[4]/P0001  & \core_dag_ilm2reg_M4_we_DO_reg[0]/NET0131  ;
  assign n7401 = ~n7390 & ~n7391 ;
  assign n7408 = n7400 & n7401 ;
  assign n7409 = n7407 & n7408 ;
  assign n7410 = n7406 & n7409 ;
  assign n7411 = n7128 & ~n7410 ;
  assign n7439 = \core_c_dec_MFTX1_E_reg/P0001  & \sport1_txctl_TX_reg[0]/P0001  ;
  assign n7440 = \core_c_dec_MFTX0_E_reg/P0001  & \sport0_txctl_TX_reg[0]/P0001  ;
  assign n7443 = ~n7439 & ~n7440 ;
  assign n7441 = \core_c_dec_MFRX1_E_reg/P0001  & \sport1_rxctl_RX_reg[0]/P0001  ;
  assign n7442 = \core_c_dec_MFRX0_E_reg/P0001  & \sport0_rxctl_RX_reg[0]/P0001  ;
  assign n7444 = ~n7441 & ~n7442 ;
  assign n7445 = n7443 & n7444 ;
  assign n7446 = n7119 & ~n7445 ;
  assign n7595 = ~n7411 & ~n7446 ;
  assign n7596 = ~n7505 & n7595 ;
  assign n7471 = ~\core_c_psq_MSTAT_reg_DO_reg[0]/P0002  & \core_eu_em_mac_em_reg_mr2rwe_DO_reg[0]/P0001  ;
  assign n7472 = \core_c_psq_MSTAT_reg_DO_reg[0]/P0002  & \core_eu_em_mac_em_reg_mr2swe_DO_reg[0]/P0001  ;
  assign n7473 = ~n7471 & ~n7472 ;
  assign n7474 = \core_c_dec_MFMR2_E_reg/P0001  & ~n7473 ;
  assign n7463 = ~\core_c_psq_MSTAT_reg_DO_reg[0]/P0002  & \core_eu_em_mac_em_reg_mx0rwe_DO_reg[0]/P0001  ;
  assign n7464 = \core_c_psq_MSTAT_reg_DO_reg[0]/P0002  & \core_eu_em_mac_em_reg_mx0swe_DO_reg[0]/P0001  ;
  assign n7465 = ~n7463 & ~n7464 ;
  assign n7466 = \core_c_dec_MFMX0_E_reg/P0001  & ~n7465 ;
  assign n7467 = ~\core_c_psq_MSTAT_reg_DO_reg[0]/P0002  & \core_eu_em_mac_em_reg_mr0rwe_DO_reg[0]/P0001  ;
  assign n7468 = \core_c_psq_MSTAT_reg_DO_reg[0]/P0002  & \core_eu_em_mac_em_reg_mr0swe_DO_reg[0]/P0001  ;
  assign n7469 = ~n7467 & ~n7468 ;
  assign n7470 = \core_c_dec_MFMR0_E_reg/P0001  & ~n7469 ;
  assign n7477 = ~n7466 & ~n7470 ;
  assign n7478 = ~n7474 & n7477 ;
  assign n7447 = ~\core_c_psq_MSTAT_reg_DO_reg[0]/P0002  & \core_eu_em_mac_em_reg_mr1rwe_DO_reg[0]/P0001  ;
  assign n7448 = \core_c_psq_MSTAT_reg_DO_reg[0]/P0002  & \core_eu_em_mac_em_reg_mr1swe_DO_reg[0]/P0001  ;
  assign n7449 = ~n7447 & ~n7448 ;
  assign n7450 = \core_c_dec_MFMR1_E_reg/P0001  & ~n7449 ;
  assign n7451 = ~\core_c_psq_MSTAT_reg_DO_reg[0]/P0002  & \core_eu_em_mac_em_reg_my0rwe_DO_reg[0]/P0001  ;
  assign n7452 = \core_c_psq_MSTAT_reg_DO_reg[0]/P0002  & \core_eu_em_mac_em_reg_my0swe_DO_reg[0]/P0001  ;
  assign n7453 = ~n7451 & ~n7452 ;
  assign n7454 = \core_c_dec_MFMY0_E_reg/P0001  & ~n7453 ;
  assign n7475 = ~n7450 & ~n7454 ;
  assign n7455 = ~\core_c_psq_MSTAT_reg_DO_reg[0]/P0002  & \core_eu_em_mac_em_reg_mx1rwe_DO_reg[0]/P0001  ;
  assign n7456 = \core_c_psq_MSTAT_reg_DO_reg[0]/P0002  & \core_eu_em_mac_em_reg_mx1swe_DO_reg[0]/P0001  ;
  assign n7457 = ~n7455 & ~n7456 ;
  assign n7458 = \core_c_dec_MFMX1_E_reg/P0001  & ~n7457 ;
  assign n7459 = ~\core_c_psq_MSTAT_reg_DO_reg[0]/P0002  & \core_eu_em_mac_em_reg_my1rwe_DO_reg[0]/P0001  ;
  assign n7460 = \core_c_psq_MSTAT_reg_DO_reg[0]/P0002  & \core_eu_em_mac_em_reg_my1swe_DO_reg[0]/P0001  ;
  assign n7461 = ~n7459 & ~n7460 ;
  assign n7462 = \core_c_dec_MFMY1_E_reg/P0001  & ~n7461 ;
  assign n7476 = ~n7458 & ~n7462 ;
  assign n7479 = n7475 & n7476 ;
  assign n7480 = n7478 & n7479 ;
  assign n7481 = n7179 & ~n7480 ;
  assign n7363 = ~\core_c_psq_MSTAT_reg_DO_reg[0]/P0002  & \core_eu_es_sht_es_reg_SBr_reg[0]/P0001  ;
  assign n7364 = \core_c_psq_MSTAT_reg_DO_reg[0]/P0002  & \core_eu_es_sht_es_reg_SBs_reg[0]/P0001  ;
  assign n7365 = ~n7363 & ~n7364 ;
  assign n7366 = \core_c_dec_MFSB_E_reg/P0001  & ~n7365 ;
  assign n7367 = ~\core_c_psq_MSTAT_reg_DO_reg[0]/P0002  & \core_eu_es_sht_es_reg_sirwe_DO_reg[0]/P0001  ;
  assign n7368 = \core_c_psq_MSTAT_reg_DO_reg[0]/P0002  & \core_eu_es_sht_es_reg_siswe_DO_reg[0]/P0001  ;
  assign n7369 = ~n7367 & ~n7368 ;
  assign n7370 = \core_c_dec_MFSI_E_reg/P0001  & ~n7369 ;
  assign n7383 = ~n7366 & ~n7370 ;
  assign n7379 = ~\core_c_psq_MSTAT_reg_DO_reg[0]/P0002  & \core_eu_es_sht_es_reg_sr0rwe_DO_reg[0]/P0001  ;
  assign n7380 = \core_c_psq_MSTAT_reg_DO_reg[0]/P0002  & \core_eu_es_sht_es_reg_sr0swe_DO_reg[0]/P0001  ;
  assign n7381 = ~n7379 & ~n7380 ;
  assign n7382 = \core_c_dec_MFSR0_E_reg/P0001  & ~n7381 ;
  assign n7371 = ~\core_c_psq_MSTAT_reg_DO_reg[0]/P0002  & \core_eu_es_sht_es_reg_serwe_DO_reg[0]/P0001  ;
  assign n7372 = \core_c_psq_MSTAT_reg_DO_reg[0]/P0002  & \core_eu_es_sht_es_reg_seswe_DO_reg[0]/P0001  ;
  assign n7373 = ~n7371 & ~n7372 ;
  assign n7374 = \core_c_dec_MFSE_E_reg/P0001  & ~n7373 ;
  assign n7375 = ~\core_c_psq_MSTAT_reg_DO_reg[0]/P0002  & \core_eu_es_sht_es_reg_sr1rwe_DO_reg[0]/P0001  ;
  assign n7376 = \core_c_psq_MSTAT_reg_DO_reg[0]/P0002  & \core_eu_es_sht_es_reg_sr1swe_DO_reg[0]/P0001  ;
  assign n7377 = ~n7375 & ~n7376 ;
  assign n7378 = \core_c_dec_MFSR1_E_reg/P0001  & ~n7377 ;
  assign n7384 = ~n7374 & ~n7378 ;
  assign n7385 = ~n7382 & n7384 ;
  assign n7386 = n7383 & n7385 ;
  assign n7387 = n7153 & ~n7386 ;
  assign n7412 = ~\core_c_psq_MSTAT_reg_DO_reg[0]/P0002  & \core_eu_ea_alu_ea_reg_ay0rwe_DO_reg[0]/P0001  ;
  assign n7413 = \core_c_psq_MSTAT_reg_DO_reg[0]/P0002  & \core_eu_ea_alu_ea_reg_ay0swe_DO_reg[0]/P0001  ;
  assign n7414 = ~n7412 & ~n7413 ;
  assign n7415 = \core_c_dec_MFAY0_E_reg/P0001  & ~n7414 ;
  assign n7432 = \core_c_dec_MFASTAT_E_reg/P0001  & \core_eu_ec_cun_AZ_reg/P0001  ;
  assign n7433 = ~n7415 & ~n7432 ;
  assign n7416 = ~\core_c_psq_MSTAT_reg_DO_reg[0]/P0002  & \core_eu_ea_alu_ea_reg_ay1rwe_DO_reg[0]/P0001  ;
  assign n7417 = \core_c_psq_MSTAT_reg_DO_reg[0]/P0002  & \core_eu_ea_alu_ea_reg_ay1swe_DO_reg[0]/P0001  ;
  assign n7418 = ~n7416 & ~n7417 ;
  assign n7419 = \core_c_dec_MFAY1_E_reg/P0001  & ~n7418 ;
  assign n7420 = ~\core_c_psq_MSTAT_reg_DO_reg[0]/P0002  & \core_eu_ea_alu_ea_reg_arrwe_DO_reg[0]/P0001  ;
  assign n7421 = \core_c_psq_MSTAT_reg_DO_reg[0]/P0002  & \core_eu_ea_alu_ea_reg_arswe_DO_reg[0]/P0001  ;
  assign n7422 = ~n7420 & ~n7421 ;
  assign n7423 = \core_c_dec_MFAR_E_reg/P0001  & ~n7422 ;
  assign n7434 = ~n7419 & ~n7423 ;
  assign n7424 = ~\core_c_psq_MSTAT_reg_DO_reg[0]/P0002  & \core_eu_ea_alu_ea_reg_ax1rwe_DO_reg[0]/P0001  ;
  assign n7425 = \core_c_psq_MSTAT_reg_DO_reg[0]/P0002  & \core_eu_ea_alu_ea_reg_ax1swe_DO_reg[0]/P0001  ;
  assign n7426 = ~n7424 & ~n7425 ;
  assign n7427 = \core_c_dec_MFAX1_E_reg/P0001  & ~n7426 ;
  assign n7428 = ~\core_c_psq_MSTAT_reg_DO_reg[0]/P0002  & \core_eu_ea_alu_ea_reg_ax0rwe_DO_reg[0]/P0001  ;
  assign n7429 = \core_c_psq_MSTAT_reg_DO_reg[0]/P0002  & \core_eu_ea_alu_ea_reg_ax0swe_DO_reg[0]/P0001  ;
  assign n7430 = ~n7428 & ~n7429 ;
  assign n7431 = \core_c_dec_MFAX0_E_reg/P0001  & ~n7430 ;
  assign n7435 = ~n7427 & ~n7431 ;
  assign n7436 = n7434 & n7435 ;
  assign n7437 = n7433 & n7436 ;
  assign n7438 = n7093 & ~n7437 ;
  assign n7597 = ~n7387 & ~n7438 ;
  assign n7598 = ~n7481 & n7597 ;
  assign n7599 = n7596 & n7598 ;
  assign n7600 = ~n7594 & n7599 ;
  assign n7601 = ~n7574 & n7600 ;
  assign n7602 = ~n7362 & n7601 ;
  assign n7603 = ~\emc_DMDoe_reg/NET0131  & ~n7602 ;
  assign n7604 = \emc_DMDoe_reg/NET0131  & \emc_DMDreg_reg[0]/P0001  ;
  assign n7605 = n7057 & ~n7604 ;
  assign n7606 = ~n7603 & n7605 ;
  assign n7607 = ~n7361 & ~n7606 ;
  assign n7608 = n6135 & n7607 ;
  assign n7624 = n6176 & ~n7608 ;
  assign n7625 = ~n7623 & n7624 ;
  assign n7626 = ~n7343 & ~n7625 ;
  assign n7627 = n7005 & ~n7626 ;
  assign n7628 = ~n7006 & ~n7627 ;
  assign n7630 = ~\core_dag_ilm1reg_M_reg[13]/NET0131  & n6496 ;
  assign n7631 = ~n7610 & ~n7630 ;
  assign n7638 = ~n6516 & ~n6521 ;
  assign n7639 = n6427 & ~n7638 ;
  assign n7640 = ~n6427 & n7638 ;
  assign n7641 = ~n7639 & ~n7640 ;
  assign n7642 = n7631 & n7641 ;
  assign n7629 = \core_dag_ilm1reg_I_reg[10]/NET0131  & n6423 ;
  assign n7632 = ~n6419 & n6461 ;
  assign n7633 = ~n6434 & ~n6457 ;
  assign n7634 = n7632 & ~n7633 ;
  assign n7635 = ~n7632 & n7633 ;
  assign n7636 = ~n7634 & ~n7635 ;
  assign n7637 = ~n7631 & n7636 ;
  assign n7643 = ~n7629 & ~n7637 ;
  assign n7644 = ~n7642 & n7643 ;
  assign n7645 = ~n6135 & n7644 ;
  assign n7652 = \DM_rd0[10]_pad  & ~n7053 ;
  assign n7646 = \DM_rdm[10]_pad  & n7016 ;
  assign n7657 = ~n7057 & ~n7646 ;
  assign n7649 = \DM_rd6[10]_pad  & n7031 ;
  assign n7650 = \DM_rd7[10]_pad  & n7034 ;
  assign n7658 = ~n7649 & ~n7650 ;
  assign n7659 = n7657 & n7658 ;
  assign n7653 = \DM_rd5[10]_pad  & n7043 ;
  assign n7648 = \DM_rd4[10]_pad  & n7028 ;
  assign n7654 = \DM_rd2[10]_pad  & n7041 ;
  assign n7647 = \DM_rd1[10]_pad  & n7022 ;
  assign n7651 = \DM_rd3[10]_pad  & n7038 ;
  assign n7655 = ~n7647 & ~n7651 ;
  assign n7656 = ~n7654 & n7655 ;
  assign n7660 = ~n7648 & n7656 ;
  assign n7661 = ~n7653 & n7660 ;
  assign n7662 = n7659 & n7661 ;
  assign n7663 = ~n7652 & n7662 ;
  assign n7664 = \regout_STD_C_reg[10]/P0001  & n6988 ;
  assign n7692 = \bdma_BCTL_reg[10]/NET0131  & n7230 ;
  assign n7691 = \emc_WSCRreg_DO_reg[10]/NET0131  & n7251 ;
  assign n7693 = \tm_tpr_reg_DO_reg[10]/NET0131  & n7293 ;
  assign n7713 = ~n7691 & ~n7693 ;
  assign n7696 = \sport0_regs_SCTLreg_DO_reg[10]/NET0131  & n7249 ;
  assign n7697 = \tm_TCR_TMP_reg[10]/NET0131  & n7289 ;
  assign n7714 = ~n7696 & ~n7697 ;
  assign n7723 = n7713 & n7714 ;
  assign n7689 = \sport1_regs_MWORDreg_DO_reg[9]/NET0131  & n7263 ;
  assign n7690 = \sport1_txctl_Wcnt_reg[2]/NET0131  & n7689 ;
  assign n7710 = \sport0_regs_MWORDreg_DO_reg[9]/NET0131  & n7276 ;
  assign n7711 = \sport0_txctl_Wcnt_reg[2]/NET0131  & n7710 ;
  assign n7724 = ~n7690 & ~n7711 ;
  assign n7725 = n7723 & n7724 ;
  assign n7728 = ~n7692 & n7725 ;
  assign n7694 = \bdma_BEAD_reg[10]/NET0131  & n7303 ;
  assign n7698 = \bdma_BIAD_reg[10]/NET0131  & n7234 ;
  assign n7729 = ~n7694 & ~n7698 ;
  assign n7730 = n7728 & n7729 ;
  assign n7707 = \bdma_BOVL_reg[10]/NET0131  & n7534 ;
  assign n7695 = \bdma_BWCOUNT_reg[10]/NET0131  & n7287 ;
  assign n7712 = \sport0_regs_AUTOreg_DO_reg[10]/NET0131  & n7295 ;
  assign n7708 = \sport1_regs_AUTOreg_DO_reg[10]/NET0131  & n7527 ;
  assign n7709 = \idma_DCTL_reg[10]/NET0131  & n7299 ;
  assign n7719 = ~n7708 & ~n7709 ;
  assign n7720 = ~n7712 & n7719 ;
  assign n7703 = \sport0_regs_FSDIVreg_DO_reg[10]/NET0131  & n7259 ;
  assign n7704 = \memc_usysr_DO_reg[10]/NET0131  & n7301 ;
  assign n7717 = ~n7703 & ~n7704 ;
  assign n7705 = \sport1_regs_SCTLreg_DO_reg[10]/NET0131  & n7281 ;
  assign n7706 = \clkc_ckr_reg_DO_reg[10]/NET0131  & n7239 ;
  assign n7718 = ~n7705 & ~n7706 ;
  assign n7721 = n7717 & n7718 ;
  assign n7699 = \idma_DOVL_reg[10]/NET0131  & n7532 ;
  assign n7700 = \sport0_regs_SCLKDIVreg_DO_reg[10]/NET0131  & n7256 ;
  assign n7715 = ~n7699 & ~n7700 ;
  assign n7701 = \sport1_regs_SCLKDIVreg_DO_reg[10]/NET0131  & n7247 ;
  assign n7702 = \sport1_regs_FSDIVreg_DO_reg[10]/NET0131  & n7273 ;
  assign n7716 = ~n7701 & ~n7702 ;
  assign n7722 = n7715 & n7716 ;
  assign n7726 = n7721 & n7722 ;
  assign n7727 = n7720 & n7726 ;
  assign n7731 = ~n7695 & n7727 ;
  assign n7732 = ~n7707 & n7731 ;
  assign n7733 = n7730 & n7732 ;
  assign n7734 = \memc_ldSREG_E_reg/NET0131  & ~n7733 ;
  assign n7794 = \core_c_dec_MFtoppcs_Eg_reg/P0001  & ~n4276 ;
  assign n7791 = \core_c_dec_IRE_reg[14]/NET0131  & ~n7216 ;
  assign n7792 = \core_c_dec_MFCNTR_E_reg/P0001  & \core_c_psq_CNTR_reg_DO_reg[10]/NET0131  ;
  assign n7793 = \core_c_dec_MFIDR_E_reg/P0001  & \sice_idr0_reg_DO_reg[10]/P0001  ;
  assign n7795 = ~n7792 & ~n7793 ;
  assign n7796 = ~n7791 & n7795 ;
  assign n7797 = ~n7794 & n7796 ;
  assign n7798 = n7215 & ~n7797 ;
  assign n7831 = \core_c_dec_MFLreg_E_reg[5]/P0001  & \core_dag_ilm2reg_L5_we_DO_reg[10]/NET0131  ;
  assign n7832 = \core_c_dec_MFLreg_E_reg[4]/P0001  & \core_dag_ilm2reg_L4_we_DO_reg[10]/NET0131  ;
  assign n7839 = ~n7831 & ~n7832 ;
  assign n7833 = \core_c_dec_MFIreg_E_reg[7]/P0001  & \core_dag_ilm2reg_I7_we_DO_reg[10]/NET0131  ;
  assign n7834 = \core_c_dec_MFIreg_E_reg[6]/P0001  & \core_dag_ilm2reg_I6_we_DO_reg[10]/NET0131  ;
  assign n7840 = ~n7833 & ~n7834 ;
  assign n7841 = n7839 & n7840 ;
  assign n7827 = \core_c_dec_MFLreg_E_reg[6]/P0001  & \core_dag_ilm2reg_L6_we_DO_reg[10]/NET0131  ;
  assign n7828 = \core_c_dec_MFLreg_E_reg[7]/P0001  & \core_dag_ilm2reg_L7_we_DO_reg[10]/NET0131  ;
  assign n7837 = ~n7827 & ~n7828 ;
  assign n7829 = \core_c_dec_MFIreg_E_reg[5]/P0001  & \core_dag_ilm2reg_I5_we_DO_reg[10]/NET0131  ;
  assign n7830 = \core_c_dec_MFMreg_E_reg[5]/P0001  & \core_dag_ilm2reg_M5_we_DO_reg[10]/NET0131  ;
  assign n7838 = ~n7829 & ~n7830 ;
  assign n7842 = n7837 & n7838 ;
  assign n7823 = \core_c_dec_MFIreg_E_reg[4]/P0001  & \core_dag_ilm2reg_I4_we_DO_reg[10]/NET0131  ;
  assign n7824 = \core_c_dec_MFMreg_E_reg[7]/P0001  & \core_dag_ilm2reg_M7_we_DO_reg[10]/NET0131  ;
  assign n7835 = ~n7823 & ~n7824 ;
  assign n7825 = \core_c_dec_MFMreg_E_reg[6]/P0001  & \core_dag_ilm2reg_M6_we_DO_reg[10]/NET0131  ;
  assign n7826 = \core_c_dec_MFMreg_E_reg[4]/P0001  & \core_dag_ilm2reg_M4_we_DO_reg[10]/NET0131  ;
  assign n7836 = ~n7825 & ~n7826 ;
  assign n7843 = n7835 & n7836 ;
  assign n7844 = n7842 & n7843 ;
  assign n7845 = n7841 & n7844 ;
  assign n7846 = n7128 & ~n7845 ;
  assign n7673 = \core_c_dec_MFMreg_E_reg[2]/P0001  & \core_dag_ilm1reg_M2_we_DO_reg[10]/NET0131  ;
  assign n7674 = \core_c_dec_MFIreg_E_reg[0]/P0001  & \core_dag_ilm1reg_I0_we_DO_reg[10]/NET0131  ;
  assign n7681 = ~n7673 & ~n7674 ;
  assign n7675 = \core_c_dec_MFLreg_E_reg[3]/P0001  & \core_dag_ilm1reg_L3_we_DO_reg[10]/NET0131  ;
  assign n7676 = \core_c_dec_MFMreg_E_reg[1]/P0001  & \core_dag_ilm1reg_M1_we_DO_reg[10]/NET0131  ;
  assign n7682 = ~n7675 & ~n7676 ;
  assign n7683 = n7681 & n7682 ;
  assign n7669 = \core_c_dec_MFIreg_E_reg[2]/P0001  & \core_dag_ilm1reg_I2_we_DO_reg[10]/NET0131  ;
  assign n7670 = \core_c_dec_MFIreg_E_reg[3]/P0001  & \core_dag_ilm1reg_I3_we_DO_reg[10]/NET0131  ;
  assign n7679 = ~n7669 & ~n7670 ;
  assign n7671 = \core_c_dec_MFIreg_E_reg[1]/P0001  & \core_dag_ilm1reg_I1_we_DO_reg[10]/NET0131  ;
  assign n7672 = \core_c_dec_MFMreg_E_reg[3]/P0001  & \core_dag_ilm1reg_M3_we_DO_reg[10]/NET0131  ;
  assign n7680 = ~n7671 & ~n7672 ;
  assign n7684 = n7679 & n7680 ;
  assign n7665 = \core_c_dec_MFMreg_E_reg[0]/P0001  & \core_dag_ilm1reg_M0_we_DO_reg[10]/NET0131  ;
  assign n7666 = \core_c_dec_MFLreg_E_reg[0]/P0001  & \core_dag_ilm1reg_L0_we_DO_reg[10]/NET0131  ;
  assign n7677 = ~n7665 & ~n7666 ;
  assign n7667 = \core_c_dec_MFLreg_E_reg[1]/P0001  & \core_dag_ilm1reg_L1_we_DO_reg[10]/NET0131  ;
  assign n7668 = \core_c_dec_MFLreg_E_reg[2]/P0001  & \core_dag_ilm1reg_L2_we_DO_reg[10]/NET0131  ;
  assign n7678 = ~n7667 & ~n7668 ;
  assign n7685 = n7677 & n7678 ;
  assign n7686 = n7684 & n7685 ;
  assign n7687 = n7683 & n7686 ;
  assign n7688 = n7068 & ~n7687 ;
  assign n7815 = \core_c_dec_MFTX1_E_reg/P0001  & \sport1_txctl_TX_reg[10]/P0001  ;
  assign n7816 = \core_c_dec_MFRX0_E_reg/P0001  & \sport0_rxctl_RX_reg[10]/P0001  ;
  assign n7819 = ~n7815 & ~n7816 ;
  assign n7817 = \core_c_dec_MFRX1_E_reg/P0001  & \sport1_rxctl_RX_reg[10]/P0001  ;
  assign n7818 = \core_c_dec_MFTX0_E_reg/P0001  & \sport0_txctl_TX_reg[10]/P0001  ;
  assign n7820 = ~n7817 & ~n7818 ;
  assign n7821 = n7819 & n7820 ;
  assign n7822 = n7119 & ~n7821 ;
  assign n7847 = ~n7688 & ~n7822 ;
  assign n7848 = ~n7846 & n7847 ;
  assign n7807 = ~\core_c_psq_MSTAT_reg_DO_reg[0]/P0002  & \core_eu_es_sht_es_reg_sr1rwe_DO_reg[10]/P0001  ;
  assign n7808 = \core_c_psq_MSTAT_reg_DO_reg[0]/P0002  & \core_eu_es_sht_es_reg_sr1swe_DO_reg[10]/P0001  ;
  assign n7809 = ~n7807 & ~n7808 ;
  assign n7810 = \core_c_dec_MFSR1_E_reg/P0001  & ~n7809 ;
  assign n7799 = ~\core_c_psq_MSTAT_reg_DO_reg[0]/P0002  & \core_eu_es_sht_es_reg_sr0rwe_DO_reg[10]/P0001  ;
  assign n7800 = \core_c_psq_MSTAT_reg_DO_reg[0]/P0002  & \core_eu_es_sht_es_reg_sr0swe_DO_reg[10]/P0001  ;
  assign n7801 = ~n7799 & ~n7800 ;
  assign n7802 = \core_c_dec_MFSR0_E_reg/P0001  & ~n7801 ;
  assign n7803 = ~\core_c_psq_MSTAT_reg_DO_reg[0]/P0002  & \core_eu_es_sht_es_reg_sirwe_DO_reg[10]/P0001  ;
  assign n7804 = \core_c_psq_MSTAT_reg_DO_reg[0]/P0002  & \core_eu_es_sht_es_reg_siswe_DO_reg[10]/P0001  ;
  assign n7805 = ~n7803 & ~n7804 ;
  assign n7806 = \core_c_dec_MFSI_E_reg/P0001  & ~n7805 ;
  assign n7811 = ~n7802 & ~n7806 ;
  assign n7812 = ~n7810 & n7811 ;
  assign n7813 = n7174 & n7812 ;
  assign n7814 = n7153 & ~n7813 ;
  assign n7755 = ~\core_c_psq_MSTAT_reg_DO_reg[0]/P0002  & \core_eu_em_mac_em_reg_mx0rwe_DO_reg[10]/P0001  ;
  assign n7756 = \core_c_psq_MSTAT_reg_DO_reg[0]/P0002  & \core_eu_em_mac_em_reg_mx0swe_DO_reg[10]/P0001  ;
  assign n7757 = ~n7755 & ~n7756 ;
  assign n7758 = \core_c_dec_MFMX0_E_reg/P0001  & ~n7757 ;
  assign n7747 = ~\core_c_psq_MSTAT_reg_DO_reg[0]/P0002  & \core_eu_em_mac_em_reg_my1rwe_DO_reg[10]/P0001  ;
  assign n7748 = \core_c_psq_MSTAT_reg_DO_reg[0]/P0002  & \core_eu_em_mac_em_reg_my1swe_DO_reg[10]/P0001  ;
  assign n7749 = ~n7747 & ~n7748 ;
  assign n7750 = \core_c_dec_MFMY1_E_reg/P0001  & ~n7749 ;
  assign n7751 = ~\core_c_psq_MSTAT_reg_DO_reg[0]/P0002  & \core_eu_em_mac_em_reg_mr0rwe_DO_reg[10]/P0001  ;
  assign n7752 = \core_c_psq_MSTAT_reg_DO_reg[0]/P0002  & \core_eu_em_mac_em_reg_mr0swe_DO_reg[10]/P0001  ;
  assign n7753 = ~n7751 & ~n7752 ;
  assign n7754 = \core_c_dec_MFMR0_E_reg/P0001  & ~n7753 ;
  assign n7761 = ~n7750 & ~n7754 ;
  assign n7762 = ~n7758 & n7761 ;
  assign n7735 = ~\core_c_psq_MSTAT_reg_DO_reg[0]/P0002  & \core_eu_em_mac_em_reg_mr1rwe_DO_reg[10]/P0001  ;
  assign n7736 = \core_c_psq_MSTAT_reg_DO_reg[0]/P0002  & \core_eu_em_mac_em_reg_mr1swe_DO_reg[10]/P0001  ;
  assign n7737 = ~n7735 & ~n7736 ;
  assign n7738 = \core_c_dec_MFMR1_E_reg/P0001  & ~n7737 ;
  assign n7759 = ~n7207 & ~n7738 ;
  assign n7739 = ~\core_c_psq_MSTAT_reg_DO_reg[0]/P0002  & \core_eu_em_mac_em_reg_mx1rwe_DO_reg[10]/P0001  ;
  assign n7740 = \core_c_psq_MSTAT_reg_DO_reg[0]/P0002  & \core_eu_em_mac_em_reg_mx1swe_DO_reg[10]/P0001  ;
  assign n7741 = ~n7739 & ~n7740 ;
  assign n7742 = \core_c_dec_MFMX1_E_reg/P0001  & ~n7741 ;
  assign n7743 = ~\core_c_psq_MSTAT_reg_DO_reg[0]/P0002  & \core_eu_em_mac_em_reg_my0rwe_DO_reg[10]/P0001  ;
  assign n7744 = \core_c_psq_MSTAT_reg_DO_reg[0]/P0002  & \core_eu_em_mac_em_reg_my0swe_DO_reg[10]/P0001  ;
  assign n7745 = ~n7743 & ~n7744 ;
  assign n7746 = \core_c_dec_MFMY0_E_reg/P0001  & ~n7745 ;
  assign n7760 = ~n7742 & ~n7746 ;
  assign n7763 = n7759 & n7760 ;
  assign n7764 = n7762 & n7763 ;
  assign n7765 = n7179 & ~n7764 ;
  assign n7766 = ~\core_c_psq_MSTAT_reg_DO_reg[0]/P0002  & \core_eu_ea_alu_ea_reg_ax0rwe_DO_reg[10]/P0001  ;
  assign n7767 = \core_c_psq_MSTAT_reg_DO_reg[0]/P0002  & \core_eu_ea_alu_ea_reg_ax0swe_DO_reg[10]/P0001  ;
  assign n7768 = ~n7766 & ~n7767 ;
  assign n7769 = \core_c_dec_MFAX0_E_reg/P0001  & ~n7768 ;
  assign n7770 = ~\core_c_psq_MSTAT_reg_DO_reg[0]/P0002  & \core_eu_ea_alu_ea_reg_ay1rwe_DO_reg[10]/P0001  ;
  assign n7771 = \core_c_psq_MSTAT_reg_DO_reg[0]/P0002  & \core_eu_ea_alu_ea_reg_ay1swe_DO_reg[10]/P0001  ;
  assign n7772 = ~n7770 & ~n7771 ;
  assign n7773 = \core_c_dec_MFAY1_E_reg/P0001  & ~n7772 ;
  assign n7786 = ~n7769 & ~n7773 ;
  assign n7782 = ~\core_c_psq_MSTAT_reg_DO_reg[0]/P0002  & \core_eu_ea_alu_ea_reg_arrwe_DO_reg[10]/P0001  ;
  assign n7783 = \core_c_psq_MSTAT_reg_DO_reg[0]/P0002  & \core_eu_ea_alu_ea_reg_arswe_DO_reg[10]/P0001  ;
  assign n7784 = ~n7782 & ~n7783 ;
  assign n7785 = \core_c_dec_MFAR_E_reg/P0001  & ~n7784 ;
  assign n7774 = ~\core_c_psq_MSTAT_reg_DO_reg[0]/P0002  & \core_eu_ea_alu_ea_reg_ay0rwe_DO_reg[10]/P0001  ;
  assign n7775 = \core_c_psq_MSTAT_reg_DO_reg[0]/P0002  & \core_eu_ea_alu_ea_reg_ay0swe_DO_reg[10]/P0001  ;
  assign n7776 = ~n7774 & ~n7775 ;
  assign n7777 = \core_c_dec_MFAY0_E_reg/P0001  & ~n7776 ;
  assign n7778 = ~\core_c_psq_MSTAT_reg_DO_reg[0]/P0002  & \core_eu_ea_alu_ea_reg_ax1rwe_DO_reg[10]/P0001  ;
  assign n7779 = \core_c_psq_MSTAT_reg_DO_reg[0]/P0002  & \core_eu_ea_alu_ea_reg_ax1swe_DO_reg[10]/P0001  ;
  assign n7780 = ~n7778 & ~n7779 ;
  assign n7781 = \core_c_dec_MFAX1_E_reg/P0001  & ~n7780 ;
  assign n7787 = ~n7777 & ~n7781 ;
  assign n7788 = ~n7785 & n7787 ;
  assign n7789 = n7786 & n7788 ;
  assign n7790 = n7093 & ~n7789 ;
  assign n7849 = ~n7765 & ~n7790 ;
  assign n7850 = ~n7814 & n7849 ;
  assign n7851 = n7848 & n7850 ;
  assign n7852 = ~n7798 & n7851 ;
  assign n7853 = ~n7734 & n7852 ;
  assign n7854 = ~n7664 & n7853 ;
  assign n7855 = ~\emc_DMDoe_reg/NET0131  & ~n7854 ;
  assign n7856 = \emc_DMDoe_reg/NET0131  & \emc_DMDreg_reg[10]/P0001  ;
  assign n7857 = n7057 & ~n7856 ;
  assign n7858 = ~n7855 & n7857 ;
  assign n7859 = ~n7663 & ~n7858 ;
  assign n7860 = n6135 & ~n7859 ;
  assign n7861 = n6176 & ~n7860 ;
  assign n7862 = ~n7645 & n7861 ;
  assign n7863 = ~n6135 & ~n6176 ;
  assign n7870 = \DM_rd0[3]_pad  & ~n7053 ;
  assign n7864 = \DM_rdm[3]_pad  & n7016 ;
  assign n7875 = ~n7057 & ~n7864 ;
  assign n7867 = \DM_rd6[3]_pad  & n7031 ;
  assign n7868 = \DM_rd7[3]_pad  & n7034 ;
  assign n7876 = ~n7867 & ~n7868 ;
  assign n7877 = n7875 & n7876 ;
  assign n7871 = \DM_rd5[3]_pad  & n7043 ;
  assign n7866 = \DM_rd4[3]_pad  & n7028 ;
  assign n7872 = \DM_rd2[3]_pad  & n7041 ;
  assign n7865 = \DM_rd1[3]_pad  & n7022 ;
  assign n7869 = \DM_rd3[3]_pad  & n7038 ;
  assign n7873 = ~n7865 & ~n7869 ;
  assign n7874 = ~n7872 & n7873 ;
  assign n7878 = ~n7866 & n7874 ;
  assign n7879 = ~n7871 & n7878 ;
  assign n7880 = n7877 & n7879 ;
  assign n7881 = ~n7870 & n7880 ;
  assign n7882 = \regout_STD_C_reg[3]/P0001  & n6988 ;
  assign n8039 = \bdma_BIAD_reg[3]/NET0131  & n7234 ;
  assign n8030 = \emc_WSCRreg_DO_reg[3]/NET0131  & n7251 ;
  assign n8031 = \sport0_regs_SCLKDIVreg_DO_reg[3]/NET0131  & n7256 ;
  assign n8056 = ~n8030 & ~n8031 ;
  assign n8032 = \sport1_regs_MWORDreg_DO_reg[3]/NET0131  & n7263 ;
  assign n8033 = \tm_tsr_reg_DO_reg[3]/NET0131  & n7540 ;
  assign n8057 = ~n8032 & ~n8033 ;
  assign n8070 = n8056 & n8057 ;
  assign n8026 = \idma_DOVL_reg[3]/NET0131  & n7532 ;
  assign n8054 = ~n7522 & ~n8026 ;
  assign n8027 = \sport0_regs_AUTOreg_DO_reg[3]/NET0131  & n7295 ;
  assign n8028 = \tm_tpr_reg_DO_reg[3]/NET0131  & n7293 ;
  assign n8055 = ~n8027 & ~n8028 ;
  assign n8071 = n8054 & n8055 ;
  assign n8072 = n8070 & n8071 ;
  assign n8076 = ~n8039 & n8072 ;
  assign n8047 = \bdma_BEAD_reg[3]/NET0131  & n7303 ;
  assign n8048 = \bdma_BCTL_reg[3]/NET0131  & n7230 ;
  assign n8077 = ~n8047 & ~n8048 ;
  assign n8078 = n8076 & n8077 ;
  assign n8044 = \bdma_BOVL_reg[3]/NET0131  & n7534 ;
  assign n8029 = \bdma_BWCOUNT_reg[3]/NET0131  & n7287 ;
  assign n8038 = \pio_pmask_reg_DO_reg[3]/NET0131  & n7297 ;
  assign n8040 = \sport0_regs_MWORDreg_DO_reg[3]/NET0131  & n7276 ;
  assign n8060 = ~n8038 & ~n8040 ;
  assign n8041 = \sport1_regs_AUTOreg_DO_reg[3]/NET0131  & n7527 ;
  assign n8042 = \tm_TCR_TMP_reg[3]/NET0131  & n7289 ;
  assign n8061 = ~n8041 & ~n8042 ;
  assign n8068 = n8060 & n8061 ;
  assign n8034 = \sport0_regs_SCTLreg_DO_reg[3]/NET0131  & n7249 ;
  assign n8035 = \emc_WSCRext_reg_DO_reg[3]/NET0131  & n7514 ;
  assign n8058 = ~n8034 & ~n8035 ;
  assign n8036 = \sport1_regs_SCLKDIVreg_DO_reg[3]/NET0131  & n7247 ;
  assign n8037 = \sport1_regs_SCTLreg_DO_reg[3]/NET0131  & n7281 ;
  assign n8059 = ~n8036 & ~n8037 ;
  assign n8069 = n8058 & n8059 ;
  assign n8073 = n8068 & n8069 ;
  assign n8050 = \idma_DCTL_reg[3]/NET0131  & n7299 ;
  assign n8051 = \PIO_out[3]_pad  & n7291 ;
  assign n8064 = ~n8050 & ~n8051 ;
  assign n8052 = \PIO_oe[3]_pad  & n7244 ;
  assign n8053 = \sport1_regs_FSDIVreg_DO_reg[3]/NET0131  & n7273 ;
  assign n8065 = ~n8052 & ~n8053 ;
  assign n8066 = n8064 & n8065 ;
  assign n8043 = \sport0_regs_FSDIVreg_DO_reg[3]/NET0131  & n7259 ;
  assign n8045 = \clkc_ckr_reg_DO_reg[3]/NET0131  & n7239 ;
  assign n8062 = ~n8043 & ~n8045 ;
  assign n8046 = \memc_usysr_DO_reg[3]/NET0131  & n7301 ;
  assign n8049 = \pio_PINT_reg[3]/NET0131  & n7271 ;
  assign n8063 = ~n8046 & ~n8049 ;
  assign n8067 = n8062 & n8063 ;
  assign n8074 = n8066 & n8067 ;
  assign n8075 = n8073 & n8074 ;
  assign n8079 = ~n8029 & n8075 ;
  assign n8080 = ~n8044 & n8079 ;
  assign n8081 = n8078 & n8080 ;
  assign n8082 = \memc_ldSREG_E_reg/NET0131  & ~n8081 ;
  assign n8086 = \core_c_dec_MFtoppcs_Eg_reg/P0001  & ~n4328 ;
  assign n8091 = \core_c_dec_MFPMOVL_E_reg/P0001  & \core_c_psq_PMOVL_regl_DO_reg[3]/NET0131  ;
  assign n8089 = \core_c_dec_MFMSTAT_E_reg/P0001  & \core_c_psq_MSTAT_reg_DO_reg[3]/NET0131  ;
  assign n8090 = \core_c_dec_MFIDR_E_reg/P0001  & \sice_idr0_reg_DO_reg[3]/P0001  ;
  assign n8094 = ~n8089 & ~n8090 ;
  assign n8095 = ~n8091 & n8094 ;
  assign n8084 = \core_c_dec_IRE_reg[7]/NET0131  & ~n7216 ;
  assign n8083 = \core_c_dec_MFCNTR_E_reg/P0001  & \core_c_psq_CNTR_reg_DO_reg[3]/NET0131  ;
  assign n8085 = \core_c_dec_MFSSTAT_E_reg/P0001  & \core_c_psq_SSTAT_reg[3]/NET0131  ;
  assign n8092 = ~n8083 & ~n8085 ;
  assign n8087 = \core_c_dec_MFDMOVL_E_reg/P0001  & \core_c_psq_DMOVL_reg_DO_reg[3]/NET0131  ;
  assign n8088 = \core_c_dec_MFIMASK_E_reg/P0001  & \core_c_psq_IMASK_reg[3]/NET0131  ;
  assign n8093 = ~n8087 & ~n8088 ;
  assign n8096 = n8092 & n8093 ;
  assign n8097 = ~n8084 & n8096 ;
  assign n8098 = n8095 & n8097 ;
  assign n8099 = ~n8086 & n8098 ;
  assign n8100 = n7215 & ~n8099 ;
  assign n8010 = \core_c_dec_MFIreg_E_reg[4]/P0001  & \core_dag_ilm2reg_I4_we_DO_reg[3]/NET0131  ;
  assign n8011 = \core_c_dec_MFMreg_E_reg[5]/P0001  & \core_dag_ilm2reg_M5_we_DO_reg[3]/NET0131  ;
  assign n8018 = ~n8010 & ~n8011 ;
  assign n8012 = \core_c_dec_MFMreg_E_reg[6]/P0001  & \core_dag_ilm2reg_M6_we_DO_reg[3]/NET0131  ;
  assign n8013 = \core_c_dec_MFMreg_E_reg[7]/P0001  & \core_dag_ilm2reg_M7_we_DO_reg[3]/NET0131  ;
  assign n8019 = ~n8012 & ~n8013 ;
  assign n8020 = n8018 & n8019 ;
  assign n8006 = \core_c_dec_MFIreg_E_reg[5]/P0001  & \core_dag_ilm2reg_I5_we_DO_reg[3]/NET0131  ;
  assign n8007 = \core_c_dec_MFIreg_E_reg[6]/P0001  & \core_dag_ilm2reg_I6_we_DO_reg[3]/NET0131  ;
  assign n8016 = ~n8006 & ~n8007 ;
  assign n8008 = \core_c_dec_MFLreg_E_reg[7]/P0001  & \core_dag_ilm2reg_L7_we_DO_reg[3]/NET0131  ;
  assign n8009 = \core_c_dec_MFMreg_E_reg[4]/P0001  & \core_dag_ilm2reg_M4_we_DO_reg[3]/NET0131  ;
  assign n8017 = ~n8008 & ~n8009 ;
  assign n8021 = n8016 & n8017 ;
  assign n8002 = \core_c_dec_MFLreg_E_reg[6]/P0001  & \core_dag_ilm2reg_L6_we_DO_reg[3]/NET0131  ;
  assign n8003 = \core_c_dec_MFIreg_E_reg[7]/P0001  & \core_dag_ilm2reg_I7_we_DO_reg[3]/NET0131  ;
  assign n8014 = ~n8002 & ~n8003 ;
  assign n8004 = \core_c_dec_MFLreg_E_reg[4]/P0001  & \core_dag_ilm2reg_L4_we_DO_reg[3]/NET0131  ;
  assign n8005 = \core_c_dec_MFLreg_E_reg[5]/P0001  & \core_dag_ilm2reg_L5_we_DO_reg[3]/NET0131  ;
  assign n8015 = ~n8004 & ~n8005 ;
  assign n8022 = n8014 & n8015 ;
  assign n8023 = n8021 & n8022 ;
  assign n8024 = n8020 & n8023 ;
  assign n8025 = n7128 & ~n8024 ;
  assign n7926 = \core_c_dec_MFMreg_E_reg[1]/P0001  & \core_dag_ilm1reg_M1_we_DO_reg[3]/NET0131  ;
  assign n7927 = \core_c_dec_MFLreg_E_reg[2]/P0001  & \core_dag_ilm1reg_L2_we_DO_reg[3]/NET0131  ;
  assign n7934 = ~n7926 & ~n7927 ;
  assign n7928 = \core_c_dec_MFLreg_E_reg[3]/P0001  & \core_dag_ilm1reg_L3_we_DO_reg[3]/NET0131  ;
  assign n7929 = \core_c_dec_MFMreg_E_reg[0]/P0001  & \core_dag_ilm1reg_M0_we_DO_reg[3]/NET0131  ;
  assign n7935 = ~n7928 & ~n7929 ;
  assign n7936 = n7934 & n7935 ;
  assign n7922 = \core_c_dec_MFMreg_E_reg[2]/P0001  & \core_dag_ilm1reg_M2_we_DO_reg[3]/NET0131  ;
  assign n7923 = \core_c_dec_MFMreg_E_reg[3]/P0001  & \core_dag_ilm1reg_M3_we_DO_reg[3]/NET0131  ;
  assign n7932 = ~n7922 & ~n7923 ;
  assign n7924 = \core_c_dec_MFLreg_E_reg[0]/P0001  & \core_dag_ilm1reg_L0_we_DO_reg[3]/NET0131  ;
  assign n7925 = \core_c_dec_MFLreg_E_reg[1]/P0001  & \core_dag_ilm1reg_L1_we_DO_reg[3]/NET0131  ;
  assign n7933 = ~n7924 & ~n7925 ;
  assign n7937 = n7932 & n7933 ;
  assign n7918 = \core_c_dec_MFIreg_E_reg[3]/P0001  & \core_dag_ilm1reg_I3_we_DO_reg[3]/NET0131  ;
  assign n7919 = \core_c_dec_MFIreg_E_reg[0]/P0001  & \core_dag_ilm1reg_I0_we_DO_reg[3]/NET0131  ;
  assign n7930 = ~n7918 & ~n7919 ;
  assign n7920 = \core_c_dec_MFIreg_E_reg[1]/P0001  & \core_dag_ilm1reg_I1_we_DO_reg[3]/NET0131  ;
  assign n7921 = \core_c_dec_MFIreg_E_reg[2]/P0001  & \core_dag_ilm1reg_I2_we_DO_reg[3]/NET0131  ;
  assign n7931 = ~n7920 & ~n7921 ;
  assign n7938 = n7930 & n7931 ;
  assign n7939 = n7937 & n7938 ;
  assign n7940 = n7936 & n7939 ;
  assign n7941 = n7068 & ~n7940 ;
  assign n7969 = \core_c_dec_MFTX1_E_reg/P0001  & \sport1_txctl_TX_reg[3]/P0001  ;
  assign n7970 = \core_c_dec_MFTX0_E_reg/P0001  & \sport0_txctl_TX_reg[3]/P0001  ;
  assign n7973 = ~n7969 & ~n7970 ;
  assign n7971 = \core_c_dec_MFRX1_E_reg/P0001  & \sport1_rxctl_RX_reg[3]/P0001  ;
  assign n7972 = \core_c_dec_MFRX0_E_reg/P0001  & \sport0_rxctl_RX_reg[3]/P0001  ;
  assign n7974 = ~n7971 & ~n7972 ;
  assign n7975 = n7973 & n7974 ;
  assign n7976 = n7119 & ~n7975 ;
  assign n8101 = ~n7941 & ~n7976 ;
  assign n8102 = ~n8025 & n8101 ;
  assign n7977 = ~\core_c_psq_MSTAT_reg_DO_reg[0]/P0002  & \core_eu_es_sht_es_reg_sirwe_DO_reg[3]/P0001  ;
  assign n7978 = \core_c_psq_MSTAT_reg_DO_reg[0]/P0002  & \core_eu_es_sht_es_reg_siswe_DO_reg[3]/P0001  ;
  assign n7979 = ~n7977 & ~n7978 ;
  assign n7980 = \core_c_dec_MFSI_E_reg/P0001  & ~n7979 ;
  assign n7981 = ~\core_c_psq_MSTAT_reg_DO_reg[0]/P0002  & \core_eu_es_sht_es_reg_SBr_reg[3]/P0001  ;
  assign n7982 = \core_c_psq_MSTAT_reg_DO_reg[0]/P0002  & \core_eu_es_sht_es_reg_SBs_reg[3]/P0001  ;
  assign n7983 = ~n7981 & ~n7982 ;
  assign n7984 = \core_c_dec_MFSB_E_reg/P0001  & ~n7983 ;
  assign n7997 = ~n7980 & ~n7984 ;
  assign n7993 = ~\core_c_psq_MSTAT_reg_DO_reg[0]/P0002  & \core_eu_es_sht_es_reg_serwe_DO_reg[3]/P0001  ;
  assign n7994 = \core_c_psq_MSTAT_reg_DO_reg[0]/P0002  & \core_eu_es_sht_es_reg_seswe_DO_reg[3]/P0001  ;
  assign n7995 = ~n7993 & ~n7994 ;
  assign n7996 = \core_c_dec_MFSE_E_reg/P0001  & ~n7995 ;
  assign n7985 = ~\core_c_psq_MSTAT_reg_DO_reg[0]/P0002  & \core_eu_es_sht_es_reg_sr0rwe_DO_reg[3]/P0001  ;
  assign n7986 = \core_c_psq_MSTAT_reg_DO_reg[0]/P0002  & \core_eu_es_sht_es_reg_sr0swe_DO_reg[3]/P0001  ;
  assign n7987 = ~n7985 & ~n7986 ;
  assign n7988 = \core_c_dec_MFSR0_E_reg/P0001  & ~n7987 ;
  assign n7989 = ~\core_c_psq_MSTAT_reg_DO_reg[0]/P0002  & \core_eu_es_sht_es_reg_sr1rwe_DO_reg[3]/P0001  ;
  assign n7990 = \core_c_psq_MSTAT_reg_DO_reg[0]/P0002  & \core_eu_es_sht_es_reg_sr1swe_DO_reg[3]/P0001  ;
  assign n7991 = ~n7989 & ~n7990 ;
  assign n7992 = \core_c_dec_MFSR1_E_reg/P0001  & ~n7991 ;
  assign n7998 = ~n7988 & ~n7992 ;
  assign n7999 = ~n7996 & n7998 ;
  assign n8000 = n7997 & n7999 ;
  assign n8001 = n7153 & ~n8000 ;
  assign n7907 = ~\core_c_psq_MSTAT_reg_DO_reg[0]/P0002  & \core_eu_em_mac_em_reg_mr0rwe_DO_reg[3]/P0001  ;
  assign n7908 = \core_c_psq_MSTAT_reg_DO_reg[0]/P0002  & \core_eu_em_mac_em_reg_mr0swe_DO_reg[3]/P0001  ;
  assign n7909 = ~n7907 & ~n7908 ;
  assign n7910 = \core_c_dec_MFMR0_E_reg/P0001  & ~n7909 ;
  assign n7899 = ~\core_c_psq_MSTAT_reg_DO_reg[0]/P0002  & \core_eu_em_mac_em_reg_mx1rwe_DO_reg[3]/P0001  ;
  assign n7900 = \core_c_psq_MSTAT_reg_DO_reg[0]/P0002  & \core_eu_em_mac_em_reg_mx1swe_DO_reg[3]/P0001  ;
  assign n7901 = ~n7899 & ~n7900 ;
  assign n7902 = \core_c_dec_MFMX1_E_reg/P0001  & ~n7901 ;
  assign n7903 = ~\core_c_psq_MSTAT_reg_DO_reg[0]/P0002  & \core_eu_em_mac_em_reg_mr2rwe_DO_reg[3]/P0001  ;
  assign n7904 = \core_c_psq_MSTAT_reg_DO_reg[0]/P0002  & \core_eu_em_mac_em_reg_mr2swe_DO_reg[3]/P0001  ;
  assign n7905 = ~n7903 & ~n7904 ;
  assign n7906 = \core_c_dec_MFMR2_E_reg/P0001  & ~n7905 ;
  assign n7913 = ~n7902 & ~n7906 ;
  assign n7914 = ~n7910 & n7913 ;
  assign n7883 = ~\core_c_psq_MSTAT_reg_DO_reg[0]/P0002  & \core_eu_em_mac_em_reg_mr1rwe_DO_reg[3]/P0001  ;
  assign n7884 = \core_c_psq_MSTAT_reg_DO_reg[0]/P0002  & \core_eu_em_mac_em_reg_mr1swe_DO_reg[3]/P0001  ;
  assign n7885 = ~n7883 & ~n7884 ;
  assign n7886 = \core_c_dec_MFMR1_E_reg/P0001  & ~n7885 ;
  assign n7887 = ~\core_c_psq_MSTAT_reg_DO_reg[0]/P0002  & \core_eu_em_mac_em_reg_mx0rwe_DO_reg[3]/P0001  ;
  assign n7888 = \core_c_psq_MSTAT_reg_DO_reg[0]/P0002  & \core_eu_em_mac_em_reg_mx0swe_DO_reg[3]/P0001  ;
  assign n7889 = ~n7887 & ~n7888 ;
  assign n7890 = \core_c_dec_MFMX0_E_reg/P0001  & ~n7889 ;
  assign n7911 = ~n7886 & ~n7890 ;
  assign n7891 = ~\core_c_psq_MSTAT_reg_DO_reg[0]/P0002  & \core_eu_em_mac_em_reg_my1rwe_DO_reg[3]/P0001  ;
  assign n7892 = \core_c_psq_MSTAT_reg_DO_reg[0]/P0002  & \core_eu_em_mac_em_reg_my1swe_DO_reg[3]/P0001  ;
  assign n7893 = ~n7891 & ~n7892 ;
  assign n7894 = \core_c_dec_MFMY1_E_reg/P0001  & ~n7893 ;
  assign n7895 = ~\core_c_psq_MSTAT_reg_DO_reg[0]/P0002  & \core_eu_em_mac_em_reg_my0rwe_DO_reg[3]/P0001  ;
  assign n7896 = \core_c_psq_MSTAT_reg_DO_reg[0]/P0002  & \core_eu_em_mac_em_reg_my0swe_DO_reg[3]/P0001  ;
  assign n7897 = ~n7895 & ~n7896 ;
  assign n7898 = \core_c_dec_MFMY0_E_reg/P0001  & ~n7897 ;
  assign n7912 = ~n7894 & ~n7898 ;
  assign n7915 = n7911 & n7912 ;
  assign n7916 = n7914 & n7915 ;
  assign n7917 = n7179 & ~n7916 ;
  assign n7942 = ~\core_c_psq_MSTAT_reg_DO_reg[0]/P0002  & \core_eu_ea_alu_ea_reg_ay0rwe_DO_reg[3]/P0001  ;
  assign n7943 = \core_c_psq_MSTAT_reg_DO_reg[0]/P0002  & \core_eu_ea_alu_ea_reg_ay0swe_DO_reg[3]/P0001  ;
  assign n7944 = ~n7942 & ~n7943 ;
  assign n7945 = \core_c_dec_MFAY0_E_reg/P0001  & ~n7944 ;
  assign n7962 = \core_c_dec_MFASTAT_E_reg/P0001  & \core_eu_ec_cun_AC_reg/P0001  ;
  assign n7963 = ~n7945 & ~n7962 ;
  assign n7946 = ~\core_c_psq_MSTAT_reg_DO_reg[0]/P0002  & \core_eu_ea_alu_ea_reg_ay1rwe_DO_reg[3]/P0001  ;
  assign n7947 = \core_c_psq_MSTAT_reg_DO_reg[0]/P0002  & \core_eu_ea_alu_ea_reg_ay1swe_DO_reg[3]/P0001  ;
  assign n7948 = ~n7946 & ~n7947 ;
  assign n7949 = \core_c_dec_MFAY1_E_reg/P0001  & ~n7948 ;
  assign n7950 = ~\core_c_psq_MSTAT_reg_DO_reg[0]/P0002  & \core_eu_ea_alu_ea_reg_arrwe_DO_reg[3]/P0001  ;
  assign n7951 = \core_c_psq_MSTAT_reg_DO_reg[0]/P0002  & \core_eu_ea_alu_ea_reg_arswe_DO_reg[3]/P0001  ;
  assign n7952 = ~n7950 & ~n7951 ;
  assign n7953 = \core_c_dec_MFAR_E_reg/P0001  & ~n7952 ;
  assign n7964 = ~n7949 & ~n7953 ;
  assign n7954 = ~\core_c_psq_MSTAT_reg_DO_reg[0]/P0002  & \core_eu_ea_alu_ea_reg_ax1rwe_DO_reg[3]/P0001  ;
  assign n7955 = \core_c_psq_MSTAT_reg_DO_reg[0]/P0002  & \core_eu_ea_alu_ea_reg_ax1swe_DO_reg[3]/P0001  ;
  assign n7956 = ~n7954 & ~n7955 ;
  assign n7957 = \core_c_dec_MFAX1_E_reg/P0001  & ~n7956 ;
  assign n7958 = ~\core_c_psq_MSTAT_reg_DO_reg[0]/P0002  & \core_eu_ea_alu_ea_reg_ax0rwe_DO_reg[3]/P0001  ;
  assign n7959 = \core_c_psq_MSTAT_reg_DO_reg[0]/P0002  & \core_eu_ea_alu_ea_reg_ax0swe_DO_reg[3]/P0001  ;
  assign n7960 = ~n7958 & ~n7959 ;
  assign n7961 = \core_c_dec_MFAX0_E_reg/P0001  & ~n7960 ;
  assign n7965 = ~n7957 & ~n7961 ;
  assign n7966 = n7964 & n7965 ;
  assign n7967 = n7963 & n7966 ;
  assign n7968 = n7093 & ~n7967 ;
  assign n8103 = ~n7917 & ~n7968 ;
  assign n8104 = ~n8001 & n8103 ;
  assign n8105 = n8102 & n8104 ;
  assign n8106 = ~n8100 & n8105 ;
  assign n8107 = ~n8082 & n8106 ;
  assign n8108 = ~n7882 & n8107 ;
  assign n8109 = ~\emc_DMDoe_reg/NET0131  & ~n8108 ;
  assign n8110 = \emc_DMDoe_reg/NET0131  & \emc_DMDreg_reg[3]/P0001  ;
  assign n8111 = n7057 & ~n8110 ;
  assign n8112 = ~n8109 & n8111 ;
  assign n8113 = ~n7881 & ~n8112 ;
  assign n8114 = n7863 & n8113 ;
  assign n8115 = \core_dag_ilm2reg_I7_we_DO_reg[10]/NET0131  & n6972 ;
  assign n8116 = \core_dag_ilm2reg_I4_we_DO_reg[10]/NET0131  & n6976 ;
  assign n8119 = ~n8115 & ~n8116 ;
  assign n8117 = \core_dag_ilm2reg_I6_we_DO_reg[10]/NET0131  & n6974 ;
  assign n8118 = \core_dag_ilm2reg_I5_we_DO_reg[10]/NET0131  & n6970 ;
  assign n8120 = ~n8117 & ~n8118 ;
  assign n8121 = n8119 & n8120 ;
  assign n8122 = n4055 & ~n8121 ;
  assign n8123 = \core_dag_ilm2reg_I4_we_DO_reg[10]/NET0131  & n6958 ;
  assign n8124 = \core_dag_ilm2reg_I7_we_DO_reg[10]/NET0131  & n6960 ;
  assign n8127 = ~n8123 & ~n8124 ;
  assign n8125 = \core_dag_ilm2reg_I6_we_DO_reg[10]/NET0131  & n6962 ;
  assign n8126 = \core_dag_ilm2reg_I5_we_DO_reg[10]/NET0131  & n6964 ;
  assign n8128 = ~n8125 & ~n8126 ;
  assign n8129 = n8127 & n8128 ;
  assign n8130 = ~n8122 & n8129 ;
  assign n8131 = n6058 & n6060 ;
  assign n8132 = \core_dag_ilm1reg_I0_we_DO_reg[10]/NET0131  & n8131 ;
  assign n8139 = ~n4055 & ~n8132 ;
  assign n8137 = \core_dag_ilm1reg_I3_we_DO_reg[10]/NET0131  & n6075 ;
  assign n8138 = n6077 & n8137 ;
  assign n8133 = \core_dag_ilm1reg_I2_we_DO_reg[10]/NET0131  & n6084 ;
  assign n8134 = n6085 & n8133 ;
  assign n8135 = \core_dag_ilm1reg_I1_we_DO_reg[10]/NET0131  & n6067 ;
  assign n8136 = n6068 & n8135 ;
  assign n8140 = ~n8134 & ~n8136 ;
  assign n8141 = ~n8138 & n8140 ;
  assign n8142 = n8139 & n8141 ;
  assign n8143 = n6097 & n8137 ;
  assign n8144 = n6095 & n8133 ;
  assign n8147 = ~n8143 & ~n8144 ;
  assign n8145 = n6091 & n8135 ;
  assign n8146 = \core_dag_ilm1reg_I0_we_DO_reg[10]/NET0131  & n6148 ;
  assign n8148 = ~n8145 & ~n8146 ;
  assign n8149 = n8147 & n8148 ;
  assign n8150 = n4055 & n8149 ;
  assign n8151 = ~n8142 & ~n8150 ;
  assign n8152 = n8130 & ~n8151 ;
  assign n8153 = n6135 & ~n6176 ;
  assign n8154 = ~n8152 & n8153 ;
  assign n8155 = ~n8114 & ~n8154 ;
  assign n8156 = ~n7862 & n8155 ;
  assign n8157 = n7005 & ~n8156 ;
  assign n8218 = ~n6326 & ~n6327 ;
  assign n8219 = ~n6370 & n8218 ;
  assign n8220 = n6370 & ~n8218 ;
  assign n8221 = ~n8219 & ~n8220 ;
  assign n8222 = ~n7631 & n8221 ;
  assign n8213 = \core_dag_ilm1reg_I_reg[3]/NET0131  & ~n6295 ;
  assign n8214 = ~n6310 & ~n6503 ;
  assign n8215 = n6310 & n6503 ;
  assign n8216 = ~n8214 & ~n8215 ;
  assign n8217 = n7631 & n8216 ;
  assign n8223 = ~n8213 & ~n8217 ;
  assign n8224 = ~n8222 & n8223 ;
  assign n8225 = n6176 & ~n8224 ;
  assign n8196 = \core_dag_ilm2reg_I_reg[10]/NET0131  & ~n6620 ;
  assign n8197 = ~\core_dag_ilm2reg_M_reg[13]/NET0131  & ~n6905 ;
  assign n8198 = ~n6714 & ~n8197 ;
  assign n8199 = ~n6699 & ~n6706 ;
  assign n8200 = ~n6850 & ~n8199 ;
  assign n8201 = n6850 & n8199 ;
  assign n8202 = ~n8200 & ~n8201 ;
  assign n8203 = ~n8198 & n8202 ;
  assign n8204 = ~n6847 & n6875 ;
  assign n8205 = ~n6857 & ~n6870 ;
  assign n8206 = ~n8204 & ~n8205 ;
  assign n8207 = n8204 & n8205 ;
  assign n8208 = ~n8206 & ~n8207 ;
  assign n8209 = n8198 & n8208 ;
  assign n8210 = ~n8203 & ~n8209 ;
  assign n8211 = ~n8196 & ~n8210 ;
  assign n8212 = ~n6176 & ~n8211 ;
  assign n8226 = n6135 & ~n8212 ;
  assign n8227 = ~n8225 & n8226 ;
  assign n8163 = ~n6111 & n8151 ;
  assign n8161 = ~n6121 & ~n8130 ;
  assign n8162 = \core_c_dec_IR_reg[14]/NET0131  & n6956 ;
  assign n8164 = ~n8161 & ~n8162 ;
  assign n8165 = ~n8163 & n8164 ;
  assign n8166 = n5949 & ~n8165 ;
  assign n8167 = \core_dag_ilm1reg_DMA_pi_DO_reg[10]/NET0131  & ~n6934 ;
  assign n8159 = \idma_DCTL_reg[10]/NET0131  & n6926 ;
  assign n8160 = \core_dag_ilm1reg_STAC_pi_DO_reg[10]/NET0131  & n6988 ;
  assign n8168 = ~n8159 & ~n8160 ;
  assign n8169 = n6924 & n8168 ;
  assign n8170 = ~n8167 & n8169 ;
  assign n8171 = ~n8166 & n8170 ;
  assign n8158 = ~\bdma_BIAD_reg[10]/NET0131  & ~n6924 ;
  assign n8172 = ~n6176 & ~n8158 ;
  assign n8173 = ~n8171 & n8172 ;
  assign n8174 = \core_dag_ilm1reg_I0_we_DO_reg[3]/NET0131  & n8131 ;
  assign n8179 = ~n4055 & ~n8174 ;
  assign n8177 = \core_dag_ilm1reg_I2_we_DO_reg[3]/NET0131  & n6084 ;
  assign n8178 = n6085 & n8177 ;
  assign n8175 = \core_dag_ilm1reg_I3_we_DO_reg[3]/NET0131  & n6140 ;
  assign n8176 = \core_dag_ilm1reg_I1_we_DO_reg[3]/NET0131  & n6142 ;
  assign n8180 = ~n8175 & ~n8176 ;
  assign n8181 = ~n8178 & n8180 ;
  assign n8182 = n8179 & n8181 ;
  assign n8183 = \core_dag_ilm1reg_I2_we_DO_reg[3]/NET0131  & n6152 ;
  assign n8184 = \core_dag_ilm1reg_I3_we_DO_reg[3]/NET0131  & n6150 ;
  assign n8188 = ~n8183 & ~n8184 ;
  assign n8185 = \core_dag_ilm1reg_I1_we_DO_reg[3]/NET0131  & n6154 ;
  assign n8186 = \core_dag_ilm1reg_I0_we_DO_reg[3]/NET0131  & n6058 ;
  assign n8187 = n6093 & n8186 ;
  assign n8189 = ~n8185 & ~n8187 ;
  assign n8190 = n8188 & n8189 ;
  assign n8191 = n4055 & n8190 ;
  assign n8192 = ~n8182 & ~n8191 ;
  assign n8193 = n6176 & n8192 ;
  assign n8194 = ~n6135 & ~n8193 ;
  assign n8195 = ~n8173 & n8194 ;
  assign n8228 = ~n7005 & ~n8195 ;
  assign n8229 = ~n8227 & n8228 ;
  assign n8230 = ~n8157 & ~n8229 ;
  assign n8239 = ~n6425 & ~n7638 ;
  assign n8240 = ~n6426 & ~n8239 ;
  assign n8241 = n6446 & ~n8240 ;
  assign n8242 = ~n6446 & n8240 ;
  assign n8243 = ~n8241 & ~n8242 ;
  assign n8244 = n7631 & n8243 ;
  assign n8231 = \core_dag_ilm1reg_I_reg[11]/NET0131  & ~n6442 ;
  assign n8232 = ~n6453 & ~n6456 ;
  assign n8233 = ~n6457 & n7632 ;
  assign n8234 = ~n6434 & ~n8233 ;
  assign n8235 = ~n8232 & ~n8234 ;
  assign n8236 = n8232 & n8234 ;
  assign n8237 = ~n8235 & ~n8236 ;
  assign n8238 = ~n7631 & n8237 ;
  assign n8245 = ~n8231 & ~n8238 ;
  assign n8246 = ~n8244 & n8245 ;
  assign n8247 = ~n6135 & n8246 ;
  assign n8254 = \DM_rd0[11]_pad  & ~n7053 ;
  assign n8248 = \DM_rdm[11]_pad  & n7016 ;
  assign n8259 = ~n7057 & ~n8248 ;
  assign n8251 = \DM_rd6[11]_pad  & n7031 ;
  assign n8252 = \DM_rd7[11]_pad  & n7034 ;
  assign n8260 = ~n8251 & ~n8252 ;
  assign n8261 = n8259 & n8260 ;
  assign n8255 = \DM_rd5[11]_pad  & n7043 ;
  assign n8250 = \DM_rd4[11]_pad  & n7028 ;
  assign n8256 = \DM_rd2[11]_pad  & n7041 ;
  assign n8249 = \DM_rd1[11]_pad  & n7022 ;
  assign n8253 = \DM_rd3[11]_pad  & n7038 ;
  assign n8257 = ~n8249 & ~n8253 ;
  assign n8258 = ~n8256 & n8257 ;
  assign n8262 = ~n8250 & n8258 ;
  assign n8263 = ~n8255 & n8262 ;
  assign n8264 = n8261 & n8263 ;
  assign n8265 = ~n8254 & n8264 ;
  assign n8266 = \regout_STD_C_reg[11]/P0001  & n6988 ;
  assign n8293 = \bdma_BCTL_reg[11]/NET0131  & n7230 ;
  assign n8291 = \tm_tpr_reg_DO_reg[11]/NET0131  & n7293 ;
  assign n8313 = ~n7522 & ~n8291 ;
  assign n8292 = \sport1_regs_SCLKDIVreg_DO_reg[11]/NET0131  & n7247 ;
  assign n8294 = \idma_DCTL_reg[11]/NET0131  & n7299 ;
  assign n8314 = ~n8292 & ~n8294 ;
  assign n8324 = n8313 & n8314 ;
  assign n8308 = \sport1_txctl_Wcnt_reg[3]/NET0131  & n7689 ;
  assign n8309 = \sport0_txctl_Wcnt_reg[3]/NET0131  & n7710 ;
  assign n8325 = ~n8308 & ~n8309 ;
  assign n8326 = n8324 & n8325 ;
  assign n8329 = ~n8293 & n8326 ;
  assign n8295 = \bdma_BIAD_reg[11]/NET0131  & n7234 ;
  assign n8298 = \bdma_BEAD_reg[11]/NET0131  & n7303 ;
  assign n8330 = ~n8295 & ~n8298 ;
  assign n8331 = n8329 & n8330 ;
  assign n8307 = \bdma_BWCOUNT_reg[11]/NET0131  & n7287 ;
  assign n8296 = \bdma_BOVL_reg[11]/NET0131  & n7534 ;
  assign n8306 = \sport1_regs_AUTOreg_DO_reg[11]/NET0131  & n7527 ;
  assign n8310 = \memc_usysr_DO_reg[11]/NET0131  & n7301 ;
  assign n8319 = ~n8306 & ~n8310 ;
  assign n8311 = \clkc_ckr_reg_DO_reg[11]/NET0131  & n7239 ;
  assign n8312 = \sport0_regs_SCLKDIVreg_DO_reg[11]/NET0131  & n7256 ;
  assign n8320 = ~n8311 & ~n8312 ;
  assign n8321 = n8319 & n8320 ;
  assign n8302 = \sport0_regs_AUTOreg_DO_reg[11]/NET0131  & n7295 ;
  assign n8303 = \emc_WSCRreg_DO_reg[11]/NET0131  & n7251 ;
  assign n8317 = ~n8302 & ~n8303 ;
  assign n8304 = \sport1_regs_FSDIVreg_DO_reg[11]/NET0131  & n7273 ;
  assign n8305 = \sport1_regs_SCTLreg_DO_reg[11]/NET0131  & n7281 ;
  assign n8318 = ~n8304 & ~n8305 ;
  assign n8322 = n8317 & n8318 ;
  assign n8297 = \idma_DOVL_reg[11]/NET0131  & n7532 ;
  assign n8299 = \sport0_regs_FSDIVreg_DO_reg[11]/NET0131  & n7259 ;
  assign n8315 = ~n8297 & ~n8299 ;
  assign n8300 = \sport0_regs_SCTLreg_DO_reg[11]/NET0131  & n7249 ;
  assign n8301 = \tm_TCR_TMP_reg[11]/NET0131  & n7289 ;
  assign n8316 = ~n8300 & ~n8301 ;
  assign n8323 = n8315 & n8316 ;
  assign n8327 = n8322 & n8323 ;
  assign n8328 = n8321 & n8327 ;
  assign n8332 = ~n8296 & n8328 ;
  assign n8333 = ~n8307 & n8332 ;
  assign n8334 = n8331 & n8333 ;
  assign n8335 = \memc_ldSREG_E_reg/NET0131  & ~n8334 ;
  assign n8395 = \core_c_dec_MFtoppcs_Eg_reg/P0001  & ~n4622 ;
  assign n8392 = \core_c_dec_IRE_reg[15]/NET0131  & ~n7216 ;
  assign n8393 = \core_c_dec_MFCNTR_E_reg/P0001  & \core_c_psq_CNTR_reg_DO_reg[11]/NET0131  ;
  assign n8394 = \core_c_dec_MFIDR_E_reg/P0001  & \sice_idr0_reg_DO_reg[11]/P0001  ;
  assign n8396 = ~n8393 & ~n8394 ;
  assign n8397 = ~n8392 & n8396 ;
  assign n8398 = ~n8395 & n8397 ;
  assign n8399 = n7215 & ~n8398 ;
  assign n8432 = \core_c_dec_MFMreg_E_reg[0]/P0001  & \core_dag_ilm1reg_M0_we_DO_reg[11]/NET0131  ;
  assign n8433 = \core_c_dec_MFLreg_E_reg[3]/P0001  & \core_dag_ilm1reg_L3_we_DO_reg[11]/NET0131  ;
  assign n8440 = ~n8432 & ~n8433 ;
  assign n8434 = \core_c_dec_MFLreg_E_reg[2]/P0001  & \core_dag_ilm1reg_L2_we_DO_reg[11]/NET0131  ;
  assign n8435 = \core_c_dec_MFMreg_E_reg[3]/P0001  & \core_dag_ilm1reg_M3_we_DO_reg[11]/NET0131  ;
  assign n8441 = ~n8434 & ~n8435 ;
  assign n8442 = n8440 & n8441 ;
  assign n8428 = \core_c_dec_MFIreg_E_reg[3]/P0001  & \core_dag_ilm1reg_I3_we_DO_reg[11]/NET0131  ;
  assign n8429 = \core_c_dec_MFLreg_E_reg[0]/P0001  & \core_dag_ilm1reg_L0_we_DO_reg[11]/NET0131  ;
  assign n8438 = ~n8428 & ~n8429 ;
  assign n8430 = \core_c_dec_MFMreg_E_reg[2]/P0001  & \core_dag_ilm1reg_M2_we_DO_reg[11]/NET0131  ;
  assign n8431 = \core_c_dec_MFIreg_E_reg[0]/P0001  & \core_dag_ilm1reg_I0_we_DO_reg[11]/NET0131  ;
  assign n8439 = ~n8430 & ~n8431 ;
  assign n8443 = n8438 & n8439 ;
  assign n8424 = \core_c_dec_MFMreg_E_reg[1]/P0001  & \core_dag_ilm1reg_M1_we_DO_reg[11]/NET0131  ;
  assign n8425 = \core_c_dec_MFIreg_E_reg[2]/P0001  & \core_dag_ilm1reg_I2_we_DO_reg[11]/NET0131  ;
  assign n8436 = ~n8424 & ~n8425 ;
  assign n8426 = \core_c_dec_MFIreg_E_reg[1]/P0001  & \core_dag_ilm1reg_I1_we_DO_reg[11]/NET0131  ;
  assign n8427 = \core_c_dec_MFLreg_E_reg[1]/P0001  & \core_dag_ilm1reg_L1_we_DO_reg[11]/NET0131  ;
  assign n8437 = ~n8426 & ~n8427 ;
  assign n8444 = n8436 & n8437 ;
  assign n8445 = n8443 & n8444 ;
  assign n8446 = n8442 & n8445 ;
  assign n8447 = n7068 & ~n8446 ;
  assign n8275 = \core_c_dec_MFLreg_E_reg[7]/P0001  & \core_dag_ilm2reg_L7_we_DO_reg[11]/NET0131  ;
  assign n8276 = \core_c_dec_MFIreg_E_reg[7]/P0001  & \core_dag_ilm2reg_I7_we_DO_reg[11]/NET0131  ;
  assign n8283 = ~n8275 & ~n8276 ;
  assign n8277 = \core_c_dec_MFMreg_E_reg[6]/P0001  & \core_dag_ilm2reg_M6_we_DO_reg[11]/NET0131  ;
  assign n8278 = \core_c_dec_MFLreg_E_reg[6]/P0001  & \core_dag_ilm2reg_L6_we_DO_reg[11]/NET0131  ;
  assign n8284 = ~n8277 & ~n8278 ;
  assign n8285 = n8283 & n8284 ;
  assign n8271 = \core_c_dec_MFLreg_E_reg[5]/P0001  & \core_dag_ilm2reg_L5_we_DO_reg[11]/NET0131  ;
  assign n8272 = \core_c_dec_MFIreg_E_reg[4]/P0001  & \core_dag_ilm2reg_I4_we_DO_reg[11]/NET0131  ;
  assign n8281 = ~n8271 & ~n8272 ;
  assign n8273 = \core_c_dec_MFLreg_E_reg[4]/P0001  & \core_dag_ilm2reg_L4_we_DO_reg[11]/NET0131  ;
  assign n8274 = \core_c_dec_MFMreg_E_reg[4]/P0001  & \core_dag_ilm2reg_M4_we_DO_reg[11]/NET0131  ;
  assign n8282 = ~n8273 & ~n8274 ;
  assign n8286 = n8281 & n8282 ;
  assign n8267 = \core_c_dec_MFMreg_E_reg[7]/P0001  & \core_dag_ilm2reg_M7_we_DO_reg[11]/NET0131  ;
  assign n8268 = \core_c_dec_MFIreg_E_reg[5]/P0001  & \core_dag_ilm2reg_I5_we_DO_reg[11]/NET0131  ;
  assign n8279 = ~n8267 & ~n8268 ;
  assign n8269 = \core_c_dec_MFIreg_E_reg[6]/P0001  & \core_dag_ilm2reg_I6_we_DO_reg[11]/NET0131  ;
  assign n8270 = \core_c_dec_MFMreg_E_reg[5]/P0001  & \core_dag_ilm2reg_M5_we_DO_reg[11]/NET0131  ;
  assign n8280 = ~n8269 & ~n8270 ;
  assign n8287 = n8279 & n8280 ;
  assign n8288 = n8286 & n8287 ;
  assign n8289 = n8285 & n8288 ;
  assign n8290 = n7128 & ~n8289 ;
  assign n8416 = \core_c_dec_MFTX1_E_reg/P0001  & \sport1_txctl_TX_reg[11]/P0001  ;
  assign n8417 = \core_c_dec_MFTX0_E_reg/P0001  & \sport0_txctl_TX_reg[11]/P0001  ;
  assign n8420 = ~n8416 & ~n8417 ;
  assign n8418 = \core_c_dec_MFRX1_E_reg/P0001  & \sport1_rxctl_RX_reg[11]/P0001  ;
  assign n8419 = \core_c_dec_MFRX0_E_reg/P0001  & \sport0_rxctl_RX_reg[11]/P0001  ;
  assign n8421 = ~n8418 & ~n8419 ;
  assign n8422 = n8420 & n8421 ;
  assign n8423 = n7119 & ~n8422 ;
  assign n8448 = ~n8290 & ~n8423 ;
  assign n8449 = ~n8447 & n8448 ;
  assign n8408 = ~\core_c_psq_MSTAT_reg_DO_reg[0]/P0002  & \core_eu_es_sht_es_reg_sr1rwe_DO_reg[11]/P0001  ;
  assign n8409 = \core_c_psq_MSTAT_reg_DO_reg[0]/P0002  & \core_eu_es_sht_es_reg_sr1swe_DO_reg[11]/P0001  ;
  assign n8410 = ~n8408 & ~n8409 ;
  assign n8411 = \core_c_dec_MFSR1_E_reg/P0001  & ~n8410 ;
  assign n8400 = ~\core_c_psq_MSTAT_reg_DO_reg[0]/P0002  & \core_eu_es_sht_es_reg_sr0rwe_DO_reg[11]/P0001  ;
  assign n8401 = \core_c_psq_MSTAT_reg_DO_reg[0]/P0002  & \core_eu_es_sht_es_reg_sr0swe_DO_reg[11]/P0001  ;
  assign n8402 = ~n8400 & ~n8401 ;
  assign n8403 = \core_c_dec_MFSR0_E_reg/P0001  & ~n8402 ;
  assign n8404 = ~\core_c_psq_MSTAT_reg_DO_reg[0]/P0002  & \core_eu_es_sht_es_reg_sirwe_DO_reg[11]/P0001  ;
  assign n8405 = \core_c_psq_MSTAT_reg_DO_reg[0]/P0002  & \core_eu_es_sht_es_reg_siswe_DO_reg[11]/P0001  ;
  assign n8406 = ~n8404 & ~n8405 ;
  assign n8407 = \core_c_dec_MFSI_E_reg/P0001  & ~n8406 ;
  assign n8412 = ~n8403 & ~n8407 ;
  assign n8413 = ~n8411 & n8412 ;
  assign n8414 = n7174 & n8413 ;
  assign n8415 = n7153 & ~n8414 ;
  assign n8356 = ~\core_c_psq_MSTAT_reg_DO_reg[0]/P0002  & \core_eu_em_mac_em_reg_mr1rwe_DO_reg[11]/P0001  ;
  assign n8357 = \core_c_psq_MSTAT_reg_DO_reg[0]/P0002  & \core_eu_em_mac_em_reg_mr1swe_DO_reg[11]/P0001  ;
  assign n8358 = ~n8356 & ~n8357 ;
  assign n8359 = \core_c_dec_MFMR1_E_reg/P0001  & ~n8358 ;
  assign n8348 = ~\core_c_psq_MSTAT_reg_DO_reg[0]/P0002  & \core_eu_em_mac_em_reg_mx1rwe_DO_reg[11]/P0001  ;
  assign n8349 = \core_c_psq_MSTAT_reg_DO_reg[0]/P0002  & \core_eu_em_mac_em_reg_mx1swe_DO_reg[11]/P0001  ;
  assign n8350 = ~n8348 & ~n8349 ;
  assign n8351 = \core_c_dec_MFMX1_E_reg/P0001  & ~n8350 ;
  assign n8352 = ~\core_c_psq_MSTAT_reg_DO_reg[0]/P0002  & \core_eu_em_mac_em_reg_mr0rwe_DO_reg[11]/P0001  ;
  assign n8353 = \core_c_psq_MSTAT_reg_DO_reg[0]/P0002  & \core_eu_em_mac_em_reg_mr0swe_DO_reg[11]/P0001  ;
  assign n8354 = ~n8352 & ~n8353 ;
  assign n8355 = \core_c_dec_MFMR0_E_reg/P0001  & ~n8354 ;
  assign n8362 = ~n8351 & ~n8355 ;
  assign n8363 = ~n8359 & n8362 ;
  assign n8336 = ~\core_c_psq_MSTAT_reg_DO_reg[0]/P0002  & \core_eu_em_mac_em_reg_my0rwe_DO_reg[11]/P0001  ;
  assign n8337 = \core_c_psq_MSTAT_reg_DO_reg[0]/P0002  & \core_eu_em_mac_em_reg_my0swe_DO_reg[11]/P0001  ;
  assign n8338 = ~n8336 & ~n8337 ;
  assign n8339 = \core_c_dec_MFMY0_E_reg/P0001  & ~n8338 ;
  assign n8360 = ~n7207 & ~n8339 ;
  assign n8340 = ~\core_c_psq_MSTAT_reg_DO_reg[0]/P0002  & \core_eu_em_mac_em_reg_my1rwe_DO_reg[11]/P0001  ;
  assign n8341 = \core_c_psq_MSTAT_reg_DO_reg[0]/P0002  & \core_eu_em_mac_em_reg_my1swe_DO_reg[11]/P0001  ;
  assign n8342 = ~n8340 & ~n8341 ;
  assign n8343 = \core_c_dec_MFMY1_E_reg/P0001  & ~n8342 ;
  assign n8344 = ~\core_c_psq_MSTAT_reg_DO_reg[0]/P0002  & \core_eu_em_mac_em_reg_mx0rwe_DO_reg[11]/P0001  ;
  assign n8345 = \core_c_psq_MSTAT_reg_DO_reg[0]/P0002  & \core_eu_em_mac_em_reg_mx0swe_DO_reg[11]/P0001  ;
  assign n8346 = ~n8344 & ~n8345 ;
  assign n8347 = \core_c_dec_MFMX0_E_reg/P0001  & ~n8346 ;
  assign n8361 = ~n8343 & ~n8347 ;
  assign n8364 = n8360 & n8361 ;
  assign n8365 = n8363 & n8364 ;
  assign n8366 = n7179 & ~n8365 ;
  assign n8367 = ~\core_c_psq_MSTAT_reg_DO_reg[0]/P0002  & \core_eu_ea_alu_ea_reg_ax0rwe_DO_reg[11]/P0001  ;
  assign n8368 = \core_c_psq_MSTAT_reg_DO_reg[0]/P0002  & \core_eu_ea_alu_ea_reg_ax0swe_DO_reg[11]/P0001  ;
  assign n8369 = ~n8367 & ~n8368 ;
  assign n8370 = \core_c_dec_MFAX0_E_reg/P0001  & ~n8369 ;
  assign n8371 = ~\core_c_psq_MSTAT_reg_DO_reg[0]/P0002  & \core_eu_ea_alu_ea_reg_ax1rwe_DO_reg[11]/P0001  ;
  assign n8372 = \core_c_psq_MSTAT_reg_DO_reg[0]/P0002  & \core_eu_ea_alu_ea_reg_ax1swe_DO_reg[11]/P0001  ;
  assign n8373 = ~n8371 & ~n8372 ;
  assign n8374 = \core_c_dec_MFAX1_E_reg/P0001  & ~n8373 ;
  assign n8387 = ~n8370 & ~n8374 ;
  assign n8383 = ~\core_c_psq_MSTAT_reg_DO_reg[0]/P0002  & \core_eu_ea_alu_ea_reg_arrwe_DO_reg[11]/P0001  ;
  assign n8384 = \core_c_psq_MSTAT_reg_DO_reg[0]/P0002  & \core_eu_ea_alu_ea_reg_arswe_DO_reg[11]/P0001  ;
  assign n8385 = ~n8383 & ~n8384 ;
  assign n8386 = \core_c_dec_MFAR_E_reg/P0001  & ~n8385 ;
  assign n8375 = ~\core_c_psq_MSTAT_reg_DO_reg[0]/P0002  & \core_eu_ea_alu_ea_reg_ay0rwe_DO_reg[11]/P0001  ;
  assign n8376 = \core_c_psq_MSTAT_reg_DO_reg[0]/P0002  & \core_eu_ea_alu_ea_reg_ay0swe_DO_reg[11]/P0001  ;
  assign n8377 = ~n8375 & ~n8376 ;
  assign n8378 = \core_c_dec_MFAY0_E_reg/P0001  & ~n8377 ;
  assign n8379 = ~\core_c_psq_MSTAT_reg_DO_reg[0]/P0002  & \core_eu_ea_alu_ea_reg_ay1rwe_DO_reg[11]/P0001  ;
  assign n8380 = \core_c_psq_MSTAT_reg_DO_reg[0]/P0002  & \core_eu_ea_alu_ea_reg_ay1swe_DO_reg[11]/P0001  ;
  assign n8381 = ~n8379 & ~n8380 ;
  assign n8382 = \core_c_dec_MFAY1_E_reg/P0001  & ~n8381 ;
  assign n8388 = ~n8378 & ~n8382 ;
  assign n8389 = ~n8386 & n8388 ;
  assign n8390 = n8387 & n8389 ;
  assign n8391 = n7093 & ~n8390 ;
  assign n8450 = ~n8366 & ~n8391 ;
  assign n8451 = ~n8415 & n8450 ;
  assign n8452 = n8449 & n8451 ;
  assign n8453 = ~n8399 & n8452 ;
  assign n8454 = ~n8335 & n8453 ;
  assign n8455 = ~n8266 & n8454 ;
  assign n8456 = ~\emc_DMDoe_reg/NET0131  & ~n8455 ;
  assign n8457 = \emc_DMDoe_reg/NET0131  & \emc_DMDreg_reg[11]/P0001  ;
  assign n8458 = n7057 & ~n8457 ;
  assign n8459 = ~n8456 & n8458 ;
  assign n8460 = ~n8265 & ~n8459 ;
  assign n8461 = n6135 & ~n8460 ;
  assign n8462 = n6176 & ~n8461 ;
  assign n8463 = ~n8247 & n8462 ;
  assign n8470 = \DM_rd0[2]_pad  & ~n7053 ;
  assign n8464 = \DM_rdm[2]_pad  & n7016 ;
  assign n8475 = ~n7057 & ~n8464 ;
  assign n8467 = \DM_rd6[2]_pad  & n7031 ;
  assign n8468 = \DM_rd7[2]_pad  & n7034 ;
  assign n8476 = ~n8467 & ~n8468 ;
  assign n8477 = n8475 & n8476 ;
  assign n8471 = \DM_rd4[2]_pad  & n7028 ;
  assign n8466 = \DM_rd5[2]_pad  & n7043 ;
  assign n8472 = \DM_rd2[2]_pad  & n7041 ;
  assign n8465 = \DM_rd1[2]_pad  & n7022 ;
  assign n8469 = \DM_rd3[2]_pad  & n7038 ;
  assign n8473 = ~n8465 & ~n8469 ;
  assign n8474 = ~n8472 & n8473 ;
  assign n8478 = ~n8466 & n8474 ;
  assign n8479 = ~n8471 & n8478 ;
  assign n8480 = n8477 & n8479 ;
  assign n8481 = ~n8470 & n8480 ;
  assign n8482 = \regout_STD_C_reg[2]/P0001  & n6988 ;
  assign n8639 = \bdma_BIAD_reg[2]/NET0131  & n7234 ;
  assign n8630 = \emc_WSCRreg_DO_reg[2]/NET0131  & n7251 ;
  assign n8631 = \sport0_regs_SCLKDIVreg_DO_reg[2]/NET0131  & n7256 ;
  assign n8656 = ~n8630 & ~n8631 ;
  assign n8632 = \sport1_regs_MWORDreg_DO_reg[2]/NET0131  & n7263 ;
  assign n8633 = \tm_tsr_reg_DO_reg[2]/NET0131  & n7540 ;
  assign n8657 = ~n8632 & ~n8633 ;
  assign n8670 = n8656 & n8657 ;
  assign n8626 = \idma_DOVL_reg[2]/NET0131  & n7532 ;
  assign n8654 = ~n7522 & ~n8626 ;
  assign n8627 = \sport0_regs_AUTOreg_DO_reg[2]/NET0131  & n7295 ;
  assign n8628 = \tm_tpr_reg_DO_reg[2]/NET0131  & n7293 ;
  assign n8655 = ~n8627 & ~n8628 ;
  assign n8671 = n8654 & n8655 ;
  assign n8672 = n8670 & n8671 ;
  assign n8676 = ~n8639 & n8672 ;
  assign n8647 = \bdma_BEAD_reg[2]/NET0131  & n7303 ;
  assign n8648 = \bdma_BCTL_reg[2]/NET0131  & n7230 ;
  assign n8677 = ~n8647 & ~n8648 ;
  assign n8678 = n8676 & n8677 ;
  assign n8644 = \bdma_BOVL_reg[2]/NET0131  & n7534 ;
  assign n8629 = \bdma_BWCOUNT_reg[2]/NET0131  & n7287 ;
  assign n8638 = \pio_pmask_reg_DO_reg[2]/NET0131  & n7297 ;
  assign n8640 = \sport0_regs_MWORDreg_DO_reg[2]/NET0131  & n7276 ;
  assign n8660 = ~n8638 & ~n8640 ;
  assign n8641 = \sport1_regs_AUTOreg_DO_reg[2]/NET0131  & n7527 ;
  assign n8642 = \tm_TCR_TMP_reg[2]/NET0131  & n7289 ;
  assign n8661 = ~n8641 & ~n8642 ;
  assign n8668 = n8660 & n8661 ;
  assign n8634 = \sport0_regs_SCTLreg_DO_reg[2]/NET0131  & n7249 ;
  assign n8635 = \emc_WSCRext_reg_DO_reg[2]/NET0131  & n7514 ;
  assign n8658 = ~n8634 & ~n8635 ;
  assign n8636 = \sport1_regs_SCLKDIVreg_DO_reg[2]/NET0131  & n7247 ;
  assign n8637 = \sport1_regs_SCTLreg_DO_reg[2]/NET0131  & n7281 ;
  assign n8659 = ~n8636 & ~n8637 ;
  assign n8669 = n8658 & n8659 ;
  assign n8673 = n8668 & n8669 ;
  assign n8650 = \idma_DCTL_reg[2]/NET0131  & n7299 ;
  assign n8651 = \PIO_out[2]_pad  & n7291 ;
  assign n8664 = ~n8650 & ~n8651 ;
  assign n8652 = \PIO_oe[2]_pad  & n7244 ;
  assign n8653 = \sport1_regs_FSDIVreg_DO_reg[2]/NET0131  & n7273 ;
  assign n8665 = ~n8652 & ~n8653 ;
  assign n8666 = n8664 & n8665 ;
  assign n8643 = \sport0_regs_FSDIVreg_DO_reg[2]/NET0131  & n7259 ;
  assign n8645 = \clkc_ckr_reg_DO_reg[2]/NET0131  & n7239 ;
  assign n8662 = ~n8643 & ~n8645 ;
  assign n8646 = \memc_usysr_DO_reg[2]/NET0131  & n7301 ;
  assign n8649 = \pio_PINT_reg[2]/NET0131  & n7271 ;
  assign n8663 = ~n8646 & ~n8649 ;
  assign n8667 = n8662 & n8663 ;
  assign n8674 = n8666 & n8667 ;
  assign n8675 = n8673 & n8674 ;
  assign n8679 = ~n8629 & n8675 ;
  assign n8680 = ~n8644 & n8679 ;
  assign n8681 = n8678 & n8680 ;
  assign n8682 = \memc_ldSREG_E_reg/NET0131  & ~n8681 ;
  assign n8686 = \core_c_dec_MFtoppcs_Eg_reg/P0001  & ~n4521 ;
  assign n8689 = \core_c_dec_MFMSTAT_E_reg/P0001  & \core_c_psq_MSTAT_reg_DO_reg[2]/NET0131  ;
  assign n8690 = \core_c_dec_MFSSTAT_E_reg/P0001  & \core_c_psq_SSTAT_reg[2]/NET0131  ;
  assign n8695 = ~n8689 & ~n8690 ;
  assign n8691 = \core_c_dec_MFCNTR_E_reg/P0001  & \core_c_psq_CNTR_reg_DO_reg[2]/NET0131  ;
  assign n8692 = \core_c_dec_MFICNTL_E_reg/P0001  & \core_c_psq_ICNTL_reg_DO_reg[2]/NET0131  ;
  assign n8696 = ~n8691 & ~n8692 ;
  assign n8697 = n8695 & n8696 ;
  assign n8687 = \core_c_dec_IRE_reg[6]/NET0131  & ~n7216 ;
  assign n8683 = \core_c_dec_MFIDR_E_reg/P0001  & \sice_idr0_reg_DO_reg[2]/P0001  ;
  assign n8684 = \core_c_dec_MFIMASK_E_reg/P0001  & \core_c_psq_IMASK_reg[2]/NET0131  ;
  assign n8693 = ~n8683 & ~n8684 ;
  assign n8685 = \core_c_dec_MFPMOVL_E_reg/P0001  & \core_c_psq_PMOVL_regl_DO_reg[2]/NET0131  ;
  assign n8688 = \core_c_dec_MFDMOVL_E_reg/P0001  & \core_c_psq_DMOVL_reg_DO_reg[2]/NET0131  ;
  assign n8694 = ~n8685 & ~n8688 ;
  assign n8698 = n8693 & n8694 ;
  assign n8699 = ~n8687 & n8698 ;
  assign n8700 = n8697 & n8699 ;
  assign n8701 = ~n8686 & n8700 ;
  assign n8702 = n7215 & ~n8701 ;
  assign n8610 = \core_c_dec_MFIreg_E_reg[7]/P0001  & \core_dag_ilm2reg_I7_we_DO_reg[2]/NET0131  ;
  assign n8611 = \core_c_dec_MFIreg_E_reg[4]/P0001  & \core_dag_ilm2reg_I4_we_DO_reg[2]/NET0131  ;
  assign n8618 = ~n8610 & ~n8611 ;
  assign n8612 = \core_c_dec_MFIreg_E_reg[5]/P0001  & \core_dag_ilm2reg_I5_we_DO_reg[2]/NET0131  ;
  assign n8613 = \core_c_dec_MFIreg_E_reg[6]/P0001  & \core_dag_ilm2reg_I6_we_DO_reg[2]/NET0131  ;
  assign n8619 = ~n8612 & ~n8613 ;
  assign n8620 = n8618 & n8619 ;
  assign n8606 = \core_c_dec_MFLreg_E_reg[4]/P0001  & \core_dag_ilm2reg_L4_we_DO_reg[2]/NET0131  ;
  assign n8607 = \core_c_dec_MFLreg_E_reg[5]/P0001  & \core_dag_ilm2reg_L5_we_DO_reg[2]/NET0131  ;
  assign n8616 = ~n8606 & ~n8607 ;
  assign n8608 = \core_c_dec_MFMreg_E_reg[6]/P0001  & \core_dag_ilm2reg_M6_we_DO_reg[2]/NET0131  ;
  assign n8609 = \core_c_dec_MFMreg_E_reg[7]/P0001  & \core_dag_ilm2reg_M7_we_DO_reg[2]/NET0131  ;
  assign n8617 = ~n8608 & ~n8609 ;
  assign n8621 = n8616 & n8617 ;
  assign n8602 = \core_c_dec_MFMreg_E_reg[5]/P0001  & \core_dag_ilm2reg_M5_we_DO_reg[2]/NET0131  ;
  assign n8603 = \core_c_dec_MFLreg_E_reg[6]/P0001  & \core_dag_ilm2reg_L6_we_DO_reg[2]/NET0131  ;
  assign n8614 = ~n8602 & ~n8603 ;
  assign n8604 = \core_c_dec_MFLreg_E_reg[7]/P0001  & \core_dag_ilm2reg_L7_we_DO_reg[2]/NET0131  ;
  assign n8605 = \core_c_dec_MFMreg_E_reg[4]/P0001  & \core_dag_ilm2reg_M4_we_DO_reg[2]/NET0131  ;
  assign n8615 = ~n8604 & ~n8605 ;
  assign n8622 = n8614 & n8615 ;
  assign n8623 = n8621 & n8622 ;
  assign n8624 = n8620 & n8623 ;
  assign n8625 = n7128 & ~n8624 ;
  assign n8516 = \core_c_dec_MFMreg_E_reg[1]/P0001  & \core_dag_ilm1reg_M1_we_DO_reg[2]/NET0131  ;
  assign n8517 = \core_c_dec_MFLreg_E_reg[2]/P0001  & \core_dag_ilm1reg_L2_we_DO_reg[2]/NET0131  ;
  assign n8524 = ~n8516 & ~n8517 ;
  assign n8518 = \core_c_dec_MFLreg_E_reg[3]/P0001  & \core_dag_ilm1reg_L3_we_DO_reg[2]/NET0131  ;
  assign n8519 = \core_c_dec_MFMreg_E_reg[0]/P0001  & \core_dag_ilm1reg_M0_we_DO_reg[2]/NET0131  ;
  assign n8525 = ~n8518 & ~n8519 ;
  assign n8526 = n8524 & n8525 ;
  assign n8512 = \core_c_dec_MFMreg_E_reg[2]/P0001  & \core_dag_ilm1reg_M2_we_DO_reg[2]/NET0131  ;
  assign n8513 = \core_c_dec_MFMreg_E_reg[3]/P0001  & \core_dag_ilm1reg_M3_we_DO_reg[2]/NET0131  ;
  assign n8522 = ~n8512 & ~n8513 ;
  assign n8514 = \core_c_dec_MFIreg_E_reg[1]/P0001  & \core_dag_ilm1reg_I1_we_DO_reg[2]/NET0131  ;
  assign n8515 = \core_c_dec_MFIreg_E_reg[2]/P0001  & \core_dag_ilm1reg_I2_we_DO_reg[2]/NET0131  ;
  assign n8523 = ~n8514 & ~n8515 ;
  assign n8527 = n8522 & n8523 ;
  assign n8508 = \core_c_dec_MFIreg_E_reg[0]/P0001  & \core_dag_ilm1reg_I0_we_DO_reg[2]/NET0131  ;
  assign n8509 = \core_c_dec_MFIreg_E_reg[3]/P0001  & \core_dag_ilm1reg_I3_we_DO_reg[2]/NET0131  ;
  assign n8520 = ~n8508 & ~n8509 ;
  assign n8510 = \core_c_dec_MFLreg_E_reg[0]/P0001  & \core_dag_ilm1reg_L0_we_DO_reg[2]/NET0131  ;
  assign n8511 = \core_c_dec_MFLreg_E_reg[1]/P0001  & \core_dag_ilm1reg_L1_we_DO_reg[2]/NET0131  ;
  assign n8521 = ~n8510 & ~n8511 ;
  assign n8528 = n8520 & n8521 ;
  assign n8529 = n8527 & n8528 ;
  assign n8530 = n8526 & n8529 ;
  assign n8531 = n7068 & ~n8530 ;
  assign n8567 = \core_c_dec_MFTX1_E_reg/P0001  & \sport1_txctl_TX_reg[2]/P0001  ;
  assign n8568 = \core_c_dec_MFTX0_E_reg/P0001  & \sport0_txctl_TX_reg[2]/P0001  ;
  assign n8571 = ~n8567 & ~n8568 ;
  assign n8569 = \core_c_dec_MFRX1_E_reg/P0001  & \sport1_rxctl_RX_reg[2]/P0001  ;
  assign n8570 = \core_c_dec_MFRX0_E_reg/P0001  & \sport0_rxctl_RX_reg[2]/P0001  ;
  assign n8572 = ~n8569 & ~n8570 ;
  assign n8573 = n8571 & n8572 ;
  assign n8574 = n7119 & ~n8573 ;
  assign n8703 = ~n8531 & ~n8574 ;
  assign n8704 = ~n8625 & n8703 ;
  assign n8575 = ~\core_c_psq_MSTAT_reg_DO_reg[0]/P0002  & \core_eu_ea_alu_ea_reg_ay0rwe_DO_reg[2]/P0001  ;
  assign n8576 = \core_c_psq_MSTAT_reg_DO_reg[0]/P0002  & \core_eu_ea_alu_ea_reg_ay0swe_DO_reg[2]/P0001  ;
  assign n8577 = ~n8575 & ~n8576 ;
  assign n8578 = \core_c_dec_MFAY0_E_reg/P0001  & ~n8577 ;
  assign n8595 = \core_c_dec_MFASTAT_E_reg/P0001  & \core_eu_ec_cun_AV_reg/P0001  ;
  assign n8596 = ~n8578 & ~n8595 ;
  assign n8579 = ~\core_c_psq_MSTAT_reg_DO_reg[0]/P0002  & \core_eu_ea_alu_ea_reg_ay1rwe_DO_reg[2]/P0001  ;
  assign n8580 = \core_c_psq_MSTAT_reg_DO_reg[0]/P0002  & \core_eu_ea_alu_ea_reg_ay1swe_DO_reg[2]/P0001  ;
  assign n8581 = ~n8579 & ~n8580 ;
  assign n8582 = \core_c_dec_MFAY1_E_reg/P0001  & ~n8581 ;
  assign n8583 = ~\core_c_psq_MSTAT_reg_DO_reg[0]/P0002  & \core_eu_ea_alu_ea_reg_arrwe_DO_reg[2]/P0001  ;
  assign n8584 = \core_c_psq_MSTAT_reg_DO_reg[0]/P0002  & \core_eu_ea_alu_ea_reg_arswe_DO_reg[2]/P0001  ;
  assign n8585 = ~n8583 & ~n8584 ;
  assign n8586 = \core_c_dec_MFAR_E_reg/P0001  & ~n8585 ;
  assign n8597 = ~n8582 & ~n8586 ;
  assign n8587 = ~\core_c_psq_MSTAT_reg_DO_reg[0]/P0002  & \core_eu_ea_alu_ea_reg_ax1rwe_DO_reg[2]/P0001  ;
  assign n8588 = \core_c_psq_MSTAT_reg_DO_reg[0]/P0002  & \core_eu_ea_alu_ea_reg_ax1swe_DO_reg[2]/P0001  ;
  assign n8589 = ~n8587 & ~n8588 ;
  assign n8590 = \core_c_dec_MFAX1_E_reg/P0001  & ~n8589 ;
  assign n8591 = ~\core_c_psq_MSTAT_reg_DO_reg[0]/P0002  & \core_eu_ea_alu_ea_reg_ax0rwe_DO_reg[2]/P0001  ;
  assign n8592 = \core_c_psq_MSTAT_reg_DO_reg[0]/P0002  & \core_eu_ea_alu_ea_reg_ax0swe_DO_reg[2]/P0001  ;
  assign n8593 = ~n8591 & ~n8592 ;
  assign n8594 = \core_c_dec_MFAX0_E_reg/P0001  & ~n8593 ;
  assign n8598 = ~n8590 & ~n8594 ;
  assign n8599 = n8597 & n8598 ;
  assign n8600 = n8596 & n8599 ;
  assign n8601 = n7093 & ~n8600 ;
  assign n8483 = ~\core_c_psq_MSTAT_reg_DO_reg[0]/P0002  & \core_eu_es_sht_es_reg_sirwe_DO_reg[2]/P0001  ;
  assign n8484 = \core_c_psq_MSTAT_reg_DO_reg[0]/P0002  & \core_eu_es_sht_es_reg_siswe_DO_reg[2]/P0001  ;
  assign n8485 = ~n8483 & ~n8484 ;
  assign n8486 = \core_c_dec_MFSI_E_reg/P0001  & ~n8485 ;
  assign n8487 = ~\core_c_psq_MSTAT_reg_DO_reg[0]/P0002  & \core_eu_es_sht_es_reg_SBr_reg[2]/P0001  ;
  assign n8488 = \core_c_psq_MSTAT_reg_DO_reg[0]/P0002  & \core_eu_es_sht_es_reg_SBs_reg[2]/P0001  ;
  assign n8489 = ~n8487 & ~n8488 ;
  assign n8490 = \core_c_dec_MFSB_E_reg/P0001  & ~n8489 ;
  assign n8503 = ~n8486 & ~n8490 ;
  assign n8499 = ~\core_c_psq_MSTAT_reg_DO_reg[0]/P0002  & \core_eu_es_sht_es_reg_serwe_DO_reg[2]/P0001  ;
  assign n8500 = \core_c_psq_MSTAT_reg_DO_reg[0]/P0002  & \core_eu_es_sht_es_reg_seswe_DO_reg[2]/P0001  ;
  assign n8501 = ~n8499 & ~n8500 ;
  assign n8502 = \core_c_dec_MFSE_E_reg/P0001  & ~n8501 ;
  assign n8491 = ~\core_c_psq_MSTAT_reg_DO_reg[0]/P0002  & \core_eu_es_sht_es_reg_sr0rwe_DO_reg[2]/P0001  ;
  assign n8492 = \core_c_psq_MSTAT_reg_DO_reg[0]/P0002  & \core_eu_es_sht_es_reg_sr0swe_DO_reg[2]/P0001  ;
  assign n8493 = ~n8491 & ~n8492 ;
  assign n8494 = \core_c_dec_MFSR0_E_reg/P0001  & ~n8493 ;
  assign n8495 = ~\core_c_psq_MSTAT_reg_DO_reg[0]/P0002  & \core_eu_es_sht_es_reg_sr1rwe_DO_reg[2]/P0001  ;
  assign n8496 = \core_c_psq_MSTAT_reg_DO_reg[0]/P0002  & \core_eu_es_sht_es_reg_sr1swe_DO_reg[2]/P0001  ;
  assign n8497 = ~n8495 & ~n8496 ;
  assign n8498 = \core_c_dec_MFSR1_E_reg/P0001  & ~n8497 ;
  assign n8504 = ~n8494 & ~n8498 ;
  assign n8505 = ~n8502 & n8504 ;
  assign n8506 = n8503 & n8505 ;
  assign n8507 = n7153 & ~n8506 ;
  assign n8556 = ~\core_c_psq_MSTAT_reg_DO_reg[0]/P0002  & \core_eu_em_mac_em_reg_mr1rwe_DO_reg[2]/P0001  ;
  assign n8557 = \core_c_psq_MSTAT_reg_DO_reg[0]/P0002  & \core_eu_em_mac_em_reg_mr1swe_DO_reg[2]/P0001  ;
  assign n8558 = ~n8556 & ~n8557 ;
  assign n8559 = \core_c_dec_MFMR1_E_reg/P0001  & ~n8558 ;
  assign n8548 = ~\core_c_psq_MSTAT_reg_DO_reg[0]/P0002  & \core_eu_em_mac_em_reg_mx0rwe_DO_reg[2]/P0001  ;
  assign n8549 = \core_c_psq_MSTAT_reg_DO_reg[0]/P0002  & \core_eu_em_mac_em_reg_mx0swe_DO_reg[2]/P0001  ;
  assign n8550 = ~n8548 & ~n8549 ;
  assign n8551 = \core_c_dec_MFMX0_E_reg/P0001  & ~n8550 ;
  assign n8552 = ~\core_c_psq_MSTAT_reg_DO_reg[0]/P0002  & \core_eu_em_mac_em_reg_mr0rwe_DO_reg[2]/P0001  ;
  assign n8553 = \core_c_psq_MSTAT_reg_DO_reg[0]/P0002  & \core_eu_em_mac_em_reg_mr0swe_DO_reg[2]/P0001  ;
  assign n8554 = ~n8552 & ~n8553 ;
  assign n8555 = \core_c_dec_MFMR0_E_reg/P0001  & ~n8554 ;
  assign n8562 = ~n8551 & ~n8555 ;
  assign n8563 = ~n8559 & n8562 ;
  assign n8532 = ~\core_c_psq_MSTAT_reg_DO_reg[0]/P0002  & \core_eu_em_mac_em_reg_mr2rwe_DO_reg[2]/P0001  ;
  assign n8533 = \core_c_psq_MSTAT_reg_DO_reg[0]/P0002  & \core_eu_em_mac_em_reg_mr2swe_DO_reg[2]/P0001  ;
  assign n8534 = ~n8532 & ~n8533 ;
  assign n8535 = \core_c_dec_MFMR2_E_reg/P0001  & ~n8534 ;
  assign n8536 = ~\core_c_psq_MSTAT_reg_DO_reg[0]/P0002  & \core_eu_em_mac_em_reg_mx1rwe_DO_reg[2]/P0001  ;
  assign n8537 = \core_c_psq_MSTAT_reg_DO_reg[0]/P0002  & \core_eu_em_mac_em_reg_mx1swe_DO_reg[2]/P0001  ;
  assign n8538 = ~n8536 & ~n8537 ;
  assign n8539 = \core_c_dec_MFMX1_E_reg/P0001  & ~n8538 ;
  assign n8560 = ~n8535 & ~n8539 ;
  assign n8540 = ~\core_c_psq_MSTAT_reg_DO_reg[0]/P0002  & \core_eu_em_mac_em_reg_my1rwe_DO_reg[2]/P0001  ;
  assign n8541 = \core_c_psq_MSTAT_reg_DO_reg[0]/P0002  & \core_eu_em_mac_em_reg_my1swe_DO_reg[2]/P0001  ;
  assign n8542 = ~n8540 & ~n8541 ;
  assign n8543 = \core_c_dec_MFMY1_E_reg/P0001  & ~n8542 ;
  assign n8544 = ~\core_c_psq_MSTAT_reg_DO_reg[0]/P0002  & \core_eu_em_mac_em_reg_my0rwe_DO_reg[2]/P0001  ;
  assign n8545 = \core_c_psq_MSTAT_reg_DO_reg[0]/P0002  & \core_eu_em_mac_em_reg_my0swe_DO_reg[2]/P0001  ;
  assign n8546 = ~n8544 & ~n8545 ;
  assign n8547 = \core_c_dec_MFMY0_E_reg/P0001  & ~n8546 ;
  assign n8561 = ~n8543 & ~n8547 ;
  assign n8564 = n8560 & n8561 ;
  assign n8565 = n8563 & n8564 ;
  assign n8566 = n7179 & ~n8565 ;
  assign n8705 = ~n8507 & ~n8566 ;
  assign n8706 = ~n8601 & n8705 ;
  assign n8707 = n8704 & n8706 ;
  assign n8708 = ~n8702 & n8707 ;
  assign n8709 = ~n8682 & n8708 ;
  assign n8710 = ~n8482 & n8709 ;
  assign n8711 = ~\emc_DMDoe_reg/NET0131  & ~n8710 ;
  assign n8712 = \emc_DMDoe_reg/NET0131  & \emc_DMDreg_reg[2]/P0001  ;
  assign n8713 = n7057 & ~n8712 ;
  assign n8714 = ~n8711 & n8713 ;
  assign n8715 = ~n8481 & ~n8714 ;
  assign n8716 = n7863 & n8715 ;
  assign n8717 = \core_dag_ilm2reg_I4_we_DO_reg[11]/NET0131  & n6976 ;
  assign n8718 = \core_dag_ilm2reg_I5_we_DO_reg[11]/NET0131  & n6970 ;
  assign n8721 = ~n8717 & ~n8718 ;
  assign n8719 = \core_dag_ilm2reg_I6_we_DO_reg[11]/NET0131  & n6974 ;
  assign n8720 = \core_dag_ilm2reg_I7_we_DO_reg[11]/NET0131  & n6972 ;
  assign n8722 = ~n8719 & ~n8720 ;
  assign n8723 = n8721 & n8722 ;
  assign n8724 = n4055 & ~n8723 ;
  assign n8725 = \core_dag_ilm2reg_I4_we_DO_reg[11]/NET0131  & n6958 ;
  assign n8726 = \core_dag_ilm2reg_I5_we_DO_reg[11]/NET0131  & n6964 ;
  assign n8729 = ~n8725 & ~n8726 ;
  assign n8727 = \core_dag_ilm2reg_I6_we_DO_reg[11]/NET0131  & n6962 ;
  assign n8728 = \core_dag_ilm2reg_I7_we_DO_reg[11]/NET0131  & n6960 ;
  assign n8730 = ~n8727 & ~n8728 ;
  assign n8731 = n8729 & n8730 ;
  assign n8732 = ~n8724 & n8731 ;
  assign n8733 = \core_dag_ilm1reg_I0_we_DO_reg[11]/NET0131  & n8131 ;
  assign n8740 = ~n4055 & ~n8733 ;
  assign n8738 = \core_dag_ilm1reg_I3_we_DO_reg[11]/NET0131  & n6075 ;
  assign n8739 = n6077 & n8738 ;
  assign n8734 = \core_dag_ilm1reg_I2_we_DO_reg[11]/NET0131  & n6084 ;
  assign n8735 = n6085 & n8734 ;
  assign n8736 = \core_dag_ilm1reg_I1_we_DO_reg[11]/NET0131  & n6067 ;
  assign n8737 = n6068 & n8736 ;
  assign n8741 = ~n8735 & ~n8737 ;
  assign n8742 = ~n8739 & n8741 ;
  assign n8743 = n8740 & n8742 ;
  assign n8744 = n6097 & n8738 ;
  assign n8745 = n6095 & n8734 ;
  assign n8748 = ~n8744 & ~n8745 ;
  assign n8746 = n6091 & n8736 ;
  assign n8747 = \core_dag_ilm1reg_I0_we_DO_reg[11]/NET0131  & n6148 ;
  assign n8749 = ~n8746 & ~n8747 ;
  assign n8750 = n8748 & n8749 ;
  assign n8751 = n4055 & n8750 ;
  assign n8752 = ~n8743 & ~n8751 ;
  assign n8753 = n8732 & ~n8752 ;
  assign n8754 = n8153 & ~n8753 ;
  assign n8755 = ~n8716 & ~n8754 ;
  assign n8756 = ~n8463 & n8755 ;
  assign n8757 = n7005 & ~n8756 ;
  assign n8805 = ~n6867 & ~n6877 ;
  assign n8806 = ~n6857 & ~n8204 ;
  assign n8807 = ~n6870 & ~n8806 ;
  assign n8808 = n8805 & ~n8807 ;
  assign n8809 = ~n8805 & n8807 ;
  assign n8810 = ~n8808 & ~n8809 ;
  assign n8811 = n8198 & n8810 ;
  assign n8798 = \core_dag_ilm2reg_I_reg[11]/NET0131  & ~n6624 ;
  assign n8799 = ~n6702 & n8199 ;
  assign n8800 = ~n6622 & ~n8799 ;
  assign n8801 = ~n6860 & ~n8800 ;
  assign n8802 = n6860 & n8800 ;
  assign n8803 = ~n8801 & ~n8802 ;
  assign n8804 = ~n8198 & n8803 ;
  assign n8812 = ~n8798 & ~n8804 ;
  assign n8813 = ~n8811 & n8812 ;
  assign n8814 = n6135 & ~n8813 ;
  assign n8820 = ~n6121 & ~n8732 ;
  assign n8818 = ~n6111 & n8752 ;
  assign n8819 = \core_c_dec_IR_reg[15]/NET0131  & n6956 ;
  assign n8821 = ~n8818 & ~n8819 ;
  assign n8822 = ~n8820 & n8821 ;
  assign n8823 = n5949 & ~n8822 ;
  assign n8824 = \core_dag_ilm1reg_DMA_pi_DO_reg[11]/NET0131  & ~n6934 ;
  assign n8816 = \core_dag_ilm1reg_STAC_pi_DO_reg[11]/NET0131  & n6988 ;
  assign n8817 = \idma_DCTL_reg[11]/NET0131  & n6926 ;
  assign n8825 = ~n8816 & ~n8817 ;
  assign n8826 = n6924 & n8825 ;
  assign n8827 = ~n8824 & n8826 ;
  assign n8828 = ~n8823 & n8827 ;
  assign n8815 = ~\bdma_BIAD_reg[11]/NET0131  & ~n6924 ;
  assign n8829 = ~n6135 & ~n8815 ;
  assign n8830 = ~n8828 & n8829 ;
  assign n8831 = ~n6176 & ~n8830 ;
  assign n8832 = ~n8814 & n8831 ;
  assign n8783 = n6339 & ~n6501 ;
  assign n8784 = ~n6339 & n6501 ;
  assign n8785 = ~n8783 & ~n8784 ;
  assign n8786 = ~n6496 & n8785 ;
  assign n8778 = ~n6343 & ~n6344 ;
  assign n8779 = n6368 & n8778 ;
  assign n8780 = ~n6368 & ~n8778 ;
  assign n8781 = ~n8779 & ~n8780 ;
  assign n8782 = n6496 & ~n8781 ;
  assign n8787 = ~\core_dag_ilm1reg_M_reg[13]/NET0131  & ~n8782 ;
  assign n8788 = ~n8786 & n8787 ;
  assign n8777 = \core_dag_ilm1reg_I_reg[2]/NET0131  & ~n6317 ;
  assign n8790 = n7612 & n8785 ;
  assign n8789 = ~n7612 & ~n8781 ;
  assign n8791 = \core_dag_ilm1reg_M_reg[13]/NET0131  & ~n8789 ;
  assign n8792 = ~n8790 & n8791 ;
  assign n8793 = ~n8777 & ~n8792 ;
  assign n8794 = ~n8788 & n8793 ;
  assign n8795 = n6135 & ~n8794 ;
  assign n8758 = \core_dag_ilm1reg_I2_we_DO_reg[2]/NET0131  & n6138 ;
  assign n8762 = ~n4055 & ~n8758 ;
  assign n8761 = \core_dag_ilm1reg_I1_we_DO_reg[2]/NET0131  & n6142 ;
  assign n8759 = \core_dag_ilm1reg_I0_we_DO_reg[2]/NET0131  & n8131 ;
  assign n8760 = \core_dag_ilm1reg_I3_we_DO_reg[2]/NET0131  & n6140 ;
  assign n8763 = ~n8759 & ~n8760 ;
  assign n8764 = ~n8761 & n8763 ;
  assign n8765 = n8762 & n8764 ;
  assign n8766 = \core_dag_ilm1reg_I2_we_DO_reg[2]/NET0131  & n6084 ;
  assign n8767 = n6095 & n8766 ;
  assign n8768 = \core_dag_ilm1reg_I1_we_DO_reg[2]/NET0131  & n6154 ;
  assign n8771 = ~n8767 & ~n8768 ;
  assign n8769 = \core_dag_ilm1reg_I0_we_DO_reg[2]/NET0131  & n6148 ;
  assign n8770 = \core_dag_ilm1reg_I3_we_DO_reg[2]/NET0131  & n6150 ;
  assign n8772 = ~n8769 & ~n8770 ;
  assign n8773 = n8771 & n8772 ;
  assign n8774 = n4055 & n8773 ;
  assign n8775 = ~n8765 & ~n8774 ;
  assign n8776 = ~n6135 & n8775 ;
  assign n8796 = n6176 & ~n8776 ;
  assign n8797 = ~n8795 & n8796 ;
  assign n8833 = ~n7005 & ~n8797 ;
  assign n8834 = ~n8832 & n8833 ;
  assign n8835 = ~n8757 & ~n8834 ;
  assign n8928 = ~n6710 & n6891 ;
  assign n8929 = n6710 & ~n6891 ;
  assign n8930 = ~n8928 & ~n8929 ;
  assign n8931 = ~n6717 & ~n8930 ;
  assign n8932 = ~n6895 & ~n6899 ;
  assign n8933 = n6880 & n8932 ;
  assign n8934 = ~n6880 & ~n8932 ;
  assign n8935 = ~n8933 & ~n8934 ;
  assign n8936 = n6713 & n8935 ;
  assign n8937 = \core_dag_ilm2reg_M_reg[13]/NET0131  & ~n8936 ;
  assign n8938 = ~n8931 & n8937 ;
  assign n8939 = \core_dag_ilm2reg_I_reg[12]/NET0131  & ~n6613 ;
  assign n8941 = ~n6905 & ~n8930 ;
  assign n8940 = n6905 & n8935 ;
  assign n8942 = ~\core_dag_ilm2reg_M_reg[13]/NET0131  & ~n8940 ;
  assign n8943 = ~n8941 & n8942 ;
  assign n8944 = ~n8939 & ~n8943 ;
  assign n8945 = ~n8938 & n8944 ;
  assign n8946 = ~n6176 & ~n8945 ;
  assign n8910 = n6350 & ~n6356 ;
  assign n8911 = ~n6350 & n6356 ;
  assign n8912 = ~n8910 & ~n8911 ;
  assign n8922 = ~n6496 & n8912 ;
  assign n8914 = ~n6360 & ~n6361 ;
  assign n8918 = n6365 & ~n8914 ;
  assign n8919 = ~n6365 & n8914 ;
  assign n8920 = ~n8918 & ~n8919 ;
  assign n8921 = n6496 & n8920 ;
  assign n8923 = ~\core_dag_ilm1reg_M_reg[13]/NET0131  & ~n8921 ;
  assign n8924 = ~n8922 & n8923 ;
  assign n8909 = \core_dag_ilm1reg_I_reg[1]/NET0131  & n6329 ;
  assign n8915 = ~n7612 & ~n8914 ;
  assign n8913 = n7612 & n8912 ;
  assign n8916 = \core_dag_ilm1reg_M_reg[13]/NET0131  & ~n8913 ;
  assign n8917 = ~n8915 & n8916 ;
  assign n8925 = ~n8909 & ~n8917 ;
  assign n8926 = ~n8924 & n8925 ;
  assign n8927 = n6176 & ~n8926 ;
  assign n8947 = n6135 & ~n8927 ;
  assign n8948 = ~n8946 & n8947 ;
  assign n8857 = \core_dag_ilm1reg_I2_we_DO_reg[12]/NET0131  & n6138 ;
  assign n8862 = ~n4055 & ~n8857 ;
  assign n8861 = \core_dag_ilm1reg_I1_we_DO_reg[12]/NET0131  & n6142 ;
  assign n8858 = \core_dag_ilm1reg_I3_we_DO_reg[12]/NET0131  & n6140 ;
  assign n8859 = \core_dag_ilm1reg_I0_we_DO_reg[12]/NET0131  & n6058 ;
  assign n8860 = n6060 & n8859 ;
  assign n8863 = ~n8858 & ~n8860 ;
  assign n8864 = ~n8861 & n8863 ;
  assign n8865 = n8862 & n8864 ;
  assign n8866 = \core_dag_ilm1reg_I0_we_DO_reg[12]/NET0131  & n6148 ;
  assign n8867 = \core_dag_ilm1reg_I1_we_DO_reg[12]/NET0131  & n6154 ;
  assign n8871 = ~n8866 & ~n8867 ;
  assign n8868 = \core_dag_ilm1reg_I2_we_DO_reg[12]/NET0131  & n6152 ;
  assign n8869 = \core_dag_ilm1reg_I3_we_DO_reg[12]/NET0131  & n6075 ;
  assign n8870 = n6097 & n8869 ;
  assign n8872 = ~n8868 & ~n8870 ;
  assign n8873 = n8871 & n8872 ;
  assign n8874 = n4055 & n8873 ;
  assign n8875 = ~n8865 & ~n8874 ;
  assign n8876 = ~n6111 & n8875 ;
  assign n8839 = \core_dag_ilm2reg_I4_we_DO_reg[12]/NET0131  & n6976 ;
  assign n8840 = \core_dag_ilm2reg_I5_we_DO_reg[12]/NET0131  & n6970 ;
  assign n8843 = ~n8839 & ~n8840 ;
  assign n8841 = \core_dag_ilm2reg_I6_we_DO_reg[12]/NET0131  & n6974 ;
  assign n8842 = \core_dag_ilm2reg_I7_we_DO_reg[12]/NET0131  & n6972 ;
  assign n8844 = ~n8841 & ~n8842 ;
  assign n8845 = n8843 & n8844 ;
  assign n8846 = n4055 & ~n8845 ;
  assign n8847 = \core_dag_ilm2reg_I7_we_DO_reg[12]/NET0131  & n6960 ;
  assign n8848 = \core_dag_ilm2reg_I4_we_DO_reg[12]/NET0131  & n6958 ;
  assign n8851 = ~n8847 & ~n8848 ;
  assign n8849 = \core_dag_ilm2reg_I6_we_DO_reg[12]/NET0131  & n6962 ;
  assign n8850 = \core_dag_ilm2reg_I5_we_DO_reg[12]/NET0131  & n6964 ;
  assign n8852 = ~n8849 & ~n8850 ;
  assign n8853 = n8851 & n8852 ;
  assign n8854 = ~n8846 & n8853 ;
  assign n8855 = ~n6121 & ~n8854 ;
  assign n8856 = \core_c_dec_IR_reg[16]/NET0131  & n6956 ;
  assign n8877 = ~n8855 & ~n8856 ;
  assign n8878 = ~n8876 & n8877 ;
  assign n8879 = n5949 & ~n8878 ;
  assign n8880 = \core_dag_ilm1reg_DMA_pi_DO_reg[12]/NET0131  & ~n6934 ;
  assign n8837 = \idma_DCTL_reg[12]/NET0131  & n6926 ;
  assign n8838 = \core_dag_ilm1reg_STAC_pi_DO_reg[12]/NET0131  & n6988 ;
  assign n8881 = ~n8837 & ~n8838 ;
  assign n8882 = n6924 & n8881 ;
  assign n8883 = ~n8880 & n8882 ;
  assign n8884 = ~n8879 & n8883 ;
  assign n8836 = ~\bdma_BIAD_reg[12]/NET0131  & ~n6924 ;
  assign n8885 = ~n6176 & ~n8836 ;
  assign n8886 = ~n8884 & n8885 ;
  assign n8887 = \core_dag_ilm1reg_I3_we_DO_reg[1]/NET0131  & n6140 ;
  assign n8893 = ~n4055 & ~n8887 ;
  assign n8891 = \core_dag_ilm1reg_I1_we_DO_reg[1]/NET0131  & n6067 ;
  assign n8892 = n6068 & n8891 ;
  assign n8888 = \core_dag_ilm1reg_I0_we_DO_reg[1]/NET0131  & n6058 ;
  assign n8889 = n6060 & n8888 ;
  assign n8890 = \core_dag_ilm1reg_I2_we_DO_reg[1]/NET0131  & n6138 ;
  assign n8894 = ~n8889 & ~n8890 ;
  assign n8895 = ~n8892 & n8894 ;
  assign n8896 = n8893 & n8895 ;
  assign n8897 = \core_dag_ilm1reg_I1_we_DO_reg[1]/NET0131  & n6154 ;
  assign n8898 = \core_dag_ilm1reg_I3_we_DO_reg[1]/NET0131  & n6150 ;
  assign n8901 = ~n8897 & ~n8898 ;
  assign n8899 = \core_dag_ilm1reg_I2_we_DO_reg[1]/NET0131  & n6152 ;
  assign n8900 = n6093 & n8888 ;
  assign n8902 = ~n8899 & ~n8900 ;
  assign n8903 = n8901 & n8902 ;
  assign n8904 = n4055 & n8903 ;
  assign n8905 = ~n8896 & ~n8904 ;
  assign n8906 = n6176 & n8905 ;
  assign n8907 = ~n6135 & ~n8906 ;
  assign n8908 = ~n8886 & n8907 ;
  assign n8949 = ~n7005 & ~n8908 ;
  assign n8950 = ~n8948 & n8949 ;
  assign n8956 = ~n6486 & ~n6490 ;
  assign n8957 = n6465 & ~n8956 ;
  assign n8958 = ~n6465 & n8956 ;
  assign n8959 = ~n8957 & ~n8958 ;
  assign n8960 = ~n7631 & n8959 ;
  assign n8951 = \core_dag_ilm1reg_I_reg[12]/NET0131  & ~n6470 ;
  assign n8952 = ~n6482 & ~n6525 ;
  assign n8953 = n6482 & n6525 ;
  assign n8954 = ~n8952 & ~n8953 ;
  assign n8955 = n7631 & ~n8954 ;
  assign n8961 = ~n8951 & ~n8955 ;
  assign n8962 = ~n8960 & n8961 ;
  assign n8963 = ~n6135 & n8962 ;
  assign n8964 = n6176 & n7005 ;
  assign n8971 = \DM_rd0[12]_pad  & ~n7053 ;
  assign n8965 = \DM_rdm[12]_pad  & n7016 ;
  assign n8976 = ~n7057 & ~n8965 ;
  assign n8968 = \DM_rd6[12]_pad  & n7031 ;
  assign n8969 = \DM_rd7[12]_pad  & n7034 ;
  assign n8977 = ~n8968 & ~n8969 ;
  assign n8978 = n8976 & n8977 ;
  assign n8972 = \DM_rd5[12]_pad  & n7043 ;
  assign n8967 = \DM_rd4[12]_pad  & n7028 ;
  assign n8973 = \DM_rd2[12]_pad  & n7041 ;
  assign n8966 = \DM_rd1[12]_pad  & n7022 ;
  assign n8970 = \DM_rd3[12]_pad  & n7038 ;
  assign n8974 = ~n8966 & ~n8970 ;
  assign n8975 = ~n8973 & n8974 ;
  assign n8979 = ~n8967 & n8975 ;
  assign n8980 = ~n8972 & n8979 ;
  assign n8981 = n8978 & n8980 ;
  assign n8982 = ~n8971 & n8981 ;
  assign n8983 = \regout_STD_C_reg[12]/P0001  & n6988 ;
  assign n9113 = \core_c_dec_MFtoppcs_Eg_reg/P0001  & ~n4694 ;
  assign n9110 = \core_c_dec_IRE_reg[16]/NET0131  & ~n7216 ;
  assign n9111 = \core_c_dec_MFCNTR_E_reg/P0001  & \core_c_psq_CNTR_reg_DO_reg[12]/NET0131  ;
  assign n9112 = \core_c_dec_MFIDR_E_reg/P0001  & \sice_idr1_reg_DO_reg[0]/P0001  ;
  assign n9114 = ~n9111 & ~n9112 ;
  assign n9115 = ~n9110 & n9114 ;
  assign n9116 = ~n9113 & n9115 ;
  assign n9117 = n7215 & ~n9116 ;
  assign n9010 = \bdma_BIAD_reg[12]/NET0131  & n7234 ;
  assign n9028 = \sport0_rxctl_SLOT1_EXT_reg[2]/NET0131  & n7710 ;
  assign n9013 = \sport1_rxctl_SLOT1_EXT_reg[2]/NET0131  & n7689 ;
  assign n9008 = \memc_usysr_DO_reg[12]/NET0131  & n7301 ;
  assign n9009 = \sport0_regs_AUTO_a_reg[12]/NET0131  & n7295 ;
  assign n9031 = ~n9008 & ~n9009 ;
  assign n9043 = ~n9013 & n9031 ;
  assign n9044 = ~n9028 & n9043 ;
  assign n9048 = ~n9010 & n9044 ;
  assign n9011 = \bdma_BCTL_reg[12]/NET0131  & n7230 ;
  assign n9022 = \bdma_BEAD_reg[12]/NET0131  & n7303 ;
  assign n9049 = ~n9011 & ~n9022 ;
  assign n9050 = n9048 & n9049 ;
  assign n9029 = \bdma_BWCOUNT_reg[12]/NET0131  & n7287 ;
  assign n9017 = \PIO_out[8]_pad  & n7291 ;
  assign n9018 = \PIO_oe[8]_pad  & n7244 ;
  assign n9034 = ~n9017 & ~n9018 ;
  assign n9019 = \tm_tpr_reg_DO_reg[12]/NET0131  & n7293 ;
  assign n9020 = \pio_PINT_reg[8]/NET0131  & n7271 ;
  assign n9035 = ~n9019 & ~n9020 ;
  assign n9041 = n9034 & n9035 ;
  assign n9012 = \emc_WSCRreg_DO_reg[12]/NET0131  & n7251 ;
  assign n9014 = \clkc_ckr_reg_DO_reg[12]/NET0131  & n7239 ;
  assign n9032 = ~n9012 & ~n9014 ;
  assign n9015 = \sport0_regs_SCTLreg_DO_reg[12]/NET0131  & n7249 ;
  assign n9016 = \sport1_regs_FSDIVreg_DO_reg[12]/NET0131  & n7273 ;
  assign n9033 = ~n9015 & ~n9016 ;
  assign n9042 = n9032 & n9033 ;
  assign n9045 = n9041 & n9042 ;
  assign n9030 = \sport1_regs_SCTLreg_DO_reg[12]/NET0131  & n7281 ;
  assign n9026 = \sport0_regs_SCLKDIVreg_DO_reg[12]/NET0131  & n7256 ;
  assign n9027 = \sport1_regs_SCLKDIVreg_DO_reg[12]/NET0131  & n7247 ;
  assign n9038 = ~n9026 & ~n9027 ;
  assign n9039 = ~n9030 & n9038 ;
  assign n9021 = \sport0_regs_FSDIVreg_DO_reg[12]/NET0131  & n7259 ;
  assign n9023 = \pio_pmask_reg_DO_reg[8]/NET0131  & n7297 ;
  assign n9036 = ~n9021 & ~n9023 ;
  assign n9024 = \tm_TCR_TMP_reg[12]/NET0131  & n7289 ;
  assign n9025 = \idma_DCTL_reg[12]/NET0131  & n7299 ;
  assign n9037 = ~n9024 & ~n9025 ;
  assign n9040 = n9036 & n9037 ;
  assign n9046 = n9039 & n9040 ;
  assign n9047 = n9045 & n9046 ;
  assign n9051 = ~n9029 & n9047 ;
  assign n9052 = n9050 & n9051 ;
  assign n9053 = \memc_ldSREG_E_reg/NET0131  & ~n9052 ;
  assign n9150 = \core_c_dec_MFLreg_E_reg[5]/P0001  & \core_dag_ilm2reg_L5_we_DO_reg[12]/NET0131  ;
  assign n9151 = \core_c_dec_MFLreg_E_reg[4]/P0001  & \core_dag_ilm2reg_L4_we_DO_reg[12]/NET0131  ;
  assign n9158 = ~n9150 & ~n9151 ;
  assign n9152 = \core_c_dec_MFIreg_E_reg[7]/P0001  & \core_dag_ilm2reg_I7_we_DO_reg[12]/NET0131  ;
  assign n9153 = \core_c_dec_MFIreg_E_reg[6]/P0001  & \core_dag_ilm2reg_I6_we_DO_reg[12]/NET0131  ;
  assign n9159 = ~n9152 & ~n9153 ;
  assign n9160 = n9158 & n9159 ;
  assign n9146 = \core_c_dec_MFMreg_E_reg[5]/P0001  & \core_dag_ilm2reg_M5_we_DO_reg[12]/NET0131  ;
  assign n9147 = \core_c_dec_MFMreg_E_reg[6]/P0001  & \core_dag_ilm2reg_M6_we_DO_reg[12]/NET0131  ;
  assign n9156 = ~n9146 & ~n9147 ;
  assign n9148 = \core_c_dec_MFIreg_E_reg[5]/P0001  & \core_dag_ilm2reg_I5_we_DO_reg[12]/NET0131  ;
  assign n9149 = \core_c_dec_MFLreg_E_reg[6]/P0001  & \core_dag_ilm2reg_L6_we_DO_reg[12]/NET0131  ;
  assign n9157 = ~n9148 & ~n9149 ;
  assign n9161 = n9156 & n9157 ;
  assign n9142 = \core_c_dec_MFIreg_E_reg[4]/P0001  & \core_dag_ilm2reg_I4_we_DO_reg[12]/NET0131  ;
  assign n9143 = \core_c_dec_MFMreg_E_reg[4]/P0001  & \core_dag_ilm2reg_M4_we_DO_reg[12]/NET0131  ;
  assign n9154 = ~n9142 & ~n9143 ;
  assign n9144 = \core_c_dec_MFLreg_E_reg[7]/P0001  & \core_dag_ilm2reg_L7_we_DO_reg[12]/NET0131  ;
  assign n9145 = \core_c_dec_MFMreg_E_reg[7]/P0001  & \core_dag_ilm2reg_M7_we_DO_reg[12]/NET0131  ;
  assign n9155 = ~n9144 & ~n9145 ;
  assign n9162 = n9154 & n9155 ;
  assign n9163 = n9161 & n9162 ;
  assign n9164 = n9160 & n9163 ;
  assign n9165 = n7128 & ~n9164 ;
  assign n8992 = \core_c_dec_MFLreg_E_reg[3]/P0001  & \core_dag_ilm1reg_L3_we_DO_reg[12]/NET0131  ;
  assign n8993 = \core_c_dec_MFIreg_E_reg[3]/P0001  & \core_dag_ilm1reg_I3_we_DO_reg[12]/NET0131  ;
  assign n9000 = ~n8992 & ~n8993 ;
  assign n8994 = \core_c_dec_MFMreg_E_reg[2]/P0001  & \core_dag_ilm1reg_M2_we_DO_reg[12]/NET0131  ;
  assign n8995 = \core_c_dec_MFLreg_E_reg[2]/P0001  & \core_dag_ilm1reg_L2_we_DO_reg[12]/NET0131  ;
  assign n9001 = ~n8994 & ~n8995 ;
  assign n9002 = n9000 & n9001 ;
  assign n8988 = \core_c_dec_MFLreg_E_reg[1]/P0001  & \core_dag_ilm1reg_L1_we_DO_reg[12]/NET0131  ;
  assign n8989 = \core_c_dec_MFIreg_E_reg[0]/P0001  & \core_dag_ilm1reg_I0_we_DO_reg[12]/NET0131  ;
  assign n8998 = ~n8988 & ~n8989 ;
  assign n8990 = \core_c_dec_MFLreg_E_reg[0]/P0001  & \core_dag_ilm1reg_L0_we_DO_reg[12]/NET0131  ;
  assign n8991 = \core_c_dec_MFMreg_E_reg[0]/P0001  & \core_dag_ilm1reg_M0_we_DO_reg[12]/NET0131  ;
  assign n8999 = ~n8990 & ~n8991 ;
  assign n9003 = n8998 & n8999 ;
  assign n8984 = \core_c_dec_MFMreg_E_reg[3]/P0001  & \core_dag_ilm1reg_M3_we_DO_reg[12]/NET0131  ;
  assign n8985 = \core_c_dec_MFIreg_E_reg[1]/P0001  & \core_dag_ilm1reg_I1_we_DO_reg[12]/NET0131  ;
  assign n8996 = ~n8984 & ~n8985 ;
  assign n8986 = \core_c_dec_MFIreg_E_reg[2]/P0001  & \core_dag_ilm1reg_I2_we_DO_reg[12]/NET0131  ;
  assign n8987 = \core_c_dec_MFMreg_E_reg[1]/P0001  & \core_dag_ilm1reg_M1_we_DO_reg[12]/NET0131  ;
  assign n8997 = ~n8986 & ~n8987 ;
  assign n9004 = n8996 & n8997 ;
  assign n9005 = n9003 & n9004 ;
  assign n9006 = n9002 & n9005 ;
  assign n9007 = n7068 & ~n9006 ;
  assign n9134 = \core_c_dec_MFTX1_E_reg/P0001  & \sport1_txctl_TX_reg[12]/P0001  ;
  assign n9135 = \core_c_dec_MFTX0_E_reg/P0001  & \sport0_txctl_TX_reg[12]/P0001  ;
  assign n9138 = ~n9134 & ~n9135 ;
  assign n9136 = \core_c_dec_MFRX1_E_reg/P0001  & \sport1_rxctl_RX_reg[12]/P0001  ;
  assign n9137 = \core_c_dec_MFRX0_E_reg/P0001  & \sport0_rxctl_RX_reg[12]/P0001  ;
  assign n9139 = ~n9136 & ~n9137 ;
  assign n9140 = n9138 & n9139 ;
  assign n9141 = n7119 & ~n9140 ;
  assign n9166 = ~n9007 & ~n9141 ;
  assign n9167 = ~n9165 & n9166 ;
  assign n9126 = ~\core_c_psq_MSTAT_reg_DO_reg[0]/P0002  & \core_eu_es_sht_es_reg_sr1rwe_DO_reg[12]/P0001  ;
  assign n9127 = \core_c_psq_MSTAT_reg_DO_reg[0]/P0002  & \core_eu_es_sht_es_reg_sr1swe_DO_reg[12]/P0001  ;
  assign n9128 = ~n9126 & ~n9127 ;
  assign n9129 = \core_c_dec_MFSR1_E_reg/P0001  & ~n9128 ;
  assign n9118 = ~\core_c_psq_MSTAT_reg_DO_reg[0]/P0002  & \core_eu_es_sht_es_reg_sr0rwe_DO_reg[12]/P0001  ;
  assign n9119 = \core_c_psq_MSTAT_reg_DO_reg[0]/P0002  & \core_eu_es_sht_es_reg_sr0swe_DO_reg[12]/P0001  ;
  assign n9120 = ~n9118 & ~n9119 ;
  assign n9121 = \core_c_dec_MFSR0_E_reg/P0001  & ~n9120 ;
  assign n9122 = ~\core_c_psq_MSTAT_reg_DO_reg[0]/P0002  & \core_eu_es_sht_es_reg_sirwe_DO_reg[12]/P0001  ;
  assign n9123 = \core_c_psq_MSTAT_reg_DO_reg[0]/P0002  & \core_eu_es_sht_es_reg_siswe_DO_reg[12]/P0001  ;
  assign n9124 = ~n9122 & ~n9123 ;
  assign n9125 = \core_c_dec_MFSI_E_reg/P0001  & ~n9124 ;
  assign n9130 = ~n9121 & ~n9125 ;
  assign n9131 = ~n9129 & n9130 ;
  assign n9132 = n7174 & n9131 ;
  assign n9133 = n7153 & ~n9132 ;
  assign n9074 = ~\core_c_psq_MSTAT_reg_DO_reg[0]/P0002  & \core_eu_em_mac_em_reg_mx0rwe_DO_reg[12]/P0001  ;
  assign n9075 = \core_c_psq_MSTAT_reg_DO_reg[0]/P0002  & \core_eu_em_mac_em_reg_mx0swe_DO_reg[12]/P0001  ;
  assign n9076 = ~n9074 & ~n9075 ;
  assign n9077 = \core_c_dec_MFMX0_E_reg/P0001  & ~n9076 ;
  assign n9066 = ~\core_c_psq_MSTAT_reg_DO_reg[0]/P0002  & \core_eu_em_mac_em_reg_my1rwe_DO_reg[12]/P0001  ;
  assign n9067 = \core_c_psq_MSTAT_reg_DO_reg[0]/P0002  & \core_eu_em_mac_em_reg_my1swe_DO_reg[12]/P0001  ;
  assign n9068 = ~n9066 & ~n9067 ;
  assign n9069 = \core_c_dec_MFMY1_E_reg/P0001  & ~n9068 ;
  assign n9070 = ~\core_c_psq_MSTAT_reg_DO_reg[0]/P0002  & \core_eu_em_mac_em_reg_mr0rwe_DO_reg[12]/P0001  ;
  assign n9071 = \core_c_psq_MSTAT_reg_DO_reg[0]/P0002  & \core_eu_em_mac_em_reg_mr0swe_DO_reg[12]/P0001  ;
  assign n9072 = ~n9070 & ~n9071 ;
  assign n9073 = \core_c_dec_MFMR0_E_reg/P0001  & ~n9072 ;
  assign n9080 = ~n9069 & ~n9073 ;
  assign n9081 = ~n9077 & n9080 ;
  assign n9054 = ~\core_c_psq_MSTAT_reg_DO_reg[0]/P0002  & \core_eu_em_mac_em_reg_mr1rwe_DO_reg[12]/P0001  ;
  assign n9055 = \core_c_psq_MSTAT_reg_DO_reg[0]/P0002  & \core_eu_em_mac_em_reg_mr1swe_DO_reg[12]/P0001  ;
  assign n9056 = ~n9054 & ~n9055 ;
  assign n9057 = \core_c_dec_MFMR1_E_reg/P0001  & ~n9056 ;
  assign n9078 = ~n7207 & ~n9057 ;
  assign n9058 = ~\core_c_psq_MSTAT_reg_DO_reg[0]/P0002  & \core_eu_em_mac_em_reg_mx1rwe_DO_reg[12]/P0001  ;
  assign n9059 = \core_c_psq_MSTAT_reg_DO_reg[0]/P0002  & \core_eu_em_mac_em_reg_mx1swe_DO_reg[12]/P0001  ;
  assign n9060 = ~n9058 & ~n9059 ;
  assign n9061 = \core_c_dec_MFMX1_E_reg/P0001  & ~n9060 ;
  assign n9062 = ~\core_c_psq_MSTAT_reg_DO_reg[0]/P0002  & \core_eu_em_mac_em_reg_my0rwe_DO_reg[12]/P0001  ;
  assign n9063 = \core_c_psq_MSTAT_reg_DO_reg[0]/P0002  & \core_eu_em_mac_em_reg_my0swe_DO_reg[12]/P0001  ;
  assign n9064 = ~n9062 & ~n9063 ;
  assign n9065 = \core_c_dec_MFMY0_E_reg/P0001  & ~n9064 ;
  assign n9079 = ~n9061 & ~n9065 ;
  assign n9082 = n9078 & n9079 ;
  assign n9083 = n9081 & n9082 ;
  assign n9084 = n7179 & ~n9083 ;
  assign n9085 = ~\core_c_psq_MSTAT_reg_DO_reg[0]/P0002  & \core_eu_ea_alu_ea_reg_ay1rwe_DO_reg[12]/P0001  ;
  assign n9086 = \core_c_psq_MSTAT_reg_DO_reg[0]/P0002  & \core_eu_ea_alu_ea_reg_ay1swe_DO_reg[12]/P0001  ;
  assign n9087 = ~n9085 & ~n9086 ;
  assign n9088 = \core_c_dec_MFAY1_E_reg/P0001  & ~n9087 ;
  assign n9089 = ~\core_c_psq_MSTAT_reg_DO_reg[0]/P0002  & \core_eu_ea_alu_ea_reg_ax0rwe_DO_reg[12]/P0001  ;
  assign n9090 = \core_c_psq_MSTAT_reg_DO_reg[0]/P0002  & \core_eu_ea_alu_ea_reg_ax0swe_DO_reg[12]/P0001  ;
  assign n9091 = ~n9089 & ~n9090 ;
  assign n9092 = \core_c_dec_MFAX0_E_reg/P0001  & ~n9091 ;
  assign n9105 = ~n9088 & ~n9092 ;
  assign n9101 = ~\core_c_psq_MSTAT_reg_DO_reg[0]/P0002  & \core_eu_ea_alu_ea_reg_arrwe_DO_reg[12]/P0001  ;
  assign n9102 = \core_c_psq_MSTAT_reg_DO_reg[0]/P0002  & \core_eu_ea_alu_ea_reg_arswe_DO_reg[12]/P0001  ;
  assign n9103 = ~n9101 & ~n9102 ;
  assign n9104 = \core_c_dec_MFAR_E_reg/P0001  & ~n9103 ;
  assign n9093 = ~\core_c_psq_MSTAT_reg_DO_reg[0]/P0002  & \core_eu_ea_alu_ea_reg_ay0rwe_DO_reg[12]/P0001  ;
  assign n9094 = \core_c_psq_MSTAT_reg_DO_reg[0]/P0002  & \core_eu_ea_alu_ea_reg_ay0swe_DO_reg[12]/P0001  ;
  assign n9095 = ~n9093 & ~n9094 ;
  assign n9096 = \core_c_dec_MFAY0_E_reg/P0001  & ~n9095 ;
  assign n9097 = ~\core_c_psq_MSTAT_reg_DO_reg[0]/P0002  & \core_eu_ea_alu_ea_reg_ax1rwe_DO_reg[12]/P0001  ;
  assign n9098 = \core_c_psq_MSTAT_reg_DO_reg[0]/P0002  & \core_eu_ea_alu_ea_reg_ax1swe_DO_reg[12]/P0001  ;
  assign n9099 = ~n9097 & ~n9098 ;
  assign n9100 = \core_c_dec_MFAX1_E_reg/P0001  & ~n9099 ;
  assign n9106 = ~n9096 & ~n9100 ;
  assign n9107 = ~n9104 & n9106 ;
  assign n9108 = n9105 & n9107 ;
  assign n9109 = n7093 & ~n9108 ;
  assign n9168 = ~n9084 & ~n9109 ;
  assign n9169 = ~n9133 & n9168 ;
  assign n9170 = n9167 & n9169 ;
  assign n9171 = ~n9053 & n9170 ;
  assign n9172 = ~n9117 & n9171 ;
  assign n9173 = ~n8983 & n9172 ;
  assign n9174 = ~\emc_DMDoe_reg/NET0131  & ~n9173 ;
  assign n9175 = \emc_DMDoe_reg/NET0131  & \emc_DMDreg_reg[12]/P0001  ;
  assign n9176 = n7057 & ~n9175 ;
  assign n9177 = ~n9174 & n9176 ;
  assign n9178 = ~n8982 & ~n9177 ;
  assign n9179 = n6135 & ~n9178 ;
  assign n9180 = n8964 & ~n9179 ;
  assign n9181 = ~n8963 & n9180 ;
  assign n9182 = n8854 & ~n8875 ;
  assign n9183 = n8153 & ~n9182 ;
  assign n9190 = \DM_rd0[1]_pad  & ~n7053 ;
  assign n9184 = \DM_rdm[1]_pad  & n7016 ;
  assign n9195 = ~n7057 & ~n9184 ;
  assign n9187 = \DM_rd6[1]_pad  & n7031 ;
  assign n9188 = \DM_rd7[1]_pad  & n7034 ;
  assign n9196 = ~n9187 & ~n9188 ;
  assign n9197 = n9195 & n9196 ;
  assign n9191 = \DM_rd5[1]_pad  & n7043 ;
  assign n9186 = \DM_rd4[1]_pad  & n7028 ;
  assign n9192 = \DM_rd2[1]_pad  & n7041 ;
  assign n9185 = \DM_rd1[1]_pad  & n7022 ;
  assign n9189 = \DM_rd3[1]_pad  & n7038 ;
  assign n9193 = ~n9185 & ~n9189 ;
  assign n9194 = ~n9192 & n9193 ;
  assign n9198 = ~n9186 & n9194 ;
  assign n9199 = ~n9191 & n9198 ;
  assign n9200 = n9197 & n9199 ;
  assign n9201 = ~n9190 & n9200 ;
  assign n9202 = \regout_STD_C_reg[1]/P0001  & n6988 ;
  assign n9359 = \bdma_BIAD_reg[1]/NET0131  & n7234 ;
  assign n9350 = \emc_WSCRreg_DO_reg[1]/NET0131  & n7251 ;
  assign n9351 = \sport1_regs_SCLKDIVreg_DO_reg[1]/NET0131  & n7247 ;
  assign n9376 = ~n9350 & ~n9351 ;
  assign n9352 = \idma_DOVL_reg[1]/NET0131  & n7532 ;
  assign n9353 = \sport0_regs_AUTOreg_DO_reg[1]/NET0131  & n7295 ;
  assign n9377 = ~n9352 & ~n9353 ;
  assign n9390 = n9376 & n9377 ;
  assign n9346 = \sport0_regs_SCTLreg_DO_reg[1]/NET0131  & n7249 ;
  assign n9374 = ~n7522 & ~n9346 ;
  assign n9347 = \tm_tsr_reg_DO_reg[1]/NET0131  & n7540 ;
  assign n9348 = \sport1_regs_MWORDreg_DO_reg[1]/NET0131  & n7263 ;
  assign n9375 = ~n9347 & ~n9348 ;
  assign n9391 = n9374 & n9375 ;
  assign n9392 = n9390 & n9391 ;
  assign n9396 = ~n9359 & n9392 ;
  assign n9367 = \bdma_BEAD_reg[1]/NET0131  & n7303 ;
  assign n9368 = \bdma_BCTL_reg[1]/NET0131  & n7230 ;
  assign n9397 = ~n9367 & ~n9368 ;
  assign n9398 = n9396 & n9397 ;
  assign n9364 = \bdma_BOVL_reg[1]/NET0131  & n7534 ;
  assign n9349 = \bdma_BWCOUNT_reg[1]/NET0131  & n7287 ;
  assign n9358 = \PIO_oe[1]_pad  & n7244 ;
  assign n9360 = \sport0_regs_MWORDreg_DO_reg[1]/NET0131  & n7276 ;
  assign n9380 = ~n9358 & ~n9360 ;
  assign n9361 = \idma_DCTL_reg[1]/NET0131  & n7299 ;
  assign n9362 = \sport1_regs_FSDIVreg_DO_reg[1]/NET0131  & n7273 ;
  assign n9381 = ~n9361 & ~n9362 ;
  assign n9388 = n9380 & n9381 ;
  assign n9354 = \sport0_regs_SCLKDIVreg_DO_reg[1]/NET0131  & n7256 ;
  assign n9355 = \emc_WSCRext_reg_DO_reg[1]/NET0131  & n7514 ;
  assign n9378 = ~n9354 & ~n9355 ;
  assign n9356 = \sport0_regs_FSDIVreg_DO_reg[1]/NET0131  & n7259 ;
  assign n9357 = \sport1_regs_AUTOreg_DO_reg[1]/NET0131  & n7527 ;
  assign n9379 = ~n9356 & ~n9357 ;
  assign n9389 = n9378 & n9379 ;
  assign n9393 = n9388 & n9389 ;
  assign n9370 = \sport1_regs_SCTLreg_DO_reg[1]/NET0131  & n7281 ;
  assign n9371 = \pio_pmask_reg_DO_reg[1]/NET0131  & n7297 ;
  assign n9384 = ~n9370 & ~n9371 ;
  assign n9372 = \PIO_out[1]_pad  & n7291 ;
  assign n9373 = \tm_TCR_TMP_reg[1]/NET0131  & n7289 ;
  assign n9385 = ~n9372 & ~n9373 ;
  assign n9386 = n9384 & n9385 ;
  assign n9363 = \memc_usysr_DO_reg[1]/NET0131  & n7301 ;
  assign n9365 = \tm_tpr_reg_DO_reg[1]/NET0131  & n7293 ;
  assign n9382 = ~n9363 & ~n9365 ;
  assign n9366 = \clkc_ckr_reg_DO_reg[1]/NET0131  & n7239 ;
  assign n9369 = \pio_PINT_reg[1]/NET0131  & n7271 ;
  assign n9383 = ~n9366 & ~n9369 ;
  assign n9387 = n9382 & n9383 ;
  assign n9394 = n9386 & n9387 ;
  assign n9395 = n9393 & n9394 ;
  assign n9399 = ~n9349 & n9395 ;
  assign n9400 = ~n9364 & n9399 ;
  assign n9401 = n9398 & n9400 ;
  assign n9402 = \memc_ldSREG_E_reg/NET0131  & ~n9401 ;
  assign n9406 = \core_c_dec_MFtoppcs_Eg_reg/P0001  & ~n4457 ;
  assign n9409 = \core_c_dec_MFMSTAT_E_reg/P0001  & \core_c_psq_MSTAT_reg_DO_reg[1]/NET0131  ;
  assign n9410 = \core_c_dec_MFSSTAT_E_reg/P0001  & \core_c_psq_SSTAT_reg[1]/NET0131  ;
  assign n9415 = ~n9409 & ~n9410 ;
  assign n9411 = \core_c_dec_MFCNTR_E_reg/P0001  & \core_c_psq_CNTR_reg_DO_reg[1]/NET0131  ;
  assign n9412 = \core_c_dec_MFICNTL_E_reg/P0001  & \core_c_psq_ICNTL_reg_DO_reg[1]/NET0131  ;
  assign n9416 = ~n9411 & ~n9412 ;
  assign n9417 = n9415 & n9416 ;
  assign n9407 = \core_c_dec_IRE_reg[5]/NET0131  & ~n7216 ;
  assign n9403 = \core_c_dec_MFDMOVL_E_reg/P0001  & \core_c_psq_DMOVL_reg_DO_reg[1]/NET0131  ;
  assign n9404 = \core_c_dec_MFIMASK_E_reg/P0001  & \core_c_psq_IMASK_reg[1]/NET0131  ;
  assign n9413 = ~n9403 & ~n9404 ;
  assign n9405 = \core_c_dec_MFPMOVL_E_reg/P0001  & \core_c_psq_PMOVL_regl_DO_reg[1]/NET0131  ;
  assign n9408 = \core_c_dec_MFIDR_E_reg/P0001  & \sice_idr0_reg_DO_reg[1]/P0001  ;
  assign n9414 = ~n9405 & ~n9408 ;
  assign n9418 = n9413 & n9414 ;
  assign n9419 = ~n9407 & n9418 ;
  assign n9420 = n9417 & n9419 ;
  assign n9421 = ~n9406 & n9420 ;
  assign n9422 = n7215 & ~n9421 ;
  assign n9330 = \core_c_dec_MFLreg_E_reg[6]/P0001  & \core_dag_ilm2reg_L6_we_DO_reg[1]/NET0131  ;
  assign n9331 = \core_c_dec_MFMreg_E_reg[5]/P0001  & \core_dag_ilm2reg_M5_we_DO_reg[1]/NET0131  ;
  assign n9338 = ~n9330 & ~n9331 ;
  assign n9332 = \core_c_dec_MFMreg_E_reg[6]/P0001  & \core_dag_ilm2reg_M6_we_DO_reg[1]/NET0131  ;
  assign n9333 = \core_c_dec_MFMreg_E_reg[7]/P0001  & \core_dag_ilm2reg_M7_we_DO_reg[1]/NET0131  ;
  assign n9339 = ~n9332 & ~n9333 ;
  assign n9340 = n9338 & n9339 ;
  assign n9326 = \core_c_dec_MFLreg_E_reg[7]/P0001  & \core_dag_ilm2reg_L7_we_DO_reg[1]/NET0131  ;
  assign n9327 = \core_c_dec_MFMreg_E_reg[4]/P0001  & \core_dag_ilm2reg_M4_we_DO_reg[1]/NET0131  ;
  assign n9336 = ~n9326 & ~n9327 ;
  assign n9328 = \core_c_dec_MFLreg_E_reg[4]/P0001  & \core_dag_ilm2reg_L4_we_DO_reg[1]/NET0131  ;
  assign n9329 = \core_c_dec_MFLreg_E_reg[5]/P0001  & \core_dag_ilm2reg_L5_we_DO_reg[1]/NET0131  ;
  assign n9337 = ~n9328 & ~n9329 ;
  assign n9341 = n9336 & n9337 ;
  assign n9322 = \core_c_dec_MFIreg_E_reg[7]/P0001  & \core_dag_ilm2reg_I7_we_DO_reg[1]/NET0131  ;
  assign n9323 = \core_c_dec_MFIreg_E_reg[4]/P0001  & \core_dag_ilm2reg_I4_we_DO_reg[1]/NET0131  ;
  assign n9334 = ~n9322 & ~n9323 ;
  assign n9324 = \core_c_dec_MFIreg_E_reg[5]/P0001  & \core_dag_ilm2reg_I5_we_DO_reg[1]/NET0131  ;
  assign n9325 = \core_c_dec_MFIreg_E_reg[6]/P0001  & \core_dag_ilm2reg_I6_we_DO_reg[1]/NET0131  ;
  assign n9335 = ~n9324 & ~n9325 ;
  assign n9342 = n9334 & n9335 ;
  assign n9343 = n9341 & n9342 ;
  assign n9344 = n9340 & n9343 ;
  assign n9345 = n7128 & ~n9344 ;
  assign n9246 = \core_c_dec_MFIreg_E_reg[0]/P0001  & \core_dag_ilm1reg_I0_we_DO_reg[1]/NET0131  ;
  assign n9247 = \core_c_dec_MFIreg_E_reg[3]/P0001  & \core_dag_ilm1reg_I3_we_DO_reg[1]/NET0131  ;
  assign n9254 = ~n9246 & ~n9247 ;
  assign n9248 = \core_c_dec_MFLreg_E_reg[0]/P0001  & \core_dag_ilm1reg_L0_we_DO_reg[1]/NET0131  ;
  assign n9249 = \core_c_dec_MFLreg_E_reg[1]/P0001  & \core_dag_ilm1reg_L1_we_DO_reg[1]/NET0131  ;
  assign n9255 = ~n9248 & ~n9249 ;
  assign n9256 = n9254 & n9255 ;
  assign n9242 = \core_c_dec_MFIreg_E_reg[1]/P0001  & \core_dag_ilm1reg_I1_we_DO_reg[1]/NET0131  ;
  assign n9243 = \core_c_dec_MFIreg_E_reg[2]/P0001  & \core_dag_ilm1reg_I2_we_DO_reg[1]/NET0131  ;
  assign n9252 = ~n9242 & ~n9243 ;
  assign n9244 = \core_c_dec_MFLreg_E_reg[3]/P0001  & \core_dag_ilm1reg_L3_we_DO_reg[1]/NET0131  ;
  assign n9245 = \core_c_dec_MFMreg_E_reg[0]/P0001  & \core_dag_ilm1reg_M0_we_DO_reg[1]/NET0131  ;
  assign n9253 = ~n9244 & ~n9245 ;
  assign n9257 = n9252 & n9253 ;
  assign n9238 = \core_c_dec_MFLreg_E_reg[2]/P0001  & \core_dag_ilm1reg_L2_we_DO_reg[1]/NET0131  ;
  assign n9239 = \core_c_dec_MFMreg_E_reg[1]/P0001  & \core_dag_ilm1reg_M1_we_DO_reg[1]/NET0131  ;
  assign n9250 = ~n9238 & ~n9239 ;
  assign n9240 = \core_c_dec_MFMreg_E_reg[2]/P0001  & \core_dag_ilm1reg_M2_we_DO_reg[1]/NET0131  ;
  assign n9241 = \core_c_dec_MFMreg_E_reg[3]/P0001  & \core_dag_ilm1reg_M3_we_DO_reg[1]/NET0131  ;
  assign n9251 = ~n9240 & ~n9241 ;
  assign n9258 = n9250 & n9251 ;
  assign n9259 = n9257 & n9258 ;
  assign n9260 = n9256 & n9259 ;
  assign n9261 = n7068 & ~n9260 ;
  assign n9287 = \core_c_dec_MFTX1_E_reg/P0001  & \sport1_txctl_TX_reg[1]/P0001  ;
  assign n9288 = \core_c_dec_MFTX0_E_reg/P0001  & \sport0_txctl_TX_reg[1]/P0001  ;
  assign n9291 = ~n9287 & ~n9288 ;
  assign n9289 = \core_c_dec_MFRX1_E_reg/P0001  & \sport1_rxctl_RX_reg[1]/P0001  ;
  assign n9290 = \core_c_dec_MFRX0_E_reg/P0001  & \sport0_rxctl_RX_reg[1]/P0001  ;
  assign n9292 = ~n9289 & ~n9290 ;
  assign n9293 = n9291 & n9292 ;
  assign n9294 = n7119 & ~n9293 ;
  assign n9423 = ~n9261 & ~n9294 ;
  assign n9424 = ~n9345 & n9423 ;
  assign n9295 = ~\core_c_psq_MSTAT_reg_DO_reg[0]/P0002  & \core_eu_ea_alu_ea_reg_arrwe_DO_reg[1]/P0001  ;
  assign n9296 = \core_c_psq_MSTAT_reg_DO_reg[0]/P0002  & \core_eu_ea_alu_ea_reg_arswe_DO_reg[1]/P0001  ;
  assign n9297 = ~n9295 & ~n9296 ;
  assign n9298 = \core_c_dec_MFAR_E_reg/P0001  & ~n9297 ;
  assign n9315 = \core_c_dec_MFASTAT_E_reg/P0001  & \core_eu_ec_cun_AN_reg/P0001  ;
  assign n9316 = ~n9298 & ~n9315 ;
  assign n9299 = ~\core_c_psq_MSTAT_reg_DO_reg[0]/P0002  & \core_eu_ea_alu_ea_reg_ay1rwe_DO_reg[1]/P0001  ;
  assign n9300 = \core_c_psq_MSTAT_reg_DO_reg[0]/P0002  & \core_eu_ea_alu_ea_reg_ay1swe_DO_reg[1]/P0001  ;
  assign n9301 = ~n9299 & ~n9300 ;
  assign n9302 = \core_c_dec_MFAY1_E_reg/P0001  & ~n9301 ;
  assign n9303 = ~\core_c_psq_MSTAT_reg_DO_reg[0]/P0002  & \core_eu_ea_alu_ea_reg_ay0rwe_DO_reg[1]/P0001  ;
  assign n9304 = \core_c_psq_MSTAT_reg_DO_reg[0]/P0002  & \core_eu_ea_alu_ea_reg_ay0swe_DO_reg[1]/P0001  ;
  assign n9305 = ~n9303 & ~n9304 ;
  assign n9306 = \core_c_dec_MFAY0_E_reg/P0001  & ~n9305 ;
  assign n9317 = ~n9302 & ~n9306 ;
  assign n9307 = ~\core_c_psq_MSTAT_reg_DO_reg[0]/P0002  & \core_eu_ea_alu_ea_reg_ax0rwe_DO_reg[1]/P0001  ;
  assign n9308 = \core_c_psq_MSTAT_reg_DO_reg[0]/P0002  & \core_eu_ea_alu_ea_reg_ax0swe_DO_reg[1]/P0001  ;
  assign n9309 = ~n9307 & ~n9308 ;
  assign n9310 = \core_c_dec_MFAX0_E_reg/P0001  & ~n9309 ;
  assign n9311 = ~\core_c_psq_MSTAT_reg_DO_reg[0]/P0002  & \core_eu_ea_alu_ea_reg_ax1rwe_DO_reg[1]/P0001  ;
  assign n9312 = \core_c_psq_MSTAT_reg_DO_reg[0]/P0002  & \core_eu_ea_alu_ea_reg_ax1swe_DO_reg[1]/P0001  ;
  assign n9313 = ~n9311 & ~n9312 ;
  assign n9314 = \core_c_dec_MFAX1_E_reg/P0001  & ~n9313 ;
  assign n9318 = ~n9310 & ~n9314 ;
  assign n9319 = n9317 & n9318 ;
  assign n9320 = n9316 & n9319 ;
  assign n9321 = n7093 & ~n9320 ;
  assign n9227 = ~\core_c_psq_MSTAT_reg_DO_reg[0]/P0002  & \core_eu_em_mac_em_reg_mr2rwe_DO_reg[1]/P0001  ;
  assign n9228 = \core_c_psq_MSTAT_reg_DO_reg[0]/P0002  & \core_eu_em_mac_em_reg_mr2swe_DO_reg[1]/P0001  ;
  assign n9229 = ~n9227 & ~n9228 ;
  assign n9230 = \core_c_dec_MFMR2_E_reg/P0001  & ~n9229 ;
  assign n9219 = ~\core_c_psq_MSTAT_reg_DO_reg[0]/P0002  & \core_eu_em_mac_em_reg_mx0rwe_DO_reg[1]/P0001  ;
  assign n9220 = \core_c_psq_MSTAT_reg_DO_reg[0]/P0002  & \core_eu_em_mac_em_reg_mx0swe_DO_reg[1]/P0001  ;
  assign n9221 = ~n9219 & ~n9220 ;
  assign n9222 = \core_c_dec_MFMX0_E_reg/P0001  & ~n9221 ;
  assign n9223 = ~\core_c_psq_MSTAT_reg_DO_reg[0]/P0002  & \core_eu_em_mac_em_reg_mr0rwe_DO_reg[1]/P0001  ;
  assign n9224 = \core_c_psq_MSTAT_reg_DO_reg[0]/P0002  & \core_eu_em_mac_em_reg_mr0swe_DO_reg[1]/P0001  ;
  assign n9225 = ~n9223 & ~n9224 ;
  assign n9226 = \core_c_dec_MFMR0_E_reg/P0001  & ~n9225 ;
  assign n9233 = ~n9222 & ~n9226 ;
  assign n9234 = ~n9230 & n9233 ;
  assign n9203 = ~\core_c_psq_MSTAT_reg_DO_reg[0]/P0002  & \core_eu_em_mac_em_reg_mr1rwe_DO_reg[1]/P0001  ;
  assign n9204 = \core_c_psq_MSTAT_reg_DO_reg[0]/P0002  & \core_eu_em_mac_em_reg_mr1swe_DO_reg[1]/P0001  ;
  assign n9205 = ~n9203 & ~n9204 ;
  assign n9206 = \core_c_dec_MFMR1_E_reg/P0001  & ~n9205 ;
  assign n9207 = ~\core_c_psq_MSTAT_reg_DO_reg[0]/P0002  & \core_eu_em_mac_em_reg_my0rwe_DO_reg[1]/P0001  ;
  assign n9208 = \core_c_psq_MSTAT_reg_DO_reg[0]/P0002  & \core_eu_em_mac_em_reg_my0swe_DO_reg[1]/P0001  ;
  assign n9209 = ~n9207 & ~n9208 ;
  assign n9210 = \core_c_dec_MFMY0_E_reg/P0001  & ~n9209 ;
  assign n9231 = ~n9206 & ~n9210 ;
  assign n9211 = ~\core_c_psq_MSTAT_reg_DO_reg[0]/P0002  & \core_eu_em_mac_em_reg_mx1rwe_DO_reg[1]/P0001  ;
  assign n9212 = \core_c_psq_MSTAT_reg_DO_reg[0]/P0002  & \core_eu_em_mac_em_reg_mx1swe_DO_reg[1]/P0001  ;
  assign n9213 = ~n9211 & ~n9212 ;
  assign n9214 = \core_c_dec_MFMX1_E_reg/P0001  & ~n9213 ;
  assign n9215 = ~\core_c_psq_MSTAT_reg_DO_reg[0]/P0002  & \core_eu_em_mac_em_reg_my1rwe_DO_reg[1]/P0001  ;
  assign n9216 = \core_c_psq_MSTAT_reg_DO_reg[0]/P0002  & \core_eu_em_mac_em_reg_my1swe_DO_reg[1]/P0001  ;
  assign n9217 = ~n9215 & ~n9216 ;
  assign n9218 = \core_c_dec_MFMY1_E_reg/P0001  & ~n9217 ;
  assign n9232 = ~n9214 & ~n9218 ;
  assign n9235 = n9231 & n9232 ;
  assign n9236 = n9234 & n9235 ;
  assign n9237 = n7179 & ~n9236 ;
  assign n9262 = ~\core_c_psq_MSTAT_reg_DO_reg[0]/P0002  & \core_eu_es_sht_es_reg_sirwe_DO_reg[1]/P0001  ;
  assign n9263 = \core_c_psq_MSTAT_reg_DO_reg[0]/P0002  & \core_eu_es_sht_es_reg_siswe_DO_reg[1]/P0001  ;
  assign n9264 = ~n9262 & ~n9263 ;
  assign n9265 = \core_c_dec_MFSI_E_reg/P0001  & ~n9264 ;
  assign n9266 = ~\core_c_psq_MSTAT_reg_DO_reg[0]/P0002  & \core_eu_es_sht_es_reg_SBr_reg[1]/P0001  ;
  assign n9267 = \core_c_psq_MSTAT_reg_DO_reg[0]/P0002  & \core_eu_es_sht_es_reg_SBs_reg[1]/P0001  ;
  assign n9268 = ~n9266 & ~n9267 ;
  assign n9269 = \core_c_dec_MFSB_E_reg/P0001  & ~n9268 ;
  assign n9282 = ~n9265 & ~n9269 ;
  assign n9278 = ~\core_c_psq_MSTAT_reg_DO_reg[0]/P0002  & \core_eu_es_sht_es_reg_sr1rwe_DO_reg[1]/P0001  ;
  assign n9279 = \core_c_psq_MSTAT_reg_DO_reg[0]/P0002  & \core_eu_es_sht_es_reg_sr1swe_DO_reg[1]/P0001  ;
  assign n9280 = ~n9278 & ~n9279 ;
  assign n9281 = \core_c_dec_MFSR1_E_reg/P0001  & ~n9280 ;
  assign n9270 = ~\core_c_psq_MSTAT_reg_DO_reg[0]/P0002  & \core_eu_es_sht_es_reg_serwe_DO_reg[1]/P0001  ;
  assign n9271 = \core_c_psq_MSTAT_reg_DO_reg[0]/P0002  & \core_eu_es_sht_es_reg_seswe_DO_reg[1]/P0001  ;
  assign n9272 = ~n9270 & ~n9271 ;
  assign n9273 = \core_c_dec_MFSE_E_reg/P0001  & ~n9272 ;
  assign n9274 = ~\core_c_psq_MSTAT_reg_DO_reg[0]/P0002  & \core_eu_es_sht_es_reg_sr0rwe_DO_reg[1]/P0001  ;
  assign n9275 = \core_c_psq_MSTAT_reg_DO_reg[0]/P0002  & \core_eu_es_sht_es_reg_sr0swe_DO_reg[1]/P0001  ;
  assign n9276 = ~n9274 & ~n9275 ;
  assign n9277 = \core_c_dec_MFSR0_E_reg/P0001  & ~n9276 ;
  assign n9283 = ~n9273 & ~n9277 ;
  assign n9284 = ~n9281 & n9283 ;
  assign n9285 = n9282 & n9284 ;
  assign n9286 = n7153 & ~n9285 ;
  assign n9425 = ~n9237 & ~n9286 ;
  assign n9426 = ~n9321 & n9425 ;
  assign n9427 = n9424 & n9426 ;
  assign n9428 = ~n9422 & n9427 ;
  assign n9429 = ~n9402 & n9428 ;
  assign n9430 = ~n9202 & n9429 ;
  assign n9431 = ~\emc_DMDoe_reg/NET0131  & ~n9430 ;
  assign n9432 = \emc_DMDoe_reg/NET0131  & \emc_DMDreg_reg[1]/P0001  ;
  assign n9433 = n7057 & ~n9432 ;
  assign n9434 = ~n9431 & n9433 ;
  assign n9435 = ~n9201 & ~n9434 ;
  assign n9436 = n7863 & n9435 ;
  assign n9437 = ~n9183 & ~n9436 ;
  assign n9438 = n7005 & ~n9437 ;
  assign n9439 = ~n9181 & ~n9438 ;
  assign n9440 = ~n8950 & n9439 ;
  assign n9477 = ~n6888 & ~n6898 ;
  assign n9478 = ~n6880 & ~n6895 ;
  assign n9479 = ~n6899 & ~n9478 ;
  assign n9480 = n9477 & ~n9479 ;
  assign n9481 = ~n9477 & n9479 ;
  assign n9482 = ~n9480 & ~n9481 ;
  assign n9483 = n6717 & ~n9482 ;
  assign n9484 = ~\core_dag_ilm2reg_M_reg[13]/NET0131  & ~n6605 ;
  assign n9485 = ~n6606 & ~n9484 ;
  assign n9486 = ~n6712 & n9485 ;
  assign n9487 = n6712 & ~n9485 ;
  assign n9488 = ~n9486 & ~n9487 ;
  assign n9489 = \core_dag_ilm2reg_M_reg[13]/NET0131  & n9488 ;
  assign n9490 = ~n9483 & n9489 ;
  assign n9491 = ~n6905 & ~n9488 ;
  assign n9492 = n6905 & ~n9482 ;
  assign n9493 = ~\core_dag_ilm2reg_M_reg[13]/NET0131  & ~n9492 ;
  assign n9494 = ~n9491 & n9493 ;
  assign n9495 = \core_dag_ilm2reg_I_reg[13]/NET0131  & n6604 ;
  assign n9496 = ~n9494 & ~n9495 ;
  assign n9497 = ~n9490 & n9496 ;
  assign n9498 = ~n6176 & ~n9497 ;
  assign n9476 = n6176 & ~n7622 ;
  assign n9499 = n6135 & ~n9476 ;
  assign n9500 = ~n9498 & n9499 ;
  assign n9446 = \core_dag_ilm2reg_I4_we_DO_reg[13]/NET0131  & n6976 ;
  assign n9447 = \core_dag_ilm2reg_I5_we_DO_reg[13]/NET0131  & n6970 ;
  assign n9450 = ~n9446 & ~n9447 ;
  assign n9448 = \core_dag_ilm2reg_I6_we_DO_reg[13]/NET0131  & n6974 ;
  assign n9449 = \core_dag_ilm2reg_I7_we_DO_reg[13]/NET0131  & n6972 ;
  assign n9451 = ~n9448 & ~n9449 ;
  assign n9452 = n9450 & n9451 ;
  assign n9453 = n4055 & ~n9452 ;
  assign n9454 = \core_dag_ilm2reg_I7_we_DO_reg[13]/NET0131  & n6960 ;
  assign n9455 = \core_dag_ilm2reg_I4_we_DO_reg[13]/NET0131  & n6958 ;
  assign n9458 = ~n9454 & ~n9455 ;
  assign n9456 = \core_dag_ilm2reg_I6_we_DO_reg[13]/NET0131  & n6962 ;
  assign n9457 = \core_dag_ilm2reg_I5_we_DO_reg[13]/NET0131  & n6964 ;
  assign n9459 = ~n9456 & ~n9457 ;
  assign n9460 = n9458 & n9459 ;
  assign n9461 = ~n9453 & n9460 ;
  assign n9462 = ~n6121 & ~n9461 ;
  assign n9444 = ~n6111 & n6160 ;
  assign n9445 = \core_c_dec_IR_reg[17]/NET0131  & n6956 ;
  assign n9463 = ~n9444 & ~n9445 ;
  assign n9464 = ~n9462 & n9463 ;
  assign n9465 = n5949 & ~n9464 ;
  assign n9466 = \core_dag_ilm1reg_DMA_pi_DO_reg[13]/NET0131  & ~n6934 ;
  assign n9442 = \core_dag_ilm1reg_STAC_pi_DO_reg[13]/NET0131  & n6988 ;
  assign n9443 = \idma_DCTL_reg[13]/NET0131  & n6926 ;
  assign n9467 = ~n9442 & ~n9443 ;
  assign n9468 = n6924 & n9467 ;
  assign n9469 = ~n9466 & n9468 ;
  assign n9470 = ~n9465 & n9469 ;
  assign n9441 = ~\bdma_BIAD_reg[13]/NET0131  & ~n6924 ;
  assign n9471 = ~n6176 & ~n9441 ;
  assign n9472 = ~n9470 & n9471 ;
  assign n9473 = n6176 & n6953 ;
  assign n9474 = ~n6135 & ~n9473 ;
  assign n9475 = ~n9472 & n9474 ;
  assign n9501 = ~n7005 & ~n9475 ;
  assign n9502 = ~n9500 & n9501 ;
  assign n9503 = ~n6160 & n9461 ;
  assign n9504 = n8153 & ~n9503 ;
  assign n9505 = n7607 & n7863 ;
  assign n9506 = ~n9504 & ~n9505 ;
  assign n9507 = n7005 & ~n9506 ;
  assign n9508 = ~n6135 & n6546 ;
  assign n9509 = n6135 & ~n7340 ;
  assign n9510 = n8964 & ~n9509 ;
  assign n9511 = ~n9508 & n9510 ;
  assign n9512 = ~n9507 & ~n9511 ;
  assign n9513 = ~n9502 & n9512 ;
  assign n9533 = ~n6135 & ~n9178 ;
  assign n9514 = \core_dag_ilm2reg_I5_we_DO_reg[1]/NET0131  & n6964 ;
  assign n9515 = \core_dag_ilm2reg_I7_we_DO_reg[1]/NET0131  & n6960 ;
  assign n9518 = ~n9514 & ~n9515 ;
  assign n9516 = \core_dag_ilm2reg_I6_we_DO_reg[1]/NET0131  & n6962 ;
  assign n9517 = \core_dag_ilm2reg_I4_we_DO_reg[1]/NET0131  & n6958 ;
  assign n9519 = ~n9516 & ~n9517 ;
  assign n9520 = n9518 & n9519 ;
  assign n9521 = ~n4055 & n9520 ;
  assign n9522 = \core_dag_ilm2reg_I4_we_DO_reg[1]/NET0131  & n6976 ;
  assign n9523 = \core_dag_ilm2reg_I5_we_DO_reg[1]/NET0131  & n6970 ;
  assign n9526 = ~n9522 & ~n9523 ;
  assign n9524 = \core_dag_ilm2reg_I6_we_DO_reg[1]/NET0131  & n6974 ;
  assign n9525 = \core_dag_ilm2reg_I7_we_DO_reg[1]/NET0131  & n6972 ;
  assign n9527 = ~n9524 & ~n9525 ;
  assign n9528 = n9526 & n9527 ;
  assign n9529 = n4055 & n9528 ;
  assign n9530 = ~n9521 & ~n9529 ;
  assign n9531 = ~n8905 & ~n9530 ;
  assign n9532 = n6135 & n9531 ;
  assign n9534 = ~n6176 & ~n9532 ;
  assign n9535 = ~n9533 & n9534 ;
  assign n9536 = ~n6135 & n8926 ;
  assign n9537 = n6135 & ~n9435 ;
  assign n9538 = n6176 & ~n9537 ;
  assign n9539 = ~n9536 & n9538 ;
  assign n9540 = ~n9535 & ~n9539 ;
  assign n9541 = n7005 & ~n9540 ;
  assign n9545 = n6596 & ~n6807 ;
  assign n9546 = ~n6596 & n6807 ;
  assign n9547 = ~n9545 & ~n9546 ;
  assign n9548 = ~n6717 & n9547 ;
  assign n9543 = ~n6811 & ~n6812 ;
  assign n9544 = n6713 & ~n9543 ;
  assign n9549 = \core_dag_ilm2reg_M_reg[13]/NET0131  & ~n9544 ;
  assign n9550 = ~n9548 & n9549 ;
  assign n9542 = \core_dag_ilm2reg_I_reg[1]/NET0131  & n6664 ;
  assign n9555 = ~n6905 & n9547 ;
  assign n9551 = n6724 & ~n9543 ;
  assign n9552 = ~n6724 & n9543 ;
  assign n9553 = ~n9551 & ~n9552 ;
  assign n9554 = n6905 & n9553 ;
  assign n9556 = ~\core_dag_ilm2reg_M_reg[13]/NET0131  & ~n9554 ;
  assign n9557 = ~n9555 & n9556 ;
  assign n9558 = ~n9542 & ~n9557 ;
  assign n9559 = ~n9550 & n9558 ;
  assign n9560 = n6135 & ~n9559 ;
  assign n9566 = ~n6121 & n9530 ;
  assign n9565 = ~n6111 & n8905 ;
  assign n9567 = \core_c_dec_IR_reg[5]/NET0131  & n6956 ;
  assign n9568 = ~n9565 & ~n9567 ;
  assign n9569 = ~n9566 & n9568 ;
  assign n9570 = n5949 & ~n9569 ;
  assign n9562 = \core_dag_ilm1reg_DMA_pi_DO_reg[1]/NET0131  & ~n6934 ;
  assign n9563 = \idma_DCTL_reg[1]/NET0131  & n6926 ;
  assign n9564 = \core_dag_ilm1reg_STAC_pi_DO_reg[1]/NET0131  & n6988 ;
  assign n9571 = ~n9563 & ~n9564 ;
  assign n9572 = n6924 & n9571 ;
  assign n9573 = ~n9562 & n9572 ;
  assign n9574 = ~n9570 & n9573 ;
  assign n9561 = ~\bdma_BIAD_reg[1]/NET0131  & ~n6924 ;
  assign n9575 = ~n6135 & ~n9561 ;
  assign n9576 = ~n9574 & n9575 ;
  assign n9577 = ~n9560 & ~n9576 ;
  assign n9578 = ~n6176 & ~n9577 ;
  assign n9580 = n6135 & n8962 ;
  assign n9579 = ~n6135 & ~n8875 ;
  assign n9581 = n6176 & ~n9579 ;
  assign n9582 = ~n9580 & n9581 ;
  assign n9583 = ~n9578 & ~n9582 ;
  assign n9584 = ~n7005 & ~n9583 ;
  assign n9585 = ~n9541 & ~n9584 ;
  assign n9605 = ~n6135 & ~n8460 ;
  assign n9586 = \core_dag_ilm2reg_I7_we_DO_reg[2]/NET0131  & n6960 ;
  assign n9587 = \core_dag_ilm2reg_I4_we_DO_reg[2]/NET0131  & n6958 ;
  assign n9590 = ~n9586 & ~n9587 ;
  assign n9588 = \core_dag_ilm2reg_I6_we_DO_reg[2]/NET0131  & n6962 ;
  assign n9589 = \core_dag_ilm2reg_I5_we_DO_reg[2]/NET0131  & n6964 ;
  assign n9591 = ~n9588 & ~n9589 ;
  assign n9592 = n9590 & n9591 ;
  assign n9593 = ~n4055 & n9592 ;
  assign n9594 = \core_dag_ilm2reg_I7_we_DO_reg[2]/NET0131  & n6972 ;
  assign n9595 = \core_dag_ilm2reg_I4_we_DO_reg[2]/NET0131  & n6976 ;
  assign n9598 = ~n9594 & ~n9595 ;
  assign n9596 = \core_dag_ilm2reg_I6_we_DO_reg[2]/NET0131  & n6974 ;
  assign n9597 = \core_dag_ilm2reg_I5_we_DO_reg[2]/NET0131  & n6970 ;
  assign n9599 = ~n9596 & ~n9597 ;
  assign n9600 = n9598 & n9599 ;
  assign n9601 = n4055 & n9600 ;
  assign n9602 = ~n9593 & ~n9601 ;
  assign n9603 = ~n8775 & ~n9602 ;
  assign n9604 = n6135 & n9603 ;
  assign n9606 = ~n6176 & ~n9604 ;
  assign n9607 = ~n9605 & n9606 ;
  assign n9608 = ~n6135 & n8794 ;
  assign n9609 = n6135 & ~n8715 ;
  assign n9610 = n6176 & ~n9609 ;
  assign n9611 = ~n9608 & n9610 ;
  assign n9612 = ~n9607 & ~n9611 ;
  assign n9613 = n7005 & ~n9612 ;
  assign n9620 = ~n6671 & ~n6799 ;
  assign n9621 = n6671 & n6799 ;
  assign n9622 = ~n9620 & ~n9621 ;
  assign n9623 = ~n8198 & n9622 ;
  assign n9614 = \core_dag_ilm2reg_I_reg[2]/NET0131  & ~n6660 ;
  assign n9615 = ~n6803 & ~n6804 ;
  assign n9616 = ~n6815 & ~n9615 ;
  assign n9617 = n6815 & n9615 ;
  assign n9618 = ~n9616 & ~n9617 ;
  assign n9619 = n8198 & n9618 ;
  assign n9624 = ~n9614 & ~n9619 ;
  assign n9625 = ~n9623 & n9624 ;
  assign n9626 = n6135 & ~n9625 ;
  assign n9632 = ~n6121 & n9602 ;
  assign n9631 = ~n6111 & n8775 ;
  assign n9633 = \core_c_dec_IR_reg[6]/NET0131  & n6956 ;
  assign n9634 = ~n9631 & ~n9633 ;
  assign n9635 = ~n9632 & n9634 ;
  assign n9636 = n5949 & ~n9635 ;
  assign n9628 = \core_dag_ilm1reg_DMA_pi_DO_reg[2]/NET0131  & ~n6934 ;
  assign n9629 = \idma_DCTL_reg[2]/NET0131  & n6926 ;
  assign n9630 = \core_dag_ilm1reg_STAC_pi_DO_reg[2]/NET0131  & n6988 ;
  assign n9637 = ~n9629 & ~n9630 ;
  assign n9638 = n6924 & n9637 ;
  assign n9639 = ~n9628 & n9638 ;
  assign n9640 = ~n9636 & n9639 ;
  assign n9627 = ~\bdma_BIAD_reg[2]/NET0131  & ~n6924 ;
  assign n9641 = ~n6135 & ~n9627 ;
  assign n9642 = ~n9640 & n9641 ;
  assign n9643 = ~n9626 & ~n9642 ;
  assign n9644 = ~n6176 & ~n9643 ;
  assign n9645 = n6135 & n8246 ;
  assign n9646 = ~n6135 & ~n8752 ;
  assign n9647 = n6176 & ~n9646 ;
  assign n9648 = ~n9645 & n9647 ;
  assign n9649 = ~n9644 & ~n9648 ;
  assign n9650 = ~n7005 & ~n9649 ;
  assign n9651 = ~n9613 & ~n9650 ;
  assign n9671 = ~n6135 & n7859 ;
  assign n9652 = \core_dag_ilm2reg_I4_we_DO_reg[3]/NET0131  & n6958 ;
  assign n9653 = \core_dag_ilm2reg_I7_we_DO_reg[3]/NET0131  & n6960 ;
  assign n9656 = ~n9652 & ~n9653 ;
  assign n9654 = \core_dag_ilm2reg_I6_we_DO_reg[3]/NET0131  & n6962 ;
  assign n9655 = \core_dag_ilm2reg_I5_we_DO_reg[3]/NET0131  & n6964 ;
  assign n9657 = ~n9654 & ~n9655 ;
  assign n9658 = n9656 & n9657 ;
  assign n9659 = ~n4055 & n9658 ;
  assign n9660 = \core_dag_ilm2reg_I4_we_DO_reg[3]/NET0131  & n6976 ;
  assign n9661 = \core_dag_ilm2reg_I5_we_DO_reg[3]/NET0131  & n6970 ;
  assign n9664 = ~n9660 & ~n9661 ;
  assign n9662 = \core_dag_ilm2reg_I6_we_DO_reg[3]/NET0131  & n6974 ;
  assign n9663 = \core_dag_ilm2reg_I7_we_DO_reg[3]/NET0131  & n6972 ;
  assign n9665 = ~n9662 & ~n9663 ;
  assign n9666 = n9664 & n9665 ;
  assign n9667 = n4055 & n9666 ;
  assign n9668 = ~n9659 & ~n9667 ;
  assign n9669 = ~n8192 & ~n9668 ;
  assign n9670 = n6135 & ~n9669 ;
  assign n9672 = ~n6176 & ~n9670 ;
  assign n9673 = ~n9671 & n9672 ;
  assign n9675 = ~n6135 & ~n8224 ;
  assign n9674 = n6135 & n8113 ;
  assign n9676 = n6176 & ~n9674 ;
  assign n9677 = ~n9675 & n9676 ;
  assign n9678 = ~n9673 & ~n9677 ;
  assign n9679 = n7005 & ~n9678 ;
  assign n9681 = n6135 & ~n7644 ;
  assign n9680 = ~n6135 & n8151 ;
  assign n9682 = n6176 & ~n9680 ;
  assign n9683 = ~n9681 & n9682 ;
  assign n9690 = ~n6673 & ~n6788 ;
  assign n9691 = n6673 & n6788 ;
  assign n9692 = ~n9690 & ~n9691 ;
  assign n9693 = ~n8198 & n9692 ;
  assign n9684 = \core_dag_ilm2reg_I_reg[3]/NET0131  & ~n6653 ;
  assign n9685 = ~n6792 & ~n6793 ;
  assign n9686 = ~n6817 & ~n9685 ;
  assign n9687 = n6817 & n9685 ;
  assign n9688 = ~n9686 & ~n9687 ;
  assign n9689 = n8198 & n9688 ;
  assign n9694 = ~n9684 & ~n9689 ;
  assign n9695 = ~n9693 & n9694 ;
  assign n9696 = n6135 & ~n9695 ;
  assign n9701 = ~n6121 & n9668 ;
  assign n9699 = ~n6111 & n8192 ;
  assign n9700 = \core_c_dec_IR_reg[7]/NET0131  & n6956 ;
  assign n9702 = ~n9699 & ~n9700 ;
  assign n9703 = ~n9701 & n9702 ;
  assign n9704 = n5949 & ~n9703 ;
  assign n9698 = \core_dag_ilm1reg_DMA_pi_DO_reg[3]/NET0131  & ~n6934 ;
  assign n9697 = \idma_DCTL_reg[3]/NET0131  & n6926 ;
  assign n9705 = \core_dag_ilm1reg_STAC_pi_DO_reg[3]/NET0131  & n6988 ;
  assign n9706 = ~n9697 & ~n9705 ;
  assign n9707 = ~n9698 & n9706 ;
  assign n9708 = ~n9704 & n9707 ;
  assign n9709 = n6924 & ~n9708 ;
  assign n9710 = \bdma_BIAD_reg[3]/NET0131  & ~n6924 ;
  assign n9711 = ~n9709 & ~n9710 ;
  assign n9712 = ~n6135 & ~n9711 ;
  assign n9713 = ~n6176 & ~n9712 ;
  assign n9714 = ~n9696 & n9713 ;
  assign n9715 = ~n9683 & ~n9714 ;
  assign n9716 = ~n7005 & ~n9715 ;
  assign n9717 = ~n9679 & ~n9716 ;
  assign n9737 = \core_dag_ilm1reg_I_reg[9]/NET0131  & n6389 ;
  assign n9738 = ~n6410 & ~n6458 ;
  assign n9739 = ~n6385 & ~n6417 ;
  assign n9740 = ~n6459 & ~n9739 ;
  assign n9741 = n9738 & ~n9740 ;
  assign n9742 = ~n9738 & n9740 ;
  assign n9743 = ~n9741 & ~n9742 ;
  assign n9744 = ~n7631 & ~n9743 ;
  assign n9745 = ~n6403 & ~n6514 ;
  assign n9746 = ~n6404 & ~n9745 ;
  assign n9747 = n6393 & ~n9746 ;
  assign n9748 = ~n6393 & n9746 ;
  assign n9749 = ~n9747 & ~n9748 ;
  assign n9750 = n7631 & n9749 ;
  assign n9751 = ~n9744 & ~n9750 ;
  assign n9752 = ~n9737 & ~n9751 ;
  assign n9753 = n6135 & ~n9752 ;
  assign n9718 = \core_dag_ilm1reg_I0_we_DO_reg[9]/NET0131  & n6058 ;
  assign n9719 = n6060 & n9718 ;
  assign n9723 = ~n4055 & ~n9719 ;
  assign n9722 = \core_dag_ilm1reg_I3_we_DO_reg[9]/NET0131  & n6140 ;
  assign n9720 = \core_dag_ilm1reg_I2_we_DO_reg[9]/NET0131  & n6138 ;
  assign n9721 = \core_dag_ilm1reg_I1_we_DO_reg[9]/NET0131  & n6142 ;
  assign n9724 = ~n9720 & ~n9721 ;
  assign n9725 = ~n9722 & n9724 ;
  assign n9726 = n9723 & n9725 ;
  assign n9727 = n6093 & n9718 ;
  assign n9728 = \core_dag_ilm1reg_I2_we_DO_reg[9]/NET0131  & n6152 ;
  assign n9731 = ~n9727 & ~n9728 ;
  assign n9729 = \core_dag_ilm1reg_I3_we_DO_reg[9]/NET0131  & n6150 ;
  assign n9730 = \core_dag_ilm1reg_I1_we_DO_reg[9]/NET0131  & n6154 ;
  assign n9732 = ~n9729 & ~n9730 ;
  assign n9733 = n9731 & n9732 ;
  assign n9734 = n4055 & n9733 ;
  assign n9735 = ~n9726 & ~n9734 ;
  assign n9736 = ~n6135 & n9735 ;
  assign n9754 = n6176 & ~n9736 ;
  assign n9755 = ~n9753 & n9754 ;
  assign n9761 = ~n6774 & ~n6820 ;
  assign n9762 = ~n6819 & ~n9761 ;
  assign n9763 = n6819 & n9761 ;
  assign n9764 = ~n9762 & ~n9763 ;
  assign n9765 = n8198 & n9764 ;
  assign n9756 = \core_dag_ilm2reg_I_reg[4]/NET0131  & n6684 ;
  assign n9757 = ~n6675 & ~n6770 ;
  assign n9758 = n6675 & n6770 ;
  assign n9759 = ~n9757 & ~n9758 ;
  assign n9760 = ~n8198 & n9759 ;
  assign n9766 = ~n9756 & ~n9760 ;
  assign n9767 = ~n9765 & n9766 ;
  assign n9768 = n6135 & ~n9767 ;
  assign n9791 = \core_dag_ilm2reg_I7_we_DO_reg[4]/NET0131  & n6960 ;
  assign n9792 = \core_dag_ilm2reg_I5_we_DO_reg[4]/NET0131  & n6964 ;
  assign n9795 = ~n9791 & ~n9792 ;
  assign n9793 = \core_dag_ilm2reg_I6_we_DO_reg[4]/NET0131  & n6962 ;
  assign n9794 = \core_dag_ilm2reg_I4_we_DO_reg[4]/NET0131  & n6958 ;
  assign n9796 = ~n9793 & ~n9794 ;
  assign n9797 = n9795 & n9796 ;
  assign n9798 = ~n4055 & n9797 ;
  assign n9799 = \core_dag_ilm2reg_I7_we_DO_reg[4]/NET0131  & n6972 ;
  assign n9800 = \core_dag_ilm2reg_I4_we_DO_reg[4]/NET0131  & n6976 ;
  assign n9803 = ~n9799 & ~n9800 ;
  assign n9801 = \core_dag_ilm2reg_I6_we_DO_reg[4]/NET0131  & n6974 ;
  assign n9802 = \core_dag_ilm2reg_I5_we_DO_reg[4]/NET0131  & n6970 ;
  assign n9804 = ~n9801 & ~n9802 ;
  assign n9805 = n9803 & n9804 ;
  assign n9806 = n4055 & n9805 ;
  assign n9807 = ~n9798 & ~n9806 ;
  assign n9808 = ~n6121 & n9807 ;
  assign n9771 = \core_dag_ilm1reg_I0_we_DO_reg[4]/NET0131  & n6058 ;
  assign n9772 = n6060 & n9771 ;
  assign n9776 = ~n4055 & ~n9772 ;
  assign n9775 = \core_dag_ilm1reg_I1_we_DO_reg[4]/NET0131  & n6142 ;
  assign n9773 = \core_dag_ilm1reg_I3_we_DO_reg[4]/NET0131  & n6140 ;
  assign n9774 = \core_dag_ilm1reg_I2_we_DO_reg[4]/NET0131  & n6138 ;
  assign n9777 = ~n9773 & ~n9774 ;
  assign n9778 = ~n9775 & n9777 ;
  assign n9779 = n9776 & n9778 ;
  assign n9780 = \core_dag_ilm1reg_I0_we_DO_reg[4]/NET0131  & n6148 ;
  assign n9781 = \core_dag_ilm1reg_I2_we_DO_reg[4]/NET0131  & n6152 ;
  assign n9784 = ~n9780 & ~n9781 ;
  assign n9782 = \core_dag_ilm1reg_I3_we_DO_reg[4]/NET0131  & n6150 ;
  assign n9783 = \core_dag_ilm1reg_I1_we_DO_reg[4]/NET0131  & n6154 ;
  assign n9785 = ~n9782 & ~n9783 ;
  assign n9786 = n9784 & n9785 ;
  assign n9787 = n4055 & n9786 ;
  assign n9788 = ~n9779 & ~n9787 ;
  assign n9789 = ~n6111 & n9788 ;
  assign n9790 = \core_c_dec_IR_reg[8]/NET0131  & n6956 ;
  assign n9809 = ~n9789 & ~n9790 ;
  assign n9810 = ~n9808 & n9809 ;
  assign n9811 = n5949 & ~n9810 ;
  assign n9770 = \core_dag_ilm1reg_DMA_pi_DO_reg[4]/NET0131  & ~n6934 ;
  assign n9769 = \idma_DCTL_reg[4]/NET0131  & n6926 ;
  assign n9812 = \core_dag_ilm1reg_STAC_pi_DO_reg[4]/NET0131  & n6988 ;
  assign n9813 = ~n9769 & ~n9812 ;
  assign n9814 = ~n9770 & n9813 ;
  assign n9815 = ~n9811 & n9814 ;
  assign n9816 = n6924 & ~n9815 ;
  assign n9817 = \bdma_BIAD_reg[4]/NET0131  & ~n6924 ;
  assign n9818 = ~n9816 & ~n9817 ;
  assign n9819 = ~n6135 & ~n9818 ;
  assign n9820 = ~n6176 & ~n9819 ;
  assign n9821 = ~n9768 & n9820 ;
  assign n9822 = ~n9755 & ~n9821 ;
  assign n9823 = ~n7005 & ~n9822 ;
  assign n10297 = ~n6304 & ~n6505 ;
  assign n10298 = n6304 & n6505 ;
  assign n10299 = ~n10297 & ~n10298 ;
  assign n10300 = n7631 & n10299 ;
  assign n10291 = \core_dag_ilm1reg_I_reg[4]/NET0131  & ~n6280 ;
  assign n10292 = ~n6308 & ~n6378 ;
  assign n10293 = ~n6372 & n10292 ;
  assign n10294 = n6372 & ~n10292 ;
  assign n10295 = ~n10293 & ~n10294 ;
  assign n10296 = ~n7631 & n10295 ;
  assign n10301 = ~n10291 & ~n10296 ;
  assign n10302 = ~n10300 & n10301 ;
  assign n10303 = n6176 & n10302 ;
  assign n10081 = \DM_rd0[9]_pad  & ~n7053 ;
  assign n10075 = \DM_rdm[9]_pad  & n7016 ;
  assign n10086 = ~n7057 & ~n10075 ;
  assign n10078 = \DM_rd6[9]_pad  & n7031 ;
  assign n10079 = \DM_rd7[9]_pad  & n7034 ;
  assign n10087 = ~n10078 & ~n10079 ;
  assign n10088 = n10086 & n10087 ;
  assign n10082 = \DM_rd4[9]_pad  & n7028 ;
  assign n10077 = \DM_rd5[9]_pad  & n7043 ;
  assign n10083 = \DM_rd2[9]_pad  & n7041 ;
  assign n10076 = \DM_rd1[9]_pad  & n7022 ;
  assign n10080 = \DM_rd3[9]_pad  & n7038 ;
  assign n10084 = ~n10076 & ~n10080 ;
  assign n10085 = ~n10083 & n10084 ;
  assign n10089 = ~n10077 & n10085 ;
  assign n10090 = ~n10082 & n10089 ;
  assign n10091 = n10088 & n10090 ;
  assign n10092 = ~n10081 & n10091 ;
  assign n10093 = \regout_STD_C_reg[9]/P0001  & n6988 ;
  assign n10234 = \bdma_BCTL_reg[9]/NET0131  & n7230 ;
  assign n10232 = \tm_tpr_reg_DO_reg[9]/NET0131  & n7293 ;
  assign n10254 = ~n7522 & ~n10232 ;
  assign n10233 = \sport0_regs_SCLKDIVreg_DO_reg[9]/NET0131  & n7256 ;
  assign n10235 = \idma_DOVL_reg[9]/NET0131  & n7532 ;
  assign n10255 = ~n10233 & ~n10235 ;
  assign n10265 = n10254 & n10255 ;
  assign n10249 = \sport0_txctl_Wcnt_reg[1]/NET0131  & n7710 ;
  assign n10250 = \sport1_txctl_Wcnt_reg[1]/NET0131  & n7689 ;
  assign n10266 = ~n10249 & ~n10250 ;
  assign n10267 = n10265 & n10266 ;
  assign n10270 = ~n10234 & n10267 ;
  assign n10236 = \bdma_BIAD_reg[9]/NET0131  & n7234 ;
  assign n10239 = \bdma_BEAD_reg[9]/NET0131  & n7303 ;
  assign n10271 = ~n10236 & ~n10239 ;
  assign n10272 = n10270 & n10271 ;
  assign n10248 = \bdma_BWCOUNT_reg[9]/NET0131  & n7287 ;
  assign n10237 = \bdma_BOVL_reg[9]/NET0131  & n7534 ;
  assign n10247 = \sport0_regs_FSDIVreg_DO_reg[9]/NET0131  & n7259 ;
  assign n10251 = \memc_usysr_DO_reg[9]/NET0131  & n7301 ;
  assign n10260 = ~n10247 & ~n10251 ;
  assign n10252 = \clkc_ckr_reg_DO_reg[9]/NET0131  & n7239 ;
  assign n10253 = \sport1_regs_AUTOreg_DO_reg[9]/NET0131  & n7527 ;
  assign n10261 = ~n10252 & ~n10253 ;
  assign n10262 = n10260 & n10261 ;
  assign n10243 = \sport0_regs_AUTOreg_DO_reg[9]/NET0131  & n7295 ;
  assign n10244 = \sport1_regs_FSDIVreg_DO_reg[9]/NET0131  & n7273 ;
  assign n10258 = ~n10243 & ~n10244 ;
  assign n10245 = \idma_DCTL_reg[9]/NET0131  & n7299 ;
  assign n10246 = \ITFS0_pad  & n7249 ;
  assign n10259 = ~n10245 & ~n10246 ;
  assign n10263 = n10258 & n10259 ;
  assign n10238 = \emc_WSCRreg_DO_reg[9]/NET0131  & n7251 ;
  assign n10240 = \ITFS1_pad  & n7281 ;
  assign n10256 = ~n10238 & ~n10240 ;
  assign n10241 = \sport1_regs_SCLKDIVreg_DO_reg[9]/NET0131  & n7247 ;
  assign n10242 = \tm_TCR_TMP_reg[9]/NET0131  & n7289 ;
  assign n10257 = ~n10241 & ~n10242 ;
  assign n10264 = n10256 & n10257 ;
  assign n10268 = n10263 & n10264 ;
  assign n10269 = n10262 & n10268 ;
  assign n10273 = ~n10237 & n10269 ;
  assign n10274 = ~n10248 & n10273 ;
  assign n10275 = n10272 & n10274 ;
  assign n10276 = \memc_ldSREG_E_reg/NET0131  & ~n10275 ;
  assign n10207 = \core_c_dec_MFtoppcs_Eg_reg/P0001  & ~n4554 ;
  assign n10209 = \core_c_dec_IRE_reg[13]/NET0131  & ~n7216 ;
  assign n10210 = \core_c_dec_MFCNTR_E_reg/P0001  & \core_c_psq_CNTR_reg_DO_reg[9]/NET0131  ;
  assign n10206 = \core_c_dec_MFIDR_E_reg/P0001  & \sice_idr0_reg_DO_reg[9]/P0001  ;
  assign n10208 = \core_c_dec_MFIMASK_E_reg/P0001  & \core_c_psq_IMASK_reg[9]/NET0131  ;
  assign n10211 = ~n10206 & ~n10208 ;
  assign n10212 = ~n10210 & n10211 ;
  assign n10213 = ~n10209 & n10212 ;
  assign n10214 = ~n10207 & n10213 ;
  assign n10215 = n7215 & ~n10214 ;
  assign n10157 = \core_c_dec_MFMreg_E_reg[5]/P0001  & \core_dag_ilm2reg_M5_we_DO_reg[9]/NET0131  ;
  assign n10158 = \core_c_dec_MFLreg_E_reg[5]/P0001  & \core_dag_ilm2reg_L5_we_DO_reg[9]/NET0131  ;
  assign n10165 = ~n10157 & ~n10158 ;
  assign n10159 = \core_c_dec_MFLreg_E_reg[4]/P0001  & \core_dag_ilm2reg_L4_we_DO_reg[9]/NET0131  ;
  assign n10160 = \core_c_dec_MFIreg_E_reg[6]/P0001  & \core_dag_ilm2reg_I6_we_DO_reg[9]/NET0131  ;
  assign n10166 = ~n10159 & ~n10160 ;
  assign n10167 = n10165 & n10166 ;
  assign n10153 = \core_c_dec_MFIreg_E_reg[4]/P0001  & \core_dag_ilm2reg_I4_we_DO_reg[9]/NET0131  ;
  assign n10154 = \core_c_dec_MFIreg_E_reg[5]/P0001  & \core_dag_ilm2reg_I5_we_DO_reg[9]/NET0131  ;
  assign n10163 = ~n10153 & ~n10154 ;
  assign n10155 = \core_c_dec_MFMreg_E_reg[7]/P0001  & \core_dag_ilm2reg_M7_we_DO_reg[9]/NET0131  ;
  assign n10156 = \core_c_dec_MFMreg_E_reg[6]/P0001  & \core_dag_ilm2reg_M6_we_DO_reg[9]/NET0131  ;
  assign n10164 = ~n10155 & ~n10156 ;
  assign n10168 = n10163 & n10164 ;
  assign n10149 = \core_c_dec_MFLreg_E_reg[6]/P0001  & \core_dag_ilm2reg_L6_we_DO_reg[9]/NET0131  ;
  assign n10150 = \core_c_dec_MFMreg_E_reg[4]/P0001  & \core_dag_ilm2reg_M4_we_DO_reg[9]/NET0131  ;
  assign n10161 = ~n10149 & ~n10150 ;
  assign n10151 = \core_c_dec_MFLreg_E_reg[7]/P0001  & \core_dag_ilm2reg_L7_we_DO_reg[9]/NET0131  ;
  assign n10152 = \core_c_dec_MFIreg_E_reg[7]/P0001  & \core_dag_ilm2reg_I7_we_DO_reg[9]/NET0131  ;
  assign n10162 = ~n10151 & ~n10152 ;
  assign n10169 = n10161 & n10162 ;
  assign n10170 = n10168 & n10169 ;
  assign n10171 = n10167 & n10170 ;
  assign n10172 = n7128 & ~n10171 ;
  assign n10133 = \core_c_dec_MFIreg_E_reg[0]/P0001  & \core_dag_ilm1reg_I0_we_DO_reg[9]/NET0131  ;
  assign n10134 = \core_c_dec_MFIreg_E_reg[3]/P0001  & \core_dag_ilm1reg_I3_we_DO_reg[9]/NET0131  ;
  assign n10141 = ~n10133 & ~n10134 ;
  assign n10135 = \core_c_dec_MFLreg_E_reg[0]/P0001  & \core_dag_ilm1reg_L0_we_DO_reg[9]/NET0131  ;
  assign n10136 = \core_c_dec_MFLreg_E_reg[1]/P0001  & \core_dag_ilm1reg_L1_we_DO_reg[9]/NET0131  ;
  assign n10142 = ~n10135 & ~n10136 ;
  assign n10143 = n10141 & n10142 ;
  assign n10129 = \core_c_dec_MFIreg_E_reg[1]/P0001  & \core_dag_ilm1reg_I1_we_DO_reg[9]/NET0131  ;
  assign n10130 = \core_c_dec_MFMreg_E_reg[2]/P0001  & \core_dag_ilm1reg_M2_we_DO_reg[9]/NET0131  ;
  assign n10139 = ~n10129 & ~n10130 ;
  assign n10131 = \core_c_dec_MFIreg_E_reg[2]/P0001  & \core_dag_ilm1reg_I2_we_DO_reg[9]/NET0131  ;
  assign n10132 = \core_c_dec_MFLreg_E_reg[2]/P0001  & \core_dag_ilm1reg_L2_we_DO_reg[9]/NET0131  ;
  assign n10140 = ~n10131 & ~n10132 ;
  assign n10144 = n10139 & n10140 ;
  assign n10125 = \core_c_dec_MFMreg_E_reg[0]/P0001  & \core_dag_ilm1reg_M0_we_DO_reg[9]/NET0131  ;
  assign n10126 = \core_c_dec_MFMreg_E_reg[3]/P0001  & \core_dag_ilm1reg_M3_we_DO_reg[9]/NET0131  ;
  assign n10137 = ~n10125 & ~n10126 ;
  assign n10127 = \core_c_dec_MFLreg_E_reg[3]/P0001  & \core_dag_ilm1reg_L3_we_DO_reg[9]/NET0131  ;
  assign n10128 = \core_c_dec_MFMreg_E_reg[1]/P0001  & \core_dag_ilm1reg_M1_we_DO_reg[9]/NET0131  ;
  assign n10138 = ~n10127 & ~n10128 ;
  assign n10145 = n10137 & n10138 ;
  assign n10146 = n10144 & n10145 ;
  assign n10147 = n10143 & n10146 ;
  assign n10148 = n7068 & ~n10147 ;
  assign n10198 = \core_c_dec_MFTX1_E_reg/P0001  & \sport1_txctl_TX_reg[9]/P0001  ;
  assign n10199 = \core_c_dec_MFRX1_E_reg/P0001  & \sport1_rxctl_RX_reg[9]/P0001  ;
  assign n10202 = ~n10198 & ~n10199 ;
  assign n10200 = \core_c_dec_MFRX0_E_reg/P0001  & \sport0_rxctl_RX_reg[9]/P0001  ;
  assign n10201 = \core_c_dec_MFTX0_E_reg/P0001  & \sport0_txctl_TX_reg[9]/P0001  ;
  assign n10203 = ~n10200 & ~n10201 ;
  assign n10204 = n10202 & n10203 ;
  assign n10205 = n7119 & ~n10204 ;
  assign n10277 = ~n10148 & ~n10205 ;
  assign n10278 = ~n10172 & n10277 ;
  assign n10224 = ~\core_c_psq_MSTAT_reg_DO_reg[0]/P0002  & \core_eu_es_sht_es_reg_sr1rwe_DO_reg[9]/P0001  ;
  assign n10225 = \core_c_psq_MSTAT_reg_DO_reg[0]/P0002  & \core_eu_es_sht_es_reg_sr1swe_DO_reg[9]/P0001  ;
  assign n10226 = ~n10224 & ~n10225 ;
  assign n10227 = \core_c_dec_MFSR1_E_reg/P0001  & ~n10226 ;
  assign n10216 = ~\core_c_psq_MSTAT_reg_DO_reg[0]/P0002  & \core_eu_es_sht_es_reg_sr0rwe_DO_reg[9]/P0001  ;
  assign n10217 = \core_c_psq_MSTAT_reg_DO_reg[0]/P0002  & \core_eu_es_sht_es_reg_sr0swe_DO_reg[9]/P0001  ;
  assign n10218 = ~n10216 & ~n10217 ;
  assign n10219 = \core_c_dec_MFSR0_E_reg/P0001  & ~n10218 ;
  assign n10220 = ~\core_c_psq_MSTAT_reg_DO_reg[0]/P0002  & \core_eu_es_sht_es_reg_sirwe_DO_reg[9]/P0001  ;
  assign n10221 = \core_c_psq_MSTAT_reg_DO_reg[0]/P0002  & \core_eu_es_sht_es_reg_siswe_DO_reg[9]/P0001  ;
  assign n10222 = ~n10220 & ~n10221 ;
  assign n10223 = \core_c_dec_MFSI_E_reg/P0001  & ~n10222 ;
  assign n10228 = ~n10219 & ~n10223 ;
  assign n10229 = ~n10227 & n10228 ;
  assign n10230 = n7174 & n10229 ;
  assign n10231 = n7153 & ~n10230 ;
  assign n10114 = ~\core_c_psq_MSTAT_reg_DO_reg[0]/P0002  & \core_eu_em_mac_em_reg_mx0rwe_DO_reg[9]/P0001  ;
  assign n10115 = \core_c_psq_MSTAT_reg_DO_reg[0]/P0002  & \core_eu_em_mac_em_reg_mx0swe_DO_reg[9]/P0001  ;
  assign n10116 = ~n10114 & ~n10115 ;
  assign n10117 = \core_c_dec_MFMX0_E_reg/P0001  & ~n10116 ;
  assign n10106 = ~\core_c_psq_MSTAT_reg_DO_reg[0]/P0002  & \core_eu_em_mac_em_reg_my1rwe_DO_reg[9]/P0001  ;
  assign n10107 = \core_c_psq_MSTAT_reg_DO_reg[0]/P0002  & \core_eu_em_mac_em_reg_my1swe_DO_reg[9]/P0001  ;
  assign n10108 = ~n10106 & ~n10107 ;
  assign n10109 = \core_c_dec_MFMY1_E_reg/P0001  & ~n10108 ;
  assign n10110 = ~\core_c_psq_MSTAT_reg_DO_reg[0]/P0002  & \core_eu_em_mac_em_reg_mr0rwe_DO_reg[9]/P0001  ;
  assign n10111 = \core_c_psq_MSTAT_reg_DO_reg[0]/P0002  & \core_eu_em_mac_em_reg_mr0swe_DO_reg[9]/P0001  ;
  assign n10112 = ~n10110 & ~n10111 ;
  assign n10113 = \core_c_dec_MFMR0_E_reg/P0001  & ~n10112 ;
  assign n10120 = ~n10109 & ~n10113 ;
  assign n10121 = ~n10117 & n10120 ;
  assign n10094 = ~\core_c_psq_MSTAT_reg_DO_reg[0]/P0002  & \core_eu_em_mac_em_reg_mr1rwe_DO_reg[9]/P0001  ;
  assign n10095 = \core_c_psq_MSTAT_reg_DO_reg[0]/P0002  & \core_eu_em_mac_em_reg_mr1swe_DO_reg[9]/P0001  ;
  assign n10096 = ~n10094 & ~n10095 ;
  assign n10097 = \core_c_dec_MFMR1_E_reg/P0001  & ~n10096 ;
  assign n10118 = ~n7207 & ~n10097 ;
  assign n10098 = ~\core_c_psq_MSTAT_reg_DO_reg[0]/P0002  & \core_eu_em_mac_em_reg_mx1rwe_DO_reg[9]/P0001  ;
  assign n10099 = \core_c_psq_MSTAT_reg_DO_reg[0]/P0002  & \core_eu_em_mac_em_reg_mx1swe_DO_reg[9]/P0001  ;
  assign n10100 = ~n10098 & ~n10099 ;
  assign n10101 = \core_c_dec_MFMX1_E_reg/P0001  & ~n10100 ;
  assign n10102 = ~\core_c_psq_MSTAT_reg_DO_reg[0]/P0002  & \core_eu_em_mac_em_reg_my0rwe_DO_reg[9]/P0001  ;
  assign n10103 = \core_c_psq_MSTAT_reg_DO_reg[0]/P0002  & \core_eu_em_mac_em_reg_my0swe_DO_reg[9]/P0001  ;
  assign n10104 = ~n10102 & ~n10103 ;
  assign n10105 = \core_c_dec_MFMY0_E_reg/P0001  & ~n10104 ;
  assign n10119 = ~n10101 & ~n10105 ;
  assign n10122 = n10118 & n10119 ;
  assign n10123 = n10121 & n10122 ;
  assign n10124 = n7179 & ~n10123 ;
  assign n10173 = ~\core_c_psq_MSTAT_reg_DO_reg[0]/P0002  & \core_eu_ea_alu_ea_reg_ay1rwe_DO_reg[9]/P0001  ;
  assign n10174 = \core_c_psq_MSTAT_reg_DO_reg[0]/P0002  & \core_eu_ea_alu_ea_reg_ay1swe_DO_reg[9]/P0001  ;
  assign n10175 = ~n10173 & ~n10174 ;
  assign n10176 = \core_c_dec_MFAY1_E_reg/P0001  & ~n10175 ;
  assign n10177 = ~\core_c_psq_MSTAT_reg_DO_reg[0]/P0002  & \core_eu_ea_alu_ea_reg_ax1rwe_DO_reg[9]/P0001  ;
  assign n10178 = \core_c_psq_MSTAT_reg_DO_reg[0]/P0002  & \core_eu_ea_alu_ea_reg_ax1swe_DO_reg[9]/P0001  ;
  assign n10179 = ~n10177 & ~n10178 ;
  assign n10180 = \core_c_dec_MFAX1_E_reg/P0001  & ~n10179 ;
  assign n10193 = ~n10176 & ~n10180 ;
  assign n10189 = ~\core_c_psq_MSTAT_reg_DO_reg[0]/P0002  & \core_eu_ea_alu_ea_reg_arrwe_DO_reg[9]/P0001  ;
  assign n10190 = \core_c_psq_MSTAT_reg_DO_reg[0]/P0002  & \core_eu_ea_alu_ea_reg_arswe_DO_reg[9]/P0001  ;
  assign n10191 = ~n10189 & ~n10190 ;
  assign n10192 = \core_c_dec_MFAR_E_reg/P0001  & ~n10191 ;
  assign n10181 = ~\core_c_psq_MSTAT_reg_DO_reg[0]/P0002  & \core_eu_ea_alu_ea_reg_ay0rwe_DO_reg[9]/P0001  ;
  assign n10182 = \core_c_psq_MSTAT_reg_DO_reg[0]/P0002  & \core_eu_ea_alu_ea_reg_ay0swe_DO_reg[9]/P0001  ;
  assign n10183 = ~n10181 & ~n10182 ;
  assign n10184 = \core_c_dec_MFAY0_E_reg/P0001  & ~n10183 ;
  assign n10185 = ~\core_c_psq_MSTAT_reg_DO_reg[0]/P0002  & \core_eu_ea_alu_ea_reg_ax0rwe_DO_reg[9]/P0001  ;
  assign n10186 = \core_c_psq_MSTAT_reg_DO_reg[0]/P0002  & \core_eu_ea_alu_ea_reg_ax0swe_DO_reg[9]/P0001  ;
  assign n10187 = ~n10185 & ~n10186 ;
  assign n10188 = \core_c_dec_MFAX0_E_reg/P0001  & ~n10187 ;
  assign n10194 = ~n10184 & ~n10188 ;
  assign n10195 = ~n10192 & n10194 ;
  assign n10196 = n10193 & n10195 ;
  assign n10197 = n7093 & ~n10196 ;
  assign n10279 = ~n10124 & ~n10197 ;
  assign n10280 = ~n10231 & n10279 ;
  assign n10281 = n10278 & n10280 ;
  assign n10282 = ~n10215 & n10281 ;
  assign n10283 = ~n10276 & n10282 ;
  assign n10284 = ~n10093 & n10283 ;
  assign n10285 = ~\emc_DMDoe_reg/NET0131  & ~n10284 ;
  assign n10286 = \emc_DMDoe_reg/NET0131  & \emc_DMDreg_reg[9]/P0001  ;
  assign n10287 = n7057 & ~n10286 ;
  assign n10288 = ~n10285 & n10287 ;
  assign n10289 = ~n10092 & ~n10288 ;
  assign n10290 = ~n6176 & ~n10289 ;
  assign n10304 = ~n6135 & ~n10290 ;
  assign n10305 = ~n10303 & n10304 ;
  assign n10071 = ~n9788 & ~n9807 ;
  assign n10072 = ~n6176 & n10071 ;
  assign n9830 = \DM_rd0[4]_pad  & ~n7053 ;
  assign n9824 = \DM_rdm[4]_pad  & n7016 ;
  assign n9835 = ~n7057 & ~n9824 ;
  assign n9827 = \DM_rd6[4]_pad  & n7031 ;
  assign n9828 = \DM_rd7[4]_pad  & n7034 ;
  assign n9836 = ~n9827 & ~n9828 ;
  assign n9837 = n9835 & n9836 ;
  assign n9831 = \DM_rd5[4]_pad  & n7043 ;
  assign n9826 = \DM_rd4[4]_pad  & n7028 ;
  assign n9832 = \DM_rd2[4]_pad  & n7041 ;
  assign n9825 = \DM_rd1[4]_pad  & n7022 ;
  assign n9829 = \DM_rd3[4]_pad  & n7038 ;
  assign n9833 = ~n9825 & ~n9829 ;
  assign n9834 = ~n9832 & n9833 ;
  assign n9838 = ~n9826 & n9834 ;
  assign n9839 = ~n9831 & n9838 ;
  assign n9840 = n9837 & n9839 ;
  assign n9841 = ~n9830 & n9840 ;
  assign n9842 = \regout_STD_C_reg[4]/P0001  & n6988 ;
  assign n9995 = \bdma_BIAD_reg[4]/NET0131  & n7234 ;
  assign n9986 = \emc_WSCRreg_DO_reg[4]/NET0131  & n7251 ;
  assign n9987 = \sport0_regs_SCLKDIVreg_DO_reg[4]/NET0131  & n7256 ;
  assign n10012 = ~n9986 & ~n9987 ;
  assign n9988 = \sport1_regs_MWORDreg_DO_reg[4]/NET0131  & n7263 ;
  assign n9989 = \tm_tsr_reg_DO_reg[4]/NET0131  & n7540 ;
  assign n10013 = ~n9988 & ~n9989 ;
  assign n10026 = n10012 & n10013 ;
  assign n9982 = \idma_DOVL_reg[4]/NET0131  & n7532 ;
  assign n10010 = ~n7522 & ~n9982 ;
  assign n9983 = \sport0_regs_AUTOreg_DO_reg[4]/NET0131  & n7295 ;
  assign n9984 = \tm_tpr_reg_DO_reg[4]/NET0131  & n7293 ;
  assign n10011 = ~n9983 & ~n9984 ;
  assign n10027 = n10010 & n10011 ;
  assign n10028 = n10026 & n10027 ;
  assign n10032 = ~n9995 & n10028 ;
  assign n10003 = \bdma_BEAD_reg[4]/NET0131  & n7303 ;
  assign n10004 = \bdma_BCTL_reg[4]/NET0131  & n7230 ;
  assign n10033 = ~n10003 & ~n10004 ;
  assign n10034 = n10032 & n10033 ;
  assign n10000 = \bdma_BOVL_reg[4]/NET0131  & n7534 ;
  assign n9985 = \bdma_BWCOUNT_reg[4]/NET0131  & n7287 ;
  assign n9994 = \pio_pmask_reg_DO_reg[4]/NET0131  & n7297 ;
  assign n9996 = \sport0_regs_MWORDreg_DO_reg[4]/NET0131  & n7276 ;
  assign n10016 = ~n9994 & ~n9996 ;
  assign n9997 = \sport1_regs_AUTOreg_DO_reg[4]/NET0131  & n7527 ;
  assign n9998 = \tm_TCR_TMP_reg[4]/NET0131  & n7289 ;
  assign n10017 = ~n9997 & ~n9998 ;
  assign n10024 = n10016 & n10017 ;
  assign n9990 = \sport0_regs_SCTLreg_DO_reg[4]/NET0131  & n7249 ;
  assign n9991 = \emc_WSCRext_reg_DO_reg[4]/NET0131  & n7514 ;
  assign n10014 = ~n9990 & ~n9991 ;
  assign n9992 = \sport1_regs_SCLKDIVreg_DO_reg[4]/NET0131  & n7247 ;
  assign n9993 = \sport1_regs_SCTLreg_DO_reg[4]/NET0131  & n7281 ;
  assign n10015 = ~n9992 & ~n9993 ;
  assign n10025 = n10014 & n10015 ;
  assign n10029 = n10024 & n10025 ;
  assign n10006 = \idma_DCTL_reg[4]/NET0131  & n7299 ;
  assign n10007 = \PIO_out[4]_pad  & n7291 ;
  assign n10020 = ~n10006 & ~n10007 ;
  assign n10008 = \PIO_oe[4]_pad  & n7244 ;
  assign n10009 = \sport1_regs_FSDIVreg_DO_reg[4]/NET0131  & n7273 ;
  assign n10021 = ~n10008 & ~n10009 ;
  assign n10022 = n10020 & n10021 ;
  assign n9999 = \sport0_regs_FSDIVreg_DO_reg[4]/NET0131  & n7259 ;
  assign n10001 = \clkc_ckr_reg_DO_reg[4]/NET0131  & n7239 ;
  assign n10018 = ~n9999 & ~n10001 ;
  assign n10002 = \memc_usysr_DO_reg[4]/NET0131  & n7301 ;
  assign n10005 = \pio_PINT_reg[4]/NET0131  & n7271 ;
  assign n10019 = ~n10002 & ~n10005 ;
  assign n10023 = n10018 & n10019 ;
  assign n10030 = n10022 & n10023 ;
  assign n10031 = n10029 & n10030 ;
  assign n10035 = ~n9985 & n10031 ;
  assign n10036 = ~n10000 & n10035 ;
  assign n10037 = n10034 & n10036 ;
  assign n10038 = \memc_ldSREG_E_reg/NET0131  & ~n10037 ;
  assign n10042 = \core_c_dec_MFtoppcs_Eg_reg/P0001  & ~n4360 ;
  assign n10047 = \core_c_dec_MFSSTAT_E_reg/P0001  & \core_c_psq_SSTAT_reg[4]/NET0131  ;
  assign n10045 = \core_c_dec_MFPMOVL_E_reg/P0001  & \core_c_psq_PMOVL_regh_DO_reg[0]/NET0131  ;
  assign n10046 = \core_c_dec_MFCNTR_E_reg/P0001  & \core_c_psq_CNTR_reg_DO_reg[4]/NET0131  ;
  assign n10050 = ~n10045 & ~n10046 ;
  assign n10051 = ~n10047 & n10050 ;
  assign n10040 = \core_c_dec_IRE_reg[8]/NET0131  & ~n7216 ;
  assign n10039 = \core_c_dec_MFICNTL_E_reg/P0001  & \core_c_psq_ICNTL_reg_DO_reg[4]/NET0131  ;
  assign n10041 = \core_c_dec_MFIDR_E_reg/P0001  & \sice_idr0_reg_DO_reg[4]/P0001  ;
  assign n10048 = ~n10039 & ~n10041 ;
  assign n10043 = \core_c_dec_MFMSTAT_E_reg/P0001  & \core_c_psq_MSTAT_reg_DO_reg[4]/NET0131  ;
  assign n10044 = \core_c_dec_MFIMASK_E_reg/P0001  & \core_c_psq_IMASK_reg[4]/NET0131  ;
  assign n10049 = ~n10043 & ~n10044 ;
  assign n10052 = n10048 & n10049 ;
  assign n10053 = ~n10040 & n10052 ;
  assign n10054 = n10051 & n10053 ;
  assign n10055 = ~n10042 & n10054 ;
  assign n10056 = n7215 & ~n10055 ;
  assign n9966 = \core_c_dec_MFLreg_E_reg[6]/P0001  & \core_dag_ilm2reg_L6_we_DO_reg[4]/NET0131  ;
  assign n9967 = \core_c_dec_MFMreg_E_reg[5]/P0001  & \core_dag_ilm2reg_M5_we_DO_reg[4]/NET0131  ;
  assign n9974 = ~n9966 & ~n9967 ;
  assign n9968 = \core_c_dec_MFMreg_E_reg[6]/P0001  & \core_dag_ilm2reg_M6_we_DO_reg[4]/NET0131  ;
  assign n9969 = \core_c_dec_MFMreg_E_reg[7]/P0001  & \core_dag_ilm2reg_M7_we_DO_reg[4]/NET0131  ;
  assign n9975 = ~n9968 & ~n9969 ;
  assign n9976 = n9974 & n9975 ;
  assign n9962 = \core_c_dec_MFLreg_E_reg[7]/P0001  & \core_dag_ilm2reg_L7_we_DO_reg[4]/NET0131  ;
  assign n9963 = \core_c_dec_MFMreg_E_reg[4]/P0001  & \core_dag_ilm2reg_M4_we_DO_reg[4]/NET0131  ;
  assign n9972 = ~n9962 & ~n9963 ;
  assign n9964 = \core_c_dec_MFIreg_E_reg[5]/P0001  & \core_dag_ilm2reg_I5_we_DO_reg[4]/NET0131  ;
  assign n9965 = \core_c_dec_MFIreg_E_reg[6]/P0001  & \core_dag_ilm2reg_I6_we_DO_reg[4]/NET0131  ;
  assign n9973 = ~n9964 & ~n9965 ;
  assign n9977 = n9972 & n9973 ;
  assign n9958 = \core_c_dec_MFIreg_E_reg[4]/P0001  & \core_dag_ilm2reg_I4_we_DO_reg[4]/NET0131  ;
  assign n9959 = \core_c_dec_MFIreg_E_reg[7]/P0001  & \core_dag_ilm2reg_I7_we_DO_reg[4]/NET0131  ;
  assign n9970 = ~n9958 & ~n9959 ;
  assign n9960 = \core_c_dec_MFLreg_E_reg[4]/P0001  & \core_dag_ilm2reg_L4_we_DO_reg[4]/NET0131  ;
  assign n9961 = \core_c_dec_MFLreg_E_reg[5]/P0001  & \core_dag_ilm2reg_L5_we_DO_reg[4]/NET0131  ;
  assign n9971 = ~n9960 & ~n9961 ;
  assign n9978 = n9970 & n9971 ;
  assign n9979 = n9977 & n9978 ;
  assign n9980 = n9976 & n9979 ;
  assign n9981 = n7128 & ~n9980 ;
  assign n9886 = \core_c_dec_MFIreg_E_reg[3]/P0001  & \core_dag_ilm1reg_I3_we_DO_reg[4]/NET0131  ;
  assign n9887 = \core_c_dec_MFIreg_E_reg[0]/P0001  & \core_dag_ilm1reg_I0_we_DO_reg[4]/NET0131  ;
  assign n9894 = ~n9886 & ~n9887 ;
  assign n9888 = \core_c_dec_MFIreg_E_reg[1]/P0001  & \core_dag_ilm1reg_I1_we_DO_reg[4]/NET0131  ;
  assign n9889 = \core_c_dec_MFIreg_E_reg[2]/P0001  & \core_dag_ilm1reg_I2_we_DO_reg[4]/NET0131  ;
  assign n9895 = ~n9888 & ~n9889 ;
  assign n9896 = n9894 & n9895 ;
  assign n9882 = \core_c_dec_MFLreg_E_reg[0]/P0001  & \core_dag_ilm1reg_L0_we_DO_reg[4]/NET0131  ;
  assign n9883 = \core_c_dec_MFLreg_E_reg[1]/P0001  & \core_dag_ilm1reg_L1_we_DO_reg[4]/NET0131  ;
  assign n9892 = ~n9882 & ~n9883 ;
  assign n9884 = \core_c_dec_MFMreg_E_reg[2]/P0001  & \core_dag_ilm1reg_M2_we_DO_reg[4]/NET0131  ;
  assign n9885 = \core_c_dec_MFMreg_E_reg[3]/P0001  & \core_dag_ilm1reg_M3_we_DO_reg[4]/NET0131  ;
  assign n9893 = ~n9884 & ~n9885 ;
  assign n9897 = n9892 & n9893 ;
  assign n9878 = \core_c_dec_MFMreg_E_reg[1]/P0001  & \core_dag_ilm1reg_M1_we_DO_reg[4]/NET0131  ;
  assign n9879 = \core_c_dec_MFLreg_E_reg[2]/P0001  & \core_dag_ilm1reg_L2_we_DO_reg[4]/NET0131  ;
  assign n9890 = ~n9878 & ~n9879 ;
  assign n9880 = \core_c_dec_MFLreg_E_reg[3]/P0001  & \core_dag_ilm1reg_L3_we_DO_reg[4]/NET0131  ;
  assign n9881 = \core_c_dec_MFMreg_E_reg[0]/P0001  & \core_dag_ilm1reg_M0_we_DO_reg[4]/NET0131  ;
  assign n9891 = ~n9880 & ~n9881 ;
  assign n9898 = n9890 & n9891 ;
  assign n9899 = n9897 & n9898 ;
  assign n9900 = n9896 & n9899 ;
  assign n9901 = n7068 & ~n9900 ;
  assign n9929 = \core_c_dec_MFTX1_E_reg/P0001  & \sport1_txctl_TX_reg[4]/P0001  ;
  assign n9930 = \core_c_dec_MFTX0_E_reg/P0001  & \sport0_txctl_TX_reg[4]/P0001  ;
  assign n9933 = ~n9929 & ~n9930 ;
  assign n9931 = \core_c_dec_MFRX1_E_reg/P0001  & \sport1_rxctl_RX_reg[4]/P0001  ;
  assign n9932 = \core_c_dec_MFRX0_E_reg/P0001  & \sport0_rxctl_RX_reg[4]/P0001  ;
  assign n9934 = ~n9931 & ~n9932 ;
  assign n9935 = n9933 & n9934 ;
  assign n9936 = n7119 & ~n9935 ;
  assign n10057 = ~n9901 & ~n9936 ;
  assign n10058 = ~n9981 & n10057 ;
  assign n9937 = ~\core_c_psq_MSTAT_reg_DO_reg[0]/P0002  & \core_eu_es_sht_es_reg_serwe_DO_reg[4]/P0001  ;
  assign n9938 = \core_c_psq_MSTAT_reg_DO_reg[0]/P0002  & \core_eu_es_sht_es_reg_seswe_DO_reg[4]/P0001  ;
  assign n9939 = ~n9937 & ~n9938 ;
  assign n9940 = \core_c_dec_MFSE_E_reg/P0001  & ~n9939 ;
  assign n9953 = ~n7169 & ~n9940 ;
  assign n9949 = ~\core_c_psq_MSTAT_reg_DO_reg[0]/P0002  & \core_eu_es_sht_es_reg_sr0rwe_DO_reg[4]/P0001  ;
  assign n9950 = \core_c_psq_MSTAT_reg_DO_reg[0]/P0002  & \core_eu_es_sht_es_reg_sr0swe_DO_reg[4]/P0001  ;
  assign n9951 = ~n9949 & ~n9950 ;
  assign n9952 = \core_c_dec_MFSR0_E_reg/P0001  & ~n9951 ;
  assign n9941 = ~\core_c_psq_MSTAT_reg_DO_reg[0]/P0002  & \core_eu_es_sht_es_reg_sirwe_DO_reg[4]/P0001  ;
  assign n9942 = \core_c_psq_MSTAT_reg_DO_reg[0]/P0002  & \core_eu_es_sht_es_reg_siswe_DO_reg[4]/P0001  ;
  assign n9943 = ~n9941 & ~n9942 ;
  assign n9944 = \core_c_dec_MFSI_E_reg/P0001  & ~n9943 ;
  assign n9945 = ~\core_c_psq_MSTAT_reg_DO_reg[0]/P0002  & \core_eu_es_sht_es_reg_sr1rwe_DO_reg[4]/P0001  ;
  assign n9946 = \core_c_psq_MSTAT_reg_DO_reg[0]/P0002  & \core_eu_es_sht_es_reg_sr1swe_DO_reg[4]/P0001  ;
  assign n9947 = ~n9945 & ~n9946 ;
  assign n9948 = \core_c_dec_MFSR1_E_reg/P0001  & ~n9947 ;
  assign n9954 = ~n9944 & ~n9948 ;
  assign n9955 = ~n9952 & n9954 ;
  assign n9956 = n9953 & n9955 ;
  assign n9957 = n7153 & ~n9956 ;
  assign n9867 = ~\core_c_psq_MSTAT_reg_DO_reg[0]/P0002  & \core_eu_em_mac_em_reg_mr0rwe_DO_reg[4]/P0001  ;
  assign n9868 = \core_c_psq_MSTAT_reg_DO_reg[0]/P0002  & \core_eu_em_mac_em_reg_mr0swe_DO_reg[4]/P0001  ;
  assign n9869 = ~n9867 & ~n9868 ;
  assign n9870 = \core_c_dec_MFMR0_E_reg/P0001  & ~n9869 ;
  assign n9859 = ~\core_c_psq_MSTAT_reg_DO_reg[0]/P0002  & \core_eu_em_mac_em_reg_mx0rwe_DO_reg[4]/P0001  ;
  assign n9860 = \core_c_psq_MSTAT_reg_DO_reg[0]/P0002  & \core_eu_em_mac_em_reg_mx0swe_DO_reg[4]/P0001  ;
  assign n9861 = ~n9859 & ~n9860 ;
  assign n9862 = \core_c_dec_MFMX0_E_reg/P0001  & ~n9861 ;
  assign n9863 = ~\core_c_psq_MSTAT_reg_DO_reg[0]/P0002  & \core_eu_em_mac_em_reg_mr2rwe_DO_reg[4]/P0001  ;
  assign n9864 = \core_c_psq_MSTAT_reg_DO_reg[0]/P0002  & \core_eu_em_mac_em_reg_mr2swe_DO_reg[4]/P0001  ;
  assign n9865 = ~n9863 & ~n9864 ;
  assign n9866 = \core_c_dec_MFMR2_E_reg/P0001  & ~n9865 ;
  assign n9873 = ~n9862 & ~n9866 ;
  assign n9874 = ~n9870 & n9873 ;
  assign n9843 = ~\core_c_psq_MSTAT_reg_DO_reg[0]/P0002  & \core_eu_em_mac_em_reg_mr1rwe_DO_reg[4]/P0001  ;
  assign n9844 = \core_c_psq_MSTAT_reg_DO_reg[0]/P0002  & \core_eu_em_mac_em_reg_mr1swe_DO_reg[4]/P0001  ;
  assign n9845 = ~n9843 & ~n9844 ;
  assign n9846 = \core_c_dec_MFMR1_E_reg/P0001  & ~n9845 ;
  assign n9847 = ~\core_c_psq_MSTAT_reg_DO_reg[0]/P0002  & \core_eu_em_mac_em_reg_mx1rwe_DO_reg[4]/P0001  ;
  assign n9848 = \core_c_psq_MSTAT_reg_DO_reg[0]/P0002  & \core_eu_em_mac_em_reg_mx1swe_DO_reg[4]/P0001  ;
  assign n9849 = ~n9847 & ~n9848 ;
  assign n9850 = \core_c_dec_MFMX1_E_reg/P0001  & ~n9849 ;
  assign n9871 = ~n9846 & ~n9850 ;
  assign n9851 = ~\core_c_psq_MSTAT_reg_DO_reg[0]/P0002  & \core_eu_em_mac_em_reg_my0rwe_DO_reg[4]/P0001  ;
  assign n9852 = \core_c_psq_MSTAT_reg_DO_reg[0]/P0002  & \core_eu_em_mac_em_reg_my0swe_DO_reg[4]/P0001  ;
  assign n9853 = ~n9851 & ~n9852 ;
  assign n9854 = \core_c_dec_MFMY0_E_reg/P0001  & ~n9853 ;
  assign n9855 = ~\core_c_psq_MSTAT_reg_DO_reg[0]/P0002  & \core_eu_em_mac_em_reg_my1rwe_DO_reg[4]/P0001  ;
  assign n9856 = \core_c_psq_MSTAT_reg_DO_reg[0]/P0002  & \core_eu_em_mac_em_reg_my1swe_DO_reg[4]/P0001  ;
  assign n9857 = ~n9855 & ~n9856 ;
  assign n9858 = \core_c_dec_MFMY1_E_reg/P0001  & ~n9857 ;
  assign n9872 = ~n9854 & ~n9858 ;
  assign n9875 = n9871 & n9872 ;
  assign n9876 = n9874 & n9875 ;
  assign n9877 = n7179 & ~n9876 ;
  assign n9902 = ~\core_c_psq_MSTAT_reg_DO_reg[0]/P0002  & \core_eu_ea_alu_ea_reg_ay0rwe_DO_reg[4]/P0001  ;
  assign n9903 = \core_c_psq_MSTAT_reg_DO_reg[0]/P0002  & \core_eu_ea_alu_ea_reg_ay0swe_DO_reg[4]/P0001  ;
  assign n9904 = ~n9902 & ~n9903 ;
  assign n9905 = \core_c_dec_MFAY0_E_reg/P0001  & ~n9904 ;
  assign n9922 = \core_c_dec_MFASTAT_E_reg/P0001  & \core_eu_ec_cun_AS_reg/P0001  ;
  assign n9923 = ~n9905 & ~n9922 ;
  assign n9906 = ~\core_c_psq_MSTAT_reg_DO_reg[0]/P0002  & \core_eu_ea_alu_ea_reg_ay1rwe_DO_reg[4]/P0001  ;
  assign n9907 = \core_c_psq_MSTAT_reg_DO_reg[0]/P0002  & \core_eu_ea_alu_ea_reg_ay1swe_DO_reg[4]/P0001  ;
  assign n9908 = ~n9906 & ~n9907 ;
  assign n9909 = \core_c_dec_MFAY1_E_reg/P0001  & ~n9908 ;
  assign n9910 = ~\core_c_psq_MSTAT_reg_DO_reg[0]/P0002  & \core_eu_ea_alu_ea_reg_arrwe_DO_reg[4]/P0001  ;
  assign n9911 = \core_c_psq_MSTAT_reg_DO_reg[0]/P0002  & \core_eu_ea_alu_ea_reg_arswe_DO_reg[4]/P0001  ;
  assign n9912 = ~n9910 & ~n9911 ;
  assign n9913 = \core_c_dec_MFAR_E_reg/P0001  & ~n9912 ;
  assign n9924 = ~n9909 & ~n9913 ;
  assign n9914 = ~\core_c_psq_MSTAT_reg_DO_reg[0]/P0002  & \core_eu_ea_alu_ea_reg_ax1rwe_DO_reg[4]/P0001  ;
  assign n9915 = \core_c_psq_MSTAT_reg_DO_reg[0]/P0002  & \core_eu_ea_alu_ea_reg_ax1swe_DO_reg[4]/P0001  ;
  assign n9916 = ~n9914 & ~n9915 ;
  assign n9917 = \core_c_dec_MFAX1_E_reg/P0001  & ~n9916 ;
  assign n9918 = ~\core_c_psq_MSTAT_reg_DO_reg[0]/P0002  & \core_eu_ea_alu_ea_reg_ax0rwe_DO_reg[4]/P0001  ;
  assign n9919 = \core_c_psq_MSTAT_reg_DO_reg[0]/P0002  & \core_eu_ea_alu_ea_reg_ax0swe_DO_reg[4]/P0001  ;
  assign n9920 = ~n9918 & ~n9919 ;
  assign n9921 = \core_c_dec_MFAX0_E_reg/P0001  & ~n9920 ;
  assign n9925 = ~n9917 & ~n9921 ;
  assign n9926 = n9924 & n9925 ;
  assign n9927 = n9923 & n9926 ;
  assign n9928 = n7093 & ~n9927 ;
  assign n10059 = ~n9877 & ~n9928 ;
  assign n10060 = ~n9957 & n10059 ;
  assign n10061 = n10058 & n10060 ;
  assign n10062 = ~n10056 & n10061 ;
  assign n10063 = ~n10038 & n10062 ;
  assign n10064 = ~n9842 & n10063 ;
  assign n10065 = ~\emc_DMDoe_reg/NET0131  & ~n10064 ;
  assign n10066 = \emc_DMDoe_reg/NET0131  & \emc_DMDreg_reg[4]/P0001  ;
  assign n10067 = n7057 & ~n10066 ;
  assign n10068 = ~n10065 & n10067 ;
  assign n10069 = ~n9841 & ~n10068 ;
  assign n10070 = n6176 & ~n10069 ;
  assign n10073 = n6135 & ~n10070 ;
  assign n10074 = ~n10072 & n10073 ;
  assign n10306 = n7005 & ~n10074 ;
  assign n10307 = ~n10305 & n10306 ;
  assign n10308 = ~n9823 & ~n10307 ;
  assign n10316 = ~n6763 & ~n6764 ;
  assign n10317 = ~n6774 & ~n6819 ;
  assign n10318 = ~n6820 & ~n10317 ;
  assign n10319 = ~n10316 & ~n10318 ;
  assign n10320 = n10316 & n10318 ;
  assign n10321 = ~n10319 & ~n10320 ;
  assign n10322 = n8198 & n10321 ;
  assign n10309 = \core_dag_ilm2reg_I_reg[5]/NET0131  & n6680 ;
  assign n10310 = ~n6675 & ~n6690 ;
  assign n10311 = ~n6686 & ~n10310 ;
  assign n10312 = ~n6759 & ~n10311 ;
  assign n10313 = n6759 & n10311 ;
  assign n10314 = ~n10312 & ~n10313 ;
  assign n10315 = ~n8198 & n10314 ;
  assign n10323 = ~n10309 & ~n10315 ;
  assign n10324 = ~n10322 & n10323 ;
  assign n10325 = ~n6176 & n10324 ;
  assign n10331 = ~n6417 & ~n6459 ;
  assign n10332 = ~n6385 & n10331 ;
  assign n10333 = n6385 & ~n10331 ;
  assign n10334 = ~n10332 & ~n10333 ;
  assign n10339 = n6496 & ~n10334 ;
  assign n10327 = ~n6413 & n6514 ;
  assign n10328 = n6413 & ~n6514 ;
  assign n10329 = ~n10327 & ~n10328 ;
  assign n10338 = ~n6496 & n10329 ;
  assign n10340 = ~\core_dag_ilm1reg_M_reg[13]/NET0131  & ~n10338 ;
  assign n10341 = ~n10339 & n10340 ;
  assign n10326 = \core_dag_ilm1reg_I_reg[8]/NET0131  & n6401 ;
  assign n10335 = ~n7612 & ~n10334 ;
  assign n10330 = n7612 & n10329 ;
  assign n10336 = \core_dag_ilm1reg_M_reg[13]/NET0131  & ~n10330 ;
  assign n10337 = ~n10335 & n10336 ;
  assign n10342 = ~n10326 & ~n10337 ;
  assign n10343 = ~n10341 & n10342 ;
  assign n10344 = n6176 & n10343 ;
  assign n10345 = ~n10325 & ~n10344 ;
  assign n10346 = n6135 & ~n10345 ;
  assign n10368 = \core_dag_ilm1reg_I1_we_DO_reg[5]/NET0131  & n6142 ;
  assign n10374 = ~n4055 & ~n10368 ;
  assign n10373 = \core_dag_ilm1reg_I3_we_DO_reg[5]/NET0131  & n6140 ;
  assign n10369 = \core_dag_ilm1reg_I0_we_DO_reg[5]/NET0131  & n6058 ;
  assign n10370 = n6060 & n10369 ;
  assign n10371 = \core_dag_ilm1reg_I2_we_DO_reg[5]/NET0131  & n6084 ;
  assign n10372 = n6085 & n10371 ;
  assign n10375 = ~n10370 & ~n10372 ;
  assign n10376 = ~n10373 & n10375 ;
  assign n10377 = n10374 & n10376 ;
  assign n10378 = n6095 & n10371 ;
  assign n10379 = \core_dag_ilm1reg_I3_we_DO_reg[5]/NET0131  & n6150 ;
  assign n10382 = ~n10378 & ~n10379 ;
  assign n10380 = \core_dag_ilm1reg_I0_we_DO_reg[5]/NET0131  & n6148 ;
  assign n10381 = \core_dag_ilm1reg_I1_we_DO_reg[5]/NET0131  & n6154 ;
  assign n10383 = ~n10380 & ~n10381 ;
  assign n10384 = n10382 & n10383 ;
  assign n10385 = n4055 & n10384 ;
  assign n10386 = ~n10377 & ~n10385 ;
  assign n10387 = ~n6111 & n10386 ;
  assign n10350 = \core_dag_ilm2reg_I4_we_DO_reg[5]/NET0131  & n6976 ;
  assign n10351 = \core_dag_ilm2reg_I7_we_DO_reg[5]/NET0131  & n6972 ;
  assign n10354 = ~n10350 & ~n10351 ;
  assign n10352 = \core_dag_ilm2reg_I6_we_DO_reg[5]/NET0131  & n6974 ;
  assign n10353 = \core_dag_ilm2reg_I5_we_DO_reg[5]/NET0131  & n6970 ;
  assign n10355 = ~n10352 & ~n10353 ;
  assign n10356 = n10354 & n10355 ;
  assign n10357 = n4055 & ~n10356 ;
  assign n10358 = \core_dag_ilm2reg_I7_we_DO_reg[5]/NET0131  & n6960 ;
  assign n10359 = \core_dag_ilm2reg_I4_we_DO_reg[5]/NET0131  & n6958 ;
  assign n10362 = ~n10358 & ~n10359 ;
  assign n10360 = \core_dag_ilm2reg_I6_we_DO_reg[5]/NET0131  & n6962 ;
  assign n10361 = \core_dag_ilm2reg_I5_we_DO_reg[5]/NET0131  & n6964 ;
  assign n10363 = ~n10360 & ~n10361 ;
  assign n10364 = n10362 & n10363 ;
  assign n10365 = ~n10357 & n10364 ;
  assign n10366 = ~n6121 & ~n10365 ;
  assign n10367 = \core_c_dec_IR_reg[9]/NET0131  & n6956 ;
  assign n10388 = ~n10366 & ~n10367 ;
  assign n10389 = ~n10387 & n10388 ;
  assign n10390 = n5949 & ~n10389 ;
  assign n10391 = \core_dag_ilm1reg_DMA_pi_DO_reg[5]/NET0131  & ~n6934 ;
  assign n10348 = \idma_DCTL_reg[5]/NET0131  & n6926 ;
  assign n10349 = \core_dag_ilm1reg_STAC_pi_DO_reg[5]/NET0131  & n6988 ;
  assign n10392 = ~n10348 & ~n10349 ;
  assign n10393 = n6924 & n10392 ;
  assign n10394 = ~n10391 & n10393 ;
  assign n10395 = ~n10390 & n10394 ;
  assign n10347 = ~\bdma_BIAD_reg[5]/NET0131  & ~n6924 ;
  assign n10396 = ~n6176 & ~n10347 ;
  assign n10397 = ~n10395 & n10396 ;
  assign n10398 = \core_dag_ilm1reg_I2_we_DO_reg[8]/NET0131  & n6084 ;
  assign n10399 = n6085 & n10398 ;
  assign n10404 = ~n4055 & ~n10399 ;
  assign n10402 = \core_dag_ilm1reg_I1_we_DO_reg[8]/NET0131  & n6067 ;
  assign n10403 = n6068 & n10402 ;
  assign n10400 = \core_dag_ilm1reg_I3_we_DO_reg[8]/NET0131  & n6140 ;
  assign n10401 = \core_dag_ilm1reg_I0_we_DO_reg[8]/NET0131  & n8131 ;
  assign n10405 = ~n10400 & ~n10401 ;
  assign n10406 = ~n10403 & n10405 ;
  assign n10407 = n10404 & n10406 ;
  assign n10408 = n6091 & n10402 ;
  assign n10409 = \core_dag_ilm1reg_I3_we_DO_reg[8]/NET0131  & n6150 ;
  assign n10412 = ~n10408 & ~n10409 ;
  assign n10410 = \core_dag_ilm1reg_I0_we_DO_reg[8]/NET0131  & n6148 ;
  assign n10411 = \core_dag_ilm1reg_I2_we_DO_reg[8]/NET0131  & n6152 ;
  assign n10413 = ~n10410 & ~n10411 ;
  assign n10414 = n10412 & n10413 ;
  assign n10415 = n4055 & n10414 ;
  assign n10416 = ~n10407 & ~n10415 ;
  assign n10417 = n6176 & n10416 ;
  assign n10418 = ~n6135 & ~n10417 ;
  assign n10419 = ~n10397 & n10418 ;
  assign n10420 = ~n7005 & ~n10419 ;
  assign n10421 = ~n10346 & n10420 ;
  assign n10422 = n10365 & ~n10386 ;
  assign n10423 = n8153 & ~n10422 ;
  assign n10430 = \DM_rd0[8]_pad  & ~n7053 ;
  assign n10424 = \DM_rdm[8]_pad  & n7016 ;
  assign n10435 = ~n7057 & ~n10424 ;
  assign n10427 = \DM_rd6[8]_pad  & n7031 ;
  assign n10428 = \DM_rd7[8]_pad  & n7034 ;
  assign n10436 = ~n10427 & ~n10428 ;
  assign n10437 = n10435 & n10436 ;
  assign n10431 = \DM_rd5[8]_pad  & n7043 ;
  assign n10426 = \DM_rd4[8]_pad  & n7028 ;
  assign n10432 = \DM_rd2[8]_pad  & n7041 ;
  assign n10425 = \DM_rd1[8]_pad  & n7022 ;
  assign n10429 = \DM_rd3[8]_pad  & n7038 ;
  assign n10433 = ~n10425 & ~n10429 ;
  assign n10434 = ~n10432 & n10433 ;
  assign n10438 = ~n10426 & n10434 ;
  assign n10439 = ~n10431 & n10438 ;
  assign n10440 = n10437 & n10439 ;
  assign n10441 = ~n10430 & n10440 ;
  assign n10442 = \regout_STD_C_reg[8]/P0001  & n6988 ;
  assign n10583 = \bdma_BCTL_reg[8]/NET0131  & n7230 ;
  assign n10581 = \tm_tpr_reg_DO_reg[8]/NET0131  & n7293 ;
  assign n10603 = ~n7522 & ~n10581 ;
  assign n10582 = \sport1_regs_FSDIVreg_DO_reg[8]/NET0131  & n7273 ;
  assign n10584 = \idma_DCTL_reg[8]/NET0131  & n7299 ;
  assign n10604 = ~n10582 & ~n10584 ;
  assign n10614 = n10603 & n10604 ;
  assign n10598 = \sport1_txctl_Wcnt_reg[0]/NET0131  & n7689 ;
  assign n10599 = \sport0_txctl_Wcnt_reg[0]/NET0131  & n7710 ;
  assign n10615 = ~n10598 & ~n10599 ;
  assign n10616 = n10614 & n10615 ;
  assign n10619 = ~n10583 & n10616 ;
  assign n10585 = \bdma_BIAD_reg[8]/NET0131  & n7234 ;
  assign n10588 = \bdma_BEAD_reg[8]/NET0131  & n7303 ;
  assign n10620 = ~n10585 & ~n10588 ;
  assign n10621 = n10619 & n10620 ;
  assign n10597 = \bdma_BWCOUNT_reg[8]/NET0131  & n7287 ;
  assign n10586 = \bdma_BOVL_reg[8]/NET0131  & n7534 ;
  assign n10596 = \IRFS1_pad  & n7281 ;
  assign n10600 = \memc_usysr_DO_reg[8]/NET0131  & n7301 ;
  assign n10609 = ~n10596 & ~n10600 ;
  assign n10601 = \clkc_ckr_reg_DO_reg[8]/NET0131  & n7239 ;
  assign n10602 = \sport0_regs_FSDIVreg_DO_reg[8]/NET0131  & n7259 ;
  assign n10610 = ~n10601 & ~n10602 ;
  assign n10611 = n10609 & n10610 ;
  assign n10592 = \sport0_regs_AUTOreg_DO_reg[8]/NET0131  & n7295 ;
  assign n10593 = \emc_WSCRreg_DO_reg[8]/NET0131  & n7251 ;
  assign n10607 = ~n10592 & ~n10593 ;
  assign n10594 = \sport1_regs_SCLKDIVreg_DO_reg[8]/NET0131  & n7247 ;
  assign n10595 = \sport1_regs_AUTOreg_DO_reg[8]/NET0131  & n7527 ;
  assign n10608 = ~n10594 & ~n10595 ;
  assign n10612 = n10607 & n10608 ;
  assign n10587 = \idma_DOVL_reg[8]/NET0131  & n7532 ;
  assign n10589 = \IRFS0_pad  & n7249 ;
  assign n10605 = ~n10587 & ~n10589 ;
  assign n10590 = \sport0_regs_SCLKDIVreg_DO_reg[8]/NET0131  & n7256 ;
  assign n10591 = \tm_TCR_TMP_reg[8]/NET0131  & n7289 ;
  assign n10606 = ~n10590 & ~n10591 ;
  assign n10613 = n10605 & n10606 ;
  assign n10617 = n10612 & n10613 ;
  assign n10618 = n10611 & n10617 ;
  assign n10622 = ~n10586 & n10618 ;
  assign n10623 = ~n10597 & n10622 ;
  assign n10624 = n10621 & n10623 ;
  assign n10625 = \memc_ldSREG_E_reg/NET0131  & ~n10624 ;
  assign n10556 = \core_c_dec_MFtoppcs_Eg_reg/P0001  & ~n4425 ;
  assign n10558 = \core_c_dec_IRE_reg[12]/NET0131  & ~n7216 ;
  assign n10559 = \core_c_dec_MFIMASK_E_reg/P0001  & \core_c_psq_IMASK_reg[8]/NET0131  ;
  assign n10555 = \core_c_dec_MFCNTR_E_reg/P0001  & \core_c_psq_CNTR_reg_DO_reg[8]/NET0131  ;
  assign n10557 = \core_c_dec_MFIDR_E_reg/P0001  & \sice_idr0_reg_DO_reg[8]/P0001  ;
  assign n10560 = ~n10555 & ~n10557 ;
  assign n10561 = ~n10559 & n10560 ;
  assign n10562 = ~n10558 & n10561 ;
  assign n10563 = ~n10556 & n10562 ;
  assign n10564 = n7215 & ~n10563 ;
  assign n10500 = \core_c_dec_MFMreg_E_reg[1]/P0001  & \core_dag_ilm1reg_M1_we_DO_reg[8]/NET0131  ;
  assign n10501 = \core_c_dec_MFIreg_E_reg[2]/P0001  & \core_dag_ilm1reg_I2_we_DO_reg[8]/NET0131  ;
  assign n10508 = ~n10500 & ~n10501 ;
  assign n10502 = \core_c_dec_MFIreg_E_reg[1]/P0001  & \core_dag_ilm1reg_I1_we_DO_reg[8]/NET0131  ;
  assign n10503 = \core_c_dec_MFLreg_E_reg[1]/P0001  & \core_dag_ilm1reg_L1_we_DO_reg[8]/NET0131  ;
  assign n10509 = ~n10502 & ~n10503 ;
  assign n10510 = n10508 & n10509 ;
  assign n10496 = \core_c_dec_MFIreg_E_reg[3]/P0001  & \core_dag_ilm1reg_I3_we_DO_reg[8]/NET0131  ;
  assign n10497 = \core_c_dec_MFLreg_E_reg[0]/P0001  & \core_dag_ilm1reg_L0_we_DO_reg[8]/NET0131  ;
  assign n10506 = ~n10496 & ~n10497 ;
  assign n10498 = \core_c_dec_MFMreg_E_reg[3]/P0001  & \core_dag_ilm1reg_M3_we_DO_reg[8]/NET0131  ;
  assign n10499 = \core_c_dec_MFMreg_E_reg[2]/P0001  & \core_dag_ilm1reg_M2_we_DO_reg[8]/NET0131  ;
  assign n10507 = ~n10498 & ~n10499 ;
  assign n10511 = n10506 & n10507 ;
  assign n10492 = \core_c_dec_MFLreg_E_reg[2]/P0001  & \core_dag_ilm1reg_L2_we_DO_reg[8]/NET0131  ;
  assign n10493 = \core_c_dec_MFMreg_E_reg[0]/P0001  & \core_dag_ilm1reg_M0_we_DO_reg[8]/NET0131  ;
  assign n10504 = ~n10492 & ~n10493 ;
  assign n10494 = \core_c_dec_MFLreg_E_reg[3]/P0001  & \core_dag_ilm1reg_L3_we_DO_reg[8]/NET0131  ;
  assign n10495 = \core_c_dec_MFIreg_E_reg[0]/P0001  & \core_dag_ilm1reg_I0_we_DO_reg[8]/NET0131  ;
  assign n10505 = ~n10494 & ~n10495 ;
  assign n10512 = n10504 & n10505 ;
  assign n10513 = n10511 & n10512 ;
  assign n10514 = n10510 & n10513 ;
  assign n10515 = n7068 & ~n10514 ;
  assign n10476 = \core_c_dec_MFLreg_E_reg[6]/P0001  & \core_dag_ilm2reg_L6_we_DO_reg[8]/NET0131  ;
  assign n10477 = \core_c_dec_MFMreg_E_reg[5]/P0001  & \core_dag_ilm2reg_M5_we_DO_reg[8]/NET0131  ;
  assign n10484 = ~n10476 & ~n10477 ;
  assign n10478 = \core_c_dec_MFMreg_E_reg[6]/P0001  & \core_dag_ilm2reg_M6_we_DO_reg[8]/NET0131  ;
  assign n10479 = \core_c_dec_MFMreg_E_reg[7]/P0001  & \core_dag_ilm2reg_M7_we_DO_reg[8]/NET0131  ;
  assign n10485 = ~n10478 & ~n10479 ;
  assign n10486 = n10484 & n10485 ;
  assign n10472 = \core_c_dec_MFLreg_E_reg[7]/P0001  & \core_dag_ilm2reg_L7_we_DO_reg[8]/NET0131  ;
  assign n10473 = \core_c_dec_MFLreg_E_reg[4]/P0001  & \core_dag_ilm2reg_L4_we_DO_reg[8]/NET0131  ;
  assign n10482 = ~n10472 & ~n10473 ;
  assign n10474 = \core_c_dec_MFMreg_E_reg[4]/P0001  & \core_dag_ilm2reg_M4_we_DO_reg[8]/NET0131  ;
  assign n10475 = \core_c_dec_MFIreg_E_reg[4]/P0001  & \core_dag_ilm2reg_I4_we_DO_reg[8]/NET0131  ;
  assign n10483 = ~n10474 & ~n10475 ;
  assign n10487 = n10482 & n10483 ;
  assign n10468 = \core_c_dec_MFIreg_E_reg[6]/P0001  & \core_dag_ilm2reg_I6_we_DO_reg[8]/NET0131  ;
  assign n10469 = \core_c_dec_MFLreg_E_reg[5]/P0001  & \core_dag_ilm2reg_L5_we_DO_reg[8]/NET0131  ;
  assign n10480 = ~n10468 & ~n10469 ;
  assign n10470 = \core_c_dec_MFIreg_E_reg[5]/P0001  & \core_dag_ilm2reg_I5_we_DO_reg[8]/NET0131  ;
  assign n10471 = \core_c_dec_MFIreg_E_reg[7]/P0001  & \core_dag_ilm2reg_I7_we_DO_reg[8]/NET0131  ;
  assign n10481 = ~n10470 & ~n10471 ;
  assign n10488 = n10480 & n10481 ;
  assign n10489 = n10487 & n10488 ;
  assign n10490 = n10486 & n10489 ;
  assign n10491 = n7128 & ~n10490 ;
  assign n10547 = \core_c_dec_MFTX1_E_reg/P0001  & \sport1_txctl_TX_reg[8]/P0001  ;
  assign n10548 = \core_c_dec_MFTX0_E_reg/P0001  & \sport0_txctl_TX_reg[8]/P0001  ;
  assign n10551 = ~n10547 & ~n10548 ;
  assign n10549 = \core_c_dec_MFRX1_E_reg/P0001  & \sport1_rxctl_RX_reg[8]/P0001  ;
  assign n10550 = \core_c_dec_MFRX0_E_reg/P0001  & \sport0_rxctl_RX_reg[8]/P0001  ;
  assign n10552 = ~n10549 & ~n10550 ;
  assign n10553 = n10551 & n10552 ;
  assign n10554 = n7119 & ~n10553 ;
  assign n10626 = ~n10491 & ~n10554 ;
  assign n10627 = ~n10515 & n10626 ;
  assign n10573 = ~\core_c_psq_MSTAT_reg_DO_reg[0]/P0002  & \core_eu_es_sht_es_reg_sr1rwe_DO_reg[8]/P0001  ;
  assign n10574 = \core_c_psq_MSTAT_reg_DO_reg[0]/P0002  & \core_eu_es_sht_es_reg_sr1swe_DO_reg[8]/P0001  ;
  assign n10575 = ~n10573 & ~n10574 ;
  assign n10576 = \core_c_dec_MFSR1_E_reg/P0001  & ~n10575 ;
  assign n10565 = ~\core_c_psq_MSTAT_reg_DO_reg[0]/P0002  & \core_eu_es_sht_es_reg_sr0rwe_DO_reg[8]/P0001  ;
  assign n10566 = \core_c_psq_MSTAT_reg_DO_reg[0]/P0002  & \core_eu_es_sht_es_reg_sr0swe_DO_reg[8]/P0001  ;
  assign n10567 = ~n10565 & ~n10566 ;
  assign n10568 = \core_c_dec_MFSR0_E_reg/P0001  & ~n10567 ;
  assign n10569 = ~\core_c_psq_MSTAT_reg_DO_reg[0]/P0002  & \core_eu_es_sht_es_reg_sirwe_DO_reg[8]/P0001  ;
  assign n10570 = \core_c_psq_MSTAT_reg_DO_reg[0]/P0002  & \core_eu_es_sht_es_reg_siswe_DO_reg[8]/P0001  ;
  assign n10571 = ~n10569 & ~n10570 ;
  assign n10572 = \core_c_dec_MFSI_E_reg/P0001  & ~n10571 ;
  assign n10577 = ~n10568 & ~n10572 ;
  assign n10578 = ~n10576 & n10577 ;
  assign n10579 = n7174 & n10578 ;
  assign n10580 = n7153 & ~n10579 ;
  assign n10443 = ~\core_c_psq_MSTAT_reg_DO_reg[0]/P0002  & \core_eu_ea_alu_ea_reg_ay1rwe_DO_reg[8]/P0001  ;
  assign n10444 = \core_c_psq_MSTAT_reg_DO_reg[0]/P0002  & \core_eu_ea_alu_ea_reg_ay1swe_DO_reg[8]/P0001  ;
  assign n10445 = ~n10443 & ~n10444 ;
  assign n10446 = \core_c_dec_MFAY1_E_reg/P0001  & ~n10445 ;
  assign n10447 = ~\core_c_psq_MSTAT_reg_DO_reg[0]/P0002  & \core_eu_ea_alu_ea_reg_ax0rwe_DO_reg[8]/P0001  ;
  assign n10448 = \core_c_psq_MSTAT_reg_DO_reg[0]/P0002  & \core_eu_ea_alu_ea_reg_ax0swe_DO_reg[8]/P0001  ;
  assign n10449 = ~n10447 & ~n10448 ;
  assign n10450 = \core_c_dec_MFAX0_E_reg/P0001  & ~n10449 ;
  assign n10463 = ~n10446 & ~n10450 ;
  assign n10459 = ~\core_c_psq_MSTAT_reg_DO_reg[0]/P0002  & \core_eu_ea_alu_ea_reg_arrwe_DO_reg[8]/P0001  ;
  assign n10460 = \core_c_psq_MSTAT_reg_DO_reg[0]/P0002  & \core_eu_ea_alu_ea_reg_arswe_DO_reg[8]/P0001  ;
  assign n10461 = ~n10459 & ~n10460 ;
  assign n10462 = \core_c_dec_MFAR_E_reg/P0001  & ~n10461 ;
  assign n10451 = ~\core_c_psq_MSTAT_reg_DO_reg[0]/P0002  & \core_eu_ea_alu_ea_reg_ay0rwe_DO_reg[8]/P0001  ;
  assign n10452 = \core_c_psq_MSTAT_reg_DO_reg[0]/P0002  & \core_eu_ea_alu_ea_reg_ay0swe_DO_reg[8]/P0001  ;
  assign n10453 = ~n10451 & ~n10452 ;
  assign n10454 = \core_c_dec_MFAY0_E_reg/P0001  & ~n10453 ;
  assign n10455 = ~\core_c_psq_MSTAT_reg_DO_reg[0]/P0002  & \core_eu_ea_alu_ea_reg_ax1rwe_DO_reg[8]/P0001  ;
  assign n10456 = \core_c_psq_MSTAT_reg_DO_reg[0]/P0002  & \core_eu_ea_alu_ea_reg_ax1swe_DO_reg[8]/P0001  ;
  assign n10457 = ~n10455 & ~n10456 ;
  assign n10458 = \core_c_dec_MFAX1_E_reg/P0001  & ~n10457 ;
  assign n10464 = ~n10454 & ~n10458 ;
  assign n10465 = ~n10462 & n10464 ;
  assign n10466 = n10463 & n10465 ;
  assign n10467 = n7093 & ~n10466 ;
  assign n10536 = ~\core_c_psq_MSTAT_reg_DO_reg[0]/P0002  & \core_eu_em_mac_em_reg_mr1rwe_DO_reg[8]/P0001  ;
  assign n10537 = \core_c_psq_MSTAT_reg_DO_reg[0]/P0002  & \core_eu_em_mac_em_reg_mr1swe_DO_reg[8]/P0001  ;
  assign n10538 = ~n10536 & ~n10537 ;
  assign n10539 = \core_c_dec_MFMR1_E_reg/P0001  & ~n10538 ;
  assign n10528 = ~\core_c_psq_MSTAT_reg_DO_reg[0]/P0002  & \core_eu_em_mac_em_reg_mx1rwe_DO_reg[8]/P0001  ;
  assign n10529 = \core_c_psq_MSTAT_reg_DO_reg[0]/P0002  & \core_eu_em_mac_em_reg_mx1swe_DO_reg[8]/P0001  ;
  assign n10530 = ~n10528 & ~n10529 ;
  assign n10531 = \core_c_dec_MFMX1_E_reg/P0001  & ~n10530 ;
  assign n10532 = ~\core_c_psq_MSTAT_reg_DO_reg[0]/P0002  & \core_eu_em_mac_em_reg_mr0rwe_DO_reg[8]/P0001  ;
  assign n10533 = \core_c_psq_MSTAT_reg_DO_reg[0]/P0002  & \core_eu_em_mac_em_reg_mr0swe_DO_reg[8]/P0001  ;
  assign n10534 = ~n10532 & ~n10533 ;
  assign n10535 = \core_c_dec_MFMR0_E_reg/P0001  & ~n10534 ;
  assign n10542 = ~n10531 & ~n10535 ;
  assign n10543 = ~n10539 & n10542 ;
  assign n10516 = ~\core_c_psq_MSTAT_reg_DO_reg[0]/P0002  & \core_eu_em_mac_em_reg_my0rwe_DO_reg[8]/P0001  ;
  assign n10517 = \core_c_psq_MSTAT_reg_DO_reg[0]/P0002  & \core_eu_em_mac_em_reg_my0swe_DO_reg[8]/P0001  ;
  assign n10518 = ~n10516 & ~n10517 ;
  assign n10519 = \core_c_dec_MFMY0_E_reg/P0001  & ~n10518 ;
  assign n10540 = ~n7207 & ~n10519 ;
  assign n10520 = ~\core_c_psq_MSTAT_reg_DO_reg[0]/P0002  & \core_eu_em_mac_em_reg_my1rwe_DO_reg[8]/P0001  ;
  assign n10521 = \core_c_psq_MSTAT_reg_DO_reg[0]/P0002  & \core_eu_em_mac_em_reg_my1swe_DO_reg[8]/P0001  ;
  assign n10522 = ~n10520 & ~n10521 ;
  assign n10523 = \core_c_dec_MFMY1_E_reg/P0001  & ~n10522 ;
  assign n10524 = ~\core_c_psq_MSTAT_reg_DO_reg[0]/P0002  & \core_eu_em_mac_em_reg_mx0rwe_DO_reg[8]/P0001  ;
  assign n10525 = \core_c_psq_MSTAT_reg_DO_reg[0]/P0002  & \core_eu_em_mac_em_reg_mx0swe_DO_reg[8]/P0001  ;
  assign n10526 = ~n10524 & ~n10525 ;
  assign n10527 = \core_c_dec_MFMX0_E_reg/P0001  & ~n10526 ;
  assign n10541 = ~n10523 & ~n10527 ;
  assign n10544 = n10540 & n10541 ;
  assign n10545 = n10543 & n10544 ;
  assign n10546 = n7179 & ~n10545 ;
  assign n10628 = ~n10467 & ~n10546 ;
  assign n10629 = ~n10580 & n10628 ;
  assign n10630 = n10627 & n10629 ;
  assign n10631 = ~n10564 & n10630 ;
  assign n10632 = ~n10625 & n10631 ;
  assign n10633 = ~n10442 & n10632 ;
  assign n10634 = ~\emc_DMDoe_reg/NET0131  & ~n10633 ;
  assign n10635 = \emc_DMDoe_reg/NET0131  & \emc_DMDreg_reg[8]/P0001  ;
  assign n10636 = n7057 & ~n10635 ;
  assign n10637 = ~n10634 & n10636 ;
  assign n10638 = ~n10441 & ~n10637 ;
  assign n10639 = n7863 & n10638 ;
  assign n10640 = ~n10423 & ~n10639 ;
  assign n10641 = n7005 & ~n10640 ;
  assign n10650 = ~n6282 & ~n6505 ;
  assign n10651 = ~n6283 & ~n10650 ;
  assign n10652 = ~n6289 & n10651 ;
  assign n10653 = n6289 & ~n10651 ;
  assign n10654 = ~n10652 & ~n10653 ;
  assign n10659 = ~n6496 & n10654 ;
  assign n10643 = ~n6293 & ~n6377 ;
  assign n10644 = ~n6308 & ~n6372 ;
  assign n10645 = ~n6378 & ~n10644 ;
  assign n10646 = n10643 & n10645 ;
  assign n10647 = ~n10643 & ~n10645 ;
  assign n10648 = ~n10646 & ~n10647 ;
  assign n10658 = n6496 & n10648 ;
  assign n10660 = ~\core_dag_ilm1reg_M_reg[13]/NET0131  & ~n10658 ;
  assign n10661 = ~n10659 & n10660 ;
  assign n10642 = \core_dag_ilm1reg_I_reg[5]/NET0131  & ~n6251 ;
  assign n10655 = n7612 & n10654 ;
  assign n10649 = ~n7612 & n10648 ;
  assign n10656 = \core_dag_ilm1reg_M_reg[13]/NET0131  & ~n10649 ;
  assign n10657 = ~n10655 & n10656 ;
  assign n10662 = ~n10642 & ~n10657 ;
  assign n10663 = ~n10661 & n10662 ;
  assign n10664 = ~n6135 & n10663 ;
  assign n10671 = \DM_rd0[5]_pad  & ~n7053 ;
  assign n10665 = \DM_rdm[5]_pad  & n7016 ;
  assign n10676 = ~n7057 & ~n10665 ;
  assign n10668 = \DM_rd6[5]_pad  & n7031 ;
  assign n10669 = \DM_rd7[5]_pad  & n7034 ;
  assign n10677 = ~n10668 & ~n10669 ;
  assign n10678 = n10676 & n10677 ;
  assign n10672 = \DM_rd5[5]_pad  & n7043 ;
  assign n10667 = \DM_rd4[5]_pad  & n7028 ;
  assign n10673 = \DM_rd2[5]_pad  & n7041 ;
  assign n10666 = \DM_rd1[5]_pad  & n7022 ;
  assign n10670 = \DM_rd3[5]_pad  & n7038 ;
  assign n10674 = ~n10666 & ~n10670 ;
  assign n10675 = ~n10673 & n10674 ;
  assign n10679 = ~n10667 & n10675 ;
  assign n10680 = ~n10672 & n10679 ;
  assign n10681 = n10678 & n10680 ;
  assign n10682 = ~n10671 & n10681 ;
  assign n10683 = \regout_STD_C_reg[5]/P0001  & n6988 ;
  assign n10727 = \bdma_BIAD_reg[5]/NET0131  & n7234 ;
  assign n10718 = \emc_WSCRreg_DO_reg[5]/NET0131  & n7251 ;
  assign n10719 = \sport0_regs_SCLKDIVreg_DO_reg[5]/NET0131  & n7256 ;
  assign n10744 = ~n10718 & ~n10719 ;
  assign n10720 = \sport1_regs_MWORDreg_DO_reg[5]/NET0131  & n7263 ;
  assign n10721 = \tm_tsr_reg_DO_reg[5]/NET0131  & n7540 ;
  assign n10745 = ~n10720 & ~n10721 ;
  assign n10758 = n10744 & n10745 ;
  assign n10711 = \idma_DOVL_reg[5]/NET0131  & n7532 ;
  assign n10742 = ~n7522 & ~n10711 ;
  assign n10712 = \sport0_regs_AUTOreg_DO_reg[5]/NET0131  & n7295 ;
  assign n10713 = \tm_tpr_reg_DO_reg[5]/NET0131  & n7293 ;
  assign n10743 = ~n10712 & ~n10713 ;
  assign n10759 = n10742 & n10743 ;
  assign n10760 = n10758 & n10759 ;
  assign n10764 = ~n10727 & n10760 ;
  assign n10735 = \bdma_BEAD_reg[5]/NET0131  & n7303 ;
  assign n10736 = \bdma_BCTL_reg[5]/NET0131  & n7230 ;
  assign n10765 = ~n10735 & ~n10736 ;
  assign n10766 = n10764 & n10765 ;
  assign n10732 = \bdma_BOVL_reg[5]/NET0131  & n7534 ;
  assign n10714 = ~\bdma_BDMA_boot_reg/NET0131_reg_syn_10  & \bdma_BWCOUNT_reg[5]/NET0131_reg_syn_2  ;
  assign n10715 = \bdma_BDMA_boot_reg/NET0131_reg_syn_10  & \bdma_BWCOUNT_reg[5]/NET0131_reg_syn_8  ;
  assign n10716 = ~n10714 & ~n10715 ;
  assign n10717 = n7287 & ~n10716 ;
  assign n10726 = \pio_pmask_reg_DO_reg[5]/NET0131  & n7297 ;
  assign n10728 = \sport0_regs_MWORDreg_DO_reg[5]/NET0131  & n7276 ;
  assign n10748 = ~n10726 & ~n10728 ;
  assign n10729 = \sport1_regs_AUTOreg_DO_reg[5]/NET0131  & n7527 ;
  assign n10730 = \tm_TCR_TMP_reg[5]/NET0131  & n7289 ;
  assign n10749 = ~n10729 & ~n10730 ;
  assign n10756 = n10748 & n10749 ;
  assign n10722 = \sport0_regs_SCTLreg_DO_reg[5]/NET0131  & n7249 ;
  assign n10723 = \emc_WSCRext_reg_DO_reg[5]/NET0131  & n7514 ;
  assign n10746 = ~n10722 & ~n10723 ;
  assign n10724 = \sport1_regs_SCLKDIVreg_DO_reg[5]/NET0131  & n7247 ;
  assign n10725 = \sport1_regs_SCTLreg_DO_reg[5]/NET0131  & n7281 ;
  assign n10747 = ~n10724 & ~n10725 ;
  assign n10757 = n10746 & n10747 ;
  assign n10761 = n10756 & n10757 ;
  assign n10738 = \idma_DCTL_reg[5]/NET0131  & n7299 ;
  assign n10739 = \PIO_out[5]_pad  & n7291 ;
  assign n10752 = ~n10738 & ~n10739 ;
  assign n10740 = \PIO_oe[5]_pad  & n7244 ;
  assign n10741 = \sport1_regs_FSDIVreg_DO_reg[5]/NET0131  & n7273 ;
  assign n10753 = ~n10740 & ~n10741 ;
  assign n10754 = n10752 & n10753 ;
  assign n10731 = \sport0_regs_FSDIVreg_DO_reg[5]/NET0131  & n7259 ;
  assign n10733 = \clkc_ckr_reg_DO_reg[5]/NET0131  & n7239 ;
  assign n10750 = ~n10731 & ~n10733 ;
  assign n10734 = \memc_usysr_DO_reg[5]/NET0131  & n7301 ;
  assign n10737 = \pio_PINT_reg[5]/NET0131  & n7271 ;
  assign n10751 = ~n10734 & ~n10737 ;
  assign n10755 = n10750 & n10751 ;
  assign n10762 = n10754 & n10755 ;
  assign n10763 = n10761 & n10762 ;
  assign n10767 = ~n10717 & n10763 ;
  assign n10768 = ~n10732 & n10767 ;
  assign n10769 = n10766 & n10768 ;
  assign n10770 = \memc_ldSREG_E_reg/NET0131  & ~n10769 ;
  assign n10772 = \core_c_dec_MFtoppcs_Eg_reg/P0001  & ~n4244 ;
  assign n10775 = \core_c_dec_MFIMASK_E_reg/P0001  & \core_c_psq_IMASK_reg[5]/NET0131  ;
  assign n10776 = \core_c_dec_MFMSTAT_E_reg/P0001  & \core_c_psq_MSTAT_reg_DO_reg[5]/NET0131  ;
  assign n10780 = ~n10775 & ~n10776 ;
  assign n10777 = \core_c_dec_MFSSTAT_E_reg/P0001  & \core_c_psq_SSTAT_reg[5]/NET0131  ;
  assign n10778 = \core_c_dec_MFIDR_E_reg/P0001  & \sice_idr0_reg_DO_reg[5]/P0001  ;
  assign n10781 = ~n10777 & ~n10778 ;
  assign n10782 = n10780 & n10781 ;
  assign n10773 = \core_c_dec_IRE_reg[9]/NET0131  & ~n7216 ;
  assign n10771 = \core_c_dec_MFPMOVL_E_reg/P0001  & \core_c_psq_PMOVL_regh_DO_reg[1]/NET0131  ;
  assign n10774 = \core_c_dec_MFCNTR_E_reg/P0001  & \core_c_psq_CNTR_reg_DO_reg[5]/NET0131  ;
  assign n10779 = ~n10771 & ~n10774 ;
  assign n10783 = ~n10773 & n10779 ;
  assign n10784 = n10782 & n10783 ;
  assign n10785 = ~n10772 & n10784 ;
  assign n10786 = n7215 & ~n10785 ;
  assign n10840 = \core_c_dec_MFIreg_E_reg[4]/P0001  & \core_dag_ilm2reg_I4_we_DO_reg[5]/NET0131  ;
  assign n10841 = \core_c_dec_MFMreg_E_reg[4]/P0001  & \core_dag_ilm2reg_M4_we_DO_reg[5]/NET0131  ;
  assign n10848 = ~n10840 & ~n10841 ;
  assign n10842 = \core_c_dec_MFLreg_E_reg[7]/P0001  & \core_dag_ilm2reg_L7_we_DO_reg[5]/NET0131  ;
  assign n10843 = \core_c_dec_MFMreg_E_reg[7]/P0001  & \core_dag_ilm2reg_M7_we_DO_reg[5]/NET0131  ;
  assign n10849 = ~n10842 & ~n10843 ;
  assign n10850 = n10848 & n10849 ;
  assign n10836 = \core_c_dec_MFMreg_E_reg[5]/P0001  & \core_dag_ilm2reg_M5_we_DO_reg[5]/NET0131  ;
  assign n10837 = \core_c_dec_MFMreg_E_reg[6]/P0001  & \core_dag_ilm2reg_M6_we_DO_reg[5]/NET0131  ;
  assign n10846 = ~n10836 & ~n10837 ;
  assign n10838 = \core_c_dec_MFIreg_E_reg[6]/P0001  & \core_dag_ilm2reg_I6_we_DO_reg[5]/NET0131  ;
  assign n10839 = \core_c_dec_MFIreg_E_reg[5]/P0001  & \core_dag_ilm2reg_I5_we_DO_reg[5]/NET0131  ;
  assign n10847 = ~n10838 & ~n10839 ;
  assign n10851 = n10846 & n10847 ;
  assign n10832 = \core_c_dec_MFIreg_E_reg[7]/P0001  & \core_dag_ilm2reg_I7_we_DO_reg[5]/NET0131  ;
  assign n10833 = \core_c_dec_MFLreg_E_reg[5]/P0001  & \core_dag_ilm2reg_L5_we_DO_reg[5]/NET0131  ;
  assign n10844 = ~n10832 & ~n10833 ;
  assign n10834 = \core_c_dec_MFLreg_E_reg[4]/P0001  & \core_dag_ilm2reg_L4_we_DO_reg[5]/NET0131  ;
  assign n10835 = \core_c_dec_MFLreg_E_reg[6]/P0001  & \core_dag_ilm2reg_L6_we_DO_reg[5]/NET0131  ;
  assign n10845 = ~n10834 & ~n10835 ;
  assign n10852 = n10844 & n10845 ;
  assign n10853 = n10851 & n10852 ;
  assign n10854 = n10850 & n10853 ;
  assign n10855 = n7128 & ~n10854 ;
  assign n10816 = \core_c_dec_MFIreg_E_reg[3]/P0001  & \core_dag_ilm1reg_I3_we_DO_reg[5]/NET0131  ;
  assign n10817 = \core_c_dec_MFIreg_E_reg[0]/P0001  & \core_dag_ilm1reg_I0_we_DO_reg[5]/NET0131  ;
  assign n10824 = ~n10816 & ~n10817 ;
  assign n10818 = \core_c_dec_MFIreg_E_reg[1]/P0001  & \core_dag_ilm1reg_I1_we_DO_reg[5]/NET0131  ;
  assign n10819 = \core_c_dec_MFIreg_E_reg[2]/P0001  & \core_dag_ilm1reg_I2_we_DO_reg[5]/NET0131  ;
  assign n10825 = ~n10818 & ~n10819 ;
  assign n10826 = n10824 & n10825 ;
  assign n10812 = \core_c_dec_MFLreg_E_reg[0]/P0001  & \core_dag_ilm1reg_L0_we_DO_reg[5]/NET0131  ;
  assign n10813 = \core_c_dec_MFMreg_E_reg[2]/P0001  & \core_dag_ilm1reg_M2_we_DO_reg[5]/NET0131  ;
  assign n10822 = ~n10812 & ~n10813 ;
  assign n10814 = \core_c_dec_MFLreg_E_reg[1]/P0001  & \core_dag_ilm1reg_L1_we_DO_reg[5]/NET0131  ;
  assign n10815 = \core_c_dec_MFLreg_E_reg[2]/P0001  & \core_dag_ilm1reg_L2_we_DO_reg[5]/NET0131  ;
  assign n10823 = ~n10814 & ~n10815 ;
  assign n10827 = n10822 & n10823 ;
  assign n10808 = \core_c_dec_MFMreg_E_reg[0]/P0001  & \core_dag_ilm1reg_M0_we_DO_reg[5]/NET0131  ;
  assign n10809 = \core_c_dec_MFMreg_E_reg[3]/P0001  & \core_dag_ilm1reg_M3_we_DO_reg[5]/NET0131  ;
  assign n10820 = ~n10808 & ~n10809 ;
  assign n10810 = \core_c_dec_MFLreg_E_reg[3]/P0001  & \core_dag_ilm1reg_L3_we_DO_reg[5]/NET0131  ;
  assign n10811 = \core_c_dec_MFMreg_E_reg[1]/P0001  & \core_dag_ilm1reg_M1_we_DO_reg[5]/NET0131  ;
  assign n10821 = ~n10810 & ~n10811 ;
  assign n10828 = n10820 & n10821 ;
  assign n10829 = n10827 & n10828 ;
  assign n10830 = n10826 & n10829 ;
  assign n10831 = n7068 & ~n10830 ;
  assign n10891 = \core_c_dec_MFTX1_E_reg/P0001  & \sport1_txctl_TX_reg[5]/P0001  ;
  assign n10892 = \core_c_dec_MFTX0_E_reg/P0001  & \sport0_txctl_TX_reg[5]/P0001  ;
  assign n10895 = ~n10891 & ~n10892 ;
  assign n10893 = \core_c_dec_MFRX1_E_reg/P0001  & \sport1_rxctl_RX_reg[5]/P0001  ;
  assign n10894 = \core_c_dec_MFRX0_E_reg/P0001  & \sport0_rxctl_RX_reg[5]/P0001  ;
  assign n10896 = ~n10893 & ~n10894 ;
  assign n10897 = n10895 & n10896 ;
  assign n10898 = n7119 & ~n10897 ;
  assign n10899 = ~n10831 & ~n10898 ;
  assign n10900 = ~n10855 & n10899 ;
  assign n10880 = ~\core_c_psq_MSTAT_reg_DO_reg[0]/P0002  & \core_eu_em_mac_em_reg_mr2rwe_DO_reg[5]/P0001  ;
  assign n10881 = \core_c_psq_MSTAT_reg_DO_reg[0]/P0002  & \core_eu_em_mac_em_reg_mr2swe_DO_reg[5]/P0001  ;
  assign n10882 = ~n10880 & ~n10881 ;
  assign n10883 = \core_c_dec_MFMR2_E_reg/P0001  & ~n10882 ;
  assign n10872 = ~\core_c_psq_MSTAT_reg_DO_reg[0]/P0002  & \core_eu_em_mac_em_reg_mx0rwe_DO_reg[5]/P0001  ;
  assign n10873 = \core_c_psq_MSTAT_reg_DO_reg[0]/P0002  & \core_eu_em_mac_em_reg_mx0swe_DO_reg[5]/P0001  ;
  assign n10874 = ~n10872 & ~n10873 ;
  assign n10875 = \core_c_dec_MFMX0_E_reg/P0001  & ~n10874 ;
  assign n10876 = ~\core_c_psq_MSTAT_reg_DO_reg[0]/P0002  & \core_eu_em_mac_em_reg_mr0rwe_DO_reg[5]/P0001  ;
  assign n10877 = \core_c_psq_MSTAT_reg_DO_reg[0]/P0002  & \core_eu_em_mac_em_reg_mr0swe_DO_reg[5]/P0001  ;
  assign n10878 = ~n10876 & ~n10877 ;
  assign n10879 = \core_c_dec_MFMR0_E_reg/P0001  & ~n10878 ;
  assign n10886 = ~n10875 & ~n10879 ;
  assign n10887 = ~n10883 & n10886 ;
  assign n10856 = ~\core_c_psq_MSTAT_reg_DO_reg[0]/P0002  & \core_eu_em_mac_em_reg_mr1rwe_DO_reg[5]/P0001  ;
  assign n10857 = \core_c_psq_MSTAT_reg_DO_reg[0]/P0002  & \core_eu_em_mac_em_reg_mr1swe_DO_reg[5]/P0001  ;
  assign n10858 = ~n10856 & ~n10857 ;
  assign n10859 = \core_c_dec_MFMR1_E_reg/P0001  & ~n10858 ;
  assign n10860 = ~\core_c_psq_MSTAT_reg_DO_reg[0]/P0002  & \core_eu_em_mac_em_reg_my0rwe_DO_reg[5]/P0001  ;
  assign n10861 = \core_c_psq_MSTAT_reg_DO_reg[0]/P0002  & \core_eu_em_mac_em_reg_my0swe_DO_reg[5]/P0001  ;
  assign n10862 = ~n10860 & ~n10861 ;
  assign n10863 = \core_c_dec_MFMY0_E_reg/P0001  & ~n10862 ;
  assign n10884 = ~n10859 & ~n10863 ;
  assign n10864 = ~\core_c_psq_MSTAT_reg_DO_reg[0]/P0002  & \core_eu_em_mac_em_reg_mx1rwe_DO_reg[5]/P0001  ;
  assign n10865 = \core_c_psq_MSTAT_reg_DO_reg[0]/P0002  & \core_eu_em_mac_em_reg_mx1swe_DO_reg[5]/P0001  ;
  assign n10866 = ~n10864 & ~n10865 ;
  assign n10867 = \core_c_dec_MFMX1_E_reg/P0001  & ~n10866 ;
  assign n10868 = ~\core_c_psq_MSTAT_reg_DO_reg[0]/P0002  & \core_eu_em_mac_em_reg_my1rwe_DO_reg[5]/P0001  ;
  assign n10869 = \core_c_psq_MSTAT_reg_DO_reg[0]/P0002  & \core_eu_em_mac_em_reg_my1swe_DO_reg[5]/P0001  ;
  assign n10870 = ~n10868 & ~n10869 ;
  assign n10871 = \core_c_dec_MFMY1_E_reg/P0001  & ~n10870 ;
  assign n10885 = ~n10867 & ~n10871 ;
  assign n10888 = n10884 & n10885 ;
  assign n10889 = n10887 & n10888 ;
  assign n10890 = n7179 & ~n10889 ;
  assign n10684 = ~\core_c_psq_MSTAT_reg_DO_reg[0]/P0002  & \core_eu_ea_alu_ea_reg_ay0rwe_DO_reg[5]/P0001  ;
  assign n10685 = \core_c_psq_MSTAT_reg_DO_reg[0]/P0002  & \core_eu_ea_alu_ea_reg_ay0swe_DO_reg[5]/P0001  ;
  assign n10686 = ~n10684 & ~n10685 ;
  assign n10687 = \core_c_dec_MFAY0_E_reg/P0001  & ~n10686 ;
  assign n10704 = \core_c_dec_MFASTAT_E_reg/P0001  & \core_eu_ec_cun_AQ_reg/P0001  ;
  assign n10705 = ~n10687 & ~n10704 ;
  assign n10688 = ~\core_c_psq_MSTAT_reg_DO_reg[0]/P0002  & \core_eu_ea_alu_ea_reg_ay1rwe_DO_reg[5]/P0001  ;
  assign n10689 = \core_c_psq_MSTAT_reg_DO_reg[0]/P0002  & \core_eu_ea_alu_ea_reg_ay1swe_DO_reg[5]/P0001  ;
  assign n10690 = ~n10688 & ~n10689 ;
  assign n10691 = \core_c_dec_MFAY1_E_reg/P0001  & ~n10690 ;
  assign n10692 = ~\core_c_psq_MSTAT_reg_DO_reg[0]/P0002  & \core_eu_ea_alu_ea_reg_arrwe_DO_reg[5]/P0001  ;
  assign n10693 = \core_c_psq_MSTAT_reg_DO_reg[0]/P0002  & \core_eu_ea_alu_ea_reg_arswe_DO_reg[5]/P0001  ;
  assign n10694 = ~n10692 & ~n10693 ;
  assign n10695 = \core_c_dec_MFAR_E_reg/P0001  & ~n10694 ;
  assign n10706 = ~n10691 & ~n10695 ;
  assign n10696 = ~\core_c_psq_MSTAT_reg_DO_reg[0]/P0002  & \core_eu_ea_alu_ea_reg_ax1rwe_DO_reg[5]/P0001  ;
  assign n10697 = \core_c_psq_MSTAT_reg_DO_reg[0]/P0002  & \core_eu_ea_alu_ea_reg_ax1swe_DO_reg[5]/P0001  ;
  assign n10698 = ~n10696 & ~n10697 ;
  assign n10699 = \core_c_dec_MFAX1_E_reg/P0001  & ~n10698 ;
  assign n10700 = ~\core_c_psq_MSTAT_reg_DO_reg[0]/P0002  & \core_eu_ea_alu_ea_reg_ax0rwe_DO_reg[5]/P0001  ;
  assign n10701 = \core_c_psq_MSTAT_reg_DO_reg[0]/P0002  & \core_eu_ea_alu_ea_reg_ax0swe_DO_reg[5]/P0001  ;
  assign n10702 = ~n10700 & ~n10701 ;
  assign n10703 = \core_c_dec_MFAX0_E_reg/P0001  & ~n10702 ;
  assign n10707 = ~n10699 & ~n10703 ;
  assign n10708 = n10706 & n10707 ;
  assign n10709 = n10705 & n10708 ;
  assign n10710 = n7093 & ~n10709 ;
  assign n10787 = ~\core_c_psq_MSTAT_reg_DO_reg[0]/P0002  & \core_eu_es_sht_es_reg_serwe_DO_reg[5]/P0001  ;
  assign n10788 = \core_c_psq_MSTAT_reg_DO_reg[0]/P0002  & \core_eu_es_sht_es_reg_seswe_DO_reg[5]/P0001  ;
  assign n10789 = ~n10787 & ~n10788 ;
  assign n10790 = \core_c_dec_MFSE_E_reg/P0001  & ~n10789 ;
  assign n10803 = ~n7169 & ~n10790 ;
  assign n10799 = ~\core_c_psq_MSTAT_reg_DO_reg[0]/P0002  & \core_eu_es_sht_es_reg_sr0rwe_DO_reg[5]/P0001  ;
  assign n10800 = \core_c_psq_MSTAT_reg_DO_reg[0]/P0002  & \core_eu_es_sht_es_reg_sr0swe_DO_reg[5]/P0001  ;
  assign n10801 = ~n10799 & ~n10800 ;
  assign n10802 = \core_c_dec_MFSR0_E_reg/P0001  & ~n10801 ;
  assign n10791 = ~\core_c_psq_MSTAT_reg_DO_reg[0]/P0002  & \core_eu_es_sht_es_reg_sirwe_DO_reg[5]/P0001  ;
  assign n10792 = \core_c_psq_MSTAT_reg_DO_reg[0]/P0002  & \core_eu_es_sht_es_reg_siswe_DO_reg[5]/P0001  ;
  assign n10793 = ~n10791 & ~n10792 ;
  assign n10794 = \core_c_dec_MFSI_E_reg/P0001  & ~n10793 ;
  assign n10795 = ~\core_c_psq_MSTAT_reg_DO_reg[0]/P0002  & \core_eu_es_sht_es_reg_sr1rwe_DO_reg[5]/P0001  ;
  assign n10796 = \core_c_psq_MSTAT_reg_DO_reg[0]/P0002  & \core_eu_es_sht_es_reg_sr1swe_DO_reg[5]/P0001  ;
  assign n10797 = ~n10795 & ~n10796 ;
  assign n10798 = \core_c_dec_MFSR1_E_reg/P0001  & ~n10797 ;
  assign n10804 = ~n10794 & ~n10798 ;
  assign n10805 = ~n10802 & n10804 ;
  assign n10806 = n10803 & n10805 ;
  assign n10807 = n7153 & ~n10806 ;
  assign n10901 = ~n10710 & ~n10807 ;
  assign n10902 = ~n10890 & n10901 ;
  assign n10903 = n10900 & n10902 ;
  assign n10904 = ~n10786 & n10903 ;
  assign n10905 = ~n10770 & n10904 ;
  assign n10906 = ~n10683 & n10905 ;
  assign n10907 = ~\emc_DMDoe_reg/NET0131  & ~n10906 ;
  assign n10908 = \emc_DMDoe_reg/NET0131  & \emc_DMDreg_reg[5]/P0001  ;
  assign n10909 = n7057 & ~n10908 ;
  assign n10910 = ~n10907 & n10909 ;
  assign n10911 = ~n10682 & ~n10910 ;
  assign n10912 = n6135 & ~n10911 ;
  assign n10913 = n8964 & ~n10912 ;
  assign n10914 = ~n10664 & n10913 ;
  assign n10915 = ~n10641 & ~n10914 ;
  assign n10916 = ~n10421 & n10915 ;
  assign n10917 = \core_dag_ilm2reg_I_reg[6]/NET0131  & ~n6647 ;
  assign n10918 = ~n6753 & ~n6778 ;
  assign n10919 = n6819 & n6821 ;
  assign n10920 = n6776 & ~n10919 ;
  assign n10921 = ~n10918 & ~n10920 ;
  assign n10922 = n10918 & n10920 ;
  assign n10923 = ~n10921 & ~n10922 ;
  assign n10924 = n8198 & n10923 ;
  assign n10925 = ~n6693 & ~n6749 ;
  assign n10926 = n6693 & n6749 ;
  assign n10927 = ~n10925 & ~n10926 ;
  assign n10928 = ~n8198 & n10927 ;
  assign n10929 = ~n10924 & ~n10928 ;
  assign n10930 = ~n10917 & ~n10929 ;
  assign n10931 = ~n6176 & n10930 ;
  assign n10942 = ~n6241 & ~n6511 ;
  assign n10943 = n6266 & ~n10942 ;
  assign n10944 = ~n6266 & n10942 ;
  assign n10945 = ~n10943 & ~n10944 ;
  assign n10950 = ~n6496 & ~n10945 ;
  assign n10933 = ~n6275 & ~n6382 ;
  assign n10934 = n6309 & ~n6372 ;
  assign n10935 = n6380 & ~n10934 ;
  assign n10936 = ~n6260 & ~n10935 ;
  assign n10937 = ~n6375 & ~n10936 ;
  assign n10938 = n10933 & n10937 ;
  assign n10939 = ~n10933 & ~n10937 ;
  assign n10940 = ~n10938 & ~n10939 ;
  assign n10949 = n6496 & n10940 ;
  assign n10951 = ~\core_dag_ilm1reg_M_reg[13]/NET0131  & ~n10949 ;
  assign n10952 = ~n10950 & n10951 ;
  assign n10932 = \core_dag_ilm1reg_I_reg[7]/NET0131  & n6262 ;
  assign n10946 = n7612 & ~n10945 ;
  assign n10941 = ~n7612 & n10940 ;
  assign n10947 = \core_dag_ilm1reg_M_reg[13]/NET0131  & ~n10941 ;
  assign n10948 = ~n10946 & n10947 ;
  assign n10953 = ~n10932 & ~n10948 ;
  assign n10954 = ~n10952 & n10953 ;
  assign n10955 = n6176 & n10954 ;
  assign n10956 = ~n10931 & ~n10955 ;
  assign n10957 = n6135 & ~n10956 ;
  assign n10979 = \core_dag_ilm1reg_I2_we_DO_reg[6]/NET0131  & n6084 ;
  assign n10980 = n6085 & n10979 ;
  assign n10984 = ~n4055 & ~n10980 ;
  assign n10983 = \core_dag_ilm1reg_I0_we_DO_reg[6]/NET0131  & n8131 ;
  assign n10981 = \core_dag_ilm1reg_I1_we_DO_reg[6]/NET0131  & n6142 ;
  assign n10982 = \core_dag_ilm1reg_I3_we_DO_reg[6]/NET0131  & n6140 ;
  assign n10985 = ~n10981 & ~n10982 ;
  assign n10986 = ~n10983 & n10985 ;
  assign n10987 = n10984 & n10986 ;
  assign n10988 = \core_dag_ilm1reg_I0_we_DO_reg[6]/NET0131  & n6148 ;
  assign n10989 = \core_dag_ilm1reg_I1_we_DO_reg[6]/NET0131  & n6154 ;
  assign n10992 = ~n10988 & ~n10989 ;
  assign n10990 = \core_dag_ilm1reg_I3_we_DO_reg[6]/NET0131  & n6150 ;
  assign n10991 = n6095 & n10979 ;
  assign n10993 = ~n10990 & ~n10991 ;
  assign n10994 = n10992 & n10993 ;
  assign n10995 = n4055 & n10994 ;
  assign n10996 = ~n10987 & ~n10995 ;
  assign n10997 = ~n6111 & n10996 ;
  assign n10961 = \core_dag_ilm2reg_I4_we_DO_reg[6]/NET0131  & n6976 ;
  assign n10962 = \core_dag_ilm2reg_I7_we_DO_reg[6]/NET0131  & n6972 ;
  assign n10965 = ~n10961 & ~n10962 ;
  assign n10963 = \core_dag_ilm2reg_I6_we_DO_reg[6]/NET0131  & n6974 ;
  assign n10964 = \core_dag_ilm2reg_I5_we_DO_reg[6]/NET0131  & n6970 ;
  assign n10966 = ~n10963 & ~n10964 ;
  assign n10967 = n10965 & n10966 ;
  assign n10968 = n4055 & ~n10967 ;
  assign n10969 = \core_dag_ilm2reg_I4_we_DO_reg[6]/NET0131  & n6958 ;
  assign n10970 = \core_dag_ilm2reg_I7_we_DO_reg[6]/NET0131  & n6960 ;
  assign n10973 = ~n10969 & ~n10970 ;
  assign n10971 = \core_dag_ilm2reg_I6_we_DO_reg[6]/NET0131  & n6962 ;
  assign n10972 = \core_dag_ilm2reg_I5_we_DO_reg[6]/NET0131  & n6964 ;
  assign n10974 = ~n10971 & ~n10972 ;
  assign n10975 = n10973 & n10974 ;
  assign n10976 = ~n10968 & n10975 ;
  assign n10977 = ~n6121 & ~n10976 ;
  assign n10978 = \core_c_dec_IR_reg[10]/NET0131  & n6956 ;
  assign n10998 = ~n10977 & ~n10978 ;
  assign n10999 = ~n10997 & n10998 ;
  assign n11000 = n5949 & ~n10999 ;
  assign n11001 = \core_dag_ilm1reg_DMA_pi_DO_reg[6]/NET0131  & ~n6934 ;
  assign n10959 = \idma_DCTL_reg[6]/NET0131  & n6926 ;
  assign n10960 = \core_dag_ilm1reg_STAC_pi_DO_reg[6]/NET0131  & n6988 ;
  assign n11002 = ~n10959 & ~n10960 ;
  assign n11003 = n6924 & n11002 ;
  assign n11004 = ~n11001 & n11003 ;
  assign n11005 = ~n11000 & n11004 ;
  assign n10958 = ~\bdma_BIAD_reg[6]/NET0131  & ~n6924 ;
  assign n11006 = ~n6176 & ~n10958 ;
  assign n11007 = ~n11005 & n11006 ;
  assign n11008 = \core_dag_ilm1reg_I2_we_DO_reg[7]/NET0131  & n6084 ;
  assign n11009 = n6085 & n11008 ;
  assign n11013 = ~n4055 & ~n11009 ;
  assign n11012 = \core_dag_ilm1reg_I0_we_DO_reg[7]/NET0131  & n8131 ;
  assign n11010 = \core_dag_ilm1reg_I3_we_DO_reg[7]/NET0131  & n6140 ;
  assign n11011 = \core_dag_ilm1reg_I1_we_DO_reg[7]/NET0131  & n6142 ;
  assign n11014 = ~n11010 & ~n11011 ;
  assign n11015 = ~n11012 & n11014 ;
  assign n11016 = n11013 & n11015 ;
  assign n11017 = \core_dag_ilm1reg_I0_we_DO_reg[7]/NET0131  & n6148 ;
  assign n11018 = \core_dag_ilm1reg_I1_we_DO_reg[7]/NET0131  & n6154 ;
  assign n11021 = ~n11017 & ~n11018 ;
  assign n11019 = \core_dag_ilm1reg_I3_we_DO_reg[7]/NET0131  & n6150 ;
  assign n11020 = n6095 & n11008 ;
  assign n11022 = ~n11019 & ~n11020 ;
  assign n11023 = n11021 & n11022 ;
  assign n11024 = n4055 & n11023 ;
  assign n11025 = ~n11016 & ~n11024 ;
  assign n11026 = n6176 & n11025 ;
  assign n11027 = ~n6135 & ~n11026 ;
  assign n11028 = ~n11007 & n11027 ;
  assign n11029 = ~n7005 & ~n11028 ;
  assign n11030 = ~n10957 & n11029 ;
  assign n11031 = n10976 & ~n10996 ;
  assign n11032 = n8153 & ~n11031 ;
  assign n11039 = \DM_rd0[7]_pad  & ~n7053 ;
  assign n11033 = \DM_rdm[7]_pad  & n7016 ;
  assign n11044 = ~n7057 & ~n11033 ;
  assign n11036 = \DM_rd6[7]_pad  & n7031 ;
  assign n11037 = \DM_rd7[7]_pad  & n7034 ;
  assign n11045 = ~n11036 & ~n11037 ;
  assign n11046 = n11044 & n11045 ;
  assign n11040 = \DM_rd5[7]_pad  & n7043 ;
  assign n11035 = \DM_rd4[7]_pad  & n7028 ;
  assign n11041 = \DM_rd2[7]_pad  & n7041 ;
  assign n11034 = \DM_rd1[7]_pad  & n7022 ;
  assign n11038 = \DM_rd3[7]_pad  & n7038 ;
  assign n11042 = ~n11034 & ~n11038 ;
  assign n11043 = ~n11041 & n11042 ;
  assign n11047 = ~n11035 & n11043 ;
  assign n11048 = ~n11040 & n11047 ;
  assign n11049 = n11046 & n11048 ;
  assign n11050 = ~n11039 & n11049 ;
  assign n11051 = \regout_STD_C_reg[7]/P0001  & n6988 ;
  assign n11092 = \bdma_BIAD_reg[7]/NET0131  & n7234 ;
  assign n11083 = \emc_WSCRreg_DO_reg[7]/NET0131  & n7251 ;
  assign n11084 = \tm_TCR_TMP_reg[7]/NET0131  & n7289 ;
  assign n11109 = ~n11083 & ~n11084 ;
  assign n11085 = \sport0_regs_SCLKDIVreg_DO_reg[7]/NET0131  & n7256 ;
  assign n11086 = \sport0_regs_AUTOreg_DO_reg[7]/NET0131  & n7295 ;
  assign n11110 = ~n11085 & ~n11086 ;
  assign n11123 = n11109 & n11110 ;
  assign n11079 = \sport1_regs_MWORDreg_DO_reg[7]/NET0131  & n7263 ;
  assign n11107 = ~n7522 & ~n11079 ;
  assign n11080 = \emc_WSCRext_reg_DO_reg[7]/NET0131  & n7514 ;
  assign n11081 = \tm_tpr_reg_DO_reg[7]/NET0131  & n7293 ;
  assign n11108 = ~n11080 & ~n11081 ;
  assign n11124 = n11107 & n11108 ;
  assign n11125 = n11123 & n11124 ;
  assign n11129 = ~n11092 & n11125 ;
  assign n11100 = \bdma_BEAD_reg[7]/NET0131  & n7303 ;
  assign n11101 = \bdma_BCTL_reg[7]/NET0131  & n7230 ;
  assign n11130 = ~n11100 & ~n11101 ;
  assign n11131 = n11129 & n11130 ;
  assign n11097 = \bdma_BOVL_reg[7]/NET0131  & n7534 ;
  assign n11082 = \bdma_BWCOUNT_reg[7]/NET0131  & n7287 ;
  assign n11091 = \pio_pmask_reg_DO_reg[7]/NET0131  & n7297 ;
  assign n11093 = \sport1_regs_SCLKDIVreg_DO_reg[7]/NET0131  & n7247 ;
  assign n11113 = ~n11091 & ~n11093 ;
  assign n11094 = \sport0_regs_MWORDreg_DO_reg[7]/NET0131  & n7276 ;
  assign n11095 = \sport0_regs_SCTLreg_DO_reg[7]/NET0131  & n7249 ;
  assign n11114 = ~n11094 & ~n11095 ;
  assign n11121 = n11113 & n11114 ;
  assign n11087 = \idma_DOVL_reg[7]/NET0131  & n7532 ;
  assign n11088 = \tm_tsr_reg_DO_reg[7]/NET0131  & n7540 ;
  assign n11111 = ~n11087 & ~n11088 ;
  assign n11089 = \sport1_regs_FSDIVreg_DO_reg[7]/NET0131  & n7273 ;
  assign n11090 = \sport0_regs_FSDIVreg_DO_reg[7]/NET0131  & n7259 ;
  assign n11112 = ~n11089 & ~n11090 ;
  assign n11122 = n11111 & n11112 ;
  assign n11126 = n11121 & n11122 ;
  assign n11103 = \sport1_regs_SCTLreg_DO_reg[7]/NET0131  & n7281 ;
  assign n11104 = \PIO_out[7]_pad  & n7291 ;
  assign n11117 = ~n11103 & ~n11104 ;
  assign n11105 = \PIO_oe[7]_pad  & n7244 ;
  assign n11106 = \idma_DCTL_reg[7]/NET0131  & n7299 ;
  assign n11118 = ~n11105 & ~n11106 ;
  assign n11119 = n11117 & n11118 ;
  assign n11096 = \sport1_regs_AUTOreg_DO_reg[7]/NET0131  & n7527 ;
  assign n11098 = \clkc_ckr_reg_DO_reg[7]/NET0131  & n7239 ;
  assign n11115 = ~n11096 & ~n11098 ;
  assign n11099 = \memc_usysr_DO_reg[7]/NET0131  & n7301 ;
  assign n11102 = \pio_PINT_reg[7]/NET0131  & n7271 ;
  assign n11116 = ~n11099 & ~n11102 ;
  assign n11120 = n11115 & n11116 ;
  assign n11127 = n11119 & n11120 ;
  assign n11128 = n11126 & n11127 ;
  assign n11132 = ~n11082 & n11128 ;
  assign n11133 = ~n11097 & n11132 ;
  assign n11134 = n11131 & n11133 ;
  assign n11135 = \memc_ldSREG_E_reg/NET0131  & ~n11134 ;
  assign n11140 = \core_c_dec_MFtoppcs_Eg_reg/P0001  & ~n4656 ;
  assign n11142 = \core_c_dec_MFIMASK_E_reg/P0001  & \core_c_psq_IMASK_reg[7]/NET0131  ;
  assign n11139 = \core_c_dec_MFSSTAT_E_reg/P0001  & \core_c_psq_SSTAT_reg[7]/NET0131  ;
  assign n11141 = \core_c_dec_MFIDR_E_reg/P0001  & \sice_idr0_reg_DO_reg[7]/P0001  ;
  assign n11144 = ~n11139 & ~n11141 ;
  assign n11145 = ~n11142 & n11144 ;
  assign n11137 = \core_c_dec_IRE_reg[11]/NET0131  & ~n7216 ;
  assign n11136 = \core_c_dec_MFPMOVL_E_reg/P0001  & \core_c_psq_PMOVL_regh_DO_reg[3]/NET0131  ;
  assign n11138 = \core_c_dec_MFCNTR_E_reg/P0001  & \core_c_psq_CNTR_reg_DO_reg[7]/NET0131  ;
  assign n11143 = ~n11136 & ~n11138 ;
  assign n11146 = ~n11137 & n11143 ;
  assign n11147 = n11145 & n11146 ;
  assign n11148 = ~n11140 & n11147 ;
  assign n11149 = n7215 & ~n11148 ;
  assign n11213 = \core_c_dec_MFLreg_E_reg[6]/P0001  & \core_dag_ilm2reg_L6_we_DO_reg[7]/NET0131  ;
  assign n11214 = \core_c_dec_MFIreg_E_reg[6]/P0001  & \core_dag_ilm2reg_I6_we_DO_reg[7]/NET0131  ;
  assign n11221 = ~n11213 & ~n11214 ;
  assign n11215 = \core_c_dec_MFIreg_E_reg[5]/P0001  & \core_dag_ilm2reg_I5_we_DO_reg[7]/NET0131  ;
  assign n11216 = \core_c_dec_MFLreg_E_reg[5]/P0001  & \core_dag_ilm2reg_L5_we_DO_reg[7]/NET0131  ;
  assign n11222 = ~n11215 & ~n11216 ;
  assign n11223 = n11221 & n11222 ;
  assign n11209 = \core_c_dec_MFIreg_E_reg[7]/P0001  & \core_dag_ilm2reg_I7_we_DO_reg[7]/NET0131  ;
  assign n11210 = \core_c_dec_MFLreg_E_reg[4]/P0001  & \core_dag_ilm2reg_L4_we_DO_reg[7]/NET0131  ;
  assign n11219 = ~n11209 & ~n11210 ;
  assign n11211 = \core_c_dec_MFMreg_E_reg[4]/P0001  & \core_dag_ilm2reg_M4_we_DO_reg[7]/NET0131  ;
  assign n11212 = \core_c_dec_MFLreg_E_reg[7]/P0001  & \core_dag_ilm2reg_L7_we_DO_reg[7]/NET0131  ;
  assign n11220 = ~n11211 & ~n11212 ;
  assign n11224 = n11219 & n11220 ;
  assign n11205 = \core_c_dec_MFMreg_E_reg[5]/P0001  & \core_dag_ilm2reg_M5_we_DO_reg[7]/NET0131  ;
  assign n11206 = \core_c_dec_MFMreg_E_reg[7]/P0001  & \core_dag_ilm2reg_M7_we_DO_reg[7]/NET0131  ;
  assign n11217 = ~n11205 & ~n11206 ;
  assign n11207 = \core_c_dec_MFMreg_E_reg[6]/P0001  & \core_dag_ilm2reg_M6_we_DO_reg[7]/NET0131  ;
  assign n11208 = \core_c_dec_MFIreg_E_reg[4]/P0001  & \core_dag_ilm2reg_I4_we_DO_reg[7]/NET0131  ;
  assign n11218 = ~n11207 & ~n11208 ;
  assign n11225 = n11217 & n11218 ;
  assign n11226 = n11224 & n11225 ;
  assign n11227 = n11223 & n11226 ;
  assign n11228 = n7128 & ~n11227 ;
  assign n11158 = \core_c_dec_MFIreg_E_reg[0]/P0001  & \core_dag_ilm1reg_I0_we_DO_reg[7]/NET0131  ;
  assign n11159 = \core_c_dec_MFIreg_E_reg[3]/P0001  & \core_dag_ilm1reg_I3_we_DO_reg[7]/NET0131  ;
  assign n11166 = ~n11158 & ~n11159 ;
  assign n11160 = \core_c_dec_MFLreg_E_reg[0]/P0001  & \core_dag_ilm1reg_L0_we_DO_reg[7]/NET0131  ;
  assign n11161 = \core_c_dec_MFLreg_E_reg[1]/P0001  & \core_dag_ilm1reg_L1_we_DO_reg[7]/NET0131  ;
  assign n11167 = ~n11160 & ~n11161 ;
  assign n11168 = n11166 & n11167 ;
  assign n11154 = \core_c_dec_MFIreg_E_reg[1]/P0001  & \core_dag_ilm1reg_I1_we_DO_reg[7]/NET0131  ;
  assign n11155 = \core_c_dec_MFLreg_E_reg[3]/P0001  & \core_dag_ilm1reg_L3_we_DO_reg[7]/NET0131  ;
  assign n11164 = ~n11154 & ~n11155 ;
  assign n11156 = \core_c_dec_MFIreg_E_reg[2]/P0001  & \core_dag_ilm1reg_I2_we_DO_reg[7]/NET0131  ;
  assign n11157 = \core_c_dec_MFMreg_E_reg[1]/P0001  & \core_dag_ilm1reg_M1_we_DO_reg[7]/NET0131  ;
  assign n11165 = ~n11156 & ~n11157 ;
  assign n11169 = n11164 & n11165 ;
  assign n11150 = \core_c_dec_MFMreg_E_reg[3]/P0001  & \core_dag_ilm1reg_M3_we_DO_reg[7]/NET0131  ;
  assign n11151 = \core_c_dec_MFMreg_E_reg[0]/P0001  & \core_dag_ilm1reg_M0_we_DO_reg[7]/NET0131  ;
  assign n11162 = ~n11150 & ~n11151 ;
  assign n11152 = \core_c_dec_MFMreg_E_reg[2]/P0001  & \core_dag_ilm1reg_M2_we_DO_reg[7]/NET0131  ;
  assign n11153 = \core_c_dec_MFLreg_E_reg[2]/P0001  & \core_dag_ilm1reg_L2_we_DO_reg[7]/NET0131  ;
  assign n11163 = ~n11152 & ~n11153 ;
  assign n11170 = n11162 & n11163 ;
  assign n11171 = n11169 & n11170 ;
  assign n11172 = n11168 & n11171 ;
  assign n11173 = n7068 & ~n11172 ;
  assign n11245 = \core_c_dec_MFTX1_E_reg/P0001  & \sport1_txctl_TX_reg[7]/P0001  ;
  assign n11246 = \core_c_dec_MFTX0_E_reg/P0001  & \sport0_txctl_TX_reg[7]/P0001  ;
  assign n11249 = ~n11245 & ~n11246 ;
  assign n11247 = \core_c_dec_MFRX1_E_reg/P0001  & \sport1_rxctl_RX_reg[7]/P0001  ;
  assign n11248 = \core_c_dec_MFRX0_E_reg/P0001  & \sport0_rxctl_RX_reg[7]/P0001  ;
  assign n11250 = ~n11247 & ~n11248 ;
  assign n11251 = n11249 & n11250 ;
  assign n11252 = n7119 & ~n11251 ;
  assign n11253 = ~n11173 & ~n11252 ;
  assign n11254 = ~n11228 & n11253 ;
  assign n11237 = ~\core_c_psq_MSTAT_reg_DO_reg[0]/P0002  & \core_eu_es_sht_es_reg_sr1rwe_DO_reg[7]/P0001  ;
  assign n11238 = \core_c_psq_MSTAT_reg_DO_reg[0]/P0002  & \core_eu_es_sht_es_reg_sr1swe_DO_reg[7]/P0001  ;
  assign n11239 = ~n11237 & ~n11238 ;
  assign n11240 = \core_c_dec_MFSR1_E_reg/P0001  & ~n11239 ;
  assign n11229 = ~\core_c_psq_MSTAT_reg_DO_reg[0]/P0002  & \core_eu_es_sht_es_reg_sr0rwe_DO_reg[7]/P0001  ;
  assign n11230 = \core_c_psq_MSTAT_reg_DO_reg[0]/P0002  & \core_eu_es_sht_es_reg_sr0swe_DO_reg[7]/P0001  ;
  assign n11231 = ~n11229 & ~n11230 ;
  assign n11232 = \core_c_dec_MFSR0_E_reg/P0001  & ~n11231 ;
  assign n11233 = ~\core_c_psq_MSTAT_reg_DO_reg[0]/P0002  & \core_eu_es_sht_es_reg_sirwe_DO_reg[7]/P0001  ;
  assign n11234 = \core_c_psq_MSTAT_reg_DO_reg[0]/P0002  & \core_eu_es_sht_es_reg_siswe_DO_reg[7]/P0001  ;
  assign n11235 = ~n11233 & ~n11234 ;
  assign n11236 = \core_c_dec_MFSI_E_reg/P0001  & ~n11235 ;
  assign n11241 = ~n11232 & ~n11236 ;
  assign n11242 = ~n11240 & n11241 ;
  assign n11243 = n7174 & n11242 ;
  assign n11244 = n7153 & ~n11243 ;
  assign n11052 = ~\core_c_psq_MSTAT_reg_DO_reg[0]/P0002  & \core_eu_ea_alu_ea_reg_ay0rwe_DO_reg[7]/P0001  ;
  assign n11053 = \core_c_psq_MSTAT_reg_DO_reg[0]/P0002  & \core_eu_ea_alu_ea_reg_ay0swe_DO_reg[7]/P0001  ;
  assign n11054 = ~n11052 & ~n11053 ;
  assign n11055 = \core_c_dec_MFAY0_E_reg/P0001  & ~n11054 ;
  assign n11072 = \core_c_dec_MFASTAT_E_reg/P0001  & \core_eu_ec_cun_SS_reg/P0001  ;
  assign n11073 = ~n11055 & ~n11072 ;
  assign n11056 = ~\core_c_psq_MSTAT_reg_DO_reg[0]/P0002  & \core_eu_ea_alu_ea_reg_ay1rwe_DO_reg[7]/P0001  ;
  assign n11057 = \core_c_psq_MSTAT_reg_DO_reg[0]/P0002  & \core_eu_ea_alu_ea_reg_ay1swe_DO_reg[7]/P0001  ;
  assign n11058 = ~n11056 & ~n11057 ;
  assign n11059 = \core_c_dec_MFAY1_E_reg/P0001  & ~n11058 ;
  assign n11060 = ~\core_c_psq_MSTAT_reg_DO_reg[0]/P0002  & \core_eu_ea_alu_ea_reg_arrwe_DO_reg[7]/P0001  ;
  assign n11061 = \core_c_psq_MSTAT_reg_DO_reg[0]/P0002  & \core_eu_ea_alu_ea_reg_arswe_DO_reg[7]/P0001  ;
  assign n11062 = ~n11060 & ~n11061 ;
  assign n11063 = \core_c_dec_MFAR_E_reg/P0001  & ~n11062 ;
  assign n11074 = ~n11059 & ~n11063 ;
  assign n11064 = ~\core_c_psq_MSTAT_reg_DO_reg[0]/P0002  & \core_eu_ea_alu_ea_reg_ax1rwe_DO_reg[7]/P0001  ;
  assign n11065 = \core_c_psq_MSTAT_reg_DO_reg[0]/P0002  & \core_eu_ea_alu_ea_reg_ax1swe_DO_reg[7]/P0001  ;
  assign n11066 = ~n11064 & ~n11065 ;
  assign n11067 = \core_c_dec_MFAX1_E_reg/P0001  & ~n11066 ;
  assign n11068 = ~\core_c_psq_MSTAT_reg_DO_reg[0]/P0002  & \core_eu_ea_alu_ea_reg_ax0rwe_DO_reg[7]/P0001  ;
  assign n11069 = \core_c_psq_MSTAT_reg_DO_reg[0]/P0002  & \core_eu_ea_alu_ea_reg_ax0swe_DO_reg[7]/P0001  ;
  assign n11070 = ~n11068 & ~n11069 ;
  assign n11071 = \core_c_dec_MFAX0_E_reg/P0001  & ~n11070 ;
  assign n11075 = ~n11067 & ~n11071 ;
  assign n11076 = n11074 & n11075 ;
  assign n11077 = n11073 & n11076 ;
  assign n11078 = n7093 & ~n11077 ;
  assign n11194 = ~\core_c_psq_MSTAT_reg_DO_reg[0]/P0002  & \core_eu_em_mac_em_reg_mr1rwe_DO_reg[7]/P0001  ;
  assign n11195 = \core_c_psq_MSTAT_reg_DO_reg[0]/P0002  & \core_eu_em_mac_em_reg_mr1swe_DO_reg[7]/P0001  ;
  assign n11196 = ~n11194 & ~n11195 ;
  assign n11197 = \core_c_dec_MFMR1_E_reg/P0001  & ~n11196 ;
  assign n11186 = ~\core_c_psq_MSTAT_reg_DO_reg[0]/P0002  & \core_eu_em_mac_em_reg_mx1rwe_DO_reg[7]/P0001  ;
  assign n11187 = \core_c_psq_MSTAT_reg_DO_reg[0]/P0002  & \core_eu_em_mac_em_reg_mx1swe_DO_reg[7]/P0001  ;
  assign n11188 = ~n11186 & ~n11187 ;
  assign n11189 = \core_c_dec_MFMX1_E_reg/P0001  & ~n11188 ;
  assign n11190 = ~\core_c_psq_MSTAT_reg_DO_reg[0]/P0002  & \core_eu_em_mac_em_reg_mr0rwe_DO_reg[7]/P0001  ;
  assign n11191 = \core_c_psq_MSTAT_reg_DO_reg[0]/P0002  & \core_eu_em_mac_em_reg_mr0swe_DO_reg[7]/P0001  ;
  assign n11192 = ~n11190 & ~n11191 ;
  assign n11193 = \core_c_dec_MFMR0_E_reg/P0001  & ~n11192 ;
  assign n11200 = ~n11189 & ~n11193 ;
  assign n11201 = ~n11197 & n11200 ;
  assign n11174 = ~\core_c_psq_MSTAT_reg_DO_reg[0]/P0002  & \core_eu_em_mac_em_reg_my0rwe_DO_reg[7]/P0001  ;
  assign n11175 = \core_c_psq_MSTAT_reg_DO_reg[0]/P0002  & \core_eu_em_mac_em_reg_my0swe_DO_reg[7]/P0001  ;
  assign n11176 = ~n11174 & ~n11175 ;
  assign n11177 = \core_c_dec_MFMY0_E_reg/P0001  & ~n11176 ;
  assign n11198 = ~n7207 & ~n11177 ;
  assign n11178 = ~\core_c_psq_MSTAT_reg_DO_reg[0]/P0002  & \core_eu_em_mac_em_reg_my1rwe_DO_reg[7]/P0001  ;
  assign n11179 = \core_c_psq_MSTAT_reg_DO_reg[0]/P0002  & \core_eu_em_mac_em_reg_my1swe_DO_reg[7]/P0001  ;
  assign n11180 = ~n11178 & ~n11179 ;
  assign n11181 = \core_c_dec_MFMY1_E_reg/P0001  & ~n11180 ;
  assign n11182 = ~\core_c_psq_MSTAT_reg_DO_reg[0]/P0002  & \core_eu_em_mac_em_reg_mx0rwe_DO_reg[7]/P0001  ;
  assign n11183 = \core_c_psq_MSTAT_reg_DO_reg[0]/P0002  & \core_eu_em_mac_em_reg_mx0swe_DO_reg[7]/P0001  ;
  assign n11184 = ~n11182 & ~n11183 ;
  assign n11185 = \core_c_dec_MFMX0_E_reg/P0001  & ~n11184 ;
  assign n11199 = ~n11181 & ~n11185 ;
  assign n11202 = n11198 & n11199 ;
  assign n11203 = n11201 & n11202 ;
  assign n11204 = n7179 & ~n11203 ;
  assign n11255 = ~n11078 & ~n11204 ;
  assign n11256 = ~n11244 & n11255 ;
  assign n11257 = n11254 & n11256 ;
  assign n11258 = ~n11149 & n11257 ;
  assign n11259 = ~n11135 & n11258 ;
  assign n11260 = ~n11051 & n11259 ;
  assign n11261 = ~\emc_DMDoe_reg/NET0131  & ~n11260 ;
  assign n11262 = \emc_DMDoe_reg/NET0131  & \emc_DMDreg_reg[7]/P0001  ;
  assign n11263 = n7057 & ~n11262 ;
  assign n11264 = ~n11261 & n11263 ;
  assign n11265 = ~n11050 & ~n11264 ;
  assign n11266 = n7863 & n11265 ;
  assign n11267 = ~n11032 & ~n11266 ;
  assign n11268 = n7005 & ~n11267 ;
  assign n11274 = ~n6260 & ~n6375 ;
  assign n11275 = ~n10935 & n11274 ;
  assign n11276 = n10935 & ~n11274 ;
  assign n11277 = ~n11275 & ~n11276 ;
  assign n11278 = ~n7631 & n11277 ;
  assign n11269 = \core_dag_ilm1reg_I_reg[6]/NET0131  & ~n6238 ;
  assign n11270 = ~n6242 & ~n6510 ;
  assign n11271 = n6242 & n6510 ;
  assign n11272 = ~n11270 & ~n11271 ;
  assign n11273 = n7631 & ~n11272 ;
  assign n11279 = ~n11269 & ~n11273 ;
  assign n11280 = ~n11278 & n11279 ;
  assign n11281 = ~n6135 & n11280 ;
  assign n11288 = \DM_rd0[6]_pad  & ~n7053 ;
  assign n11282 = \DM_rdm[6]_pad  & n7016 ;
  assign n11293 = ~n7057 & ~n11282 ;
  assign n11285 = \DM_rd6[6]_pad  & n7031 ;
  assign n11286 = \DM_rd7[6]_pad  & n7034 ;
  assign n11294 = ~n11285 & ~n11286 ;
  assign n11295 = n11293 & n11294 ;
  assign n11289 = \DM_rd5[6]_pad  & n7043 ;
  assign n11284 = \DM_rd4[6]_pad  & n7028 ;
  assign n11290 = \DM_rd2[6]_pad  & n7041 ;
  assign n11283 = \DM_rd1[6]_pad  & n7022 ;
  assign n11287 = \DM_rd3[6]_pad  & n7038 ;
  assign n11291 = ~n11283 & ~n11287 ;
  assign n11292 = ~n11290 & n11291 ;
  assign n11296 = ~n11284 & n11292 ;
  assign n11297 = ~n11289 & n11296 ;
  assign n11298 = n11295 & n11297 ;
  assign n11299 = ~n11288 & n11298 ;
  assign n11300 = \regout_STD_C_reg[6]/P0001  & n6988 ;
  assign n11322 = \core_c_dec_MFASTAT_E_reg/P0001  & ~n4174 ;
  assign n11323 = ~\core_c_psq_MSTAT_reg_DO_reg[0]/P0002  & \core_eu_ea_alu_ea_reg_ax0rwe_DO_reg[6]/P0001  ;
  assign n11324 = \core_c_psq_MSTAT_reg_DO_reg[0]/P0002  & \core_eu_ea_alu_ea_reg_ax0swe_DO_reg[6]/P0001  ;
  assign n11325 = ~n11323 & ~n11324 ;
  assign n11326 = \core_c_dec_MFAX0_E_reg/P0001  & ~n11325 ;
  assign n11327 = ~\core_c_psq_MSTAT_reg_DO_reg[0]/P0002  & \core_eu_ea_alu_ea_reg_ay0rwe_DO_reg[6]/P0001  ;
  assign n11328 = \core_c_psq_MSTAT_reg_DO_reg[0]/P0002  & \core_eu_ea_alu_ea_reg_ay0swe_DO_reg[6]/P0001  ;
  assign n11329 = ~n11327 & ~n11328 ;
  assign n11330 = \core_c_dec_MFAY0_E_reg/P0001  & ~n11329 ;
  assign n11343 = ~n11326 & ~n11330 ;
  assign n11339 = ~\core_c_psq_MSTAT_reg_DO_reg[0]/P0002  & \core_eu_ea_alu_ea_reg_arrwe_DO_reg[6]/P0001  ;
  assign n11340 = \core_c_psq_MSTAT_reg_DO_reg[0]/P0002  & \core_eu_ea_alu_ea_reg_arswe_DO_reg[6]/P0001  ;
  assign n11341 = ~n11339 & ~n11340 ;
  assign n11342 = \core_c_dec_MFAR_E_reg/P0001  & ~n11341 ;
  assign n11331 = ~\core_c_psq_MSTAT_reg_DO_reg[0]/P0002  & \core_eu_ea_alu_ea_reg_ay1rwe_DO_reg[6]/P0001  ;
  assign n11332 = \core_c_psq_MSTAT_reg_DO_reg[0]/P0002  & \core_eu_ea_alu_ea_reg_ay1swe_DO_reg[6]/P0001  ;
  assign n11333 = ~n11331 & ~n11332 ;
  assign n11334 = \core_c_dec_MFAY1_E_reg/P0001  & ~n11333 ;
  assign n11335 = ~\core_c_psq_MSTAT_reg_DO_reg[0]/P0002  & \core_eu_ea_alu_ea_reg_ax1rwe_DO_reg[6]/P0001  ;
  assign n11336 = \core_c_psq_MSTAT_reg_DO_reg[0]/P0002  & \core_eu_ea_alu_ea_reg_ax1swe_DO_reg[6]/P0001  ;
  assign n11337 = ~n11335 & ~n11336 ;
  assign n11338 = \core_c_dec_MFAX1_E_reg/P0001  & ~n11337 ;
  assign n11344 = ~n11334 & ~n11338 ;
  assign n11345 = ~n11342 & n11344 ;
  assign n11346 = n11343 & n11345 ;
  assign n11347 = ~n11322 & n11346 ;
  assign n11348 = n7093 & ~n11347 ;
  assign n11362 = \bdma_BIAD_reg[6]/NET0131  & n7234 ;
  assign n11353 = \emc_WSCRreg_DO_reg[6]/NET0131  & n7251 ;
  assign n11354 = \tm_TCR_TMP_reg[6]/NET0131  & n7289 ;
  assign n11379 = ~n11353 & ~n11354 ;
  assign n11355 = \sport0_regs_SCLKDIVreg_DO_reg[6]/NET0131  & n7256 ;
  assign n11356 = \sport0_regs_AUTOreg_DO_reg[6]/NET0131  & n7295 ;
  assign n11380 = ~n11355 & ~n11356 ;
  assign n11393 = n11379 & n11380 ;
  assign n11349 = \sport1_regs_MWORDreg_DO_reg[6]/NET0131  & n7263 ;
  assign n11377 = ~n7522 & ~n11349 ;
  assign n11350 = \emc_WSCRext_reg_DO_reg[6]/NET0131  & n7514 ;
  assign n11351 = \tm_tpr_reg_DO_reg[6]/NET0131  & n7293 ;
  assign n11378 = ~n11350 & ~n11351 ;
  assign n11394 = n11377 & n11378 ;
  assign n11395 = n11393 & n11394 ;
  assign n11399 = ~n11362 & n11395 ;
  assign n11370 = \bdma_BEAD_reg[6]/NET0131  & n7303 ;
  assign n11371 = \bdma_BCTL_reg[6]/NET0131  & n7230 ;
  assign n11400 = ~n11370 & ~n11371 ;
  assign n11401 = n11399 & n11400 ;
  assign n11367 = \bdma_BOVL_reg[6]/NET0131  & n7534 ;
  assign n11352 = \bdma_BWCOUNT_reg[6]/NET0131  & n7287 ;
  assign n11361 = \pio_pmask_reg_DO_reg[6]/NET0131  & n7297 ;
  assign n11363 = \sport1_regs_SCLKDIVreg_DO_reg[6]/NET0131  & n7247 ;
  assign n11383 = ~n11361 & ~n11363 ;
  assign n11364 = \sport0_regs_MWORDreg_DO_reg[6]/NET0131  & n7276 ;
  assign n11365 = \sport0_regs_SCTLreg_DO_reg[6]/NET0131  & n7249 ;
  assign n11384 = ~n11364 & ~n11365 ;
  assign n11391 = n11383 & n11384 ;
  assign n11357 = \idma_DOVL_reg[6]/NET0131  & n7532 ;
  assign n11358 = \tm_tsr_reg_DO_reg[6]/NET0131  & n7540 ;
  assign n11381 = ~n11357 & ~n11358 ;
  assign n11359 = \sport1_regs_FSDIVreg_DO_reg[6]/NET0131  & n7273 ;
  assign n11360 = \sport0_regs_FSDIVreg_DO_reg[6]/NET0131  & n7259 ;
  assign n11382 = ~n11359 & ~n11360 ;
  assign n11392 = n11381 & n11382 ;
  assign n11396 = n11391 & n11392 ;
  assign n11373 = \sport1_regs_SCTLreg_DO_reg[6]/NET0131  & n7281 ;
  assign n11374 = \PIO_out[6]_pad  & n7291 ;
  assign n11387 = ~n11373 & ~n11374 ;
  assign n11375 = \PIO_oe[6]_pad  & n7244 ;
  assign n11376 = \idma_DCTL_reg[6]/NET0131  & n7299 ;
  assign n11388 = ~n11375 & ~n11376 ;
  assign n11389 = n11387 & n11388 ;
  assign n11366 = \sport1_regs_AUTOreg_DO_reg[6]/NET0131  & n7527 ;
  assign n11368 = \clkc_ckr_reg_DO_reg[6]/NET0131  & n7239 ;
  assign n11385 = ~n11366 & ~n11368 ;
  assign n11369 = \memc_usysr_DO_reg[6]/NET0131  & n7301 ;
  assign n11372 = \pio_PINT_reg[6]/NET0131  & n7271 ;
  assign n11386 = ~n11369 & ~n11372 ;
  assign n11390 = n11385 & n11386 ;
  assign n11397 = n11389 & n11390 ;
  assign n11398 = n11396 & n11397 ;
  assign n11402 = ~n11352 & n11398 ;
  assign n11403 = ~n11367 & n11402 ;
  assign n11404 = n11401 & n11403 ;
  assign n11405 = \memc_ldSREG_E_reg/NET0131  & ~n11404 ;
  assign n11407 = \core_c_dec_MFtoppcs_Eg_reg/P0001  & ~n4392 ;
  assign n11410 = \core_c_dec_MFIDR_E_reg/P0001  & \sice_idr0_reg_DO_reg[6]/P0001  ;
  assign n11411 = \core_c_dec_MFMSTAT_E_reg/P0001  & \core_c_psq_MSTAT_reg_DO_reg[6]/NET0131  ;
  assign n11415 = ~n11410 & ~n11411 ;
  assign n11412 = \core_c_dec_MFSSTAT_E_reg/P0001  & \core_c_psq_SSTAT_reg[6]/NET0131  ;
  assign n11413 = \core_c_dec_MFPMOVL_E_reg/P0001  & \core_c_psq_PMOVL_regh_DO_reg[2]/NET0131  ;
  assign n11416 = ~n11412 & ~n11413 ;
  assign n11417 = n11415 & n11416 ;
  assign n11408 = \core_c_dec_IRE_reg[10]/NET0131  & ~n7216 ;
  assign n11406 = \core_c_dec_MFIMASK_E_reg/P0001  & \core_c_psq_IMASK_reg[6]/NET0131  ;
  assign n11409 = \core_c_dec_MFCNTR_E_reg/P0001  & \core_c_psq_CNTR_reg_DO_reg[6]/NET0131  ;
  assign n11414 = ~n11406 & ~n11409 ;
  assign n11418 = ~n11408 & n11414 ;
  assign n11419 = n11417 & n11418 ;
  assign n11420 = ~n11407 & n11419 ;
  assign n11421 = n7215 & ~n11420 ;
  assign n11489 = \core_c_dec_MFIreg_E_reg[7]/P0001  & \core_dag_ilm2reg_I7_we_DO_reg[6]/NET0131  ;
  assign n11490 = \core_c_dec_MFIreg_E_reg[4]/P0001  & \core_dag_ilm2reg_I4_we_DO_reg[6]/NET0131  ;
  assign n11497 = ~n11489 & ~n11490 ;
  assign n11491 = \core_c_dec_MFIreg_E_reg[5]/P0001  & \core_dag_ilm2reg_I5_we_DO_reg[6]/NET0131  ;
  assign n11492 = \core_c_dec_MFIreg_E_reg[6]/P0001  & \core_dag_ilm2reg_I6_we_DO_reg[6]/NET0131  ;
  assign n11498 = ~n11491 & ~n11492 ;
  assign n11499 = n11497 & n11498 ;
  assign n11485 = \core_c_dec_MFLreg_E_reg[4]/P0001  & \core_dag_ilm2reg_L4_we_DO_reg[6]/NET0131  ;
  assign n11486 = \core_c_dec_MFLreg_E_reg[5]/P0001  & \core_dag_ilm2reg_L5_we_DO_reg[6]/NET0131  ;
  assign n11495 = ~n11485 & ~n11486 ;
  assign n11487 = \core_c_dec_MFLreg_E_reg[7]/P0001  & \core_dag_ilm2reg_L7_we_DO_reg[6]/NET0131  ;
  assign n11488 = \core_c_dec_MFMreg_E_reg[4]/P0001  & \core_dag_ilm2reg_M4_we_DO_reg[6]/NET0131  ;
  assign n11496 = ~n11487 & ~n11488 ;
  assign n11500 = n11495 & n11496 ;
  assign n11481 = \core_c_dec_MFLreg_E_reg[6]/P0001  & \core_dag_ilm2reg_L6_we_DO_reg[6]/NET0131  ;
  assign n11482 = \core_c_dec_MFMreg_E_reg[5]/P0001  & \core_dag_ilm2reg_M5_we_DO_reg[6]/NET0131  ;
  assign n11493 = ~n11481 & ~n11482 ;
  assign n11483 = \core_c_dec_MFMreg_E_reg[6]/P0001  & \core_dag_ilm2reg_M6_we_DO_reg[6]/NET0131  ;
  assign n11484 = \core_c_dec_MFMreg_E_reg[7]/P0001  & \core_dag_ilm2reg_M7_we_DO_reg[6]/NET0131  ;
  assign n11494 = ~n11483 & ~n11484 ;
  assign n11501 = n11493 & n11494 ;
  assign n11502 = n11500 & n11501 ;
  assign n11503 = n11499 & n11502 ;
  assign n11504 = n7128 & ~n11503 ;
  assign n11465 = \core_c_dec_MFLreg_E_reg[2]/P0001  & \core_dag_ilm1reg_L2_we_DO_reg[6]/NET0131  ;
  assign n11466 = \core_c_dec_MFMreg_E_reg[1]/P0001  & \core_dag_ilm1reg_M1_we_DO_reg[6]/NET0131  ;
  assign n11473 = ~n11465 & ~n11466 ;
  assign n11467 = \core_c_dec_MFMreg_E_reg[2]/P0001  & \core_dag_ilm1reg_M2_we_DO_reg[6]/NET0131  ;
  assign n11468 = \core_c_dec_MFMreg_E_reg[3]/P0001  & \core_dag_ilm1reg_M3_we_DO_reg[6]/NET0131  ;
  assign n11474 = ~n11467 & ~n11468 ;
  assign n11475 = n11473 & n11474 ;
  assign n11461 = \core_c_dec_MFLreg_E_reg[3]/P0001  & \core_dag_ilm1reg_L3_we_DO_reg[6]/NET0131  ;
  assign n11462 = \core_c_dec_MFMreg_E_reg[0]/P0001  & \core_dag_ilm1reg_M0_we_DO_reg[6]/NET0131  ;
  assign n11471 = ~n11461 & ~n11462 ;
  assign n11463 = \core_c_dec_MFLreg_E_reg[0]/P0001  & \core_dag_ilm1reg_L0_we_DO_reg[6]/NET0131  ;
  assign n11464 = \core_c_dec_MFLreg_E_reg[1]/P0001  & \core_dag_ilm1reg_L1_we_DO_reg[6]/NET0131  ;
  assign n11472 = ~n11463 & ~n11464 ;
  assign n11476 = n11471 & n11472 ;
  assign n11457 = \core_c_dec_MFIreg_E_reg[3]/P0001  & \core_dag_ilm1reg_I3_we_DO_reg[6]/NET0131  ;
  assign n11458 = \core_c_dec_MFIreg_E_reg[0]/P0001  & \core_dag_ilm1reg_I0_we_DO_reg[6]/NET0131  ;
  assign n11469 = ~n11457 & ~n11458 ;
  assign n11459 = \core_c_dec_MFIreg_E_reg[1]/P0001  & \core_dag_ilm1reg_I1_we_DO_reg[6]/NET0131  ;
  assign n11460 = \core_c_dec_MFIreg_E_reg[2]/P0001  & \core_dag_ilm1reg_I2_we_DO_reg[6]/NET0131  ;
  assign n11470 = ~n11459 & ~n11460 ;
  assign n11477 = n11469 & n11470 ;
  assign n11478 = n11476 & n11477 ;
  assign n11479 = n11475 & n11478 ;
  assign n11480 = n7068 & ~n11479 ;
  assign n11505 = \core_c_dec_MFTX1_E_reg/P0001  & \sport1_txctl_TX_reg[6]/P0001  ;
  assign n11506 = \core_c_dec_MFTX0_E_reg/P0001  & \sport0_txctl_TX_reg[6]/P0001  ;
  assign n11509 = ~n11505 & ~n11506 ;
  assign n11507 = \core_c_dec_MFRX1_E_reg/P0001  & \sport1_rxctl_RX_reg[6]/P0001  ;
  assign n11508 = \core_c_dec_MFRX0_E_reg/P0001  & \sport0_rxctl_RX_reg[6]/P0001  ;
  assign n11510 = ~n11507 & ~n11508 ;
  assign n11511 = n11509 & n11510 ;
  assign n11512 = n7119 & ~n11511 ;
  assign n11513 = ~n11480 & ~n11512 ;
  assign n11514 = ~n11504 & n11513 ;
  assign n11301 = ~\core_c_psq_MSTAT_reg_DO_reg[0]/P0002  & \core_eu_es_sht_es_reg_serwe_DO_reg[6]/P0001  ;
  assign n11302 = \core_c_psq_MSTAT_reg_DO_reg[0]/P0002  & \core_eu_es_sht_es_reg_seswe_DO_reg[6]/P0001  ;
  assign n11303 = ~n11301 & ~n11302 ;
  assign n11304 = \core_c_dec_MFSE_E_reg/P0001  & ~n11303 ;
  assign n11317 = ~n7169 & ~n11304 ;
  assign n11313 = ~\core_c_psq_MSTAT_reg_DO_reg[0]/P0002  & \core_eu_es_sht_es_reg_sr0rwe_DO_reg[6]/P0001  ;
  assign n11314 = \core_c_psq_MSTAT_reg_DO_reg[0]/P0002  & \core_eu_es_sht_es_reg_sr0swe_DO_reg[6]/P0001  ;
  assign n11315 = ~n11313 & ~n11314 ;
  assign n11316 = \core_c_dec_MFSR0_E_reg/P0001  & ~n11315 ;
  assign n11305 = ~\core_c_psq_MSTAT_reg_DO_reg[0]/P0002  & \core_eu_es_sht_es_reg_sirwe_DO_reg[6]/P0001  ;
  assign n11306 = \core_c_psq_MSTAT_reg_DO_reg[0]/P0002  & \core_eu_es_sht_es_reg_siswe_DO_reg[6]/P0001  ;
  assign n11307 = ~n11305 & ~n11306 ;
  assign n11308 = \core_c_dec_MFSI_E_reg/P0001  & ~n11307 ;
  assign n11309 = ~\core_c_psq_MSTAT_reg_DO_reg[0]/P0002  & \core_eu_es_sht_es_reg_sr1rwe_DO_reg[6]/P0001  ;
  assign n11310 = \core_c_psq_MSTAT_reg_DO_reg[0]/P0002  & \core_eu_es_sht_es_reg_sr1swe_DO_reg[6]/P0001  ;
  assign n11311 = ~n11309 & ~n11310 ;
  assign n11312 = \core_c_dec_MFSR1_E_reg/P0001  & ~n11311 ;
  assign n11318 = ~n11308 & ~n11312 ;
  assign n11319 = ~n11316 & n11318 ;
  assign n11320 = n11317 & n11319 ;
  assign n11321 = n7153 & ~n11320 ;
  assign n11446 = ~\core_c_psq_MSTAT_reg_DO_reg[0]/P0002  & \core_eu_em_mac_em_reg_mr1rwe_DO_reg[6]/P0001  ;
  assign n11447 = \core_c_psq_MSTAT_reg_DO_reg[0]/P0002  & \core_eu_em_mac_em_reg_mr1swe_DO_reg[6]/P0001  ;
  assign n11448 = ~n11446 & ~n11447 ;
  assign n11449 = \core_c_dec_MFMR1_E_reg/P0001  & ~n11448 ;
  assign n11438 = ~\core_c_psq_MSTAT_reg_DO_reg[0]/P0002  & \core_eu_em_mac_em_reg_mx0rwe_DO_reg[6]/P0001  ;
  assign n11439 = \core_c_psq_MSTAT_reg_DO_reg[0]/P0002  & \core_eu_em_mac_em_reg_mx0swe_DO_reg[6]/P0001  ;
  assign n11440 = ~n11438 & ~n11439 ;
  assign n11441 = \core_c_dec_MFMX0_E_reg/P0001  & ~n11440 ;
  assign n11442 = ~\core_c_psq_MSTAT_reg_DO_reg[0]/P0002  & \core_eu_em_mac_em_reg_mr0rwe_DO_reg[6]/P0001  ;
  assign n11443 = \core_c_psq_MSTAT_reg_DO_reg[0]/P0002  & \core_eu_em_mac_em_reg_mr0swe_DO_reg[6]/P0001  ;
  assign n11444 = ~n11442 & ~n11443 ;
  assign n11445 = \core_c_dec_MFMR0_E_reg/P0001  & ~n11444 ;
  assign n11452 = ~n11441 & ~n11445 ;
  assign n11453 = ~n11449 & n11452 ;
  assign n11422 = ~\core_c_psq_MSTAT_reg_DO_reg[0]/P0002  & \core_eu_em_mac_em_reg_mr2rwe_DO_reg[6]/P0001  ;
  assign n11423 = \core_c_psq_MSTAT_reg_DO_reg[0]/P0002  & \core_eu_em_mac_em_reg_mr2swe_DO_reg[6]/P0001  ;
  assign n11424 = ~n11422 & ~n11423 ;
  assign n11425 = \core_c_dec_MFMR2_E_reg/P0001  & ~n11424 ;
  assign n11426 = ~\core_c_psq_MSTAT_reg_DO_reg[0]/P0002  & \core_eu_em_mac_em_reg_mx1rwe_DO_reg[6]/P0001  ;
  assign n11427 = \core_c_psq_MSTAT_reg_DO_reg[0]/P0002  & \core_eu_em_mac_em_reg_mx1swe_DO_reg[6]/P0001  ;
  assign n11428 = ~n11426 & ~n11427 ;
  assign n11429 = \core_c_dec_MFMX1_E_reg/P0001  & ~n11428 ;
  assign n11450 = ~n11425 & ~n11429 ;
  assign n11430 = ~\core_c_psq_MSTAT_reg_DO_reg[0]/P0002  & \core_eu_em_mac_em_reg_my1rwe_DO_reg[6]/P0001  ;
  assign n11431 = \core_c_psq_MSTAT_reg_DO_reg[0]/P0002  & \core_eu_em_mac_em_reg_my1swe_DO_reg[6]/P0001  ;
  assign n11432 = ~n11430 & ~n11431 ;
  assign n11433 = \core_c_dec_MFMY1_E_reg/P0001  & ~n11432 ;
  assign n11434 = ~\core_c_psq_MSTAT_reg_DO_reg[0]/P0002  & \core_eu_em_mac_em_reg_my0rwe_DO_reg[6]/P0001  ;
  assign n11435 = \core_c_psq_MSTAT_reg_DO_reg[0]/P0002  & \core_eu_em_mac_em_reg_my0swe_DO_reg[6]/P0001  ;
  assign n11436 = ~n11434 & ~n11435 ;
  assign n11437 = \core_c_dec_MFMY0_E_reg/P0001  & ~n11436 ;
  assign n11451 = ~n11433 & ~n11437 ;
  assign n11454 = n11450 & n11451 ;
  assign n11455 = n11453 & n11454 ;
  assign n11456 = n7179 & ~n11455 ;
  assign n11515 = ~n11321 & ~n11456 ;
  assign n11516 = n11514 & n11515 ;
  assign n11517 = ~n11421 & n11516 ;
  assign n11518 = ~n11405 & n11517 ;
  assign n11519 = ~n11348 & n11518 ;
  assign n11520 = ~n11300 & n11519 ;
  assign n11521 = ~\emc_DMDoe_reg/NET0131  & ~n11520 ;
  assign n11522 = \emc_DMDoe_reg/NET0131  & \emc_DMDreg_reg[6]/P0001  ;
  assign n11523 = n7057 & ~n11522 ;
  assign n11524 = ~n11521 & n11523 ;
  assign n11525 = ~n11299 & ~n11524 ;
  assign n11526 = n6135 & ~n11525 ;
  assign n11527 = n8964 & ~n11526 ;
  assign n11528 = ~n11281 & n11527 ;
  assign n11529 = ~n11268 & ~n11528 ;
  assign n11530 = ~n11030 & n11529 ;
  assign n11581 = n6176 & ~n11280 ;
  assign n11571 = ~n6743 & ~n6779 ;
  assign n11572 = ~n6778 & n10920 ;
  assign n11573 = ~n6753 & ~n11572 ;
  assign n11574 = ~n11571 & ~n11573 ;
  assign n11575 = n11571 & n11573 ;
  assign n11576 = ~n11574 & ~n11575 ;
  assign n11577 = n8198 & n11576 ;
  assign n11566 = \core_dag_ilm2reg_I_reg[7]/NET0131  & ~n6642 ;
  assign n11567 = ~n6695 & ~n6731 ;
  assign n11568 = n6695 & n6731 ;
  assign n11569 = ~n11567 & ~n11568 ;
  assign n11570 = ~n8198 & n11569 ;
  assign n11578 = ~n11566 & ~n11570 ;
  assign n11579 = ~n11577 & n11578 ;
  assign n11580 = ~n6176 & ~n11579 ;
  assign n11582 = n6135 & ~n11580 ;
  assign n11583 = ~n11581 & n11582 ;
  assign n11552 = ~n6111 & n11025 ;
  assign n11534 = \core_dag_ilm2reg_I7_we_DO_reg[7]/NET0131  & n6972 ;
  assign n11535 = \core_dag_ilm2reg_I4_we_DO_reg[7]/NET0131  & n6976 ;
  assign n11538 = ~n11534 & ~n11535 ;
  assign n11536 = \core_dag_ilm2reg_I6_we_DO_reg[7]/NET0131  & n6974 ;
  assign n11537 = \core_dag_ilm2reg_I5_we_DO_reg[7]/NET0131  & n6970 ;
  assign n11539 = ~n11536 & ~n11537 ;
  assign n11540 = n11538 & n11539 ;
  assign n11541 = n4055 & ~n11540 ;
  assign n11542 = \core_dag_ilm2reg_I4_we_DO_reg[7]/NET0131  & n6958 ;
  assign n11543 = \core_dag_ilm2reg_I7_we_DO_reg[7]/NET0131  & n6960 ;
  assign n11546 = ~n11542 & ~n11543 ;
  assign n11544 = \core_dag_ilm2reg_I6_we_DO_reg[7]/NET0131  & n6962 ;
  assign n11545 = \core_dag_ilm2reg_I5_we_DO_reg[7]/NET0131  & n6964 ;
  assign n11547 = ~n11544 & ~n11545 ;
  assign n11548 = n11546 & n11547 ;
  assign n11549 = ~n11541 & n11548 ;
  assign n11550 = ~n6121 & ~n11549 ;
  assign n11551 = \core_c_dec_IR_reg[11]/NET0131  & n6956 ;
  assign n11553 = ~n11550 & ~n11551 ;
  assign n11554 = ~n11552 & n11553 ;
  assign n11555 = n5949 & ~n11554 ;
  assign n11556 = \core_dag_ilm1reg_DMA_pi_DO_reg[7]/NET0131  & ~n6934 ;
  assign n11532 = \core_dag_ilm1reg_STAC_pi_DO_reg[7]/NET0131  & n6988 ;
  assign n11533 = \idma_DCTL_reg[7]/NET0131  & n6926 ;
  assign n11557 = ~n11532 & ~n11533 ;
  assign n11558 = n6924 & n11557 ;
  assign n11559 = ~n11556 & n11558 ;
  assign n11560 = ~n11555 & n11559 ;
  assign n11531 = ~\bdma_BIAD_reg[7]/NET0131  & ~n6924 ;
  assign n11561 = ~n6176 & ~n11531 ;
  assign n11562 = ~n11560 & n11561 ;
  assign n11563 = n6176 & n10996 ;
  assign n11564 = ~n6135 & ~n11563 ;
  assign n11565 = ~n11562 & n11564 ;
  assign n11584 = ~n7005 & ~n11565 ;
  assign n11585 = ~n11583 & n11584 ;
  assign n11591 = ~n6176 & ~n11525 ;
  assign n11592 = ~n10955 & ~n11591 ;
  assign n11593 = ~n6135 & ~n11592 ;
  assign n11586 = n6176 & ~n11265 ;
  assign n11587 = ~n11025 & n11549 ;
  assign n11588 = ~n6176 & n11587 ;
  assign n11589 = ~n11586 & ~n11588 ;
  assign n11590 = n6135 & ~n11589 ;
  assign n11594 = n7005 & ~n11590 ;
  assign n11595 = ~n11593 & n11594 ;
  assign n11596 = ~n11585 & ~n11595 ;
  assign n11597 = ~n6176 & ~n10911 ;
  assign n11598 = ~n10344 & ~n11597 ;
  assign n11599 = n7005 & ~n11598 ;
  assign n11621 = ~n6111 & n10416 ;
  assign n11603 = \core_dag_ilm2reg_I7_we_DO_reg[8]/NET0131  & n6972 ;
  assign n11604 = \core_dag_ilm2reg_I4_we_DO_reg[8]/NET0131  & n6976 ;
  assign n11607 = ~n11603 & ~n11604 ;
  assign n11605 = \core_dag_ilm2reg_I6_we_DO_reg[8]/NET0131  & n6974 ;
  assign n11606 = \core_dag_ilm2reg_I5_we_DO_reg[8]/NET0131  & n6970 ;
  assign n11608 = ~n11605 & ~n11606 ;
  assign n11609 = n11607 & n11608 ;
  assign n11610 = n4055 & ~n11609 ;
  assign n11611 = \core_dag_ilm2reg_I7_we_DO_reg[8]/NET0131  & n6960 ;
  assign n11612 = \core_dag_ilm2reg_I4_we_DO_reg[8]/NET0131  & n6958 ;
  assign n11615 = ~n11611 & ~n11612 ;
  assign n11613 = \core_dag_ilm2reg_I6_we_DO_reg[8]/NET0131  & n6962 ;
  assign n11614 = \core_dag_ilm2reg_I5_we_DO_reg[8]/NET0131  & n6964 ;
  assign n11616 = ~n11613 & ~n11614 ;
  assign n11617 = n11615 & n11616 ;
  assign n11618 = ~n11610 & n11617 ;
  assign n11619 = ~n6121 & ~n11618 ;
  assign n11620 = \core_c_dec_IR_reg[12]/NET0131  & n6956 ;
  assign n11622 = ~n11619 & ~n11620 ;
  assign n11623 = ~n11621 & n11622 ;
  assign n11624 = n5949 & ~n11623 ;
  assign n11602 = \core_dag_ilm1reg_DMA_pi_DO_reg[8]/NET0131  & ~n6934 ;
  assign n11601 = \idma_DCTL_reg[8]/NET0131  & n6926 ;
  assign n11625 = \core_dag_ilm1reg_STAC_pi_DO_reg[8]/NET0131  & n6988 ;
  assign n11626 = ~n11601 & ~n11625 ;
  assign n11627 = ~n11602 & n11626 ;
  assign n11628 = ~n11624 & n11627 ;
  assign n11629 = n6924 & ~n11628 ;
  assign n11630 = \bdma_BIAD_reg[8]/NET0131  & ~n6924 ;
  assign n11631 = ~n11629 & ~n11630 ;
  assign n11632 = ~n6176 & ~n11631 ;
  assign n11600 = n6176 & n10386 ;
  assign n11633 = ~n7005 & ~n11600 ;
  assign n11634 = ~n11632 & n11633 ;
  assign n11635 = ~n11599 & ~n11634 ;
  assign n11636 = ~n6135 & ~n11635 ;
  assign n11637 = n6176 & ~n10638 ;
  assign n11638 = ~n10416 & n11618 ;
  assign n11639 = ~n6176 & n11638 ;
  assign n11640 = ~n11637 & ~n11639 ;
  assign n11641 = n7005 & ~n11640 ;
  assign n11648 = ~n6845 & ~n6873 ;
  assign n11649 = n6825 & ~n11648 ;
  assign n11650 = ~n6825 & n11648 ;
  assign n11651 = ~n11649 & ~n11650 ;
  assign n11652 = n8198 & n11651 ;
  assign n11643 = \core_dag_ilm2reg_I_reg[8]/NET0131  & ~n6635 ;
  assign n11644 = ~n6697 & ~n6841 ;
  assign n11645 = n6697 & n6841 ;
  assign n11646 = ~n11644 & ~n11645 ;
  assign n11647 = ~n8198 & n11646 ;
  assign n11653 = ~n11643 & ~n11647 ;
  assign n11654 = ~n11652 & n11653 ;
  assign n11655 = ~n6176 & ~n11654 ;
  assign n11642 = n6176 & ~n10663 ;
  assign n11656 = ~n7005 & ~n11642 ;
  assign n11657 = ~n11655 & n11656 ;
  assign n11658 = ~n11641 & ~n11657 ;
  assign n11659 = n6135 & ~n11658 ;
  assign n11660 = ~n11636 & ~n11659 ;
  assign n11680 = ~n6135 & n9752 ;
  assign n11681 = n6135 & ~n10289 ;
  assign n11682 = n6176 & ~n11681 ;
  assign n11683 = ~n11680 & n11682 ;
  assign n11661 = n7863 & n10069 ;
  assign n11662 = \core_dag_ilm2reg_I5_we_DO_reg[9]/NET0131  & n6970 ;
  assign n11663 = \core_dag_ilm2reg_I7_we_DO_reg[9]/NET0131  & n6972 ;
  assign n11666 = ~n11662 & ~n11663 ;
  assign n11664 = \core_dag_ilm2reg_I6_we_DO_reg[9]/NET0131  & n6974 ;
  assign n11665 = \core_dag_ilm2reg_I4_we_DO_reg[9]/NET0131  & n6976 ;
  assign n11667 = ~n11664 & ~n11665 ;
  assign n11668 = n11666 & n11667 ;
  assign n11669 = n4055 & ~n11668 ;
  assign n11670 = \core_dag_ilm2reg_I4_we_DO_reg[9]/NET0131  & n6958 ;
  assign n11671 = \core_dag_ilm2reg_I7_we_DO_reg[9]/NET0131  & n6960 ;
  assign n11674 = ~n11670 & ~n11671 ;
  assign n11672 = \core_dag_ilm2reg_I6_we_DO_reg[9]/NET0131  & n6962 ;
  assign n11673 = \core_dag_ilm2reg_I5_we_DO_reg[9]/NET0131  & n6964 ;
  assign n11675 = ~n11672 & ~n11673 ;
  assign n11676 = n11674 & n11675 ;
  assign n11677 = ~n11669 & n11676 ;
  assign n11678 = ~n9735 & n11677 ;
  assign n11679 = n8153 & ~n11678 ;
  assign n11684 = ~n11661 & ~n11679 ;
  assign n11685 = ~n11683 & n11684 ;
  assign n11686 = n7005 & ~n11685 ;
  assign n11691 = ~n6121 & ~n11677 ;
  assign n11690 = ~n6111 & n9735 ;
  assign n11692 = \core_c_dec_IR_reg[13]/NET0131  & n6956 ;
  assign n11693 = ~n11690 & ~n11692 ;
  assign n11694 = ~n11691 & n11693 ;
  assign n11695 = n5949 & ~n11694 ;
  assign n11689 = \core_dag_ilm1reg_DMA_pi_DO_reg[9]/NET0131  & ~n6934 ;
  assign n11687 = \core_dag_ilm1reg_STAC_pi_DO_reg[9]/NET0131  & n6988 ;
  assign n11688 = \idma_DCTL_reg[9]/NET0131  & n6926 ;
  assign n11696 = ~n11687 & ~n11688 ;
  assign n11697 = ~n11689 & n11696 ;
  assign n11698 = ~n11695 & n11697 ;
  assign n11699 = n6924 & ~n11698 ;
  assign n11700 = \bdma_BIAD_reg[9]/NET0131  & ~n6924 ;
  assign n11701 = ~n6176 & ~n11700 ;
  assign n11702 = ~n11699 & n11701 ;
  assign n11703 = n6176 & ~n9788 ;
  assign n11704 = ~n6135 & ~n11703 ;
  assign n11705 = ~n11702 & n11704 ;
  assign n11714 = ~n6698 & ~n6703 ;
  assign n11715 = n6826 & ~n11714 ;
  assign n11716 = ~n6826 & n11714 ;
  assign n11717 = ~n11715 & ~n11716 ;
  assign n11718 = ~n8198 & n11717 ;
  assign n11706 = \core_dag_ilm2reg_I_reg[9]/NET0131  & ~n6630 ;
  assign n11707 = ~n6838 & ~n6872 ;
  assign n11708 = ~n6825 & ~n6845 ;
  assign n11709 = ~n6873 & ~n11708 ;
  assign n11710 = n11707 & ~n11709 ;
  assign n11711 = ~n11707 & n11709 ;
  assign n11712 = ~n11710 & ~n11711 ;
  assign n11713 = n8198 & n11712 ;
  assign n11719 = ~n11706 & ~n11713 ;
  assign n11720 = ~n11718 & n11719 ;
  assign n11721 = ~n6176 & n11720 ;
  assign n11722 = n6135 & ~n11721 ;
  assign n11723 = ~n10303 & n11722 ;
  assign n11724 = ~n11705 & ~n11723 ;
  assign n11725 = ~n7005 & ~n11724 ;
  assign n11726 = ~n11686 & ~n11725 ;
  assign n11731 = ~n8835 & n11660 ;
  assign n11732 = ~n11726 & n11731 ;
  assign n11728 = ~n10916 & ~n11530 ;
  assign n11729 = ~n11596 & n11728 ;
  assign n11727 = ~n9440 & ~n9513 ;
  assign n11730 = ~n8230 & n11727 ;
  assign n11733 = n11729 & n11730 ;
  assign n11734 = n11732 & n11733 ;
  assign n11735 = ~n9513 & ~n11734 ;
  assign n11739 = \memc_Dread_E_reg/NET0131  & n4117 ;
  assign n11740 = ~\core_c_dec_Long_Cg_reg/P0001  & ~\core_c_dec_Prderr_Cg_reg/NET0131  ;
  assign n11741 = n5053 & n11740 ;
  assign n11742 = ~n4117 & n11741 ;
  assign n11743 = ~\core_c_dec_IR_reg[15]/NET0131  & n6120 ;
  assign n11744 = ~\core_c_dec_IR_reg[19]/NET0131  & n6108 ;
  assign n11745 = n6026 & n6955 ;
  assign n11746 = ~n6023 & ~n11745 ;
  assign n11747 = ~n11744 & n11746 ;
  assign n11748 = ~n11743 & n11747 ;
  assign n11749 = n11742 & ~n11748 ;
  assign n11750 = n5948 & n11749 ;
  assign n11751 = ~n11739 & ~n11750 ;
  assign n11752 = \idma_DCTL_reg[14]/NET0131  & \idma_RDcyc_reg/NET0131  ;
  assign n11753 = n5068 & n11752 ;
  assign n11754 = ~n4050 & ~n5968 ;
  assign n11755 = ~n11753 & n11754 ;
  assign n11756 = ~n6922 & n11755 ;
  assign n11757 = ~n5718 & ~n11756 ;
  assign n11758 = n11751 & ~n11757 ;
  assign n11736 = \memc_Dwrite_C_reg/NET0131  & n5950 ;
  assign n11737 = ~n5950 & n6932 ;
  assign n11738 = ~n11736 & ~n11737 ;
  assign n11759 = ~n5966 & ~n5970 ;
  assign n11760 = ~n5718 & ~n11759 ;
  assign n11761 = \idma_WRcyc_reg/NET0131  & ~n5718 ;
  assign n11762 = n6925 & n11761 ;
  assign n11763 = ~n6918 & ~n11762 ;
  assign n11764 = ~n11760 & n11763 ;
  assign n11765 = n11738 & n11764 ;
  assign n11766 = n11758 & n11765 ;
  assign n11767 = n11735 & ~n11766 ;
  assign n11769 = ~n4097 & ~n11759 ;
  assign n11770 = n11763 & ~n11769 ;
  assign n11771 = ~n7602 & n11770 ;
  assign n11776 = \bdma_BRdataBUF_reg[0]/P0001  & n6918 ;
  assign n11768 = \idma_DTMP_H_reg[0]/P0001  & n11762 ;
  assign n11772 = ~n4097 & n5966 ;
  assign n11773 = \sport1_rxctl_RX_reg[0]/P0001  & n11772 ;
  assign n11774 = ~n4097 & n5970 ;
  assign n11775 = \sport0_rxctl_RX_reg[0]/P0001  & n11774 ;
  assign n11777 = ~n11773 & ~n11775 ;
  assign n11778 = ~n11768 & n11777 ;
  assign n11779 = ~n11776 & n11778 ;
  assign n11780 = ~n11771 & n11779 ;
  assign n11782 = ~n7854 & n11770 ;
  assign n11785 = \bdma_BRdataBUF_reg[10]/P0001  & n6918 ;
  assign n11781 = \idma_DTMP_H_reg[10]/P0001  & n11762 ;
  assign n11783 = \sport0_rxctl_RX_reg[10]/P0001  & n11774 ;
  assign n11784 = \sport1_rxctl_RX_reg[10]/P0001  & n11772 ;
  assign n11786 = ~n11783 & ~n11784 ;
  assign n11787 = ~n11781 & n11786 ;
  assign n11788 = ~n11785 & n11787 ;
  assign n11789 = ~n11782 & n11788 ;
  assign n11791 = ~n8455 & n11770 ;
  assign n11794 = \bdma_BRdataBUF_reg[11]/P0001  & n6918 ;
  assign n11790 = \idma_DTMP_H_reg[11]/P0001  & n11762 ;
  assign n11792 = \sport1_rxctl_RX_reg[11]/P0001  & n11772 ;
  assign n11793 = \sport0_rxctl_RX_reg[11]/P0001  & n11774 ;
  assign n11795 = ~n11792 & ~n11793 ;
  assign n11796 = ~n11790 & n11795 ;
  assign n11797 = ~n11794 & n11796 ;
  assign n11798 = ~n11791 & n11797 ;
  assign n11800 = ~n9173 & n11770 ;
  assign n11803 = \bdma_BRdataBUF_reg[12]/P0001  & n6918 ;
  assign n11799 = \idma_DTMP_H_reg[12]/P0001  & n11762 ;
  assign n11801 = \sport0_rxctl_RX_reg[12]/P0001  & n11774 ;
  assign n11802 = \sport1_rxctl_RX_reg[12]/P0001  & n11772 ;
  assign n11804 = ~n11801 & ~n11802 ;
  assign n11805 = ~n11799 & n11804 ;
  assign n11806 = ~n11803 & n11805 ;
  assign n11807 = ~n11800 & n11806 ;
  assign n11809 = ~n7335 & n11770 ;
  assign n11812 = \bdma_BRdataBUF_reg[13]/P0001  & n6918 ;
  assign n11808 = \idma_DTMP_H_reg[13]/P0001  & n11762 ;
  assign n11810 = \sport0_rxctl_RX_reg[13]/P0001  & n11774 ;
  assign n11811 = \sport1_rxctl_RX_reg[13]/P0001  & n11772 ;
  assign n11813 = ~n11810 & ~n11811 ;
  assign n11814 = ~n11808 & n11813 ;
  assign n11815 = ~n11812 & n11814 ;
  assign n11816 = ~n11809 & n11815 ;
  assign n11818 = \regout_STD_C_reg[14]/P0001  & n6988 ;
  assign n11923 = \sport0_regs_FSDIVreg_DO_reg[14]/NET0131  & n7259 ;
  assign n11924 = PM_bdry_sel_pad & n7522 ;
  assign n11935 = ~n11923 & ~n11924 ;
  assign n11925 = \memc_usysr_DO_reg[14]/NET0131  & n7301 ;
  assign n11926 = \sport0_regs_SCLKDIVreg_DO_reg[14]/NET0131  & n7256 ;
  assign n11936 = ~n11925 & ~n11926 ;
  assign n11937 = n11935 & n11936 ;
  assign n11919 = \tm_tpr_reg_DO_reg[14]/NET0131  & n7293 ;
  assign n11920 = \pio_pmask_reg_DO_reg[10]/NET0131  & n7297 ;
  assign n11933 = ~n11919 & ~n11920 ;
  assign n11921 = \sport1_regs_SCLKDIVreg_DO_reg[14]/NET0131  & n7247 ;
  assign n11922 = \sport1_regs_FSDIVreg_DO_reg[14]/NET0131  & n7273 ;
  assign n11934 = ~n11921 & ~n11922 ;
  assign n11938 = n11933 & n11934 ;
  assign n11915 = \PIO_oe[10]_pad  & n7244 ;
  assign n11916 = \tm_TCR_TMP_reg[14]/NET0131  & n7289 ;
  assign n11931 = ~n11915 & ~n11916 ;
  assign n11917 = \sport0_regs_AUTO_a_reg[14]/NET0131  & n7295 ;
  assign n11918 = \ISCLK1_pad  & n7281 ;
  assign n11932 = ~n11917 & ~n11918 ;
  assign n11939 = n11931 & n11932 ;
  assign n11943 = n11938 & n11939 ;
  assign n11944 = n11937 & n11943 ;
  assign n11911 = \bdma_BCTL_reg[14]/NET0131  & n7230 ;
  assign n11910 = \ISCLK0_pad  & n7249 ;
  assign n11912 = \clkc_ckr_reg_DO_reg[14]/NET0131  & n7239 ;
  assign n11929 = ~n11910 & ~n11912 ;
  assign n11913 = \idma_DCTL_reg[14]/NET0131  & n7299 ;
  assign n11914 = \emc_WSCRreg_DO_reg[14]/NET0131  & n7251 ;
  assign n11930 = ~n11913 & ~n11914 ;
  assign n11940 = n11929 & n11930 ;
  assign n11927 = ~n7689 & ~n7710 ;
  assign n11908 = \PIO_out[10]_pad  & n7291 ;
  assign n11909 = \pio_PINT_reg[10]/NET0131  & n7271 ;
  assign n11928 = ~n11908 & ~n11909 ;
  assign n11941 = n11927 & n11928 ;
  assign n11942 = n11940 & n11941 ;
  assign n11945 = ~n11911 & n11942 ;
  assign n11946 = n11944 & n11945 ;
  assign n11947 = \memc_ldSREG_E_reg/NET0131  & ~n11946 ;
  assign n11819 = ~\core_c_psq_MSTAT_reg_DO_reg[0]/P0002  & \core_eu_ea_alu_ea_reg_ax0rwe_DO_reg[14]/P0001  ;
  assign n11820 = \core_c_psq_MSTAT_reg_DO_reg[0]/P0002  & \core_eu_ea_alu_ea_reg_ax0swe_DO_reg[14]/P0001  ;
  assign n11821 = ~n11819 & ~n11820 ;
  assign n11822 = \core_c_dec_MFAX0_E_reg/P0001  & ~n11821 ;
  assign n11823 = ~\core_c_psq_MSTAT_reg_DO_reg[0]/P0002  & \core_eu_ea_alu_ea_reg_ax1rwe_DO_reg[14]/P0001  ;
  assign n11824 = \core_c_psq_MSTAT_reg_DO_reg[0]/P0002  & \core_eu_ea_alu_ea_reg_ax1swe_DO_reg[14]/P0001  ;
  assign n11825 = ~n11823 & ~n11824 ;
  assign n11826 = \core_c_dec_MFAX1_E_reg/P0001  & ~n11825 ;
  assign n11839 = ~n11822 & ~n11826 ;
  assign n11835 = ~\core_c_psq_MSTAT_reg_DO_reg[0]/P0002  & \core_eu_ea_alu_ea_reg_arrwe_DO_reg[14]/P0001  ;
  assign n11836 = \core_c_psq_MSTAT_reg_DO_reg[0]/P0002  & \core_eu_ea_alu_ea_reg_arswe_DO_reg[14]/P0001  ;
  assign n11837 = ~n11835 & ~n11836 ;
  assign n11838 = \core_c_dec_MFAR_E_reg/P0001  & ~n11837 ;
  assign n11827 = ~\core_c_psq_MSTAT_reg_DO_reg[0]/P0002  & \core_eu_ea_alu_ea_reg_ay0rwe_DO_reg[14]/P0001  ;
  assign n11828 = \core_c_psq_MSTAT_reg_DO_reg[0]/P0002  & \core_eu_ea_alu_ea_reg_ay0swe_DO_reg[14]/P0001  ;
  assign n11829 = ~n11827 & ~n11828 ;
  assign n11830 = \core_c_dec_MFAY0_E_reg/P0001  & ~n11829 ;
  assign n11831 = ~\core_c_psq_MSTAT_reg_DO_reg[0]/P0002  & \core_eu_ea_alu_ea_reg_ay1rwe_DO_reg[14]/P0001  ;
  assign n11832 = \core_c_psq_MSTAT_reg_DO_reg[0]/P0002  & \core_eu_ea_alu_ea_reg_ay1swe_DO_reg[14]/P0001  ;
  assign n11833 = ~n11831 & ~n11832 ;
  assign n11834 = \core_c_dec_MFAY1_E_reg/P0001  & ~n11833 ;
  assign n11840 = ~n11830 & ~n11834 ;
  assign n11841 = ~n11838 & n11840 ;
  assign n11842 = n11839 & n11841 ;
  assign n11843 = n7093 & ~n11842 ;
  assign n11905 = n7068 & ~n7078 ;
  assign n11906 = n7128 & ~n7137 ;
  assign n11907 = ~n11905 & ~n11906 ;
  assign n11891 = \core_c_dec_MFTX1_E_reg/P0001  & \sport1_txctl_TX_reg[14]/P0001  ;
  assign n11892 = \core_c_dec_MFTX0_E_reg/P0001  & \sport0_txctl_TX_reg[14]/P0001  ;
  assign n11895 = ~n11891 & ~n11892 ;
  assign n11893 = \core_c_dec_MFRX1_E_reg/P0001  & \sport1_rxctl_RX_reg[14]/P0001  ;
  assign n11894 = \core_c_dec_MFRX0_E_reg/P0001  & \sport0_rxctl_RX_reg[14]/P0001  ;
  assign n11896 = ~n11893 & ~n11894 ;
  assign n11897 = n11895 & n11896 ;
  assign n11898 = n7119 & ~n11897 ;
  assign n11901 = \core_c_dec_IRE_reg[18]/NET0131  & \core_c_dec_imm16_E_reg/P0001  ;
  assign n11899 = \core_c_dec_IRE_reg[17]/NET0131  & \core_c_dec_imm14_E_reg/P0001  ;
  assign n11900 = \core_c_dec_MFIDR_E_reg/P0001  & \sice_idr1_reg_DO_reg[2]/P0001  ;
  assign n11902 = ~n11899 & ~n11900 ;
  assign n11903 = ~n11901 & n11902 ;
  assign n11904 = n7215 & ~n11903 ;
  assign n11948 = ~n11898 & ~n11904 ;
  assign n11949 = n11907 & n11948 ;
  assign n11950 = ~n11843 & n11949 ;
  assign n11852 = ~\core_c_psq_MSTAT_reg_DO_reg[0]/P0002  & \core_eu_es_sht_es_reg_sr1rwe_DO_reg[14]/P0001  ;
  assign n11853 = \core_c_psq_MSTAT_reg_DO_reg[0]/P0002  & \core_eu_es_sht_es_reg_sr1swe_DO_reg[14]/P0001  ;
  assign n11854 = ~n11852 & ~n11853 ;
  assign n11855 = \core_c_dec_MFSR1_E_reg/P0001  & ~n11854 ;
  assign n11844 = ~\core_c_psq_MSTAT_reg_DO_reg[0]/P0002  & \core_eu_es_sht_es_reg_sr0rwe_DO_reg[14]/P0001  ;
  assign n11845 = \core_c_psq_MSTAT_reg_DO_reg[0]/P0002  & \core_eu_es_sht_es_reg_sr0swe_DO_reg[14]/P0001  ;
  assign n11846 = ~n11844 & ~n11845 ;
  assign n11847 = \core_c_dec_MFSR0_E_reg/P0001  & ~n11846 ;
  assign n11848 = ~\core_c_psq_MSTAT_reg_DO_reg[0]/P0002  & \core_eu_es_sht_es_reg_sirwe_DO_reg[14]/P0001  ;
  assign n11849 = \core_c_psq_MSTAT_reg_DO_reg[0]/P0002  & \core_eu_es_sht_es_reg_siswe_DO_reg[14]/P0001  ;
  assign n11850 = ~n11848 & ~n11849 ;
  assign n11851 = \core_c_dec_MFSI_E_reg/P0001  & ~n11850 ;
  assign n11856 = ~n11847 & ~n11851 ;
  assign n11857 = ~n11855 & n11856 ;
  assign n11858 = n7174 & n11857 ;
  assign n11859 = n7153 & ~n11858 ;
  assign n11880 = ~\core_c_psq_MSTAT_reg_DO_reg[0]/P0002  & \core_eu_em_mac_em_reg_mr1rwe_DO_reg[14]/P0001  ;
  assign n11881 = \core_c_psq_MSTAT_reg_DO_reg[0]/P0002  & \core_eu_em_mac_em_reg_mr1swe_DO_reg[14]/P0001  ;
  assign n11882 = ~n11880 & ~n11881 ;
  assign n11883 = \core_c_dec_MFMR1_E_reg/P0001  & ~n11882 ;
  assign n11872 = ~\core_c_psq_MSTAT_reg_DO_reg[0]/P0002  & \core_eu_em_mac_em_reg_mx1rwe_DO_reg[14]/P0001  ;
  assign n11873 = \core_c_psq_MSTAT_reg_DO_reg[0]/P0002  & \core_eu_em_mac_em_reg_mx1swe_DO_reg[14]/P0001  ;
  assign n11874 = ~n11872 & ~n11873 ;
  assign n11875 = \core_c_dec_MFMX1_E_reg/P0001  & ~n11874 ;
  assign n11876 = ~\core_c_psq_MSTAT_reg_DO_reg[0]/P0002  & \core_eu_em_mac_em_reg_mr0rwe_DO_reg[14]/P0001  ;
  assign n11877 = \core_c_psq_MSTAT_reg_DO_reg[0]/P0002  & \core_eu_em_mac_em_reg_mr0swe_DO_reg[14]/P0001  ;
  assign n11878 = ~n11876 & ~n11877 ;
  assign n11879 = \core_c_dec_MFMR0_E_reg/P0001  & ~n11878 ;
  assign n11886 = ~n11875 & ~n11879 ;
  assign n11887 = ~n11883 & n11886 ;
  assign n11860 = ~\core_c_psq_MSTAT_reg_DO_reg[0]/P0002  & \core_eu_em_mac_em_reg_my0rwe_DO_reg[14]/P0001  ;
  assign n11861 = \core_c_psq_MSTAT_reg_DO_reg[0]/P0002  & \core_eu_em_mac_em_reg_my0swe_DO_reg[14]/P0001  ;
  assign n11862 = ~n11860 & ~n11861 ;
  assign n11863 = \core_c_dec_MFMY0_E_reg/P0001  & ~n11862 ;
  assign n11884 = ~n7207 & ~n11863 ;
  assign n11864 = ~\core_c_psq_MSTAT_reg_DO_reg[0]/P0002  & \core_eu_em_mac_em_reg_my1rwe_DO_reg[14]/P0001  ;
  assign n11865 = \core_c_psq_MSTAT_reg_DO_reg[0]/P0002  & \core_eu_em_mac_em_reg_my1swe_DO_reg[14]/P0001  ;
  assign n11866 = ~n11864 & ~n11865 ;
  assign n11867 = \core_c_dec_MFMY1_E_reg/P0001  & ~n11866 ;
  assign n11868 = ~\core_c_psq_MSTAT_reg_DO_reg[0]/P0002  & \core_eu_em_mac_em_reg_mx0rwe_DO_reg[14]/P0001  ;
  assign n11869 = \core_c_psq_MSTAT_reg_DO_reg[0]/P0002  & \core_eu_em_mac_em_reg_mx0swe_DO_reg[14]/P0001  ;
  assign n11870 = ~n11868 & ~n11869 ;
  assign n11871 = \core_c_dec_MFMX0_E_reg/P0001  & ~n11870 ;
  assign n11885 = ~n11867 & ~n11871 ;
  assign n11888 = n11884 & n11885 ;
  assign n11889 = n11887 & n11888 ;
  assign n11890 = n7179 & ~n11889 ;
  assign n11951 = ~n11859 & ~n11890 ;
  assign n11952 = n11950 & n11951 ;
  assign n11953 = ~n11947 & n11952 ;
  assign n11954 = ~n11818 & n11953 ;
  assign n11955 = n11770 & ~n11954 ;
  assign n11958 = \bdma_BRdataBUF_reg[14]/P0001  & n6918 ;
  assign n11817 = \idma_DTMP_H_reg[14]/P0001  & n11762 ;
  assign n11956 = \sport0_rxctl_RX_reg[14]/P0001  & n11774 ;
  assign n11957 = \sport1_rxctl_RX_reg[14]/P0001  & n11772 ;
  assign n11959 = ~n11956 & ~n11957 ;
  assign n11960 = ~n11817 & n11959 ;
  assign n11961 = ~n11958 & n11960 ;
  assign n11962 = ~n11955 & n11961 ;
  assign n11964 = \regout_STD_C_reg[15]/P0001  & n6988 ;
  assign n12069 = \PIO_out[11]_pad  & n7291 ;
  assign n12067 = \tm_TCR_TMP_reg[15]/NET0131  & n7289 ;
  assign n12068 = \clkc_ckr_reg_DO_reg[15]/NET0131  & n7239 ;
  assign n12078 = ~n12067 & ~n12068 ;
  assign n12079 = ~n12069 & n12078 ;
  assign n12063 = \pio_pmask_reg_DO_reg[11]/NET0131  & n7297 ;
  assign n12064 = \sice_ICYC_en_reg/NET0131  & n7522 ;
  assign n12076 = ~n12063 & ~n12064 ;
  assign n12065 = \sport1_regs_FSDIVreg_DO_reg[15]/NET0131  & n7273 ;
  assign n12066 = \memc_usysr_DO_reg[15]/NET0131  & n7301 ;
  assign n12077 = ~n12065 & ~n12066 ;
  assign n12080 = n12076 & n12077 ;
  assign n12059 = \sport0_regs_SCTLreg_DO_reg[15]/NET0131  & n7249 ;
  assign n12060 = \sport1_regs_SCLKDIVreg_DO_reg[15]/NET0131  & n7247 ;
  assign n12074 = ~n12059 & ~n12060 ;
  assign n12061 = \pio_PINT_reg[11]/NET0131  & n7271 ;
  assign n12062 = \sport0_regs_SCLKDIVreg_DO_reg[15]/NET0131  & n7256 ;
  assign n12075 = ~n12061 & ~n12062 ;
  assign n12081 = n12074 & n12075 ;
  assign n12085 = n12080 & n12081 ;
  assign n12086 = n12079 & n12085 ;
  assign n12053 = \bdma_BCTL_reg[15]/NET0131  & n7230 ;
  assign n12055 = \tm_tpr_reg_DO_reg[15]/NET0131  & n7293 ;
  assign n12056 = \sport0_regs_AUTO_a_reg[15]/NET0131  & n7295 ;
  assign n12072 = ~n12055 & ~n12056 ;
  assign n12057 = \sport0_regs_FSDIVreg_DO_reg[15]/NET0131  & n7259 ;
  assign n12058 = \sport0_regs_MWORDreg_DO_reg[10]/NET0131  & n7276 ;
  assign n12073 = ~n12057 & ~n12058 ;
  assign n12082 = n12072 & n12073 ;
  assign n12050 = \tm_tsr_reg_DO_reg[8]/NET0131  & n7540 ;
  assign n12051 = \sport1_regs_MWORDreg_DO_reg[10]/NET0131  & n7263 ;
  assign n12070 = ~n12050 & ~n12051 ;
  assign n12052 = \sport1_regs_SCTLreg_DO_reg[15]/NET0131  & n7281 ;
  assign n12054 = \PIO_oe[11]_pad  & n7244 ;
  assign n12071 = ~n12052 & ~n12054 ;
  assign n12083 = n12070 & n12071 ;
  assign n12084 = n12082 & n12083 ;
  assign n12087 = ~n12053 & n12084 ;
  assign n12088 = n12086 & n12087 ;
  assign n12089 = \memc_ldSREG_E_reg/NET0131  & ~n12088 ;
  assign n11965 = ~\core_c_psq_MSTAT_reg_DO_reg[0]/P0002  & \core_eu_ea_alu_ea_reg_ax0rwe_DO_reg[15]/P0001  ;
  assign n11966 = \core_c_psq_MSTAT_reg_DO_reg[0]/P0002  & \core_eu_ea_alu_ea_reg_ax0swe_DO_reg[15]/P0001  ;
  assign n11967 = ~n11965 & ~n11966 ;
  assign n11968 = \core_c_dec_MFAX0_E_reg/P0001  & ~n11967 ;
  assign n11969 = ~\core_c_psq_MSTAT_reg_DO_reg[0]/P0002  & \core_eu_ea_alu_ea_reg_ax1rwe_DO_reg[15]/P0001  ;
  assign n11970 = \core_c_psq_MSTAT_reg_DO_reg[0]/P0002  & \core_eu_ea_alu_ea_reg_ax1swe_DO_reg[15]/P0001  ;
  assign n11971 = ~n11969 & ~n11970 ;
  assign n11972 = \core_c_dec_MFAX1_E_reg/P0001  & ~n11971 ;
  assign n11985 = ~n11968 & ~n11972 ;
  assign n11981 = ~\core_c_psq_MSTAT_reg_DO_reg[0]/P0002  & \core_eu_ea_alu_ea_reg_arrwe_DO_reg[15]/P0001  ;
  assign n11982 = \core_c_psq_MSTAT_reg_DO_reg[0]/P0002  & \core_eu_ea_alu_ea_reg_arswe_DO_reg[15]/P0001  ;
  assign n11983 = ~n11981 & ~n11982 ;
  assign n11984 = \core_c_dec_MFAR_E_reg/P0001  & ~n11983 ;
  assign n11973 = ~\core_c_psq_MSTAT_reg_DO_reg[0]/P0002  & \core_eu_ea_alu_ea_reg_ay0rwe_DO_reg[15]/P0001  ;
  assign n11974 = \core_c_psq_MSTAT_reg_DO_reg[0]/P0002  & \core_eu_ea_alu_ea_reg_ay0swe_DO_reg[15]/P0001  ;
  assign n11975 = ~n11973 & ~n11974 ;
  assign n11976 = \core_c_dec_MFAY0_E_reg/P0001  & ~n11975 ;
  assign n11977 = ~\core_c_psq_MSTAT_reg_DO_reg[0]/P0002  & \core_eu_ea_alu_ea_reg_ay1rwe_DO_reg[15]/P0001  ;
  assign n11978 = \core_c_psq_MSTAT_reg_DO_reg[0]/P0002  & \core_eu_ea_alu_ea_reg_ay1swe_DO_reg[15]/P0001  ;
  assign n11979 = ~n11977 & ~n11978 ;
  assign n11980 = \core_c_dec_MFAY1_E_reg/P0001  & ~n11979 ;
  assign n11986 = ~n11976 & ~n11980 ;
  assign n11987 = ~n11984 & n11986 ;
  assign n11988 = n11985 & n11987 ;
  assign n11989 = n7093 & ~n11988 ;
  assign n12037 = \core_c_dec_MFTX1_E_reg/P0001  & \sport1_txctl_TX_reg[15]/P0001  ;
  assign n12038 = \core_c_dec_MFRX1_E_reg/P0001  & \sport1_rxctl_RX_reg[15]/P0001  ;
  assign n12041 = ~n12037 & ~n12038 ;
  assign n12039 = \core_c_dec_MFTX0_E_reg/P0001  & \sport0_txctl_TX_reg[15]/P0001  ;
  assign n12040 = \core_c_dec_MFRX0_E_reg/P0001  & \sport0_rxctl_RX_reg[15]/P0001  ;
  assign n12042 = ~n12039 & ~n12040 ;
  assign n12043 = n12041 & n12042 ;
  assign n12044 = n7119 & ~n12043 ;
  assign n12046 = \core_c_dec_MFIDR_E_reg/P0001  & \sice_idr1_reg_DO_reg[3]/P0001  ;
  assign n12045 = \core_c_dec_IRE_reg[19]/NET0131  & \core_c_dec_imm16_E_reg/P0001  ;
  assign n12047 = ~n11899 & ~n12045 ;
  assign n12048 = ~n12046 & n12047 ;
  assign n12049 = n7215 & ~n12048 ;
  assign n12090 = ~n12044 & ~n12049 ;
  assign n12091 = n11907 & n12090 ;
  assign n12092 = ~n11989 & n12091 ;
  assign n11998 = ~\core_c_psq_MSTAT_reg_DO_reg[0]/P0002  & \core_eu_es_sht_es_reg_sr1rwe_DO_reg[15]/P0001  ;
  assign n11999 = \core_c_psq_MSTAT_reg_DO_reg[0]/P0002  & \core_eu_es_sht_es_reg_sr1swe_DO_reg[15]/P0001  ;
  assign n12000 = ~n11998 & ~n11999 ;
  assign n12001 = \core_c_dec_MFSR1_E_reg/P0001  & ~n12000 ;
  assign n11990 = ~\core_c_psq_MSTAT_reg_DO_reg[0]/P0002  & \core_eu_es_sht_es_reg_sr0rwe_DO_reg[15]/P0001  ;
  assign n11991 = \core_c_psq_MSTAT_reg_DO_reg[0]/P0002  & \core_eu_es_sht_es_reg_sr0swe_DO_reg[15]/P0001  ;
  assign n11992 = ~n11990 & ~n11991 ;
  assign n11993 = \core_c_dec_MFSR0_E_reg/P0001  & ~n11992 ;
  assign n11994 = ~\core_c_psq_MSTAT_reg_DO_reg[0]/P0002  & \core_eu_es_sht_es_reg_sirwe_DO_reg[15]/P0001  ;
  assign n11995 = \core_c_psq_MSTAT_reg_DO_reg[0]/P0002  & \core_eu_es_sht_es_reg_siswe_DO_reg[15]/P0001  ;
  assign n11996 = ~n11994 & ~n11995 ;
  assign n11997 = \core_c_dec_MFSI_E_reg/P0001  & ~n11996 ;
  assign n12002 = ~n11993 & ~n11997 ;
  assign n12003 = ~n12001 & n12002 ;
  assign n12004 = n7174 & n12003 ;
  assign n12005 = n7153 & ~n12004 ;
  assign n12026 = ~\core_c_psq_MSTAT_reg_DO_reg[0]/P0002  & \core_eu_em_mac_em_reg_mr1rwe_DO_reg[15]/P0001  ;
  assign n12027 = \core_c_psq_MSTAT_reg_DO_reg[0]/P0002  & \core_eu_em_mac_em_reg_mr1swe_DO_reg[15]/P0001  ;
  assign n12028 = ~n12026 & ~n12027 ;
  assign n12029 = \core_c_dec_MFMR1_E_reg/P0001  & ~n12028 ;
  assign n12018 = ~\core_c_psq_MSTAT_reg_DO_reg[0]/P0002  & \core_eu_em_mac_em_reg_mx1rwe_DO_reg[15]/P0001  ;
  assign n12019 = \core_c_psq_MSTAT_reg_DO_reg[0]/P0002  & \core_eu_em_mac_em_reg_mx1swe_DO_reg[15]/P0001  ;
  assign n12020 = ~n12018 & ~n12019 ;
  assign n12021 = \core_c_dec_MFMX1_E_reg/P0001  & ~n12020 ;
  assign n12022 = ~\core_c_psq_MSTAT_reg_DO_reg[0]/P0002  & \core_eu_em_mac_em_reg_mr0rwe_DO_reg[15]/P0001  ;
  assign n12023 = \core_c_psq_MSTAT_reg_DO_reg[0]/P0002  & \core_eu_em_mac_em_reg_mr0swe_DO_reg[15]/P0001  ;
  assign n12024 = ~n12022 & ~n12023 ;
  assign n12025 = \core_c_dec_MFMR0_E_reg/P0001  & ~n12024 ;
  assign n12032 = ~n12021 & ~n12025 ;
  assign n12033 = ~n12029 & n12032 ;
  assign n12006 = ~\core_c_psq_MSTAT_reg_DO_reg[0]/P0002  & \core_eu_em_mac_em_reg_my0rwe_DO_reg[15]/P0001  ;
  assign n12007 = \core_c_psq_MSTAT_reg_DO_reg[0]/P0002  & \core_eu_em_mac_em_reg_my0swe_DO_reg[15]/P0001  ;
  assign n12008 = ~n12006 & ~n12007 ;
  assign n12009 = \core_c_dec_MFMY0_E_reg/P0001  & ~n12008 ;
  assign n12030 = ~n7207 & ~n12009 ;
  assign n12010 = ~\core_c_psq_MSTAT_reg_DO_reg[0]/P0002  & \core_eu_em_mac_em_reg_my1rwe_DO_reg[15]/P0001  ;
  assign n12011 = \core_c_psq_MSTAT_reg_DO_reg[0]/P0002  & \core_eu_em_mac_em_reg_my1swe_DO_reg[15]/P0001  ;
  assign n12012 = ~n12010 & ~n12011 ;
  assign n12013 = \core_c_dec_MFMY1_E_reg/P0001  & ~n12012 ;
  assign n12014 = ~\core_c_psq_MSTAT_reg_DO_reg[0]/P0002  & \core_eu_em_mac_em_reg_mx0rwe_DO_reg[15]/P0001  ;
  assign n12015 = \core_c_psq_MSTAT_reg_DO_reg[0]/P0002  & \core_eu_em_mac_em_reg_mx0swe_DO_reg[15]/P0001  ;
  assign n12016 = ~n12014 & ~n12015 ;
  assign n12017 = \core_c_dec_MFMX0_E_reg/P0001  & ~n12016 ;
  assign n12031 = ~n12013 & ~n12017 ;
  assign n12034 = n12030 & n12031 ;
  assign n12035 = n12033 & n12034 ;
  assign n12036 = n7179 & ~n12035 ;
  assign n12093 = ~n12005 & ~n12036 ;
  assign n12094 = n12092 & n12093 ;
  assign n12095 = ~n12089 & n12094 ;
  assign n12096 = ~n11964 & n12095 ;
  assign n12097 = n11770 & ~n12096 ;
  assign n12100 = \bdma_BRdataBUF_reg[15]/P0001  & n6918 ;
  assign n11963 = \idma_DTMP_H_reg[15]/P0001  & n11762 ;
  assign n12098 = \sport0_rxctl_RX_reg[15]/P0001  & n11774 ;
  assign n12099 = \sport1_rxctl_RX_reg[15]/P0001  & n11772 ;
  assign n12101 = ~n12098 & ~n12099 ;
  assign n12102 = ~n11963 & n12101 ;
  assign n12103 = ~n12100 & n12102 ;
  assign n12104 = ~n12097 & n12103 ;
  assign n12106 = ~n9430 & n11770 ;
  assign n12109 = \bdma_BRdataBUF_reg[1]/P0001  & n6918 ;
  assign n12105 = \idma_DTMP_H_reg[1]/P0001  & n11762 ;
  assign n12107 = \sport1_rxctl_RX_reg[1]/P0001  & n11772 ;
  assign n12108 = \sport0_rxctl_RX_reg[1]/P0001  & n11774 ;
  assign n12110 = ~n12107 & ~n12108 ;
  assign n12111 = ~n12105 & n12110 ;
  assign n12112 = ~n12109 & n12111 ;
  assign n12113 = ~n12106 & n12112 ;
  assign n12115 = ~n8710 & n11770 ;
  assign n12118 = \bdma_BRdataBUF_reg[2]/P0001  & n6918 ;
  assign n12114 = \idma_DTMP_H_reg[2]/P0001  & n11762 ;
  assign n12116 = \sport1_rxctl_RX_reg[2]/P0001  & n11772 ;
  assign n12117 = \sport0_rxctl_RX_reg[2]/P0001  & n11774 ;
  assign n12119 = ~n12116 & ~n12117 ;
  assign n12120 = ~n12114 & n12119 ;
  assign n12121 = ~n12118 & n12120 ;
  assign n12122 = ~n12115 & n12121 ;
  assign n12124 = ~n8108 & n11770 ;
  assign n12127 = \bdma_BRdataBUF_reg[3]/P0001  & n6918 ;
  assign n12123 = \idma_DTMP_H_reg[3]/P0001  & n11762 ;
  assign n12125 = \sport1_rxctl_RX_reg[3]/P0001  & n11772 ;
  assign n12126 = \sport0_rxctl_RX_reg[3]/P0001  & n11774 ;
  assign n12128 = ~n12125 & ~n12126 ;
  assign n12129 = ~n12123 & n12128 ;
  assign n12130 = ~n12127 & n12129 ;
  assign n12131 = ~n12124 & n12130 ;
  assign n12133 = ~n10064 & n11770 ;
  assign n12136 = \bdma_BRdataBUF_reg[4]/P0001  & n6918 ;
  assign n12132 = \idma_DTMP_H_reg[4]/P0001  & n11762 ;
  assign n12134 = \sport1_rxctl_RX_reg[4]/P0001  & n11772 ;
  assign n12135 = \sport0_rxctl_RX_reg[4]/P0001  & n11774 ;
  assign n12137 = ~n12134 & ~n12135 ;
  assign n12138 = ~n12132 & n12137 ;
  assign n12139 = ~n12136 & n12138 ;
  assign n12140 = ~n12133 & n12139 ;
  assign n12142 = ~n10906 & n11770 ;
  assign n12145 = \bdma_BRdataBUF_reg[5]/P0001  & n6918 ;
  assign n12141 = \idma_DTMP_H_reg[5]/P0001  & n11762 ;
  assign n12143 = \sport1_rxctl_RX_reg[5]/P0001  & n11772 ;
  assign n12144 = \sport0_rxctl_RX_reg[5]/P0001  & n11774 ;
  assign n12146 = ~n12143 & ~n12144 ;
  assign n12147 = ~n12141 & n12146 ;
  assign n12148 = ~n12145 & n12147 ;
  assign n12149 = ~n12142 & n12148 ;
  assign n12151 = ~n11520 & n11770 ;
  assign n12154 = \bdma_BRdataBUF_reg[6]/P0001  & n6918 ;
  assign n12150 = \idma_DTMP_H_reg[6]/P0001  & n11762 ;
  assign n12152 = \sport1_rxctl_RX_reg[6]/P0001  & n11772 ;
  assign n12153 = \sport0_rxctl_RX_reg[6]/P0001  & n11774 ;
  assign n12155 = ~n12152 & ~n12153 ;
  assign n12156 = ~n12150 & n12155 ;
  assign n12157 = ~n12154 & n12156 ;
  assign n12158 = ~n12151 & n12157 ;
  assign n12163 = ~n11260 & n11770 ;
  assign n12162 = \idma_DTMP_H_reg[7]/P0001  & n11762 ;
  assign n12159 = \bdma_BRdataBUF_reg[7]/P0001  & n6918 ;
  assign n12160 = \sport1_rxctl_RX_reg[7]/P0001  & n11772 ;
  assign n12161 = \sport0_rxctl_RX_reg[7]/P0001  & n11774 ;
  assign n12164 = ~n12160 & ~n12161 ;
  assign n12165 = ~n12159 & n12164 ;
  assign n12166 = ~n12162 & n12165 ;
  assign n12167 = ~n12163 & n12166 ;
  assign n12169 = ~n10633 & n11770 ;
  assign n12172 = \bdma_BRdataBUF_reg[8]/P0001  & n6918 ;
  assign n12168 = \idma_DTMP_H_reg[8]/P0001  & n11762 ;
  assign n12170 = \sport1_rxctl_RX_reg[8]/P0001  & n11772 ;
  assign n12171 = \sport0_rxctl_RX_reg[8]/P0001  & n11774 ;
  assign n12173 = ~n12170 & ~n12171 ;
  assign n12174 = ~n12168 & n12173 ;
  assign n12175 = ~n12172 & n12174 ;
  assign n12176 = ~n12169 & n12175 ;
  assign n12178 = ~n10284 & n11770 ;
  assign n12181 = \bdma_BRdataBUF_reg[9]/P0001  & n6918 ;
  assign n12177 = \idma_DTMP_H_reg[9]/P0001  & n11762 ;
  assign n12179 = \sport0_rxctl_RX_reg[9]/P0001  & n11774 ;
  assign n12180 = \sport1_rxctl_RX_reg[9]/P0001  & n11772 ;
  assign n12182 = ~n12179 & ~n12180 ;
  assign n12183 = ~n12177 & n12182 ;
  assign n12184 = ~n12181 & n12183 ;
  assign n12185 = ~n12178 & n12184 ;
  assign n12186 = \core_c_psq_DMOVL_reg_DO_reg[2]/NET0131  & ~n5066 ;
  assign n12187 = \bdma_BOVL_reg[6]/NET0131  & n5066 ;
  assign n12188 = ~n12186 & ~n12187 ;
  assign n12189 = ~n5895 & ~n12188 ;
  assign n12190 = \idma_DOVL_reg[6]/NET0131  & n5895 ;
  assign n12191 = ~n12189 & ~n12190 ;
  assign n12192 = \core_c_psq_DMOVL_reg_DO_reg[3]/NET0131  & ~n5066 ;
  assign n12193 = \bdma_BOVL_reg[7]/NET0131  & n5066 ;
  assign n12194 = ~n12192 & ~n12193 ;
  assign n12195 = ~n5895 & ~n12194 ;
  assign n12196 = \idma_DOVL_reg[7]/NET0131  & n5895 ;
  assign n12197 = ~n12195 & ~n12196 ;
  assign n12198 = n12191 & n12197 ;
  assign n12199 = \core_c_psq_DMOVL_reg_DO_reg[0]/NET0131  & ~n5066 ;
  assign n12200 = \bdma_BOVL_reg[4]/NET0131  & n5066 ;
  assign n12201 = ~n12199 & ~n12200 ;
  assign n12202 = ~n5895 & ~n12201 ;
  assign n12203 = \idma_DOVL_reg[4]/NET0131  & n5895 ;
  assign n12204 = ~n12202 & ~n12203 ;
  assign n12205 = n12198 & n12204 ;
  assign n12206 = \core_c_psq_DMOVL_reg_DO_reg[1]/NET0131  & ~n5066 ;
  assign n12207 = \bdma_BOVL_reg[5]/NET0131  & n5066 ;
  assign n12208 = ~n12206 & ~n12207 ;
  assign n12209 = ~n5895 & ~n12208 ;
  assign n12210 = \idma_DOVL_reg[5]/NET0131  & n5895 ;
  assign n12211 = ~n12209 & ~n12210 ;
  assign n12212 = n9513 & n12211 ;
  assign n12213 = n12205 & n12212 ;
  assign n12214 = ~n11766 & n12213 ;
  assign n12215 = n12198 & ~n12204 ;
  assign n12216 = n12212 & n12215 ;
  assign n12217 = ~n11766 & n12216 ;
  assign n12218 = n9513 & ~n12211 ;
  assign n12219 = n12205 & n12218 ;
  assign n12220 = ~n11766 & n12219 ;
  assign n12221 = n12215 & n12218 ;
  assign n12222 = ~n11766 & n12221 ;
  assign n12223 = ~n12191 & n12197 ;
  assign n12224 = n12204 & n12223 ;
  assign n12225 = n12212 & n12224 ;
  assign n12226 = ~n11766 & n12225 ;
  assign n12227 = ~n12204 & n12223 ;
  assign n12228 = n12212 & n12227 ;
  assign n12229 = ~n11766 & n12228 ;
  assign n12230 = n12218 & n12224 ;
  assign n12231 = ~n11766 & n12230 ;
  assign n12232 = n12218 & n12227 ;
  assign n12233 = ~n11766 & n12232 ;
  assign n12234 = T_ICE_RSTn_pad & T_RSTn_pad ;
  assign n12235 = \clkc_DSPoff_reg/NET0131  & n12234 ;
  assign n12236 = \clkc_SlowDn_reg/NET0131  & n12234 ;
  assign n12239 = \clkc_OSCoff_reg/NET0131  & n12234 ;
  assign n12237 = ~T_CLKI_PLL_pad & T_Sel_PLL_pad ;
  assign n12238 = ~T_CLKI_OSC_pad & ~T_Sel_PLL_pad ;
  assign n12240 = ~n12237 & ~n12238 ;
  assign n12241 = ~n12239 & n12240 ;
  assign n12242 = ~n12236 & n12241 ;
  assign n12243 = \clkc_ckSTDCLK_STDCLK_reg_Q_reg/NET0131  & n12236 ;
  assign n12244 = ~n12242 & ~n12243 ;
  assign n12245 = ~n12235 & n12244 ;
  assign n12246 = \core_dag_ilm1reg_DMA_pi_DO_reg[0]/NET0131  & n5602 ;
  assign n12247 = \emc_ECS_reg[3]/NET0131  & n5592 ;
  assign n12248 = \emc_ECMcs_reg/NET0131  & n12247 ;
  assign n12249 = \sice_idr1_reg_DO_reg[4]/P0001  & n12248 ;
  assign n12250 = \emc_ECMcs_reg/NET0131  & ~n12247 ;
  assign n12251 = \emc_ECMA_reg[0]/P0001  & n12250 ;
  assign n12254 = ~n12249 & ~n12251 ;
  assign n12255 = ~n12246 & n12254 ;
  assign n12252 = \core_dag_ilm2reg_PMA_pi_DO_reg[0]/NET0131  & ~n5608 ;
  assign n12253 = \core_c_dec_IRE_reg[4]/NET0131  & n5610 ;
  assign n12256 = ~n12252 & ~n12253 ;
  assign n12257 = n12255 & n12256 ;
  assign n12258 = ~\bdma_BM_cyc_reg/P0001  & ~n12257 ;
  assign n12259 = \bdma_BEAD_reg[0]/NET0131  & \bdma_BM_cyc_reg/P0001  ;
  assign n12260 = ~n12258 & ~n12259 ;
  assign n12261 = \bdma_BEAD_reg[10]/NET0131  & \bdma_BM_cyc_reg/P0001  ;
  assign n12262 = \core_dag_ilm1reg_DMA_pi_DO_reg[10]/NET0131  & n5602 ;
  assign n12264 = \emc_ECMA_reg[10]/P0001  & \emc_ECMcs_reg/NET0131  ;
  assign n12266 = ~n12262 & ~n12264 ;
  assign n12263 = \core_dag_ilm2reg_PMA_pi_DO_reg[10]/NET0131  & ~n5608 ;
  assign n12265 = \core_c_dec_IRE_reg[14]/NET0131  & n5610 ;
  assign n12267 = ~n12263 & ~n12265 ;
  assign n12268 = n12266 & n12267 ;
  assign n12269 = ~\bdma_BM_cyc_reg/P0001  & ~n12268 ;
  assign n12270 = ~n12261 & ~n12269 ;
  assign n12271 = \bdma_BEAD_reg[12]/NET0131  & \bdma_BM_cyc_reg/P0001  ;
  assign n12273 = ~\core_c_psq_PMOVL_regl_DO_reg[3]/NET0131  & ~n5673 ;
  assign n12274 = \core_c_psq_PMOVL_regl_DO_reg[1]/NET0131  & \core_c_psq_PMOVL_regl_DO_reg[2]/NET0131  ;
  assign n12275 = n5642 & ~n12274 ;
  assign n12276 = n12273 & n12275 ;
  assign n12278 = ~\core_c_psq_PMOVL_regl_DO_reg[0]/NET0131  & n12276 ;
  assign n12277 = ~\emc_ECMA_reg[12]/P0001  & ~n12276 ;
  assign n12279 = ~PM_bdry_sel_pad & ~n12277 ;
  assign n12280 = ~n12278 & n12279 ;
  assign n12284 = ~\core_c_psq_PMOVL_regl_DO_reg[3]/NET0131  & n5643 ;
  assign n12281 = ~\core_c_psq_PMOVL_regl_DO_reg[0]/NET0131  & n5673 ;
  assign n12282 = ~\core_c_psq_PMOVL_regl_DO_reg[1]/NET0131  & ~\core_c_psq_PMOVL_regl_DO_reg[2]/NET0131  ;
  assign n12283 = ~\emc_ECMA_reg[12]/P0001  & n12282 ;
  assign n12285 = n12281 & ~n12283 ;
  assign n12286 = n12284 & n12285 ;
  assign n12287 = ~n12280 & ~n12286 ;
  assign n12288 = \emc_ECMcs_reg/NET0131  & ~n12287 ;
  assign n12272 = \core_dag_ilm1reg_DMA_pi_DO_reg[12]/NET0131  & n5602 ;
  assign n12289 = ~PM_bdry_sel_pad & ~\core_c_psq_PMOVL_regh_DO_reg[0]/NET0131  ;
  assign n12290 = PM_bdry_sel_pad & ~\core_dag_ilm2reg_PMA_pi_DO_reg[12]/NET0131  ;
  assign n12291 = ~n12289 & ~n12290 ;
  assign n12292 = ~n5608 & n12291 ;
  assign n12293 = ~n12272 & ~n12292 ;
  assign n12294 = ~n12288 & n12293 ;
  assign n12295 = ~\bdma_BM_cyc_reg/P0001  & ~n12294 ;
  assign n12296 = ~n12271 & ~n12295 ;
  assign n12298 = \core_c_psq_PMOVL_regl_DO_reg[0]/NET0131  & n5673 ;
  assign n12299 = ~\core_c_psq_PMOVL_regl_DO_reg[1]/NET0131  & n12298 ;
  assign n12300 = \core_c_psq_PMOVL_regl_DO_reg[1]/NET0131  & n12281 ;
  assign n12301 = ~n12299 & ~n12300 ;
  assign n12302 = n12284 & ~n12301 ;
  assign n12303 = ~PM_bdry_sel_pad & n12273 ;
  assign n12304 = ~\core_c_psq_PMOVL_regl_DO_reg[1]/NET0131  & n5642 ;
  assign n12305 = n12303 & n12304 ;
  assign n12306 = ~n12302 & ~n12305 ;
  assign n12307 = \emc_ECMcs_reg/NET0131  & ~n12306 ;
  assign n12297 = \core_c_psq_DMOVL_reg_DO_reg[0]/NET0131  & n5602 ;
  assign n12308 = ~PM_bdry_sel_pad & ~\core_c_psq_PMOVL_regh_DO_reg[1]/NET0131  ;
  assign n12309 = PM_bdry_sel_pad & ~\core_c_psq_PMOVL_regh_DO_reg[0]/NET0131  ;
  assign n12310 = ~n12308 & ~n12309 ;
  assign n12311 = ~n5608 & n12310 ;
  assign n12312 = ~n12297 & ~n12311 ;
  assign n12313 = ~n12307 & n12312 ;
  assign n12314 = ~\bdma_BM_cyc_reg/P0001  & ~n12313 ;
  assign n12315 = \bdma_BEAD_reg[13]/NET0131  & \bdma_BM_cyc_reg/P0001  ;
  assign n12316 = ~n12314 & ~n12315 ;
  assign n12318 = ~n12281 & ~n12299 ;
  assign n12319 = \core_c_psq_PMOVL_regl_DO_reg[2]/NET0131  & ~n12318 ;
  assign n12320 = \core_c_psq_PMOVL_regl_DO_reg[1]/NET0131  & ~\core_c_psq_PMOVL_regl_DO_reg[2]/NET0131  ;
  assign n12321 = n12298 & n12320 ;
  assign n12322 = ~n12319 & ~n12321 ;
  assign n12323 = n12284 & ~n12322 ;
  assign n12324 = n12275 & ~n12282 ;
  assign n12325 = n12303 & n12324 ;
  assign n12326 = ~n12323 & ~n12325 ;
  assign n12327 = \emc_ECMcs_reg/NET0131  & ~n12326 ;
  assign n12317 = \core_c_psq_DMOVL_reg_DO_reg[1]/NET0131  & n5602 ;
  assign n12328 = ~PM_bdry_sel_pad & ~\core_c_psq_PMOVL_regh_DO_reg[2]/NET0131  ;
  assign n12329 = PM_bdry_sel_pad & ~\core_c_psq_PMOVL_regh_DO_reg[1]/NET0131  ;
  assign n12330 = ~n12328 & ~n12329 ;
  assign n12331 = ~n5608 & n12330 ;
  assign n12332 = ~n12317 & ~n12331 ;
  assign n12333 = ~n12327 & n12332 ;
  assign n12334 = ~\bdma_BM_cyc_reg/P0001  & ~n12333 ;
  assign n12335 = \bdma_BCTL_reg[8]/NET0131  & \bdma_BM_cyc_reg/P0001  ;
  assign n12336 = ~n12334 & ~n12335 ;
  assign n12337 = \core_dag_ilm1reg_DMA_pi_DO_reg[1]/NET0131  & n5602 ;
  assign n12338 = \sice_idr1_reg_DO_reg[5]/P0001  & n12248 ;
  assign n12339 = \emc_ECMA_reg[1]/P0001  & n12250 ;
  assign n12342 = ~n12338 & ~n12339 ;
  assign n12343 = ~n12337 & n12342 ;
  assign n12340 = \core_dag_ilm2reg_PMA_pi_DO_reg[1]/NET0131  & ~n5608 ;
  assign n12341 = \core_c_dec_IRE_reg[5]/NET0131  & n5610 ;
  assign n12344 = ~n12340 & ~n12341 ;
  assign n12345 = n12343 & n12344 ;
  assign n12346 = ~\bdma_BM_cyc_reg/P0001  & ~n12345 ;
  assign n12347 = \bdma_BEAD_reg[1]/NET0131  & \bdma_BM_cyc_reg/P0001  ;
  assign n12348 = ~n12346 & ~n12347 ;
  assign n12349 = \core_dag_ilm1reg_DMA_pi_DO_reg[2]/NET0131  & n5602 ;
  assign n12350 = \sice_idr1_reg_DO_reg[6]/P0001  & n12248 ;
  assign n12351 = \emc_ECMA_reg[2]/P0001  & n12250 ;
  assign n12354 = ~n12350 & ~n12351 ;
  assign n12355 = ~n12349 & n12354 ;
  assign n12352 = \core_dag_ilm2reg_PMA_pi_DO_reg[2]/NET0131  & ~n5608 ;
  assign n12353 = \core_c_dec_IRE_reg[6]/NET0131  & n5610 ;
  assign n12356 = ~n12352 & ~n12353 ;
  assign n12357 = n12355 & n12356 ;
  assign n12358 = ~\bdma_BM_cyc_reg/P0001  & ~n12357 ;
  assign n12359 = \bdma_BEAD_reg[2]/NET0131  & \bdma_BM_cyc_reg/P0001  ;
  assign n12360 = ~n12358 & ~n12359 ;
  assign n12361 = \core_dag_ilm1reg_DMA_pi_DO_reg[3]/NET0131  & n5602 ;
  assign n12362 = \sice_idr1_reg_DO_reg[7]/P0001  & n12248 ;
  assign n12363 = \emc_ECMA_reg[3]/P0001  & n12250 ;
  assign n12366 = ~n12362 & ~n12363 ;
  assign n12367 = ~n12361 & n12366 ;
  assign n12364 = \core_dag_ilm2reg_PMA_pi_DO_reg[3]/NET0131  & ~n5608 ;
  assign n12365 = \core_c_dec_IRE_reg[7]/NET0131  & n5610 ;
  assign n12368 = ~n12364 & ~n12365 ;
  assign n12369 = n12367 & n12368 ;
  assign n12370 = ~\bdma_BM_cyc_reg/P0001  & ~n12369 ;
  assign n12371 = \bdma_BEAD_reg[3]/NET0131  & \bdma_BM_cyc_reg/P0001  ;
  assign n12372 = ~n12370 & ~n12371 ;
  assign n12373 = \core_dag_ilm1reg_DMA_pi_DO_reg[4]/NET0131  & n5602 ;
  assign n12374 = \sice_idr1_reg_DO_reg[8]/P0001  & n12248 ;
  assign n12375 = \emc_ECMA_reg[4]/P0001  & n12250 ;
  assign n12378 = ~n12374 & ~n12375 ;
  assign n12379 = ~n12373 & n12378 ;
  assign n12376 = \core_dag_ilm2reg_PMA_pi_DO_reg[4]/NET0131  & ~n5608 ;
  assign n12377 = \core_c_dec_IRE_reg[8]/NET0131  & n5610 ;
  assign n12380 = ~n12376 & ~n12377 ;
  assign n12381 = n12379 & n12380 ;
  assign n12382 = ~\bdma_BM_cyc_reg/P0001  & ~n12381 ;
  assign n12383 = \bdma_BEAD_reg[4]/NET0131  & \bdma_BM_cyc_reg/P0001  ;
  assign n12384 = ~n12382 & ~n12383 ;
  assign n12385 = \core_dag_ilm1reg_DMA_pi_DO_reg[5]/NET0131  & n5602 ;
  assign n12386 = \sice_idr1_reg_DO_reg[9]/P0001  & n12248 ;
  assign n12387 = \emc_ECMA_reg[5]/P0001  & n12250 ;
  assign n12390 = ~n12386 & ~n12387 ;
  assign n12391 = ~n12385 & n12390 ;
  assign n12388 = \core_dag_ilm2reg_PMA_pi_DO_reg[5]/NET0131  & ~n5608 ;
  assign n12389 = \core_c_dec_IRE_reg[9]/NET0131  & n5610 ;
  assign n12392 = ~n12388 & ~n12389 ;
  assign n12393 = n12391 & n12392 ;
  assign n12394 = ~\bdma_BM_cyc_reg/P0001  & ~n12393 ;
  assign n12395 = \bdma_BEAD_reg[5]/NET0131  & \bdma_BM_cyc_reg/P0001  ;
  assign n12396 = ~n12394 & ~n12395 ;
  assign n12397 = \core_dag_ilm1reg_DMA_pi_DO_reg[6]/NET0131  & n5602 ;
  assign n12398 = \sice_idr1_reg_DO_reg[10]/P0001  & n12248 ;
  assign n12399 = \emc_ECMA_reg[6]/P0001  & n12250 ;
  assign n12402 = ~n12398 & ~n12399 ;
  assign n12403 = ~n12397 & n12402 ;
  assign n12400 = \core_dag_ilm2reg_PMA_pi_DO_reg[6]/NET0131  & ~n5608 ;
  assign n12401 = \core_c_dec_IRE_reg[10]/NET0131  & n5610 ;
  assign n12404 = ~n12400 & ~n12401 ;
  assign n12405 = n12403 & n12404 ;
  assign n12406 = ~\bdma_BM_cyc_reg/P0001  & ~n12405 ;
  assign n12407 = \bdma_BEAD_reg[6]/NET0131  & \bdma_BM_cyc_reg/P0001  ;
  assign n12408 = ~n12406 & ~n12407 ;
  assign n12409 = \core_dag_ilm1reg_DMA_pi_DO_reg[7]/NET0131  & n5602 ;
  assign n12410 = \sice_idr1_reg_DO_reg[11]/P0001  & n12248 ;
  assign n12411 = \emc_ECMA_reg[7]/P0001  & n12250 ;
  assign n12414 = ~n12410 & ~n12411 ;
  assign n12415 = ~n12409 & n12414 ;
  assign n12412 = \core_dag_ilm2reg_PMA_pi_DO_reg[7]/NET0131  & ~n5608 ;
  assign n12413 = \core_c_dec_IRE_reg[11]/NET0131  & n5610 ;
  assign n12416 = ~n12412 & ~n12413 ;
  assign n12417 = n12415 & n12416 ;
  assign n12418 = ~\bdma_BM_cyc_reg/P0001  & ~n12417 ;
  assign n12419 = \bdma_BEAD_reg[7]/NET0131  & \bdma_BM_cyc_reg/P0001  ;
  assign n12420 = ~n12418 & ~n12419 ;
  assign n12421 = \bdma_BEAD_reg[8]/NET0131  & \bdma_BM_cyc_reg/P0001  ;
  assign n12422 = \core_dag_ilm1reg_DMA_pi_DO_reg[8]/NET0131  & n5602 ;
  assign n12424 = \emc_ECMA_reg[8]/P0001  & \emc_ECMcs_reg/NET0131  ;
  assign n12426 = ~n12422 & ~n12424 ;
  assign n12423 = \core_dag_ilm2reg_PMA_pi_DO_reg[8]/NET0131  & ~n5608 ;
  assign n12425 = \core_c_dec_IRE_reg[12]/NET0131  & n5610 ;
  assign n12427 = ~n12423 & ~n12425 ;
  assign n12428 = n12426 & n12427 ;
  assign n12429 = ~\bdma_BM_cyc_reg/P0001  & ~n12428 ;
  assign n12430 = ~n12421 & ~n12429 ;
  assign n12431 = \bdma_BEAD_reg[9]/NET0131  & \bdma_BM_cyc_reg/P0001  ;
  assign n12432 = \core_dag_ilm1reg_DMA_pi_DO_reg[9]/NET0131  & n5602 ;
  assign n12434 = \emc_ECMA_reg[9]/P0001  & \emc_ECMcs_reg/NET0131  ;
  assign n12436 = ~n12432 & ~n12434 ;
  assign n12433 = \core_dag_ilm2reg_PMA_pi_DO_reg[9]/NET0131  & ~n5608 ;
  assign n12435 = \core_c_dec_IRE_reg[13]/NET0131  & n5610 ;
  assign n12437 = ~n12433 & ~n12435 ;
  assign n12438 = n12436 & n12437 ;
  assign n12439 = ~\bdma_BM_cyc_reg/P0001  & ~n12438 ;
  assign n12440 = ~n12431 & ~n12439 ;
  assign n12441 = ~n5602 & ~n5610 ;
  assign n12444 = ~\emc_ECS_reg[1]/NET0131  & n5523 ;
  assign n12442 = \core_c_dec_accCM_E_reg/NET0131  & ~\core_c_dec_rdCM_E_reg/NET0131  ;
  assign n12443 = n12247 & n12442 ;
  assign n12445 = ~\bdma_BM_cyc_reg/P0001  & ~n5519 ;
  assign n12446 = ~n12443 & n12445 ;
  assign n12447 = ~n12444 & n12446 ;
  assign n12448 = n5608 & n12447 ;
  assign n12449 = n12441 & n12448 ;
  assign n12450 = ~\core_c_psq_MGNT_reg/NET0131  & ~n12449 ;
  assign n12451 = ~\core_c_psq_MGNT_reg/NET0131  & \emc_ED_oei_reg/P0001  ;
  assign n12452 = \emc_selPMDi_reg/P0001  & ~n5608 ;
  assign n12453 = \emc_selDMDi_reg/P0001  & ~n12441 ;
  assign n12456 = ~n12452 & n12453 ;
  assign n12457 = n7607 & n12456 ;
  assign n12454 = ~n12452 & ~n12453 ;
  assign n12455 = \sice_idr0_reg_DO_reg[0]/P0001  & n12454 ;
  assign n12470 = \core_c_dec_pMFMAC_Ei_reg/NET0131  & ~n6988 ;
  assign n12471 = ~n7480 & n12470 ;
  assign n12466 = \core_c_dec_pMFSHT_Ei_reg/NET0131  & ~n6988 ;
  assign n12467 = ~n7386 & n12466 ;
  assign n12468 = \core_c_dec_pMFALU_Ei_reg/NET0131  & ~n6988 ;
  assign n12469 = ~n7437 & n12468 ;
  assign n12472 = ~n12467 & ~n12469 ;
  assign n12473 = ~n12471 & n12472 ;
  assign n12474 = ~\emc_PMDoe_reg/NET0131  & ~n12473 ;
  assign n12458 = \emc_PMDoe_reg/NET0131  & \emc_PMDreg_reg[0]/P0001  ;
  assign n12459 = ~\memc_PMo_oe2_reg/P0001  & ~\memc_PMo_oe3_reg/P0001  ;
  assign n12460 = ~\memc_PMo_oe4_reg/P0001  & ~\memc_PMo_oe5_reg/P0001  ;
  assign n12461 = ~\memc_PMo_oe6_reg/P0001  & n12460 ;
  assign n12462 = ~\memc_PMo_oe7_reg/P0001  & n12461 ;
  assign n12463 = ~\memc_PMo_oe0_reg/P0001  & ~\memc_PMo_oe1_reg/P0001  ;
  assign n12464 = n12462 & n12463 ;
  assign n12465 = n12459 & n12464 ;
  assign n12475 = ~n12458 & n12465 ;
  assign n12476 = ~n12474 & n12475 ;
  assign n12477 = \memc_PMo_oe2_reg/P0001  & ~\memc_PMo_oe3_reg/P0001  ;
  assign n12478 = n12464 & n12477 ;
  assign n12480 = n12459 & n12463 ;
  assign n12481 = ~\memc_PMo_oe7_reg/P0001  & n12480 ;
  assign n12482 = \memc_PMo_oe6_reg/P0001  & n12460 ;
  assign n12483 = n12481 & n12482 ;
  assign n12484 = \memc_PMo_oe7_reg/P0001  & n12461 ;
  assign n12485 = n12480 & n12484 ;
  assign n12496 = ~n12483 & ~n12485 ;
  assign n12497 = ~n12478 & n12496 ;
  assign n12486 = ~\memc_PMo_oe6_reg/P0001  & n12481 ;
  assign n12487 = \memc_PMo_oe4_reg/P0001  & ~\memc_PMo_oe5_reg/P0001  ;
  assign n12488 = n12486 & n12487 ;
  assign n12489 = n12459 & n12462 ;
  assign n12490 = ~\memc_PMo_oe0_reg/P0001  & \memc_PMo_oe1_reg/P0001  ;
  assign n12491 = n12489 & n12490 ;
  assign n12498 = ~n12488 & ~n12491 ;
  assign n12492 = ~\memc_PMo_oe2_reg/P0001  & \memc_PMo_oe3_reg/P0001  ;
  assign n12493 = n12464 & n12492 ;
  assign n12494 = ~\memc_PMo_oe4_reg/P0001  & \memc_PMo_oe5_reg/P0001  ;
  assign n12495 = n12486 & n12494 ;
  assign n12499 = ~n12493 & ~n12495 ;
  assign n12500 = n12498 & n12499 ;
  assign n12501 = n12497 & n12500 ;
  assign n12502 = \memc_PMo_oe0_reg/P0001  & ~\memc_PMo_oe1_reg/P0001  ;
  assign n12503 = n12489 & n12502 ;
  assign n12504 = ~n12501 & ~n12503 ;
  assign n12505 = \PM_rd0[0]_pad  & ~n12504 ;
  assign n12511 = \PM_rd5[0]_pad  & n12495 ;
  assign n12509 = \PM_rd3[0]_pad  & n12493 ;
  assign n12510 = \PM_rd1[0]_pad  & n12491 ;
  assign n12515 = ~n12509 & ~n12510 ;
  assign n12516 = ~n12511 & n12515 ;
  assign n12508 = \PM_rd7[0]_pad  & n12485 ;
  assign n12507 = \PM_rd6[0]_pad  & n12483 ;
  assign n12512 = ~n12465 & ~n12507 ;
  assign n12513 = ~n12508 & n12512 ;
  assign n12479 = \PM_rd2[0]_pad  & n12478 ;
  assign n12506 = \PM_rd4[0]_pad  & n12488 ;
  assign n12514 = ~n12479 & ~n12506 ;
  assign n12517 = n12513 & n12514 ;
  assign n12518 = n12516 & n12517 ;
  assign n12519 = ~n12505 & n12518 ;
  assign n12520 = ~n12476 & ~n12519 ;
  assign n12521 = n12452 & n12520 ;
  assign n12522 = ~n12455 & ~n12521 ;
  assign n12523 = ~n12457 & n12522 ;
  assign n12524 = n12451 & ~n12523 ;
  assign n12525 = \bdma_BCTL_reg[2]/NET0131  & \bdma_BM_cyc_reg/P0001  ;
  assign n12526 = \bdma_BWdataBUF_reg[0]/P0001  & n12525 ;
  assign n12527 = ~n12524 & ~n12526 ;
  assign n12528 = \bdma_BCTL_reg[11]/NET0131  & \bdma_BM_cyc_reg/P0001  ;
  assign n12530 = n7859 & n12456 ;
  assign n12529 = \sice_idr0_reg_DO_reg[10]/P0001  & n12454 ;
  assign n12534 = ~n7789 & n12468 ;
  assign n12532 = ~n7764 & n12470 ;
  assign n12533 = ~n7813 & n12466 ;
  assign n12535 = ~n12532 & ~n12533 ;
  assign n12536 = ~n12534 & n12535 ;
  assign n12537 = ~\emc_PMDoe_reg/NET0131  & ~n12536 ;
  assign n12531 = \emc_PMDoe_reg/NET0131  & \emc_PMDreg_reg[10]/P0001  ;
  assign n12538 = n12465 & ~n12531 ;
  assign n12539 = ~n12537 & n12538 ;
  assign n12541 = \PM_rd0[10]_pad  & ~n12504 ;
  assign n12547 = \PM_rd5[10]_pad  & n12495 ;
  assign n12545 = \PM_rd3[10]_pad  & n12493 ;
  assign n12546 = \PM_rd1[10]_pad  & n12491 ;
  assign n12551 = ~n12545 & ~n12546 ;
  assign n12552 = ~n12547 & n12551 ;
  assign n12544 = \PM_rd7[10]_pad  & n12485 ;
  assign n12543 = \PM_rd6[10]_pad  & n12483 ;
  assign n12548 = ~n12465 & ~n12543 ;
  assign n12549 = ~n12544 & n12548 ;
  assign n12540 = \PM_rd2[10]_pad  & n12478 ;
  assign n12542 = \PM_rd4[10]_pad  & n12488 ;
  assign n12550 = ~n12540 & ~n12542 ;
  assign n12553 = n12549 & n12550 ;
  assign n12554 = n12552 & n12553 ;
  assign n12555 = ~n12541 & n12554 ;
  assign n12556 = ~n12539 & ~n12555 ;
  assign n12557 = n12452 & n12556 ;
  assign n12558 = ~n12529 & ~n12557 ;
  assign n12559 = ~n12530 & n12558 ;
  assign n12560 = n12451 & ~n12559 ;
  assign n12561 = ~n12528 & ~n12560 ;
  assign n12562 = \bdma_BCTL_reg[12]/NET0131  & \bdma_BM_cyc_reg/P0001  ;
  assign n12564 = n8460 & n12456 ;
  assign n12563 = \sice_idr0_reg_DO_reg[11]/P0001  & n12454 ;
  assign n12568 = ~n8390 & n12468 ;
  assign n12566 = ~n8365 & n12470 ;
  assign n12567 = ~n8414 & n12466 ;
  assign n12569 = ~n12566 & ~n12567 ;
  assign n12570 = ~n12568 & n12569 ;
  assign n12571 = ~\emc_PMDoe_reg/NET0131  & ~n12570 ;
  assign n12565 = \emc_PMDoe_reg/NET0131  & \emc_PMDreg_reg[11]/P0001  ;
  assign n12572 = n12465 & ~n12565 ;
  assign n12573 = ~n12571 & n12572 ;
  assign n12575 = \PM_rd0[11]_pad  & ~n12504 ;
  assign n12581 = \PM_rd5[11]_pad  & n12495 ;
  assign n12579 = \PM_rd3[11]_pad  & n12493 ;
  assign n12580 = \PM_rd1[11]_pad  & n12491 ;
  assign n12585 = ~n12579 & ~n12580 ;
  assign n12586 = ~n12581 & n12585 ;
  assign n12578 = \PM_rd7[11]_pad  & n12485 ;
  assign n12577 = \PM_rd6[11]_pad  & n12483 ;
  assign n12582 = ~n12465 & ~n12577 ;
  assign n12583 = ~n12578 & n12582 ;
  assign n12574 = \PM_rd2[11]_pad  & n12478 ;
  assign n12576 = \PM_rd4[11]_pad  & n12488 ;
  assign n12584 = ~n12574 & ~n12576 ;
  assign n12587 = n12583 & n12584 ;
  assign n12588 = n12586 & n12587 ;
  assign n12589 = ~n12575 & n12588 ;
  assign n12590 = ~n12573 & ~n12589 ;
  assign n12591 = n12452 & n12590 ;
  assign n12592 = ~n12563 & ~n12591 ;
  assign n12593 = ~n12564 & n12592 ;
  assign n12594 = n12451 & ~n12593 ;
  assign n12595 = ~n12562 & ~n12594 ;
  assign n12596 = \bdma_BCTL_reg[13]/NET0131  & \bdma_BM_cyc_reg/P0001  ;
  assign n12598 = n9178 & n12456 ;
  assign n12597 = \sice_idr1_reg_DO_reg[0]/P0001  & n12454 ;
  assign n12602 = ~n9108 & n12468 ;
  assign n12600 = ~n9083 & n12470 ;
  assign n12601 = ~n9132 & n12466 ;
  assign n12603 = ~n12600 & ~n12601 ;
  assign n12604 = ~n12602 & n12603 ;
  assign n12605 = ~\emc_PMDoe_reg/NET0131  & ~n12604 ;
  assign n12599 = \emc_PMDoe_reg/NET0131  & \emc_PMDreg_reg[12]/P0001  ;
  assign n12606 = n12465 & ~n12599 ;
  assign n12607 = ~n12605 & n12606 ;
  assign n12609 = \PM_rd0[12]_pad  & ~n12504 ;
  assign n12615 = \PM_rd5[12]_pad  & n12495 ;
  assign n12613 = \PM_rd3[12]_pad  & n12493 ;
  assign n12614 = \PM_rd1[12]_pad  & n12491 ;
  assign n12619 = ~n12613 & ~n12614 ;
  assign n12620 = ~n12615 & n12619 ;
  assign n12612 = \PM_rd7[12]_pad  & n12485 ;
  assign n12611 = \PM_rd6[12]_pad  & n12483 ;
  assign n12616 = ~n12465 & ~n12611 ;
  assign n12617 = ~n12612 & n12616 ;
  assign n12608 = \PM_rd2[12]_pad  & n12478 ;
  assign n12610 = \PM_rd4[12]_pad  & n12488 ;
  assign n12618 = ~n12608 & ~n12610 ;
  assign n12621 = n12617 & n12618 ;
  assign n12622 = n12620 & n12621 ;
  assign n12623 = ~n12609 & n12622 ;
  assign n12624 = ~n12607 & ~n12623 ;
  assign n12625 = n12452 & n12624 ;
  assign n12626 = ~n12597 & ~n12625 ;
  assign n12627 = ~n12598 & n12626 ;
  assign n12628 = n12451 & ~n12627 ;
  assign n12629 = ~n12596 & ~n12628 ;
  assign n12630 = \bdma_BCTL_reg[14]/NET0131  & \bdma_BM_cyc_reg/P0001  ;
  assign n12632 = n7340 & n12456 ;
  assign n12631 = \sice_idr1_reg_DO_reg[1]/P0001  & n12454 ;
  assign n12636 = ~n7117 & n12468 ;
  assign n12634 = ~n7213 & n12470 ;
  assign n12635 = ~n7177 & n12466 ;
  assign n12637 = ~n12634 & ~n12635 ;
  assign n12638 = ~n12636 & n12637 ;
  assign n12639 = ~\emc_PMDoe_reg/NET0131  & ~n12638 ;
  assign n12633 = \emc_PMDoe_reg/NET0131  & \emc_PMDreg_reg[13]/P0001  ;
  assign n12640 = n12465 & ~n12633 ;
  assign n12641 = ~n12639 & n12640 ;
  assign n12643 = \PM_rd0[13]_pad  & ~n12504 ;
  assign n12649 = \PM_rd5[13]_pad  & n12495 ;
  assign n12647 = \PM_rd3[13]_pad  & n12493 ;
  assign n12648 = \PM_rd1[13]_pad  & n12491 ;
  assign n12653 = ~n12647 & ~n12648 ;
  assign n12654 = ~n12649 & n12653 ;
  assign n12646 = \PM_rd7[13]_pad  & n12485 ;
  assign n12645 = \PM_rd6[13]_pad  & n12483 ;
  assign n12650 = ~n12465 & ~n12645 ;
  assign n12651 = ~n12646 & n12650 ;
  assign n12642 = \PM_rd2[13]_pad  & n12478 ;
  assign n12644 = \PM_rd4[13]_pad  & n12488 ;
  assign n12652 = ~n12642 & ~n12644 ;
  assign n12655 = n12651 & n12652 ;
  assign n12656 = n12654 & n12655 ;
  assign n12657 = ~n12643 & n12656 ;
  assign n12658 = ~n12641 & ~n12657 ;
  assign n12659 = n12452 & n12658 ;
  assign n12660 = ~n12631 & ~n12659 ;
  assign n12661 = ~n12632 & n12660 ;
  assign n12662 = n12451 & ~n12661 ;
  assign n12663 = ~n12630 & ~n12662 ;
  assign n12664 = \bdma_BCTL_reg[15]/NET0131  & \bdma_BM_cyc_reg/P0001  ;
  assign n12672 = \DM_rd0[14]_pad  & ~n7053 ;
  assign n12666 = \DM_rdm[14]_pad  & n7016 ;
  assign n12677 = ~n7057 & ~n12666 ;
  assign n12669 = \DM_rd6[14]_pad  & n7031 ;
  assign n12670 = \DM_rd7[14]_pad  & n7034 ;
  assign n12678 = ~n12669 & ~n12670 ;
  assign n12679 = n12677 & n12678 ;
  assign n12673 = \DM_rd5[14]_pad  & n7043 ;
  assign n12668 = \DM_rd4[14]_pad  & n7028 ;
  assign n12674 = \DM_rd2[14]_pad  & n7041 ;
  assign n12667 = \DM_rd1[14]_pad  & n7022 ;
  assign n12671 = \DM_rd3[14]_pad  & n7038 ;
  assign n12675 = ~n12667 & ~n12671 ;
  assign n12676 = ~n12674 & n12675 ;
  assign n12680 = ~n12668 & n12676 ;
  assign n12681 = ~n12673 & n12680 ;
  assign n12682 = n12679 & n12681 ;
  assign n12683 = ~n12672 & n12682 ;
  assign n12684 = ~\emc_DMDoe_reg/NET0131  & ~n11954 ;
  assign n12685 = \emc_DMDoe_reg/NET0131  & \emc_DMDreg_reg[14]/P0001  ;
  assign n12686 = n7057 & ~n12685 ;
  assign n12687 = ~n12684 & n12686 ;
  assign n12688 = ~n12683 & ~n12687 ;
  assign n12689 = n12456 & n12688 ;
  assign n12665 = \sice_idr1_reg_DO_reg[2]/P0001  & n12454 ;
  assign n12693 = ~n11889 & n12470 ;
  assign n12691 = ~n11842 & n12468 ;
  assign n12692 = ~n11858 & n12466 ;
  assign n12694 = ~n12691 & ~n12692 ;
  assign n12695 = ~n12693 & n12694 ;
  assign n12696 = ~\emc_PMDoe_reg/NET0131  & ~n12695 ;
  assign n12690 = \emc_PMDoe_reg/NET0131  & \emc_PMDreg_reg[14]/P0001  ;
  assign n12697 = n12465 & ~n12690 ;
  assign n12698 = ~n12696 & n12697 ;
  assign n12700 = \PM_rd0[14]_pad  & ~n12504 ;
  assign n12706 = \PM_rd5[14]_pad  & n12495 ;
  assign n12704 = \PM_rd3[14]_pad  & n12493 ;
  assign n12705 = \PM_rd1[14]_pad  & n12491 ;
  assign n12710 = ~n12704 & ~n12705 ;
  assign n12711 = ~n12706 & n12710 ;
  assign n12703 = \PM_rd7[14]_pad  & n12485 ;
  assign n12702 = \PM_rd6[14]_pad  & n12483 ;
  assign n12707 = ~n12465 & ~n12702 ;
  assign n12708 = ~n12703 & n12707 ;
  assign n12699 = \PM_rd2[14]_pad  & n12478 ;
  assign n12701 = \PM_rd4[14]_pad  & n12488 ;
  assign n12709 = ~n12699 & ~n12701 ;
  assign n12712 = n12708 & n12709 ;
  assign n12713 = n12711 & n12712 ;
  assign n12714 = ~n12700 & n12713 ;
  assign n12715 = ~n12698 & ~n12714 ;
  assign n12716 = n12452 & n12715 ;
  assign n12717 = ~n12665 & ~n12716 ;
  assign n12718 = ~n12689 & n12717 ;
  assign n12719 = n12451 & ~n12718 ;
  assign n12720 = ~n12664 & ~n12719 ;
  assign n12745 = \sice_idr1_reg_DO_reg[3]/P0001  & n12454 ;
  assign n12727 = \DM_rd0[15]_pad  & ~n7053 ;
  assign n12721 = \DM_rdm[15]_pad  & n7016 ;
  assign n12732 = ~n7057 & ~n12721 ;
  assign n12724 = \DM_rd6[15]_pad  & n7031 ;
  assign n12725 = \DM_rd7[15]_pad  & n7034 ;
  assign n12733 = ~n12724 & ~n12725 ;
  assign n12734 = n12732 & n12733 ;
  assign n12728 = \DM_rd5[15]_pad  & n7043 ;
  assign n12723 = \DM_rd4[15]_pad  & n7028 ;
  assign n12729 = \DM_rd2[15]_pad  & n7041 ;
  assign n12722 = \DM_rd1[15]_pad  & n7022 ;
  assign n12726 = \DM_rd3[15]_pad  & n7038 ;
  assign n12730 = ~n12722 & ~n12726 ;
  assign n12731 = ~n12729 & n12730 ;
  assign n12735 = ~n12723 & n12731 ;
  assign n12736 = ~n12728 & n12735 ;
  assign n12737 = n12734 & n12736 ;
  assign n12738 = ~n12727 & n12737 ;
  assign n12739 = ~\emc_DMDoe_reg/NET0131  & ~n12096 ;
  assign n12740 = \emc_DMDoe_reg/NET0131  & \emc_DMDreg_reg[15]/P0001  ;
  assign n12741 = n7057 & ~n12740 ;
  assign n12742 = ~n12739 & n12741 ;
  assign n12743 = ~n12738 & ~n12742 ;
  assign n12744 = n12456 & n12743 ;
  assign n12749 = ~n12035 & n12470 ;
  assign n12747 = ~n11988 & n12468 ;
  assign n12748 = ~n12004 & n12466 ;
  assign n12750 = ~n12747 & ~n12748 ;
  assign n12751 = ~n12749 & n12750 ;
  assign n12752 = ~\emc_PMDoe_reg/NET0131  & ~n12751 ;
  assign n12746 = \emc_PMDoe_reg/NET0131  & \emc_PMDreg_reg[15]/P0001  ;
  assign n12753 = n12465 & ~n12746 ;
  assign n12754 = ~n12752 & n12753 ;
  assign n12756 = \PM_rd0[15]_pad  & ~n12504 ;
  assign n12762 = \PM_rd5[15]_pad  & n12495 ;
  assign n12760 = \PM_rd3[15]_pad  & n12493 ;
  assign n12761 = \PM_rd1[15]_pad  & n12491 ;
  assign n12766 = ~n12760 & ~n12761 ;
  assign n12767 = ~n12762 & n12766 ;
  assign n12759 = \PM_rd7[15]_pad  & n12485 ;
  assign n12758 = \PM_rd6[15]_pad  & n12483 ;
  assign n12763 = ~n12465 & ~n12758 ;
  assign n12764 = ~n12759 & n12763 ;
  assign n12755 = \PM_rd2[15]_pad  & n12478 ;
  assign n12757 = \PM_rd4[15]_pad  & n12488 ;
  assign n12765 = ~n12755 & ~n12757 ;
  assign n12768 = n12764 & n12765 ;
  assign n12769 = n12767 & n12768 ;
  assign n12770 = ~n12756 & n12769 ;
  assign n12771 = ~n12754 & ~n12770 ;
  assign n12772 = n12452 & n12771 ;
  assign n12773 = ~n12744 & ~n12772 ;
  assign n12774 = ~n12745 & n12773 ;
  assign n12776 = n9435 & n12456 ;
  assign n12775 = \sice_idr0_reg_DO_reg[1]/P0001  & n12454 ;
  assign n12780 = ~n9236 & n12470 ;
  assign n12778 = ~n9285 & n12466 ;
  assign n12779 = ~n9320 & n12468 ;
  assign n12781 = ~n12778 & ~n12779 ;
  assign n12782 = ~n12780 & n12781 ;
  assign n12783 = ~\emc_PMDoe_reg/NET0131  & ~n12782 ;
  assign n12777 = \emc_PMDoe_reg/NET0131  & \emc_PMDreg_reg[1]/P0001  ;
  assign n12784 = n12465 & ~n12777 ;
  assign n12785 = ~n12783 & n12784 ;
  assign n12787 = \PM_rd0[1]_pad  & ~n12504 ;
  assign n12793 = \PM_rd5[1]_pad  & n12495 ;
  assign n12791 = \PM_rd3[1]_pad  & n12493 ;
  assign n12792 = \PM_rd1[1]_pad  & n12491 ;
  assign n12797 = ~n12791 & ~n12792 ;
  assign n12798 = ~n12793 & n12797 ;
  assign n12790 = \PM_rd7[1]_pad  & n12485 ;
  assign n12789 = \PM_rd6[1]_pad  & n12483 ;
  assign n12794 = ~n12465 & ~n12789 ;
  assign n12795 = ~n12790 & n12794 ;
  assign n12786 = \PM_rd2[1]_pad  & n12478 ;
  assign n12788 = \PM_rd4[1]_pad  & n12488 ;
  assign n12796 = ~n12786 & ~n12788 ;
  assign n12799 = n12795 & n12796 ;
  assign n12800 = n12798 & n12799 ;
  assign n12801 = ~n12787 & n12800 ;
  assign n12802 = ~n12785 & ~n12801 ;
  assign n12803 = n12452 & n12802 ;
  assign n12804 = ~n12775 & ~n12803 ;
  assign n12805 = ~n12776 & n12804 ;
  assign n12806 = n12451 & ~n12805 ;
  assign n12807 = \bdma_BWdataBUF_reg[1]/P0001  & n12525 ;
  assign n12808 = ~n12806 & ~n12807 ;
  assign n12810 = n8715 & n12456 ;
  assign n12809 = \sice_idr0_reg_DO_reg[2]/P0001  & n12454 ;
  assign n12814 = ~n8506 & n12466 ;
  assign n12812 = ~n8565 & n12470 ;
  assign n12813 = ~n8600 & n12468 ;
  assign n12815 = ~n12812 & ~n12813 ;
  assign n12816 = ~n12814 & n12815 ;
  assign n12817 = ~\emc_PMDoe_reg/NET0131  & ~n12816 ;
  assign n12811 = \emc_PMDoe_reg/NET0131  & \emc_PMDreg_reg[2]/P0001  ;
  assign n12818 = n12465 & ~n12811 ;
  assign n12819 = ~n12817 & n12818 ;
  assign n12821 = \PM_rd0[2]_pad  & ~n12504 ;
  assign n12827 = \PM_rd5[2]_pad  & n12495 ;
  assign n12825 = \PM_rd3[2]_pad  & n12493 ;
  assign n12826 = \PM_rd1[2]_pad  & n12491 ;
  assign n12831 = ~n12825 & ~n12826 ;
  assign n12832 = ~n12827 & n12831 ;
  assign n12824 = \PM_rd7[2]_pad  & n12485 ;
  assign n12823 = \PM_rd6[2]_pad  & n12483 ;
  assign n12828 = ~n12465 & ~n12823 ;
  assign n12829 = ~n12824 & n12828 ;
  assign n12820 = \PM_rd2[2]_pad  & n12478 ;
  assign n12822 = \PM_rd4[2]_pad  & n12488 ;
  assign n12830 = ~n12820 & ~n12822 ;
  assign n12833 = n12829 & n12830 ;
  assign n12834 = n12832 & n12833 ;
  assign n12835 = ~n12821 & n12834 ;
  assign n12836 = ~n12819 & ~n12835 ;
  assign n12837 = n12452 & n12836 ;
  assign n12838 = ~n12809 & ~n12837 ;
  assign n12839 = ~n12810 & n12838 ;
  assign n12840 = n12451 & ~n12839 ;
  assign n12841 = \bdma_BWdataBUF_reg[2]/P0001  & n12525 ;
  assign n12842 = ~n12840 & ~n12841 ;
  assign n12844 = n8113 & n12456 ;
  assign n12843 = \sice_idr0_reg_DO_reg[3]/P0001  & n12454 ;
  assign n12848 = ~n7916 & n12470 ;
  assign n12846 = ~n8000 & n12466 ;
  assign n12847 = ~n7967 & n12468 ;
  assign n12849 = ~n12846 & ~n12847 ;
  assign n12850 = ~n12848 & n12849 ;
  assign n12851 = ~\emc_PMDoe_reg/NET0131  & ~n12850 ;
  assign n12845 = \emc_PMDoe_reg/NET0131  & \emc_PMDreg_reg[3]/P0001  ;
  assign n12852 = n12465 & ~n12845 ;
  assign n12853 = ~n12851 & n12852 ;
  assign n12855 = \PM_rd0[3]_pad  & ~n12504 ;
  assign n12861 = \PM_rd5[3]_pad  & n12495 ;
  assign n12859 = \PM_rd3[3]_pad  & n12493 ;
  assign n12860 = \PM_rd1[3]_pad  & n12491 ;
  assign n12865 = ~n12859 & ~n12860 ;
  assign n12866 = ~n12861 & n12865 ;
  assign n12858 = \PM_rd7[3]_pad  & n12485 ;
  assign n12857 = \PM_rd6[3]_pad  & n12483 ;
  assign n12862 = ~n12465 & ~n12857 ;
  assign n12863 = ~n12858 & n12862 ;
  assign n12854 = \PM_rd2[3]_pad  & n12478 ;
  assign n12856 = \PM_rd4[3]_pad  & n12488 ;
  assign n12864 = ~n12854 & ~n12856 ;
  assign n12867 = n12863 & n12864 ;
  assign n12868 = n12866 & n12867 ;
  assign n12869 = ~n12855 & n12868 ;
  assign n12870 = ~n12853 & ~n12869 ;
  assign n12871 = n12452 & n12870 ;
  assign n12872 = ~n12843 & ~n12871 ;
  assign n12873 = ~n12844 & n12872 ;
  assign n12874 = n12451 & ~n12873 ;
  assign n12875 = \bdma_BWdataBUF_reg[3]/P0001  & n12525 ;
  assign n12876 = ~n12874 & ~n12875 ;
  assign n12878 = n10069 & n12456 ;
  assign n12877 = \sice_idr0_reg_DO_reg[4]/P0001  & n12454 ;
  assign n12882 = ~n9876 & n12470 ;
  assign n12880 = ~n9927 & n12468 ;
  assign n12881 = ~n9956 & n12466 ;
  assign n12883 = ~n12880 & ~n12881 ;
  assign n12884 = ~n12882 & n12883 ;
  assign n12885 = ~\emc_PMDoe_reg/NET0131  & ~n12884 ;
  assign n12879 = \emc_PMDoe_reg/NET0131  & \emc_PMDreg_reg[4]/P0001  ;
  assign n12886 = n12465 & ~n12879 ;
  assign n12887 = ~n12885 & n12886 ;
  assign n12889 = \PM_rd0[4]_pad  & ~n12504 ;
  assign n12895 = \PM_rd5[4]_pad  & n12495 ;
  assign n12893 = \PM_rd3[4]_pad  & n12493 ;
  assign n12894 = \PM_rd1[4]_pad  & n12491 ;
  assign n12899 = ~n12893 & ~n12894 ;
  assign n12900 = ~n12895 & n12899 ;
  assign n12892 = \PM_rd7[4]_pad  & n12485 ;
  assign n12891 = \PM_rd6[4]_pad  & n12483 ;
  assign n12896 = ~n12465 & ~n12891 ;
  assign n12897 = ~n12892 & n12896 ;
  assign n12888 = \PM_rd2[4]_pad  & n12478 ;
  assign n12890 = \PM_rd4[4]_pad  & n12488 ;
  assign n12898 = ~n12888 & ~n12890 ;
  assign n12901 = n12897 & n12898 ;
  assign n12902 = n12900 & n12901 ;
  assign n12903 = ~n12889 & n12902 ;
  assign n12904 = ~n12887 & ~n12903 ;
  assign n12905 = n12452 & n12904 ;
  assign n12906 = ~n12877 & ~n12905 ;
  assign n12907 = ~n12878 & n12906 ;
  assign n12908 = n12451 & ~n12907 ;
  assign n12909 = \bdma_BWdataBUF_reg[4]/P0001  & n12525 ;
  assign n12910 = ~n12908 & ~n12909 ;
  assign n12912 = n10911 & n12456 ;
  assign n12911 = \sice_idr0_reg_DO_reg[5]/P0001  & n12454 ;
  assign n12916 = ~n10889 & n12470 ;
  assign n12914 = ~n10709 & n12468 ;
  assign n12915 = ~n10806 & n12466 ;
  assign n12917 = ~n12914 & ~n12915 ;
  assign n12918 = ~n12916 & n12917 ;
  assign n12919 = ~\emc_PMDoe_reg/NET0131  & ~n12918 ;
  assign n12913 = \emc_PMDoe_reg/NET0131  & \emc_PMDreg_reg[5]/P0001  ;
  assign n12920 = n12465 & ~n12913 ;
  assign n12921 = ~n12919 & n12920 ;
  assign n12923 = \PM_rd0[5]_pad  & ~n12504 ;
  assign n12929 = \PM_rd5[5]_pad  & n12495 ;
  assign n12927 = \PM_rd3[5]_pad  & n12493 ;
  assign n12928 = \PM_rd1[5]_pad  & n12491 ;
  assign n12933 = ~n12927 & ~n12928 ;
  assign n12934 = ~n12929 & n12933 ;
  assign n12926 = \PM_rd7[5]_pad  & n12485 ;
  assign n12925 = \PM_rd6[5]_pad  & n12483 ;
  assign n12930 = ~n12465 & ~n12925 ;
  assign n12931 = ~n12926 & n12930 ;
  assign n12922 = \PM_rd2[5]_pad  & n12478 ;
  assign n12924 = \PM_rd4[5]_pad  & n12488 ;
  assign n12932 = ~n12922 & ~n12924 ;
  assign n12935 = n12931 & n12932 ;
  assign n12936 = n12934 & n12935 ;
  assign n12937 = ~n12923 & n12936 ;
  assign n12938 = ~n12921 & ~n12937 ;
  assign n12939 = n12452 & n12938 ;
  assign n12940 = ~n12911 & ~n12939 ;
  assign n12941 = ~n12912 & n12940 ;
  assign n12942 = n12451 & ~n12941 ;
  assign n12943 = \bdma_BWdataBUF_reg[5]/P0001  & n12525 ;
  assign n12944 = ~n12942 & ~n12943 ;
  assign n12946 = n11525 & n12456 ;
  assign n12945 = \sice_idr0_reg_DO_reg[6]/P0001  & n12454 ;
  assign n12949 = \PM_rd0[6]_pad  & ~n12504 ;
  assign n12954 = \PM_rd1[6]_pad  & n12491 ;
  assign n12951 = \PM_rd5[6]_pad  & n12495 ;
  assign n12953 = \PM_rd2[6]_pad  & n12478 ;
  assign n12958 = ~n12951 & ~n12953 ;
  assign n12959 = ~n12954 & n12958 ;
  assign n12952 = \PM_rd7[6]_pad  & n12485 ;
  assign n12947 = \PM_rd6[6]_pad  & n12483 ;
  assign n12955 = ~n12465 & ~n12947 ;
  assign n12956 = ~n12952 & n12955 ;
  assign n12948 = \PM_rd3[6]_pad  & n12493 ;
  assign n12950 = \PM_rd4[6]_pad  & n12488 ;
  assign n12957 = ~n12948 & ~n12950 ;
  assign n12960 = n12956 & n12957 ;
  assign n12961 = n12959 & n12960 ;
  assign n12962 = ~n12949 & n12961 ;
  assign n12965 = ~n11347 & n12468 ;
  assign n12964 = ~n11455 & n12470 ;
  assign n12966 = ~n11320 & n12466 ;
  assign n12967 = ~n12964 & ~n12966 ;
  assign n12968 = ~n12965 & n12967 ;
  assign n12969 = ~\emc_PMDoe_reg/NET0131  & ~n12968 ;
  assign n12963 = \emc_PMDoe_reg/NET0131  & \emc_PMDreg_reg[6]/P0001  ;
  assign n12970 = n12465 & ~n12963 ;
  assign n12971 = ~n12969 & n12970 ;
  assign n12972 = ~n12962 & ~n12971 ;
  assign n12973 = n12452 & n12972 ;
  assign n12974 = ~n12945 & ~n12973 ;
  assign n12975 = ~n12946 & n12974 ;
  assign n12976 = n12451 & ~n12975 ;
  assign n12977 = \bdma_BWdataBUF_reg[6]/P0001  & n12525 ;
  assign n12978 = ~n12976 & ~n12977 ;
  assign n12980 = n11265 & n12456 ;
  assign n12979 = \sice_idr0_reg_DO_reg[7]/P0001  & n12454 ;
  assign n12984 = ~n11203 & n12470 ;
  assign n12982 = ~n11077 & n12468 ;
  assign n12983 = ~n11243 & n12466 ;
  assign n12985 = ~n12982 & ~n12983 ;
  assign n12986 = ~n12984 & n12985 ;
  assign n12987 = ~\emc_PMDoe_reg/NET0131  & ~n12986 ;
  assign n12981 = \emc_PMDoe_reg/NET0131  & \emc_PMDreg_reg[7]/P0001  ;
  assign n12988 = n12465 & ~n12981 ;
  assign n12989 = ~n12987 & n12988 ;
  assign n12991 = \PM_rd0[7]_pad  & ~n12504 ;
  assign n12997 = \PM_rd5[7]_pad  & n12495 ;
  assign n12995 = \PM_rd3[7]_pad  & n12493 ;
  assign n12996 = \PM_rd1[7]_pad  & n12491 ;
  assign n13001 = ~n12995 & ~n12996 ;
  assign n13002 = ~n12997 & n13001 ;
  assign n12994 = \PM_rd7[7]_pad  & n12485 ;
  assign n12993 = \PM_rd6[7]_pad  & n12483 ;
  assign n12998 = ~n12465 & ~n12993 ;
  assign n12999 = ~n12994 & n12998 ;
  assign n12990 = \PM_rd2[7]_pad  & n12478 ;
  assign n12992 = \PM_rd4[7]_pad  & n12488 ;
  assign n13000 = ~n12990 & ~n12992 ;
  assign n13003 = n12999 & n13000 ;
  assign n13004 = n13002 & n13003 ;
  assign n13005 = ~n12991 & n13004 ;
  assign n13006 = ~n12989 & ~n13005 ;
  assign n13007 = n12452 & n13006 ;
  assign n13008 = ~n12979 & ~n13007 ;
  assign n13009 = ~n12980 & n13008 ;
  assign n13010 = n12451 & ~n13009 ;
  assign n13011 = \bdma_BWdataBUF_reg[7]/P0001  & n12525 ;
  assign n13012 = ~n13010 & ~n13011 ;
  assign n13013 = \bdma_BCTL_reg[9]/NET0131  & \bdma_BM_cyc_reg/P0001  ;
  assign n13015 = n10638 & n12456 ;
  assign n13014 = \sice_idr0_reg_DO_reg[8]/P0001  & n12454 ;
  assign n13019 = ~n10466 & n12468 ;
  assign n13017 = ~n10545 & n12470 ;
  assign n13018 = ~n10579 & n12466 ;
  assign n13020 = ~n13017 & ~n13018 ;
  assign n13021 = ~n13019 & n13020 ;
  assign n13022 = ~\emc_PMDoe_reg/NET0131  & ~n13021 ;
  assign n13016 = \emc_PMDoe_reg/NET0131  & \emc_PMDreg_reg[8]/P0001  ;
  assign n13023 = n12465 & ~n13016 ;
  assign n13024 = ~n13022 & n13023 ;
  assign n13026 = \PM_rd0[8]_pad  & ~n12504 ;
  assign n13032 = \PM_rd5[8]_pad  & n12495 ;
  assign n13030 = \PM_rd3[8]_pad  & n12493 ;
  assign n13031 = \PM_rd1[8]_pad  & n12491 ;
  assign n13036 = ~n13030 & ~n13031 ;
  assign n13037 = ~n13032 & n13036 ;
  assign n13029 = \PM_rd7[8]_pad  & n12485 ;
  assign n13028 = \PM_rd6[8]_pad  & n12483 ;
  assign n13033 = ~n12465 & ~n13028 ;
  assign n13034 = ~n13029 & n13033 ;
  assign n13025 = \PM_rd2[8]_pad  & n12478 ;
  assign n13027 = \PM_rd4[8]_pad  & n12488 ;
  assign n13035 = ~n13025 & ~n13027 ;
  assign n13038 = n13034 & n13035 ;
  assign n13039 = n13037 & n13038 ;
  assign n13040 = ~n13026 & n13039 ;
  assign n13041 = ~n13024 & ~n13040 ;
  assign n13042 = n12452 & n13041 ;
  assign n13043 = ~n13014 & ~n13042 ;
  assign n13044 = ~n13015 & n13043 ;
  assign n13045 = n12451 & ~n13044 ;
  assign n13046 = ~n13013 & ~n13045 ;
  assign n13047 = \bdma_BCTL_reg[10]/NET0131  & \bdma_BM_cyc_reg/P0001  ;
  assign n13049 = n10289 & n12456 ;
  assign n13048 = \sice_idr0_reg_DO_reg[9]/P0001  & n12454 ;
  assign n13053 = ~n10196 & n12468 ;
  assign n13051 = ~n10123 & n12470 ;
  assign n13052 = ~n10230 & n12466 ;
  assign n13054 = ~n13051 & ~n13052 ;
  assign n13055 = ~n13053 & n13054 ;
  assign n13056 = ~\emc_PMDoe_reg/NET0131  & ~n13055 ;
  assign n13050 = \emc_PMDoe_reg/NET0131  & \emc_PMDreg_reg[9]/P0001  ;
  assign n13057 = n12465 & ~n13050 ;
  assign n13058 = ~n13056 & n13057 ;
  assign n13060 = \PM_rd0[9]_pad  & ~n12504 ;
  assign n13066 = \PM_rd5[9]_pad  & n12495 ;
  assign n13064 = \PM_rd3[9]_pad  & n12493 ;
  assign n13065 = \PM_rd1[9]_pad  & n12491 ;
  assign n13070 = ~n13064 & ~n13065 ;
  assign n13071 = ~n13066 & n13070 ;
  assign n13063 = \PM_rd7[9]_pad  & n12485 ;
  assign n13062 = \PM_rd6[9]_pad  & n12483 ;
  assign n13067 = ~n12465 & ~n13062 ;
  assign n13068 = ~n13063 & n13067 ;
  assign n13059 = \PM_rd2[9]_pad  & n12478 ;
  assign n13061 = \PM_rd4[9]_pad  & n12488 ;
  assign n13069 = ~n13059 & ~n13061 ;
  assign n13072 = n13068 & n13069 ;
  assign n13073 = n13071 & n13072 ;
  assign n13074 = ~n13060 & n13073 ;
  assign n13075 = ~n13058 & ~n13074 ;
  assign n13076 = n12452 & n13075 ;
  assign n13077 = ~n13048 & ~n13076 ;
  assign n13078 = ~n13049 & n13077 ;
  assign n13079 = n12451 & ~n13078 ;
  assign n13080 = ~n13047 & ~n13079 ;
  assign n13081 = ~\bdma_BM_cyc_reg/P0001  & ~n12451 ;
  assign n13082 = ~n12451 & ~n12525 ;
  assign n13083 = ~\idma_DCTL_reg[14]/NET0131  & ~\idma_PCrd_1st_reg/NET0131  ;
  assign n13085 = ~\idma_DTMP_L_reg[0]/P0001  & n13083 ;
  assign n13084 = ~\idma_DTMP_H_reg[0]/P0001  & ~n13083 ;
  assign n13086 = ~\core_c_psq_PCS_reg[3]/NET0131  & ~n13084 ;
  assign n13087 = ~n13085 & n13086 ;
  assign n13088 = \idma_DTMP_H_reg[10]/P0001  & ~n13083 ;
  assign n13089 = ~\core_c_psq_PCS_reg[3]/NET0131  & ~n13088 ;
  assign n13090 = ~\core_c_psq_PCS_reg[3]/NET0131  & ~n13083 ;
  assign n13091 = \idma_DTMP_H_reg[11]/P0001  & n13090 ;
  assign n13092 = \idma_DTMP_H_reg[12]/P0001  & n13090 ;
  assign n13093 = \idma_DTMP_H_reg[13]/P0001  & ~n13083 ;
  assign n13094 = ~\core_c_psq_PCS_reg[3]/NET0131  & ~n13093 ;
  assign n13095 = \idma_DTMP_H_reg[14]/P0001  & n13090 ;
  assign n13096 = \idma_DTMP_H_reg[15]/P0001  & ~n13083 ;
  assign n13097 = ~\core_c_psq_PCS_reg[3]/NET0131  & ~n13096 ;
  assign n13099 = ~\idma_DTMP_L_reg[1]/P0001  & n13083 ;
  assign n13098 = ~\idma_DTMP_H_reg[1]/P0001  & ~n13083 ;
  assign n13100 = ~\core_c_psq_PCS_reg[3]/NET0131  & ~n13098 ;
  assign n13101 = ~n13099 & n13100 ;
  assign n13103 = \idma_DTMP_H_reg[2]/P0001  & ~n13083 ;
  assign n13102 = \idma_DTMP_L_reg[2]/P0001  & n13083 ;
  assign n13104 = ~\core_c_psq_PCS_reg[3]/NET0131  & ~n13102 ;
  assign n13105 = ~n13103 & n13104 ;
  assign n13107 = ~\idma_DTMP_L_reg[3]/P0001  & n13083 ;
  assign n13106 = ~\idma_DTMP_H_reg[3]/P0001  & ~n13083 ;
  assign n13108 = ~\core_c_psq_PCS_reg[3]/NET0131  & ~n13106 ;
  assign n13109 = ~n13107 & n13108 ;
  assign n13111 = ~\idma_DTMP_L_reg[4]/P0001  & n13083 ;
  assign n13110 = ~\idma_DTMP_H_reg[4]/P0001  & ~n13083 ;
  assign n13112 = ~\core_c_psq_PCS_reg[3]/NET0131  & ~n13110 ;
  assign n13113 = ~n13111 & n13112 ;
  assign n13115 = \idma_DTMP_H_reg[5]/P0001  & ~n13083 ;
  assign n13114 = \idma_DTMP_L_reg[5]/P0001  & n13083 ;
  assign n13116 = ~\core_c_psq_PCS_reg[3]/NET0131  & ~n13114 ;
  assign n13117 = ~n13115 & n13116 ;
  assign n13119 = ~\idma_DTMP_L_reg[6]/P0001  & n13083 ;
  assign n13118 = ~\idma_DTMP_H_reg[6]/P0001  & ~n13083 ;
  assign n13120 = ~\core_c_psq_PCS_reg[3]/NET0131  & ~n13118 ;
  assign n13121 = ~n13119 & n13120 ;
  assign n13123 = \idma_DTMP_H_reg[7]/P0001  & ~n13083 ;
  assign n13122 = \idma_DTMP_L_reg[7]/P0001  & n13083 ;
  assign n13124 = ~\core_c_psq_PCS_reg[3]/NET0131  & ~n13122 ;
  assign n13125 = ~n13123 & n13124 ;
  assign n13126 = \idma_DTMP_H_reg[8]/P0001  & n13090 ;
  assign n13127 = \idma_DTMP_H_reg[9]/P0001  & n13090 ;
  assign n13128 = ~\idma_RDCMD_reg/P0001  & ~\idma_RDcyc_reg/NET0131  ;
  assign n13129 = ~T_IMS_pad & \sice_OE_reg/P0001  ;
  assign n13130 = ~\memc_EXTC_E_reg/NET0131  & \memc_Pwrite_E_reg/NET0131  ;
  assign n13131 = ~\core_c_dec_Dummy_E_reg/NET0131  & n13130 ;
  assign n13132 = ~n4099 & ~n13131 ;
  assign n13133 = ~n4117 & n13132 ;
  assign n13134 = n6020 & ~n13133 ;
  assign n13135 = n6047 & n13133 ;
  assign n13136 = ~n5936 & ~n13133 ;
  assign n13137 = ~n13135 & ~n13136 ;
  assign n13138 = n6164 & n13137 ;
  assign n13139 = ~n13134 & n13138 ;
  assign n13141 = n6911 & n13137 ;
  assign n13140 = n6980 & n13135 ;
  assign n13142 = ~n13134 & ~n13136 ;
  assign n13143 = ~n13140 & n13142 ;
  assign n13144 = ~n13141 & n13143 ;
  assign n13145 = \bdma_CMcnt_reg[0]/NET0131  & ~\bdma_CMcnt_reg[1]/NET0131  ;
  assign n13146 = n5730 & n13145 ;
  assign n13147 = n5727 & n13146 ;
  assign n13148 = ~\bdma_BCTL_reg[2]/NET0131  & n13147 ;
  assign n13149 = ~\bdma_CMcnt_reg[0]/NET0131  & ~\bdma_CMcnt_reg[1]/NET0131  ;
  assign n13150 = n5730 & n13149 ;
  assign n13151 = \bdma_BCTL_reg[2]/NET0131  & n13150 ;
  assign n13152 = n5727 & n13151 ;
  assign n13153 = ~n13148 & ~n13152 ;
  assign n13154 = n6913 & ~n13153 ;
  assign n13156 = ~n4099 & n13130 ;
  assign n13157 = n6931 & n13156 ;
  assign n13158 = n6930 & ~n13157 ;
  assign n13159 = \core_dag_ilm2reg_PMA_pi_DO_reg[0]/NET0131  & ~n13158 ;
  assign n13160 = ~n5717 & n5880 ;
  assign n13161 = \idma_DCTL_reg[0]/NET0131  & n13160 ;
  assign n13162 = ~n6989 & ~n13161 ;
  assign n13163 = ~n13159 & n13162 ;
  assign n13164 = ~n13154 & ~n13163 ;
  assign n13155 = \bdma_BIAD_reg[0]/NET0131  & n13154 ;
  assign n13165 = ~n13137 & ~n13155 ;
  assign n13166 = ~n13164 & n13165 ;
  assign n13167 = n6968 & n13137 ;
  assign n13168 = ~n13142 & ~n13167 ;
  assign n13169 = ~n13166 & n13168 ;
  assign n13170 = ~n13144 & ~n13169 ;
  assign n13171 = ~n13139 & ~n13170 ;
  assign n13172 = n7607 & n13139 ;
  assign n13173 = ~n13171 & ~n13172 ;
  assign n13175 = n8211 & n13137 ;
  assign n13174 = n8121 & n13135 ;
  assign n13176 = n13142 & ~n13174 ;
  assign n13177 = ~n13175 & n13176 ;
  assign n13179 = \core_dag_ilm2reg_PMA_pi_DO_reg[10]/NET0131  & ~n13158 ;
  assign n13180 = \idma_DCTL_reg[10]/NET0131  & n13160 ;
  assign n13181 = ~n8160 & ~n13180 ;
  assign n13182 = ~n13179 & n13181 ;
  assign n13183 = ~n13154 & ~n13182 ;
  assign n13178 = \bdma_BIAD_reg[10]/NET0131  & n13154 ;
  assign n13184 = ~n13137 & ~n13178 ;
  assign n13185 = ~n13183 & n13184 ;
  assign n13186 = n8129 & n13137 ;
  assign n13187 = ~n13142 & ~n13186 ;
  assign n13188 = ~n13185 & n13187 ;
  assign n13189 = ~n13177 & ~n13188 ;
  assign n13190 = ~n13139 & ~n13189 ;
  assign n13191 = n7859 & n13139 ;
  assign n13192 = ~n13190 & ~n13191 ;
  assign n13194 = n8813 & n13137 ;
  assign n13193 = n8723 & n13135 ;
  assign n13195 = n13142 & ~n13193 ;
  assign n13196 = ~n13194 & n13195 ;
  assign n13198 = \core_dag_ilm2reg_PMA_pi_DO_reg[11]/NET0131  & ~n13158 ;
  assign n13199 = \idma_DCTL_reg[11]/NET0131  & n13160 ;
  assign n13200 = ~n8816 & ~n13199 ;
  assign n13201 = ~n13198 & n13200 ;
  assign n13202 = ~n13154 & ~n13201 ;
  assign n13197 = \bdma_BIAD_reg[11]/NET0131  & n13154 ;
  assign n13203 = ~n13137 & ~n13197 ;
  assign n13204 = ~n13202 & n13203 ;
  assign n13205 = n8731 & n13137 ;
  assign n13206 = ~n13142 & ~n13205 ;
  assign n13207 = ~n13204 & n13206 ;
  assign n13208 = ~n13196 & ~n13207 ;
  assign n13209 = ~n13139 & ~n13208 ;
  assign n13210 = n8460 & n13139 ;
  assign n13211 = ~n13209 & ~n13210 ;
  assign n13213 = n9559 & n13137 ;
  assign n13212 = n9528 & n13135 ;
  assign n13214 = n13142 & ~n13212 ;
  assign n13215 = ~n13213 & n13214 ;
  assign n13217 = \core_dag_ilm2reg_PMA_pi_DO_reg[1]/NET0131  & ~n13158 ;
  assign n13218 = \idma_DCTL_reg[1]/NET0131  & n13160 ;
  assign n13219 = ~n9564 & ~n13218 ;
  assign n13220 = ~n13217 & n13219 ;
  assign n13221 = ~n13154 & ~n13220 ;
  assign n13216 = \bdma_BIAD_reg[1]/NET0131  & n13154 ;
  assign n13222 = ~n13137 & ~n13216 ;
  assign n13223 = ~n13221 & n13222 ;
  assign n13224 = n9520 & n13137 ;
  assign n13225 = ~n13142 & ~n13224 ;
  assign n13226 = ~n13223 & n13225 ;
  assign n13227 = ~n13215 & ~n13226 ;
  assign n13228 = ~n13139 & ~n13227 ;
  assign n13229 = n9435 & n13139 ;
  assign n13230 = ~n13228 & ~n13229 ;
  assign n13232 = n9625 & n13137 ;
  assign n13231 = n9600 & n13135 ;
  assign n13233 = n13142 & ~n13231 ;
  assign n13234 = ~n13232 & n13233 ;
  assign n13236 = \core_dag_ilm2reg_PMA_pi_DO_reg[2]/NET0131  & ~n13158 ;
  assign n13237 = \idma_DCTL_reg[2]/NET0131  & n13160 ;
  assign n13238 = ~n9630 & ~n13237 ;
  assign n13239 = ~n13236 & n13238 ;
  assign n13240 = ~n13154 & ~n13239 ;
  assign n13235 = \bdma_BIAD_reg[2]/NET0131  & n13154 ;
  assign n13241 = ~n13137 & ~n13235 ;
  assign n13242 = ~n13240 & n13241 ;
  assign n13243 = n9592 & n13137 ;
  assign n13244 = ~n13142 & ~n13243 ;
  assign n13245 = ~n13242 & n13244 ;
  assign n13246 = ~n13234 & ~n13245 ;
  assign n13247 = ~n13139 & ~n13246 ;
  assign n13248 = n8715 & n13139 ;
  assign n13249 = ~n13247 & ~n13248 ;
  assign n13251 = \core_dag_ilm2reg_PMA_pi_DO_reg[3]/NET0131  & ~n13158 ;
  assign n13252 = \idma_DCTL_reg[3]/NET0131  & n13160 ;
  assign n13253 = ~n9705 & ~n13252 ;
  assign n13254 = ~n13251 & n13253 ;
  assign n13255 = ~n13154 & ~n13254 ;
  assign n13250 = \bdma_BIAD_reg[3]/NET0131  & n13154 ;
  assign n13256 = n13136 & ~n13250 ;
  assign n13257 = ~n13255 & n13256 ;
  assign n13259 = ~n9658 & n13134 ;
  assign n13260 = n6164 & ~n8113 ;
  assign n13261 = ~n6164 & n9695 ;
  assign n13262 = ~n13260 & ~n13261 ;
  assign n13263 = ~n13134 & n13262 ;
  assign n13264 = ~n13259 & ~n13263 ;
  assign n13265 = ~n13135 & ~n13264 ;
  assign n13258 = ~n9666 & n13135 ;
  assign n13266 = ~n13136 & ~n13258 ;
  assign n13267 = ~n13265 & n13266 ;
  assign n13268 = ~n13257 & ~n13267 ;
  assign n13271 = ~n6164 & n9767 ;
  assign n13272 = ~n13134 & n13271 ;
  assign n13270 = n9797 & n13134 ;
  assign n13273 = ~n13135 & ~n13270 ;
  assign n13274 = ~n13272 & n13273 ;
  assign n13275 = ~n9805 & n13135 ;
  assign n13276 = ~n13136 & ~n13275 ;
  assign n13277 = ~n13274 & n13276 ;
  assign n13269 = ~n10069 & n13139 ;
  assign n13279 = \core_dag_ilm2reg_PMA_pi_DO_reg[4]/NET0131  & ~n13158 ;
  assign n13280 = \idma_DCTL_reg[4]/NET0131  & n13160 ;
  assign n13281 = ~n9812 & ~n13280 ;
  assign n13282 = ~n13279 & n13281 ;
  assign n13283 = ~n13154 & ~n13282 ;
  assign n13278 = \bdma_BIAD_reg[4]/NET0131  & n13154 ;
  assign n13284 = n13136 & ~n13278 ;
  assign n13285 = ~n13283 & n13284 ;
  assign n13286 = ~n13269 & ~n13285 ;
  assign n13287 = ~n13277 & n13286 ;
  assign n13290 = ~n6164 & n10324 ;
  assign n13291 = ~n13134 & n13290 ;
  assign n13289 = n10364 & n13134 ;
  assign n13292 = ~n13135 & ~n13289 ;
  assign n13293 = ~n13291 & n13292 ;
  assign n13294 = ~n10356 & n13135 ;
  assign n13295 = ~n13136 & ~n13294 ;
  assign n13296 = ~n13293 & n13295 ;
  assign n13288 = ~n10911 & n13139 ;
  assign n13298 = \core_dag_ilm2reg_PMA_pi_DO_reg[5]/NET0131  & ~n13158 ;
  assign n13299 = \idma_DCTL_reg[5]/NET0131  & n13160 ;
  assign n13300 = ~n10349 & ~n13299 ;
  assign n13301 = ~n13298 & n13300 ;
  assign n13302 = ~n13154 & ~n13301 ;
  assign n13297 = \bdma_BIAD_reg[5]/NET0131  & n13154 ;
  assign n13303 = n13136 & ~n13297 ;
  assign n13304 = ~n13302 & n13303 ;
  assign n13305 = ~n13288 & ~n13304 ;
  assign n13306 = ~n13296 & n13305 ;
  assign n13309 = ~n6164 & n10930 ;
  assign n13310 = ~n13134 & n13309 ;
  assign n13308 = n10975 & n13134 ;
  assign n13311 = ~n13135 & ~n13308 ;
  assign n13312 = ~n13310 & n13311 ;
  assign n13313 = ~n10967 & n13135 ;
  assign n13314 = ~n13136 & ~n13313 ;
  assign n13315 = ~n13312 & n13314 ;
  assign n13307 = ~n11525 & n13139 ;
  assign n13317 = \core_dag_ilm2reg_PMA_pi_DO_reg[6]/NET0131  & ~n13158 ;
  assign n13318 = \idma_DCTL_reg[6]/NET0131  & n13160 ;
  assign n13319 = ~n10960 & ~n13318 ;
  assign n13320 = ~n13317 & n13319 ;
  assign n13321 = ~n13154 & ~n13320 ;
  assign n13316 = \bdma_BIAD_reg[6]/NET0131  & n13154 ;
  assign n13322 = n13136 & ~n13316 ;
  assign n13323 = ~n13321 & n13322 ;
  assign n13324 = ~n13307 & ~n13323 ;
  assign n13325 = ~n13315 & n13324 ;
  assign n13328 = ~n6164 & n11579 ;
  assign n13329 = ~n13134 & n13328 ;
  assign n13327 = n11548 & n13134 ;
  assign n13330 = ~n13135 & ~n13327 ;
  assign n13331 = ~n13329 & n13330 ;
  assign n13332 = ~n11540 & n13135 ;
  assign n13333 = ~n13136 & ~n13332 ;
  assign n13334 = ~n13331 & n13333 ;
  assign n13326 = ~n11265 & n13139 ;
  assign n13336 = \core_dag_ilm2reg_PMA_pi_DO_reg[7]/NET0131  & ~n13158 ;
  assign n13337 = \idma_DCTL_reg[7]/NET0131  & n13160 ;
  assign n13338 = ~n11532 & ~n13337 ;
  assign n13339 = ~n13336 & n13338 ;
  assign n13340 = ~n13154 & ~n13339 ;
  assign n13335 = \bdma_BIAD_reg[7]/NET0131  & n13154 ;
  assign n13341 = n13136 & ~n13335 ;
  assign n13342 = ~n13340 & n13341 ;
  assign n13343 = ~n13326 & ~n13342 ;
  assign n13344 = ~n13334 & n13343 ;
  assign n13347 = ~n6164 & n11654 ;
  assign n13348 = ~n13134 & n13347 ;
  assign n13346 = n11617 & n13134 ;
  assign n13349 = ~n13135 & ~n13346 ;
  assign n13350 = ~n13348 & n13349 ;
  assign n13351 = ~n11609 & n13135 ;
  assign n13352 = ~n13136 & ~n13351 ;
  assign n13353 = ~n13350 & n13352 ;
  assign n13345 = ~n10638 & n13139 ;
  assign n13355 = \core_dag_ilm2reg_PMA_pi_DO_reg[8]/NET0131  & ~n13158 ;
  assign n13356 = \idma_DCTL_reg[8]/NET0131  & n13160 ;
  assign n13357 = ~n11625 & ~n13356 ;
  assign n13358 = ~n13355 & n13357 ;
  assign n13359 = ~n13154 & ~n13358 ;
  assign n13354 = \bdma_BIAD_reg[8]/NET0131  & n13154 ;
  assign n13360 = n13136 & ~n13354 ;
  assign n13361 = ~n13359 & n13360 ;
  assign n13362 = ~n13345 & ~n13361 ;
  assign n13363 = ~n13353 & n13362 ;
  assign n13366 = ~n6164 & n11720 ;
  assign n13367 = ~n13134 & n13366 ;
  assign n13365 = n11676 & n13134 ;
  assign n13368 = ~n13135 & ~n13365 ;
  assign n13369 = ~n13367 & n13368 ;
  assign n13370 = ~n11668 & n13135 ;
  assign n13371 = ~n13136 & ~n13370 ;
  assign n13372 = ~n13369 & n13371 ;
  assign n13364 = ~n10289 & n13139 ;
  assign n13374 = \core_dag_ilm2reg_PMA_pi_DO_reg[9]/NET0131  & ~n13158 ;
  assign n13375 = \idma_DCTL_reg[9]/NET0131  & n13160 ;
  assign n13376 = ~n11687 & ~n13375 ;
  assign n13377 = ~n13374 & n13376 ;
  assign n13378 = ~n13154 & ~n13377 ;
  assign n13373 = \bdma_BIAD_reg[9]/NET0131  & n13154 ;
  assign n13379 = n13136 & ~n13373 ;
  assign n13380 = ~n13378 & n13379 ;
  assign n13381 = ~n13364 & ~n13380 ;
  assign n13382 = ~n13372 & n13381 ;
  assign n13383 = n5880 & n5882 ;
  assign n13384 = n11761 & n13383 ;
  assign n13385 = n6913 & n13148 ;
  assign n13386 = ~n7362 & n12473 ;
  assign n13387 = ~n13385 & n13386 ;
  assign n13388 = ~\bdma_BRdataBUF_reg[8]/P0001  & n13385 ;
  assign n13389 = ~n13387 & ~n13388 ;
  assign n13390 = ~n13384 & ~n13389 ;
  assign n13391 = ~\idma_DTMP_H_reg[0]/P0001  & n13384 ;
  assign n13392 = ~n13390 & ~n13391 ;
  assign n13393 = ~n7664 & n12536 ;
  assign n13394 = ~n13385 & n13393 ;
  assign n13395 = ~\bdma_BRdataBUF_reg[18]/P0001  & n13385 ;
  assign n13396 = ~n13394 & ~n13395 ;
  assign n13397 = ~n13384 & ~n13396 ;
  assign n13398 = ~\idma_DTMP_H_reg[10]/P0001  & n13384 ;
  assign n13399 = ~n13397 & ~n13398 ;
  assign n13400 = ~n8266 & n12570 ;
  assign n13401 = ~n13385 & n13400 ;
  assign n13402 = ~\bdma_BRdataBUF_reg[19]/P0001  & n13385 ;
  assign n13403 = ~n13401 & ~n13402 ;
  assign n13404 = ~n13384 & ~n13403 ;
  assign n13405 = ~\idma_DTMP_H_reg[11]/P0001  & n13384 ;
  assign n13406 = ~n13404 & ~n13405 ;
  assign n13407 = ~n8983 & n12604 ;
  assign n13408 = ~n13385 & n13407 ;
  assign n13409 = ~\bdma_BRdataBUF_reg[20]/P0001  & n13385 ;
  assign n13410 = ~n13408 & ~n13409 ;
  assign n13411 = ~n13384 & ~n13410 ;
  assign n13412 = ~\idma_DTMP_H_reg[12]/P0001  & n13384 ;
  assign n13413 = ~n13411 & ~n13412 ;
  assign n13414 = ~n7067 & n12638 ;
  assign n13415 = ~n13385 & n13414 ;
  assign n13416 = ~\bdma_BRdataBUF_reg[21]/P0001  & n13385 ;
  assign n13417 = ~n13415 & ~n13416 ;
  assign n13418 = ~n13384 & ~n13417 ;
  assign n13419 = ~\idma_DTMP_H_reg[13]/P0001  & n13384 ;
  assign n13420 = ~n13418 & ~n13419 ;
  assign n13421 = ~n11818 & n12695 ;
  assign n13422 = ~n13385 & n13421 ;
  assign n13423 = ~\bdma_BRdataBUF_reg[22]/P0001  & n13385 ;
  assign n13424 = ~n13422 & ~n13423 ;
  assign n13425 = ~n13384 & ~n13424 ;
  assign n13426 = ~\idma_DTMP_H_reg[14]/P0001  & n13384 ;
  assign n13427 = ~n13425 & ~n13426 ;
  assign n13428 = ~n11964 & n12751 ;
  assign n13429 = ~n13385 & n13428 ;
  assign n13430 = ~\bdma_BRdataBUF_reg[23]/P0001  & n13385 ;
  assign n13431 = ~n13429 & ~n13430 ;
  assign n13432 = ~n13384 & ~n13431 ;
  assign n13433 = ~\idma_DTMP_H_reg[15]/P0001  & n13384 ;
  assign n13434 = ~n13432 & ~n13433 ;
  assign n13435 = ~n9202 & n12782 ;
  assign n13436 = ~n13385 & n13435 ;
  assign n13437 = ~\bdma_BRdataBUF_reg[9]/P0001  & n13385 ;
  assign n13438 = ~n13436 & ~n13437 ;
  assign n13439 = ~n13384 & ~n13438 ;
  assign n13440 = ~\idma_DTMP_H_reg[1]/P0001  & n13384 ;
  assign n13441 = ~n13439 & ~n13440 ;
  assign n13442 = ~n8482 & n12816 ;
  assign n13443 = ~n13385 & n13442 ;
  assign n13444 = ~\bdma_BRdataBUF_reg[10]/P0001  & n13385 ;
  assign n13445 = ~n13443 & ~n13444 ;
  assign n13446 = ~n13384 & ~n13445 ;
  assign n13447 = ~\idma_DTMP_H_reg[2]/P0001  & n13384 ;
  assign n13448 = ~n13446 & ~n13447 ;
  assign n13449 = ~n7882 & n12850 ;
  assign n13450 = ~n13385 & n13449 ;
  assign n13451 = ~\bdma_BRdataBUF_reg[11]/P0001  & n13385 ;
  assign n13452 = ~n13450 & ~n13451 ;
  assign n13453 = ~n13384 & ~n13452 ;
  assign n13454 = ~\idma_DTMP_H_reg[3]/P0001  & n13384 ;
  assign n13455 = ~n13453 & ~n13454 ;
  assign n13456 = ~n9842 & n12884 ;
  assign n13457 = ~n13385 & n13456 ;
  assign n13458 = ~\bdma_BRdataBUF_reg[12]/P0001  & n13385 ;
  assign n13459 = ~n13457 & ~n13458 ;
  assign n13460 = ~n13384 & ~n13459 ;
  assign n13461 = ~\idma_DTMP_H_reg[4]/P0001  & n13384 ;
  assign n13462 = ~n13460 & ~n13461 ;
  assign n13463 = ~n10683 & n12918 ;
  assign n13464 = ~n13385 & n13463 ;
  assign n13465 = ~\bdma_BRdataBUF_reg[13]/P0001  & n13385 ;
  assign n13466 = ~n13464 & ~n13465 ;
  assign n13467 = ~n13384 & ~n13466 ;
  assign n13468 = ~\idma_DTMP_H_reg[5]/P0001  & n13384 ;
  assign n13469 = ~n13467 & ~n13468 ;
  assign n13470 = ~n11300 & n12968 ;
  assign n13471 = ~n13385 & n13470 ;
  assign n13472 = ~\bdma_BRdataBUF_reg[14]/P0001  & n13385 ;
  assign n13473 = ~n13471 & ~n13472 ;
  assign n13474 = ~n13384 & ~n13473 ;
  assign n13475 = ~\idma_DTMP_H_reg[6]/P0001  & n13384 ;
  assign n13476 = ~n13474 & ~n13475 ;
  assign n13477 = ~n11051 & n12986 ;
  assign n13478 = ~n13385 & n13477 ;
  assign n13479 = ~\bdma_BRdataBUF_reg[15]/P0001  & n13385 ;
  assign n13480 = ~n13478 & ~n13479 ;
  assign n13481 = ~n13384 & ~n13480 ;
  assign n13482 = ~\idma_DTMP_H_reg[7]/P0001  & n13384 ;
  assign n13483 = ~n13481 & ~n13482 ;
  assign n13484 = ~n10442 & n13021 ;
  assign n13485 = ~n13385 & n13484 ;
  assign n13486 = ~\bdma_BRdataBUF_reg[16]/P0001  & n13385 ;
  assign n13487 = ~n13485 & ~n13486 ;
  assign n13488 = ~n13384 & ~n13487 ;
  assign n13489 = ~\idma_DTMP_H_reg[8]/P0001  & n13384 ;
  assign n13490 = ~n13488 & ~n13489 ;
  assign n13491 = ~n10093 & n13055 ;
  assign n13492 = ~n13385 & n13491 ;
  assign n13493 = ~\bdma_BRdataBUF_reg[17]/P0001  & n13385 ;
  assign n13494 = ~n13492 & ~n13493 ;
  assign n13495 = ~n13384 & ~n13494 ;
  assign n13496 = ~\idma_DTMP_H_reg[9]/P0001  & n13384 ;
  assign n13497 = ~n13495 & ~n13496 ;
  assign n13509 = n8945 & n13137 ;
  assign n13510 = ~n13138 & n13142 ;
  assign n13511 = n8845 & ~n13137 ;
  assign n13512 = n13510 & ~n13511 ;
  assign n13513 = ~n13509 & n13512 ;
  assign n13498 = n9178 & n13139 ;
  assign n13499 = n5936 & n13134 ;
  assign n13500 = ~n8853 & n13499 ;
  assign n13502 = \core_dag_ilm2reg_PMA_pi_DO_reg[12]/NET0131  & ~n13158 ;
  assign n13503 = \idma_DCTL_reg[12]/NET0131  & n13160 ;
  assign n13504 = ~n8838 & ~n13503 ;
  assign n13505 = ~n13154 & n13504 ;
  assign n13506 = ~n13502 & n13505 ;
  assign n13501 = ~\bdma_BIAD_reg[12]/NET0131  & n13154 ;
  assign n13507 = n13136 & ~n13501 ;
  assign n13508 = ~n13506 & n13507 ;
  assign n13514 = ~n13500 & ~n13508 ;
  assign n13515 = ~n13498 & n13514 ;
  assign n13516 = ~n13513 & n13515 ;
  assign n13517 = ~PM_bdry_sel_pad & n13516 ;
  assign n13528 = n9497 & n13137 ;
  assign n13529 = n9452 & ~n13137 ;
  assign n13530 = n13510 & ~n13529 ;
  assign n13531 = ~n13528 & n13530 ;
  assign n13518 = n7340 & n13139 ;
  assign n13519 = ~n9460 & n13499 ;
  assign n13521 = \core_dag_ilm2reg_PMA_pi_DO_reg[13]/NET0131  & ~n13158 ;
  assign n13522 = \idma_DCTL_reg[13]/NET0131  & n13160 ;
  assign n13523 = ~n9442 & ~n13522 ;
  assign n13524 = ~n13154 & n13523 ;
  assign n13525 = ~n13521 & n13524 ;
  assign n13520 = ~\bdma_BIAD_reg[13]/NET0131  & n13154 ;
  assign n13526 = n13136 & ~n13520 ;
  assign n13527 = ~n13525 & n13526 ;
  assign n13532 = ~n13519 & ~n13527 ;
  assign n13533 = ~n13518 & n13532 ;
  assign n13534 = ~n13531 & n13533 ;
  assign n13535 = ~n13517 & ~n13534 ;
  assign n13536 = \core_c_psq_PMOVL_regh_DO_reg[1]/NET0131  & ~n5066 ;
  assign n13537 = \bdma_BOVL_reg[9]/NET0131  & n5066 ;
  assign n13538 = ~n13536 & ~n13537 ;
  assign n13539 = ~n5895 & ~n13538 ;
  assign n13540 = \idma_DOVL_reg[9]/NET0131  & n5895 ;
  assign n13541 = ~n13539 & ~n13540 ;
  assign n13542 = n13535 & n13541 ;
  assign n13543 = \core_c_psq_PMOVL_regh_DO_reg[3]/NET0131  & ~n5066 ;
  assign n13544 = \bdma_BOVL_reg[11]/NET0131  & n5066 ;
  assign n13545 = ~n13543 & ~n13544 ;
  assign n13546 = ~n5895 & ~n13545 ;
  assign n13547 = \idma_DOVL_reg[11]/NET0131  & n5895 ;
  assign n13548 = ~n13546 & ~n13547 ;
  assign n13549 = \core_c_psq_PMOVL_regh_DO_reg[2]/NET0131  & ~n5066 ;
  assign n13550 = \bdma_BOVL_reg[10]/NET0131  & n5066 ;
  assign n13551 = ~n13549 & ~n13550 ;
  assign n13552 = ~n5895 & ~n13551 ;
  assign n13553 = \idma_DOVL_reg[10]/NET0131  & n5895 ;
  assign n13554 = ~n13552 & ~n13553 ;
  assign n13555 = n13548 & n13554 ;
  assign n13556 = \core_c_psq_PMOVL_regh_DO_reg[0]/NET0131  & ~n5066 ;
  assign n13557 = \bdma_BOVL_reg[8]/NET0131  & n5066 ;
  assign n13558 = ~n13556 & ~n13557 ;
  assign n13559 = ~n5895 & ~n13558 ;
  assign n13560 = \idma_DOVL_reg[8]/NET0131  & n5895 ;
  assign n13561 = ~n13559 & ~n13560 ;
  assign n13562 = n13555 & n13561 ;
  assign n13563 = n13542 & n13562 ;
  assign n13574 = \core_c_dec_IR_reg[17]/NET0131  & n6119 ;
  assign n13575 = ~\core_c_dec_IR_reg[15]/NET0131  & n13574 ;
  assign n13576 = ~\core_c_dec_IR_reg[21]/NET0131  & \core_c_dec_IR_reg[22]/NET0131  ;
  assign n13577 = n6026 & n13576 ;
  assign n13578 = ~\core_c_dec_IR_reg[19]/NET0131  & n13577 ;
  assign n13579 = ~n6023 & ~n13578 ;
  assign n13580 = ~n13575 & n13579 ;
  assign n13581 = n11742 & ~n13580 ;
  assign n13582 = n13132 & n13581 ;
  assign n13568 = n5066 & n13152 ;
  assign n13569 = ~\idma_DCTL_reg[14]/NET0131  & \idma_RDcyc_reg/NET0131  ;
  assign n13570 = n5882 & n13569 ;
  assign n13571 = n5068 & n13570 ;
  assign n13572 = ~n13568 & ~n13571 ;
  assign n13573 = ~n5718 & ~n13572 ;
  assign n13583 = \memc_Pread_E_reg/NET0131  & n4117 ;
  assign n13584 = ~n13573 & ~n13583 ;
  assign n13585 = ~n13582 & n13584 ;
  assign n13564 = ~n13384 & ~n13385 ;
  assign n13565 = \memc_Pwrite_C_reg/NET0131  & n5950 ;
  assign n13566 = ~n5950 & n13156 ;
  assign n13567 = ~n13565 & ~n13566 ;
  assign n13586 = n13564 & n13567 ;
  assign n13587 = n13585 & n13586 ;
  assign n13588 = n13563 & ~n13587 ;
  assign n13589 = n13555 & ~n13561 ;
  assign n13590 = n13542 & n13589 ;
  assign n13591 = ~n13587 & n13590 ;
  assign n13592 = n13535 & ~n13541 ;
  assign n13593 = n13562 & n13592 ;
  assign n13594 = ~n13587 & n13593 ;
  assign n13595 = n13589 & n13592 ;
  assign n13596 = ~n13587 & n13595 ;
  assign n13597 = n13535 & n13548 ;
  assign n13598 = ~n13554 & n13597 ;
  assign n13599 = n13561 & n13598 ;
  assign n13600 = n13541 & n13599 ;
  assign n13601 = ~n13587 & n13600 ;
  assign n13602 = ~n13561 & n13598 ;
  assign n13603 = n13541 & n13602 ;
  assign n13604 = ~n13587 & n13603 ;
  assign n13605 = ~n13541 & n13599 ;
  assign n13606 = ~n13587 & n13605 ;
  assign n13607 = ~n13541 & n13602 ;
  assign n13608 = ~n13587 & n13607 ;
  assign n13611 = \sport0_cfg_FSi_reg/NET0131  & ~\sport0_regs_SCTLreg_DO_reg[6]/NET0131  ;
  assign n13609 = ~\sport0_cfg_FSi_reg/NET0131  & \sport0_regs_SCTLreg_DO_reg[6]/NET0131  ;
  assign n13610 = \sport0_regs_MWORDreg_DO_reg[8]/NET0131  & \sport0_regs_MWORDreg_DO_reg[9]/NET0131  ;
  assign n13612 = ~n13609 & ~n13610 ;
  assign n13613 = ~n13611 & n13612 ;
  assign n13616 = \sport1_cfg_FSi_reg/NET0131  & ~\sport1_regs_SCTLreg_DO_reg[6]/NET0131  ;
  assign n13614 = ~\sport1_cfg_FSi_reg/NET0131  & \sport1_regs_SCTLreg_DO_reg[6]/NET0131  ;
  assign n13615 = \sport1_regs_MWORDreg_DO_reg[8]/NET0131  & \sport1_regs_MWORDreg_DO_reg[9]/NET0131  ;
  assign n13617 = ~n13614 & ~n13615 ;
  assign n13618 = ~n13616 & n13617 ;
  assign n13619 = \sport0_cfg_SCLKi_h_reg/NET0131  & ~\sport0_regs_SCTLreg_DO_reg[13]/NET0131  ;
  assign n13620 = ~\sport0_cfg_SCLKi_h_reg/NET0131  & \sport0_regs_SCTLreg_DO_reg[13]/NET0131  ;
  assign n13621 = ~n13619 & ~n13620 ;
  assign n13622 = \sport1_cfg_SCLKi_h_reg/NET0131  & ~\sport1_regs_SCTLreg_DO_reg[13]/NET0131  ;
  assign n13623 = ~\sport1_cfg_SCLKi_h_reg/NET0131  & \sport1_regs_SCTLreg_DO_reg[13]/NET0131  ;
  assign n13624 = ~n13622 & ~n13623 ;
  assign n13627 = \sport0_regs_SCTLreg_DO_reg[1]/NET0131  & ~\sport0_regs_SCTLreg_DO_reg[2]/NET0131  ;
  assign n13628 = \sport0_txctl_TXSHT_reg[2]/P0001  & n13627 ;
  assign n13625 = ~\sport0_regs_SCTLreg_DO_reg[1]/NET0131  & ~\sport0_regs_SCTLreg_DO_reg[2]/NET0131  ;
  assign n13626 = \sport0_txctl_TXSHT_reg[0]/P0001  & n13625 ;
  assign n13629 = ~\sport0_regs_SCTLreg_DO_reg[0]/NET0131  & ~n13626 ;
  assign n13630 = ~n13628 & n13629 ;
  assign n13632 = \sport0_txctl_TXSHT_reg[3]/P0001  & n13627 ;
  assign n13631 = \sport0_txctl_TXSHT_reg[1]/P0001  & n13625 ;
  assign n13633 = \sport0_regs_SCTLreg_DO_reg[0]/NET0131  & ~n13631 ;
  assign n13634 = ~n13632 & n13633 ;
  assign n13635 = ~n13630 & ~n13634 ;
  assign n13643 = \sport0_regs_SCTLreg_DO_reg[0]/NET0131  & ~\sport0_txctl_TXSHT_reg[5]/P0001  ;
  assign n13641 = ~\sport0_regs_SCTLreg_DO_reg[1]/NET0131  & \sport0_regs_SCTLreg_DO_reg[2]/NET0131  ;
  assign n13642 = ~\sport0_regs_SCTLreg_DO_reg[0]/NET0131  & ~\sport0_txctl_TXSHT_reg[4]/P0001  ;
  assign n13644 = n13641 & ~n13642 ;
  assign n13645 = ~n13643 & n13644 ;
  assign n13638 = \sport0_regs_SCTLreg_DO_reg[0]/NET0131  & ~\sport0_txctl_TXSHT_reg[7]/P0001  ;
  assign n13636 = \sport0_regs_SCTLreg_DO_reg[1]/NET0131  & \sport0_regs_SCTLreg_DO_reg[2]/NET0131  ;
  assign n13637 = ~\sport0_regs_SCTLreg_DO_reg[0]/NET0131  & ~\sport0_txctl_TXSHT_reg[6]/P0001  ;
  assign n13639 = n13636 & ~n13637 ;
  assign n13640 = ~n13638 & n13639 ;
  assign n13646 = ~\sport0_regs_SCTLreg_DO_reg[3]/NET0131  & ~n13640 ;
  assign n13647 = ~n13645 & n13646 ;
  assign n13648 = ~n13635 & n13647 ;
  assign n13649 = \sport0_txctl_TXSHT_reg[13]/P0001  & n13641 ;
  assign n13652 = \sport0_regs_SCTLreg_DO_reg[0]/NET0131  & ~n13649 ;
  assign n13650 = \sport0_txctl_TXSHT_reg[11]/P0001  & n13627 ;
  assign n13651 = \sport0_txctl_TXSHT_reg[9]/P0001  & n13625 ;
  assign n13653 = ~n13650 & ~n13651 ;
  assign n13654 = n13652 & n13653 ;
  assign n13655 = \sport0_txctl_TXSHT_reg[8]/P0001  & n13625 ;
  assign n13658 = ~\sport0_regs_SCTLreg_DO_reg[0]/NET0131  & ~n13655 ;
  assign n13656 = \sport0_txctl_TXSHT_reg[12]/P0001  & n13641 ;
  assign n13657 = \sport0_txctl_TXSHT_reg[10]/P0001  & n13627 ;
  assign n13659 = ~n13656 & ~n13657 ;
  assign n13660 = n13658 & n13659 ;
  assign n13661 = ~n13654 & ~n13660 ;
  assign n13663 = \sport0_regs_SCTLreg_DO_reg[0]/NET0131  & ~\sport0_txctl_TXSHT_reg[15]/P0001  ;
  assign n13662 = ~\sport0_regs_SCTLreg_DO_reg[0]/NET0131  & ~\sport0_txctl_TXSHT_reg[14]/P0001  ;
  assign n13664 = n13636 & ~n13662 ;
  assign n13665 = ~n13663 & n13664 ;
  assign n13666 = \sport0_regs_SCTLreg_DO_reg[3]/NET0131  & ~n13665 ;
  assign n13667 = ~n13661 & n13666 ;
  assign n13668 = ~n13648 & ~n13667 ;
  assign n13669 = ~\sport0_regs_MWORDreg_DO_reg[10]/NET0131  & ~n13668 ;
  assign n13670 = \sport0_regs_MWORDreg_DO_reg[10]/NET0131  & ~\sport0_txctl_TXSHT_reg[15]/P0001  ;
  assign n13671 = ~n13669 & ~n13670 ;
  assign n13672 = ~\sport0_regs_SCTLreg_DO_reg[15]/NET0131  & n13671 ;
  assign n13673 = \sport1_regs_MWORDreg_DO_reg[10]/NET0131  & ~\sport1_txctl_TXSHT_reg[15]/P0001  ;
  assign n13676 = ~\sport1_regs_SCTLreg_DO_reg[0]/NET0131  & ~\sport1_txctl_TXSHT_reg[2]/P0001  ;
  assign n13674 = \sport1_regs_SCTLreg_DO_reg[1]/NET0131  & ~\sport1_regs_SCTLreg_DO_reg[2]/NET0131  ;
  assign n13675 = \sport1_regs_SCTLreg_DO_reg[0]/NET0131  & ~\sport1_txctl_TXSHT_reg[3]/P0001  ;
  assign n13677 = n13674 & ~n13675 ;
  assign n13678 = ~n13676 & n13677 ;
  assign n13694 = ~\sport1_regs_SCTLreg_DO_reg[3]/NET0131  & ~n13678 ;
  assign n13691 = \sport1_regs_SCTLreg_DO_reg[0]/NET0131  & ~\sport1_txctl_TXSHT_reg[1]/P0001  ;
  assign n13689 = ~\sport1_regs_SCTLreg_DO_reg[1]/NET0131  & ~\sport1_regs_SCTLreg_DO_reg[2]/NET0131  ;
  assign n13690 = ~\sport1_regs_SCTLreg_DO_reg[0]/NET0131  & ~\sport1_txctl_TXSHT_reg[0]/P0001  ;
  assign n13692 = n13689 & ~n13690 ;
  assign n13693 = ~n13691 & n13692 ;
  assign n13681 = \sport1_regs_SCTLreg_DO_reg[0]/NET0131  & ~\sport1_txctl_TXSHT_reg[7]/P0001  ;
  assign n13679 = \sport1_regs_SCTLreg_DO_reg[1]/NET0131  & \sport1_regs_SCTLreg_DO_reg[2]/NET0131  ;
  assign n13680 = ~\sport1_regs_SCTLreg_DO_reg[0]/NET0131  & ~\sport1_txctl_TXSHT_reg[6]/P0001  ;
  assign n13682 = n13679 & ~n13680 ;
  assign n13683 = ~n13681 & n13682 ;
  assign n13686 = \sport1_regs_SCTLreg_DO_reg[0]/NET0131  & ~\sport1_txctl_TXSHT_reg[5]/P0001  ;
  assign n13684 = ~\sport1_regs_SCTLreg_DO_reg[1]/NET0131  & \sport1_regs_SCTLreg_DO_reg[2]/NET0131  ;
  assign n13685 = ~\sport1_regs_SCTLreg_DO_reg[0]/NET0131  & ~\sport1_txctl_TXSHT_reg[4]/P0001  ;
  assign n13687 = n13684 & ~n13685 ;
  assign n13688 = ~n13686 & n13687 ;
  assign n13695 = ~n13683 & ~n13688 ;
  assign n13696 = ~n13693 & n13695 ;
  assign n13697 = n13694 & n13696 ;
  assign n13699 = \sport1_regs_SCTLreg_DO_reg[0]/NET0131  & ~\sport1_txctl_TXSHT_reg[15]/P0001  ;
  assign n13698 = ~\sport1_regs_SCTLreg_DO_reg[0]/NET0131  & ~\sport1_txctl_TXSHT_reg[14]/P0001  ;
  assign n13700 = n13679 & ~n13698 ;
  assign n13701 = ~n13699 & n13700 ;
  assign n13714 = \sport1_regs_SCTLreg_DO_reg[3]/NET0131  & ~n13701 ;
  assign n13711 = \sport1_regs_SCTLreg_DO_reg[0]/NET0131  & ~\sport1_txctl_TXSHT_reg[13]/P0001  ;
  assign n13710 = ~\sport1_regs_SCTLreg_DO_reg[0]/NET0131  & ~\sport1_txctl_TXSHT_reg[12]/P0001  ;
  assign n13712 = n13684 & ~n13710 ;
  assign n13713 = ~n13711 & n13712 ;
  assign n13703 = \sport1_regs_SCTLreg_DO_reg[0]/NET0131  & ~\sport1_txctl_TXSHT_reg[9]/P0001  ;
  assign n13702 = ~\sport1_regs_SCTLreg_DO_reg[0]/NET0131  & ~\sport1_txctl_TXSHT_reg[8]/P0001  ;
  assign n13704 = n13689 & ~n13702 ;
  assign n13705 = ~n13703 & n13704 ;
  assign n13707 = \sport1_regs_SCTLreg_DO_reg[0]/NET0131  & ~\sport1_txctl_TXSHT_reg[11]/P0001  ;
  assign n13706 = ~\sport1_regs_SCTLreg_DO_reg[0]/NET0131  & ~\sport1_txctl_TXSHT_reg[10]/P0001  ;
  assign n13708 = n13674 & ~n13706 ;
  assign n13709 = ~n13707 & n13708 ;
  assign n13715 = ~n13705 & ~n13709 ;
  assign n13716 = ~n13713 & n13715 ;
  assign n13717 = n13714 & n13716 ;
  assign n13718 = ~n13697 & ~n13717 ;
  assign n13719 = ~\sport1_regs_MWORDreg_DO_reg[10]/NET0131  & ~n13718 ;
  assign n13720 = ~n13673 & ~n13719 ;
  assign n13721 = ~\sport1_regs_SCTLreg_DO_reg[15]/NET0131  & n13720 ;
  assign n13723 = ~\sport0_cfg_FSi_reg/NET0131  & \sport0_regs_SCTLreg_DO_reg[7]/NET0131  ;
  assign n13722 = \sport0_cfg_FSi_reg/NET0131  & ~\sport0_regs_SCTLreg_DO_reg[7]/NET0131  ;
  assign n13724 = ~n13610 & ~n13722 ;
  assign n13725 = ~n13723 & n13724 ;
  assign n13727 = ~\sport1_cfg_FSi_reg/NET0131  & \sport1_regs_SCTLreg_DO_reg[7]/NET0131  ;
  assign n13726 = \sport1_cfg_FSi_reg/NET0131  & ~\sport1_regs_SCTLreg_DO_reg[7]/NET0131  ;
  assign n13728 = ~n13615 & ~n13726 ;
  assign n13729 = ~n13727 & n13728 ;
  assign n13730 = ~\bdma_BM_cyc_reg/P0001  & \emc_WRn_h_reg/P0001  ;
  assign n13731 = \bdma_BM_cyc_reg/P0001  & \bdma_BWRn_reg/NET0131  ;
  assign n13732 = ~n13730 & ~n13731 ;
  assign n13733 = ~T_BMODE_pad & ~T_MMAP_pad ;
  assign n13734 = \bdma_RST_pin_reg/P0001  & n13733 ;
  assign n13747 = ~n5733 & ~n13147 ;
  assign n13748 = ~n5561 & ~n5563 ;
  assign n13749 = n5560 & n5597 ;
  assign n13750 = n5587 & n13749 ;
  assign n13751 = ~n13748 & n13750 ;
  assign n13752 = ~n13747 & n13751 ;
  assign n13753 = n6915 & n13751 ;
  assign n13754 = ~n6914 & n13753 ;
  assign n13755 = ~n13752 & ~n13754 ;
  assign n13735 = ~\bdma_BWCOUNT_reg[3]/NET0131  & ~\bdma_BWCOUNT_reg[4]/NET0131  ;
  assign n13736 = ~\bdma_BWCOUNT_reg[1]/NET0131  & ~\bdma_BWCOUNT_reg[2]/NET0131  ;
  assign n13737 = ~\bdma_BWCOUNT_reg[6]/NET0131  & n13736 ;
  assign n13738 = n13735 & n13737 ;
  assign n13739 = n10716 & n13738 ;
  assign n13742 = ~\bdma_BWCOUNT_reg[7]/NET0131  & ~\bdma_BWCOUNT_reg[8]/NET0131  ;
  assign n13743 = ~\bdma_BWCOUNT_reg[9]/NET0131  & n13742 ;
  assign n13740 = ~\bdma_BWCOUNT_reg[10]/NET0131  & ~\bdma_BWCOUNT_reg[11]/NET0131  ;
  assign n13741 = ~\bdma_BWCOUNT_reg[12]/NET0131  & ~\bdma_BWCOUNT_reg[13]/NET0131  ;
  assign n13744 = n13740 & n13741 ;
  assign n13745 = n13743 & n13744 ;
  assign n13746 = n13739 & n13745 ;
  assign n13756 = \bdma_BWCOUNT_reg[0]/NET0131  & n13746 ;
  assign n13757 = ~n13755 & n13756 ;
  assign n13758 = ~n4063 & ~n13757 ;
  assign n13759 = ~n13734 & ~n13758 ;
  assign n13764 = ~\bdma_BWCOUNT_reg[0]/NET0131  & ~n13755 ;
  assign n13765 = ~\bdma_BWCOUNT_reg[1]/NET0131  & n13764 ;
  assign n13766 = ~\bdma_BWCOUNT_reg[2]/NET0131  & n13765 ;
  assign n13767 = n13735 & n13766 ;
  assign n13769 = n10716 & n13767 ;
  assign n13760 = \memc_Dwrite_E_reg/NET0131  & ~n5950 ;
  assign n13761 = ~\core_c_dec_Dummy_E_reg/NET0131  & n13760 ;
  assign n13762 = n7285 & n13761 ;
  assign n13763 = n7284 & n13762 ;
  assign n13768 = ~n10716 & ~n13767 ;
  assign n13770 = ~n13763 & ~n13768 ;
  assign n13771 = ~n13769 & n13770 ;
  assign n13772 = ~n10911 & n13763 ;
  assign n13773 = ~n13771 & ~n13772 ;
  assign n13774 = ~n13734 & ~n13773 ;
  assign n13775 = \core_c_psq_cntstk_ptr_reg[0]/NET0131  & \core_c_psq_cntstk_ptr_reg[1]/NET0131  ;
  assign n13776 = ~\core_c_psq_cntstk_ptr_reg[2]/NET0131  & n13775 ;
  assign n13777 = \core_c_dec_MTCNTR_Eg_reg/P0001  & \core_c_psq_CNTRval_reg/NET0131  ;
  assign n13778 = ~n5950 & n13777 ;
  assign n13779 = ~n13776 & n13778 ;
  assign n13780 = n13775 & n13779 ;
  assign n13781 = \core_c_psq_cntstk_cnts4x14_CNTcell_reg[0][5]/P0001  & ~n13780 ;
  assign n13782 = \core_c_psq_CNTR_reg_DO_reg[5]/NET0131  & n13780 ;
  assign n13783 = ~n13781 & ~n13782 ;
  assign n13784 = ~\core_c_psq_cntstk_ptr_reg[0]/NET0131  & ~\core_c_psq_cntstk_ptr_reg[1]/NET0131  ;
  assign n13785 = n13778 & n13784 ;
  assign n13786 = \core_c_psq_cntstk_cnts4x14_CNTcell_reg[1][5]/P0001  & ~n13785 ;
  assign n13787 = \core_c_psq_CNTR_reg_DO_reg[5]/NET0131  & n13785 ;
  assign n13788 = ~n13786 & ~n13787 ;
  assign n13789 = \core_c_psq_cntstk_ptr_reg[0]/NET0131  & ~\core_c_psq_cntstk_ptr_reg[1]/NET0131  ;
  assign n13790 = n13778 & n13789 ;
  assign n13791 = \core_c_psq_cntstk_cnts4x14_CNTcell_reg[2][5]/P0001  & ~n13790 ;
  assign n13792 = \core_c_psq_CNTR_reg_DO_reg[5]/NET0131  & n13790 ;
  assign n13793 = ~n13791 & ~n13792 ;
  assign n13794 = ~\core_c_psq_cntstk_ptr_reg[0]/NET0131  & \core_c_psq_cntstk_ptr_reg[1]/NET0131  ;
  assign n13795 = n13778 & n13794 ;
  assign n13796 = \core_c_psq_cntstk_cnts4x14_CNTcell_reg[3][5]/P0001  & ~n13795 ;
  assign n13797 = \core_c_psq_CNTR_reg_DO_reg[5]/NET0131  & n13795 ;
  assign n13798 = ~n13796 & ~n13797 ;
  assign n13799 = ~\core_c_dec_DIVQ_E_reg/P0001  & ~\core_c_dec_DIVS_E_reg/P0001  ;
  assign n13800 = ~\core_c_dec_updAF_E_reg/P0001  & n13799 ;
  assign n13801 = ~\core_c_psq_MSTAT_reg_DO_reg[0]/P0002  & ~n5950 ;
  assign n13802 = \core_c_dec_Usecond_E_reg/P0001  & n4184 ;
  assign n13803 = ~\core_c_dec_Dummy_E_reg/NET0131  & ~n13802 ;
  assign n13804 = n13801 & n13803 ;
  assign n13805 = ~n13800 & n13804 ;
  assign n13806 = ~\core_c_dec_Dummy_E_reg/NET0131  & ~n13799 ;
  assign n13807 = \core_eu_ea_alu_ea_dec_AMF_E_reg[0]/NET0131  & \core_eu_ea_alu_ea_dec_AMF_E_reg[1]/NET0131  ;
  assign n13808 = \core_eu_ea_alu_ea_dec_AMF_E_reg[2]/NET0131  & \core_eu_ea_alu_ea_dec_AMF_E_reg[3]/NET0131  ;
  assign n13809 = ~n13807 & n13808 ;
  assign n13810 = \core_eu_ea_alu_ea_dec_AMF_E_reg[3]/NET0131  & n13807 ;
  assign n13811 = \core_eu_ea_alu_ea_dec_AMF_E_reg[2]/NET0131  & n13810 ;
  assign n13825 = \core_c_dec_IRE_reg[8]/NET0131  & n12000 ;
  assign n13823 = \core_c_dec_IRE_reg[10]/NET0131  & \core_c_dec_IRE_reg[9]/NET0131  ;
  assign n13824 = ~\core_c_dec_IRE_reg[8]/NET0131  & n11992 ;
  assign n13826 = n13823 & ~n13824 ;
  assign n13827 = ~n13825 & n13826 ;
  assign n13812 = \core_c_dec_IRE_reg[10]/NET0131  & ~\core_c_dec_IRE_reg[9]/NET0131  ;
  assign n13813 = \core_c_dec_IRE_reg[8]/NET0131  & n13812 ;
  assign n13814 = ~n7206 & n13813 ;
  assign n13815 = ~\core_c_dec_IRE_reg[10]/NET0131  & ~\core_c_dec_IRE_reg[8]/NET0131  ;
  assign n13816 = \core_c_dec_IRE_reg[9]/NET0131  & n13815 ;
  assign n13817 = ~n11983 & n13816 ;
  assign n13828 = ~n13814 & ~n13817 ;
  assign n13818 = \core_c_dec_IRE_reg[8]/NET0131  & \core_c_dec_IRE_reg[9]/NET0131  ;
  assign n13819 = ~\core_c_dec_IRE_reg[10]/NET0131  & n13818 ;
  assign n13820 = ~n12024 & n13819 ;
  assign n13821 = ~\core_c_dec_IRE_reg[8]/NET0131  & n13812 ;
  assign n13822 = ~n12028 & n13821 ;
  assign n13829 = ~n13820 & ~n13822 ;
  assign n13830 = n13828 & n13829 ;
  assign n13831 = ~n13827 & n13830 ;
  assign n13834 = \core_c_dec_IRE_reg[8]/NET0131  & n11971 ;
  assign n13832 = ~\core_c_dec_IRE_reg[10]/NET0131  & ~\core_c_dec_IRE_reg[9]/NET0131  ;
  assign n13833 = ~\core_c_dec_IRE_reg[8]/NET0131  & n11967 ;
  assign n13835 = n13832 & ~n13833 ;
  assign n13836 = ~n13834 & n13835 ;
  assign n13837 = n13831 & ~n13836 ;
  assign n13838 = n13811 & ~n13837 ;
  assign n13839 = ~\core_c_dec_ALUop_E_reg/P0001  & ~\core_c_dec_DIVQ_E_reg/P0001  ;
  assign n13840 = ~\core_c_dec_DIVS_E_reg/P0001  & n13839 ;
  assign n13841 = \core_c_dec_DIVQ_E_reg/P0001  & ~\core_eu_ec_cun_AQ_reg/P0001  ;
  assign n13842 = ~n13840 & ~n13841 ;
  assign n13843 = ~\core_eu_ea_alu_ea_dec_AMF_E_reg[0]/NET0131  & ~\core_eu_ea_alu_ea_dec_AMF_E_reg[1]/NET0131  ;
  assign n13844 = \core_c_dec_DIVQ_E_reg/P0001  & n13843 ;
  assign n13845 = ~\core_eu_ea_alu_ea_dec_AMF_E_reg[2]/NET0131  & \core_eu_ea_alu_ea_dec_AMF_E_reg[3]/NET0131  ;
  assign n13846 = ~n13844 & n13845 ;
  assign n13847 = n13842 & ~n13846 ;
  assign n13848 = ~n13838 & n13847 ;
  assign n14057 = \core_c_dec_IRE_reg[8]/NET0131  & n7991 ;
  assign n14056 = ~\core_c_dec_IRE_reg[8]/NET0131  & n7987 ;
  assign n14058 = n13823 & ~n14056 ;
  assign n14059 = ~n14057 & n14058 ;
  assign n14055 = ~n7905 & n13813 ;
  assign n14060 = ~n7909 & n13819 ;
  assign n14063 = ~n14055 & ~n14060 ;
  assign n14061 = ~n7885 & n13821 ;
  assign n14062 = ~n7952 & n13816 ;
  assign n14064 = ~n14061 & ~n14062 ;
  assign n14065 = n14063 & n14064 ;
  assign n14066 = ~n14059 & n14065 ;
  assign n14067 = ~n13832 & n14066 ;
  assign n13849 = ~\core_c_dec_DIVQ_E_reg/P0001  & ~\core_eu_ea_alu_ea_dec_AMF_E_reg[0]/NET0131  ;
  assign n13850 = ~\core_eu_ea_alu_ea_dec_AMF_E_reg[2]/NET0131  & n13849 ;
  assign n13851 = \core_eu_ea_alu_ea_dec_AMF_E_reg[3]/NET0131  & ~n13850 ;
  assign n13852 = ~\core_eu_ea_alu_ea_dec_AMF_E_reg[1]/NET0131  & ~n13851 ;
  assign n13853 = ~n13840 & ~n13852 ;
  assign n14052 = \core_c_dec_IRE_reg[8]/NET0131  & ~n7956 ;
  assign n14051 = ~\core_c_dec_IRE_reg[8]/NET0131  & ~n7960 ;
  assign n14053 = n13832 & ~n14051 ;
  assign n14054 = ~n14052 & n14053 ;
  assign n14068 = n13853 & ~n14054 ;
  assign n14069 = ~n14067 & n14068 ;
  assign n14070 = n13848 & n14069 ;
  assign n14071 = ~n13848 & ~n14069 ;
  assign n14072 = ~n14070 & ~n14071 ;
  assign n13874 = \core_eu_ea_alu_ea_dec_AMF_E_reg[2]/NET0131  & ~\core_eu_ea_alu_ea_dec_AMF_E_reg[3]/NET0131  ;
  assign n13875 = ~\core_c_dec_IRE_reg[4]/NET0131  & ~\core_c_dec_IRE_reg[5]/NET0131  ;
  assign n13876 = ~\core_c_dec_IRE_reg[6]/NET0131  & ~\core_c_dec_IRE_reg[7]/NET0131  ;
  assign n13877 = n13875 & n13876 ;
  assign n13878 = \core_c_dec_cdAM_E_reg/P0001  & ~n13877 ;
  assign n14074 = \core_c_psq_MSTAT_reg_DO_reg[0]/P0002  & ~\core_eu_ea_alu_ea_reg_afswe_DO_reg[3]/P0001  ;
  assign n14033 = ~\core_c_dec_IRE_reg[11]/NET0131  & \core_c_dec_IRE_reg[12]/NET0131  ;
  assign n14073 = ~\core_c_psq_MSTAT_reg_DO_reg[0]/P0002  & ~\core_eu_ea_alu_ea_reg_afrwe_DO_reg[3]/P0001  ;
  assign n14075 = n14033 & ~n14073 ;
  assign n14076 = ~n14074 & n14075 ;
  assign n14078 = \core_c_dec_IRE_reg[11]/NET0131  & n7948 ;
  assign n14077 = ~\core_c_dec_IRE_reg[11]/NET0131  & n7944 ;
  assign n14079 = ~\core_c_dec_IRE_reg[12]/NET0131  & ~n14077 ;
  assign n14080 = ~n14078 & n14079 ;
  assign n14081 = ~n14076 & ~n14080 ;
  assign n14082 = ~n13878 & ~n14081 ;
  assign n14083 = \core_eu_ea_alu_ea_dec_piconst_DO_reg[3]/P0001  & n13878 ;
  assign n14084 = ~n14082 & ~n14083 ;
  assign n14086 = n13874 & n14084 ;
  assign n13880 = ~n13810 & ~n13840 ;
  assign n14032 = ~n13874 & n13880 ;
  assign n14085 = n14032 & ~n14084 ;
  assign n14087 = ~n13840 & ~n14085 ;
  assign n14088 = ~n14086 & n14087 ;
  assign n14089 = n14072 & n14088 ;
  assign n14131 = \core_c_dec_IRE_reg[8]/NET0131  & n8497 ;
  assign n14130 = ~\core_c_dec_IRE_reg[8]/NET0131  & n8493 ;
  assign n14132 = n13823 & ~n14130 ;
  assign n14133 = ~n14131 & n14132 ;
  assign n14129 = ~n8534 & n13813 ;
  assign n14134 = ~n8585 & n13816 ;
  assign n14137 = ~n14129 & ~n14134 ;
  assign n14135 = ~n8554 & n13819 ;
  assign n14136 = ~n8558 & n13821 ;
  assign n14138 = ~n14135 & ~n14136 ;
  assign n14139 = n14137 & n14138 ;
  assign n14140 = ~n14133 & n14139 ;
  assign n14142 = \core_c_dec_IRE_reg[8]/NET0131  & n8589 ;
  assign n14141 = ~\core_c_dec_IRE_reg[8]/NET0131  & n8593 ;
  assign n14143 = n13832 & ~n14141 ;
  assign n14144 = ~n14142 & n14143 ;
  assign n14145 = n14140 & ~n14144 ;
  assign n14146 = n13853 & ~n14145 ;
  assign n14147 = n13848 & ~n14146 ;
  assign n14148 = ~n13848 & n14146 ;
  assign n14149 = ~n14147 & ~n14148 ;
  assign n13895 = ~n13840 & ~n13874 ;
  assign n14153 = ~\core_c_psq_MSTAT_reg_DO_reg[0]/P0002  & ~\core_eu_ea_alu_ea_reg_afrwe_DO_reg[2]/P0001  ;
  assign n14154 = \core_c_psq_MSTAT_reg_DO_reg[0]/P0002  & ~\core_eu_ea_alu_ea_reg_afswe_DO_reg[2]/P0001  ;
  assign n14155 = ~n14153 & ~n14154 ;
  assign n14156 = \core_c_dec_IRE_reg[12]/NET0131  & ~n14155 ;
  assign n14152 = ~\core_c_dec_IRE_reg[12]/NET0131  & n8577 ;
  assign n14157 = ~\core_c_dec_IRE_reg[11]/NET0131  & ~n14152 ;
  assign n14158 = ~n14156 & n14157 ;
  assign n13881 = \core_c_dec_IRE_reg[11]/NET0131  & ~\core_c_dec_IRE_reg[12]/NET0131  ;
  assign n14151 = ~n8581 & n13881 ;
  assign n14159 = ~n13878 & ~n14151 ;
  assign n14160 = ~n14158 & n14159 ;
  assign n14150 = ~\core_eu_ea_alu_ea_dec_piconst_DO_reg[2]/P0001  & n13878 ;
  assign n14161 = n13880 & ~n14150 ;
  assign n14162 = ~n14160 & n14161 ;
  assign n14163 = n13895 & ~n14162 ;
  assign n14164 = n13874 & n14162 ;
  assign n14165 = ~n14163 & ~n14164 ;
  assign n14166 = ~n14149 & ~n14165 ;
  assign n14169 = \core_c_dec_IRE_reg[8]/NET0131  & n9280 ;
  assign n14168 = ~\core_c_dec_IRE_reg[8]/NET0131  & n9276 ;
  assign n14170 = n13823 & ~n14168 ;
  assign n14171 = ~n14169 & n14170 ;
  assign n14167 = ~n9229 & n13813 ;
  assign n14172 = ~n9297 & n13816 ;
  assign n14175 = ~n14167 & ~n14172 ;
  assign n14173 = ~n9225 & n13819 ;
  assign n14174 = ~n9205 & n13821 ;
  assign n14176 = ~n14173 & ~n14174 ;
  assign n14177 = n14175 & n14176 ;
  assign n14178 = ~n14171 & n14177 ;
  assign n14180 = \core_c_dec_IRE_reg[8]/NET0131  & n9313 ;
  assign n14179 = ~\core_c_dec_IRE_reg[8]/NET0131  & n9309 ;
  assign n14181 = n13832 & ~n14179 ;
  assign n14182 = ~n14180 & n14181 ;
  assign n14183 = n14178 & ~n14182 ;
  assign n14184 = n13853 & ~n14183 ;
  assign n14185 = n13848 & ~n14184 ;
  assign n14186 = ~n13848 & n14184 ;
  assign n14187 = ~n14185 & ~n14186 ;
  assign n14191 = ~\core_c_psq_MSTAT_reg_DO_reg[0]/P0002  & ~\core_eu_ea_alu_ea_reg_afrwe_DO_reg[1]/P0001  ;
  assign n14192 = \core_c_psq_MSTAT_reg_DO_reg[0]/P0002  & ~\core_eu_ea_alu_ea_reg_afswe_DO_reg[1]/P0001  ;
  assign n14193 = ~n14191 & ~n14192 ;
  assign n14194 = \core_c_dec_IRE_reg[12]/NET0131  & ~n14193 ;
  assign n14190 = ~\core_c_dec_IRE_reg[12]/NET0131  & n9305 ;
  assign n14195 = ~\core_c_dec_IRE_reg[11]/NET0131  & ~n14190 ;
  assign n14196 = ~n14194 & n14195 ;
  assign n14189 = ~n9301 & n13881 ;
  assign n14197 = ~n13878 & ~n14189 ;
  assign n14198 = ~n14196 & n14197 ;
  assign n14188 = ~\core_eu_ea_alu_ea_dec_piconst_DO_reg[1]/P0001  & n13878 ;
  assign n14199 = n13880 & ~n14188 ;
  assign n14200 = ~n14198 & n14199 ;
  assign n14201 = n13895 & ~n14200 ;
  assign n14202 = n13874 & n14200 ;
  assign n14203 = ~n14201 & ~n14202 ;
  assign n14204 = n14187 & n14203 ;
  assign n14207 = \core_c_dec_IRE_reg[8]/NET0131  & n7377 ;
  assign n14206 = ~\core_c_dec_IRE_reg[8]/NET0131  & n7381 ;
  assign n14208 = n13823 & ~n14206 ;
  assign n14209 = ~n14207 & n14208 ;
  assign n14205 = ~n7449 & n13821 ;
  assign n14210 = ~n7469 & n13819 ;
  assign n14213 = ~n14205 & ~n14210 ;
  assign n14211 = ~n7473 & n13813 ;
  assign n14212 = ~n7422 & n13816 ;
  assign n14214 = ~n14211 & ~n14212 ;
  assign n14215 = n14213 & n14214 ;
  assign n14216 = ~n14209 & n14215 ;
  assign n14217 = ~n13832 & ~n14216 ;
  assign n14219 = \core_c_dec_IRE_reg[8]/NET0131  & n7426 ;
  assign n14218 = ~\core_c_dec_IRE_reg[8]/NET0131  & n7430 ;
  assign n14220 = n13832 & ~n14218 ;
  assign n14221 = ~n14219 & n14220 ;
  assign n14222 = ~n14217 & ~n14221 ;
  assign n14223 = n13853 & ~n14222 ;
  assign n14224 = n13848 & ~n14223 ;
  assign n14225 = ~n13848 & n14223 ;
  assign n14226 = ~n14224 & ~n14225 ;
  assign n14230 = ~\core_c_psq_MSTAT_reg_DO_reg[0]/P0002  & ~\core_eu_ea_alu_ea_reg_afrwe_DO_reg[0]/P0001  ;
  assign n14231 = \core_c_psq_MSTAT_reg_DO_reg[0]/P0002  & ~\core_eu_ea_alu_ea_reg_afswe_DO_reg[0]/P0001  ;
  assign n14232 = ~n14230 & ~n14231 ;
  assign n14233 = \core_c_dec_IRE_reg[12]/NET0131  & ~n14232 ;
  assign n14229 = ~\core_c_dec_IRE_reg[12]/NET0131  & n7414 ;
  assign n14234 = ~\core_c_dec_IRE_reg[11]/NET0131  & ~n14229 ;
  assign n14235 = ~n14233 & n14234 ;
  assign n14228 = ~n7418 & n13881 ;
  assign n14236 = ~n13878 & ~n14228 ;
  assign n14237 = ~n14235 & n14236 ;
  assign n14227 = ~\core_eu_ea_alu_ea_dec_piconst_DO_reg[0]/P0001  & n13878 ;
  assign n14238 = n13880 & ~n14227 ;
  assign n14239 = ~n14237 & n14238 ;
  assign n14240 = n13895 & ~n14239 ;
  assign n14241 = n13874 & n14239 ;
  assign n14242 = ~n14240 & ~n14241 ;
  assign n14243 = ~n14226 & ~n14242 ;
  assign n14244 = ~n14187 & ~n14203 ;
  assign n14245 = \core_eu_ea_alu_ea_dec_AMF_E_reg[1]/NET0131  & \core_eu_ec_cun_AC_reg/P0001  ;
  assign n14246 = ~\core_eu_ea_alu_ea_dec_AMF_E_reg[0]/NET0131  & ~n14245 ;
  assign n14247 = ~n13807 & ~n13808 ;
  assign n14248 = ~n14246 & n14247 ;
  assign n14249 = n13807 & n13874 ;
  assign n14250 = n13842 & ~n14249 ;
  assign n14251 = ~n14248 & n14250 ;
  assign n14252 = ~n13838 & n14251 ;
  assign n14253 = ~n14244 & ~n14252 ;
  assign n14254 = n14226 & n14242 ;
  assign n14255 = ~n14253 & ~n14254 ;
  assign n14256 = ~n14243 & ~n14255 ;
  assign n14257 = ~n14204 & ~n14256 ;
  assign n14258 = ~n14166 & ~n14257 ;
  assign n14259 = ~n14089 & n14258 ;
  assign n14260 = ~n14072 & ~n14088 ;
  assign n14013 = \core_c_dec_IRE_reg[8]/NET0131  & n10797 ;
  assign n14012 = ~\core_c_dec_IRE_reg[8]/NET0131  & n10801 ;
  assign n14014 = n13823 & ~n14012 ;
  assign n14015 = ~n14013 & n14014 ;
  assign n14011 = ~n10878 & n13819 ;
  assign n14016 = ~n10858 & n13821 ;
  assign n14019 = ~n14011 & ~n14016 ;
  assign n14017 = ~n10882 & n13813 ;
  assign n14018 = ~n10694 & n13816 ;
  assign n14020 = ~n14017 & ~n14018 ;
  assign n14021 = n14019 & n14020 ;
  assign n14022 = ~n14015 & n14021 ;
  assign n14024 = \core_c_dec_IRE_reg[8]/NET0131  & n10698 ;
  assign n14023 = ~\core_c_dec_IRE_reg[8]/NET0131  & n10702 ;
  assign n14025 = n13832 & ~n14023 ;
  assign n14026 = ~n14024 & n14025 ;
  assign n14027 = n14022 & ~n14026 ;
  assign n14028 = n13853 & ~n14027 ;
  assign n14029 = ~n13848 & n14028 ;
  assign n14030 = n13848 & ~n14028 ;
  assign n14031 = ~n14029 & ~n14030 ;
  assign n14035 = \core_c_psq_MSTAT_reg_DO_reg[0]/P0002  & ~\core_eu_ea_alu_ea_reg_afswe_DO_reg[5]/P0001  ;
  assign n14034 = ~\core_c_psq_MSTAT_reg_DO_reg[0]/P0002  & ~\core_eu_ea_alu_ea_reg_afrwe_DO_reg[5]/P0001  ;
  assign n14036 = n14033 & ~n14034 ;
  assign n14037 = ~n14035 & n14036 ;
  assign n14039 = \core_c_dec_IRE_reg[11]/NET0131  & n10690 ;
  assign n14038 = ~\core_c_dec_IRE_reg[11]/NET0131  & n10686 ;
  assign n14040 = ~\core_c_dec_IRE_reg[12]/NET0131  & ~n14038 ;
  assign n14041 = ~n14039 & n14040 ;
  assign n14042 = ~n14037 & ~n14041 ;
  assign n14043 = ~n13878 & ~n14042 ;
  assign n14044 = \core_eu_ea_alu_ea_dec_piconst_DO_reg[5]/P0001  & n13878 ;
  assign n14045 = ~n14043 & ~n14044 ;
  assign n14047 = n13874 & n14045 ;
  assign n14046 = n14032 & ~n14045 ;
  assign n14048 = ~n13840 & ~n14046 ;
  assign n14049 = ~n14047 & n14048 ;
  assign n14261 = ~n14031 & n14049 ;
  assign n14262 = n14149 & n14165 ;
  assign n14263 = ~n14261 & n14262 ;
  assign n14264 = ~n14260 & ~n14263 ;
  assign n14265 = ~n14259 & n14264 ;
  assign n14092 = \core_c_dec_IRE_reg[8]/NET0131  & n9947 ;
  assign n14091 = ~\core_c_dec_IRE_reg[8]/NET0131  & n9951 ;
  assign n14093 = n13823 & ~n14091 ;
  assign n14094 = ~n14092 & n14093 ;
  assign n14090 = ~n9865 & n13813 ;
  assign n14095 = ~n9869 & n13819 ;
  assign n14098 = ~n14090 & ~n14095 ;
  assign n14096 = ~n9845 & n13821 ;
  assign n14097 = ~n9912 & n13816 ;
  assign n14099 = ~n14096 & ~n14097 ;
  assign n14100 = n14098 & n14099 ;
  assign n14101 = ~n14094 & n14100 ;
  assign n14103 = \core_c_dec_IRE_reg[8]/NET0131  & n9916 ;
  assign n14102 = ~\core_c_dec_IRE_reg[8]/NET0131  & n9920 ;
  assign n14104 = n13832 & ~n14102 ;
  assign n14105 = ~n14103 & n14104 ;
  assign n14106 = n14101 & ~n14105 ;
  assign n14107 = n13853 & ~n14106 ;
  assign n14108 = n13848 & ~n14107 ;
  assign n14109 = ~n13848 & n14107 ;
  assign n14110 = ~n14108 & ~n14109 ;
  assign n14114 = ~\core_c_psq_MSTAT_reg_DO_reg[0]/P0002  & ~\core_eu_ea_alu_ea_reg_afrwe_DO_reg[4]/P0001  ;
  assign n14115 = \core_c_psq_MSTAT_reg_DO_reg[0]/P0002  & ~\core_eu_ea_alu_ea_reg_afswe_DO_reg[4]/P0001  ;
  assign n14116 = ~n14114 & ~n14115 ;
  assign n14117 = \core_c_dec_IRE_reg[12]/NET0131  & ~n14116 ;
  assign n14113 = ~\core_c_dec_IRE_reg[12]/NET0131  & n9904 ;
  assign n14118 = ~\core_c_dec_IRE_reg[11]/NET0131  & ~n14113 ;
  assign n14119 = ~n14117 & n14118 ;
  assign n14112 = ~n9908 & n13881 ;
  assign n14120 = ~n13878 & ~n14112 ;
  assign n14121 = ~n14119 & n14120 ;
  assign n14111 = ~\core_eu_ea_alu_ea_dec_piconst_DO_reg[4]/P0001  & n13878 ;
  assign n14122 = n13880 & ~n14111 ;
  assign n14123 = ~n14121 & n14122 ;
  assign n14124 = n13895 & ~n14123 ;
  assign n14125 = n13874 & n14123 ;
  assign n14126 = ~n14124 & ~n14125 ;
  assign n14266 = ~n14110 & ~n14126 ;
  assign n14267 = ~n14261 & ~n14266 ;
  assign n14268 = ~n14265 & n14267 ;
  assign n14050 = n14031 & ~n14049 ;
  assign n14127 = n14110 & n14126 ;
  assign n14128 = ~n14089 & n14127 ;
  assign n14269 = ~n14050 & ~n14128 ;
  assign n14270 = ~n14268 & n14269 ;
  assign n13940 = \core_c_dec_IRE_reg[8]/NET0131  & n11239 ;
  assign n13939 = ~\core_c_dec_IRE_reg[8]/NET0131  & n11231 ;
  assign n13941 = n13823 & ~n13939 ;
  assign n13942 = ~n13940 & n13941 ;
  assign n13936 = ~n11192 & n13819 ;
  assign n13943 = ~n13814 & ~n13936 ;
  assign n13937 = ~n11196 & n13821 ;
  assign n13938 = ~n11062 & n13816 ;
  assign n13944 = ~n13937 & ~n13938 ;
  assign n13945 = n13943 & n13944 ;
  assign n13946 = ~n13942 & n13945 ;
  assign n13948 = \core_c_dec_IRE_reg[8]/NET0131  & n11066 ;
  assign n13947 = ~\core_c_dec_IRE_reg[8]/NET0131  & n11070 ;
  assign n13949 = n13832 & ~n13947 ;
  assign n13950 = ~n13948 & n13949 ;
  assign n13951 = n13946 & ~n13950 ;
  assign n13952 = n13853 & ~n13951 ;
  assign n13953 = ~n13848 & n13952 ;
  assign n13954 = n13848 & ~n13952 ;
  assign n13955 = ~n13953 & ~n13954 ;
  assign n13959 = ~\core_c_psq_MSTAT_reg_DO_reg[0]/P0002  & ~\core_eu_ea_alu_ea_reg_afrwe_DO_reg[7]/P0001  ;
  assign n13960 = \core_c_psq_MSTAT_reg_DO_reg[0]/P0002  & ~\core_eu_ea_alu_ea_reg_afswe_DO_reg[7]/P0001  ;
  assign n13961 = ~n13959 & ~n13960 ;
  assign n13962 = \core_c_dec_IRE_reg[12]/NET0131  & ~n13961 ;
  assign n13958 = ~\core_c_dec_IRE_reg[12]/NET0131  & n11054 ;
  assign n13963 = ~\core_c_dec_IRE_reg[11]/NET0131  & ~n13958 ;
  assign n13964 = ~n13962 & n13963 ;
  assign n13957 = ~n11058 & n13881 ;
  assign n13965 = ~n13878 & ~n13957 ;
  assign n13966 = ~n13964 & n13965 ;
  assign n13956 = ~\core_eu_ea_alu_ea_dec_piconst_DO_reg[7]/P0001  & n13878 ;
  assign n13967 = n13880 & ~n13956 ;
  assign n13968 = ~n13966 & n13967 ;
  assign n13969 = n13895 & ~n13968 ;
  assign n13970 = n13874 & n13968 ;
  assign n13971 = ~n13969 & ~n13970 ;
  assign n13972 = ~n13955 & ~n13971 ;
  assign n13975 = \core_c_dec_IRE_reg[8]/NET0131  & n11311 ;
  assign n13974 = ~\core_c_dec_IRE_reg[8]/NET0131  & n11315 ;
  assign n13976 = n13823 & ~n13974 ;
  assign n13977 = ~n13975 & n13976 ;
  assign n13973 = ~n11424 & n13813 ;
  assign n13978 = ~n11341 & n13816 ;
  assign n13981 = ~n13973 & ~n13978 ;
  assign n13979 = ~n11444 & n13819 ;
  assign n13980 = ~n11448 & n13821 ;
  assign n13982 = ~n13979 & ~n13980 ;
  assign n13983 = n13981 & n13982 ;
  assign n13984 = ~n13977 & n13983 ;
  assign n13986 = \core_c_dec_IRE_reg[8]/NET0131  & n11337 ;
  assign n13985 = ~\core_c_dec_IRE_reg[8]/NET0131  & n11325 ;
  assign n13987 = n13832 & ~n13985 ;
  assign n13988 = ~n13986 & n13987 ;
  assign n13989 = n13984 & ~n13988 ;
  assign n13990 = n13853 & ~n13989 ;
  assign n13991 = n13848 & ~n13990 ;
  assign n13992 = ~n13848 & n13990 ;
  assign n13993 = ~n13991 & ~n13992 ;
  assign n13997 = ~\core_c_psq_MSTAT_reg_DO_reg[0]/P0002  & ~\core_eu_ea_alu_ea_reg_afrwe_DO_reg[6]/P0001  ;
  assign n13998 = \core_c_psq_MSTAT_reg_DO_reg[0]/P0002  & ~\core_eu_ea_alu_ea_reg_afswe_DO_reg[6]/P0001  ;
  assign n13999 = ~n13997 & ~n13998 ;
  assign n14000 = \core_c_dec_IRE_reg[12]/NET0131  & ~n13999 ;
  assign n13996 = ~\core_c_dec_IRE_reg[12]/NET0131  & n11329 ;
  assign n14001 = ~\core_c_dec_IRE_reg[11]/NET0131  & ~n13996 ;
  assign n14002 = ~n14000 & n14001 ;
  assign n13995 = ~n11333 & n13881 ;
  assign n14003 = ~n13878 & ~n13995 ;
  assign n14004 = ~n14002 & n14003 ;
  assign n13994 = ~\core_eu_ea_alu_ea_dec_piconst_DO_reg[6]/P0001  & n13878 ;
  assign n14005 = n13880 & ~n13994 ;
  assign n14006 = ~n14004 & n14005 ;
  assign n14007 = n13895 & ~n14006 ;
  assign n14008 = n13874 & n14006 ;
  assign n14009 = ~n14007 & ~n14008 ;
  assign n14010 = ~n13993 & ~n14009 ;
  assign n14271 = ~n13972 & ~n14010 ;
  assign n14272 = ~n14270 & n14271 ;
  assign n14273 = n13955 & n13971 ;
  assign n14274 = n13993 & n14009 ;
  assign n14275 = ~n13972 & n14274 ;
  assign n14276 = ~n14273 & ~n14275 ;
  assign n14277 = ~n14272 & n14276 ;
  assign n13858 = \core_c_dec_IRE_reg[8]/NET0131  & n10226 ;
  assign n13857 = ~\core_c_dec_IRE_reg[8]/NET0131  & n10218 ;
  assign n13859 = n13823 & ~n13857 ;
  assign n13860 = ~n13858 & n13859 ;
  assign n13854 = ~n10191 & n13816 ;
  assign n13861 = ~n13814 & ~n13854 ;
  assign n13855 = ~n10112 & n13819 ;
  assign n13856 = ~n10096 & n13821 ;
  assign n13862 = ~n13855 & ~n13856 ;
  assign n13863 = n13861 & n13862 ;
  assign n13864 = ~n13860 & n13863 ;
  assign n13866 = \core_c_dec_IRE_reg[8]/NET0131  & n10179 ;
  assign n13865 = ~\core_c_dec_IRE_reg[8]/NET0131  & n10187 ;
  assign n13867 = n13832 & ~n13865 ;
  assign n13868 = ~n13866 & n13867 ;
  assign n13869 = n13864 & ~n13868 ;
  assign n13870 = n13853 & ~n13869 ;
  assign n13871 = n13848 & ~n13870 ;
  assign n13872 = ~n13848 & n13870 ;
  assign n13873 = ~n13871 & ~n13872 ;
  assign n13884 = ~\core_c_psq_MSTAT_reg_DO_reg[0]/P0002  & ~\core_eu_ea_alu_ea_reg_afrwe_DO_reg[9]/P0001  ;
  assign n13885 = \core_c_psq_MSTAT_reg_DO_reg[0]/P0002  & ~\core_eu_ea_alu_ea_reg_afswe_DO_reg[9]/P0001  ;
  assign n13886 = ~n13884 & ~n13885 ;
  assign n13887 = \core_c_dec_IRE_reg[12]/NET0131  & ~n13886 ;
  assign n13883 = ~\core_c_dec_IRE_reg[12]/NET0131  & n10183 ;
  assign n13888 = ~\core_c_dec_IRE_reg[11]/NET0131  & ~n13883 ;
  assign n13889 = ~n13887 & n13888 ;
  assign n13882 = ~n10175 & n13881 ;
  assign n13890 = ~n13878 & ~n13882 ;
  assign n13891 = ~n13889 & n13890 ;
  assign n13879 = ~\core_eu_ea_alu_ea_dec_piconst_DO_reg[9]/P0001  & n13878 ;
  assign n13892 = ~n13879 & n13880 ;
  assign n13893 = ~n13891 & n13892 ;
  assign n13894 = ~n13874 & n13893 ;
  assign n13896 = ~n13893 & ~n13895 ;
  assign n13897 = ~n13894 & ~n13896 ;
  assign n13898 = ~n13873 & n13897 ;
  assign n13903 = \core_c_dec_IRE_reg[8]/NET0131  & n10575 ;
  assign n13902 = ~\core_c_dec_IRE_reg[8]/NET0131  & n10567 ;
  assign n13904 = n13823 & ~n13902 ;
  assign n13905 = ~n13903 & n13904 ;
  assign n13899 = ~n10461 & n13816 ;
  assign n13906 = ~n13814 & ~n13899 ;
  assign n13900 = ~n10534 & n13819 ;
  assign n13901 = ~n10538 & n13821 ;
  assign n13907 = ~n13900 & ~n13901 ;
  assign n13908 = n13906 & n13907 ;
  assign n13909 = ~n13905 & n13908 ;
  assign n13911 = \core_c_dec_IRE_reg[8]/NET0131  & n10457 ;
  assign n13910 = ~\core_c_dec_IRE_reg[8]/NET0131  & n10449 ;
  assign n13912 = n13832 & ~n13910 ;
  assign n13913 = ~n13911 & n13912 ;
  assign n13914 = n13909 & ~n13913 ;
  assign n13915 = n13853 & ~n13914 ;
  assign n13916 = n13848 & ~n13915 ;
  assign n13917 = ~n13848 & n13915 ;
  assign n13918 = ~n13916 & ~n13917 ;
  assign n13922 = ~\core_c_psq_MSTAT_reg_DO_reg[0]/P0002  & ~\core_eu_ea_alu_ea_reg_afrwe_DO_reg[8]/P0001  ;
  assign n13923 = \core_c_psq_MSTAT_reg_DO_reg[0]/P0002  & ~\core_eu_ea_alu_ea_reg_afswe_DO_reg[8]/P0001  ;
  assign n13924 = ~n13922 & ~n13923 ;
  assign n13925 = \core_c_dec_IRE_reg[12]/NET0131  & ~n13924 ;
  assign n13921 = ~\core_c_dec_IRE_reg[12]/NET0131  & n10453 ;
  assign n13926 = ~\core_c_dec_IRE_reg[11]/NET0131  & ~n13921 ;
  assign n13927 = ~n13925 & n13926 ;
  assign n13920 = ~n10445 & n13881 ;
  assign n13928 = ~n13878 & ~n13920 ;
  assign n13929 = ~n13927 & n13928 ;
  assign n13919 = ~\core_eu_ea_alu_ea_dec_piconst_DO_reg[8]/P0001  & n13878 ;
  assign n13930 = n13880 & ~n13919 ;
  assign n13931 = ~n13929 & n13930 ;
  assign n13932 = n13895 & ~n13931 ;
  assign n13933 = n13874 & n13931 ;
  assign n13934 = ~n13932 & ~n13933 ;
  assign n13935 = ~n13918 & ~n13934 ;
  assign n14278 = ~n13898 & ~n13935 ;
  assign n14279 = ~n14277 & n14278 ;
  assign n14284 = \core_c_dec_IRE_reg[8]/NET0131  & n8410 ;
  assign n14283 = ~\core_c_dec_IRE_reg[8]/NET0131  & n8402 ;
  assign n14285 = n13823 & ~n14283 ;
  assign n14286 = ~n14284 & n14285 ;
  assign n14280 = ~n8354 & n13819 ;
  assign n14287 = ~n13814 & ~n14280 ;
  assign n14281 = ~n8358 & n13821 ;
  assign n14282 = ~n8385 & n13816 ;
  assign n14288 = ~n14281 & ~n14282 ;
  assign n14289 = n14287 & n14288 ;
  assign n14290 = ~n14286 & n14289 ;
  assign n14292 = \core_c_dec_IRE_reg[8]/NET0131  & n8373 ;
  assign n14291 = ~\core_c_dec_IRE_reg[8]/NET0131  & n8369 ;
  assign n14293 = n13832 & ~n14291 ;
  assign n14294 = ~n14292 & n14293 ;
  assign n14295 = n14290 & ~n14294 ;
  assign n14296 = n13853 & ~n14295 ;
  assign n14297 = ~n13848 & n14296 ;
  assign n14298 = n13848 & ~n14296 ;
  assign n14299 = ~n14297 & ~n14298 ;
  assign n14303 = ~\core_c_psq_MSTAT_reg_DO_reg[0]/P0002  & ~\core_eu_ea_alu_ea_reg_afrwe_DO_reg[11]/P0001  ;
  assign n14304 = \core_c_psq_MSTAT_reg_DO_reg[0]/P0002  & ~\core_eu_ea_alu_ea_reg_afswe_DO_reg[11]/P0001  ;
  assign n14305 = ~n14303 & ~n14304 ;
  assign n14306 = \core_c_dec_IRE_reg[12]/NET0131  & ~n14305 ;
  assign n14302 = ~\core_c_dec_IRE_reg[12]/NET0131  & n8377 ;
  assign n14307 = ~\core_c_dec_IRE_reg[11]/NET0131  & ~n14302 ;
  assign n14308 = ~n14306 & n14307 ;
  assign n14301 = ~n8381 & n13881 ;
  assign n14309 = ~n13878 & ~n14301 ;
  assign n14310 = ~n14308 & n14309 ;
  assign n14300 = ~\core_eu_ea_alu_ea_dec_piconst_DO_reg[11]/P0001  & n13878 ;
  assign n14311 = n13880 & ~n14300 ;
  assign n14312 = ~n14310 & n14311 ;
  assign n14313 = ~n13874 & n14312 ;
  assign n14314 = ~n13895 & ~n14312 ;
  assign n14315 = ~n14313 & ~n14314 ;
  assign n14316 = ~n14299 & n14315 ;
  assign n14317 = n13918 & n13934 ;
  assign n14318 = ~n14316 & n14317 ;
  assign n14319 = n13873 & ~n13897 ;
  assign n14320 = ~n14318 & ~n14319 ;
  assign n14321 = ~n14279 & n14320 ;
  assign n14326 = \core_c_dec_IRE_reg[8]/NET0131  & n7809 ;
  assign n14325 = ~\core_c_dec_IRE_reg[8]/NET0131  & n7801 ;
  assign n14327 = n13823 & ~n14325 ;
  assign n14328 = ~n14326 & n14327 ;
  assign n14322 = ~n7753 & n13819 ;
  assign n14329 = ~n13814 & ~n14322 ;
  assign n14323 = ~n7737 & n13821 ;
  assign n14324 = ~n7784 & n13816 ;
  assign n14330 = ~n14323 & ~n14324 ;
  assign n14331 = n14329 & n14330 ;
  assign n14332 = ~n14328 & n14331 ;
  assign n14334 = \core_c_dec_IRE_reg[8]/NET0131  & n7780 ;
  assign n14333 = ~\core_c_dec_IRE_reg[8]/NET0131  & n7768 ;
  assign n14335 = n13832 & ~n14333 ;
  assign n14336 = ~n14334 & n14335 ;
  assign n14337 = n14332 & ~n14336 ;
  assign n14338 = n13853 & ~n14337 ;
  assign n14339 = n13848 & ~n14338 ;
  assign n14340 = ~n13848 & n14338 ;
  assign n14341 = ~n14339 & ~n14340 ;
  assign n14345 = ~\core_c_psq_MSTAT_reg_DO_reg[0]/P0002  & ~\core_eu_ea_alu_ea_reg_afrwe_DO_reg[10]/P0001  ;
  assign n14346 = \core_c_psq_MSTAT_reg_DO_reg[0]/P0002  & ~\core_eu_ea_alu_ea_reg_afswe_DO_reg[10]/P0001  ;
  assign n14347 = ~n14345 & ~n14346 ;
  assign n14348 = \core_c_dec_IRE_reg[12]/NET0131  & ~n14347 ;
  assign n14344 = ~\core_c_dec_IRE_reg[12]/NET0131  & n7776 ;
  assign n14349 = ~\core_c_dec_IRE_reg[11]/NET0131  & ~n14344 ;
  assign n14350 = ~n14348 & n14349 ;
  assign n14343 = ~n7772 & n13881 ;
  assign n14351 = ~n13878 & ~n14343 ;
  assign n14352 = ~n14350 & n14351 ;
  assign n14342 = ~\core_eu_ea_alu_ea_dec_piconst_DO_reg[10]/P0001  & n13878 ;
  assign n14353 = n13880 & ~n14342 ;
  assign n14354 = ~n14352 & n14353 ;
  assign n14355 = ~n13874 & n14354 ;
  assign n14356 = ~n13895 & ~n14354 ;
  assign n14357 = ~n14355 & ~n14356 ;
  assign n14358 = ~n14341 & n14357 ;
  assign n14359 = ~n14316 & ~n14358 ;
  assign n14360 = ~n14321 & n14359 ;
  assign n14361 = n14299 & ~n14315 ;
  assign n14362 = n14341 & ~n14357 ;
  assign n14363 = ~n13898 & n14362 ;
  assign n14364 = ~n14361 & ~n14363 ;
  assign n14365 = ~n14360 & n14364 ;
  assign n14366 = ~n13809 & ~n14365 ;
  assign n14371 = \core_c_dec_IRE_reg[8]/NET0131  & n9128 ;
  assign n14370 = ~\core_c_dec_IRE_reg[8]/NET0131  & n9120 ;
  assign n14372 = n13823 & ~n14370 ;
  assign n14373 = ~n14371 & n14372 ;
  assign n14367 = ~n9072 & n13819 ;
  assign n14374 = ~n13814 & ~n14367 ;
  assign n14368 = ~n9056 & n13821 ;
  assign n14369 = ~n9103 & n13816 ;
  assign n14375 = ~n14368 & ~n14369 ;
  assign n14376 = n14374 & n14375 ;
  assign n14377 = ~n14373 & n14376 ;
  assign n14379 = \core_c_dec_IRE_reg[8]/NET0131  & n9099 ;
  assign n14378 = ~\core_c_dec_IRE_reg[8]/NET0131  & n9091 ;
  assign n14380 = n13832 & ~n14378 ;
  assign n14381 = ~n14379 & n14380 ;
  assign n14382 = n14377 & ~n14381 ;
  assign n14383 = n13853 & ~n14382 ;
  assign n14384 = n13848 & ~n14383 ;
  assign n14385 = ~n13848 & n14383 ;
  assign n14386 = ~n14384 & ~n14385 ;
  assign n14390 = ~\core_c_psq_MSTAT_reg_DO_reg[0]/P0002  & ~\core_eu_ea_alu_ea_reg_afrwe_DO_reg[12]/P0001  ;
  assign n14391 = \core_c_psq_MSTAT_reg_DO_reg[0]/P0002  & ~\core_eu_ea_alu_ea_reg_afswe_DO_reg[12]/P0001  ;
  assign n14392 = ~n14390 & ~n14391 ;
  assign n14393 = \core_c_dec_IRE_reg[12]/NET0131  & ~n14392 ;
  assign n14389 = ~\core_c_dec_IRE_reg[12]/NET0131  & n9095 ;
  assign n14394 = ~\core_c_dec_IRE_reg[11]/NET0131  & ~n14389 ;
  assign n14395 = ~n14393 & n14394 ;
  assign n14388 = ~n9087 & n13881 ;
  assign n14396 = ~n13878 & ~n14388 ;
  assign n14397 = ~n14395 & n14396 ;
  assign n14387 = ~\core_eu_ea_alu_ea_dec_piconst_DO_reg[12]/P0001  & n13878 ;
  assign n14398 = n13880 & ~n14387 ;
  assign n14399 = ~n14397 & n14398 ;
  assign n14400 = n13895 & ~n14399 ;
  assign n14401 = n13874 & n14399 ;
  assign n14402 = ~n14400 & ~n14401 ;
  assign n14403 = n14386 & n14402 ;
  assign n14406 = ~\core_eu_ea_alu_ea_dec_AMF_E_reg[1]/NET0131  & n13808 ;
  assign n14407 = n14403 & ~n14406 ;
  assign n14404 = n13808 & n13843 ;
  assign n14405 = ~n14403 & n14404 ;
  assign n14408 = ~n14386 & ~n14402 ;
  assign n14409 = ~n14405 & ~n14408 ;
  assign n14410 = ~n14407 & n14409 ;
  assign n14411 = n14366 & ~n14410 ;
  assign n14412 = ~n14366 & n14410 ;
  assign n14413 = ~n14411 & ~n14412 ;
  assign n14414 = ~n13806 & n14413 ;
  assign n14416 = ~n14361 & n14404 ;
  assign n14415 = n14361 & ~n14406 ;
  assign n14417 = ~n14316 & ~n14415 ;
  assign n14418 = ~n14416 & n14417 ;
  assign n14419 = n14321 & ~n14362 ;
  assign n14420 = ~n13809 & ~n14358 ;
  assign n14421 = ~n14419 & n14420 ;
  assign n14422 = ~n14418 & n14421 ;
  assign n14423 = n14418 & ~n14421 ;
  assign n14424 = ~n14422 & ~n14423 ;
  assign n14425 = n13806 & n14424 ;
  assign n14426 = ~n14414 & ~n14425 ;
  assign n14427 = n13805 & ~n14426 ;
  assign n14428 = ~\core_eu_ea_alu_ea_reg_afrwe_DO_reg[12]/P0001  & ~n13805 ;
  assign n14429 = ~n14427 & ~n14428 ;
  assign n14438 = \core_c_dec_IRE_reg[8]/NET0131  & n7156 ;
  assign n14437 = ~\core_c_dec_IRE_reg[8]/NET0131  & n7164 ;
  assign n14439 = n13823 & ~n14437 ;
  assign n14440 = ~n14438 & n14439 ;
  assign n14434 = ~n7182 & n13819 ;
  assign n14441 = ~n13814 & ~n14434 ;
  assign n14435 = ~n7202 & n13821 ;
  assign n14436 = ~n7112 & n13816 ;
  assign n14442 = ~n14435 & ~n14436 ;
  assign n14443 = n14441 & n14442 ;
  assign n14444 = ~n14440 & n14443 ;
  assign n14445 = ~n13832 & n14444 ;
  assign n14431 = \core_c_dec_IRE_reg[8]/NET0131  & ~n7100 ;
  assign n14430 = ~\core_c_dec_IRE_reg[8]/NET0131  & ~n7096 ;
  assign n14432 = n13832 & ~n14430 ;
  assign n14433 = ~n14431 & n14432 ;
  assign n14446 = n13853 & ~n14433 ;
  assign n14447 = ~n14445 & n14446 ;
  assign n14448 = n13848 & n14447 ;
  assign n14449 = ~n13848 & ~n14447 ;
  assign n14450 = ~n14448 & ~n14449 ;
  assign n14452 = \core_c_psq_MSTAT_reg_DO_reg[0]/P0002  & ~\core_eu_ea_alu_ea_reg_afswe_DO_reg[13]/P0001  ;
  assign n14451 = ~\core_c_psq_MSTAT_reg_DO_reg[0]/P0002  & ~\core_eu_ea_alu_ea_reg_afrwe_DO_reg[13]/P0001  ;
  assign n14453 = n14033 & ~n14451 ;
  assign n14454 = ~n14452 & n14453 ;
  assign n14456 = \core_c_dec_IRE_reg[11]/NET0131  & n7108 ;
  assign n14455 = ~\core_c_dec_IRE_reg[11]/NET0131  & n7104 ;
  assign n14457 = ~\core_c_dec_IRE_reg[12]/NET0131  & ~n14455 ;
  assign n14458 = ~n14456 & n14457 ;
  assign n14459 = ~n14454 & ~n14458 ;
  assign n14460 = ~n13878 & ~n14459 ;
  assign n14461 = \core_eu_ea_alu_ea_dec_piconst_DO_reg[13]/P0001  & n13878 ;
  assign n14462 = ~n14460 & ~n14461 ;
  assign n14464 = n13874 & n14462 ;
  assign n14463 = n14032 & ~n14462 ;
  assign n14465 = ~n13840 & ~n14463 ;
  assign n14466 = ~n14464 & n14465 ;
  assign n14467 = n14450 & n14466 ;
  assign n14468 = ~n14408 & ~n14467 ;
  assign n14469 = ~n14365 & n14468 ;
  assign n14470 = ~n14450 & ~n14466 ;
  assign n14471 = ~n13837 & n13853 ;
  assign n14472 = n13848 & ~n14471 ;
  assign n14473 = ~n13848 & n14471 ;
  assign n14474 = ~n14472 & ~n14473 ;
  assign n14476 = \core_c_dec_IRE_reg[11]/NET0131  & n11979 ;
  assign n14475 = ~\core_c_dec_IRE_reg[11]/NET0131  & n11975 ;
  assign n14477 = ~\core_c_dec_IRE_reg[12]/NET0131  & ~n14475 ;
  assign n14478 = ~n14476 & n14477 ;
  assign n14480 = \core_c_psq_MSTAT_reg_DO_reg[0]/P0002  & ~\core_eu_ea_alu_ea_reg_afswe_DO_reg[15]/P0001  ;
  assign n14479 = ~\core_c_psq_MSTAT_reg_DO_reg[0]/P0002  & ~\core_eu_ea_alu_ea_reg_afrwe_DO_reg[15]/P0001  ;
  assign n14481 = n14033 & ~n14479 ;
  assign n14482 = ~n14480 & n14481 ;
  assign n14483 = ~n13878 & ~n14482 ;
  assign n14484 = ~n14478 & n14483 ;
  assign n14485 = ~\core_eu_ea_alu_ea_dec_piconst_DO_reg[15]/P0001  & n13878 ;
  assign n14486 = ~n14484 & ~n14485 ;
  assign n14487 = n13880 & n14486 ;
  assign n14488 = ~n13874 & n14487 ;
  assign n14489 = ~n13895 & ~n14487 ;
  assign n14490 = ~n14488 & ~n14489 ;
  assign n14491 = ~n14474 & n14490 ;
  assign n14492 = n14403 & ~n14491 ;
  assign n14493 = ~n14470 & ~n14492 ;
  assign n14494 = ~n14469 & n14493 ;
  assign n14495 = ~n13809 & ~n14494 ;
  assign n14500 = \core_c_dec_IRE_reg[8]/NET0131  & n11854 ;
  assign n14499 = ~\core_c_dec_IRE_reg[8]/NET0131  & n11846 ;
  assign n14501 = n13823 & ~n14499 ;
  assign n14502 = ~n14500 & n14501 ;
  assign n14496 = ~n11837 & n13816 ;
  assign n14503 = ~n13814 & ~n14496 ;
  assign n14497 = ~n11878 & n13819 ;
  assign n14498 = ~n11882 & n13821 ;
  assign n14504 = ~n14497 & ~n14498 ;
  assign n14505 = n14503 & n14504 ;
  assign n14506 = ~n14502 & n14505 ;
  assign n14508 = \core_c_dec_IRE_reg[8]/NET0131  & n11825 ;
  assign n14507 = ~\core_c_dec_IRE_reg[8]/NET0131  & n11821 ;
  assign n14509 = n13832 & ~n14507 ;
  assign n14510 = ~n14508 & n14509 ;
  assign n14511 = n14506 & ~n14510 ;
  assign n14512 = n13853 & ~n14511 ;
  assign n14513 = n13848 & ~n14512 ;
  assign n14514 = ~n13848 & n14512 ;
  assign n14515 = ~n14513 & ~n14514 ;
  assign n14519 = ~\core_c_psq_MSTAT_reg_DO_reg[0]/P0002  & ~\core_eu_ea_alu_ea_reg_afrwe_DO_reg[14]/P0001  ;
  assign n14520 = \core_c_psq_MSTAT_reg_DO_reg[0]/P0002  & ~\core_eu_ea_alu_ea_reg_afswe_DO_reg[14]/P0001  ;
  assign n14521 = ~n14519 & ~n14520 ;
  assign n14522 = \core_c_dec_IRE_reg[12]/NET0131  & ~n14521 ;
  assign n14518 = ~\core_c_dec_IRE_reg[12]/NET0131  & n11829 ;
  assign n14523 = ~\core_c_dec_IRE_reg[11]/NET0131  & ~n14518 ;
  assign n14524 = ~n14522 & n14523 ;
  assign n14517 = ~n11833 & n13881 ;
  assign n14525 = ~n13878 & ~n14517 ;
  assign n14526 = ~n14524 & n14525 ;
  assign n14516 = ~\core_eu_ea_alu_ea_dec_piconst_DO_reg[14]/P0001  & n13878 ;
  assign n14527 = n13880 & ~n14516 ;
  assign n14528 = ~n14526 & n14527 ;
  assign n14529 = n13895 & ~n14528 ;
  assign n14530 = n13874 & n14528 ;
  assign n14531 = ~n14529 & ~n14530 ;
  assign n14532 = n14515 & n14531 ;
  assign n14533 = n14406 & n14532 ;
  assign n14534 = ~n14515 & ~n14531 ;
  assign n14535 = ~n14404 & ~n14532 ;
  assign n14536 = ~n14534 & n14535 ;
  assign n14537 = ~n14533 & ~n14536 ;
  assign n14538 = n14495 & ~n14537 ;
  assign n14539 = ~n14495 & n14537 ;
  assign n14540 = ~n14538 & ~n14539 ;
  assign n14541 = ~n13806 & ~n14540 ;
  assign n14543 = ~n14406 & n14470 ;
  assign n14542 = n14404 & ~n14470 ;
  assign n14544 = ~n14467 & ~n14542 ;
  assign n14545 = ~n14543 & n14544 ;
  assign n14546 = n14365 & ~n14403 ;
  assign n14547 = ~n13809 & ~n14408 ;
  assign n14548 = ~n14546 & n14547 ;
  assign n14549 = ~n14545 & n14548 ;
  assign n14550 = n14545 & ~n14548 ;
  assign n14551 = ~n14549 & ~n14550 ;
  assign n14552 = n13806 & n14551 ;
  assign n14553 = ~n14541 & ~n14552 ;
  assign n14554 = n13805 & ~n14553 ;
  assign n14555 = ~\core_eu_ea_alu_ea_reg_afrwe_DO_reg[14]/P0001  & ~n13805 ;
  assign n14556 = ~n14554 & ~n14555 ;
  assign n14557 = ~n13809 & ~n14252 ;
  assign n14559 = ~n14254 & n14404 ;
  assign n14558 = n14254 & ~n14406 ;
  assign n14560 = ~n14243 & ~n14558 ;
  assign n14561 = ~n14559 & n14560 ;
  assign n14562 = n14557 & ~n14561 ;
  assign n14563 = ~n14557 & n14561 ;
  assign n14564 = ~n14562 & ~n14563 ;
  assign n14565 = n13806 & ~n14564 ;
  assign n14566 = ~n13809 & ~n14255 ;
  assign n14567 = n14204 & n14406 ;
  assign n14568 = ~n14204 & ~n14404 ;
  assign n14569 = ~n14244 & n14568 ;
  assign n14570 = ~n14567 & ~n14569 ;
  assign n14571 = n14566 & ~n14570 ;
  assign n14572 = ~n14566 & n14570 ;
  assign n14573 = ~n14571 & ~n14572 ;
  assign n14574 = ~n13806 & n14573 ;
  assign n14575 = ~n14565 & ~n14574 ;
  assign n14576 = n13805 & ~n14575 ;
  assign n14577 = \core_eu_ea_alu_ea_reg_afrwe_DO_reg[1]/P0001  & ~n13805 ;
  assign n14578 = ~n14576 & ~n14577 ;
  assign n14579 = ~n13809 & ~n14257 ;
  assign n14581 = ~n14262 & n14404 ;
  assign n14580 = n14262 & ~n14406 ;
  assign n14582 = ~n14166 & ~n14580 ;
  assign n14583 = ~n14581 & n14582 ;
  assign n14584 = n14579 & ~n14583 ;
  assign n14585 = ~n14579 & n14583 ;
  assign n14586 = ~n14584 & ~n14585 ;
  assign n14587 = ~n13806 & ~n14586 ;
  assign n14588 = n13806 & n14573 ;
  assign n14589 = ~n14587 & ~n14588 ;
  assign n14590 = n13805 & ~n14589 ;
  assign n14591 = \core_eu_ea_alu_ea_reg_afrwe_DO_reg[2]/P0001  & ~n13805 ;
  assign n14592 = ~n14590 & ~n14591 ;
  assign n14593 = ~n13809 & ~n14265 ;
  assign n14595 = ~n14127 & n14404 ;
  assign n14594 = n14127 & ~n14406 ;
  assign n14596 = ~n14266 & ~n14594 ;
  assign n14597 = ~n14595 & n14596 ;
  assign n14598 = n14593 & ~n14597 ;
  assign n14599 = ~n14593 & n14597 ;
  assign n14600 = ~n14598 & ~n14599 ;
  assign n14601 = ~n13806 & ~n14600 ;
  assign n14602 = ~n14258 & ~n14262 ;
  assign n14603 = ~n13809 & ~n14602 ;
  assign n14605 = ~n14260 & n14404 ;
  assign n14604 = n14260 & ~n14406 ;
  assign n14606 = ~n14089 & ~n14604 ;
  assign n14607 = ~n14605 & n14606 ;
  assign n14608 = n14603 & ~n14607 ;
  assign n14609 = ~n14603 & n14607 ;
  assign n14610 = ~n14608 & ~n14609 ;
  assign n14611 = n13806 & ~n14610 ;
  assign n14612 = ~n14601 & ~n14611 ;
  assign n14613 = n13805 & ~n14612 ;
  assign n14614 = \core_eu_ea_alu_ea_reg_afrwe_DO_reg[4]/P0001  & ~n13805 ;
  assign n14615 = ~n14613 & ~n14614 ;
  assign n14616 = ~n13809 & ~n14270 ;
  assign n14618 = ~n14274 & n14404 ;
  assign n14617 = n14274 & ~n14406 ;
  assign n14619 = ~n14010 & ~n14617 ;
  assign n14620 = ~n14618 & n14619 ;
  assign n14621 = n14616 & ~n14620 ;
  assign n14622 = ~n14616 & n14620 ;
  assign n14623 = ~n14621 & ~n14622 ;
  assign n14624 = ~n13806 & ~n14623 ;
  assign n14626 = ~n14050 & n14404 ;
  assign n14625 = n14050 & ~n14406 ;
  assign n14627 = ~n14261 & ~n14625 ;
  assign n14628 = ~n14626 & n14627 ;
  assign n14629 = ~n14127 & n14265 ;
  assign n14630 = ~n13809 & ~n14266 ;
  assign n14631 = ~n14629 & n14630 ;
  assign n14632 = ~n14628 & n14631 ;
  assign n14633 = n14628 & ~n14631 ;
  assign n14634 = ~n14632 & ~n14633 ;
  assign n14635 = n13806 & ~n14634 ;
  assign n14636 = ~n14624 & ~n14635 ;
  assign n14637 = n13805 & ~n14636 ;
  assign n14638 = \core_eu_ea_alu_ea_reg_afrwe_DO_reg[6]/P0001  & ~n13805 ;
  assign n14639 = ~n14637 & ~n14638 ;
  assign n14641 = ~n14319 & n14404 ;
  assign n14640 = n14319 & ~n14406 ;
  assign n14642 = ~n13898 & ~n14640 ;
  assign n14643 = ~n14641 & n14642 ;
  assign n14644 = n14277 & ~n14317 ;
  assign n14645 = ~n13809 & ~n13935 ;
  assign n14646 = ~n14644 & n14645 ;
  assign n14647 = ~n14643 & n14646 ;
  assign n14648 = n14643 & ~n14646 ;
  assign n14649 = ~n14647 & ~n14648 ;
  assign n14650 = ~n13806 & ~n14649 ;
  assign n14651 = ~n13809 & ~n14277 ;
  assign n14653 = ~n14317 & n14404 ;
  assign n14652 = n14317 & ~n14406 ;
  assign n14654 = ~n13935 & ~n14652 ;
  assign n14655 = ~n14653 & n14654 ;
  assign n14656 = n14651 & ~n14655 ;
  assign n14657 = ~n14651 & n14655 ;
  assign n14658 = ~n14656 & ~n14657 ;
  assign n14659 = n13806 & ~n14658 ;
  assign n14660 = ~n14650 & ~n14659 ;
  assign n14661 = n13805 & ~n14660 ;
  assign n14662 = \core_eu_ea_alu_ea_reg_afrwe_DO_reg[9]/P0001  & ~n13805 ;
  assign n14663 = ~n14661 & ~n14662 ;
  assign n14664 = \core_c_psq_MSTAT_reg_DO_reg[0]/P0002  & ~n5950 ;
  assign n14665 = ~\core_c_dec_Dummy_E_reg/NET0131  & n14664 ;
  assign n14666 = ~n13802 & n14665 ;
  assign n14667 = ~n13800 & n14666 ;
  assign n14668 = ~n14426 & n14667 ;
  assign n14669 = ~\core_eu_ea_alu_ea_reg_afswe_DO_reg[12]/P0001  & ~n14667 ;
  assign n14670 = ~n14668 & ~n14669 ;
  assign n14671 = ~n14553 & n14667 ;
  assign n14672 = ~\core_eu_ea_alu_ea_reg_afswe_DO_reg[14]/P0001  & ~n14667 ;
  assign n14673 = ~n14671 & ~n14672 ;
  assign n14674 = ~n14575 & n14667 ;
  assign n14675 = \core_eu_ea_alu_ea_reg_afswe_DO_reg[1]/P0001  & ~n14667 ;
  assign n14676 = ~n14674 & ~n14675 ;
  assign n14677 = ~n14589 & n14667 ;
  assign n14678 = \core_eu_ea_alu_ea_reg_afswe_DO_reg[2]/P0001  & ~n14667 ;
  assign n14679 = ~n14677 & ~n14678 ;
  assign n14680 = ~n14612 & n14667 ;
  assign n14681 = \core_eu_ea_alu_ea_reg_afswe_DO_reg[4]/P0001  & ~n14667 ;
  assign n14682 = ~n14680 & ~n14681 ;
  assign n14683 = ~n14636 & n14667 ;
  assign n14684 = \core_eu_ea_alu_ea_reg_afswe_DO_reg[6]/P0001  & ~n14667 ;
  assign n14685 = ~n14683 & ~n14684 ;
  assign n14686 = ~n14660 & n14667 ;
  assign n14687 = \core_eu_ea_alu_ea_reg_afswe_DO_reg[9]/P0001  & ~n14667 ;
  assign n14688 = ~n14686 & ~n14687 ;
  assign n14689 = \core_c_dec_MTASTAT_E_reg/P0001  & n11525 ;
  assign n14690 = \core_c_dec_RTI_Ed_reg/P0001  & ~n4184 ;
  assign n14691 = \core_c_dec_IRE_reg[1]/NET0131  & \core_c_dec_Stkctl_Eg_reg/P0001  ;
  assign n14692 = ~n14690 & ~n14691 ;
  assign n14693 = ~\core_c_dec_IRE_reg[0]/NET0131  & ~n14690 ;
  assign n14694 = \core_c_psq_ststk_ptr_reg[0]/NET0131  & \core_c_psq_ststk_ptr_reg[1]/NET0131  ;
  assign n14695 = \core_c_psq_ststk_ptr_reg[2]/NET0131  & n14694 ;
  assign n14696 = ~n14693 & ~n14695 ;
  assign n14697 = ~n14692 & n14696 ;
  assign n14710 = ~\core_c_psq_ststk_ptr_reg[0]/NET0131  & \core_c_psq_ststk_ptr_reg[1]/NET0131  ;
  assign n14713 = ~\core_c_psq_ststk_ptr_reg[2]/NET0131  & n14710 ;
  assign n14714 = \core_c_psq_ststk_sts7x23_STcell_reg[2][6]/P0001  & n14713 ;
  assign n14698 = \core_c_psq_ststk_ptr_reg[0]/NET0131  & ~\core_c_psq_ststk_ptr_reg[1]/NET0131  ;
  assign n14708 = ~\core_c_psq_ststk_ptr_reg[2]/NET0131  & n14698 ;
  assign n14709 = \core_c_psq_ststk_sts7x23_STcell_reg[1][6]/P0001  & n14708 ;
  assign n14711 = \core_c_psq_ststk_ptr_reg[2]/NET0131  & n14710 ;
  assign n14712 = \core_c_psq_ststk_sts7x23_STcell_reg[6][6]/P0001  & n14711 ;
  assign n14717 = ~n14709 & ~n14712 ;
  assign n14718 = ~n14714 & n14717 ;
  assign n14699 = \core_c_psq_ststk_ptr_reg[2]/NET0131  & n14698 ;
  assign n14700 = \core_c_psq_ststk_sts7x23_STcell_reg[5][6]/P0001  & n14699 ;
  assign n14701 = ~\core_c_psq_ststk_ptr_reg[0]/NET0131  & ~\core_c_psq_ststk_ptr_reg[1]/NET0131  ;
  assign n14702 = ~\core_c_psq_ststk_ptr_reg[2]/NET0131  & n14701 ;
  assign n14703 = \core_c_psq_ststk_sts7x23_STcell_reg[0][6]/P0001  & n14702 ;
  assign n14715 = ~n14700 & ~n14703 ;
  assign n14704 = ~\core_c_psq_ststk_ptr_reg[2]/NET0131  & n14694 ;
  assign n14705 = \core_c_psq_ststk_sts7x23_STcell_reg[3][6]/P0001  & n14704 ;
  assign n14706 = \core_c_psq_ststk_ptr_reg[2]/NET0131  & n14701 ;
  assign n14707 = \core_c_psq_ststk_sts7x23_STcell_reg[4][6]/P0001  & n14706 ;
  assign n14716 = ~n14705 & ~n14707 ;
  assign n14719 = n14715 & n14716 ;
  assign n14720 = n14718 & n14719 ;
  assign n14721 = n14697 & ~n14720 ;
  assign n14722 = ~n14689 & ~n14721 ;
  assign n14723 = ~n5950 & ~n14722 ;
  assign n14724 = \core_eu_ec_cun_MVi_pre_C_reg/P0001  & n5950 ;
  assign n14725 = ~n14723 & ~n14724 ;
  assign n14727 = n6022 & n6026 ;
  assign n14728 = ~\core_c_dec_IR_reg[19]/NET0131  & n14727 ;
  assign n14729 = ~n4117 & ~n14728 ;
  assign n14726 = ~\core_eu_em_mac_em_reg_Sq_E_reg/P0001  & n4117 ;
  assign n14730 = ~n4121 & ~n14726 ;
  assign n14731 = ~n14729 & n14730 ;
  assign n14733 = ~\emc_EXTC_Eg_syn_reg/P0001  & n4068 ;
  assign n14734 = n5508 & ~n14733 ;
  assign n14732 = ~\memc_Dread_E_reg/NET0131  & ~\memc_IOcmd_E_reg/NET0131  ;
  assign n14735 = n5432 & ~n14732 ;
  assign n14736 = n14734 & n14735 ;
  assign n14737 = ~n12441 & n14736 ;
  assign n14738 = \emc_DMDreg_reg[8]/P0001  & ~n14737 ;
  assign n14739 = \T_ED[8]_pad  & n14737 ;
  assign n14740 = ~n14738 & ~n14739 ;
  assign n14741 = \emc_DMDreg_reg[9]/P0001  & ~n14737 ;
  assign n14742 = \T_ED[9]_pad  & n14737 ;
  assign n14743 = ~n14741 & ~n14742 ;
  assign n14744 = \memc_Pread_E_reg/NET0131  & n5434 ;
  assign n14745 = n14734 & n14744 ;
  assign n14746 = \emc_PMDreg_reg[8]/P0001  & ~n14745 ;
  assign n14747 = \T_ED[8]_pad  & n14745 ;
  assign n14748 = ~n14746 & ~n14747 ;
  assign n14749 = \emc_PMDreg_reg[9]/P0001  & ~n14745 ;
  assign n14750 = \T_ED[9]_pad  & n14745 ;
  assign n14751 = ~n14749 & ~n14750 ;
  assign n14752 = \core_c_dec_updMR_E_reg/P0001  & n13804 ;
  assign n14753 = ~\core_eu_em_mac_em_dec_emcorepi_DO_reg[3]/P0001  & \core_eu_em_mac_em_reg_mxopwe_DO_reg[15]/P0001  ;
  assign n14754 = ~\core_eu_em_mac_em_reg_myopwe_DO_reg[1]/P0001  & ~\core_eu_em_mac_em_reg_myopwe_DO_reg[2]/P0001  ;
  assign n14755 = \core_eu_em_mac_em_reg_myopwe_DO_reg[1]/P0001  & \core_eu_em_mac_em_reg_myopwe_DO_reg[2]/P0001  ;
  assign n14756 = ~n14754 & ~n14755 ;
  assign n14757 = ~\core_eu_em_mac_em_reg_myopwe_DO_reg[3]/P0001  & n14756 ;
  assign n14758 = \core_eu_em_mac_em_dec_emcorepi_DO_reg[10]/P0001  & n14757 ;
  assign n14759 = \core_eu_em_mac_em_reg_myopwe_DO_reg[3]/P0001  & n14756 ;
  assign n14760 = ~\core_eu_em_mac_em_dec_emcorepi_DO_reg[10]/P0001  & n14759 ;
  assign n14761 = ~n14758 & ~n14760 ;
  assign n14762 = ~n14753 & ~n14761 ;
  assign n14763 = ~\core_eu_em_mac_em_dec_emcorepi_DO_reg[10]/P0001  & n14757 ;
  assign n14764 = \core_eu_em_mac_em_dec_emcorepi_DO_reg[10]/P0001  & n14759 ;
  assign n14765 = ~n14763 & ~n14764 ;
  assign n14766 = n14753 & ~n14765 ;
  assign n14767 = ~n14762 & ~n14766 ;
  assign n14768 = \core_eu_em_mac_em_reg_myopwe_DO_reg[3]/P0001  & n14754 ;
  assign n14769 = ~\core_eu_em_mac_em_dec_emcorepi_DO_reg[10]/P0001  & ~n14768 ;
  assign n14770 = ~\core_eu_em_mac_em_reg_myopwe_DO_reg[3]/P0001  & n14755 ;
  assign n14771 = \core_eu_em_mac_em_dec_emcorepi_DO_reg[10]/P0001  & ~n14770 ;
  assign n14772 = ~n14769 & ~n14771 ;
  assign n14773 = ~n14753 & n14772 ;
  assign n14774 = \core_eu_em_mac_em_dec_emcorepi_DO_reg[10]/P0001  & ~n14768 ;
  assign n14775 = ~\core_eu_em_mac_em_dec_emcorepi_DO_reg[10]/P0001  & ~n14770 ;
  assign n14776 = ~n14774 & ~n14775 ;
  assign n14777 = n14753 & n14776 ;
  assign n14778 = ~n14773 & ~n14777 ;
  assign n14779 = n14767 & n14778 ;
  assign n14780 = ~\core_eu_em_mac_em_reg_myopwe_DO_reg[3]/P0001  & ~\core_eu_em_mac_em_reg_myopwe_DO_reg[4]/P0001  ;
  assign n14781 = \core_eu_em_mac_em_reg_myopwe_DO_reg[3]/P0001  & \core_eu_em_mac_em_reg_myopwe_DO_reg[4]/P0001  ;
  assign n14782 = ~n14780 & ~n14781 ;
  assign n14783 = ~\core_eu_em_mac_em_reg_myopwe_DO_reg[5]/P0001  & n14782 ;
  assign n14784 = \core_eu_em_mac_em_dec_emcorepi_DO_reg[10]/P0001  & n14783 ;
  assign n14785 = \core_eu_em_mac_em_reg_myopwe_DO_reg[5]/P0001  & n14782 ;
  assign n14786 = ~\core_eu_em_mac_em_dec_emcorepi_DO_reg[10]/P0001  & n14785 ;
  assign n14787 = ~n14784 & ~n14786 ;
  assign n14788 = ~n14753 & ~n14787 ;
  assign n14789 = ~\core_eu_em_mac_em_dec_emcorepi_DO_reg[10]/P0001  & n14783 ;
  assign n14790 = \core_eu_em_mac_em_dec_emcorepi_DO_reg[10]/P0001  & n14785 ;
  assign n14791 = ~n14789 & ~n14790 ;
  assign n14792 = n14753 & ~n14791 ;
  assign n14793 = ~n14788 & ~n14792 ;
  assign n14794 = \core_eu_em_mac_em_reg_myopwe_DO_reg[5]/P0001  & n14780 ;
  assign n14795 = ~\core_eu_em_mac_em_dec_emcorepi_DO_reg[10]/P0001  & ~n14794 ;
  assign n14796 = ~\core_eu_em_mac_em_reg_myopwe_DO_reg[5]/P0001  & n14781 ;
  assign n14797 = \core_eu_em_mac_em_dec_emcorepi_DO_reg[10]/P0001  & ~n14796 ;
  assign n14798 = ~n14795 & ~n14797 ;
  assign n14799 = ~n14753 & n14798 ;
  assign n14800 = \core_eu_em_mac_em_dec_emcorepi_DO_reg[10]/P0001  & ~n14794 ;
  assign n14801 = ~\core_eu_em_mac_em_dec_emcorepi_DO_reg[10]/P0001  & ~n14796 ;
  assign n14802 = ~n14800 & ~n14801 ;
  assign n14803 = n14753 & n14802 ;
  assign n14804 = ~n14799 & ~n14803 ;
  assign n14805 = n14793 & n14804 ;
  assign n14806 = n14779 & n14805 ;
  assign n14807 = \core_eu_em_mac_em_reg_myopwe_DO_reg[5]/P0001  & \core_eu_em_mac_em_reg_myopwe_DO_reg[6]/P0001  ;
  assign n14808 = ~\core_eu_em_mac_em_reg_myopwe_DO_reg[5]/P0001  & ~\core_eu_em_mac_em_reg_myopwe_DO_reg[6]/P0001  ;
  assign n14809 = ~n14807 & ~n14808 ;
  assign n14810 = ~\core_eu_em_mac_em_reg_myopwe_DO_reg[7]/P0001  & n14809 ;
  assign n14811 = \core_eu_em_mac_em_dec_emcorepi_DO_reg[10]/P0001  & n14810 ;
  assign n14812 = \core_eu_em_mac_em_reg_myopwe_DO_reg[7]/P0001  & n14809 ;
  assign n14813 = ~\core_eu_em_mac_em_dec_emcorepi_DO_reg[10]/P0001  & n14812 ;
  assign n14814 = ~n14811 & ~n14813 ;
  assign n14815 = ~n14753 & ~n14814 ;
  assign n14816 = \core_eu_em_mac_em_dec_emcorepi_DO_reg[10]/P0001  & n14812 ;
  assign n14817 = ~\core_eu_em_mac_em_dec_emcorepi_DO_reg[10]/P0001  & n14810 ;
  assign n14818 = ~n14816 & ~n14817 ;
  assign n14819 = n14753 & ~n14818 ;
  assign n14820 = ~n14815 & ~n14819 ;
  assign n14821 = \core_eu_em_mac_em_reg_myopwe_DO_reg[7]/P0001  & n14808 ;
  assign n14822 = ~\core_eu_em_mac_em_dec_emcorepi_DO_reg[10]/P0001  & ~n14821 ;
  assign n14823 = ~\core_eu_em_mac_em_reg_myopwe_DO_reg[7]/P0001  & n14807 ;
  assign n14824 = \core_eu_em_mac_em_dec_emcorepi_DO_reg[10]/P0001  & ~n14823 ;
  assign n14825 = ~n14822 & ~n14824 ;
  assign n14826 = ~n14753 & n14825 ;
  assign n14827 = ~\core_eu_em_mac_em_dec_emcorepi_DO_reg[10]/P0001  & ~n14823 ;
  assign n14828 = \core_eu_em_mac_em_dec_emcorepi_DO_reg[10]/P0001  & ~n14821 ;
  assign n14829 = ~n14827 & ~n14828 ;
  assign n14830 = n14753 & n14829 ;
  assign n14831 = ~n14826 & ~n14830 ;
  assign n14832 = n14820 & n14831 ;
  assign n14833 = n14806 & n14832 ;
  assign n14834 = \core_eu_em_mac_em_reg_myopwe_DO_reg[0]/P0001  & \core_eu_em_mac_em_reg_myopwe_DO_reg[1]/P0001  ;
  assign n14835 = ~\core_eu_em_mac_em_dec_emcorepi_DO_reg[10]/P0001  & n14834 ;
  assign n14836 = \core_eu_em_mac_em_reg_myopwe_DO_reg[0]/P0001  & ~\core_eu_em_mac_em_reg_myopwe_DO_reg[1]/P0001  ;
  assign n14837 = \core_eu_em_mac_em_dec_emcorepi_DO_reg[10]/P0001  & n14836 ;
  assign n14838 = ~n14835 & ~n14837 ;
  assign n14839 = ~n14753 & ~n14838 ;
  assign n14840 = \core_eu_em_mac_em_dec_emcorepi_DO_reg[10]/P0001  & n14834 ;
  assign n14841 = ~\core_eu_em_mac_em_dec_emcorepi_DO_reg[10]/P0001  & n14836 ;
  assign n14842 = ~n14840 & ~n14841 ;
  assign n14843 = n14753 & ~n14842 ;
  assign n14844 = ~n14839 & ~n14843 ;
  assign n14845 = ~\core_eu_em_mac_em_dec_emcorepi_DO_reg[10]/P0001  & ~\core_eu_em_mac_em_reg_myopwe_DO_reg[0]/P0001  ;
  assign n14846 = \core_eu_em_mac_em_reg_myopwe_DO_reg[1]/P0001  & n14845 ;
  assign n14847 = ~n14753 & n14846 ;
  assign n14848 = \core_eu_em_mac_em_dec_emcorepi_DO_reg[10]/P0001  & ~\core_eu_em_mac_em_reg_myopwe_DO_reg[0]/P0001  ;
  assign n14849 = \core_eu_em_mac_em_reg_myopwe_DO_reg[1]/P0001  & n14848 ;
  assign n14850 = n14753 & n14849 ;
  assign n14851 = ~n14847 & ~n14850 ;
  assign n14852 = n14844 & n14851 ;
  assign n14853 = n14833 & n14852 ;
  assign n14854 = ~\core_eu_em_mac_em_reg_myopwe_DO_reg[7]/P0001  & ~\core_eu_em_mac_em_reg_myopwe_DO_reg[8]/P0001  ;
  assign n14855 = \core_eu_em_mac_em_reg_myopwe_DO_reg[7]/P0001  & \core_eu_em_mac_em_reg_myopwe_DO_reg[8]/P0001  ;
  assign n14856 = ~n14854 & ~n14855 ;
  assign n14857 = ~\core_eu_em_mac_em_reg_myopwe_DO_reg[9]/P0001  & n14856 ;
  assign n14858 = \core_eu_em_mac_em_dec_emcorepi_DO_reg[10]/P0001  & n14857 ;
  assign n14859 = \core_eu_em_mac_em_reg_myopwe_DO_reg[9]/P0001  & n14856 ;
  assign n14860 = ~\core_eu_em_mac_em_dec_emcorepi_DO_reg[10]/P0001  & n14859 ;
  assign n14861 = ~n14858 & ~n14860 ;
  assign n14862 = ~n14753 & ~n14861 ;
  assign n14863 = ~\core_eu_em_mac_em_dec_emcorepi_DO_reg[10]/P0001  & n14857 ;
  assign n14864 = \core_eu_em_mac_em_dec_emcorepi_DO_reg[10]/P0001  & n14859 ;
  assign n14865 = ~n14863 & ~n14864 ;
  assign n14866 = n14753 & ~n14865 ;
  assign n14867 = ~n14862 & ~n14866 ;
  assign n14868 = \core_eu_em_mac_em_reg_myopwe_DO_reg[9]/P0001  & n14854 ;
  assign n14869 = ~\core_eu_em_mac_em_dec_emcorepi_DO_reg[10]/P0001  & ~n14868 ;
  assign n14870 = ~\core_eu_em_mac_em_reg_myopwe_DO_reg[9]/P0001  & n14855 ;
  assign n14871 = \core_eu_em_mac_em_dec_emcorepi_DO_reg[10]/P0001  & ~n14870 ;
  assign n14872 = ~n14869 & ~n14871 ;
  assign n14873 = ~n14753 & n14872 ;
  assign n14874 = \core_eu_em_mac_em_dec_emcorepi_DO_reg[10]/P0001  & ~n14868 ;
  assign n14875 = ~\core_eu_em_mac_em_dec_emcorepi_DO_reg[10]/P0001  & ~n14870 ;
  assign n14876 = ~n14874 & ~n14875 ;
  assign n14877 = n14753 & n14876 ;
  assign n14878 = ~n14873 & ~n14877 ;
  assign n14879 = n14867 & n14878 ;
  assign n14880 = ~\core_eu_em_mac_em_reg_myopwe_DO_reg[10]/P0001  & ~\core_eu_em_mac_em_reg_myopwe_DO_reg[9]/P0001  ;
  assign n14881 = \core_eu_em_mac_em_reg_myopwe_DO_reg[10]/P0001  & \core_eu_em_mac_em_reg_myopwe_DO_reg[9]/P0001  ;
  assign n14882 = ~n14880 & ~n14881 ;
  assign n14883 = ~\core_eu_em_mac_em_reg_myopwe_DO_reg[11]/P0001  & n14882 ;
  assign n14884 = \core_eu_em_mac_em_dec_emcorepi_DO_reg[10]/P0001  & n14883 ;
  assign n14885 = \core_eu_em_mac_em_reg_myopwe_DO_reg[11]/P0001  & n14882 ;
  assign n14886 = ~\core_eu_em_mac_em_dec_emcorepi_DO_reg[10]/P0001  & n14885 ;
  assign n14887 = ~n14884 & ~n14886 ;
  assign n14888 = ~n14753 & ~n14887 ;
  assign n14889 = ~\core_eu_em_mac_em_dec_emcorepi_DO_reg[10]/P0001  & n14883 ;
  assign n14890 = \core_eu_em_mac_em_dec_emcorepi_DO_reg[10]/P0001  & n14885 ;
  assign n14891 = ~n14889 & ~n14890 ;
  assign n14892 = n14753 & ~n14891 ;
  assign n14893 = ~n14888 & ~n14892 ;
  assign n14894 = \core_eu_em_mac_em_reg_myopwe_DO_reg[11]/P0001  & n14880 ;
  assign n14895 = ~\core_eu_em_mac_em_dec_emcorepi_DO_reg[10]/P0001  & ~n14894 ;
  assign n14896 = ~\core_eu_em_mac_em_reg_myopwe_DO_reg[11]/P0001  & n14881 ;
  assign n14897 = \core_eu_em_mac_em_dec_emcorepi_DO_reg[10]/P0001  & ~n14896 ;
  assign n14898 = ~n14895 & ~n14897 ;
  assign n14899 = ~n14753 & n14898 ;
  assign n14900 = \core_eu_em_mac_em_dec_emcorepi_DO_reg[10]/P0001  & ~n14894 ;
  assign n14901 = ~\core_eu_em_mac_em_dec_emcorepi_DO_reg[10]/P0001  & ~n14896 ;
  assign n14902 = ~n14900 & ~n14901 ;
  assign n14903 = n14753 & n14902 ;
  assign n14904 = ~n14899 & ~n14903 ;
  assign n14905 = n14893 & n14904 ;
  assign n14906 = n14879 & n14905 ;
  assign n14907 = \core_eu_em_mac_em_reg_myopwe_DO_reg[11]/P0001  & \core_eu_em_mac_em_reg_myopwe_DO_reg[12]/P0001  ;
  assign n14908 = ~\core_eu_em_mac_em_reg_myopwe_DO_reg[11]/P0001  & ~\core_eu_em_mac_em_reg_myopwe_DO_reg[12]/P0001  ;
  assign n14909 = ~n14907 & ~n14908 ;
  assign n14910 = ~\core_eu_em_mac_em_reg_myopwe_DO_reg[13]/P0001  & n14909 ;
  assign n14911 = \core_eu_em_mac_em_dec_emcorepi_DO_reg[10]/P0001  & n14910 ;
  assign n14912 = \core_eu_em_mac_em_reg_myopwe_DO_reg[13]/P0001  & n14909 ;
  assign n14913 = ~\core_eu_em_mac_em_dec_emcorepi_DO_reg[10]/P0001  & n14912 ;
  assign n14914 = ~n14911 & ~n14913 ;
  assign n14915 = ~n14753 & ~n14914 ;
  assign n14916 = \core_eu_em_mac_em_dec_emcorepi_DO_reg[10]/P0001  & n14912 ;
  assign n14917 = ~\core_eu_em_mac_em_dec_emcorepi_DO_reg[10]/P0001  & n14910 ;
  assign n14918 = ~n14916 & ~n14917 ;
  assign n14919 = n14753 & ~n14918 ;
  assign n14920 = ~n14915 & ~n14919 ;
  assign n14921 = \core_eu_em_mac_em_reg_myopwe_DO_reg[13]/P0001  & n14908 ;
  assign n14922 = ~\core_eu_em_mac_em_dec_emcorepi_DO_reg[10]/P0001  & ~n14921 ;
  assign n14923 = ~\core_eu_em_mac_em_reg_myopwe_DO_reg[13]/P0001  & n14907 ;
  assign n14924 = \core_eu_em_mac_em_dec_emcorepi_DO_reg[10]/P0001  & ~n14923 ;
  assign n14925 = ~n14922 & ~n14924 ;
  assign n14926 = ~n14753 & n14925 ;
  assign n14927 = ~\core_eu_em_mac_em_dec_emcorepi_DO_reg[10]/P0001  & ~n14923 ;
  assign n14928 = \core_eu_em_mac_em_dec_emcorepi_DO_reg[10]/P0001  & ~n14921 ;
  assign n14929 = ~n14927 & ~n14928 ;
  assign n14930 = n14753 & n14929 ;
  assign n14931 = ~n14926 & ~n14930 ;
  assign n14932 = n14920 & n14931 ;
  assign n14933 = n14906 & n14932 ;
  assign n14936 = \core_c_dec_MACop_E_reg/P0001  & ~n9229 ;
  assign n14937 = ~\core_c_psq_MSTAT_reg_DO_reg[4]/NET0131  & ~n14936 ;
  assign n14934 = \core_c_dec_MACop_E_reg/P0001  & ~n7473 ;
  assign n14935 = \core_c_psq_MSTAT_reg_DO_reg[4]/NET0131  & ~n14934 ;
  assign n14938 = ~\core_eu_em_mac_em_dec_emcorepi_DO_reg[1]/P0001  & ~n14935 ;
  assign n14939 = ~n14937 & n14938 ;
  assign n14940 = ~\core_eu_em_mac_em_reg_myopwe_DO_reg[13]/P0001  & ~\core_eu_em_mac_em_reg_myopwe_DO_reg[14]/P0001  ;
  assign n14941 = \core_eu_em_mac_em_reg_myopwe_DO_reg[13]/P0001  & \core_eu_em_mac_em_reg_myopwe_DO_reg[14]/P0001  ;
  assign n14942 = ~n14940 & ~n14941 ;
  assign n14943 = ~\core_eu_em_mac_em_reg_myopwe_DO_reg[15]/P0001  & n14942 ;
  assign n14944 = \core_eu_em_mac_em_dec_emcorepi_DO_reg[10]/P0001  & n14943 ;
  assign n14945 = \core_eu_em_mac_em_reg_myopwe_DO_reg[15]/P0001  & n14942 ;
  assign n14946 = ~\core_eu_em_mac_em_dec_emcorepi_DO_reg[10]/P0001  & n14945 ;
  assign n14947 = ~n14944 & ~n14946 ;
  assign n14948 = ~n14753 & ~n14947 ;
  assign n14949 = ~\core_eu_em_mac_em_dec_emcorepi_DO_reg[10]/P0001  & n14943 ;
  assign n14950 = \core_eu_em_mac_em_dec_emcorepi_DO_reg[10]/P0001  & n14945 ;
  assign n14951 = ~n14949 & ~n14950 ;
  assign n14952 = n14753 & ~n14951 ;
  assign n14953 = ~n14948 & ~n14952 ;
  assign n14954 = \core_eu_em_mac_em_reg_myopwe_DO_reg[15]/P0001  & n14940 ;
  assign n14955 = ~\core_eu_em_mac_em_dec_emcorepi_DO_reg[10]/P0001  & ~n14954 ;
  assign n14956 = ~\core_eu_em_mac_em_reg_myopwe_DO_reg[15]/P0001  & n14941 ;
  assign n14957 = \core_eu_em_mac_em_dec_emcorepi_DO_reg[10]/P0001  & ~n14956 ;
  assign n14958 = ~n14955 & ~n14957 ;
  assign n14959 = ~n14753 & n14958 ;
  assign n14960 = \core_eu_em_mac_em_dec_emcorepi_DO_reg[10]/P0001  & ~n14954 ;
  assign n14961 = ~\core_eu_em_mac_em_dec_emcorepi_DO_reg[10]/P0001  & ~n14956 ;
  assign n14962 = ~n14960 & ~n14961 ;
  assign n14963 = n14753 & n14962 ;
  assign n14964 = ~n14959 & ~n14963 ;
  assign n14965 = n14953 & n14964 ;
  assign n14966 = \core_eu_em_mac_em_dec_emcorepi_DO_reg[2]/P0001  & \core_eu_em_mac_em_reg_myopwe_DO_reg[15]/P0001  ;
  assign n14967 = \core_eu_em_mac_em_dec_emcorepi_DO_reg[10]/P0001  & n14966 ;
  assign n14968 = ~n14753 & n14967 ;
  assign n14969 = ~\core_eu_em_mac_em_dec_emcorepi_DO_reg[10]/P0001  & n14966 ;
  assign n14970 = n14753 & n14969 ;
  assign n14971 = ~n14968 & ~n14970 ;
  assign n14972 = n14965 & n14971 ;
  assign n14973 = ~n14939 & n14972 ;
  assign n14974 = n14939 & ~n14972 ;
  assign n14975 = ~n14973 & ~n14974 ;
  assign n14976 = ~\core_eu_em_mac_em_reg_mxopwe_DO_reg[15]/P0001  & ~n14967 ;
  assign n14977 = \core_eu_em_mac_em_reg_mxopwe_DO_reg[15]/P0001  & ~n14969 ;
  assign n14978 = ~n14976 & ~n14977 ;
  assign n14979 = n14965 & ~n14978 ;
  assign n14980 = ~n14965 & n14978 ;
  assign n14983 = ~\core_c_psq_MSTAT_reg_DO_reg[4]/NET0131  & ~n14934 ;
  assign n14981 = \core_c_dec_MACop_E_reg/P0001  & ~n12028 ;
  assign n14982 = \core_c_psq_MSTAT_reg_DO_reg[4]/NET0131  & ~n14981 ;
  assign n14984 = ~\core_eu_em_mac_em_dec_emcorepi_DO_reg[1]/P0001  & ~n14982 ;
  assign n14985 = ~n14983 & n14984 ;
  assign n14986 = ~n14980 & ~n14985 ;
  assign n14987 = ~n14979 & ~n14986 ;
  assign n14988 = ~n14975 & ~n14987 ;
  assign n14989 = ~n14933 & ~n14988 ;
  assign n14990 = ~n14879 & ~n14905 ;
  assign n14991 = ~n14932 & n14990 ;
  assign n14992 = ~n14933 & ~n14991 ;
  assign n14993 = \core_c_dec_MACop_E_reg/P0001  & ~\core_c_psq_MSTAT_reg_DO_reg[4]/NET0131  ;
  assign n14994 = ~n8534 & n14993 ;
  assign n14995 = \core_c_psq_MSTAT_reg_DO_reg[4]/NET0131  & n14936 ;
  assign n14996 = ~n14994 & ~n14995 ;
  assign n14997 = ~\core_eu_em_mac_em_dec_emcorepi_DO_reg[1]/P0001  & ~n14996 ;
  assign n14998 = n14972 & ~n14997 ;
  assign n14999 = ~n14972 & n14997 ;
  assign n15000 = ~n14998 & ~n14999 ;
  assign n15001 = ~n14974 & ~n15000 ;
  assign n15002 = n14974 & ~n14997 ;
  assign n15003 = ~n15001 & ~n15002 ;
  assign n15004 = n14992 & ~n15003 ;
  assign n15005 = ~n14992 & n15003 ;
  assign n15006 = ~n15004 & ~n15005 ;
  assign n15007 = ~n14989 & ~n15006 ;
  assign n15008 = n14989 & n15006 ;
  assign n15009 = ~n15007 & ~n15008 ;
  assign n15010 = ~n14979 & ~n14980 ;
  assign n15011 = n14985 & ~n15010 ;
  assign n15012 = ~n14985 & n15010 ;
  assign n15013 = ~n15011 & ~n15012 ;
  assign n15014 = ~\core_eu_em_mac_em_reg_mxopwe_DO_reg[14]/P0001  & ~n14967 ;
  assign n15015 = \core_eu_em_mac_em_reg_mxopwe_DO_reg[14]/P0001  & ~n14969 ;
  assign n15016 = ~n15014 & ~n15015 ;
  assign n15017 = ~\core_eu_em_mac_em_reg_mxopwe_DO_reg[15]/P0001  & n14958 ;
  assign n15018 = \core_eu_em_mac_em_reg_mxopwe_DO_reg[15]/P0001  & n14962 ;
  assign n15019 = ~n15017 & ~n15018 ;
  assign n15020 = n14953 & n15019 ;
  assign n15021 = ~n15016 & n15020 ;
  assign n15022 = n15016 & ~n15020 ;
  assign n15025 = ~\core_c_psq_MSTAT_reg_DO_reg[4]/NET0131  & ~n14981 ;
  assign n15023 = \core_c_dec_MACop_E_reg/P0001  & ~n11882 ;
  assign n15024 = \core_c_psq_MSTAT_reg_DO_reg[4]/NET0131  & ~n15023 ;
  assign n15026 = ~\core_eu_em_mac_em_dec_emcorepi_DO_reg[1]/P0001  & ~n15024 ;
  assign n15027 = ~n15025 & n15026 ;
  assign n15028 = ~n15022 & ~n15027 ;
  assign n15029 = ~n15021 & ~n15028 ;
  assign n15030 = n15013 & ~n15029 ;
  assign n15031 = ~n14933 & ~n15030 ;
  assign n15032 = n14975 & n14987 ;
  assign n15033 = ~n14988 & ~n15032 ;
  assign n15034 = n14992 & n15033 ;
  assign n15035 = ~n14992 & ~n15033 ;
  assign n15036 = ~n15034 & ~n15035 ;
  assign n15037 = ~n15031 & n15036 ;
  assign n15038 = ~n14991 & ~n15032 ;
  assign n15039 = ~n15036 & n15038 ;
  assign n15040 = ~n15037 & ~n15039 ;
  assign n15041 = n15009 & ~n15040 ;
  assign n15042 = ~n14853 & ~n15041 ;
  assign n15043 = ~n14933 & ~n15001 ;
  assign n15044 = \core_c_dec_MACop_E_reg/P0001  & \core_c_psq_MSTAT_reg_DO_reg[4]/NET0131  ;
  assign n15045 = ~n8534 & n15044 ;
  assign n15046 = \core_c_dec_MACop_E_reg/P0001  & ~n7905 ;
  assign n15047 = ~\core_c_psq_MSTAT_reg_DO_reg[4]/NET0131  & n15046 ;
  assign n15048 = ~n15045 & ~n15047 ;
  assign n15049 = ~\core_eu_em_mac_em_dec_emcorepi_DO_reg[1]/P0001  & ~n15048 ;
  assign n15050 = n14972 & ~n15049 ;
  assign n15051 = ~n14972 & n15049 ;
  assign n15052 = ~n15050 & ~n15051 ;
  assign n15053 = ~n14999 & ~n15052 ;
  assign n15054 = n14999 & n15048 ;
  assign n15055 = ~n15053 & ~n15054 ;
  assign n15056 = n14992 & ~n15055 ;
  assign n15057 = ~n14992 & n15055 ;
  assign n15058 = ~n15056 & ~n15057 ;
  assign n15059 = ~n15043 & ~n15058 ;
  assign n15060 = n15043 & n15058 ;
  assign n15061 = ~n15059 & ~n15060 ;
  assign n15062 = ~n14991 & ~n15002 ;
  assign n15063 = n15006 & n15062 ;
  assign n15064 = ~n15007 & ~n15063 ;
  assign n15065 = n15061 & ~n15064 ;
  assign n15066 = ~n15061 & n15064 ;
  assign n15067 = ~n15065 & ~n15066 ;
  assign n15068 = n14853 & ~n15067 ;
  assign n15069 = ~n14853 & n15067 ;
  assign n15070 = ~n15068 & ~n15069 ;
  assign n15071 = ~n15042 & n15070 ;
  assign n15072 = ~n15041 & n15069 ;
  assign n15073 = ~n15071 & ~n15072 ;
  assign n15074 = n15031 & ~n15036 ;
  assign n15075 = ~n15037 & ~n15074 ;
  assign n15076 = ~n15021 & ~n15022 ;
  assign n15077 = n15027 & ~n15076 ;
  assign n15078 = ~n15027 & n15076 ;
  assign n15079 = ~n15077 & ~n15078 ;
  assign n15080 = ~\core_eu_em_mac_em_reg_mxopwe_DO_reg[13]/P0001  & ~n14967 ;
  assign n15081 = \core_eu_em_mac_em_reg_mxopwe_DO_reg[13]/P0001  & ~n14969 ;
  assign n15082 = ~n15080 & ~n15081 ;
  assign n15084 = \core_eu_em_mac_em_reg_mxopwe_DO_reg[15]/P0001  & ~n14951 ;
  assign n15083 = ~\core_eu_em_mac_em_reg_mxopwe_DO_reg[15]/P0001  & ~n14947 ;
  assign n15085 = ~\core_eu_em_mac_em_reg_mxopwe_DO_reg[14]/P0001  & n14958 ;
  assign n15086 = \core_eu_em_mac_em_reg_mxopwe_DO_reg[14]/P0001  & n14962 ;
  assign n15087 = ~n15085 & ~n15086 ;
  assign n15088 = ~n15083 & n15087 ;
  assign n15089 = ~n15084 & n15088 ;
  assign n15090 = ~n15082 & n15089 ;
  assign n15091 = n15082 & ~n15089 ;
  assign n15094 = ~\core_c_psq_MSTAT_reg_DO_reg[4]/NET0131  & ~n15023 ;
  assign n15092 = \core_c_dec_MACop_E_reg/P0001  & ~n7202 ;
  assign n15093 = \core_c_psq_MSTAT_reg_DO_reg[4]/NET0131  & ~n15092 ;
  assign n15095 = ~\core_eu_em_mac_em_dec_emcorepi_DO_reg[1]/P0001  & ~n15093 ;
  assign n15096 = ~n15094 & n15095 ;
  assign n15097 = ~n15091 & ~n15096 ;
  assign n15098 = ~n15090 & ~n15097 ;
  assign n15099 = n15079 & ~n15098 ;
  assign n15100 = ~n14933 & ~n15099 ;
  assign n15101 = ~n15013 & n15029 ;
  assign n15102 = ~n15030 & ~n15101 ;
  assign n15103 = n14992 & ~n15102 ;
  assign n15104 = ~n14992 & n15102 ;
  assign n15105 = ~n15103 & ~n15104 ;
  assign n15106 = ~n15100 & ~n15105 ;
  assign n15107 = ~n14991 & ~n15101 ;
  assign n15108 = n15105 & n15107 ;
  assign n15109 = ~n15106 & ~n15108 ;
  assign n15110 = n15075 & ~n15109 ;
  assign n15111 = ~n14853 & ~n15110 ;
  assign n15112 = ~n15009 & n15040 ;
  assign n15113 = ~n15041 & ~n15112 ;
  assign n15114 = n14853 & n15113 ;
  assign n15115 = ~n14853 & ~n15113 ;
  assign n15116 = ~n15114 & ~n15115 ;
  assign n15117 = ~n15111 & ~n15116 ;
  assign n15118 = ~n15112 & n15116 ;
  assign n15119 = ~n15117 & ~n15118 ;
  assign n15120 = n15073 & ~n15119 ;
  assign n15121 = ~n15073 & n15119 ;
  assign n15122 = ~n15120 & ~n15121 ;
  assign n15123 = n15100 & n15105 ;
  assign n15124 = ~n15106 & ~n15123 ;
  assign n15125 = ~\core_eu_em_mac_em_reg_mxopwe_DO_reg[15]/P0001  & n14925 ;
  assign n15126 = \core_eu_em_mac_em_reg_mxopwe_DO_reg[15]/P0001  & n14929 ;
  assign n15127 = ~n15125 & ~n15126 ;
  assign n15128 = n14920 & n15127 ;
  assign n15129 = ~n14906 & ~n15128 ;
  assign n15130 = ~n14990 & ~n15129 ;
  assign n15131 = ~n14906 & ~n14990 ;
  assign n15132 = ~n14932 & n15131 ;
  assign n15133 = n14932 & ~n15131 ;
  assign n15134 = ~n15132 & ~n15133 ;
  assign n15135 = n15130 & ~n15134 ;
  assign n15136 = ~n15090 & ~n15091 ;
  assign n15137 = n15096 & ~n15136 ;
  assign n15138 = ~n15096 & n15136 ;
  assign n15139 = ~n15137 & ~n15138 ;
  assign n15142 = ~\core_c_psq_MSTAT_reg_DO_reg[4]/NET0131  & ~n15092 ;
  assign n15140 = \core_c_dec_MACop_E_reg/P0001  & ~n9056 ;
  assign n15141 = \core_c_psq_MSTAT_reg_DO_reg[4]/NET0131  & ~n15140 ;
  assign n15143 = ~\core_eu_em_mac_em_dec_emcorepi_DO_reg[1]/P0001  & ~n15141 ;
  assign n15144 = ~n15142 & n15143 ;
  assign n15146 = \core_eu_em_mac_em_reg_mxopwe_DO_reg[14]/P0001  & ~n14951 ;
  assign n15145 = ~\core_eu_em_mac_em_reg_mxopwe_DO_reg[14]/P0001  & ~n14947 ;
  assign n15147 = ~\core_eu_em_mac_em_reg_mxopwe_DO_reg[13]/P0001  & n14958 ;
  assign n15148 = \core_eu_em_mac_em_reg_mxopwe_DO_reg[13]/P0001  & n14962 ;
  assign n15149 = ~n15147 & ~n15148 ;
  assign n15150 = ~n15145 & n15149 ;
  assign n15151 = ~n15146 & n15150 ;
  assign n15152 = n15144 & ~n15151 ;
  assign n15153 = ~n15144 & n15151 ;
  assign n15154 = ~\core_eu_em_mac_em_reg_mxopwe_DO_reg[12]/P0001  & n14967 ;
  assign n15155 = \core_eu_em_mac_em_reg_mxopwe_DO_reg[12]/P0001  & n14969 ;
  assign n15156 = ~n15154 & ~n15155 ;
  assign n15157 = ~n15153 & ~n15156 ;
  assign n15158 = ~n15152 & ~n15157 ;
  assign n15159 = n15139 & n15158 ;
  assign n15160 = ~n15135 & ~n15159 ;
  assign n15161 = ~n15079 & n15098 ;
  assign n15162 = ~n15099 & ~n15161 ;
  assign n15163 = n14992 & ~n15162 ;
  assign n15164 = ~n14992 & n15162 ;
  assign n15165 = ~n15163 & ~n15164 ;
  assign n15166 = ~n15160 & ~n15165 ;
  assign n15167 = ~n14991 & ~n15161 ;
  assign n15168 = n15165 & n15167 ;
  assign n15169 = ~n15166 & ~n15168 ;
  assign n15170 = n15124 & ~n15169 ;
  assign n15171 = ~n14853 & ~n15170 ;
  assign n15172 = ~n15075 & n15109 ;
  assign n15173 = ~n15110 & ~n15172 ;
  assign n15174 = n14853 & n15173 ;
  assign n15175 = ~n14853 & ~n15173 ;
  assign n15176 = ~n15174 & ~n15175 ;
  assign n15177 = ~n15171 & ~n15176 ;
  assign n15178 = ~n15172 & n15176 ;
  assign n15179 = ~n15177 & ~n15178 ;
  assign n15180 = n15111 & n15113 ;
  assign n15181 = ~n15117 & ~n15180 ;
  assign n15182 = n15179 & ~n15181 ;
  assign n15183 = ~n15179 & n15181 ;
  assign n15184 = n15160 & n15165 ;
  assign n15185 = ~n15166 & ~n15184 ;
  assign n15187 = \core_eu_em_mac_em_reg_mxopwe_DO_reg[15]/P0001  & ~n14918 ;
  assign n15186 = ~\core_eu_em_mac_em_reg_mxopwe_DO_reg[15]/P0001  & ~n14914 ;
  assign n15188 = ~\core_eu_em_mac_em_reg_mxopwe_DO_reg[14]/P0001  & n14925 ;
  assign n15189 = \core_eu_em_mac_em_reg_mxopwe_DO_reg[14]/P0001  & n14929 ;
  assign n15190 = ~n15188 & ~n15189 ;
  assign n15191 = ~n15186 & n15190 ;
  assign n15192 = ~n15187 & n15191 ;
  assign n15193 = ~n14906 & ~n15192 ;
  assign n15194 = ~n14990 & ~n15193 ;
  assign n15195 = ~n15128 & n15131 ;
  assign n15196 = n15128 & ~n15131 ;
  assign n15197 = ~n15195 & ~n15196 ;
  assign n15198 = n15194 & ~n15197 ;
  assign n15199 = ~\core_eu_em_mac_em_reg_mxopwe_DO_reg[11]/P0001  & ~n14967 ;
  assign n15200 = \core_eu_em_mac_em_reg_mxopwe_DO_reg[11]/P0001  & ~n14969 ;
  assign n15201 = ~n15199 & ~n15200 ;
  assign n15203 = \core_eu_em_mac_em_reg_mxopwe_DO_reg[13]/P0001  & ~n14951 ;
  assign n15202 = ~\core_eu_em_mac_em_reg_mxopwe_DO_reg[13]/P0001  & ~n14947 ;
  assign n15204 = ~\core_eu_em_mac_em_reg_mxopwe_DO_reg[12]/P0001  & n14958 ;
  assign n15205 = \core_eu_em_mac_em_reg_mxopwe_DO_reg[12]/P0001  & n14962 ;
  assign n15206 = ~n15204 & ~n15205 ;
  assign n15207 = ~n15202 & n15206 ;
  assign n15208 = ~n15203 & n15207 ;
  assign n15209 = n15201 & ~n15208 ;
  assign n15210 = ~n15201 & n15208 ;
  assign n15213 = ~\core_c_psq_MSTAT_reg_DO_reg[4]/NET0131  & ~n15140 ;
  assign n15211 = \core_c_dec_MACop_E_reg/P0001  & ~n8358 ;
  assign n15212 = \core_c_psq_MSTAT_reg_DO_reg[4]/NET0131  & ~n15211 ;
  assign n15214 = ~\core_eu_em_mac_em_dec_emcorepi_DO_reg[1]/P0001  & ~n15212 ;
  assign n15215 = ~n15213 & n15214 ;
  assign n15216 = ~n15210 & n15215 ;
  assign n15217 = ~n15209 & ~n15216 ;
  assign n15218 = ~n15152 & ~n15153 ;
  assign n15219 = ~n15156 & n15218 ;
  assign n15220 = n15156 & ~n15218 ;
  assign n15221 = ~n15219 & ~n15220 ;
  assign n15222 = n15217 & ~n15221 ;
  assign n15223 = ~n15198 & ~n15222 ;
  assign n15224 = ~n15130 & n15134 ;
  assign n15225 = ~n15135 & ~n15224 ;
  assign n15226 = ~n15139 & ~n15158 ;
  assign n15227 = ~n15159 & ~n15226 ;
  assign n15228 = n15225 & n15227 ;
  assign n15229 = ~n15225 & ~n15227 ;
  assign n15230 = ~n15228 & ~n15229 ;
  assign n15231 = ~n15223 & n15230 ;
  assign n15232 = ~n15224 & ~n15226 ;
  assign n15233 = ~n15230 & n15232 ;
  assign n15234 = ~n15231 & ~n15233 ;
  assign n15235 = n15185 & ~n15234 ;
  assign n15236 = ~n14853 & ~n15235 ;
  assign n15237 = ~n15124 & n15169 ;
  assign n15238 = ~n15170 & ~n15237 ;
  assign n15239 = n14853 & n15238 ;
  assign n15240 = ~n14853 & ~n15238 ;
  assign n15241 = ~n15239 & ~n15240 ;
  assign n15242 = ~n15236 & ~n15241 ;
  assign n15243 = n15236 & n15238 ;
  assign n15244 = ~n15242 & ~n15243 ;
  assign n15245 = n15171 & n15173 ;
  assign n15246 = ~n15177 & ~n15245 ;
  assign n15247 = ~n15244 & ~n15246 ;
  assign n15248 = n15223 & ~n15230 ;
  assign n15249 = ~n15231 & ~n15248 ;
  assign n15250 = ~n15209 & ~n15210 ;
  assign n15251 = n15215 & n15250 ;
  assign n15252 = ~n15215 & ~n15250 ;
  assign n15253 = ~n15251 & ~n15252 ;
  assign n15256 = ~\core_c_psq_MSTAT_reg_DO_reg[4]/NET0131  & ~n15211 ;
  assign n15254 = \core_c_dec_MACop_E_reg/P0001  & ~n7737 ;
  assign n15255 = \core_c_psq_MSTAT_reg_DO_reg[4]/NET0131  & ~n15254 ;
  assign n15257 = ~\core_eu_em_mac_em_dec_emcorepi_DO_reg[1]/P0001  & ~n15255 ;
  assign n15258 = ~n15256 & n15257 ;
  assign n15260 = \core_eu_em_mac_em_reg_mxopwe_DO_reg[12]/P0001  & ~n14951 ;
  assign n15259 = ~\core_eu_em_mac_em_reg_mxopwe_DO_reg[12]/P0001  & ~n14947 ;
  assign n15261 = ~\core_eu_em_mac_em_reg_mxopwe_DO_reg[11]/P0001  & n14958 ;
  assign n15262 = \core_eu_em_mac_em_reg_mxopwe_DO_reg[11]/P0001  & n14962 ;
  assign n15263 = ~n15261 & ~n15262 ;
  assign n15264 = ~n15259 & n15263 ;
  assign n15265 = ~n15260 & n15264 ;
  assign n15266 = n15258 & ~n15265 ;
  assign n15267 = ~n15258 & n15265 ;
  assign n15268 = ~\core_eu_em_mac_em_reg_mxopwe_DO_reg[10]/P0001  & n14967 ;
  assign n15269 = \core_eu_em_mac_em_reg_mxopwe_DO_reg[10]/P0001  & n14969 ;
  assign n15270 = ~n15268 & ~n15269 ;
  assign n15271 = ~n15267 & ~n15270 ;
  assign n15272 = ~n15266 & ~n15271 ;
  assign n15273 = ~n15253 & n15272 ;
  assign n15275 = \core_eu_em_mac_em_reg_mxopwe_DO_reg[14]/P0001  & ~n14918 ;
  assign n15274 = ~\core_eu_em_mac_em_reg_mxopwe_DO_reg[14]/P0001  & ~n14914 ;
  assign n15276 = ~\core_eu_em_mac_em_reg_mxopwe_DO_reg[13]/P0001  & n14925 ;
  assign n15277 = \core_eu_em_mac_em_reg_mxopwe_DO_reg[13]/P0001  & n14929 ;
  assign n15278 = ~n15276 & ~n15277 ;
  assign n15279 = ~n15274 & n15278 ;
  assign n15280 = ~n15275 & n15279 ;
  assign n15281 = n14879 & n15280 ;
  assign n15282 = ~\core_eu_em_mac_em_reg_mxopwe_DO_reg[15]/P0001  & n14898 ;
  assign n15283 = \core_eu_em_mac_em_reg_mxopwe_DO_reg[15]/P0001  & n14902 ;
  assign n15284 = ~n15282 & ~n15283 ;
  assign n15285 = n14893 & n15284 ;
  assign n15286 = ~n15281 & ~n15285 ;
  assign n15287 = ~n14879 & ~n15280 ;
  assign n15288 = ~n15286 & ~n15287 ;
  assign n15289 = n15131 & ~n15192 ;
  assign n15290 = ~n15131 & n15192 ;
  assign n15291 = ~n15289 & ~n15290 ;
  assign n15292 = n15288 & ~n15291 ;
  assign n15293 = ~n15273 & ~n15292 ;
  assign n15294 = ~n15194 & n15197 ;
  assign n15295 = ~n15198 & ~n15294 ;
  assign n15296 = ~n15217 & n15221 ;
  assign n15297 = ~n15222 & ~n15296 ;
  assign n15298 = n15295 & n15297 ;
  assign n15299 = ~n15295 & ~n15297 ;
  assign n15300 = ~n15298 & ~n15299 ;
  assign n15301 = ~n15293 & n15300 ;
  assign n15302 = ~n15294 & ~n15296 ;
  assign n15303 = ~n15300 & n15302 ;
  assign n15304 = ~n15301 & ~n15303 ;
  assign n15305 = n15249 & ~n15304 ;
  assign n15306 = ~n14853 & ~n15305 ;
  assign n15307 = ~n15185 & n15234 ;
  assign n15308 = ~n15235 & ~n15307 ;
  assign n15309 = n14853 & n15308 ;
  assign n15310 = ~n14853 & ~n15308 ;
  assign n15311 = ~n15309 & ~n15310 ;
  assign n15312 = ~n15306 & ~n15311 ;
  assign n15313 = ~n15307 & n15311 ;
  assign n15314 = ~n15312 & ~n15313 ;
  assign n15315 = ~n15237 & n15241 ;
  assign n15316 = ~n15242 & ~n15315 ;
  assign n15317 = n15246 & ~n15316 ;
  assign n15318 = n15314 & ~n15317 ;
  assign n15319 = ~n15247 & ~n15318 ;
  assign n16061 = \core_eu_em_mac_em_reg_mxopwe_DO_reg[1]/P0001  & ~n14791 ;
  assign n16060 = ~\core_eu_em_mac_em_reg_mxopwe_DO_reg[1]/P0001  & ~n14787 ;
  assign n16062 = ~\core_eu_em_mac_em_reg_mxopwe_DO_reg[0]/P0001  & n14798 ;
  assign n16063 = \core_eu_em_mac_em_reg_mxopwe_DO_reg[0]/P0001  & n14802 ;
  assign n16064 = ~n16062 & ~n16063 ;
  assign n16065 = ~n16060 & n16064 ;
  assign n16066 = ~n16061 & n16065 ;
  assign n16068 = \core_eu_em_mac_em_reg_mxopwe_DO_reg[3]/P0001  & ~n14765 ;
  assign n16067 = ~\core_eu_em_mac_em_reg_mxopwe_DO_reg[3]/P0001  & ~n14761 ;
  assign n16069 = ~\core_eu_em_mac_em_reg_mxopwe_DO_reg[2]/P0001  & n14772 ;
  assign n16070 = \core_eu_em_mac_em_reg_mxopwe_DO_reg[2]/P0001  & n14776 ;
  assign n16071 = ~n16069 & ~n16070 ;
  assign n16072 = ~n16067 & n16071 ;
  assign n16073 = ~n16068 & n16072 ;
  assign n16074 = ~n16066 & ~n16073 ;
  assign n15994 = \core_eu_em_mac_em_reg_mxopwe_DO_reg[2]/P0001  & ~n14791 ;
  assign n15993 = ~\core_eu_em_mac_em_reg_mxopwe_DO_reg[2]/P0001  & ~n14787 ;
  assign n15995 = ~\core_eu_em_mac_em_reg_mxopwe_DO_reg[1]/P0001  & n14798 ;
  assign n15996 = \core_eu_em_mac_em_reg_mxopwe_DO_reg[1]/P0001  & n14802 ;
  assign n15997 = ~n15995 & ~n15996 ;
  assign n15998 = ~n15993 & n15997 ;
  assign n15999 = ~n15994 & n15998 ;
  assign n15981 = ~\core_eu_em_mac_em_reg_mxopwe_DO_reg[0]/P0001  & ~n14814 ;
  assign n15982 = \core_eu_em_mac_em_reg_mxopwe_DO_reg[0]/P0001  & ~n14818 ;
  assign n15983 = ~n15981 & ~n15982 ;
  assign n15985 = \core_eu_em_mac_em_reg_mxopwe_DO_reg[4]/P0001  & ~n14765 ;
  assign n15984 = ~\core_eu_em_mac_em_reg_mxopwe_DO_reg[4]/P0001  & ~n14761 ;
  assign n15986 = ~\core_eu_em_mac_em_reg_mxopwe_DO_reg[3]/P0001  & n14772 ;
  assign n15987 = \core_eu_em_mac_em_reg_mxopwe_DO_reg[3]/P0001  & n14776 ;
  assign n15988 = ~n15986 & ~n15987 ;
  assign n15989 = ~n15984 & n15988 ;
  assign n15990 = ~n15985 & n15989 ;
  assign n15991 = ~n15983 & ~n15990 ;
  assign n15992 = n15983 & n15990 ;
  assign n16075 = ~n15991 & ~n15992 ;
  assign n16076 = n15999 & ~n16075 ;
  assign n16077 = ~n15999 & n16075 ;
  assign n16078 = ~n16076 & ~n16077 ;
  assign n16079 = ~n16074 & ~n16078 ;
  assign n16080 = ~n11444 & n14993 ;
  assign n16081 = ~n10878 & n15044 ;
  assign n16082 = ~n16080 & ~n16081 ;
  assign n16083 = ~\core_eu_em_mac_em_dec_emcorepi_DO_reg[1]/P0001  & ~n16082 ;
  assign n16085 = \core_eu_em_mac_em_reg_mxopwe_DO_reg[5]/P0001  & ~n14842 ;
  assign n16084 = ~\core_eu_em_mac_em_reg_mxopwe_DO_reg[5]/P0001  & ~n14838 ;
  assign n16086 = ~\core_eu_em_mac_em_reg_mxopwe_DO_reg[4]/P0001  & n14846 ;
  assign n16087 = \core_eu_em_mac_em_reg_mxopwe_DO_reg[4]/P0001  & n14849 ;
  assign n16088 = ~n16086 & ~n16087 ;
  assign n16089 = ~n16084 & n16088 ;
  assign n16090 = ~n16085 & n16089 ;
  assign n16091 = ~n16083 & n16090 ;
  assign n16092 = n16083 & ~n16090 ;
  assign n16093 = ~n14798 & ~n16092 ;
  assign n16094 = ~n16091 & ~n16093 ;
  assign n16018 = \core_eu_em_mac_em_reg_mxopwe_DO_reg[6]/P0001  & ~n14842 ;
  assign n16017 = ~\core_eu_em_mac_em_reg_mxopwe_DO_reg[6]/P0001  & ~n14838 ;
  assign n16019 = ~\core_eu_em_mac_em_reg_mxopwe_DO_reg[5]/P0001  & n14846 ;
  assign n16020 = \core_eu_em_mac_em_reg_mxopwe_DO_reg[5]/P0001  & n14849 ;
  assign n16021 = ~n16019 & ~n16020 ;
  assign n16022 = ~n16017 & n16021 ;
  assign n16023 = ~n16018 & n16022 ;
  assign n16011 = ~n11192 & n14993 ;
  assign n16012 = ~n11444 & n15044 ;
  assign n16013 = ~n16011 & ~n16012 ;
  assign n16014 = ~\core_eu_em_mac_em_dec_emcorepi_DO_reg[1]/P0001  & ~n16013 ;
  assign n16015 = ~n14814 & n16014 ;
  assign n16016 = n14814 & ~n16014 ;
  assign n16095 = ~n16015 & ~n16016 ;
  assign n16096 = n16023 & n16095 ;
  assign n16097 = ~n16023 & ~n16095 ;
  assign n16098 = ~n16096 & ~n16097 ;
  assign n16099 = ~n16094 & n16098 ;
  assign n16100 = ~n16079 & ~n16099 ;
  assign n16000 = ~n15992 & ~n15999 ;
  assign n16001 = ~n15991 & ~n16000 ;
  assign n15921 = \core_eu_em_mac_em_reg_mxopwe_DO_reg[1]/P0001  & ~n14818 ;
  assign n15920 = ~\core_eu_em_mac_em_reg_mxopwe_DO_reg[1]/P0001  & ~n14814 ;
  assign n15922 = ~\core_eu_em_mac_em_reg_mxopwe_DO_reg[0]/P0001  & n14825 ;
  assign n15923 = \core_eu_em_mac_em_reg_mxopwe_DO_reg[0]/P0001  & n14829 ;
  assign n15924 = ~n15922 & ~n15923 ;
  assign n15925 = ~n15920 & n15924 ;
  assign n15926 = ~n15921 & n15925 ;
  assign n15905 = \core_eu_em_mac_em_reg_mxopwe_DO_reg[5]/P0001  & ~n14765 ;
  assign n15904 = ~\core_eu_em_mac_em_reg_mxopwe_DO_reg[5]/P0001  & ~n14761 ;
  assign n15906 = ~\core_eu_em_mac_em_reg_mxopwe_DO_reg[4]/P0001  & n14772 ;
  assign n15907 = \core_eu_em_mac_em_reg_mxopwe_DO_reg[4]/P0001  & n14776 ;
  assign n15908 = ~n15906 & ~n15907 ;
  assign n15909 = ~n15904 & n15908 ;
  assign n15910 = ~n15905 & n15909 ;
  assign n15912 = \core_eu_em_mac_em_reg_mxopwe_DO_reg[3]/P0001  & ~n14791 ;
  assign n15911 = ~\core_eu_em_mac_em_reg_mxopwe_DO_reg[3]/P0001  & ~n14787 ;
  assign n15913 = ~\core_eu_em_mac_em_reg_mxopwe_DO_reg[2]/P0001  & n14798 ;
  assign n15914 = \core_eu_em_mac_em_reg_mxopwe_DO_reg[2]/P0001  & n14802 ;
  assign n15915 = ~n15913 & ~n15914 ;
  assign n15916 = ~n15911 & n15915 ;
  assign n15917 = ~n15912 & n15916 ;
  assign n15918 = ~n15910 & ~n15917 ;
  assign n15919 = n15910 & n15917 ;
  assign n16002 = ~n15918 & ~n15919 ;
  assign n16003 = n15926 & ~n16002 ;
  assign n16004 = ~n15926 & n16002 ;
  assign n16005 = ~n16003 & ~n16004 ;
  assign n16006 = n16001 & ~n16005 ;
  assign n16101 = ~n16001 & n16005 ;
  assign n16102 = ~n16006 & ~n16101 ;
  assign n15946 = ~n10534 & n14993 ;
  assign n15947 = ~n11192 & n15044 ;
  assign n15948 = ~n15946 & ~n15947 ;
  assign n15949 = ~\core_eu_em_mac_em_dec_emcorepi_DO_reg[1]/P0001  & ~n15948 ;
  assign n15939 = \core_eu_em_mac_em_reg_mxopwe_DO_reg[7]/P0001  & ~n14842 ;
  assign n15938 = ~\core_eu_em_mac_em_reg_mxopwe_DO_reg[7]/P0001  & ~n14838 ;
  assign n15940 = ~\core_eu_em_mac_em_reg_mxopwe_DO_reg[6]/P0001  & n14846 ;
  assign n15941 = \core_eu_em_mac_em_reg_mxopwe_DO_reg[6]/P0001  & n14849 ;
  assign n15942 = ~n15940 & ~n15941 ;
  assign n15943 = ~n15938 & n15942 ;
  assign n15944 = ~n15939 & n15943 ;
  assign n15945 = ~n14825 & n15944 ;
  assign n15950 = n14825 & ~n15944 ;
  assign n16007 = ~n15945 & ~n15950 ;
  assign n16008 = n15949 & n16007 ;
  assign n16009 = ~n15949 & ~n16007 ;
  assign n16010 = ~n16008 & ~n16009 ;
  assign n16024 = ~n16016 & ~n16023 ;
  assign n16025 = ~n16015 & ~n16024 ;
  assign n16026 = ~n16010 & n16025 ;
  assign n16103 = n16010 & ~n16025 ;
  assign n16104 = ~n16026 & ~n16103 ;
  assign n16105 = n16102 & ~n16104 ;
  assign n16106 = ~n16102 & n16104 ;
  assign n16107 = ~n16105 & ~n16106 ;
  assign n16108 = ~n16100 & ~n16107 ;
  assign n16109 = n16100 & n16107 ;
  assign n16110 = ~n16108 & ~n16109 ;
  assign n16111 = \core_eu_em_mac_em_reg_mxopwe_DO_reg[0]/P0001  & ~n14791 ;
  assign n16112 = ~\core_eu_em_mac_em_reg_mxopwe_DO_reg[0]/P0001  & ~n14787 ;
  assign n16113 = ~n16111 & ~n16112 ;
  assign n16115 = \core_eu_em_mac_em_reg_mxopwe_DO_reg[2]/P0001  & ~n14765 ;
  assign n16114 = ~\core_eu_em_mac_em_reg_mxopwe_DO_reg[2]/P0001  & ~n14761 ;
  assign n16116 = ~\core_eu_em_mac_em_reg_mxopwe_DO_reg[1]/P0001  & n14772 ;
  assign n16117 = \core_eu_em_mac_em_reg_mxopwe_DO_reg[1]/P0001  & n14776 ;
  assign n16118 = ~n16116 & ~n16117 ;
  assign n16119 = ~n16114 & n16118 ;
  assign n16120 = ~n16115 & n16119 ;
  assign n16121 = ~n16113 & ~n16120 ;
  assign n16122 = n16066 & n16073 ;
  assign n16123 = ~n16074 & ~n16122 ;
  assign n16124 = ~n16121 & ~n16123 ;
  assign n16125 = ~n10878 & n14993 ;
  assign n16126 = ~n9869 & n15044 ;
  assign n16127 = ~n16125 & ~n16126 ;
  assign n16128 = ~\core_eu_em_mac_em_dec_emcorepi_DO_reg[1]/P0001  & ~n16127 ;
  assign n16129 = ~n14787 & n16128 ;
  assign n16130 = n14787 & ~n16128 ;
  assign n16132 = \core_eu_em_mac_em_reg_mxopwe_DO_reg[4]/P0001  & ~n14842 ;
  assign n16131 = ~\core_eu_em_mac_em_reg_mxopwe_DO_reg[4]/P0001  & ~n14838 ;
  assign n16133 = ~\core_eu_em_mac_em_reg_mxopwe_DO_reg[3]/P0001  & n14846 ;
  assign n16134 = \core_eu_em_mac_em_reg_mxopwe_DO_reg[3]/P0001  & n14849 ;
  assign n16135 = ~n16133 & ~n16134 ;
  assign n16136 = ~n16131 & n16135 ;
  assign n16137 = ~n16132 & n16136 ;
  assign n16138 = ~n16130 & ~n16137 ;
  assign n16139 = ~n16129 & ~n16138 ;
  assign n16140 = ~n16091 & ~n16092 ;
  assign n16141 = n14798 & ~n16140 ;
  assign n16142 = ~n14798 & n16140 ;
  assign n16143 = ~n16141 & ~n16142 ;
  assign n16144 = n16139 & n16143 ;
  assign n16145 = ~n16124 & ~n16144 ;
  assign n16146 = n16074 & n16078 ;
  assign n16147 = ~n16079 & ~n16146 ;
  assign n16148 = n16094 & ~n16098 ;
  assign n16149 = ~n16099 & ~n16148 ;
  assign n16150 = n16147 & n16149 ;
  assign n16151 = ~n16147 & ~n16149 ;
  assign n16152 = ~n16150 & ~n16151 ;
  assign n16153 = ~n16145 & n16152 ;
  assign n16154 = ~n16146 & ~n16148 ;
  assign n16155 = ~n16152 & n16154 ;
  assign n16156 = ~n16153 & ~n16155 ;
  assign n16157 = ~n16110 & n16156 ;
  assign n16158 = n16110 & ~n16156 ;
  assign n16159 = ~n16157 & ~n16158 ;
  assign n16160 = n16145 & ~n16152 ;
  assign n16161 = ~n16153 & ~n16160 ;
  assign n16162 = ~n9869 & n14993 ;
  assign n16163 = ~n7909 & n15044 ;
  assign n16164 = ~n16162 & ~n16163 ;
  assign n16165 = ~\core_eu_em_mac_em_dec_emcorepi_DO_reg[1]/P0001  & ~n16164 ;
  assign n16167 = ~\core_eu_em_mac_em_reg_mxopwe_DO_reg[3]/P0001  & ~n14838 ;
  assign n16166 = \core_eu_em_mac_em_reg_mxopwe_DO_reg[3]/P0001  & ~n14842 ;
  assign n16168 = \core_eu_em_mac_em_reg_mxopwe_DO_reg[2]/P0001  & n14849 ;
  assign n16169 = ~\core_eu_em_mac_em_reg_mxopwe_DO_reg[2]/P0001  & n14846 ;
  assign n16170 = ~n16168 & ~n16169 ;
  assign n16171 = ~n16166 & n16170 ;
  assign n16172 = ~n16167 & n16171 ;
  assign n16173 = ~n16165 & n16172 ;
  assign n16174 = n16165 & ~n16172 ;
  assign n16175 = ~n14772 & ~n16174 ;
  assign n16176 = ~n16173 & ~n16175 ;
  assign n16177 = ~n16129 & ~n16130 ;
  assign n16178 = ~n16137 & n16177 ;
  assign n16179 = n16137 & ~n16177 ;
  assign n16180 = ~n16178 & ~n16179 ;
  assign n16181 = ~n16176 & ~n16180 ;
  assign n16182 = n16113 & n16120 ;
  assign n16183 = ~n16121 & ~n16182 ;
  assign n16184 = ~n16181 & n16183 ;
  assign n16185 = ~n16139 & ~n16143 ;
  assign n16186 = ~n16144 & ~n16185 ;
  assign n16187 = n16121 & n16123 ;
  assign n16188 = ~n16124 & ~n16187 ;
  assign n16189 = n16186 & n16188 ;
  assign n16190 = ~n16186 & ~n16188 ;
  assign n16191 = ~n16189 & ~n16190 ;
  assign n16192 = ~n16184 & n16191 ;
  assign n16193 = ~n16185 & ~n16187 ;
  assign n16194 = ~n16191 & n16193 ;
  assign n16195 = ~n16192 & ~n16194 ;
  assign n16196 = ~n16161 & n16195 ;
  assign n16197 = n16161 & ~n16195 ;
  assign n16198 = ~n7909 & n14993 ;
  assign n16199 = \core_c_dec_MACop_E_reg/P0001  & ~n8554 ;
  assign n16200 = \core_c_psq_MSTAT_reg_DO_reg[4]/NET0131  & n16199 ;
  assign n16201 = ~n16198 & ~n16200 ;
  assign n16202 = ~\core_eu_em_mac_em_dec_emcorepi_DO_reg[1]/P0001  & ~n16201 ;
  assign n16204 = \core_eu_em_mac_em_reg_mxopwe_DO_reg[2]/P0001  & ~n14842 ;
  assign n16203 = ~\core_eu_em_mac_em_reg_mxopwe_DO_reg[2]/P0001  & ~n14838 ;
  assign n16205 = ~\core_eu_em_mac_em_reg_mxopwe_DO_reg[1]/P0001  & n14846 ;
  assign n16206 = \core_eu_em_mac_em_reg_mxopwe_DO_reg[1]/P0001  & n14849 ;
  assign n16207 = ~n16205 & ~n16206 ;
  assign n16208 = ~n16203 & n16207 ;
  assign n16209 = ~n16204 & n16208 ;
  assign n16210 = ~n16202 & n16209 ;
  assign n16211 = n16202 & ~n16209 ;
  assign n16212 = n14761 & ~n16211 ;
  assign n16213 = ~n16210 & ~n16212 ;
  assign n16214 = ~n16173 & ~n16174 ;
  assign n16215 = n14772 & ~n16214 ;
  assign n16216 = ~n14772 & n16214 ;
  assign n16217 = ~n16215 & ~n16216 ;
  assign n16218 = ~n16213 & n16217 ;
  assign n16220 = \core_eu_em_mac_em_reg_mxopwe_DO_reg[1]/P0001  & ~n14765 ;
  assign n16219 = ~\core_eu_em_mac_em_reg_mxopwe_DO_reg[1]/P0001  & ~n14761 ;
  assign n16221 = ~\core_eu_em_mac_em_reg_mxopwe_DO_reg[0]/P0001  & n14772 ;
  assign n16222 = \core_eu_em_mac_em_reg_mxopwe_DO_reg[0]/P0001  & n14776 ;
  assign n16223 = ~n16221 & ~n16222 ;
  assign n16224 = ~n16219 & n16223 ;
  assign n16225 = ~n16220 & n16224 ;
  assign n16226 = ~n16218 & ~n16225 ;
  assign n16227 = n16176 & n16180 ;
  assign n16228 = ~n16181 & ~n16227 ;
  assign n16229 = n16183 & n16228 ;
  assign n16230 = ~n16183 & ~n16228 ;
  assign n16231 = ~n16229 & ~n16230 ;
  assign n16232 = ~n16226 & n16231 ;
  assign n16233 = ~n16227 & ~n16231 ;
  assign n16234 = ~n16232 & ~n16233 ;
  assign n16235 = n16184 & ~n16191 ;
  assign n16236 = ~n16192 & ~n16235 ;
  assign n16237 = n16234 & ~n16236 ;
  assign n16238 = ~n16234 & n16236 ;
  assign n16239 = ~n16237 & ~n16238 ;
  assign n16240 = n16226 & ~n16231 ;
  assign n16241 = ~n16232 & ~n16240 ;
  assign n16242 = ~n9225 & n15044 ;
  assign n16243 = ~\core_c_psq_MSTAT_reg_DO_reg[4]/NET0131  & n16199 ;
  assign n16244 = ~n16242 & ~n16243 ;
  assign n16245 = ~\core_eu_em_mac_em_dec_emcorepi_DO_reg[1]/P0001  & ~n16244 ;
  assign n16247 = \core_eu_em_mac_em_reg_mxopwe_DO_reg[1]/P0001  & ~n14842 ;
  assign n16246 = ~\core_eu_em_mac_em_reg_mxopwe_DO_reg[1]/P0001  & ~n14838 ;
  assign n16248 = ~\core_eu_em_mac_em_reg_mxopwe_DO_reg[0]/P0001  & n14846 ;
  assign n16249 = \core_eu_em_mac_em_reg_mxopwe_DO_reg[0]/P0001  & n14849 ;
  assign n16250 = ~n16248 & ~n16249 ;
  assign n16251 = ~n16246 & n16250 ;
  assign n16252 = ~n16247 & n16251 ;
  assign n16253 = n16245 & ~n16252 ;
  assign n16254 = ~n16245 & n16252 ;
  assign n16255 = n14846 & ~n16254 ;
  assign n16256 = ~n16253 & ~n16255 ;
  assign n16257 = ~n16210 & ~n16211 ;
  assign n16258 = n14761 & n16257 ;
  assign n16259 = ~n14761 & ~n16257 ;
  assign n16260 = ~n16258 & ~n16259 ;
  assign n16261 = n16256 & n16260 ;
  assign n16262 = \core_eu_em_mac_em_reg_mxopwe_DO_reg[0]/P0001  & ~n14765 ;
  assign n16263 = ~\core_eu_em_mac_em_reg_mxopwe_DO_reg[0]/P0001  & ~n14761 ;
  assign n16264 = ~n16262 & ~n16263 ;
  assign n16265 = ~n16261 & ~n16264 ;
  assign n16266 = n16213 & ~n16217 ;
  assign n16267 = ~n16218 & ~n16266 ;
  assign n16268 = n16225 & ~n16267 ;
  assign n16269 = ~n16225 & n16267 ;
  assign n16270 = ~n16268 & ~n16269 ;
  assign n16271 = ~n16265 & n16270 ;
  assign n16272 = ~n16266 & ~n16270 ;
  assign n16273 = ~n16271 & ~n16272 ;
  assign n16274 = ~n16241 & n16273 ;
  assign n16275 = n16241 & ~n16273 ;
  assign n16276 = ~n16274 & ~n16275 ;
  assign n16277 = ~n16253 & ~n16254 ;
  assign n16278 = n14846 & n16277 ;
  assign n16279 = ~n14846 & ~n16277 ;
  assign n16280 = ~n16278 & ~n16279 ;
  assign n16281 = \core_eu_em_mac_em_reg_mxopwe_DO_reg[0]/P0001  & n14842 ;
  assign n16282 = ~n14838 & ~n16281 ;
  assign n16283 = ~n7469 & n15044 ;
  assign n16284 = ~n9225 & n14993 ;
  assign n16285 = ~n16283 & ~n16284 ;
  assign n16286 = ~\core_eu_em_mac_em_dec_emcorepi_DO_reg[1]/P0001  & ~n16285 ;
  assign n16287 = \core_eu_em_mac_em_reg_mxopwe_DO_reg[0]/P0001  & ~n14842 ;
  assign n16288 = n14838 & ~n16287 ;
  assign n16289 = n16286 & ~n16288 ;
  assign n16290 = ~n16282 & ~n16289 ;
  assign n16291 = n16280 & ~n16290 ;
  assign n16292 = ~n16256 & ~n16260 ;
  assign n16293 = ~n16261 & ~n16292 ;
  assign n16294 = ~n16264 & n16293 ;
  assign n16295 = n16264 & ~n16293 ;
  assign n16296 = ~n16294 & ~n16295 ;
  assign n16297 = n16291 & n16296 ;
  assign n16299 = n16265 & ~n16270 ;
  assign n16298 = n16264 & n16292 ;
  assign n16300 = ~n16271 & ~n16298 ;
  assign n16301 = ~n16299 & n16300 ;
  assign n16302 = n16297 & ~n16301 ;
  assign n16303 = n16270 & n16298 ;
  assign n16304 = ~n16302 & ~n16303 ;
  assign n16305 = n16276 & ~n16304 ;
  assign n16306 = ~n16274 & ~n16305 ;
  assign n16307 = n16239 & ~n16306 ;
  assign n16308 = ~n16237 & ~n16307 ;
  assign n16309 = ~n16197 & ~n16308 ;
  assign n16310 = ~n16196 & ~n16309 ;
  assign n16311 = n16159 & ~n16310 ;
  assign n16312 = ~n16157 & ~n16311 ;
  assign n16027 = ~n16006 & ~n16026 ;
  assign n15927 = ~n15919 & ~n15926 ;
  assign n15928 = ~n15918 & ~n15927 ;
  assign n15717 = \core_eu_em_mac_em_reg_mxopwe_DO_reg[2]/P0001  & ~n14818 ;
  assign n15716 = ~\core_eu_em_mac_em_reg_mxopwe_DO_reg[2]/P0001  & ~n14814 ;
  assign n15718 = ~\core_eu_em_mac_em_reg_mxopwe_DO_reg[1]/P0001  & n14825 ;
  assign n15719 = \core_eu_em_mac_em_reg_mxopwe_DO_reg[1]/P0001  & n14829 ;
  assign n15720 = ~n15718 & ~n15719 ;
  assign n15721 = ~n15716 & n15720 ;
  assign n15722 = ~n15717 & n15721 ;
  assign n15701 = \core_eu_em_mac_em_reg_mxopwe_DO_reg[6]/P0001  & ~n14765 ;
  assign n15700 = ~\core_eu_em_mac_em_reg_mxopwe_DO_reg[6]/P0001  & ~n14761 ;
  assign n15702 = ~\core_eu_em_mac_em_reg_mxopwe_DO_reg[5]/P0001  & n14772 ;
  assign n15703 = \core_eu_em_mac_em_reg_mxopwe_DO_reg[5]/P0001  & n14776 ;
  assign n15704 = ~n15702 & ~n15703 ;
  assign n15705 = ~n15700 & n15704 ;
  assign n15706 = ~n15701 & n15705 ;
  assign n15708 = \core_eu_em_mac_em_reg_mxopwe_DO_reg[4]/P0001  & ~n14791 ;
  assign n15707 = ~\core_eu_em_mac_em_reg_mxopwe_DO_reg[4]/P0001  & ~n14787 ;
  assign n15709 = ~\core_eu_em_mac_em_reg_mxopwe_DO_reg[3]/P0001  & n14798 ;
  assign n15710 = \core_eu_em_mac_em_reg_mxopwe_DO_reg[3]/P0001  & n14802 ;
  assign n15711 = ~n15709 & ~n15710 ;
  assign n15712 = ~n15707 & n15711 ;
  assign n15713 = ~n15708 & n15712 ;
  assign n15714 = ~n15706 & ~n15713 ;
  assign n15715 = n15706 & n15713 ;
  assign n15929 = ~n15714 & ~n15715 ;
  assign n15930 = n15722 & ~n15929 ;
  assign n15931 = ~n15722 & n15929 ;
  assign n15932 = ~n15930 & ~n15931 ;
  assign n15933 = n15928 & ~n15932 ;
  assign n16028 = ~n15928 & n15932 ;
  assign n16029 = ~n15933 & ~n16028 ;
  assign n15730 = ~n10112 & n14993 ;
  assign n15731 = ~n10534 & n15044 ;
  assign n15732 = ~n15730 & ~n15731 ;
  assign n15733 = ~\core_eu_em_mac_em_dec_emcorepi_DO_reg[1]/P0001  & ~n15732 ;
  assign n15735 = \core_eu_em_mac_em_reg_mxopwe_DO_reg[8]/P0001  & ~n14842 ;
  assign n15734 = ~\core_eu_em_mac_em_reg_mxopwe_DO_reg[8]/P0001  & ~n14838 ;
  assign n15736 = ~\core_eu_em_mac_em_reg_mxopwe_DO_reg[7]/P0001  & n14846 ;
  assign n15737 = \core_eu_em_mac_em_reg_mxopwe_DO_reg[7]/P0001  & n14849 ;
  assign n15738 = ~n15736 & ~n15737 ;
  assign n15739 = ~n15734 & n15738 ;
  assign n15740 = ~n15735 & n15739 ;
  assign n15741 = ~n15733 & n15740 ;
  assign n15742 = n15733 & ~n15740 ;
  assign n15934 = ~n15741 & ~n15742 ;
  assign n15935 = n14861 & ~n15934 ;
  assign n15936 = ~n14861 & n15934 ;
  assign n15937 = ~n15935 & ~n15936 ;
  assign n15951 = ~n15949 & ~n15950 ;
  assign n15952 = ~n15945 & ~n15951 ;
  assign n15953 = ~n15937 & ~n15952 ;
  assign n16030 = n15937 & n15952 ;
  assign n16031 = ~n15953 & ~n16030 ;
  assign n16032 = n16029 & n16031 ;
  assign n16033 = ~n16029 & ~n16031 ;
  assign n16034 = ~n16032 & ~n16033 ;
  assign n16035 = ~n16027 & n16034 ;
  assign n16313 = n16027 & ~n16034 ;
  assign n16314 = ~n16035 & ~n16313 ;
  assign n16315 = ~n16101 & ~n16103 ;
  assign n16316 = n16107 & n16315 ;
  assign n16317 = ~n16108 & ~n16316 ;
  assign n16318 = n16314 & ~n16317 ;
  assign n16319 = ~n16314 & n16317 ;
  assign n16320 = ~n16318 & ~n16319 ;
  assign n16321 = \core_eu_em_mac_em_reg_mxopwe_DO_reg[0]/P0001  & ~n14865 ;
  assign n16322 = ~\core_eu_em_mac_em_reg_mxopwe_DO_reg[0]/P0001  & ~n14861 ;
  assign n16323 = ~n16321 & ~n16322 ;
  assign n16324 = ~n16320 & n16323 ;
  assign n16325 = n16320 & ~n16323 ;
  assign n16326 = ~n16324 & ~n16325 ;
  assign n16327 = ~n16312 & n16326 ;
  assign n16328 = ~n16318 & ~n16323 ;
  assign n16041 = \core_eu_em_mac_em_reg_mxopwe_DO_reg[1]/P0001  & ~n14865 ;
  assign n16040 = ~\core_eu_em_mac_em_reg_mxopwe_DO_reg[1]/P0001  & ~n14861 ;
  assign n16042 = ~\core_eu_em_mac_em_reg_mxopwe_DO_reg[0]/P0001  & n14872 ;
  assign n16043 = \core_eu_em_mac_em_reg_mxopwe_DO_reg[0]/P0001  & n14876 ;
  assign n16044 = ~n16042 & ~n16043 ;
  assign n16045 = ~n16040 & n16044 ;
  assign n16046 = ~n16041 & n16045 ;
  assign n15954 = ~n15933 & ~n15953 ;
  assign n15723 = ~n15715 & ~n15722 ;
  assign n15724 = ~n15714 & ~n15723 ;
  assign n15485 = \core_eu_em_mac_em_reg_mxopwe_DO_reg[3]/P0001  & ~n14818 ;
  assign n15484 = ~\core_eu_em_mac_em_reg_mxopwe_DO_reg[3]/P0001  & ~n14814 ;
  assign n15486 = ~\core_eu_em_mac_em_reg_mxopwe_DO_reg[2]/P0001  & n14825 ;
  assign n15487 = \core_eu_em_mac_em_reg_mxopwe_DO_reg[2]/P0001  & n14829 ;
  assign n15488 = ~n15486 & ~n15487 ;
  assign n15489 = ~n15484 & n15488 ;
  assign n15490 = ~n15485 & n15489 ;
  assign n15469 = \core_eu_em_mac_em_reg_mxopwe_DO_reg[5]/P0001  & ~n14791 ;
  assign n15468 = ~\core_eu_em_mac_em_reg_mxopwe_DO_reg[5]/P0001  & ~n14787 ;
  assign n15470 = ~\core_eu_em_mac_em_reg_mxopwe_DO_reg[4]/P0001  & n14798 ;
  assign n15471 = \core_eu_em_mac_em_reg_mxopwe_DO_reg[4]/P0001  & n14802 ;
  assign n15472 = ~n15470 & ~n15471 ;
  assign n15473 = ~n15468 & n15472 ;
  assign n15474 = ~n15469 & n15473 ;
  assign n15476 = \core_eu_em_mac_em_reg_mxopwe_DO_reg[7]/P0001  & ~n14765 ;
  assign n15475 = ~\core_eu_em_mac_em_reg_mxopwe_DO_reg[7]/P0001  & ~n14761 ;
  assign n15477 = ~\core_eu_em_mac_em_reg_mxopwe_DO_reg[6]/P0001  & n14772 ;
  assign n15478 = \core_eu_em_mac_em_reg_mxopwe_DO_reg[6]/P0001  & n14776 ;
  assign n15479 = ~n15477 & ~n15478 ;
  assign n15480 = ~n15475 & n15479 ;
  assign n15481 = ~n15476 & n15480 ;
  assign n15482 = ~n15474 & ~n15481 ;
  assign n15483 = n15474 & n15481 ;
  assign n15725 = ~n15482 & ~n15483 ;
  assign n15726 = n15490 & ~n15725 ;
  assign n15727 = ~n15490 & n15725 ;
  assign n15728 = ~n15726 & ~n15727 ;
  assign n15729 = n15724 & ~n15728 ;
  assign n15955 = ~n15724 & n15728 ;
  assign n15956 = ~n15729 & ~n15955 ;
  assign n15743 = n14861 & ~n15742 ;
  assign n15744 = ~n15741 & ~n15743 ;
  assign n15498 = ~n10112 & n15044 ;
  assign n15321 = \core_c_dec_MACop_E_reg/P0001  & ~n7753 ;
  assign n15499 = ~\core_c_psq_MSTAT_reg_DO_reg[4]/NET0131  & n15321 ;
  assign n15500 = ~n15498 & ~n15499 ;
  assign n15501 = ~\core_eu_em_mac_em_dec_emcorepi_DO_reg[1]/P0001  & ~n15500 ;
  assign n15503 = \core_eu_em_mac_em_reg_mxopwe_DO_reg[9]/P0001  & ~n14842 ;
  assign n15502 = ~\core_eu_em_mac_em_reg_mxopwe_DO_reg[9]/P0001  & ~n14838 ;
  assign n15504 = ~\core_eu_em_mac_em_reg_mxopwe_DO_reg[8]/P0001  & n14846 ;
  assign n15505 = \core_eu_em_mac_em_reg_mxopwe_DO_reg[8]/P0001  & n14849 ;
  assign n15506 = ~n15504 & ~n15505 ;
  assign n15507 = ~n15502 & n15506 ;
  assign n15508 = ~n15503 & n15507 ;
  assign n15509 = ~n15501 & n15508 ;
  assign n15510 = n15501 & ~n15508 ;
  assign n15745 = ~n15509 & ~n15510 ;
  assign n15746 = n14872 & n15745 ;
  assign n15747 = ~n14872 & ~n15745 ;
  assign n15748 = ~n15746 & ~n15747 ;
  assign n15749 = ~n15744 & ~n15748 ;
  assign n15957 = n15744 & n15748 ;
  assign n15958 = ~n15749 & ~n15957 ;
  assign n15959 = n15956 & n15958 ;
  assign n15960 = ~n15956 & ~n15958 ;
  assign n15961 = ~n15959 & ~n15960 ;
  assign n15962 = ~n15954 & n15961 ;
  assign n15979 = n15954 & ~n15961 ;
  assign n15980 = ~n15962 & ~n15979 ;
  assign n16036 = ~n16028 & ~n16030 ;
  assign n16037 = ~n16034 & n16036 ;
  assign n16038 = ~n16035 & ~n16037 ;
  assign n16039 = n15980 & ~n16038 ;
  assign n16329 = ~n15980 & n16038 ;
  assign n16330 = ~n16039 & ~n16329 ;
  assign n16331 = n16046 & ~n16330 ;
  assign n16332 = ~n16046 & n16330 ;
  assign n16333 = ~n16331 & ~n16332 ;
  assign n16334 = ~n16328 & n16333 ;
  assign n16335 = ~n16329 & ~n16333 ;
  assign n16336 = ~n16334 & ~n16335 ;
  assign n16047 = ~n16039 & ~n16046 ;
  assign n15531 = \core_eu_em_mac_em_reg_mxopwe_DO_reg[0]/P0001  & ~n14891 ;
  assign n15532 = ~\core_eu_em_mac_em_reg_mxopwe_DO_reg[0]/P0001  & ~n14887 ;
  assign n15533 = ~n15531 & ~n15532 ;
  assign n15535 = \core_eu_em_mac_em_reg_mxopwe_DO_reg[2]/P0001  & ~n14865 ;
  assign n15534 = ~\core_eu_em_mac_em_reg_mxopwe_DO_reg[2]/P0001  & ~n14861 ;
  assign n15536 = ~\core_eu_em_mac_em_reg_mxopwe_DO_reg[1]/P0001  & n14872 ;
  assign n15537 = \core_eu_em_mac_em_reg_mxopwe_DO_reg[1]/P0001  & n14876 ;
  assign n15538 = ~n15536 & ~n15537 ;
  assign n15539 = ~n15534 & n15538 ;
  assign n15540 = ~n15535 & n15539 ;
  assign n15541 = ~n15533 & ~n15540 ;
  assign n15900 = n15533 & n15540 ;
  assign n15901 = ~n15541 & ~n15900 ;
  assign n15750 = ~n15729 & ~n15749 ;
  assign n15491 = ~n15483 & ~n15490 ;
  assign n15492 = ~n15482 & ~n15491 ;
  assign n15371 = \core_eu_em_mac_em_reg_mxopwe_DO_reg[4]/P0001  & ~n14818 ;
  assign n15370 = ~\core_eu_em_mac_em_reg_mxopwe_DO_reg[4]/P0001  & ~n14814 ;
  assign n15372 = ~\core_eu_em_mac_em_reg_mxopwe_DO_reg[3]/P0001  & n14825 ;
  assign n15373 = \core_eu_em_mac_em_reg_mxopwe_DO_reg[3]/P0001  & n14829 ;
  assign n15374 = ~n15372 & ~n15373 ;
  assign n15375 = ~n15370 & n15374 ;
  assign n15376 = ~n15371 & n15375 ;
  assign n15355 = \core_eu_em_mac_em_reg_mxopwe_DO_reg[6]/P0001  & ~n14791 ;
  assign n15354 = ~\core_eu_em_mac_em_reg_mxopwe_DO_reg[6]/P0001  & ~n14787 ;
  assign n15356 = ~\core_eu_em_mac_em_reg_mxopwe_DO_reg[5]/P0001  & n14798 ;
  assign n15357 = \core_eu_em_mac_em_reg_mxopwe_DO_reg[5]/P0001  & n14802 ;
  assign n15358 = ~n15356 & ~n15357 ;
  assign n15359 = ~n15354 & n15358 ;
  assign n15360 = ~n15355 & n15359 ;
  assign n15362 = \core_eu_em_mac_em_reg_mxopwe_DO_reg[8]/P0001  & ~n14765 ;
  assign n15361 = ~\core_eu_em_mac_em_reg_mxopwe_DO_reg[8]/P0001  & ~n14761 ;
  assign n15363 = ~\core_eu_em_mac_em_reg_mxopwe_DO_reg[7]/P0001  & n14772 ;
  assign n15364 = \core_eu_em_mac_em_reg_mxopwe_DO_reg[7]/P0001  & n14776 ;
  assign n15365 = ~n15363 & ~n15364 ;
  assign n15366 = ~n15361 & n15365 ;
  assign n15367 = ~n15362 & n15366 ;
  assign n15368 = ~n15360 & ~n15367 ;
  assign n15369 = n15360 & n15367 ;
  assign n15493 = ~n15368 & ~n15369 ;
  assign n15494 = n15376 & ~n15493 ;
  assign n15495 = ~n15376 & n15493 ;
  assign n15496 = ~n15494 & ~n15495 ;
  assign n15497 = n15492 & ~n15496 ;
  assign n15751 = ~n15492 & n15496 ;
  assign n15752 = ~n15497 & ~n15751 ;
  assign n15511 = ~n14872 & ~n15510 ;
  assign n15512 = ~n15509 & ~n15511 ;
  assign n15320 = ~n8354 & n14993 ;
  assign n15322 = \core_c_psq_MSTAT_reg_DO_reg[4]/NET0131  & n15321 ;
  assign n15323 = ~n15320 & ~n15322 ;
  assign n15324 = ~\core_eu_em_mac_em_dec_emcorepi_DO_reg[1]/P0001  & ~n15323 ;
  assign n15326 = \core_eu_em_mac_em_reg_mxopwe_DO_reg[10]/P0001  & ~n14842 ;
  assign n15325 = ~\core_eu_em_mac_em_reg_mxopwe_DO_reg[10]/P0001  & ~n14838 ;
  assign n15327 = ~\core_eu_em_mac_em_reg_mxopwe_DO_reg[9]/P0001  & n14846 ;
  assign n15328 = \core_eu_em_mac_em_reg_mxopwe_DO_reg[9]/P0001  & n14849 ;
  assign n15329 = ~n15327 & ~n15328 ;
  assign n15330 = ~n15325 & n15329 ;
  assign n15331 = ~n15326 & n15330 ;
  assign n15332 = ~n15324 & n15331 ;
  assign n15333 = n15324 & ~n15331 ;
  assign n15513 = ~n15332 & ~n15333 ;
  assign n15514 = n14887 & ~n15513 ;
  assign n15515 = ~n14887 & n15513 ;
  assign n15516 = ~n15514 & ~n15515 ;
  assign n15517 = ~n15512 & ~n15516 ;
  assign n15753 = n15512 & n15516 ;
  assign n15754 = ~n15517 & ~n15753 ;
  assign n15755 = n15752 & n15754 ;
  assign n15756 = ~n15752 & ~n15754 ;
  assign n15757 = ~n15755 & ~n15756 ;
  assign n15758 = ~n15750 & n15757 ;
  assign n15902 = n15750 & ~n15757 ;
  assign n15903 = ~n15758 & ~n15902 ;
  assign n15963 = ~n15955 & ~n15957 ;
  assign n15964 = ~n15961 & n15963 ;
  assign n15965 = ~n15962 & ~n15964 ;
  assign n15966 = n15903 & ~n15965 ;
  assign n16048 = ~n15903 & n15965 ;
  assign n16049 = ~n15966 & ~n16048 ;
  assign n16050 = ~n15901 & ~n16049 ;
  assign n16051 = n15901 & n16049 ;
  assign n16052 = ~n16050 & ~n16051 ;
  assign n16053 = ~n16047 & n16052 ;
  assign n16337 = n16047 & ~n16052 ;
  assign n16338 = ~n16053 & ~n16337 ;
  assign n16339 = ~n16336 & n16338 ;
  assign n16341 = n16328 & ~n16333 ;
  assign n16340 = n16319 & n16323 ;
  assign n16342 = ~n16334 & ~n16340 ;
  assign n16343 = ~n16341 & n16342 ;
  assign n16344 = ~n16339 & ~n16343 ;
  assign n16345 = n16327 & n16344 ;
  assign n16346 = n16336 & ~n16338 ;
  assign n16347 = n16333 & n16340 ;
  assign n16348 = ~n16339 & n16347 ;
  assign n16349 = ~n16346 & ~n16348 ;
  assign n16350 = ~n16345 & n16349 ;
  assign n15334 = n14887 & ~n15333 ;
  assign n15335 = ~n15332 & ~n15334 ;
  assign n15336 = ~n9072 & n14993 ;
  assign n15337 = ~n8354 & n15044 ;
  assign n15338 = ~n15336 & ~n15337 ;
  assign n15339 = ~\core_eu_em_mac_em_dec_emcorepi_DO_reg[1]/P0001  & ~n15338 ;
  assign n15341 = \core_eu_em_mac_em_reg_mxopwe_DO_reg[11]/P0001  & ~n14842 ;
  assign n15340 = ~\core_eu_em_mac_em_reg_mxopwe_DO_reg[11]/P0001  & ~n14838 ;
  assign n15342 = ~\core_eu_em_mac_em_reg_mxopwe_DO_reg[10]/P0001  & n14846 ;
  assign n15343 = \core_eu_em_mac_em_reg_mxopwe_DO_reg[10]/P0001  & n14849 ;
  assign n15344 = ~n15342 & ~n15343 ;
  assign n15345 = ~n15340 & n15344 ;
  assign n15346 = ~n15341 & n15345 ;
  assign n15347 = n15339 & ~n15346 ;
  assign n15348 = ~n15339 & n15346 ;
  assign n15349 = ~n15347 & ~n15348 ;
  assign n15350 = n14898 & n15349 ;
  assign n15351 = ~n14898 & ~n15349 ;
  assign n15352 = ~n15350 & ~n15351 ;
  assign n15353 = ~n15335 & ~n15352 ;
  assign n15377 = ~n15369 & ~n15376 ;
  assign n15378 = ~n15368 & ~n15377 ;
  assign n15380 = \core_eu_em_mac_em_reg_mxopwe_DO_reg[7]/P0001  & ~n14791 ;
  assign n15379 = ~\core_eu_em_mac_em_reg_mxopwe_DO_reg[7]/P0001  & ~n14787 ;
  assign n15381 = ~\core_eu_em_mac_em_reg_mxopwe_DO_reg[6]/P0001  & n14798 ;
  assign n15382 = \core_eu_em_mac_em_reg_mxopwe_DO_reg[6]/P0001  & n14802 ;
  assign n15383 = ~n15381 & ~n15382 ;
  assign n15384 = ~n15379 & n15383 ;
  assign n15385 = ~n15380 & n15384 ;
  assign n15387 = \core_eu_em_mac_em_reg_mxopwe_DO_reg[9]/P0001  & ~n14765 ;
  assign n15386 = ~\core_eu_em_mac_em_reg_mxopwe_DO_reg[9]/P0001  & ~n14761 ;
  assign n15388 = ~\core_eu_em_mac_em_reg_mxopwe_DO_reg[8]/P0001  & n14772 ;
  assign n15389 = \core_eu_em_mac_em_reg_mxopwe_DO_reg[8]/P0001  & n14776 ;
  assign n15390 = ~n15388 & ~n15389 ;
  assign n15391 = ~n15386 & n15390 ;
  assign n15392 = ~n15387 & n15391 ;
  assign n15393 = n15385 & n15392 ;
  assign n15394 = ~n15385 & ~n15392 ;
  assign n15395 = ~n15393 & ~n15394 ;
  assign n15397 = \core_eu_em_mac_em_reg_mxopwe_DO_reg[5]/P0001  & ~n14818 ;
  assign n15396 = ~\core_eu_em_mac_em_reg_mxopwe_DO_reg[5]/P0001  & ~n14814 ;
  assign n15398 = ~\core_eu_em_mac_em_reg_mxopwe_DO_reg[4]/P0001  & n14825 ;
  assign n15399 = \core_eu_em_mac_em_reg_mxopwe_DO_reg[4]/P0001  & n14829 ;
  assign n15400 = ~n15398 & ~n15399 ;
  assign n15401 = ~n15396 & n15400 ;
  assign n15402 = ~n15397 & n15401 ;
  assign n15403 = ~n15395 & n15402 ;
  assign n15404 = n15395 & ~n15402 ;
  assign n15405 = ~n15403 & ~n15404 ;
  assign n15406 = n15378 & ~n15405 ;
  assign n15407 = ~n15353 & ~n15406 ;
  assign n15408 = ~n15393 & ~n15402 ;
  assign n15409 = ~n15394 & ~n15408 ;
  assign n15411 = \core_eu_em_mac_em_reg_mxopwe_DO_reg[10]/P0001  & ~n14765 ;
  assign n15410 = ~\core_eu_em_mac_em_reg_mxopwe_DO_reg[10]/P0001  & ~n14761 ;
  assign n15412 = ~\core_eu_em_mac_em_reg_mxopwe_DO_reg[9]/P0001  & n14772 ;
  assign n15413 = \core_eu_em_mac_em_reg_mxopwe_DO_reg[9]/P0001  & n14776 ;
  assign n15414 = ~n15412 & ~n15413 ;
  assign n15415 = ~n15410 & n15414 ;
  assign n15416 = ~n15411 & n15415 ;
  assign n15418 = \core_eu_em_mac_em_reg_mxopwe_DO_reg[8]/P0001  & ~n14791 ;
  assign n15417 = ~\core_eu_em_mac_em_reg_mxopwe_DO_reg[8]/P0001  & ~n14787 ;
  assign n15419 = ~\core_eu_em_mac_em_reg_mxopwe_DO_reg[7]/P0001  & n14798 ;
  assign n15420 = \core_eu_em_mac_em_reg_mxopwe_DO_reg[7]/P0001  & n14802 ;
  assign n15421 = ~n15419 & ~n15420 ;
  assign n15422 = ~n15417 & n15421 ;
  assign n15423 = ~n15418 & n15422 ;
  assign n15424 = n15416 & n15423 ;
  assign n15425 = ~n15416 & ~n15423 ;
  assign n15426 = ~n15424 & ~n15425 ;
  assign n15428 = \core_eu_em_mac_em_reg_mxopwe_DO_reg[6]/P0001  & ~n14818 ;
  assign n15427 = ~\core_eu_em_mac_em_reg_mxopwe_DO_reg[6]/P0001  & ~n14814 ;
  assign n15429 = ~\core_eu_em_mac_em_reg_mxopwe_DO_reg[5]/P0001  & n14825 ;
  assign n15430 = \core_eu_em_mac_em_reg_mxopwe_DO_reg[5]/P0001  & n14829 ;
  assign n15431 = ~n15429 & ~n15430 ;
  assign n15432 = ~n15427 & n15431 ;
  assign n15433 = ~n15428 & n15432 ;
  assign n15434 = ~n15426 & n15433 ;
  assign n15435 = n15426 & ~n15433 ;
  assign n15436 = ~n15434 & ~n15435 ;
  assign n15437 = n15409 & ~n15436 ;
  assign n15438 = ~n15409 & n15436 ;
  assign n15439 = ~n15437 & ~n15438 ;
  assign n15440 = ~n14898 & ~n15347 ;
  assign n15441 = ~n15348 & ~n15440 ;
  assign n15442 = ~n7182 & n14993 ;
  assign n15443 = ~n9072 & n15044 ;
  assign n15444 = ~n15442 & ~n15443 ;
  assign n15445 = ~\core_eu_em_mac_em_dec_emcorepi_DO_reg[1]/P0001  & ~n15444 ;
  assign n15447 = \core_eu_em_mac_em_reg_mxopwe_DO_reg[12]/P0001  & ~n14842 ;
  assign n15446 = ~\core_eu_em_mac_em_reg_mxopwe_DO_reg[12]/P0001  & ~n14838 ;
  assign n15448 = ~\core_eu_em_mac_em_reg_mxopwe_DO_reg[11]/P0001  & n14846 ;
  assign n15449 = \core_eu_em_mac_em_reg_mxopwe_DO_reg[11]/P0001  & n14849 ;
  assign n15450 = ~n15448 & ~n15449 ;
  assign n15451 = ~n15446 & n15450 ;
  assign n15452 = ~n15447 & n15451 ;
  assign n15453 = n15445 & ~n15452 ;
  assign n15454 = ~n15445 & n15452 ;
  assign n15455 = ~n15453 & ~n15454 ;
  assign n15456 = n14914 & ~n15455 ;
  assign n15457 = ~n14914 & n15455 ;
  assign n15458 = ~n15456 & ~n15457 ;
  assign n15459 = ~n15441 & ~n15458 ;
  assign n15460 = n15441 & n15458 ;
  assign n15461 = ~n15459 & ~n15460 ;
  assign n15462 = n15439 & n15461 ;
  assign n15463 = ~n15439 & ~n15461 ;
  assign n15464 = ~n15462 & ~n15463 ;
  assign n15465 = ~n15407 & n15464 ;
  assign n15466 = n15407 & ~n15464 ;
  assign n15467 = ~n15465 & ~n15466 ;
  assign n15518 = ~n15497 & ~n15517 ;
  assign n15519 = ~n15378 & n15405 ;
  assign n15520 = ~n15406 & ~n15519 ;
  assign n15521 = n15335 & n15352 ;
  assign n15522 = ~n15353 & ~n15521 ;
  assign n15523 = n15520 & n15522 ;
  assign n15524 = ~n15520 & ~n15522 ;
  assign n15525 = ~n15523 & ~n15524 ;
  assign n15526 = n15518 & n15525 ;
  assign n15527 = ~n15519 & ~n15521 ;
  assign n15528 = ~n15525 & ~n15527 ;
  assign n15529 = ~n15526 & ~n15528 ;
  assign n15530 = n15467 & n15529 ;
  assign n15543 = \core_eu_em_mac_em_reg_mxopwe_DO_reg[1]/P0001  & ~n14891 ;
  assign n15542 = ~\core_eu_em_mac_em_reg_mxopwe_DO_reg[1]/P0001  & ~n14887 ;
  assign n15544 = ~\core_eu_em_mac_em_reg_mxopwe_DO_reg[0]/P0001  & n14898 ;
  assign n15545 = \core_eu_em_mac_em_reg_mxopwe_DO_reg[0]/P0001  & n14902 ;
  assign n15546 = ~n15544 & ~n15545 ;
  assign n15547 = ~n15542 & n15546 ;
  assign n15548 = ~n15543 & n15547 ;
  assign n15550 = \core_eu_em_mac_em_reg_mxopwe_DO_reg[3]/P0001  & ~n14865 ;
  assign n15549 = ~\core_eu_em_mac_em_reg_mxopwe_DO_reg[3]/P0001  & ~n14861 ;
  assign n15551 = ~\core_eu_em_mac_em_reg_mxopwe_DO_reg[2]/P0001  & n14872 ;
  assign n15552 = \core_eu_em_mac_em_reg_mxopwe_DO_reg[2]/P0001  & n14876 ;
  assign n15553 = ~n15551 & ~n15552 ;
  assign n15554 = ~n15549 & n15553 ;
  assign n15555 = ~n15550 & n15554 ;
  assign n15556 = ~n15548 & ~n15555 ;
  assign n15557 = n15548 & n15555 ;
  assign n15558 = ~n15556 & ~n15557 ;
  assign n15559 = n15541 & n15558 ;
  assign n15560 = ~\core_eu_em_mac_em_reg_mxopwe_DO_reg[0]/P0001  & ~n14914 ;
  assign n15561 = \core_eu_em_mac_em_reg_mxopwe_DO_reg[0]/P0001  & ~n14918 ;
  assign n15562 = ~n15560 & ~n15561 ;
  assign n15564 = \core_eu_em_mac_em_reg_mxopwe_DO_reg[2]/P0001  & ~n14891 ;
  assign n15563 = ~\core_eu_em_mac_em_reg_mxopwe_DO_reg[2]/P0001  & ~n14887 ;
  assign n15565 = ~\core_eu_em_mac_em_reg_mxopwe_DO_reg[1]/P0001  & n14898 ;
  assign n15566 = \core_eu_em_mac_em_reg_mxopwe_DO_reg[1]/P0001  & n14902 ;
  assign n15567 = ~n15565 & ~n15566 ;
  assign n15568 = ~n15563 & n15567 ;
  assign n15569 = ~n15564 & n15568 ;
  assign n15570 = n15562 & n15569 ;
  assign n15571 = ~n15562 & ~n15569 ;
  assign n15572 = ~n15570 & ~n15571 ;
  assign n15574 = \core_eu_em_mac_em_reg_mxopwe_DO_reg[4]/P0001  & ~n14865 ;
  assign n15573 = ~\core_eu_em_mac_em_reg_mxopwe_DO_reg[4]/P0001  & ~n14861 ;
  assign n15575 = ~\core_eu_em_mac_em_reg_mxopwe_DO_reg[3]/P0001  & n14872 ;
  assign n15576 = \core_eu_em_mac_em_reg_mxopwe_DO_reg[3]/P0001  & n14876 ;
  assign n15577 = ~n15575 & ~n15576 ;
  assign n15578 = ~n15573 & n15577 ;
  assign n15579 = ~n15574 & n15578 ;
  assign n15580 = ~n15572 & n15579 ;
  assign n15581 = n15572 & ~n15579 ;
  assign n15582 = ~n15580 & ~n15581 ;
  assign n15583 = n15556 & n15582 ;
  assign n15584 = ~n15556 & ~n15582 ;
  assign n15585 = ~n15583 & ~n15584 ;
  assign n15586 = ~n15559 & ~n15585 ;
  assign n15587 = ~n15530 & ~n15586 ;
  assign n15588 = ~n15437 & ~n15459 ;
  assign n15589 = ~n15424 & ~n15433 ;
  assign n15590 = ~n15425 & ~n15589 ;
  assign n15592 = \core_eu_em_mac_em_reg_mxopwe_DO_reg[9]/P0001  & ~n14791 ;
  assign n15591 = ~\core_eu_em_mac_em_reg_mxopwe_DO_reg[9]/P0001  & ~n14787 ;
  assign n15593 = ~\core_eu_em_mac_em_reg_mxopwe_DO_reg[8]/P0001  & n14798 ;
  assign n15594 = \core_eu_em_mac_em_reg_mxopwe_DO_reg[8]/P0001  & n14802 ;
  assign n15595 = ~n15593 & ~n15594 ;
  assign n15596 = ~n15591 & n15595 ;
  assign n15597 = ~n15592 & n15596 ;
  assign n15599 = \core_eu_em_mac_em_reg_mxopwe_DO_reg[11]/P0001  & ~n14765 ;
  assign n15598 = ~\core_eu_em_mac_em_reg_mxopwe_DO_reg[11]/P0001  & ~n14761 ;
  assign n15600 = ~\core_eu_em_mac_em_reg_mxopwe_DO_reg[10]/P0001  & n14772 ;
  assign n15601 = \core_eu_em_mac_em_reg_mxopwe_DO_reg[10]/P0001  & n14776 ;
  assign n15602 = ~n15600 & ~n15601 ;
  assign n15603 = ~n15598 & n15602 ;
  assign n15604 = ~n15599 & n15603 ;
  assign n15605 = n15597 & n15604 ;
  assign n15606 = ~n15597 & ~n15604 ;
  assign n15607 = ~n15605 & ~n15606 ;
  assign n15609 = \core_eu_em_mac_em_reg_mxopwe_DO_reg[7]/P0001  & ~n14818 ;
  assign n15608 = ~\core_eu_em_mac_em_reg_mxopwe_DO_reg[7]/P0001  & ~n14814 ;
  assign n15610 = ~\core_eu_em_mac_em_reg_mxopwe_DO_reg[6]/P0001  & n14825 ;
  assign n15611 = \core_eu_em_mac_em_reg_mxopwe_DO_reg[6]/P0001  & n14829 ;
  assign n15612 = ~n15610 & ~n15611 ;
  assign n15613 = ~n15608 & n15612 ;
  assign n15614 = ~n15609 & n15613 ;
  assign n15615 = ~n15607 & n15614 ;
  assign n15616 = n15607 & ~n15614 ;
  assign n15617 = ~n15615 & ~n15616 ;
  assign n15618 = n15590 & ~n15617 ;
  assign n15619 = ~n15590 & n15617 ;
  assign n15620 = ~n15618 & ~n15619 ;
  assign n15621 = ~n11878 & n14993 ;
  assign n15622 = ~n7182 & n15044 ;
  assign n15623 = ~n15621 & ~n15622 ;
  assign n15624 = ~\core_eu_em_mac_em_dec_emcorepi_DO_reg[1]/P0001  & ~n15623 ;
  assign n15625 = ~n14925 & ~n15624 ;
  assign n15626 = n14925 & n15624 ;
  assign n15627 = ~n15625 & ~n15626 ;
  assign n15629 = \core_eu_em_mac_em_reg_mxopwe_DO_reg[13]/P0001  & ~n14842 ;
  assign n15628 = ~\core_eu_em_mac_em_reg_mxopwe_DO_reg[13]/P0001  & ~n14838 ;
  assign n15630 = ~\core_eu_em_mac_em_reg_mxopwe_DO_reg[12]/P0001  & n14846 ;
  assign n15631 = \core_eu_em_mac_em_reg_mxopwe_DO_reg[12]/P0001  & n14849 ;
  assign n15632 = ~n15630 & ~n15631 ;
  assign n15633 = ~n15628 & n15632 ;
  assign n15634 = ~n15629 & n15633 ;
  assign n15635 = ~n15627 & n15634 ;
  assign n15636 = n15627 & ~n15634 ;
  assign n15637 = ~n15635 & ~n15636 ;
  assign n15638 = n14914 & ~n15453 ;
  assign n15639 = ~n15454 & ~n15638 ;
  assign n15640 = ~n15637 & ~n15639 ;
  assign n15641 = n15637 & n15639 ;
  assign n15642 = ~n15640 & ~n15641 ;
  assign n15643 = n15620 & n15642 ;
  assign n15644 = ~n15620 & ~n15642 ;
  assign n15645 = ~n15643 & ~n15644 ;
  assign n15646 = ~n15588 & n15645 ;
  assign n15647 = n15588 & ~n15645 ;
  assign n15648 = ~n15646 & ~n15647 ;
  assign n15649 = ~n15438 & ~n15460 ;
  assign n15650 = ~n15464 & n15649 ;
  assign n15651 = ~n15465 & ~n15650 ;
  assign n15652 = n15648 & ~n15651 ;
  assign n15653 = ~n15648 & n15651 ;
  assign n15654 = ~n15652 & ~n15653 ;
  assign n15655 = ~n15570 & ~n15579 ;
  assign n15656 = ~n15571 & ~n15655 ;
  assign n15658 = \core_eu_em_mac_em_reg_mxopwe_DO_reg[5]/P0001  & ~n14865 ;
  assign n15657 = ~\core_eu_em_mac_em_reg_mxopwe_DO_reg[5]/P0001  & ~n14861 ;
  assign n15659 = ~\core_eu_em_mac_em_reg_mxopwe_DO_reg[4]/P0001  & n14872 ;
  assign n15660 = \core_eu_em_mac_em_reg_mxopwe_DO_reg[4]/P0001  & n14876 ;
  assign n15661 = ~n15659 & ~n15660 ;
  assign n15662 = ~n15657 & n15661 ;
  assign n15663 = ~n15658 & n15662 ;
  assign n15665 = \core_eu_em_mac_em_reg_mxopwe_DO_reg[1]/P0001  & ~n14918 ;
  assign n15664 = ~\core_eu_em_mac_em_reg_mxopwe_DO_reg[1]/P0001  & ~n14914 ;
  assign n15666 = ~\core_eu_em_mac_em_reg_mxopwe_DO_reg[0]/P0001  & n14925 ;
  assign n15667 = \core_eu_em_mac_em_reg_mxopwe_DO_reg[0]/P0001  & n14929 ;
  assign n15668 = ~n15666 & ~n15667 ;
  assign n15669 = ~n15664 & n15668 ;
  assign n15670 = ~n15665 & n15669 ;
  assign n15671 = n15663 & n15670 ;
  assign n15672 = ~n15663 & ~n15670 ;
  assign n15673 = ~n15671 & ~n15672 ;
  assign n15675 = \core_eu_em_mac_em_reg_mxopwe_DO_reg[3]/P0001  & ~n14891 ;
  assign n15674 = ~\core_eu_em_mac_em_reg_mxopwe_DO_reg[3]/P0001  & ~n14887 ;
  assign n15676 = ~\core_eu_em_mac_em_reg_mxopwe_DO_reg[2]/P0001  & n14898 ;
  assign n15677 = \core_eu_em_mac_em_reg_mxopwe_DO_reg[2]/P0001  & n14902 ;
  assign n15678 = ~n15676 & ~n15677 ;
  assign n15679 = ~n15674 & n15678 ;
  assign n15680 = ~n15675 & n15679 ;
  assign n15681 = ~n15673 & n15680 ;
  assign n15682 = n15673 & ~n15680 ;
  assign n15683 = ~n15681 & ~n15682 ;
  assign n15684 = n15656 & ~n15683 ;
  assign n15685 = ~n15656 & n15683 ;
  assign n15686 = ~n15684 & ~n15685 ;
  assign n15687 = ~n15583 & ~n15686 ;
  assign n15688 = n15583 & n15686 ;
  assign n15689 = ~n15687 & ~n15688 ;
  assign n15690 = n15654 & n15689 ;
  assign n15691 = ~n15654 & ~n15689 ;
  assign n15692 = ~n15690 & ~n15691 ;
  assign n15693 = n15587 & ~n15692 ;
  assign n15694 = ~n15587 & n15692 ;
  assign n15695 = ~n15693 & ~n15694 ;
  assign n15696 = ~n15541 & ~n15558 ;
  assign n15697 = ~n15559 & ~n15696 ;
  assign n15698 = ~n15518 & ~n15525 ;
  assign n15699 = ~n15526 & ~n15698 ;
  assign n15759 = ~n15751 & ~n15753 ;
  assign n15760 = ~n15757 & n15759 ;
  assign n15761 = ~n15758 & ~n15760 ;
  assign n15762 = ~n15699 & ~n15761 ;
  assign n15763 = n15697 & ~n15762 ;
  assign n15764 = ~n15467 & ~n15529 ;
  assign n15765 = ~n15530 & ~n15764 ;
  assign n15766 = n15559 & n15582 ;
  assign n15767 = ~n15586 & ~n15766 ;
  assign n15768 = n15765 & n15767 ;
  assign n15769 = ~n15765 & ~n15767 ;
  assign n15770 = ~n15768 & ~n15769 ;
  assign n15771 = ~n15763 & n15770 ;
  assign n15772 = ~n15764 & ~n15766 ;
  assign n15773 = ~n15770 & n15772 ;
  assign n15774 = ~n15771 & ~n15773 ;
  assign n15775 = n15695 & ~n15774 ;
  assign n15776 = ~n15652 & ~n15687 ;
  assign n15777 = ~\core_c_psq_MSTAT_reg_DO_reg[4]/NET0131  & \core_eu_em_mac_em_dec_emcorepi_DO_reg[0]/P0001  ;
  assign n15778 = \core_eu_em_mac_em_reg_mxopwe_DO_reg[0]/P0001  & ~n14951 ;
  assign n15779 = ~\core_eu_em_mac_em_reg_mxopwe_DO_reg[0]/P0001  & ~n14947 ;
  assign n15780 = ~n15778 & ~n15779 ;
  assign n15781 = n15777 & ~n15780 ;
  assign n15782 = ~n15777 & n15780 ;
  assign n15783 = ~n15781 & ~n15782 ;
  assign n15784 = ~n15671 & ~n15680 ;
  assign n15785 = ~n15672 & ~n15784 ;
  assign n15787 = \core_eu_em_mac_em_reg_mxopwe_DO_reg[4]/P0001  & ~n14891 ;
  assign n15786 = ~\core_eu_em_mac_em_reg_mxopwe_DO_reg[4]/P0001  & ~n14887 ;
  assign n15788 = ~\core_eu_em_mac_em_reg_mxopwe_DO_reg[3]/P0001  & n14898 ;
  assign n15789 = \core_eu_em_mac_em_reg_mxopwe_DO_reg[3]/P0001  & n14902 ;
  assign n15790 = ~n15788 & ~n15789 ;
  assign n15791 = ~n15786 & n15790 ;
  assign n15792 = ~n15787 & n15791 ;
  assign n15794 = \core_eu_em_mac_em_reg_mxopwe_DO_reg[6]/P0001  & ~n14865 ;
  assign n15793 = ~\core_eu_em_mac_em_reg_mxopwe_DO_reg[6]/P0001  & ~n14861 ;
  assign n15795 = ~\core_eu_em_mac_em_reg_mxopwe_DO_reg[5]/P0001  & n14872 ;
  assign n15796 = \core_eu_em_mac_em_reg_mxopwe_DO_reg[5]/P0001  & n14876 ;
  assign n15797 = ~n15795 & ~n15796 ;
  assign n15798 = ~n15793 & n15797 ;
  assign n15799 = ~n15794 & n15798 ;
  assign n15800 = n15792 & n15799 ;
  assign n15801 = ~n15792 & ~n15799 ;
  assign n15802 = ~n15800 & ~n15801 ;
  assign n15804 = \core_eu_em_mac_em_reg_mxopwe_DO_reg[2]/P0001  & ~n14918 ;
  assign n15803 = ~\core_eu_em_mac_em_reg_mxopwe_DO_reg[2]/P0001  & ~n14914 ;
  assign n15805 = ~\core_eu_em_mac_em_reg_mxopwe_DO_reg[1]/P0001  & n14925 ;
  assign n15806 = \core_eu_em_mac_em_reg_mxopwe_DO_reg[1]/P0001  & n14929 ;
  assign n15807 = ~n15805 & ~n15806 ;
  assign n15808 = ~n15803 & n15807 ;
  assign n15809 = ~n15804 & n15808 ;
  assign n15810 = ~n15802 & n15809 ;
  assign n15811 = n15802 & ~n15809 ;
  assign n15812 = ~n15810 & ~n15811 ;
  assign n15813 = ~n15785 & n15812 ;
  assign n15814 = n15785 & ~n15812 ;
  assign n15815 = ~n15813 & ~n15814 ;
  assign n15816 = n15783 & n15815 ;
  assign n15817 = ~n15783 & ~n15815 ;
  assign n15818 = ~n15816 & ~n15817 ;
  assign n15819 = ~n15685 & ~n15818 ;
  assign n15820 = n15685 & n15818 ;
  assign n15821 = ~n15819 & ~n15820 ;
  assign n15822 = ~n15618 & ~n15640 ;
  assign n15823 = ~n15605 & ~n15614 ;
  assign n15824 = ~n15606 & ~n15823 ;
  assign n15826 = \core_eu_em_mac_em_reg_mxopwe_DO_reg[10]/P0001  & ~n14791 ;
  assign n15825 = ~\core_eu_em_mac_em_reg_mxopwe_DO_reg[10]/P0001  & ~n14787 ;
  assign n15827 = ~\core_eu_em_mac_em_reg_mxopwe_DO_reg[9]/P0001  & n14798 ;
  assign n15828 = \core_eu_em_mac_em_reg_mxopwe_DO_reg[9]/P0001  & n14802 ;
  assign n15829 = ~n15827 & ~n15828 ;
  assign n15830 = ~n15825 & n15829 ;
  assign n15831 = ~n15826 & n15830 ;
  assign n15833 = \core_eu_em_mac_em_reg_mxopwe_DO_reg[12]/P0001  & ~n14765 ;
  assign n15832 = ~\core_eu_em_mac_em_reg_mxopwe_DO_reg[12]/P0001  & ~n14761 ;
  assign n15834 = ~\core_eu_em_mac_em_reg_mxopwe_DO_reg[11]/P0001  & n14772 ;
  assign n15835 = \core_eu_em_mac_em_reg_mxopwe_DO_reg[11]/P0001  & n14776 ;
  assign n15836 = ~n15834 & ~n15835 ;
  assign n15837 = ~n15832 & n15836 ;
  assign n15838 = ~n15833 & n15837 ;
  assign n15839 = n15831 & n15838 ;
  assign n15840 = ~n15831 & ~n15838 ;
  assign n15841 = ~n15839 & ~n15840 ;
  assign n15843 = \core_eu_em_mac_em_reg_mxopwe_DO_reg[8]/P0001  & ~n14818 ;
  assign n15842 = ~\core_eu_em_mac_em_reg_mxopwe_DO_reg[8]/P0001  & ~n14814 ;
  assign n15844 = ~\core_eu_em_mac_em_reg_mxopwe_DO_reg[7]/P0001  & n14825 ;
  assign n15845 = \core_eu_em_mac_em_reg_mxopwe_DO_reg[7]/P0001  & n14829 ;
  assign n15846 = ~n15844 & ~n15845 ;
  assign n15847 = ~n15842 & n15846 ;
  assign n15848 = ~n15843 & n15847 ;
  assign n15849 = ~n15841 & n15848 ;
  assign n15850 = n15841 & ~n15848 ;
  assign n15851 = ~n15849 & ~n15850 ;
  assign n15852 = n15824 & ~n15851 ;
  assign n15853 = ~n15824 & n15851 ;
  assign n15854 = ~n15852 & ~n15853 ;
  assign n15855 = ~n15625 & ~n15634 ;
  assign n15856 = ~n15626 & ~n15855 ;
  assign n15857 = ~n12024 & n14993 ;
  assign n15858 = ~n11878 & n15044 ;
  assign n15859 = ~n15857 & ~n15858 ;
  assign n15860 = ~\core_eu_em_mac_em_dec_emcorepi_DO_reg[1]/P0001  & ~n15859 ;
  assign n15862 = \core_eu_em_mac_em_reg_mxopwe_DO_reg[14]/P0001  & ~n14842 ;
  assign n15861 = ~\core_eu_em_mac_em_reg_mxopwe_DO_reg[14]/P0001  & ~n14838 ;
  assign n15863 = ~\core_eu_em_mac_em_reg_mxopwe_DO_reg[13]/P0001  & n14846 ;
  assign n15864 = \core_eu_em_mac_em_reg_mxopwe_DO_reg[13]/P0001  & n14849 ;
  assign n15865 = ~n15863 & ~n15864 ;
  assign n15866 = ~n15861 & n15865 ;
  assign n15867 = ~n15862 & n15866 ;
  assign n15868 = ~n15860 & n15867 ;
  assign n15869 = n15860 & ~n15867 ;
  assign n15870 = ~n15868 & ~n15869 ;
  assign n15871 = n14947 & n15870 ;
  assign n15872 = ~n14947 & ~n15870 ;
  assign n15873 = ~n15871 & ~n15872 ;
  assign n15874 = n15856 & n15873 ;
  assign n15875 = ~n15856 & ~n15873 ;
  assign n15876 = ~n15874 & ~n15875 ;
  assign n15877 = n15854 & n15876 ;
  assign n15878 = ~n15854 & ~n15876 ;
  assign n15879 = ~n15877 & ~n15878 ;
  assign n15880 = ~n15822 & n15879 ;
  assign n15881 = n15822 & ~n15879 ;
  assign n15882 = ~n15880 & ~n15881 ;
  assign n15883 = ~n15619 & ~n15641 ;
  assign n15884 = ~n15645 & n15883 ;
  assign n15885 = ~n15646 & ~n15884 ;
  assign n15886 = n15882 & ~n15885 ;
  assign n15887 = ~n15882 & n15885 ;
  assign n15888 = ~n15886 & ~n15887 ;
  assign n15889 = n15821 & n15888 ;
  assign n15890 = ~n15821 & ~n15888 ;
  assign n15891 = ~n15889 & ~n15890 ;
  assign n15892 = ~n15776 & n15891 ;
  assign n15893 = n15776 & ~n15891 ;
  assign n15894 = ~n15892 & ~n15893 ;
  assign n15895 = ~n15653 & ~n15688 ;
  assign n15896 = ~n15692 & n15895 ;
  assign n15897 = ~n15694 & ~n15896 ;
  assign n15898 = n15894 & ~n15897 ;
  assign n15899 = ~n15775 & ~n15898 ;
  assign n15967 = n15901 & ~n15966 ;
  assign n15968 = n15699 & n15761 ;
  assign n15969 = ~n15762 & ~n15968 ;
  assign n15970 = n15697 & ~n15969 ;
  assign n15971 = ~n15697 & n15969 ;
  assign n15972 = ~n15970 & ~n15971 ;
  assign n15973 = ~n15967 & ~n15972 ;
  assign n15974 = ~n15968 & n15972 ;
  assign n15975 = ~n15973 & ~n15974 ;
  assign n15976 = n15763 & ~n15770 ;
  assign n15977 = ~n15771 & ~n15976 ;
  assign n15978 = ~n15975 & n15977 ;
  assign n16054 = ~n16048 & ~n16052 ;
  assign n16055 = ~n16053 & ~n16054 ;
  assign n16056 = n15967 & n15972 ;
  assign n16057 = ~n15973 & ~n16056 ;
  assign n16058 = ~n16055 & n16057 ;
  assign n16059 = ~n15978 & ~n16058 ;
  assign n16351 = n15899 & n16059 ;
  assign n16352 = ~n16350 & n16351 ;
  assign n16355 = n15975 & ~n15977 ;
  assign n16356 = n16055 & ~n16057 ;
  assign n16357 = ~n15978 & n16356 ;
  assign n16358 = ~n16355 & ~n16357 ;
  assign n16359 = n15899 & ~n16358 ;
  assign n16353 = ~n15695 & n15774 ;
  assign n16354 = ~n15898 & n16353 ;
  assign n16360 = ~n15894 & n15897 ;
  assign n16361 = ~n16354 & ~n16360 ;
  assign n16362 = ~n16359 & n16361 ;
  assign n16363 = ~n16352 & n16362 ;
  assign n16364 = ~n14779 & ~n14805 ;
  assign n16366 = \core_eu_em_mac_em_reg_mxopwe_DO_reg[15]/P0001  & ~n14818 ;
  assign n16365 = ~\core_eu_em_mac_em_reg_mxopwe_DO_reg[15]/P0001  & ~n14814 ;
  assign n16367 = ~\core_eu_em_mac_em_reg_mxopwe_DO_reg[14]/P0001  & n14825 ;
  assign n16368 = \core_eu_em_mac_em_reg_mxopwe_DO_reg[14]/P0001  & n14829 ;
  assign n16369 = ~n16367 & ~n16368 ;
  assign n16370 = ~n16365 & n16369 ;
  assign n16371 = ~n16366 & n16370 ;
  assign n16372 = ~n14806 & ~n16371 ;
  assign n16373 = ~n16364 & ~n16372 ;
  assign n16374 = ~n14806 & ~n16364 ;
  assign n16375 = ~\core_eu_em_mac_em_reg_mxopwe_DO_reg[15]/P0001  & n14825 ;
  assign n16376 = \core_eu_em_mac_em_reg_mxopwe_DO_reg[15]/P0001  & n14829 ;
  assign n16377 = ~n16375 & ~n16376 ;
  assign n16378 = n14820 & n16377 ;
  assign n16379 = n16374 & ~n16378 ;
  assign n16380 = ~n16374 & n16378 ;
  assign n16381 = ~n16379 & ~n16380 ;
  assign n16382 = n16373 & ~n16381 ;
  assign n16383 = ~n14852 & ~n16382 ;
  assign n16384 = ~n14806 & ~n16378 ;
  assign n16385 = ~n16364 & ~n16384 ;
  assign n16386 = ~n14832 & n16374 ;
  assign n16387 = n14832 & ~n16374 ;
  assign n16388 = ~n16386 & ~n16387 ;
  assign n16389 = ~n16385 & n16388 ;
  assign n16390 = n16385 & ~n16388 ;
  assign n16391 = ~n16389 & ~n16390 ;
  assign n16392 = ~n14852 & n16391 ;
  assign n16393 = n14852 & ~n16391 ;
  assign n16394 = ~n16392 & ~n16393 ;
  assign n16395 = ~n16383 & n16394 ;
  assign n16396 = ~n16382 & n16392 ;
  assign n16397 = ~n16395 & ~n16396 ;
  assign n16398 = ~\core_eu_em_mac_em_reg_mxopwe_DO_reg[15]/P0001  & n14798 ;
  assign n16399 = \core_eu_em_mac_em_reg_mxopwe_DO_reg[15]/P0001  & n14802 ;
  assign n16400 = ~n16398 & ~n16399 ;
  assign n16401 = n14793 & n16400 ;
  assign n16402 = n14779 & n16401 ;
  assign n16404 = \core_eu_em_mac_em_reg_mxopwe_DO_reg[14]/P0001  & ~n14818 ;
  assign n16403 = ~\core_eu_em_mac_em_reg_mxopwe_DO_reg[14]/P0001  & ~n14814 ;
  assign n16405 = ~\core_eu_em_mac_em_reg_mxopwe_DO_reg[13]/P0001  & n14825 ;
  assign n16406 = \core_eu_em_mac_em_reg_mxopwe_DO_reg[13]/P0001  & n14829 ;
  assign n16407 = ~n16405 & ~n16406 ;
  assign n16408 = ~n16403 & n16407 ;
  assign n16409 = ~n16404 & n16408 ;
  assign n16410 = ~n16402 & ~n16409 ;
  assign n16411 = ~n14779 & ~n16401 ;
  assign n16412 = ~n16410 & ~n16411 ;
  assign n16413 = ~n16371 & n16374 ;
  assign n16414 = n16371 & ~n16374 ;
  assign n16415 = ~n16413 & ~n16414 ;
  assign n16416 = n16412 & ~n16415 ;
  assign n16417 = ~n14852 & ~n16416 ;
  assign n16418 = ~n16373 & n16381 ;
  assign n16419 = ~n16382 & ~n16418 ;
  assign n16420 = n14852 & ~n16419 ;
  assign n16421 = n16383 & ~n16418 ;
  assign n16422 = ~n16420 & ~n16421 ;
  assign n16423 = ~n16417 & n16422 ;
  assign n16424 = ~n16418 & ~n16422 ;
  assign n16425 = ~n16423 & ~n16424 ;
  assign n16426 = n16397 & ~n16425 ;
  assign n16428 = ~\core_eu_em_mac_em_reg_mxopwe_DO_reg[13]/P0001  & ~n14861 ;
  assign n16427 = \core_eu_em_mac_em_reg_mxopwe_DO_reg[13]/P0001  & ~n14865 ;
  assign n16429 = ~\core_eu_em_mac_em_reg_mxopwe_DO_reg[12]/P0001  & n14872 ;
  assign n16430 = \core_eu_em_mac_em_reg_mxopwe_DO_reg[12]/P0001  & n14876 ;
  assign n16431 = ~n16429 & ~n16430 ;
  assign n16432 = ~n16427 & n16431 ;
  assign n16433 = ~n16428 & n16432 ;
  assign n16435 = \core_eu_em_mac_em_reg_mxopwe_DO_reg[11]/P0001  & ~n14891 ;
  assign n16434 = ~\core_eu_em_mac_em_reg_mxopwe_DO_reg[11]/P0001  & ~n14887 ;
  assign n16436 = ~\core_eu_em_mac_em_reg_mxopwe_DO_reg[10]/P0001  & n14898 ;
  assign n16437 = \core_eu_em_mac_em_reg_mxopwe_DO_reg[10]/P0001  & n14902 ;
  assign n16438 = ~n16436 & ~n16437 ;
  assign n16439 = ~n16434 & n16438 ;
  assign n16440 = ~n16435 & n16439 ;
  assign n16441 = n16433 & n16440 ;
  assign n16443 = \core_eu_em_mac_em_reg_mxopwe_DO_reg[9]/P0001  & ~n14918 ;
  assign n16442 = ~\core_eu_em_mac_em_reg_mxopwe_DO_reg[9]/P0001  & ~n14914 ;
  assign n16444 = ~\core_eu_em_mac_em_reg_mxopwe_DO_reg[8]/P0001  & n14925 ;
  assign n16445 = \core_eu_em_mac_em_reg_mxopwe_DO_reg[8]/P0001  & n14929 ;
  assign n16446 = ~n16444 & ~n16445 ;
  assign n16447 = ~n16442 & n16446 ;
  assign n16448 = ~n16443 & n16447 ;
  assign n16449 = ~n16441 & ~n16448 ;
  assign n16450 = ~n16433 & ~n16440 ;
  assign n16451 = ~n16449 & ~n16450 ;
  assign n16453 = \core_eu_em_mac_em_reg_mxopwe_DO_reg[14]/P0001  & ~n14865 ;
  assign n16452 = ~\core_eu_em_mac_em_reg_mxopwe_DO_reg[14]/P0001  & ~n14861 ;
  assign n16454 = ~\core_eu_em_mac_em_reg_mxopwe_DO_reg[13]/P0001  & n14872 ;
  assign n16455 = \core_eu_em_mac_em_reg_mxopwe_DO_reg[13]/P0001  & n14876 ;
  assign n16456 = ~n16454 & ~n16455 ;
  assign n16457 = ~n16452 & n16456 ;
  assign n16458 = ~n16453 & n16457 ;
  assign n16460 = \core_eu_em_mac_em_reg_mxopwe_DO_reg[12]/P0001  & ~n14891 ;
  assign n16459 = ~\core_eu_em_mac_em_reg_mxopwe_DO_reg[12]/P0001  & ~n14887 ;
  assign n16461 = ~\core_eu_em_mac_em_reg_mxopwe_DO_reg[11]/P0001  & n14898 ;
  assign n16462 = \core_eu_em_mac_em_reg_mxopwe_DO_reg[11]/P0001  & n14902 ;
  assign n16463 = ~n16461 & ~n16462 ;
  assign n16464 = ~n16459 & n16463 ;
  assign n16465 = ~n16460 & n16464 ;
  assign n16466 = n16458 & n16465 ;
  assign n16467 = ~n16458 & ~n16465 ;
  assign n16468 = ~n16466 & ~n16467 ;
  assign n16470 = \core_eu_em_mac_em_reg_mxopwe_DO_reg[10]/P0001  & ~n14918 ;
  assign n16469 = ~\core_eu_em_mac_em_reg_mxopwe_DO_reg[10]/P0001  & ~n14914 ;
  assign n16471 = ~\core_eu_em_mac_em_reg_mxopwe_DO_reg[9]/P0001  & n14925 ;
  assign n16472 = \core_eu_em_mac_em_reg_mxopwe_DO_reg[9]/P0001  & n14929 ;
  assign n16473 = ~n16471 & ~n16472 ;
  assign n16474 = ~n16469 & n16473 ;
  assign n16475 = ~n16470 & n16474 ;
  assign n16476 = ~n16468 & n16475 ;
  assign n16477 = n16468 & ~n16475 ;
  assign n16478 = ~n16476 & ~n16477 ;
  assign n16479 = n16451 & ~n16478 ;
  assign n16480 = ~\core_eu_em_mac_em_reg_mxopwe_DO_reg[6]/P0001  & ~n14967 ;
  assign n16481 = \core_eu_em_mac_em_reg_mxopwe_DO_reg[6]/P0001  & ~n14969 ;
  assign n16482 = ~n16480 & ~n16481 ;
  assign n16484 = \core_eu_em_mac_em_reg_mxopwe_DO_reg[8]/P0001  & ~n14951 ;
  assign n16483 = ~\core_eu_em_mac_em_reg_mxopwe_DO_reg[8]/P0001  & ~n14947 ;
  assign n16485 = ~\core_eu_em_mac_em_reg_mxopwe_DO_reg[7]/P0001  & n14958 ;
  assign n16486 = \core_eu_em_mac_em_reg_mxopwe_DO_reg[7]/P0001  & n14962 ;
  assign n16487 = ~n16485 & ~n16486 ;
  assign n16488 = ~n16483 & n16487 ;
  assign n16489 = ~n16484 & n16488 ;
  assign n16490 = ~n16482 & n16489 ;
  assign n16491 = n16482 & ~n16489 ;
  assign n16492 = ~n16490 & ~n16491 ;
  assign n16495 = \core_c_dec_MACop_E_reg/P0001  & ~n11196 ;
  assign n16496 = ~\core_c_psq_MSTAT_reg_DO_reg[4]/NET0131  & ~n16495 ;
  assign n16493 = \core_c_dec_MACop_E_reg/P0001  & ~n11448 ;
  assign n16494 = \core_c_psq_MSTAT_reg_DO_reg[4]/NET0131  & ~n16493 ;
  assign n16497 = ~\core_eu_em_mac_em_dec_emcorepi_DO_reg[1]/P0001  & ~n16494 ;
  assign n16498 = ~n16496 & n16497 ;
  assign n16499 = ~n16492 & n16498 ;
  assign n16500 = n16492 & ~n16498 ;
  assign n16501 = ~n16499 & ~n16500 ;
  assign n16502 = ~\core_eu_em_mac_em_reg_mxopwe_DO_reg[5]/P0001  & ~n14967 ;
  assign n16503 = \core_eu_em_mac_em_reg_mxopwe_DO_reg[5]/P0001  & ~n14969 ;
  assign n16504 = ~n16502 & ~n16503 ;
  assign n16506 = \core_eu_em_mac_em_reg_mxopwe_DO_reg[7]/P0001  & ~n14951 ;
  assign n16505 = ~\core_eu_em_mac_em_reg_mxopwe_DO_reg[7]/P0001  & ~n14947 ;
  assign n16507 = ~\core_eu_em_mac_em_reg_mxopwe_DO_reg[6]/P0001  & n14958 ;
  assign n16508 = \core_eu_em_mac_em_reg_mxopwe_DO_reg[6]/P0001  & n14962 ;
  assign n16509 = ~n16507 & ~n16508 ;
  assign n16510 = ~n16505 & n16509 ;
  assign n16511 = ~n16506 & n16510 ;
  assign n16512 = ~n16504 & n16511 ;
  assign n16513 = n16504 & ~n16511 ;
  assign n16516 = ~\core_c_psq_MSTAT_reg_DO_reg[4]/NET0131  & ~n16493 ;
  assign n16514 = \core_c_dec_MACop_E_reg/P0001  & ~n10858 ;
  assign n16515 = \core_c_psq_MSTAT_reg_DO_reg[4]/NET0131  & ~n16514 ;
  assign n16517 = ~\core_eu_em_mac_em_dec_emcorepi_DO_reg[1]/P0001  & ~n16515 ;
  assign n16518 = ~n16516 & n16517 ;
  assign n16519 = ~n16513 & ~n16518 ;
  assign n16520 = ~n16512 & ~n16519 ;
  assign n16521 = n16501 & ~n16520 ;
  assign n16522 = ~n16479 & ~n16521 ;
  assign n16523 = ~n16490 & n16498 ;
  assign n16524 = ~n16491 & ~n16523 ;
  assign n16526 = \core_c_dec_MACop_E_reg/P0001  & ~n10538 ;
  assign n16527 = ~\core_c_psq_MSTAT_reg_DO_reg[4]/NET0131  & ~n16526 ;
  assign n16525 = \core_c_psq_MSTAT_reg_DO_reg[4]/NET0131  & ~n16495 ;
  assign n16528 = ~\core_eu_em_mac_em_dec_emcorepi_DO_reg[1]/P0001  & ~n16525 ;
  assign n16529 = ~n16527 & n16528 ;
  assign n16531 = \core_eu_em_mac_em_reg_mxopwe_DO_reg[9]/P0001  & ~n14951 ;
  assign n16530 = ~\core_eu_em_mac_em_reg_mxopwe_DO_reg[9]/P0001  & ~n14947 ;
  assign n16532 = ~\core_eu_em_mac_em_reg_mxopwe_DO_reg[8]/P0001  & n14958 ;
  assign n16533 = \core_eu_em_mac_em_reg_mxopwe_DO_reg[8]/P0001  & n14962 ;
  assign n16534 = ~n16532 & ~n16533 ;
  assign n16535 = ~n16530 & n16534 ;
  assign n16536 = ~n16531 & n16535 ;
  assign n16537 = n16529 & ~n16536 ;
  assign n16538 = ~n16529 & n16536 ;
  assign n16539 = ~n16537 & ~n16538 ;
  assign n16540 = ~\core_eu_em_mac_em_reg_mxopwe_DO_reg[7]/P0001  & n14967 ;
  assign n16541 = \core_eu_em_mac_em_reg_mxopwe_DO_reg[7]/P0001  & n14969 ;
  assign n16542 = ~n16540 & ~n16541 ;
  assign n16543 = n16539 & n16542 ;
  assign n16544 = ~n16539 & ~n16542 ;
  assign n16545 = ~n16543 & ~n16544 ;
  assign n16546 = n16524 & n16545 ;
  assign n16547 = ~n16524 & ~n16545 ;
  assign n16548 = ~n16546 & ~n16547 ;
  assign n16549 = ~n16466 & ~n16475 ;
  assign n16550 = ~n16467 & ~n16549 ;
  assign n16552 = \core_eu_em_mac_em_reg_mxopwe_DO_reg[13]/P0001  & ~n14891 ;
  assign n16551 = ~\core_eu_em_mac_em_reg_mxopwe_DO_reg[13]/P0001  & ~n14887 ;
  assign n16553 = ~\core_eu_em_mac_em_reg_mxopwe_DO_reg[12]/P0001  & n14898 ;
  assign n16554 = \core_eu_em_mac_em_reg_mxopwe_DO_reg[12]/P0001  & n14902 ;
  assign n16555 = ~n16553 & ~n16554 ;
  assign n16556 = ~n16551 & n16555 ;
  assign n16557 = ~n16552 & n16556 ;
  assign n16559 = \core_eu_em_mac_em_reg_mxopwe_DO_reg[15]/P0001  & ~n14865 ;
  assign n16558 = ~\core_eu_em_mac_em_reg_mxopwe_DO_reg[15]/P0001  & ~n14861 ;
  assign n16560 = ~\core_eu_em_mac_em_reg_mxopwe_DO_reg[14]/P0001  & n14872 ;
  assign n16561 = \core_eu_em_mac_em_reg_mxopwe_DO_reg[14]/P0001  & n14876 ;
  assign n16562 = ~n16560 & ~n16561 ;
  assign n16563 = ~n16558 & n16562 ;
  assign n16564 = ~n16559 & n16563 ;
  assign n16565 = n16557 & n16564 ;
  assign n16566 = ~n16557 & ~n16564 ;
  assign n16567 = ~n16565 & ~n16566 ;
  assign n16569 = \core_eu_em_mac_em_reg_mxopwe_DO_reg[11]/P0001  & ~n14918 ;
  assign n16568 = ~\core_eu_em_mac_em_reg_mxopwe_DO_reg[11]/P0001  & ~n14914 ;
  assign n16570 = ~\core_eu_em_mac_em_reg_mxopwe_DO_reg[10]/P0001  & n14925 ;
  assign n16571 = \core_eu_em_mac_em_reg_mxopwe_DO_reg[10]/P0001  & n14929 ;
  assign n16572 = ~n16570 & ~n16571 ;
  assign n16573 = ~n16568 & n16572 ;
  assign n16574 = ~n16569 & n16573 ;
  assign n16575 = ~n16567 & n16574 ;
  assign n16576 = n16567 & ~n16574 ;
  assign n16577 = ~n16575 & ~n16576 ;
  assign n16578 = n16550 & ~n16577 ;
  assign n16579 = ~n16550 & n16577 ;
  assign n16580 = ~n16578 & ~n16579 ;
  assign n16581 = n16548 & ~n16580 ;
  assign n16582 = ~n16548 & n16580 ;
  assign n16583 = ~n16581 & ~n16582 ;
  assign n16584 = ~n16522 & ~n16583 ;
  assign n16585 = n16522 & n16583 ;
  assign n16586 = ~n16584 & ~n16585 ;
  assign n16587 = ~n16512 & ~n16513 ;
  assign n16588 = n16518 & ~n16587 ;
  assign n16589 = ~n16518 & n16587 ;
  assign n16590 = ~n16588 & ~n16589 ;
  assign n16593 = ~\core_c_psq_MSTAT_reg_DO_reg[4]/NET0131  & ~n16514 ;
  assign n16591 = \core_c_dec_MACop_E_reg/P0001  & ~n9845 ;
  assign n16592 = \core_c_psq_MSTAT_reg_DO_reg[4]/NET0131  & ~n16591 ;
  assign n16594 = ~\core_eu_em_mac_em_dec_emcorepi_DO_reg[1]/P0001  & ~n16592 ;
  assign n16595 = ~n16593 & n16594 ;
  assign n16597 = \core_eu_em_mac_em_reg_mxopwe_DO_reg[6]/P0001  & ~n14951 ;
  assign n16596 = ~\core_eu_em_mac_em_reg_mxopwe_DO_reg[6]/P0001  & ~n14947 ;
  assign n16598 = ~\core_eu_em_mac_em_reg_mxopwe_DO_reg[5]/P0001  & n14958 ;
  assign n16599 = \core_eu_em_mac_em_reg_mxopwe_DO_reg[5]/P0001  & n14962 ;
  assign n16600 = ~n16598 & ~n16599 ;
  assign n16601 = ~n16596 & n16600 ;
  assign n16602 = ~n16597 & n16601 ;
  assign n16603 = n16595 & ~n16602 ;
  assign n16604 = ~n16595 & n16602 ;
  assign n16605 = ~\core_eu_em_mac_em_reg_mxopwe_DO_reg[4]/P0001  & n14967 ;
  assign n16606 = \core_eu_em_mac_em_reg_mxopwe_DO_reg[4]/P0001  & n14969 ;
  assign n16607 = ~n16605 & ~n16606 ;
  assign n16608 = ~n16604 & ~n16607 ;
  assign n16609 = ~n16603 & ~n16608 ;
  assign n16610 = n16590 & n16609 ;
  assign n16612 = \core_eu_em_mac_em_reg_mxopwe_DO_reg[10]/P0001  & ~n14891 ;
  assign n16611 = ~\core_eu_em_mac_em_reg_mxopwe_DO_reg[10]/P0001  & ~n14887 ;
  assign n16613 = ~\core_eu_em_mac_em_reg_mxopwe_DO_reg[9]/P0001  & n14898 ;
  assign n16614 = \core_eu_em_mac_em_reg_mxopwe_DO_reg[9]/P0001  & n14902 ;
  assign n16615 = ~n16613 & ~n16614 ;
  assign n16616 = ~n16611 & n16615 ;
  assign n16617 = ~n16612 & n16616 ;
  assign n16619 = \core_eu_em_mac_em_reg_mxopwe_DO_reg[12]/P0001  & ~n14865 ;
  assign n16618 = ~\core_eu_em_mac_em_reg_mxopwe_DO_reg[12]/P0001  & ~n14861 ;
  assign n16620 = ~\core_eu_em_mac_em_reg_mxopwe_DO_reg[11]/P0001  & n14872 ;
  assign n16621 = \core_eu_em_mac_em_reg_mxopwe_DO_reg[11]/P0001  & n14876 ;
  assign n16622 = ~n16620 & ~n16621 ;
  assign n16623 = ~n16618 & n16622 ;
  assign n16624 = ~n16619 & n16623 ;
  assign n16625 = n16617 & n16624 ;
  assign n16627 = \core_eu_em_mac_em_reg_mxopwe_DO_reg[8]/P0001  & ~n14918 ;
  assign n16626 = ~\core_eu_em_mac_em_reg_mxopwe_DO_reg[8]/P0001  & ~n14914 ;
  assign n16628 = ~\core_eu_em_mac_em_reg_mxopwe_DO_reg[7]/P0001  & n14925 ;
  assign n16629 = \core_eu_em_mac_em_reg_mxopwe_DO_reg[7]/P0001  & n14929 ;
  assign n16630 = ~n16628 & ~n16629 ;
  assign n16631 = ~n16626 & n16630 ;
  assign n16632 = ~n16627 & n16631 ;
  assign n16633 = ~n16625 & ~n16632 ;
  assign n16634 = ~n16617 & ~n16624 ;
  assign n16635 = ~n16633 & ~n16634 ;
  assign n16636 = ~n16441 & ~n16450 ;
  assign n16637 = n16448 & ~n16636 ;
  assign n16638 = ~n16448 & n16636 ;
  assign n16639 = ~n16637 & ~n16638 ;
  assign n16640 = n16635 & ~n16639 ;
  assign n16641 = ~n16610 & ~n16640 ;
  assign n16642 = ~n16451 & n16478 ;
  assign n16643 = ~n16479 & ~n16642 ;
  assign n16644 = ~n16501 & n16520 ;
  assign n16645 = ~n16521 & ~n16644 ;
  assign n16646 = n16643 & n16645 ;
  assign n16647 = ~n16643 & ~n16645 ;
  assign n16648 = ~n16646 & ~n16647 ;
  assign n16649 = ~n16641 & n16648 ;
  assign n16650 = ~n16642 & ~n16644 ;
  assign n16651 = ~n16648 & n16650 ;
  assign n16652 = ~n16649 & ~n16651 ;
  assign n16653 = n16586 & ~n16652 ;
  assign n16654 = ~n16426 & ~n16653 ;
  assign n16655 = ~n16546 & ~n16578 ;
  assign n16656 = ~n16565 & ~n16574 ;
  assign n16657 = ~n16566 & ~n16656 ;
  assign n16658 = ~\core_eu_em_mac_em_reg_mxopwe_DO_reg[15]/P0001  & n14872 ;
  assign n16659 = \core_eu_em_mac_em_reg_mxopwe_DO_reg[15]/P0001  & n14876 ;
  assign n16660 = ~n16658 & ~n16659 ;
  assign n16661 = n14867 & n16660 ;
  assign n16663 = \core_eu_em_mac_em_reg_mxopwe_DO_reg[14]/P0001  & ~n14891 ;
  assign n16662 = ~\core_eu_em_mac_em_reg_mxopwe_DO_reg[14]/P0001  & ~n14887 ;
  assign n16664 = ~\core_eu_em_mac_em_reg_mxopwe_DO_reg[13]/P0001  & n14898 ;
  assign n16665 = \core_eu_em_mac_em_reg_mxopwe_DO_reg[13]/P0001  & n14902 ;
  assign n16666 = ~n16664 & ~n16665 ;
  assign n16667 = ~n16662 & n16666 ;
  assign n16668 = ~n16663 & n16667 ;
  assign n16669 = n16661 & n16668 ;
  assign n16670 = ~n16661 & ~n16668 ;
  assign n16671 = ~n16669 & ~n16670 ;
  assign n16673 = \core_eu_em_mac_em_reg_mxopwe_DO_reg[12]/P0001  & ~n14918 ;
  assign n16672 = ~\core_eu_em_mac_em_reg_mxopwe_DO_reg[12]/P0001  & ~n14914 ;
  assign n16674 = ~\core_eu_em_mac_em_reg_mxopwe_DO_reg[11]/P0001  & n14925 ;
  assign n16675 = \core_eu_em_mac_em_reg_mxopwe_DO_reg[11]/P0001  & n14929 ;
  assign n16676 = ~n16674 & ~n16675 ;
  assign n16677 = ~n16672 & n16676 ;
  assign n16678 = ~n16673 & n16677 ;
  assign n16679 = ~n16671 & n16678 ;
  assign n16680 = n16671 & ~n16678 ;
  assign n16681 = ~n16679 & ~n16680 ;
  assign n16682 = ~n16657 & n16681 ;
  assign n16683 = n16657 & ~n16681 ;
  assign n16684 = ~n16682 & ~n16683 ;
  assign n16685 = ~\core_eu_em_mac_em_reg_mxopwe_DO_reg[8]/P0001  & ~n14967 ;
  assign n16686 = \core_eu_em_mac_em_reg_mxopwe_DO_reg[8]/P0001  & ~n14969 ;
  assign n16687 = ~n16685 & ~n16686 ;
  assign n16689 = \core_eu_em_mac_em_reg_mxopwe_DO_reg[10]/P0001  & ~n14951 ;
  assign n16688 = ~\core_eu_em_mac_em_reg_mxopwe_DO_reg[10]/P0001  & ~n14947 ;
  assign n16690 = ~\core_eu_em_mac_em_reg_mxopwe_DO_reg[9]/P0001  & n14958 ;
  assign n16691 = \core_eu_em_mac_em_reg_mxopwe_DO_reg[9]/P0001  & n14962 ;
  assign n16692 = ~n16690 & ~n16691 ;
  assign n16693 = ~n16688 & n16692 ;
  assign n16694 = ~n16689 & n16693 ;
  assign n16695 = ~n16687 & n16694 ;
  assign n16696 = n16687 & ~n16694 ;
  assign n16697 = ~n16695 & ~n16696 ;
  assign n16699 = \core_c_dec_MACop_E_reg/P0001  & ~n10096 ;
  assign n16700 = ~\core_c_psq_MSTAT_reg_DO_reg[4]/NET0131  & ~n16699 ;
  assign n16698 = \core_c_psq_MSTAT_reg_DO_reg[4]/NET0131  & ~n16526 ;
  assign n16701 = ~\core_eu_em_mac_em_dec_emcorepi_DO_reg[1]/P0001  & ~n16698 ;
  assign n16702 = ~n16700 & n16701 ;
  assign n16703 = n16697 & n16702 ;
  assign n16704 = ~n16697 & ~n16702 ;
  assign n16705 = ~n16703 & ~n16704 ;
  assign n16706 = ~n16538 & ~n16542 ;
  assign n16707 = ~n16537 & ~n16706 ;
  assign n16708 = n16705 & ~n16707 ;
  assign n16709 = ~n16705 & n16707 ;
  assign n16710 = ~n16708 & ~n16709 ;
  assign n16711 = n16684 & n16710 ;
  assign n16712 = ~n16684 & ~n16710 ;
  assign n16713 = ~n16711 & ~n16712 ;
  assign n16714 = ~n16655 & n16713 ;
  assign n16715 = n16655 & ~n16713 ;
  assign n16716 = ~n16714 & ~n16715 ;
  assign n16717 = ~n16547 & ~n16579 ;
  assign n16718 = n16583 & n16717 ;
  assign n16719 = ~n16584 & ~n16718 ;
  assign n16720 = ~n16716 & n16719 ;
  assign n16721 = n16716 & ~n16719 ;
  assign n16722 = ~n16720 & ~n16721 ;
  assign n16723 = ~n16389 & ~n16394 ;
  assign n16724 = ~n16395 & ~n16723 ;
  assign n16725 = ~n14832 & n16364 ;
  assign n16726 = ~n14833 & ~n16725 ;
  assign n16727 = ~n14852 & n16390 ;
  assign n16728 = n16726 & ~n16727 ;
  assign n16729 = ~n16726 & n16727 ;
  assign n16730 = ~n16728 & ~n16729 ;
  assign n16731 = n16724 & ~n16730 ;
  assign n16732 = ~n16724 & n16730 ;
  assign n16733 = ~n16731 & ~n16732 ;
  assign n16734 = n16722 & n16733 ;
  assign n16735 = ~n16722 & ~n16733 ;
  assign n16736 = ~n16734 & ~n16735 ;
  assign n16737 = ~n16654 & n16736 ;
  assign n16738 = n16654 & ~n16736 ;
  assign n16739 = ~n16737 & ~n16738 ;
  assign n16740 = n16417 & n16419 ;
  assign n16741 = ~n16423 & ~n16740 ;
  assign n16743 = \core_eu_em_mac_em_reg_mxopwe_DO_reg[15]/P0001  & ~n14791 ;
  assign n16742 = ~\core_eu_em_mac_em_reg_mxopwe_DO_reg[15]/P0001  & ~n14787 ;
  assign n16744 = ~\core_eu_em_mac_em_reg_mxopwe_DO_reg[14]/P0001  & n14798 ;
  assign n16745 = \core_eu_em_mac_em_reg_mxopwe_DO_reg[14]/P0001  & n14802 ;
  assign n16746 = ~n16744 & ~n16745 ;
  assign n16747 = ~n16742 & n16746 ;
  assign n16748 = ~n16743 & n16747 ;
  assign n16749 = n14779 & n16748 ;
  assign n16751 = \core_eu_em_mac_em_reg_mxopwe_DO_reg[13]/P0001  & ~n14818 ;
  assign n16750 = ~\core_eu_em_mac_em_reg_mxopwe_DO_reg[13]/P0001  & ~n14814 ;
  assign n16752 = ~\core_eu_em_mac_em_reg_mxopwe_DO_reg[12]/P0001  & n14825 ;
  assign n16753 = \core_eu_em_mac_em_reg_mxopwe_DO_reg[12]/P0001  & n14829 ;
  assign n16754 = ~n16752 & ~n16753 ;
  assign n16755 = ~n16750 & n16754 ;
  assign n16756 = ~n16751 & n16755 ;
  assign n16757 = ~n16749 & ~n16756 ;
  assign n16758 = ~n14779 & ~n16748 ;
  assign n16759 = ~n16757 & ~n16758 ;
  assign n16760 = ~n16402 & ~n16411 ;
  assign n16761 = n16409 & ~n16760 ;
  assign n16762 = ~n16409 & n16760 ;
  assign n16763 = ~n16761 & ~n16762 ;
  assign n16764 = n16759 & ~n16763 ;
  assign n16765 = ~n14852 & ~n16764 ;
  assign n16766 = ~n16412 & n16415 ;
  assign n16767 = ~n16416 & ~n16766 ;
  assign n16768 = ~n14852 & n16767 ;
  assign n16769 = n14852 & ~n16767 ;
  assign n16770 = ~n16768 & ~n16769 ;
  assign n16771 = ~n16765 & n16770 ;
  assign n16772 = ~n16766 & ~n16770 ;
  assign n16773 = ~n16771 & ~n16772 ;
  assign n16774 = n16741 & ~n16773 ;
  assign n16775 = n16641 & ~n16648 ;
  assign n16776 = ~n16649 & ~n16775 ;
  assign n16777 = ~\core_eu_em_mac_em_reg_mxopwe_DO_reg[3]/P0001  & ~n14967 ;
  assign n16778 = \core_eu_em_mac_em_reg_mxopwe_DO_reg[3]/P0001  & ~n14969 ;
  assign n16779 = ~n16777 & ~n16778 ;
  assign n16781 = \core_eu_em_mac_em_reg_mxopwe_DO_reg[5]/P0001  & ~n14951 ;
  assign n16780 = ~\core_eu_em_mac_em_reg_mxopwe_DO_reg[5]/P0001  & ~n14947 ;
  assign n16782 = ~\core_eu_em_mac_em_reg_mxopwe_DO_reg[4]/P0001  & n14958 ;
  assign n16783 = \core_eu_em_mac_em_reg_mxopwe_DO_reg[4]/P0001  & n14962 ;
  assign n16784 = ~n16782 & ~n16783 ;
  assign n16785 = ~n16780 & n16784 ;
  assign n16786 = ~n16781 & n16785 ;
  assign n16787 = ~n16779 & n16786 ;
  assign n16788 = n16779 & ~n16786 ;
  assign n16791 = ~\core_c_psq_MSTAT_reg_DO_reg[4]/NET0131  & ~n16591 ;
  assign n16789 = \core_c_dec_MACop_E_reg/P0001  & ~n7885 ;
  assign n16790 = \core_c_psq_MSTAT_reg_DO_reg[4]/NET0131  & ~n16789 ;
  assign n16792 = ~\core_eu_em_mac_em_dec_emcorepi_DO_reg[1]/P0001  & ~n16790 ;
  assign n16793 = ~n16791 & n16792 ;
  assign n16794 = ~n16788 & ~n16793 ;
  assign n16795 = ~n16787 & ~n16794 ;
  assign n16796 = ~n16603 & ~n16604 ;
  assign n16797 = ~n16607 & n16796 ;
  assign n16798 = n16607 & ~n16796 ;
  assign n16799 = ~n16797 & ~n16798 ;
  assign n16800 = ~n16795 & ~n16799 ;
  assign n16802 = \core_eu_em_mac_em_reg_mxopwe_DO_reg[11]/P0001  & ~n14865 ;
  assign n16801 = ~\core_eu_em_mac_em_reg_mxopwe_DO_reg[11]/P0001  & ~n14861 ;
  assign n16803 = ~\core_eu_em_mac_em_reg_mxopwe_DO_reg[10]/P0001  & n14872 ;
  assign n16804 = \core_eu_em_mac_em_reg_mxopwe_DO_reg[10]/P0001  & n14876 ;
  assign n16805 = ~n16803 & ~n16804 ;
  assign n16806 = ~n16801 & n16805 ;
  assign n16807 = ~n16802 & n16806 ;
  assign n16809 = \core_eu_em_mac_em_reg_mxopwe_DO_reg[9]/P0001  & ~n14891 ;
  assign n16808 = ~\core_eu_em_mac_em_reg_mxopwe_DO_reg[9]/P0001  & ~n14887 ;
  assign n16810 = ~\core_eu_em_mac_em_reg_mxopwe_DO_reg[8]/P0001  & n14898 ;
  assign n16811 = \core_eu_em_mac_em_reg_mxopwe_DO_reg[8]/P0001  & n14902 ;
  assign n16812 = ~n16810 & ~n16811 ;
  assign n16813 = ~n16808 & n16812 ;
  assign n16814 = ~n16809 & n16813 ;
  assign n16815 = n16807 & n16814 ;
  assign n16817 = \core_eu_em_mac_em_reg_mxopwe_DO_reg[7]/P0001  & ~n14918 ;
  assign n16816 = ~\core_eu_em_mac_em_reg_mxopwe_DO_reg[7]/P0001  & ~n14914 ;
  assign n16818 = ~\core_eu_em_mac_em_reg_mxopwe_DO_reg[6]/P0001  & n14925 ;
  assign n16819 = \core_eu_em_mac_em_reg_mxopwe_DO_reg[6]/P0001  & n14929 ;
  assign n16820 = ~n16818 & ~n16819 ;
  assign n16821 = ~n16816 & n16820 ;
  assign n16822 = ~n16817 & n16821 ;
  assign n16823 = ~n16815 & ~n16822 ;
  assign n16824 = ~n16807 & ~n16814 ;
  assign n16825 = ~n16823 & ~n16824 ;
  assign n16826 = ~n16625 & ~n16634 ;
  assign n16827 = n16632 & ~n16826 ;
  assign n16828 = ~n16632 & n16826 ;
  assign n16829 = ~n16827 & ~n16828 ;
  assign n16830 = n16825 & ~n16829 ;
  assign n16831 = ~n16800 & ~n16830 ;
  assign n16832 = ~n16635 & n16639 ;
  assign n16833 = ~n16640 & ~n16832 ;
  assign n16834 = ~n16590 & ~n16609 ;
  assign n16835 = ~n16610 & ~n16834 ;
  assign n16836 = n16833 & ~n16835 ;
  assign n16837 = ~n16833 & n16835 ;
  assign n16838 = ~n16836 & ~n16837 ;
  assign n16839 = ~n16831 & ~n16838 ;
  assign n16840 = ~n16832 & ~n16834 ;
  assign n16841 = n16838 & n16840 ;
  assign n16842 = ~n16839 & ~n16841 ;
  assign n16843 = n16776 & ~n16842 ;
  assign n16844 = ~n16774 & ~n16843 ;
  assign n16845 = ~n16397 & n16425 ;
  assign n16846 = ~n16426 & ~n16845 ;
  assign n16847 = ~n16586 & n16652 ;
  assign n16848 = ~n16653 & ~n16847 ;
  assign n16849 = n16846 & n16848 ;
  assign n16850 = ~n16846 & ~n16848 ;
  assign n16851 = ~n16849 & ~n16850 ;
  assign n16852 = n16844 & n16851 ;
  assign n16853 = ~n16845 & ~n16847 ;
  assign n16854 = ~n16851 & ~n16853 ;
  assign n16855 = ~n16852 & ~n16854 ;
  assign n16856 = n16739 & n16855 ;
  assign n16857 = ~n16844 & ~n16851 ;
  assign n16858 = ~n16852 & ~n16857 ;
  assign n16859 = n16831 & n16838 ;
  assign n16860 = ~n16839 & ~n16859 ;
  assign n16862 = \core_eu_em_mac_em_reg_mxopwe_DO_reg[10]/P0001  & ~n14865 ;
  assign n16861 = ~\core_eu_em_mac_em_reg_mxopwe_DO_reg[10]/P0001  & ~n14861 ;
  assign n16863 = ~\core_eu_em_mac_em_reg_mxopwe_DO_reg[9]/P0001  & n14872 ;
  assign n16864 = \core_eu_em_mac_em_reg_mxopwe_DO_reg[9]/P0001  & n14876 ;
  assign n16865 = ~n16863 & ~n16864 ;
  assign n16866 = ~n16861 & n16865 ;
  assign n16867 = ~n16862 & n16866 ;
  assign n16869 = \core_eu_em_mac_em_reg_mxopwe_DO_reg[8]/P0001  & ~n14891 ;
  assign n16868 = ~\core_eu_em_mac_em_reg_mxopwe_DO_reg[8]/P0001  & ~n14887 ;
  assign n16870 = ~\core_eu_em_mac_em_reg_mxopwe_DO_reg[7]/P0001  & n14898 ;
  assign n16871 = \core_eu_em_mac_em_reg_mxopwe_DO_reg[7]/P0001  & n14902 ;
  assign n16872 = ~n16870 & ~n16871 ;
  assign n16873 = ~n16868 & n16872 ;
  assign n16874 = ~n16869 & n16873 ;
  assign n16875 = n16867 & n16874 ;
  assign n16877 = \core_eu_em_mac_em_reg_mxopwe_DO_reg[6]/P0001  & ~n14918 ;
  assign n16876 = ~\core_eu_em_mac_em_reg_mxopwe_DO_reg[6]/P0001  & ~n14914 ;
  assign n16878 = ~\core_eu_em_mac_em_reg_mxopwe_DO_reg[5]/P0001  & n14925 ;
  assign n16879 = \core_eu_em_mac_em_reg_mxopwe_DO_reg[5]/P0001  & n14929 ;
  assign n16880 = ~n16878 & ~n16879 ;
  assign n16881 = ~n16876 & n16880 ;
  assign n16882 = ~n16877 & n16881 ;
  assign n16883 = ~n16875 & ~n16882 ;
  assign n16884 = ~n16867 & ~n16874 ;
  assign n16885 = ~n16883 & ~n16884 ;
  assign n16886 = ~n16815 & ~n16824 ;
  assign n16887 = n16822 & ~n16886 ;
  assign n16888 = ~n16822 & n16886 ;
  assign n16889 = ~n16887 & ~n16888 ;
  assign n16890 = n16885 & ~n16889 ;
  assign n16891 = ~n16787 & ~n16788 ;
  assign n16892 = n16793 & ~n16891 ;
  assign n16893 = ~n16793 & n16891 ;
  assign n16894 = ~n16892 & ~n16893 ;
  assign n16897 = ~\core_c_psq_MSTAT_reg_DO_reg[4]/NET0131  & ~n16789 ;
  assign n16895 = \core_c_dec_MACop_E_reg/P0001  & ~n8558 ;
  assign n16896 = \core_c_psq_MSTAT_reg_DO_reg[4]/NET0131  & ~n16895 ;
  assign n16898 = ~\core_eu_em_mac_em_dec_emcorepi_DO_reg[1]/P0001  & ~n16896 ;
  assign n16899 = ~n16897 & n16898 ;
  assign n16901 = \core_eu_em_mac_em_reg_mxopwe_DO_reg[4]/P0001  & ~n14951 ;
  assign n16900 = ~\core_eu_em_mac_em_reg_mxopwe_DO_reg[4]/P0001  & ~n14947 ;
  assign n16902 = ~\core_eu_em_mac_em_reg_mxopwe_DO_reg[3]/P0001  & n14958 ;
  assign n16903 = \core_eu_em_mac_em_reg_mxopwe_DO_reg[3]/P0001  & n14962 ;
  assign n16904 = ~n16902 & ~n16903 ;
  assign n16905 = ~n16900 & n16904 ;
  assign n16906 = ~n16901 & n16905 ;
  assign n16907 = n16899 & ~n16906 ;
  assign n16908 = ~n16899 & n16906 ;
  assign n16909 = ~\core_eu_em_mac_em_reg_mxopwe_DO_reg[2]/P0001  & n14967 ;
  assign n16910 = \core_eu_em_mac_em_reg_mxopwe_DO_reg[2]/P0001  & n14969 ;
  assign n16911 = ~n16909 & ~n16910 ;
  assign n16912 = ~n16908 & ~n16911 ;
  assign n16913 = ~n16907 & ~n16912 ;
  assign n16914 = n16894 & n16913 ;
  assign n16915 = ~n16890 & ~n16914 ;
  assign n16916 = ~n16825 & n16829 ;
  assign n16917 = ~n16830 & ~n16916 ;
  assign n16918 = n16795 & n16799 ;
  assign n16919 = ~n16800 & ~n16918 ;
  assign n16920 = n16917 & ~n16919 ;
  assign n16921 = ~n16917 & n16919 ;
  assign n16922 = ~n16920 & ~n16921 ;
  assign n16923 = n16915 & ~n16922 ;
  assign n16924 = ~n16916 & ~n16918 ;
  assign n16925 = n16922 & ~n16924 ;
  assign n16926 = ~n16923 & ~n16925 ;
  assign n16927 = n16860 & n16926 ;
  assign n16929 = \core_eu_em_mac_em_reg_mxopwe_DO_reg[12]/P0001  & ~n14818 ;
  assign n16928 = ~\core_eu_em_mac_em_reg_mxopwe_DO_reg[12]/P0001  & ~n14814 ;
  assign n16930 = ~\core_eu_em_mac_em_reg_mxopwe_DO_reg[11]/P0001  & n14825 ;
  assign n16931 = \core_eu_em_mac_em_reg_mxopwe_DO_reg[11]/P0001  & n14829 ;
  assign n16932 = ~n16930 & ~n16931 ;
  assign n16933 = ~n16928 & n16932 ;
  assign n16934 = ~n16929 & n16933 ;
  assign n16936 = \core_eu_em_mac_em_reg_mxopwe_DO_reg[14]/P0001  & ~n14791 ;
  assign n16935 = ~\core_eu_em_mac_em_reg_mxopwe_DO_reg[14]/P0001  & ~n14787 ;
  assign n16937 = ~\core_eu_em_mac_em_reg_mxopwe_DO_reg[13]/P0001  & n14798 ;
  assign n16938 = \core_eu_em_mac_em_reg_mxopwe_DO_reg[13]/P0001  & n14802 ;
  assign n16939 = ~n16937 & ~n16938 ;
  assign n16940 = ~n16935 & n16939 ;
  assign n16941 = ~n16936 & n16940 ;
  assign n16942 = n16934 & n16941 ;
  assign n16943 = ~\core_eu_em_mac_em_reg_mxopwe_DO_reg[15]/P0001  & n14772 ;
  assign n16944 = \core_eu_em_mac_em_reg_mxopwe_DO_reg[15]/P0001  & n14776 ;
  assign n16945 = ~n16943 & ~n16944 ;
  assign n16946 = n14767 & n16945 ;
  assign n16947 = ~n16942 & ~n16946 ;
  assign n16948 = ~n16934 & ~n16941 ;
  assign n16949 = ~n16947 & ~n16948 ;
  assign n16950 = ~n16749 & ~n16758 ;
  assign n16951 = n16756 & ~n16950 ;
  assign n16952 = ~n16756 & n16950 ;
  assign n16953 = ~n16951 & ~n16952 ;
  assign n16954 = n16949 & ~n16953 ;
  assign n16955 = ~n14852 & ~n16954 ;
  assign n16956 = ~n16759 & n16763 ;
  assign n16957 = ~n16764 & ~n16956 ;
  assign n16958 = n14852 & ~n16957 ;
  assign n16959 = n16765 & ~n16956 ;
  assign n16960 = ~n16958 & ~n16959 ;
  assign n16961 = ~n16955 & n16960 ;
  assign n16962 = ~n16956 & ~n16960 ;
  assign n16963 = ~n16961 & ~n16962 ;
  assign n16964 = ~n16764 & n16768 ;
  assign n16965 = ~n16771 & ~n16964 ;
  assign n16966 = ~n16963 & n16965 ;
  assign n16967 = ~n16927 & ~n16966 ;
  assign n16968 = ~n16741 & n16773 ;
  assign n16969 = ~n16774 & ~n16968 ;
  assign n16970 = ~n16776 & n16842 ;
  assign n16971 = ~n16843 & ~n16970 ;
  assign n16972 = n16969 & n16971 ;
  assign n16973 = ~n16969 & ~n16971 ;
  assign n16974 = ~n16972 & ~n16973 ;
  assign n16975 = ~n16967 & n16974 ;
  assign n16976 = ~n16968 & ~n16970 ;
  assign n16977 = ~n16974 & n16976 ;
  assign n16978 = ~n16975 & ~n16977 ;
  assign n16979 = ~n16858 & ~n16978 ;
  assign n16980 = ~n16856 & ~n16979 ;
  assign n16981 = ~n16683 & ~n16709 ;
  assign n16982 = ~n16669 & ~n16678 ;
  assign n16983 = ~n16670 & ~n16982 ;
  assign n16985 = \core_eu_em_mac_em_reg_mxopwe_DO_reg[13]/P0001  & ~n14918 ;
  assign n16984 = ~\core_eu_em_mac_em_reg_mxopwe_DO_reg[13]/P0001  & ~n14914 ;
  assign n16986 = ~\core_eu_em_mac_em_reg_mxopwe_DO_reg[12]/P0001  & n14925 ;
  assign n16987 = \core_eu_em_mac_em_reg_mxopwe_DO_reg[12]/P0001  & n14929 ;
  assign n16988 = ~n16986 & ~n16987 ;
  assign n16989 = ~n16984 & n16988 ;
  assign n16990 = ~n16985 & n16989 ;
  assign n16991 = n14879 & n16990 ;
  assign n16992 = ~n14879 & ~n16990 ;
  assign n16993 = ~n16991 & ~n16992 ;
  assign n16995 = ~\core_eu_em_mac_em_reg_mxopwe_DO_reg[15]/P0001  & ~n14887 ;
  assign n16994 = \core_eu_em_mac_em_reg_mxopwe_DO_reg[15]/P0001  & ~n14891 ;
  assign n16996 = ~\core_eu_em_mac_em_reg_mxopwe_DO_reg[14]/P0001  & n14898 ;
  assign n16997 = \core_eu_em_mac_em_reg_mxopwe_DO_reg[14]/P0001  & n14902 ;
  assign n16998 = ~n16996 & ~n16997 ;
  assign n16999 = ~n16994 & n16998 ;
  assign n17000 = ~n16995 & n16999 ;
  assign n17001 = ~n16993 & n17000 ;
  assign n17002 = n16993 & ~n17000 ;
  assign n17003 = ~n17001 & ~n17002 ;
  assign n17004 = n16983 & ~n17003 ;
  assign n17005 = ~n16983 & n17003 ;
  assign n17006 = ~n17004 & ~n17005 ;
  assign n17007 = ~\core_eu_em_mac_em_reg_mxopwe_DO_reg[9]/P0001  & ~n14967 ;
  assign n17008 = \core_eu_em_mac_em_reg_mxopwe_DO_reg[9]/P0001  & ~n14969 ;
  assign n17009 = ~n17007 & ~n17008 ;
  assign n17011 = \core_eu_em_mac_em_reg_mxopwe_DO_reg[11]/P0001  & ~n14951 ;
  assign n17010 = ~\core_eu_em_mac_em_reg_mxopwe_DO_reg[11]/P0001  & ~n14947 ;
  assign n17012 = ~\core_eu_em_mac_em_reg_mxopwe_DO_reg[10]/P0001  & n14958 ;
  assign n17013 = \core_eu_em_mac_em_reg_mxopwe_DO_reg[10]/P0001  & n14962 ;
  assign n17014 = ~n17012 & ~n17013 ;
  assign n17015 = ~n17010 & n17014 ;
  assign n17016 = ~n17011 & n17015 ;
  assign n17017 = n17009 & ~n17016 ;
  assign n17018 = ~n17009 & n17016 ;
  assign n17019 = ~n17017 & ~n17018 ;
  assign n17021 = ~\core_c_psq_MSTAT_reg_DO_reg[4]/NET0131  & ~n15254 ;
  assign n17020 = \core_c_psq_MSTAT_reg_DO_reg[4]/NET0131  & ~n16699 ;
  assign n17022 = ~\core_eu_em_mac_em_dec_emcorepi_DO_reg[1]/P0001  & ~n17020 ;
  assign n17023 = ~n17021 & n17022 ;
  assign n17024 = ~n17019 & n17023 ;
  assign n17025 = n17019 & ~n17023 ;
  assign n17026 = ~n17024 & ~n17025 ;
  assign n17027 = ~n16696 & ~n16702 ;
  assign n17028 = ~n16695 & ~n17027 ;
  assign n17029 = n17026 & ~n17028 ;
  assign n17030 = ~n17026 & n17028 ;
  assign n17031 = ~n17029 & ~n17030 ;
  assign n17032 = n17006 & n17031 ;
  assign n17033 = ~n17006 & ~n17031 ;
  assign n17034 = ~n17032 & ~n17033 ;
  assign n17035 = ~n16981 & n17034 ;
  assign n17036 = n16981 & ~n17034 ;
  assign n17037 = ~n17035 & ~n17036 ;
  assign n17038 = ~n16682 & ~n16708 ;
  assign n17039 = ~n16713 & n17038 ;
  assign n17040 = ~n16714 & ~n17039 ;
  assign n17041 = n17037 & ~n17040 ;
  assign n17042 = ~n14853 & ~n17041 ;
  assign n17043 = ~n17004 & ~n17029 ;
  assign n17044 = ~n16991 & ~n17000 ;
  assign n17045 = ~n16992 & ~n17044 ;
  assign n17046 = ~n15281 & ~n15287 ;
  assign n17047 = n15285 & ~n17046 ;
  assign n17048 = ~n15285 & n17046 ;
  assign n17049 = ~n17047 & ~n17048 ;
  assign n17050 = ~n17045 & n17049 ;
  assign n17051 = n17045 & ~n17049 ;
  assign n17052 = ~n17050 & ~n17051 ;
  assign n17053 = ~n15266 & ~n15267 ;
  assign n17054 = ~n15270 & n17053 ;
  assign n17055 = n15270 & ~n17053 ;
  assign n17056 = ~n17054 & ~n17055 ;
  assign n17057 = ~n17018 & n17023 ;
  assign n17058 = ~n17017 & ~n17057 ;
  assign n17059 = n17056 & ~n17058 ;
  assign n17060 = ~n17056 & n17058 ;
  assign n17061 = ~n17059 & ~n17060 ;
  assign n17062 = n17052 & n17061 ;
  assign n17063 = ~n17052 & ~n17061 ;
  assign n17064 = ~n17062 & ~n17063 ;
  assign n17065 = n17043 & ~n17064 ;
  assign n17066 = ~n17043 & n17064 ;
  assign n17067 = ~n17065 & ~n17066 ;
  assign n17068 = ~n17005 & ~n17030 ;
  assign n17069 = ~n17034 & n17068 ;
  assign n17070 = ~n17035 & ~n17069 ;
  assign n17071 = n17067 & ~n17070 ;
  assign n17072 = ~n17067 & n17070 ;
  assign n17073 = ~n17071 & ~n17072 ;
  assign n17074 = n14853 & n17073 ;
  assign n17075 = ~n14853 & ~n17073 ;
  assign n17076 = ~n17074 & ~n17075 ;
  assign n17077 = ~n17042 & ~n17076 ;
  assign n17078 = n17042 & n17073 ;
  assign n17079 = ~n17077 & ~n17078 ;
  assign n17080 = ~n16721 & ~n16732 ;
  assign n17081 = ~n17037 & n17040 ;
  assign n17082 = ~n17041 & ~n17081 ;
  assign n17083 = n14853 & n17082 ;
  assign n17084 = ~n14853 & ~n17082 ;
  assign n17085 = ~n17083 & ~n17084 ;
  assign n17086 = ~n17080 & ~n17085 ;
  assign n17087 = n17080 & n17085 ;
  assign n17088 = ~n17086 & ~n17087 ;
  assign n17089 = ~n16720 & ~n16731 ;
  assign n17090 = ~n16736 & n17089 ;
  assign n17091 = ~n16737 & ~n17090 ;
  assign n17092 = n17088 & ~n17091 ;
  assign n17093 = ~n17079 & ~n17092 ;
  assign n17094 = ~n17081 & n17085 ;
  assign n17095 = ~n17086 & ~n17094 ;
  assign n17096 = n17091 & n17095 ;
  assign n17097 = ~n17093 & ~n17096 ;
  assign n17098 = n16980 & ~n17097 ;
  assign n17100 = \core_eu_em_mac_em_reg_mxopwe_DO_reg[13]/P0001  & ~n14791 ;
  assign n17099 = ~\core_eu_em_mac_em_reg_mxopwe_DO_reg[13]/P0001  & ~n14787 ;
  assign n17101 = ~\core_eu_em_mac_em_reg_mxopwe_DO_reg[12]/P0001  & n14798 ;
  assign n17102 = \core_eu_em_mac_em_reg_mxopwe_DO_reg[12]/P0001  & n14802 ;
  assign n17103 = ~n17101 & ~n17102 ;
  assign n17104 = ~n17099 & n17103 ;
  assign n17105 = ~n17100 & n17104 ;
  assign n17107 = \core_eu_em_mac_em_reg_mxopwe_DO_reg[15]/P0001  & ~n14765 ;
  assign n17106 = ~\core_eu_em_mac_em_reg_mxopwe_DO_reg[15]/P0001  & ~n14761 ;
  assign n17108 = ~\core_eu_em_mac_em_reg_mxopwe_DO_reg[14]/P0001  & n14772 ;
  assign n17109 = \core_eu_em_mac_em_reg_mxopwe_DO_reg[14]/P0001  & n14776 ;
  assign n17110 = ~n17108 & ~n17109 ;
  assign n17111 = ~n17106 & n17110 ;
  assign n17112 = ~n17107 & n17111 ;
  assign n17113 = n17105 & n17112 ;
  assign n17115 = \core_eu_em_mac_em_reg_mxopwe_DO_reg[11]/P0001  & ~n14818 ;
  assign n17114 = ~\core_eu_em_mac_em_reg_mxopwe_DO_reg[11]/P0001  & ~n14814 ;
  assign n17116 = ~\core_eu_em_mac_em_reg_mxopwe_DO_reg[10]/P0001  & n14825 ;
  assign n17117 = \core_eu_em_mac_em_reg_mxopwe_DO_reg[10]/P0001  & n14829 ;
  assign n17118 = ~n17116 & ~n17117 ;
  assign n17119 = ~n17114 & n17118 ;
  assign n17120 = ~n17115 & n17119 ;
  assign n17121 = ~n17113 & ~n17120 ;
  assign n17122 = ~n17105 & ~n17112 ;
  assign n17123 = ~n17121 & ~n17122 ;
  assign n17124 = ~n16942 & ~n16948 ;
  assign n17125 = n16946 & ~n17124 ;
  assign n17126 = ~n16946 & n17124 ;
  assign n17127 = ~n17125 & ~n17126 ;
  assign n17128 = n17123 & ~n17127 ;
  assign n17129 = ~n14852 & ~n17128 ;
  assign n17130 = ~n16949 & n16953 ;
  assign n17131 = ~n16954 & ~n17130 ;
  assign n17132 = ~n14852 & n17131 ;
  assign n17133 = n14852 & ~n17131 ;
  assign n17134 = ~n17132 & ~n17133 ;
  assign n17135 = ~n17129 & n17134 ;
  assign n17136 = ~n17128 & n17132 ;
  assign n17137 = ~n17135 & ~n17136 ;
  assign n17139 = \core_eu_em_mac_em_reg_mxopwe_DO_reg[12]/P0001  & ~n14791 ;
  assign n17138 = ~\core_eu_em_mac_em_reg_mxopwe_DO_reg[12]/P0001  & ~n14787 ;
  assign n17140 = ~\core_eu_em_mac_em_reg_mxopwe_DO_reg[11]/P0001  & n14798 ;
  assign n17141 = \core_eu_em_mac_em_reg_mxopwe_DO_reg[11]/P0001  & n14802 ;
  assign n17142 = ~n17140 & ~n17141 ;
  assign n17143 = ~n17138 & n17142 ;
  assign n17144 = ~n17139 & n17143 ;
  assign n17146 = \core_eu_em_mac_em_reg_mxopwe_DO_reg[14]/P0001  & ~n14765 ;
  assign n17145 = ~\core_eu_em_mac_em_reg_mxopwe_DO_reg[14]/P0001  & ~n14761 ;
  assign n17147 = ~\core_eu_em_mac_em_reg_mxopwe_DO_reg[13]/P0001  & n14772 ;
  assign n17148 = \core_eu_em_mac_em_reg_mxopwe_DO_reg[13]/P0001  & n14776 ;
  assign n17149 = ~n17147 & ~n17148 ;
  assign n17150 = ~n17145 & n17149 ;
  assign n17151 = ~n17146 & n17150 ;
  assign n17152 = n17144 & n17151 ;
  assign n17154 = \core_eu_em_mac_em_reg_mxopwe_DO_reg[10]/P0001  & ~n14818 ;
  assign n17153 = ~\core_eu_em_mac_em_reg_mxopwe_DO_reg[10]/P0001  & ~n14814 ;
  assign n17155 = ~\core_eu_em_mac_em_reg_mxopwe_DO_reg[9]/P0001  & n14825 ;
  assign n17156 = \core_eu_em_mac_em_reg_mxopwe_DO_reg[9]/P0001  & n14829 ;
  assign n17157 = ~n17155 & ~n17156 ;
  assign n17158 = ~n17153 & n17157 ;
  assign n17159 = ~n17154 & n17158 ;
  assign n17160 = ~n17152 & ~n17159 ;
  assign n17161 = ~n17144 & ~n17151 ;
  assign n17162 = ~n17160 & ~n17161 ;
  assign n17163 = ~n17113 & ~n17122 ;
  assign n17164 = n17120 & ~n17163 ;
  assign n17165 = ~n17120 & n17163 ;
  assign n17166 = ~n17164 & ~n17165 ;
  assign n17167 = n17162 & ~n17166 ;
  assign n17168 = ~\core_eu_em_mac_em_reg_mxopwe_DO_reg[15]/P0001  & n14846 ;
  assign n17169 = \core_eu_em_mac_em_reg_mxopwe_DO_reg[15]/P0001  & n14849 ;
  assign n17170 = ~n17168 & ~n17169 ;
  assign n17171 = n14844 & n17170 ;
  assign n17172 = n14967 & ~n17171 ;
  assign n17173 = n14852 & ~n17172 ;
  assign n17174 = ~n17167 & ~n17173 ;
  assign n17175 = ~n17123 & n17127 ;
  assign n17176 = ~n17128 & ~n17175 ;
  assign n17177 = n14852 & ~n17176 ;
  assign n17178 = ~n14852 & n17176 ;
  assign n17179 = ~n17177 & ~n17178 ;
  assign n17180 = n17174 & n17179 ;
  assign n17181 = n14852 & n17175 ;
  assign n17182 = ~n17180 & ~n17181 ;
  assign n17183 = n17137 & n17182 ;
  assign n17185 = \core_eu_em_mac_em_reg_mxopwe_DO_reg[9]/P0001  & ~n14865 ;
  assign n17184 = ~\core_eu_em_mac_em_reg_mxopwe_DO_reg[9]/P0001  & ~n14861 ;
  assign n17186 = ~\core_eu_em_mac_em_reg_mxopwe_DO_reg[8]/P0001  & n14872 ;
  assign n17187 = \core_eu_em_mac_em_reg_mxopwe_DO_reg[8]/P0001  & n14876 ;
  assign n17188 = ~n17186 & ~n17187 ;
  assign n17189 = ~n17184 & n17188 ;
  assign n17190 = ~n17185 & n17189 ;
  assign n17192 = \core_eu_em_mac_em_reg_mxopwe_DO_reg[5]/P0001  & ~n14918 ;
  assign n17191 = ~\core_eu_em_mac_em_reg_mxopwe_DO_reg[5]/P0001  & ~n14914 ;
  assign n17193 = ~\core_eu_em_mac_em_reg_mxopwe_DO_reg[4]/P0001  & n14925 ;
  assign n17194 = \core_eu_em_mac_em_reg_mxopwe_DO_reg[4]/P0001  & n14929 ;
  assign n17195 = ~n17193 & ~n17194 ;
  assign n17196 = ~n17191 & n17195 ;
  assign n17197 = ~n17192 & n17196 ;
  assign n17198 = n17190 & n17197 ;
  assign n17200 = \core_eu_em_mac_em_reg_mxopwe_DO_reg[7]/P0001  & ~n14891 ;
  assign n17199 = ~\core_eu_em_mac_em_reg_mxopwe_DO_reg[7]/P0001  & ~n14887 ;
  assign n17201 = ~\core_eu_em_mac_em_reg_mxopwe_DO_reg[6]/P0001  & n14898 ;
  assign n17202 = \core_eu_em_mac_em_reg_mxopwe_DO_reg[6]/P0001  & n14902 ;
  assign n17203 = ~n17201 & ~n17202 ;
  assign n17204 = ~n17199 & n17203 ;
  assign n17205 = ~n17200 & n17204 ;
  assign n17206 = ~n17198 & ~n17205 ;
  assign n17207 = ~n17190 & ~n17197 ;
  assign n17208 = ~n17206 & ~n17207 ;
  assign n17209 = ~n16875 & ~n16884 ;
  assign n17210 = n16882 & ~n17209 ;
  assign n17211 = ~n16882 & n17209 ;
  assign n17212 = ~n17210 & ~n17211 ;
  assign n17213 = n17208 & ~n17212 ;
  assign n17214 = ~n16907 & ~n16908 ;
  assign n17215 = ~n16911 & n17214 ;
  assign n17216 = n16911 & ~n17214 ;
  assign n17217 = ~n17215 & ~n17216 ;
  assign n17220 = ~\core_c_psq_MSTAT_reg_DO_reg[4]/NET0131  & ~n16895 ;
  assign n17218 = \core_c_dec_MACop_E_reg/P0001  & ~n9205 ;
  assign n17219 = \core_c_psq_MSTAT_reg_DO_reg[4]/NET0131  & ~n17218 ;
  assign n17221 = ~\core_eu_em_mac_em_dec_emcorepi_DO_reg[1]/P0001  & ~n17219 ;
  assign n17222 = ~n17220 & n17221 ;
  assign n17224 = \core_eu_em_mac_em_reg_mxopwe_DO_reg[3]/P0001  & ~n14951 ;
  assign n17223 = ~\core_eu_em_mac_em_reg_mxopwe_DO_reg[3]/P0001  & ~n14947 ;
  assign n17225 = ~\core_eu_em_mac_em_reg_mxopwe_DO_reg[2]/P0001  & n14958 ;
  assign n17226 = \core_eu_em_mac_em_reg_mxopwe_DO_reg[2]/P0001  & n14962 ;
  assign n17227 = ~n17225 & ~n17226 ;
  assign n17228 = ~n17223 & n17227 ;
  assign n17229 = ~n17224 & n17228 ;
  assign n17230 = n17222 & ~n17229 ;
  assign n17231 = ~n17222 & n17229 ;
  assign n17232 = ~\core_eu_em_mac_em_reg_mxopwe_DO_reg[1]/P0001  & n14967 ;
  assign n17233 = \core_eu_em_mac_em_reg_mxopwe_DO_reg[1]/P0001  & n14969 ;
  assign n17234 = ~n17232 & ~n17233 ;
  assign n17235 = ~n17231 & ~n17234 ;
  assign n17236 = ~n17230 & ~n17235 ;
  assign n17237 = ~n17217 & n17236 ;
  assign n17238 = ~n17213 & ~n17237 ;
  assign n17239 = ~n16885 & n16889 ;
  assign n17240 = ~n16890 & ~n17239 ;
  assign n17241 = ~n16894 & ~n16913 ;
  assign n17242 = ~n16914 & ~n17241 ;
  assign n17243 = n17240 & n17242 ;
  assign n17244 = ~n17240 & ~n17242 ;
  assign n17245 = ~n17243 & ~n17244 ;
  assign n17246 = ~n17238 & n17245 ;
  assign n17247 = n17238 & ~n17245 ;
  assign n17248 = ~n17246 & ~n17247 ;
  assign n17250 = \core_eu_em_mac_em_reg_mxopwe_DO_reg[6]/P0001  & ~n14891 ;
  assign n17249 = ~\core_eu_em_mac_em_reg_mxopwe_DO_reg[6]/P0001  & ~n14887 ;
  assign n17251 = ~\core_eu_em_mac_em_reg_mxopwe_DO_reg[5]/P0001  & n14898 ;
  assign n17252 = \core_eu_em_mac_em_reg_mxopwe_DO_reg[5]/P0001  & n14902 ;
  assign n17253 = ~n17251 & ~n17252 ;
  assign n17254 = ~n17249 & n17253 ;
  assign n17255 = ~n17250 & n17254 ;
  assign n17257 = \core_eu_em_mac_em_reg_mxopwe_DO_reg[8]/P0001  & ~n14865 ;
  assign n17256 = ~\core_eu_em_mac_em_reg_mxopwe_DO_reg[8]/P0001  & ~n14861 ;
  assign n17258 = ~\core_eu_em_mac_em_reg_mxopwe_DO_reg[7]/P0001  & n14872 ;
  assign n17259 = \core_eu_em_mac_em_reg_mxopwe_DO_reg[7]/P0001  & n14876 ;
  assign n17260 = ~n17258 & ~n17259 ;
  assign n17261 = ~n17256 & n17260 ;
  assign n17262 = ~n17257 & n17261 ;
  assign n17263 = n17255 & n17262 ;
  assign n17265 = \core_eu_em_mac_em_reg_mxopwe_DO_reg[4]/P0001  & ~n14918 ;
  assign n17264 = ~\core_eu_em_mac_em_reg_mxopwe_DO_reg[4]/P0001  & ~n14914 ;
  assign n17266 = ~\core_eu_em_mac_em_reg_mxopwe_DO_reg[3]/P0001  & n14925 ;
  assign n17267 = \core_eu_em_mac_em_reg_mxopwe_DO_reg[3]/P0001  & n14929 ;
  assign n17268 = ~n17266 & ~n17267 ;
  assign n17269 = ~n17264 & n17268 ;
  assign n17270 = ~n17265 & n17269 ;
  assign n17271 = ~n17263 & ~n17270 ;
  assign n17272 = ~n17255 & ~n17262 ;
  assign n17273 = ~n17271 & ~n17272 ;
  assign n17274 = ~n17198 & ~n17207 ;
  assign n17275 = n17205 & ~n17274 ;
  assign n17276 = ~n17205 & n17274 ;
  assign n17277 = ~n17275 & ~n17276 ;
  assign n17278 = n17273 & ~n17277 ;
  assign n17279 = ~n17230 & ~n17231 ;
  assign n17280 = ~n17234 & n17279 ;
  assign n17281 = n17234 & ~n17279 ;
  assign n17282 = ~n17280 & ~n17281 ;
  assign n17285 = ~\core_c_psq_MSTAT_reg_DO_reg[4]/NET0131  & ~n17218 ;
  assign n17283 = \core_c_dec_MACop_E_reg/P0001  & ~n7449 ;
  assign n17284 = \core_c_psq_MSTAT_reg_DO_reg[4]/NET0131  & ~n17283 ;
  assign n17286 = ~\core_eu_em_mac_em_dec_emcorepi_DO_reg[1]/P0001  & ~n17284 ;
  assign n17287 = ~n17285 & n17286 ;
  assign n17289 = \core_eu_em_mac_em_reg_mxopwe_DO_reg[2]/P0001  & ~n14951 ;
  assign n17288 = ~\core_eu_em_mac_em_reg_mxopwe_DO_reg[2]/P0001  & ~n14947 ;
  assign n17290 = ~\core_eu_em_mac_em_reg_mxopwe_DO_reg[1]/P0001  & n14958 ;
  assign n17291 = \core_eu_em_mac_em_reg_mxopwe_DO_reg[1]/P0001  & n14962 ;
  assign n17292 = ~n17290 & ~n17291 ;
  assign n17293 = ~n17288 & n17292 ;
  assign n17294 = ~n17289 & n17293 ;
  assign n17295 = n17287 & ~n17294 ;
  assign n17296 = ~n17287 & n17294 ;
  assign n17297 = ~\core_eu_em_mac_em_reg_mxopwe_DO_reg[0]/P0001  & n14967 ;
  assign n17298 = \core_eu_em_mac_em_reg_mxopwe_DO_reg[0]/P0001  & n14969 ;
  assign n17299 = ~n17297 & ~n17298 ;
  assign n17300 = ~n17296 & ~n17299 ;
  assign n17301 = ~n17295 & ~n17300 ;
  assign n17302 = ~n17282 & n17301 ;
  assign n17303 = ~n17278 & ~n17302 ;
  assign n17304 = ~n17208 & n17212 ;
  assign n17305 = ~n17213 & ~n17304 ;
  assign n17306 = n17217 & ~n17236 ;
  assign n17307 = ~n17237 & ~n17306 ;
  assign n17308 = n17305 & n17307 ;
  assign n17309 = ~n17305 & ~n17307 ;
  assign n17310 = ~n17308 & ~n17309 ;
  assign n17311 = ~n17303 & n17310 ;
  assign n17312 = ~n17304 & ~n17306 ;
  assign n17313 = ~n17310 & n17312 ;
  assign n17314 = ~n17311 & ~n17313 ;
  assign n17315 = n17248 & ~n17314 ;
  assign n17316 = ~n17183 & ~n17315 ;
  assign n17317 = ~n16915 & n16922 ;
  assign n17318 = ~n16923 & ~n17317 ;
  assign n17319 = ~n17239 & ~n17241 ;
  assign n17320 = ~n17245 & n17319 ;
  assign n17321 = ~n17246 & ~n17320 ;
  assign n17322 = ~n17318 & ~n17321 ;
  assign n17323 = n17318 & n17321 ;
  assign n17324 = ~n17322 & ~n17323 ;
  assign n17325 = n16955 & n16957 ;
  assign n17326 = ~n16961 & ~n17325 ;
  assign n17327 = ~n17130 & ~n17134 ;
  assign n17328 = ~n17135 & ~n17327 ;
  assign n17329 = ~n17326 & n17328 ;
  assign n17330 = n17326 & ~n17328 ;
  assign n17331 = ~n17329 & ~n17330 ;
  assign n17332 = n17324 & n17331 ;
  assign n17333 = ~n17324 & ~n17331 ;
  assign n17334 = ~n17332 & ~n17333 ;
  assign n17335 = ~n17316 & ~n17334 ;
  assign n17336 = n17316 & n17334 ;
  assign n17337 = ~n17335 & ~n17336 ;
  assign n17338 = n17303 & ~n17310 ;
  assign n17339 = ~n17311 & ~n17338 ;
  assign n17340 = \core_c_psq_MSTAT_reg_DO_reg[4]/NET0131  & \core_eu_em_mac_em_dec_emcorepi_DO_reg[0]/P0001  ;
  assign n17341 = ~\core_c_psq_MSTAT_reg_DO_reg[4]/NET0131  & ~\core_eu_em_mac_em_dec_emcorepi_DO_reg[1]/P0001  ;
  assign n17342 = n17283 & n17341 ;
  assign n17343 = ~n17340 & ~n17342 ;
  assign n17345 = ~\core_eu_em_mac_em_reg_mxopwe_DO_reg[1]/P0001  & ~n14947 ;
  assign n17344 = \core_eu_em_mac_em_reg_mxopwe_DO_reg[1]/P0001  & ~n14951 ;
  assign n17346 = ~\core_eu_em_mac_em_reg_mxopwe_DO_reg[0]/P0001  & n14958 ;
  assign n17347 = \core_eu_em_mac_em_reg_mxopwe_DO_reg[0]/P0001  & n14962 ;
  assign n17348 = ~n17346 & ~n17347 ;
  assign n17349 = ~n17344 & n17348 ;
  assign n17350 = ~n17345 & n17349 ;
  assign n17351 = ~n17343 & ~n17350 ;
  assign n17352 = ~n17295 & ~n17296 ;
  assign n17353 = ~n17299 & n17352 ;
  assign n17354 = n17299 & ~n17352 ;
  assign n17355 = ~n17353 & ~n17354 ;
  assign n17356 = ~n17351 & ~n17355 ;
  assign n17358 = \core_eu_em_mac_em_reg_mxopwe_DO_reg[5]/P0001  & ~n14891 ;
  assign n17357 = ~\core_eu_em_mac_em_reg_mxopwe_DO_reg[5]/P0001  & ~n14887 ;
  assign n17359 = ~\core_eu_em_mac_em_reg_mxopwe_DO_reg[4]/P0001  & n14898 ;
  assign n17360 = \core_eu_em_mac_em_reg_mxopwe_DO_reg[4]/P0001  & n14902 ;
  assign n17361 = ~n17359 & ~n17360 ;
  assign n17362 = ~n17357 & n17361 ;
  assign n17363 = ~n17358 & n17362 ;
  assign n17365 = \core_eu_em_mac_em_reg_mxopwe_DO_reg[7]/P0001  & ~n14865 ;
  assign n17364 = ~\core_eu_em_mac_em_reg_mxopwe_DO_reg[7]/P0001  & ~n14861 ;
  assign n17366 = ~\core_eu_em_mac_em_reg_mxopwe_DO_reg[6]/P0001  & n14872 ;
  assign n17367 = \core_eu_em_mac_em_reg_mxopwe_DO_reg[6]/P0001  & n14876 ;
  assign n17368 = ~n17366 & ~n17367 ;
  assign n17369 = ~n17364 & n17368 ;
  assign n17370 = ~n17365 & n17369 ;
  assign n17371 = n17363 & n17370 ;
  assign n17373 = \core_eu_em_mac_em_reg_mxopwe_DO_reg[3]/P0001  & ~n14918 ;
  assign n17372 = ~\core_eu_em_mac_em_reg_mxopwe_DO_reg[3]/P0001  & ~n14914 ;
  assign n17374 = ~\core_eu_em_mac_em_reg_mxopwe_DO_reg[2]/P0001  & n14925 ;
  assign n17375 = \core_eu_em_mac_em_reg_mxopwe_DO_reg[2]/P0001  & n14929 ;
  assign n17376 = ~n17374 & ~n17375 ;
  assign n17377 = ~n17372 & n17376 ;
  assign n17378 = ~n17373 & n17377 ;
  assign n17379 = ~n17371 & ~n17378 ;
  assign n17380 = ~n17363 & ~n17370 ;
  assign n17381 = ~n17379 & ~n17380 ;
  assign n17382 = ~n17263 & ~n17272 ;
  assign n17383 = n17270 & ~n17382 ;
  assign n17384 = ~n17270 & n17382 ;
  assign n17385 = ~n17383 & ~n17384 ;
  assign n17386 = n17381 & ~n17385 ;
  assign n17387 = ~n17356 & ~n17386 ;
  assign n17388 = ~n17273 & n17277 ;
  assign n17389 = ~n17278 & ~n17388 ;
  assign n17390 = n17282 & ~n17301 ;
  assign n17391 = ~n17302 & ~n17390 ;
  assign n17392 = n17389 & ~n17391 ;
  assign n17393 = ~n17389 & n17391 ;
  assign n17394 = ~n17392 & ~n17393 ;
  assign n17395 = n17387 & ~n17394 ;
  assign n17396 = ~n17388 & ~n17390 ;
  assign n17397 = n17394 & ~n17396 ;
  assign n17398 = ~n17395 & ~n17397 ;
  assign n17399 = n17339 & n17398 ;
  assign n17400 = ~n17174 & ~n17179 ;
  assign n17401 = ~n17180 & ~n17400 ;
  assign n17403 = \core_eu_em_mac_em_reg_mxopwe_DO_reg[11]/P0001  & ~n14791 ;
  assign n17402 = ~\core_eu_em_mac_em_reg_mxopwe_DO_reg[11]/P0001  & ~n14787 ;
  assign n17404 = ~\core_eu_em_mac_em_reg_mxopwe_DO_reg[10]/P0001  & n14798 ;
  assign n17405 = \core_eu_em_mac_em_reg_mxopwe_DO_reg[10]/P0001  & n14802 ;
  assign n17406 = ~n17404 & ~n17405 ;
  assign n17407 = ~n17402 & n17406 ;
  assign n17408 = ~n17403 & n17407 ;
  assign n17410 = \core_eu_em_mac_em_reg_mxopwe_DO_reg[13]/P0001  & ~n14765 ;
  assign n17409 = ~\core_eu_em_mac_em_reg_mxopwe_DO_reg[13]/P0001  & ~n14761 ;
  assign n17411 = ~\core_eu_em_mac_em_reg_mxopwe_DO_reg[12]/P0001  & n14772 ;
  assign n17412 = \core_eu_em_mac_em_reg_mxopwe_DO_reg[12]/P0001  & n14776 ;
  assign n17413 = ~n17411 & ~n17412 ;
  assign n17414 = ~n17409 & n17413 ;
  assign n17415 = ~n17410 & n17414 ;
  assign n17416 = n17408 & n17415 ;
  assign n17418 = \core_eu_em_mac_em_reg_mxopwe_DO_reg[9]/P0001  & ~n14818 ;
  assign n17417 = ~\core_eu_em_mac_em_reg_mxopwe_DO_reg[9]/P0001  & ~n14814 ;
  assign n17419 = ~\core_eu_em_mac_em_reg_mxopwe_DO_reg[8]/P0001  & n14825 ;
  assign n17420 = \core_eu_em_mac_em_reg_mxopwe_DO_reg[8]/P0001  & n14829 ;
  assign n17421 = ~n17419 & ~n17420 ;
  assign n17422 = ~n17417 & n17421 ;
  assign n17423 = ~n17418 & n17422 ;
  assign n17424 = ~n17416 & ~n17423 ;
  assign n17425 = ~n17408 & ~n17415 ;
  assign n17426 = ~n17424 & ~n17425 ;
  assign n17427 = ~n17152 & ~n17161 ;
  assign n17428 = n17159 & ~n17427 ;
  assign n17429 = ~n17159 & n17427 ;
  assign n17430 = ~n17428 & ~n17429 ;
  assign n17431 = n17426 & ~n17430 ;
  assign n17432 = ~n14967 & n17171 ;
  assign n17433 = ~n17172 & ~n17432 ;
  assign n17435 = \core_eu_em_mac_em_reg_mxopwe_DO_reg[15]/P0001  & ~n14842 ;
  assign n17434 = ~\core_eu_em_mac_em_reg_mxopwe_DO_reg[15]/P0001  & ~n14838 ;
  assign n17436 = ~\core_eu_em_mac_em_reg_mxopwe_DO_reg[14]/P0001  & n14846 ;
  assign n17437 = \core_eu_em_mac_em_reg_mxopwe_DO_reg[14]/P0001  & n14849 ;
  assign n17438 = ~n17436 & ~n17437 ;
  assign n17439 = ~n17434 & n17438 ;
  assign n17440 = ~n17435 & n17439 ;
  assign n17441 = n14958 & ~n17440 ;
  assign n17442 = ~n14958 & n17440 ;
  assign n17443 = \core_c_dec_MACop_E_reg/P0001  & ~\core_eu_em_mac_em_dec_emcorepi_DO_reg[1]/P0001  ;
  assign n17444 = \core_c_psq_MSTAT_reg_DO_reg[4]/NET0131  & n17443 ;
  assign n17445 = ~n12024 & n17444 ;
  assign n17446 = ~n17442 & n17445 ;
  assign n17447 = ~n17441 & ~n17446 ;
  assign n17448 = ~n17433 & n17447 ;
  assign n17449 = ~n17431 & ~n17448 ;
  assign n17450 = ~n17162 & n17166 ;
  assign n17451 = ~n17167 & ~n17450 ;
  assign n17452 = ~n14852 & n17172 ;
  assign n17453 = ~n17173 & ~n17452 ;
  assign n17454 = n17451 & n17453 ;
  assign n17455 = ~n17451 & ~n17453 ;
  assign n17456 = ~n17454 & ~n17455 ;
  assign n17457 = n17449 & n17456 ;
  assign n17458 = ~n17450 & ~n17452 ;
  assign n17459 = ~n17456 & ~n17458 ;
  assign n17460 = ~n17457 & ~n17459 ;
  assign n17461 = ~n17401 & n17460 ;
  assign n17462 = ~n17399 & ~n17461 ;
  assign n17463 = ~n17248 & n17314 ;
  assign n17464 = ~n17315 & ~n17463 ;
  assign n17465 = ~n17137 & ~n17182 ;
  assign n17466 = ~n17183 & ~n17465 ;
  assign n17467 = n17464 & ~n17466 ;
  assign n17468 = ~n17464 & n17466 ;
  assign n17469 = ~n17467 & ~n17468 ;
  assign n17470 = ~n17462 & ~n17469 ;
  assign n17471 = ~n17463 & ~n17465 ;
  assign n17472 = n17469 & n17471 ;
  assign n17473 = ~n17470 & ~n17472 ;
  assign n17474 = ~n17337 & ~n17473 ;
  assign n17475 = n17462 & n17469 ;
  assign n17476 = ~n17470 & ~n17475 ;
  assign n17477 = ~n17449 & ~n17456 ;
  assign n17478 = ~n17457 & ~n17477 ;
  assign n17479 = ~n14947 & ~n15868 ;
  assign n17480 = ~n15869 & ~n17479 ;
  assign n17481 = ~n17441 & ~n17442 ;
  assign n17482 = n17445 & n17481 ;
  assign n17483 = ~n17445 & ~n17481 ;
  assign n17484 = ~n17482 & ~n17483 ;
  assign n17485 = n17480 & ~n17484 ;
  assign n17486 = ~n15839 & ~n15848 ;
  assign n17487 = ~n15840 & ~n17486 ;
  assign n17488 = ~n17416 & ~n17425 ;
  assign n17489 = n17423 & ~n17488 ;
  assign n17490 = ~n17423 & n17488 ;
  assign n17491 = ~n17489 & ~n17490 ;
  assign n17492 = n17487 & ~n17491 ;
  assign n17493 = ~n17485 & ~n17492 ;
  assign n17494 = ~n17426 & n17430 ;
  assign n17495 = ~n17431 & ~n17494 ;
  assign n17496 = n17433 & ~n17447 ;
  assign n17497 = ~n17448 & ~n17496 ;
  assign n17498 = n17495 & n17497 ;
  assign n17499 = ~n17495 & ~n17497 ;
  assign n17500 = ~n17498 & ~n17499 ;
  assign n17501 = n17493 & n17500 ;
  assign n17502 = ~n17494 & ~n17496 ;
  assign n17503 = ~n17500 & ~n17502 ;
  assign n17504 = ~n17501 & ~n17503 ;
  assign n17505 = ~n17478 & n17504 ;
  assign n17506 = ~n17387 & n17394 ;
  assign n17507 = ~n17395 & ~n17506 ;
  assign n17508 = n17343 & n17350 ;
  assign n17509 = ~n17351 & ~n17508 ;
  assign n17510 = ~n15781 & ~n17509 ;
  assign n17511 = ~n15800 & ~n15809 ;
  assign n17512 = ~n15801 & ~n17511 ;
  assign n17513 = ~n17371 & ~n17380 ;
  assign n17514 = n17378 & ~n17513 ;
  assign n17515 = ~n17378 & n17513 ;
  assign n17516 = ~n17514 & ~n17515 ;
  assign n17517 = n17512 & ~n17516 ;
  assign n17518 = ~n17510 & ~n17517 ;
  assign n17519 = ~n17381 & n17385 ;
  assign n17520 = ~n17386 & ~n17519 ;
  assign n17521 = n17351 & n17355 ;
  assign n17522 = ~n17356 & ~n17521 ;
  assign n17523 = n17520 & n17522 ;
  assign n17524 = ~n17520 & ~n17522 ;
  assign n17525 = ~n17523 & ~n17524 ;
  assign n17526 = n17518 & n17525 ;
  assign n17527 = ~n17519 & ~n17521 ;
  assign n17528 = ~n17525 & ~n17527 ;
  assign n17529 = ~n17526 & ~n17528 ;
  assign n17530 = ~n17507 & n17529 ;
  assign n17531 = ~n17505 & ~n17530 ;
  assign n17532 = n17401 & ~n17460 ;
  assign n17533 = ~n17461 & ~n17532 ;
  assign n17534 = ~n17339 & ~n17398 ;
  assign n17535 = ~n17399 & ~n17534 ;
  assign n17536 = n17533 & n17535 ;
  assign n17537 = ~n17533 & ~n17535 ;
  assign n17538 = ~n17536 & ~n17537 ;
  assign n17539 = n17531 & n17538 ;
  assign n17540 = ~n17532 & ~n17534 ;
  assign n17541 = ~n17538 & ~n17540 ;
  assign n17542 = ~n17539 & ~n17541 ;
  assign n17543 = n17476 & n17542 ;
  assign n17544 = ~n17474 & ~n17543 ;
  assign n17545 = ~n17322 & ~n17330 ;
  assign n17546 = ~n16860 & ~n16926 ;
  assign n17547 = ~n16927 & ~n17546 ;
  assign n17548 = n16963 & ~n16965 ;
  assign n17549 = ~n16966 & ~n17548 ;
  assign n17550 = n17547 & n17549 ;
  assign n17551 = ~n17547 & ~n17549 ;
  assign n17552 = ~n17550 & ~n17551 ;
  assign n17553 = ~n17545 & ~n17552 ;
  assign n17554 = n17545 & n17552 ;
  assign n17555 = ~n17553 & ~n17554 ;
  assign n17556 = ~n17323 & ~n17329 ;
  assign n17557 = ~n17334 & ~n17556 ;
  assign n17558 = ~n17336 & ~n17557 ;
  assign n17559 = ~n17555 & n17558 ;
  assign n17560 = ~n17546 & ~n17548 ;
  assign n17561 = ~n17552 & ~n17560 ;
  assign n17562 = ~n17554 & ~n17561 ;
  assign n17563 = n16967 & ~n16974 ;
  assign n17564 = ~n16975 & ~n17563 ;
  assign n17565 = n17562 & n17564 ;
  assign n17566 = ~n17559 & ~n17565 ;
  assign n17567 = n17544 & n17566 ;
  assign n17568 = n17098 & n17567 ;
  assign n17569 = ~n17531 & ~n17538 ;
  assign n17570 = ~n17539 & ~n17569 ;
  assign n17571 = ~n17493 & ~n17500 ;
  assign n17572 = ~n17501 & ~n17571 ;
  assign n17573 = ~n15852 & ~n15874 ;
  assign n17574 = ~n17487 & n17491 ;
  assign n17575 = ~n17492 & ~n17574 ;
  assign n17576 = ~n17480 & n17484 ;
  assign n17577 = ~n17485 & ~n17576 ;
  assign n17578 = n17575 & ~n17577 ;
  assign n17579 = ~n17575 & n17577 ;
  assign n17580 = ~n17578 & ~n17579 ;
  assign n17581 = ~n17573 & ~n17580 ;
  assign n17582 = ~n17574 & ~n17576 ;
  assign n17583 = n17580 & n17582 ;
  assign n17584 = ~n17581 & ~n17583 ;
  assign n17585 = ~n17572 & ~n17584 ;
  assign n17586 = ~n17518 & ~n17525 ;
  assign n17587 = ~n17526 & ~n17586 ;
  assign n17588 = n15783 & ~n15814 ;
  assign n17589 = ~n17512 & n17516 ;
  assign n17590 = ~n17517 & ~n17589 ;
  assign n17591 = n15781 & n17509 ;
  assign n17592 = ~n17510 & ~n17591 ;
  assign n17593 = n17590 & ~n17592 ;
  assign n17594 = ~n17590 & n17592 ;
  assign n17595 = ~n17593 & ~n17594 ;
  assign n17596 = ~n17588 & ~n17595 ;
  assign n17597 = ~n17589 & ~n17591 ;
  assign n17598 = n17595 & n17597 ;
  assign n17599 = ~n17596 & ~n17598 ;
  assign n17600 = ~n17587 & ~n17599 ;
  assign n17601 = ~n17585 & ~n17600 ;
  assign n17602 = n17478 & ~n17504 ;
  assign n17603 = ~n17505 & ~n17602 ;
  assign n17604 = n17507 & ~n17529 ;
  assign n17605 = ~n17530 & ~n17604 ;
  assign n17606 = n17603 & n17605 ;
  assign n17607 = ~n17603 & ~n17605 ;
  assign n17608 = ~n17606 & ~n17607 ;
  assign n17609 = n17601 & n17608 ;
  assign n17610 = ~n17602 & ~n17604 ;
  assign n17611 = ~n17608 & ~n17610 ;
  assign n17612 = ~n17609 & ~n17611 ;
  assign n17613 = ~n17570 & n17612 ;
  assign n17614 = ~n17601 & ~n17608 ;
  assign n17615 = ~n17609 & ~n17614 ;
  assign n17616 = n17573 & n17580 ;
  assign n17617 = ~n17581 & ~n17616 ;
  assign n17618 = ~n15853 & ~n15875 ;
  assign n17619 = ~n15879 & n17618 ;
  assign n17620 = ~n15880 & ~n17619 ;
  assign n17621 = n17617 & ~n17620 ;
  assign n17623 = n17588 & n17595 ;
  assign n17622 = ~n15783 & n15813 ;
  assign n17624 = ~n17596 & ~n17622 ;
  assign n17625 = ~n17623 & n17624 ;
  assign n17626 = ~n17621 & ~n17625 ;
  assign n17627 = n17572 & n17584 ;
  assign n17628 = ~n17585 & ~n17627 ;
  assign n17629 = n17587 & n17599 ;
  assign n17630 = ~n17600 & ~n17629 ;
  assign n17631 = n17628 & ~n17630 ;
  assign n17632 = ~n17628 & n17630 ;
  assign n17633 = ~n17631 & ~n17632 ;
  assign n17634 = ~n17626 & ~n17633 ;
  assign n17635 = ~n17627 & ~n17629 ;
  assign n17636 = n17633 & n17635 ;
  assign n17637 = ~n17634 & ~n17636 ;
  assign n17638 = ~n17615 & ~n17637 ;
  assign n17639 = ~n17613 & ~n17638 ;
  assign n17640 = n17626 & n17633 ;
  assign n17641 = ~n17634 & ~n17640 ;
  assign n17642 = ~n15819 & ~n15886 ;
  assign n17643 = ~n17617 & n17620 ;
  assign n17644 = ~n17621 & ~n17643 ;
  assign n17645 = ~n17595 & n17622 ;
  assign n17646 = ~n17625 & ~n17645 ;
  assign n17647 = n17644 & n17646 ;
  assign n17648 = ~n17644 & ~n17646 ;
  assign n17649 = ~n17647 & ~n17648 ;
  assign n17650 = ~n17642 & n17649 ;
  assign n17651 = ~n17643 & ~n17645 ;
  assign n17652 = ~n17649 & n17651 ;
  assign n17653 = ~n17650 & ~n17652 ;
  assign n17654 = n17641 & ~n17653 ;
  assign n17655 = n17642 & ~n17649 ;
  assign n17656 = ~n17650 & ~n17655 ;
  assign n17657 = ~n15820 & ~n15887 ;
  assign n17658 = ~n15891 & n17657 ;
  assign n17659 = ~n15892 & ~n17658 ;
  assign n17660 = n17656 & ~n17659 ;
  assign n17661 = ~n17654 & ~n17660 ;
  assign n17662 = n17639 & n17661 ;
  assign n17663 = n17568 & n17662 ;
  assign n17664 = ~n16363 & n17663 ;
  assign n17676 = ~n17476 & ~n17542 ;
  assign n17677 = n17337 & n17473 ;
  assign n17678 = ~n17676 & ~n17677 ;
  assign n17679 = ~n17474 & ~n17678 ;
  assign n17680 = n17566 & n17679 ;
  assign n17681 = ~n17562 & ~n17564 ;
  assign n17682 = n17555 & ~n17558 ;
  assign n17683 = ~n17565 & n17682 ;
  assign n17684 = ~n17681 & ~n17683 ;
  assign n17685 = ~n17680 & n17684 ;
  assign n17686 = n17098 & ~n17685 ;
  assign n17667 = ~n17641 & n17653 ;
  assign n17668 = ~n17656 & n17659 ;
  assign n17669 = ~n17667 & ~n17668 ;
  assign n17670 = ~n17654 & ~n17669 ;
  assign n17671 = n17639 & n17670 ;
  assign n17665 = n17615 & n17637 ;
  assign n17666 = ~n17613 & n17665 ;
  assign n17672 = n17570 & ~n17612 ;
  assign n17673 = ~n17666 & ~n17672 ;
  assign n17674 = ~n17671 & n17673 ;
  assign n17675 = n17568 & ~n17674 ;
  assign n17687 = ~n16739 & ~n16855 ;
  assign n17688 = n16858 & n16978 ;
  assign n17689 = ~n16856 & n17688 ;
  assign n17690 = ~n17687 & ~n17689 ;
  assign n17691 = ~n17097 & ~n17690 ;
  assign n17692 = ~n17088 & n17091 ;
  assign n17693 = ~n17095 & ~n17692 ;
  assign n17694 = ~n17079 & ~n17693 ;
  assign n17695 = ~n17691 & ~n17694 ;
  assign n17696 = ~n17675 & n17695 ;
  assign n17697 = ~n17686 & n17696 ;
  assign n17698 = ~n17664 & n17697 ;
  assign n17699 = ~n17051 & ~n17060 ;
  assign n17700 = n15253 & ~n15272 ;
  assign n17701 = ~n15273 & ~n17700 ;
  assign n17702 = ~n15288 & n15291 ;
  assign n17703 = ~n15292 & ~n17702 ;
  assign n17704 = n17701 & ~n17703 ;
  assign n17705 = ~n17701 & n17703 ;
  assign n17706 = ~n17704 & ~n17705 ;
  assign n17707 = ~n17699 & ~n17706 ;
  assign n17708 = n17699 & n17706 ;
  assign n17709 = ~n17707 & ~n17708 ;
  assign n17710 = ~n17050 & ~n17059 ;
  assign n17711 = ~n17064 & n17710 ;
  assign n17712 = ~n17066 & ~n17711 ;
  assign n17713 = n17709 & ~n17712 ;
  assign n17714 = ~n14853 & ~n17713 ;
  assign n17715 = n15293 & ~n15300 ;
  assign n17716 = ~n15301 & ~n17715 ;
  assign n17717 = ~n17700 & ~n17702 ;
  assign n17718 = n17706 & n17717 ;
  assign n17719 = ~n17707 & ~n17718 ;
  assign n17720 = ~n17716 & n17719 ;
  assign n17721 = n17716 & ~n17719 ;
  assign n17722 = ~n17720 & ~n17721 ;
  assign n17723 = n14853 & n17722 ;
  assign n17724 = ~n14853 & ~n17722 ;
  assign n17725 = ~n17723 & ~n17724 ;
  assign n17726 = ~n17714 & ~n17725 ;
  assign n17727 = n17714 & n17722 ;
  assign n17728 = ~n17726 & ~n17727 ;
  assign n17729 = ~n14853 & ~n17071 ;
  assign n17730 = ~n17709 & n17712 ;
  assign n17731 = ~n17713 & ~n17730 ;
  assign n17732 = n14853 & n17731 ;
  assign n17733 = ~n14853 & ~n17731 ;
  assign n17734 = ~n17732 & ~n17733 ;
  assign n17735 = ~n17729 & ~n17734 ;
  assign n17736 = n17729 & n17731 ;
  assign n17737 = ~n17735 & ~n17736 ;
  assign n17738 = ~n17728 & ~n17737 ;
  assign n17739 = ~n17730 & n17734 ;
  assign n17740 = ~n17735 & ~n17739 ;
  assign n17741 = n17728 & ~n17740 ;
  assign n17742 = ~n17072 & n17076 ;
  assign n17743 = ~n17077 & ~n17742 ;
  assign n17744 = ~n17741 & n17743 ;
  assign n17745 = ~n17738 & ~n17744 ;
  assign n17746 = n15306 & n15308 ;
  assign n17747 = ~n15312 & ~n17746 ;
  assign n17748 = ~n17720 & n17725 ;
  assign n17749 = ~n17726 & ~n17748 ;
  assign n17750 = ~n14853 & ~n17721 ;
  assign n17751 = ~n15249 & n15304 ;
  assign n17752 = ~n15305 & ~n17751 ;
  assign n17753 = n14853 & n17752 ;
  assign n17754 = ~n14853 & ~n17752 ;
  assign n17755 = ~n17753 & ~n17754 ;
  assign n17756 = ~n17750 & ~n17755 ;
  assign n17757 = n17750 & n17752 ;
  assign n17758 = ~n17756 & ~n17757 ;
  assign n17759 = ~n17749 & n17758 ;
  assign n17760 = ~n17747 & ~n17759 ;
  assign n17761 = ~n17751 & n17755 ;
  assign n17762 = ~n17756 & ~n17761 ;
  assign n17763 = n17749 & n17762 ;
  assign n17764 = ~n17760 & ~n17763 ;
  assign n17765 = ~n17745 & ~n17764 ;
  assign n17766 = ~n17698 & n17765 ;
  assign n17770 = ~n17728 & n17740 ;
  assign n17771 = n17738 & n17743 ;
  assign n17772 = ~n17770 & ~n17771 ;
  assign n17773 = ~n17764 & ~n17772 ;
  assign n17767 = n17747 & ~n17762 ;
  assign n17768 = n17749 & ~n17758 ;
  assign n17769 = ~n17767 & n17768 ;
  assign n17774 = ~n17747 & n17762 ;
  assign n17775 = ~n17769 & ~n17774 ;
  assign n17776 = ~n17773 & n17775 ;
  assign n17777 = ~n17766 & n17776 ;
  assign n17778 = ~n15314 & n17777 ;
  assign n17779 = ~n15244 & ~n17778 ;
  assign n17780 = ~n15319 & n17779 ;
  assign n17781 = ~n15246 & n15316 ;
  assign n17782 = n15247 & n15314 ;
  assign n17783 = ~n17781 & ~n17782 ;
  assign n17784 = ~n17780 & n17783 ;
  assign n17785 = ~n15183 & ~n17784 ;
  assign n17786 = ~n15182 & ~n17785 ;
  assign n17787 = n15122 & ~n17786 ;
  assign n17788 = ~n15122 & n17786 ;
  assign n17789 = ~n17787 & ~n17788 ;
  assign n17790 = \core_c_psq_MSTAT_reg_DO_reg[4]/NET0131  & ~n17789 ;
  assign n17791 = ~n15182 & ~n15183 ;
  assign n17792 = n17784 & n17791 ;
  assign n17793 = ~n17784 & ~n17791 ;
  assign n17794 = ~n17792 & ~n17793 ;
  assign n17795 = ~\core_c_psq_MSTAT_reg_DO_reg[4]/NET0131  & n17794 ;
  assign n17796 = ~n17790 & ~n17795 ;
  assign n17797 = n14752 & ~n17796 ;
  assign n17798 = ~\core_c_psq_MSTAT_reg_DO_reg[0]/P0002  & n5951 ;
  assign n17799 = \core_c_dec_MTMR2_E_reg/P0001  & n17798 ;
  assign n17800 = ~\core_eu_em_mac_em_reg_mr2rwe_DO_reg[2]/P0001  & ~n17799 ;
  assign n17801 = ~\core_c_dec_Dummy_E_reg/NET0131  & \core_c_dec_MTMR2_E_reg/P0001  ;
  assign n17802 = ~\core_c_dec_Dummy_E_reg/NET0131  & \core_c_dec_MTMR1_E_reg/P0001  ;
  assign n17803 = \core_c_dec_satMR_E_reg/P0001  & ~n4174 ;
  assign n17804 = ~\core_c_dec_Dummy_E_reg/NET0131  & n17803 ;
  assign n17805 = ~n17802 & ~n17804 ;
  assign n17806 = ~\core_c_dec_updMR_E_reg/P0001  & n17805 ;
  assign n17807 = ~n17801 & n17806 ;
  assign n17808 = ~\core_c_psq_MSTAT_reg_DO_reg[0]/P0002  & ~n17807 ;
  assign n17809 = n13801 & ~n17805 ;
  assign n17810 = ~n17799 & ~n17809 ;
  assign n17811 = n17808 & ~n17810 ;
  assign n17812 = ~\core_c_dec_accPM_E_reg/P0001  & ~n8715 ;
  assign n17813 = \core_c_dec_accPM_E_reg/P0001  & ~n12836 ;
  assign n17814 = ~n17812 & ~n17813 ;
  assign n17815 = ~n17809 & n17814 ;
  assign n17816 = n17811 & ~n17815 ;
  assign n17817 = ~n17800 & ~n17816 ;
  assign n17818 = ~\core_c_dec_accPM_E_reg/P0001  & ~n12743 ;
  assign n17819 = \core_c_dec_accPM_E_reg/P0001  & ~n12771 ;
  assign n17820 = ~n17818 & ~n17819 ;
  assign n17821 = \core_c_dec_MTMR1_E_reg/P0001  & ~n17803 ;
  assign n17822 = n17820 & n17821 ;
  assign n17823 = n17798 & n17822 ;
  assign n17824 = ~n17817 & ~n17823 ;
  assign n17825 = ~\core_eu_em_mac_em_reg_mr2rwe_DO_reg[2]/P0001  & ~n17808 ;
  assign n17826 = ~n17824 & ~n17825 ;
  assign n17827 = n17798 & n17803 ;
  assign n17828 = \core_eu_em_mac_em_reg_mr2rwe_DO_reg[7]/P0001  & n17827 ;
  assign n17829 = ~n14752 & ~n17828 ;
  assign n17830 = ~n17826 & n17829 ;
  assign n17831 = ~n17797 & ~n17830 ;
  assign n17832 = ~\core_c_dec_MTSR1_E_reg/P0001  & ~\core_c_dec_updSR_E_reg/P0001  ;
  assign n17833 = n13804 & ~n17832 ;
  assign n17834 = ~\core_c_dec_accPM_E_reg/P0001  & ~n7340 ;
  assign n17835 = \core_c_dec_accPM_E_reg/P0001  & ~n12658 ;
  assign n17836 = ~n17834 & ~n17835 ;
  assign n17837 = \core_c_dec_MTSR1_E_reg/P0001  & ~n17836 ;
  assign n17838 = \core_c_dec_IRE_reg[13]/NET0131  & \core_c_dec_IRE_reg[14]/NET0131  ;
  assign n17839 = \core_c_dec_SHTop_E_reg/P0001  & ~n17838 ;
  assign n17937 = ~n11996 & n13832 ;
  assign n17938 = n13831 & ~n17937 ;
  assign n17939 = \core_c_dec_IRE_reg[13]/NET0131  & ~\core_c_dec_IRE_reg[14]/NET0131  ;
  assign n17940 = ~n17938 & n17939 ;
  assign n17840 = ~\core_c_dec_IRE_reg[13]/NET0131  & \core_c_dec_IRE_reg[14]/NET0131  ;
  assign n17941 = ~\core_c_dec_IRE_reg[12]/NET0131  & \core_eu_ec_cun_AC_reg/P0001  ;
  assign n17942 = \core_eu_ec_cun_AV_reg/P0001  & n17941 ;
  assign n17943 = n17840 & n17942 ;
  assign n17944 = ~n17940 & ~n17943 ;
  assign n17945 = n17839 & ~n17944 ;
  assign n17841 = n7373 & n9272 ;
  assign n17851 = n8501 & n17841 ;
  assign n17853 = n7995 & n17851 ;
  assign n17863 = n9939 & n17853 ;
  assign n17884 = n10789 & n17863 ;
  assign n17885 = n11303 & n17884 ;
  assign n17886 = ~n11303 & ~n17884 ;
  assign n17887 = ~n17885 & ~n17886 ;
  assign n17888 = n17840 & ~n17887 ;
  assign n17890 = ~\core_c_dec_imSHT_E_reg/P0001  & ~n11303 ;
  assign n17889 = \core_c_dec_IRE_reg[6]/NET0131  & \core_c_dec_imSHT_E_reg/P0001  ;
  assign n17891 = ~n17840 & ~n17889 ;
  assign n17892 = ~n17890 & n17891 ;
  assign n17893 = ~n17888 & ~n17892 ;
  assign n17904 = ~n10789 & ~n17863 ;
  assign n17905 = ~n17884 & ~n17904 ;
  assign n17906 = n17840 & ~n17905 ;
  assign n17908 = ~\core_c_dec_imSHT_E_reg/P0001  & ~n10789 ;
  assign n17907 = \core_c_dec_IRE_reg[5]/NET0131  & \core_c_dec_imSHT_E_reg/P0001  ;
  assign n17909 = ~n17840 & ~n17907 ;
  assign n17910 = ~n17908 & n17909 ;
  assign n17911 = ~n17906 & ~n17910 ;
  assign n17946 = n17893 & n17911 ;
  assign n17895 = ~\core_c_dec_imSHT_E_reg/P0001  & ~n7172 ;
  assign n17894 = \core_c_dec_IRE_reg[7]/NET0131  & \core_c_dec_imSHT_E_reg/P0001  ;
  assign n17896 = ~n17840 & ~n17894 ;
  assign n17897 = ~n17895 & n17896 ;
  assign n17899 = n7172 & ~n17885 ;
  assign n17898 = ~n7172 & n17885 ;
  assign n17900 = n17840 & ~n17898 ;
  assign n17901 = ~n17899 & n17900 ;
  assign n17902 = ~n17897 & ~n17901 ;
  assign n17947 = n17839 & n17902 ;
  assign n17948 = n17946 & n17947 ;
  assign n17949 = ~\core_c_dec_IRE_reg[12]/NET0131  & n17948 ;
  assign n17842 = ~n7373 & ~n9272 ;
  assign n17843 = ~n17841 & ~n17842 ;
  assign n17844 = n17840 & ~n17843 ;
  assign n17846 = ~\core_c_dec_imSHT_E_reg/P0001  & ~n9272 ;
  assign n17845 = \core_c_dec_IRE_reg[1]/NET0131  & \core_c_dec_imSHT_E_reg/P0001  ;
  assign n17847 = ~n17840 & ~n17845 ;
  assign n17848 = ~n17846 & n17847 ;
  assign n17849 = ~n17844 & ~n17848 ;
  assign n17850 = n17839 & n17849 ;
  assign n17852 = ~n7995 & ~n17851 ;
  assign n17854 = ~n17852 & ~n17853 ;
  assign n17855 = n17840 & ~n17854 ;
  assign n17857 = ~\core_c_dec_imSHT_E_reg/P0001  & ~n7995 ;
  assign n17856 = \core_c_dec_IRE_reg[3]/NET0131  & \core_c_dec_imSHT_E_reg/P0001  ;
  assign n17858 = ~n17840 & ~n17856 ;
  assign n17859 = ~n17857 & n17858 ;
  assign n17860 = ~n17855 & ~n17859 ;
  assign n17861 = n17839 & n17860 ;
  assign n17862 = ~n17850 & ~n17861 ;
  assign n17864 = ~n9939 & ~n17853 ;
  assign n17865 = ~n17863 & ~n17864 ;
  assign n17866 = n17840 & ~n17865 ;
  assign n17868 = ~\core_c_dec_imSHT_E_reg/P0001  & ~n9939 ;
  assign n17867 = \core_c_dec_IRE_reg[4]/NET0131  & \core_c_dec_imSHT_E_reg/P0001  ;
  assign n17869 = ~n17840 & ~n17867 ;
  assign n17870 = ~n17868 & n17869 ;
  assign n17871 = ~n17866 & ~n17870 ;
  assign n17873 = ~n8501 & ~n17841 ;
  assign n17874 = ~n17851 & ~n17873 ;
  assign n17875 = n17840 & ~n17874 ;
  assign n17877 = ~\core_c_dec_imSHT_E_reg/P0001  & ~n8501 ;
  assign n17876 = \core_c_dec_IRE_reg[2]/NET0131  & \core_c_dec_imSHT_E_reg/P0001  ;
  assign n17878 = ~n17840 & ~n17876 ;
  assign n17879 = ~n17877 & n17878 ;
  assign n17880 = ~n17875 & ~n17879 ;
  assign n17881 = n17839 & n17880 ;
  assign n17950 = n17871 & n17881 ;
  assign n17951 = n17862 & n17950 ;
  assign n17952 = n17949 & n17951 ;
  assign n17926 = \core_c_dec_imSHT_E_reg/P0001  & ~n17840 ;
  assign n17927 = n7373 & ~n17926 ;
  assign n17928 = ~\core_c_dec_IRE_reg[0]/NET0131  & n17926 ;
  assign n17929 = ~n17927 & ~n17928 ;
  assign n17931 = n17839 & n17929 ;
  assign n17903 = ~n17893 & ~n17902 ;
  assign n17918 = \core_c_dec_IRE_reg[12]/NET0131  & n17839 ;
  assign n17919 = ~n17911 & n17918 ;
  assign n17920 = n17903 & n17919 ;
  assign n17872 = n17839 & n17871 ;
  assign n17882 = ~n17872 & ~n17881 ;
  assign n17953 = n17850 & ~n17860 ;
  assign n17954 = n17882 & n17953 ;
  assign n17955 = n17920 & n17954 ;
  assign n17956 = ~n17931 & n17955 ;
  assign n17957 = \core_c_dec_IRE_reg[12]/NET0131  & n17948 ;
  assign n17958 = n17950 & n17953 ;
  assign n17959 = n17957 & n17958 ;
  assign n17960 = n17929 & n17959 ;
  assign n17961 = n17839 & n17960 ;
  assign n17962 = ~n17956 & ~n17961 ;
  assign n17963 = ~n17952 & n17962 ;
  assign n17964 = n17945 & ~n17963 ;
  assign n17916 = n17872 & ~n17880 ;
  assign n17917 = n17862 & n17916 ;
  assign n17970 = n17917 & n17957 ;
  assign n17971 = n17931 & ~n17944 ;
  assign n17972 = n17970 & n17971 ;
  assign n17973 = ~n17871 & n17881 ;
  assign n17974 = n17849 & n17861 ;
  assign n17975 = n17973 & n17974 ;
  assign n17965 = ~n17929 & n17945 ;
  assign n17976 = n17949 & n17965 ;
  assign n17977 = n17975 & n17976 ;
  assign n17978 = ~n17972 & ~n17977 ;
  assign n17979 = n17931 & n17949 ;
  assign n17980 = n17958 & n17979 ;
  assign n17981 = ~n17931 & n17959 ;
  assign n17982 = ~n17980 & ~n17981 ;
  assign n17983 = n17945 & ~n17982 ;
  assign n17984 = n17978 & ~n17983 ;
  assign n17966 = ~n17849 & n17861 ;
  assign n17985 = n17966 & n17973 ;
  assign n17986 = n17920 & n17985 ;
  assign n17987 = n17965 & n17986 ;
  assign n17988 = n17984 & ~n17987 ;
  assign n17967 = n17950 & n17966 ;
  assign n17968 = n17957 & n17967 ;
  assign n17996 = n17931 & n17968 ;
  assign n17997 = n17979 & n17985 ;
  assign n17998 = ~n17996 & ~n17997 ;
  assign n17999 = n17945 & ~n17998 ;
  assign n17989 = ~n17931 & n17949 ;
  assign n17990 = n17953 & n17973 ;
  assign n17991 = n17989 & n17990 ;
  assign n17992 = n17951 & n17957 ;
  assign n17993 = ~n17931 & n17992 ;
  assign n17994 = ~n17991 & ~n17993 ;
  assign n17995 = n17945 & ~n17994 ;
  assign n17969 = n17965 & n17968 ;
  assign n18000 = n17862 & n17973 ;
  assign n18001 = n17920 & n18000 ;
  assign n18002 = n17971 & n18001 ;
  assign n18003 = ~n17969 & ~n18002 ;
  assign n18004 = ~n17995 & n18003 ;
  assign n18005 = ~n17999 & n18004 ;
  assign n18006 = n17988 & n18005 ;
  assign n18007 = ~n17964 & n18006 ;
  assign n18028 = n17916 & n17966 ;
  assign n18139 = n17989 & n18028 ;
  assign n18140 = n17945 & n18139 ;
  assign n18141 = n17955 & n17971 ;
  assign n18142 = ~n18140 & ~n18141 ;
  assign n18143 = n17965 & n17970 ;
  assign n18066 = n17950 & n17974 ;
  assign n18067 = n17957 & n18066 ;
  assign n18144 = n17971 & n18067 ;
  assign n18145 = ~n18143 & ~n18144 ;
  assign n18146 = n18142 & n18145 ;
  assign n17912 = ~\core_c_dec_IRE_reg[12]/NET0131  & ~n17911 ;
  assign n17913 = n17903 & n17912 ;
  assign n17914 = n17839 & ~n17913 ;
  assign n18035 = n17882 & n17966 ;
  assign n18157 = ~n17914 & n18035 ;
  assign n18158 = n17920 & n18028 ;
  assign n18159 = ~n18157 & ~n18158 ;
  assign n18160 = ~n10793 & n13832 ;
  assign n18161 = n14022 & ~n18160 ;
  assign n18162 = n17839 & ~n18161 ;
  assign n18163 = ~n17929 & n18162 ;
  assign n18164 = ~n9943 & n13832 ;
  assign n18165 = n14101 & ~n18164 ;
  assign n18166 = n17931 & ~n18165 ;
  assign n18167 = ~n18163 & ~n18166 ;
  assign n18168 = ~n18159 & ~n18167 ;
  assign n18131 = ~n17914 & n18000 ;
  assign n18132 = n17920 & n17951 ;
  assign n18133 = ~n18131 & ~n18132 ;
  assign n18169 = ~n10222 & n13832 ;
  assign n18170 = n13864 & ~n18169 ;
  assign n18171 = n17839 & ~n18170 ;
  assign n18172 = ~n17929 & n18171 ;
  assign n18173 = ~n18133 & n18172 ;
  assign n18199 = ~n18168 & ~n18173 ;
  assign n18178 = n17920 & n17958 ;
  assign n18179 = ~n17914 & n17990 ;
  assign n18180 = ~n18178 & ~n18179 ;
  assign n18181 = ~n11235 & n13832 ;
  assign n18182 = n13946 & ~n18181 ;
  assign n18183 = n17839 & ~n18182 ;
  assign n18184 = ~n17929 & n18183 ;
  assign n18185 = ~n11307 & n13832 ;
  assign n18186 = n13984 & ~n18185 ;
  assign n18187 = n17839 & ~n18186 ;
  assign n18188 = n17929 & n18187 ;
  assign n18189 = ~n18184 & ~n18188 ;
  assign n18190 = ~n18180 & ~n18189 ;
  assign n17883 = n17862 & n17882 ;
  assign n18191 = n17883 & n17920 ;
  assign n18192 = n17945 & n18191 ;
  assign n18077 = n17882 & n17974 ;
  assign n18193 = ~n17958 & ~n18077 ;
  assign n18194 = n17976 & ~n18193 ;
  assign n18195 = ~n18192 & ~n18194 ;
  assign n18200 = ~n18190 & n18195 ;
  assign n18201 = n18199 & n18200 ;
  assign n18094 = n17920 & n17967 ;
  assign n18095 = ~n17914 & n17985 ;
  assign n18096 = ~n18094 & ~n18095 ;
  assign n18097 = ~n9264 & n13832 ;
  assign n18098 = n14178 & ~n18097 ;
  assign n18099 = n17839 & ~n18098 ;
  assign n18100 = ~n17929 & n18099 ;
  assign n18101 = ~n7369 & n13832 ;
  assign n18102 = ~n14217 & ~n18101 ;
  assign n18103 = n17931 & ~n18102 ;
  assign n18104 = ~n18100 & ~n18103 ;
  assign n18105 = ~n18096 & ~n18104 ;
  assign n18020 = n17916 & n17953 ;
  assign n18106 = n17920 & n18020 ;
  assign n18107 = ~n17914 & n17954 ;
  assign n18108 = ~n18106 & ~n18107 ;
  assign n18109 = ~n8406 & n13832 ;
  assign n18110 = n14290 & ~n18109 ;
  assign n18111 = n17839 & ~n18110 ;
  assign n18112 = ~n17929 & n18111 ;
  assign n18113 = ~n7805 & n13832 ;
  assign n18114 = n14332 & ~n18113 ;
  assign n18115 = n17839 & ~n18114 ;
  assign n18116 = n17929 & n18115 ;
  assign n18117 = ~n18112 & ~n18116 ;
  assign n18118 = ~n18108 & ~n18117 ;
  assign n18197 = ~n18105 & ~n18118 ;
  assign n18119 = ~n17914 & n18077 ;
  assign n18045 = n17916 & n17974 ;
  assign n18120 = n17920 & n18045 ;
  assign n18121 = ~n18119 & ~n18120 ;
  assign n18122 = ~n7979 & n13832 ;
  assign n18123 = n14066 & ~n18122 ;
  assign n18124 = n17839 & ~n18123 ;
  assign n18125 = ~n17929 & n18124 ;
  assign n18126 = ~n8485 & n13832 ;
  assign n18127 = n14140 & ~n18126 ;
  assign n18128 = n17931 & ~n18127 ;
  assign n18129 = ~n18125 & ~n18128 ;
  assign n18130 = ~n18121 & ~n18129 ;
  assign n18134 = ~n10571 & n13832 ;
  assign n18135 = n13909 & ~n18134 ;
  assign n18136 = n17931 & ~n18135 ;
  assign n18137 = ~n18133 & n18136 ;
  assign n18198 = ~n18130 & ~n18137 ;
  assign n18202 = n18197 & n18198 ;
  assign n18205 = n18201 & n18202 ;
  assign n18206 = n18146 & n18205 ;
  assign n18150 = n17979 & n17990 ;
  assign n18151 = n17989 & n18000 ;
  assign n18152 = ~n18150 & ~n18151 ;
  assign n18147 = n17967 & n17979 ;
  assign n18148 = n17931 & n17986 ;
  assign n18149 = ~n18147 & ~n18148 ;
  assign n18153 = n17920 & n18077 ;
  assign n18154 = n18149 & ~n18153 ;
  assign n18155 = n18152 & n18154 ;
  assign n18156 = n17945 & ~n18155 ;
  assign n18174 = ~n11850 & n13832 ;
  assign n18175 = n14506 & ~n18174 ;
  assign n18089 = n17920 & n17975 ;
  assign n18090 = n17949 & n18066 ;
  assign n18091 = ~n18089 & ~n18090 ;
  assign n18176 = n17931 & ~n18091 ;
  assign n18177 = ~n18175 & n18176 ;
  assign n18088 = n17839 & ~n17938 ;
  assign n18092 = ~n17931 & ~n18091 ;
  assign n18093 = n18088 & n18092 ;
  assign n17915 = n17883 & ~n17914 ;
  assign n17921 = n17917 & n17920 ;
  assign n17922 = ~n17915 & ~n17921 ;
  assign n17923 = ~n7160 & n13832 ;
  assign n17924 = n14444 & ~n17923 ;
  assign n17925 = n17839 & ~n17924 ;
  assign n17930 = n17925 & ~n17929 ;
  assign n17932 = ~n9124 & n13832 ;
  assign n17933 = n14377 & ~n17932 ;
  assign n17934 = n17931 & ~n17933 ;
  assign n17935 = ~n17930 & ~n17934 ;
  assign n17936 = ~n17922 & ~n17935 ;
  assign n18138 = \core_c_dec_IRE_reg[11]/NET0131  & ~n7156 ;
  assign n18196 = ~n17936 & ~n18138 ;
  assign n18203 = ~n18093 & n18196 ;
  assign n18204 = ~n18177 & n18203 ;
  assign n18207 = ~n18156 & n18204 ;
  assign n18208 = n18206 & n18207 ;
  assign n18027 = n17985 & n17989 ;
  assign n18029 = n17957 & n18028 ;
  assign n18030 = ~n17931 & n18029 ;
  assign n18031 = ~n18027 & ~n18030 ;
  assign n18032 = n17945 & ~n18031 ;
  assign n18033 = n17949 & n17975 ;
  assign n18034 = n17971 & n18033 ;
  assign n18036 = n17949 & n18035 ;
  assign n18037 = n17945 & n18036 ;
  assign n18038 = ~n18034 & ~n18037 ;
  assign n18039 = n17917 & n17949 ;
  assign n18040 = n17971 & n18039 ;
  assign n18041 = n18038 & ~n18040 ;
  assign n18042 = ~n18032 & n18041 ;
  assign n18043 = n17967 & n17989 ;
  assign n18021 = n17957 & n18020 ;
  assign n18044 = ~n17931 & n18021 ;
  assign n18046 = n17979 & n18045 ;
  assign n18047 = ~n18044 & ~n18046 ;
  assign n18048 = ~n18043 & n18047 ;
  assign n18049 = n17945 & ~n18048 ;
  assign n18050 = n18042 & ~n18049 ;
  assign n18008 = \core_c_dec_IRE_reg[12]/NET0131  & ~n17893 ;
  assign n18009 = n17902 & n17945 ;
  assign n18010 = n18008 & n18009 ;
  assign n18011 = ~n17871 & n17945 ;
  assign n18012 = n17957 & n18011 ;
  assign n18013 = ~n17946 & ~n18008 ;
  assign n18014 = n18009 & n18013 ;
  assign n18015 = ~n18012 & ~n18014 ;
  assign n18016 = ~n18010 & n18015 ;
  assign n18017 = n17883 & n17949 ;
  assign n18018 = n17945 & n18017 ;
  assign n18019 = n18016 & ~n18018 ;
  assign n18022 = n17931 & n18021 ;
  assign n18023 = ~n17944 & n18022 ;
  assign n18024 = n18019 & ~n18023 ;
  assign n18051 = n17957 & n18045 ;
  assign n18052 = n17965 & n18051 ;
  assign n18053 = n17971 & n18029 ;
  assign n18054 = ~n18052 & ~n18053 ;
  assign n18055 = n17920 & n18035 ;
  assign n18056 = n17920 & n17990 ;
  assign n18057 = ~n18055 & ~n18056 ;
  assign n18058 = n17965 & ~n18057 ;
  assign n18059 = n18054 & ~n18058 ;
  assign n18025 = n17945 & n17949 ;
  assign n18026 = n17954 & n18025 ;
  assign n18060 = n17965 & n18001 ;
  assign n18061 = ~n18026 & ~n18060 ;
  assign n18062 = n18059 & n18061 ;
  assign n18063 = n18024 & n18062 ;
  assign n18064 = n18050 & n18063 ;
  assign n18068 = ~n18039 & ~n18067 ;
  assign n18069 = n17965 & ~n18068 ;
  assign n18071 = n17979 & n18028 ;
  assign n18070 = n17989 & n18045 ;
  assign n18072 = n17949 & n18020 ;
  assign n18073 = ~n18070 & ~n18072 ;
  assign n18074 = ~n18071 & n18073 ;
  assign n18075 = n17945 & ~n18074 ;
  assign n18076 = ~n18069 & ~n18075 ;
  assign n18065 = n17971 & ~n18057 ;
  assign n18078 = n17949 & n18077 ;
  assign n18079 = ~n18051 & ~n18078 ;
  assign n18080 = n17931 & ~n18079 ;
  assign n18081 = n17949 & n18000 ;
  assign n18082 = ~n17992 & ~n18081 ;
  assign n18083 = n17931 & ~n18082 ;
  assign n18084 = ~n18080 & ~n18083 ;
  assign n18085 = n17945 & ~n18084 ;
  assign n18086 = ~n18065 & ~n18085 ;
  assign n18087 = n18076 & n18086 ;
  assign n18209 = n18064 & n18087 ;
  assign n18210 = n18208 & n18209 ;
  assign n18211 = n18007 & n18210 ;
  assign n18212 = ~\core_c_dec_MTSR1_E_reg/P0001  & n18211 ;
  assign n18213 = ~n17837 & ~n18212 ;
  assign n18214 = n17833 & ~n18213 ;
  assign n18215 = ~\core_eu_es_sht_es_reg_sr1rwe_DO_reg[13]/P0001  & ~n17833 ;
  assign n18216 = ~n18214 & ~n18215 ;
  assign n18217 = \core_c_psq_TRAP_Eg_reg/NET0131  & ~n4112 ;
  assign n18218 = ~\core_c_dec_IRE_reg[0]/NET0131  & n14691 ;
  assign n18219 = ~n5950 & n18218 ;
  assign n18220 = ~n18217 & ~n18219 ;
  assign n18221 = n14713 & ~n18220 ;
  assign n18222 = \core_c_psq_ststk_sts7x23_STcell_reg[3][0]/P0001  & ~n18221 ;
  assign n18223 = \core_eu_ec_cun_AZ_reg/P0001  & n18221 ;
  assign n18224 = ~n18222 & ~n18223 ;
  assign n18225 = \core_dag_ilm1reg_DMA_pi_DO_reg[4]/NET0131  & n5944 ;
  assign n18226 = n13761 & n18225 ;
  assign n18227 = ~\memc_MMR_web_reg/NET0131  & n18226 ;
  assign n18228 = n7237 & n7283 ;
  assign n18229 = n18227 & n18228 ;
  assign n18230 = n7226 & n7283 ;
  assign n18231 = n18227 & n18230 ;
  assign n18232 = n12688 & n18231 ;
  assign n18233 = ~n18229 & ~n18232 ;
  assign n18234 = \sport0_regs_SCTLreg_DO_reg[12]/NET0131  & n18233 ;
  assign n18235 = n12688 & n18226 ;
  assign n18236 = n18230 & n18235 ;
  assign n18237 = n18229 & ~n18236 ;
  assign n18238 = n9178 & n18237 ;
  assign n18239 = ~n18234 & ~n18238 ;
  assign n18240 = n14708 & ~n18220 ;
  assign n18241 = \core_c_psq_ststk_sts7x23_STcell_reg[2][9]/P0001  & ~n18240 ;
  assign n18242 = \core_c_psq_MSTAT_reg_DO_reg[1]/NET0131  & n18240 ;
  assign n18243 = ~n18241 & ~n18242 ;
  assign n18244 = \core_c_psq_ststk_sts7x23_STcell_reg[2][8]/P0001  & ~n18240 ;
  assign n18245 = \core_c_psq_MSTAT_reg_DO_reg[0]/P0002  & n18240 ;
  assign n18246 = ~n18244 & ~n18245 ;
  assign n18247 = \core_c_psq_ststk_sts7x23_STcell_reg[2][7]/P0001  & ~n18240 ;
  assign n18248 = \core_eu_ec_cun_SS_reg/P0001  & n18240 ;
  assign n18249 = ~n18247 & ~n18248 ;
  assign n18250 = \core_c_psq_ststk_sts7x23_STcell_reg[2][6]/P0001  & ~n18240 ;
  assign n18251 = ~n4174 & n18240 ;
  assign n18252 = ~n18250 & ~n18251 ;
  assign n18253 = \core_c_psq_ststk_sts7x23_STcell_reg[2][5]/P0001  & ~n18240 ;
  assign n18254 = \core_eu_ec_cun_AQ_reg/P0001  & n18240 ;
  assign n18255 = ~n18253 & ~n18254 ;
  assign n18256 = \core_c_psq_ststk_sts7x23_STcell_reg[2][4]/P0001  & ~n18240 ;
  assign n18257 = \core_eu_ec_cun_AS_reg/P0001  & n18240 ;
  assign n18258 = ~n18256 & ~n18257 ;
  assign n18259 = \core_c_psq_ststk_sts7x23_STcell_reg[2][3]/P0001  & ~n18240 ;
  assign n18260 = \core_eu_ec_cun_AC_reg/P0001  & n18240 ;
  assign n18261 = ~n18259 & ~n18260 ;
  assign n18262 = \core_c_dec_updMR_E_reg/P0001  & n14666 ;
  assign n18271 = \core_c_dec_MTMR0_E_reg/P0001  & n14665 ;
  assign n18274 = ~\core_c_dec_accPM_E_reg/P0001  & ~n11525 ;
  assign n18275 = \core_c_dec_accPM_E_reg/P0001  & ~n12972 ;
  assign n18276 = ~n18274 & ~n18275 ;
  assign n18277 = n18271 & ~n18276 ;
  assign n18272 = ~\core_eu_em_mac_em_reg_mr0swe_DO_reg[6]/P0001  & ~n18271 ;
  assign n18263 = ~\core_c_dec_Dummy_E_reg/NET0131  & \core_c_dec_MTMR0_E_reg/P0001  ;
  assign n18264 = ~n17804 & ~n18263 ;
  assign n18265 = ~\core_c_dec_updMR_E_reg/P0001  & n18264 ;
  assign n18266 = \core_c_psq_MSTAT_reg_DO_reg[0]/P0002  & ~n18265 ;
  assign n18268 = n14665 & n17803 ;
  assign n18273 = n18266 & ~n18268 ;
  assign n18278 = ~n18272 & n18273 ;
  assign n18279 = ~n18277 & n18278 ;
  assign n18267 = \core_eu_em_mac_em_reg_mr0swe_DO_reg[6]/P0001  & ~n18266 ;
  assign n18269 = ~\core_eu_em_mac_em_reg_mr2swe_DO_reg[7]/P0001  & n18268 ;
  assign n18270 = n18266 & n18269 ;
  assign n18280 = ~n18267 & ~n18270 ;
  assign n18281 = ~n18279 & n18280 ;
  assign n18282 = ~n18262 & ~n18281 ;
  assign n18283 = ~n16239 & n16306 ;
  assign n18284 = ~n16307 & ~n18283 ;
  assign n18285 = ~\core_c_psq_MSTAT_reg_DO_reg[4]/NET0131  & ~n18284 ;
  assign n18286 = ~n16196 & ~n16197 ;
  assign n18287 = ~n16308 & n18286 ;
  assign n18288 = n16308 & ~n18286 ;
  assign n18289 = ~n18287 & ~n18288 ;
  assign n18290 = \core_c_psq_MSTAT_reg_DO_reg[4]/NET0131  & ~n18289 ;
  assign n18291 = ~n18285 & ~n18290 ;
  assign n18292 = n18262 & n18291 ;
  assign n18293 = ~n18282 & ~n18292 ;
  assign n18294 = \core_c_psq_ststk_sts7x23_STcell_reg[2][2]/P0001  & ~n18240 ;
  assign n18295 = \core_eu_ec_cun_AV_reg/P0001  & n18240 ;
  assign n18296 = ~n18294 & ~n18295 ;
  assign n18297 = \core_c_psq_ststk_sts7x23_STcell_reg[2][24]/P0001  & ~n18240 ;
  assign n18298 = \core_c_psq_IMASK_reg[9]/NET0131  & n18240 ;
  assign n18299 = ~n18297 & ~n18298 ;
  assign n18300 = \core_c_psq_ststk_sts7x23_STcell_reg[2][23]/P0001  & ~n18240 ;
  assign n18301 = \core_c_psq_IMASK_reg[8]/NET0131  & n18240 ;
  assign n18302 = ~n18300 & ~n18301 ;
  assign n18303 = \core_c_psq_ststk_sts7x23_STcell_reg[2][22]/P0001  & ~n18240 ;
  assign n18304 = \core_c_psq_IMASK_reg[7]/NET0131  & n18240 ;
  assign n18305 = ~n18303 & ~n18304 ;
  assign n18306 = \core_c_psq_ststk_sts7x23_STcell_reg[2][21]/P0001  & ~n18240 ;
  assign n18307 = \core_c_psq_IMASK_reg[6]/NET0131  & n18240 ;
  assign n18308 = ~n18306 & ~n18307 ;
  assign n18309 = \core_c_psq_ststk_sts7x23_STcell_reg[2][20]/P0001  & ~n18240 ;
  assign n18310 = \core_c_psq_IMASK_reg[5]/NET0131  & n18240 ;
  assign n18311 = ~n18309 & ~n18310 ;
  assign n18312 = \core_c_psq_ststk_sts7x23_STcell_reg[2][1]/P0001  & ~n18240 ;
  assign n18313 = \core_eu_ec_cun_AN_reg/P0001  & n18240 ;
  assign n18314 = ~n18312 & ~n18313 ;
  assign n18315 = \core_c_psq_ststk_sts7x23_STcell_reg[2][19]/P0001  & ~n18240 ;
  assign n18316 = \core_c_psq_IMASK_reg[4]/NET0131  & n18240 ;
  assign n18317 = ~n18315 & ~n18316 ;
  assign n18318 = \core_c_psq_ststk_sts7x23_STcell_reg[2][18]/P0001  & ~n18240 ;
  assign n18319 = \core_c_psq_IMASK_reg[3]/NET0131  & n18240 ;
  assign n18320 = ~n18318 & ~n18319 ;
  assign n18321 = \core_c_psq_ststk_sts7x23_STcell_reg[2][17]/P0001  & ~n18240 ;
  assign n18322 = \core_c_psq_IMASK_reg[2]/NET0131  & n18240 ;
  assign n18323 = ~n18321 & ~n18322 ;
  assign n18324 = n14752 & ~n18291 ;
  assign n18326 = ~\core_c_psq_MSTAT_reg_DO_reg[0]/P0002  & ~n18265 ;
  assign n18325 = n13801 & ~n17804 ;
  assign n18327 = n18263 & n18325 ;
  assign n18328 = n18326 & n18327 ;
  assign n18329 = n18276 & n18328 ;
  assign n18330 = n13801 & ~n18264 ;
  assign n18331 = \core_eu_em_mac_em_reg_mr0rwe_DO_reg[6]/P0001  & ~n18330 ;
  assign n18332 = ~\core_eu_em_mac_em_reg_mr2rwe_DO_reg[7]/P0001  & n17827 ;
  assign n18333 = n18326 & n18332 ;
  assign n18334 = ~n14752 & ~n18333 ;
  assign n18335 = ~n18331 & n18334 ;
  assign n18336 = ~n18329 & n18335 ;
  assign n18337 = ~n18324 & ~n18336 ;
  assign n18338 = \core_c_psq_ststk_sts7x23_STcell_reg[2][16]/P0001  & ~n18240 ;
  assign n18339 = \core_c_psq_IMASK_reg[1]/NET0131  & n18240 ;
  assign n18340 = ~n18338 & ~n18339 ;
  assign n18341 = \core_c_psq_ststk_sts7x23_STcell_reg[2][15]/P0001  & ~n18240 ;
  assign n18342 = \core_c_psq_IMASK_reg[0]/NET0131  & n18240 ;
  assign n18343 = ~n18341 & ~n18342 ;
  assign n18344 = \core_c_psq_ststk_sts7x23_STcell_reg[2][14]/P0001  & ~n18240 ;
  assign n18345 = \core_c_psq_MSTAT_reg_DO_reg[6]/NET0131  & n18240 ;
  assign n18346 = ~n18344 & ~n18345 ;
  assign n18347 = \core_c_psq_ststk_sts7x23_STcell_reg[2][13]/P0001  & ~n18240 ;
  assign n18348 = \core_c_psq_MSTAT_reg_DO_reg[5]/NET0131  & n18240 ;
  assign n18349 = ~n18347 & ~n18348 ;
  assign n18350 = \core_c_psq_ststk_sts7x23_STcell_reg[2][12]/P0001  & ~n18240 ;
  assign n18351 = \core_c_psq_MSTAT_reg_DO_reg[4]/NET0131  & n18240 ;
  assign n18352 = ~n18350 & ~n18351 ;
  assign n18353 = \core_c_psq_ststk_sts7x23_STcell_reg[2][11]/P0001  & ~n18240 ;
  assign n18354 = \core_c_psq_MSTAT_reg_DO_reg[3]/NET0131  & n18240 ;
  assign n18355 = ~n18353 & ~n18354 ;
  assign n18356 = \core_c_psq_ststk_sts7x23_STcell_reg[2][10]/P0001  & ~n18240 ;
  assign n18357 = \core_c_psq_MSTAT_reg_DO_reg[2]/NET0131  & n18240 ;
  assign n18358 = ~n18356 & ~n18357 ;
  assign n18359 = \core_c_psq_ststk_sts7x23_STcell_reg[2][0]/P0001  & ~n18240 ;
  assign n18360 = \core_eu_ec_cun_AZ_reg/P0001  & n18240 ;
  assign n18361 = ~n18359 & ~n18360 ;
  assign n18362 = n14702 & ~n18220 ;
  assign n18363 = \core_c_psq_ststk_sts7x23_STcell_reg[1][9]/P0001  & ~n18362 ;
  assign n18364 = \core_c_psq_MSTAT_reg_DO_reg[1]/NET0131  & n18362 ;
  assign n18365 = ~n18363 & ~n18364 ;
  assign n18366 = \core_c_psq_ststk_sts7x23_STcell_reg[1][8]/P0001  & ~n18362 ;
  assign n18367 = \core_c_psq_MSTAT_reg_DO_reg[0]/P0002  & n18362 ;
  assign n18368 = ~n18366 & ~n18367 ;
  assign n18369 = ~\sport0_txctl_TX_reg[0]/P0001  & ~\sport0_txctl_TX_reg[1]/P0001  ;
  assign n18370 = ~\sport0_txctl_TX_reg[2]/P0001  & n18369 ;
  assign n18371 = ~\sport0_txctl_TX_reg[3]/P0001  & n18370 ;
  assign n18372 = ~\sport0_txctl_TX_reg[4]/P0001  & n18371 ;
  assign n18373 = ~\sport0_txctl_TX_reg[5]/P0001  & n18372 ;
  assign n18374 = ~\sport0_txctl_TX_reg[6]/P0001  & n18373 ;
  assign n18375 = ~\sport0_txctl_TX_reg[7]/P0001  & n18374 ;
  assign n18376 = ~\sport0_txctl_TX_reg[8]/P0001  & n18375 ;
  assign n18377 = \sport0_txctl_TX_reg[15]/P0001  & ~n18376 ;
  assign n18378 = \sport0_txctl_TX_reg[9]/P0001  & n18377 ;
  assign n18379 = ~\sport0_txctl_TX_reg[9]/P0001  & ~n18377 ;
  assign n18380 = ~n18378 & ~n18379 ;
  assign n18381 = \sport0_txctl_TX_reg[15]/P0001  & ~n18372 ;
  assign n18382 = ~\sport0_txctl_TX_reg[5]/P0001  & ~n18381 ;
  assign n18383 = \sport0_txctl_TX_reg[5]/P0001  & n18381 ;
  assign n18384 = ~n18382 & ~n18383 ;
  assign n18385 = ~\sport0_regs_SCTLreg_DO_reg[4]/NET0131  & n18384 ;
  assign n18386 = ~\sport0_txctl_TX_reg[15]/P0001  & \sport0_txctl_TX_reg[1]/P0001  ;
  assign n18387 = \sport0_txctl_TX_reg[0]/P0001  & \sport0_txctl_TX_reg[1]/P0001  ;
  assign n18388 = \sport0_txctl_TX_reg[15]/P0001  & ~n18369 ;
  assign n18389 = ~n18387 & n18388 ;
  assign n18390 = ~n18386 & ~n18389 ;
  assign n18391 = ~\sport0_regs_SCTLreg_DO_reg[4]/NET0131  & ~n18390 ;
  assign n18392 = \sport0_txctl_TX_reg[0]/P0001  & n18391 ;
  assign n18393 = \sport0_txctl_TX_reg[2]/P0001  & ~n18388 ;
  assign n18394 = ~\sport0_txctl_TX_reg[2]/P0001  & n18388 ;
  assign n18395 = ~n18393 & ~n18394 ;
  assign n18396 = n18392 & ~n18395 ;
  assign n18397 = \sport0_txctl_TX_reg[15]/P0001  & ~n18370 ;
  assign n18398 = \sport0_txctl_TX_reg[3]/P0001  & ~n18397 ;
  assign n18399 = ~\sport0_txctl_TX_reg[3]/P0001  & n18397 ;
  assign n18400 = ~n18398 & ~n18399 ;
  assign n18401 = n18396 & ~n18400 ;
  assign n18402 = ~\sport0_txctl_TX_reg[15]/P0001  & \sport0_txctl_TX_reg[4]/P0001  ;
  assign n18403 = \sport0_txctl_TX_reg[4]/P0001  & ~n18371 ;
  assign n18404 = n18381 & ~n18403 ;
  assign n18405 = ~n18402 & ~n18404 ;
  assign n18406 = n18401 & ~n18405 ;
  assign n18407 = ~n18385 & ~n18406 ;
  assign n18408 = \sport0_txctl_TX_reg[15]/P0001  & ~n18373 ;
  assign n18409 = \sport0_txctl_TX_reg[6]/P0001  & n18408 ;
  assign n18410 = ~\sport0_txctl_TX_reg[6]/P0001  & ~n18408 ;
  assign n18411 = ~n18409 & ~n18410 ;
  assign n18412 = ~n18407 & n18411 ;
  assign n18413 = \sport0_txctl_TX_reg[15]/P0001  & ~n18374 ;
  assign n18414 = \sport0_txctl_TX_reg[7]/P0001  & n18413 ;
  assign n18415 = ~\sport0_txctl_TX_reg[7]/P0001  & ~n18413 ;
  assign n18416 = ~n18414 & ~n18415 ;
  assign n18417 = n18412 & n18416 ;
  assign n18418 = \sport0_txctl_TX_reg[15]/P0001  & ~n18375 ;
  assign n18419 = \sport0_txctl_TX_reg[8]/P0001  & n18418 ;
  assign n18420 = ~\sport0_txctl_TX_reg[8]/P0001  & ~n18418 ;
  assign n18421 = ~n18419 & ~n18420 ;
  assign n18422 = n18417 & n18421 ;
  assign n18423 = n18380 & n18422 ;
  assign n18424 = ~\sport0_txctl_TX_reg[9]/P0001  & n18376 ;
  assign n18425 = \sport0_txctl_TX_reg[15]/P0001  & ~n18424 ;
  assign n18426 = ~\sport0_txctl_TX_reg[10]/P0001  & ~n18425 ;
  assign n18427 = \sport0_txctl_TX_reg[10]/P0001  & \sport0_txctl_TX_reg[15]/P0001  ;
  assign n18428 = ~n18424 & n18427 ;
  assign n18429 = ~n18426 & ~n18428 ;
  assign n18430 = n18423 & n18429 ;
  assign n18431 = ~n18425 & ~n18427 ;
  assign n18432 = \sport0_txctl_TX_reg[11]/P0001  & ~n18431 ;
  assign n18433 = ~\sport0_txctl_TX_reg[11]/P0001  & n18431 ;
  assign n18434 = ~n18432 & ~n18433 ;
  assign n18435 = n18430 & n18434 ;
  assign n18436 = ~\sport0_txctl_TX_reg[10]/P0001  & ~\sport0_txctl_TX_reg[11]/P0001  ;
  assign n18437 = \sport0_txctl_TX_reg[15]/P0001  & ~n18436 ;
  assign n18438 = ~n18425 & ~n18437 ;
  assign n18439 = \sport0_txctl_TX_reg[12]/P0001  & ~n18438 ;
  assign n18440 = ~\sport0_txctl_TX_reg[12]/P0001  & n18438 ;
  assign n18441 = ~n18439 & ~n18440 ;
  assign n18442 = n18435 & n18441 ;
  assign n18443 = ~n18435 & ~n18441 ;
  assign n18444 = ~n18442 & ~n18443 ;
  assign n18445 = \sport0_regs_SCTLreg_DO_reg[4]/NET0131  & n18444 ;
  assign n18451 = \sport0_regs_SCTLreg_DO_reg[4]/NET0131  & ~n18384 ;
  assign n18452 = n18442 & ~n18451 ;
  assign n18446 = ~\sport0_txctl_TX_reg[12]/P0001  & n18436 ;
  assign n18447 = n18424 & n18446 ;
  assign n18448 = \sport0_txctl_TX_reg[13]/P0001  & \sport0_txctl_TX_reg[15]/P0001  ;
  assign n18449 = ~n18447 & n18448 ;
  assign n18450 = \sport0_txctl_TX_reg[14]/P0001  & ~n18449 ;
  assign n18453 = ~\sport0_txctl_TX_reg[13]/P0001  & ~\sport0_txctl_TX_reg[15]/P0001  ;
  assign n18454 = ~\sport0_txctl_TX_reg[14]/P0001  & ~n18453 ;
  assign n18455 = ~n18450 & ~n18454 ;
  assign n18456 = ~n18452 & n18455 ;
  assign n18457 = ~n18445 & n18456 ;
  assign n18458 = n18430 & ~n18451 ;
  assign n18459 = n18434 & ~n18458 ;
  assign n18460 = ~n18434 & n18458 ;
  assign n18461 = ~n18459 & ~n18460 ;
  assign n18462 = ~\sport0_regs_SCTLreg_DO_reg[4]/NET0131  & ~n18461 ;
  assign n18463 = ~n18423 & ~n18429 ;
  assign n18464 = ~n18430 & ~n18463 ;
  assign n18465 = \sport0_regs_SCTLreg_DO_reg[4]/NET0131  & n18464 ;
  assign n18466 = ~n18462 & ~n18465 ;
  assign n18467 = n18457 & n18466 ;
  assign n18468 = \sport0_regs_SCTLreg_DO_reg[4]/NET0131  & ~n18461 ;
  assign n18469 = ~n18444 & n18456 ;
  assign n18470 = ~n18468 & n18469 ;
  assign n18471 = n18467 & n18470 ;
  assign n18472 = ~\sport0_regs_SCTLreg_DO_reg[4]/NET0131  & n18464 ;
  assign n18473 = n18422 & ~n18451 ;
  assign n18474 = n18380 & ~n18473 ;
  assign n18475 = ~n18380 & n18473 ;
  assign n18476 = ~n18474 & ~n18475 ;
  assign n18477 = \sport0_regs_SCTLreg_DO_reg[4]/NET0131  & ~n18476 ;
  assign n18478 = ~n18472 & ~n18477 ;
  assign n18479 = n18457 & n18478 ;
  assign n18480 = n18471 & n18479 ;
  assign n18481 = ~n18467 & n18470 ;
  assign n18482 = ~n18480 & ~n18481 ;
  assign n18483 = n18407 & ~n18411 ;
  assign n18484 = ~n18412 & ~n18483 ;
  assign n18485 = ~\sport0_regs_SCTLreg_DO_reg[4]/NET0131  & ~n18484 ;
  assign n18486 = ~n18385 & ~n18451 ;
  assign n18487 = n18406 & n18486 ;
  assign n18488 = ~n18406 & ~n18486 ;
  assign n18489 = ~n18487 & ~n18488 ;
  assign n18490 = \sport0_regs_SCTLreg_DO_reg[4]/NET0131  & ~n18489 ;
  assign n18491 = ~n18485 & ~n18490 ;
  assign n18492 = n18457 & n18491 ;
  assign n18493 = n18412 & ~n18451 ;
  assign n18494 = n18416 & ~n18493 ;
  assign n18495 = ~n18416 & n18493 ;
  assign n18496 = ~n18494 & ~n18495 ;
  assign n18497 = ~\sport0_regs_SCTLreg_DO_reg[4]/NET0131  & ~n18496 ;
  assign n18498 = \sport0_regs_SCTLreg_DO_reg[4]/NET0131  & n18484 ;
  assign n18499 = ~n18497 & ~n18498 ;
  assign n18500 = n18457 & n18499 ;
  assign n18501 = n18492 & n18500 ;
  assign n18502 = \sport0_regs_SCTLreg_DO_reg[4]/NET0131  & ~n18496 ;
  assign n18503 = ~n18417 & ~n18421 ;
  assign n18504 = ~n18422 & ~n18503 ;
  assign n18505 = ~\sport0_regs_SCTLreg_DO_reg[4]/NET0131  & n18504 ;
  assign n18506 = ~n18502 & ~n18505 ;
  assign n18507 = n18457 & n18506 ;
  assign n18508 = ~n18501 & n18507 ;
  assign n18509 = ~\sport0_regs_SCTLreg_DO_reg[4]/NET0131  & ~n18476 ;
  assign n18510 = \sport0_regs_SCTLreg_DO_reg[4]/NET0131  & n18504 ;
  assign n18511 = ~n18509 & ~n18510 ;
  assign n18512 = n18457 & n18511 ;
  assign n18513 = n18479 & n18512 ;
  assign n18514 = n18471 & n18513 ;
  assign n18515 = ~n18508 & n18514 ;
  assign n18516 = ~n18482 & ~n18515 ;
  assign n18517 = \sport0_txctl_ldTX_cmp_reg/P0001  & ~n18516 ;
  assign n18518 = \core_c_dec_MTTX0_E_reg/P0001  & n5951 ;
  assign n18519 = ~\auctl_T0Sack_reg/NET0131  & ~n18518 ;
  assign n18521 = n10069 & ~n18519 ;
  assign n18520 = \sport0_txctl_TX_reg[4]/P0001  & n18519 ;
  assign n18522 = ~\sport0_txctl_ldTX_cmp_reg/P0001  & ~n18520 ;
  assign n18523 = ~n18521 & n18522 ;
  assign n18524 = ~n18517 & ~n18523 ;
  assign n18525 = \core_c_psq_ststk_sts7x23_STcell_reg[1][7]/P0001  & ~n18362 ;
  assign n18526 = \core_eu_ec_cun_SS_reg/P0001  & n18362 ;
  assign n18527 = ~n18525 & ~n18526 ;
  assign n18528 = \core_c_psq_ststk_sts7x23_STcell_reg[1][6]/P0001  & ~n18362 ;
  assign n18529 = ~n4174 & n18362 ;
  assign n18530 = ~n18528 & ~n18529 ;
  assign n18531 = \core_c_psq_ststk_sts7x23_STcell_reg[1][5]/P0001  & ~n18362 ;
  assign n18532 = \core_eu_ec_cun_AQ_reg/P0001  & n18362 ;
  assign n18533 = ~n18531 & ~n18532 ;
  assign n18534 = \core_c_psq_ststk_sts7x23_STcell_reg[1][4]/P0001  & ~n18362 ;
  assign n18535 = \core_eu_ec_cun_AS_reg/P0001  & n18362 ;
  assign n18536 = ~n18534 & ~n18535 ;
  assign n18537 = \core_c_psq_ststk_sts7x23_STcell_reg[1][3]/P0001  & ~n18362 ;
  assign n18538 = \core_eu_ec_cun_AC_reg/P0001  & n18362 ;
  assign n18539 = ~n18537 & ~n18538 ;
  assign n18540 = \core_c_psq_ststk_sts7x23_STcell_reg[1][2]/P0001  & ~n18362 ;
  assign n18541 = \core_eu_ec_cun_AV_reg/P0001  & n18362 ;
  assign n18542 = ~n18540 & ~n18541 ;
  assign n18543 = \core_c_psq_ststk_sts7x23_STcell_reg[1][24]/P0001  & ~n18362 ;
  assign n18544 = \core_c_psq_IMASK_reg[9]/NET0131  & n18362 ;
  assign n18545 = ~n18543 & ~n18544 ;
  assign n18546 = \core_c_psq_ststk_sts7x23_STcell_reg[1][23]/P0001  & ~n18362 ;
  assign n18547 = \core_c_psq_IMASK_reg[8]/NET0131  & n18362 ;
  assign n18548 = ~n18546 & ~n18547 ;
  assign n18549 = \core_c_psq_ststk_sts7x23_STcell_reg[1][22]/P0001  & ~n18362 ;
  assign n18550 = \core_c_psq_IMASK_reg[7]/NET0131  & n18362 ;
  assign n18551 = ~n18549 & ~n18550 ;
  assign n18552 = \core_c_psq_ststk_sts7x23_STcell_reg[1][21]/P0001  & ~n18362 ;
  assign n18553 = \core_c_psq_IMASK_reg[6]/NET0131  & n18362 ;
  assign n18554 = ~n18552 & ~n18553 ;
  assign n18555 = \core_c_psq_ststk_sts7x23_STcell_reg[1][20]/P0001  & ~n18362 ;
  assign n18556 = \core_c_psq_IMASK_reg[5]/NET0131  & n18362 ;
  assign n18557 = ~n18555 & ~n18556 ;
  assign n18558 = \core_c_psq_ststk_sts7x23_STcell_reg[1][1]/P0001  & ~n18362 ;
  assign n18559 = \core_eu_ec_cun_AN_reg/P0001  & n18362 ;
  assign n18560 = ~n18558 & ~n18559 ;
  assign n18561 = \core_c_psq_ststk_sts7x23_STcell_reg[1][19]/P0001  & ~n18362 ;
  assign n18562 = \core_c_psq_IMASK_reg[4]/NET0131  & n18362 ;
  assign n18563 = ~n18561 & ~n18562 ;
  assign n18564 = \core_c_psq_ststk_sts7x23_STcell_reg[1][18]/P0001  & ~n18362 ;
  assign n18565 = \core_c_psq_IMASK_reg[3]/NET0131  & n18362 ;
  assign n18566 = ~n18564 & ~n18565 ;
  assign n18567 = \core_c_psq_ststk_sts7x23_STcell_reg[1][17]/P0001  & ~n18362 ;
  assign n18568 = \core_c_psq_IMASK_reg[2]/NET0131  & n18362 ;
  assign n18569 = ~n18567 & ~n18568 ;
  assign n18570 = \core_c_psq_ststk_sts7x23_STcell_reg[1][16]/P0001  & ~n18362 ;
  assign n18571 = \core_c_psq_IMASK_reg[1]/NET0131  & n18362 ;
  assign n18572 = ~n18570 & ~n18571 ;
  assign n18573 = \core_c_psq_ststk_sts7x23_STcell_reg[1][15]/P0001  & ~n18362 ;
  assign n18574 = \core_c_psq_IMASK_reg[0]/NET0131  & n18362 ;
  assign n18575 = ~n18573 & ~n18574 ;
  assign n18576 = \core_c_psq_ststk_sts7x23_STcell_reg[1][14]/P0001  & ~n18362 ;
  assign n18577 = \core_c_psq_MSTAT_reg_DO_reg[6]/NET0131  & n18362 ;
  assign n18578 = ~n18576 & ~n18577 ;
  assign n18579 = \core_c_psq_ststk_sts7x23_STcell_reg[1][13]/P0001  & ~n18362 ;
  assign n18580 = \core_c_psq_MSTAT_reg_DO_reg[5]/NET0131  & n18362 ;
  assign n18581 = ~n18579 & ~n18580 ;
  assign n18582 = \core_c_psq_ststk_sts7x23_STcell_reg[1][12]/P0001  & ~n18362 ;
  assign n18583 = \core_c_psq_MSTAT_reg_DO_reg[4]/NET0131  & n18362 ;
  assign n18584 = ~n18582 & ~n18583 ;
  assign n18585 = \core_c_psq_ststk_sts7x23_STcell_reg[1][11]/P0001  & ~n18362 ;
  assign n18586 = \core_c_psq_MSTAT_reg_DO_reg[3]/NET0131  & n18362 ;
  assign n18587 = ~n18585 & ~n18586 ;
  assign n18588 = \core_c_psq_ststk_sts7x23_STcell_reg[1][10]/P0001  & ~n18362 ;
  assign n18589 = \core_c_psq_MSTAT_reg_DO_reg[2]/NET0131  & n18362 ;
  assign n18590 = ~n18588 & ~n18589 ;
  assign n18591 = \core_c_psq_ststk_sts7x23_STcell_reg[1][0]/P0001  & ~n18362 ;
  assign n18592 = \core_eu_ec_cun_AZ_reg/P0001  & n18362 ;
  assign n18593 = ~n18591 & ~n18592 ;
  assign n18594 = n14695 & ~n18220 ;
  assign n18595 = \core_c_psq_ststk_sts7x23_STcell_reg[0][9]/P0001  & ~n18594 ;
  assign n18596 = \core_c_psq_MSTAT_reg_DO_reg[1]/NET0131  & n18594 ;
  assign n18597 = ~n18595 & ~n18596 ;
  assign n18598 = \core_c_psq_ststk_sts7x23_STcell_reg[0][8]/P0001  & ~n18594 ;
  assign n18599 = \core_c_psq_MSTAT_reg_DO_reg[0]/P0002  & n18594 ;
  assign n18600 = ~n18598 & ~n18599 ;
  assign n18601 = \core_c_psq_ststk_sts7x23_STcell_reg[0][7]/P0001  & ~n18594 ;
  assign n18602 = \core_eu_ec_cun_SS_reg/P0001  & n18594 ;
  assign n18603 = ~n18601 & ~n18602 ;
  assign n18604 = \core_c_psq_ststk_sts7x23_STcell_reg[0][6]/P0001  & ~n18594 ;
  assign n18605 = ~n4174 & n18594 ;
  assign n18606 = ~n18604 & ~n18605 ;
  assign n18607 = \core_c_psq_ststk_sts7x23_STcell_reg[0][5]/P0001  & ~n18594 ;
  assign n18608 = \core_eu_ec_cun_AQ_reg/P0001  & n18594 ;
  assign n18609 = ~n18607 & ~n18608 ;
  assign n18610 = \core_c_psq_ststk_sts7x23_STcell_reg[0][4]/P0001  & ~n18594 ;
  assign n18611 = \core_eu_ec_cun_AS_reg/P0001  & n18594 ;
  assign n18612 = ~n18610 & ~n18611 ;
  assign n18613 = \core_c_psq_ststk_sts7x23_STcell_reg[0][3]/P0001  & ~n18594 ;
  assign n18614 = \core_eu_ec_cun_AC_reg/P0001  & n18594 ;
  assign n18615 = ~n18613 & ~n18614 ;
  assign n18616 = \core_c_psq_ststk_sts7x23_STcell_reg[0][2]/P0001  & ~n18594 ;
  assign n18617 = \core_eu_ec_cun_AV_reg/P0001  & n18594 ;
  assign n18618 = ~n18616 & ~n18617 ;
  assign n18619 = \core_c_psq_ststk_sts7x23_STcell_reg[0][24]/P0001  & ~n18594 ;
  assign n18620 = \core_c_psq_IMASK_reg[9]/NET0131  & n18594 ;
  assign n18621 = ~n18619 & ~n18620 ;
  assign n18622 = \core_c_psq_ststk_sts7x23_STcell_reg[0][23]/P0001  & ~n18594 ;
  assign n18623 = \core_c_psq_IMASK_reg[8]/NET0131  & n18594 ;
  assign n18624 = ~n18622 & ~n18623 ;
  assign n18625 = \core_c_psq_ststk_sts7x23_STcell_reg[0][22]/P0001  & ~n18594 ;
  assign n18626 = \core_c_psq_IMASK_reg[7]/NET0131  & n18594 ;
  assign n18627 = ~n18625 & ~n18626 ;
  assign n18628 = \core_c_psq_ststk_sts7x23_STcell_reg[0][21]/P0001  & ~n18594 ;
  assign n18629 = \core_c_psq_IMASK_reg[6]/NET0131  & n18594 ;
  assign n18630 = ~n18628 & ~n18629 ;
  assign n18631 = \core_c_psq_ststk_sts7x23_STcell_reg[0][20]/P0001  & ~n18594 ;
  assign n18632 = \core_c_psq_IMASK_reg[5]/NET0131  & n18594 ;
  assign n18633 = ~n18631 & ~n18632 ;
  assign n18634 = \core_c_psq_ststk_sts7x23_STcell_reg[0][1]/P0001  & ~n18594 ;
  assign n18635 = \core_eu_ec_cun_AN_reg/P0001  & n18594 ;
  assign n18636 = ~n18634 & ~n18635 ;
  assign n18637 = \core_c_psq_ststk_sts7x23_STcell_reg[0][19]/P0001  & ~n18594 ;
  assign n18638 = \core_c_psq_IMASK_reg[4]/NET0131  & n18594 ;
  assign n18639 = ~n18637 & ~n18638 ;
  assign n18640 = \core_c_psq_ststk_sts7x23_STcell_reg[0][18]/P0001  & ~n18594 ;
  assign n18641 = \core_c_psq_IMASK_reg[3]/NET0131  & n18594 ;
  assign n18642 = ~n18640 & ~n18641 ;
  assign n18643 = \core_c_psq_ststk_sts7x23_STcell_reg[0][17]/P0001  & ~n18594 ;
  assign n18644 = \core_c_psq_IMASK_reg[2]/NET0131  & n18594 ;
  assign n18645 = ~n18643 & ~n18644 ;
  assign n18646 = \core_c_psq_ststk_sts7x23_STcell_reg[0][16]/P0001  & ~n18594 ;
  assign n18647 = \core_c_psq_IMASK_reg[1]/NET0131  & n18594 ;
  assign n18648 = ~n18646 & ~n18647 ;
  assign n18649 = \core_c_psq_ststk_sts7x23_STcell_reg[0][15]/P0001  & ~n18594 ;
  assign n18650 = \core_c_psq_IMASK_reg[0]/NET0131  & n18594 ;
  assign n18651 = ~n18649 & ~n18650 ;
  assign n18652 = n7284 & n18227 ;
  assign n18653 = ~n18232 & ~n18652 ;
  assign n18654 = \sport0_regs_FSDIVreg_DO_reg[9]/NET0131  & n18653 ;
  assign n18655 = ~n18236 & n18652 ;
  assign n18656 = n10289 & n18655 ;
  assign n18657 = ~n18654 & ~n18656 ;
  assign n18658 = \core_c_psq_ststk_sts7x23_STcell_reg[0][14]/P0001  & ~n18594 ;
  assign n18659 = \core_c_psq_MSTAT_reg_DO_reg[6]/NET0131  & n18594 ;
  assign n18660 = ~n18658 & ~n18659 ;
  assign n18661 = \core_c_psq_ststk_sts7x23_STcell_reg[0][13]/P0001  & ~n18594 ;
  assign n18662 = \core_c_psq_MSTAT_reg_DO_reg[5]/NET0131  & n18594 ;
  assign n18663 = ~n18661 & ~n18662 ;
  assign n18664 = \core_c_psq_ststk_sts7x23_STcell_reg[0][12]/P0001  & ~n18594 ;
  assign n18665 = \core_c_psq_MSTAT_reg_DO_reg[4]/NET0131  & n18594 ;
  assign n18666 = ~n18664 & ~n18665 ;
  assign n18667 = \core_c_psq_ststk_sts7x23_STcell_reg[0][11]/P0001  & ~n18594 ;
  assign n18668 = \core_c_psq_MSTAT_reg_DO_reg[3]/NET0131  & n18594 ;
  assign n18669 = ~n18667 & ~n18668 ;
  assign n18670 = \sport0_regs_FSDIVreg_DO_reg[8]/NET0131  & n18653 ;
  assign n18671 = n10638 & n18655 ;
  assign n18672 = ~n18670 & ~n18671 ;
  assign n18673 = \core_c_psq_ststk_sts7x23_STcell_reg[0][10]/P0001  & ~n18594 ;
  assign n18674 = \core_c_psq_MSTAT_reg_DO_reg[2]/NET0131  & n18594 ;
  assign n18675 = ~n18673 & ~n18674 ;
  assign n18676 = \core_c_psq_ststk_sts7x23_STcell_reg[0][0]/P0001  & ~n18594 ;
  assign n18677 = \core_eu_ec_cun_AZ_reg/P0001  & n18594 ;
  assign n18678 = ~n18676 & ~n18677 ;
  assign n18679 = n14694 & ~n18220 ;
  assign n18680 = ~n5950 & ~n14692 ;
  assign n18681 = n14696 & n18680 ;
  assign n18682 = n14701 & n18220 ;
  assign n18683 = n18681 & n18682 ;
  assign n18684 = ~n18679 & ~n18683 ;
  assign n18685 = \core_c_psq_ststk_ptr_reg[2]/NET0131  & n18684 ;
  assign n18686 = ~\core_c_psq_ststk_ptr_reg[2]/NET0131  & ~n18684 ;
  assign n18687 = ~n18685 & ~n18686 ;
  assign n18688 = ~n14711 & ~n18220 ;
  assign n18689 = ~n18681 & ~n18688 ;
  assign n18690 = ~\core_c_psq_ststk_ptr_reg[0]/NET0131  & ~n18689 ;
  assign n18691 = \core_c_psq_ststk_ptr_reg[0]/NET0131  & n18689 ;
  assign n18692 = ~n18690 & ~n18691 ;
  assign n18693 = \sport0_regs_FSDIVreg_DO_reg[14]/NET0131  & n18653 ;
  assign n18694 = n12688 & n18655 ;
  assign n18695 = ~n18693 & ~n18694 ;
  assign n18696 = ~n13806 & ~n14551 ;
  assign n18697 = n13806 & ~n14413 ;
  assign n18698 = ~n18696 & ~n18697 ;
  assign n18699 = n14667 & ~n18698 ;
  assign n18700 = \core_eu_ea_alu_ea_reg_afswe_DO_reg[13]/P0001  & ~n14667 ;
  assign n18701 = ~n18699 & ~n18700 ;
  assign n18702 = \sport0_regs_FSDIVreg_DO_reg[13]/NET0131  & n18653 ;
  assign n18703 = n7340 & n18655 ;
  assign n18704 = ~n18702 & ~n18703 ;
  assign n18705 = \sport0_regs_FSDIVreg_DO_reg[15]/NET0131  & n18653 ;
  assign n18706 = n12743 & n18655 ;
  assign n18707 = ~n18705 & ~n18706 ;
  assign n18708 = \sport0_regs_FSDIVreg_DO_reg[12]/NET0131  & n18653 ;
  assign n18709 = n9178 & n18655 ;
  assign n18710 = ~n18708 & ~n18709 ;
  assign n18711 = \sport0_regs_FSDIVreg_DO_reg[11]/NET0131  & n18653 ;
  assign n18712 = n8460 & n18655 ;
  assign n18713 = ~n18711 & ~n18712 ;
  assign n18714 = \sport0_regs_FSDIVreg_DO_reg[10]/NET0131  & n18653 ;
  assign n18715 = n7859 & n18655 ;
  assign n18716 = ~n18714 & ~n18715 ;
  assign n18717 = n14666 & ~n17832 ;
  assign n18718 = \core_c_dec_MTSR1_E_reg/P0001  & ~n18276 ;
  assign n18793 = n17954 & n17979 ;
  assign n18794 = ~n18151 & ~n18793 ;
  assign n18795 = n17945 & ~n18794 ;
  assign n18796 = n18015 & ~n18795 ;
  assign n18797 = ~n18018 & n18796 ;
  assign n18798 = ~n17964 & ~n18085 ;
  assign n18799 = n18797 & n18798 ;
  assign n18800 = ~n18060 & n18799 ;
  assign n18722 = n17931 & ~n18161 ;
  assign n18723 = ~n17922 & n18722 ;
  assign n18732 = n17931 & n18090 ;
  assign n18733 = ~n18182 & n18732 ;
  assign n18814 = ~n18723 & ~n18733 ;
  assign n18739 = n18147 & ~n18170 ;
  assign n18740 = n17839 & ~n18127 ;
  assign n18741 = ~n17929 & n18740 ;
  assign n18742 = n17931 & ~n18098 ;
  assign n18743 = ~n18741 & ~n18742 ;
  assign n18744 = ~n18133 & ~n18743 ;
  assign n18815 = ~n18739 & ~n18744 ;
  assign n18819 = n18814 & n18815 ;
  assign n18754 = n17929 & n18183 ;
  assign n18755 = n18089 & n18754 ;
  assign n18756 = ~n17929 & n18187 ;
  assign n18757 = n17921 & n18756 ;
  assign n18803 = ~n18755 & ~n18757 ;
  assign n18763 = n17929 & n18124 ;
  assign n18764 = n18106 & n18763 ;
  assign n18765 = n17839 & ~n18175 ;
  assign n18766 = ~n17929 & n18765 ;
  assign n18767 = n18055 & n18766 ;
  assign n18804 = ~n18764 & ~n18767 ;
  assign n18805 = n18803 & n18804 ;
  assign n18772 = \core_c_dec_IRE_reg[11]/NET0131  & ~n11311 ;
  assign n18801 = ~n18002 & ~n18772 ;
  assign n18748 = n17839 & ~n17933 ;
  assign n18749 = ~n17929 & n18748 ;
  assign n18750 = n18153 & n18749 ;
  assign n18751 = n17839 & ~n18102 ;
  assign n18752 = ~n17929 & n18751 ;
  assign n18753 = n18178 & n18752 ;
  assign n18802 = ~n18750 & ~n18753 ;
  assign n18806 = n18801 & n18802 ;
  assign n18812 = n18805 & n18806 ;
  assign n18813 = n17978 & n18054 ;
  assign n18820 = n18812 & n18813 ;
  assign n18824 = n18819 & n18820 ;
  assign n18734 = ~n17991 & ~n17997 ;
  assign n18735 = n17945 & ~n18734 ;
  assign n18736 = ~n17968 & ~n17993 ;
  assign n18737 = n17945 & ~n18736 ;
  assign n18738 = ~n18735 & ~n18737 ;
  assign n18745 = n17839 & ~n18165 ;
  assign n18746 = ~n17929 & n18745 ;
  assign n18747 = ~n18108 & n18746 ;
  assign n18758 = n17839 & ~n18135 ;
  assign n18759 = ~n17929 & n18758 ;
  assign n18760 = ~n18091 & n18759 ;
  assign n18816 = ~n18747 & ~n18760 ;
  assign n18768 = n18139 & n18765 ;
  assign n18769 = n18043 & n18115 ;
  assign n18817 = ~n18768 & ~n18769 ;
  assign n18818 = n18816 & n18817 ;
  assign n18825 = n18738 & n18818 ;
  assign n18826 = n18824 & n18825 ;
  assign n18774 = n17929 & n18055 ;
  assign n18775 = ~n18071 & ~n18774 ;
  assign n18776 = ~n17924 & ~n18775 ;
  assign n18777 = ~n17933 & n18070 ;
  assign n18778 = ~n18776 & ~n18777 ;
  assign n18779 = n17839 & ~n18778 ;
  assign n18792 = n18148 & ~n18170 ;
  assign n18783 = n17965 & n18021 ;
  assign n18784 = n18179 & n18752 ;
  assign n18809 = ~n18783 & ~n18784 ;
  assign n18810 = ~n18792 & n18809 ;
  assign n18761 = ~n17929 & n17986 ;
  assign n18762 = n18115 & n18761 ;
  assign n18770 = n17959 & n18112 ;
  assign n18807 = ~n18762 & ~n18770 ;
  assign n18771 = n17915 & n18756 ;
  assign n18773 = n18107 & n18763 ;
  assign n18808 = ~n18771 & ~n18773 ;
  assign n18811 = n18807 & n18808 ;
  assign n18821 = n18810 & n18811 ;
  assign n18719 = n17931 & n18153 ;
  assign n18720 = ~n18046 & ~n18719 ;
  assign n18721 = n18111 & ~n18720 ;
  assign n18780 = n17931 & n18056 ;
  assign n18781 = ~n17980 & ~n18780 ;
  assign n18782 = n18088 & ~n18781 ;
  assign n18822 = ~n18721 & ~n18782 ;
  assign n18823 = n18821 & n18822 ;
  assign n18827 = ~n18779 & n18823 ;
  assign n18828 = n18826 & n18827 ;
  assign n18724 = ~n18032 & n18145 ;
  assign n18725 = n18020 & n18025 ;
  assign n18726 = n18724 & ~n18725 ;
  assign n18727 = n18038 & ~n18141 ;
  assign n18728 = ~n18040 & ~n18069 ;
  assign n18729 = n18195 & n18728 ;
  assign n18730 = n18727 & n18729 ;
  assign n18731 = n18726 & n18730 ;
  assign n18785 = n17965 & n18056 ;
  assign n18786 = n17945 & n18150 ;
  assign n18787 = ~n17929 & n18026 ;
  assign n18788 = ~n18010 & ~n18023 ;
  assign n18789 = ~n18787 & n18788 ;
  assign n18790 = ~n18786 & n18789 ;
  assign n18791 = ~n18785 & n18790 ;
  assign n18829 = n18731 & n18791 ;
  assign n18830 = n18828 & n18829 ;
  assign n18831 = n18800 & n18830 ;
  assign n18832 = ~\core_c_dec_MTSR1_E_reg/P0001  & n18831 ;
  assign n18833 = ~n18718 & ~n18832 ;
  assign n18834 = n18717 & ~n18833 ;
  assign n18835 = ~\core_eu_es_sht_es_reg_sr1swe_DO_reg[6]/P0001  & ~n18717 ;
  assign n18836 = ~n18834 & ~n18835 ;
  assign n18837 = \core_c_dec_updMR_E_reg/P0001  & n4118 ;
  assign n18838 = ~n6023 & ~n6108 ;
  assign n18839 = n6022 & n6117 ;
  assign n18840 = ~n13577 & ~n18839 ;
  assign n18841 = ~n14728 & n18840 ;
  assign n18842 = n18838 & n18841 ;
  assign n18843 = ~\core_c_dec_IR_reg[15]/NET0131  & ~\core_c_dec_IR_reg[16]/NET0131  ;
  assign n18844 = ~\core_c_dec_IR_reg[13]/NET0131  & ~\core_c_dec_IR_reg[14]/NET0131  ;
  assign n18845 = n18843 & n18844 ;
  assign n18846 = ~\core_c_dec_IR_reg[17]/NET0131  & ~n18845 ;
  assign n18847 = ~n18842 & n18846 ;
  assign n18848 = ~n4117 & n18847 ;
  assign n18849 = \core_c_dec_IR_reg[18]/NET0131  & ~n6023 ;
  assign n18850 = n4116 & ~n18849 ;
  assign n18851 = n18848 & n18850 ;
  assign n18852 = ~n18837 & ~n18851 ;
  assign n18853 = n13805 & ~n18698 ;
  assign n18854 = \core_eu_ea_alu_ea_reg_afrwe_DO_reg[13]/P0001  & ~n13805 ;
  assign n18855 = ~n18853 & ~n18854 ;
  assign n18856 = \sice_ICYC_reg[0]/NET0131  & \sice_ICYC_reg[1]/NET0131  ;
  assign n18857 = \sice_ICYC_reg[2]/NET0131  & n18856 ;
  assign n18858 = \sice_ICYC_reg[3]/NET0131  & n18857 ;
  assign n18859 = \sice_ICYC_reg[4]/NET0131  & n18858 ;
  assign n18860 = \sice_ICYC_reg[5]/NET0131  & n18859 ;
  assign n18861 = \sice_ICYC_reg[6]/NET0131  & n18860 ;
  assign n18862 = ~\sice_ICYC_reg[7]/NET0131  & ~n18861 ;
  assign n18863 = \sice_ICYC_reg[7]/NET0131  & n18861 ;
  assign n18864 = ~n18862 & ~n18863 ;
  assign n18865 = \sice_IIRC_reg[0]/NET0131  & \sice_IIRC_reg[1]/NET0131  ;
  assign n18866 = \sice_IIRC_reg[2]/NET0131  & n18865 ;
  assign n18867 = \sice_IIRC_reg[3]/NET0131  & n18866 ;
  assign n18868 = \sice_IIRC_reg[4]/NET0131  & n18867 ;
  assign n18869 = \sice_IIRC_reg[5]/NET0131  & n18868 ;
  assign n18870 = \sice_IIRC_reg[6]/NET0131  & n18869 ;
  assign n18871 = \sice_IIRC_reg[7]/NET0131  & n18870 ;
  assign n18872 = ~\sice_IIRC_reg[7]/NET0131  & ~n18870 ;
  assign n18873 = ~n18871 & ~n18872 ;
  assign n18874 = \core_eu_em_mac_em_dec_emcorepi_DO_reg[3]/P0001  & ~n18848 ;
  assign n18875 = \core_c_dec_IR_reg[14]/NET0131  & ~n18843 ;
  assign n18876 = n18848 & n18875 ;
  assign n18877 = ~n18874 & ~n18876 ;
  assign n18878 = \core_eu_em_mac_em_dec_emcorepi_DO_reg[2]/P0001  & ~n18848 ;
  assign n18879 = \core_c_dec_IR_reg[13]/NET0131  & ~n18843 ;
  assign n18880 = n18848 & n18879 ;
  assign n18881 = ~n18878 & ~n18880 ;
  assign n18882 = n17833 & ~n18833 ;
  assign n18883 = ~\core_eu_es_sht_es_reg_sr1rwe_DO_reg[6]/P0001  & ~n17833 ;
  assign n18884 = ~n18882 & ~n18883 ;
  assign n18885 = ~\core_c_dec_MTSR0_E_reg/P0001  & ~\core_c_dec_updSR_E_reg/P0001  ;
  assign n18886 = n14666 & ~n18885 ;
  assign n18887 = \core_c_dec_MTSR0_E_reg/P0001  & ~n18276 ;
  assign n18921 = ~n18079 & n18749 ;
  assign n18912 = ~n17955 & ~n18072 ;
  assign n18917 = n18763 & ~n18912 ;
  assign n18918 = ~n18039 & ~n18191 ;
  assign n18919 = ~n18722 & ~n18756 ;
  assign n18920 = ~n18918 & ~n18919 ;
  assign n18929 = ~n18917 & ~n18920 ;
  assign n18930 = ~n18921 & n18929 ;
  assign n18907 = ~n17952 & ~n18001 ;
  assign n18908 = ~n18743 & ~n18907 ;
  assign n18909 = ~n18029 & ~n18036 ;
  assign n18910 = n18766 & ~n18909 ;
  assign n18927 = ~n18908 & ~n18910 ;
  assign n18913 = n18746 & ~n18912 ;
  assign n18914 = ~n18033 & ~n18067 ;
  assign n18915 = ~n18754 & ~n18759 ;
  assign n18916 = ~n18914 & ~n18915 ;
  assign n18928 = ~n18913 & ~n18916 ;
  assign n18931 = n18927 & n18928 ;
  assign n18888 = ~n17960 & ~n18150 ;
  assign n18889 = n18088 & ~n18888 ;
  assign n18905 = n17931 & ~n18110 ;
  assign n18906 = ~n18079 & n18905 ;
  assign n18911 = \core_c_dec_IRE_reg[11]/NET0131  & ~n11315 ;
  assign n18925 = ~n18018 & ~n18911 ;
  assign n18926 = ~n18906 & n18925 ;
  assign n18932 = ~n18889 & n18926 ;
  assign n18936 = n18931 & n18932 ;
  assign n18937 = n18930 & n18936 ;
  assign n18900 = n17959 & n17965 ;
  assign n18901 = ~n17972 & ~n18900 ;
  assign n18902 = ~n18143 & ~n18783 ;
  assign n18903 = n18901 & n18902 ;
  assign n18904 = n18789 & n18903 ;
  assign n18890 = n17971 & ~n18082 ;
  assign n18891 = ~n17995 & ~n18890 ;
  assign n18892 = n18796 & n18891 ;
  assign n18893 = n17958 & n17989 ;
  assign n18894 = ~n17931 & n18056 ;
  assign n18895 = ~n18893 & ~n18894 ;
  assign n18896 = n18751 & ~n18895 ;
  assign n18897 = ~n17931 & n17968 ;
  assign n18898 = ~n18027 & ~n18897 ;
  assign n18899 = n18115 & ~n18898 ;
  assign n18933 = ~n18896 & ~n18899 ;
  assign n18922 = n17931 & ~n18909 ;
  assign n18923 = ~n17924 & n18922 ;
  assign n18924 = ~n17998 & n18171 ;
  assign n18934 = ~n18923 & ~n18924 ;
  assign n18935 = n18933 & n18934 ;
  assign n18938 = n18892 & n18935 ;
  assign n18939 = n18904 & n18938 ;
  assign n18940 = n18937 & n18939 ;
  assign n18941 = ~\core_c_dec_MTSR0_E_reg/P0001  & n18940 ;
  assign n18942 = ~n18887 & ~n18941 ;
  assign n18943 = n18886 & ~n18942 ;
  assign n18944 = ~\core_eu_es_sht_es_reg_sr0swe_DO_reg[6]/P0001  & ~n18886 ;
  assign n18945 = ~n18943 & ~n18944 ;
  assign n18946 = n7270 & n18227 ;
  assign n18947 = \sport1_regs_MWORDreg_DO_reg[7]/NET0131  & ~n18946 ;
  assign n18948 = ~n12688 & n18946 ;
  assign n18949 = n11265 & n18948 ;
  assign n18950 = ~n18947 & ~n18949 ;
  assign n18951 = \sport1_regs_MWORDreg_DO_reg[6]/NET0131  & ~n18946 ;
  assign n18952 = n11525 & n18948 ;
  assign n18953 = ~n18951 & ~n18952 ;
  assign n18954 = \sport1_regs_MWORDreg_DO_reg[5]/NET0131  & ~n18946 ;
  assign n18955 = n10911 & n18948 ;
  assign n18956 = ~n18954 & ~n18955 ;
  assign n18957 = ~n7340 & n18946 ;
  assign n18958 = ~\sport1_regs_MWORDreg_DO_reg[8]/NET0131  & ~n18946 ;
  assign n18959 = ~n18957 & ~n18958 ;
  assign n18960 = \sport1_regs_MWORDreg_DO_reg[4]/NET0131  & ~n18946 ;
  assign n18961 = n10069 & n18948 ;
  assign n18962 = ~n18960 & ~n18961 ;
  assign n18963 = \sport1_regs_MWORDreg_DO_reg[1]/NET0131  & ~n18946 ;
  assign n18964 = n9435 & n18948 ;
  assign n18965 = ~n18963 & ~n18964 ;
  assign n18966 = \sport1_regs_MWORDreg_DO_reg[0]/NET0131  & ~n18946 ;
  assign n18967 = n7607 & n18948 ;
  assign n18968 = ~n18966 & ~n18967 ;
  assign n18969 = ~n7340 & n18231 ;
  assign n18970 = ~\sport0_regs_MWORDreg_DO_reg[8]/NET0131  & ~n18231 ;
  assign n18971 = ~n18969 & ~n18970 ;
  assign n18972 = ~\core_c_dec_accPM_E_reg/P0001  & ~n9435 ;
  assign n18973 = \core_c_dec_accPM_E_reg/P0001  & ~n12802 ;
  assign n18974 = ~n18972 & ~n18973 ;
  assign n18975 = \core_c_dec_MTSR0_E_reg/P0001  & ~n18974 ;
  assign n18983 = ~n18022 & ~n18793 ;
  assign n18984 = n18765 & ~n18983 ;
  assign n18985 = ~n17998 & ~n18165 ;
  assign n19002 = ~n18984 & ~n18985 ;
  assign n18986 = ~n17933 & n18083 ;
  assign n18989 = n18162 & ~n18898 ;
  assign n19003 = ~n18986 & ~n18989 ;
  assign n19004 = n19002 & n19003 ;
  assign n18978 = \core_c_dec_IRE_reg[11]/NET0131  & ~n9276 ;
  assign n18994 = ~n18143 & ~n18978 ;
  assign n18995 = n18901 & n18994 ;
  assign n18976 = n17930 & ~n18082 ;
  assign n18977 = ~n18129 & ~n18914 ;
  assign n18996 = ~n18976 & ~n18977 ;
  assign n19000 = n18995 & n18996 ;
  assign n18980 = n17954 & n17989 ;
  assign n18981 = ~n18044 & ~n18980 ;
  assign n18982 = n18088 & ~n18981 ;
  assign n19001 = n18019 & ~n18982 ;
  assign n19005 = n19000 & n19001 ;
  assign n18987 = ~n17961 & ~n18150 ;
  assign n18988 = ~n18114 & ~n18987 ;
  assign n18979 = ~n18079 & ~n18189 ;
  assign n18990 = ~n18104 & ~n18918 ;
  assign n18997 = ~n18979 & ~n18990 ;
  assign n18991 = ~n18136 & ~n18172 ;
  assign n18992 = ~n18909 & ~n18991 ;
  assign n18993 = n17991 & n18111 ;
  assign n18998 = ~n18992 & ~n18993 ;
  assign n18999 = n18997 & n18998 ;
  assign n19006 = ~n18988 & n18999 ;
  assign n19007 = n19005 & n19006 ;
  assign n19008 = n19004 & n19007 ;
  assign n19009 = ~\core_c_dec_MTSR0_E_reg/P0001  & n19008 ;
  assign n19010 = ~n18975 & ~n19009 ;
  assign n19011 = n18886 & ~n19010 ;
  assign n19012 = ~\core_eu_es_sht_es_reg_sr0swe_DO_reg[1]/P0001  & ~n18886 ;
  assign n19013 = ~n19011 & ~n19012 ;
  assign n19014 = \sport0_regs_MWORDreg_DO_reg[7]/NET0131  & ~n18231 ;
  assign n19015 = ~n12688 & n18231 ;
  assign n19016 = n11265 & n19015 ;
  assign n19017 = ~n19014 & ~n19016 ;
  assign n19018 = \sport0_regs_MWORDreg_DO_reg[6]/NET0131  & ~n18231 ;
  assign n19019 = n11525 & n19015 ;
  assign n19020 = ~n19018 & ~n19019 ;
  assign n19021 = \sport0_regs_MWORDreg_DO_reg[5]/NET0131  & ~n18231 ;
  assign n19022 = n10911 & n19015 ;
  assign n19023 = ~n19021 & ~n19022 ;
  assign n19024 = n10069 & ~n18236 ;
  assign n19025 = n18231 & ~n19024 ;
  assign n19026 = ~\sport0_regs_MWORDreg_DO_reg[4]/NET0131  & ~n18231 ;
  assign n19027 = ~n19025 & ~n19026 ;
  assign n19028 = \sport0_regs_MWORDreg_DO_reg[1]/NET0131  & ~n18231 ;
  assign n19029 = n9435 & n19015 ;
  assign n19030 = ~n19028 & ~n19029 ;
  assign n19031 = \sport0_regs_MWORDreg_DO_reg[0]/NET0131  & ~n18231 ;
  assign n19032 = n7607 & n19015 ;
  assign n19033 = ~n19031 & ~n19032 ;
  assign n19034 = n13804 & ~n18885 ;
  assign n19035 = ~n18942 & n19034 ;
  assign n19036 = ~\core_eu_es_sht_es_reg_sr0rwe_DO_reg[6]/P0001  & ~n19034 ;
  assign n19037 = ~n19035 & ~n19036 ;
  assign n19038 = \memc_Dread_E_reg/NET0131  & n5435 ;
  assign n19039 = ~\memc_IOcmd_E_reg/NET0131  & ~n19038 ;
  assign n19040 = ~PM_bdry_sel_pad & ~\core_dag_ilm2reg_PMA_pi_DO_reg[12]/NET0131  ;
  assign n19041 = \core_dag_ilm2reg_PMA_pi_DO_reg[13]/NET0131  & ~n19040 ;
  assign n19042 = \core_c_dec_Double_E_reg/P0001  & \core_c_psq_PMOVL_regh_DO_reg[3]/NET0131  ;
  assign n19043 = n19041 & n19042 ;
  assign n19044 = \core_c_psq_PCS_reg[3]/NET0131  & ~n4068 ;
  assign n19045 = ~n5697 & ~n5712 ;
  assign n19046 = ~\core_c_psq_PCS_reg[3]/NET0131  & ~n19045 ;
  assign n19047 = ~n19044 & ~n19046 ;
  assign n19048 = ~\core_c_psq_ECYC_reg/P0001  & ~n14733 ;
  assign n19049 = ~n19047 & n19048 ;
  assign n19050 = ~n19043 & n19049 ;
  assign n19051 = ~n14733 & n19043 ;
  assign n19052 = n5560 & n19051 ;
  assign n19053 = n5598 & n19052 ;
  assign n19054 = ~n19050 & ~n19053 ;
  assign n19055 = ~n19039 & ~n19054 ;
  assign n19056 = ~n4117 & ~n14733 ;
  assign n19057 = \emc_DMDoe_reg/NET0131  & ~n19056 ;
  assign n19058 = n19054 & n19057 ;
  assign n19059 = ~n19055 & ~n19058 ;
  assign n19060 = ~n19010 & n19034 ;
  assign n19061 = ~\core_eu_es_sht_es_reg_sr0rwe_DO_reg[1]/P0001  & ~n19034 ;
  assign n19062 = ~n19060 & ~n19061 ;
  assign n19063 = ~\sport1_regs_MWORDreg_DO_reg[9]/NET0131  & ~n18946 ;
  assign n19064 = ~n18948 & ~n19063 ;
  assign n19065 = \sport0_regs_MWORDreg_DO_reg[9]/NET0131  & ~n18231 ;
  assign n19066 = ~n18232 & ~n19065 ;
  assign n19088 = \sport1_cfg_SCLKi_cnt_reg[1]/NET0131  & ~\sport1_regs_SCLKDIVreg_DO_reg[1]/NET0131  ;
  assign n19089 = ~\sport1_cfg_SCLKi_cnt_reg[13]/NET0131  & \sport1_regs_SCLKDIVreg_DO_reg[13]/NET0131  ;
  assign n19109 = ~n19088 & ~n19089 ;
  assign n19090 = \sport1_cfg_SCLKi_cnt_reg[9]/NET0131  & ~\sport1_regs_SCLKDIVreg_DO_reg[9]/NET0131  ;
  assign n19091 = ~\sport1_cfg_SCLKi_cnt_reg[0]/NET0131  & \sport1_regs_SCLKDIVreg_DO_reg[0]/NET0131  ;
  assign n19110 = ~n19090 & ~n19091 ;
  assign n19117 = n19109 & n19110 ;
  assign n19084 = ~\sport1_cfg_SCLKi_cnt_reg[1]/NET0131  & \sport1_regs_SCLKDIVreg_DO_reg[1]/NET0131  ;
  assign n19085 = \sport1_cfg_SCLKi_cnt_reg[0]/NET0131  & ~\sport1_regs_SCLKDIVreg_DO_reg[0]/NET0131  ;
  assign n19107 = ~n19084 & ~n19085 ;
  assign n19086 = ~\sport1_cfg_SCLKi_cnt_reg[14]/NET0131  & \sport1_regs_SCLKDIVreg_DO_reg[14]/NET0131  ;
  assign n19087 = \sport1_cfg_SCLKi_cnt_reg[14]/NET0131  & ~\sport1_regs_SCLKDIVreg_DO_reg[14]/NET0131  ;
  assign n19108 = ~n19086 & ~n19087 ;
  assign n19118 = n19107 & n19108 ;
  assign n19125 = n19117 & n19118 ;
  assign n19096 = ~\sport1_cfg_SCLKi_cnt_reg[8]/NET0131  & \sport1_regs_SCLKDIVreg_DO_reg[8]/NET0131  ;
  assign n19097 = \sport1_cfg_SCLKi_cnt_reg[8]/NET0131  & ~\sport1_regs_SCLKDIVreg_DO_reg[8]/NET0131  ;
  assign n19113 = ~n19096 & ~n19097 ;
  assign n19098 = \sport1_cfg_SCLKi_cnt_reg[3]/NET0131  & ~\sport1_regs_SCLKDIVreg_DO_reg[3]/NET0131  ;
  assign n19099 = ~\sport1_cfg_SCLKi_cnt_reg[3]/NET0131  & \sport1_regs_SCLKDIVreg_DO_reg[3]/NET0131  ;
  assign n19114 = ~n19098 & ~n19099 ;
  assign n19115 = n19113 & n19114 ;
  assign n19092 = ~\sport1_cfg_SCLKi_cnt_reg[12]/NET0131  & \sport1_regs_SCLKDIVreg_DO_reg[12]/NET0131  ;
  assign n19093 = \sport1_cfg_SCLKi_cnt_reg[6]/NET0131  & ~\sport1_regs_SCLKDIVreg_DO_reg[6]/NET0131  ;
  assign n19111 = ~n19092 & ~n19093 ;
  assign n19094 = \sport1_cfg_SCLKi_cnt_reg[12]/NET0131  & ~\sport1_regs_SCLKDIVreg_DO_reg[12]/NET0131  ;
  assign n19095 = ~\sport1_cfg_SCLKi_cnt_reg[4]/NET0131  & \sport1_regs_SCLKDIVreg_DO_reg[4]/NET0131  ;
  assign n19112 = ~n19094 & ~n19095 ;
  assign n19116 = n19111 & n19112 ;
  assign n19126 = n19115 & n19116 ;
  assign n19127 = n19125 & n19126 ;
  assign n19069 = ~\sport1_cfg_SCLKi_cnt_reg[6]/NET0131  & \sport1_regs_SCLKDIVreg_DO_reg[6]/NET0131  ;
  assign n19070 = \sport1_cfg_SCLKi_cnt_reg[2]/NET0131  & ~\sport1_regs_SCLKDIVreg_DO_reg[2]/NET0131  ;
  assign n19101 = ~n19069 & ~n19070 ;
  assign n19071 = \sport1_cfg_SCLKi_cnt_reg[15]/NET0131  & ~\sport1_regs_SCLKDIVreg_DO_reg[15]/NET0131  ;
  assign n19072 = \sport1_cfg_SCLKi_cnt_reg[13]/NET0131  & ~\sport1_regs_SCLKDIVreg_DO_reg[13]/NET0131  ;
  assign n19102 = ~n19071 & ~n19072 ;
  assign n19121 = n19101 & n19102 ;
  assign n19081 = ~\sport1_cfg_SCLKi_cnt_reg[7]/NET0131  & ~\sport1_regs_SCLKDIVreg_DO_reg[7]/NET0131  ;
  assign n19082 = \sport1_cfg_SCLKi_cnt_reg[7]/NET0131  & \sport1_regs_SCLKDIVreg_DO_reg[7]/NET0131  ;
  assign n19083 = ~n19081 & ~n19082 ;
  assign n19067 = ~\sport1_cfg_SCLKi_cnt_reg[15]/NET0131  & \sport1_regs_SCLKDIVreg_DO_reg[15]/NET0131  ;
  assign n19068 = ~\sport1_cfg_SCLKi_cnt_reg[5]/NET0131  & \sport1_regs_SCLKDIVreg_DO_reg[5]/NET0131  ;
  assign n19100 = ~n19067 & ~n19068 ;
  assign n19122 = ~n19083 & n19100 ;
  assign n19123 = n19121 & n19122 ;
  assign n19077 = ~\sport1_cfg_SCLKi_cnt_reg[9]/NET0131  & \sport1_regs_SCLKDIVreg_DO_reg[9]/NET0131  ;
  assign n19078 = \sport1_cfg_SCLKi_cnt_reg[4]/NET0131  & ~\sport1_regs_SCLKDIVreg_DO_reg[4]/NET0131  ;
  assign n19105 = ~n19077 & ~n19078 ;
  assign n19079 = ~\sport1_cfg_SCLKi_cnt_reg[2]/NET0131  & \sport1_regs_SCLKDIVreg_DO_reg[2]/NET0131  ;
  assign n19080 = \sport1_cfg_SCLKi_cnt_reg[11]/NET0131  & ~\sport1_regs_SCLKDIVreg_DO_reg[11]/NET0131  ;
  assign n19106 = ~n19079 & ~n19080 ;
  assign n19119 = n19105 & n19106 ;
  assign n19073 = \sport1_cfg_SCLKi_cnt_reg[10]/NET0131  & ~\sport1_regs_SCLKDIVreg_DO_reg[10]/NET0131  ;
  assign n19074 = ~\sport1_cfg_SCLKi_cnt_reg[11]/NET0131  & \sport1_regs_SCLKDIVreg_DO_reg[11]/NET0131  ;
  assign n19103 = ~n19073 & ~n19074 ;
  assign n19075 = ~\sport1_cfg_SCLKi_cnt_reg[10]/NET0131  & \sport1_regs_SCLKDIVreg_DO_reg[10]/NET0131  ;
  assign n19076 = \sport1_cfg_SCLKi_cnt_reg[5]/NET0131  & ~\sport1_regs_SCLKDIVreg_DO_reg[5]/NET0131  ;
  assign n19104 = ~n19075 & ~n19076 ;
  assign n19120 = n19103 & n19104 ;
  assign n19124 = n19119 & n19120 ;
  assign n19128 = n19123 & n19124 ;
  assign n19129 = n19127 & n19128 ;
  assign n19130 = \sport1_cfg_SP_ENg_reg/NET0131  & ~n19129 ;
  assign n19131 = ~\sport1_cfg_SCLKi_h_reg/NET0131  & ~n19130 ;
  assign n19132 = \sport1_cfg_SCLKi_h_reg/NET0131  & n19130 ;
  assign n19133 = ~n19131 & ~n19132 ;
  assign n19155 = \sport0_cfg_SCLKi_cnt_reg[13]/NET0131  & ~\sport0_regs_SCLKDIVreg_DO_reg[13]/NET0131  ;
  assign n19156 = ~\sport0_cfg_SCLKi_cnt_reg[5]/NET0131  & \sport0_regs_SCLKDIVreg_DO_reg[5]/NET0131  ;
  assign n19176 = ~n19155 & ~n19156 ;
  assign n19157 = \sport0_cfg_SCLKi_cnt_reg[1]/NET0131  & ~\sport0_regs_SCLKDIVreg_DO_reg[1]/NET0131  ;
  assign n19158 = ~\sport0_cfg_SCLKi_cnt_reg[12]/NET0131  & \sport0_regs_SCLKDIVreg_DO_reg[12]/NET0131  ;
  assign n19177 = ~n19157 & ~n19158 ;
  assign n19184 = n19176 & n19177 ;
  assign n19151 = ~\sport0_cfg_SCLKi_cnt_reg[13]/NET0131  & \sport0_regs_SCLKDIVreg_DO_reg[13]/NET0131  ;
  assign n19152 = \sport0_cfg_SCLKi_cnt_reg[12]/NET0131  & ~\sport0_regs_SCLKDIVreg_DO_reg[12]/NET0131  ;
  assign n19174 = ~n19151 & ~n19152 ;
  assign n19153 = ~\sport0_cfg_SCLKi_cnt_reg[6]/NET0131  & \sport0_regs_SCLKDIVreg_DO_reg[6]/NET0131  ;
  assign n19154 = \sport0_cfg_SCLKi_cnt_reg[6]/NET0131  & ~\sport0_regs_SCLKDIVreg_DO_reg[6]/NET0131  ;
  assign n19175 = ~n19153 & ~n19154 ;
  assign n19185 = n19174 & n19175 ;
  assign n19192 = n19184 & n19185 ;
  assign n19163 = ~\sport0_cfg_SCLKi_cnt_reg[0]/NET0131  & \sport0_regs_SCLKDIVreg_DO_reg[0]/NET0131  ;
  assign n19164 = \sport0_cfg_SCLKi_cnt_reg[0]/NET0131  & ~\sport0_regs_SCLKDIVreg_DO_reg[0]/NET0131  ;
  assign n19180 = ~n19163 & ~n19164 ;
  assign n19165 = \sport0_cfg_SCLKi_cnt_reg[15]/NET0131  & ~\sport0_regs_SCLKDIVreg_DO_reg[15]/NET0131  ;
  assign n19166 = ~\sport0_cfg_SCLKi_cnt_reg[15]/NET0131  & \sport0_regs_SCLKDIVreg_DO_reg[15]/NET0131  ;
  assign n19181 = ~n19165 & ~n19166 ;
  assign n19182 = n19180 & n19181 ;
  assign n19159 = ~\sport0_cfg_SCLKi_cnt_reg[4]/NET0131  & \sport0_regs_SCLKDIVreg_DO_reg[4]/NET0131  ;
  assign n19160 = \sport0_cfg_SCLKi_cnt_reg[10]/NET0131  & ~\sport0_regs_SCLKDIVreg_DO_reg[10]/NET0131  ;
  assign n19178 = ~n19159 & ~n19160 ;
  assign n19161 = \sport0_cfg_SCLKi_cnt_reg[4]/NET0131  & ~\sport0_regs_SCLKDIVreg_DO_reg[4]/NET0131  ;
  assign n19162 = ~\sport0_cfg_SCLKi_cnt_reg[8]/NET0131  & \sport0_regs_SCLKDIVreg_DO_reg[8]/NET0131  ;
  assign n19179 = ~n19161 & ~n19162 ;
  assign n19183 = n19178 & n19179 ;
  assign n19193 = n19182 & n19183 ;
  assign n19194 = n19192 & n19193 ;
  assign n19136 = ~\sport0_cfg_SCLKi_cnt_reg[10]/NET0131  & \sport0_regs_SCLKDIVreg_DO_reg[10]/NET0131  ;
  assign n19137 = \sport0_cfg_SCLKi_cnt_reg[14]/NET0131  & ~\sport0_regs_SCLKDIVreg_DO_reg[14]/NET0131  ;
  assign n19168 = ~n19136 & ~n19137 ;
  assign n19138 = \sport0_cfg_SCLKi_cnt_reg[7]/NET0131  & ~\sport0_regs_SCLKDIVreg_DO_reg[7]/NET0131  ;
  assign n19139 = \sport0_cfg_SCLKi_cnt_reg[5]/NET0131  & ~\sport0_regs_SCLKDIVreg_DO_reg[5]/NET0131  ;
  assign n19169 = ~n19138 & ~n19139 ;
  assign n19188 = n19168 & n19169 ;
  assign n19148 = ~\sport0_cfg_SCLKi_cnt_reg[11]/NET0131  & ~\sport0_regs_SCLKDIVreg_DO_reg[11]/NET0131  ;
  assign n19149 = \sport0_cfg_SCLKi_cnt_reg[11]/NET0131  & \sport0_regs_SCLKDIVreg_DO_reg[11]/NET0131  ;
  assign n19150 = ~n19148 & ~n19149 ;
  assign n19134 = ~\sport0_cfg_SCLKi_cnt_reg[7]/NET0131  & \sport0_regs_SCLKDIVreg_DO_reg[7]/NET0131  ;
  assign n19135 = ~\sport0_cfg_SCLKi_cnt_reg[9]/NET0131  & \sport0_regs_SCLKDIVreg_DO_reg[9]/NET0131  ;
  assign n19167 = ~n19134 & ~n19135 ;
  assign n19189 = ~n19150 & n19167 ;
  assign n19190 = n19188 & n19189 ;
  assign n19144 = ~\sport0_cfg_SCLKi_cnt_reg[1]/NET0131  & \sport0_regs_SCLKDIVreg_DO_reg[1]/NET0131  ;
  assign n19145 = \sport0_cfg_SCLKi_cnt_reg[8]/NET0131  & ~\sport0_regs_SCLKDIVreg_DO_reg[8]/NET0131  ;
  assign n19172 = ~n19144 & ~n19145 ;
  assign n19146 = ~\sport0_cfg_SCLKi_cnt_reg[14]/NET0131  & \sport0_regs_SCLKDIVreg_DO_reg[14]/NET0131  ;
  assign n19147 = \sport0_cfg_SCLKi_cnt_reg[3]/NET0131  & ~\sport0_regs_SCLKDIVreg_DO_reg[3]/NET0131  ;
  assign n19173 = ~n19146 & ~n19147 ;
  assign n19186 = n19172 & n19173 ;
  assign n19140 = \sport0_cfg_SCLKi_cnt_reg[2]/NET0131  & ~\sport0_regs_SCLKDIVreg_DO_reg[2]/NET0131  ;
  assign n19141 = ~\sport0_cfg_SCLKi_cnt_reg[3]/NET0131  & \sport0_regs_SCLKDIVreg_DO_reg[3]/NET0131  ;
  assign n19170 = ~n19140 & ~n19141 ;
  assign n19142 = ~\sport0_cfg_SCLKi_cnt_reg[2]/NET0131  & \sport0_regs_SCLKDIVreg_DO_reg[2]/NET0131  ;
  assign n19143 = \sport0_cfg_SCLKi_cnt_reg[9]/NET0131  & ~\sport0_regs_SCLKDIVreg_DO_reg[9]/NET0131  ;
  assign n19171 = ~n19142 & ~n19143 ;
  assign n19187 = n19170 & n19171 ;
  assign n19191 = n19186 & n19187 ;
  assign n19195 = n19190 & n19191 ;
  assign n19196 = n19194 & n19195 ;
  assign n19197 = \sport0_cfg_SP_ENg_reg/NET0131  & ~n19196 ;
  assign n19198 = ~\sport0_cfg_SCLKi_h_reg/NET0131  & ~n19197 ;
  assign n19199 = \sport0_cfg_SCLKi_h_reg/NET0131  & n19197 ;
  assign n19200 = ~n19198 & ~n19199 ;
  assign n19201 = \core_c_dec_MTASTAT_E_reg/P0001  & n5951 ;
  assign n19202 = ~n18681 & ~n19201 ;
  assign n19203 = ~n5950 & n13803 ;
  assign n19204 = \core_c_dec_ALUop_E_reg/P0001  & n19203 ;
  assign n19205 = n19202 & ~n19204 ;
  assign n19206 = \core_c_dec_ALUop_E_reg/P0001  & n13803 ;
  assign n19207 = ~n14494 & ~n14534 ;
  assign n19208 = ~n14532 & ~n19207 ;
  assign n19210 = n14474 & ~n14490 ;
  assign n19211 = n19208 & ~n19210 ;
  assign n19209 = ~n14491 & ~n19208 ;
  assign n19212 = ~n13809 & ~n19209 ;
  assign n19213 = ~n19211 & n19212 ;
  assign n19214 = \core_c_psq_MSTAT_reg_DO_reg[3]/NET0131  & n19213 ;
  assign n19215 = ~n13809 & ~n19208 ;
  assign n19217 = n14404 & ~n19210 ;
  assign n19216 = ~n14406 & n19210 ;
  assign n19218 = ~n14491 & ~n19216 ;
  assign n19219 = ~n19217 & n19218 ;
  assign n19220 = n19215 & ~n19219 ;
  assign n19221 = ~n19215 & n19219 ;
  assign n19222 = ~n19220 & ~n19221 ;
  assign n19223 = n19214 & n19222 ;
  assign n19224 = ~n19214 & ~n19222 ;
  assign n19225 = ~n19223 & ~n19224 ;
  assign n19226 = n19206 & ~n19225 ;
  assign n19227 = \core_c_dec_MTASTAT_E_reg/P0001  & n9435 ;
  assign n19234 = \core_c_psq_ststk_sts7x23_STcell_reg[6][1]/P0001  & n14711 ;
  assign n19232 = \core_c_psq_ststk_sts7x23_STcell_reg[1][1]/P0001  & n14708 ;
  assign n19233 = \core_c_psq_ststk_sts7x23_STcell_reg[5][1]/P0001  & n14699 ;
  assign n19237 = ~n19232 & ~n19233 ;
  assign n19238 = ~n19234 & n19237 ;
  assign n19228 = \core_c_psq_ststk_sts7x23_STcell_reg[2][1]/P0001  & n14713 ;
  assign n19229 = \core_c_psq_ststk_sts7x23_STcell_reg[0][1]/P0001  & n14702 ;
  assign n19235 = ~n19228 & ~n19229 ;
  assign n19230 = \core_c_psq_ststk_sts7x23_STcell_reg[3][1]/P0001  & n14704 ;
  assign n19231 = \core_c_psq_ststk_sts7x23_STcell_reg[4][1]/P0001  & n14706 ;
  assign n19236 = ~n19230 & ~n19231 ;
  assign n19239 = n19235 & n19236 ;
  assign n19240 = n19238 & n19239 ;
  assign n19241 = n14697 & ~n19240 ;
  assign n19242 = ~n19227 & ~n19241 ;
  assign n19243 = ~n19226 & n19242 ;
  assign n19245 = \core_c_psq_MSTAT_reg_DO_reg[2]/NET0131  & \core_eu_ec_cun_AV_reg/P0001  ;
  assign n19246 = ~n19213 & ~n19245 ;
  assign n19247 = n19206 & ~n19246 ;
  assign n19244 = \core_c_dec_MTASTAT_E_reg/P0001  & n8715 ;
  assign n19254 = \core_c_psq_ststk_sts7x23_STcell_reg[6][2]/P0001  & n14711 ;
  assign n19252 = \core_c_psq_ststk_sts7x23_STcell_reg[1][2]/P0001  & n14708 ;
  assign n19253 = \core_c_psq_ststk_sts7x23_STcell_reg[5][2]/P0001  & n14699 ;
  assign n19257 = ~n19252 & ~n19253 ;
  assign n19258 = ~n19254 & n19257 ;
  assign n19248 = \core_c_psq_ststk_sts7x23_STcell_reg[2][2]/P0001  & n14713 ;
  assign n19249 = \core_c_psq_ststk_sts7x23_STcell_reg[0][2]/P0001  & n14702 ;
  assign n19255 = ~n19248 & ~n19249 ;
  assign n19250 = \core_c_psq_ststk_sts7x23_STcell_reg[3][2]/P0001  & n14704 ;
  assign n19251 = \core_c_psq_ststk_sts7x23_STcell_reg[4][2]/P0001  & n14706 ;
  assign n19256 = ~n19250 & ~n19251 ;
  assign n19259 = n19255 & n19256 ;
  assign n19260 = n19258 & n19259 ;
  assign n19261 = n14697 & ~n19260 ;
  assign n19262 = ~n19244 & ~n19261 ;
  assign n19263 = ~n19247 & n19262 ;
  assign n19264 = ~n19243 & ~n19263 ;
  assign n19265 = n19243 & n19263 ;
  assign n19266 = ~n19264 & ~n19265 ;
  assign n19270 = ~\core_c_dec_IR_reg[0]/NET0131  & ~\core_c_dec_IR_reg[1]/NET0131  ;
  assign n19271 = n6091 & n19270 ;
  assign n19272 = n19266 & n19271 ;
  assign n19267 = \core_c_dec_IR_reg[0]/NET0131  & ~\core_c_dec_IR_reg[1]/NET0131  ;
  assign n19268 = n6091 & n19267 ;
  assign n19269 = ~n19266 & n19268 ;
  assign n19301 = \core_c_dec_IR_reg[0]/NET0131  & \core_c_dec_IR_reg[1]/NET0131  ;
  assign n19302 = n6091 & n19301 ;
  assign n19303 = n19263 & n19302 ;
  assign n19298 = ~\core_c_dec_IR_reg[0]/NET0131  & \core_c_dec_IR_reg[1]/NET0131  ;
  assign n19299 = n6091 & n19298 ;
  assign n19300 = ~n19263 & n19299 ;
  assign n19273 = n6095 & n19267 ;
  assign n19274 = ~n14491 & n19207 ;
  assign n19275 = ~n14467 & n14532 ;
  assign n19276 = ~n19210 & ~n19275 ;
  assign n19277 = ~n19274 & n19276 ;
  assign n19278 = ~n13809 & ~n19277 ;
  assign n19279 = n19206 & n19278 ;
  assign n19286 = \core_c_psq_ststk_sts7x23_STcell_reg[2][3]/P0001  & n14713 ;
  assign n19284 = \core_c_psq_ststk_sts7x23_STcell_reg[1][3]/P0001  & n14708 ;
  assign n19285 = \core_c_psq_ststk_sts7x23_STcell_reg[6][3]/P0001  & n14711 ;
  assign n19289 = ~n19284 & ~n19285 ;
  assign n19290 = ~n19286 & n19289 ;
  assign n19280 = \core_c_psq_ststk_sts7x23_STcell_reg[5][3]/P0001  & n14699 ;
  assign n19281 = \core_c_psq_ststk_sts7x23_STcell_reg[0][3]/P0001  & n14702 ;
  assign n19287 = ~n19280 & ~n19281 ;
  assign n19282 = \core_c_psq_ststk_sts7x23_STcell_reg[3][3]/P0001  & n14704 ;
  assign n19283 = \core_c_psq_ststk_sts7x23_STcell_reg[4][3]/P0001  & n14706 ;
  assign n19288 = ~n19282 & ~n19283 ;
  assign n19291 = n19287 & n19288 ;
  assign n19292 = n19290 & n19291 ;
  assign n19293 = n14697 & ~n19292 ;
  assign n19294 = \core_c_dec_MTASTAT_E_reg/P0001  & n8113 ;
  assign n19295 = ~n19293 & ~n19294 ;
  assign n19296 = ~n19279 & n19295 ;
  assign n19297 = n19273 & n19296 ;
  assign n19304 = n6095 & n19270 ;
  assign n19305 = ~n19296 & n19304 ;
  assign n19306 = ~n19297 & ~n19305 ;
  assign n19307 = ~n19300 & n19306 ;
  assign n19308 = ~n19303 & n19307 ;
  assign n19309 = ~n19269 & n19308 ;
  assign n19310 = ~n19272 & n19309 ;
  assign n19311 = ~n19205 & ~n19310 ;
  assign n19312 = \core_eu_ea_alu_ea_dec_AMF_E_reg[4]/NET0131  & n19206 ;
  assign n19313 = ~n5950 & n13811 ;
  assign n19314 = n19312 & n19313 ;
  assign n19315 = n19202 & ~n19314 ;
  assign n19316 = ~\core_eu_ec_cun_AS_reg/P0001  & ~n19301 ;
  assign n19317 = \core_eu_ec_cun_AS_reg/P0001  & ~n19298 ;
  assign n19318 = ~n19316 & ~n19317 ;
  assign n19319 = n19315 & n19318 ;
  assign n19328 = \core_c_psq_ststk_sts7x23_STcell_reg[1][4]/P0001  & n14708 ;
  assign n19326 = \core_c_psq_ststk_sts7x23_STcell_reg[2][4]/P0001  & n14713 ;
  assign n19327 = \core_c_psq_ststk_sts7x23_STcell_reg[3][4]/P0001  & n14704 ;
  assign n19331 = ~n19326 & ~n19327 ;
  assign n19332 = ~n19328 & n19331 ;
  assign n19322 = \core_c_psq_ststk_sts7x23_STcell_reg[5][4]/P0001  & n14699 ;
  assign n19323 = \core_c_psq_ststk_sts7x23_STcell_reg[0][4]/P0001  & n14702 ;
  assign n19329 = ~n19322 & ~n19323 ;
  assign n19324 = \core_c_psq_ststk_sts7x23_STcell_reg[6][4]/P0001  & n14711 ;
  assign n19325 = \core_c_psq_ststk_sts7x23_STcell_reg[4][4]/P0001  & n14706 ;
  assign n19330 = ~n19324 & ~n19325 ;
  assign n19333 = n19329 & n19330 ;
  assign n19334 = n19332 & n19333 ;
  assign n19335 = n14697 & ~n19334 ;
  assign n19320 = n13838 & n19312 ;
  assign n19321 = \core_c_dec_MTASTAT_E_reg/P0001  & n10069 ;
  assign n19336 = ~n19320 & ~n19321 ;
  assign n19337 = ~n19335 & n19336 ;
  assign n19339 = ~n19301 & n19337 ;
  assign n19338 = ~n19298 & ~n19337 ;
  assign n19340 = ~n19315 & ~n19338 ;
  assign n19341 = ~n19339 & n19340 ;
  assign n19342 = ~n19319 & ~n19341 ;
  assign n19343 = n6095 & ~n19342 ;
  assign n19344 = \core_eu_ec_cun_AC_reg/P0001  & n19304 ;
  assign n19345 = ~\core_eu_ec_cun_AV_reg/P0001  & n19302 ;
  assign n19350 = ~n19344 & ~n19345 ;
  assign n19346 = \core_eu_ec_cun_AV_reg/P0001  & n19299 ;
  assign n19347 = ~n4137 & n19268 ;
  assign n19351 = ~n19346 & ~n19347 ;
  assign n19348 = n4137 & n19271 ;
  assign n19349 = ~\core_eu_ec_cun_AC_reg/P0001  & n19273 ;
  assign n19352 = ~n19348 & ~n19349 ;
  assign n19353 = n19351 & n19352 ;
  assign n19354 = n19350 & n19353 ;
  assign n19355 = n19205 & ~n19354 ;
  assign n19356 = n6097 & n19301 ;
  assign n19357 = ~n4117 & ~n19356 ;
  assign n19358 = ~n19355 & n19357 ;
  assign n19359 = ~n19343 & n19358 ;
  assign n19360 = ~n19311 & n19359 ;
  assign n19361 = ~\core_eu_ec_cun_condOK_CE_reg/P0001  & n4117 ;
  assign n19362 = n4149 & ~n19361 ;
  assign n19363 = ~n19360 & n19362 ;
  assign n19364 = n15314 & ~n17777 ;
  assign n19365 = ~n17778 & ~n19364 ;
  assign n19366 = n15244 & n19365 ;
  assign n19367 = ~n15244 & ~n19365 ;
  assign n19368 = ~n19366 & ~n19367 ;
  assign n19369 = \core_c_psq_MSTAT_reg_DO_reg[4]/NET0131  & ~n19368 ;
  assign n19370 = ~n17767 & ~n17774 ;
  assign n19371 = ~n17698 & ~n17745 ;
  assign n19372 = n17772 & ~n19371 ;
  assign n19373 = ~n17759 & ~n19372 ;
  assign n19374 = ~n17768 & ~n19373 ;
  assign n19375 = n19370 & ~n19374 ;
  assign n19376 = ~n19370 & n19374 ;
  assign n19377 = ~n19375 & ~n19376 ;
  assign n19378 = ~\core_c_psq_MSTAT_reg_DO_reg[4]/NET0131  & n19377 ;
  assign n19379 = ~n19369 & ~n19378 ;
  assign n19380 = n18262 & ~n19379 ;
  assign n19381 = n14664 & ~n17805 ;
  assign n19382 = \core_eu_em_mac_em_reg_mr1swe_DO_reg[15]/P0001  & ~n19381 ;
  assign n19383 = \core_c_psq_MSTAT_reg_DO_reg[0]/P0002  & ~n17806 ;
  assign n19384 = \core_eu_em_mac_em_reg_mr2swe_DO_reg[7]/P0001  & n18268 ;
  assign n19385 = n14665 & n17822 ;
  assign n19386 = ~n19384 & ~n19385 ;
  assign n19387 = n19383 & ~n19386 ;
  assign n19388 = ~n19382 & ~n19387 ;
  assign n19389 = ~n18262 & ~n19388 ;
  assign n19390 = \core_eu_em_mac_em_reg_mr1swe_DO_reg[15]/P0001  & ~n19383 ;
  assign n19391 = ~n19389 & ~n19390 ;
  assign n19392 = ~n19380 & n19391 ;
  assign n19393 = n14752 & ~n19379 ;
  assign n19394 = \core_eu_em_mac_em_reg_mr1rwe_DO_reg[15]/P0001  & ~n17809 ;
  assign n19395 = ~\core_c_psq_MSTAT_reg_DO_reg[0]/P0002  & ~n17806 ;
  assign n19396 = ~n17823 & ~n17828 ;
  assign n19397 = n19395 & ~n19396 ;
  assign n19398 = ~n19394 & ~n19397 ;
  assign n19399 = ~n14752 & ~n19398 ;
  assign n19400 = \core_eu_em_mac_em_reg_mr1rwe_DO_reg[15]/P0001  & ~n19395 ;
  assign n19401 = ~n19399 & ~n19400 ;
  assign n19402 = ~n19393 & n19401 ;
  assign n19403 = \core_c_psq_MSTAT_reg_DO_reg[4]/NET0131  & ~n17794 ;
  assign n19404 = ~n15317 & ~n17781 ;
  assign n19405 = n17779 & n19404 ;
  assign n19406 = ~n17779 & ~n19404 ;
  assign n19407 = ~n19405 & ~n19406 ;
  assign n19408 = ~\core_c_psq_MSTAT_reg_DO_reg[4]/NET0131  & n19407 ;
  assign n19409 = ~n19403 & ~n19408 ;
  assign n19410 = ~\sport0_cfg_SCLKi_cnt_reg[0]/NET0131  & ~\sport0_cfg_SCLKi_cnt_reg[1]/NET0131  ;
  assign n19411 = \sport0_cfg_SCLKi_cnt_reg[0]/NET0131  & \sport0_cfg_SCLKi_cnt_reg[1]/NET0131  ;
  assign n19412 = ~n19410 & ~n19411 ;
  assign n19413 = n19197 & n19412 ;
  assign n19414 = n17698 & ~n17743 ;
  assign n19415 = ~n17698 & n17743 ;
  assign n19416 = ~n19414 & ~n19415 ;
  assign n19417 = n17737 & n19416 ;
  assign n19418 = ~n17737 & ~n19416 ;
  assign n19419 = ~n19417 & ~n19418 ;
  assign n19420 = \core_c_psq_MSTAT_reg_DO_reg[4]/NET0131  & ~n19419 ;
  assign n19421 = ~n16363 & n17662 ;
  assign n19422 = n17674 & ~n19421 ;
  assign n19423 = n17567 & ~n19422 ;
  assign n19424 = n17685 & ~n19423 ;
  assign n19425 = n16980 & ~n19424 ;
  assign n19426 = n17690 & ~n19425 ;
  assign n19427 = ~n17692 & n19426 ;
  assign n19428 = ~n17092 & ~n19427 ;
  assign n19429 = n17079 & ~n19428 ;
  assign n19430 = ~n17079 & n19428 ;
  assign n19431 = ~n19429 & ~n19430 ;
  assign n19432 = n17095 & n19431 ;
  assign n19433 = ~n17095 & ~n19431 ;
  assign n19434 = ~n19432 & ~n19433 ;
  assign n19435 = ~\core_c_psq_MSTAT_reg_DO_reg[4]/NET0131  & n19434 ;
  assign n19436 = ~n19420 & ~n19435 ;
  assign n19437 = ~\sport1_cfg_SCLKi_cnt_reg[0]/NET0131  & ~\sport1_cfg_SCLKi_cnt_reg[1]/NET0131  ;
  assign n19438 = \sport1_cfg_SCLKi_cnt_reg[0]/NET0131  & \sport1_cfg_SCLKi_cnt_reg[1]/NET0131  ;
  assign n19439 = ~n19437 & ~n19438 ;
  assign n19440 = n19130 & n19439 ;
  assign n19468 = \clkc_OUTcnt_reg[0]/NET0131  & \clkc_OUTcnt_reg[1]/NET0131  ;
  assign n19469 = \clkc_OUTcnt_reg[2]/NET0131  & n19468 ;
  assign n19470 = \clkc_OUTcnt_reg[3]/NET0131  & n19469 ;
  assign n19471 = \clkc_OUTcnt_reg[4]/NET0131  & n19470 ;
  assign n19472 = \clkc_OUTcnt_reg[5]/NET0131  & n19471 ;
  assign n19474 = \clkc_OUTcnt_reg[6]/NET0131  & n19472 ;
  assign n19441 = \clkc_OUTcnt_reg[0]/NET0131  & ~\clkc_ckr_reg_DO_reg[8]/NET0131  ;
  assign n19442 = ~\clkc_OUTcnt_reg[6]/NET0131  & \clkc_ckr_reg_DO_reg[14]/NET0131  ;
  assign n19443 = ~\clkc_OUTcnt_reg[2]/NET0131  & \clkc_ckr_reg_DO_reg[10]/NET0131  ;
  assign n19455 = ~n19442 & ~n19443 ;
  assign n19444 = ~\clkc_OUTcnt_reg[3]/NET0131  & \clkc_ckr_reg_DO_reg[11]/NET0131  ;
  assign n19445 = ~\clkc_OUTcnt_reg[0]/NET0131  & \clkc_ckr_reg_DO_reg[8]/NET0131  ;
  assign n19456 = ~n19444 & ~n19445 ;
  assign n19446 = \clkc_OUTcnt_reg[3]/NET0131  & ~\clkc_ckr_reg_DO_reg[11]/NET0131  ;
  assign n19447 = \clkc_OUTcnt_reg[2]/NET0131  & ~\clkc_ckr_reg_DO_reg[10]/NET0131  ;
  assign n19457 = ~n19446 & ~n19447 ;
  assign n19463 = n19456 & n19457 ;
  assign n19464 = n19455 & n19463 ;
  assign n19454 = \clkc_OUTcnt_reg[6]/NET0131  & ~\clkc_ckr_reg_DO_reg[14]/NET0131  ;
  assign n19452 = ~\clkc_OUTcnt_reg[5]/NET0131  & \clkc_ckr_reg_DO_reg[13]/NET0131  ;
  assign n19453 = \clkc_OUTcnt_reg[4]/NET0131  & ~\clkc_ckr_reg_DO_reg[12]/NET0131  ;
  assign n19460 = ~n19452 & ~n19453 ;
  assign n19461 = ~n19454 & n19460 ;
  assign n19448 = ~\clkc_OUTcnt_reg[4]/NET0131  & \clkc_ckr_reg_DO_reg[12]/NET0131  ;
  assign n19449 = \clkc_OUTcnt_reg[1]/NET0131  & ~\clkc_ckr_reg_DO_reg[9]/NET0131  ;
  assign n19458 = ~n19448 & ~n19449 ;
  assign n19450 = \clkc_OUTcnt_reg[5]/NET0131  & ~\clkc_ckr_reg_DO_reg[13]/NET0131  ;
  assign n19451 = ~\clkc_OUTcnt_reg[1]/NET0131  & \clkc_ckr_reg_DO_reg[9]/NET0131  ;
  assign n19459 = ~n19450 & ~n19451 ;
  assign n19462 = n19458 & n19459 ;
  assign n19465 = n19461 & n19462 ;
  assign n19466 = n19464 & n19465 ;
  assign n19467 = ~n19441 & n19466 ;
  assign n19473 = ~\clkc_OUTcnt_reg[6]/NET0131  & ~n19472 ;
  assign n19475 = ~n19467 & ~n19473 ;
  assign n19476 = ~n19474 & n19475 ;
  assign n19477 = \core_c_psq_INT_en_reg/NET0131  & ~n4094 ;
  assign n19478 = \core_c_psq_Iact_E_reg[4]/NET0131  & ~n19477 ;
  assign n19481 = \core_c_psq_IMASK_reg[9]/NET0131  & \core_c_psq_Iflag_reg[8]/NET0131  ;
  assign n19482 = ~\core_c_psq_Iflag_reg[10]/NET0131  & ~n19481 ;
  assign n19483 = ~\core_c_psq_PCS_reg[3]/NET0131  & ~n19482 ;
  assign n19484 = n19477 & ~n19483 ;
  assign n19485 = \core_c_psq_IMASK_reg[8]/NET0131  & \core_c_psq_Iflag_reg[9]/NET0131  ;
  assign n19486 = ~\core_c_psq_PCS_reg[3]/NET0131  & n19485 ;
  assign n19487 = n19484 & ~n19486 ;
  assign n19479 = \core_c_psq_IMASK_reg[4]/NET0131  & \core_c_psq_Iflag_reg[5]/NET0131  ;
  assign n19480 = ~\core_c_psq_PCS_reg[3]/NET0131  & n19479 ;
  assign n19488 = \core_c_psq_IMASK_reg[7]/NET0131  & \core_c_psq_Iflag_reg[6]/NET0131  ;
  assign n19489 = ~\core_c_psq_PCS_reg[3]/NET0131  & n19488 ;
  assign n19490 = \core_c_psq_IMASK_reg[5]/NET0131  & \core_c_psq_Iflag_reg[4]/NET0131  ;
  assign n19491 = ~\core_c_psq_PCS_reg[3]/NET0131  & n19490 ;
  assign n19492 = \core_c_psq_IMASK_reg[6]/NET0131  & \core_c_psq_Iflag_reg[7]/NET0131  ;
  assign n19493 = ~\core_c_psq_PCS_reg[3]/NET0131  & n19492 ;
  assign n19494 = ~n19491 & ~n19493 ;
  assign n19495 = ~n19489 & n19494 ;
  assign n19496 = n19480 & n19495 ;
  assign n19497 = n19487 & n19496 ;
  assign n19498 = ~n19478 & ~n19497 ;
  assign n19499 = \core_c_dec_MTMR1_E_reg/P0001  & n14665 ;
  assign n19502 = ~\core_c_dec_accPM_E_reg/P0001  & ~n10289 ;
  assign n19503 = \core_c_dec_accPM_E_reg/P0001  & ~n13075 ;
  assign n19504 = ~n19502 & ~n19503 ;
  assign n19505 = n19499 & ~n19504 ;
  assign n19500 = ~\core_eu_em_mac_em_reg_mr1swe_DO_reg[9]/P0001  & ~n19499 ;
  assign n19501 = ~n18268 & n19383 ;
  assign n19506 = ~n19500 & n19501 ;
  assign n19507 = ~n19505 & n19506 ;
  assign n19508 = n18269 & n19383 ;
  assign n19509 = \core_eu_em_mac_em_reg_mr1swe_DO_reg[9]/P0001  & ~n19383 ;
  assign n19510 = ~n19508 & ~n19509 ;
  assign n19511 = ~n19507 & n19510 ;
  assign n19512 = ~n18262 & ~n19511 ;
  assign n19513 = ~n17092 & ~n17692 ;
  assign n19514 = n19426 & n19513 ;
  assign n19515 = ~n19426 & ~n19513 ;
  assign n19516 = ~n19514 & ~n19515 ;
  assign n19517 = \core_c_psq_MSTAT_reg_DO_reg[4]/NET0131  & ~n19516 ;
  assign n19518 = ~n16856 & ~n17687 ;
  assign n19519 = ~n16979 & ~n19424 ;
  assign n19520 = ~n17688 & ~n19519 ;
  assign n19521 = n19518 & ~n19520 ;
  assign n19522 = ~n19518 & n19520 ;
  assign n19523 = ~n19521 & ~n19522 ;
  assign n19524 = ~\core_c_psq_MSTAT_reg_DO_reg[4]/NET0131  & n19523 ;
  assign n19525 = ~n19517 & ~n19524 ;
  assign n19526 = n18262 & ~n19525 ;
  assign n19527 = ~n19512 & ~n19526 ;
  assign n19529 = \core_c_dec_IR_reg[16]/NET0131  & n6028 ;
  assign n19530 = ~n6119 & ~n19529 ;
  assign n19531 = ~n4117 & n19530 ;
  assign n19528 = ~\core_c_dec_SHTop_E_reg/P0001  & n4117 ;
  assign n19532 = n4116 & ~n19528 ;
  assign n19533 = ~n19531 & n19532 ;
  assign n19534 = \sport0_cfg_SCLKi_cnt_reg[2]/NET0131  & n19411 ;
  assign n19535 = \sport0_cfg_SCLKi_cnt_reg[3]/NET0131  & n19534 ;
  assign n19536 = \sport0_cfg_SCLKi_cnt_reg[4]/NET0131  & n19535 ;
  assign n19537 = ~\sport0_cfg_SCLKi_cnt_reg[5]/NET0131  & ~n19536 ;
  assign n19538 = \sport0_cfg_SCLKi_cnt_reg[5]/NET0131  & n19536 ;
  assign n19539 = ~n19537 & ~n19538 ;
  assign n19540 = n19197 & n19539 ;
  assign n19541 = ~\sport0_cfg_SCLKi_cnt_reg[2]/NET0131  & ~n19411 ;
  assign n19542 = ~n19534 & ~n19541 ;
  assign n19543 = n19197 & n19542 ;
  assign n19544 = \sport0_cfg_SCLKi_cnt_reg[6]/NET0131  & n19538 ;
  assign n19545 = \sport0_cfg_SCLKi_cnt_reg[7]/NET0131  & n19544 ;
  assign n19546 = \sport0_cfg_SCLKi_cnt_reg[8]/NET0131  & n19545 ;
  assign n19547 = \sport0_cfg_SCLKi_cnt_reg[9]/NET0131  & n19546 ;
  assign n19548 = \sport0_cfg_SCLKi_cnt_reg[10]/NET0131  & n19547 ;
  assign n19549 = \sport0_cfg_SCLKi_cnt_reg[11]/NET0131  & n19548 ;
  assign n19550 = \sport0_cfg_SCLKi_cnt_reg[12]/NET0131  & n19549 ;
  assign n19552 = \sport0_cfg_SCLKi_cnt_reg[13]/NET0131  & n19550 ;
  assign n19551 = ~\sport0_cfg_SCLKi_cnt_reg[13]/NET0131  & ~n19550 ;
  assign n19553 = n19197 & ~n19551 ;
  assign n19554 = ~n19552 & n19553 ;
  assign n19555 = ~\sport0_cfg_SCLKi_cnt_reg[0]/NET0131  & n19197 ;
  assign n19557 = ~\core_c_dec_accPM_E_reg/P0001  & ~n7607 ;
  assign n19558 = \core_c_dec_accPM_E_reg/P0001  & ~n12520 ;
  assign n19559 = ~n19557 & ~n19558 ;
  assign n19560 = n19499 & ~n19559 ;
  assign n19556 = ~\core_eu_em_mac_em_reg_mr1swe_DO_reg[0]/P0001  & ~n19499 ;
  assign n19561 = n19501 & ~n19556 ;
  assign n19562 = ~n19560 & n19561 ;
  assign n19563 = \core_eu_em_mac_em_reg_mr1swe_DO_reg[0]/P0001  & ~n19383 ;
  assign n19564 = ~n19508 & ~n19563 ;
  assign n19565 = ~n19562 & n19564 ;
  assign n19566 = ~n18262 & ~n19565 ;
  assign n19567 = ~n17660 & ~n17668 ;
  assign n19568 = n16363 & n19567 ;
  assign n19569 = ~n16363 & ~n19567 ;
  assign n19570 = ~n19568 & ~n19569 ;
  assign n19594 = \core_c_psq_MSTAT_reg_DO_reg[4]/NET0131  & ~n19570 ;
  assign n19586 = ~n15898 & ~n16360 ;
  assign n19580 = n16059 & ~n16350 ;
  assign n19581 = n16358 & ~n19580 ;
  assign n19587 = ~n15775 & ~n19581 ;
  assign n19588 = ~n16353 & ~n19587 ;
  assign n19589 = n19586 & ~n19588 ;
  assign n19590 = ~n19586 & n19588 ;
  assign n19591 = ~n19589 & ~n19590 ;
  assign n19595 = ~\core_c_psq_MSTAT_reg_DO_reg[4]/NET0131  & n19591 ;
  assign n19596 = ~n19594 & ~n19595 ;
  assign n19579 = ~n15775 & ~n16353 ;
  assign n19582 = ~n19579 & n19581 ;
  assign n19583 = n19579 & ~n19581 ;
  assign n19584 = ~n19582 & ~n19583 ;
  assign n19585 = ~\core_c_psq_MSTAT_reg_DO_reg[4]/NET0131  & n19584 ;
  assign n19592 = \core_c_psq_MSTAT_reg_DO_reg[4]/NET0131  & n19591 ;
  assign n19593 = ~n19585 & ~n19592 ;
  assign n19602 = ~n15978 & ~n16355 ;
  assign n19603 = ~n16058 & ~n16350 ;
  assign n19604 = ~n16356 & ~n19603 ;
  assign n19605 = n19602 & ~n19604 ;
  assign n19606 = ~n19602 & n19604 ;
  assign n19607 = ~n19605 & ~n19606 ;
  assign n19634 = ~\core_c_psq_MSTAT_reg_DO_reg[4]/NET0131  & n19607 ;
  assign n19635 = \core_c_psq_MSTAT_reg_DO_reg[4]/NET0131  & n19584 ;
  assign n19636 = ~n19634 & ~n19635 ;
  assign n19597 = ~n16058 & ~n16356 ;
  assign n19598 = n16350 & ~n19597 ;
  assign n19599 = ~n16350 & n19597 ;
  assign n19600 = ~n19598 & ~n19599 ;
  assign n19601 = ~\core_c_psq_MSTAT_reg_DO_reg[4]/NET0131  & ~n19600 ;
  assign n19608 = \core_c_psq_MSTAT_reg_DO_reg[4]/NET0131  & ~n19607 ;
  assign n19609 = ~n19601 & ~n19608 ;
  assign n19610 = n16327 & ~n16343 ;
  assign n19611 = ~n16347 & ~n19610 ;
  assign n19612 = ~n16339 & ~n16346 ;
  assign n19613 = ~n19611 & n19612 ;
  assign n19614 = n19611 & ~n19612 ;
  assign n19615 = ~n19613 & ~n19614 ;
  assign n19637 = \core_c_psq_MSTAT_reg_DO_reg[4]/NET0131  & ~n19615 ;
  assign n19638 = ~n16343 & ~n16347 ;
  assign n19639 = ~n16327 & n19638 ;
  assign n19640 = n16327 & ~n19638 ;
  assign n19641 = ~n19639 & ~n19640 ;
  assign n19642 = ~\core_c_psq_MSTAT_reg_DO_reg[4]/NET0131  & n19641 ;
  assign n19643 = ~n19637 & ~n19642 ;
  assign n19616 = ~\core_c_psq_MSTAT_reg_DO_reg[4]/NET0131  & n19615 ;
  assign n19617 = \core_c_psq_MSTAT_reg_DO_reg[4]/NET0131  & n19600 ;
  assign n19618 = ~n19616 & ~n19617 ;
  assign n19644 = \core_c_psq_MSTAT_reg_DO_reg[4]/NET0131  & ~n19641 ;
  assign n19629 = n16312 & ~n16326 ;
  assign n19630 = ~n16327 & ~n19629 ;
  assign n19645 = ~\core_c_psq_MSTAT_reg_DO_reg[4]/NET0131  & n19630 ;
  assign n19646 = ~n19644 & ~n19645 ;
  assign n19631 = \core_c_psq_MSTAT_reg_DO_reg[4]/NET0131  & ~n19630 ;
  assign n19620 = ~n16159 & n16310 ;
  assign n19621 = ~n16311 & ~n19620 ;
  assign n19632 = ~\core_c_psq_MSTAT_reg_DO_reg[4]/NET0131  & ~n19621 ;
  assign n19633 = ~n19631 & ~n19632 ;
  assign n19619 = ~\core_c_psq_MSTAT_reg_DO_reg[4]/NET0131  & n18289 ;
  assign n19622 = \core_c_psq_MSTAT_reg_DO_reg[4]/NET0131  & n19621 ;
  assign n19623 = ~n19619 & ~n19622 ;
  assign n19624 = ~n16276 & n16304 ;
  assign n19625 = ~n16305 & ~n19624 ;
  assign n19626 = ~\core_c_psq_MSTAT_reg_DO_reg[4]/NET0131  & n19625 ;
  assign n19627 = \core_c_psq_MSTAT_reg_DO_reg[4]/NET0131  & n18284 ;
  assign n19628 = ~n19626 & ~n19627 ;
  assign n19654 = ~n16301 & ~n16303 ;
  assign n19655 = ~n16297 & n19654 ;
  assign n19656 = n16297 & ~n19654 ;
  assign n19657 = ~n19655 & ~n19656 ;
  assign n19668 = ~\core_c_psq_MSTAT_reg_DO_reg[4]/NET0131  & ~n19657 ;
  assign n19669 = \core_c_psq_MSTAT_reg_DO_reg[4]/NET0131  & n19625 ;
  assign n19670 = ~n19668 & ~n19669 ;
  assign n19658 = \core_c_psq_MSTAT_reg_DO_reg[4]/NET0131  & ~n19657 ;
  assign n19659 = ~n16291 & ~n16296 ;
  assign n19660 = ~n16297 & ~n19659 ;
  assign n19661 = ~\core_c_psq_MSTAT_reg_DO_reg[4]/NET0131  & n19660 ;
  assign n19662 = ~n19658 & ~n19661 ;
  assign n19663 = ~n16280 & n16290 ;
  assign n19664 = ~n16291 & ~n19663 ;
  assign n19671 = ~\core_c_psq_MSTAT_reg_DO_reg[4]/NET0131  & n19664 ;
  assign n19672 = \core_c_psq_MSTAT_reg_DO_reg[4]/NET0131  & n19660 ;
  assign n19673 = ~n19671 & ~n19672 ;
  assign n19665 = \core_c_psq_MSTAT_reg_DO_reg[4]/NET0131  & ~n19664 ;
  assign n19647 = \core_eu_em_mac_em_reg_mxopwe_DO_reg[0]/P0001  & \core_eu_em_mac_em_reg_myopwe_DO_reg[0]/P0001  ;
  assign n19648 = ~n16286 & n19647 ;
  assign n19649 = n16286 & ~n19647 ;
  assign n19650 = ~n19648 & ~n19649 ;
  assign n19666 = ~\core_c_psq_MSTAT_reg_DO_reg[4]/NET0131  & n19650 ;
  assign n19667 = ~n19665 & ~n19666 ;
  assign n19651 = \core_c_psq_MSTAT_reg_DO_reg[4]/NET0131  & ~n19650 ;
  assign n19652 = ~n7469 & n17341 ;
  assign n19653 = ~n19651 & ~n19652 ;
  assign n19674 = \core_eu_em_mac_em_dec_emcorepi_DO_reg[0]/P0001  & ~\memc_usysr_DO_reg[10]/NET0131  ;
  assign n19675 = n19653 & n19674 ;
  assign n19676 = ~n19667 & n19675 ;
  assign n19677 = n19673 & n19676 ;
  assign n19678 = n19662 & n19677 ;
  assign n19679 = n19670 & n19678 ;
  assign n19680 = n19628 & n19679 ;
  assign n19681 = ~n18291 & n19680 ;
  assign n19682 = n19623 & n19681 ;
  assign n19683 = ~n19633 & n19682 ;
  assign n19684 = n19646 & n19683 ;
  assign n19685 = n19618 & n19684 ;
  assign n19686 = ~n19643 & n19685 ;
  assign n19687 = ~n19609 & n19686 ;
  assign n19688 = n19636 & n19687 ;
  assign n19689 = n19593 & n19688 ;
  assign n19690 = n19596 & n19689 ;
  assign n19571 = ~\core_c_psq_MSTAT_reg_DO_reg[4]/NET0131  & n19570 ;
  assign n19572 = ~n17654 & ~n17667 ;
  assign n19573 = ~n16363 & ~n17660 ;
  assign n19574 = ~n17668 & ~n19573 ;
  assign n19575 = n19572 & ~n19574 ;
  assign n19576 = ~n19572 & n19574 ;
  assign n19577 = ~n19575 & ~n19576 ;
  assign n19578 = \core_c_psq_MSTAT_reg_DO_reg[4]/NET0131  & ~n19577 ;
  assign n19691 = ~n19571 & ~n19578 ;
  assign n19692 = ~n19690 & n19691 ;
  assign n19693 = n18262 & n19692 ;
  assign n19694 = ~n19566 & ~n19693 ;
  assign n19695 = \core_c_dec_Post2_E_reg/P0001  & n4117 ;
  assign n19701 = ~n13574 & ~n13577 ;
  assign n19702 = ~n6023 & n19701 ;
  assign n19696 = ~\core_c_dec_IR_reg[16]/NET0131  & \core_c_dec_IR_reg[17]/NET0131  ;
  assign n19697 = ~\core_c_dec_IR_reg[18]/NET0131  & \core_c_dec_IR_reg[19]/NET0131  ;
  assign n19698 = n6027 & n19697 ;
  assign n19699 = n19696 & n19698 ;
  assign n19700 = \core_c_dec_IR_reg[4]/NET0131  & n19699 ;
  assign n19703 = n6121 & ~n19700 ;
  assign n19704 = n19702 & n19703 ;
  assign n19705 = ~n4117 & ~n19704 ;
  assign n19706 = ~n19695 & ~n19705 ;
  assign n19707 = n4116 & ~n19706 ;
  assign n19708 = \core_c_dec_MTSR1_E_reg/P0001  & ~n17820 ;
  assign n19744 = n18120 & n18745 ;
  assign n19733 = n17920 & n18066 ;
  assign n19734 = ~n17914 & n17975 ;
  assign n19735 = ~n19733 & ~n19734 ;
  assign n19745 = ~n18102 & ~n19735 ;
  assign n19748 = ~n19744 & ~n19745 ;
  assign n19746 = ~n18159 & n18187 ;
  assign n19747 = ~n18180 & n18758 ;
  assign n19749 = ~n19746 & ~n19747 ;
  assign n19750 = n19748 & n19749 ;
  assign n19751 = n17931 & ~n19750 ;
  assign n19725 = ~n18147 & ~n18153 ;
  assign n19726 = ~n18176 & n19725 ;
  assign n19727 = n18084 & n19726 ;
  assign n19728 = n17945 & ~n19727 ;
  assign n19730 = n18059 & n18195 ;
  assign n19731 = n18142 & n19730 ;
  assign n19764 = ~n19728 & n19731 ;
  assign n19765 = ~n19751 & n19764 ;
  assign n19716 = n18076 & n18145 ;
  assign n19719 = ~n18159 & n18184 ;
  assign n19720 = ~n17929 & n18088 ;
  assign n19721 = n17929 & n18765 ;
  assign n19722 = ~n19720 & ~n19721 ;
  assign n19723 = ~n17922 & ~n19722 ;
  assign n19755 = ~n19719 & ~n19723 ;
  assign n19724 = ~n18121 & n18163 ;
  assign n19729 = n17965 & ~n18091 ;
  assign n19756 = ~n19724 & ~n19729 ;
  assign n19759 = n19755 & n19756 ;
  assign n19717 = n17931 & ~n18108 ;
  assign n19718 = ~n17933 & n19717 ;
  assign n19709 = n18119 & n18166 ;
  assign n19742 = n17930 & n18106 ;
  assign n19743 = \core_c_dec_IRE_reg[11]/NET0131  & ~n12000 ;
  assign n19752 = ~n19742 & ~n19743 ;
  assign n19753 = ~n18065 & n19752 ;
  assign n19754 = ~n19709 & n19753 ;
  assign n19760 = ~n19718 & n19754 ;
  assign n19761 = n19759 & n19760 ;
  assign n19738 = n18171 & ~n18180 ;
  assign n19739 = n17925 & n18107 ;
  assign n19740 = ~n19738 & ~n19739 ;
  assign n19741 = ~n17931 & ~n19740 ;
  assign n19737 = ~n18096 & ~n18129 ;
  assign n19732 = ~n18117 & ~n18133 ;
  assign n19736 = n18100 & ~n19735 ;
  assign n19757 = ~n19732 & ~n19736 ;
  assign n19758 = ~n19737 & n19757 ;
  assign n19762 = ~n19741 & n19758 ;
  assign n19763 = n19761 & n19762 ;
  assign n19766 = n19716 & n19763 ;
  assign n19767 = n19765 & n19766 ;
  assign n19713 = n18790 & n18797 ;
  assign n19710 = ~n17931 & n18001 ;
  assign n19711 = ~n18148 & ~n19710 ;
  assign n19712 = n17945 & ~n19711 ;
  assign n19714 = n18050 & ~n19712 ;
  assign n19715 = n19713 & n19714 ;
  assign n19768 = n18007 & n19715 ;
  assign n19769 = n19767 & n19768 ;
  assign n19770 = ~\core_c_dec_MTSR1_E_reg/P0001  & n19769 ;
  assign n19771 = ~n19708 & ~n19770 ;
  assign n19772 = n18717 & ~n19771 ;
  assign n19773 = ~\core_eu_es_sht_es_reg_sr1swe_DO_reg[15]/P0001  & ~n18717 ;
  assign n19774 = ~n19772 & ~n19773 ;
  assign n19775 = n14752 & n19525 ;
  assign n19776 = n17802 & n18325 ;
  assign n19777 = n19504 & n19776 ;
  assign n19778 = \core_eu_em_mac_em_reg_mr1rwe_DO_reg[9]/P0001  & ~n17809 ;
  assign n19779 = n18332 & n19395 ;
  assign n19780 = ~n14752 & ~n19779 ;
  assign n19781 = ~n19778 & n19780 ;
  assign n19782 = ~n19777 & n19781 ;
  assign n19783 = ~n19775 & ~n19782 ;
  assign n19784 = \core_c_dec_MTSR0_E_reg/P0001  & ~n17836 ;
  assign n19787 = n17976 & n18077 ;
  assign n19788 = ~n18037 & ~n19787 ;
  assign n19789 = ~n18032 & ~n18085 ;
  assign n19790 = n19788 & n19789 ;
  assign n19791 = n18902 & n19790 ;
  assign n19792 = n18054 & n19713 ;
  assign n19793 = n18738 & n19792 ;
  assign n19794 = n19791 & n19793 ;
  assign n19804 = ~n18043 & ~n18761 ;
  assign n19805 = n18099 & ~n19804 ;
  assign n19808 = n17931 & ~n18914 ;
  assign n19809 = ~n18175 & n19808 ;
  assign n19833 = ~n19805 & ~n19809 ;
  assign n19815 = n18745 & ~n18775 ;
  assign n19817 = ~n17931 & n18055 ;
  assign n19818 = ~n18139 & ~n19817 ;
  assign n19819 = n18162 & ~n19818 ;
  assign n19834 = ~n19815 & ~n19819 ;
  assign n19835 = n19833 & n19834 ;
  assign n19795 = n18070 & n18124 ;
  assign n19799 = n18056 & ~n18189 ;
  assign n19816 = \core_c_dec_IRE_reg[11]/NET0131  & ~n7164 ;
  assign n19821 = ~n19799 & ~n19816 ;
  assign n19800 = ~n18129 & n18153 ;
  assign n19814 = n17986 & n18103 ;
  assign n19822 = ~n19800 & ~n19814 ;
  assign n19823 = n19821 & n19822 ;
  assign n19824 = ~n19795 & n19823 ;
  assign n19796 = ~n18117 & ~n18912 ;
  assign n19797 = ~n18914 & n19720 ;
  assign n19825 = ~n19796 & ~n19797 ;
  assign n19831 = n19824 & n19825 ;
  assign n19785 = n17931 & ~n18918 ;
  assign n19786 = ~n17933 & n19785 ;
  assign n19801 = ~n17929 & n17952 ;
  assign n19802 = ~n19710 & ~n19801 ;
  assign n19803 = n18171 & ~n19802 ;
  assign n19832 = ~n19786 & ~n19803 ;
  assign n19836 = n19831 & n19832 ;
  assign n19820 = n18136 & ~n18907 ;
  assign n19811 = n17945 & n17959 ;
  assign n19812 = ~n17972 & ~n19811 ;
  assign n19813 = n18147 & n18751 ;
  assign n19828 = n19812 & ~n19813 ;
  assign n19829 = ~n19820 & n19828 ;
  assign n19798 = n17980 & n18187 ;
  assign n19806 = n18046 & n18740 ;
  assign n19826 = ~n19798 & ~n19806 ;
  assign n19807 = n17930 & ~n18918 ;
  assign n19810 = n18183 & n18893 ;
  assign n19827 = ~n19807 & ~n19810 ;
  assign n19830 = n19826 & n19827 ;
  assign n19837 = n19829 & n19830 ;
  assign n19838 = n19836 & n19837 ;
  assign n19839 = n19835 & n19838 ;
  assign n19840 = n19794 & n19839 ;
  assign n19841 = ~\core_c_dec_MTSR0_E_reg/P0001  & n19840 ;
  assign n19842 = ~n19784 & ~n19841 ;
  assign n19843 = n18886 & ~n19842 ;
  assign n19844 = ~\core_eu_es_sht_es_reg_sr0swe_DO_reg[13]/P0001  & ~n18886 ;
  assign n19845 = ~n19843 & ~n19844 ;
  assign n19846 = ~\core_c_dec_accPM_E_reg/P0001  & ~n7859 ;
  assign n19847 = \core_c_dec_accPM_E_reg/P0001  & ~n12556 ;
  assign n19848 = ~n19846 & ~n19847 ;
  assign n19849 = \core_c_dec_MTSR0_E_reg/P0001  & ~n19848 ;
  assign n19850 = ~n17938 & n18080 ;
  assign n19859 = n18754 & ~n18912 ;
  assign n19867 = n18055 & ~n18743 ;
  assign n19866 = n18056 & n18746 ;
  assign n19876 = \core_c_dec_IRE_reg[11]/NET0131  & ~n7801 ;
  assign n19878 = ~n19866 & ~n19876 ;
  assign n19879 = ~n19867 & n19878 ;
  assign n19880 = ~n19859 & n19879 ;
  assign n19886 = ~n19850 & n19880 ;
  assign n19851 = n17925 & ~n17998 ;
  assign n19856 = ~n17931 & n18153 ;
  assign n19857 = ~n18070 & ~n19856 ;
  assign n19858 = n18751 & ~n19857 ;
  assign n19887 = ~n19851 & ~n19858 ;
  assign n19890 = n19886 & n19887 ;
  assign n19877 = n18139 & n18740 ;
  assign n19870 = ~n18749 & ~n18905 ;
  assign n19871 = ~n18914 & ~n19870 ;
  assign n19872 = n18071 & n18099 ;
  assign n19883 = ~n19871 & ~n19872 ;
  assign n19884 = ~n19877 & n19883 ;
  assign n19861 = n18745 & n18893 ;
  assign n19862 = ~n17929 & n18115 ;
  assign n19863 = n17931 & ~n18170 ;
  assign n19864 = ~n19862 & ~n19863 ;
  assign n19865 = ~n18918 & ~n19864 ;
  assign n19881 = ~n19861 & ~n19865 ;
  assign n19868 = ~n18907 & ~n18919 ;
  assign n19869 = n18759 & ~n18912 ;
  assign n19882 = ~n19868 & ~n19869 ;
  assign n19885 = n19881 & n19882 ;
  assign n19891 = n19884 & n19885 ;
  assign n19892 = n19890 & n19891 ;
  assign n19852 = ~n17959 & ~n18030 ;
  assign n19853 = n17945 & ~n19852 ;
  assign n19854 = ~n18143 & ~n19853 ;
  assign n19855 = n18891 & n19854 ;
  assign n19875 = n18765 & ~n18898 ;
  assign n19860 = n18124 & ~n18781 ;
  assign n19873 = ~n17972 & ~n18783 ;
  assign n19874 = n19788 & n19873 ;
  assign n19888 = ~n19860 & n19874 ;
  assign n19889 = ~n19875 & n19888 ;
  assign n19893 = n19855 & n19889 ;
  assign n19894 = n19892 & n19893 ;
  assign n19895 = n19792 & n19894 ;
  assign n19896 = ~\core_c_dec_MTSR0_E_reg/P0001  & n19895 ;
  assign n19897 = ~n19849 & ~n19896 ;
  assign n19898 = n18886 & ~n19897 ;
  assign n19899 = ~\core_eu_es_sht_es_reg_sr0swe_DO_reg[10]/P0001  & ~n18886 ;
  assign n19900 = ~n19898 & ~n19899 ;
  assign n19901 = n19034 & ~n19842 ;
  assign n19902 = ~\core_eu_es_sht_es_reg_sr0rwe_DO_reg[13]/P0001  & ~n19034 ;
  assign n19903 = ~n19901 & ~n19902 ;
  assign n19904 = \core_c_dec_MACop_E_reg/P0001  & n4117 ;
  assign n19905 = ~n18848 & ~n19904 ;
  assign n19906 = n4116 & ~n19905 ;
  assign n19907 = n19034 & ~n19897 ;
  assign n19908 = ~\core_eu_es_sht_es_reg_sr0rwe_DO_reg[10]/P0001  & ~n19034 ;
  assign n19909 = ~n19907 & ~n19908 ;
  assign n19910 = n5730 & n13751 ;
  assign n19911 = \bdma_CMcnt_reg[0]/NET0131  & n19910 ;
  assign n19912 = \bdma_CMcnt_reg[1]/NET0131  & ~n19911 ;
  assign n19913 = n13146 & n13751 ;
  assign n19914 = ~n19912 & ~n19913 ;
  assign n19915 = ~n13752 & ~n19914 ;
  assign n19916 = ~\bdma_CMcnt_reg[0]/NET0131  & ~n19910 ;
  assign n19917 = ~n13752 & ~n19911 ;
  assign n19918 = ~n19916 & n19917 ;
  assign n19921 = ~n6917 & n13747 ;
  assign n19922 = ~\bdma_BCTL_reg[2]/NET0131  & n5533 ;
  assign n19923 = n5554 & n19922 ;
  assign n19924 = ~n19921 & n19923 ;
  assign n19919 = ~n6921 & ~n13151 ;
  assign n19920 = ~\bdma_BMcyc_del_reg/P0001  & ~n19919 ;
  assign n19925 = ~\bdma_BSreq_reg/NET0131  & ~n19920 ;
  assign n19926 = ~n19924 & n19925 ;
  assign n19927 = n17833 & ~n19771 ;
  assign n19928 = ~\core_eu_es_sht_es_reg_sr1rwe_DO_reg[15]/P0001  & ~n17833 ;
  assign n19929 = ~n19927 & ~n19928 ;
  assign n19933 = ~\sport0_regs_SCTLreg_DO_reg[11]/NET0131  & ~\sport0_regs_SCTLreg_DO_reg[12]/NET0131  ;
  assign n19934 = ~\ITFS0_pad  & \T_TFS0_pad  ;
  assign n19935 = \ITFS0_pad  & ~n13725 ;
  assign n19936 = ~n19934 & ~n19935 ;
  assign n19937 = \sport0_regs_SCTLreg_DO_reg[7]/NET0131  & ~n19936 ;
  assign n19938 = ~\sport0_regs_SCTLreg_DO_reg[7]/NET0131  & n19936 ;
  assign n19939 = ~n19937 & ~n19938 ;
  assign n19940 = \sport0_cfg_SP_ENg_reg/NET0131  & ~\sport0_cfg_TFSgi_d_reg/NET0131  ;
  assign n19941 = n19939 & n19940 ;
  assign n19942 = n19933 & ~n19941 ;
  assign n19944 = \sport0_cfg_TFSg_d3_reg/NET0131  & \sport0_regs_SCTLreg_DO_reg[11]/NET0131  ;
  assign n19943 = \sport0_cfg_TFSg_d2_reg/NET0131  & ~\sport0_regs_SCTLreg_DO_reg[11]/NET0131  ;
  assign n19945 = \sport0_regs_SCTLreg_DO_reg[12]/NET0131  & ~n19943 ;
  assign n19946 = ~n19944 & n19945 ;
  assign n19931 = ~\sport0_cfg_TFSg_d1_reg/NET0131  & \sport0_regs_SCTLreg_DO_reg[11]/NET0131  ;
  assign n19932 = ~\sport0_regs_SCTLreg_DO_reg[12]/NET0131  & n19931 ;
  assign n19947 = \sport0_txctl_TCS_reg[0]/NET0131  & ~n19932 ;
  assign n19948 = ~n19946 & n19947 ;
  assign n19949 = ~n19942 & n19948 ;
  assign n19950 = ~\sport0_txctl_TCS_reg[2]/NET0131  & ~n19949 ;
  assign n19930 = \sport0_txctl_TCS_reg[0]/NET0131  & \sport0_txctl_TCS_reg[2]/NET0131  ;
  assign n19951 = ~\sport0_txctl_TCS_reg[1]/NET0131  & ~n19930 ;
  assign n19952 = ~n19950 & n19951 ;
  assign n19953 = ~\sport0_txctl_TCS_reg[0]/NET0131  & \sport0_txctl_TCS_reg[1]/NET0131  ;
  assign n19954 = ~\sport0_txctl_TCS_reg[2]/NET0131  & n19953 ;
  assign n19955 = ~\sport0_txctl_Bcnt_reg[0]/NET0131  & ~\sport0_txctl_Bcnt_reg[1]/NET0131  ;
  assign n19956 = ~\sport0_txctl_Bcnt_reg[2]/NET0131  & n19955 ;
  assign n19957 = ~\sport0_txctl_Bcnt_reg[3]/NET0131  & n19956 ;
  assign n19958 = ~\sport0_txctl_Bcnt_reg[4]/NET0131  & n19957 ;
  assign n19959 = n19954 & ~n19958 ;
  assign n19960 = ~n19952 & ~n19959 ;
  assign n19961 = \sport0_txctl_TXSHT_reg[14]/P0001  & ~n19960 ;
  assign n19962 = \sport0_txctl_TX_reg[15]/P0001  & n19960 ;
  assign n19963 = ~n19961 & ~n19962 ;
  assign n19964 = n14752 & ~n19692 ;
  assign n19965 = n19559 & n19776 ;
  assign n19966 = \core_eu_em_mac_em_reg_mr1rwe_DO_reg[0]/P0001  & ~n17809 ;
  assign n19967 = n19780 & ~n19966 ;
  assign n19968 = ~n19965 & n19967 ;
  assign n19969 = ~n19964 & ~n19968 ;
  assign n19970 = ~\core_c_dec_accPM_E_reg/P0001  & ~n11265 ;
  assign n19971 = \core_c_dec_accPM_E_reg/P0001  & ~n13006 ;
  assign n19972 = ~n19970 & ~n19971 ;
  assign n19973 = \core_c_dec_MTSR1_E_reg/P0001  & ~n19972 ;
  assign n19984 = ~n17981 & n18720 ;
  assign n19985 = n18748 & ~n19984 ;
  assign n19993 = ~n18091 & ~n18991 ;
  assign n19994 = n18100 & ~n18180 ;
  assign n20011 = ~n19993 & ~n19994 ;
  assign n19998 = ~n18108 & n18166 ;
  assign n20002 = ~n17922 & ~n18189 ;
  assign n20012 = ~n19998 & ~n20002 ;
  assign n20013 = n20011 & n20012 ;
  assign n20022 = ~n18085 & n20013 ;
  assign n20023 = ~n19985 & n20022 ;
  assign n19978 = ~n17931 & n17986 ;
  assign n19979 = ~n18043 & ~n19978 ;
  assign n19980 = n18111 & ~n19979 ;
  assign n19981 = n18765 & ~n18775 ;
  assign n20016 = ~n19980 & ~n19981 ;
  assign n19988 = ~n18069 & ~n18725 ;
  assign n19989 = n18115 & ~n18149 ;
  assign n20017 = n19988 & ~n19989 ;
  assign n20020 = n20016 & n20017 ;
  assign n19974 = n18125 & n18132 ;
  assign n20000 = \core_c_dec_IRE_reg[11]/NET0131  & ~n11239 ;
  assign n20003 = ~n19974 & ~n20000 ;
  assign n19983 = n18103 & n18178 ;
  assign n20001 = n18106 & n18163 ;
  assign n20004 = ~n19983 & ~n20001 ;
  assign n20005 = n20003 & n20004 ;
  assign n20006 = ~n18040 & ~n18783 ;
  assign n20009 = n20005 & n20006 ;
  assign n19982 = n18128 & ~n18133 ;
  assign n20010 = n18054 & ~n19982 ;
  assign n20014 = n20009 & n20010 ;
  assign n19995 = n18125 & n18131 ;
  assign n19986 = n18103 & n18179 ;
  assign n19987 = n18107 & n18163 ;
  assign n20007 = ~n19986 & ~n19987 ;
  assign n20008 = ~n19995 & n20007 ;
  assign n20015 = n18727 & n20008 ;
  assign n20021 = n20014 & n20015 ;
  assign n20024 = n20020 & n20021 ;
  assign n20027 = n20023 & n20024 ;
  assign n20028 = n18791 & n20027 ;
  assign n19975 = ~n18060 & n18797 ;
  assign n19976 = ~n17964 & n18195 ;
  assign n19977 = n19975 & n19976 ;
  assign n19999 = n18724 & ~n18735 ;
  assign n19996 = ~n18002 & ~n18737 ;
  assign n19997 = n17978 & n19996 ;
  assign n19992 = n18088 & ~n19818 ;
  assign n19990 = n17925 & ~n19857 ;
  assign n19991 = n17945 & ~n18781 ;
  assign n20018 = ~n19990 & ~n19991 ;
  assign n20019 = ~n19992 & n20018 ;
  assign n20025 = n19997 & n20019 ;
  assign n20026 = n19999 & n20025 ;
  assign n20029 = n19977 & n20026 ;
  assign n20030 = n20028 & n20029 ;
  assign n20031 = ~\core_c_dec_MTSR1_E_reg/P0001  & n20030 ;
  assign n20032 = ~n19973 & ~n20031 ;
  assign n20033 = n18717 & ~n20032 ;
  assign n20034 = ~\core_eu_es_sht_es_reg_sr1swe_DO_reg[7]/P0001  & ~n18717 ;
  assign n20035 = ~n20033 & ~n20034 ;
  assign n20036 = ~\bdma_BSreq_reg/NET0131  & n5534 ;
  assign n20037 = \bdma_BWcnt_reg[0]/NET0131  & \bdma_BWcnt_reg[1]/NET0131  ;
  assign n20038 = n20036 & n20037 ;
  assign n20039 = \bdma_BWcnt_reg[2]/NET0131  & n20038 ;
  assign n20040 = \bdma_BWcnt_reg[3]/NET0131  & n20039 ;
  assign n20041 = ~\bdma_BWcnt_reg[4]/NET0131  & ~n20040 ;
  assign n20042 = \bdma_BWcnt_reg[4]/NET0131  & n20040 ;
  assign n20043 = ~n20041 & ~n20042 ;
  assign n20044 = ~n13750 & n20043 ;
  assign n20045 = ~n13806 & ~n14424 ;
  assign n20046 = ~n13809 & ~n14321 ;
  assign n20048 = ~n14362 & n14404 ;
  assign n20047 = n14362 & ~n14406 ;
  assign n20049 = ~n14358 & ~n20047 ;
  assign n20050 = ~n20048 & n20049 ;
  assign n20051 = n20046 & ~n20050 ;
  assign n20052 = ~n20046 & n20050 ;
  assign n20053 = ~n20051 & ~n20052 ;
  assign n20054 = n13806 & ~n20053 ;
  assign n20055 = ~n20045 & ~n20054 ;
  assign n20056 = n14667 & ~n20055 ;
  assign n20057 = \core_eu_ea_alu_ea_reg_afswe_DO_reg[11]/P0001  & ~n14667 ;
  assign n20058 = ~n20056 & ~n20057 ;
  assign n20059 = n13805 & ~n20055 ;
  assign n20060 = \core_eu_ea_alu_ea_reg_afrwe_DO_reg[11]/P0001  & ~n13805 ;
  assign n20061 = ~n20059 & ~n20060 ;
  assign n20065 = \idma_IAL_reg/P0001  & ~\idma_ISn_reg/P0001  ;
  assign n20066 = \idma_IADi_reg[15]/P0001  & n20065 ;
  assign n20067 = n7530 & n18226 ;
  assign n20068 = ~n20066 & ~n20067 ;
  assign n20069 = ~\idma_IADi_reg[15]/P0001  & n20065 ;
  assign n20070 = ~\core_dag_ilm1reg_DMA_pi_DO_reg[2]/NET0131  & ~\core_dag_ilm1reg_DMA_pi_DO_reg[3]/NET0131  ;
  assign n20071 = n7261 & n20070 ;
  assign n20072 = n13762 & n20071 ;
  assign n20073 = ~n20069 & ~n20072 ;
  assign n20074 = n20068 & n20073 ;
  assign n20062 = ~\idma_DCTL_reg[14]/NET0131  & \idma_RDCMD_d1_reg/P0001  ;
  assign n20063 = ~\idma_RDCMD_reg/P0001  & n20062 ;
  assign n20064 = ~\idma_PCrd_1st_reg/NET0131  & n20063 ;
  assign n20075 = \idma_PCrd_1st_reg/NET0131  & ~n20063 ;
  assign n20076 = ~n20064 & ~n20075 ;
  assign n20077 = n20074 & n20076 ;
  assign n20078 = ~\core_c_dec_accPM_E_reg/P0001  & ~n10069 ;
  assign n20079 = \core_c_dec_accPM_E_reg/P0001  & ~n12904 ;
  assign n20080 = ~n20078 & ~n20079 ;
  assign n20081 = \core_c_dec_MTSR1_E_reg/P0001  & ~n20080 ;
  assign n20106 = n18054 & n18790 ;
  assign n20107 = n18738 & n20106 ;
  assign n20103 = ~n18091 & ~n18919 ;
  assign n20098 = n18046 & n18171 ;
  assign n20100 = n18043 & n18758 ;
  assign n20126 = ~n20098 & ~n20100 ;
  assign n20127 = ~n20103 & n20126 ;
  assign n20092 = n17925 & n17980 ;
  assign n20089 = n18153 & n19863 ;
  assign n20099 = n18106 & ~n18743 ;
  assign n20115 = ~n20089 & ~n20099 ;
  assign n20102 = n18132 & n18752 ;
  assign n20111 = n17986 & n18754 ;
  assign n20116 = ~n20102 & ~n20111 ;
  assign n20117 = n20115 & n20116 ;
  assign n20124 = ~n20092 & n20117 ;
  assign n20093 = n18147 & ~n18182 ;
  assign n20096 = ~n18746 & ~n18763 ;
  assign n20097 = ~n17922 & ~n20096 ;
  assign n20125 = ~n20093 & ~n20097 ;
  assign n20128 = n20124 & n20125 ;
  assign n20135 = n20127 & n20128 ;
  assign n20084 = ~n18141 & ~n18783 ;
  assign n20085 = ~n17977 & ~n18900 ;
  assign n20086 = n20084 & n20085 ;
  assign n20087 = n19988 & n20086 ;
  assign n20112 = n17945 & ~n17962 ;
  assign n20136 = n20087 & ~n20112 ;
  assign n20137 = n20135 & n20136 ;
  assign n20104 = n17931 & ~n18907 ;
  assign n20105 = ~n17938 & n20104 ;
  assign n20108 = n18038 & ~n19787 ;
  assign n20131 = ~n20105 & n20108 ;
  assign n20109 = n18748 & ~n19818 ;
  assign n20113 = n18765 & ~n18895 ;
  assign n20132 = ~n20109 & ~n20113 ;
  assign n20133 = n20131 & n20132 ;
  assign n20091 = n17951 & n17976 ;
  assign n20094 = n18758 & n18761 ;
  assign n20120 = ~n20091 & ~n20094 ;
  assign n20095 = n18131 & n18752 ;
  assign n20110 = ~n17924 & n18780 ;
  assign n20121 = ~n20095 & ~n20110 ;
  assign n20122 = n20120 & n20121 ;
  assign n20083 = \core_c_dec_IRE_reg[11]/NET0131  & ~n9947 ;
  assign n20114 = ~n18192 & ~n20083 ;
  assign n20118 = ~n17972 & n20114 ;
  assign n20088 = n18107 & ~n18743 ;
  assign n20119 = ~n18040 & ~n20088 ;
  assign n20123 = n20118 & n20119 ;
  assign n20129 = n20122 & n20123 ;
  assign n20082 = n18115 & ~n19857 ;
  assign n20101 = n18111 & ~n18775 ;
  assign n20130 = ~n20082 & ~n20101 ;
  assign n20134 = n20129 & n20130 ;
  assign n20138 = n20133 & n20134 ;
  assign n20139 = n20137 & n20138 ;
  assign n20090 = n18145 & n19789 ;
  assign n20140 = n19975 & n20090 ;
  assign n20141 = n20139 & n20140 ;
  assign n20142 = n20107 & n20141 ;
  assign n20143 = ~\core_c_dec_MTSR1_E_reg/P0001  & n20142 ;
  assign n20144 = ~n20081 & ~n20143 ;
  assign n20145 = n18717 & ~n20144 ;
  assign n20146 = ~\core_eu_es_sht_es_reg_sr1swe_DO_reg[4]/P0001  & ~n18717 ;
  assign n20147 = ~n20145 & ~n20146 ;
  assign n20148 = ~\core_c_dec_accPM_E_reg/P0001  & ~n12688 ;
  assign n20149 = \core_c_dec_accPM_E_reg/P0001  & ~n12715 ;
  assign n20150 = ~n20148 & ~n20149 ;
  assign n20151 = \core_c_dec_MTSR1_E_reg/P0001  & ~n20150 ;
  assign n20153 = ~n17922 & n18766 ;
  assign n20154 = n18106 & n18905 ;
  assign n20174 = \core_c_dec_IRE_reg[11]/NET0131  & ~n11854 ;
  assign n20178 = ~n20154 & ~n20174 ;
  assign n20179 = ~n20153 & n20178 ;
  assign n20155 = ~n18159 & ~n18919 ;
  assign n20156 = ~n18121 & n18746 ;
  assign n20180 = ~n20155 & ~n20156 ;
  assign n20183 = n20179 & n20180 ;
  assign n20152 = ~n17938 & n18176 ;
  assign n20184 = n18059 & ~n20152 ;
  assign n20185 = n20183 & n20184 ;
  assign n20176 = ~n18092 & n19725 ;
  assign n20177 = n17945 & ~n20176 ;
  assign n20175 = ~n18108 & n18749 ;
  assign n20157 = ~n18096 & ~n18743 ;
  assign n20158 = ~n18133 & n19862 ;
  assign n20181 = ~n20157 & ~n20158 ;
  assign n20182 = ~n20175 & n20181 ;
  assign n20186 = ~n20177 & n20182 ;
  assign n20187 = n20185 & n20186 ;
  assign n20188 = n18006 & n20187 ;
  assign n20160 = ~n17922 & ~n17924 ;
  assign n20162 = n18107 & ~n18110 ;
  assign n20165 = n17931 & ~n20162 ;
  assign n20166 = ~n20160 & n20165 ;
  assign n20164 = ~n18180 & ~n18182 ;
  assign n20161 = ~n18121 & ~n18123 ;
  assign n20163 = ~n18133 & ~n18170 ;
  assign n20167 = ~n20161 & ~n20163 ;
  assign n20168 = ~n20164 & n20167 ;
  assign n20169 = n20166 & n20168 ;
  assign n20170 = n18751 & ~n19735 ;
  assign n20171 = ~n17931 & ~n19747 ;
  assign n20172 = ~n20170 & n20171 ;
  assign n20173 = ~n20169 & ~n20172 ;
  assign n20189 = n18087 & ~n20173 ;
  assign n20190 = n20188 & n20189 ;
  assign n20159 = n18146 & n19976 ;
  assign n20191 = n19715 & n20159 ;
  assign n20192 = n20190 & n20191 ;
  assign n20193 = ~\core_c_dec_MTSR1_E_reg/P0001  & n20192 ;
  assign n20194 = ~n20151 & ~n20193 ;
  assign n20195 = n18717 & ~n20194 ;
  assign n20196 = ~\core_eu_es_sht_es_reg_sr1swe_DO_reg[14]/P0001  & ~n18717 ;
  assign n20197 = ~n20195 & ~n20196 ;
  assign n20198 = n17833 & ~n20032 ;
  assign n20199 = ~\core_eu_es_sht_es_reg_sr1rwe_DO_reg[7]/P0001  & ~n17833 ;
  assign n20200 = ~n20198 & ~n20199 ;
  assign n20205 = ~n5581 & n13749 ;
  assign n20208 = ~n5586 & n20205 ;
  assign n20209 = ~n5582 & n20208 ;
  assign n20206 = n5586 & n20205 ;
  assign n20207 = ~n12444 & n20206 ;
  assign n20201 = ~n5581 & ~n5586 ;
  assign n20202 = ~n5519 & ~n5587 ;
  assign n20203 = ~n20201 & n20202 ;
  assign n20204 = n5605 & n20203 ;
  assign n20210 = ~n13750 & ~n20204 ;
  assign n20211 = ~n20207 & n20210 ;
  assign n20212 = ~n20209 & n20211 ;
  assign n20213 = ~n5523 & n5583 ;
  assign n20214 = \emc_RWcnt_reg[0]/P0001  & ~n20213 ;
  assign n20215 = \emc_RWcnt_reg[1]/P0001  & n20214 ;
  assign n20216 = \emc_RWcnt_reg[2]/P0001  & n20215 ;
  assign n20217 = \emc_RWcnt_reg[3]/P0001  & n20216 ;
  assign n20218 = \emc_RWcnt_reg[4]/P0001  & n20217 ;
  assign n20219 = ~\emc_RWcnt_reg[5]/P0001  & ~n20218 ;
  assign n20220 = \emc_RWcnt_reg[5]/P0001  & n20218 ;
  assign n20221 = ~n20219 & ~n20220 ;
  assign n20222 = n20212 & n20221 ;
  assign n20223 = ~\emc_RWcnt_reg[4]/P0001  & ~n20217 ;
  assign n20224 = ~n20218 & ~n20223 ;
  assign n20225 = n20212 & n20224 ;
  assign n20226 = n17833 & ~n20144 ;
  assign n20227 = ~\core_eu_es_sht_es_reg_sr1rwe_DO_reg[4]/P0001  & ~n17833 ;
  assign n20228 = ~n20226 & ~n20227 ;
  assign n20229 = n17833 & ~n20194 ;
  assign n20230 = ~\core_eu_es_sht_es_reg_sr1rwe_DO_reg[14]/P0001  & ~n17833 ;
  assign n20231 = ~n20229 & ~n20230 ;
  assign n20232 = \sport1_cfg_SCLKi_cnt_reg[2]/NET0131  & n19438 ;
  assign n20233 = \sport1_cfg_SCLKi_cnt_reg[3]/NET0131  & n20232 ;
  assign n20234 = \sport1_cfg_SCLKi_cnt_reg[4]/NET0131  & n20233 ;
  assign n20235 = \sport1_cfg_SCLKi_cnt_reg[5]/NET0131  & n20234 ;
  assign n20236 = \sport1_cfg_SCLKi_cnt_reg[6]/NET0131  & n20235 ;
  assign n20237 = \sport1_cfg_SCLKi_cnt_reg[7]/NET0131  & n20236 ;
  assign n20238 = \sport1_cfg_SCLKi_cnt_reg[8]/NET0131  & n20237 ;
  assign n20240 = \sport1_cfg_SCLKi_cnt_reg[9]/NET0131  & n20238 ;
  assign n20239 = ~\sport1_cfg_SCLKi_cnt_reg[9]/NET0131  & ~n20238 ;
  assign n20241 = n19130 & ~n20239 ;
  assign n20242 = ~n20240 & n20241 ;
  assign n20243 = ~\sport1_cfg_SCLKi_cnt_reg[5]/NET0131  & ~n20234 ;
  assign n20244 = ~n20235 & ~n20243 ;
  assign n20245 = n19130 & n20244 ;
  assign n20246 = ~\sport1_cfg_SCLKi_cnt_reg[2]/NET0131  & ~n19438 ;
  assign n20247 = ~n20232 & ~n20246 ;
  assign n20248 = n19130 & n20247 ;
  assign n20249 = \sport1_cfg_SCLKi_cnt_reg[10]/NET0131  & n20240 ;
  assign n20250 = \sport1_cfg_SCLKi_cnt_reg[11]/NET0131  & n20249 ;
  assign n20251 = \sport1_cfg_SCLKi_cnt_reg[12]/NET0131  & n20250 ;
  assign n20253 = \sport1_cfg_SCLKi_cnt_reg[13]/NET0131  & n20251 ;
  assign n20252 = ~\sport1_cfg_SCLKi_cnt_reg[13]/NET0131  & ~n20251 ;
  assign n20254 = n19130 & ~n20252 ;
  assign n20255 = ~n20253 & n20254 ;
  assign n20256 = ~\sport1_cfg_SCLKi_cnt_reg[0]/NET0131  & n19130 ;
  assign n20257 = ~\core_c_dec_accPM_E_reg/P0001  & ~n10911 ;
  assign n20258 = \core_c_dec_accPM_E_reg/P0001  & ~n12938 ;
  assign n20259 = ~n20257 & ~n20258 ;
  assign n20260 = \core_c_dec_MTSR0_E_reg/P0001  & ~n20259 ;
  assign n20274 = n18797 & n18904 ;
  assign n20270 = ~n17933 & n18922 ;
  assign n20267 = ~n17998 & n18758 ;
  assign n20268 = n18171 & ~n18898 ;
  assign n20283 = ~n20267 & ~n20268 ;
  assign n20284 = ~n20270 & n20283 ;
  assign n20273 = ~n18129 & ~n18912 ;
  assign n20269 = ~n18104 & ~n18907 ;
  assign n20271 = n17991 & n18088 ;
  assign n20279 = ~n20269 & ~n20271 ;
  assign n20280 = ~n20273 & n20279 ;
  assign n20262 = ~n18167 & ~n18918 ;
  assign n20263 = n17930 & ~n18909 ;
  assign n20277 = ~n20262 & ~n20263 ;
  assign n20265 = ~n18189 & ~n18914 ;
  assign n20266 = ~n18079 & ~n18117 ;
  assign n20278 = ~n20265 & ~n20266 ;
  assign n20281 = n20277 & n20278 ;
  assign n20261 = n18765 & ~n18888 ;
  assign n20264 = \core_c_dec_IRE_reg[11]/NET0131  & ~n10801 ;
  assign n20272 = n17965 & n17992 ;
  assign n20275 = ~n20264 & ~n20272 ;
  assign n20276 = ~n18890 & n20275 ;
  assign n20282 = ~n20261 & n20276 ;
  assign n20285 = n20281 & n20282 ;
  assign n20286 = n20280 & n20285 ;
  assign n20287 = n20284 & n20286 ;
  assign n20288 = n20274 & n20287 ;
  assign n20289 = ~\core_c_dec_MTSR0_E_reg/P0001  & n20288 ;
  assign n20290 = ~n20260 & ~n20289 ;
  assign n20291 = n18886 & ~n20290 ;
  assign n20292 = ~\core_eu_es_sht_es_reg_sr0swe_DO_reg[5]/P0001  & ~n18886 ;
  assign n20293 = ~n20291 & ~n20292 ;
  assign n20294 = \core_c_dec_MTSR0_E_reg/P0001  & ~n19559 ;
  assign n20298 = n18765 & ~n18981 ;
  assign n20302 = n17925 & ~n18983 ;
  assign n20321 = ~n20298 & ~n20302 ;
  assign n20303 = n18171 & ~n18888 ;
  assign n20306 = ~n17998 & n18124 ;
  assign n20322 = ~n20303 & ~n20306 ;
  assign n20323 = n20321 & n20322 ;
  assign n20301 = n17991 & n18115 ;
  assign n20305 = n18754 & ~n18909 ;
  assign n20316 = ~n20301 & ~n20305 ;
  assign n20307 = n18752 & ~n18918 ;
  assign n20308 = n17929 & n18088 ;
  assign n20309 = ~n17965 & ~n20308 ;
  assign n20310 = ~n17970 & ~n18017 ;
  assign n20311 = ~n20309 & ~n20310 ;
  assign n20317 = ~n20307 & ~n20311 ;
  assign n20318 = n20316 & n20317 ;
  assign n20295 = n18759 & ~n18909 ;
  assign n20297 = ~n18082 & ~n19870 ;
  assign n20314 = ~n20295 & ~n20297 ;
  assign n20299 = ~n18079 & ~n18919 ;
  assign n20300 = ~n18743 & ~n18914 ;
  assign n20315 = ~n20299 & ~n20300 ;
  assign n20319 = n20314 & n20315 ;
  assign n20296 = n18745 & ~n18898 ;
  assign n20304 = \core_c_dec_IRE_reg[11]/NET0131  & ~n7381 ;
  assign n20312 = ~n18900 & ~n20304 ;
  assign n20313 = n18016 & n20312 ;
  assign n20320 = ~n20296 & n20313 ;
  assign n20324 = n20319 & n20320 ;
  assign n20325 = n20318 & n20324 ;
  assign n20326 = n20323 & n20325 ;
  assign n20327 = ~\core_c_dec_MTSR0_E_reg/P0001  & n20326 ;
  assign n20328 = ~n20294 & ~n20327 ;
  assign n20329 = n18886 & ~n20328 ;
  assign n20330 = ~\core_eu_es_sht_es_reg_sr0swe_DO_reg[0]/P0001  & ~n18886 ;
  assign n20331 = ~n20329 & ~n20330 ;
  assign n20332 = n19034 & ~n20290 ;
  assign n20333 = ~\core_eu_es_sht_es_reg_sr0rwe_DO_reg[5]/P0001  & ~n19034 ;
  assign n20334 = ~n20332 & ~n20333 ;
  assign n20335 = n19034 & ~n20328 ;
  assign n20336 = ~\core_eu_es_sht_es_reg_sr0rwe_DO_reg[0]/P0001  & ~n19034 ;
  assign n20337 = ~n20335 & ~n20336 ;
  assign n20338 = ~\sport0_cfg_SCLKi_cnt_reg[9]/NET0131  & ~n19546 ;
  assign n20339 = n19197 & ~n19547 ;
  assign n20340 = ~n20338 & n20339 ;
  assign n20341 = \emc_PMcst_reg/NET0131  & n14733 ;
  assign n20342 = \core_c_psq_PMOVL_regh_DO_reg[3]/NET0131  & ~n4068 ;
  assign n20343 = n19041 & n20342 ;
  assign n20344 = \memc_Pread_E_reg/NET0131  & n20343 ;
  assign n20345 = n19049 & n20344 ;
  assign n20351 = ~n20341 & ~n20345 ;
  assign n20346 = \memc_Pwrite_E_reg/NET0131  & n20343 ;
  assign n20347 = n19049 & n20346 ;
  assign n20348 = \emc_PMcst_reg/NET0131  & ~n5593 ;
  assign n20349 = ~n5604 & n20348 ;
  assign n20350 = ~n19049 & n20349 ;
  assign n20352 = ~n20347 & ~n20350 ;
  assign n20353 = n20351 & n20352 ;
  assign n20358 = ~\tm_TCR_TMP_reg[1]/NET0131  & ~\tm_TCR_TMP_reg[2]/NET0131  ;
  assign n20359 = ~\tm_TCR_TMP_reg[3]/NET0131  & n20358 ;
  assign n20360 = ~\tm_TCR_TMP_reg[0]/NET0131  & n20359 ;
  assign n20361 = ~\tm_TCR_TMP_reg[4]/NET0131  & ~\tm_TCR_TMP_reg[5]/NET0131  ;
  assign n20362 = ~\tm_TCR_TMP_reg[6]/NET0131  & ~\tm_TCR_TMP_reg[7]/NET0131  ;
  assign n20363 = n20361 & n20362 ;
  assign n20364 = n20360 & n20363 ;
  assign n20367 = ~\tm_TCR_TMP_reg[14]/NET0131  & ~\tm_TCR_TMP_reg[15]/NET0131  ;
  assign n20368 = ~\tm_TCR_TMP_reg[8]/NET0131  & ~\tm_TCR_TMP_reg[9]/NET0131  ;
  assign n20369 = n20367 & n20368 ;
  assign n20365 = ~\tm_TCR_TMP_reg[10]/NET0131  & ~\tm_TCR_TMP_reg[11]/NET0131  ;
  assign n20366 = ~\tm_TCR_TMP_reg[12]/NET0131  & ~\tm_TCR_TMP_reg[13]/NET0131  ;
  assign n20370 = n20365 & n20366 ;
  assign n20371 = n20369 & n20370 ;
  assign n20372 = n20364 & n20371 ;
  assign n20356 = ~\T_TMODE[0]_pad  & \tm_WR_TSR_TMP_GEN1_reg/P0001  ;
  assign n20357 = ~\tm_WR_TSR_TMP_GEN2_reg/P0001  & n20356 ;
  assign n20354 = ~\T_TMODE[0]_pad  & \tm_WR_TCR_TMP_GEN1_reg/P0001  ;
  assign n20355 = ~\tm_WR_TCR_TMP_GEN2_reg/P0001  & n20354 ;
  assign n20373 = \tm_MSTAT5_syn_reg/NET0131  & ~n20355 ;
  assign n20374 = ~n20357 & n20373 ;
  assign n20375 = n20372 & n20374 ;
  assign n20376 = \core_c_dec_updAF_E_reg/P0001  & n4118 ;
  assign n20377 = n5664 & ~n18842 ;
  assign n20378 = n4116 & n18849 ;
  assign n20379 = n20377 & n20378 ;
  assign n20380 = ~n20376 & ~n20379 ;
  assign n20381 = ~\idma_WRcnt_reg[0]/NET0131  & ~\idma_WRcnt_reg[1]/NET0131  ;
  assign n20382 = ~\idma_WRcnt_reg[2]/NET0131  & n20381 ;
  assign n20383 = \idma_WRtrue_reg/NET0131  & ~n20382 ;
  assign n20384 = ~\idma_WRCMD_d1_reg/P0001  & \idma_WRCMD_reg/P0001  ;
  assign n20385 = ~n20383 & ~n20384 ;
  assign n20386 = ~\idma_DCTL_reg[14]/NET0131  & ~\idma_PM_1st_reg/NET0131  ;
  assign n20387 = ~\idma_ISn_reg/P0001  & ~\idma_IWRn_reg/P0001  ;
  assign n20388 = \idma_WRtrue_reg/NET0131  & n20387 ;
  assign n20389 = \auctl_DSack_reg/NET0131  & ~n20386 ;
  assign n20390 = ~\idma_RDcnt_reg[0]/NET0131  & ~\idma_RDcnt_reg[1]/NET0131  ;
  assign n20391 = ~\idma_RDcnt_reg[2]/NET0131  & n20386 ;
  assign n20392 = n20390 & n20391 ;
  assign n20393 = ~n20389 & ~n20392 ;
  assign n20394 = \idma_RDcyc_reg/NET0131  & ~n20393 ;
  assign n20395 = ~n20388 & ~n20394 ;
  assign n20396 = ~n20386 & ~n20395 ;
  assign n20397 = \core_eu_em_mac_em_dec_emcorepi_DO_reg[0]/P0001  & ~n18848 ;
  assign n20398 = n18843 & n18848 ;
  assign n20399 = ~n20397 & ~n20398 ;
  assign n20400 = n7226 & n20070 ;
  assign n20401 = n18226 & n20400 ;
  assign n20402 = ~\memc_MMR_web_reg/NET0131  & n20401 ;
  assign n20403 = ~n10289 & n20402 ;
  assign n20404 = ~\sport0_regs_AUTOreg_DO_reg[9]/NET0131  & ~n20402 ;
  assign n20405 = ~n20403 & ~n20404 ;
  assign n20406 = ~\sport1_rxctl_Wcnt_reg[4]/NET0131  & ~\sport1_rxctl_Wcnt_reg[5]/NET0131  ;
  assign n20407 = ~\sport1_rxctl_Wcnt_reg[6]/NET0131  & n20406 ;
  assign n20408 = ~\sport1_rxctl_Wcnt_reg[7]/NET0131  & n20407 ;
  assign n20411 = \sport1_rxctl_Wcnt_reg[0]/NET0131  & \sport1_rxctl_Wcnt_reg[1]/NET0131  ;
  assign n20412 = ~\sport1_rxctl_Wcnt_reg[2]/NET0131  & \sport1_rxctl_Wcnt_reg[3]/NET0131  ;
  assign n20413 = n20411 & n20412 ;
  assign n20409 = \sport1_rxctl_Bcnt_reg[1]/NET0131  & ~\sport1_rxctl_Bcnt_reg[2]/NET0131  ;
  assign n20410 = ~\sport1_rxctl_Bcnt_reg[3]/NET0131  & ~\sport1_rxctl_Bcnt_reg[4]/NET0131  ;
  assign n20414 = n20409 & n20410 ;
  assign n20415 = n20413 & n20414 ;
  assign n20416 = n20408 & n20415 ;
  assign n20417 = ~\sport1_rxctl_Bcnt_reg[0]/NET0131  & n20416 ;
  assign n20418 = \sport1_regs_SCTLreg_DO_reg[15]/NET0131  & ~n13720 ;
  assign n20419 = ~\T_RD1_pad  & ~\sport1_regs_SCTLreg_DO_reg[15]/NET0131  ;
  assign n20420 = ~n20418 & ~n20419 ;
  assign n20421 = n20417 & ~n20420 ;
  assign n20422 = ~\sport1_rxctl_SLOT1_EXT_reg[2]/NET0131  & ~n20417 ;
  assign n20423 = ~n20421 & ~n20422 ;
  assign n20424 = \sport1_rxctl_Bcnt_reg[0]/NET0131  & n20416 ;
  assign n20425 = ~n20420 & n20424 ;
  assign n20426 = ~\sport1_rxctl_SLOT1_EXT_reg[3]/NET0131  & ~n20424 ;
  assign n20427 = ~n20425 & ~n20426 ;
  assign n20428 = ~\sport0_rxctl_Wcnt_reg[4]/NET0131  & ~\sport0_rxctl_Wcnt_reg[5]/NET0131  ;
  assign n20429 = ~\sport0_rxctl_Wcnt_reg[6]/NET0131  & n20428 ;
  assign n20430 = ~\sport0_rxctl_Wcnt_reg[7]/NET0131  & n20429 ;
  assign n20433 = \sport0_rxctl_Wcnt_reg[0]/NET0131  & \sport0_rxctl_Wcnt_reg[1]/NET0131  ;
  assign n20434 = ~\sport0_rxctl_Wcnt_reg[2]/NET0131  & \sport0_rxctl_Wcnt_reg[3]/NET0131  ;
  assign n20435 = n20433 & n20434 ;
  assign n20431 = \sport0_rxctl_Bcnt_reg[1]/NET0131  & ~\sport0_rxctl_Bcnt_reg[2]/NET0131  ;
  assign n20432 = ~\sport0_rxctl_Bcnt_reg[3]/NET0131  & ~\sport0_rxctl_Bcnt_reg[4]/NET0131  ;
  assign n20436 = n20431 & n20432 ;
  assign n20437 = n20435 & n20436 ;
  assign n20438 = n20430 & n20437 ;
  assign n20439 = ~\sport0_rxctl_Bcnt_reg[0]/NET0131  & n20438 ;
  assign n20440 = \sport0_regs_SCTLreg_DO_reg[15]/NET0131  & ~n13671 ;
  assign n20441 = ~\T_RD0_pad  & ~\sport0_regs_SCTLreg_DO_reg[15]/NET0131  ;
  assign n20442 = ~n20440 & ~n20441 ;
  assign n20443 = n20439 & ~n20442 ;
  assign n20444 = ~\sport0_rxctl_SLOT1_EXT_reg[2]/NET0131  & ~n20439 ;
  assign n20445 = ~n20443 & ~n20444 ;
  assign n20446 = \sport0_rxctl_Bcnt_reg[0]/NET0131  & n20438 ;
  assign n20447 = ~n20442 & n20446 ;
  assign n20448 = ~\sport0_rxctl_SLOT1_EXT_reg[3]/NET0131  & ~n20446 ;
  assign n20449 = ~n20447 & ~n20448 ;
  assign n20450 = ~n10638 & n20402 ;
  assign n20451 = ~\sport0_regs_AUTOreg_DO_reg[8]/NET0131  & ~n20402 ;
  assign n20452 = ~n20450 & ~n20451 ;
  assign n20453 = ~IACKn_pad & \idma_IRDn_reg/P0001  ;
  assign n20454 = \idma_IWRn_reg/P0001  & n20453 ;
  assign n20456 = \idma_WRtrue_reg/NET0131  & ~n20454 ;
  assign n20457 = ~\idma_WRcnt_reg[0]/NET0131  & n20456 ;
  assign n20458 = \idma_WRcnt_reg[1]/NET0131  & ~n20457 ;
  assign n20455 = n20384 & ~n20454 ;
  assign n20459 = n20381 & n20456 ;
  assign n20460 = ~n20455 & ~n20459 ;
  assign n20461 = ~n20458 & n20460 ;
  assign n20462 = ~\memc_usysr_DO_reg[8]/NET0131  & n20455 ;
  assign n20463 = ~n20461 & ~n20462 ;
  assign n20464 = ~\core_c_dec_IR_reg[5]/NET0131  & ~\core_c_dec_IR_reg[6]/NET0131  ;
  assign n20465 = ~\core_c_dec_IR_reg[4]/NET0131  & ~\core_c_dec_IR_reg[7]/NET0131  ;
  assign n20466 = n20464 & n20465 ;
  assign n20467 = n14728 & ~n20466 ;
  assign n20468 = n5664 & n20467 ;
  assign n20469 = \core_eu_ea_alu_ea_dec_piconst_DO_reg[9]/P0001  & ~n20468 ;
  assign n20470 = ~\core_c_dec_IR_reg[11]/NET0131  & \core_c_dec_IR_reg[12]/NET0131  ;
  assign n20471 = ~\core_c_dec_IR_reg[7]/NET0131  & n20470 ;
  assign n20475 = \core_c_dec_IR_reg[4]/NET0131  & \core_c_dec_IR_reg[5]/NET0131  ;
  assign n20476 = ~n20471 & n20475 ;
  assign n20472 = \core_c_dec_IR_reg[4]/NET0131  & ~\core_c_dec_IR_reg[5]/NET0131  ;
  assign n20473 = \core_c_dec_IR_reg[6]/NET0131  & n20472 ;
  assign n20474 = n20471 & n20473 ;
  assign n20477 = \core_c_dec_IR_reg[5]/NET0131  & ~\core_c_dec_IR_reg[6]/NET0131  ;
  assign n20478 = \core_c_dec_IR_reg[4]/NET0131  & n20477 ;
  assign n20479 = ~n20474 & ~n20478 ;
  assign n20480 = ~n20476 & n20479 ;
  assign n20481 = n20468 & ~n20480 ;
  assign n20482 = ~n20469 & ~n20481 ;
  assign n20483 = \core_eu_ea_alu_ea_dec_piconst_DO_reg[8]/P0001  & ~n20468 ;
  assign n20484 = \core_c_dec_IR_reg[4]/NET0131  & n20464 ;
  assign n20485 = n20471 & n20484 ;
  assign n20486 = \core_c_dec_IR_reg[5]/NET0131  & \core_c_dec_IR_reg[6]/NET0131  ;
  assign n20487 = \core_c_dec_IR_reg[4]/NET0131  & n20486 ;
  assign n20488 = ~n20476 & ~n20487 ;
  assign n20489 = ~n20485 & n20488 ;
  assign n20490 = n20468 & ~n20489 ;
  assign n20491 = ~n20483 & ~n20490 ;
  assign n20492 = \core_eu_ea_alu_ea_dec_piconst_DO_reg[7]/P0001  & ~n20468 ;
  assign n20493 = \core_c_dec_IR_reg[11]/NET0131  & ~\core_c_dec_IR_reg[12]/NET0131  ;
  assign n20494 = \core_c_dec_IR_reg[7]/NET0131  & n20493 ;
  assign n20496 = n20473 & n20494 ;
  assign n20495 = n20475 & ~n20494 ;
  assign n20497 = ~n20478 & ~n20495 ;
  assign n20498 = ~n20496 & n20497 ;
  assign n20499 = n20468 & ~n20498 ;
  assign n20500 = ~n20492 & ~n20499 ;
  assign n20501 = \core_eu_ea_alu_ea_dec_piconst_DO_reg[6]/P0001  & ~n20468 ;
  assign n20502 = n20484 & n20494 ;
  assign n20503 = ~n20487 & ~n20495 ;
  assign n20504 = ~n20502 & n20503 ;
  assign n20505 = n20468 & ~n20504 ;
  assign n20506 = ~n20501 & ~n20505 ;
  assign n20507 = \core_eu_ea_alu_ea_dec_piconst_DO_reg[5]/P0001  & ~n20468 ;
  assign n20508 = ~\core_c_dec_IR_reg[12]/NET0131  & ~\core_c_dec_IR_reg[7]/NET0131  ;
  assign n20509 = \core_c_dec_IR_reg[11]/NET0131  & n20508 ;
  assign n20511 = n20473 & n20509 ;
  assign n20510 = n20475 & ~n20509 ;
  assign n20512 = ~n20478 & ~n20510 ;
  assign n20513 = ~n20511 & n20512 ;
  assign n20514 = n20468 & ~n20513 ;
  assign n20515 = ~n20507 & ~n20514 ;
  assign n20516 = \core_eu_ea_alu_ea_dec_piconst_DO_reg[4]/P0001  & ~n20468 ;
  assign n20517 = n20484 & n20509 ;
  assign n20518 = ~n20487 & ~n20510 ;
  assign n20519 = ~n20517 & n20518 ;
  assign n20520 = n20468 & ~n20519 ;
  assign n20521 = ~n20516 & ~n20520 ;
  assign n20522 = \core_eu_ea_alu_ea_dec_piconst_DO_reg[3]/P0001  & ~n20468 ;
  assign n20523 = ~\core_c_dec_IR_reg[11]/NET0131  & ~\core_c_dec_IR_reg[12]/NET0131  ;
  assign n20524 = \core_c_dec_IR_reg[7]/NET0131  & n20523 ;
  assign n20526 = n20473 & n20524 ;
  assign n20525 = n20475 & ~n20524 ;
  assign n20527 = ~n20478 & ~n20525 ;
  assign n20528 = ~n20526 & n20527 ;
  assign n20529 = n20468 & ~n20528 ;
  assign n20530 = ~n20522 & ~n20529 ;
  assign n20531 = \core_eu_ea_alu_ea_dec_piconst_DO_reg[2]/P0001  & ~n20468 ;
  assign n20532 = n20484 & n20524 ;
  assign n20533 = ~n20487 & ~n20525 ;
  assign n20534 = ~n20532 & n20533 ;
  assign n20535 = n20468 & ~n20534 ;
  assign n20536 = ~n20531 & ~n20535 ;
  assign n20537 = \core_eu_ea_alu_ea_dec_piconst_DO_reg[1]/P0001  & ~n20468 ;
  assign n20538 = ~\core_c_dec_IR_reg[11]/NET0131  & n20508 ;
  assign n20540 = n20473 & n20538 ;
  assign n20539 = n20475 & ~n20538 ;
  assign n20541 = ~n20478 & ~n20539 ;
  assign n20542 = ~n20540 & n20541 ;
  assign n20543 = n20468 & ~n20542 ;
  assign n20544 = ~n20537 & ~n20543 ;
  assign n20545 = \core_eu_ea_alu_ea_dec_piconst_DO_reg[11]/P0001  & ~n20468 ;
  assign n20546 = \core_c_dec_IR_reg[7]/NET0131  & n20470 ;
  assign n20548 = n20473 & n20546 ;
  assign n20547 = n20475 & ~n20546 ;
  assign n20549 = ~n20478 & ~n20547 ;
  assign n20550 = ~n20548 & n20549 ;
  assign n20551 = n20468 & ~n20550 ;
  assign n20552 = ~n20545 & ~n20551 ;
  assign n20553 = \core_eu_ea_alu_ea_dec_piconst_DO_reg[10]/P0001  & ~n20468 ;
  assign n20554 = n20484 & n20546 ;
  assign n20555 = ~n20487 & ~n20547 ;
  assign n20556 = ~n20554 & n20555 ;
  assign n20557 = n20468 & ~n20556 ;
  assign n20558 = ~n20553 & ~n20557 ;
  assign n20559 = \core_eu_ea_alu_ea_dec_piconst_DO_reg[0]/P0001  & ~n20468 ;
  assign n20560 = n20484 & n20538 ;
  assign n20561 = ~n20487 & ~n20539 ;
  assign n20562 = ~n20560 & n20561 ;
  assign n20563 = n20468 & ~n20562 ;
  assign n20564 = ~n20559 & ~n20563 ;
  assign n20565 = ~n8460 & n20402 ;
  assign n20566 = ~\sport0_regs_AUTOreg_DO_reg[11]/NET0131  & ~n20402 ;
  assign n20567 = ~n20565 & ~n20566 ;
  assign n20568 = ~n7859 & n20402 ;
  assign n20569 = ~\sport0_regs_AUTOreg_DO_reg[10]/NET0131  & ~n20402 ;
  assign n20570 = ~n20568 & ~n20569 ;
  assign n20571 = ~\core_c_dec_DU_Eg_reg/P0001  & ~\core_c_dec_MpopLP_Eg_reg/P0001  ;
  assign n20572 = ~\core_c_psq_Eqend_Ed_reg/P0001  & n20571 ;
  assign n20573 = ~\core_c_psq_lpstk_ptr_reg[2]/NET0131  & n4849 ;
  assign n20574 = \core_c_dec_DU_Eg_reg/P0001  & ~n5950 ;
  assign n20575 = ~n20573 & n20574 ;
  assign n20576 = ~n20572 & n20575 ;
  assign n20577 = ~\core_c_dec_MpopLP_Eg_reg/P0001  & ~n4842 ;
  assign n20578 = ~n5950 & ~n20577 ;
  assign n20579 = ~\core_c_psq_lpstk_ptr_reg[2]/NET0131  & n20578 ;
  assign n20580 = ~n20572 & n20579 ;
  assign n20581 = ~n20576 & ~n20580 ;
  assign n20582 = ~n4847 & ~n4851 ;
  assign n20583 = n20574 & ~n20582 ;
  assign n20584 = ~n20575 & n20582 ;
  assign n20585 = ~n20583 & ~n20584 ;
  assign n20586 = ~n20581 & ~n20585 ;
  assign n20587 = \core_c_psq_lpstk_ptr_reg[1]/NET0131  & n20581 ;
  assign n20588 = ~n20586 & ~n20587 ;
  assign n20589 = \core_c_psq_lpstk_ptr_reg[0]/NET0131  & ~n20581 ;
  assign n20590 = ~\core_c_psq_lpstk_ptr_reg[0]/NET0131  & n20581 ;
  assign n20591 = ~n20589 & ~n20590 ;
  assign n20592 = \core_c_psq_Iact_E_reg[7]/NET0131  & ~n19477 ;
  assign n20593 = n19487 & n19489 ;
  assign n20594 = ~n20592 & ~n20593 ;
  assign n20595 = n4849 & n20576 ;
  assign n20596 = \core_c_psq_lpstk_ptr_reg[2]/NET0131  & ~n20595 ;
  assign n20597 = n4845 & ~n20572 ;
  assign n20598 = ~n20575 & n20597 ;
  assign n20599 = n20578 & n20598 ;
  assign n20600 = ~n20596 & ~n20599 ;
  assign n20601 = n6164 & ~n10638 ;
  assign n20602 = ~n13347 & ~n20601 ;
  assign n20603 = ~n6047 & n20602 ;
  assign n20604 = n11609 & ~n20603 ;
  assign n20605 = n6029 & ~n20604 ;
  assign n20606 = \core_c_dec_IR_reg[18]/NET0131  & ~\core_c_dec_IR_reg[19]/NET0131  ;
  assign n20607 = n6118 & n20606 ;
  assign n20608 = \core_c_dec_IR_reg[12]/NET0131  & n20607 ;
  assign n20609 = ~n4094 & ~n20608 ;
  assign n20610 = ~n20605 & n20609 ;
  assign n20611 = ~\core_c_psq_Taddr_Eb_reg[8]/P0001  & n4094 ;
  assign n20612 = ~n20610 & ~n20611 ;
  assign n20613 = n6164 & ~n11265 ;
  assign n20614 = ~n13328 & ~n20613 ;
  assign n20615 = ~n6047 & n20614 ;
  assign n20616 = n11540 & ~n20615 ;
  assign n20617 = n6029 & ~n20616 ;
  assign n20618 = \core_c_dec_IR_reg[11]/NET0131  & n20607 ;
  assign n20619 = ~n4094 & ~n20618 ;
  assign n20620 = ~n20617 & n20619 ;
  assign n20621 = ~\core_c_psq_Taddr_Eb_reg[7]/P0001  & n4094 ;
  assign n20622 = ~n20620 & ~n20621 ;
  assign n20623 = n6164 & ~n11525 ;
  assign n20624 = ~n13309 & ~n20623 ;
  assign n20625 = ~n6047 & n20624 ;
  assign n20626 = n10967 & ~n20625 ;
  assign n20627 = n6029 & ~n20626 ;
  assign n20628 = \core_c_dec_IR_reg[10]/NET0131  & n20607 ;
  assign n20629 = ~n4094 & ~n20628 ;
  assign n20630 = ~n20627 & n20629 ;
  assign n20631 = ~\core_c_psq_Taddr_Eb_reg[6]/P0001  & n4094 ;
  assign n20632 = ~n20630 & ~n20631 ;
  assign n20633 = n6164 & ~n10911 ;
  assign n20634 = ~n13290 & ~n20633 ;
  assign n20635 = ~n6047 & n20634 ;
  assign n20636 = n10356 & ~n20635 ;
  assign n20637 = n6029 & ~n20636 ;
  assign n20638 = \core_c_dec_IR_reg[9]/NET0131  & n20607 ;
  assign n20639 = ~n4094 & ~n20638 ;
  assign n20640 = ~n20637 & n20639 ;
  assign n20641 = ~\core_c_psq_Taddr_Eb_reg[5]/P0001  & n4094 ;
  assign n20642 = ~n20640 & ~n20641 ;
  assign n20643 = n6164 & ~n10069 ;
  assign n20644 = ~n13271 & ~n20643 ;
  assign n20645 = ~n6047 & n20644 ;
  assign n20646 = n9805 & ~n20645 ;
  assign n20647 = n6029 & ~n20646 ;
  assign n20648 = \core_c_dec_IR_reg[8]/NET0131  & n20607 ;
  assign n20649 = ~n4094 & ~n20648 ;
  assign n20650 = ~n20647 & n20649 ;
  assign n20651 = ~\core_c_psq_Taddr_Eb_reg[4]/P0001  & n4094 ;
  assign n20652 = ~n20650 & ~n20651 ;
  assign n20653 = ~n6047 & n13262 ;
  assign n20654 = n9666 & ~n20653 ;
  assign n20655 = n6029 & ~n20654 ;
  assign n20656 = \core_c_dec_IR_reg[7]/NET0131  & n20607 ;
  assign n20657 = ~n4094 & ~n20656 ;
  assign n20658 = ~n20655 & n20657 ;
  assign n20659 = ~\core_c_psq_Taddr_Eb_reg[3]/P0001  & n4094 ;
  assign n20660 = ~n20658 & ~n20659 ;
  assign n20661 = ~n6164 & ~n9625 ;
  assign n20662 = n6164 & n8715 ;
  assign n20663 = ~n20661 & ~n20662 ;
  assign n20664 = ~n6047 & ~n20663 ;
  assign n20665 = n9600 & ~n20664 ;
  assign n20666 = n6029 & ~n20665 ;
  assign n20667 = \core_c_dec_IR_reg[6]/NET0131  & n20607 ;
  assign n20668 = ~n4094 & ~n20667 ;
  assign n20669 = ~n20666 & n20668 ;
  assign n20670 = ~\core_c_psq_Taddr_Eb_reg[2]/P0001  & n4094 ;
  assign n20671 = ~n20669 & ~n20670 ;
  assign n20672 = ~n6164 & ~n9559 ;
  assign n20673 = n6164 & n9435 ;
  assign n20674 = ~n20672 & ~n20673 ;
  assign n20675 = ~n6047 & ~n20674 ;
  assign n20676 = n9528 & ~n20675 ;
  assign n20677 = n6029 & ~n20676 ;
  assign n20678 = \core_c_dec_IR_reg[5]/NET0131  & n20607 ;
  assign n20679 = ~n4094 & ~n20678 ;
  assign n20680 = ~n20677 & n20679 ;
  assign n20681 = ~\core_c_psq_Taddr_Eb_reg[1]/P0001  & n4094 ;
  assign n20682 = ~n20680 & ~n20681 ;
  assign n20683 = ~n6164 & ~n9497 ;
  assign n20684 = n6164 & n7340 ;
  assign n20685 = ~n20683 & ~n20684 ;
  assign n20686 = ~n6047 & ~n20685 ;
  assign n20687 = n9452 & ~n20686 ;
  assign n20688 = n6029 & ~n20687 ;
  assign n20689 = \core_c_dec_IR_reg[17]/NET0131  & n20607 ;
  assign n20690 = ~n4094 & ~n20689 ;
  assign n20691 = ~n20688 & n20690 ;
  assign n20692 = ~\core_c_psq_Taddr_Eb_reg[13]/P0001  & n4094 ;
  assign n20693 = ~n20691 & ~n20692 ;
  assign n20694 = ~n6164 & ~n8945 ;
  assign n20695 = n6164 & n9178 ;
  assign n20696 = ~n20694 & ~n20695 ;
  assign n20697 = ~n6047 & ~n20696 ;
  assign n20698 = n8845 & ~n20697 ;
  assign n20699 = n6029 & ~n20698 ;
  assign n20700 = \core_c_dec_IR_reg[16]/NET0131  & n20607 ;
  assign n20701 = ~n4094 & ~n20700 ;
  assign n20702 = ~n20699 & n20701 ;
  assign n20703 = ~\core_c_psq_Taddr_Eb_reg[12]/P0001  & n4094 ;
  assign n20704 = ~n20702 & ~n20703 ;
  assign n20705 = ~n6164 & ~n8813 ;
  assign n20706 = n6164 & n8460 ;
  assign n20707 = ~n20705 & ~n20706 ;
  assign n20708 = ~n6047 & ~n20707 ;
  assign n20709 = n8723 & ~n20708 ;
  assign n20710 = n6029 & ~n20709 ;
  assign n20711 = \core_c_dec_IR_reg[15]/NET0131  & n20607 ;
  assign n20712 = ~n4094 & ~n20711 ;
  assign n20713 = ~n20710 & n20712 ;
  assign n20714 = ~\core_c_psq_Taddr_Eb_reg[11]/P0001  & n4094 ;
  assign n20715 = ~n20713 & ~n20714 ;
  assign n20716 = n6164 & ~n7859 ;
  assign n20717 = ~n6164 & n8211 ;
  assign n20718 = ~n20716 & ~n20717 ;
  assign n20719 = ~n6047 & n20718 ;
  assign n20720 = n8121 & ~n20719 ;
  assign n20721 = n6029 & ~n20720 ;
  assign n20722 = \core_c_dec_IR_reg[14]/NET0131  & n20607 ;
  assign n20723 = ~n4094 & ~n20722 ;
  assign n20724 = ~n20721 & n20723 ;
  assign n20725 = ~\core_c_psq_Taddr_Eb_reg[10]/P0001  & n4094 ;
  assign n20726 = ~n20724 & ~n20725 ;
  assign n20727 = ~n6164 & ~n6911 ;
  assign n20728 = n6164 & n7607 ;
  assign n20729 = ~n20727 & ~n20728 ;
  assign n20730 = ~n6047 & ~n20729 ;
  assign n20731 = n6980 & ~n20730 ;
  assign n20732 = n6029 & ~n20731 ;
  assign n20733 = \core_c_dec_IR_reg[4]/NET0131  & n20607 ;
  assign n20734 = ~n4094 & ~n20733 ;
  assign n20735 = ~n20732 & n20734 ;
  assign n20736 = ~\core_c_psq_Taddr_Eb_reg[0]/P0001  & n4094 ;
  assign n20737 = ~n20735 & ~n20736 ;
  assign n20738 = \sice_ICYC_reg[8]/NET0131  & n18863 ;
  assign n20739 = \sice_ICYC_reg[9]/NET0131  & n20738 ;
  assign n20740 = \sice_ICYC_reg[10]/NET0131  & n20739 ;
  assign n20741 = \sice_ICYC_reg[11]/NET0131  & n20740 ;
  assign n20742 = \sice_ICYC_reg[12]/NET0131  & n20741 ;
  assign n20743 = \sice_ICYC_reg[13]/NET0131  & n20742 ;
  assign n20744 = \sice_ICYC_reg[14]/NET0131  & n20743 ;
  assign n20745 = \sice_ICYC_reg[15]/NET0131  & n20744 ;
  assign n20746 = \sice_ICYC_reg[16]/NET0131  & n20745 ;
  assign n20747 = \sice_ICYC_reg[17]/NET0131  & n20746 ;
  assign n20748 = \sice_ICYC_reg[18]/NET0131  & n20747 ;
  assign n20749 = \sice_ICYC_reg[19]/NET0131  & n20748 ;
  assign n20750 = \sice_ICYC_reg[20]/NET0131  & n20749 ;
  assign n20751 = ~\sice_ICYC_reg[21]/NET0131  & ~n20750 ;
  assign n20752 = \sice_ICYC_reg[21]/NET0131  & n20750 ;
  assign n20753 = ~n20751 & ~n20752 ;
  assign n20754 = n6164 & ~n10289 ;
  assign n20755 = ~n13366 & ~n20754 ;
  assign n20756 = ~n6047 & n20755 ;
  assign n20757 = n11668 & ~n20756 ;
  assign n20758 = n6029 & ~n20757 ;
  assign n20759 = \core_c_dec_IR_reg[13]/NET0131  & n20607 ;
  assign n20760 = ~n4094 & ~n20759 ;
  assign n20761 = ~n20758 & n20760 ;
  assign n20762 = ~\core_c_psq_Taddr_Eb_reg[9]/P0001  & n4094 ;
  assign n20763 = ~n20761 & ~n20762 ;
  assign n20766 = ~\bdma_BEAD_reg[0]/NET0131  & ~n13147 ;
  assign n20767 = n13751 & ~n20766 ;
  assign n20769 = \bdma_BEAD_reg[1]/NET0131  & n20767 ;
  assign n20764 = n13762 & n20070 ;
  assign n20765 = n7237 & n20764 ;
  assign n20768 = ~\bdma_BEAD_reg[1]/NET0131  & ~n20767 ;
  assign n20770 = ~n20765 & ~n20768 ;
  assign n20771 = ~n20769 & n20770 ;
  assign n20772 = n9435 & n20765 ;
  assign n20773 = ~n20771 & ~n20772 ;
  assign n20774 = ~n13147 & n13751 ;
  assign n20775 = \bdma_BEAD_reg[0]/NET0131  & ~n20774 ;
  assign n20776 = ~\bdma_BEAD_reg[0]/NET0131  & n20774 ;
  assign n20777 = ~n20775 & ~n20776 ;
  assign n20778 = ~n20765 & ~n20777 ;
  assign n20779 = n7607 & n20765 ;
  assign n20780 = ~n20778 & ~n20779 ;
  assign n20781 = \clkc_CLKOUT_reg/NET0131  & ~n19467 ;
  assign n20782 = ~\clkc_CLKOUT_reg/NET0131  & n19467 ;
  assign n20783 = ~n20781 & ~n20782 ;
  assign n20784 = ~\sice_ICYC_reg[22]/NET0131  & ~n20752 ;
  assign n20785 = \sice_ICYC_reg[22]/NET0131  & n20752 ;
  assign n20786 = ~n20784 & ~n20785 ;
  assign n20787 = n7513 & n18226 ;
  assign n20788 = ~\memc_MMR_web_reg/NET0131  & n20787 ;
  assign n20789 = ~n11265 & n20788 ;
  assign n20790 = ~\tm_tsr_reg_DO_reg[7]/NET0131  & ~n20788 ;
  assign n20791 = ~n20789 & ~n20790 ;
  assign n20792 = ~n11525 & n20788 ;
  assign n20793 = ~\tm_tsr_reg_DO_reg[6]/NET0131  & ~n20788 ;
  assign n20794 = ~n20792 & ~n20793 ;
  assign n20795 = ~n10911 & n20788 ;
  assign n20796 = ~\tm_tsr_reg_DO_reg[5]/NET0131  & ~n20788 ;
  assign n20797 = ~n20795 & ~n20796 ;
  assign n20798 = ~n8113 & n20788 ;
  assign n20799 = ~\tm_tsr_reg_DO_reg[3]/NET0131  & ~n20788 ;
  assign n20800 = ~n20798 & ~n20799 ;
  assign n20801 = ~n8715 & n20788 ;
  assign n20802 = ~\tm_tsr_reg_DO_reg[2]/NET0131  & ~n20788 ;
  assign n20803 = ~n20801 & ~n20802 ;
  assign n20804 = ~n10069 & n20788 ;
  assign n20805 = ~\tm_tsr_reg_DO_reg[4]/NET0131  & ~n20788 ;
  assign n20806 = ~n20804 & ~n20805 ;
  assign n20807 = ~n9435 & n20788 ;
  assign n20808 = ~\tm_tsr_reg_DO_reg[1]/NET0131  & ~n20788 ;
  assign n20809 = ~n20807 & ~n20808 ;
  assign n20810 = ~n7607 & n20788 ;
  assign n20811 = ~\tm_tsr_reg_DO_reg[0]/NET0131  & ~n20788 ;
  assign n20812 = ~n20810 & ~n20811 ;
  assign n20813 = ~n12743 & n20788 ;
  assign n20814 = ~\tm_tsr_reg_DO_reg[8]/NET0131  & ~n20788 ;
  assign n20815 = ~n20813 & ~n20814 ;
  assign n20816 = ~\memc_usysr_DO_reg[7]/NET0131  & n20455 ;
  assign n20817 = \idma_WRcnt_reg[0]/NET0131  & ~n20456 ;
  assign n20818 = ~n20455 & ~n20457 ;
  assign n20819 = ~n20817 & n20818 ;
  assign n20820 = ~n20816 & ~n20819 ;
  assign n20822 = ~\idma_DCTL_reg[14]/NET0131  & ~n20454 ;
  assign n20823 = ~\idma_PM_1st_reg/NET0131  & n20822 ;
  assign n20825 = \idma_RDcyc_reg/NET0131  & n20823 ;
  assign n20826 = ~\idma_RDcnt_reg[0]/NET0131  & n20825 ;
  assign n20827 = \idma_RDcnt_reg[1]/NET0131  & ~n20826 ;
  assign n20821 = ~\idma_RDCMD_d1_reg/P0001  & \idma_RDCMD_reg/P0001  ;
  assign n20824 = n20821 & n20823 ;
  assign n20828 = n20390 & n20825 ;
  assign n20829 = ~n20824 & ~n20828 ;
  assign n20830 = ~n20827 & n20829 ;
  assign n20831 = ~\memc_usysr_DO_reg[5]/NET0131  & n20824 ;
  assign n20832 = ~n20830 & ~n20831 ;
  assign n20833 = ~\memc_usysr_DO_reg[4]/NET0131  & n20824 ;
  assign n20834 = \idma_RDcnt_reg[0]/NET0131  & ~n20825 ;
  assign n20835 = ~n20824 & ~n20826 ;
  assign n20836 = ~n20834 & n20835 ;
  assign n20837 = ~n20833 & ~n20836 ;
  assign n20838 = \core_c_dec_updAR_E_reg/P0001  & n4118 ;
  assign n20839 = n18850 & n20377 ;
  assign n20840 = ~n20838 & ~n20839 ;
  assign n20841 = ~\sice_ICYC_reg[3]/NET0131  & ~n18857 ;
  assign n20842 = ~n18858 & ~n20841 ;
  assign n20843 = ~\sice_IIRC_reg[3]/NET0131  & ~n18866 ;
  assign n20844 = ~n18867 & ~n20843 ;
  assign n20845 = \clkc_oscntr_reg_DO_reg[0]/NET0131  & \clkc_oscntr_reg_DO_reg[1]/NET0131  ;
  assign n20846 = \clkc_oscntr_reg_DO_reg[2]/NET0131  & ~n20845 ;
  assign n20847 = \clkc_oscntr_reg_DO_reg[2]/NET0131  & \clkc_oscntr_reg_DO_reg[3]/NET0131  ;
  assign n20848 = ~\clkc_oscntr_reg_DO_reg[2]/NET0131  & ~\clkc_oscntr_reg_DO_reg[3]/NET0131  ;
  assign n20849 = ~n20847 & ~n20848 ;
  assign n20850 = ~n20846 & ~n20849 ;
  assign n20851 = n20846 & n20849 ;
  assign n20852 = ~n20850 & ~n20851 ;
  assign n20853 = \sice_IIRC_reg[8]/NET0131  & n18871 ;
  assign n20854 = \sice_IIRC_reg[9]/NET0131  & n20853 ;
  assign n20855 = \sice_IIRC_reg[10]/NET0131  & n20854 ;
  assign n20856 = \sice_IIRC_reg[11]/NET0131  & n20855 ;
  assign n20857 = \sice_IIRC_reg[12]/NET0131  & n20856 ;
  assign n20858 = \sice_IIRC_reg[13]/NET0131  & n20857 ;
  assign n20859 = \sice_IIRC_reg[14]/NET0131  & n20858 ;
  assign n20860 = ~\sice_IIRC_reg[14]/NET0131  & ~n20858 ;
  assign n20861 = ~n20859 & ~n20860 ;
  assign n20862 = ~\sice_ICYC_reg[14]/NET0131  & ~n20743 ;
  assign n20863 = ~n20744 & ~n20862 ;
  assign n20864 = \core_c_dec_updMF_E_reg/P0001  & n14666 ;
  assign n20865 = \core_eu_em_mac_em_reg_mfswe_DO_reg[9]/P0001  & ~n20864 ;
  assign n20866 = ~n19525 & n20864 ;
  assign n20867 = ~n20865 & ~n20866 ;
  assign n20876 = \sport0_regs_SCTLreg_DO_reg[4]/NET0131  & ~\sport0_rxctl_RX_reg[5]/P0001  ;
  assign n20877 = ~\sport0_regs_SCTLreg_DO_reg[4]/NET0131  & \sport0_rxctl_RX_reg[5]/P0001  ;
  assign n20878 = ~n20876 & ~n20877 ;
  assign n20879 = \sport0_rxctl_RX_reg[6]/P0001  & ~n20878 ;
  assign n20880 = ~\sport0_regs_SCTLreg_DO_reg[4]/NET0131  & ~n20879 ;
  assign n20881 = \sport0_rxctl_RX_reg[4]/P0001  & n20879 ;
  assign n20882 = \sport0_regs_SCTLreg_DO_reg[4]/NET0131  & ~n20881 ;
  assign n20886 = \sport0_regs_SCTLreg_DO_reg[4]/NET0131  & ~\sport0_rxctl_RX_reg[1]/P0001  ;
  assign n20887 = ~\sport0_regs_SCTLreg_DO_reg[4]/NET0131  & \sport0_rxctl_RX_reg[1]/P0001  ;
  assign n20888 = ~n20886 & ~n20887 ;
  assign n20889 = ~\sport0_rxctl_RX_reg[4]/P0001  & n20888 ;
  assign n20885 = ~\sport0_rxctl_RX_reg[2]/P0001  & \sport0_rxctl_RX_reg[4]/P0001  ;
  assign n20890 = ~n20878 & ~n20885 ;
  assign n20891 = ~n20889 & n20890 ;
  assign n20883 = \sport0_rxctl_RX_reg[0]/P0001  & \sport0_rxctl_RX_reg[4]/P0001  ;
  assign n20884 = n20878 & n20883 ;
  assign n20892 = \sport0_rxctl_RX_reg[6]/P0001  & ~n20884 ;
  assign n20893 = ~n20891 & n20892 ;
  assign n20894 = n20882 & ~n20893 ;
  assign n20897 = ~\sport0_rxctl_RX_reg[0]/P0001  & ~n20878 ;
  assign n20898 = ~\sport0_rxctl_RX_reg[4]/P0001  & ~n20897 ;
  assign n20895 = ~n20878 & ~n20888 ;
  assign n20896 = \sport0_rxctl_RX_reg[4]/P0001  & n20895 ;
  assign n20899 = \sport0_rxctl_RX_reg[6]/P0001  & ~n20896 ;
  assign n20900 = ~n20898 & n20899 ;
  assign n20901 = ~n20882 & ~n20900 ;
  assign n20902 = ~n20894 & ~n20901 ;
  assign n20903 = n20880 & ~n20902 ;
  assign n20904 = \sport0_rxctl_RX_reg[4]/P0001  & n20878 ;
  assign n20905 = n20888 & n20904 ;
  assign n20907 = \sport0_rxctl_RX_reg[0]/P0001  & n20878 ;
  assign n20906 = \sport0_rxctl_RX_reg[2]/P0001  & ~n20878 ;
  assign n20908 = ~\sport0_rxctl_RX_reg[4]/P0001  & ~n20906 ;
  assign n20909 = ~n20907 & n20908 ;
  assign n20910 = ~n20905 & ~n20909 ;
  assign n20911 = \sport0_rxctl_RX_reg[6]/P0001  & ~n20910 ;
  assign n20912 = \sport0_regs_SCTLreg_DO_reg[4]/NET0131  & ~\sport0_rxctl_RX_reg[3]/P0001  ;
  assign n20913 = ~\sport0_regs_SCTLreg_DO_reg[4]/NET0131  & \sport0_rxctl_RX_reg[3]/P0001  ;
  assign n20914 = ~n20912 & ~n20913 ;
  assign n20915 = \sport0_rxctl_RX_reg[6]/P0001  & ~n20914 ;
  assign n20916 = \sport0_rxctl_RX_reg[4]/P0001  & ~n20878 ;
  assign n20917 = ~n20915 & n20916 ;
  assign n20918 = ~n20911 & ~n20917 ;
  assign n20919 = n20882 & ~n20918 ;
  assign n20920 = ~n20882 & n20893 ;
  assign n20921 = ~n20919 & ~n20920 ;
  assign n20922 = n20903 & n20921 ;
  assign n20925 = n20878 & ~n20888 ;
  assign n20926 = ~n20878 & ~n20914 ;
  assign n20927 = \sport0_rxctl_RX_reg[6]/P0001  & n20926 ;
  assign n20928 = ~n20925 & ~n20927 ;
  assign n20929 = ~\sport0_rxctl_RX_reg[4]/P0001  & ~n20928 ;
  assign n20923 = ~n20878 & ~n20883 ;
  assign n20924 = ~\sport0_rxctl_RX_reg[6]/P0001  & ~n20923 ;
  assign n20930 = \sport0_rxctl_RX_reg[2]/P0001  & n20878 ;
  assign n20931 = \sport0_rxctl_RX_reg[4]/P0001  & n20930 ;
  assign n20932 = ~n20924 & ~n20931 ;
  assign n20933 = ~n20929 & n20932 ;
  assign n20934 = n20882 & ~n20933 ;
  assign n20935 = ~n20882 & n20918 ;
  assign n20936 = ~n20934 & ~n20935 ;
  assign n20937 = ~n20922 & n20936 ;
  assign n20940 = n20882 & n20900 ;
  assign n20941 = n20879 & ~n20883 ;
  assign n20942 = ~n20882 & n20941 ;
  assign n20943 = ~n20940 & ~n20942 ;
  assign n20938 = ~\sport0_regs_SCTLreg_DO_reg[4]/NET0131  & ~n20881 ;
  assign n20939 = n20879 & ~n20938 ;
  assign n20944 = ~n20902 & ~n20939 ;
  assign n20945 = n20943 & n20944 ;
  assign n20946 = n20921 & n20945 ;
  assign n20947 = ~n20936 & n20946 ;
  assign n20948 = ~\sport0_regs_SCTLreg_DO_reg[4]/NET0131  & n20947 ;
  assign n20949 = ~n20937 & ~n20948 ;
  assign n20950 = ~n20880 & n20902 ;
  assign n20951 = ~n20903 & ~n20950 ;
  assign n20952 = \sport0_rxctl_RX_reg[6]/P0001  & n20876 ;
  assign n20953 = ~n20938 & ~n20952 ;
  assign n20954 = n20943 & n20953 ;
  assign n20955 = n20951 & n20954 ;
  assign n20956 = n20921 & n20955 ;
  assign n20957 = n20949 & n20956 ;
  assign n20958 = ~\sport0_rxctl_RX_reg[7]/P0001  & ~n20957 ;
  assign n20959 = ~\sport0_rxctl_RX_reg[6]/P0001  & ~n20895 ;
  assign n20960 = n20878 & n20914 ;
  assign n20961 = \sport0_rxctl_RX_reg[4]/P0001  & ~n20960 ;
  assign n20962 = ~n20959 & n20961 ;
  assign n20963 = ~\sport0_rxctl_RX_reg[6]/P0001  & ~n20897 ;
  assign n20964 = ~n20930 & ~n20963 ;
  assign n20965 = ~\sport0_rxctl_RX_reg[4]/P0001  & ~n20964 ;
  assign n20966 = ~n20962 & ~n20965 ;
  assign n20967 = n20882 & n20966 ;
  assign n20968 = ~n20882 & n20933 ;
  assign n20969 = ~n20967 & ~n20968 ;
  assign n20970 = \sport0_rxctl_RX_reg[4]/P0001  & n20952 ;
  assign n20971 = ~n20969 & ~n20970 ;
  assign n20972 = n20947 & ~n20971 ;
  assign n20973 = ~n20947 & n20971 ;
  assign n20974 = ~\sport0_regs_SCTLreg_DO_reg[4]/NET0131  & ~n20973 ;
  assign n20975 = ~n20972 & n20974 ;
  assign n20976 = ~n20967 & ~n20975 ;
  assign n20978 = n20958 & ~n20976 ;
  assign n20875 = \sport0_regs_SCTLreg_DO_reg[5]/NET0131  & \sport0_rxctl_ldRX_cmp_reg/P0001  ;
  assign n20977 = ~n20958 & n20976 ;
  assign n20979 = n20875 & ~n20977 ;
  assign n20980 = ~n20978 & n20979 ;
  assign n20981 = ~\sport0_rxctl_ldRX_cmp_reg/P0001  & n10911 ;
  assign n20868 = \sport0_rxctl_a_sync1_reg/P0001  & ~\sport0_rxctl_a_sync2_reg/P0001  ;
  assign n20873 = ~\sport0_regs_SCTLreg_DO_reg[5]/NET0131  & \sport0_rxctl_ldRX_cmp_reg/P0001  ;
  assign n20874 = \sport0_rxctl_RX_reg[5]/P0001  & n20873 ;
  assign n20982 = ~n20868 & ~n20874 ;
  assign n20983 = ~n20981 & n20982 ;
  assign n20984 = ~n20980 & n20983 ;
  assign n20869 = \core_c_dec_MTRX0_E_reg/P0001  & n5951 ;
  assign n20870 = ~n20868 & ~n20869 ;
  assign n20871 = ~\sport0_rxctl_ldRX_cmp_reg/P0001  & n20870 ;
  assign n20872 = ~\sport0_rxctl_RXSHT_reg[5]/P0001  & n20868 ;
  assign n20985 = ~n20871 & ~n20872 ;
  assign n20986 = ~n20984 & n20985 ;
  assign n20987 = \sport0_rxctl_RX_reg[5]/P0001  & n20871 ;
  assign n20988 = ~n20986 & ~n20987 ;
  assign n20989 = ~\clkc_OUTcnt_reg[0]/NET0131  & ~n19466 ;
  assign n20990 = \core_c_dec_updMF_E_reg/P0001  & n13804 ;
  assign n20991 = \core_eu_em_mac_em_reg_mfrwe_DO_reg[9]/P0001  & ~n20990 ;
  assign n20992 = ~n19525 & n20990 ;
  assign n20993 = ~n20991 & ~n20992 ;
  assign n20994 = \core_c_dec_MTSR1_E_reg/P0001  & ~n18974 ;
  assign n21005 = n18139 & n18171 ;
  assign n21006 = n18043 & n18162 ;
  assign n21029 = ~n21005 & ~n21006 ;
  assign n21007 = n18046 & n18187 ;
  assign n21010 = n17945 & n17960 ;
  assign n21030 = ~n21007 & ~n21010 ;
  assign n21033 = n21029 & n21030 ;
  assign n21001 = ~n17922 & ~n18104 ;
  assign n21002 = n17930 & ~n18907 ;
  assign n21027 = ~n21001 & ~n21002 ;
  assign n21003 = ~n18091 & n18125 ;
  assign n21004 = ~n18912 & n19720 ;
  assign n21028 = ~n21003 & ~n21004 ;
  assign n21034 = n21027 & n21028 ;
  assign n21040 = n21033 & n21034 ;
  assign n20998 = ~n18069 & n19873 ;
  assign n20999 = n20085 & n20998 ;
  assign n21017 = n18111 & n18893 ;
  assign n21013 = n18070 & n18183 ;
  assign n21014 = ~n18127 & n18732 ;
  assign n21031 = ~n21013 & ~n21014 ;
  assign n21032 = ~n21017 & n21031 ;
  assign n21041 = n20999 & n21032 ;
  assign n21042 = n21040 & n21041 ;
  assign n21011 = n18115 & ~n18781 ;
  assign n21008 = ~n17933 & n20104 ;
  assign n21009 = n18758 & ~n18775 ;
  assign n21037 = ~n21008 & ~n21009 ;
  assign n21038 = ~n21011 & n21037 ;
  assign n21019 = \core_c_dec_IRE_reg[11]/NET0131  & ~n9280 ;
  assign n21020 = ~n18192 & ~n21019 ;
  assign n20995 = n18153 & ~n18189 ;
  assign n21012 = n18055 & n18172 ;
  assign n21021 = ~n20995 & ~n21012 ;
  assign n21024 = n21020 & n21021 ;
  assign n21025 = ~n18040 & n21024 ;
  assign n21000 = n18147 & n18745 ;
  assign n21018 = n17986 & ~n18167 ;
  assign n21015 = n18089 & n18128 ;
  assign n21016 = n18056 & n18112 ;
  assign n21022 = ~n21015 & ~n21016 ;
  assign n21023 = ~n21018 & n21022 ;
  assign n21026 = ~n21000 & n21023 ;
  assign n21035 = n21025 & n21026 ;
  assign n20996 = n17931 & ~n18912 ;
  assign n20997 = ~n18175 & n20996 ;
  assign n21036 = n20108 & ~n20997 ;
  assign n21039 = n21035 & n21036 ;
  assign n21043 = n21038 & n21039 ;
  assign n21044 = n21042 & n21043 ;
  assign n21045 = n20090 & n21044 ;
  assign n21046 = n19793 & n21045 ;
  assign n21047 = ~\core_c_dec_MTSR1_E_reg/P0001  & n21046 ;
  assign n21048 = ~n20994 & ~n21047 ;
  assign n21049 = n18717 & ~n21048 ;
  assign n21050 = ~\core_eu_es_sht_es_reg_sr1swe_DO_reg[1]/P0001  & ~n18717 ;
  assign n21051 = ~n21049 & ~n21050 ;
  assign n21052 = ~\clkc_OUTcnt_reg[5]/NET0131  & ~n19471 ;
  assign n21053 = ~n19472 & ~n21052 ;
  assign n21054 = ~n19467 & n21053 ;
  assign n21055 = n17833 & ~n21048 ;
  assign n21056 = ~\core_eu_es_sht_es_reg_sr1rwe_DO_reg[1]/P0001  & ~n17833 ;
  assign n21057 = ~n21055 & ~n21056 ;
  assign n21058 = ~\clkc_OUTcnt_reg[2]/NET0131  & ~n19468 ;
  assign n21059 = ~n19469 & ~n21058 ;
  assign n21060 = ~n19467 & n21059 ;
  assign n21063 = n18271 & ~n20259 ;
  assign n21062 = ~\core_eu_em_mac_em_reg_mr0swe_DO_reg[5]/P0001  & ~n18271 ;
  assign n21064 = n18273 & ~n21062 ;
  assign n21065 = ~n21063 & n21064 ;
  assign n21061 = \core_eu_em_mac_em_reg_mr0swe_DO_reg[5]/P0001  & ~n18266 ;
  assign n21066 = ~n18270 & ~n21061 ;
  assign n21067 = ~n21065 & n21066 ;
  assign n21068 = ~n18262 & ~n21067 ;
  assign n21069 = n18262 & ~n19628 ;
  assign n21070 = ~n21068 & ~n21069 ;
  assign n21071 = n14752 & n19628 ;
  assign n21072 = n18328 & n20259 ;
  assign n21073 = \core_eu_em_mac_em_reg_mr0rwe_DO_reg[5]/P0001  & ~n18330 ;
  assign n21074 = n18334 & ~n21073 ;
  assign n21075 = ~n21072 & n21074 ;
  assign n21076 = ~n21071 & ~n21075 ;
  assign n21077 = \core_c_dec_MTSR1_E_reg/P0001  & ~n17814 ;
  assign n21079 = ~n18034 & ~n18192 ;
  assign n21080 = ~n18040 & n21079 ;
  assign n21081 = n18145 & n21080 ;
  assign n21082 = ~n20112 & n21081 ;
  assign n21083 = n19790 & n21082 ;
  assign n21084 = n19793 & n21083 ;
  assign n21091 = n18147 & n18162 ;
  assign n21092 = n18766 & ~n18907 ;
  assign n21111 = ~n21091 & ~n21092 ;
  assign n21095 = ~n18912 & n20308 ;
  assign n21102 = ~n18108 & n18752 ;
  assign n21112 = ~n21095 & ~n21102 ;
  assign n21113 = n21111 & n21112 ;
  assign n21087 = ~n18091 & ~n20096 ;
  assign n21088 = n18071 & n18171 ;
  assign n21109 = ~n21087 & ~n21088 ;
  assign n21089 = n17980 & n18111 ;
  assign n21090 = ~n17922 & ~n18743 ;
  assign n21110 = ~n21089 & ~n21090 ;
  assign n21114 = n21109 & n21110 ;
  assign n21120 = n21113 & n21114 ;
  assign n21121 = n20999 & n21120 ;
  assign n21099 = ~n17924 & n20104 ;
  assign n21096 = n18187 & ~n19804 ;
  assign n21098 = n18115 & ~n19818 ;
  assign n21117 = ~n21096 & ~n21098 ;
  assign n21118 = ~n21099 & n21117 ;
  assign n21103 = ~n18182 & n18719 ;
  assign n21078 = n18171 & n18774 ;
  assign n21097 = n17965 & n18072 ;
  assign n21106 = ~n21078 & ~n21097 ;
  assign n21107 = ~n21103 & n21106 ;
  assign n21086 = n18046 & n18183 ;
  assign n21101 = n17986 & n18722 ;
  assign n21093 = n18056 & n18905 ;
  assign n21100 = \core_c_dec_IRE_reg[11]/NET0131  & ~n8497 ;
  assign n21104 = ~n21093 & ~n21100 ;
  assign n21105 = ~n21101 & n21104 ;
  assign n21108 = ~n21086 & n21105 ;
  assign n21115 = n21107 & n21108 ;
  assign n21085 = n18758 & ~n19857 ;
  assign n21094 = n18748 & ~n18895 ;
  assign n21116 = ~n21085 & ~n21094 ;
  assign n21119 = n21115 & n21116 ;
  assign n21122 = n21118 & n21119 ;
  assign n21123 = n21121 & n21122 ;
  assign n21124 = n21084 & n21123 ;
  assign n21125 = ~\core_c_dec_MTSR1_E_reg/P0001  & n21124 ;
  assign n21126 = ~n21077 & ~n21125 ;
  assign n21127 = n18717 & ~n21126 ;
  assign n21128 = ~\core_eu_es_sht_es_reg_sr1swe_DO_reg[2]/P0001  & ~n18717 ;
  assign n21129 = ~n21127 & ~n21128 ;
  assign n21130 = n17833 & ~n21126 ;
  assign n21131 = ~\core_eu_es_sht_es_reg_sr1rwe_DO_reg[2]/P0001  & ~n17833 ;
  assign n21132 = ~n21130 & ~n21131 ;
  assign n21133 = \core_c_dec_Call_Ed_reg/P0001  & ~n4184 ;
  assign n21134 = ~\core_c_dec_DU_Eg_reg/P0001  & ~\core_c_dec_MTtoppcs_Eg_reg/P0001  ;
  assign n21135 = ~n21133 & n21134 ;
  assign n21136 = ~n5950 & ~n21135 ;
  assign n21137 = ~n18217 & ~n21136 ;
  assign n21138 = ~\core_c_psq_pcstk_ptr_reg[4]/NET0131  & n4215 ;
  assign n21139 = ~n21137 & n21138 ;
  assign n21140 = ~\core_c_psq_SSTAT_reg[1]/NET0131  & ~n21139 ;
  assign n21141 = \core_c_dec_MTSR0_E_reg/P0001  & ~n17814 ;
  assign n21145 = ~n18110 & ~n18987 ;
  assign n21146 = ~n18909 & ~n19864 ;
  assign n21148 = ~n18079 & ~n18915 ;
  assign n21161 = ~n21146 & ~n21148 ;
  assign n21150 = n17991 & n18748 ;
  assign n21152 = n18752 & ~n18912 ;
  assign n21162 = ~n21150 & ~n21152 ;
  assign n21163 = n21161 & n21162 ;
  assign n21143 = ~n18082 & n18766 ;
  assign n21151 = \core_c_dec_IRE_reg[11]/NET0131  & ~n8493 ;
  assign n21160 = ~n21143 & ~n21151 ;
  assign n21164 = n18019 & n21160 ;
  assign n21170 = n21163 & n21164 ;
  assign n21171 = ~n21145 & n21170 ;
  assign n21155 = n18745 & ~n18914 ;
  assign n21156 = n18740 & ~n18918 ;
  assign n21157 = ~n21155 & ~n21156 ;
  assign n21158 = ~n18026 & n21157 ;
  assign n21159 = ~n17931 & ~n21158 ;
  assign n21154 = n18088 & ~n18983 ;
  assign n21149 = ~n18123 & n19808 ;
  assign n21153 = ~n17924 & n18083 ;
  assign n21167 = ~n21149 & ~n21153 ;
  assign n21168 = ~n21154 & n21167 ;
  assign n21142 = n18187 & ~n18898 ;
  assign n21165 = n18903 & ~n21142 ;
  assign n21144 = ~n18098 & n19785 ;
  assign n21147 = ~n17998 & n18162 ;
  assign n21166 = ~n21144 & ~n21147 ;
  assign n21169 = n21165 & n21166 ;
  assign n21172 = n21168 & n21169 ;
  assign n21173 = ~n21159 & n21172 ;
  assign n21174 = n21171 & n21173 ;
  assign n21175 = ~\core_c_dec_MTSR0_E_reg/P0001  & n21174 ;
  assign n21176 = ~n21141 & ~n21175 ;
  assign n21177 = n18886 & ~n21176 ;
  assign n21178 = ~\core_eu_es_sht_es_reg_sr0swe_DO_reg[2]/P0001  & ~n18886 ;
  assign n21179 = ~n21177 & ~n21178 ;
  assign n21180 = \core_c_dec_MTSR0_E_reg/P0001  & ~n20150 ;
  assign n21184 = n18740 & ~n19804 ;
  assign n21185 = n18099 & ~n18149 ;
  assign n21219 = ~n21184 & ~n21185 ;
  assign n21201 = n18183 & ~n18781 ;
  assign n21202 = ~n17924 & n19785 ;
  assign n21220 = ~n21201 & ~n21202 ;
  assign n21221 = n21219 & n21220 ;
  assign n21195 = n17952 & n19862 ;
  assign n21197 = n17952 & n19863 ;
  assign n21207 = ~n21195 & ~n21197 ;
  assign n21198 = n18039 & n18766 ;
  assign n21199 = n17965 & n18067 ;
  assign n21208 = ~n21198 & ~n21199 ;
  assign n21209 = n21207 & n21208 ;
  assign n21196 = n18191 & n18766 ;
  assign n21191 = n18055 & n18722 ;
  assign n21194 = n18153 & ~n20096 ;
  assign n21204 = ~n21191 & ~n21194 ;
  assign n21205 = ~n21196 & n21204 ;
  assign n21182 = n18001 & ~n19864 ;
  assign n21188 = \core_c_dec_IRE_reg[11]/NET0131  & ~n11846 ;
  assign n21203 = ~n21182 & ~n21188 ;
  assign n21206 = ~n19811 & n21203 ;
  assign n21210 = n21205 & n21206 ;
  assign n21217 = n21209 & n21210 ;
  assign n21181 = n18187 & ~n19818 ;
  assign n21183 = n18758 & ~n18895 ;
  assign n21218 = ~n21181 & ~n21183 ;
  assign n21222 = n21217 & n21218 ;
  assign n21190 = ~n18914 & n20308 ;
  assign n21192 = ~n18091 & n18752 ;
  assign n21213 = ~n21190 & ~n21192 ;
  assign n21193 = n18070 & n18745 ;
  assign n21200 = n18071 & n18162 ;
  assign n21214 = ~n21193 & ~n21200 ;
  assign n21215 = n21213 & n21214 ;
  assign n21186 = n18905 & ~n18912 ;
  assign n21211 = n17978 & ~n21186 ;
  assign n21187 = n18749 & ~n18912 ;
  assign n21189 = n18046 & n18124 ;
  assign n21212 = ~n21187 & ~n21189 ;
  assign n21216 = n21211 & n21212 ;
  assign n21223 = n21215 & n21216 ;
  assign n21224 = n21222 & n21223 ;
  assign n21225 = n21221 & n21224 ;
  assign n21226 = n19794 & n21225 ;
  assign n21227 = ~\core_c_dec_MTSR0_E_reg/P0001  & n21226 ;
  assign n21228 = ~n21180 & ~n21227 ;
  assign n21229 = n18886 & ~n21228 ;
  assign n21230 = ~\core_eu_es_sht_es_reg_sr0swe_DO_reg[14]/P0001  & ~n18886 ;
  assign n21231 = ~n21229 & ~n21230 ;
  assign n21232 = n19034 & ~n21176 ;
  assign n21233 = ~\core_eu_es_sht_es_reg_sr0rwe_DO_reg[2]/P0001  & ~n19034 ;
  assign n21234 = ~n21232 & ~n21233 ;
  assign n21235 = n19034 & ~n21228 ;
  assign n21236 = ~\core_eu_es_sht_es_reg_sr0rwe_DO_reg[14]/P0001  & ~n19034 ;
  assign n21237 = ~n21235 & ~n21236 ;
  assign n21238 = \core_c_psq_PCS_reg[14]/NET0131  & \emc_eRDY_reg/NET0131  ;
  assign n21239 = \core_c_psq_PCS_reg[1]/NET0131  & n4068 ;
  assign n21240 = n4105 & n21239 ;
  assign n21241 = ~n21238 & ~n21240 ;
  assign n21242 = n4094 & n21241 ;
  assign n21244 = ~n5046 & ~n21242 ;
  assign n21243 = ~\core_c_psq_Eqend_D_reg/P0001  & n21242 ;
  assign n21245 = n4116 & ~n21243 ;
  assign n21246 = ~n21244 & n21245 ;
  assign n21247 = \core_c_dec_MpopLP_Eg_reg/P0001  & n4117 ;
  assign n21248 = \core_c_dec_IR_reg[16]/NET0131  & \core_c_dec_IR_reg[17]/NET0131  ;
  assign n21249 = n6027 & n6116 ;
  assign n21250 = n21248 & n21249 ;
  assign n21251 = n11742 & n21250 ;
  assign n21252 = \core_c_dec_IR_reg[3]/NET0131  & n21251 ;
  assign n21253 = ~n21247 & ~n21252 ;
  assign n21254 = n4116 & ~n21253 ;
  assign n21255 = \core_c_dec_Call_Ed_reg/P0001  & n4117 ;
  assign n21256 = ~n6029 & ~n20607 ;
  assign n21257 = n11742 & ~n21256 ;
  assign n21258 = ~\core_c_dec_IR_reg[4]/NET0131  & ~n20607 ;
  assign n21259 = n21257 & ~n21258 ;
  assign n21260 = ~n21255 & ~n21259 ;
  assign n21261 = n4116 & ~n21260 ;
  assign n21262 = \core_c_dec_ALUop_E_reg/P0001  & n4117 ;
  assign n21263 = ~n20377 & ~n21262 ;
  assign n21264 = n4116 & ~n21263 ;
  assign n21265 = ~\bdma_BWcnt_reg[3]/NET0131  & ~n20039 ;
  assign n21266 = ~n20040 & ~n21265 ;
  assign n21267 = ~n13750 & n21266 ;
  assign n21268 = n13762 & n20400 ;
  assign n21270 = ~n10069 & n21268 ;
  assign n21271 = ~n10911 & ~n11265 ;
  assign n21272 = ~n11525 & n21271 ;
  assign n21273 = n21270 & n21272 ;
  assign n21269 = n11265 & n21268 ;
  assign n21274 = \bdma_BCTL_reg[7]/NET0131  & ~n21268 ;
  assign n21275 = ~n21269 & ~n21274 ;
  assign n21276 = ~n21273 & n21275 ;
  assign n21277 = n11525 & n21268 ;
  assign n21278 = \bdma_BCTL_reg[6]/NET0131  & ~n21268 ;
  assign n21279 = ~n21277 & ~n21278 ;
  assign n21280 = ~n21273 & n21279 ;
  assign n21281 = n10911 & n21268 ;
  assign n21282 = \bdma_BCTL_reg[5]/NET0131  & ~n21268 ;
  assign n21283 = ~n21281 & ~n21282 ;
  assign n21284 = ~n21273 & n21283 ;
  assign n21285 = ~\bdma_BCTL_reg[4]/NET0131  & ~n21268 ;
  assign n21286 = ~n21270 & ~n21285 ;
  assign n21287 = ~n21273 & ~n21286 ;
  assign n21288 = ~\clkc_OUTcnt_reg[0]/NET0131  & ~\clkc_OUTcnt_reg[1]/NET0131  ;
  assign n21289 = ~n19468 & ~n21288 ;
  assign n21290 = ~n19467 & n21289 ;
  assign n21291 = n7270 & n13762 ;
  assign n21292 = \pio_PIO_RES_OUT_reg[8]/P0001  & ~\pio_PIO_RES_reg[8]/NET0131  ;
  assign n21293 = ~\pio_PIO_RES_OUT_reg[8]/P0001  & \pio_PIO_RES_reg[8]/NET0131  ;
  assign n21294 = ~n21292 & ~n21293 ;
  assign n21295 = ~\PIO_oe[8]_pad  & \pio_pmask_reg_DO_reg[8]/NET0131  ;
  assign n21296 = ~n21294 & n21295 ;
  assign n21297 = ~\pio_PINT_reg[8]/NET0131  & ~n21296 ;
  assign n21298 = ~n21291 & n21297 ;
  assign n21299 = ~n9178 & n21291 ;
  assign n21300 = ~n21298 & ~n21299 ;
  assign n21301 = ~\tm_WR_TSR_KEEP_TO_TMCLK_p_reg/NET0131  & ~\tm_WR_TSR_p_reg/P0001  ;
  assign n21302 = ~\emc_RWcnt_reg[3]/P0001  & ~n20216 ;
  assign n21303 = ~n20217 & ~n21302 ;
  assign n21304 = n20212 & n21303 ;
  assign n21305 = ~\emc_RWcnt_reg[2]/P0001  & ~n20215 ;
  assign n21306 = ~n20216 & ~n21305 ;
  assign n21307 = n20212 & n21306 ;
  assign n21308 = ~\emc_RWcnt_reg[1]/P0001  & ~n20214 ;
  assign n21309 = ~n20215 & ~n21308 ;
  assign n21310 = n20212 & n21309 ;
  assign n21311 = ~\emc_RWcnt_reg[0]/P0001  & n20213 ;
  assign n21312 = ~n20214 & ~n21311 ;
  assign n21313 = n20212 & n21312 ;
  assign n21314 = \core_c_dec_MACop_E_reg/P0001  & n19203 ;
  assign n21315 = n19202 & ~n21314 ;
  assign n21316 = ~\sport0_txctl_ldTX_cmp_reg/P0001  & ~n18519 ;
  assign n21317 = n10289 & n21316 ;
  assign n21318 = ~\sport0_txctl_ldTX_cmp_reg/P0001  & n18519 ;
  assign n21319 = \sport0_txctl_TX_reg[9]/P0001  & n21318 ;
  assign n21320 = ~\sport0_txctl_TX_reg[15]/P0001  & \sport0_txctl_ldTX_cmp_reg/P0001  ;
  assign n21321 = ~n21319 & ~n21320 ;
  assign n21322 = ~n21317 & n21321 ;
  assign n21323 = n10638 & n21316 ;
  assign n21324 = \sport0_txctl_TX_reg[8]/P0001  & n21318 ;
  assign n21325 = ~n21320 & ~n21324 ;
  assign n21326 = ~n21323 & n21325 ;
  assign n21327 = n11265 & n21316 ;
  assign n21328 = \sport0_txctl_TX_reg[7]/P0001  & n21318 ;
  assign n21329 = ~n21320 & ~n21328 ;
  assign n21330 = ~n21327 & n21329 ;
  assign n21331 = \pio_PIO_RES_OUT_reg[9]/P0001  & ~\pio_PIO_RES_reg[9]/NET0131  ;
  assign n21332 = ~\pio_PIO_RES_OUT_reg[9]/P0001  & \pio_PIO_RES_reg[9]/NET0131  ;
  assign n21333 = ~n21331 & ~n21332 ;
  assign n21334 = ~\PIO_oe[9]_pad  & \pio_pmask_reg_DO_reg[9]/NET0131  ;
  assign n21335 = ~n21333 & n21334 ;
  assign n21336 = ~\pio_PINT_reg[9]/NET0131  & ~n21335 ;
  assign n21337 = ~n21291 & n21336 ;
  assign n21338 = ~n7340 & n21291 ;
  assign n21339 = ~n21337 & ~n21338 ;
  assign n21341 = n12743 & n21316 ;
  assign n21340 = \sport0_txctl_TX_reg[15]/P0001  & n21318 ;
  assign n21342 = ~n21320 & ~n21340 ;
  assign n21343 = ~n21341 & n21342 ;
  assign n21344 = n7340 & n21316 ;
  assign n21345 = \sport0_txctl_TX_reg[13]/P0001  & n21318 ;
  assign n21346 = ~n21320 & ~n21345 ;
  assign n21347 = ~n21344 & n21346 ;
  assign n21348 = n12688 & n21316 ;
  assign n21349 = \sport0_txctl_TX_reg[14]/P0001  & n21318 ;
  assign n21350 = ~n21320 & ~n21349 ;
  assign n21351 = ~n21348 & n21350 ;
  assign n21352 = n9178 & n21316 ;
  assign n21353 = \sport0_txctl_TX_reg[12]/P0001  & n21318 ;
  assign n21354 = ~n21320 & ~n21353 ;
  assign n21355 = ~n21352 & n21354 ;
  assign n21356 = n8460 & n21316 ;
  assign n21357 = \sport0_txctl_TX_reg[11]/P0001  & n21318 ;
  assign n21358 = ~n21320 & ~n21357 ;
  assign n21359 = ~n21356 & n21358 ;
  assign n21360 = n7859 & n21316 ;
  assign n21361 = \sport0_txctl_TX_reg[10]/P0001  & n21318 ;
  assign n21362 = ~n21320 & ~n21361 ;
  assign n21363 = ~n21360 & n21362 ;
  assign n21364 = \core_eu_em_mac_em_reg_mfswe_DO_reg[0]/P0001  & ~n20864 ;
  assign n21365 = n19692 & n20864 ;
  assign n21366 = ~n21364 & ~n21365 ;
  assign n21367 = ~\sport0_regs_SCTLreg_DO_reg[5]/NET0131  & ~n20870 ;
  assign n21368 = ~n20875 & ~n21367 ;
  assign n21369 = \sport0_cfg_SP_ENg_reg/NET0131  & \sport0_regs_AUTOreg_DO_reg[0]/NET0131  ;
  assign n21370 = ~n21368 & n21369 ;
  assign n21371 = ~\sport0_rxctl_RSreq_reg/NET0131  & ~n21370 ;
  assign n21372 = \core_eu_em_mac_em_reg_mfrwe_DO_reg[0]/P0001  & ~n20990 ;
  assign n21373 = n19692 & n20990 ;
  assign n21374 = ~n21372 & ~n21373 ;
  assign n21375 = ~\IRFS1_pad  & \T_RFS1_pad  ;
  assign n21376 = \IRFS1_pad  & ~n13618 ;
  assign n21377 = ~n21375 & ~n21376 ;
  assign n21378 = ~\sport1_regs_SCTLreg_DO_reg[6]/NET0131  & n21377 ;
  assign n21379 = \sport1_regs_SCTLreg_DO_reg[6]/NET0131  & ~n21377 ;
  assign n21380 = ~n21378 & ~n21379 ;
  assign n21381 = ~\sport1_cfg_RFSgi_d_reg/NET0131  & \sport1_cfg_SP_ENg_reg/NET0131  ;
  assign n21382 = n21380 & n21381 ;
  assign n21383 = ~\IRFS0_pad  & \T_RFS0_pad  ;
  assign n21384 = \IRFS0_pad  & ~n13613 ;
  assign n21385 = ~n21383 & ~n21384 ;
  assign n21386 = ~\sport0_regs_SCTLreg_DO_reg[6]/NET0131  & n21385 ;
  assign n21387 = \sport0_regs_SCTLreg_DO_reg[6]/NET0131  & ~n21385 ;
  assign n21388 = ~n21386 & ~n21387 ;
  assign n21389 = ~\sport0_cfg_RFSgi_d_reg/NET0131  & \sport0_cfg_SP_ENg_reg/NET0131  ;
  assign n21390 = n21388 & n21389 ;
  assign n21391 = \core_c_psq_Iact_E_reg[9]/NET0131  & ~n4116 ;
  assign n21392 = ~\core_c_psq_IFC_reg[7]/NET0131  & ~n21391 ;
  assign n21393 = \core_c_psq_ICNTL_reg_DO_reg[2]/NET0131  & ~n21392 ;
  assign n21394 = \core_c_psq_ICNTL_reg_DO_reg[2]/NET0131  & \core_c_psq_T_IRQ2_s1_reg/P0001  ;
  assign n21395 = \core_c_psq_irq2_de_OUT_reg/P0001  & ~n21394 ;
  assign n21396 = ~\core_c_psq_IFC_reg[15]/NET0131  & ~\core_c_psq_Iflag_reg[9]/NET0131  ;
  assign n21397 = \core_c_psq_ICNTL_reg_DO_reg[2]/NET0131  & ~n21396 ;
  assign n21398 = ~n21395 & ~n21397 ;
  assign n21399 = ~n21393 & ~n21398 ;
  assign n21400 = ~\core_c_psq_ICNTL_reg_DO_reg[1]/NET0131  & \core_c_psq_irq1_de_OUT_reg/P0001  ;
  assign n21405 = \core_c_psq_Iact_E_reg[2]/NET0131  & ~n4116 ;
  assign n21406 = ~\core_c_psq_IFC_reg[2]/NET0131  & ~n21405 ;
  assign n21401 = ~\core_c_psq_T_IRQ1_s1_reg/P0001  & \core_c_psq_irq1_de_OUT_reg/P0001  ;
  assign n21402 = ~\core_c_psq_IFC_reg[10]/NET0131  & ~n21401 ;
  assign n21403 = ~\memc_usysr_DO_reg[11]/NET0131  & ~n21402 ;
  assign n21404 = ~\core_c_psq_Iflag_reg[12]/NET0131  & ~n21403 ;
  assign n21407 = \core_c_psq_ICNTL_reg_DO_reg[1]/NET0131  & ~n21404 ;
  assign n21408 = n21406 & n21407 ;
  assign n21409 = ~n21400 & ~n21408 ;
  assign n21410 = ~\core_c_psq_ICNTL_reg_DO_reg[0]/NET0131  & \core_c_psq_irq0_de_OUT_reg/P0001  ;
  assign n21415 = \core_c_psq_Iact_E_reg[1]/NET0131  & ~n4116 ;
  assign n21416 = ~\core_c_psq_IFC_reg[1]/NET0131  & ~n21415 ;
  assign n21411 = ~\core_c_psq_T_IRQ0_s1_reg/P0001  & \core_c_psq_irq0_de_OUT_reg/P0001  ;
  assign n21412 = ~\core_c_psq_IFC_reg[9]/NET0131  & ~n21411 ;
  assign n21413 = ~\memc_usysr_DO_reg[11]/NET0131  & ~n21412 ;
  assign n21414 = ~\core_c_psq_Iflag_reg[11]/NET0131  & ~n21413 ;
  assign n21417 = \core_c_psq_ICNTL_reg_DO_reg[0]/NET0131  & ~n21414 ;
  assign n21418 = n21416 & n21417 ;
  assign n21419 = ~n21410 & ~n21418 ;
  assign n21420 = \core_c_dec_updSR_E_reg/P0001  & n4118 ;
  assign n21421 = n4116 & ~n4117 ;
  assign n21422 = \core_c_dec_IR_reg[13]/NET0131  & \core_c_dec_IR_reg[14]/NET0131  ;
  assign n21423 = ~n19530 & ~n21422 ;
  assign n21424 = n21421 & n21423 ;
  assign n21425 = ~n21420 & ~n21424 ;
  assign n21427 = n6115 & n19698 ;
  assign n21428 = ~\core_c_psq_PCS_reg[3]/NET0131  & n21427 ;
  assign n21429 = n11742 & n21428 ;
  assign n21426 = \core_c_dec_Nseq_Ed_reg/P0001  & n4117 ;
  assign n21430 = ~n21257 & ~n21426 ;
  assign n21431 = ~n21429 & n21430 ;
  assign n21432 = n4116 & ~n21431 ;
  assign n21434 = ~\core_c_dec_IR_reg[4]/NET0131  & n21429 ;
  assign n21433 = \core_c_dec_Nrti_Ed_reg/P0001  & n4117 ;
  assign n21435 = ~n21257 & ~n21433 ;
  assign n21436 = ~n21434 & n21435 ;
  assign n21437 = n4116 & ~n21436 ;
  assign n21438 = \pio_PIO_RES_OUT_reg[5]/P0001  & ~\pio_PIO_RES_reg[5]/NET0131  ;
  assign n21439 = ~\pio_PIO_RES_OUT_reg[5]/P0001  & \pio_PIO_RES_reg[5]/NET0131  ;
  assign n21440 = ~n21438 & ~n21439 ;
  assign n21441 = ~\PIO_oe[5]_pad  & \pio_pmask_reg_DO_reg[5]/NET0131  ;
  assign n21442 = ~n21440 & n21441 ;
  assign n21443 = ~\pio_PINT_reg[5]/NET0131  & ~n21442 ;
  assign n21444 = ~n21291 & n21443 ;
  assign n21445 = ~n10911 & n21291 ;
  assign n21446 = ~n21444 & ~n21445 ;
  assign n21447 = \pio_PIO_RES_OUT_reg[4]/P0001  & ~\pio_PIO_RES_reg[4]/NET0131  ;
  assign n21448 = ~\pio_PIO_RES_OUT_reg[4]/P0001  & \pio_PIO_RES_reg[4]/NET0131  ;
  assign n21449 = ~n21447 & ~n21448 ;
  assign n21450 = ~\PIO_oe[4]_pad  & \pio_pmask_reg_DO_reg[4]/NET0131  ;
  assign n21451 = ~n21449 & n21450 ;
  assign n21452 = ~\pio_PINT_reg[4]/NET0131  & ~n21451 ;
  assign n21453 = ~n21291 & n21452 ;
  assign n21454 = ~n10069 & n21291 ;
  assign n21455 = ~n21453 & ~n21454 ;
  assign n21456 = \pio_PIO_RES_OUT_reg[11]/P0001  & ~\pio_PIO_RES_reg[11]/NET0131  ;
  assign n21457 = ~\pio_PIO_RES_OUT_reg[11]/P0001  & \pio_PIO_RES_reg[11]/NET0131  ;
  assign n21458 = ~n21456 & ~n21457 ;
  assign n21459 = ~\PIO_oe[11]_pad  & \pio_pmask_reg_DO_reg[11]/NET0131  ;
  assign n21460 = ~n21458 & n21459 ;
  assign n21461 = ~\pio_PINT_reg[11]/NET0131  & ~n21460 ;
  assign n21462 = ~n21291 & n21461 ;
  assign n21463 = ~n12743 & n21291 ;
  assign n21464 = ~n21462 & ~n21463 ;
  assign n21465 = \pio_PIO_RES_OUT_reg[2]/P0001  & ~\pio_PIO_RES_reg[2]/NET0131  ;
  assign n21466 = ~\pio_PIO_RES_OUT_reg[2]/P0001  & \pio_PIO_RES_reg[2]/NET0131  ;
  assign n21467 = ~n21465 & ~n21466 ;
  assign n21468 = ~\PIO_oe[2]_pad  & \pio_pmask_reg_DO_reg[2]/NET0131  ;
  assign n21469 = ~n21467 & n21468 ;
  assign n21470 = ~\pio_PINT_reg[2]/NET0131  & ~n21469 ;
  assign n21471 = ~n21291 & n21470 ;
  assign n21472 = ~n8715 & n21291 ;
  assign n21473 = ~n21471 & ~n21472 ;
  assign n21474 = \pio_PIO_RES_OUT_reg[10]/P0001  & ~\pio_PIO_RES_reg[10]/NET0131  ;
  assign n21475 = ~\pio_PIO_RES_OUT_reg[10]/P0001  & \pio_PIO_RES_reg[10]/NET0131  ;
  assign n21476 = ~n21474 & ~n21475 ;
  assign n21477 = ~\PIO_oe[10]_pad  & \pio_pmask_reg_DO_reg[10]/NET0131  ;
  assign n21478 = ~n21476 & n21477 ;
  assign n21479 = ~\pio_PINT_reg[10]/NET0131  & ~n21478 ;
  assign n21480 = ~n21291 & n21479 ;
  assign n21481 = ~n12688 & n21291 ;
  assign n21482 = ~n21480 & ~n21481 ;
  assign n21483 = \pio_PIO_RES_OUT_reg[0]/P0001  & ~\pio_PIO_RES_reg[0]/NET0131  ;
  assign n21484 = ~\pio_PIO_RES_OUT_reg[0]/P0001  & \pio_PIO_RES_reg[0]/NET0131  ;
  assign n21485 = ~n21483 & ~n21484 ;
  assign n21486 = ~\PIO_oe[0]_pad  & \pio_pmask_reg_DO_reg[0]/NET0131  ;
  assign n21487 = ~n21485 & n21486 ;
  assign n21488 = ~\pio_PINT_reg[0]/NET0131  & ~n21487 ;
  assign n21489 = ~n21291 & n21488 ;
  assign n21490 = ~n7607 & n21291 ;
  assign n21491 = ~n21489 & ~n21490 ;
  assign n21492 = \core_c_psq_Iact_E_reg[5]/NET0131  & ~n19477 ;
  assign n21493 = ~n19488 & n19491 ;
  assign n21494 = ~n19493 & n21493 ;
  assign n21495 = n19487 & n21494 ;
  assign n21496 = ~n21492 & ~n21495 ;
  assign n21497 = \pio_PIO_RES_OUT_reg[1]/P0001  & ~\pio_PIO_RES_reg[1]/NET0131  ;
  assign n21498 = ~\pio_PIO_RES_OUT_reg[1]/P0001  & \pio_PIO_RES_reg[1]/NET0131  ;
  assign n21499 = ~n21497 & ~n21498 ;
  assign n21500 = ~\PIO_oe[1]_pad  & \pio_pmask_reg_DO_reg[1]/NET0131  ;
  assign n21501 = ~n21499 & n21500 ;
  assign n21502 = ~\pio_PINT_reg[1]/NET0131  & ~n21501 ;
  assign n21503 = ~n21291 & n21502 ;
  assign n21504 = ~n9435 & n21291 ;
  assign n21505 = ~n21503 & ~n21504 ;
  assign n21506 = \pio_PIO_RES_OUT_reg[3]/P0001  & ~\pio_PIO_RES_reg[3]/NET0131  ;
  assign n21507 = ~\pio_PIO_RES_OUT_reg[3]/P0001  & \pio_PIO_RES_reg[3]/NET0131  ;
  assign n21508 = ~n21506 & ~n21507 ;
  assign n21509 = ~\PIO_oe[3]_pad  & \pio_pmask_reg_DO_reg[3]/NET0131  ;
  assign n21510 = ~n21508 & n21509 ;
  assign n21511 = ~\pio_PINT_reg[3]/NET0131  & ~n21510 ;
  assign n21512 = ~n21291 & n21511 ;
  assign n21513 = ~n8113 & n21291 ;
  assign n21514 = ~n21512 & ~n21513 ;
  assign n21515 = \pio_PIO_RES_OUT_reg[6]/P0001  & ~\pio_PIO_RES_reg[6]/NET0131  ;
  assign n21516 = ~\pio_PIO_RES_OUT_reg[6]/P0001  & \pio_PIO_RES_reg[6]/NET0131  ;
  assign n21517 = ~n21515 & ~n21516 ;
  assign n21518 = ~\PIO_oe[6]_pad  & \pio_pmask_reg_DO_reg[6]/NET0131  ;
  assign n21519 = ~n21517 & n21518 ;
  assign n21520 = ~\pio_PINT_reg[6]/NET0131  & ~n21519 ;
  assign n21521 = ~n21291 & n21520 ;
  assign n21522 = ~n11525 & n21291 ;
  assign n21523 = ~n21521 & ~n21522 ;
  assign n21524 = \core_eu_ea_alu_ea_dec_piconst_DO_reg[15]/P0001  & ~n20468 ;
  assign n21525 = \core_c_dec_IR_reg[4]/NET0131  & n14728 ;
  assign n21526 = n5664 & n21525 ;
  assign n21527 = \core_c_dec_IR_reg[11]/NET0131  & \core_c_dec_IR_reg[12]/NET0131  ;
  assign n21528 = \core_c_dec_IR_reg[7]/NET0131  & n21527 ;
  assign n21530 = ~\core_c_dec_IR_reg[5]/NET0131  & \core_c_dec_IR_reg[6]/NET0131  ;
  assign n21531 = n21528 & n21530 ;
  assign n21529 = \core_c_dec_IR_reg[5]/NET0131  & ~n21528 ;
  assign n21532 = ~n20477 & ~n21529 ;
  assign n21533 = ~n21531 & n21532 ;
  assign n21534 = n21526 & ~n21533 ;
  assign n21535 = ~n21524 & ~n21534 ;
  assign n21536 = \core_eu_ea_alu_ea_dec_piconst_DO_reg[14]/P0001  & ~n20468 ;
  assign n21537 = n20464 & n21528 ;
  assign n21538 = ~n20486 & ~n21529 ;
  assign n21539 = ~n21537 & n21538 ;
  assign n21540 = n21526 & ~n21539 ;
  assign n21541 = ~n21536 & ~n21540 ;
  assign n21542 = \core_eu_ea_alu_ea_dec_piconst_DO_reg[13]/P0001  & ~n20468 ;
  assign n21543 = ~\core_c_dec_IR_reg[7]/NET0131  & n21527 ;
  assign n21545 = n21530 & n21543 ;
  assign n21544 = \core_c_dec_IR_reg[5]/NET0131  & ~n21543 ;
  assign n21546 = ~n20477 & ~n21544 ;
  assign n21547 = ~n21545 & n21546 ;
  assign n21548 = n21526 & ~n21547 ;
  assign n21549 = ~n21542 & ~n21548 ;
  assign n21550 = \core_eu_ea_alu_ea_dec_piconst_DO_reg[12]/P0001  & ~n20468 ;
  assign n21551 = n20464 & n21543 ;
  assign n21552 = ~n20486 & ~n21544 ;
  assign n21553 = ~n21551 & n21552 ;
  assign n21554 = n21526 & ~n21553 ;
  assign n21555 = ~n21550 & ~n21554 ;
  assign n21559 = ~\core_c_dec_IR_reg[17]/NET0131  & n5615 ;
  assign n21560 = n19698 & n21559 ;
  assign n21556 = n6027 & n20606 ;
  assign n21557 = ~n4117 & n21556 ;
  assign n21558 = n6115 & n21557 ;
  assign n21561 = ~n20377 & ~n21558 ;
  assign n21562 = ~n21560 & n21561 ;
  assign n21565 = ~\sport0_rxctl_ldRX_cmp_reg/P0001  & n10069 ;
  assign n21566 = ~\sport0_rxctl_RX_reg[7]/P0001  & ~n20956 ;
  assign n21568 = ~n20949 & n21566 ;
  assign n21567 = n20949 & ~n21566 ;
  assign n21569 = n20875 & ~n21567 ;
  assign n21570 = ~n21568 & n21569 ;
  assign n21564 = \sport0_rxctl_RX_reg[4]/P0001  & n20873 ;
  assign n21571 = ~n20868 & ~n21564 ;
  assign n21572 = ~n21570 & n21571 ;
  assign n21573 = ~n21565 & n21572 ;
  assign n21563 = ~\sport0_rxctl_RXSHT_reg[4]/P0001  & n20868 ;
  assign n21574 = ~n20871 & ~n21563 ;
  assign n21575 = ~n21573 & n21574 ;
  assign n21576 = \sport0_rxctl_RX_reg[4]/P0001  & n20871 ;
  assign n21577 = ~n21575 & ~n21576 ;
  assign n21578 = n5692 & ~n5936 ;
  assign n21579 = ~n19705 & n21578 ;
  assign n21580 = \pio_PIO_RES_OUT_reg[7]/P0001  & ~\pio_PIO_RES_reg[7]/NET0131  ;
  assign n21581 = ~\pio_PIO_RES_OUT_reg[7]/P0001  & \pio_PIO_RES_reg[7]/NET0131  ;
  assign n21582 = ~n21580 & ~n21581 ;
  assign n21583 = ~\PIO_oe[7]_pad  & \pio_pmask_reg_DO_reg[7]/NET0131  ;
  assign n21584 = ~n21582 & n21583 ;
  assign n21585 = ~\pio_PINT_reg[7]/NET0131  & ~n21584 ;
  assign n21586 = ~n21291 & n21585 ;
  assign n21587 = ~n11265 & n21291 ;
  assign n21588 = ~n21586 & ~n21587 ;
  assign n21589 = ~\core_c_dec_IR_reg[4]/NET0131  & n19699 ;
  assign n21590 = n6111 & ~n21589 ;
  assign n21591 = ~n4117 & ~n21590 ;
  assign n21592 = n21578 & ~n21591 ;
  assign n21593 = \core_c_psq_SSTAT_reg[4]/NET0131  & ~n18217 ;
  assign n21594 = ~n18680 & n21593 ;
  assign n21595 = ~n14695 & ~n14702 ;
  assign n21596 = ~n14693 & ~n21595 ;
  assign n21597 = n18680 & n21596 ;
  assign n21598 = ~n21594 & ~n21597 ;
  assign n21599 = \emc_PMDoe_reg/NET0131  & ~n19049 ;
  assign n21600 = ~n19056 & n21599 ;
  assign n21601 = ~n20345 & ~n21600 ;
  assign n21602 = ~n14698 & ~n14710 ;
  assign n21603 = ~n18220 & n21602 ;
  assign n21604 = ~n18688 & ~n21602 ;
  assign n21605 = ~n21603 & ~n21604 ;
  assign n21606 = n4851 & n20576 ;
  assign n21607 = \core_c_psq_lpstk_lps4x22_LPcell_reg[3][9]/P0001  & ~n21606 ;
  assign n21608 = \core_c_dec_IRE_reg[5]/NET0131  & n21606 ;
  assign n21609 = ~n21607 & ~n21608 ;
  assign n21610 = \core_c_psq_lpstk_lps4x22_LPcell_reg[3][8]/P0001  & ~n21606 ;
  assign n21611 = \core_c_dec_IRE_reg[4]/NET0131  & n21606 ;
  assign n21612 = ~n21610 & ~n21611 ;
  assign n21613 = \core_c_psq_lpstk_lps4x22_LPcell_reg[3][7]/P0001  & ~n21606 ;
  assign n21614 = \core_c_dec_IRE_reg[3]/NET0131  & n21606 ;
  assign n21615 = ~n21613 & ~n21614 ;
  assign n21616 = \core_c_psq_lpstk_lps4x22_LPcell_reg[3][6]/P0001  & ~n21606 ;
  assign n21617 = \core_c_dec_IRE_reg[2]/NET0131  & n21606 ;
  assign n21618 = ~n21616 & ~n21617 ;
  assign n21619 = \core_c_psq_lpstk_lps4x22_LPcell_reg[3][5]/P0001  & ~n21606 ;
  assign n21620 = \core_c_dec_IRE_reg[1]/NET0131  & n21606 ;
  assign n21621 = ~n21619 & ~n21620 ;
  assign n21622 = \core_c_psq_lpstk_lps4x22_LPcell_reg[3][4]/P0001  & ~n21606 ;
  assign n21623 = \core_c_dec_IRE_reg[0]/NET0131  & n21606 ;
  assign n21624 = ~n21622 & ~n21623 ;
  assign n21625 = \core_c_psq_lpstk_lps4x22_LPcell_reg[3][21]/P0001  & ~n21606 ;
  assign n21626 = \core_c_dec_IRE_reg[17]/NET0131  & n21606 ;
  assign n21627 = ~n21625 & ~n21626 ;
  assign n21628 = \core_c_psq_lpstk_lps4x22_LPcell_reg[3][20]/P0001  & ~n21606 ;
  assign n21629 = \core_c_dec_IRE_reg[16]/NET0131  & n21606 ;
  assign n21630 = ~n21628 & ~n21629 ;
  assign n21631 = \core_c_psq_lpstk_lps4x22_LPcell_reg[3][19]/P0001  & ~n21606 ;
  assign n21632 = \core_c_dec_IRE_reg[15]/NET0131  & n21606 ;
  assign n21633 = ~n21631 & ~n21632 ;
  assign n21634 = \core_c_psq_lpstk_lps4x22_LPcell_reg[3][18]/P0001  & ~n21606 ;
  assign n21635 = \core_c_dec_IRE_reg[14]/NET0131  & n21606 ;
  assign n21636 = ~n21634 & ~n21635 ;
  assign n21637 = \core_c_psq_lpstk_lps4x22_LPcell_reg[3][17]/P0001  & ~n21606 ;
  assign n21638 = \core_c_dec_IRE_reg[13]/NET0131  & n21606 ;
  assign n21639 = ~n21637 & ~n21638 ;
  assign n21640 = \core_c_psq_lpstk_lps4x22_LPcell_reg[3][16]/P0001  & ~n21606 ;
  assign n21641 = \core_c_dec_IRE_reg[12]/NET0131  & n21606 ;
  assign n21642 = ~n21640 & ~n21641 ;
  assign n21643 = \core_c_psq_lpstk_lps4x22_LPcell_reg[3][15]/P0001  & ~n21606 ;
  assign n21644 = \core_c_dec_IRE_reg[11]/NET0131  & n21606 ;
  assign n21645 = ~n21643 & ~n21644 ;
  assign n21646 = \core_c_psq_lpstk_lps4x22_LPcell_reg[3][14]/P0001  & ~n21606 ;
  assign n21647 = \core_c_dec_IRE_reg[10]/NET0131  & n21606 ;
  assign n21648 = ~n21646 & ~n21647 ;
  assign n21649 = \core_c_psq_lpstk_lps4x22_LPcell_reg[3][13]/P0001  & ~n21606 ;
  assign n21650 = \core_c_dec_IRE_reg[9]/NET0131  & n21606 ;
  assign n21651 = ~n21649 & ~n21650 ;
  assign n21652 = \core_c_psq_lpstk_lps4x22_LPcell_reg[3][12]/P0001  & ~n21606 ;
  assign n21653 = \core_c_dec_IRE_reg[8]/NET0131  & n21606 ;
  assign n21654 = ~n21652 & ~n21653 ;
  assign n21655 = \core_c_psq_lpstk_lps4x22_LPcell_reg[3][11]/P0001  & ~n21606 ;
  assign n21656 = \core_c_dec_IRE_reg[7]/NET0131  & n21606 ;
  assign n21657 = ~n21655 & ~n21656 ;
  assign n21658 = \core_c_psq_lpstk_lps4x22_LPcell_reg[3][10]/P0001  & ~n21606 ;
  assign n21659 = \core_c_dec_IRE_reg[6]/NET0131  & n21606 ;
  assign n21660 = ~n21658 & ~n21659 ;
  assign n21661 = ~\core_c_dec_accPM_E_reg/P0001  & ~n8113 ;
  assign n21662 = \core_c_dec_accPM_E_reg/P0001  & ~n12870 ;
  assign n21663 = ~n21661 & ~n21662 ;
  assign n21664 = \core_c_dec_MTSR1_E_reg/P0001  & ~n21663 ;
  assign n21680 = n18043 & n18183 ;
  assign n21678 = ~n18091 & ~n18167 ;
  assign n21679 = ~n18104 & ~n18108 ;
  assign n21688 = ~n21678 & ~n21679 ;
  assign n21689 = ~n21680 & n21688 ;
  assign n21665 = n18088 & n19801 ;
  assign n21671 = n18046 & n18758 ;
  assign n21686 = ~n21665 & ~n21671 ;
  assign n21673 = ~n17922 & ~n18129 ;
  assign n21674 = n18147 & n18187 ;
  assign n21687 = ~n21673 & ~n21674 ;
  assign n21690 = n21686 & n21687 ;
  assign n21696 = n21689 & n21690 ;
  assign n21697 = n20087 & n21696 ;
  assign n21677 = ~n17933 & ~n18781 ;
  assign n21669 = n17925 & ~n18895 ;
  assign n21675 = ~n18175 & n20104 ;
  assign n21693 = ~n21669 & ~n21675 ;
  assign n21694 = ~n21677 & n21693 ;
  assign n21666 = n18111 & ~n19818 ;
  assign n21670 = \core_c_dec_IRE_reg[11]/NET0131  & ~n7991 ;
  assign n21672 = n18001 & n19720 ;
  assign n21682 = ~n21670 & ~n21672 ;
  assign n21676 = n17986 & ~n18189 ;
  assign n21681 = n18136 & n18153 ;
  assign n21683 = ~n21676 & ~n21681 ;
  assign n21684 = n21682 & n21683 ;
  assign n21685 = ~n17972 & n21684 ;
  assign n21691 = ~n21666 & n21685 ;
  assign n21667 = n18171 & ~n19857 ;
  assign n21668 = n18115 & ~n18775 ;
  assign n21692 = ~n21667 & ~n21668 ;
  assign n21695 = n21691 & n21692 ;
  assign n21698 = n21694 & n21695 ;
  assign n21699 = n21697 & n21698 ;
  assign n21700 = n21084 & n21699 ;
  assign n21701 = ~\core_c_dec_MTSR1_E_reg/P0001  & n21700 ;
  assign n21702 = ~n21664 & ~n21701 ;
  assign n21703 = n18717 & ~n21702 ;
  assign n21704 = ~\core_eu_es_sht_es_reg_sr1swe_DO_reg[3]/P0001  & ~n18717 ;
  assign n21705 = ~n21703 & ~n21704 ;
  assign n21706 = n4847 & n20576 ;
  assign n21707 = \core_c_psq_lpstk_lps4x22_LPcell_reg[2][9]/P0001  & ~n21706 ;
  assign n21708 = \core_c_dec_IRE_reg[5]/NET0131  & n21706 ;
  assign n21709 = ~n21707 & ~n21708 ;
  assign n21710 = \core_c_psq_lpstk_lps4x22_LPcell_reg[2][8]/P0001  & ~n21706 ;
  assign n21711 = \core_c_dec_IRE_reg[4]/NET0131  & n21706 ;
  assign n21712 = ~n21710 & ~n21711 ;
  assign n21713 = \core_c_psq_lpstk_lps4x22_LPcell_reg[2][7]/P0001  & ~n21706 ;
  assign n21714 = \core_c_dec_IRE_reg[3]/NET0131  & n21706 ;
  assign n21715 = ~n21713 & ~n21714 ;
  assign n21716 = \core_c_psq_lpstk_lps4x22_LPcell_reg[2][6]/P0001  & ~n21706 ;
  assign n21717 = \core_c_dec_IRE_reg[2]/NET0131  & n21706 ;
  assign n21718 = ~n21716 & ~n21717 ;
  assign n21719 = \core_c_psq_lpstk_lps4x22_LPcell_reg[2][5]/P0001  & ~n21706 ;
  assign n21720 = \core_c_dec_IRE_reg[1]/NET0131  & n21706 ;
  assign n21721 = ~n21719 & ~n21720 ;
  assign n21722 = \core_c_psq_lpstk_lps4x22_LPcell_reg[2][4]/P0001  & ~n21706 ;
  assign n21723 = \core_c_dec_IRE_reg[0]/NET0131  & n21706 ;
  assign n21724 = ~n21722 & ~n21723 ;
  assign n21725 = \core_c_psq_lpstk_lps4x22_LPcell_reg[2][21]/P0001  & ~n21706 ;
  assign n21726 = \core_c_dec_IRE_reg[17]/NET0131  & n21706 ;
  assign n21727 = ~n21725 & ~n21726 ;
  assign n21728 = \core_c_psq_lpstk_lps4x22_LPcell_reg[2][20]/P0001  & ~n21706 ;
  assign n21729 = \core_c_dec_IRE_reg[16]/NET0131  & n21706 ;
  assign n21730 = ~n21728 & ~n21729 ;
  assign n21731 = \core_c_psq_lpstk_lps4x22_LPcell_reg[2][19]/P0001  & ~n21706 ;
  assign n21732 = \core_c_dec_IRE_reg[15]/NET0131  & n21706 ;
  assign n21733 = ~n21731 & ~n21732 ;
  assign n21734 = \core_c_psq_lpstk_lps4x22_LPcell_reg[2][18]/P0001  & ~n21706 ;
  assign n21735 = \core_c_dec_IRE_reg[14]/NET0131  & n21706 ;
  assign n21736 = ~n21734 & ~n21735 ;
  assign n21737 = \core_c_psq_lpstk_lps4x22_LPcell_reg[2][17]/P0001  & ~n21706 ;
  assign n21738 = \core_c_dec_IRE_reg[13]/NET0131  & n21706 ;
  assign n21739 = ~n21737 & ~n21738 ;
  assign n21740 = \core_c_psq_lpstk_lps4x22_LPcell_reg[2][16]/P0001  & ~n21706 ;
  assign n21741 = \core_c_dec_IRE_reg[12]/NET0131  & n21706 ;
  assign n21742 = ~n21740 & ~n21741 ;
  assign n21743 = \core_c_psq_lpstk_lps4x22_LPcell_reg[2][15]/P0001  & ~n21706 ;
  assign n21744 = \core_c_dec_IRE_reg[11]/NET0131  & n21706 ;
  assign n21745 = ~n21743 & ~n21744 ;
  assign n21746 = \core_c_psq_lpstk_lps4x22_LPcell_reg[2][14]/P0001  & ~n21706 ;
  assign n21747 = \core_c_dec_IRE_reg[10]/NET0131  & n21706 ;
  assign n21748 = ~n21746 & ~n21747 ;
  assign n21749 = \core_c_psq_lpstk_lps4x22_LPcell_reg[2][13]/P0001  & ~n21706 ;
  assign n21750 = \core_c_dec_IRE_reg[9]/NET0131  & n21706 ;
  assign n21751 = ~n21749 & ~n21750 ;
  assign n21752 = \core_c_psq_lpstk_lps4x22_LPcell_reg[2][12]/P0001  & ~n21706 ;
  assign n21753 = \core_c_dec_IRE_reg[8]/NET0131  & n21706 ;
  assign n21754 = ~n21752 & ~n21753 ;
  assign n21755 = \core_c_psq_lpstk_lps4x22_LPcell_reg[2][11]/P0001  & ~n21706 ;
  assign n21756 = \core_c_dec_IRE_reg[7]/NET0131  & n21706 ;
  assign n21757 = ~n21755 & ~n21756 ;
  assign n21758 = \core_c_psq_lpstk_lps4x22_LPcell_reg[2][10]/P0001  & ~n21706 ;
  assign n21759 = \core_c_dec_IRE_reg[6]/NET0131  & n21706 ;
  assign n21760 = ~n21758 & ~n21759 ;
  assign n21761 = n20575 & n20597 ;
  assign n21762 = \core_c_psq_lpstk_lps4x22_LPcell_reg[1][9]/P0001  & ~n21761 ;
  assign n21763 = \core_c_dec_IRE_reg[5]/NET0131  & n21761 ;
  assign n21764 = ~n21762 & ~n21763 ;
  assign n21765 = \core_c_psq_lpstk_lps4x22_LPcell_reg[1][8]/P0001  & ~n21761 ;
  assign n21766 = \core_c_dec_IRE_reg[4]/NET0131  & n21761 ;
  assign n21767 = ~n21765 & ~n21766 ;
  assign n21768 = \core_c_psq_lpstk_lps4x22_LPcell_reg[1][7]/P0001  & ~n21761 ;
  assign n21769 = \core_c_dec_IRE_reg[3]/NET0131  & n21761 ;
  assign n21770 = ~n21768 & ~n21769 ;
  assign n21771 = \core_c_psq_lpstk_lps4x22_LPcell_reg[1][6]/P0001  & ~n21761 ;
  assign n21772 = \core_c_dec_IRE_reg[2]/NET0131  & n21761 ;
  assign n21773 = ~n21771 & ~n21772 ;
  assign n21774 = \core_c_psq_lpstk_lps4x22_LPcell_reg[1][5]/P0001  & ~n21761 ;
  assign n21775 = \core_c_dec_IRE_reg[1]/NET0131  & n21761 ;
  assign n21776 = ~n21774 & ~n21775 ;
  assign n21777 = \core_c_psq_lpstk_lps4x22_LPcell_reg[1][4]/P0001  & ~n21761 ;
  assign n21778 = \core_c_dec_IRE_reg[0]/NET0131  & n21761 ;
  assign n21779 = ~n21777 & ~n21778 ;
  assign n21780 = \core_c_psq_lpstk_lps4x22_LPcell_reg[1][21]/P0001  & ~n21761 ;
  assign n21781 = \core_c_dec_IRE_reg[17]/NET0131  & n21761 ;
  assign n21782 = ~n21780 & ~n21781 ;
  assign n21783 = \core_c_psq_lpstk_lps4x22_LPcell_reg[1][20]/P0001  & ~n21761 ;
  assign n21784 = \core_c_dec_IRE_reg[16]/NET0131  & n21761 ;
  assign n21785 = ~n21783 & ~n21784 ;
  assign n21786 = \core_c_psq_lpstk_lps4x22_LPcell_reg[1][19]/P0001  & ~n21761 ;
  assign n21787 = \core_c_dec_IRE_reg[15]/NET0131  & n21761 ;
  assign n21788 = ~n21786 & ~n21787 ;
  assign n21789 = \core_c_psq_lpstk_lps4x22_LPcell_reg[1][18]/P0001  & ~n21761 ;
  assign n21790 = \core_c_dec_IRE_reg[14]/NET0131  & n21761 ;
  assign n21791 = ~n21789 & ~n21790 ;
  assign n21792 = \core_c_psq_lpstk_lps4x22_LPcell_reg[1][17]/P0001  & ~n21761 ;
  assign n21793 = \core_c_dec_IRE_reg[13]/NET0131  & n21761 ;
  assign n21794 = ~n21792 & ~n21793 ;
  assign n21795 = \core_c_psq_lpstk_lps4x22_LPcell_reg[1][16]/P0001  & ~n21761 ;
  assign n21796 = \core_c_dec_IRE_reg[12]/NET0131  & n21761 ;
  assign n21797 = ~n21795 & ~n21796 ;
  assign n21798 = n13806 & ~n14649 ;
  assign n21799 = ~n13806 & ~n20053 ;
  assign n21800 = ~n21798 & ~n21799 ;
  assign n21801 = n14667 & ~n21800 ;
  assign n21802 = \core_eu_ea_alu_ea_reg_afswe_DO_reg[10]/P0001  & ~n14667 ;
  assign n21803 = ~n21801 & ~n21802 ;
  assign n21804 = \core_c_psq_lpstk_lps4x22_LPcell_reg[1][15]/P0001  & ~n21761 ;
  assign n21805 = \core_c_dec_IRE_reg[11]/NET0131  & n21761 ;
  assign n21806 = ~n21804 & ~n21805 ;
  assign n21807 = \core_c_psq_lpstk_lps4x22_LPcell_reg[1][14]/P0001  & ~n21761 ;
  assign n21808 = \core_c_dec_IRE_reg[10]/NET0131  & n21761 ;
  assign n21809 = ~n21807 & ~n21808 ;
  assign n21810 = \core_c_psq_lpstk_lps4x22_LPcell_reg[1][12]/P0001  & ~n21761 ;
  assign n21811 = \core_c_dec_IRE_reg[8]/NET0131  & n21761 ;
  assign n21812 = ~n21810 & ~n21811 ;
  assign n21813 = \core_c_psq_lpstk_lps4x22_LPcell_reg[1][11]/P0001  & ~n21761 ;
  assign n21814 = \core_c_dec_IRE_reg[7]/NET0131  & n21761 ;
  assign n21815 = ~n21813 & ~n21814 ;
  assign n21816 = \core_c_psq_lpstk_lps4x22_LPcell_reg[1][10]/P0001  & ~n21761 ;
  assign n21817 = \core_c_dec_IRE_reg[6]/NET0131  & n21761 ;
  assign n21818 = ~n21816 & ~n21817 ;
  assign n21819 = \core_c_psq_lpstk_lps4x22_LPcell_reg[0][9]/P0001  & ~n20595 ;
  assign n21820 = \core_c_dec_IRE_reg[5]/NET0131  & n20595 ;
  assign n21821 = ~n21819 & ~n21820 ;
  assign n21822 = \core_c_psq_lpstk_lps4x22_LPcell_reg[0][8]/P0001  & ~n20595 ;
  assign n21823 = \core_c_dec_IRE_reg[4]/NET0131  & n20595 ;
  assign n21824 = ~n21822 & ~n21823 ;
  assign n21825 = \core_c_psq_lpstk_lps4x22_LPcell_reg[0][6]/P0001  & ~n20595 ;
  assign n21826 = \core_c_dec_IRE_reg[2]/NET0131  & n20595 ;
  assign n21827 = ~n21825 & ~n21826 ;
  assign n21828 = \core_c_psq_lpstk_lps4x22_LPcell_reg[0][5]/P0001  & ~n20595 ;
  assign n21829 = \core_c_dec_IRE_reg[1]/NET0131  & n20595 ;
  assign n21830 = ~n21828 & ~n21829 ;
  assign n21831 = \core_c_psq_lpstk_lps4x22_LPcell_reg[0][4]/P0001  & ~n20595 ;
  assign n21832 = \core_c_dec_IRE_reg[0]/NET0131  & n20595 ;
  assign n21833 = ~n21831 & ~n21832 ;
  assign n21834 = n13805 & ~n21800 ;
  assign n21835 = \core_eu_ea_alu_ea_reg_afrwe_DO_reg[10]/P0001  & ~n13805 ;
  assign n21836 = ~n21834 & ~n21835 ;
  assign n21837 = \core_c_psq_lpstk_lps4x22_LPcell_reg[0][21]/P0001  & ~n20595 ;
  assign n21838 = \core_c_dec_IRE_reg[17]/NET0131  & n20595 ;
  assign n21839 = ~n21837 & ~n21838 ;
  assign n21840 = \core_c_psq_lpstk_lps4x22_LPcell_reg[0][20]/P0001  & ~n20595 ;
  assign n21841 = \core_c_dec_IRE_reg[16]/NET0131  & n20595 ;
  assign n21842 = ~n21840 & ~n21841 ;
  assign n21843 = \core_c_psq_lpstk_lps4x22_LPcell_reg[0][19]/P0001  & ~n20595 ;
  assign n21844 = \core_c_dec_IRE_reg[15]/NET0131  & n20595 ;
  assign n21845 = ~n21843 & ~n21844 ;
  assign n21846 = \core_c_psq_lpstk_lps4x22_LPcell_reg[0][18]/P0001  & ~n20595 ;
  assign n21847 = \core_c_dec_IRE_reg[14]/NET0131  & n20595 ;
  assign n21848 = ~n21846 & ~n21847 ;
  assign n21849 = \core_c_psq_lpstk_lps4x22_LPcell_reg[0][17]/P0001  & ~n20595 ;
  assign n21850 = \core_c_dec_IRE_reg[13]/NET0131  & n20595 ;
  assign n21851 = ~n21849 & ~n21850 ;
  assign n21852 = \core_c_psq_lpstk_lps4x22_LPcell_reg[0][15]/P0001  & ~n20595 ;
  assign n21853 = \core_c_dec_IRE_reg[11]/NET0131  & n20595 ;
  assign n21854 = ~n21852 & ~n21853 ;
  assign n21855 = \core_c_psq_lpstk_lps4x22_LPcell_reg[0][14]/P0001  & ~n20595 ;
  assign n21856 = \core_c_dec_IRE_reg[10]/NET0131  & n20595 ;
  assign n21857 = ~n21855 & ~n21856 ;
  assign n21858 = \core_c_psq_lpstk_lps4x22_LPcell_reg[0][13]/P0001  & ~n20595 ;
  assign n21859 = \core_c_dec_IRE_reg[9]/NET0131  & n20595 ;
  assign n21860 = ~n21858 & ~n21859 ;
  assign n21861 = \core_c_psq_lpstk_lps4x22_LPcell_reg[0][12]/P0001  & ~n20595 ;
  assign n21862 = \core_c_dec_IRE_reg[8]/NET0131  & n20595 ;
  assign n21863 = ~n21861 & ~n21862 ;
  assign n21864 = \core_c_psq_lpstk_lps4x22_LPcell_reg[0][11]/P0001  & ~n20595 ;
  assign n21865 = \core_c_dec_IRE_reg[7]/NET0131  & n20595 ;
  assign n21866 = ~n21864 & ~n21865 ;
  assign n21867 = \core_c_psq_lpstk_lps4x22_LPcell_reg[0][10]/P0001  & ~n20595 ;
  assign n21868 = \core_c_dec_IRE_reg[6]/NET0131  & n20595 ;
  assign n21869 = ~n21867 & ~n21868 ;
  assign n21870 = ~n13789 & ~n13794 ;
  assign n21871 = n13779 & n21870 ;
  assign n21872 = ~n13778 & ~n21870 ;
  assign n21873 = ~n21871 & ~n21872 ;
  assign n21874 = \core_c_psq_Iact_E_reg[4]/NET0131  & ~n4116 ;
  assign n21875 = \core_c_psq_T_IRQE1_reg/P0001  & ~\core_c_psq_T_IRQE1_s1_reg/P0001  ;
  assign n21876 = ~\core_c_psq_IFC_reg[12]/NET0131  & ~\core_c_psq_Iflag_reg[4]/NET0131  ;
  assign n21877 = ~n21875 & n21876 ;
  assign n21878 = ~\core_c_psq_IFC_reg[4]/NET0131  & ~n21877 ;
  assign n21879 = ~n21874 & n21878 ;
  assign n21880 = n14711 & ~n18220 ;
  assign n21881 = ~\core_c_psq_SSTAT_reg[5]/NET0131  & ~n21880 ;
  assign n21882 = \core_c_psq_lpstk_lps4x22_LPcell_reg[0][16]/P0001  & ~n20595 ;
  assign n21883 = \core_c_dec_IRE_reg[12]/NET0131  & n20595 ;
  assign n21884 = ~n21882 & ~n21883 ;
  assign n21885 = \bdma_DM_2nd_reg/NET0131  & ~n13753 ;
  assign n21886 = ~\bdma_DM_2nd_reg/NET0131  & n13753 ;
  assign n21887 = ~n21885 & ~n21886 ;
  assign n21888 = \core_c_psq_lpstk_lps4x22_LPcell_reg[0][7]/P0001  & ~n20595 ;
  assign n21889 = \core_c_dec_IRE_reg[3]/NET0131  & n20595 ;
  assign n21890 = ~n21888 & ~n21889 ;
  assign n21891 = ~\memc_MMR_web_reg/NET0131  & n13762 ;
  assign n21892 = n18230 & n21891 ;
  assign n21893 = ~n7340 & n21892 ;
  assign n21894 = ~\pio_pmask_reg_DO_reg[9]/NET0131  & ~n21892 ;
  assign n21895 = ~n21893 & ~n21894 ;
  assign n21896 = n18228 & n21891 ;
  assign n21897 = ~n9178 & n21896 ;
  assign n21898 = ~\PIO_oe[8]_pad  & ~n21896 ;
  assign n21899 = ~n21897 & ~n21898 ;
  assign n21900 = n17833 & ~n21702 ;
  assign n21901 = ~\core_eu_es_sht_es_reg_sr1rwe_DO_reg[3]/P0001  & ~n17833 ;
  assign n21902 = ~n21900 & ~n21901 ;
  assign n21903 = \core_c_psq_lpstk_lps4x22_LPcell_reg[1][13]/P0001  & ~n21761 ;
  assign n21904 = \core_c_dec_IRE_reg[9]/NET0131  & n21761 ;
  assign n21905 = ~n21903 & ~n21904 ;
  assign n21906 = n7526 & n18227 ;
  assign n21907 = ~n10289 & n21906 ;
  assign n21908 = ~\memc_usysr_DO_reg[9]/NET0131  & ~n21906 ;
  assign n21909 = ~n21907 & ~n21908 ;
  assign n21910 = ~n10638 & n21906 ;
  assign n21911 = ~\memc_usysr_DO_reg[8]/NET0131  & ~n21906 ;
  assign n21912 = ~n21910 & ~n21911 ;
  assign n21913 = ~n7340 & n21906 ;
  assign n21914 = ~\memc_usysr_DO_reg[13]/NET0131  & ~n21906 ;
  assign n21915 = ~n21913 & ~n21914 ;
  assign n21916 = ~n8460 & n21906 ;
  assign n21917 = ~\memc_usysr_DO_reg[11]/NET0131  & ~n21906 ;
  assign n21918 = ~n21916 & ~n21917 ;
  assign n21919 = ~n7859 & n21906 ;
  assign n21920 = ~\memc_usysr_DO_reg[10]/NET0131  & ~n21906 ;
  assign n21921 = ~n21919 & ~n21920 ;
  assign n21922 = n7232 & n18227 ;
  assign n21923 = n20070 & n21922 ;
  assign n21924 = ~n10289 & n21923 ;
  assign n21925 = ~\sport1_regs_SCLKDIVreg_DO_reg[9]/NET0131  & ~n21923 ;
  assign n21926 = ~n21924 & ~n21925 ;
  assign n21927 = ~n10638 & n21923 ;
  assign n21928 = ~\sport1_regs_SCLKDIVreg_DO_reg[8]/NET0131  & ~n21923 ;
  assign n21929 = ~n21927 & ~n21928 ;
  assign n21930 = \core_c_dec_MTSR0_E_reg/P0001  & ~n21663 ;
  assign n21933 = n17931 & ~n21157 ;
  assign n21937 = n17925 & n17991 ;
  assign n21939 = n18125 & ~n18918 ;
  assign n21947 = ~n21937 & ~n21939 ;
  assign n21940 = ~n18082 & n19720 ;
  assign n21943 = n18163 & ~n18914 ;
  assign n21948 = ~n21940 & ~n21943 ;
  assign n21949 = n21947 & n21948 ;
  assign n21955 = n18024 & n21949 ;
  assign n21956 = ~n21933 & n21955 ;
  assign n21942 = n18183 & ~n18898 ;
  assign n21938 = n18748 & ~n18888 ;
  assign n21941 = ~n17998 & n18187 ;
  assign n21952 = ~n21938 & ~n21941 ;
  assign n21953 = ~n21942 & n21952 ;
  assign n21931 = ~n18117 & ~n18909 ;
  assign n21936 = \core_c_dec_IRE_reg[11]/NET0131  & ~n7987 ;
  assign n21944 = ~n18026 & ~n21936 ;
  assign n21945 = ~n21931 & n21944 ;
  assign n21932 = ~n18079 & ~n18991 ;
  assign n21934 = ~n18104 & ~n18912 ;
  assign n21946 = ~n21932 & ~n21934 ;
  assign n21950 = n21945 & n21946 ;
  assign n21935 = n18083 & ~n18175 ;
  assign n21951 = n18903 & ~n21935 ;
  assign n21954 = n21950 & n21951 ;
  assign n21957 = n21953 & n21954 ;
  assign n21958 = n21956 & n21957 ;
  assign n21959 = ~\core_c_dec_MTSR0_E_reg/P0001  & n21958 ;
  assign n21960 = ~n21930 & ~n21959 ;
  assign n21961 = n18886 & ~n21960 ;
  assign n21962 = ~\core_eu_es_sht_es_reg_sr0swe_DO_reg[3]/P0001  & ~n18886 ;
  assign n21963 = ~n21961 & ~n21962 ;
  assign n21964 = ~n7340 & n21923 ;
  assign n21965 = ~\sport1_regs_SCLKDIVreg_DO_reg[13]/NET0131  & ~n21923 ;
  assign n21966 = ~n21964 & ~n21965 ;
  assign n21967 = ~n9178 & n21923 ;
  assign n21968 = ~\sport1_regs_SCLKDIVreg_DO_reg[12]/NET0131  & ~n21923 ;
  assign n21969 = ~n21967 & ~n21968 ;
  assign n21970 = ~n8460 & n21923 ;
  assign n21971 = ~\sport1_regs_SCLKDIVreg_DO_reg[11]/NET0131  & ~n21923 ;
  assign n21972 = ~n21970 & ~n21971 ;
  assign n21973 = ~n7859 & n21923 ;
  assign n21974 = ~\sport1_regs_SCLKDIVreg_DO_reg[10]/NET0131  & ~n21923 ;
  assign n21975 = ~n21973 & ~n21974 ;
  assign n21976 = n7526 & n21891 ;
  assign n21977 = ~n10638 & n21976 ;
  assign n21978 = ~\sport1_regs_AUTOreg_DO_reg[8]/NET0131  & ~n21976 ;
  assign n21979 = ~n21977 & ~n21978 ;
  assign n21980 = ~n10289 & n21976 ;
  assign n21981 = ~\sport1_regs_AUTOreg_DO_reg[9]/NET0131  & ~n21976 ;
  assign n21982 = ~n21980 & ~n21981 ;
  assign n21983 = ~n8460 & n21976 ;
  assign n21984 = ~\sport1_regs_AUTOreg_DO_reg[11]/NET0131  & ~n21976 ;
  assign n21985 = ~n21983 & ~n21984 ;
  assign n21986 = ~n7859 & n21976 ;
  assign n21987 = ~\sport1_regs_AUTOreg_DO_reg[10]/NET0131  & ~n21976 ;
  assign n21988 = ~n21986 & ~n21987 ;
  assign n21989 = ~\core_c_dec_MTAY0_E_reg/P0001  & n13799 ;
  assign n21990 = n14665 & ~n21989 ;
  assign n21991 = ~\core_c_dec_Double_E_reg/P0001  & ~\core_c_dec_accPM_E_reg/P0001  ;
  assign n21992 = ~n10289 & n21991 ;
  assign n21993 = ~n13075 & ~n21991 ;
  assign n21994 = ~n21992 & ~n21993 ;
  assign n21995 = ~n13806 & ~n21994 ;
  assign n21996 = n10453 & n13806 ;
  assign n21997 = ~n21995 & ~n21996 ;
  assign n21998 = n21990 & ~n21997 ;
  assign n21999 = ~\core_eu_ea_alu_ea_reg_ay0swe_DO_reg[9]/P0001  & ~n21990 ;
  assign n22000 = ~n21998 & ~n21999 ;
  assign n22001 = n13041 & ~n21991 ;
  assign n22002 = n10638 & n21991 ;
  assign n22003 = ~n22001 & ~n22002 ;
  assign n22004 = ~n13806 & n22003 ;
  assign n22005 = n11054 & n13806 ;
  assign n22006 = ~n22004 & ~n22005 ;
  assign n22007 = n21990 & ~n22006 ;
  assign n22008 = ~\core_eu_ea_alu_ea_reg_ay0swe_DO_reg[8]/P0001  & ~n21990 ;
  assign n22009 = ~n22007 & ~n22008 ;
  assign n22010 = ~n11265 & n21991 ;
  assign n22011 = ~n13006 & ~n21991 ;
  assign n22012 = ~n22010 & ~n22011 ;
  assign n22013 = ~n13806 & ~n22012 ;
  assign n22014 = n11329 & n13806 ;
  assign n22015 = ~n22013 & ~n22014 ;
  assign n22016 = n21990 & ~n22015 ;
  assign n22017 = ~\core_eu_ea_alu_ea_reg_ay0swe_DO_reg[7]/P0001  & ~n21990 ;
  assign n22018 = ~n22016 & ~n22017 ;
  assign n22019 = ~n11525 & n21991 ;
  assign n22020 = ~n12972 & ~n21991 ;
  assign n22021 = ~n22019 & ~n22020 ;
  assign n22022 = ~n13806 & ~n22021 ;
  assign n22023 = n10686 & n13806 ;
  assign n22024 = ~n22022 & ~n22023 ;
  assign n22025 = n21990 & ~n22024 ;
  assign n22026 = ~\core_eu_ea_alu_ea_reg_ay0swe_DO_reg[6]/P0001  & ~n21990 ;
  assign n22027 = ~n22025 & ~n22026 ;
  assign n22028 = ~n10911 & n21991 ;
  assign n22029 = ~n12938 & ~n21991 ;
  assign n22030 = ~n22028 & ~n22029 ;
  assign n22031 = ~n13806 & ~n22030 ;
  assign n22032 = n9904 & n13806 ;
  assign n22033 = ~n22031 & ~n22032 ;
  assign n22034 = n21990 & ~n22033 ;
  assign n22035 = ~\core_eu_ea_alu_ea_reg_ay0swe_DO_reg[5]/P0001  & ~n21990 ;
  assign n22036 = ~n22034 & ~n22035 ;
  assign n22037 = ~n10069 & n21991 ;
  assign n22038 = ~n12904 & ~n21991 ;
  assign n22039 = ~n22037 & ~n22038 ;
  assign n22040 = ~n13806 & ~n22039 ;
  assign n22041 = n7944 & n13806 ;
  assign n22042 = ~n22040 & ~n22041 ;
  assign n22043 = n21990 & ~n22042 ;
  assign n22044 = ~\core_eu_ea_alu_ea_reg_ay0swe_DO_reg[4]/P0001  & ~n21990 ;
  assign n22045 = ~n22043 & ~n22044 ;
  assign n22046 = ~n8113 & n21991 ;
  assign n22047 = ~n12870 & ~n21991 ;
  assign n22048 = ~n22046 & ~n22047 ;
  assign n22049 = ~n13806 & ~n22048 ;
  assign n22050 = n8577 & n13806 ;
  assign n22051 = ~n22049 & ~n22050 ;
  assign n22052 = n21990 & ~n22051 ;
  assign n22053 = ~\core_eu_ea_alu_ea_reg_ay0swe_DO_reg[3]/P0001  & ~n21990 ;
  assign n22054 = ~n22052 & ~n22053 ;
  assign n22055 = ~n8715 & n21991 ;
  assign n22056 = ~n12836 & ~n21991 ;
  assign n22057 = ~n22055 & ~n22056 ;
  assign n22058 = ~n13806 & ~n22057 ;
  assign n22059 = n9305 & n13806 ;
  assign n22060 = ~n22058 & ~n22059 ;
  assign n22061 = n21990 & ~n22060 ;
  assign n22062 = ~\core_eu_ea_alu_ea_reg_ay0swe_DO_reg[2]/P0001  & ~n21990 ;
  assign n22063 = ~n22061 & ~n22062 ;
  assign n22064 = ~n12743 & n21991 ;
  assign n22065 = ~n12771 & ~n21991 ;
  assign n22066 = ~n22064 & ~n22065 ;
  assign n22067 = ~n13806 & ~n22066 ;
  assign n22068 = n11829 & n13806 ;
  assign n22069 = ~n22067 & ~n22068 ;
  assign n22070 = n21990 & ~n22069 ;
  assign n22071 = ~\core_eu_ea_alu_ea_reg_ay0swe_DO_reg[15]/P0001  & ~n21990 ;
  assign n22072 = ~n22070 & ~n22071 ;
  assign n22073 = ~n12688 & n21991 ;
  assign n22074 = ~n12715 & ~n21991 ;
  assign n22075 = ~n22073 & ~n22074 ;
  assign n22076 = ~n13806 & ~n22075 ;
  assign n22077 = n7104 & n13806 ;
  assign n22078 = ~n22076 & ~n22077 ;
  assign n22079 = n21990 & ~n22078 ;
  assign n22080 = ~\core_eu_ea_alu_ea_reg_ay0swe_DO_reg[14]/P0001  & ~n21990 ;
  assign n22081 = ~n22079 & ~n22080 ;
  assign n22082 = ~n7340 & n21991 ;
  assign n22083 = ~n12658 & ~n21991 ;
  assign n22084 = ~n22082 & ~n22083 ;
  assign n22085 = ~n13806 & ~n22084 ;
  assign n22086 = n9095 & n13806 ;
  assign n22087 = ~n22085 & ~n22086 ;
  assign n22088 = n21990 & ~n22087 ;
  assign n22089 = ~\core_eu_ea_alu_ea_reg_ay0swe_DO_reg[13]/P0001  & ~n21990 ;
  assign n22090 = ~n22088 & ~n22089 ;
  assign n22091 = n12624 & ~n21991 ;
  assign n22092 = n9178 & n21991 ;
  assign n22093 = ~n22091 & ~n22092 ;
  assign n22094 = ~n13806 & n22093 ;
  assign n22095 = n8377 & n13806 ;
  assign n22096 = ~n22094 & ~n22095 ;
  assign n22097 = n21990 & ~n22096 ;
  assign n22098 = ~\core_eu_ea_alu_ea_reg_ay0swe_DO_reg[12]/P0001  & ~n21990 ;
  assign n22099 = ~n22097 & ~n22098 ;
  assign n22100 = n19034 & ~n21960 ;
  assign n22101 = ~\core_eu_es_sht_es_reg_sr0rwe_DO_reg[3]/P0001  & ~n19034 ;
  assign n22102 = ~n22100 & ~n22101 ;
  assign n22103 = n12590 & ~n21991 ;
  assign n22104 = n8460 & n21991 ;
  assign n22105 = ~n22103 & ~n22104 ;
  assign n22106 = ~n13806 & n22105 ;
  assign n22107 = n7776 & n13806 ;
  assign n22108 = ~n22106 & ~n22107 ;
  assign n22109 = n21990 & ~n22108 ;
  assign n22110 = ~\core_eu_ea_alu_ea_reg_ay0swe_DO_reg[11]/P0001  & ~n21990 ;
  assign n22111 = ~n22109 & ~n22110 ;
  assign n22112 = ~n7859 & n21991 ;
  assign n22113 = ~n12556 & ~n21991 ;
  assign n22114 = ~n22112 & ~n22113 ;
  assign n22115 = ~n13806 & ~n22114 ;
  assign n22116 = n10183 & n13806 ;
  assign n22117 = ~n22115 & ~n22116 ;
  assign n22118 = n21990 & ~n22117 ;
  assign n22119 = ~\core_eu_ea_alu_ea_reg_ay0swe_DO_reg[10]/P0001  & ~n21990 ;
  assign n22120 = ~n22118 & ~n22119 ;
  assign n22121 = ~n7340 & n21896 ;
  assign n22122 = ~\PIO_oe[9]_pad  & ~n21896 ;
  assign n22123 = ~n22121 & ~n22122 ;
  assign n22124 = n7283 & n21922 ;
  assign n22125 = ~n10289 & n22124 ;
  assign n22126 = ~\sport0_regs_SCLKDIVreg_DO_reg[9]/NET0131  & ~n22124 ;
  assign n22127 = ~n22125 & ~n22126 ;
  assign n22128 = ~n10638 & n22124 ;
  assign n22129 = ~\sport0_regs_SCLKDIVreg_DO_reg[8]/NET0131  & ~n22124 ;
  assign n22130 = ~n22128 & ~n22129 ;
  assign n22131 = ~n7340 & n22124 ;
  assign n22132 = ~\sport0_regs_SCLKDIVreg_DO_reg[13]/NET0131  & ~n22124 ;
  assign n22133 = ~n22131 & ~n22132 ;
  assign n22134 = ~n9178 & n22124 ;
  assign n22135 = ~\sport0_regs_SCLKDIVreg_DO_reg[12]/NET0131  & ~n22124 ;
  assign n22136 = ~n22134 & ~n22135 ;
  assign n22137 = ~n8460 & n22124 ;
  assign n22138 = ~\sport0_regs_SCLKDIVreg_DO_reg[11]/NET0131  & ~n22124 ;
  assign n22139 = ~n22137 & ~n22138 ;
  assign n22140 = ~n7859 & n22124 ;
  assign n22141 = ~\sport0_regs_SCLKDIVreg_DO_reg[10]/NET0131  & ~n22124 ;
  assign n22142 = ~n22140 & ~n22141 ;
  assign n22143 = ~n9178 & n21892 ;
  assign n22144 = ~\pio_pmask_reg_DO_reg[8]/NET0131  & ~n21892 ;
  assign n22145 = ~n22143 & ~n22144 ;
  assign n22146 = ~n9178 & n20401 ;
  assign n22147 = ~\sport0_regs_AUTO_a_reg[12]/NET0131  & ~n20401 ;
  assign n22148 = ~n22146 & ~n22147 ;
  assign n22149 = ~n9435 & n21991 ;
  assign n22150 = ~n12802 & ~n21991 ;
  assign n22151 = ~n22149 & ~n22150 ;
  assign n22152 = ~n13806 & n22151 ;
  assign n22153 = ~n7414 & n13806 ;
  assign n22154 = ~n22152 & ~n22153 ;
  assign n22155 = n21990 & ~n22154 ;
  assign n22156 = \core_eu_ea_alu_ea_reg_ay0swe_DO_reg[1]/P0001  & ~n21990 ;
  assign n22157 = ~n22155 & ~n22156 ;
  assign n22158 = n17798 & ~n21989 ;
  assign n22159 = ~n21997 & n22158 ;
  assign n22160 = ~\core_eu_ea_alu_ea_reg_ay0rwe_DO_reg[9]/P0001  & ~n22158 ;
  assign n22161 = ~n22159 & ~n22160 ;
  assign n22162 = ~n22006 & n22158 ;
  assign n22163 = ~\core_eu_ea_alu_ea_reg_ay0rwe_DO_reg[8]/P0001  & ~n22158 ;
  assign n22164 = ~n22162 & ~n22163 ;
  assign n22165 = ~n22015 & n22158 ;
  assign n22166 = ~\core_eu_ea_alu_ea_reg_ay0rwe_DO_reg[7]/P0001  & ~n22158 ;
  assign n22167 = ~n22165 & ~n22166 ;
  assign n22168 = ~n22024 & n22158 ;
  assign n22169 = ~\core_eu_ea_alu_ea_reg_ay0rwe_DO_reg[6]/P0001  & ~n22158 ;
  assign n22170 = ~n22168 & ~n22169 ;
  assign n22171 = ~n22033 & n22158 ;
  assign n22172 = ~\core_eu_ea_alu_ea_reg_ay0rwe_DO_reg[5]/P0001  & ~n22158 ;
  assign n22173 = ~n22171 & ~n22172 ;
  assign n22174 = ~n22042 & n22158 ;
  assign n22175 = ~\core_eu_ea_alu_ea_reg_ay0rwe_DO_reg[4]/P0001  & ~n22158 ;
  assign n22176 = ~n22174 & ~n22175 ;
  assign n22177 = ~n22051 & n22158 ;
  assign n22178 = ~\core_eu_ea_alu_ea_reg_ay0rwe_DO_reg[3]/P0001  & ~n22158 ;
  assign n22179 = ~n22177 & ~n22178 ;
  assign n22180 = ~n22060 & n22158 ;
  assign n22181 = ~\core_eu_ea_alu_ea_reg_ay0rwe_DO_reg[2]/P0001  & ~n22158 ;
  assign n22182 = ~n22180 & ~n22181 ;
  assign n22183 = ~n22154 & n22158 ;
  assign n22184 = \core_eu_ea_alu_ea_reg_ay0rwe_DO_reg[1]/P0001  & ~n22158 ;
  assign n22185 = ~n22183 & ~n22184 ;
  assign n22186 = ~n22069 & n22158 ;
  assign n22187 = ~\core_eu_ea_alu_ea_reg_ay0rwe_DO_reg[15]/P0001  & ~n22158 ;
  assign n22188 = ~n22186 & ~n22187 ;
  assign n22189 = ~n22078 & n22158 ;
  assign n22190 = ~\core_eu_ea_alu_ea_reg_ay0rwe_DO_reg[14]/P0001  & ~n22158 ;
  assign n22191 = ~n22189 & ~n22190 ;
  assign n22192 = ~n22087 & n22158 ;
  assign n22193 = ~\core_eu_ea_alu_ea_reg_ay0rwe_DO_reg[13]/P0001  & ~n22158 ;
  assign n22194 = ~n22192 & ~n22193 ;
  assign n22195 = ~n22096 & n22158 ;
  assign n22196 = ~\core_eu_ea_alu_ea_reg_ay0rwe_DO_reg[12]/P0001  & ~n22158 ;
  assign n22197 = ~n22195 & ~n22196 ;
  assign n22198 = ~n22108 & n22158 ;
  assign n22199 = ~\core_eu_ea_alu_ea_reg_ay0rwe_DO_reg[11]/P0001  & ~n22158 ;
  assign n22200 = ~n22198 & ~n22199 ;
  assign n22201 = ~n22117 & n22158 ;
  assign n22202 = ~\core_eu_ea_alu_ea_reg_ay0rwe_DO_reg[10]/P0001  & ~n22158 ;
  assign n22203 = ~n22201 & ~n22202 ;
  assign n22204 = ~n12743 & n22124 ;
  assign n22205 = ~\sport0_regs_SCLKDIVreg_DO_reg[15]/NET0131  & ~n22124 ;
  assign n22206 = ~n22204 & ~n22205 ;
  assign n22207 = ~n8113 & n22124 ;
  assign n22208 = ~\sport0_regs_SCLKDIVreg_DO_reg[3]/NET0131  & ~n22124 ;
  assign n22209 = ~n22207 & ~n22208 ;
  assign n22210 = ~n10911 & n22124 ;
  assign n22211 = ~\sport0_regs_SCLKDIVreg_DO_reg[5]/NET0131  & ~n22124 ;
  assign n22212 = ~n22210 & ~n22211 ;
  assign n22213 = ~n12743 & n20401 ;
  assign n22214 = ~\sport0_regs_AUTO_a_reg[15]/NET0131  & ~n20401 ;
  assign n22215 = ~n22213 & ~n22214 ;
  assign n22216 = ~n11265 & n21892 ;
  assign n22217 = ~\pio_pmask_reg_DO_reg[7]/NET0131  & ~n21892 ;
  assign n22218 = ~n22216 & ~n22217 ;
  assign n22219 = ~n11525 & n21892 ;
  assign n22220 = ~\pio_pmask_reg_DO_reg[6]/NET0131  & ~n21892 ;
  assign n22221 = ~n22219 & ~n22220 ;
  assign n22222 = ~n8113 & n21892 ;
  assign n22223 = ~\pio_pmask_reg_DO_reg[3]/NET0131  & ~n21892 ;
  assign n22224 = ~n22222 & ~n22223 ;
  assign n22225 = ~n12743 & n21892 ;
  assign n22226 = ~\pio_pmask_reg_DO_reg[11]/NET0131  & ~n21892 ;
  assign n22227 = ~n22225 & ~n22226 ;
  assign n22228 = ~\sice_ICYC_reg[18]/NET0131  & ~n20747 ;
  assign n22229 = ~n20748 & ~n22228 ;
  assign n22230 = ~n8715 & n21892 ;
  assign n22231 = ~\pio_pmask_reg_DO_reg[2]/NET0131  & ~n21892 ;
  assign n22232 = ~n22230 & ~n22231 ;
  assign n22233 = ~n7607 & n21892 ;
  assign n22234 = ~\pio_pmask_reg_DO_reg[0]/NET0131  & ~n21892 ;
  assign n22235 = ~n22233 & ~n22234 ;
  assign n22236 = ~n11265 & n21896 ;
  assign n22237 = ~\PIO_oe[7]_pad  & ~n21896 ;
  assign n22238 = ~n22236 & ~n22237 ;
  assign n22239 = ~n11525 & n21896 ;
  assign n22240 = ~\PIO_oe[6]_pad  & ~n21896 ;
  assign n22241 = ~n22239 & ~n22240 ;
  assign n22242 = ~n10069 & n21896 ;
  assign n22243 = ~\PIO_oe[4]_pad  & ~n21896 ;
  assign n22244 = ~n22242 & ~n22243 ;
  assign n22245 = ~n8715 & n21896 ;
  assign n22246 = ~\PIO_oe[2]_pad  & ~n21896 ;
  assign n22247 = ~n22245 & ~n22246 ;
  assign n22248 = ~n9435 & n21896 ;
  assign n22249 = ~\PIO_oe[1]_pad  & ~n21896 ;
  assign n22250 = ~n22248 & ~n22249 ;
  assign n22251 = ~n12743 & n21896 ;
  assign n22252 = ~\PIO_oe[11]_pad  & ~n21896 ;
  assign n22253 = ~n22251 & ~n22252 ;
  assign n22254 = ~n11265 & n21906 ;
  assign n22255 = ~\memc_usysr_DO_reg[7]/NET0131  & ~n21906 ;
  assign n22256 = ~n22254 & ~n22255 ;
  assign n22257 = ~n12688 & n21892 ;
  assign n22258 = ~\pio_pmask_reg_DO_reg[10]/NET0131  & ~n21892 ;
  assign n22259 = ~n22257 & ~n22258 ;
  assign n22260 = ~n10911 & n21892 ;
  assign n22261 = ~\pio_pmask_reg_DO_reg[5]/NET0131  & ~n21892 ;
  assign n22262 = ~n22260 & ~n22261 ;
  assign n22263 = ~n10911 & n21906 ;
  assign n22264 = ~\memc_usysr_DO_reg[5]/NET0131  & ~n21906 ;
  assign n22265 = ~n22263 & ~n22264 ;
  assign n22266 = ~n11525 & n21906 ;
  assign n22267 = ~\memc_usysr_DO_reg[6]/NET0131  & ~n21906 ;
  assign n22268 = ~n22266 & ~n22267 ;
  assign n22269 = ~n10069 & n21906 ;
  assign n22270 = ~\memc_usysr_DO_reg[4]/NET0131  & ~n21906 ;
  assign n22271 = ~n22269 & ~n22270 ;
  assign n22272 = ~n8715 & n21906 ;
  assign n22273 = ~\memc_usysr_DO_reg[2]/NET0131  & ~n21906 ;
  assign n22274 = ~n22272 & ~n22273 ;
  assign n22275 = ~n9435 & n21906 ;
  assign n22276 = ~\memc_usysr_DO_reg[1]/NET0131  & ~n21906 ;
  assign n22277 = ~n22275 & ~n22276 ;
  assign n22278 = ~n12743 & n21906 ;
  assign n22279 = ~\memc_usysr_DO_reg[15]/NET0131  & ~n21906 ;
  assign n22280 = ~n22278 & ~n22279 ;
  assign n22281 = ~n12688 & n21906 ;
  assign n22282 = ~\memc_usysr_DO_reg[14]/NET0131  & ~n21906 ;
  assign n22283 = ~n22281 & ~n22282 ;
  assign n22284 = ~n7607 & n21906 ;
  assign n22285 = ~\memc_usysr_DO_reg[0]/NET0131  & ~n21906 ;
  assign n22286 = ~n22284 & ~n22285 ;
  assign n22287 = \idma_RDcyc_reg/NET0131  & n20393 ;
  assign n22288 = ~n20821 & ~n22287 ;
  assign n22289 = n7261 & n7525 ;
  assign n22290 = n18226 & n22289 ;
  assign n22291 = ~\memc_MMR_web_reg/NET0131  & n22290 ;
  assign n22292 = ~n8460 & n22291 ;
  assign n22293 = ~\tm_tcr_reg_DO_reg[11]/NET0131  & ~n22291 ;
  assign n22294 = ~n22292 & ~n22293 ;
  assign n22295 = ~n8113 & n21896 ;
  assign n22296 = ~\PIO_oe[3]_pad  & ~n21896 ;
  assign n22297 = ~n22295 & ~n22296 ;
  assign n22298 = n7513 & n21891 ;
  assign n22299 = ~n11265 & n22298 ;
  assign n22300 = ~\emc_WSCRext_reg_DO_reg[7]/NET0131  & ~n22298 ;
  assign n22301 = ~n22299 & ~n22300 ;
  assign n22302 = ~n11525 & n22298 ;
  assign n22303 = ~\emc_WSCRext_reg_DO_reg[6]/NET0131  & ~n22298 ;
  assign n22304 = ~n22302 & ~n22303 ;
  assign n22305 = ~n10911 & n22298 ;
  assign n22306 = ~\emc_WSCRext_reg_DO_reg[5]/NET0131  & ~n22298 ;
  assign n22307 = ~n22305 & ~n22306 ;
  assign n22308 = ~n10069 & n22298 ;
  assign n22309 = ~\emc_WSCRext_reg_DO_reg[4]/NET0131  & ~n22298 ;
  assign n22310 = ~n22308 & ~n22309 ;
  assign n22311 = ~n8113 & n22298 ;
  assign n22312 = ~\emc_WSCRext_reg_DO_reg[3]/NET0131  & ~n22298 ;
  assign n22313 = ~n22311 & ~n22312 ;
  assign n22314 = ~n8715 & n22298 ;
  assign n22315 = ~\emc_WSCRext_reg_DO_reg[2]/NET0131  & ~n22298 ;
  assign n22316 = ~n22314 & ~n22315 ;
  assign n22317 = ~n9435 & n22298 ;
  assign n22318 = ~\emc_WSCRext_reg_DO_reg[1]/NET0131  & ~n22298 ;
  assign n22319 = ~n22317 & ~n22318 ;
  assign n22320 = ~n7607 & n22298 ;
  assign n22321 = ~\emc_WSCRext_reg_DO_reg[0]/NET0131  & ~n22298 ;
  assign n22322 = ~n22320 & ~n22321 ;
  assign n22323 = ~n11265 & n21923 ;
  assign n22324 = ~\sport1_regs_SCLKDIVreg_DO_reg[7]/NET0131  & ~n21923 ;
  assign n22325 = ~n22323 & ~n22324 ;
  assign n22326 = ~n11525 & n21923 ;
  assign n22327 = ~\sport1_regs_SCLKDIVreg_DO_reg[6]/NET0131  & ~n21923 ;
  assign n22328 = ~n22326 & ~n22327 ;
  assign n22329 = ~n10911 & n21923 ;
  assign n22330 = ~\sport1_regs_SCLKDIVreg_DO_reg[5]/NET0131  & ~n21923 ;
  assign n22331 = ~n22329 & ~n22330 ;
  assign n22332 = ~n10069 & n21923 ;
  assign n22333 = ~\sport1_regs_SCLKDIVreg_DO_reg[4]/NET0131  & ~n21923 ;
  assign n22334 = ~n22332 & ~n22333 ;
  assign n22335 = ~n8113 & n21923 ;
  assign n22336 = ~\sport1_regs_SCLKDIVreg_DO_reg[3]/NET0131  & ~n21923 ;
  assign n22337 = ~n22335 & ~n22336 ;
  assign n22338 = ~n8715 & n21923 ;
  assign n22339 = ~\sport1_regs_SCLKDIVreg_DO_reg[2]/NET0131  & ~n21923 ;
  assign n22340 = ~n22338 & ~n22339 ;
  assign n22341 = ~n9435 & n21923 ;
  assign n22342 = ~\sport1_regs_SCLKDIVreg_DO_reg[1]/NET0131  & ~n21923 ;
  assign n22343 = ~n22341 & ~n22342 ;
  assign n22344 = ~n12743 & n21923 ;
  assign n22345 = ~\sport1_regs_SCLKDIVreg_DO_reg[15]/NET0131  & ~n21923 ;
  assign n22346 = ~n22344 & ~n22345 ;
  assign n22347 = ~n12688 & n21923 ;
  assign n22348 = ~\sport1_regs_SCLKDIVreg_DO_reg[14]/NET0131  & ~n21923 ;
  assign n22349 = ~n22347 & ~n22348 ;
  assign n22350 = ~n7607 & n21923 ;
  assign n22351 = ~\sport1_regs_SCLKDIVreg_DO_reg[0]/NET0131  & ~n21923 ;
  assign n22352 = ~n22350 & ~n22351 ;
  assign n22353 = ~n11265 & n21976 ;
  assign n22354 = ~\sport1_regs_AUTOreg_DO_reg[7]/NET0131  & ~n21976 ;
  assign n22355 = ~n22353 & ~n22354 ;
  assign n22356 = ~n11525 & n21976 ;
  assign n22357 = ~\sport1_regs_AUTOreg_DO_reg[6]/NET0131  & ~n21976 ;
  assign n22358 = ~n22356 & ~n22357 ;
  assign n22359 = ~n10911 & n21976 ;
  assign n22360 = ~\sport1_regs_AUTOreg_DO_reg[5]/NET0131  & ~n21976 ;
  assign n22361 = ~n22359 & ~n22360 ;
  assign n22362 = ~n10069 & n21976 ;
  assign n22363 = ~\sport1_regs_AUTOreg_DO_reg[4]/NET0131  & ~n21976 ;
  assign n22364 = ~n22362 & ~n22363 ;
  assign n22365 = ~n8113 & n21976 ;
  assign n22366 = ~\sport1_regs_AUTOreg_DO_reg[3]/NET0131  & ~n21976 ;
  assign n22367 = ~n22365 & ~n22366 ;
  assign n22368 = ~n8715 & n21976 ;
  assign n22369 = ~\sport1_regs_AUTOreg_DO_reg[2]/NET0131  & ~n21976 ;
  assign n22370 = ~n22368 & ~n22369 ;
  assign n22371 = ~n9435 & n21976 ;
  assign n22372 = ~\sport1_regs_AUTOreg_DO_reg[1]/NET0131  & ~n21976 ;
  assign n22373 = ~n22371 & ~n22372 ;
  assign n22374 = ~n7607 & n21976 ;
  assign n22375 = ~\sport1_regs_AUTOreg_DO_reg[0]/NET0131  & ~n21976 ;
  assign n22376 = ~n22374 & ~n22375 ;
  assign n22377 = ~n10911 & n21896 ;
  assign n22378 = ~\PIO_oe[5]_pad  & ~n21896 ;
  assign n22379 = ~n22377 & ~n22378 ;
  assign n22380 = ~n10069 & n21892 ;
  assign n22381 = ~\pio_pmask_reg_DO_reg[4]/NET0131  & ~n21892 ;
  assign n22382 = ~n22380 & ~n22381 ;
  assign n22383 = ~n7607 & n21896 ;
  assign n22384 = ~\PIO_oe[0]_pad  & ~n21896 ;
  assign n22385 = ~n22383 & ~n22384 ;
  assign n22386 = \sport0_regs_AUTO_a_reg[14]/NET0131  & ~n20401 ;
  assign n22387 = n18235 & n20400 ;
  assign n22388 = ~n22386 & ~n22387 ;
  assign n22389 = ~n9435 & n21892 ;
  assign n22390 = ~\pio_pmask_reg_DO_reg[1]/NET0131  & ~n21892 ;
  assign n22391 = ~n22389 & ~n22390 ;
  assign n22392 = ~n8113 & n21906 ;
  assign n22393 = ~\memc_usysr_DO_reg[3]/NET0131  & ~n21906 ;
  assign n22394 = ~n22392 & ~n22393 ;
  assign n22395 = ~n12688 & n21896 ;
  assign n22396 = ~\PIO_oe[10]_pad  & ~n21896 ;
  assign n22397 = ~n22395 & ~n22396 ;
  assign n22398 = \tm_tcr_reg_DO_reg[10]/NET0131  & n20355 ;
  assign n22399 = ~\T_TMODE[0]_pad  & \core_c_psq_MSTAT_reg_DO_reg[5]/NET0131  ;
  assign n22400 = n20372 & n22399 ;
  assign n22402 = ~\tm_TSR_TMP_reg[1]/NET0131  & ~\tm_TSR_TMP_reg[2]/NET0131  ;
  assign n22403 = ~\tm_TSR_TMP_reg[0]/NET0131  & ~\tm_TSR_TMP_reg[3]/NET0131  ;
  assign n22404 = n22402 & n22403 ;
  assign n22405 = ~\tm_TSR_TMP_reg[4]/NET0131  & ~\tm_TSR_TMP_reg[5]/NET0131  ;
  assign n22406 = ~\tm_TSR_TMP_reg[6]/NET0131  & ~\tm_TSR_TMP_reg[7]/NET0131  ;
  assign n22407 = n22405 & n22406 ;
  assign n22408 = n22404 & n22407 ;
  assign n22409 = \core_c_psq_MSTAT_reg_DO_reg[5]/NET0131  & n22408 ;
  assign n22410 = ~\T_TMODE[0]_pad  & ~n22409 ;
  assign n22411 = ~\core_c_psq_PCS_reg[3]/NET0131  & ~n22410 ;
  assign n22412 = ~\tm_TCR_TMP_reg[10]/NET0131  & ~n22411 ;
  assign n22413 = ~\T_TMODE[0]_pad  & ~n20364 ;
  assign n22414 = \tm_TCR_TMP_reg[8]/NET0131  & n22413 ;
  assign n22415 = \tm_TCR_TMP_reg[9]/NET0131  & n22414 ;
  assign n22416 = ~\tm_TCR_TMP_reg[10]/NET0131  & ~n22415 ;
  assign n22417 = \tm_TCR_TMP_reg[10]/NET0131  & n22415 ;
  assign n22418 = ~n22416 & ~n22417 ;
  assign n22419 = ~\tm_TCR_TMP_reg[9]/NET0131  & ~n22414 ;
  assign n22420 = ~n22415 & ~n22419 ;
  assign n22421 = ~\tm_TCR_TMP_reg[8]/NET0131  & ~n22413 ;
  assign n22422 = ~n22414 & ~n22421 ;
  assign n22423 = ~n22420 & ~n22422 ;
  assign n22425 = n22418 & ~n22423 ;
  assign n22424 = ~n22418 & n22423 ;
  assign n22426 = n22411 & ~n22424 ;
  assign n22427 = ~n22425 & n22426 ;
  assign n22428 = ~n22412 & ~n22427 ;
  assign n22429 = ~n22400 & ~n22428 ;
  assign n22401 = ~\tm_tpr_reg_DO_reg[10]/NET0131  & n22400 ;
  assign n22430 = ~n20355 & ~n22401 ;
  assign n22431 = ~n22429 & n22430 ;
  assign n22432 = ~n22398 & ~n22431 ;
  assign n22433 = ~n11265 & n22124 ;
  assign n22434 = ~\sport0_regs_SCLKDIVreg_DO_reg[7]/NET0131  & ~n22124 ;
  assign n22435 = ~n22433 & ~n22434 ;
  assign n22436 = ~n11525 & n22124 ;
  assign n22437 = ~\sport0_regs_SCLKDIVreg_DO_reg[6]/NET0131  & ~n22124 ;
  assign n22438 = ~n22436 & ~n22437 ;
  assign n22439 = ~n10069 & n22124 ;
  assign n22440 = ~\sport0_regs_SCLKDIVreg_DO_reg[4]/NET0131  & ~n22124 ;
  assign n22441 = ~n22439 & ~n22440 ;
  assign n22442 = ~n8715 & n22124 ;
  assign n22443 = ~\sport0_regs_SCLKDIVreg_DO_reg[2]/NET0131  & ~n22124 ;
  assign n22444 = ~n22442 & ~n22443 ;
  assign n22445 = ~n9435 & n22124 ;
  assign n22446 = ~\sport0_regs_SCLKDIVreg_DO_reg[1]/NET0131  & ~n22124 ;
  assign n22447 = ~n22445 & ~n22446 ;
  assign n22448 = ~n12688 & n22124 ;
  assign n22449 = ~\sport0_regs_SCLKDIVreg_DO_reg[14]/NET0131  & ~n22124 ;
  assign n22450 = ~n22448 & ~n22449 ;
  assign n22451 = ~n7607 & n22124 ;
  assign n22452 = ~\sport0_regs_SCLKDIVreg_DO_reg[0]/NET0131  & ~n22124 ;
  assign n22453 = ~n22451 & ~n22452 ;
  assign n22454 = \core_c_psq_Iact_E_reg[8]/NET0131  & ~n19477 ;
  assign n22455 = n19484 & n19486 ;
  assign n22456 = ~n22454 & ~n22455 ;
  assign n22457 = n7237 & n18227 ;
  assign n22458 = n7269 & n22457 ;
  assign n22459 = ~n10289 & n22458 ;
  assign n22460 = ~\clkc_ckr_reg_DO_reg[9]/NET0131  & ~n22458 ;
  assign n22461 = ~n22459 & ~n22460 ;
  assign n22462 = ~n10638 & n22458 ;
  assign n22463 = ~\clkc_ckr_reg_DO_reg[8]/NET0131  & ~n22458 ;
  assign n22464 = ~n22462 & ~n22463 ;
  assign n22465 = ~n7340 & n22458 ;
  assign n22466 = ~\clkc_ckr_reg_DO_reg[13]/NET0131  & ~n22458 ;
  assign n22467 = ~n22465 & ~n22466 ;
  assign n22468 = ~n9178 & n22458 ;
  assign n22469 = ~\clkc_ckr_reg_DO_reg[12]/NET0131  & ~n22458 ;
  assign n22470 = ~n22468 & ~n22469 ;
  assign n22471 = ~n7859 & n22458 ;
  assign n22472 = ~\clkc_ckr_reg_DO_reg[10]/NET0131  & ~n22458 ;
  assign n22473 = ~n22471 & ~n22472 ;
  assign n22474 = ~n8460 & n22458 ;
  assign n22475 = ~\clkc_ckr_reg_DO_reg[11]/NET0131  & ~n22458 ;
  assign n22476 = ~n22474 & ~n22475 ;
  assign n22477 = n7525 & n21922 ;
  assign n22478 = ~n8460 & n22477 ;
  assign n22479 = ~\tm_tpr_reg_DO_reg[11]/NET0131  & ~n22477 ;
  assign n22480 = ~n22478 & ~n22479 ;
  assign n22481 = ~n7859 & n22477 ;
  assign n22482 = ~\tm_tpr_reg_DO_reg[10]/NET0131  & ~n22477 ;
  assign n22483 = ~n22481 & ~n22482 ;
  assign n22484 = n7525 & n22457 ;
  assign n22485 = ~n10289 & n22484 ;
  assign n22486 = ~\emc_WSCRreg_DO_reg[9]/NET0131  & ~n22484 ;
  assign n22487 = ~n22485 & ~n22486 ;
  assign n22488 = ~n10638 & n22484 ;
  assign n22489 = ~\emc_WSCRreg_DO_reg[8]/NET0131  & ~n22484 ;
  assign n22490 = ~n22488 & ~n22489 ;
  assign n22491 = ~n7340 & n22484 ;
  assign n22492 = ~\emc_WSCRreg_DO_reg[13]/NET0131  & ~n22484 ;
  assign n22493 = ~n22491 & ~n22492 ;
  assign n22494 = ~n9178 & n22484 ;
  assign n22495 = ~\emc_WSCRreg_DO_reg[12]/NET0131  & ~n22484 ;
  assign n22496 = ~n22494 & ~n22495 ;
  assign n22497 = ~n8460 & n22484 ;
  assign n22498 = ~\emc_WSCRreg_DO_reg[11]/NET0131  & ~n22484 ;
  assign n22499 = ~n22497 & ~n22498 ;
  assign n22500 = ~n7859 & n22484 ;
  assign n22501 = ~\emc_WSCRreg_DO_reg[10]/NET0131  & ~n22484 ;
  assign n22502 = ~n22500 & ~n22501 ;
  assign n22503 = ~\sice_ICYC_reg[10]/NET0131  & ~n20739 ;
  assign n22504 = ~n20740 & ~n22503 ;
  assign n22505 = ~\sice_IIRC_reg[10]/NET0131  & ~n20854 ;
  assign n22506 = ~n20855 & ~n22505 ;
  assign n22507 = \emc_PMDreg_reg[7]/P0001  & ~n14745 ;
  assign n22508 = \T_ED[7]_pad  & n14745 ;
  assign n22509 = ~n22507 & ~n22508 ;
  assign n22510 = \emc_PMDreg_reg[6]/P0001  & ~n14745 ;
  assign n22511 = \T_ED[6]_pad  & n14745 ;
  assign n22512 = ~n22510 & ~n22511 ;
  assign n22513 = \emc_PMDreg_reg[5]/P0001  & ~n14745 ;
  assign n22514 = \T_ED[5]_pad  & n14745 ;
  assign n22515 = ~n22513 & ~n22514 ;
  assign n22516 = \emc_PMDreg_reg[4]/P0001  & ~n14745 ;
  assign n22517 = \T_ED[4]_pad  & n14745 ;
  assign n22518 = ~n22516 & ~n22517 ;
  assign n22519 = \emc_PMDreg_reg[3]/P0001  & ~n14745 ;
  assign n22520 = \T_ED[3]_pad  & n14745 ;
  assign n22521 = ~n22519 & ~n22520 ;
  assign n22522 = \emc_PMDreg_reg[2]/P0001  & ~n14745 ;
  assign n22523 = \T_ED[2]_pad  & n14745 ;
  assign n22524 = ~n22522 & ~n22523 ;
  assign n22525 = \emc_PMDreg_reg[1]/P0001  & ~n14745 ;
  assign n22526 = \T_ED[1]_pad  & n14745 ;
  assign n22527 = ~n22525 & ~n22526 ;
  assign n22528 = \emc_PMDreg_reg[15]/P0001  & ~n14745 ;
  assign n22529 = \T_ED[15]_pad  & n14745 ;
  assign n22530 = ~n22528 & ~n22529 ;
  assign n22531 = \emc_PMDreg_reg[14]/P0001  & ~n14745 ;
  assign n22532 = \T_ED[14]_pad  & n14745 ;
  assign n22533 = ~n22531 & ~n22532 ;
  assign n22534 = \emc_PMDreg_reg[13]/P0001  & ~n14745 ;
  assign n22535 = \T_ED[13]_pad  & n14745 ;
  assign n22536 = ~n22534 & ~n22535 ;
  assign n22537 = \emc_PMDreg_reg[12]/P0001  & ~n14745 ;
  assign n22538 = \T_ED[12]_pad  & n14745 ;
  assign n22539 = ~n22537 & ~n22538 ;
  assign n22540 = \emc_PMDreg_reg[11]/P0001  & ~n14745 ;
  assign n22541 = \T_ED[11]_pad  & n14745 ;
  assign n22542 = ~n22540 & ~n22541 ;
  assign n22543 = \emc_PMDreg_reg[10]/P0001  & ~n14745 ;
  assign n22544 = \T_ED[10]_pad  & n14745 ;
  assign n22545 = ~n22543 & ~n22544 ;
  assign n22546 = \emc_PMDreg_reg[0]/P0001  & ~n14745 ;
  assign n22547 = \T_ED[0]_pad  & n14745 ;
  assign n22548 = ~n22546 & ~n22547 ;
  assign n22549 = ~n11265 & n22458 ;
  assign n22550 = ~\clkc_ckr_reg_DO_reg[7]/NET0131  & ~n22458 ;
  assign n22551 = ~n22549 & ~n22550 ;
  assign n22552 = ~n11525 & n22458 ;
  assign n22553 = ~\clkc_ckr_reg_DO_reg[6]/NET0131  & ~n22458 ;
  assign n22554 = ~n22552 & ~n22553 ;
  assign n22555 = ~n10911 & n22458 ;
  assign n22556 = ~\clkc_ckr_reg_DO_reg[5]/NET0131  & ~n22458 ;
  assign n22557 = ~n22555 & ~n22556 ;
  assign n22558 = ~n10069 & n22458 ;
  assign n22559 = ~\clkc_ckr_reg_DO_reg[4]/NET0131  & ~n22458 ;
  assign n22560 = ~n22558 & ~n22559 ;
  assign n22561 = ~n8113 & n22458 ;
  assign n22562 = ~\clkc_ckr_reg_DO_reg[3]/NET0131  & ~n22458 ;
  assign n22563 = ~n22561 & ~n22562 ;
  assign n22564 = ~n8715 & n22458 ;
  assign n22565 = ~\clkc_ckr_reg_DO_reg[2]/NET0131  & ~n22458 ;
  assign n22566 = ~n22564 & ~n22565 ;
  assign n22567 = ~n9435 & n22458 ;
  assign n22568 = ~\clkc_ckr_reg_DO_reg[1]/NET0131  & ~n22458 ;
  assign n22569 = ~n22567 & ~n22568 ;
  assign n22570 = ~n12743 & n22458 ;
  assign n22571 = ~\clkc_ckr_reg_DO_reg[15]/NET0131  & ~n22458 ;
  assign n22572 = ~n22570 & ~n22571 ;
  assign n22573 = ~n12688 & n22458 ;
  assign n22574 = ~\clkc_ckr_reg_DO_reg[14]/NET0131  & ~n22458 ;
  assign n22575 = ~n22573 & ~n22574 ;
  assign n22576 = ~n7607 & n22458 ;
  assign n22577 = ~\clkc_ckr_reg_DO_reg[0]/NET0131  & ~n22458 ;
  assign n22578 = ~n22576 & ~n22577 ;
  assign n22579 = ~\sice_ICYC_reg[17]/NET0131  & ~n20746 ;
  assign n22580 = ~n20747 & ~n22579 ;
  assign n22581 = \sice_IIRC_reg[15]/NET0131  & n20859 ;
  assign n22582 = \sice_IIRC_reg[16]/NET0131  & n22581 ;
  assign n22583 = ~\sice_IIRC_reg[17]/NET0131  & ~n22582 ;
  assign n22584 = \sice_IIRC_reg[17]/NET0131  & n22582 ;
  assign n22585 = ~n22583 & ~n22584 ;
  assign n22586 = ~\sice_IIRC_reg[13]/NET0131  & ~n20857 ;
  assign n22587 = ~n20858 & ~n22586 ;
  assign n22588 = ~\sice_ICYC_reg[13]/NET0131  & ~n20742 ;
  assign n22589 = ~n20743 & ~n22588 ;
  assign n22590 = ~n11265 & n22477 ;
  assign n22591 = ~\tm_tpr_reg_DO_reg[7]/NET0131  & ~n22477 ;
  assign n22592 = ~n22590 & ~n22591 ;
  assign n22593 = ~n11525 & n22477 ;
  assign n22594 = ~\tm_tpr_reg_DO_reg[6]/NET0131  & ~n22477 ;
  assign n22595 = ~n22593 & ~n22594 ;
  assign n22596 = ~n10911 & n22477 ;
  assign n22597 = ~\tm_tpr_reg_DO_reg[5]/NET0131  & ~n22477 ;
  assign n22598 = ~n22596 & ~n22597 ;
  assign n22599 = ~n8113 & n22477 ;
  assign n22600 = ~\tm_tpr_reg_DO_reg[3]/NET0131  & ~n22477 ;
  assign n22601 = ~n22599 & ~n22600 ;
  assign n22602 = ~n8715 & n22477 ;
  assign n22603 = ~\tm_tpr_reg_DO_reg[2]/NET0131  & ~n22477 ;
  assign n22604 = ~n22602 & ~n22603 ;
  assign n22605 = ~n9435 & n22477 ;
  assign n22606 = ~\tm_tpr_reg_DO_reg[1]/NET0131  & ~n22477 ;
  assign n22607 = ~n22605 & ~n22606 ;
  assign n22608 = ~n10069 & n22477 ;
  assign n22609 = ~\tm_tpr_reg_DO_reg[4]/NET0131  & ~n22477 ;
  assign n22610 = ~n22608 & ~n22609 ;
  assign n22611 = ~n12743 & n22477 ;
  assign n22612 = ~\tm_tpr_reg_DO_reg[15]/NET0131  & ~n22477 ;
  assign n22613 = ~n22611 & ~n22612 ;
  assign n22614 = ~n12688 & n22477 ;
  assign n22615 = ~\tm_tpr_reg_DO_reg[14]/NET0131  & ~n22477 ;
  assign n22616 = ~n22614 & ~n22615 ;
  assign n22617 = ~n7607 & n22477 ;
  assign n22618 = ~\tm_tpr_reg_DO_reg[0]/NET0131  & ~n22477 ;
  assign n22619 = ~n22617 & ~n22618 ;
  assign n22620 = ~n11265 & n22484 ;
  assign n22621 = ~\emc_WSCRreg_DO_reg[7]/NET0131  & ~n22484 ;
  assign n22622 = ~n22620 & ~n22621 ;
  assign n22623 = ~n11525 & n22484 ;
  assign n22624 = ~\emc_WSCRreg_DO_reg[6]/NET0131  & ~n22484 ;
  assign n22625 = ~n22623 & ~n22624 ;
  assign n22626 = ~n10911 & n22484 ;
  assign n22627 = ~\emc_WSCRreg_DO_reg[5]/NET0131  & ~n22484 ;
  assign n22628 = ~n22626 & ~n22627 ;
  assign n22629 = ~n10069 & n22484 ;
  assign n22630 = ~\emc_WSCRreg_DO_reg[4]/NET0131  & ~n22484 ;
  assign n22631 = ~n22629 & ~n22630 ;
  assign n22632 = ~n8113 & n22484 ;
  assign n22633 = ~\emc_WSCRreg_DO_reg[3]/NET0131  & ~n22484 ;
  assign n22634 = ~n22632 & ~n22633 ;
  assign n22635 = ~n8715 & n22484 ;
  assign n22636 = ~\emc_WSCRreg_DO_reg[2]/NET0131  & ~n22484 ;
  assign n22637 = ~n22635 & ~n22636 ;
  assign n22638 = ~n9435 & n22484 ;
  assign n22639 = ~\emc_WSCRreg_DO_reg[1]/NET0131  & ~n22484 ;
  assign n22640 = ~n22638 & ~n22639 ;
  assign n22641 = ~n12688 & n22484 ;
  assign n22642 = ~\emc_WSCRreg_DO_reg[14]/NET0131  & ~n22484 ;
  assign n22643 = ~n22641 & ~n22642 ;
  assign n22644 = ~n7607 & n22484 ;
  assign n22645 = ~\emc_WSCRreg_DO_reg[0]/NET0131  & ~n22484 ;
  assign n22646 = ~n22644 & ~n22645 ;
  assign n22650 = ~\sport1_regs_SCTLreg_DO_reg[11]/NET0131  & ~\sport1_regs_SCTLreg_DO_reg[12]/NET0131  ;
  assign n22651 = ~\ITFS1_pad  & \T_TFS1_pad  ;
  assign n22652 = \ITFS1_pad  & ~n13729 ;
  assign n22653 = ~n22651 & ~n22652 ;
  assign n22654 = \sport1_regs_SCTLreg_DO_reg[7]/NET0131  & ~n22653 ;
  assign n22655 = ~\sport1_regs_SCTLreg_DO_reg[7]/NET0131  & n22653 ;
  assign n22656 = ~n22654 & ~n22655 ;
  assign n22657 = \sport1_cfg_SP_ENg_reg/NET0131  & ~\sport1_cfg_TFSgi_d_reg/NET0131  ;
  assign n22658 = n22656 & n22657 ;
  assign n22659 = n22650 & ~n22658 ;
  assign n22661 = \sport1_cfg_TFSg_d3_reg/NET0131  & \sport1_regs_SCTLreg_DO_reg[11]/NET0131  ;
  assign n22660 = \sport1_cfg_TFSg_d2_reg/NET0131  & ~\sport1_regs_SCTLreg_DO_reg[11]/NET0131  ;
  assign n22662 = \sport1_regs_SCTLreg_DO_reg[12]/NET0131  & ~n22660 ;
  assign n22663 = ~n22661 & n22662 ;
  assign n22648 = ~\sport1_cfg_TFSg_d1_reg/NET0131  & \sport1_regs_SCTLreg_DO_reg[11]/NET0131  ;
  assign n22649 = ~\sport1_regs_SCTLreg_DO_reg[12]/NET0131  & n22648 ;
  assign n22664 = \sport1_txctl_TCS_reg[0]/NET0131  & ~n22649 ;
  assign n22665 = ~n22663 & n22664 ;
  assign n22666 = ~n22659 & n22665 ;
  assign n22667 = ~\sport1_txctl_TCS_reg[2]/NET0131  & ~n22666 ;
  assign n22647 = \sport1_txctl_TCS_reg[0]/NET0131  & \sport1_txctl_TCS_reg[2]/NET0131  ;
  assign n22668 = ~\sport1_txctl_TCS_reg[1]/NET0131  & ~n22647 ;
  assign n22669 = ~n22667 & n22668 ;
  assign n22670 = ~\sport1_txctl_TCS_reg[0]/NET0131  & \sport1_txctl_TCS_reg[1]/NET0131  ;
  assign n22671 = ~\sport1_txctl_TCS_reg[2]/NET0131  & n22670 ;
  assign n22672 = ~\sport1_txctl_Bcnt_reg[0]/NET0131  & ~\sport1_txctl_Bcnt_reg[1]/NET0131  ;
  assign n22673 = ~\sport1_txctl_Bcnt_reg[2]/NET0131  & n22672 ;
  assign n22674 = ~\sport1_txctl_Bcnt_reg[3]/NET0131  & n22673 ;
  assign n22675 = ~\sport1_txctl_Bcnt_reg[4]/NET0131  & n22674 ;
  assign n22676 = n22671 & ~n22675 ;
  assign n22677 = ~n22669 & ~n22676 ;
  assign n22678 = \sport1_txctl_TXSHT_reg[9]/P0001  & ~n22677 ;
  assign n22679 = \sport1_txctl_TX_reg[10]/P0001  & n22677 ;
  assign n22680 = ~n22678 & ~n22679 ;
  assign n22683 = n18271 & ~n20080 ;
  assign n22682 = ~\core_eu_em_mac_em_reg_mr0swe_DO_reg[4]/P0001  & ~n18271 ;
  assign n22684 = n18273 & ~n22682 ;
  assign n22685 = ~n22683 & n22684 ;
  assign n22681 = \core_eu_em_mac_em_reg_mr0swe_DO_reg[4]/P0001  & ~n18266 ;
  assign n22686 = ~n18270 & ~n22681 ;
  assign n22687 = ~n22685 & n22686 ;
  assign n22688 = ~n18262 & ~n22687 ;
  assign n22689 = n18262 & ~n19670 ;
  assign n22690 = ~n22688 & ~n22689 ;
  assign n22691 = n14752 & n19670 ;
  assign n22692 = n18328 & n20080 ;
  assign n22693 = \core_eu_em_mac_em_reg_mr0rwe_DO_reg[4]/P0001  & ~n18330 ;
  assign n22694 = n18334 & ~n22693 ;
  assign n22695 = ~n22692 & n22694 ;
  assign n22696 = ~n22691 & ~n22695 ;
  assign n22698 = \sport0_txctl_ldTX_cmp_reg/P0001  & n18514 ;
  assign n22697 = \sport0_txctl_TX_reg[6]/P0001  & n21318 ;
  assign n22699 = n11525 & n21316 ;
  assign n22700 = ~n22697 & ~n22699 ;
  assign n22701 = ~n22698 & n22700 ;
  assign n22702 = ~n15120 & ~n15183 ;
  assign n22703 = ~n15319 & n22702 ;
  assign n22704 = ~n17777 & n22703 ;
  assign n22706 = ~n17783 & n22702 ;
  assign n22705 = ~n15120 & n15182 ;
  assign n22707 = ~n15121 & ~n22705 ;
  assign n22708 = ~n22706 & n22707 ;
  assign n22709 = ~n22704 & n22708 ;
  assign n22710 = ~n14933 & ~n15053 ;
  assign n22711 = ~n9865 & n14993 ;
  assign n22712 = \core_c_psq_MSTAT_reg_DO_reg[4]/NET0131  & n15046 ;
  assign n22713 = ~n22711 & ~n22712 ;
  assign n22714 = ~\core_eu_em_mac_em_dec_emcorepi_DO_reg[1]/P0001  & ~n22713 ;
  assign n22715 = ~n14972 & n22714 ;
  assign n22716 = n14972 & ~n22714 ;
  assign n22717 = ~n22715 & ~n22716 ;
  assign n22718 = ~n15051 & ~n22717 ;
  assign n22719 = n15051 & n22713 ;
  assign n22720 = ~n22718 & ~n22719 ;
  assign n22721 = n14992 & ~n22720 ;
  assign n22722 = ~n14992 & n22720 ;
  assign n22723 = ~n22721 & ~n22722 ;
  assign n22724 = ~n22710 & ~n22723 ;
  assign n22725 = n22710 & n22723 ;
  assign n22726 = ~n22724 & ~n22725 ;
  assign n22727 = ~n14991 & ~n15054 ;
  assign n22728 = n15058 & n22727 ;
  assign n22729 = ~n15059 & ~n22728 ;
  assign n22730 = n22726 & ~n22729 ;
  assign n22731 = ~n14853 & ~n22730 ;
  assign n22732 = ~n14933 & ~n22718 ;
  assign n22733 = ~n10882 & n14993 ;
  assign n22734 = ~n9865 & n15044 ;
  assign n22735 = ~n22733 & ~n22734 ;
  assign n22736 = ~\core_eu_em_mac_em_dec_emcorepi_DO_reg[1]/P0001  & ~n22735 ;
  assign n22737 = ~n14972 & n22736 ;
  assign n22738 = n14972 & ~n22736 ;
  assign n22739 = ~n22737 & ~n22738 ;
  assign n22740 = ~n22715 & ~n22739 ;
  assign n22741 = n22715 & n22735 ;
  assign n22742 = ~n22740 & ~n22741 ;
  assign n22743 = n14992 & ~n22742 ;
  assign n22744 = ~n14992 & n22742 ;
  assign n22745 = ~n22743 & ~n22744 ;
  assign n22746 = n22732 & ~n22745 ;
  assign n22747 = ~n22732 & n22745 ;
  assign n22748 = ~n22746 & ~n22747 ;
  assign n22749 = ~n14991 & ~n22719 ;
  assign n22750 = n22723 & n22749 ;
  assign n22751 = ~n22724 & ~n22750 ;
  assign n22752 = ~n22748 & ~n22751 ;
  assign n22753 = n22748 & n22751 ;
  assign n22754 = ~n22752 & ~n22753 ;
  assign n22755 = n14853 & n22754 ;
  assign n22756 = ~n14853 & ~n22754 ;
  assign n22757 = ~n22755 & ~n22756 ;
  assign n22758 = ~n22731 & ~n22757 ;
  assign n22759 = n22731 & n22754 ;
  assign n22760 = ~n22758 & ~n22759 ;
  assign n22761 = ~n14853 & n15065 ;
  assign n22762 = ~n22726 & n22729 ;
  assign n22763 = ~n22730 & ~n22762 ;
  assign n22764 = n22761 & n22763 ;
  assign n22765 = ~n22761 & ~n22763 ;
  assign n22766 = ~n22764 & ~n22765 ;
  assign n22767 = ~n22760 & n22766 ;
  assign n22768 = n14853 & ~n22729 ;
  assign n22769 = n22765 & ~n22768 ;
  assign n22770 = n22760 & ~n22769 ;
  assign n22771 = ~n15066 & ~n15070 ;
  assign n22772 = ~n15071 & ~n22771 ;
  assign n22773 = ~n22770 & n22772 ;
  assign n22774 = ~n22767 & ~n22773 ;
  assign n22775 = ~n22709 & ~n22774 ;
  assign n22776 = ~n22760 & n22769 ;
  assign n22777 = n22767 & n22772 ;
  assign n22778 = ~n22776 & ~n22777 ;
  assign n22779 = ~n22775 & n22778 ;
  assign n22780 = ~n14853 & ~n22752 ;
  assign n22781 = ~n14933 & ~n22740 ;
  assign n22782 = ~n11424 & n14993 ;
  assign n22783 = ~n10882 & n15044 ;
  assign n22784 = ~n22782 & ~n22783 ;
  assign n22785 = ~\core_eu_em_mac_em_dec_emcorepi_DO_reg[1]/P0001  & ~n22784 ;
  assign n22786 = ~n14972 & n22785 ;
  assign n22787 = n14972 & ~n22785 ;
  assign n22788 = ~n22786 & ~n22787 ;
  assign n22789 = ~n22737 & ~n22788 ;
  assign n22790 = n22737 & n22784 ;
  assign n22791 = ~n22789 & ~n22790 ;
  assign n22792 = n14992 & ~n22791 ;
  assign n22793 = ~n14992 & n22791 ;
  assign n22794 = ~n22792 & ~n22793 ;
  assign n22795 = n22781 & ~n22794 ;
  assign n22796 = ~n22781 & n22794 ;
  assign n22797 = ~n22795 & ~n22796 ;
  assign n22798 = ~n14991 & ~n22741 ;
  assign n22799 = n22745 & ~n22798 ;
  assign n22800 = ~n22746 & ~n22799 ;
  assign n22801 = ~n22797 & n22800 ;
  assign n22802 = n22797 & ~n22800 ;
  assign n22803 = ~n22801 & ~n22802 ;
  assign n22804 = n14853 & n22803 ;
  assign n22805 = ~n14853 & ~n22803 ;
  assign n22806 = ~n22804 & ~n22805 ;
  assign n22807 = ~n22780 & ~n22806 ;
  assign n22808 = ~n22802 & n22806 ;
  assign n22809 = ~n22807 & ~n22808 ;
  assign n22810 = ~n14933 & ~n22789 ;
  assign n22811 = ~n7206 & n14993 ;
  assign n22812 = ~n11424 & n15044 ;
  assign n22813 = ~n22811 & ~n22812 ;
  assign n22814 = ~\core_eu_em_mac_em_dec_emcorepi_DO_reg[1]/P0001  & ~n22813 ;
  assign n22816 = n14972 & n22814 ;
  assign n22815 = ~n14972 & ~n22814 ;
  assign n22817 = ~n22786 & ~n22815 ;
  assign n22818 = ~n22816 & n22817 ;
  assign n22819 = n22786 & ~n22814 ;
  assign n22820 = ~n22818 & ~n22819 ;
  assign n22821 = n14992 & ~n22820 ;
  assign n22822 = ~n14992 & n22820 ;
  assign n22823 = ~n22821 & ~n22822 ;
  assign n22824 = ~n22810 & n22823 ;
  assign n22825 = n22810 & ~n22823 ;
  assign n22826 = ~n22824 & ~n22825 ;
  assign n22827 = ~n14991 & ~n22790 ;
  assign n22828 = n22794 & ~n22827 ;
  assign n22829 = ~n22795 & ~n22828 ;
  assign n22830 = ~n22826 & n22829 ;
  assign n22831 = n22826 & ~n22829 ;
  assign n22832 = ~n22830 & ~n22831 ;
  assign n22833 = ~n14853 & n22801 ;
  assign n22834 = ~n22832 & n22833 ;
  assign n22835 = n22832 & ~n22833 ;
  assign n22836 = ~n22834 & ~n22835 ;
  assign n22837 = ~n22809 & n22836 ;
  assign n22838 = ~n22753 & n22757 ;
  assign n22839 = ~n22758 & ~n22838 ;
  assign n22840 = n22780 & n22803 ;
  assign n22841 = ~n22807 & ~n22840 ;
  assign n22842 = ~n22839 & n22841 ;
  assign n22843 = ~n22837 & ~n22842 ;
  assign n22844 = ~n22779 & n22843 ;
  assign n22845 = n22809 & ~n22836 ;
  assign n22846 = n22839 & ~n22841 ;
  assign n22847 = ~n22837 & n22846 ;
  assign n22848 = ~n22845 & ~n22847 ;
  assign n22849 = ~n22844 & n22848 ;
  assign n22850 = ~n7206 & n17443 ;
  assign n22851 = ~n14991 & ~n22819 ;
  assign n22852 = n22823 & ~n22851 ;
  assign n22853 = ~n22825 & ~n22852 ;
  assign n22854 = n22815 & ~n22853 ;
  assign n22855 = ~n22815 & n22853 ;
  assign n22856 = ~n22854 & ~n22855 ;
  assign n22857 = n22850 & n22856 ;
  assign n22858 = ~n22850 & ~n22856 ;
  assign n22859 = ~n22857 & ~n22858 ;
  assign n22860 = ~n22830 & n22833 ;
  assign n22861 = ~n22831 & ~n22833 ;
  assign n22862 = ~n22860 & ~n22861 ;
  assign n22863 = n22859 & ~n22862 ;
  assign n22864 = ~n22859 & n22862 ;
  assign n22865 = ~n22863 & ~n22864 ;
  assign n22866 = ~n14991 & ~n22818 ;
  assign n22867 = ~n14992 & n22818 ;
  assign n22868 = ~n22866 & ~n22867 ;
  assign n22869 = n22865 & ~n22868 ;
  assign n22870 = ~n22865 & n22868 ;
  assign n22871 = ~n22869 & ~n22870 ;
  assign n22872 = n22849 & n22871 ;
  assign n22873 = ~n22849 & ~n22871 ;
  assign n22874 = ~n22872 & ~n22873 ;
  assign n22875 = \core_c_psq_MSTAT_reg_DO_reg[4]/NET0131  & ~n22874 ;
  assign n22876 = ~n22837 & ~n22845 ;
  assign n22877 = ~n22779 & ~n22842 ;
  assign n22878 = ~n22846 & ~n22877 ;
  assign n22879 = n22876 & ~n22878 ;
  assign n22880 = ~n22876 & n22878 ;
  assign n22881 = ~n22879 & ~n22880 ;
  assign n22882 = ~\core_c_psq_MSTAT_reg_DO_reg[4]/NET0131  & n22881 ;
  assign n22883 = ~n22875 & ~n22882 ;
  assign n22884 = \core_c_dec_MTSR0_E_reg/P0001  & ~n20080 ;
  assign n22896 = ~n17998 & n18183 ;
  assign n22894 = n17925 & ~n18888 ;
  assign n22895 = ~n17938 & n18083 ;
  assign n22906 = ~n22894 & ~n22895 ;
  assign n22907 = ~n22896 & n22906 ;
  assign n22897 = n17991 & n18765 ;
  assign n22891 = n18746 & ~n18918 ;
  assign n22893 = ~n18743 & ~n18912 ;
  assign n22902 = ~n22891 & ~n22893 ;
  assign n22903 = ~n22897 & n22902 ;
  assign n22886 = n18752 & ~n18907 ;
  assign n22887 = ~n18914 & ~n18919 ;
  assign n22900 = ~n22886 & ~n22887 ;
  assign n22889 = n18763 & ~n18918 ;
  assign n22890 = ~n18079 & ~n19864 ;
  assign n22901 = ~n22889 & ~n22890 ;
  assign n22904 = n22900 & n22901 ;
  assign n22892 = n18758 & ~n18898 ;
  assign n22885 = ~n18909 & ~n19870 ;
  assign n22888 = \core_c_dec_IRE_reg[11]/NET0131  & ~n9951 ;
  assign n22898 = ~n20272 & ~n22888 ;
  assign n22899 = ~n22885 & n22898 ;
  assign n22905 = ~n22892 & n22899 ;
  assign n22908 = n22904 & n22905 ;
  assign n22909 = n22903 & n22908 ;
  assign n22910 = n22907 & n22909 ;
  assign n22911 = n20274 & n22910 ;
  assign n22912 = ~\core_c_dec_MTSR0_E_reg/P0001  & n22911 ;
  assign n22913 = ~n22884 & ~n22912 ;
  assign n22914 = n18886 & ~n22913 ;
  assign n22915 = ~\core_eu_es_sht_es_reg_sr0swe_DO_reg[4]/P0001  & ~n18886 ;
  assign n22916 = ~n22914 & ~n22915 ;
  assign n22917 = n19034 & ~n22913 ;
  assign n22918 = ~\core_eu_es_sht_es_reg_sr0rwe_DO_reg[4]/P0001  & ~n19034 ;
  assign n22919 = ~n22917 & ~n22918 ;
  assign n22920 = \core_c_psq_MSTAT_reg_DO_reg[4]/NET0131  & n22881 ;
  assign n22921 = ~n22842 & ~n22846 ;
  assign n22922 = ~n22779 & n22921 ;
  assign n22923 = n22779 & ~n22921 ;
  assign n22924 = ~n22922 & ~n22923 ;
  assign n22925 = ~\core_c_psq_MSTAT_reg_DO_reg[4]/NET0131  & n22924 ;
  assign n22926 = ~n22920 & ~n22925 ;
  assign n22927 = \core_eu_em_mac_em_reg_mrovfwe_DO_reg[0]/P0001  & ~n21314 ;
  assign n22928 = ~n19379 & n21314 ;
  assign n22929 = ~n22927 & ~n22928 ;
  assign n22930 = \core_c_dec_satMR_E_reg/P0001  & n4117 ;
  assign n22931 = n19696 & n21557 ;
  assign n22932 = ~n22930 & ~n22931 ;
  assign n22933 = n4116 & ~n22932 ;
  assign n22934 = \core_c_dec_DIVS_E_reg/P0001  & n4117 ;
  assign n22935 = ~n21558 & ~n22934 ;
  assign n22936 = n4116 & ~n22935 ;
  assign n22938 = n19499 & ~n19972 ;
  assign n22937 = ~\core_eu_em_mac_em_reg_mr1swe_DO_reg[7]/P0001  & ~n19499 ;
  assign n22939 = n19501 & ~n22937 ;
  assign n22940 = ~n22938 & n22939 ;
  assign n22941 = \core_eu_em_mac_em_reg_mr1swe_DO_reg[7]/P0001  & ~n19383 ;
  assign n22942 = ~n19508 & ~n22941 ;
  assign n22943 = ~n22940 & n22942 ;
  assign n22944 = ~n18262 & ~n22943 ;
  assign n22945 = ~n16979 & ~n17688 ;
  assign n22946 = ~n19424 & n22945 ;
  assign n22947 = n19424 & ~n22945 ;
  assign n22948 = ~n22946 & ~n22947 ;
  assign n22949 = \core_c_psq_MSTAT_reg_DO_reg[4]/NET0131  & ~n22948 ;
  assign n22950 = n17544 & ~n19422 ;
  assign n22951 = ~n17679 & ~n22950 ;
  assign n22952 = ~n17559 & ~n22951 ;
  assign n22953 = ~n17682 & ~n22952 ;
  assign n22954 = ~n17565 & ~n17681 ;
  assign n22955 = n22953 & n22954 ;
  assign n22956 = ~n22953 & ~n22954 ;
  assign n22957 = ~n22955 & ~n22956 ;
  assign n22958 = ~\core_c_psq_MSTAT_reg_DO_reg[4]/NET0131  & n22957 ;
  assign n22959 = ~n22949 & ~n22958 ;
  assign n22960 = n18262 & n22959 ;
  assign n22961 = ~n22944 & ~n22960 ;
  assign n22962 = n7340 & n20401 ;
  assign n22964 = \core_c_psq_lpstk_lps4x22_LPcell_reg[0][3]/P0001  & n4845 ;
  assign n22965 = \core_c_psq_lpstk_lps4x22_LPcell_reg[1][3]/P0001  & n4847 ;
  assign n22968 = ~n22964 & ~n22965 ;
  assign n22966 = \core_c_psq_lpstk_lps4x22_LPcell_reg[2][3]/P0001  & n4851 ;
  assign n22967 = \core_c_psq_lpstk_lps4x22_LPcell_reg[3][3]/P0001  & n4849 ;
  assign n22969 = ~n22966 & ~n22967 ;
  assign n22970 = n22968 & n22969 ;
  assign n22971 = ~n4117 & n22970 ;
  assign n22963 = ~\core_eu_ec_cun_TERM_E_reg[3]/P0001  & n4117 ;
  assign n22972 = n4150 & ~n22963 ;
  assign n22973 = ~n22971 & n22972 ;
  assign n22975 = \core_c_psq_lpstk_lps4x22_LPcell_reg[0][2]/P0001  & n4845 ;
  assign n22976 = \core_c_psq_lpstk_lps4x22_LPcell_reg[1][2]/P0001  & n4847 ;
  assign n22979 = ~n22975 & ~n22976 ;
  assign n22977 = \core_c_psq_lpstk_lps4x22_LPcell_reg[2][2]/P0001  & n4851 ;
  assign n22978 = \core_c_psq_lpstk_lps4x22_LPcell_reg[3][2]/P0001  & n4849 ;
  assign n22980 = ~n22977 & ~n22978 ;
  assign n22981 = n22979 & n22980 ;
  assign n22982 = ~n4117 & n22981 ;
  assign n22974 = ~\core_eu_ec_cun_TERM_E_reg[2]/P0001  & n4117 ;
  assign n22983 = n4150 & ~n22974 ;
  assign n22984 = ~n22982 & n22983 ;
  assign n22986 = n19499 & ~n20150 ;
  assign n22985 = ~\core_eu_em_mac_em_reg_mr1swe_DO_reg[14]/P0001  & ~n19499 ;
  assign n22987 = n19501 & ~n22985 ;
  assign n22988 = ~n22986 & n22987 ;
  assign n22989 = \core_eu_em_mac_em_reg_mr1swe_DO_reg[14]/P0001  & ~n19383 ;
  assign n22990 = ~n19508 & ~n22989 ;
  assign n22991 = ~n22988 & n22990 ;
  assign n22992 = ~n18262 & ~n22991 ;
  assign n22993 = ~n17759 & ~n17768 ;
  assign n22994 = ~n19372 & n22993 ;
  assign n22995 = n19372 & ~n22993 ;
  assign n22996 = ~n22994 & ~n22995 ;
  assign n22997 = ~\core_c_psq_MSTAT_reg_DO_reg[4]/NET0131  & n22996 ;
  assign n22998 = \core_c_psq_MSTAT_reg_DO_reg[4]/NET0131  & n19377 ;
  assign n22999 = ~n22997 & ~n22998 ;
  assign n23000 = n18262 & ~n22999 ;
  assign n23001 = ~n22992 & ~n23000 ;
  assign n23002 = \core_c_dec_BR_Ed_reg/P0001  & n4117 ;
  assign n23003 = ~n21257 & ~n23002 ;
  assign n23004 = n4116 & ~n23003 ;
  assign n23005 = \core_c_dec_imSHT_E_reg/P0001  & n4117 ;
  assign n23006 = n6119 & n21559 ;
  assign n23007 = ~n23005 & ~n23006 ;
  assign n23008 = n4116 & ~n23007 ;
  assign n23009 = \core_c_dec_Stkctl_Eg_reg/P0001  & n4117 ;
  assign n23010 = ~n21251 & ~n23009 ;
  assign n23011 = n4116 & ~n23010 ;
  assign n23012 = n14752 & ~n22959 ;
  assign n23013 = n19776 & n19972 ;
  assign n23014 = \core_eu_em_mac_em_reg_mr1rwe_DO_reg[7]/P0001  & ~n17809 ;
  assign n23015 = n19780 & ~n23014 ;
  assign n23016 = ~n23013 & n23015 ;
  assign n23017 = ~n23012 & ~n23016 ;
  assign n23020 = \clkc_CTR_cnt_reg[0]/NET0131  & \clkc_CTR_cnt_reg[1]/NET0131  ;
  assign n23021 = ~\clkc_RSTtext_reg/P0001  & n23020 ;
  assign n23018 = ~\sice_GOICE_1_reg/NET0131  & ~\sice_GOICE_2_reg/NET0131  ;
  assign n23019 = ~\sice_GOICE_s1_reg/NET0131  & ~n23018 ;
  assign n23022 = n4149 & ~n23019 ;
  assign n23023 = n23021 & n23022 ;
  assign n23024 = ~\bdma_BWcnt_reg[2]/NET0131  & ~n20038 ;
  assign n23025 = ~n20039 & ~n23024 ;
  assign n23026 = ~n13750 & n23025 ;
  assign n23027 = \sice_IAR_reg[0]/NET0131  & ~\sice_IAR_reg[3]/NET0131  ;
  assign n23028 = ~\sice_IAR_reg[1]/NET0131  & ~\sice_IAR_reg[2]/NET0131  ;
  assign n23029 = n23027 & n23028 ;
  assign n23030 = T_IMS_pad & ~\sice_ICS_reg[1]/NET0131  ;
  assign n23031 = \sice_ICS_reg[0]/NET0131  & \sice_ICS_reg[2]/NET0131  ;
  assign n23032 = n23030 & n23031 ;
  assign n23033 = n23029 & n23032 ;
  assign n23034 = ~\sice_IRST_reg/NET0131  & \sice_SPC_reg[18]/P0001  ;
  assign n23035 = n23033 & n23034 ;
  assign n23036 = ~\sice_CLR_I_reg/NET0131  & \sice_SPC_reg[21]/P0001  ;
  assign n23037 = n23033 & n23036 ;
  assign n23044 = n18500 & n18507 ;
  assign n23045 = \sport0_regs_SCTLreg_DO_reg[4]/NET0131  & ~n18492 ;
  assign n23046 = n23044 & n23045 ;
  assign n23047 = n18514 & n23046 ;
  assign n23049 = n18500 & n18512 ;
  assign n23050 = ~n18507 & ~n23049 ;
  assign n23053 = n18507 & n18514 ;
  assign n23061 = n18501 & n23053 ;
  assign n23054 = ~n18500 & n23053 ;
  assign n23055 = ~n18396 & n18400 ;
  assign n23056 = ~n18401 & ~n23055 ;
  assign n23057 = \sport0_regs_SCTLreg_DO_reg[4]/NET0131  & n23056 ;
  assign n23039 = ~n18401 & n18405 ;
  assign n23040 = ~n18406 & ~n23039 ;
  assign n23058 = ~\sport0_regs_SCTLreg_DO_reg[4]/NET0131  & n23040 ;
  assign n23059 = ~n23057 & ~n23058 ;
  assign n23060 = n18457 & ~n23059 ;
  assign n23062 = ~n23054 & n23060 ;
  assign n23063 = ~n23061 & n23062 ;
  assign n23038 = ~\sport0_regs_SCTLreg_DO_reg[4]/NET0131  & n18489 ;
  assign n23041 = \sport0_regs_SCTLreg_DO_reg[4]/NET0131  & n23040 ;
  assign n23042 = ~n23038 & ~n23041 ;
  assign n23064 = n18500 & n23042 ;
  assign n23065 = n18492 & ~n23064 ;
  assign n23066 = n23053 & n23065 ;
  assign n23067 = ~n23063 & ~n23066 ;
  assign n23051 = n18480 & ~n18512 ;
  assign n23052 = ~n18507 & n18514 ;
  assign n23068 = ~n23051 & ~n23052 ;
  assign n23069 = ~n23067 & n23068 ;
  assign n23070 = ~n23050 & ~n23069 ;
  assign n23071 = n18479 & ~n23070 ;
  assign n23072 = n18471 & ~n23071 ;
  assign n23073 = ~n18481 & ~n23072 ;
  assign n23074 = n18479 & ~n23073 ;
  assign n23075 = n18512 & n23072 ;
  assign n23076 = ~n23074 & ~n23075 ;
  assign n23077 = ~n23047 & ~n23076 ;
  assign n23043 = n18457 & ~n23042 ;
  assign n23048 = ~n23043 & n23047 ;
  assign n23078 = n18467 & ~n18470 ;
  assign n23079 = ~n23048 & ~n23078 ;
  assign n23080 = ~n23077 & n23079 ;
  assign n23081 = ~\sport0_regs_SCTLreg_DO_reg[4]/NET0131  & ~n23080 ;
  assign n23082 = \sport0_regs_SCTLreg_DO_reg[4]/NET0131  & n23080 ;
  assign n23083 = ~n23081 & ~n23082 ;
  assign n23084 = \sport0_txctl_ldTX_cmp_reg/P0001  & ~n23083 ;
  assign n23085 = ~\sport0_txctl_ldTX_cmp_reg/P0001  & n8113 ;
  assign n23086 = ~n23084 & ~n23085 ;
  assign n23087 = ~n21318 & ~n23086 ;
  assign n23088 = \sport0_txctl_TX_reg[3]/P0001  & n21318 ;
  assign n23089 = ~n23087 & ~n23088 ;
  assign n23090 = ~\sice_CLR_M_reg/NET0131  & \sice_SPC_reg[22]/P0001  ;
  assign n23091 = n23033 & n23090 ;
  assign n23092 = \clkc_OSCoff_set_reg/P0001  & \clkc_SLEEP_reg/NET0131  ;
  assign n23093 = ~\clkc_OSCoff_reg/NET0131  & ~n23092 ;
  assign n23102 = \pio_PINT_reg[5]/NET0131  & \pio_pmask_reg_DO_reg[5]/NET0131  ;
  assign n23103 = \pio_PINT_reg[11]/NET0131  & \pio_pmask_reg_DO_reg[11]/NET0131  ;
  assign n23110 = ~n23102 & ~n23103 ;
  assign n23104 = \pio_PINT_reg[2]/NET0131  & \pio_pmask_reg_DO_reg[2]/NET0131  ;
  assign n23105 = \pio_PINT_reg[9]/NET0131  & \pio_pmask_reg_DO_reg[9]/NET0131  ;
  assign n23111 = ~n23104 & ~n23105 ;
  assign n23112 = n23110 & n23111 ;
  assign n23098 = \pio_PINT_reg[6]/NET0131  & \pio_pmask_reg_DO_reg[6]/NET0131  ;
  assign n23099 = \pio_PINT_reg[10]/NET0131  & \pio_pmask_reg_DO_reg[10]/NET0131  ;
  assign n23108 = ~n23098 & ~n23099 ;
  assign n23100 = \pio_PINT_reg[4]/NET0131  & \pio_pmask_reg_DO_reg[4]/NET0131  ;
  assign n23101 = \pio_PINT_reg[0]/NET0131  & \pio_pmask_reg_DO_reg[0]/NET0131  ;
  assign n23109 = ~n23100 & ~n23101 ;
  assign n23113 = n23108 & n23109 ;
  assign n23094 = \pio_PINT_reg[3]/NET0131  & \pio_pmask_reg_DO_reg[3]/NET0131  ;
  assign n23095 = \pio_PINT_reg[8]/NET0131  & \pio_pmask_reg_DO_reg[8]/NET0131  ;
  assign n23106 = ~n23094 & ~n23095 ;
  assign n23096 = \pio_PINT_reg[7]/NET0131  & \pio_pmask_reg_DO_reg[7]/NET0131  ;
  assign n23097 = \pio_PINT_reg[1]/NET0131  & \pio_pmask_reg_DO_reg[1]/NET0131  ;
  assign n23107 = ~n23096 & ~n23097 ;
  assign n23114 = n23106 & n23107 ;
  assign n23115 = n23113 & n23114 ;
  assign n23116 = n23112 & n23115 ;
  assign n23117 = n4149 & ~n20357 ;
  assign n23118 = ~\tm_WR_TCR_KEEP_TO_TMCLK_p_reg/NET0131  & ~\tm_WR_TCR_p_reg/P0001  ;
  assign n23119 = n14752 & n22999 ;
  assign n23120 = n19776 & n20150 ;
  assign n23121 = \core_eu_em_mac_em_reg_mr1rwe_DO_reg[14]/P0001  & ~n17809 ;
  assign n23122 = n19780 & ~n23121 ;
  assign n23123 = ~n23120 & n23122 ;
  assign n23124 = ~n23119 & ~n23123 ;
  assign n23126 = \core_c_psq_lpstk_lps4x22_LPcell_reg[3][1]/P0001  & n4849 ;
  assign n23127 = \core_c_psq_lpstk_lps4x22_LPcell_reg[2][1]/P0001  & n4851 ;
  assign n23130 = ~n23126 & ~n23127 ;
  assign n23128 = \core_c_psq_lpstk_lps4x22_LPcell_reg[1][1]/P0001  & n4847 ;
  assign n23129 = \core_c_psq_lpstk_lps4x22_LPcell_reg[0][1]/P0001  & n4845 ;
  assign n23131 = ~n23128 & ~n23129 ;
  assign n23132 = n23130 & n23131 ;
  assign n23133 = ~n4117 & n23132 ;
  assign n23125 = ~\core_eu_ec_cun_TERM_E_reg[1]/P0001  & n4117 ;
  assign n23134 = n4150 & ~n23125 ;
  assign n23135 = ~n23133 & n23134 ;
  assign n23137 = \core_c_psq_lpstk_lps4x22_LPcell_reg[0][0]/P0001  & n4845 ;
  assign n23138 = \core_c_psq_lpstk_lps4x22_LPcell_reg[1][0]/P0001  & n4847 ;
  assign n23141 = ~n23137 & ~n23138 ;
  assign n23139 = \core_c_psq_lpstk_lps4x22_LPcell_reg[2][0]/P0001  & n4851 ;
  assign n23140 = \core_c_psq_lpstk_lps4x22_LPcell_reg[3][0]/P0001  & n4849 ;
  assign n23142 = ~n23139 & ~n23140 ;
  assign n23143 = n23141 & n23142 ;
  assign n23144 = ~n4117 & n23143 ;
  assign n23136 = ~\core_eu_ec_cun_TERM_E_reg[0]/P0001  & n4117 ;
  assign n23145 = n4150 & ~n23136 ;
  assign n23146 = ~n23144 & n23145 ;
  assign n23152 = n18481 & n18507 ;
  assign n23157 = \sport0_regs_SCTLreg_DO_reg[4]/NET0131  & n18390 ;
  assign n23158 = ~n18392 & n18395 ;
  assign n23159 = ~n18396 & ~n23158 ;
  assign n23160 = ~\sport0_regs_SCTLreg_DO_reg[4]/NET0131  & ~n23159 ;
  assign n23161 = ~n23157 & ~n23160 ;
  assign n23162 = n18457 & n23161 ;
  assign n23163 = ~n23061 & ~n23162 ;
  assign n23147 = \sport0_regs_SCTLreg_DO_reg[4]/NET0131  & ~n18395 ;
  assign n23148 = ~\sport0_regs_SCTLreg_DO_reg[4]/NET0131  & n23056 ;
  assign n23149 = ~n23147 & ~n23148 ;
  assign n23150 = n18457 & ~n23149 ;
  assign n23164 = n23061 & ~n23150 ;
  assign n23165 = ~n23163 & ~n23164 ;
  assign n23166 = ~n23054 & ~n23165 ;
  assign n23156 = n23054 & ~n23060 ;
  assign n23167 = ~n23052 & ~n23156 ;
  assign n23168 = ~n23166 & n23167 ;
  assign n23155 = n23043 & n23052 ;
  assign n23169 = ~n23051 & ~n23155 ;
  assign n23170 = ~n23168 & n23169 ;
  assign n23154 = ~n18492 & n23051 ;
  assign n23171 = n18479 & ~n23154 ;
  assign n23172 = ~n23170 & n23171 ;
  assign n23153 = ~n18479 & ~n18500 ;
  assign n23173 = n18471 & ~n23153 ;
  assign n23174 = ~n23172 & n23173 ;
  assign n23175 = ~n23152 & ~n23174 ;
  assign n23176 = ~n23047 & ~n23175 ;
  assign n23151 = n23047 & ~n23150 ;
  assign n23177 = ~n18470 & n18512 ;
  assign n23178 = ~n23151 & ~n23177 ;
  assign n23179 = ~n23176 & n23178 ;
  assign n23180 = ~\sport0_regs_SCTLreg_DO_reg[4]/NET0131  & ~n23179 ;
  assign n23181 = \sport0_regs_SCTLreg_DO_reg[4]/NET0131  & n23179 ;
  assign n23182 = ~n23180 & ~n23181 ;
  assign n23183 = \sport0_txctl_ldTX_cmp_reg/P0001  & ~n23182 ;
  assign n23184 = ~\sport0_txctl_ldTX_cmp_reg/P0001  & n9435 ;
  assign n23185 = ~n23183 & ~n23184 ;
  assign n23186 = ~n21318 & ~n23185 ;
  assign n23187 = \sport0_txctl_TX_reg[1]/P0001  & n21318 ;
  assign n23188 = ~n23186 & ~n23187 ;
  assign n23191 = ~\sport0_rxctl_ldRX_cmp_reg/P0001  & n8113 ;
  assign n23192 = ~n20903 & ~n20921 ;
  assign n23193 = ~n20922 & ~n23192 ;
  assign n23194 = ~\sport0_rxctl_RX_reg[7]/P0001  & ~n20955 ;
  assign n23196 = ~n23193 & n23194 ;
  assign n23195 = n23193 & ~n23194 ;
  assign n23197 = n20875 & ~n23195 ;
  assign n23198 = ~n23196 & n23197 ;
  assign n23190 = \sport0_rxctl_RX_reg[3]/P0001  & n20873 ;
  assign n23199 = ~n20868 & ~n23190 ;
  assign n23200 = ~n23198 & n23199 ;
  assign n23201 = ~n23191 & n23200 ;
  assign n23189 = ~\sport0_rxctl_RXSHT_reg[3]/P0001  & n20868 ;
  assign n23202 = ~n20871 & ~n23189 ;
  assign n23203 = ~n23201 & n23202 ;
  assign n23204 = \sport0_rxctl_RX_reg[3]/P0001  & n20871 ;
  assign n23205 = ~n23203 & ~n23204 ;
  assign n23207 = ~n18276 & n19499 ;
  assign n23206 = ~\core_eu_em_mac_em_reg_mr1swe_DO_reg[6]/P0001  & ~n19499 ;
  assign n23208 = n19501 & ~n23206 ;
  assign n23209 = ~n23207 & n23208 ;
  assign n23210 = \core_eu_em_mac_em_reg_mr1swe_DO_reg[6]/P0001  & ~n19383 ;
  assign n23211 = ~n19508 & ~n23210 ;
  assign n23212 = ~n23209 & n23211 ;
  assign n23213 = ~n18262 & ~n23212 ;
  assign n23214 = \core_c_psq_MSTAT_reg_DO_reg[4]/NET0131  & ~n22957 ;
  assign n23215 = ~n17559 & ~n17682 ;
  assign n23216 = n22951 & ~n23215 ;
  assign n23217 = ~n22951 & n23215 ;
  assign n23218 = ~n23216 & ~n23217 ;
  assign n23219 = ~\core_c_psq_MSTAT_reg_DO_reg[4]/NET0131  & n23218 ;
  assign n23220 = ~n23214 & ~n23219 ;
  assign n23221 = n18262 & ~n23220 ;
  assign n23222 = ~n23213 & ~n23221 ;
  assign n23223 = n14752 & n23220 ;
  assign n23224 = n18276 & n19776 ;
  assign n23225 = \core_eu_em_mac_em_reg_mr1rwe_DO_reg[6]/P0001  & ~n17809 ;
  assign n23226 = n19780 & ~n23225 ;
  assign n23227 = ~n23224 & n23226 ;
  assign n23228 = ~n23223 & ~n23227 ;
  assign n23229 = \core_c_dec_IDLE_Eg_reg/P0001  & n4118 ;
  assign n23231 = n11741 & n21421 ;
  assign n23230 = n6024 & n21249 ;
  assign n23232 = ~\core_c_dec_IR_reg[4]/NET0131  & n23230 ;
  assign n23233 = n23231 & n23232 ;
  assign n23234 = ~n23229 & ~n23233 ;
  assign n23235 = n4117 & n5696 ;
  assign n23236 = \memc_ldSREG_E_reg/NET0131  & n23235 ;
  assign n23237 = n11751 & ~n11753 ;
  assign n23238 = n11734 & ~n23235 ;
  assign n23239 = ~n23237 & n23238 ;
  assign n23240 = ~n23236 & ~n23239 ;
  assign n23241 = ~\core_c_dec_MTMSTAT_Eg_reg/P0001  & ~\core_c_dec_Modctl_Eg_reg/P0001  ;
  assign n23242 = ~n14697 & n23241 ;
  assign n23243 = ~n5950 & ~n23242 ;
  assign n23245 = ~n14273 & n14404 ;
  assign n23244 = n14273 & ~n14406 ;
  assign n23246 = ~n13972 & ~n23244 ;
  assign n23247 = ~n23245 & n23246 ;
  assign n23248 = n14270 & ~n14274 ;
  assign n23249 = ~n13809 & ~n14010 ;
  assign n23250 = ~n23248 & n23249 ;
  assign n23251 = ~n23247 & n23250 ;
  assign n23252 = n23247 & ~n23250 ;
  assign n23253 = ~n23251 & ~n23252 ;
  assign n23254 = n13806 & ~n23253 ;
  assign n23255 = ~n13806 & ~n14658 ;
  assign n23256 = ~n23254 & ~n23255 ;
  assign n23257 = n14667 & ~n23256 ;
  assign n23258 = \core_eu_ea_alu_ea_reg_afswe_DO_reg[8]/P0001  & ~n14667 ;
  assign n23259 = ~n23257 & ~n23258 ;
  assign n23260 = n13805 & ~n23256 ;
  assign n23261 = \core_eu_ea_alu_ea_reg_afrwe_DO_reg[8]/P0001  & ~n13805 ;
  assign n23262 = ~n23260 & ~n23261 ;
  assign n23263 = ~n22669 & ~n22671 ;
  assign n23264 = n22671 & n22675 ;
  assign n23265 = ~n23263 & ~n23264 ;
  assign n23268 = ~\sport1_txctl_Wcnt_reg[4]/NET0131  & ~\sport1_txctl_Wcnt_reg[5]/NET0131  ;
  assign n23269 = ~\sport1_txctl_Wcnt_reg[6]/NET0131  & ~\sport1_txctl_Wcnt_reg[7]/NET0131  ;
  assign n23270 = n23268 & n23269 ;
  assign n23266 = ~\sport1_txctl_Wcnt_reg[0]/NET0131  & ~\sport1_txctl_Wcnt_reg[1]/NET0131  ;
  assign n23267 = ~\sport1_txctl_Wcnt_reg[2]/NET0131  & ~\sport1_txctl_Wcnt_reg[3]/NET0131  ;
  assign n23271 = n23266 & n23267 ;
  assign n23272 = n23270 & n23271 ;
  assign n23273 = ~n23263 & ~n23272 ;
  assign n23274 = ~n23265 & ~n23273 ;
  assign n23275 = ~n19952 & ~n19954 ;
  assign n23276 = n19954 & n19958 ;
  assign n23277 = ~n23275 & ~n23276 ;
  assign n23280 = ~\sport0_txctl_Wcnt_reg[4]/NET0131  & ~\sport0_txctl_Wcnt_reg[5]/NET0131  ;
  assign n23281 = ~\sport0_txctl_Wcnt_reg[6]/NET0131  & ~\sport0_txctl_Wcnt_reg[7]/NET0131  ;
  assign n23282 = n23280 & n23281 ;
  assign n23278 = ~\sport0_txctl_Wcnt_reg[0]/NET0131  & ~\sport0_txctl_Wcnt_reg[1]/NET0131  ;
  assign n23279 = ~\sport0_txctl_Wcnt_reg[2]/NET0131  & ~\sport0_txctl_Wcnt_reg[3]/NET0131  ;
  assign n23283 = n23278 & n23279 ;
  assign n23284 = n23282 & n23283 ;
  assign n23285 = ~n23275 & ~n23284 ;
  assign n23286 = ~n23277 & ~n23285 ;
  assign n23287 = \core_c_psq_SSTAT_reg[6]/NET0131  & ~n20574 ;
  assign n23288 = ~n20578 & ~n23287 ;
  assign n23289 = ~n4845 & n20579 ;
  assign n23290 = ~n23288 & ~n23289 ;
  assign n23291 = \core_c_psq_IFA_reg[0]/P0001  & ~n21242 ;
  assign n23292 = \core_c_psq_DRA_reg[0]/P0001  & n21242 ;
  assign n23293 = ~n23291 & ~n23292 ;
  assign n23294 = \core_c_psq_IFA_reg[9]/P0001  & ~n21242 ;
  assign n23295 = \core_c_psq_DRA_reg[9]/P0001  & n21242 ;
  assign n23296 = ~n23294 & ~n23295 ;
  assign n23297 = \core_c_psq_IFA_reg[8]/P0001  & ~n21242 ;
  assign n23298 = \core_c_psq_DRA_reg[8]/P0001  & n21242 ;
  assign n23299 = ~n23297 & ~n23298 ;
  assign n23300 = \core_c_psq_IFA_reg[7]/P0001  & ~n21242 ;
  assign n23301 = \core_c_psq_DRA_reg[7]/P0001  & n21242 ;
  assign n23302 = ~n23300 & ~n23301 ;
  assign n23303 = \core_c_psq_IFA_reg[6]/P0001  & ~n21242 ;
  assign n23304 = \core_c_psq_DRA_reg[6]/P0001  & n21242 ;
  assign n23305 = ~n23303 & ~n23304 ;
  assign n23306 = \core_c_psq_IFA_reg[5]/P0001  & ~n21242 ;
  assign n23307 = \core_c_psq_DRA_reg[5]/P0001  & n21242 ;
  assign n23308 = ~n23306 & ~n23307 ;
  assign n23309 = \core_c_psq_IFA_reg[4]/P0001  & ~n21242 ;
  assign n23310 = \core_c_psq_DRA_reg[4]/P0001  & n21242 ;
  assign n23311 = ~n23309 & ~n23310 ;
  assign n23312 = \core_c_psq_IFA_reg[3]/P0001  & ~n21242 ;
  assign n23313 = \core_c_psq_DRA_reg[3]/P0001  & n21242 ;
  assign n23314 = ~n23312 & ~n23313 ;
  assign n23315 = \core_c_psq_IFA_reg[2]/P0001  & ~n21242 ;
  assign n23316 = \core_c_psq_DRA_reg[2]/P0001  & n21242 ;
  assign n23317 = ~n23315 & ~n23316 ;
  assign n23318 = \core_c_psq_IFA_reg[1]/P0001  & ~n21242 ;
  assign n23319 = \core_c_psq_DRA_reg[1]/P0001  & n21242 ;
  assign n23320 = ~n23318 & ~n23319 ;
  assign n23321 = \core_c_psq_IFA_reg[12]/P0001  & ~n21242 ;
  assign n23322 = \core_c_psq_DRA_reg[12]/P0001  & n21242 ;
  assign n23323 = ~n23321 & ~n23322 ;
  assign n23324 = \core_c_psq_IFA_reg[11]/P0001  & ~n21242 ;
  assign n23325 = \core_c_psq_DRA_reg[11]/P0001  & n21242 ;
  assign n23326 = ~n23324 & ~n23325 ;
  assign n23327 = \core_c_psq_IFA_reg[10]/P0001  & ~n21242 ;
  assign n23328 = \core_c_psq_DRA_reg[10]/P0001  & n21242 ;
  assign n23329 = ~n23327 & ~n23328 ;
  assign n23330 = \core_c_psq_IFA_reg[13]/P0001  & ~n21242 ;
  assign n23331 = \core_c_psq_DRA_reg[13]/P0001  & n21242 ;
  assign n23332 = ~n23330 & ~n23331 ;
  assign n23333 = \core_c_dec_Post1_E_reg/P0001  & n4118 ;
  assign n23334 = n21421 & ~n21590 ;
  assign n23335 = ~n23333 & ~n23334 ;
  assign n23336 = ~n4117 & ~n19702 ;
  assign n23337 = \core_dag_ilm2reg_PMA_pi_DO_reg[13]/NET0131  & ~n23336 ;
  assign n23338 = ~n20687 & n23336 ;
  assign n23339 = ~n23337 & ~n23338 ;
  assign n23340 = \core_dag_ilm2reg_PMA_pi_DO_reg[12]/NET0131  & ~n23336 ;
  assign n23341 = ~n20698 & n23336 ;
  assign n23342 = ~n23340 & ~n23341 ;
  assign n23343 = ~n4057 & ~n5950 ;
  assign n23344 = ~\core_c_dec_accPM_E_reg/P0001  & \core_dag_ilm1reg_DMA_pi_DO_reg[9]/NET0131  ;
  assign n23345 = \core_c_dec_accPM_E_reg/P0001  & \core_dag_ilm2reg_PMA_pi_DO_reg[9]/NET0131  ;
  assign n23346 = ~n23344 & ~n23345 ;
  assign n23347 = n23343 & ~n23346 ;
  assign n23348 = \core_dag_ilm1reg_STAC_pi_DO_reg[9]/NET0131  & ~n23343 ;
  assign n23349 = ~n23347 & ~n23348 ;
  assign n23350 = ~\core_c_dec_accPM_E_reg/P0001  & \core_dag_ilm1reg_DMA_pi_DO_reg[8]/NET0131  ;
  assign n23351 = \core_c_dec_accPM_E_reg/P0001  & \core_dag_ilm2reg_PMA_pi_DO_reg[8]/NET0131  ;
  assign n23352 = ~n23350 & ~n23351 ;
  assign n23353 = n23343 & ~n23352 ;
  assign n23354 = \core_dag_ilm1reg_STAC_pi_DO_reg[8]/NET0131  & ~n23343 ;
  assign n23355 = ~n23353 & ~n23354 ;
  assign n23356 = ~\core_c_dec_accPM_E_reg/P0001  & \core_dag_ilm1reg_DMA_pi_DO_reg[7]/NET0131  ;
  assign n23357 = \core_c_dec_accPM_E_reg/P0001  & \core_dag_ilm2reg_PMA_pi_DO_reg[7]/NET0131  ;
  assign n23358 = ~n23356 & ~n23357 ;
  assign n23359 = n23343 & ~n23358 ;
  assign n23360 = \core_dag_ilm1reg_STAC_pi_DO_reg[7]/NET0131  & ~n23343 ;
  assign n23361 = ~n23359 & ~n23360 ;
  assign n23362 = ~\core_c_dec_accPM_E_reg/P0001  & \core_dag_ilm1reg_DMA_pi_DO_reg[6]/NET0131  ;
  assign n23363 = \core_c_dec_accPM_E_reg/P0001  & \core_dag_ilm2reg_PMA_pi_DO_reg[6]/NET0131  ;
  assign n23364 = ~n23362 & ~n23363 ;
  assign n23365 = n23343 & ~n23364 ;
  assign n23366 = \core_dag_ilm1reg_STAC_pi_DO_reg[6]/NET0131  & ~n23343 ;
  assign n23367 = ~n23365 & ~n23366 ;
  assign n23368 = ~\core_c_dec_accPM_E_reg/P0001  & \core_dag_ilm1reg_DMA_pi_DO_reg[5]/NET0131  ;
  assign n23369 = \core_c_dec_accPM_E_reg/P0001  & \core_dag_ilm2reg_PMA_pi_DO_reg[5]/NET0131  ;
  assign n23370 = ~n23368 & ~n23369 ;
  assign n23371 = n23343 & ~n23370 ;
  assign n23372 = \core_dag_ilm1reg_STAC_pi_DO_reg[5]/NET0131  & ~n23343 ;
  assign n23373 = ~n23371 & ~n23372 ;
  assign n23374 = ~\core_c_dec_accPM_E_reg/P0001  & \core_dag_ilm1reg_DMA_pi_DO_reg[13]/NET0131  ;
  assign n23375 = \core_c_dec_accPM_E_reg/P0001  & \core_dag_ilm2reg_PMA_pi_DO_reg[13]/NET0131  ;
  assign n23376 = ~n23374 & ~n23375 ;
  assign n23377 = n23343 & ~n23376 ;
  assign n23378 = \core_dag_ilm1reg_STAC_pi_DO_reg[13]/NET0131  & ~n23343 ;
  assign n23379 = ~n23377 & ~n23378 ;
  assign n23380 = ~\core_c_dec_accPM_E_reg/P0001  & \core_dag_ilm1reg_DMA_pi_DO_reg[12]/NET0131  ;
  assign n23381 = \core_c_dec_accPM_E_reg/P0001  & \core_dag_ilm2reg_PMA_pi_DO_reg[12]/NET0131  ;
  assign n23382 = ~n23380 & ~n23381 ;
  assign n23383 = n23343 & ~n23382 ;
  assign n23384 = \core_dag_ilm1reg_STAC_pi_DO_reg[12]/NET0131  & ~n23343 ;
  assign n23385 = ~n23383 & ~n23384 ;
  assign n23386 = ~\core_c_dec_accPM_E_reg/P0001  & \core_dag_ilm1reg_DMA_pi_DO_reg[11]/NET0131  ;
  assign n23387 = \core_c_dec_accPM_E_reg/P0001  & \core_dag_ilm2reg_PMA_pi_DO_reg[11]/NET0131  ;
  assign n23388 = ~n23386 & ~n23387 ;
  assign n23389 = n23343 & ~n23388 ;
  assign n23390 = \core_dag_ilm1reg_STAC_pi_DO_reg[11]/NET0131  & ~n23343 ;
  assign n23391 = ~n23389 & ~n23390 ;
  assign n23392 = ~\core_c_dec_accPM_E_reg/P0001  & \core_dag_ilm1reg_DMA_pi_DO_reg[10]/NET0131  ;
  assign n23393 = \core_c_dec_accPM_E_reg/P0001  & \core_dag_ilm2reg_PMA_pi_DO_reg[10]/NET0131  ;
  assign n23394 = ~n23392 & ~n23393 ;
  assign n23395 = n23343 & ~n23394 ;
  assign n23396 = \core_dag_ilm1reg_STAC_pi_DO_reg[10]/NET0131  & ~n23343 ;
  assign n23397 = ~n23395 & ~n23396 ;
  assign n23398 = n5429 & ~n14733 ;
  assign n23399 = \emc_IOcst_reg/NET0131  & ~n23398 ;
  assign n23400 = ~n19049 & n23399 ;
  assign n23401 = \memc_IOcmd_E_reg/NET0131  & ~n4068 ;
  assign n23402 = n19049 & n23401 ;
  assign n23403 = ~n23400 & ~n23402 ;
  assign n23404 = \core_eu_em_mac_em_reg_mfswe_DO_reg[15]/P0001  & ~n20864 ;
  assign n23405 = ~n19379 & n20864 ;
  assign n23406 = ~n23404 & ~n23405 ;
  assign n23407 = \sice_IAR_reg[1]/NET0131  & \sice_IAR_reg[2]/NET0131  ;
  assign n23408 = ~\sice_IAR_reg[0]/NET0131  & ~\sice_IAR_reg[3]/NET0131  ;
  assign n23409 = n23407 & n23408 ;
  assign n23410 = n23032 & n23409 ;
  assign n23411 = \sice_ICYC_en_reg/NET0131  & ~n23410 ;
  assign n23412 = \sice_SPC_reg[23]/P0001  & n23410 ;
  assign n23413 = ~n23411 & ~n23412 ;
  assign n23414 = \core_eu_em_mac_em_reg_mfrwe_DO_reg[15]/P0001  & ~n20990 ;
  assign n23415 = ~n19379 & n20990 ;
  assign n23416 = ~n23414 & ~n23415 ;
  assign n23417 = n20845 & n20847 ;
  assign n23418 = \clkc_oscntr_reg_DO_reg[4]/NET0131  & n23417 ;
  assign n23419 = \clkc_oscntr_reg_DO_reg[5]/NET0131  & n23418 ;
  assign n23420 = \clkc_oscntr_reg_DO_reg[6]/NET0131  & n23419 ;
  assign n23421 = \clkc_oscntr_reg_DO_reg[7]/NET0131  & n23420 ;
  assign n23422 = \clkc_oscntr_reg_DO_reg[8]/NET0131  & n23421 ;
  assign n23423 = ~\clkc_oscntr_reg_DO_reg[9]/NET0131  & ~n23422 ;
  assign n23424 = \clkc_oscntr_reg_DO_reg[9]/NET0131  & n23422 ;
  assign n23425 = ~n23423 & ~n23424 ;
  assign n23426 = \core_eu_em_mac_em_reg_mfswe_DO_reg[6]/P0001  & ~n20864 ;
  assign n23427 = n20864 & ~n23220 ;
  assign n23428 = ~n23426 & ~n23427 ;
  assign n23429 = \sport1_rxctl_a_sync1_reg/P0001  & ~\sport1_rxctl_a_sync2_reg/P0001  ;
  assign n23430 = \core_c_dec_MTRX1_E_reg/P0001  & n5951 ;
  assign n23431 = \sport1_rxctl_RX_reg[9]/P0001  & ~n23430 ;
  assign n23432 = n10289 & n23430 ;
  assign n23433 = ~n23431 & ~n23432 ;
  assign n23434 = ~n23429 & ~n23433 ;
  assign n23435 = \sport1_rxctl_RXSHT_reg[9]/P0001  & n23429 ;
  assign n23436 = ~n23434 & ~n23435 ;
  assign n23437 = \sport1_rxctl_RX_reg[8]/P0001  & ~n23430 ;
  assign n23438 = n10638 & n23430 ;
  assign n23439 = ~n23437 & ~n23438 ;
  assign n23440 = ~n23429 & ~n23439 ;
  assign n23441 = \sport1_rxctl_RXSHT_reg[8]/P0001  & n23429 ;
  assign n23442 = ~n23440 & ~n23441 ;
  assign n23443 = \sport1_rxctl_RX_reg[7]/P0001  & ~n23430 ;
  assign n23444 = n11265 & n23430 ;
  assign n23445 = ~n23443 & ~n23444 ;
  assign n23446 = ~n23429 & ~n23445 ;
  assign n23447 = \sport1_rxctl_RXSHT_reg[7]/P0001  & n23429 ;
  assign n23448 = ~n23446 & ~n23447 ;
  assign n23449 = \sport1_rxctl_RX_reg[4]/P0001  & ~n23430 ;
  assign n23450 = n10069 & n23430 ;
  assign n23451 = ~n23449 & ~n23450 ;
  assign n23452 = ~n23429 & ~n23451 ;
  assign n23453 = \sport1_rxctl_RXSHT_reg[4]/P0001  & n23429 ;
  assign n23454 = ~n23452 & ~n23453 ;
  assign n23455 = \sport1_rxctl_RX_reg[6]/P0001  & ~n23430 ;
  assign n23456 = n11525 & n23430 ;
  assign n23457 = ~n23455 & ~n23456 ;
  assign n23458 = ~n23429 & ~n23457 ;
  assign n23459 = \sport1_rxctl_RXSHT_reg[6]/P0001  & n23429 ;
  assign n23460 = ~n23458 & ~n23459 ;
  assign n23461 = \sport1_rxctl_RX_reg[3]/P0001  & ~n23430 ;
  assign n23462 = n8113 & n23430 ;
  assign n23463 = ~n23461 & ~n23462 ;
  assign n23464 = ~n23429 & ~n23463 ;
  assign n23465 = \sport1_rxctl_RXSHT_reg[3]/P0001  & n23429 ;
  assign n23466 = ~n23464 & ~n23465 ;
  assign n23467 = \sport1_rxctl_RX_reg[5]/P0001  & ~n23430 ;
  assign n23468 = n10911 & n23430 ;
  assign n23469 = ~n23467 & ~n23468 ;
  assign n23470 = ~n23429 & ~n23469 ;
  assign n23471 = \sport1_rxctl_RXSHT_reg[5]/P0001  & n23429 ;
  assign n23472 = ~n23470 & ~n23471 ;
  assign n23473 = \core_eu_em_mac_em_reg_mfrwe_DO_reg[6]/P0001  & ~n20990 ;
  assign n23474 = n20990 & ~n23220 ;
  assign n23475 = ~n23473 & ~n23474 ;
  assign n23476 = \sport1_rxctl_RX_reg[2]/P0001  & ~n23430 ;
  assign n23477 = n8715 & n23430 ;
  assign n23478 = ~n23476 & ~n23477 ;
  assign n23479 = ~n23429 & ~n23478 ;
  assign n23480 = \sport1_rxctl_RXSHT_reg[2]/P0001  & n23429 ;
  assign n23481 = ~n23479 & ~n23480 ;
  assign n23482 = \sport1_rxctl_RX_reg[1]/P0001  & ~n23430 ;
  assign n23483 = n9435 & n23430 ;
  assign n23484 = ~n23482 & ~n23483 ;
  assign n23485 = ~n23429 & ~n23484 ;
  assign n23486 = \sport1_rxctl_RXSHT_reg[1]/P0001  & n23429 ;
  assign n23487 = ~n23485 & ~n23486 ;
  assign n23488 = \sport1_rxctl_RX_reg[15]/P0001  & ~n23430 ;
  assign n23489 = n12743 & n23430 ;
  assign n23490 = ~n23488 & ~n23489 ;
  assign n23491 = ~n23429 & ~n23490 ;
  assign n23492 = \sport1_rxctl_RXSHT_reg[15]/P0001  & n23429 ;
  assign n23493 = ~n23491 & ~n23492 ;
  assign n23494 = \sport1_rxctl_RX_reg[14]/P0001  & ~n23430 ;
  assign n23495 = n12688 & n23430 ;
  assign n23496 = ~n23494 & ~n23495 ;
  assign n23497 = ~n23429 & ~n23496 ;
  assign n23498 = \sport1_rxctl_RXSHT_reg[14]/P0001  & n23429 ;
  assign n23499 = ~n23497 & ~n23498 ;
  assign n23500 = \sport1_rxctl_RX_reg[13]/P0001  & ~n23430 ;
  assign n23501 = n7340 & n23430 ;
  assign n23502 = ~n23500 & ~n23501 ;
  assign n23503 = ~n23429 & ~n23502 ;
  assign n23504 = \sport1_rxctl_RXSHT_reg[13]/P0001  & n23429 ;
  assign n23505 = ~n23503 & ~n23504 ;
  assign n23506 = \sport1_rxctl_RX_reg[12]/P0001  & ~n23430 ;
  assign n23507 = n9178 & n23430 ;
  assign n23508 = ~n23506 & ~n23507 ;
  assign n23509 = ~n23429 & ~n23508 ;
  assign n23510 = \sport1_rxctl_RXSHT_reg[12]/P0001  & n23429 ;
  assign n23511 = ~n23509 & ~n23510 ;
  assign n23512 = \sport1_rxctl_RX_reg[11]/P0001  & ~n23430 ;
  assign n23513 = n8460 & n23430 ;
  assign n23514 = ~n23512 & ~n23513 ;
  assign n23515 = ~n23429 & ~n23514 ;
  assign n23516 = \sport1_rxctl_RXSHT_reg[11]/P0001  & n23429 ;
  assign n23517 = ~n23515 & ~n23516 ;
  assign n23518 = \sport1_rxctl_RX_reg[10]/P0001  & ~n23430 ;
  assign n23519 = n7859 & n23430 ;
  assign n23520 = ~n23518 & ~n23519 ;
  assign n23521 = ~n23429 & ~n23520 ;
  assign n23522 = \sport1_rxctl_RXSHT_reg[10]/P0001  & n23429 ;
  assign n23523 = ~n23521 & ~n23522 ;
  assign n23524 = \sport1_rxctl_RX_reg[0]/P0001  & ~n23430 ;
  assign n23525 = n7607 & n23430 ;
  assign n23526 = ~n23524 & ~n23525 ;
  assign n23527 = ~n23429 & ~n23526 ;
  assign n23528 = \sport1_rxctl_RXSHT_reg[0]/P0001  & n23429 ;
  assign n23529 = ~n23527 & ~n23528 ;
  assign n23530 = \core_c_psq_Iact_E_reg[10]/NET0131  & ~n4116 ;
  assign n23531 = \core_c_psq_T_PWRDN_reg/P0001  & ~\core_c_psq_T_PWRDN_s1_reg/P0001  ;
  assign n23532 = ~\core_c_psq_Iflag_reg[10]/NET0131  & ~\sport0_regs_AUTO_a_reg[13]/NET0131  ;
  assign n23533 = ~n23531 & n23532 ;
  assign n23534 = ~n23530 & ~n23533 ;
  assign n23535 = ~\sice_ICYC_reg[9]/NET0131  & ~n20738 ;
  assign n23536 = ~n20739 & ~n23535 ;
  assign n23537 = ~\sice_IIRC_reg[6]/NET0131  & ~n18869 ;
  assign n23538 = ~n18870 & ~n23537 ;
  assign n23539 = ~\sice_IIRC_reg[9]/NET0131  & ~n20853 ;
  assign n23540 = ~n20854 & ~n23539 ;
  assign n23541 = ~\sice_ICYC_reg[6]/NET0131  & ~n18860 ;
  assign n23542 = ~n18861 & ~n23541 ;
  assign n23543 = \emc_DMDreg_reg[7]/P0001  & ~n14737 ;
  assign n23544 = \T_ED[7]_pad  & n14737 ;
  assign n23545 = ~n23543 & ~n23544 ;
  assign n23546 = \emc_DMDreg_reg[6]/P0001  & ~n14737 ;
  assign n23547 = \T_ED[6]_pad  & n14737 ;
  assign n23548 = ~n23546 & ~n23547 ;
  assign n23549 = \emc_DMDreg_reg[5]/P0001  & ~n14737 ;
  assign n23550 = \T_ED[5]_pad  & n14737 ;
  assign n23551 = ~n23549 & ~n23550 ;
  assign n23552 = \emc_DMDreg_reg[4]/P0001  & ~n14737 ;
  assign n23553 = \T_ED[4]_pad  & n14737 ;
  assign n23554 = ~n23552 & ~n23553 ;
  assign n23555 = \emc_DMDreg_reg[3]/P0001  & ~n14737 ;
  assign n23556 = \T_ED[3]_pad  & n14737 ;
  assign n23557 = ~n23555 & ~n23556 ;
  assign n23558 = \emc_DMDreg_reg[2]/P0001  & ~n14737 ;
  assign n23559 = \T_ED[2]_pad  & n14737 ;
  assign n23560 = ~n23558 & ~n23559 ;
  assign n23561 = \emc_DMDreg_reg[1]/P0001  & ~n14737 ;
  assign n23562 = \T_ED[1]_pad  & n14737 ;
  assign n23563 = ~n23561 & ~n23562 ;
  assign n23564 = \emc_DMDreg_reg[15]/P0001  & ~n14737 ;
  assign n23565 = \T_ED[15]_pad  & n14737 ;
  assign n23566 = ~n23564 & ~n23565 ;
  assign n23567 = \emc_DMDreg_reg[14]/P0001  & ~n14737 ;
  assign n23568 = \T_ED[14]_pad  & n14737 ;
  assign n23569 = ~n23567 & ~n23568 ;
  assign n23570 = \emc_DMDreg_reg[13]/P0001  & ~n14737 ;
  assign n23571 = \T_ED[13]_pad  & n14737 ;
  assign n23572 = ~n23570 & ~n23571 ;
  assign n23573 = \emc_DMDreg_reg[12]/P0001  & ~n14737 ;
  assign n23574 = \T_ED[12]_pad  & n14737 ;
  assign n23575 = ~n23573 & ~n23574 ;
  assign n23576 = \emc_DMDreg_reg[11]/P0001  & ~n14737 ;
  assign n23577 = \T_ED[11]_pad  & n14737 ;
  assign n23578 = ~n23576 & ~n23577 ;
  assign n23579 = \emc_DMDreg_reg[10]/P0001  & ~n14737 ;
  assign n23580 = \T_ED[10]_pad  & n14737 ;
  assign n23581 = ~n23579 & ~n23580 ;
  assign n23582 = \emc_DMDreg_reg[0]/P0001  & ~n14737 ;
  assign n23583 = \T_ED[0]_pad  & n14737 ;
  assign n23584 = ~n23582 & ~n23583 ;
  assign n23590 = n9272 & ~n9939 ;
  assign n23591 = ~n10789 & ~n11303 ;
  assign n23592 = n23590 & n23591 ;
  assign n23585 = \core_c_dec_SHTop_E_reg/P0001  & n17838 ;
  assign n23587 = n14033 & n23585 ;
  assign n23588 = ~n7172 & ~n7373 ;
  assign n23589 = n7995 & n8501 ;
  assign n23593 = n23588 & n23589 ;
  assign n23594 = n23587 & n23593 ;
  assign n23595 = n23592 & n23594 ;
  assign n23586 = ~\core_c_dec_IRE_reg[12]/NET0131  & n23585 ;
  assign n23596 = ~\core_c_dec_MTSE_E_reg/P0001  & ~n23586 ;
  assign n23597 = ~n23595 & n23596 ;
  assign n23598 = n13804 & ~n23597 ;
  assign n23599 = \core_c_dec_MTSE_E_reg/P0001  & ~n19559 ;
  assign n23600 = n17938 & n23585 ;
  assign n23601 = ~n18123 & n23600 ;
  assign n23602 = ~n17938 & n23585 ;
  assign n23603 = n18123 & n23602 ;
  assign n23604 = ~n23601 & ~n23603 ;
  assign n23605 = ~n18127 & n23600 ;
  assign n23606 = n18127 & n23602 ;
  assign n23607 = ~n23605 & ~n23606 ;
  assign n23611 = n17938 & ~n18102 ;
  assign n23612 = ~n17938 & n18102 ;
  assign n23613 = ~n23611 & ~n23612 ;
  assign n23608 = ~n17938 & n18098 ;
  assign n23609 = ~n18098 & ~n23602 ;
  assign n23610 = ~n23608 & ~n23609 ;
  assign n23614 = n23585 & n23610 ;
  assign n23615 = ~n23613 & n23614 ;
  assign n23616 = n23607 & ~n23615 ;
  assign n23617 = n23604 & ~n23616 ;
  assign n23618 = ~n18165 & n23600 ;
  assign n23619 = n18165 & n23602 ;
  assign n23620 = ~n23618 & ~n23619 ;
  assign n23621 = ~n23617 & n23620 ;
  assign n23623 = n17938 & n18161 ;
  assign n23622 = ~n17938 & ~n18161 ;
  assign n23624 = n23585 & ~n23622 ;
  assign n23625 = ~n23623 & n23624 ;
  assign n23626 = ~n23621 & ~n23625 ;
  assign n23628 = n17938 & n18186 ;
  assign n23627 = ~n17938 & ~n18186 ;
  assign n23629 = n23585 & ~n23627 ;
  assign n23630 = ~n23628 & n23629 ;
  assign n23631 = ~n23626 & ~n23630 ;
  assign n23632 = ~n18182 & n23600 ;
  assign n23633 = n18182 & n23602 ;
  assign n23634 = ~n23632 & ~n23633 ;
  assign n23635 = ~n23631 & n23634 ;
  assign n23636 = ~n18135 & n23600 ;
  assign n23637 = n18135 & n23602 ;
  assign n23638 = ~n23636 & ~n23637 ;
  assign n23639 = ~n23635 & n23638 ;
  assign n23640 = ~n18170 & n23600 ;
  assign n23641 = n18170 & n23602 ;
  assign n23642 = ~n23640 & ~n23641 ;
  assign n23643 = ~n23639 & n23642 ;
  assign n23644 = ~n18114 & n23600 ;
  assign n23645 = n18114 & n23602 ;
  assign n23646 = ~n23644 & ~n23645 ;
  assign n23647 = ~n23643 & n23646 ;
  assign n23648 = ~n18110 & n23600 ;
  assign n23649 = n18110 & n23602 ;
  assign n23650 = ~n23648 & ~n23649 ;
  assign n23651 = ~n23647 & n23650 ;
  assign n23652 = ~n17933 & n23600 ;
  assign n23653 = n17933 & n23602 ;
  assign n23654 = ~n23652 & ~n23653 ;
  assign n23655 = ~n23651 & n23654 ;
  assign n23656 = ~n17924 & n23600 ;
  assign n23657 = n17924 & n23602 ;
  assign n23658 = ~n23656 & ~n23657 ;
  assign n23659 = ~n23655 & n23658 ;
  assign n23660 = ~n18175 & n23600 ;
  assign n23661 = n18175 & n23602 ;
  assign n23662 = ~n23660 & ~n23661 ;
  assign n23663 = ~n23659 & n23662 ;
  assign n23664 = \core_eu_ec_cun_AV_reg/P0001  & n13881 ;
  assign n23665 = n23585 & n23664 ;
  assign n23667 = \core_eu_ec_cun_SS_reg/P0001  & n23602 ;
  assign n23666 = ~\core_eu_ec_cun_SS_reg/P0001  & n17938 ;
  assign n23668 = n23587 & ~n23666 ;
  assign n23669 = ~n23667 & n23668 ;
  assign n23670 = ~n23665 & ~n23669 ;
  assign n23671 = ~n23663 & n23670 ;
  assign n23672 = ~\core_c_dec_MTSE_E_reg/P0001  & n23671 ;
  assign n23673 = ~n23599 & ~n23672 ;
  assign n23674 = n23598 & ~n23673 ;
  assign n23675 = ~\core_eu_es_sht_es_reg_serwe_DO_reg[0]/P0001  & ~n23598 ;
  assign n23676 = ~n23674 & ~n23675 ;
  assign n23677 = n14666 & ~n23597 ;
  assign n23678 = ~n23673 & n23677 ;
  assign n23679 = ~\core_eu_es_sht_es_reg_seswe_DO_reg[0]/P0001  & ~n23677 ;
  assign n23680 = ~n23678 & ~n23679 ;
  assign n23681 = ~n13806 & n23253 ;
  assign n23682 = n13806 & n14623 ;
  assign n23683 = ~n23681 & ~n23682 ;
  assign n23684 = n14667 & ~n23683 ;
  assign n23685 = ~\core_eu_ea_alu_ea_reg_afswe_DO_reg[7]/P0001  & ~n14667 ;
  assign n23686 = ~n23684 & ~n23685 ;
  assign n23687 = n13805 & ~n23683 ;
  assign n23688 = ~\core_eu_ea_alu_ea_reg_afrwe_DO_reg[7]/P0001  & ~n13805 ;
  assign n23689 = ~n23687 & ~n23688 ;
  assign n23690 = n4149 & ~n20355 ;
  assign n23691 = n12234 & ~n23019 ;
  assign n23692 = ~\core_c_dec_cdAM_E_reg/P0001  & n4117 ;
  assign n23693 = n4116 & ~n14729 ;
  assign n23694 = ~n23692 & n23693 ;
  assign n23695 = \tm_tcr_reg_DO_reg[9]/NET0131  & n20355 ;
  assign n23699 = n22411 & n22423 ;
  assign n23697 = n22411 & ~n22422 ;
  assign n23698 = \tm_TCR_TMP_reg[9]/NET0131  & ~n23697 ;
  assign n23700 = ~n22400 & ~n23698 ;
  assign n23701 = ~n23699 & n23700 ;
  assign n23696 = ~\tm_tpr_reg_DO_reg[9]/NET0131  & n22400 ;
  assign n23702 = ~n20355 & ~n23696 ;
  assign n23703 = ~n23701 & n23702 ;
  assign n23704 = ~n23695 & ~n23703 ;
  assign n23705 = n13776 & n13778 ;
  assign n23706 = ~\core_c_psq_SSTAT_reg[3]/NET0131  & ~n23705 ;
  assign n23707 = \core_c_dec_DIVQ_E_reg/P0001  & n4117 ;
  assign n23708 = ~n21560 & ~n23707 ;
  assign n23709 = n4116 & ~n23708 ;
  assign n23710 = \bdma_BWcnt_reg[0]/NET0131  & n20036 ;
  assign n23711 = ~\bdma_BWcnt_reg[1]/NET0131  & ~n23710 ;
  assign n23712 = ~n20038 & ~n23711 ;
  assign n23713 = ~n13750 & n23712 ;
  assign n23716 = n4071 & n6929 ;
  assign n23717 = n4112 & n23716 ;
  assign n23714 = ~\clkc_SlowDn_reg/NET0131  & ~\clkc_SlowDn_s1_reg/P0001  ;
  assign n23715 = ~\clkc_SlowDn_s2_reg/P0001  & n23714 ;
  assign n23718 = ~n23018 & n23715 ;
  assign n23719 = n23717 & n23718 ;
  assign n23720 = \core_c_dec_NOP_E_reg/P0001  & n4117 ;
  assign n23721 = \core_c_dec_IR_reg[15]/NET0131  & ~\core_c_dec_IR_reg[16]/NET0131  ;
  assign n23722 = n21249 & n23721 ;
  assign n23723 = n5664 & n23722 ;
  assign n23724 = ~n23720 & ~n23723 ;
  assign n23725 = n4116 & ~n23724 ;
  assign n23726 = n23264 & ~n23272 ;
  assign n23727 = ~n23429 & ~n23430 ;
  assign n23728 = \sport1_cfg_SP_ENg_reg/NET0131  & \sport1_regs_AUTOreg_DO_reg[0]/NET0131  ;
  assign n23729 = ~n23727 & n23728 ;
  assign n23730 = ~\sport1_rxctl_RSreq_reg/NET0131  & ~n23729 ;
  assign n23731 = \emc_eRDY_reg/NET0131  & n4118 ;
  assign n23732 = ~\T_TMODE[1]_pad  & n5581 ;
  assign n23733 = n5560 & n23732 ;
  assign n23734 = \T_TMODE[1]_pad  & ~n5581 ;
  assign n23735 = n5605 & n23734 ;
  assign n23736 = ~n23733 & ~n23735 ;
  assign n23737 = ~\emc_eRDY_reg/NET0131  & ~n5586 ;
  assign n23738 = ~n23736 & n23737 ;
  assign n23739 = ~n23731 & ~n23738 ;
  assign n23740 = ~\sport0_regs_SCTLreg_DO_reg[5]/NET0131  & n20868 ;
  assign n23741 = ~n20875 & ~n23740 ;
  assign n23742 = \sport0_cfg_SP_ENg_reg/NET0131  & ~n23741 ;
  assign n23743 = \sport0_regs_SCTLreg_DO_reg[5]/NET0131  & \sport0_txctl_b_sync1_reg/P0001  ;
  assign n23744 = n23276 & ~n23284 ;
  assign n23745 = \memc_LDaST_Eg_reg/NET0131  & n4117 ;
  assign n23746 = n5946 & ~n11748 ;
  assign n23747 = n13130 & ~n13580 ;
  assign n23748 = ~n23746 & ~n23747 ;
  assign n23749 = n6931 & ~n23748 ;
  assign n23750 = n11741 & n23749 ;
  assign n23751 = ~n23745 & ~n23750 ;
  assign n23752 = \memc_selMIO_E_reg/P0001  & n23235 ;
  assign n23753 = ~n23238 & ~n23752 ;
  assign n23754 = \core_c_dec_MTSI_E_reg/P0001  & n14665 ;
  assign n23755 = ~\core_c_dec_accPM_E_reg/P0001  & ~n8460 ;
  assign n23756 = \core_c_dec_accPM_E_reg/P0001  & ~n12590 ;
  assign n23757 = ~n23755 & ~n23756 ;
  assign n23758 = n23754 & ~n23757 ;
  assign n23759 = ~\core_eu_es_sht_es_reg_siswe_DO_reg[11]/P0001  & ~n23754 ;
  assign n23760 = ~n23758 & ~n23759 ;
  assign n23761 = n6106 & ~n7859 ;
  assign n23762 = ~n6106 & n7644 ;
  assign n23763 = ~n23761 & ~n23762 ;
  assign n23764 = ~n6084 & n23763 ;
  assign n23765 = ~n8133 & ~n23764 ;
  assign n23766 = \core_c_dec_MTMY1_E_reg/P0001  & n14665 ;
  assign n23767 = ~n21994 & n23766 ;
  assign n23768 = ~\core_eu_em_mac_em_reg_my1swe_DO_reg[9]/P0001  & ~n23766 ;
  assign n23769 = ~n23767 & ~n23768 ;
  assign n23770 = \core_eu_em_mac_em_reg_my1swe_DO_reg[8]/P0001  & ~n23766 ;
  assign n23771 = ~n22003 & n23766 ;
  assign n23772 = ~n23770 & ~n23771 ;
  assign n23773 = ~n22084 & n23766 ;
  assign n23774 = ~\core_eu_em_mac_em_reg_my1swe_DO_reg[13]/P0001  & ~n23766 ;
  assign n23775 = ~n23773 & ~n23774 ;
  assign n23776 = \core_eu_em_mac_em_reg_my1swe_DO_reg[12]/P0001  & ~n23766 ;
  assign n23777 = ~n22093 & n23766 ;
  assign n23778 = ~n23776 & ~n23777 ;
  assign n23779 = \core_eu_em_mac_em_reg_my1swe_DO_reg[11]/P0001  & ~n23766 ;
  assign n23780 = ~n22105 & n23766 ;
  assign n23781 = ~n23779 & ~n23780 ;
  assign n23782 = \core_c_dec_MTMY1_E_reg/P0001  & n17798 ;
  assign n23783 = ~n21994 & n23782 ;
  assign n23784 = ~\core_eu_em_mac_em_reg_my1rwe_DO_reg[9]/P0001  & ~n23782 ;
  assign n23785 = ~n23783 & ~n23784 ;
  assign n23786 = ~n22084 & n23782 ;
  assign n23787 = ~\core_eu_em_mac_em_reg_my1rwe_DO_reg[13]/P0001  & ~n23782 ;
  assign n23788 = ~n23786 & ~n23787 ;
  assign n23789 = \core_eu_em_mac_em_reg_my1rwe_DO_reg[12]/P0001  & ~n23782 ;
  assign n23790 = ~n22093 & n23782 ;
  assign n23791 = ~n23789 & ~n23790 ;
  assign n23792 = \core_eu_em_mac_em_reg_my1rwe_DO_reg[11]/P0001  & ~n23782 ;
  assign n23793 = ~n22105 & n23782 ;
  assign n23794 = ~n23792 & ~n23793 ;
  assign n23795 = ~n22114 & n23782 ;
  assign n23796 = ~\core_eu_em_mac_em_reg_my1rwe_DO_reg[10]/P0001  & ~n23782 ;
  assign n23797 = ~n23795 & ~n23796 ;
  assign n23798 = \core_c_dec_MTMY0_E_reg/P0001  & n14665 ;
  assign n23799 = ~n21994 & n23798 ;
  assign n23800 = ~\core_eu_em_mac_em_reg_my0swe_DO_reg[9]/P0001  & ~n23798 ;
  assign n23801 = ~n23799 & ~n23800 ;
  assign n23802 = \core_eu_em_mac_em_reg_my0swe_DO_reg[8]/P0001  & ~n23798 ;
  assign n23803 = ~n22003 & n23798 ;
  assign n23804 = ~n23802 & ~n23803 ;
  assign n23805 = \core_eu_em_mac_em_reg_my0swe_DO_reg[12]/P0001  & ~n23798 ;
  assign n23806 = ~n22093 & n23798 ;
  assign n23807 = ~n23805 & ~n23806 ;
  assign n23808 = \core_eu_em_mac_em_reg_my0swe_DO_reg[11]/P0001  & ~n23798 ;
  assign n23809 = ~n22105 & n23798 ;
  assign n23810 = ~n23808 & ~n23809 ;
  assign n23811 = ~n22114 & n23798 ;
  assign n23812 = ~\core_eu_em_mac_em_reg_my0swe_DO_reg[10]/P0001  & ~n23798 ;
  assign n23813 = ~n23811 & ~n23812 ;
  assign n23814 = \core_c_dec_MTMY0_E_reg/P0001  & n17798 ;
  assign n23815 = ~n21994 & n23814 ;
  assign n23816 = ~\core_eu_em_mac_em_reg_my0rwe_DO_reg[9]/P0001  & ~n23814 ;
  assign n23817 = ~n23815 & ~n23816 ;
  assign n23818 = \core_eu_em_mac_em_reg_my0rwe_DO_reg[8]/P0001  & ~n23814 ;
  assign n23819 = ~n22003 & n23814 ;
  assign n23820 = ~n23818 & ~n23819 ;
  assign n23821 = \core_eu_em_mac_em_reg_my0rwe_DO_reg[12]/P0001  & ~n23814 ;
  assign n23822 = ~n22093 & n23814 ;
  assign n23823 = ~n23821 & ~n23822 ;
  assign n23824 = ~n22114 & n23814 ;
  assign n23825 = ~\core_eu_em_mac_em_reg_my0rwe_DO_reg[10]/P0001  & ~n23814 ;
  assign n23826 = ~n23824 & ~n23825 ;
  assign n23827 = n7530 & n13762 ;
  assign n23828 = ~n10289 & n23827 ;
  assign n23829 = ~\bdma_BOVL_reg[9]/NET0131  & ~n23827 ;
  assign n23830 = ~n23828 & ~n23829 ;
  assign n23831 = ~n10638 & n23827 ;
  assign n23832 = ~\bdma_BOVL_reg[8]/NET0131  & ~n23827 ;
  assign n23833 = ~n23831 & ~n23832 ;
  assign n23834 = ~n8460 & n23827 ;
  assign n23835 = ~\bdma_BOVL_reg[11]/NET0131  & ~n23827 ;
  assign n23836 = ~n23834 & ~n23835 ;
  assign n23837 = ~n7859 & n23827 ;
  assign n23838 = ~\bdma_BOVL_reg[10]/NET0131  & ~n23827 ;
  assign n23839 = ~n23837 & ~n23838 ;
  assign n23840 = ~n10289 & n21268 ;
  assign n23841 = ~\bdma_BCTL_reg[9]/NET0131  & ~n21268 ;
  assign n23842 = ~n23840 & ~n23841 ;
  assign n23843 = ~n10638 & n21268 ;
  assign n23844 = ~\bdma_BCTL_reg[8]/NET0131  & ~n21268 ;
  assign n23845 = ~n23843 & ~n23844 ;
  assign n23846 = ~n7340 & n21268 ;
  assign n23847 = ~\bdma_BCTL_reg[13]/NET0131  & ~n21268 ;
  assign n23848 = ~n23846 & ~n23847 ;
  assign n23849 = ~n9178 & n21268 ;
  assign n23850 = ~\bdma_BCTL_reg[12]/NET0131  & ~n21268 ;
  assign n23851 = ~n23849 & ~n23850 ;
  assign n23852 = ~n8460 & n21268 ;
  assign n23853 = ~\bdma_BCTL_reg[11]/NET0131  & ~n21268 ;
  assign n23854 = ~n23852 & ~n23853 ;
  assign n23855 = ~n7859 & n21268 ;
  assign n23856 = ~\bdma_BCTL_reg[10]/NET0131  & ~n21268 ;
  assign n23857 = ~n23855 & ~n23856 ;
  assign n23858 = ~\core_c_dec_accPM_E_reg/P0001  & ~n10638 ;
  assign n23859 = \core_c_dec_accPM_E_reg/P0001  & ~n13041 ;
  assign n23860 = ~n23858 & ~n23859 ;
  assign n23861 = n23754 & ~n23860 ;
  assign n23862 = ~\core_eu_es_sht_es_reg_siswe_DO_reg[8]/P0001  & ~n23754 ;
  assign n23863 = ~n23861 & ~n23862 ;
  assign n23864 = \core_c_dec_MTTX1_E_reg/P0001  & n5951 ;
  assign n23865 = ~\auctl_T1Sack_reg/NET0131  & ~n23864 ;
  assign n23866 = n10289 & ~n23865 ;
  assign n23867 = \sport1_txctl_TX_reg[9]/P0001  & n23865 ;
  assign n23868 = ~n23866 & ~n23867 ;
  assign n23869 = n10638 & ~n23865 ;
  assign n23870 = \sport1_txctl_TX_reg[8]/P0001  & n23865 ;
  assign n23871 = ~n23869 & ~n23870 ;
  assign n23872 = n9178 & ~n23865 ;
  assign n23873 = \sport1_txctl_TX_reg[12]/P0001  & n23865 ;
  assign n23874 = ~n23872 & ~n23873 ;
  assign n23875 = n8460 & ~n23865 ;
  assign n23876 = \sport1_txctl_TX_reg[11]/P0001  & n23865 ;
  assign n23877 = ~n23875 & ~n23876 ;
  assign n23878 = n7859 & ~n23865 ;
  assign n23879 = \sport1_txctl_TX_reg[10]/P0001  & n23865 ;
  assign n23880 = ~n23878 & ~n23879 ;
  assign n23881 = \core_eu_em_mac_em_reg_my1rwe_DO_reg[8]/P0001  & ~n23782 ;
  assign n23882 = ~n22003 & n23782 ;
  assign n23883 = ~n23881 & ~n23882 ;
  assign n23884 = n6106 & ~n8113 ;
  assign n23885 = ~n6106 & n8224 ;
  assign n23886 = ~n23884 & ~n23885 ;
  assign n23887 = ~n6084 & n23886 ;
  assign n23888 = ~n8177 & ~n23887 ;
  assign n23889 = \core_c_dec_MTAY1_E_reg/P0001  & n14665 ;
  assign n23890 = ~n21994 & n23889 ;
  assign n23891 = ~\core_eu_ea_alu_ea_reg_ay1swe_DO_reg[9]/P0001  & ~n23889 ;
  assign n23892 = ~n23890 & ~n23891 ;
  assign n23893 = \core_eu_ea_alu_ea_reg_ay1swe_DO_reg[8]/P0001  & ~n23889 ;
  assign n23894 = ~n22003 & n23889 ;
  assign n23895 = ~n23893 & ~n23894 ;
  assign n23896 = ~n22084 & n23889 ;
  assign n23897 = ~\core_eu_ea_alu_ea_reg_ay1swe_DO_reg[13]/P0001  & ~n23889 ;
  assign n23898 = ~n23896 & ~n23897 ;
  assign n23899 = \core_eu_ea_alu_ea_reg_ay1swe_DO_reg[12]/P0001  & ~n23889 ;
  assign n23900 = ~n22093 & n23889 ;
  assign n23901 = ~n23899 & ~n23900 ;
  assign n23902 = \core_eu_ea_alu_ea_reg_ay1swe_DO_reg[11]/P0001  & ~n23889 ;
  assign n23903 = ~n22105 & n23889 ;
  assign n23904 = ~n23902 & ~n23903 ;
  assign n23905 = ~n22114 & n23889 ;
  assign n23906 = ~\core_eu_ea_alu_ea_reg_ay1swe_DO_reg[10]/P0001  & ~n23889 ;
  assign n23907 = ~n23905 & ~n23906 ;
  assign n23908 = \core_c_dec_MTAX1_E_reg/P0001  & n14665 ;
  assign n23909 = ~n19504 & n23908 ;
  assign n23910 = ~\core_eu_ea_alu_ea_reg_ax1swe_DO_reg[9]/P0001  & ~n23908 ;
  assign n23911 = ~n23909 & ~n23910 ;
  assign n23912 = ~n23860 & n23908 ;
  assign n23913 = ~\core_eu_ea_alu_ea_reg_ax1swe_DO_reg[8]/P0001  & ~n23908 ;
  assign n23914 = ~n23912 & ~n23913 ;
  assign n23915 = ~n17836 & n23908 ;
  assign n23916 = ~\core_eu_ea_alu_ea_reg_ax1swe_DO_reg[13]/P0001  & ~n23908 ;
  assign n23917 = ~n23915 & ~n23916 ;
  assign n23918 = ~\core_c_dec_accPM_E_reg/P0001  & ~n9178 ;
  assign n23919 = \core_c_dec_accPM_E_reg/P0001  & ~n12624 ;
  assign n23920 = ~n23918 & ~n23919 ;
  assign n23921 = n23908 & ~n23920 ;
  assign n23922 = ~\core_eu_ea_alu_ea_reg_ax1swe_DO_reg[12]/P0001  & ~n23908 ;
  assign n23923 = ~n23921 & ~n23922 ;
  assign n23924 = ~n23757 & n23908 ;
  assign n23925 = ~\core_eu_ea_alu_ea_reg_ax1swe_DO_reg[11]/P0001  & ~n23908 ;
  assign n23926 = ~n23924 & ~n23925 ;
  assign n23927 = ~n19848 & n23908 ;
  assign n23928 = ~\core_eu_ea_alu_ea_reg_ax1swe_DO_reg[10]/P0001  & ~n23908 ;
  assign n23929 = ~n23927 & ~n23928 ;
  assign n23930 = \core_c_dec_MTAX0_E_reg/P0001  & n14665 ;
  assign n23931 = ~n19504 & n23930 ;
  assign n23932 = ~\core_eu_ea_alu_ea_reg_ax0swe_DO_reg[9]/P0001  & ~n23930 ;
  assign n23933 = ~n23931 & ~n23932 ;
  assign n23934 = ~n23860 & n23930 ;
  assign n23935 = ~\core_eu_ea_alu_ea_reg_ax0swe_DO_reg[8]/P0001  & ~n23930 ;
  assign n23936 = ~n23934 & ~n23935 ;
  assign n23937 = ~n17836 & n23930 ;
  assign n23938 = ~\core_eu_ea_alu_ea_reg_ax0swe_DO_reg[13]/P0001  & ~n23930 ;
  assign n23939 = ~n23937 & ~n23938 ;
  assign n23940 = ~n23920 & n23930 ;
  assign n23941 = ~\core_eu_ea_alu_ea_reg_ax0swe_DO_reg[12]/P0001  & ~n23930 ;
  assign n23942 = ~n23940 & ~n23941 ;
  assign n23943 = ~n23757 & n23930 ;
  assign n23944 = ~\core_eu_ea_alu_ea_reg_ax0swe_DO_reg[11]/P0001  & ~n23930 ;
  assign n23945 = ~n23943 & ~n23944 ;
  assign n23946 = ~n19848 & n23930 ;
  assign n23947 = ~\core_eu_ea_alu_ea_reg_ax0swe_DO_reg[10]/P0001  & ~n23930 ;
  assign n23948 = ~n23946 & ~n23947 ;
  assign n23949 = \core_eu_em_mac_em_reg_my0rwe_DO_reg[11]/P0001  & ~n23814 ;
  assign n23950 = ~n22105 & n23814 ;
  assign n23951 = ~n23949 & ~n23950 ;
  assign n23952 = ~n22084 & n23814 ;
  assign n23953 = ~\core_eu_em_mac_em_reg_my0rwe_DO_reg[13]/P0001  & ~n23814 ;
  assign n23954 = ~n23952 & ~n23953 ;
  assign n23955 = ~\core_c_dec_Dummy_E_reg/NET0131  & \core_c_dec_MTIreg_E_reg[7]/P0001  ;
  assign n23956 = ~n5999 & ~n23955 ;
  assign n23957 = ~n5994 & n23956 ;
  assign n23958 = ~n6000 & ~n23957 ;
  assign n23959 = \core_dag_ilm2reg_I7_we_DO_reg[9]/NET0131  & ~n23958 ;
  assign n23960 = ~n6000 & n20755 ;
  assign n23961 = ~n23959 & ~n23960 ;
  assign n23962 = \core_dag_ilm2reg_I7_we_DO_reg[6]/NET0131  & ~n23958 ;
  assign n23963 = ~n6000 & n20624 ;
  assign n23964 = ~n23962 & ~n23963 ;
  assign n23965 = \core_dag_ilm2reg_I7_we_DO_reg[5]/NET0131  & ~n23958 ;
  assign n23966 = ~n6000 & n20634 ;
  assign n23967 = ~n23965 & ~n23966 ;
  assign n23968 = \core_dag_ilm2reg_I7_we_DO_reg[13]/NET0131  & ~n23958 ;
  assign n23969 = ~n6000 & ~n20685 ;
  assign n23970 = ~n23968 & ~n23969 ;
  assign n23971 = \core_dag_ilm2reg_I7_we_DO_reg[12]/NET0131  & ~n23958 ;
  assign n23972 = ~n6000 & ~n20696 ;
  assign n23973 = ~n23971 & ~n23972 ;
  assign n23974 = ~n6008 & n20755 ;
  assign n23975 = \core_dag_ilm2reg_I6_we_DO_reg[9]/NET0131  & n6008 ;
  assign n23976 = ~n23974 & ~n23975 ;
  assign n23977 = ~n6008 & n20602 ;
  assign n23978 = \core_dag_ilm2reg_I6_we_DO_reg[8]/NET0131  & n6008 ;
  assign n23979 = ~n23977 & ~n23978 ;
  assign n23980 = ~n6008 & n20614 ;
  assign n23981 = \core_dag_ilm2reg_I6_we_DO_reg[7]/NET0131  & n6008 ;
  assign n23982 = ~n23980 & ~n23981 ;
  assign n23983 = ~n6008 & n20624 ;
  assign n23984 = \core_dag_ilm2reg_I6_we_DO_reg[6]/NET0131  & n6008 ;
  assign n23985 = ~n23983 & ~n23984 ;
  assign n23986 = ~n6008 & n20634 ;
  assign n23987 = \core_dag_ilm2reg_I6_we_DO_reg[5]/NET0131  & n6008 ;
  assign n23988 = ~n23986 & ~n23987 ;
  assign n23989 = ~n6008 & ~n20685 ;
  assign n23990 = \core_dag_ilm2reg_I6_we_DO_reg[13]/NET0131  & n6008 ;
  assign n23991 = ~n23989 & ~n23990 ;
  assign n23992 = ~n6008 & ~n20696 ;
  assign n23993 = \core_dag_ilm2reg_I6_we_DO_reg[12]/NET0131  & n6008 ;
  assign n23994 = ~n23992 & ~n23993 ;
  assign n23995 = ~n6008 & ~n20707 ;
  assign n23996 = \core_dag_ilm2reg_I6_we_DO_reg[11]/NET0131  & n6008 ;
  assign n23997 = ~n23995 & ~n23996 ;
  assign n23998 = ~n6008 & n20718 ;
  assign n23999 = \core_dag_ilm2reg_I6_we_DO_reg[10]/NET0131  & n6008 ;
  assign n24000 = ~n23998 & ~n23999 ;
  assign n24001 = ~\core_c_dec_Dummy_E_reg/NET0131  & \core_c_dec_MTIreg_E_reg[5]/P0001  ;
  assign n24002 = ~n6014 & ~n24001 ;
  assign n24003 = ~n6011 & n24002 ;
  assign n24004 = ~n6015 & ~n24003 ;
  assign n24005 = \core_dag_ilm2reg_I5_we_DO_reg[9]/NET0131  & ~n24004 ;
  assign n24006 = ~n6015 & n20755 ;
  assign n24007 = ~n24005 & ~n24006 ;
  assign n24008 = \core_dag_ilm2reg_I5_we_DO_reg[6]/NET0131  & ~n24004 ;
  assign n24009 = ~n6015 & n20624 ;
  assign n24010 = ~n24008 & ~n24009 ;
  assign n24011 = \core_dag_ilm2reg_I5_we_DO_reg[5]/NET0131  & ~n24004 ;
  assign n24012 = ~n6015 & n20634 ;
  assign n24013 = ~n24011 & ~n24012 ;
  assign n24014 = \core_dag_ilm2reg_I5_we_DO_reg[13]/NET0131  & ~n24004 ;
  assign n24015 = ~n6015 & ~n20685 ;
  assign n24016 = ~n24014 & ~n24015 ;
  assign n24017 = \core_dag_ilm2reg_I5_we_DO_reg[12]/NET0131  & ~n24004 ;
  assign n24018 = ~n6015 & ~n20696 ;
  assign n24019 = ~n24017 & ~n24018 ;
  assign n24020 = ~\core_c_dec_Dummy_E_reg/NET0131  & \core_c_dec_MTIreg_E_reg[4]/P0001  ;
  assign n24021 = ~n5963 & ~n24020 ;
  assign n24022 = ~n5958 & n24021 ;
  assign n24023 = ~n5964 & ~n24022 ;
  assign n24024 = \core_dag_ilm2reg_I4_we_DO_reg[9]/NET0131  & ~n24023 ;
  assign n24025 = ~n5964 & n20755 ;
  assign n24026 = ~n24024 & ~n24025 ;
  assign n24027 = \core_dag_ilm2reg_I4_we_DO_reg[8]/NET0131  & ~n24023 ;
  assign n24028 = n20602 & n24023 ;
  assign n24029 = ~n24027 & ~n24028 ;
  assign n24030 = \core_dag_ilm2reg_I4_we_DO_reg[7]/NET0131  & ~n24023 ;
  assign n24031 = n20614 & n24023 ;
  assign n24032 = ~n24030 & ~n24031 ;
  assign n24033 = \core_dag_ilm2reg_I4_we_DO_reg[6]/NET0131  & ~n24023 ;
  assign n24034 = ~n5964 & n20624 ;
  assign n24035 = ~n24033 & ~n24034 ;
  assign n24036 = \core_dag_ilm2reg_I4_we_DO_reg[5]/NET0131  & ~n24023 ;
  assign n24037 = ~n5964 & n20634 ;
  assign n24038 = ~n24036 & ~n24037 ;
  assign n24039 = \core_dag_ilm2reg_I4_we_DO_reg[13]/NET0131  & ~n24023 ;
  assign n24040 = ~n5964 & ~n20685 ;
  assign n24041 = ~n24039 & ~n24040 ;
  assign n24042 = \core_dag_ilm2reg_I4_we_DO_reg[12]/NET0131  & ~n24023 ;
  assign n24043 = ~n5964 & ~n20696 ;
  assign n24044 = ~n24042 & ~n24043 ;
  assign n24045 = ~n20707 & n24023 ;
  assign n24046 = \core_dag_ilm2reg_I4_we_DO_reg[11]/NET0131  & ~n24023 ;
  assign n24047 = ~n24045 & ~n24046 ;
  assign n24048 = ~n20718 & n24023 ;
  assign n24049 = ~\core_dag_ilm2reg_I4_we_DO_reg[10]/NET0131  & ~n24023 ;
  assign n24050 = ~n24048 & ~n24049 ;
  assign n24051 = ~n19504 & n23754 ;
  assign n24052 = ~\core_eu_es_sht_es_reg_siswe_DO_reg[9]/P0001  & ~n23754 ;
  assign n24053 = ~n24051 & ~n24052 ;
  assign n24054 = n23754 & ~n23920 ;
  assign n24055 = ~\core_eu_es_sht_es_reg_siswe_DO_reg[12]/P0001  & ~n23754 ;
  assign n24056 = ~n24054 & ~n24055 ;
  assign n24057 = ~n22084 & n23798 ;
  assign n24058 = ~\core_eu_em_mac_em_reg_my0swe_DO_reg[13]/P0001  & ~n23798 ;
  assign n24059 = ~n24057 & ~n24058 ;
  assign n24060 = n6106 & ~n10638 ;
  assign n24061 = ~n6106 & n10343 ;
  assign n24062 = ~n24060 & ~n24061 ;
  assign n24063 = ~n6075 & n24062 ;
  assign n24064 = \core_dag_ilm1reg_I3_we_DO_reg[8]/NET0131  & n6075 ;
  assign n24065 = ~n24063 & ~n24064 ;
  assign n24066 = n6106 & ~n10911 ;
  assign n24067 = ~n6106 & n10663 ;
  assign n24068 = ~n24066 & ~n24067 ;
  assign n24069 = ~n6075 & ~n24068 ;
  assign n24070 = ~\core_dag_ilm1reg_I3_we_DO_reg[5]/NET0131  & n6075 ;
  assign n24071 = ~n24069 & ~n24070 ;
  assign n24072 = n6106 & ~n9435 ;
  assign n24073 = ~n6106 & n8926 ;
  assign n24074 = ~n24072 & ~n24073 ;
  assign n24075 = ~n6075 & ~n24074 ;
  assign n24076 = ~\core_dag_ilm1reg_I3_we_DO_reg[1]/NET0131  & n6075 ;
  assign n24077 = ~n24075 & ~n24076 ;
  assign n24078 = n6106 & ~n7340 ;
  assign n24079 = ~n6106 & n6546 ;
  assign n24080 = ~n24078 & ~n24079 ;
  assign n24081 = ~n6075 & n24080 ;
  assign n24082 = \core_dag_ilm1reg_I3_we_DO_reg[13]/NET0131  & n6075 ;
  assign n24083 = ~n24081 & ~n24082 ;
  assign n24084 = ~n6106 & ~n8962 ;
  assign n24085 = n6106 & n9178 ;
  assign n24086 = ~n24084 & ~n24085 ;
  assign n24087 = ~n6075 & ~n24086 ;
  assign n24088 = ~n8869 & ~n24087 ;
  assign n24089 = ~n6106 & ~n8246 ;
  assign n24090 = n6106 & n8460 ;
  assign n24091 = ~n24089 & ~n24090 ;
  assign n24092 = ~n6075 & ~n24091 ;
  assign n24093 = ~n8738 & ~n24092 ;
  assign n24094 = ~n6075 & n23763 ;
  assign n24095 = ~n8137 & ~n24094 ;
  assign n24096 = ~n6106 & ~n9752 ;
  assign n24097 = n6106 & n10289 ;
  assign n24098 = ~n24096 & ~n24097 ;
  assign n24099 = ~n6084 & ~n24098 ;
  assign n24100 = \core_dag_ilm1reg_I2_we_DO_reg[9]/NET0131  & n6084 ;
  assign n24101 = ~n24099 & ~n24100 ;
  assign n24102 = ~n6084 & n24062 ;
  assign n24103 = ~n10398 & ~n24102 ;
  assign n24104 = ~n6106 & ~n10954 ;
  assign n24105 = n6106 & n11265 ;
  assign n24106 = ~n24104 & ~n24105 ;
  assign n24107 = ~n6084 & ~n24106 ;
  assign n24108 = ~n11008 & ~n24107 ;
  assign n24109 = ~n6106 & ~n11280 ;
  assign n24110 = n6106 & n11525 ;
  assign n24111 = ~n24109 & ~n24110 ;
  assign n24112 = ~n6084 & ~n24111 ;
  assign n24113 = ~n10979 & ~n24112 ;
  assign n24114 = ~n6084 & n24068 ;
  assign n24115 = ~n10371 & ~n24114 ;
  assign n24116 = ~n6106 & ~n10302 ;
  assign n24117 = n6106 & n10069 ;
  assign n24118 = ~n24116 & ~n24117 ;
  assign n24119 = ~n6084 & ~n24118 ;
  assign n24120 = \core_dag_ilm1reg_I2_we_DO_reg[4]/NET0131  & n6084 ;
  assign n24121 = ~n24119 & ~n24120 ;
  assign n24122 = ~n6106 & ~n8794 ;
  assign n24123 = n6106 & n8715 ;
  assign n24124 = ~n24122 & ~n24123 ;
  assign n24125 = ~n6084 & ~n24124 ;
  assign n24126 = ~n8766 & ~n24125 ;
  assign n24127 = ~n6084 & ~n24074 ;
  assign n24128 = ~\core_dag_ilm1reg_I2_we_DO_reg[1]/NET0131  & n6084 ;
  assign n24129 = ~n24127 & ~n24128 ;
  assign n24130 = ~n6084 & n24080 ;
  assign n24131 = \core_dag_ilm1reg_I2_we_DO_reg[13]/NET0131  & n6084 ;
  assign n24132 = ~n24130 & ~n24131 ;
  assign n24133 = ~n6084 & ~n24086 ;
  assign n24134 = \core_dag_ilm1reg_I2_we_DO_reg[12]/NET0131  & n6084 ;
  assign n24135 = ~n24133 & ~n24134 ;
  assign n24136 = ~n6084 & ~n24091 ;
  assign n24137 = ~n8734 & ~n24136 ;
  assign n24138 = n7340 & ~n23865 ;
  assign n24139 = \sport1_txctl_TX_reg[13]/P0001  & n23865 ;
  assign n24140 = ~n24138 & ~n24139 ;
  assign n24141 = ~n6106 & ~n7622 ;
  assign n24142 = n6106 & n7607 ;
  assign n24143 = ~n24141 & ~n24142 ;
  assign n24144 = ~n6084 & ~n24143 ;
  assign n24145 = \core_dag_ilm1reg_I2_we_DO_reg[0]/NET0131  & n6084 ;
  assign n24146 = ~n24144 & ~n24145 ;
  assign n24147 = ~n6067 & n24062 ;
  assign n24148 = ~n10402 & ~n24147 ;
  assign n24149 = \core_dag_ilm1reg_I1_we_DO_reg[5]/NET0131  & n6067 ;
  assign n24150 = ~n6067 & n24068 ;
  assign n24151 = ~n24149 & ~n24150 ;
  assign n24152 = ~n6067 & n24074 ;
  assign n24153 = ~n8891 & ~n24152 ;
  assign n24154 = \core_dag_ilm1reg_I1_we_DO_reg[13]/NET0131  & n6067 ;
  assign n24155 = ~n6067 & n24080 ;
  assign n24156 = ~n24154 & ~n24155 ;
  assign n24157 = ~n6067 & n24086 ;
  assign n24158 = ~\core_dag_ilm1reg_I1_we_DO_reg[12]/NET0131  & n6067 ;
  assign n24159 = ~n24157 & ~n24158 ;
  assign n24160 = ~n6067 & ~n24091 ;
  assign n24161 = ~n8736 & ~n24160 ;
  assign n24162 = ~n6067 & n23763 ;
  assign n24163 = ~n8135 & ~n24162 ;
  assign n24164 = ~n6058 & ~n24098 ;
  assign n24165 = ~n9718 & ~n24164 ;
  assign n24166 = \core_dag_ilm1reg_I0_we_DO_reg[8]/NET0131  & n6058 ;
  assign n24167 = ~n6058 & n24062 ;
  assign n24168 = ~n24166 & ~n24167 ;
  assign n24169 = ~n6058 & ~n24106 ;
  assign n24170 = \core_dag_ilm1reg_I0_we_DO_reg[7]/NET0131  & n6058 ;
  assign n24171 = ~n24169 & ~n24170 ;
  assign n24172 = ~n6058 & ~n24111 ;
  assign n24173 = \core_dag_ilm1reg_I0_we_DO_reg[6]/NET0131  & n6058 ;
  assign n24174 = ~n24172 & ~n24173 ;
  assign n24175 = ~n6058 & n24068 ;
  assign n24176 = ~n10369 & ~n24175 ;
  assign n24177 = ~n6058 & ~n24118 ;
  assign n24178 = ~n9771 & ~n24177 ;
  assign n24179 = ~n6058 & n23886 ;
  assign n24180 = ~n8186 & ~n24179 ;
  assign n24181 = ~n6058 & ~n24124 ;
  assign n24182 = \core_dag_ilm1reg_I0_we_DO_reg[2]/NET0131  & n6058 ;
  assign n24183 = ~n24181 & ~n24182 ;
  assign n24184 = ~n6058 & n24074 ;
  assign n24185 = ~n8888 & ~n24184 ;
  assign n24186 = ~n6058 & n24080 ;
  assign n24187 = ~n6136 & ~n24186 ;
  assign n24188 = ~n6058 & ~n24086 ;
  assign n24189 = ~n8859 & ~n24188 ;
  assign n24190 = \core_dag_ilm1reg_I0_we_DO_reg[11]/NET0131  & n6058 ;
  assign n24191 = ~n6058 & ~n24091 ;
  assign n24192 = ~n24190 & ~n24191 ;
  assign n24193 = \core_dag_ilm1reg_I0_we_DO_reg[10]/NET0131  & n6058 ;
  assign n24194 = ~n6058 & n23763 ;
  assign n24195 = ~n24193 & ~n24194 ;
  assign n24196 = ~n6058 & ~n24143 ;
  assign n24197 = ~n6936 & ~n24196 ;
  assign n24198 = ~n22114 & n23766 ;
  assign n24199 = ~\core_eu_em_mac_em_reg_my1swe_DO_reg[10]/P0001  & ~n23766 ;
  assign n24200 = ~n24198 & ~n24199 ;
  assign n24201 = ~n17836 & n23754 ;
  assign n24202 = ~\core_eu_es_sht_es_reg_siswe_DO_reg[13]/P0001  & ~n23754 ;
  assign n24203 = ~n24201 & ~n24202 ;
  assign n24204 = ~n19848 & n23754 ;
  assign n24205 = ~\core_eu_es_sht_es_reg_siswe_DO_reg[10]/P0001  & ~n23754 ;
  assign n24206 = ~n24204 & ~n24205 ;
  assign n24207 = \core_dag_ilm2reg_I7_we_DO_reg[4]/NET0131  & ~n23958 ;
  assign n24208 = ~n6000 & n20644 ;
  assign n24209 = ~n24207 & ~n24208 ;
  assign n24210 = \core_dag_ilm2reg_I7_we_DO_reg[3]/NET0131  & ~n23958 ;
  assign n24211 = ~n6000 & n13262 ;
  assign n24212 = ~n24210 & ~n24211 ;
  assign n24213 = \core_dag_ilm2reg_I7_we_DO_reg[2]/NET0131  & ~n23958 ;
  assign n24214 = ~n6000 & ~n20663 ;
  assign n24215 = ~n24213 & ~n24214 ;
  assign n24216 = \core_dag_ilm2reg_I7_we_DO_reg[1]/NET0131  & ~n23958 ;
  assign n24217 = ~n6000 & ~n20674 ;
  assign n24218 = ~n24216 & ~n24217 ;
  assign n24219 = \core_dag_ilm2reg_I7_we_DO_reg[0]/NET0131  & ~n23958 ;
  assign n24220 = ~n6000 & ~n20729 ;
  assign n24221 = ~n24219 & ~n24220 ;
  assign n24222 = ~n6008 & n20644 ;
  assign n24223 = \core_dag_ilm2reg_I6_we_DO_reg[4]/NET0131  & n6008 ;
  assign n24224 = ~n24222 & ~n24223 ;
  assign n24225 = ~n6008 & n13262 ;
  assign n24226 = \core_dag_ilm2reg_I6_we_DO_reg[3]/NET0131  & n6008 ;
  assign n24227 = ~n24225 & ~n24226 ;
  assign n24228 = ~n6008 & ~n20663 ;
  assign n24229 = \core_dag_ilm2reg_I6_we_DO_reg[2]/NET0131  & n6008 ;
  assign n24230 = ~n24228 & ~n24229 ;
  assign n24231 = ~n6008 & ~n20674 ;
  assign n24232 = \core_dag_ilm2reg_I6_we_DO_reg[1]/NET0131  & n6008 ;
  assign n24233 = ~n24231 & ~n24232 ;
  assign n24234 = ~n6008 & ~n20729 ;
  assign n24235 = \core_dag_ilm2reg_I6_we_DO_reg[0]/NET0131  & n6008 ;
  assign n24236 = ~n24234 & ~n24235 ;
  assign n24237 = \core_dag_ilm2reg_I5_we_DO_reg[4]/NET0131  & ~n24004 ;
  assign n24238 = ~n6015 & n20644 ;
  assign n24239 = ~n24237 & ~n24238 ;
  assign n24240 = \core_dag_ilm2reg_I5_we_DO_reg[3]/NET0131  & ~n24004 ;
  assign n24241 = ~n6015 & n13262 ;
  assign n24242 = ~n24240 & ~n24241 ;
  assign n24243 = \core_dag_ilm2reg_I5_we_DO_reg[2]/NET0131  & ~n24004 ;
  assign n24244 = ~n6015 & ~n20663 ;
  assign n24245 = ~n24243 & ~n24244 ;
  assign n24246 = \core_dag_ilm2reg_I5_we_DO_reg[1]/NET0131  & ~n24004 ;
  assign n24247 = ~n6015 & ~n20674 ;
  assign n24248 = ~n24246 & ~n24247 ;
  assign n24249 = \core_dag_ilm2reg_I5_we_DO_reg[0]/NET0131  & ~n24004 ;
  assign n24250 = ~n6015 & ~n20729 ;
  assign n24251 = ~n24249 & ~n24250 ;
  assign n24252 = \core_dag_ilm2reg_I4_we_DO_reg[4]/NET0131  & ~n24023 ;
  assign n24253 = ~n5964 & n20644 ;
  assign n24254 = ~n24252 & ~n24253 ;
  assign n24255 = \core_dag_ilm2reg_I4_we_DO_reg[3]/NET0131  & ~n24023 ;
  assign n24256 = ~n5964 & n13262 ;
  assign n24257 = ~n24255 & ~n24256 ;
  assign n24258 = \core_dag_ilm2reg_I4_we_DO_reg[2]/NET0131  & ~n24023 ;
  assign n24259 = ~n5964 & ~n20663 ;
  assign n24260 = ~n24258 & ~n24259 ;
  assign n24261 = \core_dag_ilm2reg_I4_we_DO_reg[1]/NET0131  & ~n24023 ;
  assign n24262 = ~n5964 & ~n20674 ;
  assign n24263 = ~n24261 & ~n24262 ;
  assign n24264 = \core_dag_ilm2reg_I4_we_DO_reg[0]/NET0131  & ~n24023 ;
  assign n24265 = ~n5964 & ~n20729 ;
  assign n24266 = ~n24264 & ~n24265 ;
  assign n24267 = n23027 & n23407 ;
  assign n24268 = ~\sice_ICYC_clr_reg/NET0131  & \sice_SPC_reg[23]/P0001  ;
  assign n24269 = n23032 & n24268 ;
  assign n24270 = n24267 & n24269 ;
  assign n24271 = \core_c_psq_Iact_E_reg[9]/NET0131  & ~n19477 ;
  assign n24272 = ~\core_c_psq_Iflag_reg[10]/NET0131  & ~\core_c_psq_PCS_reg[3]/NET0131  ;
  assign n24273 = n19481 & n24272 ;
  assign n24274 = n19477 & n24273 ;
  assign n24275 = ~n24271 & ~n24274 ;
  assign n24276 = ~n22021 & n23782 ;
  assign n24277 = ~\core_eu_em_mac_em_reg_my1rwe_DO_reg[6]/P0001  & ~n23782 ;
  assign n24278 = ~n24276 & ~n24277 ;
  assign n24279 = \core_c_psq_lpstk_lps4x22_LPcell_reg[3][3]/P0001  & ~n4851 ;
  assign n24280 = \core_c_psq_PMOVL_regl_DO_reg[3]/NET0131  & n4851 ;
  assign n24281 = ~n24279 & ~n24280 ;
  assign n24282 = \core_c_psq_lpstk_lps4x22_LPcell_reg[3][2]/P0001  & ~n4851 ;
  assign n24283 = \core_c_psq_PMOVL_regl_DO_reg[2]/NET0131  & n4851 ;
  assign n24284 = ~n24282 & ~n24283 ;
  assign n24285 = \core_c_psq_lpstk_lps4x22_LPcell_reg[3][1]/P0001  & ~n4851 ;
  assign n24286 = \core_c_psq_PMOVL_regl_DO_reg[1]/NET0131  & n4851 ;
  assign n24287 = ~n24285 & ~n24286 ;
  assign n24288 = \core_c_psq_lpstk_lps4x22_LPcell_reg[3][0]/P0001  & ~n4851 ;
  assign n24289 = \core_c_psq_PMOVL_regl_DO_reg[0]/NET0131  & n4851 ;
  assign n24290 = ~n24288 & ~n24289 ;
  assign n24291 = \core_c_psq_lpstk_lps4x22_LPcell_reg[2][3]/P0001  & ~n4847 ;
  assign n24292 = \core_c_psq_PMOVL_regl_DO_reg[3]/NET0131  & n4847 ;
  assign n24293 = ~n24291 & ~n24292 ;
  assign n24294 = \core_c_psq_lpstk_lps4x22_LPcell_reg[2][1]/P0001  & ~n4847 ;
  assign n24295 = \core_c_psq_PMOVL_regl_DO_reg[1]/NET0131  & n4847 ;
  assign n24296 = ~n24294 & ~n24295 ;
  assign n24297 = \core_c_psq_lpstk_lps4x22_LPcell_reg[1][2]/P0001  & ~n4845 ;
  assign n24298 = \core_c_psq_PMOVL_regl_DO_reg[2]/NET0131  & n4845 ;
  assign n24299 = ~n24297 & ~n24298 ;
  assign n24300 = \core_c_psq_lpstk_lps4x22_LPcell_reg[1][0]/P0001  & ~n4845 ;
  assign n24301 = \core_c_psq_PMOVL_regl_DO_reg[0]/NET0131  & n4845 ;
  assign n24302 = ~n24300 & ~n24301 ;
  assign n24303 = \core_c_psq_lpstk_lps4x22_LPcell_reg[0][3]/P0001  & ~n4849 ;
  assign n24304 = \core_c_psq_PMOVL_regl_DO_reg[3]/NET0131  & n4849 ;
  assign n24305 = ~n24303 & ~n24304 ;
  assign n24306 = \core_c_psq_lpstk_lps4x22_LPcell_reg[0][2]/P0001  & ~n4849 ;
  assign n24307 = \core_c_psq_PMOVL_regl_DO_reg[2]/NET0131  & n4849 ;
  assign n24308 = ~n24306 & ~n24307 ;
  assign n24309 = \core_c_psq_lpstk_lps4x22_LPcell_reg[0][1]/P0001  & ~n4849 ;
  assign n24310 = \core_c_psq_PMOVL_regl_DO_reg[1]/NET0131  & n4849 ;
  assign n24311 = ~n24309 & ~n24310 ;
  assign n24312 = \core_c_psq_lpstk_lps4x22_LPcell_reg[2][2]/P0001  & ~n4847 ;
  assign n24313 = \core_c_psq_PMOVL_regl_DO_reg[2]/NET0131  & n4847 ;
  assign n24314 = ~n24312 & ~n24313 ;
  assign n24315 = \core_c_psq_cntstk_cnts4x14_CNTcell_reg[3][8]/P0001  & ~n13794 ;
  assign n24316 = \core_c_psq_CNTR_reg_DO_reg[8]/NET0131  & n13794 ;
  assign n24317 = ~n24315 & ~n24316 ;
  assign n24318 = \core_c_psq_cntstk_cnts4x14_CNTcell_reg[3][7]/P0001  & ~n13794 ;
  assign n24319 = \core_c_psq_CNTR_reg_DO_reg[7]/NET0131  & n13794 ;
  assign n24320 = ~n24318 & ~n24319 ;
  assign n24321 = \core_c_psq_cntstk_cnts4x14_CNTcell_reg[3][6]/P0001  & ~n13794 ;
  assign n24322 = \core_c_psq_CNTR_reg_DO_reg[6]/NET0131  & n13794 ;
  assign n24323 = ~n24321 & ~n24322 ;
  assign n24324 = \core_c_psq_cntstk_cnts4x14_CNTcell_reg[3][4]/P0001  & ~n13794 ;
  assign n24325 = \core_c_psq_CNTR_reg_DO_reg[4]/NET0131  & n13794 ;
  assign n24326 = ~n24324 & ~n24325 ;
  assign n24327 = \core_c_psq_cntstk_cnts4x14_CNTcell_reg[3][3]/P0001  & ~n13794 ;
  assign n24328 = \core_c_psq_CNTR_reg_DO_reg[3]/NET0131  & n13794 ;
  assign n24329 = ~n24327 & ~n24328 ;
  assign n24330 = \core_c_psq_cntstk_cnts4x14_CNTcell_reg[3][2]/P0001  & ~n13794 ;
  assign n24331 = \core_c_psq_CNTR_reg_DO_reg[2]/NET0131  & n13794 ;
  assign n24332 = ~n24330 & ~n24331 ;
  assign n24333 = \core_c_psq_cntstk_cnts4x14_CNTcell_reg[3][13]/P0001  & ~n13794 ;
  assign n24334 = \core_c_psq_CNTR_reg_DO_reg[13]/NET0131  & n13794 ;
  assign n24335 = ~n24333 & ~n24334 ;
  assign n24336 = \core_c_psq_cntstk_cnts4x14_CNTcell_reg[3][12]/P0001  & ~n13794 ;
  assign n24337 = \core_c_psq_CNTR_reg_DO_reg[12]/NET0131  & n13794 ;
  assign n24338 = ~n24336 & ~n24337 ;
  assign n24339 = \core_c_psq_cntstk_cnts4x14_CNTcell_reg[3][11]/P0001  & ~n13794 ;
  assign n24340 = \core_c_psq_CNTR_reg_DO_reg[11]/NET0131  & n13794 ;
  assign n24341 = ~n24339 & ~n24340 ;
  assign n24342 = \core_c_psq_cntstk_cnts4x14_CNTcell_reg[3][10]/P0001  & ~n13794 ;
  assign n24343 = \core_c_psq_CNTR_reg_DO_reg[10]/NET0131  & n13794 ;
  assign n24344 = ~n24342 & ~n24343 ;
  assign n24345 = \core_c_psq_cntstk_cnts4x14_CNTcell_reg[3][0]/P0001  & ~n13794 ;
  assign n24346 = \core_c_psq_CNTR_reg_DO_reg[0]/NET0131  & n13794 ;
  assign n24347 = ~n24345 & ~n24346 ;
  assign n24348 = \core_c_psq_cntstk_cnts4x14_CNTcell_reg[2][6]/P0001  & ~n13789 ;
  assign n24349 = \core_c_psq_CNTR_reg_DO_reg[6]/NET0131  & n13789 ;
  assign n24350 = ~n24348 & ~n24349 ;
  assign n24351 = \core_c_psq_cntstk_cnts4x14_CNTcell_reg[2][3]/P0001  & ~n13789 ;
  assign n24352 = \core_c_psq_CNTR_reg_DO_reg[3]/NET0131  & n13789 ;
  assign n24353 = ~n24351 & ~n24352 ;
  assign n24354 = \core_c_psq_cntstk_cnts4x14_CNTcell_reg[2][2]/P0001  & ~n13789 ;
  assign n24355 = \core_c_psq_CNTR_reg_DO_reg[2]/NET0131  & n13789 ;
  assign n24356 = ~n24354 & ~n24355 ;
  assign n24357 = \core_c_psq_cntstk_cnts4x14_CNTcell_reg[2][13]/P0001  & ~n13789 ;
  assign n24358 = \core_c_psq_CNTR_reg_DO_reg[13]/NET0131  & n13789 ;
  assign n24359 = ~n24357 & ~n24358 ;
  assign n24360 = \core_c_psq_cntstk_cnts4x14_CNTcell_reg[2][11]/P0001  & ~n13789 ;
  assign n24361 = \core_c_psq_CNTR_reg_DO_reg[11]/NET0131  & n13789 ;
  assign n24362 = ~n24360 & ~n24361 ;
  assign n24363 = \core_c_psq_cntstk_cnts4x14_CNTcell_reg[2][0]/P0001  & ~n13789 ;
  assign n24364 = \core_c_psq_CNTR_reg_DO_reg[0]/NET0131  & n13789 ;
  assign n24365 = ~n24363 & ~n24364 ;
  assign n24366 = \core_c_psq_cntstk_cnts4x14_CNTcell_reg[1][8]/P0001  & ~n13784 ;
  assign n24367 = \core_c_psq_CNTR_reg_DO_reg[8]/NET0131  & n13784 ;
  assign n24368 = ~n24366 & ~n24367 ;
  assign n24369 = \core_c_psq_cntstk_cnts4x14_CNTcell_reg[1][7]/P0001  & ~n13784 ;
  assign n24370 = \core_c_psq_CNTR_reg_DO_reg[7]/NET0131  & n13784 ;
  assign n24371 = ~n24369 & ~n24370 ;
  assign n24372 = \core_c_psq_cntstk_cnts4x14_CNTcell_reg[1][6]/P0001  & ~n13784 ;
  assign n24373 = \core_c_psq_CNTR_reg_DO_reg[6]/NET0131  & n13784 ;
  assign n24374 = ~n24372 & ~n24373 ;
  assign n24375 = \core_c_psq_cntstk_cnts4x14_CNTcell_reg[1][3]/P0001  & ~n13784 ;
  assign n24376 = \core_c_psq_CNTR_reg_DO_reg[3]/NET0131  & n13784 ;
  assign n24377 = ~n24375 & ~n24376 ;
  assign n24378 = \core_c_psq_cntstk_cnts4x14_CNTcell_reg[1][2]/P0001  & ~n13784 ;
  assign n24379 = \core_c_psq_CNTR_reg_DO_reg[2]/NET0131  & n13784 ;
  assign n24380 = ~n24378 & ~n24379 ;
  assign n24381 = \core_c_psq_cntstk_cnts4x14_CNTcell_reg[1][1]/P0001  & ~n13784 ;
  assign n24382 = \core_c_psq_CNTR_reg_DO_reg[1]/NET0131  & n13784 ;
  assign n24383 = ~n24381 & ~n24382 ;
  assign n24384 = \core_c_psq_cntstk_cnts4x14_CNTcell_reg[1][13]/P0001  & ~n13784 ;
  assign n24385 = \core_c_psq_CNTR_reg_DO_reg[13]/NET0131  & n13784 ;
  assign n24386 = ~n24384 & ~n24385 ;
  assign n24387 = \core_c_psq_cntstk_cnts4x14_CNTcell_reg[1][11]/P0001  & ~n13784 ;
  assign n24388 = \core_c_psq_CNTR_reg_DO_reg[11]/NET0131  & n13784 ;
  assign n24389 = ~n24387 & ~n24388 ;
  assign n24390 = \core_c_psq_cntstk_cnts4x14_CNTcell_reg[1][10]/P0001  & ~n13784 ;
  assign n24391 = \core_c_psq_CNTR_reg_DO_reg[10]/NET0131  & n13784 ;
  assign n24392 = ~n24390 & ~n24391 ;
  assign n24393 = \core_c_psq_cntstk_cnts4x14_CNTcell_reg[0][9]/P0001  & ~n13775 ;
  assign n24394 = \core_c_psq_CNTR_reg_DO_reg[9]/NET0131  & n13775 ;
  assign n24395 = ~n24393 & ~n24394 ;
  assign n24396 = ~n18276 & n23754 ;
  assign n24397 = ~\core_eu_es_sht_es_reg_siswe_DO_reg[6]/P0001  & ~n23754 ;
  assign n24398 = ~n24396 & ~n24397 ;
  assign n24399 = ~n22048 & n23814 ;
  assign n24400 = ~\core_eu_em_mac_em_reg_my0rwe_DO_reg[3]/P0001  & ~n23814 ;
  assign n24401 = ~n24399 & ~n24400 ;
  assign n24402 = \core_c_dec_MTPMOVL_E_reg/P0001  & n5951 ;
  assign n24403 = n7607 & n8113 ;
  assign n24404 = n8715 & n9435 ;
  assign n24405 = n24403 & n24404 ;
  assign n24406 = n24402 & ~n24405 ;
  assign n24407 = ~\core_c_psq_PMOVL_regl_DO_reg[3]/NET0131  & ~n24406 ;
  assign n24408 = ~n8113 & n24402 ;
  assign n24409 = ~n24407 & ~n24408 ;
  assign n24410 = ~\core_c_psq_PMOVL_regl_DO_reg[2]/NET0131  & ~n24406 ;
  assign n24411 = ~n8715 & n24402 ;
  assign n24412 = ~n24410 & ~n24411 ;
  assign n24413 = ~n9435 & n24406 ;
  assign n24414 = ~\core_c_psq_PMOVL_regl_DO_reg[1]/NET0131  & ~n24406 ;
  assign n24415 = ~n24413 & ~n24414 ;
  assign n24416 = ~n7607 & n24406 ;
  assign n24417 = ~\core_c_psq_PMOVL_regl_DO_reg[0]/NET0131  & ~n24406 ;
  assign n24418 = ~n24416 & ~n24417 ;
  assign n24419 = n10069 & n10911 ;
  assign n24420 = n11265 & n24419 ;
  assign n24421 = n11525 & n24420 ;
  assign n24422 = n24402 & ~n24421 ;
  assign n24423 = ~\core_c_psq_PMOVL_regh_DO_reg[3]/NET0131  & ~n24422 ;
  assign n24424 = ~n11265 & n24402 ;
  assign n24425 = ~n24423 & ~n24424 ;
  assign n24426 = ~n11525 & n24422 ;
  assign n24427 = ~\core_c_psq_PMOVL_regh_DO_reg[2]/NET0131  & ~n24422 ;
  assign n24428 = ~n24426 & ~n24427 ;
  assign n24429 = ~\core_c_psq_PMOVL_regh_DO_reg[1]/NET0131  & ~n24422 ;
  assign n24430 = ~n10911 & n24402 ;
  assign n24431 = ~n24429 & ~n24430 ;
  assign n24432 = ~n19972 & n23754 ;
  assign n24433 = ~\core_eu_es_sht_es_reg_siswe_DO_reg[7]/P0001  & ~n23754 ;
  assign n24434 = ~n24432 & ~n24433 ;
  assign n24435 = \core_c_psq_cntstk_cnts4x14_CNTcell_reg[1][4]/P0001  & ~n13784 ;
  assign n24436 = \core_c_psq_CNTR_reg_DO_reg[4]/NET0131  & n13784 ;
  assign n24437 = ~n24435 & ~n24436 ;
  assign n24438 = \core_c_psq_cntstk_cnts4x14_CNTcell_reg[0][11]/P0001  & ~n13775 ;
  assign n24439 = \core_c_psq_CNTR_reg_DO_reg[11]/NET0131  & n13775 ;
  assign n24440 = ~n24438 & ~n24439 ;
  assign n24441 = n6117 & n13576 ;
  assign n24442 = ~n6107 & ~n24441 ;
  assign n24443 = ~n4117 & n24442 ;
  assign n24444 = ~\core_c_dec_imm16_E_reg/P0001  & n4117 ;
  assign n24445 = ~n24443 & ~n24444 ;
  assign n24446 = ~n10069 & n24422 ;
  assign n24447 = ~\core_c_psq_PMOVL_regh_DO_reg[0]/NET0131  & ~n24422 ;
  assign n24448 = ~n24446 & ~n24447 ;
  assign n24449 = \core_c_psq_lpstk_lps4x22_LPcell_reg[2][0]/P0001  & ~n4847 ;
  assign n24450 = \core_c_psq_PMOVL_regl_DO_reg[0]/NET0131  & n4847 ;
  assign n24451 = ~n24449 & ~n24450 ;
  assign n24452 = \core_c_psq_cntstk_cnts4x14_CNTcell_reg[0][12]/P0001  & ~n13775 ;
  assign n24453 = \core_c_psq_CNTR_reg_DO_reg[12]/NET0131  & n13775 ;
  assign n24454 = ~n24452 & ~n24453 ;
  assign n24455 = \core_c_psq_lpstk_lps4x22_LPcell_reg[0][0]/P0001  & ~n4849 ;
  assign n24456 = \core_c_psq_PMOVL_regl_DO_reg[0]/NET0131  & n4849 ;
  assign n24457 = ~n24455 & ~n24456 ;
  assign n24458 = ~n22012 & n23766 ;
  assign n24459 = ~\core_eu_em_mac_em_reg_my1swe_DO_reg[7]/P0001  & ~n23766 ;
  assign n24460 = ~n24458 & ~n24459 ;
  assign n24461 = ~n22021 & n23766 ;
  assign n24462 = ~\core_eu_em_mac_em_reg_my1swe_DO_reg[6]/P0001  & ~n23766 ;
  assign n24463 = ~n24461 & ~n24462 ;
  assign n24464 = ~n22030 & n23766 ;
  assign n24465 = ~\core_eu_em_mac_em_reg_my1swe_DO_reg[5]/P0001  & ~n23766 ;
  assign n24466 = ~n24464 & ~n24465 ;
  assign n24467 = ~n22039 & n23766 ;
  assign n24468 = ~\core_eu_em_mac_em_reg_my1swe_DO_reg[4]/P0001  & ~n23766 ;
  assign n24469 = ~n24467 & ~n24468 ;
  assign n24470 = ~n22048 & n23766 ;
  assign n24471 = ~\core_eu_em_mac_em_reg_my1swe_DO_reg[3]/P0001  & ~n23766 ;
  assign n24472 = ~n24470 & ~n24471 ;
  assign n24473 = ~n22057 & n23766 ;
  assign n24474 = ~\core_eu_em_mac_em_reg_my1swe_DO_reg[2]/P0001  & ~n23766 ;
  assign n24475 = ~n24473 & ~n24474 ;
  assign n24476 = ~n22151 & n23766 ;
  assign n24477 = ~\core_eu_em_mac_em_reg_my1swe_DO_reg[1]/P0001  & ~n23766 ;
  assign n24478 = ~n24476 & ~n24477 ;
  assign n24479 = ~n22066 & n23766 ;
  assign n24480 = ~\core_eu_em_mac_em_reg_my1swe_DO_reg[15]/P0001  & ~n23766 ;
  assign n24481 = ~n24479 & ~n24480 ;
  assign n24482 = ~n22075 & n23766 ;
  assign n24483 = ~\core_eu_em_mac_em_reg_my1swe_DO_reg[14]/P0001  & ~n23766 ;
  assign n24484 = ~n24482 & ~n24483 ;
  assign n24485 = ~n22012 & n23782 ;
  assign n24486 = ~\core_eu_em_mac_em_reg_my1rwe_DO_reg[7]/P0001  & ~n23782 ;
  assign n24487 = ~n24485 & ~n24486 ;
  assign n24488 = ~n22039 & n23782 ;
  assign n24489 = ~\core_eu_em_mac_em_reg_my1rwe_DO_reg[4]/P0001  & ~n23782 ;
  assign n24490 = ~n24488 & ~n24489 ;
  assign n24491 = ~n22048 & n23782 ;
  assign n24492 = ~\core_eu_em_mac_em_reg_my1rwe_DO_reg[3]/P0001  & ~n23782 ;
  assign n24493 = ~n24491 & ~n24492 ;
  assign n24494 = ~n22151 & n23782 ;
  assign n24495 = ~\core_eu_em_mac_em_reg_my1rwe_DO_reg[1]/P0001  & ~n23782 ;
  assign n24496 = ~n24494 & ~n24495 ;
  assign n24497 = ~n22066 & n23782 ;
  assign n24498 = ~\core_eu_em_mac_em_reg_my1rwe_DO_reg[15]/P0001  & ~n23782 ;
  assign n24499 = ~n24497 & ~n24498 ;
  assign n24500 = ~n22075 & n23782 ;
  assign n24501 = ~\core_eu_em_mac_em_reg_my1rwe_DO_reg[14]/P0001  & ~n23782 ;
  assign n24502 = ~n24500 & ~n24501 ;
  assign n24503 = ~n22039 & n23798 ;
  assign n24504 = ~\core_eu_em_mac_em_reg_my0swe_DO_reg[4]/P0001  & ~n23798 ;
  assign n24505 = ~n24503 & ~n24504 ;
  assign n24506 = ~n22021 & n23798 ;
  assign n24507 = ~\core_eu_em_mac_em_reg_my0swe_DO_reg[6]/P0001  & ~n23798 ;
  assign n24508 = ~n24506 & ~n24507 ;
  assign n24509 = ~n22048 & n23798 ;
  assign n24510 = ~\core_eu_em_mac_em_reg_my0swe_DO_reg[3]/P0001  & ~n23798 ;
  assign n24511 = ~n24509 & ~n24510 ;
  assign n24512 = ~n22151 & n23798 ;
  assign n24513 = ~\core_eu_em_mac_em_reg_my0swe_DO_reg[1]/P0001  & ~n23798 ;
  assign n24514 = ~n24512 & ~n24513 ;
  assign n24515 = ~n7607 & n21991 ;
  assign n24516 = ~n12520 & ~n21991 ;
  assign n24517 = ~n24515 & ~n24516 ;
  assign n24518 = n23798 & ~n24517 ;
  assign n24519 = ~\core_eu_em_mac_em_reg_my0swe_DO_reg[0]/P0001  & ~n23798 ;
  assign n24520 = ~n24518 & ~n24519 ;
  assign n24521 = ~n22012 & n23814 ;
  assign n24522 = ~\core_eu_em_mac_em_reg_my0rwe_DO_reg[7]/P0001  & ~n23814 ;
  assign n24523 = ~n24521 & ~n24522 ;
  assign n24524 = ~n22030 & n23814 ;
  assign n24525 = ~\core_eu_em_mac_em_reg_my0rwe_DO_reg[5]/P0001  & ~n23814 ;
  assign n24526 = ~n24524 & ~n24525 ;
  assign n24527 = ~n22039 & n23814 ;
  assign n24528 = ~\core_eu_em_mac_em_reg_my0rwe_DO_reg[4]/P0001  & ~n23814 ;
  assign n24529 = ~n24527 & ~n24528 ;
  assign n24530 = ~n22057 & n23814 ;
  assign n24531 = ~\core_eu_em_mac_em_reg_my0rwe_DO_reg[2]/P0001  & ~n23814 ;
  assign n24532 = ~n24530 & ~n24531 ;
  assign n24533 = \core_c_psq_lpstk_lps4x22_LPcell_reg[1][3]/P0001  & ~n4845 ;
  assign n24534 = \core_c_psq_PMOVL_regl_DO_reg[3]/NET0131  & n4845 ;
  assign n24535 = ~n24533 & ~n24534 ;
  assign n24536 = ~n22075 & n23814 ;
  assign n24537 = ~\core_eu_em_mac_em_reg_my0rwe_DO_reg[14]/P0001  & ~n23814 ;
  assign n24538 = ~n24536 & ~n24537 ;
  assign n24539 = n23814 & ~n24517 ;
  assign n24540 = ~\core_eu_em_mac_em_reg_my0rwe_DO_reg[0]/P0001  & ~n23814 ;
  assign n24541 = ~n24539 & ~n24540 ;
  assign n24542 = \core_c_psq_cntstk_cnts4x14_CNTcell_reg[1][9]/P0001  & ~n13784 ;
  assign n24543 = \core_c_psq_CNTR_reg_DO_reg[9]/NET0131  & n13784 ;
  assign n24544 = ~n24542 & ~n24543 ;
  assign n24545 = ~n11265 & n23827 ;
  assign n24546 = ~\bdma_BOVL_reg[7]/NET0131  & ~n23827 ;
  assign n24547 = ~n24545 & ~n24546 ;
  assign n24548 = ~n11525 & n23827 ;
  assign n24549 = ~\bdma_BOVL_reg[6]/NET0131  & ~n23827 ;
  assign n24550 = ~n24548 & ~n24549 ;
  assign n24551 = ~n10911 & n23827 ;
  assign n24552 = ~\bdma_BOVL_reg[5]/NET0131  & ~n23827 ;
  assign n24553 = ~n24551 & ~n24552 ;
  assign n24554 = ~n10069 & n23827 ;
  assign n24555 = ~\bdma_BOVL_reg[4]/NET0131  & ~n23827 ;
  assign n24556 = ~n24554 & ~n24555 ;
  assign n24557 = ~n8113 & n23827 ;
  assign n24558 = ~\bdma_BOVL_reg[3]/NET0131  & ~n23827 ;
  assign n24559 = ~n24557 & ~n24558 ;
  assign n24560 = ~n8715 & n23827 ;
  assign n24561 = ~\bdma_BOVL_reg[2]/NET0131  & ~n23827 ;
  assign n24562 = ~n24560 & ~n24561 ;
  assign n24563 = ~n9435 & n23827 ;
  assign n24564 = ~\bdma_BOVL_reg[1]/NET0131  & ~n23827 ;
  assign n24565 = ~n24563 & ~n24564 ;
  assign n24566 = ~n7607 & n23827 ;
  assign n24567 = ~\bdma_BOVL_reg[0]/NET0131  & ~n23827 ;
  assign n24568 = ~n24566 & ~n24567 ;
  assign n24569 = ~n8113 & n21268 ;
  assign n24570 = ~\bdma_BCTL_reg[3]/NET0131  & ~n21268 ;
  assign n24571 = ~n24569 & ~n24570 ;
  assign n24572 = ~n8715 & n21268 ;
  assign n24573 = ~\bdma_BCTL_reg[2]/NET0131  & ~n21268 ;
  assign n24574 = ~n24572 & ~n24573 ;
  assign n24575 = ~n9435 & n21268 ;
  assign n24576 = ~\bdma_BCTL_reg[1]/NET0131  & ~n21268 ;
  assign n24577 = ~n24575 & ~n24576 ;
  assign n24578 = ~n12743 & n21268 ;
  assign n24579 = ~\bdma_BCTL_reg[15]/NET0131  & ~n21268 ;
  assign n24580 = ~n24578 & ~n24579 ;
  assign n24581 = ~n12688 & n21268 ;
  assign n24582 = ~\bdma_BCTL_reg[14]/NET0131  & ~n21268 ;
  assign n24583 = ~n24581 & ~n24582 ;
  assign n24584 = ~n7607 & n21268 ;
  assign n24585 = ~\bdma_BCTL_reg[0]/NET0131  & ~n21268 ;
  assign n24586 = ~n24584 & ~n24585 ;
  assign n24587 = \core_c_psq_cntstk_cnts4x14_CNTcell_reg[2][10]/P0001  & ~n13789 ;
  assign n24588 = \core_c_psq_CNTR_reg_DO_reg[10]/NET0131  & n13789 ;
  assign n24589 = ~n24587 & ~n24588 ;
  assign n24590 = \core_c_psq_cntstk_cnts4x14_CNTcell_reg[2][12]/P0001  & ~n13789 ;
  assign n24591 = \core_c_psq_CNTR_reg_DO_reg[12]/NET0131  & n13789 ;
  assign n24592 = ~n24590 & ~n24591 ;
  assign n24593 = \core_c_psq_cntstk_cnts4x14_CNTcell_reg[0][13]/P0001  & ~n13775 ;
  assign n24594 = \core_c_psq_CNTR_reg_DO_reg[13]/NET0131  & n13775 ;
  assign n24595 = ~n24593 & ~n24594 ;
  assign n24596 = ~\sice_ICYC_reg[5]/NET0131  & ~n18859 ;
  assign n24597 = ~n18860 & ~n24596 ;
  assign n24598 = \core_c_psq_lpstk_lps4x22_LPcell_reg[1][1]/P0001  & ~n4845 ;
  assign n24599 = \core_c_psq_PMOVL_regl_DO_reg[1]/NET0131  & n4845 ;
  assign n24600 = ~n24598 & ~n24599 ;
  assign n24601 = \core_c_psq_cntstk_cnts4x14_CNTcell_reg[2][1]/P0001  & ~n13789 ;
  assign n24602 = \core_c_psq_CNTR_reg_DO_reg[1]/NET0131  & n13789 ;
  assign n24603 = ~n24601 & ~n24602 ;
  assign n24604 = \core_c_psq_cntstk_cnts4x14_CNTcell_reg[2][4]/P0001  & ~n13789 ;
  assign n24605 = \core_c_psq_CNTR_reg_DO_reg[4]/NET0131  & n13789 ;
  assign n24606 = ~n24604 & ~n24605 ;
  assign n24607 = n23766 & ~n24517 ;
  assign n24608 = ~\core_eu_em_mac_em_reg_my1swe_DO_reg[0]/P0001  & ~n23766 ;
  assign n24609 = ~n24607 & ~n24608 ;
  assign n24610 = \core_c_psq_cntstk_cnts4x14_CNTcell_reg[0][10]/P0001  & ~n13775 ;
  assign n24611 = \core_c_psq_CNTR_reg_DO_reg[10]/NET0131  & n13775 ;
  assign n24612 = ~n24610 & ~n24611 ;
  assign n24613 = \core_c_psq_cntstk_cnts4x14_CNTcell_reg[0][1]/P0001  & ~n13775 ;
  assign n24614 = \core_c_psq_CNTR_reg_DO_reg[1]/NET0131  & n13775 ;
  assign n24615 = ~n24613 & ~n24614 ;
  assign n24616 = \core_c_psq_cntstk_cnts4x14_CNTcell_reg[2][7]/P0001  & ~n13789 ;
  assign n24617 = \core_c_psq_CNTR_reg_DO_reg[7]/NET0131  & n13789 ;
  assign n24618 = ~n24616 & ~n24617 ;
  assign n24619 = \core_c_psq_cntstk_cnts4x14_CNTcell_reg[2][8]/P0001  & ~n13789 ;
  assign n24620 = \core_c_psq_CNTR_reg_DO_reg[8]/NET0131  & n13789 ;
  assign n24621 = ~n24619 & ~n24620 ;
  assign n24622 = \core_c_psq_cntstk_cnts4x14_CNTcell_reg[0][7]/P0001  & ~n13775 ;
  assign n24623 = \core_c_psq_CNTR_reg_DO_reg[7]/NET0131  & n13775 ;
  assign n24624 = ~n24622 & ~n24623 ;
  assign n24625 = \core_c_psq_cntstk_cnts4x14_CNTcell_reg[2][9]/P0001  & ~n13789 ;
  assign n24626 = \core_c_psq_CNTR_reg_DO_reg[9]/NET0131  & n13789 ;
  assign n24627 = ~n24625 & ~n24626 ;
  assign n24628 = ~n20150 & n23754 ;
  assign n24629 = ~\core_eu_es_sht_es_reg_siswe_DO_reg[14]/P0001  & ~n23754 ;
  assign n24630 = ~n24628 & ~n24629 ;
  assign n24631 = ~n17814 & n23754 ;
  assign n24632 = ~\core_eu_es_sht_es_reg_siswe_DO_reg[2]/P0001  & ~n23754 ;
  assign n24633 = ~n24631 & ~n24632 ;
  assign n24634 = \core_c_psq_cntstk_cnts4x14_CNTcell_reg[0][8]/P0001  & ~n13775 ;
  assign n24635 = \core_c_psq_CNTR_reg_DO_reg[8]/NET0131  & n13775 ;
  assign n24636 = ~n24634 & ~n24635 ;
  assign n24637 = ~n18974 & n23754 ;
  assign n24638 = ~\core_eu_es_sht_es_reg_siswe_DO_reg[1]/P0001  & ~n23754 ;
  assign n24639 = ~n24637 & ~n24638 ;
  assign n24640 = \core_c_psq_cntstk_cnts4x14_CNTcell_reg[0][2]/P0001  & ~n13775 ;
  assign n24641 = \core_c_psq_CNTR_reg_DO_reg[2]/NET0131  & n13775 ;
  assign n24642 = ~n24640 & ~n24641 ;
  assign n24643 = \memc_Dwrite_E_reg/NET0131  & n4117 ;
  assign n24645 = \core_c_dec_IR_reg[15]/NET0131  & n6120 ;
  assign n24646 = \core_c_dec_IR_reg[19]/NET0131  & n6108 ;
  assign n24644 = \core_c_dec_IR_reg[20]/NET0131  & n6956 ;
  assign n24647 = ~n6107 & ~n24644 ;
  assign n24648 = ~n24646 & n24647 ;
  assign n24649 = ~n24645 & n24648 ;
  assign n24650 = n11742 & ~n24649 ;
  assign n24651 = ~n24643 & ~n24650 ;
  assign n24652 = \core_c_psq_cntstk_cnts4x14_CNTcell_reg[3][1]/P0001  & ~n13794 ;
  assign n24653 = \core_c_psq_CNTR_reg_DO_reg[1]/NET0131  & n13794 ;
  assign n24654 = ~n24652 & ~n24653 ;
  assign n24655 = ~n21663 & n23754 ;
  assign n24656 = ~\core_eu_es_sht_es_reg_siswe_DO_reg[3]/P0001  & ~n23754 ;
  assign n24657 = ~n24655 & ~n24656 ;
  assign n24658 = \core_c_psq_cntstk_cnts4x14_CNTcell_reg[1][12]/P0001  & ~n13784 ;
  assign n24659 = \core_c_psq_CNTR_reg_DO_reg[12]/NET0131  & n13784 ;
  assign n24660 = ~n24658 & ~n24659 ;
  assign n24661 = n11265 & ~n23865 ;
  assign n24662 = \sport1_txctl_TX_reg[7]/P0001  & n23865 ;
  assign n24663 = ~n24661 & ~n24662 ;
  assign n24664 = \core_c_psq_cntstk_cnts4x14_CNTcell_reg[1][0]/P0001  & ~n13784 ;
  assign n24665 = \core_c_psq_CNTR_reg_DO_reg[0]/NET0131  & n13784 ;
  assign n24666 = ~n24664 & ~n24665 ;
  assign n24667 = n11525 & ~n23865 ;
  assign n24668 = \sport1_txctl_TX_reg[6]/P0001  & n23865 ;
  assign n24669 = ~n24667 & ~n24668 ;
  assign n24670 = n10911 & ~n23865 ;
  assign n24671 = \sport1_txctl_TX_reg[5]/P0001  & n23865 ;
  assign n24672 = ~n24670 & ~n24671 ;
  assign n24673 = n10069 & ~n23865 ;
  assign n24674 = \sport1_txctl_TX_reg[4]/P0001  & n23865 ;
  assign n24675 = ~n24673 & ~n24674 ;
  assign n24676 = n8113 & ~n23865 ;
  assign n24677 = \sport1_txctl_TX_reg[3]/P0001  & n23865 ;
  assign n24678 = ~n24676 & ~n24677 ;
  assign n24679 = n8715 & ~n23865 ;
  assign n24680 = \sport1_txctl_TX_reg[2]/P0001  & n23865 ;
  assign n24681 = ~n24679 & ~n24680 ;
  assign n24682 = n9435 & ~n23865 ;
  assign n24683 = \sport1_txctl_TX_reg[1]/P0001  & n23865 ;
  assign n24684 = ~n24682 & ~n24683 ;
  assign n24685 = n12743 & ~n23865 ;
  assign n24686 = \sport1_txctl_TX_reg[15]/P0001  & n23865 ;
  assign n24687 = ~n24685 & ~n24686 ;
  assign n24688 = n12688 & ~n23865 ;
  assign n24689 = \sport1_txctl_TX_reg[14]/P0001  & n23865 ;
  assign n24690 = ~n24688 & ~n24689 ;
  assign n24691 = n7607 & ~n23865 ;
  assign n24692 = \sport1_txctl_TX_reg[0]/P0001  & n23865 ;
  assign n24693 = ~n24691 & ~n24692 ;
  assign n24694 = ~n20080 & n23754 ;
  assign n24695 = ~\core_eu_es_sht_es_reg_siswe_DO_reg[4]/P0001  & ~n23754 ;
  assign n24696 = ~n24694 & ~n24695 ;
  assign n24697 = \core_c_psq_cntstk_cnts4x14_CNTcell_reg[0][3]/P0001  & ~n13775 ;
  assign n24698 = \core_c_psq_CNTR_reg_DO_reg[3]/NET0131  & n13775 ;
  assign n24699 = ~n24697 & ~n24698 ;
  assign n24700 = \core_c_psq_cntstk_cnts4x14_CNTcell_reg[0][4]/P0001  & ~n13775 ;
  assign n24701 = \core_c_psq_CNTR_reg_DO_reg[4]/NET0131  & n13775 ;
  assign n24702 = ~n24700 & ~n24701 ;
  assign n24703 = ~n22021 & n23814 ;
  assign n24704 = ~\core_eu_em_mac_em_reg_my0rwe_DO_reg[6]/P0001  & ~n23814 ;
  assign n24705 = ~n24703 & ~n24704 ;
  assign n24706 = ~n22030 & n23798 ;
  assign n24707 = ~\core_eu_em_mac_em_reg_my0swe_DO_reg[5]/P0001  & ~n23798 ;
  assign n24708 = ~n24706 & ~n24707 ;
  assign n24709 = \core_eu_ec_cun_updateMV_C_reg/P0001  & n5950 ;
  assign n24710 = ~n21314 & ~n24709 ;
  assign n24711 = \core_c_psq_MSTAT_reg_DO_reg[4]/NET0131  & ~n22924 ;
  assign n24712 = ~n22770 & ~n22776 ;
  assign n24713 = ~n22766 & ~n22772 ;
  assign n24714 = n22766 & n22772 ;
  assign n24715 = n22709 & ~n24714 ;
  assign n24716 = ~n24713 & ~n24715 ;
  assign n24717 = n24712 & ~n24716 ;
  assign n24718 = ~n24712 & n24716 ;
  assign n24719 = ~n24717 & ~n24718 ;
  assign n24720 = ~\core_c_psq_MSTAT_reg_DO_reg[4]/NET0131  & n24719 ;
  assign n24721 = ~n24711 & ~n24720 ;
  assign n24722 = ~n22012 & n23889 ;
  assign n24723 = ~\core_eu_ea_alu_ea_reg_ay1swe_DO_reg[7]/P0001  & ~n23889 ;
  assign n24724 = ~n24722 & ~n24723 ;
  assign n24725 = ~n22021 & n23889 ;
  assign n24726 = ~\core_eu_ea_alu_ea_reg_ay1swe_DO_reg[6]/P0001  & ~n23889 ;
  assign n24727 = ~n24725 & ~n24726 ;
  assign n24728 = ~n22030 & n23889 ;
  assign n24729 = ~\core_eu_ea_alu_ea_reg_ay1swe_DO_reg[5]/P0001  & ~n23889 ;
  assign n24730 = ~n24728 & ~n24729 ;
  assign n24731 = ~n22039 & n23889 ;
  assign n24732 = ~\core_eu_ea_alu_ea_reg_ay1swe_DO_reg[4]/P0001  & ~n23889 ;
  assign n24733 = ~n24731 & ~n24732 ;
  assign n24734 = ~n22048 & n23889 ;
  assign n24735 = ~\core_eu_ea_alu_ea_reg_ay1swe_DO_reg[3]/P0001  & ~n23889 ;
  assign n24736 = ~n24734 & ~n24735 ;
  assign n24737 = ~n22057 & n23889 ;
  assign n24738 = ~\core_eu_ea_alu_ea_reg_ay1swe_DO_reg[2]/P0001  & ~n23889 ;
  assign n24739 = ~n24737 & ~n24738 ;
  assign n24740 = ~n22151 & n23889 ;
  assign n24741 = ~\core_eu_ea_alu_ea_reg_ay1swe_DO_reg[1]/P0001  & ~n23889 ;
  assign n24742 = ~n24740 & ~n24741 ;
  assign n24743 = ~n22066 & n23889 ;
  assign n24744 = ~\core_eu_ea_alu_ea_reg_ay1swe_DO_reg[15]/P0001  & ~n23889 ;
  assign n24745 = ~n24743 & ~n24744 ;
  assign n24746 = ~n22075 & n23889 ;
  assign n24747 = ~\core_eu_ea_alu_ea_reg_ay1swe_DO_reg[14]/P0001  & ~n23889 ;
  assign n24748 = ~n24746 & ~n24747 ;
  assign n24749 = n23889 & ~n24517 ;
  assign n24750 = ~\core_eu_ea_alu_ea_reg_ay1swe_DO_reg[0]/P0001  & ~n23889 ;
  assign n24751 = ~n24749 & ~n24750 ;
  assign n24752 = ~n19972 & n23908 ;
  assign n24753 = ~\core_eu_ea_alu_ea_reg_ax1swe_DO_reg[7]/P0001  & ~n23908 ;
  assign n24754 = ~n24752 & ~n24753 ;
  assign n24755 = ~n18276 & n23908 ;
  assign n24756 = ~\core_eu_ea_alu_ea_reg_ax1swe_DO_reg[6]/P0001  & ~n23908 ;
  assign n24757 = ~n24755 & ~n24756 ;
  assign n24758 = ~n20259 & n23908 ;
  assign n24759 = ~\core_eu_ea_alu_ea_reg_ax1swe_DO_reg[5]/P0001  & ~n23908 ;
  assign n24760 = ~n24758 & ~n24759 ;
  assign n24761 = ~n20080 & n23908 ;
  assign n24762 = ~\core_eu_ea_alu_ea_reg_ax1swe_DO_reg[4]/P0001  & ~n23908 ;
  assign n24763 = ~n24761 & ~n24762 ;
  assign n24764 = ~n21663 & n23908 ;
  assign n24765 = ~\core_eu_ea_alu_ea_reg_ax1swe_DO_reg[3]/P0001  & ~n23908 ;
  assign n24766 = ~n24764 & ~n24765 ;
  assign n24767 = ~n17814 & n23908 ;
  assign n24768 = ~\core_eu_ea_alu_ea_reg_ax1swe_DO_reg[2]/P0001  & ~n23908 ;
  assign n24769 = ~n24767 & ~n24768 ;
  assign n24770 = ~n18974 & n23908 ;
  assign n24771 = ~\core_eu_ea_alu_ea_reg_ax1swe_DO_reg[1]/P0001  & ~n23908 ;
  assign n24772 = ~n24770 & ~n24771 ;
  assign n24773 = ~n17820 & n23908 ;
  assign n24774 = ~\core_eu_ea_alu_ea_reg_ax1swe_DO_reg[15]/P0001  & ~n23908 ;
  assign n24775 = ~n24773 & ~n24774 ;
  assign n24776 = ~n20150 & n23908 ;
  assign n24777 = ~\core_eu_ea_alu_ea_reg_ax1swe_DO_reg[14]/P0001  & ~n23908 ;
  assign n24778 = ~n24776 & ~n24777 ;
  assign n24779 = ~n19559 & n23908 ;
  assign n24780 = ~\core_eu_ea_alu_ea_reg_ax1swe_DO_reg[0]/P0001  & ~n23908 ;
  assign n24781 = ~n24779 & ~n24780 ;
  assign n24782 = ~n19972 & n23930 ;
  assign n24783 = ~\core_eu_ea_alu_ea_reg_ax0swe_DO_reg[7]/P0001  & ~n23930 ;
  assign n24784 = ~n24782 & ~n24783 ;
  assign n24785 = ~n18276 & n23930 ;
  assign n24786 = ~\core_eu_ea_alu_ea_reg_ax0swe_DO_reg[6]/P0001  & ~n23930 ;
  assign n24787 = ~n24785 & ~n24786 ;
  assign n24788 = ~n20259 & n23930 ;
  assign n24789 = ~\core_eu_ea_alu_ea_reg_ax0swe_DO_reg[5]/P0001  & ~n23930 ;
  assign n24790 = ~n24788 & ~n24789 ;
  assign n24791 = ~n20080 & n23930 ;
  assign n24792 = ~\core_eu_ea_alu_ea_reg_ax0swe_DO_reg[4]/P0001  & ~n23930 ;
  assign n24793 = ~n24791 & ~n24792 ;
  assign n24794 = ~n21663 & n23930 ;
  assign n24795 = ~\core_eu_ea_alu_ea_reg_ax0swe_DO_reg[3]/P0001  & ~n23930 ;
  assign n24796 = ~n24794 & ~n24795 ;
  assign n24797 = ~n17814 & n23930 ;
  assign n24798 = ~\core_eu_ea_alu_ea_reg_ax0swe_DO_reg[2]/P0001  & ~n23930 ;
  assign n24799 = ~n24797 & ~n24798 ;
  assign n24800 = ~n18974 & n23930 ;
  assign n24801 = ~\core_eu_ea_alu_ea_reg_ax0swe_DO_reg[1]/P0001  & ~n23930 ;
  assign n24802 = ~n24800 & ~n24801 ;
  assign n24803 = ~n17820 & n23930 ;
  assign n24804 = ~\core_eu_ea_alu_ea_reg_ax0swe_DO_reg[15]/P0001  & ~n23930 ;
  assign n24805 = ~n24803 & ~n24804 ;
  assign n24806 = ~n20150 & n23930 ;
  assign n24807 = ~\core_eu_ea_alu_ea_reg_ax0swe_DO_reg[14]/P0001  & ~n23930 ;
  assign n24808 = ~n24806 & ~n24807 ;
  assign n24809 = ~n19559 & n23930 ;
  assign n24810 = ~\core_eu_ea_alu_ea_reg_ax0swe_DO_reg[0]/P0001  & ~n23930 ;
  assign n24811 = ~n24809 & ~n24810 ;
  assign n24812 = ~n22066 & n23798 ;
  assign n24813 = ~\core_eu_em_mac_em_reg_my0swe_DO_reg[15]/P0001  & ~n23798 ;
  assign n24814 = ~n24812 & ~n24813 ;
  assign n24815 = n19698 & n21248 ;
  assign n24816 = n23231 & n24815 ;
  assign n24817 = \core_c_dec_Modctl_Eg_reg/P0001  & n4118 ;
  assign n24818 = ~n24816 & ~n24817 ;
  assign n24819 = ~n22066 & n23814 ;
  assign n24820 = ~\core_eu_em_mac_em_reg_my0rwe_DO_reg[15]/P0001  & ~n23814 ;
  assign n24821 = ~n24819 & ~n24820 ;
  assign n24822 = \core_c_psq_cntstk_cnts4x14_CNTcell_reg[0][0]/P0001  & ~n13775 ;
  assign n24823 = \core_c_psq_CNTR_reg_DO_reg[0]/NET0131  & n13775 ;
  assign n24824 = ~n24822 & ~n24823 ;
  assign n24825 = ~n22151 & n23814 ;
  assign n24826 = ~\core_eu_em_mac_em_reg_my0rwe_DO_reg[1]/P0001  & ~n23814 ;
  assign n24827 = ~n24825 & ~n24826 ;
  assign n24828 = \core_c_psq_cntstk_cnts4x14_CNTcell_reg[3][9]/P0001  & ~n13794 ;
  assign n24829 = \core_c_psq_CNTR_reg_DO_reg[9]/NET0131  & n13794 ;
  assign n24830 = ~n24828 & ~n24829 ;
  assign n24831 = ~n20259 & n23754 ;
  assign n24832 = ~\core_eu_es_sht_es_reg_siswe_DO_reg[5]/P0001  & ~n23754 ;
  assign n24833 = ~n24831 & ~n24832 ;
  assign n24834 = \core_c_psq_cntstk_cnts4x14_CNTcell_reg[0][6]/P0001  & ~n13775 ;
  assign n24835 = \core_c_psq_CNTR_reg_DO_reg[6]/NET0131  & n13775 ;
  assign n24836 = ~n24834 & ~n24835 ;
  assign n24837 = ~n22075 & n23798 ;
  assign n24838 = ~\core_eu_em_mac_em_reg_my0swe_DO_reg[14]/P0001  & ~n23798 ;
  assign n24839 = ~n24837 & ~n24838 ;
  assign n24840 = ~n22057 & n23798 ;
  assign n24841 = ~\core_eu_em_mac_em_reg_my0swe_DO_reg[2]/P0001  & ~n23798 ;
  assign n24842 = ~n24840 & ~n24841 ;
  assign n24843 = ~n22012 & n23798 ;
  assign n24844 = ~\core_eu_em_mac_em_reg_my0swe_DO_reg[7]/P0001  & ~n23798 ;
  assign n24845 = ~n24843 & ~n24844 ;
  assign n24846 = n23782 & ~n24517 ;
  assign n24847 = ~\core_eu_em_mac_em_reg_my1rwe_DO_reg[0]/P0001  & ~n23782 ;
  assign n24848 = ~n24846 & ~n24847 ;
  assign n24849 = ~n22057 & n23782 ;
  assign n24850 = ~\core_eu_em_mac_em_reg_my1rwe_DO_reg[2]/P0001  & ~n23782 ;
  assign n24851 = ~n24849 & ~n24850 ;
  assign n24852 = ~n17820 & n23754 ;
  assign n24853 = ~\core_eu_es_sht_es_reg_siswe_DO_reg[15]/P0001  & ~n23754 ;
  assign n24854 = ~n24852 & ~n24853 ;
  assign n24855 = ~n19559 & n23754 ;
  assign n24856 = ~\core_eu_es_sht_es_reg_siswe_DO_reg[0]/P0001  & ~n23754 ;
  assign n24857 = ~n24855 & ~n24856 ;
  assign n24858 = ~n22030 & n23782 ;
  assign n24859 = ~\core_eu_em_mac_em_reg_my1rwe_DO_reg[5]/P0001  & ~n23782 ;
  assign n24860 = ~n24858 & ~n24859 ;
  assign n24861 = \sice_IDONE_reg/NET0131  & n5950 ;
  assign n24862 = ~\core_c_dec_NOP_E_reg/P0001  & n19203 ;
  assign n24863 = ~n24861 & ~n24862 ;
  assign n24864 = ~\sice_IIRC_reg[2]/NET0131  & ~n18865 ;
  assign n24865 = ~n18866 & ~n24864 ;
  assign n24866 = ~\clkc_oscntr_reg_DO_reg[2]/NET0131  & n20845 ;
  assign n24867 = ~n20846 & ~n24866 ;
  assign n24868 = ~\sice_ICYC_reg[2]/NET0131  & ~n18856 ;
  assign n24869 = ~n18857 & ~n24868 ;
  assign n24870 = \core_c_dec_MTAY1_E_reg/P0001  & n17798 ;
  assign n24871 = ~n21994 & n24870 ;
  assign n24872 = ~\core_eu_ea_alu_ea_reg_ay1rwe_DO_reg[9]/P0001  & ~n24870 ;
  assign n24873 = ~n24871 & ~n24872 ;
  assign n24874 = \core_eu_ea_alu_ea_reg_ay1rwe_DO_reg[8]/P0001  & ~n24870 ;
  assign n24875 = ~n22003 & n24870 ;
  assign n24876 = ~n24874 & ~n24875 ;
  assign n24877 = ~n22012 & n24870 ;
  assign n24878 = ~\core_eu_ea_alu_ea_reg_ay1rwe_DO_reg[7]/P0001  & ~n24870 ;
  assign n24879 = ~n24877 & ~n24878 ;
  assign n24880 = ~n22021 & n24870 ;
  assign n24881 = ~\core_eu_ea_alu_ea_reg_ay1rwe_DO_reg[6]/P0001  & ~n24870 ;
  assign n24882 = ~n24880 & ~n24881 ;
  assign n24883 = ~n22030 & n24870 ;
  assign n24884 = ~\core_eu_ea_alu_ea_reg_ay1rwe_DO_reg[5]/P0001  & ~n24870 ;
  assign n24885 = ~n24883 & ~n24884 ;
  assign n24886 = ~n22039 & n24870 ;
  assign n24887 = ~\core_eu_ea_alu_ea_reg_ay1rwe_DO_reg[4]/P0001  & ~n24870 ;
  assign n24888 = ~n24886 & ~n24887 ;
  assign n24889 = ~n22048 & n24870 ;
  assign n24890 = ~\core_eu_ea_alu_ea_reg_ay1rwe_DO_reg[3]/P0001  & ~n24870 ;
  assign n24891 = ~n24889 & ~n24890 ;
  assign n24892 = ~n22057 & n24870 ;
  assign n24893 = ~\core_eu_ea_alu_ea_reg_ay1rwe_DO_reg[2]/P0001  & ~n24870 ;
  assign n24894 = ~n24892 & ~n24893 ;
  assign n24895 = ~n22151 & n24870 ;
  assign n24896 = ~\core_eu_ea_alu_ea_reg_ay1rwe_DO_reg[1]/P0001  & ~n24870 ;
  assign n24897 = ~n24895 & ~n24896 ;
  assign n24898 = ~n22066 & n24870 ;
  assign n24899 = ~\core_eu_ea_alu_ea_reg_ay1rwe_DO_reg[15]/P0001  & ~n24870 ;
  assign n24900 = ~n24898 & ~n24899 ;
  assign n24901 = ~n22075 & n24870 ;
  assign n24902 = ~\core_eu_ea_alu_ea_reg_ay1rwe_DO_reg[14]/P0001  & ~n24870 ;
  assign n24903 = ~n24901 & ~n24902 ;
  assign n24904 = ~n22084 & n24870 ;
  assign n24905 = ~\core_eu_ea_alu_ea_reg_ay1rwe_DO_reg[13]/P0001  & ~n24870 ;
  assign n24906 = ~n24904 & ~n24905 ;
  assign n24907 = \core_eu_ea_alu_ea_reg_ay1rwe_DO_reg[12]/P0001  & ~n24870 ;
  assign n24908 = ~n22093 & n24870 ;
  assign n24909 = ~n24907 & ~n24908 ;
  assign n24910 = \core_eu_ea_alu_ea_reg_ay1rwe_DO_reg[11]/P0001  & ~n24870 ;
  assign n24911 = ~n22105 & n24870 ;
  assign n24912 = ~n24910 & ~n24911 ;
  assign n24913 = ~n22114 & n24870 ;
  assign n24914 = ~\core_eu_ea_alu_ea_reg_ay1rwe_DO_reg[10]/P0001  & ~n24870 ;
  assign n24915 = ~n24913 & ~n24914 ;
  assign n24916 = ~n24517 & n24870 ;
  assign n24917 = ~\core_eu_ea_alu_ea_reg_ay1rwe_DO_reg[0]/P0001  & ~n24870 ;
  assign n24918 = ~n24916 & ~n24917 ;
  assign n24920 = n19499 & ~n23860 ;
  assign n24919 = ~\core_eu_em_mac_em_reg_mr1swe_DO_reg[8]/P0001  & ~n19499 ;
  assign n24921 = n19501 & ~n24919 ;
  assign n24922 = ~n24920 & n24921 ;
  assign n24923 = \core_eu_em_mac_em_reg_mr1swe_DO_reg[8]/P0001  & ~n19383 ;
  assign n24924 = ~n19508 & ~n24923 ;
  assign n24925 = ~n24922 & n24924 ;
  assign n24926 = ~n18262 & ~n24925 ;
  assign n24927 = ~\core_c_psq_MSTAT_reg_DO_reg[4]/NET0131  & n22948 ;
  assign n24928 = \core_c_psq_MSTAT_reg_DO_reg[4]/NET0131  & n19523 ;
  assign n24929 = ~n24927 & ~n24928 ;
  assign n24930 = n18262 & ~n24929 ;
  assign n24931 = ~n24926 & ~n24930 ;
  assign n24934 = ~\sport0_rxctl_ldRX_cmp_reg/P0001  & n8715 ;
  assign n24935 = ~\sport0_rxctl_RX_reg[7]/P0001  & ~n20954 ;
  assign n24937 = ~n20951 & n24935 ;
  assign n24936 = n20951 & ~n24935 ;
  assign n24938 = n20875 & ~n24936 ;
  assign n24939 = ~n24937 & n24938 ;
  assign n24933 = \sport0_rxctl_RX_reg[2]/P0001  & n20873 ;
  assign n24940 = ~n20868 & ~n24933 ;
  assign n24941 = ~n24939 & n24940 ;
  assign n24942 = ~n24934 & n24941 ;
  assign n24932 = ~\sport0_rxctl_RXSHT_reg[2]/P0001  & n20868 ;
  assign n24943 = ~n20871 & ~n24932 ;
  assign n24944 = ~n24942 & n24943 ;
  assign n24945 = \sport0_rxctl_RX_reg[2]/P0001  & n20871 ;
  assign n24946 = ~n24944 & ~n24945 ;
  assign n24948 = ~n17836 & n19499 ;
  assign n24947 = ~\core_eu_em_mac_em_reg_mr1swe_DO_reg[13]/P0001  & ~n19499 ;
  assign n24949 = n19501 & ~n24947 ;
  assign n24950 = ~n24948 & n24949 ;
  assign n24951 = \core_eu_em_mac_em_reg_mr1swe_DO_reg[13]/P0001  & ~n19383 ;
  assign n24952 = ~n19508 & ~n24951 ;
  assign n24953 = ~n24950 & n24952 ;
  assign n24954 = ~n18262 & ~n24953 ;
  assign n24955 = ~n17741 & ~n17770 ;
  assign n24956 = ~n17737 & ~n19414 ;
  assign n24957 = ~n19415 & ~n24956 ;
  assign n24958 = n24955 & n24957 ;
  assign n24959 = ~n24955 & ~n24957 ;
  assign n24960 = ~n24958 & ~n24959 ;
  assign n24961 = ~\core_c_psq_MSTAT_reg_DO_reg[4]/NET0131  & ~n24960 ;
  assign n24962 = \core_c_psq_MSTAT_reg_DO_reg[4]/NET0131  & n22996 ;
  assign n24963 = ~n24961 & ~n24962 ;
  assign n24964 = n18262 & ~n24963 ;
  assign n24965 = ~n24954 & ~n24964 ;
  assign n24966 = ~\clkc_oscntr_reg_DO_reg[5]/NET0131  & ~n23418 ;
  assign n24967 = ~n23419 & ~n24966 ;
  assign n24968 = \clkc_CTR_cnt_reg[0]/NET0131  & ~\clkc_CTR_cnt_reg[1]/NET0131  ;
  assign n24971 = n18271 & ~n21663 ;
  assign n24970 = ~\core_eu_em_mac_em_reg_mr0swe_DO_reg[3]/P0001  & ~n18271 ;
  assign n24972 = n18273 & ~n24970 ;
  assign n24973 = ~n24971 & n24972 ;
  assign n24969 = \core_eu_em_mac_em_reg_mr0swe_DO_reg[3]/P0001  & ~n18266 ;
  assign n24974 = ~n18270 & ~n24969 ;
  assign n24975 = ~n24973 & n24974 ;
  assign n24976 = ~n18262 & ~n24975 ;
  assign n24977 = n18262 & ~n19662 ;
  assign n24978 = ~n24976 & ~n24977 ;
  assign n24979 = n14752 & n19662 ;
  assign n24980 = n18328 & n21663 ;
  assign n24981 = \core_eu_em_mac_em_reg_mr0rwe_DO_reg[3]/P0001  & ~n18330 ;
  assign n24982 = n18334 & ~n24981 ;
  assign n24983 = ~n24980 & n24982 ;
  assign n24984 = ~n24979 & ~n24983 ;
  assign n24985 = ~n13806 & ~n14634 ;
  assign n24986 = n13806 & ~n14600 ;
  assign n24987 = ~n24985 & ~n24986 ;
  assign n24988 = n14667 & ~n24987 ;
  assign n24989 = \core_eu_ea_alu_ea_reg_afswe_DO_reg[5]/P0001  & ~n14667 ;
  assign n24990 = ~n24988 & ~n24989 ;
  assign n24991 = n13805 & ~n24987 ;
  assign n24992 = \core_eu_ea_alu_ea_reg_afrwe_DO_reg[5]/P0001  & ~n13805 ;
  assign n24993 = ~n24991 & ~n24992 ;
  assign n24995 = n19499 & ~n23920 ;
  assign n24994 = ~\core_eu_em_mac_em_reg_mr1swe_DO_reg[12]/P0001  & ~n19499 ;
  assign n24996 = n19501 & ~n24994 ;
  assign n24997 = ~n24995 & n24996 ;
  assign n24998 = \core_eu_em_mac_em_reg_mr1swe_DO_reg[12]/P0001  & ~n19383 ;
  assign n24999 = ~n19508 & ~n24998 ;
  assign n25000 = ~n24997 & n24999 ;
  assign n25001 = ~n18262 & ~n25000 ;
  assign n25002 = \core_c_psq_MSTAT_reg_DO_reg[4]/NET0131  & n24960 ;
  assign n25003 = ~\core_c_psq_MSTAT_reg_DO_reg[4]/NET0131  & n19419 ;
  assign n25004 = ~n25002 & ~n25003 ;
  assign n25005 = n18262 & n25004 ;
  assign n25006 = ~n25001 & ~n25005 ;
  assign n25007 = ~n6107 & ~n6956 ;
  assign n25008 = ~n6120 & n25007 ;
  assign n25009 = n18838 & n25008 ;
  assign n25010 = ~\sice_IAR_reg[1]/NET0131  & \sice_IAR_reg[2]/NET0131  ;
  assign n25011 = \sice_IAR_reg[0]/NET0131  & \sice_IAR_reg[3]/NET0131  ;
  assign n25012 = n25010 & n25011 ;
  assign n25013 = n23032 & n25012 ;
  assign n25014 = n14752 & n24929 ;
  assign n25015 = n19776 & n23860 ;
  assign n25016 = \core_eu_em_mac_em_reg_mr1rwe_DO_reg[8]/P0001  & ~n17809 ;
  assign n25017 = n19780 & ~n25016 ;
  assign n25018 = ~n25015 & n25017 ;
  assign n25019 = ~n25014 & ~n25018 ;
  assign n25020 = \core_c_dec_EXIT_E_reg/P0001  & n4118 ;
  assign n25021 = \core_c_psq_PCS_reg[3]/NET0131  & n21427 ;
  assign n25022 = n21421 & n25021 ;
  assign n25023 = ~n25020 & ~n25022 ;
  assign n25024 = n13150 & n19923 ;
  assign n25025 = n23407 & n25011 ;
  assign n25026 = n23032 & n25025 ;
  assign n25027 = n14752 & n24963 ;
  assign n25028 = n17836 & n19776 ;
  assign n25029 = \core_eu_em_mac_em_reg_mr1rwe_DO_reg[13]/P0001  & ~n17809 ;
  assign n25030 = n19780 & ~n25029 ;
  assign n25031 = ~n25028 & n25030 ;
  assign n25032 = ~n25027 & ~n25031 ;
  assign n25033 = \sice_IAR_reg[1]/NET0131  & ~\sice_IAR_reg[2]/NET0131  ;
  assign n25034 = n25011 & n25033 ;
  assign n25035 = n23032 & n25034 ;
  assign n25036 = n14752 & ~n25004 ;
  assign n25037 = n19776 & n23920 ;
  assign n25038 = \core_eu_em_mac_em_reg_mr1rwe_DO_reg[12]/P0001  & ~n17809 ;
  assign n25039 = n19780 & ~n25038 ;
  assign n25040 = ~n25037 & n25039 ;
  assign n25041 = ~n25036 & ~n25040 ;
  assign n25042 = ~\clkc_RSTtext_reg/P0001  & n12234 ;
  assign n25043 = n23020 & n25042 ;
  assign n25044 = n20573 & n20574 ;
  assign n25045 = ~\core_c_psq_SSTAT_reg[7]/NET0131  & ~n25044 ;
  assign n25047 = ~n4117 & n19701 ;
  assign n25046 = ~\core_c_dec_accPM_E_reg/P0001  & n4117 ;
  assign n25048 = n4116 & ~n25046 ;
  assign n25049 = ~n25047 & n25048 ;
  assign n25050 = \core_c_dec_RET_Ed_reg/P0001  & n4117 ;
  assign n25051 = ~n21429 & ~n25050 ;
  assign n25052 = n4116 & ~n25051 ;
  assign n25053 = ~\sice_IAR_reg[0]/NET0131  & \sice_IAR_reg[3]/NET0131  ;
  assign n25054 = n25010 & n25053 ;
  assign n25055 = n23032 & n25054 ;
  assign n25056 = \sport0_cfg_SP_ENg_reg/NET0131  & ~\sport0_txctl_TCS_reg[1]/NET0131  ;
  assign n25057 = ~n19960 & n25056 ;
  assign n25058 = \sport0_regs_AUTOreg_DO_reg[1]/NET0131  & n25057 ;
  assign n25059 = ~\sport0_txctl_TSreqi_reg/NET0131  & ~n25058 ;
  assign n25060 = ~\bdma_BWcnt_reg[0]/NET0131  & ~n20036 ;
  assign n25061 = ~n23710 & ~n25060 ;
  assign n25062 = ~n13750 & n25061 ;
  assign n25063 = \core_c_psq_MSTAT_reg_DO_reg[4]/NET0131  & ~n24719 ;
  assign n25064 = ~n24713 & ~n24714 ;
  assign n25065 = n22709 & ~n25064 ;
  assign n25066 = ~n22709 & n25064 ;
  assign n25067 = ~n25065 & ~n25066 ;
  assign n25068 = ~\core_c_psq_MSTAT_reg_DO_reg[4]/NET0131  & n25067 ;
  assign n25069 = ~n25063 & ~n25068 ;
  assign n25070 = \sport1_cfg_SP_ENg_reg/NET0131  & ~\sport1_txctl_TCS_reg[1]/NET0131  ;
  assign n25071 = ~n22677 & n25070 ;
  assign n25072 = \sport1_regs_AUTOreg_DO_reg[1]/NET0131  & n25071 ;
  assign n25073 = ~\sport1_txctl_TSreqi_reg/NET0131  & ~n25072 ;
  assign n25074 = n23028 & n25011 ;
  assign n25075 = n23032 & n25074 ;
  assign n25076 = ~\bdma_BWcnt_reg[2]/NET0131  & ~\bdma_BWcnt_reg[3]/NET0131  ;
  assign n25077 = ~\bdma_BWcnt_reg[4]/NET0131  & n25076 ;
  assign n25078 = n12525 & n20037 ;
  assign n25079 = n25077 & n25078 ;
  assign n25080 = ~\core_c_dec_IR_reg[15]/NET0131  & n19696 ;
  assign n25081 = n21249 & n25080 ;
  assign n25082 = n11741 & n25081 ;
  assign n25083 = ~\sice_IAR_reg[1]/NET0131  & n23408 ;
  assign n25084 = \sice_IAR_reg[2]/NET0131  & n25083 ;
  assign n25085 = n23032 & n25084 ;
  assign n25086 = \core_c_psq_MSTAT_reg_DO_reg[4]/NET0131  & ~n19407 ;
  assign n25087 = ~\core_c_psq_MSTAT_reg_DO_reg[4]/NET0131  & n19368 ;
  assign n25088 = ~n25086 & ~n25087 ;
  assign n25089 = \core_c_psq_T_IRQ1p_reg/P0001  & \core_c_psq_irq1_de_OUT_reg/P0001  ;
  assign n25090 = ~\core_c_psq_T_IRQ1p_reg/P0001  & ~\core_c_psq_irq1_de_OUT_reg/P0001  ;
  assign n25091 = \core_c_psq_irq1_de_IN_syn_reg/P0001  & ~n25090 ;
  assign n25092 = ~n25089 & ~n25091 ;
  assign n25093 = \core_c_psq_T_IRQ0p_reg/P0001  & \core_c_psq_irq0_de_OUT_reg/P0001  ;
  assign n25094 = ~\core_c_psq_T_IRQ0p_reg/P0001  & ~\core_c_psq_irq0_de_OUT_reg/P0001  ;
  assign n25095 = \core_c_psq_irq0_de_IN_syn_reg/P0001  & ~n25094 ;
  assign n25096 = ~n25093 & ~n25095 ;
  assign n25097 = \core_c_dec_MTIFC_Eg_reg/P0001  & ~n5950 ;
  assign n25098 = n8460 & n25097 ;
  assign n25099 = \core_c_psq_IFC_reg[10]/NET0131  & ~\core_c_psq_IFC_reg[11]/NET0131  ;
  assign n25100 = ~n25097 & n25099 ;
  assign n25101 = ~n25098 & ~n25100 ;
  assign n25102 = \core_c_psq_T_IRQ2p_reg/P0001  & \core_c_psq_irq2_de_OUT_reg/P0001  ;
  assign n25103 = ~\core_c_psq_T_IRQ2p_reg/P0001  & ~\core_c_psq_irq2_de_OUT_reg/P0001  ;
  assign n25104 = \core_c_psq_irq2_de_IN_syn_reg/P0001  & ~n25103 ;
  assign n25105 = ~n25102 & ~n25104 ;
  assign n25106 = n10289 & n25097 ;
  assign n25107 = \core_c_psq_IFC_reg[8]/NET0131  & ~\core_c_psq_IFC_reg[9]/NET0131  ;
  assign n25108 = ~n25097 & n25107 ;
  assign n25109 = ~n25106 & ~n25108 ;
  assign n25110 = \core_c_psq_T_IRQL1p_reg/P0001  & \core_c_psq_irql1_de_OUT_reg/P0001  ;
  assign n25111 = ~\core_c_psq_T_IRQL1p_reg/P0001  & ~\core_c_psq_irql1_de_OUT_reg/P0001  ;
  assign n25112 = \core_c_psq_irql1_de_IN_syn_reg/P0001  & ~n25111 ;
  assign n25113 = ~n25110 & ~n25112 ;
  assign n25114 = \core_c_dec_MTMX1_E_reg/P0001  & n17798 ;
  assign n25115 = ~n17836 & n25114 ;
  assign n25116 = ~\core_eu_em_mac_em_reg_mx1rwe_DO_reg[13]/P0001  & ~n25114 ;
  assign n25117 = ~n25115 & ~n25116 ;
  assign n25118 = \core_c_dec_MTMX0_E_reg/P0001  & n17798 ;
  assign n25119 = ~n19848 & n25118 ;
  assign n25120 = ~\core_eu_em_mac_em_reg_mx0rwe_DO_reg[10]/P0001  & ~n25118 ;
  assign n25121 = ~n25119 & ~n25120 ;
  assign n25122 = ~n23920 & n25118 ;
  assign n25123 = ~\core_eu_em_mac_em_reg_mx0rwe_DO_reg[12]/P0001  & ~n25118 ;
  assign n25124 = ~n25122 & ~n25123 ;
  assign n25125 = \core_c_dec_MTMX0_E_reg/P0001  & n14665 ;
  assign n25126 = ~n23920 & n25125 ;
  assign n25127 = ~\core_eu_em_mac_em_reg_mx0swe_DO_reg[12]/P0001  & ~n25125 ;
  assign n25128 = ~n25126 & ~n25127 ;
  assign n25129 = ~n23920 & n25114 ;
  assign n25130 = ~\core_eu_em_mac_em_reg_mx1rwe_DO_reg[12]/P0001  & ~n25114 ;
  assign n25131 = ~n25129 & ~n25130 ;
  assign n25132 = \core_c_dec_MTMX1_E_reg/P0001  & n14665 ;
  assign n25133 = ~n19504 & n25132 ;
  assign n25134 = ~\core_eu_em_mac_em_reg_mx1swe_DO_reg[9]/P0001  & ~n25132 ;
  assign n25135 = ~n25133 & ~n25134 ;
  assign n25136 = ~n17836 & n25132 ;
  assign n25137 = ~\core_eu_em_mac_em_reg_mx1swe_DO_reg[13]/P0001  & ~n25132 ;
  assign n25138 = ~n25136 & ~n25137 ;
  assign n25139 = ~n23920 & n25132 ;
  assign n25140 = ~\core_eu_em_mac_em_reg_mx1swe_DO_reg[12]/P0001  & ~n25132 ;
  assign n25141 = ~n25139 & ~n25140 ;
  assign n25142 = ~n19848 & n25132 ;
  assign n25143 = ~\core_eu_em_mac_em_reg_mx1swe_DO_reg[10]/P0001  & ~n25132 ;
  assign n25144 = ~n25142 & ~n25143 ;
  assign n25145 = ~n23860 & n25114 ;
  assign n25146 = ~\core_eu_em_mac_em_reg_mx1rwe_DO_reg[8]/P0001  & ~n25114 ;
  assign n25147 = ~n25145 & ~n25146 ;
  assign n25148 = ~n23860 & n25125 ;
  assign n25149 = ~\core_eu_em_mac_em_reg_mx0swe_DO_reg[8]/P0001  & ~n25125 ;
  assign n25150 = ~n25148 & ~n25149 ;
  assign n25151 = ~n17836 & n25125 ;
  assign n25152 = ~\core_eu_em_mac_em_reg_mx0swe_DO_reg[13]/P0001  & ~n25125 ;
  assign n25153 = ~n25151 & ~n25152 ;
  assign n25154 = ~n23757 & n25125 ;
  assign n25155 = ~\core_eu_em_mac_em_reg_mx0swe_DO_reg[11]/P0001  & ~n25125 ;
  assign n25156 = ~n25154 & ~n25155 ;
  assign n25157 = ~n23860 & n25118 ;
  assign n25158 = ~\core_eu_em_mac_em_reg_mx0rwe_DO_reg[8]/P0001  & ~n25118 ;
  assign n25159 = ~n25157 & ~n25158 ;
  assign n25160 = ~n17836 & n25118 ;
  assign n25161 = ~\core_eu_em_mac_em_reg_mx0rwe_DO_reg[13]/P0001  & ~n25118 ;
  assign n25162 = ~n25160 & ~n25161 ;
  assign n25163 = ~n19504 & n25118 ;
  assign n25164 = ~\core_eu_em_mac_em_reg_mx0rwe_DO_reg[9]/P0001  & ~n25118 ;
  assign n25165 = ~n25163 & ~n25164 ;
  assign n25166 = ~n23757 & n25118 ;
  assign n25167 = ~\core_eu_em_mac_em_reg_mx0rwe_DO_reg[11]/P0001  & ~n25118 ;
  assign n25168 = ~n25166 & ~n25167 ;
  assign n25169 = ~n23757 & n25132 ;
  assign n25170 = ~\core_eu_em_mac_em_reg_mx1swe_DO_reg[11]/P0001  & ~n25132 ;
  assign n25171 = ~n25169 & ~n25170 ;
  assign n25172 = ~n19848 & n25125 ;
  assign n25173 = ~\core_eu_em_mac_em_reg_mx0swe_DO_reg[10]/P0001  & ~n25125 ;
  assign n25174 = ~n25172 & ~n25173 ;
  assign n25175 = ~n19504 & n25125 ;
  assign n25176 = ~\core_eu_em_mac_em_reg_mx0swe_DO_reg[9]/P0001  & ~n25125 ;
  assign n25177 = ~n25175 & ~n25176 ;
  assign n25178 = ~n23860 & n25132 ;
  assign n25179 = ~\core_eu_em_mac_em_reg_mx1swe_DO_reg[8]/P0001  & ~n25132 ;
  assign n25180 = ~n25178 & ~n25179 ;
  assign n25181 = ~n23757 & n25114 ;
  assign n25182 = ~\core_eu_em_mac_em_reg_mx1rwe_DO_reg[11]/P0001  & ~n25114 ;
  assign n25183 = ~n25181 & ~n25182 ;
  assign n25184 = ~n19848 & n25114 ;
  assign n25185 = ~\core_eu_em_mac_em_reg_mx1rwe_DO_reg[10]/P0001  & ~n25114 ;
  assign n25186 = ~n25184 & ~n25185 ;
  assign n25187 = ~n19504 & n25114 ;
  assign n25188 = ~\core_eu_em_mac_em_reg_mx1rwe_DO_reg[9]/P0001  & ~n25114 ;
  assign n25189 = ~n25187 & ~n25188 ;
  assign n25190 = n4099 & ~n5950 ;
  assign n25191 = \memc_Pwrite_E_reg/NET0131  & ~n12918 ;
  assign n25192 = ~\memc_Pwrite_E_reg/NET0131  & ~n10905 ;
  assign n25193 = ~n25191 & ~n25192 ;
  assign n25194 = n25190 & ~n25193 ;
  assign n25195 = \regout_STD_C_reg[5]/P0001  & ~n25190 ;
  assign n25196 = ~n25194 & ~n25195 ;
  assign n25197 = ~n17814 & n25132 ;
  assign n25198 = ~\core_eu_em_mac_em_reg_mx1swe_DO_reg[2]/P0001  & ~n25132 ;
  assign n25199 = ~n25197 & ~n25198 ;
  assign n25200 = ~\core_c_psq_PCS_reg[10]/NET0131  & n4094 ;
  assign n25201 = ~T_BRn_pad & ~n25200 ;
  assign n25202 = \core_c_psq_MREQ_reg/NET0131  & n5679 ;
  assign n25203 = n4112 & n25202 ;
  assign n25204 = n25200 & n25203 ;
  assign n25205 = ~n25201 & ~n25204 ;
  assign n25206 = \core_c_dec_IRE_reg[6]/NET0131  & \core_c_dec_Stkctl_Eg_reg/P0001  ;
  assign n25207 = ~n5950 & n25206 ;
  assign n25208 = \core_c_psq_INT_en_reg/NET0131  & ~n25207 ;
  assign n25209 = \core_c_dec_IRE_reg[5]/NET0131  & n25207 ;
  assign n25210 = ~n25208 & ~n25209 ;
  assign n25211 = \memc_Pwrite_E_reg/NET0131  & ~n12751 ;
  assign n25212 = ~\memc_Pwrite_E_reg/NET0131  & ~n12095 ;
  assign n25213 = ~n25211 & ~n25212 ;
  assign n25214 = n25190 & ~n25213 ;
  assign n25215 = \regout_STD_C_reg[15]/P0001  & ~n25190 ;
  assign n25216 = ~n25214 & ~n25215 ;
  assign n25217 = n10638 & n25097 ;
  assign n25218 = ~\core_c_psq_IFC_reg[8]/NET0131  & \core_c_psq_IFC_reg[9]/NET0131  ;
  assign n25219 = ~n25097 & n25218 ;
  assign n25220 = ~n25217 & ~n25219 ;
  assign n25221 = n11265 & n25097 ;
  assign n25222 = \core_c_psq_IFC_reg[6]/NET0131  & ~\core_c_psq_IFC_reg[7]/NET0131  ;
  assign n25223 = ~n25097 & n25222 ;
  assign n25224 = ~n25221 & ~n25223 ;
  assign n25225 = \core_c_dec_MTDMOVL_E_reg/P0001  & n5951 ;
  assign n25226 = ~n8113 & n25225 ;
  assign n25227 = ~\core_c_psq_DMOVL_reg_DO_reg[3]/NET0131  & ~n25225 ;
  assign n25228 = ~n25226 & ~n25227 ;
  assign n25229 = ~n8715 & n25225 ;
  assign n25230 = ~\core_c_psq_DMOVL_reg_DO_reg[2]/NET0131  & ~n25225 ;
  assign n25231 = ~n25229 & ~n25230 ;
  assign n25232 = ~n9435 & n25225 ;
  assign n25233 = ~\core_c_psq_DMOVL_reg_DO_reg[1]/NET0131  & ~n25225 ;
  assign n25234 = ~n25232 & ~n25233 ;
  assign n25235 = ~n7607 & n25225 ;
  assign n25236 = ~\core_c_psq_DMOVL_reg_DO_reg[0]/NET0131  & ~n25225 ;
  assign n25237 = ~n25235 & ~n25236 ;
  assign n25238 = \memc_Pwrite_E_reg/NET0131  & ~n12638 ;
  assign n25239 = ~\memc_Pwrite_E_reg/NET0131  & ~n7334 ;
  assign n25240 = ~n25238 & ~n25239 ;
  assign n25241 = n25190 & ~n25240 ;
  assign n25242 = \regout_STD_C_reg[13]/P0001  & ~n25190 ;
  assign n25243 = ~n25241 & ~n25242 ;
  assign n25244 = \core_c_dec_IR_reg[19]/NET0131  & n14727 ;
  assign n25245 = ~n4117 & n25244 ;
  assign n25246 = \core_c_dec_imm14_E_reg/P0001  & n4117 ;
  assign n25247 = ~n25245 & ~n25246 ;
  assign n25248 = \core_c_dec_DU_Eg_reg/P0001  & n4118 ;
  assign n25249 = \core_c_dec_IR_reg[19]/NET0131  & n6118 ;
  assign n25250 = n23231 & n25249 ;
  assign n25251 = ~n25248 & ~n25250 ;
  assign n25252 = ~n20259 & n25114 ;
  assign n25253 = ~\core_eu_em_mac_em_reg_mx1rwe_DO_reg[5]/P0001  & ~n25114 ;
  assign n25254 = ~n25252 & ~n25253 ;
  assign n25255 = ~n20259 & n25118 ;
  assign n25256 = ~\core_eu_em_mac_em_reg_mx0rwe_DO_reg[5]/P0001  & ~n25118 ;
  assign n25257 = ~n25255 & ~n25256 ;
  assign n25258 = ~n20150 & n25125 ;
  assign n25259 = ~\core_eu_em_mac_em_reg_mx0swe_DO_reg[14]/P0001  & ~n25125 ;
  assign n25260 = ~n25258 & ~n25259 ;
  assign n25261 = ~n19972 & n25132 ;
  assign n25262 = ~\core_eu_em_mac_em_reg_mx1swe_DO_reg[7]/P0001  & ~n25132 ;
  assign n25263 = ~n25261 & ~n25262 ;
  assign n25264 = ~n20259 & n25132 ;
  assign n25265 = ~\core_eu_em_mac_em_reg_mx1swe_DO_reg[5]/P0001  & ~n25132 ;
  assign n25266 = ~n25264 & ~n25265 ;
  assign n25267 = ~n21663 & n25132 ;
  assign n25268 = ~\core_eu_em_mac_em_reg_mx1swe_DO_reg[3]/P0001  & ~n25132 ;
  assign n25269 = ~n25267 & ~n25268 ;
  assign n25270 = ~n18974 & n25132 ;
  assign n25271 = ~\core_eu_em_mac_em_reg_mx1swe_DO_reg[1]/P0001  & ~n25132 ;
  assign n25272 = ~n25270 & ~n25271 ;
  assign n25273 = ~n18276 & n25114 ;
  assign n25274 = ~\core_eu_em_mac_em_reg_mx1rwe_DO_reg[6]/P0001  & ~n25114 ;
  assign n25275 = ~n25273 & ~n25274 ;
  assign n25276 = ~n21663 & n25114 ;
  assign n25277 = ~\core_eu_em_mac_em_reg_mx1rwe_DO_reg[3]/P0001  & ~n25114 ;
  assign n25278 = ~n25276 & ~n25277 ;
  assign n25279 = ~n17814 & n25114 ;
  assign n25280 = ~\core_eu_em_mac_em_reg_mx1rwe_DO_reg[2]/P0001  & ~n25114 ;
  assign n25281 = ~n25279 & ~n25280 ;
  assign n25282 = ~n17820 & n25114 ;
  assign n25283 = ~\core_eu_em_mac_em_reg_mx1rwe_DO_reg[15]/P0001  & ~n25114 ;
  assign n25284 = ~n25282 & ~n25283 ;
  assign n25285 = ~n19559 & n25114 ;
  assign n25286 = ~\core_eu_em_mac_em_reg_mx1rwe_DO_reg[0]/P0001  & ~n25114 ;
  assign n25287 = ~n25285 & ~n25286 ;
  assign n25288 = ~n19972 & n25125 ;
  assign n25289 = ~\core_eu_em_mac_em_reg_mx0swe_DO_reg[7]/P0001  & ~n25125 ;
  assign n25290 = ~n25288 & ~n25289 ;
  assign n25291 = ~n18276 & n25125 ;
  assign n25292 = ~\core_eu_em_mac_em_reg_mx0swe_DO_reg[6]/P0001  & ~n25125 ;
  assign n25293 = ~n25291 & ~n25292 ;
  assign n25294 = ~n21663 & n25125 ;
  assign n25295 = ~\core_eu_em_mac_em_reg_mx0swe_DO_reg[3]/P0001  & ~n25125 ;
  assign n25296 = ~n25294 & ~n25295 ;
  assign n25297 = ~n17814 & n25125 ;
  assign n25298 = ~\core_eu_em_mac_em_reg_mx0swe_DO_reg[2]/P0001  & ~n25125 ;
  assign n25299 = ~n25297 & ~n25298 ;
  assign n25300 = ~n18276 & n25118 ;
  assign n25301 = ~\core_eu_em_mac_em_reg_mx0rwe_DO_reg[6]/P0001  & ~n25118 ;
  assign n25302 = ~n25300 & ~n25301 ;
  assign n25303 = ~n21663 & n25118 ;
  assign n25304 = ~\core_eu_em_mac_em_reg_mx0rwe_DO_reg[3]/P0001  & ~n25118 ;
  assign n25305 = ~n25303 & ~n25304 ;
  assign n25306 = ~n17814 & n25118 ;
  assign n25307 = ~\core_eu_em_mac_em_reg_mx0rwe_DO_reg[2]/P0001  & ~n25118 ;
  assign n25308 = ~n25306 & ~n25307 ;
  assign n25309 = ~n20150 & n25118 ;
  assign n25310 = ~\core_eu_em_mac_em_reg_mx0rwe_DO_reg[14]/P0001  & ~n25118 ;
  assign n25311 = ~n25309 & ~n25310 ;
  assign n25312 = ~n19559 & n25118 ;
  assign n25313 = ~\core_eu_em_mac_em_reg_mx0rwe_DO_reg[0]/P0001  & ~n25118 ;
  assign n25314 = ~n25312 & ~n25313 ;
  assign n25315 = \core_c_dec_RTI_Ed_reg/P0001  & n4118 ;
  assign n25316 = \core_c_dec_IR_reg[4]/NET0131  & n4116 ;
  assign n25317 = n21429 & n25316 ;
  assign n25318 = ~n25315 & ~n25317 ;
  assign n25319 = \memc_Pwrite_E_reg/NET0131  & ~n13055 ;
  assign n25320 = ~\memc_Pwrite_E_reg/NET0131  & ~n10283 ;
  assign n25321 = ~n25319 & ~n25320 ;
  assign n25322 = n25190 & ~n25321 ;
  assign n25323 = \regout_STD_C_reg[9]/P0001  & ~n25190 ;
  assign n25324 = ~n25322 & ~n25323 ;
  assign n25325 = \memc_Pwrite_E_reg/NET0131  & ~n12850 ;
  assign n25326 = ~\memc_Pwrite_E_reg/NET0131  & ~n8107 ;
  assign n25327 = ~n25325 & ~n25326 ;
  assign n25328 = n25190 & ~n25327 ;
  assign n25329 = \regout_STD_C_reg[3]/P0001  & ~n25190 ;
  assign n25330 = ~n25328 & ~n25329 ;
  assign n25331 = \memc_Pwrite_E_reg/NET0131  & ~n12570 ;
  assign n25332 = ~\memc_Pwrite_E_reg/NET0131  & ~n8454 ;
  assign n25333 = ~n25331 & ~n25332 ;
  assign n25334 = n25190 & ~n25333 ;
  assign n25335 = \regout_STD_C_reg[11]/P0001  & ~n25190 ;
  assign n25336 = ~n25334 & ~n25335 ;
  assign n25337 = ~n18974 & n25125 ;
  assign n25338 = ~\core_eu_em_mac_em_reg_mx0swe_DO_reg[1]/P0001  & ~n25125 ;
  assign n25339 = ~n25337 & ~n25338 ;
  assign n25340 = n7859 & n25097 ;
  assign n25341 = ~\core_c_psq_IFC_reg[10]/NET0131  & \core_c_psq_IFC_reg[11]/NET0131  ;
  assign n25342 = ~n25097 & n25341 ;
  assign n25343 = ~n25340 & ~n25342 ;
  assign n25344 = ~n20150 & n25114 ;
  assign n25345 = ~\core_eu_em_mac_em_reg_mx1rwe_DO_reg[14]/P0001  & ~n25114 ;
  assign n25346 = ~n25344 & ~n25345 ;
  assign n25347 = ~n20080 & n25132 ;
  assign n25348 = ~\core_eu_em_mac_em_reg_mx1swe_DO_reg[4]/P0001  & ~n25132 ;
  assign n25349 = ~n25347 & ~n25348 ;
  assign n25350 = ~n19559 & n25125 ;
  assign n25351 = ~\core_eu_em_mac_em_reg_mx0swe_DO_reg[0]/P0001  & ~n25125 ;
  assign n25352 = ~n25350 & ~n25351 ;
  assign n25353 = n8113 & n25097 ;
  assign n25354 = \core_c_psq_IFC_reg[2]/NET0131  & ~\core_c_psq_IFC_reg[3]/NET0131  ;
  assign n25355 = ~n25097 & n25354 ;
  assign n25356 = ~n25353 & ~n25355 ;
  assign n25357 = n10911 & n25097 ;
  assign n25358 = \core_c_psq_IFC_reg[4]/NET0131  & ~\core_c_psq_IFC_reg[5]/NET0131  ;
  assign n25359 = ~n25097 & n25358 ;
  assign n25360 = ~n25357 & ~n25359 ;
  assign n25361 = ~n17820 & n25125 ;
  assign n25362 = ~\core_eu_em_mac_em_reg_mx0swe_DO_reg[15]/P0001  & ~n25125 ;
  assign n25363 = ~n25361 & ~n25362 ;
  assign n25364 = \memc_Pwrite_E_reg/NET0131  & ~n12695 ;
  assign n25365 = ~\memc_Pwrite_E_reg/NET0131  & ~n11953 ;
  assign n25366 = ~n25364 & ~n25365 ;
  assign n25367 = n25190 & ~n25366 ;
  assign n25368 = \regout_STD_C_reg[14]/P0001  & ~n25190 ;
  assign n25369 = ~n25367 & ~n25368 ;
  assign n25370 = ~n17820 & n25118 ;
  assign n25371 = ~\core_eu_em_mac_em_reg_mx0rwe_DO_reg[15]/P0001  & ~n25118 ;
  assign n25372 = ~n25370 & ~n25371 ;
  assign n25373 = \memc_Pwrite_E_reg/NET0131  & ~n12782 ;
  assign n25374 = ~\memc_Pwrite_E_reg/NET0131  & ~n9429 ;
  assign n25375 = ~n25373 & ~n25374 ;
  assign n25376 = n25190 & ~n25375 ;
  assign n25377 = \regout_STD_C_reg[1]/P0001  & ~n25190 ;
  assign n25378 = ~n25376 & ~n25377 ;
  assign n25379 = ~n19972 & n25118 ;
  assign n25380 = ~\core_eu_em_mac_em_reg_mx0rwe_DO_reg[7]/P0001  & ~n25118 ;
  assign n25381 = ~n25379 & ~n25380 ;
  assign n25382 = ~n20080 & n25125 ;
  assign n25383 = ~\core_eu_em_mac_em_reg_mx0swe_DO_reg[4]/P0001  & ~n25125 ;
  assign n25384 = ~n25382 & ~n25383 ;
  assign n25385 = ~n18974 & n25114 ;
  assign n25386 = ~\core_eu_em_mac_em_reg_mx1rwe_DO_reg[1]/P0001  & ~n25114 ;
  assign n25387 = ~n25385 & ~n25386 ;
  assign n25388 = \memc_Pwrite_E_reg/NET0131  & ~n13021 ;
  assign n25389 = ~\memc_Pwrite_E_reg/NET0131  & ~n10632 ;
  assign n25390 = ~n25388 & ~n25389 ;
  assign n25391 = n25190 & ~n25390 ;
  assign n25392 = \regout_STD_C_reg[8]/P0001  & ~n25190 ;
  assign n25393 = ~n25391 & ~n25392 ;
  assign n25394 = \memc_Pwrite_E_reg/NET0131  & ~n12884 ;
  assign n25395 = ~\memc_Pwrite_E_reg/NET0131  & ~n10063 ;
  assign n25396 = ~n25394 & ~n25395 ;
  assign n25397 = n25190 & ~n25396 ;
  assign n25398 = \regout_STD_C_reg[4]/P0001  & ~n25190 ;
  assign n25399 = ~n25397 & ~n25398 ;
  assign n25400 = ~n18276 & n25132 ;
  assign n25401 = ~\core_eu_em_mac_em_reg_mx1swe_DO_reg[6]/P0001  & ~n25132 ;
  assign n25402 = ~n25400 & ~n25401 ;
  assign n25403 = ~n20150 & n25132 ;
  assign n25404 = ~\core_eu_em_mac_em_reg_mx1swe_DO_reg[14]/P0001  & ~n25132 ;
  assign n25405 = ~n25403 & ~n25404 ;
  assign n25406 = \memc_Pwrite_E_reg/NET0131  & ~n12473 ;
  assign n25407 = ~\memc_Pwrite_E_reg/NET0131  & ~n7601 ;
  assign n25408 = ~n25406 & ~n25407 ;
  assign n25409 = n25190 & ~n25408 ;
  assign n25410 = \regout_STD_C_reg[0]/P0001  & ~n25190 ;
  assign n25411 = ~n25409 & ~n25410 ;
  assign n25412 = \memc_Pwrite_E_reg/NET0131  & ~n12986 ;
  assign n25413 = ~\memc_Pwrite_E_reg/NET0131  & ~n11259 ;
  assign n25414 = ~n25412 & ~n25413 ;
  assign n25415 = n25190 & ~n25414 ;
  assign n25416 = \regout_STD_C_reg[7]/P0001  & ~n25190 ;
  assign n25417 = ~n25415 & ~n25416 ;
  assign n25418 = n9435 & n25097 ;
  assign n25419 = \core_c_psq_IFC_reg[0]/NET0131  & ~\core_c_psq_IFC_reg[1]/NET0131  ;
  assign n25420 = ~n25097 & n25419 ;
  assign n25421 = ~n25418 & ~n25420 ;
  assign n25422 = \memc_Pwrite_E_reg/NET0131  & ~n12604 ;
  assign n25423 = ~\memc_Pwrite_E_reg/NET0131  & ~n9172 ;
  assign n25424 = ~n25422 & ~n25423 ;
  assign n25425 = n25190 & ~n25424 ;
  assign n25426 = \regout_STD_C_reg[12]/P0001  & ~n25190 ;
  assign n25427 = ~n25425 & ~n25426 ;
  assign n25428 = \memc_Pwrite_E_reg/NET0131  & ~n12816 ;
  assign n25429 = ~\memc_Pwrite_E_reg/NET0131  & ~n8709 ;
  assign n25430 = ~n25428 & ~n25429 ;
  assign n25431 = n25190 & ~n25430 ;
  assign n25432 = \regout_STD_C_reg[2]/P0001  & ~n25190 ;
  assign n25433 = ~n25431 & ~n25432 ;
  assign n25434 = ~n19559 & n25132 ;
  assign n25435 = ~\core_eu_em_mac_em_reg_mx1swe_DO_reg[0]/P0001  & ~n25132 ;
  assign n25436 = ~n25434 & ~n25435 ;
  assign n25437 = \memc_Pwrite_E_reg/NET0131  & ~n12536 ;
  assign n25438 = ~\memc_Pwrite_E_reg/NET0131  & ~n7853 ;
  assign n25439 = ~n25437 & ~n25438 ;
  assign n25440 = n25190 & ~n25439 ;
  assign n25441 = \regout_STD_C_reg[10]/P0001  & ~n25190 ;
  assign n25442 = ~n25440 & ~n25441 ;
  assign n25443 = ~n20080 & n25118 ;
  assign n25444 = ~\core_eu_em_mac_em_reg_mx0rwe_DO_reg[4]/P0001  & ~n25118 ;
  assign n25445 = ~n25443 & ~n25444 ;
  assign n25446 = \memc_Pwrite_E_reg/NET0131  & ~n12968 ;
  assign n25447 = ~\memc_Pwrite_E_reg/NET0131  & ~n11519 ;
  assign n25448 = ~n25446 & ~n25447 ;
  assign n25449 = n25190 & ~n25448 ;
  assign n25450 = \regout_STD_C_reg[6]/P0001  & ~n25190 ;
  assign n25451 = ~n25449 & ~n25450 ;
  assign n25452 = ~n20080 & n25114 ;
  assign n25453 = ~\core_eu_em_mac_em_reg_mx1rwe_DO_reg[4]/P0001  & ~n25114 ;
  assign n25454 = ~n25452 & ~n25453 ;
  assign n25455 = ~n19972 & n25114 ;
  assign n25456 = ~\core_eu_em_mac_em_reg_mx1rwe_DO_reg[7]/P0001  & ~n25114 ;
  assign n25457 = ~n25455 & ~n25456 ;
  assign n25458 = ~n20259 & n25125 ;
  assign n25459 = ~\core_eu_em_mac_em_reg_mx0swe_DO_reg[5]/P0001  & ~n25125 ;
  assign n25460 = ~n25458 & ~n25459 ;
  assign n25461 = ~n17820 & n25132 ;
  assign n25462 = ~\core_eu_em_mac_em_reg_mx1swe_DO_reg[15]/P0001  & ~n25132 ;
  assign n25463 = ~n25461 & ~n25462 ;
  assign n25464 = ~n18974 & n25118 ;
  assign n25465 = ~\core_eu_em_mac_em_reg_mx0rwe_DO_reg[1]/P0001  & ~n25118 ;
  assign n25466 = ~n25464 & ~n25465 ;
  assign n25467 = \memc_Pwrite_E_reg/NET0131  & n4117 ;
  assign n25468 = \core_c_dec_IR_reg[15]/NET0131  & n13574 ;
  assign n25469 = \core_c_dec_IR_reg[19]/NET0131  & n13577 ;
  assign n25470 = ~n25468 & ~n25469 ;
  assign n25471 = n11742 & ~n25470 ;
  assign n25472 = ~n25467 & ~n25471 ;
  assign n25473 = n11525 & n25097 ;
  assign n25474 = ~\core_c_psq_IFC_reg[6]/NET0131  & \core_c_psq_IFC_reg[7]/NET0131  ;
  assign n25475 = ~n25097 & n25474 ;
  assign n25476 = ~n25473 & ~n25475 ;
  assign n25477 = n10069 & n25097 ;
  assign n25478 = ~\core_c_psq_IFC_reg[4]/NET0131  & \core_c_psq_IFC_reg[5]/NET0131  ;
  assign n25479 = ~n25097 & n25478 ;
  assign n25480 = ~n25477 & ~n25479 ;
  assign n25481 = n8715 & n25097 ;
  assign n25482 = ~\core_c_psq_IFC_reg[2]/NET0131  & \core_c_psq_IFC_reg[3]/NET0131  ;
  assign n25483 = ~n25097 & n25482 ;
  assign n25484 = ~n25481 & ~n25483 ;
  assign n25485 = n7607 & n25097 ;
  assign n25486 = ~\core_c_psq_IFC_reg[0]/NET0131  & \core_c_psq_IFC_reg[1]/NET0131  ;
  assign n25487 = ~n25097 & n25486 ;
  assign n25488 = ~n25485 & ~n25487 ;
  assign n25489 = \core_c_psq_MSTAT_reg_DO_reg[5]/NET0131  & ~n22408 ;
  assign n25490 = ~\T_TMODE[0]_pad  & ~n25489 ;
  assign n25491 = ~n20357 & ~n25490 ;
  assign n25492 = ~\T_TMODE[0]_pad  & ~n22404 ;
  assign n25493 = ~\core_c_psq_PCS_reg[3]/NET0131  & ~n25492 ;
  assign n25494 = ~\tm_TSR_TMP_reg[4]/NET0131  & n25493 ;
  assign n25495 = ~\tm_TSR_TMP_reg[5]/NET0131  & n25494 ;
  assign n25496 = ~\tm_TSR_TMP_reg[6]/NET0131  & n25495 ;
  assign n25497 = \tm_TSR_TMP_reg[7]/NET0131  & ~n25496 ;
  assign n25498 = ~\tm_TSR_TMP_reg[7]/NET0131  & n25496 ;
  assign n25499 = ~n25497 & ~n25498 ;
  assign n25500 = n25491 & ~n25499 ;
  assign n25501 = \tm_tsr_reg_DO_reg[7]/NET0131  & ~n25491 ;
  assign n25502 = ~n25500 & ~n25501 ;
  assign n25503 = \core_c_dec_MTSI_E_reg/P0001  & n17798 ;
  assign n25504 = ~n19504 & n25503 ;
  assign n25505 = ~\core_eu_es_sht_es_reg_sirwe_DO_reg[9]/P0001  & ~n25503 ;
  assign n25506 = ~n25504 & ~n25505 ;
  assign n25507 = ~n17836 & n25503 ;
  assign n25508 = ~\core_eu_es_sht_es_reg_sirwe_DO_reg[13]/P0001  & ~n25503 ;
  assign n25509 = ~n25507 & ~n25508 ;
  assign n25510 = ~n23860 & n25503 ;
  assign n25511 = ~\core_eu_es_sht_es_reg_sirwe_DO_reg[8]/P0001  & ~n25503 ;
  assign n25512 = ~n25510 & ~n25511 ;
  assign n25513 = ~n18276 & n25503 ;
  assign n25514 = ~\core_eu_es_sht_es_reg_sirwe_DO_reg[6]/P0001  & ~n25503 ;
  assign n25515 = ~n25513 & ~n25514 ;
  assign n25516 = ~n17814 & n25503 ;
  assign n25517 = ~\core_eu_es_sht_es_reg_sirwe_DO_reg[2]/P0001  & ~n25503 ;
  assign n25518 = ~n25516 & ~n25517 ;
  assign n25519 = ~n23757 & n25503 ;
  assign n25520 = ~\core_eu_es_sht_es_reg_sirwe_DO_reg[11]/P0001  & ~n25503 ;
  assign n25521 = ~n25519 & ~n25520 ;
  assign n25522 = ~n19559 & n25503 ;
  assign n25523 = ~\core_eu_es_sht_es_reg_sirwe_DO_reg[0]/P0001  & ~n25503 ;
  assign n25524 = ~n25522 & ~n25523 ;
  assign n25525 = ~n20259 & n25503 ;
  assign n25526 = ~\core_eu_es_sht_es_reg_sirwe_DO_reg[5]/P0001  & ~n25503 ;
  assign n25527 = ~n25525 & ~n25526 ;
  assign n25528 = \core_c_dec_MTAX0_E_reg/P0001  & n17798 ;
  assign n25529 = ~n23860 & n25528 ;
  assign n25530 = ~\core_eu_ea_alu_ea_reg_ax0rwe_DO_reg[8]/P0001  & ~n25528 ;
  assign n25531 = ~n25529 & ~n25530 ;
  assign n25532 = ~n17820 & n25503 ;
  assign n25533 = ~\core_eu_es_sht_es_reg_sirwe_DO_reg[15]/P0001  & ~n25503 ;
  assign n25534 = ~n25532 & ~n25533 ;
  assign n25535 = \core_c_dec_MTAX1_E_reg/P0001  & n17798 ;
  assign n25536 = ~n19504 & n25535 ;
  assign n25537 = ~\core_eu_ea_alu_ea_reg_ax1rwe_DO_reg[9]/P0001  & ~n25535 ;
  assign n25538 = ~n25536 & ~n25537 ;
  assign n25539 = ~n23860 & n25535 ;
  assign n25540 = ~\core_eu_ea_alu_ea_reg_ax1rwe_DO_reg[8]/P0001  & ~n25535 ;
  assign n25541 = ~n25539 & ~n25540 ;
  assign n25542 = ~n19972 & n25535 ;
  assign n25543 = ~\core_eu_ea_alu_ea_reg_ax1rwe_DO_reg[7]/P0001  & ~n25535 ;
  assign n25544 = ~n25542 & ~n25543 ;
  assign n25545 = ~n18276 & n25535 ;
  assign n25546 = ~\core_eu_ea_alu_ea_reg_ax1rwe_DO_reg[6]/P0001  & ~n25535 ;
  assign n25547 = ~n25545 & ~n25546 ;
  assign n25548 = ~n20259 & n25535 ;
  assign n25549 = ~\core_eu_ea_alu_ea_reg_ax1rwe_DO_reg[5]/P0001  & ~n25535 ;
  assign n25550 = ~n25548 & ~n25549 ;
  assign n25551 = ~n20080 & n25535 ;
  assign n25552 = ~\core_eu_ea_alu_ea_reg_ax1rwe_DO_reg[4]/P0001  & ~n25535 ;
  assign n25553 = ~n25551 & ~n25552 ;
  assign n25554 = ~n21663 & n25535 ;
  assign n25555 = ~\core_eu_ea_alu_ea_reg_ax1rwe_DO_reg[3]/P0001  & ~n25535 ;
  assign n25556 = ~n25554 & ~n25555 ;
  assign n25557 = ~n17814 & n25535 ;
  assign n25558 = ~\core_eu_ea_alu_ea_reg_ax1rwe_DO_reg[2]/P0001  & ~n25535 ;
  assign n25559 = ~n25557 & ~n25558 ;
  assign n25560 = ~n18974 & n25535 ;
  assign n25561 = ~\core_eu_ea_alu_ea_reg_ax1rwe_DO_reg[1]/P0001  & ~n25535 ;
  assign n25562 = ~n25560 & ~n25561 ;
  assign n25563 = ~n17820 & n25535 ;
  assign n25564 = ~\core_eu_ea_alu_ea_reg_ax1rwe_DO_reg[15]/P0001  & ~n25535 ;
  assign n25565 = ~n25563 & ~n25564 ;
  assign n25566 = ~n20150 & n25535 ;
  assign n25567 = ~\core_eu_ea_alu_ea_reg_ax1rwe_DO_reg[14]/P0001  & ~n25535 ;
  assign n25568 = ~n25566 & ~n25567 ;
  assign n25569 = ~n17836 & n25535 ;
  assign n25570 = ~\core_eu_ea_alu_ea_reg_ax1rwe_DO_reg[13]/P0001  & ~n25535 ;
  assign n25571 = ~n25569 & ~n25570 ;
  assign n25572 = ~n23920 & n25535 ;
  assign n25573 = ~\core_eu_ea_alu_ea_reg_ax1rwe_DO_reg[12]/P0001  & ~n25535 ;
  assign n25574 = ~n25572 & ~n25573 ;
  assign n25575 = ~n23757 & n25535 ;
  assign n25576 = ~\core_eu_ea_alu_ea_reg_ax1rwe_DO_reg[11]/P0001  & ~n25535 ;
  assign n25577 = ~n25575 & ~n25576 ;
  assign n25578 = ~n19848 & n25535 ;
  assign n25579 = ~\core_eu_ea_alu_ea_reg_ax1rwe_DO_reg[10]/P0001  & ~n25535 ;
  assign n25580 = ~n25578 & ~n25579 ;
  assign n25581 = ~n19559 & n25535 ;
  assign n25582 = ~\core_eu_ea_alu_ea_reg_ax1rwe_DO_reg[0]/P0001  & ~n25535 ;
  assign n25583 = ~n25581 & ~n25582 ;
  assign n25584 = ~n19504 & n25528 ;
  assign n25585 = ~\core_eu_ea_alu_ea_reg_ax0rwe_DO_reg[9]/P0001  & ~n25528 ;
  assign n25586 = ~n25584 & ~n25585 ;
  assign n25587 = ~n19972 & n25528 ;
  assign n25588 = ~\core_eu_ea_alu_ea_reg_ax0rwe_DO_reg[7]/P0001  & ~n25528 ;
  assign n25589 = ~n25587 & ~n25588 ;
  assign n25590 = ~n18276 & n25528 ;
  assign n25591 = ~\core_eu_ea_alu_ea_reg_ax0rwe_DO_reg[6]/P0001  & ~n25528 ;
  assign n25592 = ~n25590 & ~n25591 ;
  assign n25593 = ~n20259 & n25528 ;
  assign n25594 = ~\core_eu_ea_alu_ea_reg_ax0rwe_DO_reg[5]/P0001  & ~n25528 ;
  assign n25595 = ~n25593 & ~n25594 ;
  assign n25596 = ~n20080 & n25528 ;
  assign n25597 = ~\core_eu_ea_alu_ea_reg_ax0rwe_DO_reg[4]/P0001  & ~n25528 ;
  assign n25598 = ~n25596 & ~n25597 ;
  assign n25599 = ~n21663 & n25528 ;
  assign n25600 = ~\core_eu_ea_alu_ea_reg_ax0rwe_DO_reg[3]/P0001  & ~n25528 ;
  assign n25601 = ~n25599 & ~n25600 ;
  assign n25602 = ~n17814 & n25528 ;
  assign n25603 = ~\core_eu_ea_alu_ea_reg_ax0rwe_DO_reg[2]/P0001  & ~n25528 ;
  assign n25604 = ~n25602 & ~n25603 ;
  assign n25605 = ~n18974 & n25528 ;
  assign n25606 = ~\core_eu_ea_alu_ea_reg_ax0rwe_DO_reg[1]/P0001  & ~n25528 ;
  assign n25607 = ~n25605 & ~n25606 ;
  assign n25608 = ~n17836 & n25528 ;
  assign n25609 = ~\core_eu_ea_alu_ea_reg_ax0rwe_DO_reg[13]/P0001  & ~n25528 ;
  assign n25610 = ~n25608 & ~n25609 ;
  assign n25611 = ~n23920 & n25528 ;
  assign n25612 = ~\core_eu_ea_alu_ea_reg_ax0rwe_DO_reg[12]/P0001  & ~n25528 ;
  assign n25613 = ~n25611 & ~n25612 ;
  assign n25614 = ~n23757 & n25528 ;
  assign n25615 = ~\core_eu_ea_alu_ea_reg_ax0rwe_DO_reg[11]/P0001  & ~n25528 ;
  assign n25616 = ~n25614 & ~n25615 ;
  assign n25617 = ~n19848 & n25528 ;
  assign n25618 = ~\core_eu_ea_alu_ea_reg_ax0rwe_DO_reg[10]/P0001  & ~n25528 ;
  assign n25619 = ~n25617 & ~n25618 ;
  assign n25620 = ~n19559 & n25528 ;
  assign n25621 = ~\core_eu_ea_alu_ea_reg_ax0rwe_DO_reg[0]/P0001  & ~n25528 ;
  assign n25622 = ~n25620 & ~n25621 ;
  assign n25623 = ~n19972 & n25503 ;
  assign n25624 = ~\core_eu_es_sht_es_reg_sirwe_DO_reg[7]/P0001  & ~n25503 ;
  assign n25625 = ~n25623 & ~n25624 ;
  assign n25626 = ~n20080 & n25503 ;
  assign n25627 = ~\core_eu_es_sht_es_reg_sirwe_DO_reg[4]/P0001  & ~n25503 ;
  assign n25628 = ~n25626 & ~n25627 ;
  assign n25629 = ~n21663 & n25503 ;
  assign n25630 = ~\core_eu_es_sht_es_reg_sirwe_DO_reg[3]/P0001  & ~n25503 ;
  assign n25631 = ~n25629 & ~n25630 ;
  assign n25632 = ~n18974 & n25503 ;
  assign n25633 = ~\core_eu_es_sht_es_reg_sirwe_DO_reg[1]/P0001  & ~n25503 ;
  assign n25634 = ~n25632 & ~n25633 ;
  assign n25635 = ~n20150 & n25503 ;
  assign n25636 = ~\core_eu_es_sht_es_reg_sirwe_DO_reg[14]/P0001  & ~n25503 ;
  assign n25637 = ~n25635 & ~n25636 ;
  assign n25638 = ~n23920 & n25503 ;
  assign n25639 = ~\core_eu_es_sht_es_reg_sirwe_DO_reg[12]/P0001  & ~n25503 ;
  assign n25640 = ~n25638 & ~n25639 ;
  assign n25641 = ~n19848 & n25503 ;
  assign n25642 = ~\core_eu_es_sht_es_reg_sirwe_DO_reg[10]/P0001  & ~n25503 ;
  assign n25643 = ~n25641 & ~n25642 ;
  assign n25644 = ~n20150 & n25528 ;
  assign n25645 = ~\core_eu_ea_alu_ea_reg_ax0rwe_DO_reg[14]/P0001  & ~n25528 ;
  assign n25646 = ~n25644 & ~n25645 ;
  assign n25647 = ~n17820 & n25528 ;
  assign n25648 = ~\core_eu_ea_alu_ea_reg_ax0rwe_DO_reg[15]/P0001  & ~n25528 ;
  assign n25649 = ~n25647 & ~n25648 ;
  assign n25650 = \PIO_oe[8]_pad  & \PIO_oe[9]_pad  ;
  assign n25651 = \memc_MMR_web_reg/NET0131  & n25650 ;
  assign n25652 = \pio_PIO_RES_reg[9]/NET0131  & ~n25651 ;
  assign n25653 = \pio_PIO_RES_OUT_reg[9]/P0001  & n25651 ;
  assign n25654 = ~n25652 & ~n25653 ;
  assign n25655 = \PIO_oe[0]_pad  & \PIO_oe[1]_pad  ;
  assign n25656 = \memc_MMR_web_reg/NET0131  & n25655 ;
  assign n25657 = \pio_PIO_RES_reg[1]/NET0131  & ~n25656 ;
  assign n25658 = \pio_PIO_RES_OUT_reg[1]/P0001  & n25656 ;
  assign n25659 = ~n25657 & ~n25658 ;
  assign n25660 = \PIO_oe[10]_pad  & \PIO_oe[11]_pad  ;
  assign n25661 = \memc_MMR_web_reg/NET0131  & n25660 ;
  assign n25662 = \pio_PIO_RES_reg[11]/NET0131  & ~n25661 ;
  assign n25663 = \pio_PIO_RES_OUT_reg[11]/P0001  & n25661 ;
  assign n25664 = ~n25662 & ~n25663 ;
  assign n25665 = \PIO_oe[2]_pad  & \PIO_oe[3]_pad  ;
  assign n25666 = \memc_MMR_web_reg/NET0131  & n25665 ;
  assign n25667 = \pio_PIO_RES_reg[3]/NET0131  & ~n25666 ;
  assign n25668 = \pio_PIO_RES_OUT_reg[3]/P0001  & n25666 ;
  assign n25669 = ~n25667 & ~n25668 ;
  assign n25670 = \PIO_oe[6]_pad  & \PIO_oe[7]_pad  ;
  assign n25671 = \memc_MMR_web_reg/NET0131  & n25670 ;
  assign n25672 = \pio_PIO_RES_reg[7]/NET0131  & ~n25671 ;
  assign n25673 = \pio_PIO_RES_OUT_reg[7]/P0001  & n25671 ;
  assign n25674 = ~n25672 & ~n25673 ;
  assign n25675 = \pio_PIO_RES_reg[8]/NET0131  & ~n25651 ;
  assign n25676 = \pio_PIO_RES_OUT_reg[8]/P0001  & n25651 ;
  assign n25677 = ~n25675 & ~n25676 ;
  assign n25678 = \PIO_oe[4]_pad  & \PIO_oe[5]_pad  ;
  assign n25679 = \memc_MMR_web_reg/NET0131  & n25678 ;
  assign n25680 = \pio_PIO_RES_reg[5]/NET0131  & ~n25679 ;
  assign n25681 = \pio_PIO_RES_OUT_reg[5]/P0001  & n25679 ;
  assign n25682 = ~n25680 & ~n25681 ;
  assign n25683 = PWDACK_pad & ~\clkc_SLEEP_reg/NET0131  ;
  assign n25684 = \core_c_psq_PCS_reg[7]/NET0131  & n25683 ;
  assign n25685 = \clkc_oscntr_reg_DO_reg[0]/NET0131  & ~n25684 ;
  assign n25686 = ~\clkc_oscntr_reg_DO_reg[0]/NET0131  & n25684 ;
  assign n25687 = ~n25685 & ~n25686 ;
  assign n25688 = \core_c_dec_IR_reg[1]/NET0131  & ~n6023 ;
  assign n25689 = \core_c_dec_IR_reg[5]/NET0131  & n6023 ;
  assign n25690 = ~n25688 & ~n25689 ;
  assign n25691 = ~n4117 & ~n25690 ;
  assign n25692 = \core_dag_ilm2reg_M_E_reg[1]/NET0131  & n4117 ;
  assign n25693 = ~n25691 & ~n25692 ;
  assign n25694 = \core_c_dec_IR_reg[0]/NET0131  & ~n6023 ;
  assign n25695 = \core_c_dec_IR_reg[4]/NET0131  & n6023 ;
  assign n25696 = ~n25694 & ~n25695 ;
  assign n25697 = ~n4117 & ~n25696 ;
  assign n25698 = \core_dag_ilm2reg_M_E_reg[0]/NET0131  & n4117 ;
  assign n25699 = ~n25697 & ~n25698 ;
  assign n25700 = ~n13585 & n13593 ;
  assign n25701 = n13563 & ~n13585 ;
  assign n25702 = ~n13585 & n13590 ;
  assign n25703 = ~n13585 & n13600 ;
  assign n25704 = \tm_tcr_reg_DO_reg[8]/NET0131  & n20355 ;
  assign n25706 = \tm_TCR_TMP_reg[8]/NET0131  & ~n22411 ;
  assign n25707 = ~n22400 & ~n25706 ;
  assign n25708 = ~n23697 & n25707 ;
  assign n25705 = ~\tm_tpr_reg_DO_reg[8]/NET0131  & n22400 ;
  assign n25709 = ~n20355 & ~n25705 ;
  assign n25710 = ~n25708 & n25709 ;
  assign n25711 = ~n25704 & ~n25710 ;
  assign n25712 = ~n11758 & n12232 ;
  assign n25713 = ~n11758 & n12230 ;
  assign n25714 = ~n11758 & n12228 ;
  assign n25715 = ~n11758 & n12225 ;
  assign n25716 = ~n11758 & n12221 ;
  assign n25717 = ~n11758 & n12219 ;
  assign n25718 = ~n11758 & n12216 ;
  assign n25719 = ~n11758 & n12213 ;
  assign n25720 = n11735 & ~n11758 ;
  assign n25721 = ~n13585 & n13607 ;
  assign n25722 = ~n13585 & n13595 ;
  assign n25723 = ~n13585 & n13603 ;
  assign n25724 = ~n13585 & n13605 ;
  assign n25725 = ~n4117 & n6023 ;
  assign n25726 = \core_c_dec_Double_E_reg/P0001  & n4117 ;
  assign n25727 = ~n25725 & ~n25726 ;
  assign n25728 = n4116 & ~n25727 ;
  assign n25730 = ~\core_eu_ec_cun_COND_E_reg[0]/P0001  & n4117 ;
  assign n25729 = ~\core_c_dec_IR_reg[0]/NET0131  & ~n4117 ;
  assign n25731 = n4150 & ~n25729 ;
  assign n25732 = ~n25730 & n25731 ;
  assign n25733 = \core_eu_ec_cun_COND_E_reg[1]/P0001  & n4117 ;
  assign n25734 = \core_c_dec_IR_reg[1]/NET0131  & ~n4117 ;
  assign n25735 = ~n25733 & ~n25734 ;
  assign n25736 = n4150 & ~n25735 ;
  assign n25737 = ~\clkc_Awake_reg/NET0131  & n25042 ;
  assign n25738 = \sport1_cfg_SP_ENg_reg/NET0131  & n23429 ;
  assign n25739 = ~n11739 & ~n11749 ;
  assign n25740 = ~n13581 & ~n13583 ;
  assign n25741 = ~n22981 & n23132 ;
  assign n25745 = n22970 & n23143 ;
  assign n25746 = n25741 & n25745 ;
  assign n25747 = ~n19266 & n25746 ;
  assign n25742 = n22970 & ~n23143 ;
  assign n25743 = n25741 & n25742 ;
  assign n25744 = n19266 & n25743 ;
  assign n25752 = ~n22981 & ~n23132 ;
  assign n25755 = n25742 & n25752 ;
  assign n25756 = ~n19263 & n25755 ;
  assign n25753 = n25745 & n25752 ;
  assign n25754 = n19263 & n25753 ;
  assign n25748 = n22981 & n23132 ;
  assign n25749 = ~n22970 & n23143 ;
  assign n25750 = n25748 & n25749 ;
  assign n25751 = n19296 & n25750 ;
  assign n25757 = ~n22970 & ~n23143 ;
  assign n25758 = n25748 & n25757 ;
  assign n25759 = ~n19296 & n25758 ;
  assign n25760 = ~n25751 & ~n25759 ;
  assign n25761 = ~n25754 & n25760 ;
  assign n25762 = ~n25756 & n25761 ;
  assign n25763 = ~n25744 & n25762 ;
  assign n25764 = ~n25747 & n25763 ;
  assign n25765 = ~n19205 & ~n25764 ;
  assign n25778 = ~n19315 & ~n19337 ;
  assign n25779 = \core_eu_ec_cun_AS_reg/P0001  & n19315 ;
  assign n25780 = ~n25778 & ~n25779 ;
  assign n25782 = ~n23143 & n25780 ;
  assign n25781 = n23143 & ~n25780 ;
  assign n25783 = ~n22970 & n22981 ;
  assign n25784 = ~n23132 & n25783 ;
  assign n25785 = ~n25781 & n25784 ;
  assign n25786 = ~n25782 & n25785 ;
  assign n25767 = \core_eu_ec_cun_AV_reg/P0001  & ~n25755 ;
  assign n25768 = ~\core_eu_ec_cun_AV_reg/P0001  & ~n25753 ;
  assign n25769 = ~n25767 & ~n25768 ;
  assign n25766 = n4137 & n25743 ;
  assign n25770 = ~n4137 & n25746 ;
  assign n25773 = ~n25766 & ~n25770 ;
  assign n25771 = ~\core_eu_ec_cun_AC_reg/P0001  & n25750 ;
  assign n25772 = \core_eu_ec_cun_AC_reg/P0001  & n25758 ;
  assign n25774 = ~n25771 & ~n25772 ;
  assign n25775 = n25773 & n25774 ;
  assign n25776 = ~n25769 & n25775 ;
  assign n25777 = n19205 & ~n25776 ;
  assign n25787 = ~n4117 & ~n25777 ;
  assign n25788 = ~n25786 & n25787 ;
  assign n25789 = ~n25765 & n25788 ;
  assign n25790 = ~\core_eu_ec_cun_termOK_CE_reg/P0001  & n4117 ;
  assign n25791 = n4149 & ~n25790 ;
  assign n25792 = ~n25789 & n25791 ;
  assign n25793 = ~\T_PIOin[3]_pad  & ~\pio_PIO_RES_reg[3]/NET0131  ;
  assign n25794 = \T_PIOin[3]_pad  & \pio_PIO_RES_reg[3]/NET0131  ;
  assign n25795 = ~\pio_PIO_IN_P_reg[3]/P0001  & ~n25794 ;
  assign n25796 = ~n25793 & ~n25795 ;
  assign n25797 = ~\T_PIOin[1]_pad  & ~\pio_PIO_RES_reg[1]/NET0131  ;
  assign n25798 = \T_PIOin[1]_pad  & \pio_PIO_RES_reg[1]/NET0131  ;
  assign n25799 = ~\pio_PIO_IN_P_reg[1]/P0001  & ~n25798 ;
  assign n25800 = ~n25797 & ~n25799 ;
  assign n25801 = ~\T_PIOin[10]_pad  & ~\pio_PIO_RES_reg[10]/NET0131  ;
  assign n25802 = \T_PIOin[10]_pad  & \pio_PIO_RES_reg[10]/NET0131  ;
  assign n25803 = ~\pio_PIO_IN_P_reg[10]/P0001  & ~n25802 ;
  assign n25804 = ~n25801 & ~n25803 ;
  assign n25806 = ~\core_c_dec_Long_Cg_reg/P0001  & n5950 ;
  assign n25805 = ~\core_c_dec_Long_Eg_reg/P0001  & ~n5950 ;
  assign n25807 = n4116 & ~n25805 ;
  assign n25808 = ~n25806 & n25807 ;
  assign n25809 = ~\auctl_T0Sack_reg/NET0131  & n4050 ;
  assign n25810 = ~n4097 & n25809 ;
  assign n25811 = ~\auctl_R1Sack_reg/NET0131  & n11772 ;
  assign n25812 = ~\T_PIOin[8]_pad  & ~\pio_PIO_RES_reg[8]/NET0131  ;
  assign n25813 = \T_PIOin[8]_pad  & \pio_PIO_RES_reg[8]/NET0131  ;
  assign n25814 = ~\pio_PIO_IN_P_reg[8]/P0001  & ~n25813 ;
  assign n25815 = ~n25812 & ~n25814 ;
  assign n25816 = ~\T_PIOin[5]_pad  & ~\pio_PIO_RES_reg[5]/NET0131  ;
  assign n25817 = \T_PIOin[5]_pad  & \pio_PIO_RES_reg[5]/NET0131  ;
  assign n25818 = ~\pio_PIO_IN_P_reg[5]/P0001  & ~n25817 ;
  assign n25819 = ~n25816 & ~n25818 ;
  assign n25820 = ~\T_PIOin[6]_pad  & ~\pio_PIO_RES_reg[6]/NET0131  ;
  assign n25821 = \T_PIOin[6]_pad  & \pio_PIO_RES_reg[6]/NET0131  ;
  assign n25822 = ~\pio_PIO_IN_P_reg[6]/P0001  & ~n25821 ;
  assign n25823 = ~n25820 & ~n25822 ;
  assign n25824 = ~\T_PIOin[11]_pad  & ~\pio_PIO_RES_reg[11]/NET0131  ;
  assign n25825 = \T_PIOin[11]_pad  & \pio_PIO_RES_reg[11]/NET0131  ;
  assign n25826 = ~\pio_PIO_IN_P_reg[11]/P0001  & ~n25825 ;
  assign n25827 = ~n25824 & ~n25826 ;
  assign n25828 = ~\auctl_R0Sack_reg/NET0131  & n11774 ;
  assign n25829 = ~\auctl_T1Sack_reg/NET0131  & n5968 ;
  assign n25830 = ~n4097 & n25829 ;
  assign n25831 = \tm_tcr_reg_DO_reg[15]/NET0131  & n20355 ;
  assign n25833 = ~\tm_TCR_TMP_reg[11]/NET0131  & ~n22417 ;
  assign n25834 = n22424 & n25833 ;
  assign n25835 = \tm_TCR_TMP_reg[11]/NET0131  & n22417 ;
  assign n25836 = ~n22423 & n25835 ;
  assign n25837 = ~\T_TMODE[0]_pad  & ~n25836 ;
  assign n25838 = ~n25834 & n25837 ;
  assign n25839 = n22411 & ~n25838 ;
  assign n25840 = ~\tm_TCR_TMP_reg[12]/NET0131  & n25839 ;
  assign n25841 = ~\tm_TCR_TMP_reg[13]/NET0131  & n25840 ;
  assign n25842 = ~\tm_TCR_TMP_reg[14]/NET0131  & n25841 ;
  assign n25843 = ~\tm_TCR_TMP_reg[15]/NET0131  & ~n25842 ;
  assign n25844 = \tm_TCR_TMP_reg[15]/NET0131  & n25842 ;
  assign n25845 = ~n25843 & ~n25844 ;
  assign n25846 = ~n22400 & ~n25845 ;
  assign n25832 = ~\tm_tpr_reg_DO_reg[15]/NET0131  & n22400 ;
  assign n25847 = ~n20355 & ~n25832 ;
  assign n25848 = ~n25846 & n25847 ;
  assign n25849 = ~n25831 & ~n25848 ;
  assign n25850 = ~\T_TMODE[1]_pad  & \core_c_dec_PPclr_reg/P0001  ;
  assign n25851 = \core_eu_ec_cun_COND_E_reg[2]/P0001  & n4117 ;
  assign n25852 = \core_c_dec_IR_reg[2]/NET0131  & ~n4117 ;
  assign n25853 = ~n25851 & ~n25852 ;
  assign n25854 = n4150 & ~n25853 ;
  assign n25855 = ~\T_PIOin[4]_pad  & ~\pio_PIO_RES_reg[4]/NET0131  ;
  assign n25856 = \T_PIOin[4]_pad  & \pio_PIO_RES_reg[4]/NET0131  ;
  assign n25857 = ~\pio_PIO_IN_P_reg[4]/P0001  & ~n25856 ;
  assign n25858 = ~n25855 & ~n25857 ;
  assign n25859 = ~\T_PIOin[7]_pad  & ~\pio_PIO_RES_reg[7]/NET0131  ;
  assign n25860 = \T_PIOin[7]_pad  & \pio_PIO_RES_reg[7]/NET0131  ;
  assign n25861 = ~\pio_PIO_IN_P_reg[7]/P0001  & ~n25860 ;
  assign n25862 = ~n25859 & ~n25861 ;
  assign n25863 = \core_eu_ec_cun_COND_E_reg[3]/P0001  & n4117 ;
  assign n25864 = \core_c_dec_IR_reg[3]/NET0131  & ~n4117 ;
  assign n25865 = ~n25863 & ~n25864 ;
  assign n25866 = n4150 & ~n25865 ;
  assign n25867 = ~\T_PIOin[9]_pad  & ~\pio_PIO_RES_reg[9]/NET0131  ;
  assign n25868 = \T_PIOin[9]_pad  & \pio_PIO_RES_reg[9]/NET0131  ;
  assign n25869 = ~\pio_PIO_IN_P_reg[9]/P0001  & ~n25868 ;
  assign n25870 = ~n25867 & ~n25869 ;
  assign n25874 = n18470 & ~n23047 ;
  assign n25883 = ~n23060 & n23061 ;
  assign n25882 = ~n23061 & ~n23150 ;
  assign n25884 = ~n23054 & ~n25882 ;
  assign n25885 = ~n25883 & n25884 ;
  assign n25881 = n23043 & n23054 ;
  assign n25886 = ~n23052 & ~n25881 ;
  assign n25887 = ~n25885 & n25886 ;
  assign n25880 = ~n18492 & n23052 ;
  assign n25888 = ~n23051 & ~n25880 ;
  assign n25889 = ~n25887 & n25888 ;
  assign n25878 = ~n18500 & n23051 ;
  assign n25876 = n18471 & ~n18479 ;
  assign n25879 = ~n18481 & ~n25876 ;
  assign n25890 = ~n25878 & n25879 ;
  assign n25891 = ~n25889 & n25890 ;
  assign n25875 = ~n18467 & n18512 ;
  assign n25877 = n18507 & n25876 ;
  assign n25892 = ~n25875 & ~n25877 ;
  assign n25893 = ~n25891 & n25892 ;
  assign n25894 = n25874 & ~n25893 ;
  assign n25873 = ~n18470 & n18479 ;
  assign n25895 = n23047 & ~n23060 ;
  assign n25896 = ~n25873 & ~n25895 ;
  assign n25897 = ~n25894 & n25896 ;
  assign n25898 = \sport0_txctl_ldTX_cmp_reg/P0001  & ~n25897 ;
  assign n25871 = \sport0_txctl_TX_reg[2]/P0001  & n21318 ;
  assign n25872 = n8715 & n21316 ;
  assign n25899 = ~n25871 & ~n25872 ;
  assign n25900 = ~n25898 & n25899 ;
  assign n25901 = ~\T_PIOin[2]_pad  & ~\pio_PIO_RES_reg[2]/NET0131  ;
  assign n25902 = \T_PIOin[2]_pad  & \pio_PIO_RES_reg[2]/NET0131  ;
  assign n25903 = ~\pio_PIO_IN_P_reg[2]/P0001  & ~n25902 ;
  assign n25904 = ~n25901 & ~n25903 ;
  assign n25905 = \T_TMODE[1]_pad  & n20206 ;
  assign n25906 = \T_TMODE[1]_pad  & n5518 ;
  assign n25907 = n5592 & n25906 ;
  assign n25908 = \emc_ECMcs_reg/NET0131  & ~n25907 ;
  assign n25909 = ~n25905 & ~n25908 ;
  assign n25910 = ~\T_PIOin[0]_pad  & ~\pio_PIO_RES_reg[0]/NET0131  ;
  assign n25911 = \T_PIOin[0]_pad  & \pio_PIO_RES_reg[0]/NET0131  ;
  assign n25912 = ~\pio_PIO_IN_P_reg[0]/P0001  & ~n25911 ;
  assign n25913 = ~n25910 & ~n25912 ;
  assign n25914 = \core_c_psq_Eqend_Ed_reg/P0001  & n4094 ;
  assign n25915 = \core_c_psq_Eqend_D_reg/P0001  & ~n4094 ;
  assign n25916 = n11741 & n25915 ;
  assign n25917 = ~n25914 & ~n25916 ;
  assign n25918 = n4116 & ~n25917 ;
  assign n25927 = ~\sport0_txctl_TX_reg[0]/P0001  & ~n18391 ;
  assign n25928 = ~n18392 & ~n25927 ;
  assign n25929 = ~n23061 & n25928 ;
  assign n25926 = n23061 & n23161 ;
  assign n25930 = ~n23054 & ~n25926 ;
  assign n25931 = ~n25929 & n25930 ;
  assign n25932 = n23054 & n23149 ;
  assign n25933 = ~n23052 & ~n25932 ;
  assign n25934 = ~n25931 & n25933 ;
  assign n25925 = n23052 & ~n23059 ;
  assign n25935 = ~n23051 & ~n25925 ;
  assign n25936 = ~n25934 & n25935 ;
  assign n25924 = n23042 & n23051 ;
  assign n25937 = n18457 & ~n25924 ;
  assign n25938 = ~n25936 & n25937 ;
  assign n25939 = n25879 & ~n25938 ;
  assign n25922 = ~n18467 & n18500 ;
  assign n25923 = ~n18492 & n25876 ;
  assign n25940 = ~n25922 & ~n25923 ;
  assign n25941 = ~n25939 & n25940 ;
  assign n25942 = n25874 & ~n25941 ;
  assign n25920 = ~n18470 & n18507 ;
  assign n25921 = n23047 & ~n23162 ;
  assign n25943 = ~n25920 & ~n25921 ;
  assign n25944 = ~n25942 & n25943 ;
  assign n25945 = \sport0_txctl_ldTX_cmp_reg/P0001  & ~n25944 ;
  assign n25919 = \sport0_txctl_TX_reg[0]/P0001  & n21318 ;
  assign n25946 = n7607 & n21316 ;
  assign n25947 = ~n25919 & ~n25946 ;
  assign n25948 = ~n25945 & n25947 ;
  assign n25949 = \core_c_dec_IRE_reg[3]/NET0131  & ~\core_c_psq_PCS_reg[7]/NET0131  ;
  assign n25950 = n4115 & n25949 ;
  assign n25951 = PWDACK_pad & ~\clkc_Awake_reg/NET0131  ;
  assign n25952 = \core_c_psq_PCS_reg[7]/NET0131  & n25951 ;
  assign n25953 = ~n25950 & ~n25952 ;
  assign n25954 = \core_c_dec_MTLreg_E_reg[4]/P0001  & n5951 ;
  assign n25955 = \core_c_dec_MTLreg_E_reg[5]/P0001  & n5951 ;
  assign n25956 = \core_c_dec_rdCM_E_reg/NET0131  & n4117 ;
  assign n25957 = ~\core_c_dec_IR_reg[20]/NET0131  & n5888 ;
  assign n25958 = ~n25956 & ~n25957 ;
  assign n25959 = \core_c_dec_MTLreg_E_reg[7]/P0001  & n5951 ;
  assign n25960 = ~\core_c_psq_PCS_reg[7]/NET0131  & n11736 ;
  assign n25961 = ~n13760 & ~n25960 ;
  assign n25962 = \memc_usysr_DO_reg[11]/NET0131  & \sport1_regs_MWORDreg_DO_reg[9]/NET0131  ;
  assign n25963 = ~\sport1_txctl_SP_EN_D1_reg/P0001  & n25962 ;
  assign n25964 = ~\sport1_txctl_TSreqi_reg/NET0131  & ~n25963 ;
  assign n25965 = \core_c_dec_MTLreg_E_reg[6]/P0001  & n5951 ;
  assign n25966 = \memc_usysr_DO_reg[12]/NET0131  & \sport0_regs_MWORDreg_DO_reg[9]/NET0131  ;
  assign n25967 = ~\sport0_txctl_SP_EN_D1_reg/P0001  & n25966 ;
  assign n25968 = ~\sport0_txctl_TSreqi_reg/NET0131  & ~n25967 ;
  assign n25969 = ~IACKn_pad & \sice_RCS_reg[0]/NET0131  ;
  assign n25970 = ~\sice_RCS_reg[1]/NET0131  & n25969 ;
  assign n25971 = ~\sice_RCS_reg[0]/NET0131  & \sice_RCS_reg[1]/NET0131  ;
  assign n25972 = ~n25970 & ~n25971 ;
  assign n25973 = \core_c_dec_MTLreg_E_reg[2]/P0001  & n5951 ;
  assign n25974 = \core_c_dec_MTLreg_E_reg[1]/P0001  & n5951 ;
  assign n25975 = \core_c_dec_MTLreg_E_reg[0]/P0001  & n5951 ;
  assign n25976 = \core_c_dec_MTLreg_E_reg[3]/P0001  & n5951 ;
  assign n25977 = \core_c_psq_Iact_E_reg[10]/NET0131  & ~n19477 ;
  assign n25978 = \core_c_psq_Iflag_reg[10]/NET0131  & ~\core_c_psq_PCS_reg[3]/NET0131  ;
  assign n25979 = n19477 & n25978 ;
  assign n25980 = ~n25977 & ~n25979 ;
  assign n25981 = \clkc_SLEEP_reg/NET0131  & \core_c_psq_PCS_reg[7]/NET0131  ;
  assign n25982 = ~n25950 & ~n25981 ;
  assign n25983 = ~n13806 & ~n14610 ;
  assign n25984 = n13806 & ~n14586 ;
  assign n25985 = ~n25983 & ~n25984 ;
  assign n25986 = n14667 & ~n25985 ;
  assign n25987 = \core_eu_ea_alu_ea_reg_afswe_DO_reg[3]/P0001  & ~n14667 ;
  assign n25988 = ~n25986 & ~n25987 ;
  assign n25989 = \core_c_dec_MTICNTL_Eg_reg/P0001  & ~n5950 ;
  assign n25990 = ~n10069 & n25989 ;
  assign n25991 = ~\core_c_psq_ICNTL_reg_DO_reg[4]/NET0131  & ~n25989 ;
  assign n25992 = ~n25990 & ~n25991 ;
  assign n25993 = ~n8715 & n25989 ;
  assign n25994 = ~\core_c_psq_ICNTL_reg_DO_reg[2]/NET0131  & ~n25989 ;
  assign n25995 = ~n25993 & ~n25994 ;
  assign n25996 = n13805 & ~n25985 ;
  assign n25997 = \core_eu_ea_alu_ea_reg_afrwe_DO_reg[3]/P0001  & ~n13805 ;
  assign n25998 = ~n25996 & ~n25997 ;
  assign n25999 = \memc_STI_Cg_reg/NET0131  & n5950 ;
  assign n26000 = ~n5946 & ~n13130 ;
  assign n26001 = n5951 & ~n26000 ;
  assign n26002 = ~n25999 & ~n26001 ;
  assign n26004 = n19499 & ~n20259 ;
  assign n26003 = ~\core_eu_em_mac_em_reg_mr1swe_DO_reg[5]/P0001  & ~n19499 ;
  assign n26005 = n19501 & ~n26003 ;
  assign n26006 = ~n26004 & n26005 ;
  assign n26007 = \core_eu_em_mac_em_reg_mr1swe_DO_reg[5]/P0001  & ~n19383 ;
  assign n26008 = ~n19508 & ~n26007 ;
  assign n26009 = ~n26006 & n26008 ;
  assign n26010 = ~n18262 & ~n26009 ;
  assign n26011 = ~n17543 & ~n19422 ;
  assign n26012 = ~n17676 & ~n26011 ;
  assign n26013 = ~n17474 & ~n17677 ;
  assign n26014 = ~n26012 & n26013 ;
  assign n26015 = n26012 & ~n26013 ;
  assign n26016 = ~n26014 & ~n26015 ;
  assign n26017 = ~\core_c_psq_MSTAT_reg_DO_reg[4]/NET0131  & n26016 ;
  assign n26018 = \core_c_psq_MSTAT_reg_DO_reg[4]/NET0131  & n23218 ;
  assign n26019 = ~n26017 & ~n26018 ;
  assign n26020 = n18262 & ~n26019 ;
  assign n26021 = ~n26010 & ~n26020 ;
  assign n26022 = \tm_TSR_TMP_reg[6]/NET0131  & ~n25495 ;
  assign n26023 = ~n25496 & ~n26022 ;
  assign n26024 = n25491 & ~n26023 ;
  assign n26025 = \tm_tsr_reg_DO_reg[6]/NET0131  & ~n25491 ;
  assign n26026 = ~n26024 & ~n26025 ;
  assign n26027 = \memc_Pwrite_E_reg/NET0131  & ~n5950 ;
  assign n26028 = ~\core_c_psq_PCS_reg[7]/NET0131  & n13565 ;
  assign n26029 = ~n26027 & ~n26028 ;
  assign n26030 = \core_c_psq_PCS_reg[7]/NET0131  & ~\core_c_psq_TRAP_R_L_reg/NET0131  ;
  assign n26031 = \clkc_STBY_reg/NET0131  & n26030 ;
  assign n26032 = ~\core_c_dec_IRE_reg[3]/NET0131  & ~\core_c_psq_PCS_reg[7]/NET0131  ;
  assign n26033 = n4115 & n26032 ;
  assign n26034 = ~n26031 & ~n26033 ;
  assign n26035 = n14752 & n26019 ;
  assign n26036 = n19776 & n20259 ;
  assign n26037 = \core_eu_em_mac_em_reg_mr1rwe_DO_reg[5]/P0001  & ~n17809 ;
  assign n26038 = n19780 & ~n26037 ;
  assign n26039 = ~n26036 & n26038 ;
  assign n26040 = ~n26035 & ~n26039 ;
  assign n26041 = ~\sice_IIRC_reg[0]/NET0131  & ~\sice_IIRC_reg[1]/NET0131  ;
  assign n26042 = ~n18865 & ~n26041 ;
  assign n26043 = ~\sice_ICYC_reg[0]/NET0131  & ~\sice_ICYC_reg[1]/NET0131  ;
  assign n26044 = ~n18856 & ~n26043 ;
  assign n26045 = ~\clkc_oscntr_reg_DO_reg[0]/NET0131  & ~\clkc_oscntr_reg_DO_reg[1]/NET0131  ;
  assign n26046 = ~n20845 & ~n26045 ;
  assign n26047 = \core_eu_em_mac_em_reg_mfswe_DO_reg[5]/P0001  & ~n20864 ;
  assign n26048 = n20864 & ~n26019 ;
  assign n26049 = ~n26047 & ~n26048 ;
  assign n26050 = n12743 & n25097 ;
  assign n26051 = n19045 & n25202 ;
  assign n26052 = n5524 & n5575 ;
  assign n26053 = n12688 & n25097 ;
  assign n26054 = ~\clkc_SIDLE_s2_reg/NET0131  & ~\clkc_STBY_reg/NET0131  ;
  assign n26055 = n12241 & ~n26054 ;
  assign n26056 = \core_eu_em_mac_em_reg_mfrwe_DO_reg[5]/P0001  & ~n20990 ;
  assign n26057 = n20990 & ~n26019 ;
  assign n26058 = ~n26056 & ~n26057 ;
  assign n26059 = \core_c_dec_MTMreg_E_reg[6]/P0001  & n5951 ;
  assign n26060 = \core_c_dec_MTMreg_E_reg[5]/P0001  & n5951 ;
  assign n26061 = ~\core_c_psq_PCS_reg[3]/NET0131  & n4098 ;
  assign n26062 = ~\auctl_DSack_reg/NET0131  & n5068 ;
  assign n26063 = ~n26061 & n26062 ;
  assign n26064 = ~T_IMS_pad & \sice_ICS_reg[1]/NET0131  ;
  assign n26065 = ~\sice_ICS_reg[2]/NET0131  & n26064 ;
  assign n26066 = n7340 & n25097 ;
  assign n26067 = ~\auctl_BSack_reg/NET0131  & n5644 ;
  assign n26068 = ~\auctl_DSack_reg/NET0131  & ~\auctl_RST_reg/P0001  ;
  assign n26069 = \clkc_DSPoff_reg/NET0131  & \clkc_SLEEP_reg/NET0131  ;
  assign n26070 = \sport0_regs_AUTO_a_reg[15]/NET0131  & n26069 ;
  assign n26071 = n9178 & n25097 ;
  assign n26072 = \core_eu_ec_cun_mven_FFout_reg/NET0131  & n12245 ;
  assign n26073 = n4149 & ~n26072 ;
  assign n26074 = \core_c_dec_MTMreg_E_reg[7]/P0001  & n5951 ;
  assign n26075 = \core_c_dec_MTMreg_E_reg[4]/P0001  & n5951 ;
  assign n26076 = \core_c_dec_MTMreg_E_reg[1]/P0001  & n5951 ;
  assign n26077 = \core_c_dec_MTMreg_E_reg[3]/P0001  & n5951 ;
  assign n26078 = ~\auctl_BSack_reg/NET0131  & ~\auctl_RST_reg/P0001  ;
  assign n26079 = \core_c_dec_MTMreg_E_reg[2]/P0001  & n5951 ;
  assign n26080 = \core_c_dec_MTMreg_E_reg[0]/P0001  & n5951 ;
  assign n26081 = ~\core_c_psq_PCS2or3_reg/NET0131  & ~\core_c_psq_PCS_reg[4]/NET0131  ;
  assign n26082 = \auctl_STEAL_reg/NET0131  & ~n26081 ;
  assign n26083 = ~\clkc_SIDLE_s1_reg/NET0131  & \clkc_SIDLE_s2_reg/NET0131  ;
  assign n26084 = \core_c_psq_PCS_reg[7]/NET0131  & ~n26083 ;
  assign n26085 = \bdma_RST_pin_reg/P0001  & ~n13733 ;
  assign n26086 = \core_c_dec_IRE_reg[3]/NET0131  & n4117 ;
  assign n26087 = ~n25864 & ~n26086 ;
  assign n26088 = T_BMODE_pad & ~T_MMAP_pad ;
  assign n26089 = \bdma_RST_pin_reg/P0001  & ~n26088 ;
  assign n26090 = \bdma_RST_pin_reg/P0001  & n26088 ;
  assign n26091 = \core_c_dec_IRE_reg[2]/NET0131  & n4117 ;
  assign n26092 = ~n25852 & ~n26091 ;
  assign n26093 = ~\bdma_BDMAmode_reg/NET0131  & ~n4116 ;
  assign n26094 = n4149 & ~n26093 ;
  assign n26095 = ~\core_c_dec_Dummy_E_reg/NET0131  & n4117 ;
  assign n26096 = ~n11742 & ~n26095 ;
  assign n26097 = ~\core_c_dec_accPM_E_reg/P0001  & \core_dag_ilm1reg_DMA_pi_DO_reg[2]/NET0131  ;
  assign n26098 = \core_c_dec_accPM_E_reg/P0001  & \core_dag_ilm2reg_PMA_pi_DO_reg[2]/NET0131  ;
  assign n26099 = ~n26097 & ~n26098 ;
  assign n26100 = \core_c_dec_IR_reg[0]/NET0131  & ~n4117 ;
  assign n26101 = \core_c_dec_IRE_reg[0]/NET0131  & n4117 ;
  assign n26102 = ~n26100 & ~n26101 ;
  assign n26103 = \core_c_dec_IRE_reg[1]/NET0131  & n4117 ;
  assign n26104 = ~n25734 & ~n26103 ;
  assign n26105 = ~\core_c_dec_accPM_E_reg/P0001  & \core_dag_ilm1reg_DMA_pi_DO_reg[3]/NET0131  ;
  assign n26106 = \core_c_dec_accPM_E_reg/P0001  & \core_dag_ilm2reg_PMA_pi_DO_reg[3]/NET0131  ;
  assign n26107 = ~n26105 & ~n26106 ;
  assign n26108 = ~\core_c_dec_accPM_E_reg/P0001  & \core_dag_ilm1reg_DMA_pi_DO_reg[4]/NET0131  ;
  assign n26109 = \core_c_dec_accPM_E_reg/P0001  & \core_dag_ilm2reg_PMA_pi_DO_reg[4]/NET0131  ;
  assign n26110 = ~n26108 & ~n26109 ;
  assign n26111 = ~\core_c_dec_accPM_E_reg/P0001  & \core_dag_ilm1reg_DMA_pi_DO_reg[0]/NET0131  ;
  assign n26112 = \core_c_dec_accPM_E_reg/P0001  & \core_dag_ilm2reg_PMA_pi_DO_reg[0]/NET0131  ;
  assign n26113 = ~n26111 & ~n26112 ;
  assign n26114 = ~\core_c_dec_accPM_E_reg/P0001  & \core_dag_ilm1reg_DMA_pi_DO_reg[1]/NET0131  ;
  assign n26115 = \core_c_dec_accPM_E_reg/P0001  & \core_dag_ilm2reg_PMA_pi_DO_reg[1]/NET0131  ;
  assign n26116 = ~n26114 & ~n26115 ;
  assign n26117 = ~\tm_tsr_reg_DO_reg[8]/NET0131  & ~n12245 ;
  assign n26118 = \tm_tsr_reg_DO_reg[8]/NET0131  & ~n12241 ;
  assign n26119 = ~n26117 & ~n26118 ;
  assign n26120 = ~\clkc_DSPoff_reg/NET0131  & \clkc_SLEEP_reg/NET0131  ;
  assign n26121 = ~\clkc_Cnt4096_reg/NET0131  & \clkc_DSPoff_reg/NET0131  ;
  assign n26122 = ~n26120 & ~n26121 ;
  assign n26123 = \sport1_txctl_TXSHT_reg[13]/P0001  & ~n22677 ;
  assign n26124 = \sport1_txctl_TX_reg[14]/P0001  & n22677 ;
  assign n26125 = ~n26123 & ~n26124 ;
  assign n26126 = n4094 & n4116 ;
  assign n26127 = ~n5635 & ~n26126 ;
  assign n26128 = \core_c_psq_IFA_reg[12]/P0001  & n26126 ;
  assign n26129 = ~n26127 & ~n26128 ;
  assign n26130 = ~n5419 & ~n26126 ;
  assign n26131 = \core_c_psq_IFA_reg[9]/P0001  & n26126 ;
  assign n26132 = ~n26130 & ~n26131 ;
  assign n26133 = ~n5338 & ~n26126 ;
  assign n26134 = \core_c_psq_IFA_reg[6]/P0001  & n26126 ;
  assign n26135 = ~n26133 & ~n26134 ;
  assign n26136 = ~n5311 & ~n26126 ;
  assign n26137 = \core_c_psq_IFA_reg[5]/P0001  & n26126 ;
  assign n26138 = ~n26136 & ~n26137 ;
  assign n26139 = ~n5208 & ~n26126 ;
  assign n26140 = \core_c_psq_IFA_reg[2]/P0001  & n26126 ;
  assign n26141 = ~n26139 & ~n26140 ;
  assign n26142 = ~n5169 & ~n26126 ;
  assign n26143 = \core_c_psq_IFA_reg[1]/P0001  & n26126 ;
  assign n26144 = ~n26142 & ~n26143 ;
  assign n26145 = ~n5142 & ~n26126 ;
  assign n26146 = \core_c_psq_IFA_reg[11]/P0001  & n26126 ;
  assign n26147 = ~n26145 & ~n26146 ;
  assign n26148 = ~n5064 & ~n26126 ;
  assign n26149 = \core_c_psq_IFA_reg[0]/P0001  & n26126 ;
  assign n26150 = ~n26148 & ~n26149 ;
  assign n26151 = \core_c_psq_DRA_reg[7]/P0001  & ~n4094 ;
  assign n26152 = \core_c_psq_EXA_reg[7]/P0001  & n4094 ;
  assign n26153 = ~n26151 & ~n26152 ;
  assign n26154 = \core_c_psq_DRA_reg[6]/P0001  & ~n4094 ;
  assign n26155 = \core_c_psq_EXA_reg[6]/P0001  & n4094 ;
  assign n26156 = ~n26154 & ~n26155 ;
  assign n26157 = \core_c_psq_DRA_reg[3]/P0001  & ~n4094 ;
  assign n26158 = \core_c_psq_EXA_reg[3]/P0001  & n4094 ;
  assign n26159 = ~n26157 & ~n26158 ;
  assign n26160 = \core_c_psq_DRA_reg[2]/P0001  & ~n4094 ;
  assign n26161 = \core_c_psq_EXA_reg[2]/P0001  & n4094 ;
  assign n26162 = ~n26160 & ~n26161 ;
  assign n26163 = \core_c_psq_DRA_reg[13]/P0001  & ~n4094 ;
  assign n26164 = \core_c_psq_EXA_reg[13]/P0001  & n4094 ;
  assign n26165 = ~n26163 & ~n26164 ;
  assign n26166 = \core_c_psq_DRA_reg[12]/P0001  & ~n4094 ;
  assign n26167 = \core_c_psq_EXA_reg[12]/P0001  & n4094 ;
  assign n26168 = ~n26166 & ~n26167 ;
  assign n26169 = \core_c_dec_accCM_E_reg/NET0131  & n4117 ;
  assign n26170 = ~n5888 & ~n26169 ;
  assign n26171 = ~n5245 & ~n26126 ;
  assign n26172 = \core_c_psq_IFA_reg[3]/P0001  & n26126 ;
  assign n26173 = ~n26171 & ~n26172 ;
  assign n26174 = \core_c_psq_DRA_reg[0]/P0001  & ~n4094 ;
  assign n26175 = \core_c_psq_EXA_reg[0]/P0001  & n4094 ;
  assign n26176 = ~n26174 & ~n26175 ;
  assign n26177 = n4829 & ~n5950 ;
  assign n26178 = \core_c_dec_Prderr_Cg_reg/NET0131  & n5950 ;
  assign n26179 = ~n26177 & ~n26178 ;
  assign n26180 = \core_c_psq_DRA_reg[9]/P0001  & ~n4094 ;
  assign n26181 = \core_c_psq_EXA_reg[9]/P0001  & n4094 ;
  assign n26182 = ~n26180 & ~n26181 ;
  assign n26183 = \core_c_dec_IR_reg[18]/NET0131  & ~n4117 ;
  assign n26184 = \core_c_dec_IRE_reg[18]/NET0131  & n4117 ;
  assign n26185 = ~n26183 & ~n26184 ;
  assign n26186 = \core_c_dec_IR_reg[19]/NET0131  & ~n4117 ;
  assign n26187 = \core_c_dec_IRE_reg[19]/NET0131  & n4117 ;
  assign n26188 = ~n26186 & ~n26187 ;
  assign n26189 = ~n5365 & ~n26126 ;
  assign n26190 = \core_c_psq_IFA_reg[7]/P0001  & n26126 ;
  assign n26191 = ~n26189 & ~n26190 ;
  assign n26192 = \sport1_txctl_TXSHT_reg[14]/P0001  & ~n22677 ;
  assign n26193 = \sport1_txctl_TX_reg[15]/P0001  & n22677 ;
  assign n26194 = ~n26192 & ~n26193 ;
  assign n26195 = ~n4117 & ~n6033 ;
  assign n26196 = \core_dag_ilm2reg_IL_E_reg[1]/P0001  & n4117 ;
  assign n26197 = ~n26195 & ~n26196 ;
  assign n26198 = ~n4117 & ~n6036 ;
  assign n26199 = \core_dag_ilm2reg_IL_E_reg[0]/P0001  & n4117 ;
  assign n26200 = ~n26198 & ~n26199 ;
  assign n26201 = n4099 & ~n5981 ;
  assign n26202 = \core_dag_ilm1reg_STEALI_E_reg[2]/P0001  & ~n4099 ;
  assign n26203 = ~n26201 & ~n26202 ;
  assign n26204 = n4099 & ~n5974 ;
  assign n26205 = \core_dag_ilm1reg_STEALI_E_reg[1]/P0001  & ~n4099 ;
  assign n26206 = ~n26204 & ~n26205 ;
  assign n26207 = n4099 & ~n5989 ;
  assign n26208 = \core_dag_ilm1reg_STEALI_E_reg[0]/P0001  & ~n4099 ;
  assign n26209 = ~n26207 & ~n26208 ;
  assign n26210 = \sport1_txctl_TXSHT_reg[12]/P0001  & ~n22677 ;
  assign n26211 = \sport1_txctl_TX_reg[13]/P0001  & n22677 ;
  assign n26212 = ~n26210 & ~n26211 ;
  assign n26213 = \core_c_psq_DRA_reg[1]/P0001  & ~n4094 ;
  assign n26214 = \core_c_psq_EXA_reg[1]/P0001  & n4094 ;
  assign n26215 = ~n26213 & ~n26214 ;
  assign n26216 = \core_c_psq_DRA_reg[10]/P0001  & ~n4094 ;
  assign n26217 = \core_c_psq_EXA_reg[10]/P0001  & n4094 ;
  assign n26218 = ~n26216 & ~n26217 ;
  assign n26219 = \core_c_psq_DRA_reg[11]/P0001  & ~n4094 ;
  assign n26220 = \core_c_psq_EXA_reg[11]/P0001  & n4094 ;
  assign n26221 = ~n26219 & ~n26220 ;
  assign n26222 = \core_c_psq_DRA_reg[5]/P0001  & ~n4094 ;
  assign n26223 = \core_c_psq_EXA_reg[5]/P0001  & n4094 ;
  assign n26224 = ~n26222 & ~n26223 ;
  assign n26225 = \core_c_psq_DRA_reg[4]/P0001  & ~n4094 ;
  assign n26226 = \core_c_psq_EXA_reg[4]/P0001  & n4094 ;
  assign n26227 = ~n26225 & ~n26226 ;
  assign n26228 = \core_c_psq_DRA_reg[8]/P0001  & ~n4094 ;
  assign n26229 = \core_c_psq_EXA_reg[8]/P0001  & n4094 ;
  assign n26230 = ~n26228 & ~n26229 ;
  assign n26231 = ~n5113 & ~n26126 ;
  assign n26232 = \core_c_psq_IFA_reg[10]/P0001  & n26126 ;
  assign n26233 = ~n26231 & ~n26232 ;
  assign n26234 = ~n5660 & ~n26126 ;
  assign n26235 = \core_c_psq_IFA_reg[13]/P0001  & n26126 ;
  assign n26236 = ~n26234 & ~n26235 ;
  assign n26237 = ~n5279 & ~n26126 ;
  assign n26238 = \core_c_psq_IFA_reg[4]/P0001  & n26126 ;
  assign n26239 = ~n26237 & ~n26238 ;
  assign n26240 = ~n5392 & ~n26126 ;
  assign n26241 = \core_c_psq_IFA_reg[8]/P0001  & n26126 ;
  assign n26242 = ~n26240 & ~n26241 ;
  assign n26245 = ~\sport0_rxctl_ldRX_cmp_reg/P0001  & n9435 ;
  assign n26246 = ~n20938 & ~n20943 ;
  assign n26247 = ~n20880 & ~n26246 ;
  assign n26248 = ~\sport0_rxctl_RX_reg[7]/P0001  & ~n20953 ;
  assign n26250 = ~n26247 & n26248 ;
  assign n26249 = n26247 & ~n26248 ;
  assign n26251 = n20875 & ~n26249 ;
  assign n26252 = ~n26250 & n26251 ;
  assign n26244 = \sport0_rxctl_RX_reg[1]/P0001  & n20873 ;
  assign n26253 = ~n20868 & ~n26244 ;
  assign n26254 = ~n26252 & n26253 ;
  assign n26255 = ~n26245 & n26254 ;
  assign n26243 = ~\sport0_rxctl_RXSHT_reg[1]/P0001  & n20868 ;
  assign n26256 = ~n20871 & ~n26243 ;
  assign n26257 = ~n26255 & n26256 ;
  assign n26258 = \sport0_rxctl_RX_reg[1]/P0001  & n20871 ;
  assign n26259 = ~n26257 & ~n26258 ;
  assign n26260 = \core_c_dec_MTSE_E_reg/P0001  & ~n18974 ;
  assign n26261 = ~n23630 & n23634 ;
  assign n26262 = n23620 & ~n23625 ;
  assign n26264 = n23610 & n23613 ;
  assign n26263 = n23604 & n23607 ;
  assign n26265 = n23585 & n26263 ;
  assign n26266 = ~n26264 & n26265 ;
  assign n26267 = n26262 & ~n26266 ;
  assign n26268 = n26261 & ~n26267 ;
  assign n26269 = n23638 & n23642 ;
  assign n26270 = ~n26268 & n26269 ;
  assign n26271 = n23646 & n23650 ;
  assign n26272 = ~n26270 & n26271 ;
  assign n26273 = n23654 & n23658 ;
  assign n26274 = ~n26272 & n26273 ;
  assign n26275 = n23662 & n23670 ;
  assign n26276 = ~n26274 & n26275 ;
  assign n26277 = ~\core_c_dec_MTSE_E_reg/P0001  & ~n26276 ;
  assign n26278 = ~n26260 & ~n26277 ;
  assign n26279 = n23677 & ~n26278 ;
  assign n26280 = ~\core_eu_es_sht_es_reg_seswe_DO_reg[1]/P0001  & ~n23677 ;
  assign n26281 = ~n26279 & ~n26280 ;
  assign n26282 = n23598 & ~n26278 ;
  assign n26283 = ~\core_eu_es_sht_es_reg_serwe_DO_reg[1]/P0001  & ~n23598 ;
  assign n26284 = ~n26282 & ~n26283 ;
  assign n26285 = ~\clkc_CTR_cnt_reg[0]/NET0131  & \clkc_CTR_cnt_reg[1]/NET0131  ;
  assign n26286 = ~n24968 & ~n26285 ;
  assign n26287 = ~\auctl_R0Sack_reg/NET0131  & ~\auctl_RST_reg/P0001  ;
  assign n26288 = ~\auctl_RST_reg/P0001  & ~\auctl_T0Sack_reg/NET0131  ;
  assign n26289 = ~\auctl_R1Sack_reg/NET0131  & ~\auctl_RST_reg/P0001  ;
  assign n26290 = \sice_ICYC_en_syn_reg/P0001  & n12245 ;
  assign n26291 = ~\auctl_RST_reg/P0001  & ~\auctl_T1Sack_reg/NET0131  ;
  assign n26292 = n4116 & n4149 ;
  assign n26294 = ~\sice_ICS_reg[0]/NET0131  & ~\sice_ICS_reg[1]/NET0131  ;
  assign n26293 = \sice_ICS_reg[0]/NET0131  & \sice_ICS_reg[1]/NET0131  ;
  assign n26295 = T_IMS_pad & ~n26293 ;
  assign n26296 = ~n26294 & n26295 ;
  assign n26297 = \sice_ICS_reg[2]/NET0131  & ~n26296 ;
  assign n26298 = \sice_ICS_reg[0]/NET0131  & ~\sice_ICS_reg[2]/NET0131  ;
  assign n26299 = ~n23030 & ~n26064 ;
  assign n26300 = n26298 & n26299 ;
  assign n26301 = ~n26297 & ~n26300 ;
  assign n26302 = n12234 & ~n26301 ;
  assign n26304 = n19499 & ~n20080 ;
  assign n26303 = ~\core_eu_em_mac_em_reg_mr1swe_DO_reg[4]/P0001  & ~n19499 ;
  assign n26305 = n19501 & ~n26303 ;
  assign n26306 = ~n26304 & n26305 ;
  assign n26307 = \core_eu_em_mac_em_reg_mr1swe_DO_reg[4]/P0001  & ~n19383 ;
  assign n26308 = ~n19508 & ~n26307 ;
  assign n26309 = ~n26306 & n26308 ;
  assign n26310 = ~n18262 & ~n26309 ;
  assign n26311 = \core_c_psq_MSTAT_reg_DO_reg[4]/NET0131  & n26016 ;
  assign n26312 = ~n17543 & ~n17676 ;
  assign n26313 = n19422 & ~n26312 ;
  assign n26314 = ~n19422 & n26312 ;
  assign n26315 = ~n26313 & ~n26314 ;
  assign n26316 = ~\core_c_psq_MSTAT_reg_DO_reg[4]/NET0131  & n26315 ;
  assign n26317 = ~n26311 & ~n26316 ;
  assign n26318 = n18262 & ~n26317 ;
  assign n26319 = ~n26310 & ~n26318 ;
  assign n26320 = ~\clkc_ckr_reg_DO_reg[15]/NET0131  & n12245 ;
  assign n26321 = n14752 & n26317 ;
  assign n26322 = n19776 & n20080 ;
  assign n26323 = \core_eu_em_mac_em_reg_mr1rwe_DO_reg[4]/P0001  & ~n17809 ;
  assign n26324 = n19780 & ~n26323 ;
  assign n26325 = ~n26322 & n26324 ;
  assign n26326 = ~n26321 & ~n26325 ;
  assign n26327 = ~T_ISn_pad & ~T_IWRn_pad ;
  assign n26329 = T_IMS_pad & ~n23031 ;
  assign n26331 = \sice_ICS_reg[1]/NET0131  & n26329 ;
  assign n26328 = ~\sice_ICS_reg[2]/NET0131  & n26294 ;
  assign n26330 = ~\sice_ICS_reg[1]/NET0131  & ~n26329 ;
  assign n26332 = ~n26328 & ~n26330 ;
  assign n26333 = ~n26331 & n26332 ;
  assign n26334 = n12234 & n26333 ;
  assign n26335 = ~\sice_ICS_reg[1]/NET0131  & n26298 ;
  assign n26336 = ~T_IMS_pad & ~n26335 ;
  assign n26337 = n12234 & n26336 ;
  assign n26338 = ~\sice_ICYC_clr_reg/NET0131  & n4149 ;
  assign n26357 = \core_c_dec_updSR_E_reg/P0001  & n13803 ;
  assign n26362 = ~\core_c_dec_Dummy_E_reg/NET0131  & \core_c_dec_MTSR1_E_reg/P0001  ;
  assign n26363 = ~n26357 & ~n26362 ;
  assign n26356 = \core_c_dec_IR_reg[10]/NET0131  & \core_c_dec_IR_reg[9]/NET0131  ;
  assign n26364 = \core_c_dec_IR_reg[8]/NET0131  & n26356 ;
  assign n26365 = ~n26363 & n26364 ;
  assign n26358 = n18846 & n21525 ;
  assign n26359 = \core_c_dec_IR_reg[8]/NET0131  & ~n26358 ;
  assign n26360 = n26356 & ~n26359 ;
  assign n26361 = n26357 & n26360 ;
  assign n26350 = \core_c_dec_updAR_E_reg/P0001  & ~n13802 ;
  assign n26351 = ~\core_c_dec_MTAR_E_reg/P0001  & ~n26350 ;
  assign n26352 = ~\core_c_dec_IR_reg[10]/NET0131  & ~\core_c_dec_IR_reg[8]/NET0131  ;
  assign n26353 = \core_c_dec_IR_reg[9]/NET0131  & n26352 ;
  assign n26354 = ~\core_c_dec_Dummy_E_reg/NET0131  & n26353 ;
  assign n26355 = ~n26351 & n26354 ;
  assign n26339 = ~\core_c_dec_IR_reg[10]/NET0131  & \core_c_dec_IR_reg[8]/NET0131  ;
  assign n26340 = ~n18264 & n26339 ;
  assign n26341 = ~\core_c_dec_Dummy_E_reg/NET0131  & \core_c_dec_IR_reg[10]/NET0131  ;
  assign n26342 = ~\core_c_dec_IR_reg[8]/NET0131  & \core_c_dec_MTSR0_E_reg/P0001  ;
  assign n26343 = n26341 & n26342 ;
  assign n26344 = ~n26340 & ~n26343 ;
  assign n26345 = \core_c_dec_IR_reg[9]/NET0131  & ~n26344 ;
  assign n26346 = \core_c_dec_IR_reg[10]/NET0131  & ~\core_c_dec_IR_reg[9]/NET0131  ;
  assign n26347 = \core_c_dec_IR_reg[8]/NET0131  & n17801 ;
  assign n26348 = n17805 & ~n26347 ;
  assign n26349 = n26346 & ~n26348 ;
  assign n26366 = ~n26345 & ~n26349 ;
  assign n26367 = ~n26355 & n26366 ;
  assign n26368 = ~n26361 & n26367 ;
  assign n26369 = ~n26365 & n26368 ;
  assign n26370 = n18847 & ~n26369 ;
  assign n26371 = \core_c_dec_IR_reg[9]/NET0131  & n26339 ;
  assign n26372 = n18263 & n26371 ;
  assign n26373 = ~\core_c_dec_IR_reg[8]/NET0131  & ~\core_c_dec_IR_reg[9]/NET0131  ;
  assign n26374 = \core_c_dec_MTMR1_E_reg/P0001  & n26341 ;
  assign n26375 = n26373 & n26374 ;
  assign n26376 = ~n26372 & ~n26375 ;
  assign n26377 = n26370 & ~n26376 ;
  assign n26378 = ~n5689 & n26377 ;
  assign n26379 = ~n5689 & n26346 ;
  assign n26380 = \core_c_dec_IR_reg[8]/NET0131  & n26379 ;
  assign n26381 = n17802 & n26380 ;
  assign n26382 = n26370 & n26381 ;
  assign n26383 = ~n26378 & ~n26382 ;
  assign n26384 = n26346 & n26347 ;
  assign n26385 = n18847 & n26384 ;
  assign n26386 = \core_c_dec_accPM_E_reg/P0001  & n26385 ;
  assign n26387 = ~n5689 & n26386 ;
  assign n26388 = n26383 & ~n26387 ;
  assign n26389 = n26383 & n26387 ;
  assign n26390 = ~\core_c_dec_accPM_E_reg/P0001  & ~n5689 ;
  assign n26391 = n26385 & n26390 ;
  assign n26392 = ~n26386 & ~n26391 ;
  assign n26393 = n26382 & n26392 ;
  assign n26394 = ~n26389 & ~n26393 ;
  assign n26395 = ~n26378 & n26394 ;
  assign n26396 = ~n26388 & n26395 ;
  assign n26397 = \sport0_txctl_TXSHT_reg[12]/P0001  & ~n19960 ;
  assign n26398 = \sport0_txctl_TX_reg[13]/P0001  & n19960 ;
  assign n26399 = ~n26397 & ~n26398 ;
  assign n26407 = ~\sice_DBR1_reg[10]/P0001  & ~\sice_DMR1_reg[10]/NET0131  ;
  assign n26408 = \core_dag_ilm2reg_PMA_pi_DO_reg[10]/NET0131  & n26407 ;
  assign n26425 = ~\core_c_psq_PMOVL_regh_DO_reg[3]/NET0131  & ~\sice_DBR1_reg[17]/P0001  ;
  assign n26426 = \core_c_psq_PMOVL_regh_DO_reg[3]/NET0131  & \sice_DBR1_reg[17]/P0001  ;
  assign n26427 = ~n26425 & ~n26426 ;
  assign n26478 = ~n26408 & ~n26427 ;
  assign n26444 = \sice_DBR1_reg[10]/P0001  & ~\sice_DMR1_reg[10]/NET0131  ;
  assign n26445 = ~\core_dag_ilm2reg_PMA_pi_DO_reg[10]/NET0131  & n26444 ;
  assign n26470 = \sice_DBR1_reg[11]/P0001  & ~\sice_DMR1_reg[11]/NET0131  ;
  assign n26471 = ~\core_dag_ilm2reg_PMA_pi_DO_reg[11]/NET0131  & n26470 ;
  assign n26479 = ~n26445 & ~n26471 ;
  assign n26480 = n26478 & n26479 ;
  assign n26409 = \core_c_psq_PMOVL_regh_DO_reg[2]/NET0131  & ~\sice_DBR1_reg[16]/P0001  ;
  assign n26410 = ~\core_c_psq_PMOVL_regh_DO_reg[2]/NET0131  & \sice_DBR1_reg[16]/P0001  ;
  assign n26411 = ~n26409 & ~n26410 ;
  assign n26412 = ~\sice_DMR1_reg[16]/NET0131  & ~n26411 ;
  assign n26405 = ~\sice_DBR1_reg[11]/P0001  & ~\sice_DMR1_reg[11]/NET0131  ;
  assign n26406 = \core_dag_ilm2reg_PMA_pi_DO_reg[11]/NET0131  & n26405 ;
  assign n26476 = ~\sice_DBR1_reg[18]/P0001  & \sice_DMR1_reg[17]/NET0131  ;
  assign n26477 = ~n26406 & n26476 ;
  assign n26481 = ~n26412 & n26477 ;
  assign n26414 = \core_dag_ilm2reg_PMA_pi_DO_reg[1]/NET0131  & \sice_DBR1_reg[1]/P0001  ;
  assign n26413 = ~\core_dag_ilm2reg_PMA_pi_DO_reg[1]/NET0131  & ~\sice_DBR1_reg[1]/P0001  ;
  assign n26415 = ~\sice_DMR1_reg[1]/NET0131  & ~n26413 ;
  assign n26416 = ~n26414 & n26415 ;
  assign n26418 = \core_dag_ilm2reg_PMA_pi_DO_reg[3]/NET0131  & \sice_DBR1_reg[3]/P0001  ;
  assign n26417 = ~\core_dag_ilm2reg_PMA_pi_DO_reg[3]/NET0131  & ~\sice_DBR1_reg[3]/P0001  ;
  assign n26419 = ~\sice_DMR1_reg[3]/NET0131  & ~n26417 ;
  assign n26420 = ~n26418 & n26419 ;
  assign n26482 = ~n26416 & ~n26420 ;
  assign n26492 = n26481 & n26482 ;
  assign n26493 = n26480 & n26492 ;
  assign n26459 = \core_dag_ilm2reg_PMA_pi_DO_reg[0]/NET0131  & \sice_DBR1_reg[0]/P0001  ;
  assign n26458 = ~\core_dag_ilm2reg_PMA_pi_DO_reg[0]/NET0131  & ~\sice_DBR1_reg[0]/P0001  ;
  assign n26460 = ~\sice_DMR1_reg[0]/NET0131  & ~n26458 ;
  assign n26461 = ~n26459 & n26460 ;
  assign n26463 = \core_dag_ilm2reg_PMA_pi_DO_reg[6]/NET0131  & \sice_DBR1_reg[6]/P0001  ;
  assign n26462 = ~\core_dag_ilm2reg_PMA_pi_DO_reg[6]/NET0131  & ~\sice_DBR1_reg[6]/P0001  ;
  assign n26464 = ~\sice_DMR1_reg[6]/NET0131  & ~n26462 ;
  assign n26465 = ~n26463 & n26464 ;
  assign n26487 = ~n26461 & ~n26465 ;
  assign n26466 = \core_dag_ilm2reg_PMA_pi_DO_reg[9]/NET0131  & ~\sice_DBR1_reg[9]/P0001  ;
  assign n26467 = ~\core_dag_ilm2reg_PMA_pi_DO_reg[9]/NET0131  & \sice_DBR1_reg[9]/P0001  ;
  assign n26468 = ~n26466 & ~n26467 ;
  assign n26469 = ~\sice_DMR1_reg[9]/NET0131  & ~n26468 ;
  assign n26473 = \core_dag_ilm2reg_PMA_pi_DO_reg[7]/NET0131  & \sice_DBR1_reg[7]/P0001  ;
  assign n26472 = ~\core_dag_ilm2reg_PMA_pi_DO_reg[7]/NET0131  & ~\sice_DBR1_reg[7]/P0001  ;
  assign n26474 = ~\sice_DMR1_reg[7]/NET0131  & ~n26472 ;
  assign n26475 = ~n26473 & n26474 ;
  assign n26488 = ~n26469 & ~n26475 ;
  assign n26489 = n26487 & n26488 ;
  assign n26441 = \core_dag_ilm2reg_PMA_pi_DO_reg[13]/NET0131  & \sice_DBR1_reg[13]/P0001  ;
  assign n26440 = ~\core_dag_ilm2reg_PMA_pi_DO_reg[13]/NET0131  & ~\sice_DBR1_reg[13]/P0001  ;
  assign n26442 = ~\sice_DMR1_reg[13]/NET0131  & ~n26440 ;
  assign n26443 = ~n26441 & n26442 ;
  assign n26446 = \core_dag_ilm2reg_PMA_pi_DO_reg[5]/NET0131  & ~\sice_DBR1_reg[5]/P0001  ;
  assign n26447 = ~\core_dag_ilm2reg_PMA_pi_DO_reg[5]/NET0131  & \sice_DBR1_reg[5]/P0001  ;
  assign n26448 = ~n26446 & ~n26447 ;
  assign n26449 = ~\sice_DMR1_reg[5]/NET0131  & ~n26448 ;
  assign n26485 = ~n26443 & ~n26449 ;
  assign n26451 = \core_dag_ilm2reg_PMA_pi_DO_reg[12]/NET0131  & \sice_DBR1_reg[12]/P0001  ;
  assign n26450 = ~\core_dag_ilm2reg_PMA_pi_DO_reg[12]/NET0131  & ~\sice_DBR1_reg[12]/P0001  ;
  assign n26452 = ~\sice_DMR1_reg[12]/NET0131  & ~n26450 ;
  assign n26453 = ~n26451 & n26452 ;
  assign n26454 = \core_dag_ilm2reg_PMA_pi_DO_reg[8]/NET0131  & ~\sice_DBR1_reg[8]/P0001  ;
  assign n26455 = ~\core_dag_ilm2reg_PMA_pi_DO_reg[8]/NET0131  & \sice_DBR1_reg[8]/P0001  ;
  assign n26456 = ~n26454 & ~n26455 ;
  assign n26457 = ~\sice_DMR1_reg[8]/NET0131  & ~n26456 ;
  assign n26486 = ~n26453 & ~n26457 ;
  assign n26490 = n26485 & n26486 ;
  assign n26422 = \core_c_psq_PMOVL_regh_DO_reg[1]/NET0131  & \sice_DBR1_reg[15]/P0001  ;
  assign n26421 = ~\core_c_psq_PMOVL_regh_DO_reg[1]/NET0131  & ~\sice_DBR1_reg[15]/P0001  ;
  assign n26423 = ~\sice_DMR1_reg[15]/NET0131  & ~n26421 ;
  assign n26424 = ~n26422 & n26423 ;
  assign n26429 = \core_dag_ilm2reg_PMA_pi_DO_reg[2]/NET0131  & \sice_DBR1_reg[2]/P0001  ;
  assign n26428 = ~\core_dag_ilm2reg_PMA_pi_DO_reg[2]/NET0131  & ~\sice_DBR1_reg[2]/P0001  ;
  assign n26430 = ~\sice_DMR1_reg[2]/NET0131  & ~n26428 ;
  assign n26431 = ~n26429 & n26430 ;
  assign n26483 = ~n26424 & ~n26431 ;
  assign n26432 = \core_c_psq_PMOVL_regh_DO_reg[0]/NET0131  & ~\sice_DBR1_reg[14]/P0001  ;
  assign n26433 = ~\core_c_psq_PMOVL_regh_DO_reg[0]/NET0131  & \sice_DBR1_reg[14]/P0001  ;
  assign n26434 = ~n26432 & ~n26433 ;
  assign n26435 = ~\sice_DMR1_reg[14]/NET0131  & ~n26434 ;
  assign n26437 = \core_dag_ilm2reg_PMA_pi_DO_reg[4]/NET0131  & \sice_DBR1_reg[4]/P0001  ;
  assign n26436 = ~\core_dag_ilm2reg_PMA_pi_DO_reg[4]/NET0131  & ~\sice_DBR1_reg[4]/P0001  ;
  assign n26438 = ~\sice_DMR1_reg[4]/NET0131  & ~n26436 ;
  assign n26439 = ~n26437 & n26438 ;
  assign n26484 = ~n26435 & ~n26439 ;
  assign n26491 = n26483 & n26484 ;
  assign n26494 = n26490 & n26491 ;
  assign n26495 = n26489 & n26494 ;
  assign n26496 = n26493 & n26495 ;
  assign n26501 = ~\sice_DBR2_reg[5]/P0001  & ~\sice_DMR2_reg[5]/NET0131  ;
  assign n26502 = \core_dag_ilm2reg_PMA_pi_DO_reg[5]/NET0131  & n26501 ;
  assign n26503 = ~\sice_DBR2_reg[10]/P0001  & ~\sice_DMR2_reg[10]/NET0131  ;
  assign n26504 = \core_dag_ilm2reg_PMA_pi_DO_reg[10]/NET0131  & n26503 ;
  assign n26570 = ~n26502 & ~n26504 ;
  assign n26545 = \sice_DBR2_reg[10]/P0001  & ~\sice_DMR2_reg[10]/NET0131  ;
  assign n26546 = ~\core_dag_ilm2reg_PMA_pi_DO_reg[10]/NET0131  & n26545 ;
  assign n26547 = \sice_DBR2_reg[5]/P0001  & ~\sice_DMR2_reg[5]/NET0131  ;
  assign n26548 = ~\core_dag_ilm2reg_PMA_pi_DO_reg[5]/NET0131  & n26547 ;
  assign n26571 = ~n26546 & ~n26548 ;
  assign n26572 = n26570 & n26571 ;
  assign n26498 = \core_dag_ilm2reg_PMA_pi_DO_reg[9]/NET0131  & \sice_DBR2_reg[9]/P0001  ;
  assign n26497 = ~\core_dag_ilm2reg_PMA_pi_DO_reg[9]/NET0131  & ~\sice_DBR2_reg[9]/P0001  ;
  assign n26499 = ~\sice_DMR2_reg[9]/NET0131  & ~n26497 ;
  assign n26500 = ~n26498 & n26499 ;
  assign n26566 = ~\core_c_psq_PMOVL_regh_DO_reg[3]/NET0131  & \sice_DBR2_reg[17]/P0001  ;
  assign n26565 = \core_c_psq_PMOVL_regh_DO_reg[3]/NET0131  & ~\sice_DBR2_reg[17]/P0001  ;
  assign n26567 = ~\sice_DBR2_reg[18]/P0001  & \sice_DMR2_reg[17]/NET0131  ;
  assign n26568 = ~n26565 & n26567 ;
  assign n26569 = ~n26566 & n26568 ;
  assign n26573 = ~n26500 & n26569 ;
  assign n26505 = \core_dag_ilm2reg_PMA_pi_DO_reg[11]/NET0131  & ~\sice_DBR2_reg[11]/P0001  ;
  assign n26506 = ~\core_dag_ilm2reg_PMA_pi_DO_reg[11]/NET0131  & \sice_DBR2_reg[11]/P0001  ;
  assign n26507 = ~n26505 & ~n26506 ;
  assign n26508 = ~\sice_DMR2_reg[11]/NET0131  & ~n26507 ;
  assign n26509 = \core_dag_ilm2reg_PMA_pi_DO_reg[4]/NET0131  & ~\sice_DBR2_reg[4]/P0001  ;
  assign n26510 = ~\core_dag_ilm2reg_PMA_pi_DO_reg[4]/NET0131  & \sice_DBR2_reg[4]/P0001  ;
  assign n26511 = ~n26509 & ~n26510 ;
  assign n26512 = ~\sice_DMR2_reg[4]/NET0131  & ~n26511 ;
  assign n26574 = ~n26508 & ~n26512 ;
  assign n26584 = n26573 & n26574 ;
  assign n26585 = n26572 & n26584 ;
  assign n26549 = \core_dag_ilm2reg_PMA_pi_DO_reg[7]/NET0131  & ~\sice_DBR2_reg[7]/P0001  ;
  assign n26550 = ~\core_dag_ilm2reg_PMA_pi_DO_reg[7]/NET0131  & \sice_DBR2_reg[7]/P0001  ;
  assign n26551 = ~n26549 & ~n26550 ;
  assign n26552 = ~\sice_DMR2_reg[7]/NET0131  & ~n26551 ;
  assign n26553 = \core_dag_ilm2reg_PMA_pi_DO_reg[2]/NET0131  & ~\sice_DBR2_reg[2]/P0001  ;
  assign n26554 = ~\core_dag_ilm2reg_PMA_pi_DO_reg[2]/NET0131  & \sice_DBR2_reg[2]/P0001  ;
  assign n26555 = ~n26553 & ~n26554 ;
  assign n26556 = ~\sice_DMR2_reg[2]/NET0131  & ~n26555 ;
  assign n26579 = ~n26552 & ~n26556 ;
  assign n26558 = \core_dag_ilm2reg_PMA_pi_DO_reg[0]/NET0131  & \sice_DBR2_reg[0]/P0001  ;
  assign n26557 = ~\core_dag_ilm2reg_PMA_pi_DO_reg[0]/NET0131  & ~\sice_DBR2_reg[0]/P0001  ;
  assign n26559 = ~\sice_DMR2_reg[0]/NET0131  & ~n26557 ;
  assign n26560 = ~n26558 & n26559 ;
  assign n26562 = \core_dag_ilm2reg_PMA_pi_DO_reg[13]/NET0131  & \sice_DBR2_reg[13]/P0001  ;
  assign n26561 = ~\core_dag_ilm2reg_PMA_pi_DO_reg[13]/NET0131  & ~\sice_DBR2_reg[13]/P0001  ;
  assign n26563 = ~\sice_DMR2_reg[13]/NET0131  & ~n26561 ;
  assign n26564 = ~n26562 & n26563 ;
  assign n26580 = ~n26560 & ~n26564 ;
  assign n26581 = n26579 & n26580 ;
  assign n26529 = \core_dag_ilm2reg_PMA_pi_DO_reg[3]/NET0131  & ~\sice_DBR2_reg[3]/P0001  ;
  assign n26530 = ~\core_dag_ilm2reg_PMA_pi_DO_reg[3]/NET0131  & \sice_DBR2_reg[3]/P0001  ;
  assign n26531 = ~n26529 & ~n26530 ;
  assign n26532 = ~\sice_DMR2_reg[3]/NET0131  & ~n26531 ;
  assign n26534 = \core_dag_ilm2reg_PMA_pi_DO_reg[12]/NET0131  & \sice_DBR2_reg[12]/P0001  ;
  assign n26533 = ~\core_dag_ilm2reg_PMA_pi_DO_reg[12]/NET0131  & ~\sice_DBR2_reg[12]/P0001  ;
  assign n26535 = ~\sice_DMR2_reg[12]/NET0131  & ~n26533 ;
  assign n26536 = ~n26534 & n26535 ;
  assign n26577 = ~n26532 & ~n26536 ;
  assign n26538 = \core_dag_ilm2reg_PMA_pi_DO_reg[1]/NET0131  & \sice_DBR2_reg[1]/P0001  ;
  assign n26537 = ~\core_dag_ilm2reg_PMA_pi_DO_reg[1]/NET0131  & ~\sice_DBR2_reg[1]/P0001  ;
  assign n26539 = ~\sice_DMR2_reg[1]/NET0131  & ~n26537 ;
  assign n26540 = ~n26538 & n26539 ;
  assign n26542 = \core_c_psq_PMOVL_regh_DO_reg[2]/NET0131  & \sice_DBR2_reg[16]/P0001  ;
  assign n26541 = ~\core_c_psq_PMOVL_regh_DO_reg[2]/NET0131  & ~\sice_DBR2_reg[16]/P0001  ;
  assign n26543 = ~\sice_DMR2_reg[16]/NET0131  & ~n26541 ;
  assign n26544 = ~n26542 & n26543 ;
  assign n26578 = ~n26540 & ~n26544 ;
  assign n26582 = n26577 & n26578 ;
  assign n26514 = \core_c_psq_PMOVL_regh_DO_reg[0]/NET0131  & \sice_DBR2_reg[14]/P0001  ;
  assign n26513 = ~\core_c_psq_PMOVL_regh_DO_reg[0]/NET0131  & ~\sice_DBR2_reg[14]/P0001  ;
  assign n26515 = ~\sice_DMR2_reg[14]/NET0131  & ~n26513 ;
  assign n26516 = ~n26514 & n26515 ;
  assign n26517 = \core_dag_ilm2reg_PMA_pi_DO_reg[8]/NET0131  & ~\sice_DBR2_reg[8]/P0001  ;
  assign n26518 = ~\core_dag_ilm2reg_PMA_pi_DO_reg[8]/NET0131  & \sice_DBR2_reg[8]/P0001  ;
  assign n26519 = ~n26517 & ~n26518 ;
  assign n26520 = ~\sice_DMR2_reg[8]/NET0131  & ~n26519 ;
  assign n26575 = ~n26516 & ~n26520 ;
  assign n26522 = \core_c_psq_PMOVL_regh_DO_reg[1]/NET0131  & \sice_DBR2_reg[15]/P0001  ;
  assign n26521 = ~\core_c_psq_PMOVL_regh_DO_reg[1]/NET0131  & ~\sice_DBR2_reg[15]/P0001  ;
  assign n26523 = ~\sice_DMR2_reg[15]/NET0131  & ~n26521 ;
  assign n26524 = ~n26522 & n26523 ;
  assign n26526 = \core_dag_ilm2reg_PMA_pi_DO_reg[6]/NET0131  & \sice_DBR2_reg[6]/P0001  ;
  assign n26525 = ~\core_dag_ilm2reg_PMA_pi_DO_reg[6]/NET0131  & ~\sice_DBR2_reg[6]/P0001  ;
  assign n26527 = ~\sice_DMR2_reg[6]/NET0131  & ~n26525 ;
  assign n26528 = ~n26526 & n26527 ;
  assign n26576 = ~n26524 & ~n26528 ;
  assign n26583 = n26575 & n26576 ;
  assign n26586 = n26582 & n26583 ;
  assign n26587 = n26581 & n26586 ;
  assign n26588 = n26585 & n26587 ;
  assign n26589 = ~n26496 & ~n26588 ;
  assign n26590 = ~\core_c_dec_Dummy_E_reg/NET0131  & \memc_accPM_E_reg/NET0131  ;
  assign n26591 = ~n26589 & n26590 ;
  assign n26592 = ~\core_dag_ilm1reg_DMA_pi_DO_reg[10]/NET0131  & n26545 ;
  assign n26593 = ~\core_dag_ilm1reg_DMA_pi_DO_reg[5]/NET0131  & n26547 ;
  assign n26663 = ~n26592 & ~n26593 ;
  assign n26645 = \core_dag_ilm1reg_DMA_pi_DO_reg[10]/NET0131  & n26503 ;
  assign n26646 = \core_dag_ilm1reg_DMA_pi_DO_reg[5]/NET0131  & n26501 ;
  assign n26664 = ~n26645 & ~n26646 ;
  assign n26665 = n26663 & n26664 ;
  assign n26594 = \core_dag_ilm1reg_DMA_pi_DO_reg[3]/NET0131  & ~\sice_DBR2_reg[3]/P0001  ;
  assign n26595 = ~\core_dag_ilm1reg_DMA_pi_DO_reg[3]/NET0131  & \sice_DBR2_reg[3]/P0001  ;
  assign n26596 = ~n26594 & ~n26595 ;
  assign n26597 = ~\sice_DMR2_reg[3]/NET0131  & ~n26596 ;
  assign n26630 = ~\core_c_psq_DMOVL_reg_DO_reg[3]/NET0131  & \sice_DBR2_reg[17]/P0001  ;
  assign n26659 = \sice_DBR2_reg[18]/P0001  & \sice_DMR2_reg[17]/NET0131  ;
  assign n26660 = ~n26630 & n26659 ;
  assign n26631 = ~\core_c_dec_Dummy_E_reg/NET0131  & \memc_accDM_E_reg/NET0131  ;
  assign n26632 = \core_c_psq_DMOVL_reg_DO_reg[3]/NET0131  & ~\sice_DBR2_reg[17]/P0001  ;
  assign n26661 = n26631 & ~n26632 ;
  assign n26662 = n26660 & n26661 ;
  assign n26666 = ~n26597 & n26662 ;
  assign n26599 = \core_dag_ilm1reg_DMA_pi_DO_reg[1]/NET0131  & \sice_DBR2_reg[1]/P0001  ;
  assign n26598 = ~\core_dag_ilm1reg_DMA_pi_DO_reg[1]/NET0131  & ~\sice_DBR2_reg[1]/P0001  ;
  assign n26600 = ~\sice_DMR2_reg[1]/NET0131  & ~n26598 ;
  assign n26601 = ~n26599 & n26600 ;
  assign n26602 = \core_dag_ilm1reg_DMA_pi_DO_reg[11]/NET0131  & ~\sice_DBR2_reg[11]/P0001  ;
  assign n26603 = ~\core_dag_ilm1reg_DMA_pi_DO_reg[11]/NET0131  & \sice_DBR2_reg[11]/P0001  ;
  assign n26604 = ~n26602 & ~n26603 ;
  assign n26605 = ~\sice_DMR2_reg[11]/NET0131  & ~n26604 ;
  assign n26667 = ~n26601 & ~n26605 ;
  assign n26677 = n26666 & n26667 ;
  assign n26678 = n26665 & n26677 ;
  assign n26642 = \core_dag_ilm1reg_DMA_pi_DO_reg[13]/NET0131  & \sice_DBR2_reg[13]/P0001  ;
  assign n26641 = ~\core_dag_ilm1reg_DMA_pi_DO_reg[13]/NET0131  & ~\sice_DBR2_reg[13]/P0001  ;
  assign n26643 = ~\sice_DMR2_reg[13]/NET0131  & ~n26641 ;
  assign n26644 = ~n26642 & n26643 ;
  assign n26647 = \core_dag_ilm1reg_DMA_pi_DO_reg[7]/NET0131  & ~\sice_DBR2_reg[7]/P0001  ;
  assign n26648 = ~\core_dag_ilm1reg_DMA_pi_DO_reg[7]/NET0131  & \sice_DBR2_reg[7]/P0001  ;
  assign n26649 = ~n26647 & ~n26648 ;
  assign n26650 = ~\sice_DMR2_reg[7]/NET0131  & ~n26649 ;
  assign n26672 = ~n26644 & ~n26650 ;
  assign n26652 = \core_dag_ilm1reg_DMA_pi_DO_reg[2]/NET0131  & \sice_DBR2_reg[2]/P0001  ;
  assign n26651 = ~\core_dag_ilm1reg_DMA_pi_DO_reg[2]/NET0131  & ~\sice_DBR2_reg[2]/P0001  ;
  assign n26653 = ~\sice_DMR2_reg[2]/NET0131  & ~n26651 ;
  assign n26654 = ~n26652 & n26653 ;
  assign n26656 = \core_dag_ilm1reg_DMA_pi_DO_reg[4]/NET0131  & \sice_DBR2_reg[4]/P0001  ;
  assign n26655 = ~\core_dag_ilm1reg_DMA_pi_DO_reg[4]/NET0131  & ~\sice_DBR2_reg[4]/P0001  ;
  assign n26657 = ~\sice_DMR2_reg[4]/NET0131  & ~n26655 ;
  assign n26658 = ~n26656 & n26657 ;
  assign n26673 = ~n26654 & ~n26658 ;
  assign n26674 = n26672 & n26673 ;
  assign n26623 = \core_dag_ilm1reg_DMA_pi_DO_reg[9]/NET0131  & \sice_DBR2_reg[9]/P0001  ;
  assign n26622 = ~\core_dag_ilm1reg_DMA_pi_DO_reg[9]/NET0131  & ~\sice_DBR2_reg[9]/P0001  ;
  assign n26624 = ~\sice_DMR2_reg[9]/NET0131  & ~n26622 ;
  assign n26625 = ~n26623 & n26624 ;
  assign n26627 = \core_dag_ilm1reg_DMA_pi_DO_reg[0]/NET0131  & \sice_DBR2_reg[0]/P0001  ;
  assign n26626 = ~\core_dag_ilm1reg_DMA_pi_DO_reg[0]/NET0131  & ~\sice_DBR2_reg[0]/P0001  ;
  assign n26628 = ~\sice_DMR2_reg[0]/NET0131  & ~n26626 ;
  assign n26629 = ~n26627 & n26628 ;
  assign n26670 = ~n26625 & ~n26629 ;
  assign n26634 = \core_c_psq_DMOVL_reg_DO_reg[1]/NET0131  & \sice_DBR2_reg[15]/P0001  ;
  assign n26633 = ~\core_c_psq_DMOVL_reg_DO_reg[1]/NET0131  & ~\sice_DBR2_reg[15]/P0001  ;
  assign n26635 = ~\sice_DMR2_reg[15]/NET0131  & ~n26633 ;
  assign n26636 = ~n26634 & n26635 ;
  assign n26637 = \core_c_psq_DMOVL_reg_DO_reg[0]/NET0131  & ~\sice_DBR2_reg[14]/P0001  ;
  assign n26638 = ~\core_c_psq_DMOVL_reg_DO_reg[0]/NET0131  & \sice_DBR2_reg[14]/P0001  ;
  assign n26639 = ~n26637 & ~n26638 ;
  assign n26640 = ~\sice_DMR2_reg[14]/NET0131  & ~n26639 ;
  assign n26671 = ~n26636 & ~n26640 ;
  assign n26675 = n26670 & n26671 ;
  assign n26607 = \core_dag_ilm1reg_DMA_pi_DO_reg[12]/NET0131  & \sice_DBR2_reg[12]/P0001  ;
  assign n26606 = ~\core_dag_ilm1reg_DMA_pi_DO_reg[12]/NET0131  & ~\sice_DBR2_reg[12]/P0001  ;
  assign n26608 = ~\sice_DMR2_reg[12]/NET0131  & ~n26606 ;
  assign n26609 = ~n26607 & n26608 ;
  assign n26611 = \core_dag_ilm1reg_DMA_pi_DO_reg[6]/NET0131  & \sice_DBR2_reg[6]/P0001  ;
  assign n26610 = ~\core_dag_ilm1reg_DMA_pi_DO_reg[6]/NET0131  & ~\sice_DBR2_reg[6]/P0001  ;
  assign n26612 = ~\sice_DMR2_reg[6]/NET0131  & ~n26610 ;
  assign n26613 = ~n26611 & n26612 ;
  assign n26668 = ~n26609 & ~n26613 ;
  assign n26615 = \core_dag_ilm1reg_DMA_pi_DO_reg[8]/NET0131  & \sice_DBR2_reg[8]/P0001  ;
  assign n26614 = ~\core_dag_ilm1reg_DMA_pi_DO_reg[8]/NET0131  & ~\sice_DBR2_reg[8]/P0001  ;
  assign n26616 = ~\sice_DMR2_reg[8]/NET0131  & ~n26614 ;
  assign n26617 = ~n26615 & n26616 ;
  assign n26618 = \core_c_psq_DMOVL_reg_DO_reg[2]/NET0131  & ~\sice_DBR2_reg[16]/P0001  ;
  assign n26619 = ~\core_c_psq_DMOVL_reg_DO_reg[2]/NET0131  & \sice_DBR2_reg[16]/P0001  ;
  assign n26620 = ~n26618 & ~n26619 ;
  assign n26621 = ~\sice_DMR2_reg[16]/NET0131  & ~n26620 ;
  assign n26669 = ~n26617 & ~n26621 ;
  assign n26676 = n26668 & n26669 ;
  assign n26679 = n26675 & n26676 ;
  assign n26680 = n26674 & n26679 ;
  assign n26681 = n26678 & n26680 ;
  assign n26683 = ~\core_dag_ilm1reg_DMA_pi_DO_reg[10]/NET0131  & n26444 ;
  assign n26704 = ~\core_dag_ilm1reg_DMA_pi_DO_reg[11]/NET0131  & n26470 ;
  assign n26752 = ~n26683 & ~n26704 ;
  assign n26717 = ~\core_c_psq_DMOVL_reg_DO_reg[3]/NET0131  & ~\sice_DBR1_reg[17]/P0001  ;
  assign n26718 = \core_c_psq_DMOVL_reg_DO_reg[3]/NET0131  & \sice_DBR1_reg[17]/P0001  ;
  assign n26719 = ~n26717 & ~n26718 ;
  assign n26744 = \core_dag_ilm1reg_DMA_pi_DO_reg[11]/NET0131  & n26405 ;
  assign n26753 = ~n26719 & ~n26744 ;
  assign n26754 = n26752 & n26753 ;
  assign n26684 = \core_dag_ilm1reg_DMA_pi_DO_reg[2]/NET0131  & ~\sice_DBR1_reg[2]/P0001  ;
  assign n26685 = ~\core_dag_ilm1reg_DMA_pi_DO_reg[2]/NET0131  & \sice_DBR1_reg[2]/P0001  ;
  assign n26686 = ~n26684 & ~n26685 ;
  assign n26687 = ~\sice_DMR1_reg[2]/NET0131  & ~n26686 ;
  assign n26682 = \core_dag_ilm1reg_DMA_pi_DO_reg[10]/NET0131  & n26407 ;
  assign n26749 = \sice_DBR1_reg[18]/P0001  & \sice_DMR1_reg[17]/NET0131  ;
  assign n26750 = n26631 & n26749 ;
  assign n26751 = ~n26682 & n26750 ;
  assign n26755 = ~n26687 & n26751 ;
  assign n26689 = \core_c_psq_DMOVL_reg_DO_reg[2]/NET0131  & \sice_DBR1_reg[16]/P0001  ;
  assign n26688 = ~\core_c_psq_DMOVL_reg_DO_reg[2]/NET0131  & ~\sice_DBR1_reg[16]/P0001  ;
  assign n26690 = ~\sice_DMR1_reg[16]/NET0131  & ~n26688 ;
  assign n26691 = ~n26689 & n26690 ;
  assign n26693 = \core_dag_ilm1reg_DMA_pi_DO_reg[5]/NET0131  & \sice_DBR1_reg[5]/P0001  ;
  assign n26692 = ~\core_dag_ilm1reg_DMA_pi_DO_reg[5]/NET0131  & ~\sice_DBR1_reg[5]/P0001  ;
  assign n26694 = ~\sice_DMR1_reg[5]/NET0131  & ~n26692 ;
  assign n26695 = ~n26693 & n26694 ;
  assign n26756 = ~n26691 & ~n26695 ;
  assign n26766 = n26755 & n26756 ;
  assign n26767 = n26754 & n26766 ;
  assign n26733 = \core_dag_ilm1reg_DMA_pi_DO_reg[8]/NET0131  & \sice_DBR1_reg[8]/P0001  ;
  assign n26732 = ~\core_dag_ilm1reg_DMA_pi_DO_reg[8]/NET0131  & ~\sice_DBR1_reg[8]/P0001  ;
  assign n26734 = ~\sice_DMR1_reg[8]/NET0131  & ~n26732 ;
  assign n26735 = ~n26733 & n26734 ;
  assign n26737 = \core_dag_ilm1reg_DMA_pi_DO_reg[4]/NET0131  & \sice_DBR1_reg[4]/P0001  ;
  assign n26736 = ~\core_dag_ilm1reg_DMA_pi_DO_reg[4]/NET0131  & ~\sice_DBR1_reg[4]/P0001  ;
  assign n26738 = ~\sice_DMR1_reg[4]/NET0131  & ~n26736 ;
  assign n26739 = ~n26737 & n26738 ;
  assign n26761 = ~n26735 & ~n26739 ;
  assign n26740 = \core_dag_ilm1reg_DMA_pi_DO_reg[6]/NET0131  & ~\sice_DBR1_reg[6]/P0001  ;
  assign n26741 = ~\core_dag_ilm1reg_DMA_pi_DO_reg[6]/NET0131  & \sice_DBR1_reg[6]/P0001  ;
  assign n26742 = ~n26740 & ~n26741 ;
  assign n26743 = ~\sice_DMR1_reg[6]/NET0131  & ~n26742 ;
  assign n26746 = \core_dag_ilm1reg_DMA_pi_DO_reg[0]/NET0131  & \sice_DBR1_reg[0]/P0001  ;
  assign n26745 = ~\core_dag_ilm1reg_DMA_pi_DO_reg[0]/NET0131  & ~\sice_DBR1_reg[0]/P0001  ;
  assign n26747 = ~\sice_DMR1_reg[0]/NET0131  & ~n26745 ;
  assign n26748 = ~n26746 & n26747 ;
  assign n26762 = ~n26743 & ~n26748 ;
  assign n26763 = n26761 & n26762 ;
  assign n26714 = \core_dag_ilm1reg_DMA_pi_DO_reg[13]/NET0131  & \sice_DBR1_reg[13]/P0001  ;
  assign n26713 = ~\core_dag_ilm1reg_DMA_pi_DO_reg[13]/NET0131  & ~\sice_DBR1_reg[13]/P0001  ;
  assign n26715 = ~\sice_DMR1_reg[13]/NET0131  & ~n26713 ;
  assign n26716 = ~n26714 & n26715 ;
  assign n26720 = \core_c_psq_DMOVL_reg_DO_reg[1]/NET0131  & ~\sice_DBR1_reg[15]/P0001  ;
  assign n26721 = ~\core_c_psq_DMOVL_reg_DO_reg[1]/NET0131  & \sice_DBR1_reg[15]/P0001  ;
  assign n26722 = ~n26720 & ~n26721 ;
  assign n26723 = ~\sice_DMR1_reg[15]/NET0131  & ~n26722 ;
  assign n26759 = ~n26716 & ~n26723 ;
  assign n26725 = \core_c_psq_DMOVL_reg_DO_reg[0]/NET0131  & \sice_DBR1_reg[14]/P0001  ;
  assign n26724 = ~\core_c_psq_DMOVL_reg_DO_reg[0]/NET0131  & ~\sice_DBR1_reg[14]/P0001  ;
  assign n26726 = ~\sice_DMR1_reg[14]/NET0131  & ~n26724 ;
  assign n26727 = ~n26725 & n26726 ;
  assign n26728 = \core_dag_ilm1reg_DMA_pi_DO_reg[3]/NET0131  & ~\sice_DBR1_reg[3]/P0001  ;
  assign n26729 = ~\core_dag_ilm1reg_DMA_pi_DO_reg[3]/NET0131  & \sice_DBR1_reg[3]/P0001  ;
  assign n26730 = ~n26728 & ~n26729 ;
  assign n26731 = ~\sice_DMR1_reg[3]/NET0131  & ~n26730 ;
  assign n26760 = ~n26727 & ~n26731 ;
  assign n26764 = n26759 & n26760 ;
  assign n26697 = \core_dag_ilm1reg_DMA_pi_DO_reg[7]/NET0131  & \sice_DBR1_reg[7]/P0001  ;
  assign n26696 = ~\core_dag_ilm1reg_DMA_pi_DO_reg[7]/NET0131  & ~\sice_DBR1_reg[7]/P0001  ;
  assign n26698 = ~\sice_DMR1_reg[7]/NET0131  & ~n26696 ;
  assign n26699 = ~n26697 & n26698 ;
  assign n26701 = \core_dag_ilm1reg_DMA_pi_DO_reg[12]/NET0131  & \sice_DBR1_reg[12]/P0001  ;
  assign n26700 = ~\core_dag_ilm1reg_DMA_pi_DO_reg[12]/NET0131  & ~\sice_DBR1_reg[12]/P0001  ;
  assign n26702 = ~\sice_DMR1_reg[12]/NET0131  & ~n26700 ;
  assign n26703 = ~n26701 & n26702 ;
  assign n26757 = ~n26699 & ~n26703 ;
  assign n26705 = \core_dag_ilm1reg_DMA_pi_DO_reg[1]/NET0131  & ~\sice_DBR1_reg[1]/P0001  ;
  assign n26706 = ~\core_dag_ilm1reg_DMA_pi_DO_reg[1]/NET0131  & \sice_DBR1_reg[1]/P0001  ;
  assign n26707 = ~n26705 & ~n26706 ;
  assign n26708 = ~\sice_DMR1_reg[1]/NET0131  & ~n26707 ;
  assign n26710 = \core_dag_ilm1reg_DMA_pi_DO_reg[9]/NET0131  & \sice_DBR1_reg[9]/P0001  ;
  assign n26709 = ~\core_dag_ilm1reg_DMA_pi_DO_reg[9]/NET0131  & ~\sice_DBR1_reg[9]/P0001  ;
  assign n26711 = ~\sice_DMR1_reg[9]/NET0131  & ~n26709 ;
  assign n26712 = ~n26710 & n26711 ;
  assign n26758 = ~n26708 & ~n26712 ;
  assign n26765 = n26757 & n26758 ;
  assign n26768 = n26764 & n26765 ;
  assign n26769 = n26763 & n26768 ;
  assign n26770 = n26767 & n26769 ;
  assign n26771 = ~n26681 & ~n26770 ;
  assign n26772 = ~n26591 & n26771 ;
  assign n26773 = \sice_ITR_reg[2]/NET0131  & ~n26772 ;
  assign n26864 = \core_c_psq_DRA_reg[6]/P0001  & ~\sice_IBR2_reg[6]/P0001  ;
  assign n26865 = ~\core_c_psq_DRA_reg[6]/P0001  & \sice_IBR2_reg[6]/P0001  ;
  assign n26866 = ~n26864 & ~n26865 ;
  assign n26867 = ~\sice_IMR2_reg[6]/NET0131  & ~n26866 ;
  assign n26933 = ~\core_c_psq_PMOVL_regl_DO_reg[3]/NET0131  & \sice_IBR2_reg[17]/P0001  ;
  assign n26932 = \core_c_psq_PMOVL_regl_DO_reg[3]/NET0131  & ~\sice_IBR2_reg[17]/P0001  ;
  assign n26934 = \sice_IMR2_reg[17]/NET0131  & \sice_ITR_reg[1]/NET0131  ;
  assign n26935 = ~n26932 & n26934 ;
  assign n26936 = ~n26933 & n26935 ;
  assign n26937 = ~n26867 & n26936 ;
  assign n26869 = \core_c_psq_DRA_reg[12]/P0001  & \sice_IBR2_reg[12]/P0001  ;
  assign n26868 = ~\core_c_psq_DRA_reg[12]/P0001  & ~\sice_IBR2_reg[12]/P0001  ;
  assign n26870 = ~\sice_IMR2_reg[12]/NET0131  & ~n26868 ;
  assign n26871 = ~n26869 & n26870 ;
  assign n26872 = \core_c_psq_DRA_reg[9]/P0001  & ~\sice_IBR2_reg[9]/P0001  ;
  assign n26873 = ~\core_c_psq_DRA_reg[9]/P0001  & \sice_IBR2_reg[9]/P0001  ;
  assign n26874 = ~n26872 & ~n26873 ;
  assign n26875 = ~\sice_IMR2_reg[9]/NET0131  & ~n26874 ;
  assign n26938 = ~n26871 & ~n26875 ;
  assign n26877 = \core_c_psq_DRA_reg[4]/P0001  & \sice_IBR2_reg[4]/P0001  ;
  assign n26876 = ~\core_c_psq_DRA_reg[4]/P0001  & ~\sice_IBR2_reg[4]/P0001  ;
  assign n26878 = ~\sice_IMR2_reg[4]/NET0131  & ~n26876 ;
  assign n26879 = ~n26877 & n26878 ;
  assign n26881 = \core_c_psq_PMOVL_regl_DO_reg[2]/NET0131  & \sice_IBR2_reg[16]/P0001  ;
  assign n26880 = ~\core_c_psq_PMOVL_regl_DO_reg[2]/NET0131  & ~\sice_IBR2_reg[16]/P0001  ;
  assign n26882 = ~\sice_IMR2_reg[16]/NET0131  & ~n26880 ;
  assign n26883 = ~n26881 & n26882 ;
  assign n26939 = ~n26879 & ~n26883 ;
  assign n26949 = n26938 & n26939 ;
  assign n26950 = n26937 & n26949 ;
  assign n26916 = \core_c_psq_DRA_reg[11]/P0001  & ~\sice_IBR2_reg[11]/P0001  ;
  assign n26917 = ~\core_c_psq_DRA_reg[11]/P0001  & \sice_IBR2_reg[11]/P0001  ;
  assign n26918 = ~n26916 & ~n26917 ;
  assign n26919 = ~\sice_IMR2_reg[11]/NET0131  & ~n26918 ;
  assign n26921 = \core_c_psq_DRA_reg[3]/P0001  & \sice_IBR2_reg[3]/P0001  ;
  assign n26920 = ~\core_c_psq_DRA_reg[3]/P0001  & ~\sice_IBR2_reg[3]/P0001  ;
  assign n26922 = ~\sice_IMR2_reg[3]/NET0131  & ~n26920 ;
  assign n26923 = ~n26921 & n26922 ;
  assign n26944 = ~n26919 & ~n26923 ;
  assign n26924 = \core_c_psq_PMOVL_regl_DO_reg[1]/NET0131  & ~\sice_IBR2_reg[15]/P0001  ;
  assign n26925 = ~\core_c_psq_PMOVL_regl_DO_reg[1]/NET0131  & \sice_IBR2_reg[15]/P0001  ;
  assign n26926 = ~n26924 & ~n26925 ;
  assign n26927 = ~\sice_IMR2_reg[15]/NET0131  & ~n26926 ;
  assign n26929 = \core_c_psq_DRA_reg[10]/P0001  & \sice_IBR2_reg[10]/P0001  ;
  assign n26928 = ~\core_c_psq_DRA_reg[10]/P0001  & ~\sice_IBR2_reg[10]/P0001  ;
  assign n26930 = ~\sice_IMR2_reg[10]/NET0131  & ~n26928 ;
  assign n26931 = ~n26929 & n26930 ;
  assign n26945 = ~n26927 & ~n26931 ;
  assign n26946 = n26944 & n26945 ;
  assign n26900 = \core_c_psq_DRA_reg[13]/P0001  & ~\sice_IBR2_reg[13]/P0001  ;
  assign n26901 = ~\core_c_psq_DRA_reg[13]/P0001  & \sice_IBR2_reg[13]/P0001  ;
  assign n26902 = ~n26900 & ~n26901 ;
  assign n26903 = ~\sice_IMR2_reg[13]/NET0131  & ~n26902 ;
  assign n26905 = \core_c_psq_DRA_reg[5]/P0001  & \sice_IBR2_reg[5]/P0001  ;
  assign n26904 = ~\core_c_psq_DRA_reg[5]/P0001  & ~\sice_IBR2_reg[5]/P0001  ;
  assign n26906 = ~\sice_IMR2_reg[5]/NET0131  & ~n26904 ;
  assign n26907 = ~n26905 & n26906 ;
  assign n26942 = ~n26903 & ~n26907 ;
  assign n26909 = \core_c_psq_PMOVL_regl_DO_reg[0]/NET0131  & \sice_IBR2_reg[14]/P0001  ;
  assign n26908 = ~\core_c_psq_PMOVL_regl_DO_reg[0]/NET0131  & ~\sice_IBR2_reg[14]/P0001  ;
  assign n26910 = ~\sice_IMR2_reg[14]/NET0131  & ~n26908 ;
  assign n26911 = ~n26909 & n26910 ;
  assign n26912 = \core_c_psq_DRA_reg[7]/P0001  & ~\sice_IBR2_reg[7]/P0001  ;
  assign n26913 = ~\core_c_psq_DRA_reg[7]/P0001  & \sice_IBR2_reg[7]/P0001  ;
  assign n26914 = ~n26912 & ~n26913 ;
  assign n26915 = ~\sice_IMR2_reg[7]/NET0131  & ~n26914 ;
  assign n26943 = ~n26911 & ~n26915 ;
  assign n26947 = n26942 & n26943 ;
  assign n26884 = \core_c_psq_DRA_reg[1]/P0001  & ~\sice_IBR2_reg[1]/P0001  ;
  assign n26885 = ~\core_c_psq_DRA_reg[1]/P0001  & \sice_IBR2_reg[1]/P0001  ;
  assign n26886 = ~n26884 & ~n26885 ;
  assign n26887 = ~\sice_IMR2_reg[1]/NET0131  & ~n26886 ;
  assign n26888 = \core_c_psq_DRA_reg[2]/P0001  & ~\sice_IBR2_reg[2]/P0001  ;
  assign n26889 = ~\core_c_psq_DRA_reg[2]/P0001  & \sice_IBR2_reg[2]/P0001  ;
  assign n26890 = ~n26888 & ~n26889 ;
  assign n26891 = ~\sice_IMR2_reg[2]/NET0131  & ~n26890 ;
  assign n26940 = ~n26887 & ~n26891 ;
  assign n26892 = \core_c_psq_DRA_reg[0]/P0001  & ~\sice_IBR2_reg[0]/P0001  ;
  assign n26893 = ~\core_c_psq_DRA_reg[0]/P0001  & \sice_IBR2_reg[0]/P0001  ;
  assign n26894 = ~n26892 & ~n26893 ;
  assign n26895 = ~\sice_IMR2_reg[0]/NET0131  & ~n26894 ;
  assign n26897 = \core_c_psq_DRA_reg[8]/P0001  & \sice_IBR2_reg[8]/P0001  ;
  assign n26896 = ~\core_c_psq_DRA_reg[8]/P0001  & ~\sice_IBR2_reg[8]/P0001  ;
  assign n26898 = ~\sice_IMR2_reg[8]/NET0131  & ~n26896 ;
  assign n26899 = ~n26897 & n26898 ;
  assign n26941 = ~n26895 & ~n26899 ;
  assign n26948 = n26940 & n26941 ;
  assign n26951 = n26947 & n26948 ;
  assign n26952 = n26946 & n26951 ;
  assign n26953 = n26950 & n26952 ;
  assign n26774 = \core_c_psq_PMOVL_regl_DO_reg[2]/NET0131  & ~\sice_IBR1_reg[16]/P0001  ;
  assign n26775 = ~\core_c_psq_PMOVL_regl_DO_reg[2]/NET0131  & \sice_IBR1_reg[16]/P0001  ;
  assign n26776 = ~n26774 & ~n26775 ;
  assign n26777 = ~\sice_IMR1_reg[16]/NET0131  & ~n26776 ;
  assign n26843 = ~\core_c_psq_PMOVL_regl_DO_reg[3]/NET0131  & \sice_IBR1_reg[17]/P0001  ;
  assign n26842 = \core_c_psq_PMOVL_regl_DO_reg[3]/NET0131  & ~\sice_IBR1_reg[17]/P0001  ;
  assign n26844 = \sice_IMR1_reg[17]/NET0131  & \sice_ITR_reg[1]/NET0131  ;
  assign n26845 = ~n26842 & n26844 ;
  assign n26846 = ~n26843 & n26845 ;
  assign n26847 = ~n26777 & n26846 ;
  assign n26778 = \core_c_psq_DRA_reg[13]/P0001  & ~\sice_IBR1_reg[13]/P0001  ;
  assign n26779 = ~\core_c_psq_DRA_reg[13]/P0001  & \sice_IBR1_reg[13]/P0001  ;
  assign n26780 = ~n26778 & ~n26779 ;
  assign n26781 = ~\sice_IMR1_reg[13]/NET0131  & ~n26780 ;
  assign n26783 = \core_c_psq_DRA_reg[6]/P0001  & \sice_IBR1_reg[6]/P0001  ;
  assign n26782 = ~\core_c_psq_DRA_reg[6]/P0001  & ~\sice_IBR1_reg[6]/P0001  ;
  assign n26784 = ~\sice_IMR1_reg[6]/NET0131  & ~n26782 ;
  assign n26785 = ~n26783 & n26784 ;
  assign n26848 = ~n26781 & ~n26785 ;
  assign n26786 = \core_c_psq_DRA_reg[12]/P0001  & ~\sice_IBR1_reg[12]/P0001  ;
  assign n26787 = ~\core_c_psq_DRA_reg[12]/P0001  & \sice_IBR1_reg[12]/P0001  ;
  assign n26788 = ~n26786 & ~n26787 ;
  assign n26789 = ~\sice_IMR1_reg[12]/NET0131  & ~n26788 ;
  assign n26791 = \core_c_psq_DRA_reg[8]/P0001  & \sice_IBR1_reg[8]/P0001  ;
  assign n26790 = ~\core_c_psq_DRA_reg[8]/P0001  & ~\sice_IBR1_reg[8]/P0001  ;
  assign n26792 = ~\sice_IMR1_reg[8]/NET0131  & ~n26790 ;
  assign n26793 = ~n26791 & n26792 ;
  assign n26849 = ~n26789 & ~n26793 ;
  assign n26859 = n26848 & n26849 ;
  assign n26860 = n26847 & n26859 ;
  assign n26826 = \core_c_psq_DRA_reg[3]/P0001  & ~\sice_IBR1_reg[3]/P0001  ;
  assign n26827 = ~\core_c_psq_DRA_reg[3]/P0001  & \sice_IBR1_reg[3]/P0001  ;
  assign n26828 = ~n26826 & ~n26827 ;
  assign n26829 = ~\sice_IMR1_reg[3]/NET0131  & ~n26828 ;
  assign n26831 = \core_c_psq_DRA_reg[0]/P0001  & \sice_IBR1_reg[0]/P0001  ;
  assign n26830 = ~\core_c_psq_DRA_reg[0]/P0001  & ~\sice_IBR1_reg[0]/P0001  ;
  assign n26832 = ~\sice_IMR1_reg[0]/NET0131  & ~n26830 ;
  assign n26833 = ~n26831 & n26832 ;
  assign n26854 = ~n26829 & ~n26833 ;
  assign n26834 = \core_c_psq_DRA_reg[9]/P0001  & ~\sice_IBR1_reg[9]/P0001  ;
  assign n26835 = ~\core_c_psq_DRA_reg[9]/P0001  & \sice_IBR1_reg[9]/P0001  ;
  assign n26836 = ~n26834 & ~n26835 ;
  assign n26837 = ~\sice_IMR1_reg[9]/NET0131  & ~n26836 ;
  assign n26839 = \core_c_psq_DRA_reg[2]/P0001  & \sice_IBR1_reg[2]/P0001  ;
  assign n26838 = ~\core_c_psq_DRA_reg[2]/P0001  & ~\sice_IBR1_reg[2]/P0001  ;
  assign n26840 = ~\sice_IMR1_reg[2]/NET0131  & ~n26838 ;
  assign n26841 = ~n26839 & n26840 ;
  assign n26855 = ~n26837 & ~n26841 ;
  assign n26856 = n26854 & n26855 ;
  assign n26811 = \core_c_psq_DRA_reg[1]/P0001  & \sice_IBR1_reg[1]/P0001  ;
  assign n26810 = ~\core_c_psq_DRA_reg[1]/P0001  & ~\sice_IBR1_reg[1]/P0001  ;
  assign n26812 = ~\sice_IMR1_reg[1]/NET0131  & ~n26810 ;
  assign n26813 = ~n26811 & n26812 ;
  assign n26815 = \core_c_psq_DRA_reg[4]/P0001  & \sice_IBR1_reg[4]/P0001  ;
  assign n26814 = ~\core_c_psq_DRA_reg[4]/P0001  & ~\sice_IBR1_reg[4]/P0001  ;
  assign n26816 = ~\sice_IMR1_reg[4]/NET0131  & ~n26814 ;
  assign n26817 = ~n26815 & n26816 ;
  assign n26852 = ~n26813 & ~n26817 ;
  assign n26819 = \core_c_psq_DRA_reg[11]/P0001  & \sice_IBR1_reg[11]/P0001  ;
  assign n26818 = ~\core_c_psq_DRA_reg[11]/P0001  & ~\sice_IBR1_reg[11]/P0001  ;
  assign n26820 = ~\sice_IMR1_reg[11]/NET0131  & ~n26818 ;
  assign n26821 = ~n26819 & n26820 ;
  assign n26822 = \core_c_psq_PMOVL_regl_DO_reg[0]/NET0131  & ~\sice_IBR1_reg[14]/P0001  ;
  assign n26823 = ~\core_c_psq_PMOVL_regl_DO_reg[0]/NET0131  & \sice_IBR1_reg[14]/P0001  ;
  assign n26824 = ~n26822 & ~n26823 ;
  assign n26825 = ~\sice_IMR1_reg[14]/NET0131  & ~n26824 ;
  assign n26853 = ~n26821 & ~n26825 ;
  assign n26857 = n26852 & n26853 ;
  assign n26795 = \core_c_psq_DRA_reg[5]/P0001  & \sice_IBR1_reg[5]/P0001  ;
  assign n26794 = ~\core_c_psq_DRA_reg[5]/P0001  & ~\sice_IBR1_reg[5]/P0001  ;
  assign n26796 = ~\sice_IMR1_reg[5]/NET0131  & ~n26794 ;
  assign n26797 = ~n26795 & n26796 ;
  assign n26798 = \core_c_psq_DRA_reg[10]/P0001  & ~\sice_IBR1_reg[10]/P0001  ;
  assign n26799 = ~\core_c_psq_DRA_reg[10]/P0001  & \sice_IBR1_reg[10]/P0001  ;
  assign n26800 = ~n26798 & ~n26799 ;
  assign n26801 = ~\sice_IMR1_reg[10]/NET0131  & ~n26800 ;
  assign n26850 = ~n26797 & ~n26801 ;
  assign n26803 = \core_c_psq_PMOVL_regl_DO_reg[1]/NET0131  & \sice_IBR1_reg[15]/P0001  ;
  assign n26802 = ~\core_c_psq_PMOVL_regl_DO_reg[1]/NET0131  & ~\sice_IBR1_reg[15]/P0001  ;
  assign n26804 = ~\sice_IMR1_reg[15]/NET0131  & ~n26802 ;
  assign n26805 = ~n26803 & n26804 ;
  assign n26806 = \core_c_psq_DRA_reg[7]/P0001  & ~\sice_IBR1_reg[7]/P0001  ;
  assign n26807 = ~\core_c_psq_DRA_reg[7]/P0001  & \sice_IBR1_reg[7]/P0001  ;
  assign n26808 = ~n26806 & ~n26807 ;
  assign n26809 = ~\sice_IMR1_reg[7]/NET0131  & ~n26808 ;
  assign n26851 = ~n26805 & ~n26809 ;
  assign n26858 = n26850 & n26851 ;
  assign n26861 = n26857 & n26858 ;
  assign n26862 = n26856 & n26861 ;
  assign n26863 = n26860 & n26862 ;
  assign n26400 = ~\core_c_psq_PCS_reg[0]/NET0131  & ~\core_c_psq_PCS_reg[15]/NET0131  ;
  assign n26401 = ~\core_c_psq_PCS_reg[1]/NET0131  & \sice_GOICE_syn_reg/P0001  ;
  assign n26402 = n26400 & n26401 ;
  assign n26403 = \core_c_dec_IR_reg[4]/NET0131  & \sice_ITR_reg[0]/NET0131  ;
  assign n26404 = n23230 & n26403 ;
  assign n26954 = ~n26402 & ~n26404 ;
  assign n26955 = ~n26863 & n26954 ;
  assign n26956 = ~n26953 & n26955 ;
  assign n26957 = ~n26773 & n26956 ;
  assign n26958 = ~n4093 & ~n26957 ;
  assign n26959 = n11741 & n26958 ;
  assign n26960 = ~\sice_HALT_E_reg/P0001  & ~n26959 ;
  assign n26961 = n12234 & n23717 ;
  assign n26962 = ~n26960 & n26961 ;
  assign n26964 = n26388 & ~n26391 ;
  assign n26963 = n26377 & n26390 ;
  assign n26965 = ~n26389 & ~n26963 ;
  assign n26966 = ~n26964 & n26965 ;
  assign n26967 = \sice_UpdDR_sd1_reg/P0001  & ~\sice_UpdDR_sd2_reg/P0001  ;
  assign n26968 = n23408 & n25033 ;
  assign n26969 = n26967 & n26968 ;
  assign n26970 = ~\core_c_dec_Dummy_E_reg/NET0131  & \core_c_dec_MTIDR_E_reg/P0001  ;
  assign n26971 = ~\core_c_dec_rdCM_E_reg/NET0131  & ~n26970 ;
  assign n26972 = ~n5950 & ~n26971 ;
  assign n26973 = ~n26969 & ~n26972 ;
  assign n26975 = n12743 & n26970 ;
  assign n26976 = \T_TMODE[1]_pad  & \emc_ECMDreg_reg[15]/P0001  ;
  assign n26977 = ~\idma_CMo_oe3_reg/P0001  & ~\idma_CMo_oe4_reg/P0001  ;
  assign n26978 = ~\idma_CMo_oe5_reg/P0001  & n26977 ;
  assign n26979 = ~\idma_CMo_oe6_reg/P0001  & n26978 ;
  assign n26986 = ~\idma_CMo_oe1_reg/P0001  & ~\idma_CMo_oe2_reg/P0001  ;
  assign n26991 = n26979 & n26986 ;
  assign n26992 = ~\idma_CM_oe_reg/P0001  & \idma_CMo_oe0_reg/P0001  ;
  assign n26993 = ~\idma_CMo_oe7_reg/P0001  & n26992 ;
  assign n26994 = n26991 & n26993 ;
  assign n26980 = ~\idma_CM_oe_reg/P0001  & ~\idma_CMo_oe0_reg/P0001  ;
  assign n26996 = \idma_CMo_oe7_reg/P0001  & n26980 ;
  assign n26997 = n26991 & n26996 ;
  assign n27013 = ~n26994 & ~n26997 ;
  assign n26981 = ~\idma_CMo_oe7_reg/P0001  & n26980 ;
  assign n26982 = n26979 & n26981 ;
  assign n26999 = ~\idma_CMo_oe1_reg/P0001  & \idma_CMo_oe2_reg/P0001  ;
  assign n27000 = n26982 & n26999 ;
  assign n26987 = n26981 & n26986 ;
  assign n27002 = ~\idma_CMo_oe6_reg/P0001  & n26987 ;
  assign n27003 = \idma_CMo_oe5_reg/P0001  & n26977 ;
  assign n27004 = n27002 & n27003 ;
  assign n27014 = ~n27000 & ~n27004 ;
  assign n27015 = n27013 & n27014 ;
  assign n27006 = ~\idma_CMo_oe5_reg/P0001  & n27002 ;
  assign n27010 = \idma_CMo_oe3_reg/P0001  & ~\idma_CMo_oe4_reg/P0001  ;
  assign n27011 = n27006 & n27010 ;
  assign n27007 = ~\idma_CMo_oe3_reg/P0001  & \idma_CMo_oe4_reg/P0001  ;
  assign n27008 = n27006 & n27007 ;
  assign n26983 = \idma_CMo_oe1_reg/P0001  & ~\idma_CMo_oe2_reg/P0001  ;
  assign n26984 = n26982 & n26983 ;
  assign n26988 = \idma_CMo_oe6_reg/P0001  & n26978 ;
  assign n26989 = n26987 & n26988 ;
  assign n27012 = ~n26984 & ~n26989 ;
  assign n27016 = ~n27008 & n27012 ;
  assign n27017 = ~n27011 & n27016 ;
  assign n27018 = n27015 & n27017 ;
  assign n27019 = \CM_rdm[15]_pad  & n27018 ;
  assign n26995 = \CM_rd0[15]_pad  & n26994 ;
  assign n26998 = \CM_rd7[15]_pad  & n26997 ;
  assign n27022 = ~n26995 & ~n26998 ;
  assign n27001 = \CM_rd2[15]_pad  & n27000 ;
  assign n27005 = \CM_rd5[15]_pad  & n27004 ;
  assign n27023 = ~n27001 & ~n27005 ;
  assign n27024 = n27022 & n27023 ;
  assign n27020 = \CM_rd3[15]_pad  & n27011 ;
  assign n27009 = \CM_rd4[15]_pad  & n27008 ;
  assign n26985 = \CM_rd1[15]_pad  & n26984 ;
  assign n26990 = \CM_rd6[15]_pad  & n26989 ;
  assign n27021 = ~n26985 & ~n26990 ;
  assign n27025 = ~n27009 & n27021 ;
  assign n27026 = ~n27020 & n27025 ;
  assign n27027 = n27024 & n27026 ;
  assign n27028 = ~n27019 & n27027 ;
  assign n27029 = ~\T_TMODE[1]_pad  & ~n27028 ;
  assign n27030 = ~n26976 & ~n27029 ;
  assign n27031 = \core_c_dec_rdCM_E_reg/NET0131  & ~n27030 ;
  assign n27032 = ~n26975 & ~n27031 ;
  assign n27033 = ~n26973 & ~n27032 ;
  assign n26974 = \sice_idr1_reg_DO_reg[3]/P0001  & n26973 ;
  assign n27034 = \sice_SPC_reg[15]/P0001  & n26969 ;
  assign n27035 = ~n26974 & ~n27034 ;
  assign n27036 = ~n27033 & n27035 ;
  assign n27038 = ~n18974 & n19499 ;
  assign n27037 = ~\core_eu_em_mac_em_reg_mr1swe_DO_reg[1]/P0001  & ~n19499 ;
  assign n27039 = n19501 & ~n27037 ;
  assign n27040 = ~n27038 & n27039 ;
  assign n27041 = \core_eu_em_mac_em_reg_mr1swe_DO_reg[1]/P0001  & ~n19383 ;
  assign n27042 = ~n19508 & ~n27041 ;
  assign n27043 = ~n27040 & n27042 ;
  assign n27044 = ~n18262 & ~n27043 ;
  assign n27045 = ~\core_c_psq_MSTAT_reg_DO_reg[4]/NET0131  & n19577 ;
  assign n27046 = ~n17638 & ~n17665 ;
  assign n27047 = ~n16363 & n17661 ;
  assign n27048 = ~n17670 & ~n27047 ;
  assign n27049 = ~n27046 & n27048 ;
  assign n27050 = n27046 & ~n27048 ;
  assign n27051 = ~n27049 & ~n27050 ;
  assign n27052 = \core_c_psq_MSTAT_reg_DO_reg[4]/NET0131  & n27051 ;
  assign n27053 = ~n27045 & ~n27052 ;
  assign n27054 = n18262 & ~n27053 ;
  assign n27055 = ~n27044 & ~n27054 ;
  assign n27057 = n12688 & n26970 ;
  assign n27058 = \T_TMODE[1]_pad  & \emc_ECMDreg_reg[14]/P0001  ;
  assign n27066 = \CM_rdm[14]_pad  & n27018 ;
  assign n27061 = \CM_rd0[14]_pad  & n26994 ;
  assign n27062 = \CM_rd7[14]_pad  & n26997 ;
  assign n27069 = ~n27061 & ~n27062 ;
  assign n27063 = \CM_rd2[14]_pad  & n27000 ;
  assign n27064 = \CM_rd5[14]_pad  & n27004 ;
  assign n27070 = ~n27063 & ~n27064 ;
  assign n27071 = n27069 & n27070 ;
  assign n27067 = \CM_rd3[14]_pad  & n27011 ;
  assign n27065 = \CM_rd4[14]_pad  & n27008 ;
  assign n27059 = \CM_rd1[14]_pad  & n26984 ;
  assign n27060 = \CM_rd6[14]_pad  & n26989 ;
  assign n27068 = ~n27059 & ~n27060 ;
  assign n27072 = ~n27065 & n27068 ;
  assign n27073 = ~n27067 & n27072 ;
  assign n27074 = n27071 & n27073 ;
  assign n27075 = ~n27066 & n27074 ;
  assign n27076 = ~\T_TMODE[1]_pad  & ~n27075 ;
  assign n27077 = ~n27058 & ~n27076 ;
  assign n27078 = \core_c_dec_rdCM_E_reg/NET0131  & ~n27077 ;
  assign n27079 = ~n27057 & ~n27078 ;
  assign n27080 = ~n26973 & ~n27079 ;
  assign n27056 = \sice_idr1_reg_DO_reg[2]/P0001  & n26973 ;
  assign n27081 = \sice_SPC_reg[14]/P0001  & n26969 ;
  assign n27082 = ~n27056 & ~n27081 ;
  assign n27083 = ~n27080 & n27082 ;
  assign n27085 = n11265 & n26970 ;
  assign n27086 = \T_TMODE[1]_pad  & \emc_ECMDreg_reg[7]/P0001  ;
  assign n27094 = \CM_rdm[7]_pad  & n27018 ;
  assign n27089 = \CM_rd0[7]_pad  & n26994 ;
  assign n27090 = \CM_rd7[7]_pad  & n26997 ;
  assign n27097 = ~n27089 & ~n27090 ;
  assign n27091 = \CM_rd2[7]_pad  & n27000 ;
  assign n27092 = \CM_rd5[7]_pad  & n27004 ;
  assign n27098 = ~n27091 & ~n27092 ;
  assign n27099 = n27097 & n27098 ;
  assign n27095 = \CM_rd3[7]_pad  & n27011 ;
  assign n27093 = \CM_rd4[7]_pad  & n27008 ;
  assign n27087 = \CM_rd1[7]_pad  & n26984 ;
  assign n27088 = \CM_rd6[7]_pad  & n26989 ;
  assign n27096 = ~n27087 & ~n27088 ;
  assign n27100 = ~n27093 & n27096 ;
  assign n27101 = ~n27095 & n27100 ;
  assign n27102 = n27099 & n27101 ;
  assign n27103 = ~n27094 & n27102 ;
  assign n27104 = ~\T_TMODE[1]_pad  & ~n27103 ;
  assign n27105 = ~n27086 & ~n27104 ;
  assign n27106 = \core_c_dec_rdCM_E_reg/NET0131  & ~n27105 ;
  assign n27107 = ~n27085 & ~n27106 ;
  assign n27108 = ~n26973 & ~n27107 ;
  assign n27084 = \sice_idr0_reg_DO_reg[7]/P0001  & n26973 ;
  assign n27109 = \sice_SPC_reg[7]/P0001  & n26969 ;
  assign n27110 = ~n27084 & ~n27109 ;
  assign n27111 = ~n27108 & n27110 ;
  assign n27113 = n11525 & n26970 ;
  assign n27114 = \T_TMODE[1]_pad  & \emc_ECMDreg_reg[6]/P0001  ;
  assign n27122 = \CM_rdm[6]_pad  & n27018 ;
  assign n27117 = \CM_rd0[6]_pad  & n26994 ;
  assign n27118 = \CM_rd7[6]_pad  & n26997 ;
  assign n27125 = ~n27117 & ~n27118 ;
  assign n27119 = \CM_rd2[6]_pad  & n27000 ;
  assign n27120 = \CM_rd5[6]_pad  & n27004 ;
  assign n27126 = ~n27119 & ~n27120 ;
  assign n27127 = n27125 & n27126 ;
  assign n27123 = \CM_rd3[6]_pad  & n27011 ;
  assign n27121 = \CM_rd4[6]_pad  & n27008 ;
  assign n27115 = \CM_rd1[6]_pad  & n26984 ;
  assign n27116 = \CM_rd6[6]_pad  & n26989 ;
  assign n27124 = ~n27115 & ~n27116 ;
  assign n27128 = ~n27121 & n27124 ;
  assign n27129 = ~n27123 & n27128 ;
  assign n27130 = n27127 & n27129 ;
  assign n27131 = ~n27122 & n27130 ;
  assign n27132 = ~\T_TMODE[1]_pad  & ~n27131 ;
  assign n27133 = ~n27114 & ~n27132 ;
  assign n27134 = \core_c_dec_rdCM_E_reg/NET0131  & ~n27133 ;
  assign n27135 = ~n27113 & ~n27134 ;
  assign n27136 = ~n26973 & ~n27135 ;
  assign n27112 = \sice_idr0_reg_DO_reg[6]/P0001  & n26973 ;
  assign n27137 = \sice_SPC_reg[6]/P0001  & n26969 ;
  assign n27138 = ~n27112 & ~n27137 ;
  assign n27139 = ~n27136 & n27138 ;
  assign n27141 = n10911 & n26970 ;
  assign n27142 = \T_TMODE[1]_pad  & \emc_ECMDreg_reg[5]/P0001  ;
  assign n27150 = \CM_rdm[5]_pad  & n27018 ;
  assign n27145 = \CM_rd0[5]_pad  & n26994 ;
  assign n27146 = \CM_rd7[5]_pad  & n26997 ;
  assign n27153 = ~n27145 & ~n27146 ;
  assign n27147 = \CM_rd2[5]_pad  & n27000 ;
  assign n27148 = \CM_rd5[5]_pad  & n27004 ;
  assign n27154 = ~n27147 & ~n27148 ;
  assign n27155 = n27153 & n27154 ;
  assign n27151 = \CM_rd3[5]_pad  & n27011 ;
  assign n27149 = \CM_rd4[5]_pad  & n27008 ;
  assign n27143 = \CM_rd1[5]_pad  & n26984 ;
  assign n27144 = \CM_rd6[5]_pad  & n26989 ;
  assign n27152 = ~n27143 & ~n27144 ;
  assign n27156 = ~n27149 & n27152 ;
  assign n27157 = ~n27151 & n27156 ;
  assign n27158 = n27155 & n27157 ;
  assign n27159 = ~n27150 & n27158 ;
  assign n27160 = ~\T_TMODE[1]_pad  & ~n27159 ;
  assign n27161 = ~n27142 & ~n27160 ;
  assign n27162 = \core_c_dec_rdCM_E_reg/NET0131  & ~n27161 ;
  assign n27163 = ~n27141 & ~n27162 ;
  assign n27164 = ~n26973 & ~n27163 ;
  assign n27140 = \sice_idr0_reg_DO_reg[5]/P0001  & n26973 ;
  assign n27165 = \sice_SPC_reg[5]/P0001  & n26969 ;
  assign n27166 = ~n27140 & ~n27165 ;
  assign n27167 = ~n27164 & n27166 ;
  assign n27169 = n10069 & n26970 ;
  assign n27170 = \T_TMODE[1]_pad  & \emc_ECMDreg_reg[4]/P0001  ;
  assign n27178 = \CM_rdm[4]_pad  & n27018 ;
  assign n27173 = \CM_rd0[4]_pad  & n26994 ;
  assign n27174 = \CM_rd7[4]_pad  & n26997 ;
  assign n27181 = ~n27173 & ~n27174 ;
  assign n27175 = \CM_rd2[4]_pad  & n27000 ;
  assign n27176 = \CM_rd5[4]_pad  & n27004 ;
  assign n27182 = ~n27175 & ~n27176 ;
  assign n27183 = n27181 & n27182 ;
  assign n27179 = \CM_rd3[4]_pad  & n27011 ;
  assign n27177 = \CM_rd4[4]_pad  & n27008 ;
  assign n27171 = \CM_rd1[4]_pad  & n26984 ;
  assign n27172 = \CM_rd6[4]_pad  & n26989 ;
  assign n27180 = ~n27171 & ~n27172 ;
  assign n27184 = ~n27177 & n27180 ;
  assign n27185 = ~n27179 & n27184 ;
  assign n27186 = n27183 & n27185 ;
  assign n27187 = ~n27178 & n27186 ;
  assign n27188 = ~\T_TMODE[1]_pad  & ~n27187 ;
  assign n27189 = ~n27170 & ~n27188 ;
  assign n27190 = \core_c_dec_rdCM_E_reg/NET0131  & ~n27189 ;
  assign n27191 = ~n27169 & ~n27190 ;
  assign n27192 = ~n26973 & ~n27191 ;
  assign n27168 = \sice_idr0_reg_DO_reg[4]/P0001  & n26973 ;
  assign n27193 = \sice_SPC_reg[4]/P0001  & n26969 ;
  assign n27194 = ~n27168 & ~n27193 ;
  assign n27195 = ~n27192 & n27194 ;
  assign n27197 = n8113 & n26970 ;
  assign n27198 = \T_TMODE[1]_pad  & \emc_ECMDreg_reg[3]/P0001  ;
  assign n27206 = \CM_rdm[3]_pad  & n27018 ;
  assign n27201 = \CM_rd0[3]_pad  & n26994 ;
  assign n27202 = \CM_rd7[3]_pad  & n26997 ;
  assign n27209 = ~n27201 & ~n27202 ;
  assign n27203 = \CM_rd2[3]_pad  & n27000 ;
  assign n27204 = \CM_rd5[3]_pad  & n27004 ;
  assign n27210 = ~n27203 & ~n27204 ;
  assign n27211 = n27209 & n27210 ;
  assign n27207 = \CM_rd3[3]_pad  & n27011 ;
  assign n27205 = \CM_rd4[3]_pad  & n27008 ;
  assign n27199 = \CM_rd1[3]_pad  & n26984 ;
  assign n27200 = \CM_rd6[3]_pad  & n26989 ;
  assign n27208 = ~n27199 & ~n27200 ;
  assign n27212 = ~n27205 & n27208 ;
  assign n27213 = ~n27207 & n27212 ;
  assign n27214 = n27211 & n27213 ;
  assign n27215 = ~n27206 & n27214 ;
  assign n27216 = ~\T_TMODE[1]_pad  & ~n27215 ;
  assign n27217 = ~n27198 & ~n27216 ;
  assign n27218 = \core_c_dec_rdCM_E_reg/NET0131  & ~n27217 ;
  assign n27219 = ~n27197 & ~n27218 ;
  assign n27220 = ~n26973 & ~n27219 ;
  assign n27196 = \sice_idr0_reg_DO_reg[3]/P0001  & n26973 ;
  assign n27221 = \sice_SPC_reg[3]/P0001  & n26969 ;
  assign n27222 = ~n27196 & ~n27221 ;
  assign n27223 = ~n27220 & n27222 ;
  assign n27225 = n8715 & n26970 ;
  assign n27226 = \T_TMODE[1]_pad  & \emc_ECMDreg_reg[2]/P0001  ;
  assign n27234 = \CM_rdm[2]_pad  & n27018 ;
  assign n27229 = \CM_rd0[2]_pad  & n26994 ;
  assign n27230 = \CM_rd7[2]_pad  & n26997 ;
  assign n27237 = ~n27229 & ~n27230 ;
  assign n27231 = \CM_rd2[2]_pad  & n27000 ;
  assign n27232 = \CM_rd5[2]_pad  & n27004 ;
  assign n27238 = ~n27231 & ~n27232 ;
  assign n27239 = n27237 & n27238 ;
  assign n27235 = \CM_rd3[2]_pad  & n27011 ;
  assign n27233 = \CM_rd4[2]_pad  & n27008 ;
  assign n27227 = \CM_rd1[2]_pad  & n26984 ;
  assign n27228 = \CM_rd6[2]_pad  & n26989 ;
  assign n27236 = ~n27227 & ~n27228 ;
  assign n27240 = ~n27233 & n27236 ;
  assign n27241 = ~n27235 & n27240 ;
  assign n27242 = n27239 & n27241 ;
  assign n27243 = ~n27234 & n27242 ;
  assign n27244 = ~\T_TMODE[1]_pad  & ~n27243 ;
  assign n27245 = ~n27226 & ~n27244 ;
  assign n27246 = \core_c_dec_rdCM_E_reg/NET0131  & ~n27245 ;
  assign n27247 = ~n27225 & ~n27246 ;
  assign n27248 = ~n26973 & ~n27247 ;
  assign n27224 = \sice_idr0_reg_DO_reg[2]/P0001  & n26973 ;
  assign n27249 = \sice_SPC_reg[2]/P0001  & n26969 ;
  assign n27250 = ~n27224 & ~n27249 ;
  assign n27251 = ~n27248 & n27250 ;
  assign n27253 = n9435 & n26970 ;
  assign n27254 = \T_TMODE[1]_pad  & \emc_ECMDreg_reg[1]/P0001  ;
  assign n27262 = \CM_rdm[1]_pad  & n27018 ;
  assign n27257 = \CM_rd0[1]_pad  & n26994 ;
  assign n27258 = \CM_rd7[1]_pad  & n26997 ;
  assign n27265 = ~n27257 & ~n27258 ;
  assign n27259 = \CM_rd2[1]_pad  & n27000 ;
  assign n27260 = \CM_rd5[1]_pad  & n27004 ;
  assign n27266 = ~n27259 & ~n27260 ;
  assign n27267 = n27265 & n27266 ;
  assign n27263 = \CM_rd3[1]_pad  & n27011 ;
  assign n27261 = \CM_rd4[1]_pad  & n27008 ;
  assign n27255 = \CM_rd1[1]_pad  & n26984 ;
  assign n27256 = \CM_rd6[1]_pad  & n26989 ;
  assign n27264 = ~n27255 & ~n27256 ;
  assign n27268 = ~n27261 & n27264 ;
  assign n27269 = ~n27263 & n27268 ;
  assign n27270 = n27267 & n27269 ;
  assign n27271 = ~n27262 & n27270 ;
  assign n27272 = ~\T_TMODE[1]_pad  & ~n27271 ;
  assign n27273 = ~n27254 & ~n27272 ;
  assign n27274 = \core_c_dec_rdCM_E_reg/NET0131  & ~n27273 ;
  assign n27275 = ~n27253 & ~n27274 ;
  assign n27276 = ~n26973 & ~n27275 ;
  assign n27252 = \sice_idr0_reg_DO_reg[1]/P0001  & n26973 ;
  assign n27277 = \sice_SPC_reg[1]/P0001  & n26969 ;
  assign n27278 = ~n27252 & ~n27277 ;
  assign n27279 = ~n27276 & n27278 ;
  assign n27281 = n7607 & n26970 ;
  assign n27282 = \T_TMODE[1]_pad  & \emc_ECMDreg_reg[0]/P0001  ;
  assign n27290 = \CM_rdm[0]_pad  & n27018 ;
  assign n27285 = \CM_rd0[0]_pad  & n26994 ;
  assign n27286 = \CM_rd7[0]_pad  & n26997 ;
  assign n27293 = ~n27285 & ~n27286 ;
  assign n27287 = \CM_rd2[0]_pad  & n27000 ;
  assign n27288 = \CM_rd5[0]_pad  & n27004 ;
  assign n27294 = ~n27287 & ~n27288 ;
  assign n27295 = n27293 & n27294 ;
  assign n27291 = \CM_rd3[0]_pad  & n27011 ;
  assign n27289 = \CM_rd4[0]_pad  & n27008 ;
  assign n27283 = \CM_rd1[0]_pad  & n26984 ;
  assign n27284 = \CM_rd6[0]_pad  & n26989 ;
  assign n27292 = ~n27283 & ~n27284 ;
  assign n27296 = ~n27289 & n27292 ;
  assign n27297 = ~n27291 & n27296 ;
  assign n27298 = n27295 & n27297 ;
  assign n27299 = ~n27290 & n27298 ;
  assign n27300 = ~\T_TMODE[1]_pad  & ~n27299 ;
  assign n27301 = ~n27282 & ~n27300 ;
  assign n27302 = \core_c_dec_rdCM_E_reg/NET0131  & ~n27301 ;
  assign n27303 = ~n27281 & ~n27302 ;
  assign n27304 = ~n26973 & ~n27303 ;
  assign n27280 = \sice_idr0_reg_DO_reg[0]/P0001  & n26973 ;
  assign n27305 = \sice_SPC_reg[0]/P0001  & n26969 ;
  assign n27306 = ~n27280 & ~n27305 ;
  assign n27307 = ~n27304 & n27306 ;
  assign n27308 = n14752 & n27053 ;
  assign n27309 = n18974 & n19776 ;
  assign n27310 = \core_eu_em_mac_em_reg_mr1rwe_DO_reg[1]/P0001  & ~n17809 ;
  assign n27311 = n19780 & ~n27310 ;
  assign n27312 = ~n27309 & n27311 ;
  assign n27313 = ~n27308 & ~n27312 ;
  assign n27315 = n7340 & n26970 ;
  assign n27316 = \T_TMODE[1]_pad  & \emc_ECMDreg_reg[13]/P0001  ;
  assign n27324 = \CM_rdm[13]_pad  & n27018 ;
  assign n27319 = \CM_rd0[13]_pad  & n26994 ;
  assign n27320 = \CM_rd7[13]_pad  & n26997 ;
  assign n27327 = ~n27319 & ~n27320 ;
  assign n27321 = \CM_rd2[13]_pad  & n27000 ;
  assign n27322 = \CM_rd5[13]_pad  & n27004 ;
  assign n27328 = ~n27321 & ~n27322 ;
  assign n27329 = n27327 & n27328 ;
  assign n27325 = \CM_rd3[13]_pad  & n27011 ;
  assign n27323 = \CM_rd4[13]_pad  & n27008 ;
  assign n27317 = \CM_rd1[13]_pad  & n26984 ;
  assign n27318 = \CM_rd6[13]_pad  & n26989 ;
  assign n27326 = ~n27317 & ~n27318 ;
  assign n27330 = ~n27323 & n27326 ;
  assign n27331 = ~n27325 & n27330 ;
  assign n27332 = n27329 & n27331 ;
  assign n27333 = ~n27324 & n27332 ;
  assign n27334 = ~\T_TMODE[1]_pad  & ~n27333 ;
  assign n27335 = ~n27316 & ~n27334 ;
  assign n27336 = \core_c_dec_rdCM_E_reg/NET0131  & ~n27335 ;
  assign n27337 = ~n27315 & ~n27336 ;
  assign n27338 = ~n26973 & ~n27337 ;
  assign n27314 = \sice_idr1_reg_DO_reg[1]/P0001  & n26973 ;
  assign n27339 = \sice_SPC_reg[13]/P0001  & n26969 ;
  assign n27340 = ~n27314 & ~n27339 ;
  assign n27341 = ~n27338 & n27340 ;
  assign n27343 = n9178 & n26970 ;
  assign n27344 = \T_TMODE[1]_pad  & \emc_ECMDreg_reg[12]/P0001  ;
  assign n27352 = \CM_rdm[12]_pad  & n27018 ;
  assign n27347 = \CM_rd0[12]_pad  & n26994 ;
  assign n27348 = \CM_rd7[12]_pad  & n26997 ;
  assign n27355 = ~n27347 & ~n27348 ;
  assign n27349 = \CM_rd2[12]_pad  & n27000 ;
  assign n27350 = \CM_rd5[12]_pad  & n27004 ;
  assign n27356 = ~n27349 & ~n27350 ;
  assign n27357 = n27355 & n27356 ;
  assign n27353 = \CM_rd3[12]_pad  & n27011 ;
  assign n27351 = \CM_rd4[12]_pad  & n27008 ;
  assign n27345 = \CM_rd1[12]_pad  & n26984 ;
  assign n27346 = \CM_rd6[12]_pad  & n26989 ;
  assign n27354 = ~n27345 & ~n27346 ;
  assign n27358 = ~n27351 & n27354 ;
  assign n27359 = ~n27353 & n27358 ;
  assign n27360 = n27357 & n27359 ;
  assign n27361 = ~n27352 & n27360 ;
  assign n27362 = ~\T_TMODE[1]_pad  & ~n27361 ;
  assign n27363 = ~n27344 & ~n27362 ;
  assign n27364 = \core_c_dec_rdCM_E_reg/NET0131  & ~n27363 ;
  assign n27365 = ~n27343 & ~n27364 ;
  assign n27366 = ~n26973 & ~n27365 ;
  assign n27342 = \sice_idr1_reg_DO_reg[0]/P0001  & n26973 ;
  assign n27367 = \sice_SPC_reg[12]/P0001  & n26969 ;
  assign n27368 = ~n27342 & ~n27367 ;
  assign n27369 = ~n27366 & n27368 ;
  assign n27371 = n10638 & n26970 ;
  assign n27372 = \T_TMODE[1]_pad  & \emc_ECMDreg_reg[8]/P0001  ;
  assign n27380 = \CM_rdm[8]_pad  & n27018 ;
  assign n27375 = \CM_rd0[8]_pad  & n26994 ;
  assign n27376 = \CM_rd7[8]_pad  & n26997 ;
  assign n27383 = ~n27375 & ~n27376 ;
  assign n27377 = \CM_rd2[8]_pad  & n27000 ;
  assign n27378 = \CM_rd5[8]_pad  & n27004 ;
  assign n27384 = ~n27377 & ~n27378 ;
  assign n27385 = n27383 & n27384 ;
  assign n27381 = \CM_rd3[8]_pad  & n27011 ;
  assign n27379 = \CM_rd4[8]_pad  & n27008 ;
  assign n27373 = \CM_rd1[8]_pad  & n26984 ;
  assign n27374 = \CM_rd6[8]_pad  & n26989 ;
  assign n27382 = ~n27373 & ~n27374 ;
  assign n27386 = ~n27379 & n27382 ;
  assign n27387 = ~n27381 & n27386 ;
  assign n27388 = n27385 & n27387 ;
  assign n27389 = ~n27380 & n27388 ;
  assign n27390 = ~\T_TMODE[1]_pad  & ~n27389 ;
  assign n27391 = ~n27372 & ~n27390 ;
  assign n27392 = \core_c_dec_rdCM_E_reg/NET0131  & ~n27391 ;
  assign n27393 = ~n27371 & ~n27392 ;
  assign n27394 = ~n26973 & ~n27393 ;
  assign n27370 = \sice_idr0_reg_DO_reg[8]/P0001  & n26973 ;
  assign n27395 = \sice_SPC_reg[8]/P0001  & n26969 ;
  assign n27396 = ~n27370 & ~n27395 ;
  assign n27397 = ~n27394 & n27396 ;
  assign n27399 = n10289 & n26970 ;
  assign n27400 = \T_TMODE[1]_pad  & \emc_ECMDreg_reg[9]/P0001  ;
  assign n27408 = \CM_rdm[9]_pad  & n27018 ;
  assign n27403 = \CM_rd0[9]_pad  & n26994 ;
  assign n27404 = \CM_rd7[9]_pad  & n26997 ;
  assign n27411 = ~n27403 & ~n27404 ;
  assign n27405 = \CM_rd2[9]_pad  & n27000 ;
  assign n27406 = \CM_rd5[9]_pad  & n27004 ;
  assign n27412 = ~n27405 & ~n27406 ;
  assign n27413 = n27411 & n27412 ;
  assign n27409 = \CM_rd3[9]_pad  & n27011 ;
  assign n27407 = \CM_rd4[9]_pad  & n27008 ;
  assign n27401 = \CM_rd1[9]_pad  & n26984 ;
  assign n27402 = \CM_rd6[9]_pad  & n26989 ;
  assign n27410 = ~n27401 & ~n27402 ;
  assign n27414 = ~n27407 & n27410 ;
  assign n27415 = ~n27409 & n27414 ;
  assign n27416 = n27413 & n27415 ;
  assign n27417 = ~n27408 & n27416 ;
  assign n27418 = ~\T_TMODE[1]_pad  & ~n27417 ;
  assign n27419 = ~n27400 & ~n27418 ;
  assign n27420 = \core_c_dec_rdCM_E_reg/NET0131  & ~n27419 ;
  assign n27421 = ~n27399 & ~n27420 ;
  assign n27422 = ~n26973 & ~n27421 ;
  assign n27398 = \sice_idr0_reg_DO_reg[9]/P0001  & n26973 ;
  assign n27423 = \sice_SPC_reg[9]/P0001  & n26969 ;
  assign n27424 = ~n27398 & ~n27423 ;
  assign n27425 = ~n27422 & n27424 ;
  assign n27427 = n8460 & n26970 ;
  assign n27428 = \T_TMODE[1]_pad  & \emc_ECMDreg_reg[11]/P0001  ;
  assign n27436 = \CM_rdm[11]_pad  & n27018 ;
  assign n27431 = \CM_rd0[11]_pad  & n26994 ;
  assign n27432 = \CM_rd7[11]_pad  & n26997 ;
  assign n27439 = ~n27431 & ~n27432 ;
  assign n27433 = \CM_rd2[11]_pad  & n27000 ;
  assign n27434 = \CM_rd5[11]_pad  & n27004 ;
  assign n27440 = ~n27433 & ~n27434 ;
  assign n27441 = n27439 & n27440 ;
  assign n27437 = \CM_rd3[11]_pad  & n27011 ;
  assign n27435 = \CM_rd4[11]_pad  & n27008 ;
  assign n27429 = \CM_rd1[11]_pad  & n26984 ;
  assign n27430 = \CM_rd6[11]_pad  & n26989 ;
  assign n27438 = ~n27429 & ~n27430 ;
  assign n27442 = ~n27435 & n27438 ;
  assign n27443 = ~n27437 & n27442 ;
  assign n27444 = n27441 & n27443 ;
  assign n27445 = ~n27436 & n27444 ;
  assign n27446 = ~\T_TMODE[1]_pad  & ~n27445 ;
  assign n27447 = ~n27428 & ~n27446 ;
  assign n27448 = \core_c_dec_rdCM_E_reg/NET0131  & ~n27447 ;
  assign n27449 = ~n27427 & ~n27448 ;
  assign n27450 = ~n26973 & ~n27449 ;
  assign n27426 = \sice_idr0_reg_DO_reg[11]/P0001  & n26973 ;
  assign n27451 = \sice_SPC_reg[11]/P0001  & n26969 ;
  assign n27452 = ~n27426 & ~n27451 ;
  assign n27453 = ~n27450 & n27452 ;
  assign n27455 = n7859 & n26970 ;
  assign n27456 = \T_TMODE[1]_pad  & \emc_ECMDreg_reg[10]/P0001  ;
  assign n27464 = \CM_rdm[10]_pad  & n27018 ;
  assign n27459 = \CM_rd0[10]_pad  & n26994 ;
  assign n27460 = \CM_rd7[10]_pad  & n26997 ;
  assign n27467 = ~n27459 & ~n27460 ;
  assign n27461 = \CM_rd2[10]_pad  & n27000 ;
  assign n27462 = \CM_rd5[10]_pad  & n27004 ;
  assign n27468 = ~n27461 & ~n27462 ;
  assign n27469 = n27467 & n27468 ;
  assign n27465 = \CM_rd3[10]_pad  & n27011 ;
  assign n27463 = \CM_rd4[10]_pad  & n27008 ;
  assign n27457 = \CM_rd1[10]_pad  & n26984 ;
  assign n27458 = \CM_rd6[10]_pad  & n26989 ;
  assign n27466 = ~n27457 & ~n27458 ;
  assign n27470 = ~n27463 & n27466 ;
  assign n27471 = ~n27465 & n27470 ;
  assign n27472 = n27469 & n27471 ;
  assign n27473 = ~n27464 & n27472 ;
  assign n27474 = ~\T_TMODE[1]_pad  & ~n27473 ;
  assign n27475 = ~n27456 & ~n27474 ;
  assign n27476 = \core_c_dec_rdCM_E_reg/NET0131  & ~n27475 ;
  assign n27477 = ~n27455 & ~n27476 ;
  assign n27478 = ~n26973 & ~n27477 ;
  assign n27454 = \sice_idr0_reg_DO_reg[10]/P0001  & n26973 ;
  assign n27479 = \sice_SPC_reg[10]/P0001  & n26969 ;
  assign n27480 = ~n27454 & ~n27479 ;
  assign n27481 = ~n27478 & n27480 ;
  assign n27482 = \core_c_dec_MTSE_E_reg/P0001  & ~n17814 ;
  assign n27483 = n26262 & n26263 ;
  assign n27484 = n26261 & n26269 ;
  assign n27485 = ~n27483 & n27484 ;
  assign n27486 = n26271 & n26273 ;
  assign n27487 = ~n27485 & n27486 ;
  assign n27488 = n26275 & ~n27487 ;
  assign n27489 = ~\core_c_dec_MTSE_E_reg/P0001  & ~n27488 ;
  assign n27490 = ~n27482 & ~n27489 ;
  assign n27491 = n23677 & ~n27490 ;
  assign n27492 = ~\core_eu_es_sht_es_reg_seswe_DO_reg[2]/P0001  & ~n23677 ;
  assign n27493 = ~n27491 & ~n27492 ;
  assign n27494 = n23598 & ~n27490 ;
  assign n27495 = ~\core_eu_es_sht_es_reg_serwe_DO_reg[2]/P0001  & ~n23598 ;
  assign n27496 = ~n27494 & ~n27495 ;
  assign n27498 = n13569 & ~n27028 ;
  assign n27499 = ~n5882 & n13569 ;
  assign n27500 = \idma_IADi_reg[7]/P0001  & ~n27499 ;
  assign n27501 = ~n13570 & ~n27500 ;
  assign n27502 = ~n27498 & n27501 ;
  assign n27497 = ~n13006 & n13570 ;
  assign n27503 = ~n11752 & ~n27497 ;
  assign n27504 = ~n27502 & n27503 ;
  assign n27505 = n11265 & n11752 ;
  assign n27506 = ~n27504 & ~n27505 ;
  assign n27507 = ~n12972 & n13570 ;
  assign n27508 = n13569 & ~n27075 ;
  assign n27509 = \idma_IADi_reg[6]/P0001  & ~n27499 ;
  assign n27510 = ~n13570 & ~n27509 ;
  assign n27511 = ~n27508 & n27510 ;
  assign n27512 = ~n11752 & ~n27511 ;
  assign n27513 = ~n27507 & n27512 ;
  assign n27514 = n11525 & n11752 ;
  assign n27515 = ~n27513 & ~n27514 ;
  assign n27517 = n13569 & ~n27333 ;
  assign n27518 = \idma_IADi_reg[5]/P0001  & ~n27499 ;
  assign n27519 = ~n13570 & ~n27518 ;
  assign n27520 = ~n27517 & n27519 ;
  assign n27516 = ~n12938 & n13570 ;
  assign n27521 = ~n11752 & ~n27516 ;
  assign n27522 = ~n27520 & n27521 ;
  assign n27523 = n10911 & n11752 ;
  assign n27524 = ~n27522 & ~n27523 ;
  assign n27526 = n13569 & ~n27361 ;
  assign n27527 = \idma_IADi_reg[4]/P0001  & ~n27499 ;
  assign n27528 = ~n13570 & ~n27527 ;
  assign n27529 = ~n27526 & n27528 ;
  assign n27525 = ~n12904 & n13570 ;
  assign n27530 = ~n11752 & ~n27525 ;
  assign n27531 = ~n27529 & n27530 ;
  assign n27532 = n10069 & n11752 ;
  assign n27533 = ~n27531 & ~n27532 ;
  assign n27535 = n13569 & ~n27445 ;
  assign n27536 = \idma_IADi_reg[3]/P0001  & ~n27499 ;
  assign n27537 = ~n13570 & ~n27536 ;
  assign n27538 = ~n27535 & n27537 ;
  assign n27534 = ~n12870 & n13570 ;
  assign n27539 = ~n11752 & ~n27534 ;
  assign n27540 = ~n27538 & n27539 ;
  assign n27541 = n8113 & n11752 ;
  assign n27542 = ~n27540 & ~n27541 ;
  assign n27544 = n13569 & ~n27473 ;
  assign n27545 = \idma_IADi_reg[2]/P0001  & ~n27499 ;
  assign n27546 = ~n13570 & ~n27545 ;
  assign n27547 = ~n27544 & n27546 ;
  assign n27543 = ~n12836 & n13570 ;
  assign n27548 = ~n11752 & ~n27543 ;
  assign n27549 = ~n27547 & n27548 ;
  assign n27550 = n8715 & n11752 ;
  assign n27551 = ~n27549 & ~n27550 ;
  assign n27553 = n13569 & ~n27417 ;
  assign n27554 = \idma_IADi_reg[1]/P0001  & ~n27499 ;
  assign n27555 = ~n13570 & ~n27554 ;
  assign n27556 = ~n27553 & n27555 ;
  assign n27552 = ~n12802 & n13570 ;
  assign n27557 = ~n11752 & ~n27552 ;
  assign n27558 = ~n27556 & n27557 ;
  assign n27559 = n9435 & n11752 ;
  assign n27560 = ~n27558 & ~n27559 ;
  assign n27568 = \CM_rdm[23]_pad  & n27018 ;
  assign n27563 = \CM_rd0[23]_pad  & n26994 ;
  assign n27564 = \CM_rd7[23]_pad  & n26997 ;
  assign n27571 = ~n27563 & ~n27564 ;
  assign n27565 = \CM_rd2[23]_pad  & n27000 ;
  assign n27566 = \CM_rd5[23]_pad  & n27004 ;
  assign n27572 = ~n27565 & ~n27566 ;
  assign n27573 = n27571 & n27572 ;
  assign n27569 = \CM_rd3[23]_pad  & n27011 ;
  assign n27567 = \CM_rd4[23]_pad  & n27008 ;
  assign n27561 = \CM_rd1[23]_pad  & n26984 ;
  assign n27562 = \CM_rd6[23]_pad  & n26989 ;
  assign n27570 = ~n27561 & ~n27562 ;
  assign n27574 = ~n27567 & n27570 ;
  assign n27575 = ~n27569 & n27574 ;
  assign n27576 = n27573 & n27575 ;
  assign n27577 = ~n27568 & n27576 ;
  assign n27578 = n27499 & ~n27577 ;
  assign n27579 = \idma_IADi_reg[15]/P0001  & ~n27499 ;
  assign n27580 = ~n27578 & ~n27579 ;
  assign n27581 = ~n13570 & ~n27580 ;
  assign n27582 = n12771 & n13570 ;
  assign n27583 = ~n27581 & ~n27582 ;
  assign n27584 = ~n11752 & ~n27583 ;
  assign n27585 = n11752 & n12743 ;
  assign n27586 = ~n27584 & ~n27585 ;
  assign n27594 = \CM_rdm[22]_pad  & n27018 ;
  assign n27589 = \CM_rd0[22]_pad  & n26994 ;
  assign n27590 = \CM_rd7[22]_pad  & n26997 ;
  assign n27597 = ~n27589 & ~n27590 ;
  assign n27591 = \CM_rd2[22]_pad  & n27000 ;
  assign n27592 = \CM_rd5[22]_pad  & n27004 ;
  assign n27598 = ~n27591 & ~n27592 ;
  assign n27599 = n27597 & n27598 ;
  assign n27595 = \CM_rd3[22]_pad  & n27011 ;
  assign n27593 = \CM_rd4[22]_pad  & n27008 ;
  assign n27587 = \CM_rd1[22]_pad  & n26984 ;
  assign n27588 = \CM_rd6[22]_pad  & n26989 ;
  assign n27596 = ~n27587 & ~n27588 ;
  assign n27600 = ~n27593 & n27596 ;
  assign n27601 = ~n27595 & n27600 ;
  assign n27602 = n27599 & n27601 ;
  assign n27603 = ~n27594 & n27602 ;
  assign n27604 = n27499 & ~n27603 ;
  assign n27605 = \idma_IADi_reg[14]/P0001  & ~n27499 ;
  assign n27606 = ~n27604 & ~n27605 ;
  assign n27607 = ~n13570 & ~n27606 ;
  assign n27608 = n12715 & n13570 ;
  assign n27609 = ~n27607 & ~n27608 ;
  assign n27610 = ~n11752 & ~n27609 ;
  assign n27611 = n11752 & n12688 ;
  assign n27612 = ~n27610 & ~n27611 ;
  assign n27614 = n13569 & ~n27389 ;
  assign n27615 = \idma_IADi_reg[0]/P0001  & ~n27499 ;
  assign n27616 = ~n13570 & ~n27615 ;
  assign n27617 = ~n27614 & n27616 ;
  assign n27613 = ~n12520 & n13570 ;
  assign n27618 = ~n11752 & ~n27613 ;
  assign n27619 = ~n27617 & n27618 ;
  assign n27620 = n7607 & n11752 ;
  assign n27621 = ~n27619 & ~n27620 ;
  assign n27622 = \tm_TSR_TMP_reg[5]/NET0131  & ~n25494 ;
  assign n27623 = ~n25495 & ~n27622 ;
  assign n27624 = n25491 & ~n27623 ;
  assign n27625 = \tm_tsr_reg_DO_reg[5]/NET0131  & ~n25491 ;
  assign n27626 = ~n27624 & ~n27625 ;
  assign n27634 = \CM_rdm[17]_pad  & n27018 ;
  assign n27629 = \CM_rd0[17]_pad  & n26994 ;
  assign n27630 = \CM_rd7[17]_pad  & n26997 ;
  assign n27637 = ~n27629 & ~n27630 ;
  assign n27631 = \CM_rd2[17]_pad  & n27000 ;
  assign n27632 = \CM_rd5[17]_pad  & n27004 ;
  assign n27638 = ~n27631 & ~n27632 ;
  assign n27639 = n27637 & n27638 ;
  assign n27635 = \CM_rd3[17]_pad  & n27011 ;
  assign n27633 = \CM_rd4[17]_pad  & n27008 ;
  assign n27627 = \CM_rd1[17]_pad  & n26984 ;
  assign n27628 = \CM_rd6[17]_pad  & n26989 ;
  assign n27636 = ~n27627 & ~n27628 ;
  assign n27640 = ~n27633 & n27636 ;
  assign n27641 = ~n27635 & n27640 ;
  assign n27642 = n27639 & n27641 ;
  assign n27643 = ~n27634 & n27642 ;
  assign n27644 = n27499 & ~n27643 ;
  assign n27645 = \idma_IADi_reg[9]/P0001  & ~n27499 ;
  assign n27646 = ~n27644 & ~n27645 ;
  assign n27647 = ~n13570 & ~n27646 ;
  assign n27648 = n13075 & n13570 ;
  assign n27649 = ~n27647 & ~n27648 ;
  assign n27650 = ~n11752 & ~n27649 ;
  assign n27651 = n10289 & n11752 ;
  assign n27652 = ~n27650 & ~n27651 ;
  assign n27660 = \CM_rdm[16]_pad  & n27018 ;
  assign n27655 = \CM_rd0[16]_pad  & n26994 ;
  assign n27656 = \CM_rd7[16]_pad  & n26997 ;
  assign n27663 = ~n27655 & ~n27656 ;
  assign n27657 = \CM_rd2[16]_pad  & n27000 ;
  assign n27658 = \CM_rd5[16]_pad  & n27004 ;
  assign n27664 = ~n27657 & ~n27658 ;
  assign n27665 = n27663 & n27664 ;
  assign n27661 = \CM_rd3[16]_pad  & n27011 ;
  assign n27659 = \CM_rd4[16]_pad  & n27008 ;
  assign n27653 = \CM_rd1[16]_pad  & n26984 ;
  assign n27654 = \CM_rd6[16]_pad  & n26989 ;
  assign n27662 = ~n27653 & ~n27654 ;
  assign n27666 = ~n27659 & n27662 ;
  assign n27667 = ~n27661 & n27666 ;
  assign n27668 = n27665 & n27667 ;
  assign n27669 = ~n27660 & n27668 ;
  assign n27670 = n27499 & ~n27669 ;
  assign n27671 = \idma_IADi_reg[8]/P0001  & ~n27499 ;
  assign n27672 = ~n27670 & ~n27671 ;
  assign n27673 = ~n13570 & ~n27672 ;
  assign n27674 = n13041 & n13570 ;
  assign n27675 = ~n27673 & ~n27674 ;
  assign n27676 = ~n11752 & ~n27675 ;
  assign n27677 = n10638 & n11752 ;
  assign n27678 = ~n27676 & ~n27677 ;
  assign n27686 = \CM_rdm[21]_pad  & n27018 ;
  assign n27681 = \CM_rd0[21]_pad  & n26994 ;
  assign n27682 = \CM_rd7[21]_pad  & n26997 ;
  assign n27689 = ~n27681 & ~n27682 ;
  assign n27683 = \CM_rd2[21]_pad  & n27000 ;
  assign n27684 = \CM_rd5[21]_pad  & n27004 ;
  assign n27690 = ~n27683 & ~n27684 ;
  assign n27691 = n27689 & n27690 ;
  assign n27687 = \CM_rd3[21]_pad  & n27011 ;
  assign n27685 = \CM_rd4[21]_pad  & n27008 ;
  assign n27679 = \CM_rd1[21]_pad  & n26984 ;
  assign n27680 = \CM_rd6[21]_pad  & n26989 ;
  assign n27688 = ~n27679 & ~n27680 ;
  assign n27692 = ~n27685 & n27688 ;
  assign n27693 = ~n27687 & n27692 ;
  assign n27694 = n27691 & n27693 ;
  assign n27695 = ~n27686 & n27694 ;
  assign n27696 = n27499 & ~n27695 ;
  assign n27697 = \idma_IADi_reg[13]/P0001  & ~n27499 ;
  assign n27698 = ~n27696 & ~n27697 ;
  assign n27699 = ~n13570 & ~n27698 ;
  assign n27700 = n12658 & n13570 ;
  assign n27701 = ~n27699 & ~n27700 ;
  assign n27702 = ~n11752 & ~n27701 ;
  assign n27703 = n7340 & n11752 ;
  assign n27704 = ~n27702 & ~n27703 ;
  assign n27712 = \CM_rdm[20]_pad  & n27018 ;
  assign n27707 = \CM_rd0[20]_pad  & n26994 ;
  assign n27708 = \CM_rd7[20]_pad  & n26997 ;
  assign n27715 = ~n27707 & ~n27708 ;
  assign n27709 = \CM_rd2[20]_pad  & n27000 ;
  assign n27710 = \CM_rd5[20]_pad  & n27004 ;
  assign n27716 = ~n27709 & ~n27710 ;
  assign n27717 = n27715 & n27716 ;
  assign n27713 = \CM_rd3[20]_pad  & n27011 ;
  assign n27711 = \CM_rd4[20]_pad  & n27008 ;
  assign n27705 = \CM_rd1[20]_pad  & n26984 ;
  assign n27706 = \CM_rd6[20]_pad  & n26989 ;
  assign n27714 = ~n27705 & ~n27706 ;
  assign n27718 = ~n27711 & n27714 ;
  assign n27719 = ~n27713 & n27718 ;
  assign n27720 = n27717 & n27719 ;
  assign n27721 = ~n27712 & n27720 ;
  assign n27722 = n27499 & ~n27721 ;
  assign n27723 = \idma_IADi_reg[12]/P0001  & ~n27499 ;
  assign n27724 = ~n27722 & ~n27723 ;
  assign n27725 = ~n13570 & ~n27724 ;
  assign n27726 = n12624 & n13570 ;
  assign n27727 = ~n27725 & ~n27726 ;
  assign n27728 = ~n11752 & ~n27727 ;
  assign n27729 = n9178 & n11752 ;
  assign n27730 = ~n27728 & ~n27729 ;
  assign n27738 = \CM_rdm[19]_pad  & n27018 ;
  assign n27733 = \CM_rd0[19]_pad  & n26994 ;
  assign n27734 = \CM_rd7[19]_pad  & n26997 ;
  assign n27741 = ~n27733 & ~n27734 ;
  assign n27735 = \CM_rd2[19]_pad  & n27000 ;
  assign n27736 = \CM_rd5[19]_pad  & n27004 ;
  assign n27742 = ~n27735 & ~n27736 ;
  assign n27743 = n27741 & n27742 ;
  assign n27739 = \CM_rd3[19]_pad  & n27011 ;
  assign n27737 = \CM_rd4[19]_pad  & n27008 ;
  assign n27731 = \CM_rd1[19]_pad  & n26984 ;
  assign n27732 = \CM_rd6[19]_pad  & n26989 ;
  assign n27740 = ~n27731 & ~n27732 ;
  assign n27744 = ~n27737 & n27740 ;
  assign n27745 = ~n27739 & n27744 ;
  assign n27746 = n27743 & n27745 ;
  assign n27747 = ~n27738 & n27746 ;
  assign n27748 = n27499 & ~n27747 ;
  assign n27749 = \idma_IADi_reg[11]/P0001  & ~n27499 ;
  assign n27750 = ~n27748 & ~n27749 ;
  assign n27751 = ~n13570 & ~n27750 ;
  assign n27752 = n12590 & n13570 ;
  assign n27753 = ~n27751 & ~n27752 ;
  assign n27754 = ~n11752 & ~n27753 ;
  assign n27755 = n8460 & n11752 ;
  assign n27756 = ~n27754 & ~n27755 ;
  assign n27764 = \CM_rdm[18]_pad  & n27018 ;
  assign n27759 = \CM_rd0[18]_pad  & n26994 ;
  assign n27760 = \CM_rd7[18]_pad  & n26997 ;
  assign n27767 = ~n27759 & ~n27760 ;
  assign n27761 = \CM_rd2[18]_pad  & n27000 ;
  assign n27762 = \CM_rd5[18]_pad  & n27004 ;
  assign n27768 = ~n27761 & ~n27762 ;
  assign n27769 = n27767 & n27768 ;
  assign n27765 = \CM_rd3[18]_pad  & n27011 ;
  assign n27763 = \CM_rd4[18]_pad  & n27008 ;
  assign n27757 = \CM_rd1[18]_pad  & n26984 ;
  assign n27758 = \CM_rd6[18]_pad  & n26989 ;
  assign n27766 = ~n27757 & ~n27758 ;
  assign n27770 = ~n27763 & n27766 ;
  assign n27771 = ~n27765 & n27770 ;
  assign n27772 = n27769 & n27771 ;
  assign n27773 = ~n27764 & n27772 ;
  assign n27774 = n27499 & ~n27773 ;
  assign n27775 = \idma_IADi_reg[10]/P0001  & ~n27499 ;
  assign n27776 = ~n27774 & ~n27775 ;
  assign n27777 = ~n13570 & ~n27776 ;
  assign n27778 = n12556 & n13570 ;
  assign n27779 = ~n27777 & ~n27778 ;
  assign n27780 = ~n11752 & ~n27779 ;
  assign n27781 = n7859 & n11752 ;
  assign n27782 = ~n27780 & ~n27781 ;
  assign n27783 = ~n6931 & ~n6988 ;
  assign n27784 = ~n13567 & ~n27783 ;
  assign n27785 = n13564 & ~n27784 ;
  assign n27786 = n13597 & ~n27785 ;
  assign n27788 = ~n17814 & n19499 ;
  assign n27787 = ~\core_eu_em_mac_em_reg_mr1swe_DO_reg[2]/P0001  & ~n19499 ;
  assign n27789 = n19501 & ~n27787 ;
  assign n27790 = ~n27788 & n27789 ;
  assign n27791 = \core_eu_em_mac_em_reg_mr1swe_DO_reg[2]/P0001  & ~n19383 ;
  assign n27792 = ~n19508 & ~n27791 ;
  assign n27793 = ~n27790 & n27792 ;
  assign n27794 = ~n18262 & ~n27793 ;
  assign n27795 = ~\core_c_psq_MSTAT_reg_DO_reg[4]/NET0131  & ~n27051 ;
  assign n27796 = ~n17613 & ~n17672 ;
  assign n27797 = ~n17638 & ~n27048 ;
  assign n27798 = ~n17665 & ~n27797 ;
  assign n27799 = n27796 & ~n27798 ;
  assign n27800 = ~n27796 & n27798 ;
  assign n27801 = ~n27799 & ~n27800 ;
  assign n27802 = \core_c_psq_MSTAT_reg_DO_reg[4]/NET0131  & ~n27801 ;
  assign n27803 = ~n27795 & ~n27802 ;
  assign n27804 = n18262 & n27803 ;
  assign n27805 = ~n27794 & ~n27804 ;
  assign n27807 = n19499 & ~n21663 ;
  assign n27806 = ~\core_eu_em_mac_em_reg_mr1swe_DO_reg[3]/P0001  & ~n19499 ;
  assign n27808 = n19501 & ~n27806 ;
  assign n27809 = ~n27807 & n27808 ;
  assign n27810 = \core_eu_em_mac_em_reg_mr1swe_DO_reg[3]/P0001  & ~n19383 ;
  assign n27811 = ~n19508 & ~n27810 ;
  assign n27812 = ~n27809 & n27811 ;
  assign n27813 = ~n18262 & ~n27812 ;
  assign n27814 = ~\core_c_psq_MSTAT_reg_DO_reg[4]/NET0131  & n27801 ;
  assign n27815 = \core_c_psq_MSTAT_reg_DO_reg[4]/NET0131  & n26315 ;
  assign n27816 = ~n27814 & ~n27815 ;
  assign n27817 = n18262 & ~n27816 ;
  assign n27818 = ~n27813 & ~n27817 ;
  assign n27819 = n14752 & n27816 ;
  assign n27820 = n19776 & n21663 ;
  assign n27821 = \core_eu_em_mac_em_reg_mr1rwe_DO_reg[3]/P0001  & ~n17809 ;
  assign n27822 = n19780 & ~n27821 ;
  assign n27823 = ~n27820 & n27822 ;
  assign n27824 = ~n27819 & ~n27823 ;
  assign n27825 = n14752 & ~n27803 ;
  assign n27826 = n17814 & n19776 ;
  assign n27827 = \core_eu_em_mac_em_reg_mr1rwe_DO_reg[2]/P0001  & ~n17809 ;
  assign n27828 = n19780 & ~n27827 ;
  assign n27829 = ~n27826 & n27828 ;
  assign n27830 = ~n27825 & ~n27829 ;
  assign n27833 = n18271 & ~n20150 ;
  assign n27832 = ~\core_eu_em_mac_em_reg_mr0swe_DO_reg[14]/P0001  & ~n18271 ;
  assign n27834 = n18273 & ~n27832 ;
  assign n27835 = ~n27833 & n27834 ;
  assign n27831 = \core_eu_em_mac_em_reg_mr0swe_DO_reg[14]/P0001  & ~n18266 ;
  assign n27836 = ~n18270 & ~n27831 ;
  assign n27837 = ~n27835 & n27836 ;
  assign n27838 = ~n18262 & ~n27837 ;
  assign n27839 = n18262 & ~n19593 ;
  assign n27840 = ~n27838 & ~n27839 ;
  assign n27841 = n14752 & n19593 ;
  assign n27842 = n18328 & n20150 ;
  assign n27843 = \core_eu_em_mac_em_reg_mr0rwe_DO_reg[14]/P0001  & ~n18330 ;
  assign n27844 = n18334 & ~n27843 ;
  assign n27845 = ~n27842 & n27844 ;
  assign n27846 = ~n27841 & ~n27845 ;
  assign n27849 = ~n17814 & n18271 ;
  assign n27848 = ~\core_eu_em_mac_em_reg_mr0swe_DO_reg[2]/P0001  & ~n18271 ;
  assign n27850 = n18273 & ~n27848 ;
  assign n27851 = ~n27849 & n27850 ;
  assign n27847 = \core_eu_em_mac_em_reg_mr0swe_DO_reg[2]/P0001  & ~n18266 ;
  assign n27852 = ~n18270 & ~n27847 ;
  assign n27853 = ~n27851 & n27852 ;
  assign n27854 = ~n18262 & ~n27853 ;
  assign n27855 = n18262 & ~n19673 ;
  assign n27856 = ~n27854 & ~n27855 ;
  assign n27857 = n14752 & n19673 ;
  assign n27858 = n17814 & n18328 ;
  assign n27859 = \core_eu_em_mac_em_reg_mr0rwe_DO_reg[2]/P0001  & ~n18330 ;
  assign n27860 = n18334 & ~n27859 ;
  assign n27861 = ~n27858 & n27860 ;
  assign n27862 = ~n27857 & ~n27861 ;
  assign n27865 = ~n17820 & n18271 ;
  assign n27864 = ~\core_eu_em_mac_em_reg_mr0swe_DO_reg[15]/P0001  & ~n18271 ;
  assign n27866 = n18273 & ~n27864 ;
  assign n27867 = ~n27865 & n27866 ;
  assign n27863 = \core_eu_em_mac_em_reg_mr0swe_DO_reg[15]/P0001  & ~n18266 ;
  assign n27868 = ~n18270 & ~n27863 ;
  assign n27869 = ~n27867 & n27868 ;
  assign n27870 = ~n18262 & ~n27869 ;
  assign n27871 = n18262 & ~n19596 ;
  assign n27872 = ~n27870 & ~n27871 ;
  assign n27873 = ~n13806 & n14564 ;
  assign n27874 = n11975 & n13806 ;
  assign n27875 = ~n27873 & ~n27874 ;
  assign n27876 = n14667 & ~n27875 ;
  assign n27877 = ~\core_eu_ea_alu_ea_reg_afswe_DO_reg[0]/P0001  & ~n14667 ;
  assign n27878 = ~n27876 & ~n27877 ;
  assign n27879 = n13805 & ~n27875 ;
  assign n27880 = ~\core_eu_ea_alu_ea_reg_afrwe_DO_reg[0]/P0001  & ~n13805 ;
  assign n27881 = ~n27879 & ~n27880 ;
  assign n27882 = n14752 & n19596 ;
  assign n27883 = n17820 & n18328 ;
  assign n27884 = \core_eu_em_mac_em_reg_mr0rwe_DO_reg[15]/P0001  & ~n18330 ;
  assign n27885 = n18334 & ~n27884 ;
  assign n27886 = ~n27883 & n27885 ;
  assign n27887 = ~n27882 & ~n27886 ;
  assign n27888 = \tm_tcr_reg_DO_reg[7]/NET0131  & n20355 ;
  assign n27890 = ~\T_TMODE[0]_pad  & ~n20360 ;
  assign n27893 = ~\tm_TCR_TMP_reg[4]/NET0131  & ~n27890 ;
  assign n27894 = ~\tm_TCR_TMP_reg[5]/NET0131  & n27893 ;
  assign n27895 = n22411 & n27894 ;
  assign n27896 = ~\tm_TCR_TMP_reg[6]/NET0131  & n27895 ;
  assign n27897 = \tm_TCR_TMP_reg[7]/NET0131  & ~n27896 ;
  assign n27891 = n20363 & ~n27890 ;
  assign n27892 = n22411 & n27891 ;
  assign n27898 = ~n22400 & ~n27892 ;
  assign n27899 = ~n27897 & n27898 ;
  assign n27889 = ~\tm_tpr_reg_DO_reg[7]/NET0131  & n22400 ;
  assign n27900 = ~n20355 & ~n27889 ;
  assign n27901 = ~n27899 & n27900 ;
  assign n27902 = ~n27888 & ~n27901 ;
  assign n27903 = n23407 & n25053 ;
  assign n27904 = n23032 & n27903 ;
  assign n27905 = n25749 & n25752 ;
  assign n27906 = n4186 & n27905 ;
  assign n27909 = \core_c_dec_BR_Ed_reg/P0001  & ~\core_c_dec_IRE_reg[0]/NET0131  ;
  assign n27910 = \core_c_dec_IRE_reg[1]/NET0131  & n27909 ;
  assign n27911 = n6071 & n27910 ;
  assign n27907 = \core_c_dec_IRE_reg[2]/NET0131  & \core_c_dec_Stkctl_Eg_reg/P0001  ;
  assign n27908 = ~\core_c_dec_MTCNTR_Eg_reg/P0001  & ~\core_c_dec_MTOWRCNTR_Eg_reg/P0001  ;
  assign n27912 = ~n27907 & n27908 ;
  assign n27913 = ~n27911 & n27912 ;
  assign n27914 = ~n27906 & n27913 ;
  assign n27915 = ~n5950 & ~n27914 ;
  assign n27916 = \core_c_psq_CE_reg/NET0131  & ~n27915 ;
  assign n27918 = n4842 & n27905 ;
  assign n27917 = \core_c_psq_CE_reg/NET0131  & n27911 ;
  assign n27919 = ~n27907 & ~n27917 ;
  assign n27920 = ~n27918 & n27919 ;
  assign n27921 = ~\core_c_psq_cntstk_ptr_reg[2]/NET0131  & ~n27920 ;
  assign n27922 = ~\core_c_psq_CNTR_reg_DO_reg[0]/NET0131  & ~\core_c_psq_CNTR_reg_DO_reg[1]/NET0131  ;
  assign n27923 = ~\core_c_psq_CNTR_reg_DO_reg[2]/NET0131  & n27922 ;
  assign n27924 = ~\core_c_psq_CNTR_reg_DO_reg[3]/NET0131  & n27923 ;
  assign n27925 = ~\core_c_psq_CNTR_reg_DO_reg[4]/NET0131  & n27924 ;
  assign n27926 = ~\core_c_psq_CNTR_reg_DO_reg[5]/NET0131  & n27925 ;
  assign n27927 = ~\core_c_psq_CNTR_reg_DO_reg[6]/NET0131  & n27926 ;
  assign n27928 = ~\core_c_psq_CNTR_reg_DO_reg[7]/NET0131  & n27927 ;
  assign n27929 = ~\core_c_psq_CNTR_reg_DO_reg[8]/NET0131  & n27928 ;
  assign n27930 = ~\core_c_psq_CNTR_reg_DO_reg[9]/NET0131  & n27929 ;
  assign n27931 = ~\core_c_psq_CNTR_reg_DO_reg[10]/NET0131  & n27930 ;
  assign n27932 = ~\core_c_psq_CNTR_reg_DO_reg[11]/NET0131  & n27931 ;
  assign n27933 = ~\core_c_psq_CNTR_reg_DO_reg[12]/NET0131  & n27932 ;
  assign n27934 = \core_c_psq_CNTR_reg_DO_reg[12]/NET0131  & ~n27932 ;
  assign n27935 = ~n27933 & ~n27934 ;
  assign n27936 = ~n27921 & ~n27935 ;
  assign n27937 = \core_c_psq_cntstk_cnts4x14_CNTcell_reg[3][12]/P0001  & n13775 ;
  assign n27938 = \core_c_psq_cntstk_cnts4x14_CNTcell_reg[1][12]/P0001  & n13789 ;
  assign n27941 = ~n27937 & ~n27938 ;
  assign n27939 = \core_c_psq_cntstk_cnts4x14_CNTcell_reg[2][12]/P0001  & n13794 ;
  assign n27940 = \core_c_psq_cntstk_cnts4x14_CNTcell_reg[0][12]/P0001  & n13784 ;
  assign n27942 = ~n27939 & ~n27940 ;
  assign n27943 = n27941 & n27942 ;
  assign n27944 = n27921 & ~n27943 ;
  assign n27945 = ~n27936 & ~n27944 ;
  assign n27946 = n27908 & ~n27945 ;
  assign n27947 = n9178 & ~n27908 ;
  assign n27948 = ~n27946 & ~n27947 ;
  assign n27949 = \core_c_psq_CNTR_reg_DO_reg[10]/NET0131  & ~n27930 ;
  assign n27950 = ~n27931 & ~n27949 ;
  assign n27951 = ~n27921 & ~n27950 ;
  assign n27952 = \core_c_psq_cntstk_cnts4x14_CNTcell_reg[3][10]/P0001  & n13775 ;
  assign n27953 = \core_c_psq_cntstk_cnts4x14_CNTcell_reg[0][10]/P0001  & n13784 ;
  assign n27956 = ~n27952 & ~n27953 ;
  assign n27954 = \core_c_psq_cntstk_cnts4x14_CNTcell_reg[1][10]/P0001  & n13789 ;
  assign n27955 = \core_c_psq_cntstk_cnts4x14_CNTcell_reg[2][10]/P0001  & n13794 ;
  assign n27957 = ~n27954 & ~n27955 ;
  assign n27958 = n27956 & n27957 ;
  assign n27959 = n27921 & ~n27958 ;
  assign n27960 = ~n27951 & ~n27959 ;
  assign n27961 = n27908 & ~n27960 ;
  assign n27962 = n7859 & ~n27908 ;
  assign n27963 = ~n27961 & ~n27962 ;
  assign n28144 = n27948 & n27963 ;
  assign n27964 = \core_c_psq_CNTR_reg_DO_reg[8]/NET0131  & ~n27928 ;
  assign n27965 = ~n27929 & ~n27964 ;
  assign n27966 = ~n27921 & ~n27965 ;
  assign n27967 = \core_c_psq_cntstk_cnts4x14_CNTcell_reg[3][8]/P0001  & n13775 ;
  assign n27968 = \core_c_psq_cntstk_cnts4x14_CNTcell_reg[2][8]/P0001  & n13794 ;
  assign n27971 = ~n27967 & ~n27968 ;
  assign n27969 = \core_c_psq_cntstk_cnts4x14_CNTcell_reg[1][8]/P0001  & n13789 ;
  assign n27970 = \core_c_psq_cntstk_cnts4x14_CNTcell_reg[0][8]/P0001  & n13784 ;
  assign n27972 = ~n27969 & ~n27970 ;
  assign n27973 = n27971 & n27972 ;
  assign n27974 = n27921 & ~n27973 ;
  assign n27975 = ~n27966 & ~n27974 ;
  assign n27976 = n27908 & ~n27975 ;
  assign n27977 = n10638 & ~n27908 ;
  assign n27978 = ~n27976 & ~n27977 ;
  assign n27979 = \core_c_psq_CNTR_reg_DO_reg[4]/NET0131  & ~n27924 ;
  assign n27980 = ~n27925 & ~n27979 ;
  assign n27981 = ~n27921 & ~n27980 ;
  assign n27982 = \core_c_psq_cntstk_cnts4x14_CNTcell_reg[2][4]/P0001  & n13794 ;
  assign n27983 = \core_c_psq_cntstk_cnts4x14_CNTcell_reg[1][4]/P0001  & n13789 ;
  assign n27986 = ~n27982 & ~n27983 ;
  assign n27984 = \core_c_psq_cntstk_cnts4x14_CNTcell_reg[3][4]/P0001  & n13775 ;
  assign n27985 = \core_c_psq_cntstk_cnts4x14_CNTcell_reg[0][4]/P0001  & n13784 ;
  assign n27987 = ~n27984 & ~n27985 ;
  assign n27988 = n27986 & n27987 ;
  assign n27989 = n27921 & ~n27988 ;
  assign n27990 = ~n27981 & ~n27989 ;
  assign n27991 = n27908 & ~n27990 ;
  assign n27992 = n10069 & ~n27908 ;
  assign n27993 = ~n27991 & ~n27992 ;
  assign n28145 = n27978 & n27993 ;
  assign n27994 = n9435 & ~n27908 ;
  assign n28003 = \core_c_psq_CNTR_reg_DO_reg[0]/NET0131  & \core_c_psq_CNTR_reg_DO_reg[1]/NET0131  ;
  assign n28004 = ~n27922 & ~n28003 ;
  assign n28005 = ~n27921 & n28004 ;
  assign n27995 = \core_c_psq_cntstk_cnts4x14_CNTcell_reg[0][1]/P0001  & n13784 ;
  assign n27996 = \core_c_psq_cntstk_cnts4x14_CNTcell_reg[3][1]/P0001  & n13775 ;
  assign n27999 = ~n27995 & ~n27996 ;
  assign n27997 = \core_c_psq_cntstk_cnts4x14_CNTcell_reg[2][1]/P0001  & n13794 ;
  assign n27998 = \core_c_psq_cntstk_cnts4x14_CNTcell_reg[1][1]/P0001  & n13789 ;
  assign n28000 = ~n27997 & ~n27998 ;
  assign n28001 = n27999 & n28000 ;
  assign n28002 = n27921 & n28001 ;
  assign n28006 = n27908 & ~n28002 ;
  assign n28007 = ~n28005 & n28006 ;
  assign n28008 = ~n27994 & ~n28007 ;
  assign n28009 = \core_c_psq_CNTR_reg_DO_reg[9]/NET0131  & ~n27929 ;
  assign n28010 = ~n27930 & ~n28009 ;
  assign n28011 = ~n27921 & ~n28010 ;
  assign n28012 = \core_c_psq_cntstk_cnts4x14_CNTcell_reg[3][9]/P0001  & n13775 ;
  assign n28013 = \core_c_psq_cntstk_cnts4x14_CNTcell_reg[2][9]/P0001  & n13794 ;
  assign n28016 = ~n28012 & ~n28013 ;
  assign n28014 = \core_c_psq_cntstk_cnts4x14_CNTcell_reg[1][9]/P0001  & n13789 ;
  assign n28015 = \core_c_psq_cntstk_cnts4x14_CNTcell_reg[0][9]/P0001  & n13784 ;
  assign n28017 = ~n28014 & ~n28015 ;
  assign n28018 = n28016 & n28017 ;
  assign n28019 = n27921 & ~n28018 ;
  assign n28020 = ~n28011 & ~n28019 ;
  assign n28021 = n27908 & ~n28020 ;
  assign n28022 = n10289 & ~n27908 ;
  assign n28023 = ~n28021 & ~n28022 ;
  assign n28146 = n28008 & n28023 ;
  assign n28153 = n28145 & n28146 ;
  assign n28154 = n28144 & n28153 ;
  assign n28084 = \core_c_psq_CNTR_reg_DO_reg[7]/NET0131  & ~n27927 ;
  assign n28085 = ~n27928 & ~n28084 ;
  assign n28086 = ~n27921 & ~n28085 ;
  assign n28087 = \core_c_psq_cntstk_cnts4x14_CNTcell_reg[2][7]/P0001  & n13794 ;
  assign n28088 = \core_c_psq_cntstk_cnts4x14_CNTcell_reg[1][7]/P0001  & n13789 ;
  assign n28091 = ~n28087 & ~n28088 ;
  assign n28089 = \core_c_psq_cntstk_cnts4x14_CNTcell_reg[0][7]/P0001  & n13784 ;
  assign n28090 = \core_c_psq_cntstk_cnts4x14_CNTcell_reg[3][7]/P0001  & n13775 ;
  assign n28092 = ~n28089 & ~n28090 ;
  assign n28093 = n28091 & n28092 ;
  assign n28094 = n27921 & ~n28093 ;
  assign n28095 = ~n28086 & ~n28094 ;
  assign n28096 = n27908 & ~n28095 ;
  assign n28097 = n11265 & ~n27908 ;
  assign n28098 = ~n28096 & ~n28097 ;
  assign n28099 = \core_c_psq_CNTR_reg_DO_reg[6]/NET0131  & ~n27926 ;
  assign n28100 = ~n27927 & ~n28099 ;
  assign n28101 = ~n27921 & ~n28100 ;
  assign n28102 = \core_c_psq_cntstk_cnts4x14_CNTcell_reg[3][6]/P0001  & n13775 ;
  assign n28103 = \core_c_psq_cntstk_cnts4x14_CNTcell_reg[0][6]/P0001  & n13784 ;
  assign n28106 = ~n28102 & ~n28103 ;
  assign n28104 = \core_c_psq_cntstk_cnts4x14_CNTcell_reg[1][6]/P0001  & n13789 ;
  assign n28105 = \core_c_psq_cntstk_cnts4x14_CNTcell_reg[2][6]/P0001  & n13794 ;
  assign n28107 = ~n28104 & ~n28105 ;
  assign n28108 = n28106 & n28107 ;
  assign n28109 = n27921 & ~n28108 ;
  assign n28110 = ~n28101 & ~n28109 ;
  assign n28111 = n27908 & ~n28110 ;
  assign n28112 = n11525 & ~n27908 ;
  assign n28113 = ~n28111 & ~n28112 ;
  assign n28149 = n28098 & n28113 ;
  assign n28114 = \core_c_psq_CNTR_reg_DO_reg[5]/NET0131  & ~n27925 ;
  assign n28115 = ~n27926 & ~n28114 ;
  assign n28116 = ~n27921 & ~n28115 ;
  assign n28117 = \core_c_psq_cntstk_cnts4x14_CNTcell_reg[3][5]/P0001  & n13775 ;
  assign n28118 = \core_c_psq_cntstk_cnts4x14_CNTcell_reg[0][5]/P0001  & n13784 ;
  assign n28121 = ~n28117 & ~n28118 ;
  assign n28119 = \core_c_psq_cntstk_cnts4x14_CNTcell_reg[2][5]/P0001  & n13794 ;
  assign n28120 = \core_c_psq_cntstk_cnts4x14_CNTcell_reg[1][5]/P0001  & n13789 ;
  assign n28122 = ~n28119 & ~n28120 ;
  assign n28123 = n28121 & n28122 ;
  assign n28124 = n27921 & ~n28123 ;
  assign n28125 = ~n28116 & ~n28124 ;
  assign n28126 = n27908 & ~n28125 ;
  assign n28127 = n10911 & ~n27908 ;
  assign n28128 = ~n28126 & ~n28127 ;
  assign n28129 = \core_c_psq_CNTR_reg_DO_reg[11]/NET0131  & ~n27931 ;
  assign n28130 = ~n27932 & ~n28129 ;
  assign n28131 = ~n27921 & ~n28130 ;
  assign n28132 = \core_c_psq_cntstk_cnts4x14_CNTcell_reg[3][11]/P0001  & n13775 ;
  assign n28133 = \core_c_psq_cntstk_cnts4x14_CNTcell_reg[0][11]/P0001  & n13784 ;
  assign n28136 = ~n28132 & ~n28133 ;
  assign n28134 = \core_c_psq_cntstk_cnts4x14_CNTcell_reg[1][11]/P0001  & n13789 ;
  assign n28135 = \core_c_psq_cntstk_cnts4x14_CNTcell_reg[2][11]/P0001  & n13794 ;
  assign n28137 = ~n28134 & ~n28135 ;
  assign n28138 = n28136 & n28137 ;
  assign n28139 = n27921 & ~n28138 ;
  assign n28140 = ~n28131 & ~n28139 ;
  assign n28141 = n27908 & ~n28140 ;
  assign n28142 = n8460 & ~n27908 ;
  assign n28143 = ~n28141 & ~n28142 ;
  assign n28150 = n28128 & n28143 ;
  assign n28151 = n28149 & n28150 ;
  assign n28024 = \core_c_psq_CNTR_reg_DO_reg[3]/NET0131  & ~n27923 ;
  assign n28025 = ~n27924 & ~n28024 ;
  assign n28026 = ~n27921 & ~n28025 ;
  assign n28027 = \core_c_psq_cntstk_cnts4x14_CNTcell_reg[2][3]/P0001  & n13794 ;
  assign n28028 = \core_c_psq_cntstk_cnts4x14_CNTcell_reg[1][3]/P0001  & n13789 ;
  assign n28031 = ~n28027 & ~n28028 ;
  assign n28029 = \core_c_psq_cntstk_cnts4x14_CNTcell_reg[3][3]/P0001  & n13775 ;
  assign n28030 = \core_c_psq_cntstk_cnts4x14_CNTcell_reg[0][3]/P0001  & n13784 ;
  assign n28032 = ~n28029 & ~n28030 ;
  assign n28033 = n28031 & n28032 ;
  assign n28034 = n27921 & ~n28033 ;
  assign n28035 = ~n28026 & ~n28034 ;
  assign n28036 = n27908 & ~n28035 ;
  assign n28037 = n8113 & ~n27908 ;
  assign n28038 = ~n28036 & ~n28037 ;
  assign n28039 = n7340 & ~n27908 ;
  assign n28044 = \core_c_psq_cntstk_cnts4x14_CNTcell_reg[0][13]/P0001  & n13784 ;
  assign n28045 = \core_c_psq_cntstk_cnts4x14_CNTcell_reg[3][13]/P0001  & n13775 ;
  assign n28048 = ~n28044 & ~n28045 ;
  assign n28046 = \core_c_psq_cntstk_cnts4x14_CNTcell_reg[2][13]/P0001  & n13794 ;
  assign n28047 = \core_c_psq_cntstk_cnts4x14_CNTcell_reg[1][13]/P0001  & n13789 ;
  assign n28049 = ~n28046 & ~n28047 ;
  assign n28050 = n28048 & n28049 ;
  assign n28051 = n27921 & n28050 ;
  assign n28040 = \core_c_psq_CNTR_reg_DO_reg[13]/NET0131  & ~n27933 ;
  assign n28041 = ~\core_c_psq_CNTR_reg_DO_reg[13]/NET0131  & n27933 ;
  assign n28042 = ~n28040 & ~n28041 ;
  assign n28043 = ~n27921 & n28042 ;
  assign n28052 = n27908 & ~n28043 ;
  assign n28053 = ~n28051 & n28052 ;
  assign n28054 = ~n28039 & ~n28053 ;
  assign n28147 = n28038 & n28054 ;
  assign n28055 = \core_c_psq_CNTR_reg_DO_reg[2]/NET0131  & ~n27922 ;
  assign n28056 = ~n27923 & ~n28055 ;
  assign n28057 = ~n27921 & ~n28056 ;
  assign n28058 = \core_c_psq_cntstk_cnts4x14_CNTcell_reg[2][2]/P0001  & n13794 ;
  assign n28059 = \core_c_psq_cntstk_cnts4x14_CNTcell_reg[1][2]/P0001  & n13789 ;
  assign n28062 = ~n28058 & ~n28059 ;
  assign n28060 = \core_c_psq_cntstk_cnts4x14_CNTcell_reg[3][2]/P0001  & n13775 ;
  assign n28061 = \core_c_psq_cntstk_cnts4x14_CNTcell_reg[0][2]/P0001  & n13784 ;
  assign n28063 = ~n28060 & ~n28061 ;
  assign n28064 = n28062 & n28063 ;
  assign n28065 = n27921 & ~n28064 ;
  assign n28066 = ~n28057 & ~n28065 ;
  assign n28067 = n27908 & ~n28066 ;
  assign n28068 = n8715 & ~n27908 ;
  assign n28069 = ~n28067 & ~n28068 ;
  assign n28072 = \core_c_psq_cntstk_cnts4x14_CNTcell_reg[0][0]/P0001  & n13784 ;
  assign n28073 = \core_c_psq_cntstk_cnts4x14_CNTcell_reg[2][0]/P0001  & n13794 ;
  assign n28076 = ~n28072 & ~n28073 ;
  assign n28074 = \core_c_psq_cntstk_cnts4x14_CNTcell_reg[1][0]/P0001  & n13789 ;
  assign n28075 = \core_c_psq_cntstk_cnts4x14_CNTcell_reg[3][0]/P0001  & n13775 ;
  assign n28077 = ~n28074 & ~n28075 ;
  assign n28078 = n28076 & n28077 ;
  assign n28079 = n27921 & ~n28078 ;
  assign n28071 = ~\core_c_psq_CNTR_reg_DO_reg[0]/NET0131  & ~n27921 ;
  assign n28080 = n27908 & ~n28071 ;
  assign n28081 = ~n28079 & n28080 ;
  assign n28070 = ~n7607 & ~n27908 ;
  assign n28082 = n27915 & ~n28070 ;
  assign n28083 = ~n28081 & n28082 ;
  assign n28148 = n28069 & n28083 ;
  assign n28152 = n28147 & n28148 ;
  assign n28155 = n28151 & n28152 ;
  assign n28156 = n28154 & n28155 ;
  assign n28157 = ~n27916 & ~n28156 ;
  assign n28158 = ~n27103 & n27499 ;
  assign n28159 = ~n27500 & ~n28158 ;
  assign n28160 = \idma_PM_1st_reg/NET0131  & ~n20394 ;
  assign n28161 = ~\idma_PM_1st_reg/NET0131  & ~n20388 ;
  assign n28162 = n20822 & ~n28161 ;
  assign n28163 = ~n28160 & n28162 ;
  assign n28164 = ~n13570 & n28163 ;
  assign n28165 = ~n28159 & n28164 ;
  assign n28166 = \idma_DTMP_L_reg[7]/P0001  & ~n28163 ;
  assign n28167 = ~n28165 & ~n28166 ;
  assign n28168 = ~n27187 & n27499 ;
  assign n28169 = ~n27527 & ~n28168 ;
  assign n28170 = n28164 & ~n28169 ;
  assign n28171 = \idma_DTMP_L_reg[4]/P0001  & ~n28163 ;
  assign n28172 = ~n28170 & ~n28171 ;
  assign n28173 = ~n27215 & n27499 ;
  assign n28174 = ~n27536 & ~n28173 ;
  assign n28175 = n28164 & ~n28174 ;
  assign n28176 = \idma_DTMP_L_reg[3]/P0001  & ~n28163 ;
  assign n28177 = ~n28175 & ~n28176 ;
  assign n28178 = ~n27131 & n27499 ;
  assign n28179 = ~n27509 & ~n28178 ;
  assign n28180 = n28164 & ~n28179 ;
  assign n28181 = \idma_DTMP_L_reg[6]/P0001  & ~n28163 ;
  assign n28182 = ~n28180 & ~n28181 ;
  assign n28183 = ~n27243 & n27499 ;
  assign n28184 = ~n27545 & ~n28183 ;
  assign n28185 = n28164 & ~n28184 ;
  assign n28186 = \idma_DTMP_L_reg[2]/P0001  & ~n28163 ;
  assign n28187 = ~n28185 & ~n28186 ;
  assign n28188 = ~n27159 & n27499 ;
  assign n28189 = ~n27518 & ~n28188 ;
  assign n28190 = n28164 & ~n28189 ;
  assign n28191 = \idma_DTMP_L_reg[5]/P0001  & ~n28163 ;
  assign n28192 = ~n28190 & ~n28191 ;
  assign n28193 = ~n27271 & n27499 ;
  assign n28194 = ~n27554 & ~n28193 ;
  assign n28195 = n28164 & ~n28194 ;
  assign n28196 = \idma_DTMP_L_reg[1]/P0001  & ~n28163 ;
  assign n28197 = ~n28195 & ~n28196 ;
  assign n28198 = ~n27299 & n27499 ;
  assign n28199 = ~n27615 & ~n28198 ;
  assign n28200 = n28164 & ~n28199 ;
  assign n28201 = \idma_DTMP_L_reg[0]/P0001  & ~n28163 ;
  assign n28202 = ~n28200 & ~n28201 ;
  assign n28203 = n23027 & n25033 ;
  assign n28204 = n26967 & n28203 ;
  assign n28205 = ~\core_c_dec_IR_reg[9]/NET0131  & ~n28204 ;
  assign n28206 = ~\sice_SPC_reg[9]/P0001  & n28204 ;
  assign n28207 = ~n28205 & ~n28206 ;
  assign n28208 = n21242 & ~n28207 ;
  assign n28209 = ~n21242 & n27419 ;
  assign n28210 = ~n28208 & ~n28209 ;
  assign n28211 = ~\core_c_dec_IR_reg[8]/NET0131  & ~n28204 ;
  assign n28212 = ~\sice_SPC_reg[8]/P0001  & n28204 ;
  assign n28213 = ~n28211 & ~n28212 ;
  assign n28214 = n21242 & ~n28213 ;
  assign n28215 = ~n21242 & n27391 ;
  assign n28216 = ~n28214 & ~n28215 ;
  assign n28217 = ~\core_c_dec_IR_reg[7]/NET0131  & ~n28204 ;
  assign n28218 = ~\sice_SPC_reg[7]/P0001  & n28204 ;
  assign n28219 = ~n28217 & ~n28218 ;
  assign n28220 = n21242 & ~n28219 ;
  assign n28221 = ~n21242 & n27105 ;
  assign n28222 = ~n28220 & ~n28221 ;
  assign n28223 = ~\core_c_dec_IR_reg[6]/NET0131  & ~n28204 ;
  assign n28224 = ~\sice_SPC_reg[6]/P0001  & n28204 ;
  assign n28225 = ~n28223 & ~n28224 ;
  assign n28226 = n21242 & ~n28225 ;
  assign n28227 = ~n21242 & n27133 ;
  assign n28228 = ~n28226 & ~n28227 ;
  assign n28229 = ~\core_c_dec_IR_reg[5]/NET0131  & ~n28204 ;
  assign n28230 = ~\sice_SPC_reg[5]/P0001  & n28204 ;
  assign n28231 = ~n28229 & ~n28230 ;
  assign n28232 = n21242 & ~n28231 ;
  assign n28233 = ~n21242 & n27161 ;
  assign n28234 = ~n28232 & ~n28233 ;
  assign n28235 = ~\core_c_dec_IR_reg[4]/NET0131  & ~n28204 ;
  assign n28236 = ~\sice_SPC_reg[4]/P0001  & n28204 ;
  assign n28237 = ~n28235 & ~n28236 ;
  assign n28238 = n21242 & ~n28237 ;
  assign n28239 = ~n21242 & n27189 ;
  assign n28240 = ~n28238 & ~n28239 ;
  assign n28241 = ~\core_c_dec_IR_reg[3]/NET0131  & ~n28204 ;
  assign n28242 = ~\sice_SPC_reg[3]/P0001  & n28204 ;
  assign n28243 = ~n28241 & ~n28242 ;
  assign n28244 = n21242 & ~n28243 ;
  assign n28245 = ~n21242 & n27217 ;
  assign n28246 = ~n28244 & ~n28245 ;
  assign n28247 = ~\core_c_dec_IR_reg[2]/NET0131  & ~n28204 ;
  assign n28248 = ~\sice_SPC_reg[2]/P0001  & n28204 ;
  assign n28249 = ~n28247 & ~n28248 ;
  assign n28250 = n21242 & ~n28249 ;
  assign n28251 = ~n21242 & n27245 ;
  assign n28252 = ~n28250 & ~n28251 ;
  assign n28253 = ~\core_c_dec_IR_reg[23]/NET0131  & ~n28204 ;
  assign n28254 = ~\sice_SPC_reg[23]/P0001  & n28204 ;
  assign n28255 = ~n28253 & ~n28254 ;
  assign n28256 = n21242 & ~n28255 ;
  assign n28257 = \T_TMODE[1]_pad  & \emc_ECMDreg_reg[23]/P0001  ;
  assign n28258 = ~\T_TMODE[1]_pad  & ~n27577 ;
  assign n28259 = ~n28257 & ~n28258 ;
  assign n28260 = ~n21242 & n28259 ;
  assign n28261 = ~n28256 & ~n28260 ;
  assign n28262 = ~\core_c_dec_IR_reg[22]/NET0131  & ~n28204 ;
  assign n28263 = ~\sice_SPC_reg[22]/P0001  & n28204 ;
  assign n28264 = ~n28262 & ~n28263 ;
  assign n28265 = n21242 & ~n28264 ;
  assign n28266 = \T_TMODE[1]_pad  & \emc_ECMDreg_reg[22]/P0001  ;
  assign n28267 = ~\T_TMODE[1]_pad  & ~n27603 ;
  assign n28268 = ~n28266 & ~n28267 ;
  assign n28269 = ~n21242 & n28268 ;
  assign n28270 = ~n28265 & ~n28269 ;
  assign n28271 = ~\core_c_dec_IR_reg[21]/NET0131  & ~n28204 ;
  assign n28272 = ~\sice_SPC_reg[21]/P0001  & n28204 ;
  assign n28273 = ~n28271 & ~n28272 ;
  assign n28274 = n21242 & ~n28273 ;
  assign n28275 = \T_TMODE[1]_pad  & \emc_ECMDreg_reg[21]/P0001  ;
  assign n28276 = ~\T_TMODE[1]_pad  & ~n27695 ;
  assign n28277 = ~n28275 & ~n28276 ;
  assign n28278 = ~n21242 & n28277 ;
  assign n28279 = ~n28274 & ~n28278 ;
  assign n28280 = ~\core_c_dec_IR_reg[20]/NET0131  & ~n28204 ;
  assign n28281 = ~\sice_SPC_reg[20]/P0001  & n28204 ;
  assign n28282 = ~n28280 & ~n28281 ;
  assign n28283 = n21242 & ~n28282 ;
  assign n28284 = \T_TMODE[1]_pad  & \emc_ECMDreg_reg[20]/P0001  ;
  assign n28285 = ~\T_TMODE[1]_pad  & ~n27721 ;
  assign n28286 = ~n28284 & ~n28285 ;
  assign n28287 = ~n21242 & n28286 ;
  assign n28288 = ~n28283 & ~n28287 ;
  assign n28289 = ~\core_c_dec_IR_reg[19]/NET0131  & ~n28204 ;
  assign n28290 = ~\sice_SPC_reg[19]/P0001  & n28204 ;
  assign n28291 = ~n28289 & ~n28290 ;
  assign n28292 = n21242 & ~n28291 ;
  assign n28293 = \T_TMODE[1]_pad  & \emc_ECMDreg_reg[19]/P0001  ;
  assign n28294 = ~\T_TMODE[1]_pad  & ~n27747 ;
  assign n28295 = ~n28293 & ~n28294 ;
  assign n28296 = ~n21242 & n28295 ;
  assign n28297 = ~n28292 & ~n28296 ;
  assign n28298 = ~\core_c_dec_IR_reg[18]/NET0131  & ~n28204 ;
  assign n28299 = ~\sice_SPC_reg[18]/P0001  & n28204 ;
  assign n28300 = ~n28298 & ~n28299 ;
  assign n28301 = n21242 & ~n28300 ;
  assign n28302 = \T_TMODE[1]_pad  & \emc_ECMDreg_reg[18]/P0001  ;
  assign n28303 = ~\T_TMODE[1]_pad  & ~n27773 ;
  assign n28304 = ~n28302 & ~n28303 ;
  assign n28305 = ~n21242 & n28304 ;
  assign n28306 = ~n28301 & ~n28305 ;
  assign n28307 = ~\core_c_dec_IR_reg[17]/NET0131  & ~n28204 ;
  assign n28308 = ~\sice_SPC_reg[17]/P0001  & n28204 ;
  assign n28309 = ~n28307 & ~n28308 ;
  assign n28310 = n21242 & ~n28309 ;
  assign n28311 = \T_TMODE[1]_pad  & \emc_ECMDreg_reg[17]/P0001  ;
  assign n28312 = ~\T_TMODE[1]_pad  & ~n27643 ;
  assign n28313 = ~n28311 & ~n28312 ;
  assign n28314 = ~n21242 & n28313 ;
  assign n28315 = ~n28310 & ~n28314 ;
  assign n28316 = ~\core_c_dec_IR_reg[16]/NET0131  & ~n28204 ;
  assign n28317 = ~\sice_SPC_reg[16]/P0001  & n28204 ;
  assign n28318 = ~n28316 & ~n28317 ;
  assign n28319 = n21242 & ~n28318 ;
  assign n28320 = \T_TMODE[1]_pad  & \emc_ECMDreg_reg[16]/P0001  ;
  assign n28321 = ~\T_TMODE[1]_pad  & ~n27669 ;
  assign n28322 = ~n28320 & ~n28321 ;
  assign n28323 = ~n21242 & n28322 ;
  assign n28324 = ~n28319 & ~n28323 ;
  assign n28325 = ~\core_c_dec_IR_reg[15]/NET0131  & ~n28204 ;
  assign n28326 = ~\sice_SPC_reg[15]/P0001  & n28204 ;
  assign n28327 = ~n28325 & ~n28326 ;
  assign n28328 = n21242 & ~n28327 ;
  assign n28329 = ~n21242 & n27030 ;
  assign n28330 = ~n28328 & ~n28329 ;
  assign n28331 = ~\core_c_dec_IR_reg[14]/NET0131  & ~n28204 ;
  assign n28332 = ~\sice_SPC_reg[14]/P0001  & n28204 ;
  assign n28333 = ~n28331 & ~n28332 ;
  assign n28334 = n21242 & ~n28333 ;
  assign n28335 = ~n21242 & n27077 ;
  assign n28336 = ~n28334 & ~n28335 ;
  assign n28337 = ~\core_c_dec_IR_reg[13]/NET0131  & ~n28204 ;
  assign n28338 = ~\sice_SPC_reg[13]/P0001  & n28204 ;
  assign n28339 = ~n28337 & ~n28338 ;
  assign n28340 = n21242 & ~n28339 ;
  assign n28341 = ~n21242 & n27335 ;
  assign n28342 = ~n28340 & ~n28341 ;
  assign n28343 = ~\core_c_dec_IR_reg[12]/NET0131  & ~n28204 ;
  assign n28344 = ~\sice_SPC_reg[12]/P0001  & n28204 ;
  assign n28345 = ~n28343 & ~n28344 ;
  assign n28346 = n21242 & ~n28345 ;
  assign n28347 = ~n21242 & n27363 ;
  assign n28348 = ~n28346 & ~n28347 ;
  assign n28349 = ~\core_c_dec_IR_reg[11]/NET0131  & ~n28204 ;
  assign n28350 = ~\sice_SPC_reg[11]/P0001  & n28204 ;
  assign n28351 = ~n28349 & ~n28350 ;
  assign n28352 = n21242 & ~n28351 ;
  assign n28353 = ~n21242 & n27447 ;
  assign n28354 = ~n28352 & ~n28353 ;
  assign n28355 = ~\core_c_dec_IR_reg[10]/NET0131  & ~n28204 ;
  assign n28356 = ~\sice_SPC_reg[10]/P0001  & n28204 ;
  assign n28357 = ~n28355 & ~n28356 ;
  assign n28358 = n21242 & ~n28357 ;
  assign n28359 = ~n21242 & n27475 ;
  assign n28360 = ~n28358 & ~n28359 ;
  assign n28361 = \sice_SPC_reg[21]/P0001  & n26969 ;
  assign n28362 = \core_c_dec_rdCM_E_reg/NET0131  & ~n28277 ;
  assign n28363 = ~n28361 & ~n28362 ;
  assign n28364 = \sice_SPC_reg[20]/P0001  & n26969 ;
  assign n28365 = \core_c_dec_rdCM_E_reg/NET0131  & ~n28286 ;
  assign n28366 = ~n28364 & ~n28365 ;
  assign n28367 = \sice_SPC_reg[19]/P0001  & n26969 ;
  assign n28368 = \core_c_dec_rdCM_E_reg/NET0131  & ~n28295 ;
  assign n28369 = ~n28367 & ~n28368 ;
  assign n28370 = \sice_SPC_reg[18]/P0001  & n26969 ;
  assign n28371 = \core_c_dec_rdCM_E_reg/NET0131  & ~n28304 ;
  assign n28372 = ~n28370 & ~n28371 ;
  assign n28373 = \sice_SPC_reg[17]/P0001  & n26969 ;
  assign n28374 = \core_c_dec_rdCM_E_reg/NET0131  & ~n28313 ;
  assign n28375 = ~n28373 & ~n28374 ;
  assign n28376 = \sice_SPC_reg[16]/P0001  & n26969 ;
  assign n28377 = \core_c_dec_rdCM_E_reg/NET0131  & ~n28322 ;
  assign n28378 = ~n28376 & ~n28377 ;
  assign n28379 = \sice_SPC_reg[23]/P0001  & n26969 ;
  assign n28380 = \core_c_dec_rdCM_E_reg/NET0131  & ~n28259 ;
  assign n28381 = ~n28379 & ~n28380 ;
  assign n28382 = \sice_SPC_reg[22]/P0001  & n26969 ;
  assign n28383 = \core_c_dec_rdCM_E_reg/NET0131  & ~n28268 ;
  assign n28384 = ~n28382 & ~n28383 ;
  assign n28385 = ~\auctl_BSack_reg/NET0131  & \bdma_BWdataBUF_h_reg[8]/P0001  ;
  assign n28386 = n6921 & n10638 ;
  assign n28387 = n12520 & n13152 ;
  assign n28388 = ~n5727 & n13151 ;
  assign n28389 = ~n27389 & n28388 ;
  assign n28390 = ~n28387 & ~n28389 ;
  assign n28391 = ~n28386 & n28390 ;
  assign n28392 = \auctl_BSack_reg/NET0131  & ~n28391 ;
  assign n28393 = ~n28385 & ~n28392 ;
  assign n28394 = ~\auctl_BSack_reg/NET0131  & \bdma_BWdataBUF_h_reg[9]/P0001  ;
  assign n28395 = n6921 & n10289 ;
  assign n28396 = n12802 & n13152 ;
  assign n28397 = ~n27417 & n28388 ;
  assign n28398 = ~n28396 & ~n28397 ;
  assign n28399 = ~n28395 & n28398 ;
  assign n28400 = \auctl_BSack_reg/NET0131  & ~n28399 ;
  assign n28401 = ~n28394 & ~n28400 ;
  assign n28402 = ~\auctl_BSack_reg/NET0131  & \bdma_BWdataBUF_h_reg[15]/P0001  ;
  assign n28403 = n6921 & n12743 ;
  assign n28404 = n13006 & n13152 ;
  assign n28405 = ~n27028 & n28388 ;
  assign n28406 = ~n28404 & ~n28405 ;
  assign n28407 = ~n28403 & n28406 ;
  assign n28408 = \auctl_BSack_reg/NET0131  & ~n28407 ;
  assign n28409 = ~n28402 & ~n28408 ;
  assign n28410 = ~\auctl_BSack_reg/NET0131  & \bdma_BWdataBUF_h_reg[14]/P0001  ;
  assign n28413 = n12972 & n13152 ;
  assign n28411 = n6921 & n12688 ;
  assign n28412 = ~n27075 & n28388 ;
  assign n28414 = ~n28411 & ~n28412 ;
  assign n28415 = ~n28413 & n28414 ;
  assign n28416 = \auctl_BSack_reg/NET0131  & ~n28415 ;
  assign n28417 = ~n28410 & ~n28416 ;
  assign n28418 = ~\auctl_BSack_reg/NET0131  & \bdma_BWdataBUF_h_reg[13]/P0001  ;
  assign n28419 = n6921 & n7340 ;
  assign n28420 = n12938 & n13152 ;
  assign n28421 = ~n27333 & n28388 ;
  assign n28422 = ~n28420 & ~n28421 ;
  assign n28423 = ~n28419 & n28422 ;
  assign n28424 = \auctl_BSack_reg/NET0131  & ~n28423 ;
  assign n28425 = ~n28418 & ~n28424 ;
  assign n28426 = ~\auctl_BSack_reg/NET0131  & \bdma_BWdataBUF_h_reg[12]/P0001  ;
  assign n28427 = n6921 & n9178 ;
  assign n28428 = n12904 & n13152 ;
  assign n28429 = ~n27361 & n28388 ;
  assign n28430 = ~n28428 & ~n28429 ;
  assign n28431 = ~n28427 & n28430 ;
  assign n28432 = \auctl_BSack_reg/NET0131  & ~n28431 ;
  assign n28433 = ~n28426 & ~n28432 ;
  assign n28434 = ~\auctl_BSack_reg/NET0131  & \bdma_BWdataBUF_h_reg[11]/P0001  ;
  assign n28435 = n6921 & n8460 ;
  assign n28436 = n12870 & n13152 ;
  assign n28437 = ~n27445 & n28388 ;
  assign n28438 = ~n28436 & ~n28437 ;
  assign n28439 = ~n28435 & n28438 ;
  assign n28440 = \auctl_BSack_reg/NET0131  & ~n28439 ;
  assign n28441 = ~n28434 & ~n28440 ;
  assign n28442 = ~\auctl_BSack_reg/NET0131  & \bdma_BWdataBUF_h_reg[10]/P0001  ;
  assign n28443 = n6921 & n7859 ;
  assign n28444 = n12836 & n13152 ;
  assign n28445 = ~n27473 & n28388 ;
  assign n28446 = ~n28444 & ~n28445 ;
  assign n28447 = ~n28443 & n28446 ;
  assign n28448 = \auctl_BSack_reg/NET0131  & ~n28447 ;
  assign n28449 = ~n28442 & ~n28448 ;
  assign n28450 = ~\core_c_dec_IR_reg[1]/NET0131  & ~n28204 ;
  assign n28451 = ~\sice_SPC_reg[1]/P0001  & n28204 ;
  assign n28452 = ~n28450 & ~n28451 ;
  assign n28453 = n21242 & ~n28452 ;
  assign n28454 = ~n21242 & n27273 ;
  assign n28455 = ~n28453 & ~n28454 ;
  assign n28456 = ~\core_c_dec_IR_reg[0]/NET0131  & ~n28204 ;
  assign n28457 = ~\sice_SPC_reg[0]/P0001  & n28204 ;
  assign n28458 = ~n28456 & ~n28457 ;
  assign n28459 = n21242 & ~n28458 ;
  assign n28460 = ~n21242 & n27301 ;
  assign n28461 = ~n28459 & ~n28460 ;
  assign n28462 = ~\auctl_BSack_reg/NET0131  & \bdma_BWdataBUF_h_reg[7]/P0001  ;
  assign n28463 = n6921 & n11265 ;
  assign n28464 = ~n27103 & n28388 ;
  assign n28465 = ~n28463 & ~n28464 ;
  assign n28466 = \auctl_BSack_reg/NET0131  & ~n28465 ;
  assign n28467 = ~n28462 & ~n28466 ;
  assign n28468 = ~\auctl_BSack_reg/NET0131  & \bdma_BWdataBUF_h_reg[6]/P0001  ;
  assign n28469 = n6921 & n11525 ;
  assign n28470 = ~n27131 & n28388 ;
  assign n28471 = ~n28469 & ~n28470 ;
  assign n28472 = \auctl_BSack_reg/NET0131  & ~n28471 ;
  assign n28473 = ~n28468 & ~n28472 ;
  assign n28474 = ~\auctl_BSack_reg/NET0131  & \bdma_BWdataBUF_h_reg[5]/P0001  ;
  assign n28475 = n6921 & n10911 ;
  assign n28476 = ~n27159 & n28388 ;
  assign n28477 = ~n28475 & ~n28476 ;
  assign n28478 = \auctl_BSack_reg/NET0131  & ~n28477 ;
  assign n28479 = ~n28474 & ~n28478 ;
  assign n28480 = ~\auctl_BSack_reg/NET0131  & \bdma_BWdataBUF_h_reg[4]/P0001  ;
  assign n28481 = n6921 & n10069 ;
  assign n28482 = ~n27187 & n28388 ;
  assign n28483 = ~n28481 & ~n28482 ;
  assign n28484 = \auctl_BSack_reg/NET0131  & ~n28483 ;
  assign n28485 = ~n28480 & ~n28484 ;
  assign n28486 = ~\auctl_BSack_reg/NET0131  & \bdma_BWdataBUF_h_reg[3]/P0001  ;
  assign n28487 = n6921 & n8113 ;
  assign n28488 = ~n27215 & n28388 ;
  assign n28489 = ~n28487 & ~n28488 ;
  assign n28490 = \auctl_BSack_reg/NET0131  & ~n28489 ;
  assign n28491 = ~n28486 & ~n28490 ;
  assign n28492 = ~\auctl_BSack_reg/NET0131  & \bdma_BWdataBUF_h_reg[2]/P0001  ;
  assign n28493 = n6921 & n8715 ;
  assign n28494 = ~n27243 & n28388 ;
  assign n28495 = ~n28493 & ~n28494 ;
  assign n28496 = \auctl_BSack_reg/NET0131  & ~n28495 ;
  assign n28497 = ~n28492 & ~n28496 ;
  assign n28498 = ~\auctl_BSack_reg/NET0131  & \bdma_BWdataBUF_h_reg[23]/P0001  ;
  assign n28499 = n12771 & n13152 ;
  assign n28500 = ~n27577 & n28388 ;
  assign n28501 = ~n28499 & ~n28500 ;
  assign n28502 = \auctl_BSack_reg/NET0131  & ~n28501 ;
  assign n28503 = ~n28498 & ~n28502 ;
  assign n28504 = ~\auctl_BSack_reg/NET0131  & \bdma_BWdataBUF_h_reg[22]/P0001  ;
  assign n28505 = n12715 & n13152 ;
  assign n28506 = ~n27603 & n28388 ;
  assign n28507 = ~n28505 & ~n28506 ;
  assign n28508 = \auctl_BSack_reg/NET0131  & ~n28507 ;
  assign n28509 = ~n28504 & ~n28508 ;
  assign n28510 = ~\auctl_BSack_reg/NET0131  & \bdma_BWdataBUF_h_reg[21]/P0001  ;
  assign n28511 = n12658 & n13152 ;
  assign n28512 = ~n27695 & n28388 ;
  assign n28513 = ~n28511 & ~n28512 ;
  assign n28514 = \auctl_BSack_reg/NET0131  & ~n28513 ;
  assign n28515 = ~n28510 & ~n28514 ;
  assign n28516 = ~\auctl_BSack_reg/NET0131  & \bdma_BWdataBUF_h_reg[20]/P0001  ;
  assign n28517 = n12624 & n13152 ;
  assign n28518 = ~n27721 & n28388 ;
  assign n28519 = ~n28517 & ~n28518 ;
  assign n28520 = \auctl_BSack_reg/NET0131  & ~n28519 ;
  assign n28521 = ~n28516 & ~n28520 ;
  assign n28522 = ~\auctl_BSack_reg/NET0131  & \bdma_BWdataBUF_h_reg[1]/P0001  ;
  assign n28523 = n6921 & n9435 ;
  assign n28524 = ~n27271 & n28388 ;
  assign n28525 = ~n28523 & ~n28524 ;
  assign n28526 = \auctl_BSack_reg/NET0131  & ~n28525 ;
  assign n28527 = ~n28522 & ~n28526 ;
  assign n28528 = n18262 & n19409 ;
  assign n28529 = ~n18262 & ~n19384 ;
  assign n28530 = n14664 & n17801 ;
  assign n28531 = ~\core_eu_em_mac_em_reg_mr2swe_DO_reg[1]/P0001  & ~n28530 ;
  assign n28532 = \core_c_psq_MSTAT_reg_DO_reg[0]/P0002  & ~n17807 ;
  assign n28533 = ~n19381 & ~n28530 ;
  assign n28534 = n28532 & ~n28533 ;
  assign n28535 = n18974 & ~n19381 ;
  assign n28536 = n28534 & ~n28535 ;
  assign n28537 = ~n28531 & ~n28536 ;
  assign n28538 = ~n19385 & ~n28537 ;
  assign n28539 = ~\core_eu_em_mac_em_reg_mr2swe_DO_reg[1]/P0001  & ~n28532 ;
  assign n28540 = ~n28538 & ~n28539 ;
  assign n28541 = n28529 & ~n28540 ;
  assign n28542 = ~n28528 & ~n28541 ;
  assign n28543 = ~\core_c_dec_MACop_E_reg/P0001  & ~n18847 ;
  assign n28544 = n4117 & ~n5689 ;
  assign n28545 = ~n28543 & ~n28544 ;
  assign n28546 = n5689 & ~n13832 ;
  assign n28547 = ~\core_c_dec_IR_reg[10]/NET0131  & ~\core_c_dec_IR_reg[9]/NET0131  ;
  assign n28548 = ~n5689 & ~n28547 ;
  assign n28549 = ~n28546 & ~n28548 ;
  assign n28550 = n28545 & ~n28549 ;
  assign n28558 = ~n5689 & n26353 ;
  assign n28559 = n26370 & n28558 ;
  assign n28561 = ~\core_c_dec_MTAR_E_reg/P0001  & ~n19214 ;
  assign n28562 = ~n14586 & n28561 ;
  assign n28560 = \core_c_dec_MTAR_E_reg/P0001  & n17814 ;
  assign n28563 = ~\core_c_dec_MTAR_E_reg/P0001  & ~n19278 ;
  assign n28564 = n19214 & n28563 ;
  assign n28565 = ~n28560 & ~n28564 ;
  assign n28566 = ~n28562 & n28565 ;
  assign n28567 = n28559 & ~n28566 ;
  assign n28568 = \core_eu_em_mac_em_reg_s2_reg/P0000_reg_syn_2  & n26395 ;
  assign n28569 = ~n26388 & ~n28568 ;
  assign n28570 = ~n26396 & n26966 ;
  assign n28571 = ~\core_eu_em_mac_em_reg_s0_reg/P0000_reg_syn_2  & n26396 ;
  assign n28572 = ~n28570 & ~n28571 ;
  assign n28573 = \core_eu_em_mac_em_reg_s1_reg/P0000_reg_syn_2  & n26396 ;
  assign n28574 = n26394 & ~n28573 ;
  assign n28575 = ~n28572 & ~n28574 ;
  assign n28576 = n17820 & n28575 ;
  assign n28577 = n28572 & n28574 ;
  assign n28579 = ~n8715 & n28577 ;
  assign n28578 = ~n12836 & ~n28577 ;
  assign n28580 = ~n28575 & ~n28578 ;
  assign n28581 = ~n28579 & n28580 ;
  assign n28582 = ~n28576 & ~n28581 ;
  assign n28583 = n28569 & ~n28582 ;
  assign n28600 = n17804 & n26370 ;
  assign n28601 = n7206 & n28600 ;
  assign n28586 = ~\core_c_dec_IR_reg[8]/NET0131  & n26379 ;
  assign n28592 = ~n5689 & n26371 ;
  assign n28602 = ~n28586 & ~n28592 ;
  assign n28603 = n28601 & ~n28602 ;
  assign n28604 = ~n7206 & n26379 ;
  assign n28605 = n28600 & n28604 ;
  assign n28606 = \core_c_dec_IR_reg[8]/NET0131  & n28605 ;
  assign n28607 = ~n28603 & ~n28606 ;
  assign n28596 = ~n26370 & n26380 ;
  assign n28597 = n5689 & n13813 ;
  assign n28598 = ~n28596 & ~n28597 ;
  assign n28599 = ~n8534 & ~n28598 ;
  assign n28587 = ~n26370 & n28586 ;
  assign n28588 = n5689 & n13821 ;
  assign n28589 = ~n28587 & ~n28588 ;
  assign n28590 = ~n8558 & ~n28589 ;
  assign n28591 = n5689 & n13819 ;
  assign n28593 = ~n26370 & n28592 ;
  assign n28594 = ~n28591 & ~n28593 ;
  assign n28595 = ~n8554 & ~n28594 ;
  assign n28608 = ~n28590 & ~n28595 ;
  assign n28609 = ~n28599 & n28608 ;
  assign n28610 = n28607 & n28609 ;
  assign n28611 = n28572 & n28610 ;
  assign n28584 = ~n28569 & n28574 ;
  assign n28585 = ~n8715 & ~n28572 ;
  assign n28612 = n28584 & ~n28585 ;
  assign n28613 = ~n28611 & n28612 ;
  assign n28615 = \core_c_dec_IR_reg[8]/NET0131  & ~\core_c_dec_MTSR1_E_reg/P0001  ;
  assign n28553 = ~n5689 & n26356 ;
  assign n28626 = n26370 & n28553 ;
  assign n28627 = n28615 & n28626 ;
  assign n28628 = ~n21124 & n28627 ;
  assign n28632 = n5689 & n13816 ;
  assign n28633 = ~n26370 & n28558 ;
  assign n28634 = ~n28632 & ~n28633 ;
  assign n28635 = ~n8585 & ~n28634 ;
  assign n28614 = ~\core_c_dec_IR_reg[8]/NET0131  & ~\core_c_dec_MTSR0_E_reg/P0001  ;
  assign n28616 = ~n28614 & ~n28615 ;
  assign n28617 = n26370 & n28616 ;
  assign n28618 = \core_c_dec_accPM_E_reg/P0001  & n28553 ;
  assign n28619 = n28617 & n28618 ;
  assign n28620 = n12836 & n28619 ;
  assign n28629 = ~\core_c_dec_accPM_E_reg/P0001  & n28553 ;
  assign n28630 = n28617 & n28629 ;
  assign n28631 = n8715 & n28630 ;
  assign n28638 = ~n28620 & ~n28631 ;
  assign n28639 = ~n28635 & n28638 ;
  assign n28636 = n28614 & n28626 ;
  assign n28637 = ~n21174 & n28636 ;
  assign n28551 = \core_c_dec_IRE_reg[8]/NET0131  & n5689 ;
  assign n28552 = n13823 & n28551 ;
  assign n28554 = ~n26370 & n28553 ;
  assign n28555 = \core_c_dec_IR_reg[8]/NET0131  & n28554 ;
  assign n28556 = ~n28552 & ~n28555 ;
  assign n28557 = ~n8497 & ~n28556 ;
  assign n28621 = ~\core_c_dec_IR_reg[8]/NET0131  & n28554 ;
  assign n28622 = ~\core_c_dec_IRE_reg[8]/NET0131  & n13823 ;
  assign n28623 = n5689 & n28622 ;
  assign n28624 = ~n28621 & ~n28623 ;
  assign n28625 = ~n8493 & ~n28624 ;
  assign n28640 = ~n28557 & ~n28625 ;
  assign n28641 = ~n28637 & n28640 ;
  assign n28642 = n28639 & n28641 ;
  assign n28643 = ~n28628 & n28642 ;
  assign n28644 = ~n28613 & n28643 ;
  assign n28645 = ~n28583 & n28644 ;
  assign n28646 = ~n28567 & n28645 ;
  assign n28647 = n28550 & ~n28646 ;
  assign n28655 = ~n5689 & n18847 ;
  assign n28657 = ~\core_c_dec_Dummy_E_reg/NET0131  & n28547 ;
  assign n28654 = \core_c_dec_IR_reg[8]/NET0131  & ~\core_c_dec_MTMX1_E_reg/P0001  ;
  assign n28656 = ~\core_c_dec_IR_reg[8]/NET0131  & ~\core_c_dec_MTMX0_E_reg/P0001  ;
  assign n28658 = ~n28654 & ~n28656 ;
  assign n28659 = n28657 & n28658 ;
  assign n28660 = n28655 & n28659 ;
  assign n28664 = n17814 & n28660 ;
  assign n28648 = \core_c_dec_MACop_E_reg/P0001  & n5689 ;
  assign n28649 = ~n18848 & ~n28648 ;
  assign n28651 = \core_c_dec_IR_reg[8]/NET0131  & ~n5689 ;
  assign n28652 = ~n28551 & ~n28651 ;
  assign n28661 = n8538 & ~n28652 ;
  assign n28653 = n8550 & n28652 ;
  assign n28662 = ~n28653 & ~n28660 ;
  assign n28663 = ~n28661 & n28662 ;
  assign n28665 = ~n28649 & ~n28663 ;
  assign n28666 = ~n28664 & n28665 ;
  assign n28650 = ~\core_eu_em_mac_em_reg_mxopwe_DO_reg[2]/P0001  & n28649 ;
  assign n28667 = ~n28550 & ~n28650 ;
  assign n28668 = ~n28666 & n28667 ;
  assign n28669 = ~n28647 & ~n28668 ;
  assign n28670 = ~\auctl_BSack_reg/NET0131  & \bdma_BWdataBUF_h_reg[19]/P0001  ;
  assign n28671 = n12590 & n13152 ;
  assign n28672 = ~n27747 & n28388 ;
  assign n28673 = ~n28671 & ~n28672 ;
  assign n28674 = \auctl_BSack_reg/NET0131  & ~n28673 ;
  assign n28675 = ~n28670 & ~n28674 ;
  assign n28676 = ~\auctl_BSack_reg/NET0131  & \bdma_BWdataBUF_h_reg[18]/P0001  ;
  assign n28677 = n12556 & n13152 ;
  assign n28678 = ~n27773 & n28388 ;
  assign n28679 = ~n28677 & ~n28678 ;
  assign n28680 = \auctl_BSack_reg/NET0131  & ~n28679 ;
  assign n28681 = ~n28676 & ~n28680 ;
  assign n28682 = ~\auctl_BSack_reg/NET0131  & \bdma_BWdataBUF_h_reg[17]/P0001  ;
  assign n28683 = n13075 & n13152 ;
  assign n28684 = ~n27643 & n28388 ;
  assign n28685 = ~n28683 & ~n28684 ;
  assign n28686 = \auctl_BSack_reg/NET0131  & ~n28685 ;
  assign n28687 = ~n28682 & ~n28686 ;
  assign n28688 = ~\auctl_BSack_reg/NET0131  & \bdma_BWdataBUF_h_reg[16]/P0001  ;
  assign n28689 = n13041 & n13152 ;
  assign n28690 = ~n27669 & n28388 ;
  assign n28691 = ~n28689 & ~n28690 ;
  assign n28692 = \auctl_BSack_reg/NET0131  & ~n28691 ;
  assign n28693 = ~n28688 & ~n28692 ;
  assign n28694 = ~\auctl_BSack_reg/NET0131  & \bdma_BWdataBUF_h_reg[0]/P0001  ;
  assign n28695 = n6921 & n7607 ;
  assign n28696 = ~n27299 & n28388 ;
  assign n28697 = ~n28695 & ~n28696 ;
  assign n28698 = \auctl_BSack_reg/NET0131  & ~n28697 ;
  assign n28699 = ~n28694 & ~n28698 ;
  assign n28700 = \core_c_dec_IR_reg[12]/NET0131  & ~n5689 ;
  assign n28701 = \core_c_dec_IRE_reg[12]/NET0131  & n5689 ;
  assign n28702 = ~n28700 & ~n28701 ;
  assign n28703 = \core_c_dec_IR_reg[11]/NET0131  & ~n5689 ;
  assign n28704 = \core_c_dec_IRE_reg[11]/NET0131  & n5689 ;
  assign n28705 = ~n28703 & ~n28704 ;
  assign n28706 = ~n28702 & ~n28705 ;
  assign n28708 = \core_c_dec_IR_reg[11]/NET0131  & ~\core_c_dec_MTMY1_E_reg/P0001  ;
  assign n28707 = ~\core_c_dec_IR_reg[11]/NET0131  & ~\core_c_dec_MTMY0_E_reg/P0001  ;
  assign n28709 = ~\core_c_dec_Dummy_E_reg/NET0131  & ~\core_c_dec_IR_reg[12]/NET0131  ;
  assign n28710 = ~n28707 & n28709 ;
  assign n28711 = ~n28708 & n28710 ;
  assign n28712 = ~n26358 & n28711 ;
  assign n28713 = n28655 & n28712 ;
  assign n28714 = ~n28706 & ~n28713 ;
  assign n28715 = ~n5689 & ~n21525 ;
  assign n28716 = ~\core_eu_em_mac_em_reg_Sq_E_reg/P0001  & n5689 ;
  assign n28717 = ~n28715 & ~n28716 ;
  assign n28718 = n28714 & n28717 ;
  assign n28719 = n28550 & n28718 ;
  assign n28720 = ~n28544 & n28718 ;
  assign n28721 = n28660 & n28720 ;
  assign n28722 = ~n4117 & n28713 ;
  assign n28723 = ~\core_c_dec_Double_E_reg/P0001  & n28722 ;
  assign n28724 = ~n28721 & ~n28723 ;
  assign n28725 = ~\core_c_dec_accPM_E_reg/P0001  & ~n28724 ;
  assign n28731 = n8715 & n28725 ;
  assign n28726 = \core_c_dec_accPM_E_reg/P0001  & n28721 ;
  assign n28727 = ~n21991 & n28722 ;
  assign n28728 = ~n28726 & ~n28727 ;
  assign n28729 = ~n28725 & ~n28728 ;
  assign n28730 = n12836 & n28729 ;
  assign n28733 = ~n28544 & ~n28717 ;
  assign n28734 = n28714 & n28733 ;
  assign n28741 = ~n28702 & n28734 ;
  assign n28742 = ~\core_c_psq_MSTAT_reg_DO_reg[0]/P0002  & ~\core_eu_em_mac_em_reg_mfrwe_DO_reg[2]/P0001  ;
  assign n28743 = \core_c_psq_MSTAT_reg_DO_reg[0]/P0002  & ~\core_eu_em_mac_em_reg_mfswe_DO_reg[2]/P0001  ;
  assign n28744 = ~n28742 & ~n28743 ;
  assign n28745 = n28741 & n28744 ;
  assign n28735 = n28702 & n28734 ;
  assign n28732 = n8546 & n28705 ;
  assign n28736 = n8542 & ~n28705 ;
  assign n28737 = ~n28732 & ~n28736 ;
  assign n28738 = n28735 & n28737 ;
  assign n28739 = n28549 & n28720 ;
  assign n28740 = n28663 & n28739 ;
  assign n28746 = ~n28738 & ~n28740 ;
  assign n28747 = ~n28745 & n28746 ;
  assign n28748 = ~n28730 & n28747 ;
  assign n28749 = ~n28731 & n28748 ;
  assign n28750 = ~n28543 & ~n28749 ;
  assign n28751 = \core_eu_em_mac_em_reg_myopwe_DO_reg[2]/P0001  & ~n28545 ;
  assign n28752 = ~n28750 & ~n28751 ;
  assign n28753 = ~n28719 & ~n28752 ;
  assign n28754 = ~n28646 & n28719 ;
  assign n28755 = ~n28753 & ~n28754 ;
  assign n28756 = \tm_tcr_reg_DO_reg[14]/NET0131  & n20355 ;
  assign n28758 = \tm_TCR_TMP_reg[14]/NET0131  & ~n25841 ;
  assign n28759 = ~n22400 & ~n25842 ;
  assign n28760 = ~n28758 & n28759 ;
  assign n28757 = ~\tm_tpr_reg_DO_reg[14]/NET0131  & n22400 ;
  assign n28761 = ~n20355 & ~n28757 ;
  assign n28762 = ~n28760 & n28761 ;
  assign n28763 = ~n28756 & ~n28762 ;
  assign n28764 = n14752 & n19409 ;
  assign n28765 = ~\core_eu_em_mac_em_reg_mr2rwe_DO_reg[1]/P0001  & ~n17799 ;
  assign n28766 = ~n17809 & n18974 ;
  assign n28767 = n17811 & ~n28766 ;
  assign n28768 = ~n28765 & ~n28767 ;
  assign n28769 = ~n17823 & ~n28768 ;
  assign n28770 = ~\core_eu_em_mac_em_reg_mr2rwe_DO_reg[1]/P0001  & ~n17808 ;
  assign n28771 = ~n28769 & ~n28770 ;
  assign n28772 = n17829 & ~n28771 ;
  assign n28773 = ~n28764 & ~n28772 ;
  assign n28775 = \sport0_regs_SCTLreg_DO_reg[5]/NET0131  & ~n20953 ;
  assign n28774 = ~\sport0_regs_SCTLreg_DO_reg[5]/NET0131  & \sport0_rxctl_RX_reg[0]/P0001  ;
  assign n28776 = \sport0_rxctl_ldRX_cmp_reg/P0001  & ~n28774 ;
  assign n28777 = ~n28775 & n28776 ;
  assign n28778 = n7607 & n20869 ;
  assign n28779 = \sport0_rxctl_RX_reg[0]/P0001  & ~n20869 ;
  assign n28780 = ~\sport0_rxctl_ldRX_cmp_reg/P0001  & ~n28779 ;
  assign n28781 = ~n28778 & n28780 ;
  assign n28782 = ~n28777 & ~n28781 ;
  assign n28783 = ~n20868 & ~n28782 ;
  assign n28784 = ~\sport0_rxctl_RXSHT_reg[0]/P0001  & n20868 ;
  assign n28785 = ~n28783 & ~n28784 ;
  assign n28786 = ~\sport1_cfg_SP_ENg_D1_reg/P0001  & \sport1_cfg_SP_ENg_reg/NET0131  ;
  assign n28787 = \sport1_regs_FSDIVreg_DO_reg[15]/NET0131  & n28786 ;
  assign n28856 = \sport1_cfg_FSi_cnt_reg[0]/NET0131  & \sport1_cfg_SP_ENg_reg/NET0131  ;
  assign n28857 = \sport1_cfg_FSi_cnt_reg[1]/NET0131  & n28856 ;
  assign n28858 = \sport1_cfg_FSi_cnt_reg[2]/NET0131  & n28857 ;
  assign n28859 = \sport1_cfg_FSi_cnt_reg[3]/NET0131  & n28858 ;
  assign n28860 = \sport1_cfg_FSi_cnt_reg[4]/NET0131  & n28859 ;
  assign n28861 = \sport1_cfg_FSi_cnt_reg[5]/NET0131  & n28860 ;
  assign n28862 = \sport1_cfg_FSi_cnt_reg[6]/NET0131  & n28861 ;
  assign n28863 = \sport1_cfg_FSi_cnt_reg[7]/NET0131  & n28862 ;
  assign n28864 = \sport1_cfg_FSi_cnt_reg[8]/NET0131  & n28863 ;
  assign n28865 = \sport1_cfg_FSi_cnt_reg[9]/NET0131  & n28864 ;
  assign n28866 = \sport1_cfg_FSi_cnt_reg[10]/NET0131  & n28865 ;
  assign n28867 = \sport1_cfg_FSi_cnt_reg[11]/NET0131  & n28866 ;
  assign n28868 = \sport1_cfg_FSi_cnt_reg[12]/NET0131  & n28867 ;
  assign n28869 = \sport1_cfg_FSi_cnt_reg[13]/NET0131  & n28868 ;
  assign n28870 = \sport1_cfg_FSi_cnt_reg[14]/NET0131  & n28869 ;
  assign n28872 = \sport1_cfg_FSi_cnt_reg[15]/NET0131  & n28870 ;
  assign n28788 = ~\IRFS1_pad  & ~\ITFS1_pad  ;
  assign n28809 = \sport1_cfg_FSi_cnt_reg[11]/NET0131  & ~\sport1_regs_FSDIVreg_DO_reg[11]/NET0131  ;
  assign n28810 = \sport1_cfg_FSi_cnt_reg[14]/NET0131  & ~\sport1_regs_FSDIVreg_DO_reg[14]/NET0131  ;
  assign n28831 = ~n28809 & ~n28810 ;
  assign n28811 = ~\sport1_cfg_FSi_cnt_reg[9]/NET0131  & \sport1_regs_FSDIVreg_DO_reg[9]/NET0131  ;
  assign n28812 = \sport1_cfg_FSi_cnt_reg[2]/NET0131  & ~\sport1_regs_FSDIVreg_DO_reg[2]/NET0131  ;
  assign n28832 = ~n28811 & ~n28812 ;
  assign n28839 = n28831 & n28832 ;
  assign n28805 = \sport1_cfg_FSi_cnt_reg[1]/NET0131  & ~\sport1_regs_FSDIVreg_DO_reg[1]/NET0131  ;
  assign n28806 = \sport1_cfg_FSi_cnt_reg[7]/NET0131  & ~\sport1_regs_FSDIVreg_DO_reg[7]/NET0131  ;
  assign n28829 = ~n28805 & ~n28806 ;
  assign n28807 = \sport1_cfg_FSi_cnt_reg[3]/NET0131  & ~\sport1_regs_FSDIVreg_DO_reg[3]/NET0131  ;
  assign n28808 = \sport1_cfg_FSi_cnt_reg[9]/NET0131  & ~\sport1_regs_FSDIVreg_DO_reg[9]/NET0131  ;
  assign n28830 = ~n28807 & ~n28808 ;
  assign n28840 = n28829 & n28830 ;
  assign n28847 = n28839 & n28840 ;
  assign n28817 = \sport1_cfg_FSi_cnt_reg[13]/NET0131  & ~\sport1_regs_FSDIVreg_DO_reg[13]/NET0131  ;
  assign n28818 = ~\sport1_cfg_FSi_cnt_reg[15]/NET0131  & \sport1_regs_FSDIVreg_DO_reg[15]/NET0131  ;
  assign n28835 = ~n28817 & ~n28818 ;
  assign n28819 = \sport1_cfg_FSi_cnt_reg[12]/NET0131  & ~\sport1_regs_FSDIVreg_DO_reg[12]/NET0131  ;
  assign n28820 = ~\sport1_cfg_FSi_cnt_reg[6]/NET0131  & \sport1_regs_FSDIVreg_DO_reg[6]/NET0131  ;
  assign n28836 = ~n28819 & ~n28820 ;
  assign n28837 = n28835 & n28836 ;
  assign n28813 = ~\sport1_cfg_FSi_cnt_reg[7]/NET0131  & \sport1_regs_FSDIVreg_DO_reg[7]/NET0131  ;
  assign n28814 = ~\sport1_cfg_FSi_cnt_reg[14]/NET0131  & \sport1_regs_FSDIVreg_DO_reg[14]/NET0131  ;
  assign n28833 = ~n28813 & ~n28814 ;
  assign n28815 = ~\sport1_cfg_FSi_cnt_reg[13]/NET0131  & \sport1_regs_FSDIVreg_DO_reg[13]/NET0131  ;
  assign n28816 = \sport1_cfg_FSi_cnt_reg[6]/NET0131  & ~\sport1_regs_FSDIVreg_DO_reg[6]/NET0131  ;
  assign n28834 = ~n28815 & ~n28816 ;
  assign n28838 = n28833 & n28834 ;
  assign n28848 = n28837 & n28838 ;
  assign n28849 = n28847 & n28848 ;
  assign n28793 = \sport1_cfg_FSi_cnt_reg[5]/NET0131  & ~\sport1_regs_FSDIVreg_DO_reg[5]/NET0131  ;
  assign n28794 = ~\sport1_cfg_FSi_cnt_reg[8]/NET0131  & \sport1_regs_FSDIVreg_DO_reg[8]/NET0131  ;
  assign n28823 = ~n28793 & ~n28794 ;
  assign n28795 = ~\sport1_cfg_FSi_cnt_reg[5]/NET0131  & \sport1_regs_FSDIVreg_DO_reg[5]/NET0131  ;
  assign n28796 = ~\sport1_cfg_FSi_cnt_reg[10]/NET0131  & \sport1_regs_FSDIVreg_DO_reg[10]/NET0131  ;
  assign n28824 = ~n28795 & ~n28796 ;
  assign n28843 = n28823 & n28824 ;
  assign n28789 = \sport1_cfg_FSi_cnt_reg[8]/NET0131  & ~\sport1_regs_FSDIVreg_DO_reg[8]/NET0131  ;
  assign n28790 = ~\sport1_cfg_FSi_cnt_reg[0]/NET0131  & \sport1_regs_FSDIVreg_DO_reg[0]/NET0131  ;
  assign n28821 = ~n28789 & ~n28790 ;
  assign n28791 = ~\sport1_cfg_FSi_cnt_reg[11]/NET0131  & \sport1_regs_FSDIVreg_DO_reg[11]/NET0131  ;
  assign n28792 = \sport1_cfg_FSi_cnt_reg[4]/NET0131  & ~\sport1_regs_FSDIVreg_DO_reg[4]/NET0131  ;
  assign n28822 = ~n28791 & ~n28792 ;
  assign n28844 = n28821 & n28822 ;
  assign n28845 = n28843 & n28844 ;
  assign n28801 = ~\sport1_cfg_FSi_cnt_reg[1]/NET0131  & \sport1_regs_FSDIVreg_DO_reg[1]/NET0131  ;
  assign n28802 = ~\sport1_cfg_FSi_cnt_reg[12]/NET0131  & \sport1_regs_FSDIVreg_DO_reg[12]/NET0131  ;
  assign n28827 = ~n28801 & ~n28802 ;
  assign n28803 = \sport1_cfg_FSi_cnt_reg[15]/NET0131  & ~\sport1_regs_FSDIVreg_DO_reg[15]/NET0131  ;
  assign n28804 = \sport1_cfg_FSi_cnt_reg[0]/NET0131  & ~\sport1_regs_FSDIVreg_DO_reg[0]/NET0131  ;
  assign n28828 = ~n28803 & ~n28804 ;
  assign n28841 = n28827 & n28828 ;
  assign n28797 = ~\sport1_cfg_FSi_cnt_reg[4]/NET0131  & \sport1_regs_FSDIVreg_DO_reg[4]/NET0131  ;
  assign n28798 = ~\sport1_cfg_FSi_cnt_reg[3]/NET0131  & \sport1_regs_FSDIVreg_DO_reg[3]/NET0131  ;
  assign n28825 = ~n28797 & ~n28798 ;
  assign n28799 = \sport1_cfg_FSi_cnt_reg[10]/NET0131  & ~\sport1_regs_FSDIVreg_DO_reg[10]/NET0131  ;
  assign n28800 = ~\sport1_cfg_FSi_cnt_reg[2]/NET0131  & \sport1_regs_FSDIVreg_DO_reg[2]/NET0131  ;
  assign n28826 = ~n28799 & ~n28800 ;
  assign n28842 = n28825 & n28826 ;
  assign n28846 = n28841 & n28842 ;
  assign n28850 = n28845 & n28846 ;
  assign n28851 = n28849 & n28850 ;
  assign n28852 = ~n28788 & ~n28851 ;
  assign n28853 = \memc_usysr_DO_reg[11]/NET0131  & \sport1_cfg_SP_ENg_reg/NET0131  ;
  assign n28854 = ~n28852 & n28853 ;
  assign n28855 = ~n28786 & ~n28854 ;
  assign n28871 = ~\sport1_cfg_FSi_cnt_reg[15]/NET0131  & ~n28870 ;
  assign n28873 = n28855 & ~n28871 ;
  assign n28874 = ~n28872 & n28873 ;
  assign n28875 = ~n28787 & ~n28874 ;
  assign n28876 = ~\sport0_cfg_SP_ENg_D1_reg/P0001  & \sport0_cfg_SP_ENg_reg/NET0131  ;
  assign n28877 = \sport0_regs_FSDIVreg_DO_reg[15]/NET0131  & n28876 ;
  assign n28946 = \sport0_cfg_FSi_cnt_reg[0]/NET0131  & \sport0_cfg_SP_ENg_reg/NET0131  ;
  assign n28947 = \sport0_cfg_FSi_cnt_reg[1]/NET0131  & n28946 ;
  assign n28948 = \sport0_cfg_FSi_cnt_reg[2]/NET0131  & n28947 ;
  assign n28949 = \sport0_cfg_FSi_cnt_reg[3]/NET0131  & n28948 ;
  assign n28950 = \sport0_cfg_FSi_cnt_reg[4]/NET0131  & n28949 ;
  assign n28951 = \sport0_cfg_FSi_cnt_reg[5]/NET0131  & n28950 ;
  assign n28952 = \sport0_cfg_FSi_cnt_reg[6]/NET0131  & n28951 ;
  assign n28953 = \sport0_cfg_FSi_cnt_reg[7]/NET0131  & n28952 ;
  assign n28954 = \sport0_cfg_FSi_cnt_reg[8]/NET0131  & n28953 ;
  assign n28955 = \sport0_cfg_FSi_cnt_reg[9]/NET0131  & n28954 ;
  assign n28956 = \sport0_cfg_FSi_cnt_reg[10]/NET0131  & n28955 ;
  assign n28957 = \sport0_cfg_FSi_cnt_reg[11]/NET0131  & n28956 ;
  assign n28958 = \sport0_cfg_FSi_cnt_reg[12]/NET0131  & n28957 ;
  assign n28959 = \sport0_cfg_FSi_cnt_reg[13]/NET0131  & n28958 ;
  assign n28960 = \sport0_cfg_FSi_cnt_reg[14]/NET0131  & n28959 ;
  assign n28962 = \sport0_cfg_FSi_cnt_reg[15]/NET0131  & n28960 ;
  assign n28878 = ~\IRFS0_pad  & ~\ITFS0_pad  ;
  assign n28899 = \sport0_cfg_FSi_cnt_reg[11]/NET0131  & ~\sport0_regs_FSDIVreg_DO_reg[11]/NET0131  ;
  assign n28900 = \sport0_cfg_FSi_cnt_reg[14]/NET0131  & ~\sport0_regs_FSDIVreg_DO_reg[14]/NET0131  ;
  assign n28921 = ~n28899 & ~n28900 ;
  assign n28901 = ~\sport0_cfg_FSi_cnt_reg[9]/NET0131  & \sport0_regs_FSDIVreg_DO_reg[9]/NET0131  ;
  assign n28902 = \sport0_cfg_FSi_cnt_reg[3]/NET0131  & ~\sport0_regs_FSDIVreg_DO_reg[3]/NET0131  ;
  assign n28922 = ~n28901 & ~n28902 ;
  assign n28929 = n28921 & n28922 ;
  assign n28895 = \sport0_cfg_FSi_cnt_reg[2]/NET0131  & ~\sport0_regs_FSDIVreg_DO_reg[2]/NET0131  ;
  assign n28896 = \sport0_cfg_FSi_cnt_reg[7]/NET0131  & ~\sport0_regs_FSDIVreg_DO_reg[7]/NET0131  ;
  assign n28919 = ~n28895 & ~n28896 ;
  assign n28897 = \sport0_cfg_FSi_cnt_reg[0]/NET0131  & ~\sport0_regs_FSDIVreg_DO_reg[0]/NET0131  ;
  assign n28898 = \sport0_cfg_FSi_cnt_reg[9]/NET0131  & ~\sport0_regs_FSDIVreg_DO_reg[9]/NET0131  ;
  assign n28920 = ~n28897 & ~n28898 ;
  assign n28930 = n28919 & n28920 ;
  assign n28937 = n28929 & n28930 ;
  assign n28907 = \sport0_cfg_FSi_cnt_reg[13]/NET0131  & ~\sport0_regs_FSDIVreg_DO_reg[13]/NET0131  ;
  assign n28908 = ~\sport0_cfg_FSi_cnt_reg[15]/NET0131  & \sport0_regs_FSDIVreg_DO_reg[15]/NET0131  ;
  assign n28925 = ~n28907 & ~n28908 ;
  assign n28909 = \sport0_cfg_FSi_cnt_reg[12]/NET0131  & ~\sport0_regs_FSDIVreg_DO_reg[12]/NET0131  ;
  assign n28910 = ~\sport0_cfg_FSi_cnt_reg[6]/NET0131  & \sport0_regs_FSDIVreg_DO_reg[6]/NET0131  ;
  assign n28926 = ~n28909 & ~n28910 ;
  assign n28927 = n28925 & n28926 ;
  assign n28903 = ~\sport0_cfg_FSi_cnt_reg[7]/NET0131  & \sport0_regs_FSDIVreg_DO_reg[7]/NET0131  ;
  assign n28904 = ~\sport0_cfg_FSi_cnt_reg[14]/NET0131  & \sport0_regs_FSDIVreg_DO_reg[14]/NET0131  ;
  assign n28923 = ~n28903 & ~n28904 ;
  assign n28905 = ~\sport0_cfg_FSi_cnt_reg[13]/NET0131  & \sport0_regs_FSDIVreg_DO_reg[13]/NET0131  ;
  assign n28906 = \sport0_cfg_FSi_cnt_reg[6]/NET0131  & ~\sport0_regs_FSDIVreg_DO_reg[6]/NET0131  ;
  assign n28924 = ~n28905 & ~n28906 ;
  assign n28928 = n28923 & n28924 ;
  assign n28938 = n28927 & n28928 ;
  assign n28939 = n28937 & n28938 ;
  assign n28883 = \sport0_cfg_FSi_cnt_reg[5]/NET0131  & ~\sport0_regs_FSDIVreg_DO_reg[5]/NET0131  ;
  assign n28884 = ~\sport0_cfg_FSi_cnt_reg[8]/NET0131  & \sport0_regs_FSDIVreg_DO_reg[8]/NET0131  ;
  assign n28913 = ~n28883 & ~n28884 ;
  assign n28885 = ~\sport0_cfg_FSi_cnt_reg[5]/NET0131  & \sport0_regs_FSDIVreg_DO_reg[5]/NET0131  ;
  assign n28886 = ~\sport0_cfg_FSi_cnt_reg[10]/NET0131  & \sport0_regs_FSDIVreg_DO_reg[10]/NET0131  ;
  assign n28914 = ~n28885 & ~n28886 ;
  assign n28933 = n28913 & n28914 ;
  assign n28879 = \sport0_cfg_FSi_cnt_reg[8]/NET0131  & ~\sport0_regs_FSDIVreg_DO_reg[8]/NET0131  ;
  assign n28880 = ~\sport0_cfg_FSi_cnt_reg[1]/NET0131  & \sport0_regs_FSDIVreg_DO_reg[1]/NET0131  ;
  assign n28911 = ~n28879 & ~n28880 ;
  assign n28881 = ~\sport0_cfg_FSi_cnt_reg[11]/NET0131  & \sport0_regs_FSDIVreg_DO_reg[11]/NET0131  ;
  assign n28882 = \sport0_cfg_FSi_cnt_reg[4]/NET0131  & ~\sport0_regs_FSDIVreg_DO_reg[4]/NET0131  ;
  assign n28912 = ~n28881 & ~n28882 ;
  assign n28934 = n28911 & n28912 ;
  assign n28935 = n28933 & n28934 ;
  assign n28891 = ~\sport0_cfg_FSi_cnt_reg[2]/NET0131  & \sport0_regs_FSDIVreg_DO_reg[2]/NET0131  ;
  assign n28892 = ~\sport0_cfg_FSi_cnt_reg[12]/NET0131  & \sport0_regs_FSDIVreg_DO_reg[12]/NET0131  ;
  assign n28917 = ~n28891 & ~n28892 ;
  assign n28893 = \sport0_cfg_FSi_cnt_reg[15]/NET0131  & ~\sport0_regs_FSDIVreg_DO_reg[15]/NET0131  ;
  assign n28894 = \sport0_cfg_FSi_cnt_reg[1]/NET0131  & ~\sport0_regs_FSDIVreg_DO_reg[1]/NET0131  ;
  assign n28918 = ~n28893 & ~n28894 ;
  assign n28931 = n28917 & n28918 ;
  assign n28887 = ~\sport0_cfg_FSi_cnt_reg[4]/NET0131  & \sport0_regs_FSDIVreg_DO_reg[4]/NET0131  ;
  assign n28888 = ~\sport0_cfg_FSi_cnt_reg[0]/NET0131  & \sport0_regs_FSDIVreg_DO_reg[0]/NET0131  ;
  assign n28915 = ~n28887 & ~n28888 ;
  assign n28889 = \sport0_cfg_FSi_cnt_reg[10]/NET0131  & ~\sport0_regs_FSDIVreg_DO_reg[10]/NET0131  ;
  assign n28890 = ~\sport0_cfg_FSi_cnt_reg[3]/NET0131  & \sport0_regs_FSDIVreg_DO_reg[3]/NET0131  ;
  assign n28916 = ~n28889 & ~n28890 ;
  assign n28932 = n28915 & n28916 ;
  assign n28936 = n28931 & n28932 ;
  assign n28940 = n28935 & n28936 ;
  assign n28941 = n28939 & n28940 ;
  assign n28942 = ~n28878 & ~n28941 ;
  assign n28943 = \memc_usysr_DO_reg[12]/NET0131  & \sport0_cfg_SP_ENg_reg/NET0131  ;
  assign n28944 = ~n28942 & n28943 ;
  assign n28945 = ~n28876 & ~n28944 ;
  assign n28961 = ~\sport0_cfg_FSi_cnt_reg[15]/NET0131  & ~n28960 ;
  assign n28963 = n28945 & ~n28961 ;
  assign n28964 = ~n28962 & n28963 ;
  assign n28965 = ~n28877 & ~n28964 ;
  assign n28968 = ~n17836 & n18271 ;
  assign n28967 = ~\core_eu_em_mac_em_reg_mr0swe_DO_reg[13]/P0001  & ~n18271 ;
  assign n28969 = n18273 & ~n28967 ;
  assign n28970 = ~n28968 & n28969 ;
  assign n28966 = \core_eu_em_mac_em_reg_mr0swe_DO_reg[13]/P0001  & ~n18266 ;
  assign n28971 = ~n18270 & ~n28966 ;
  assign n28972 = ~n28970 & n28971 ;
  assign n28973 = ~n18262 & ~n28972 ;
  assign n28974 = n18262 & ~n19636 ;
  assign n28975 = ~n28973 & ~n28974 ;
  assign n28976 = n14752 & n19636 ;
  assign n28977 = n17836 & n18328 ;
  assign n28978 = \core_eu_em_mac_em_reg_mr0rwe_DO_reg[13]/P0001  & ~n18330 ;
  assign n28979 = n18334 & ~n28978 ;
  assign n28980 = ~n28977 & n28979 ;
  assign n28981 = ~n28976 & ~n28980 ;
  assign n28982 = ~n26301 & n26333 ;
  assign n28983 = \sport1_txctl_TXSHT_reg[11]/P0001  & ~n22677 ;
  assign n28984 = \sport1_txctl_TX_reg[12]/P0001  & n22677 ;
  assign n28985 = ~n28983 & ~n28984 ;
  assign n28988 = ~n14623 & n28561 ;
  assign n28987 = \core_c_dec_MTAR_E_reg/P0001  & n18276 ;
  assign n28989 = ~n28564 & ~n28987 ;
  assign n28990 = ~n28988 & n28989 ;
  assign n28991 = n28559 & ~n28990 ;
  assign n28992 = n28572 & ~n28574 ;
  assign n28993 = n12972 & n28992 ;
  assign n28994 = ~n28576 & ~n28993 ;
  assign n28995 = n28569 & ~n28994 ;
  assign n29010 = ~n11424 & ~n28598 ;
  assign n29008 = ~n11444 & ~n28594 ;
  assign n29009 = ~n11448 & ~n28589 ;
  assign n29011 = ~n29008 & ~n29009 ;
  assign n29012 = ~n29010 & n29011 ;
  assign n29013 = n28607 & n29012 ;
  assign n29014 = n28572 & n29013 ;
  assign n29007 = ~n11525 & ~n28572 ;
  assign n29015 = n28584 & ~n29007 ;
  assign n29016 = ~n29014 & n29015 ;
  assign n28998 = ~n11525 & n28572 ;
  assign n28996 = ~n12972 & ~n28572 ;
  assign n28997 = n28569 & n28574 ;
  assign n28999 = ~n28996 & n28997 ;
  assign n29000 = ~n28998 & n28999 ;
  assign n29004 = ~n11315 & ~n28624 ;
  assign n28986 = ~n11311 & ~n28556 ;
  assign n29002 = ~n18940 & n28636 ;
  assign n29019 = ~n28986 & ~n29002 ;
  assign n29020 = ~n29004 & n29019 ;
  assign n29006 = ~n18831 & n28627 ;
  assign n29005 = n12972 & n28619 ;
  assign n29001 = ~n11341 & ~n28634 ;
  assign n29003 = n11525 & n28630 ;
  assign n29017 = ~n29001 & ~n29003 ;
  assign n29018 = ~n29005 & n29017 ;
  assign n29021 = ~n29006 & n29018 ;
  assign n29022 = n29020 & n29021 ;
  assign n29023 = ~n29000 & n29022 ;
  assign n29024 = ~n29016 & n29023 ;
  assign n29025 = ~n28995 & n29024 ;
  assign n29026 = ~n28991 & n29025 ;
  assign n29027 = n28550 & ~n29026 ;
  assign n29033 = n18276 & n28660 ;
  assign n29030 = n11428 & ~n28652 ;
  assign n29029 = n11440 & n28652 ;
  assign n29031 = ~n28660 & ~n29029 ;
  assign n29032 = ~n29030 & n29031 ;
  assign n29034 = ~n28649 & ~n29032 ;
  assign n29035 = ~n29033 & n29034 ;
  assign n29028 = ~\core_eu_em_mac_em_reg_mxopwe_DO_reg[6]/P0001  & n28649 ;
  assign n29036 = ~n28550 & ~n29028 ;
  assign n29037 = ~n29035 & n29036 ;
  assign n29038 = ~n29027 & ~n29037 ;
  assign n29039 = ~n14634 & n28561 ;
  assign n29040 = \core_c_dec_MTAR_E_reg/P0001  & n20259 ;
  assign n29041 = ~n28564 & ~n29040 ;
  assign n29042 = ~n29039 & n29041 ;
  assign n29043 = n28559 & ~n29042 ;
  assign n29090 = ~n10911 & n28577 ;
  assign n29089 = ~n12938 & ~n28577 ;
  assign n29091 = ~n28575 & ~n29089 ;
  assign n29092 = ~n29090 & n29091 ;
  assign n29093 = ~n28576 & ~n29092 ;
  assign n29094 = n28569 & ~n29093 ;
  assign n29100 = ~n10878 & ~n28594 ;
  assign n29098 = ~n10882 & ~n28598 ;
  assign n29099 = ~n10858 & ~n28589 ;
  assign n29101 = ~n29098 & ~n29099 ;
  assign n29102 = ~n29100 & n29101 ;
  assign n29103 = n28607 & n29102 ;
  assign n29104 = n28572 & n29103 ;
  assign n29097 = ~n10911 & ~n28572 ;
  assign n29105 = n28584 & ~n29097 ;
  assign n29106 = ~n29104 & n29105 ;
  assign n29047 = ~n18002 & n20107 ;
  assign n29059 = n18071 & n18748 ;
  assign n29057 = ~n17922 & ~n18167 ;
  assign n29058 = ~n18108 & ~n18129 ;
  assign n29069 = ~n29057 & ~n29058 ;
  assign n29070 = ~n29059 & n29069 ;
  assign n29051 = ~n18114 & n18719 ;
  assign n29054 = n17934 & n18055 ;
  assign n29053 = \core_c_dec_IRE_reg[11]/NET0131  & ~n10797 ;
  assign n29065 = ~n18192 & ~n29053 ;
  assign n29066 = ~n29054 & n29065 ;
  assign n29067 = ~n29051 & n29066 ;
  assign n29050 = ~n18091 & ~n18189 ;
  assign n29056 = ~n18104 & ~n18133 ;
  assign n29068 = ~n29050 & ~n29056 ;
  assign n29071 = n29067 & n29068 ;
  assign n29046 = n18088 & ~n18895 ;
  assign n29072 = n18041 & ~n29046 ;
  assign n29079 = n29071 & n29072 ;
  assign n29080 = n29070 & n29079 ;
  assign n29060 = n18765 & ~n18781 ;
  assign n29061 = n18171 & ~n19979 ;
  assign n29075 = ~n29060 & ~n29061 ;
  assign n29062 = ~n18135 & ~n18149 ;
  assign n29063 = ~n17981 & ~n18046 ;
  assign n29064 = n18115 & ~n29063 ;
  assign n29076 = ~n29062 & ~n29064 ;
  assign n29077 = n29075 & n29076 ;
  assign n29048 = n17925 & ~n19818 ;
  assign n29049 = ~n18069 & ~n19787 ;
  assign n29073 = ~n29048 & n29049 ;
  assign n29052 = n17978 & n20084 ;
  assign n29055 = n18111 & ~n19857 ;
  assign n29074 = n29052 & ~n29055 ;
  assign n29078 = n29073 & n29074 ;
  assign n29081 = n29077 & n29078 ;
  assign n29082 = n18726 & n29081 ;
  assign n29083 = n29080 & n29082 ;
  assign n29084 = n18800 & n29083 ;
  assign n29085 = n29047 & n29084 ;
  assign n29086 = n28627 & ~n29085 ;
  assign n29096 = n12938 & n28619 ;
  assign n29045 = ~n10694 & ~n28634 ;
  assign n29095 = n10911 & n28630 ;
  assign n29107 = ~n29045 & ~n29095 ;
  assign n29108 = ~n29096 & n29107 ;
  assign n29088 = ~n20288 & n28636 ;
  assign n29044 = ~n10801 & ~n28624 ;
  assign n29087 = ~n10797 & ~n28556 ;
  assign n29109 = ~n29044 & ~n29087 ;
  assign n29110 = ~n29088 & n29109 ;
  assign n29111 = n29108 & n29110 ;
  assign n29112 = ~n29086 & n29111 ;
  assign n29113 = ~n29106 & n29112 ;
  assign n29114 = ~n29094 & n29113 ;
  assign n29115 = ~n29043 & n29114 ;
  assign n29116 = n28550 & ~n29115 ;
  assign n29122 = n20259 & n28660 ;
  assign n29119 = n10866 & ~n28652 ;
  assign n29118 = n10874 & n28652 ;
  assign n29120 = ~n28660 & ~n29118 ;
  assign n29121 = ~n29119 & n29120 ;
  assign n29123 = ~n28649 & ~n29121 ;
  assign n29124 = ~n29122 & n29123 ;
  assign n29117 = ~\core_eu_em_mac_em_reg_mxopwe_DO_reg[5]/P0001  & n28649 ;
  assign n29125 = ~n28550 & ~n29117 ;
  assign n29126 = ~n29124 & n29125 ;
  assign n29127 = ~n29116 & ~n29126 ;
  assign n29130 = ~n14600 & n28561 ;
  assign n29129 = \core_c_dec_MTAR_E_reg/P0001  & n20080 ;
  assign n29131 = ~n28564 & ~n29129 ;
  assign n29132 = ~n29130 & n29131 ;
  assign n29133 = n28559 & ~n29132 ;
  assign n29134 = n12904 & n28992 ;
  assign n29135 = ~n28576 & ~n29134 ;
  assign n29136 = n28569 & ~n29135 ;
  assign n29150 = ~n9865 & ~n28598 ;
  assign n29148 = ~n9845 & ~n28589 ;
  assign n29149 = ~n9869 & ~n28594 ;
  assign n29151 = ~n29148 & ~n29149 ;
  assign n29152 = ~n29150 & n29151 ;
  assign n29153 = n28607 & n29152 ;
  assign n29154 = n28572 & n29153 ;
  assign n29147 = ~n10069 & ~n28572 ;
  assign n29155 = n28584 & ~n29147 ;
  assign n29156 = ~n29154 & n29155 ;
  assign n29138 = ~n10069 & n28572 ;
  assign n29137 = ~n12904 & ~n28572 ;
  assign n29139 = n28997 & ~n29137 ;
  assign n29140 = ~n29138 & n29139 ;
  assign n29146 = ~n9951 & ~n28624 ;
  assign n29141 = ~n9947 & ~n28556 ;
  assign n29143 = ~n22911 & n28636 ;
  assign n29159 = ~n29141 & ~n29143 ;
  assign n29160 = ~n29146 & n29159 ;
  assign n29128 = ~n20142 & n28627 ;
  assign n29145 = n12904 & n28619 ;
  assign n29142 = ~n9912 & ~n28634 ;
  assign n29144 = n10069 & n28630 ;
  assign n29157 = ~n29142 & ~n29144 ;
  assign n29158 = ~n29145 & n29157 ;
  assign n29161 = ~n29128 & n29158 ;
  assign n29162 = n29160 & n29161 ;
  assign n29163 = ~n29140 & n29162 ;
  assign n29164 = ~n29156 & n29163 ;
  assign n29165 = ~n29136 & n29164 ;
  assign n29166 = ~n29133 & n29165 ;
  assign n29167 = n28550 & ~n29166 ;
  assign n29173 = n20080 & n28660 ;
  assign n29170 = n9849 & ~n28652 ;
  assign n29169 = n9861 & n28652 ;
  assign n29171 = ~n28660 & ~n29169 ;
  assign n29172 = ~n29170 & n29171 ;
  assign n29174 = ~n28649 & ~n29172 ;
  assign n29175 = ~n29173 & n29174 ;
  assign n29168 = ~\core_eu_em_mac_em_reg_mxopwe_DO_reg[4]/P0001  & n28649 ;
  assign n29176 = ~n28550 & ~n29168 ;
  assign n29177 = ~n29175 & n29176 ;
  assign n29178 = ~n29167 & ~n29177 ;
  assign n29181 = n14573 & n28561 ;
  assign n29180 = \core_c_dec_MTAR_E_reg/P0001  & n18974 ;
  assign n29182 = ~n28564 & ~n29180 ;
  assign n29183 = ~n29181 & n29182 ;
  assign n29184 = n28559 & ~n29183 ;
  assign n29186 = ~n9435 & n28577 ;
  assign n29185 = ~n12802 & ~n28577 ;
  assign n29187 = ~n28575 & ~n29185 ;
  assign n29188 = ~n29186 & n29187 ;
  assign n29189 = ~n28576 & ~n29188 ;
  assign n29190 = n28569 & ~n29189 ;
  assign n29200 = ~n9205 & ~n28589 ;
  assign n29198 = ~n9225 & ~n28594 ;
  assign n29199 = ~n9229 & ~n28598 ;
  assign n29201 = ~n29198 & ~n29199 ;
  assign n29202 = ~n29200 & n29201 ;
  assign n29203 = n28607 & n29202 ;
  assign n29204 = n28572 & n29203 ;
  assign n29197 = ~n9435 & ~n28572 ;
  assign n29205 = n28584 & ~n29197 ;
  assign n29206 = ~n29204 & n29205 ;
  assign n29192 = ~n21046 & n28627 ;
  assign n29193 = ~n9297 & ~n28634 ;
  assign n29194 = n12802 & n28619 ;
  assign n29207 = ~n29193 & ~n29194 ;
  assign n29195 = n9435 & n28630 ;
  assign n29196 = ~n19008 & n28636 ;
  assign n29208 = ~n29195 & ~n29196 ;
  assign n29209 = n29207 & n29208 ;
  assign n29179 = ~n9280 & ~n28556 ;
  assign n29191 = ~n9276 & ~n28624 ;
  assign n29210 = ~n29179 & ~n29191 ;
  assign n29211 = n29209 & n29210 ;
  assign n29212 = ~n29192 & n29211 ;
  assign n29213 = ~n29206 & n29212 ;
  assign n29214 = ~n29190 & n29213 ;
  assign n29215 = ~n29184 & n29214 ;
  assign n29216 = n28550 & ~n29215 ;
  assign n29222 = n18974 & n28660 ;
  assign n29219 = n9213 & ~n28652 ;
  assign n29218 = n9221 & n28652 ;
  assign n29220 = ~n28660 & ~n29218 ;
  assign n29221 = ~n29219 & n29220 ;
  assign n29223 = ~n28649 & ~n29221 ;
  assign n29224 = ~n29222 & n29223 ;
  assign n29217 = ~\core_eu_em_mac_em_reg_mxopwe_DO_reg[1]/P0001  & n28649 ;
  assign n29225 = ~n28550 & ~n29217 ;
  assign n29226 = ~n29224 & n29225 ;
  assign n29227 = ~n29216 & ~n29226 ;
  assign n29228 = \sport0_cfg_SCLKi_cnt_reg[14]/NET0131  & n19552 ;
  assign n29230 = \sport0_cfg_SCLKi_cnt_reg[15]/NET0131  & n29228 ;
  assign n29229 = ~\sport0_cfg_SCLKi_cnt_reg[15]/NET0131  & ~n29228 ;
  assign n29231 = n19197 & ~n29229 ;
  assign n29232 = ~n29230 & n29231 ;
  assign n29287 = \core_c_dec_MTAR_E_reg/P0001  & n17820 ;
  assign n29288 = n19214 & n19278 ;
  assign n29289 = ~n19224 & ~n29288 ;
  assign n29290 = ~\core_c_dec_MTAR_E_reg/P0001  & ~n29289 ;
  assign n29291 = ~n29287 & ~n29290 ;
  assign n29292 = n28559 & ~n29291 ;
  assign n29306 = n13006 & n28992 ;
  assign n29307 = ~n28576 & ~n29306 ;
  assign n29308 = n28569 & ~n29307 ;
  assign n29293 = ~n12028 & ~n28589 ;
  assign n29297 = ~n28605 & ~n29293 ;
  assign n29296 = ~n12024 & ~n28594 ;
  assign n29294 = n28592 & n28601 ;
  assign n29295 = ~n7206 & ~n28598 ;
  assign n29298 = ~n29294 & ~n29295 ;
  assign n29299 = ~n29296 & n29298 ;
  assign n29300 = n29297 & n29299 ;
  assign n29301 = n28577 & ~n29300 ;
  assign n29302 = n11265 & ~n28572 ;
  assign n29303 = n28574 & n29302 ;
  assign n29304 = ~n29301 & ~n29303 ;
  assign n29305 = ~n28569 & ~n29304 ;
  assign n29310 = ~n12743 & n28572 ;
  assign n29309 = ~n12771 & ~n28572 ;
  assign n29311 = n28997 & ~n29309 ;
  assign n29312 = ~n29310 & n29311 ;
  assign n29317 = n12743 & n28630 ;
  assign n29313 = n12771 & n28619 ;
  assign n29316 = ~n11983 & ~n28634 ;
  assign n29319 = ~n29313 & ~n29316 ;
  assign n29320 = ~n29317 & n29319 ;
  assign n29314 = ~n12000 & ~n28556 ;
  assign n29315 = ~n11992 & ~n28624 ;
  assign n29321 = ~n29314 & ~n29315 ;
  assign n29322 = n29320 & n29321 ;
  assign n29244 = ~n18091 & ~n18104 ;
  assign n29245 = n18071 & n18187 ;
  assign n29271 = ~n29244 & ~n29245 ;
  assign n29246 = n18112 & ~n18907 ;
  assign n29247 = ~n18127 & n18147 ;
  assign n29272 = ~n29246 & ~n29247 ;
  assign n29273 = n29271 & n29272 ;
  assign n29236 = n17980 & ~n18135 ;
  assign n29237 = n18171 & n18893 ;
  assign n29269 = ~n29236 & ~n29237 ;
  assign n29240 = n18139 & n18183 ;
  assign n29243 = n18046 & n18745 ;
  assign n29270 = ~n29240 & ~n29243 ;
  assign n29274 = n29269 & n29270 ;
  assign n29280 = n29273 & n29274 ;
  assign n29281 = n18724 & n29280 ;
  assign n29248 = n17979 & n18077 ;
  assign n29249 = ~n17981 & ~n29248 ;
  assign n29250 = ~n18083 & n29249 ;
  assign n29251 = n17945 & ~n29250 ;
  assign n29252 = n17978 & ~n29251 ;
  assign n29259 = n18162 & ~n19857 ;
  assign n29238 = n18124 & ~n19804 ;
  assign n29239 = ~n18783 & ~n21010 ;
  assign n29277 = ~n29238 & n29239 ;
  assign n29278 = ~n29259 & n29277 ;
  assign n29233 = ~n18127 & n18148 ;
  assign n29234 = n18039 & ~n19722 ;
  assign n29265 = ~n29233 & ~n29234 ;
  assign n29241 = ~n17935 & n18072 ;
  assign n29242 = n17971 & n18051 ;
  assign n29266 = ~n29241 & ~n29242 ;
  assign n29267 = n29265 & n29266 ;
  assign n29254 = n18056 & ~n18991 ;
  assign n29256 = n18191 & ~n19722 ;
  assign n29261 = ~n29254 & ~n29256 ;
  assign n29257 = n18153 & n18166 ;
  assign n29258 = ~n17935 & n17955 ;
  assign n29262 = ~n29257 & ~n29258 ;
  assign n29263 = n29261 & n29262 ;
  assign n29253 = n18055 & ~n18189 ;
  assign n29255 = \core_c_dec_IRE_reg[11]/NET0131  & ~n11992 ;
  assign n29260 = ~n29253 & ~n29255 ;
  assign n29264 = ~n21199 & n29260 ;
  assign n29268 = n29263 & n29264 ;
  assign n29275 = n29267 & n29268 ;
  assign n29235 = ~n18114 & n20104 ;
  assign n29276 = n20108 & ~n29235 ;
  assign n29279 = n29275 & n29276 ;
  assign n29282 = n29278 & n29279 ;
  assign n29283 = n29252 & n29282 ;
  assign n29284 = n29281 & n29283 ;
  assign n29285 = n19793 & n29284 ;
  assign n29286 = n28636 & ~n29285 ;
  assign n29318 = ~n19769 & n28627 ;
  assign n29323 = ~n29286 & ~n29318 ;
  assign n29324 = n29322 & n29323 ;
  assign n29325 = ~n29312 & n29324 ;
  assign n29326 = ~n29305 & n29325 ;
  assign n29327 = ~n29308 & n29326 ;
  assign n29328 = ~n29292 & n29327 ;
  assign n29329 = n28550 & ~n29328 ;
  assign n29335 = n17820 & n28660 ;
  assign n29332 = n12020 & ~n28652 ;
  assign n29331 = n12016 & n28652 ;
  assign n29333 = ~n28660 & ~n29331 ;
  assign n29334 = ~n29332 & n29333 ;
  assign n29336 = ~n28649 & ~n29334 ;
  assign n29337 = ~n29335 & n29336 ;
  assign n29330 = ~\core_eu_em_mac_em_reg_mxopwe_DO_reg[15]/P0001  & n28649 ;
  assign n29338 = ~n28550 & ~n29330 ;
  assign n29339 = ~n29337 & n29338 ;
  assign n29340 = ~n29329 & ~n29339 ;
  assign n29341 = \sport0_txctl_TXSHT_reg[11]/P0001  & ~n19960 ;
  assign n29342 = \sport0_txctl_TX_reg[12]/P0001  & n19960 ;
  assign n29343 = ~n29341 & ~n29342 ;
  assign n29345 = n9435 & n28725 ;
  assign n29344 = n12802 & n28729 ;
  assign n29351 = ~\core_c_psq_MSTAT_reg_DO_reg[0]/P0002  & ~\core_eu_em_mac_em_reg_mfrwe_DO_reg[1]/P0001  ;
  assign n29352 = \core_c_psq_MSTAT_reg_DO_reg[0]/P0002  & ~\core_eu_em_mac_em_reg_mfswe_DO_reg[1]/P0001  ;
  assign n29353 = ~n29351 & ~n29352 ;
  assign n29354 = n28741 & n29353 ;
  assign n29346 = n9209 & n28705 ;
  assign n29347 = n9217 & ~n28705 ;
  assign n29348 = ~n29346 & ~n29347 ;
  assign n29349 = n28735 & n29348 ;
  assign n29350 = n28739 & n29221 ;
  assign n29355 = ~n29349 & ~n29350 ;
  assign n29356 = ~n29354 & n29355 ;
  assign n29357 = ~n29344 & n29356 ;
  assign n29358 = ~n29345 & n29357 ;
  assign n29359 = ~n28543 & ~n29358 ;
  assign n29360 = \core_eu_em_mac_em_reg_myopwe_DO_reg[1]/P0001  & ~n28545 ;
  assign n29361 = ~n29359 & ~n29360 ;
  assign n29362 = ~n28719 & ~n29361 ;
  assign n29363 = n28719 & ~n29215 ;
  assign n29364 = ~n29362 & ~n29363 ;
  assign n29366 = n10069 & n28725 ;
  assign n29365 = n12904 & n28729 ;
  assign n29372 = ~\core_c_psq_MSTAT_reg_DO_reg[0]/P0002  & ~\core_eu_em_mac_em_reg_mfrwe_DO_reg[4]/P0001  ;
  assign n29373 = \core_c_psq_MSTAT_reg_DO_reg[0]/P0002  & ~\core_eu_em_mac_em_reg_mfswe_DO_reg[4]/P0001  ;
  assign n29374 = ~n29372 & ~n29373 ;
  assign n29375 = n28741 & n29374 ;
  assign n29367 = n9853 & n28705 ;
  assign n29368 = n9857 & ~n28705 ;
  assign n29369 = ~n29367 & ~n29368 ;
  assign n29370 = n28735 & n29369 ;
  assign n29371 = n28739 & n29172 ;
  assign n29376 = ~n29370 & ~n29371 ;
  assign n29377 = ~n29375 & n29376 ;
  assign n29378 = ~n29365 & n29377 ;
  assign n29379 = ~n29366 & n29378 ;
  assign n29380 = ~n28543 & ~n29379 ;
  assign n29381 = \core_eu_em_mac_em_reg_myopwe_DO_reg[4]/P0001  & ~n28545 ;
  assign n29382 = ~n29380 & ~n29381 ;
  assign n29383 = ~n28719 & ~n29382 ;
  assign n29384 = n28719 & ~n29166 ;
  assign n29385 = ~n29383 & ~n29384 ;
  assign n29387 = n11525 & n28725 ;
  assign n29386 = n12972 & n28729 ;
  assign n29393 = ~\core_c_psq_MSTAT_reg_DO_reg[0]/P0002  & ~\core_eu_em_mac_em_reg_mfrwe_DO_reg[6]/P0001  ;
  assign n29394 = \core_c_psq_MSTAT_reg_DO_reg[0]/P0002  & ~\core_eu_em_mac_em_reg_mfswe_DO_reg[6]/P0001  ;
  assign n29395 = ~n29393 & ~n29394 ;
  assign n29396 = n28741 & n29395 ;
  assign n29388 = n11436 & n28705 ;
  assign n29389 = n11432 & ~n28705 ;
  assign n29390 = ~n29388 & ~n29389 ;
  assign n29391 = n28735 & n29390 ;
  assign n29392 = n28739 & n29032 ;
  assign n29397 = ~n29391 & ~n29392 ;
  assign n29398 = ~n29396 & n29397 ;
  assign n29399 = ~n29386 & n29398 ;
  assign n29400 = ~n29387 & n29399 ;
  assign n29401 = ~n28543 & ~n29400 ;
  assign n29402 = \core_eu_em_mac_em_reg_myopwe_DO_reg[6]/P0001  & ~n28545 ;
  assign n29403 = ~n29401 & ~n29402 ;
  assign n29404 = ~n28719 & ~n29403 ;
  assign n29405 = n28719 & ~n29026 ;
  assign n29406 = ~n29404 & ~n29405 ;
  assign n29407 = \sport1_cfg_SCLKi_cnt_reg[14]/NET0131  & n20253 ;
  assign n29409 = \sport1_cfg_SCLKi_cnt_reg[15]/NET0131  & n29407 ;
  assign n29408 = ~\sport1_cfg_SCLKi_cnt_reg[15]/NET0131  & ~n29407 ;
  assign n29410 = n19130 & ~n29408 ;
  assign n29411 = ~n29409 & n29410 ;
  assign n29413 = n10911 & n28725 ;
  assign n29412 = n12938 & n28729 ;
  assign n29419 = ~\core_c_psq_MSTAT_reg_DO_reg[0]/P0002  & ~\core_eu_em_mac_em_reg_mfrwe_DO_reg[5]/P0001  ;
  assign n29420 = \core_c_psq_MSTAT_reg_DO_reg[0]/P0002  & ~\core_eu_em_mac_em_reg_mfswe_DO_reg[5]/P0001  ;
  assign n29421 = ~n29419 & ~n29420 ;
  assign n29422 = n28741 & n29421 ;
  assign n29414 = n10862 & n28705 ;
  assign n29415 = n10870 & ~n28705 ;
  assign n29416 = ~n29414 & ~n29415 ;
  assign n29417 = n28735 & n29416 ;
  assign n29418 = n28739 & n29121 ;
  assign n29423 = ~n29417 & ~n29418 ;
  assign n29424 = ~n29422 & n29423 ;
  assign n29425 = ~n29412 & n29424 ;
  assign n29426 = ~n29413 & n29425 ;
  assign n29427 = ~n28543 & ~n29426 ;
  assign n29428 = \core_eu_em_mac_em_reg_myopwe_DO_reg[5]/P0001  & ~n28545 ;
  assign n29429 = ~n29427 & ~n29428 ;
  assign n29430 = ~n28719 & ~n29429 ;
  assign n29431 = n28719 & ~n29115 ;
  assign n29432 = ~n29430 & ~n29431 ;
  assign n29433 = n12771 & n28729 ;
  assign n29434 = n12743 & n28725 ;
  assign n29440 = ~\core_c_psq_MSTAT_reg_DO_reg[0]/P0002  & ~\core_eu_em_mac_em_reg_mfrwe_DO_reg[15]/P0001  ;
  assign n29441 = \core_c_psq_MSTAT_reg_DO_reg[0]/P0002  & ~\core_eu_em_mac_em_reg_mfswe_DO_reg[15]/P0001  ;
  assign n29442 = ~n29440 & ~n29441 ;
  assign n29443 = n28741 & n29442 ;
  assign n29435 = n12008 & n28705 ;
  assign n29436 = n12012 & ~n28705 ;
  assign n29437 = ~n29435 & ~n29436 ;
  assign n29438 = n28735 & n29437 ;
  assign n29439 = n28739 & n29334 ;
  assign n29444 = ~n29438 & ~n29439 ;
  assign n29445 = ~n29443 & n29444 ;
  assign n29446 = ~n29434 & n29445 ;
  assign n29447 = ~n29433 & n29446 ;
  assign n29448 = ~n28543 & ~n29447 ;
  assign n29449 = \core_eu_em_mac_em_reg_myopwe_DO_reg[15]/P0001  & ~n28545 ;
  assign n29450 = ~n29448 & ~n29449 ;
  assign n29451 = ~n28719 & ~n29450 ;
  assign n29452 = n28719 & ~n29328 ;
  assign n29453 = ~n29451 & ~n29452 ;
  assign n29454 = \core_eu_es_sht_es_reg_serwe_DO_reg[7]/P0001  & ~n23598 ;
  assign n29455 = \core_c_dec_MTSE_E_reg/P0001  & n19972 ;
  assign n29456 = ~n23587 & ~n23662 ;
  assign n29457 = ~n23665 & ~n29456 ;
  assign n29458 = ~\core_c_dec_MTSE_E_reg/P0001  & n29457 ;
  assign n29459 = ~n29455 & ~n29458 ;
  assign n29460 = n23598 & ~n29459 ;
  assign n29461 = ~n29454 & ~n29460 ;
  assign n29462 = \core_eu_es_sht_es_reg_serwe_DO_reg[6]/P0001  & ~n23598 ;
  assign n29463 = \core_c_dec_MTSE_E_reg/P0001  & n18276 ;
  assign n29464 = ~n29458 & ~n29463 ;
  assign n29465 = n23598 & ~n29464 ;
  assign n29466 = ~n29462 & ~n29465 ;
  assign n29469 = n18271 & ~n23920 ;
  assign n29468 = ~\core_eu_em_mac_em_reg_mr0swe_DO_reg[12]/P0001  & ~n18271 ;
  assign n29470 = n18273 & ~n29468 ;
  assign n29471 = ~n29469 & n29470 ;
  assign n29467 = \core_eu_em_mac_em_reg_mr0swe_DO_reg[12]/P0001  & ~n18266 ;
  assign n29472 = ~n18270 & ~n29467 ;
  assign n29473 = ~n29471 & n29472 ;
  assign n29474 = ~n18262 & ~n29473 ;
  assign n29475 = n18262 & n19609 ;
  assign n29476 = ~n29474 & ~n29475 ;
  assign n29477 = \core_c_dec_MTSE_E_reg/P0001  & ~n20080 ;
  assign n29478 = n23587 & n23662 ;
  assign n29479 = n29457 & ~n29478 ;
  assign n29480 = ~n23669 & ~n29479 ;
  assign n29481 = ~\core_c_dec_MTSE_E_reg/P0001  & n29480 ;
  assign n29482 = ~n29477 & ~n29481 ;
  assign n29483 = n23598 & ~n29482 ;
  assign n29484 = ~\core_eu_es_sht_es_reg_serwe_DO_reg[4]/P0001  & ~n23598 ;
  assign n29485 = ~n29483 & ~n29484 ;
  assign n29486 = \core_eu_es_sht_es_reg_serwe_DO_reg[5]/P0001  & ~n23598 ;
  assign n29487 = \core_c_dec_MTSE_E_reg/P0001  & n20259 ;
  assign n29488 = ~n29458 & ~n29487 ;
  assign n29489 = n23598 & ~n29488 ;
  assign n29490 = ~n29486 & ~n29489 ;
  assign n29491 = \core_c_dec_MTSE_E_reg/P0001  & ~n21663 ;
  assign n29492 = n27484 & n27486 ;
  assign n29493 = n26275 & ~n29492 ;
  assign n29494 = ~\core_c_dec_MTSE_E_reg/P0001  & ~n29493 ;
  assign n29495 = ~n29491 & ~n29494 ;
  assign n29496 = n23598 & ~n29495 ;
  assign n29497 = ~\core_eu_es_sht_es_reg_serwe_DO_reg[3]/P0001  & ~n23598 ;
  assign n29498 = ~n29496 & ~n29497 ;
  assign n29499 = n14752 & ~n19609 ;
  assign n29500 = n18328 & n23920 ;
  assign n29501 = \core_eu_em_mac_em_reg_mr0rwe_DO_reg[12]/P0001  & ~n18330 ;
  assign n29502 = n18334 & ~n29501 ;
  assign n29503 = ~n29500 & n29502 ;
  assign n29504 = ~n29499 & ~n29503 ;
  assign n29505 = \core_eu_es_sht_es_reg_seswe_DO_reg[6]/P0001  & ~n23677 ;
  assign n29506 = n23677 & ~n29464 ;
  assign n29507 = ~n29505 & ~n29506 ;
  assign n29508 = \core_eu_es_sht_es_reg_seswe_DO_reg[7]/P0001  & ~n23677 ;
  assign n29509 = n23677 & ~n29459 ;
  assign n29510 = ~n29508 & ~n29509 ;
  assign n29511 = \core_eu_es_sht_es_reg_seswe_DO_reg[5]/P0001  & ~n23677 ;
  assign n29512 = n23677 & ~n29488 ;
  assign n29513 = ~n29511 & ~n29512 ;
  assign n29514 = n23677 & ~n29482 ;
  assign n29515 = ~\core_eu_es_sht_es_reg_seswe_DO_reg[4]/P0001  & ~n23677 ;
  assign n29516 = ~n29514 & ~n29515 ;
  assign n29517 = n23677 & ~n29495 ;
  assign n29518 = ~\core_eu_es_sht_es_reg_seswe_DO_reg[3]/P0001  & ~n23677 ;
  assign n29519 = ~n29517 & ~n29518 ;
  assign n29558 = ~n14649 & n28561 ;
  assign n29557 = \core_c_dec_MTAR_E_reg/P0001  & n19504 ;
  assign n29559 = ~n28564 & ~n29557 ;
  assign n29560 = ~n29558 & n29559 ;
  assign n29561 = n28559 & ~n29560 ;
  assign n29562 = n28607 & ~n29295 ;
  assign n29563 = ~n10096 & ~n28589 ;
  assign n29564 = ~n10112 & ~n28594 ;
  assign n29565 = ~n29563 & ~n29564 ;
  assign n29566 = n29562 & n29565 ;
  assign n29567 = n28577 & ~n29566 ;
  assign n29568 = ~n29303 & ~n29567 ;
  assign n29569 = ~n28569 & ~n29568 ;
  assign n29629 = ~n13075 & ~n28572 ;
  assign n29628 = ~n10289 & n28572 ;
  assign n29630 = n28997 & ~n29628 ;
  assign n29631 = ~n29629 & n29630 ;
  assign n29572 = n10289 & n28630 ;
  assign n29570 = ~n10191 & ~n28634 ;
  assign n29571 = n13075 & n28619 ;
  assign n29632 = ~n29570 & ~n29571 ;
  assign n29633 = ~n29572 & n29632 ;
  assign n29573 = ~n10218 & ~n28624 ;
  assign n29574 = ~n10226 & ~n28556 ;
  assign n29634 = ~n29573 & ~n29574 ;
  assign n29635 = n29633 & n29634 ;
  assign n29521 = n19855 & n19873 ;
  assign n29522 = n19713 & n29521 ;
  assign n29533 = ~n18079 & n18765 ;
  assign n29534 = n18758 & ~n18918 ;
  assign n29535 = n18115 & ~n18914 ;
  assign n29536 = ~n29534 & ~n29535 ;
  assign n29537 = n17839 & ~n29536 ;
  assign n29538 = ~n29533 & ~n29537 ;
  assign n29539 = n17929 & ~n29538 ;
  assign n29529 = n18740 & ~n18781 ;
  assign n29530 = n17925 & ~n18898 ;
  assign n29548 = ~n29529 & ~n29530 ;
  assign n29531 = n18099 & ~n19818 ;
  assign n29540 = n18124 & ~n18895 ;
  assign n29549 = ~n29531 & ~n29540 ;
  assign n29550 = n29548 & n29549 ;
  assign n29528 = n18172 & ~n18918 ;
  assign n29524 = n18112 & ~n18914 ;
  assign n29527 = ~n18079 & n19720 ;
  assign n29544 = ~n29524 & ~n29527 ;
  assign n29545 = ~n29528 & n29544 ;
  assign n29532 = \core_c_dec_IRE_reg[11]/NET0131  & ~n10218 ;
  assign n29541 = ~n18037 & ~n29532 ;
  assign n29542 = ~n18053 & n29541 ;
  assign n29520 = ~n18167 & ~n18907 ;
  assign n29523 = ~n18189 & ~n18912 ;
  assign n29543 = ~n29520 & ~n29523 ;
  assign n29546 = n29542 & n29543 ;
  assign n29525 = n18751 & ~n18775 ;
  assign n29526 = ~n17998 & n18748 ;
  assign n29547 = ~n29525 & ~n29526 ;
  assign n29551 = n29546 & n29547 ;
  assign n29552 = n29545 & n29551 ;
  assign n29553 = n29550 & n29552 ;
  assign n29554 = ~n29539 & n29553 ;
  assign n29555 = n29522 & n29554 ;
  assign n29556 = n28636 & ~n29555 ;
  assign n29579 = ~n18065 & ~n18735 ;
  assign n29588 = ~n18114 & n18732 ;
  assign n29578 = ~n18104 & ~n18159 ;
  assign n29582 = n18070 & n18088 ;
  assign n29612 = ~n29578 & ~n29582 ;
  assign n29613 = ~n29588 & n29612 ;
  assign n29620 = n19996 & n29613 ;
  assign n29621 = n29579 & n29620 ;
  assign n29580 = n17925 & ~n19979 ;
  assign n29581 = n18107 & ~n18189 ;
  assign n29594 = ~n18129 & n18179 ;
  assign n29605 = ~n29581 & ~n29594 ;
  assign n29595 = n18131 & ~n18167 ;
  assign n29596 = n17915 & n18172 ;
  assign n29606 = ~n29595 & ~n29596 ;
  assign n29607 = n29605 & n29606 ;
  assign n29616 = ~n29580 & n29607 ;
  assign n29589 = ~n17980 & ~n18071 ;
  assign n29590 = n17945 & ~n29589 ;
  assign n29597 = n18765 & ~n29063 ;
  assign n29617 = ~n29590 & ~n29597 ;
  assign n29618 = n29616 & n29617 ;
  assign n29575 = ~n18091 & n18112 ;
  assign n29610 = ~n18140 & ~n29575 ;
  assign n29576 = n18147 & n18748 ;
  assign n29577 = ~n17922 & n18136 ;
  assign n29611 = ~n29576 & ~n29577 ;
  assign n29614 = n29610 & n29611 ;
  assign n29583 = \core_c_dec_IRE_reg[11]/NET0131  & ~n10226 ;
  assign n29584 = n18106 & ~n18189 ;
  assign n29598 = ~n29583 & ~n29584 ;
  assign n29585 = n18132 & ~n18167 ;
  assign n29586 = n17921 & n18172 ;
  assign n29599 = ~n29585 & ~n29586 ;
  assign n29603 = n29598 & n29599 ;
  assign n29604 = ~n18058 & ~n18783 ;
  assign n29608 = n29603 & n29604 ;
  assign n29587 = n18089 & n18116 ;
  assign n29591 = ~n18129 & n18178 ;
  assign n29600 = ~n29587 & ~n29591 ;
  assign n29592 = n18153 & ~n19722 ;
  assign n29593 = n17934 & n17986 ;
  assign n29601 = ~n29592 & ~n29593 ;
  assign n29602 = n29600 & n29601 ;
  assign n29609 = n17978 & n29602 ;
  assign n29615 = n29608 & n29609 ;
  assign n29619 = n29614 & n29615 ;
  assign n29622 = n29618 & n29619 ;
  assign n29623 = n29621 & n29622 ;
  assign n29624 = n18731 & n20106 ;
  assign n29625 = n29623 & n29624 ;
  assign n29626 = n18800 & n29625 ;
  assign n29627 = n28627 & ~n29626 ;
  assign n29636 = ~n29556 & ~n29627 ;
  assign n29637 = n29635 & n29636 ;
  assign n29638 = ~n29631 & n29637 ;
  assign n29639 = ~n29308 & n29638 ;
  assign n29640 = ~n29569 & n29639 ;
  assign n29641 = ~n29561 & n29640 ;
  assign n29642 = n28719 & ~n29641 ;
  assign n29645 = n13075 & ~n28728 ;
  assign n29646 = ~\core_c_psq_MSTAT_reg_DO_reg[0]/P0002  & ~\core_eu_em_mac_em_reg_mfrwe_DO_reg[9]/P0001  ;
  assign n29647 = \core_c_psq_MSTAT_reg_DO_reg[0]/P0002  & ~\core_eu_em_mac_em_reg_mfswe_DO_reg[9]/P0001  ;
  assign n29648 = ~n29646 & ~n29647 ;
  assign n29649 = n28741 & n29648 ;
  assign n29659 = \core_eu_em_mac_em_reg_myopwe_DO_reg[9]/P0001  & ~n28545 ;
  assign n29660 = ~n29649 & ~n29659 ;
  assign n29651 = n10100 & ~n28652 ;
  assign n29650 = n10116 & n28652 ;
  assign n29652 = ~n28660 & ~n29650 ;
  assign n29653 = ~n29651 & n29652 ;
  assign n29654 = n28739 & n29653 ;
  assign n29655 = n10104 & n28705 ;
  assign n29656 = n10108 & ~n28705 ;
  assign n29657 = ~n29655 & ~n29656 ;
  assign n29658 = n28735 & n29657 ;
  assign n29661 = ~n29654 & ~n29658 ;
  assign n29662 = n29660 & n29661 ;
  assign n29663 = ~n28725 & n29662 ;
  assign n29664 = ~n29645 & n29663 ;
  assign n29643 = ~n28543 & n28725 ;
  assign n29644 = ~n10289 & n29643 ;
  assign n29665 = ~\core_eu_em_mac_em_reg_myopwe_DO_reg[9]/P0001  & n28543 ;
  assign n29666 = ~n28719 & ~n29665 ;
  assign n29667 = ~n29644 & n29666 ;
  assign n29668 = ~n29664 & n29667 ;
  assign n29669 = ~n29642 & ~n29668 ;
  assign n29672 = ~n14551 & n28561 ;
  assign n29671 = \core_c_dec_MTAR_E_reg/P0001  & n17836 ;
  assign n29673 = ~n28564 & ~n29671 ;
  assign n29674 = ~n29672 & n29673 ;
  assign n29675 = n28559 & ~n29674 ;
  assign n29676 = ~n7202 & ~n28589 ;
  assign n29677 = ~n7182 & ~n28594 ;
  assign n29678 = ~n29676 & ~n29677 ;
  assign n29679 = n29562 & n29678 ;
  assign n29680 = n28577 & ~n29679 ;
  assign n29681 = ~n29303 & ~n29680 ;
  assign n29682 = ~n28569 & ~n29681 ;
  assign n29684 = ~n7340 & n28572 ;
  assign n29683 = ~n12658 & ~n28572 ;
  assign n29685 = n28997 & ~n29683 ;
  assign n29686 = ~n29684 & n29685 ;
  assign n29692 = ~n19840 & n28636 ;
  assign n29670 = ~n18211 & n28627 ;
  assign n29689 = n7340 & n28630 ;
  assign n29687 = n12658 & n28619 ;
  assign n29688 = ~n7112 & ~n28634 ;
  assign n29693 = ~n29687 & ~n29688 ;
  assign n29694 = ~n29689 & n29693 ;
  assign n29690 = ~n7164 & ~n28624 ;
  assign n29691 = ~n7156 & ~n28556 ;
  assign n29695 = ~n29690 & ~n29691 ;
  assign n29696 = n29694 & n29695 ;
  assign n29697 = ~n29670 & n29696 ;
  assign n29698 = ~n29692 & n29697 ;
  assign n29699 = ~n29686 & n29698 ;
  assign n29700 = ~n29308 & n29699 ;
  assign n29701 = ~n29682 & n29700 ;
  assign n29702 = ~n29675 & n29701 ;
  assign n29703 = n28719 & ~n29702 ;
  assign n29706 = n7340 & n28725 ;
  assign n29707 = n28725 & ~n28727 ;
  assign n29708 = \core_eu_em_mac_em_reg_myopwe_DO_reg[13]/P0001  & n28544 ;
  assign n29710 = n7186 & ~n28652 ;
  assign n29709 = n7194 & n28652 ;
  assign n29711 = ~n28660 & ~n29709 ;
  assign n29712 = ~n29710 & n29711 ;
  assign n29713 = n28739 & n29712 ;
  assign n29722 = ~n29708 & ~n29713 ;
  assign n29714 = n7198 & n28705 ;
  assign n29715 = n7190 & ~n28705 ;
  assign n29716 = ~n29714 & ~n29715 ;
  assign n29717 = n28735 & n29716 ;
  assign n29718 = ~\core_c_psq_MSTAT_reg_DO_reg[0]/P0002  & ~\core_eu_em_mac_em_reg_mfrwe_DO_reg[13]/P0001  ;
  assign n29719 = \core_c_psq_MSTAT_reg_DO_reg[0]/P0002  & ~\core_eu_em_mac_em_reg_mfswe_DO_reg[13]/P0001  ;
  assign n29720 = ~n29718 & ~n29719 ;
  assign n29721 = n28741 & n29720 ;
  assign n29723 = ~n29717 & ~n29721 ;
  assign n29724 = n29722 & n29723 ;
  assign n29725 = ~n29707 & ~n29724 ;
  assign n29705 = n12658 & n28729 ;
  assign n29726 = ~n28543 & ~n29705 ;
  assign n29727 = ~n29725 & n29726 ;
  assign n29728 = ~n29706 & n29727 ;
  assign n29704 = ~\core_eu_em_mac_em_reg_myopwe_DO_reg[13]/P0001  & n28543 ;
  assign n29729 = ~n28719 & ~n29704 ;
  assign n29730 = ~n29728 & n29729 ;
  assign n29731 = ~n29703 & ~n29730 ;
  assign n29734 = ~n14424 & n28561 ;
  assign n29733 = \core_c_dec_MTAR_E_reg/P0001  & n23757 ;
  assign n29735 = ~n28564 & ~n29733 ;
  assign n29736 = ~n29734 & n29735 ;
  assign n29737 = n28559 & ~n29736 ;
  assign n29738 = ~n8354 & ~n28594 ;
  assign n29739 = ~n8358 & ~n28589 ;
  assign n29740 = ~n29738 & ~n29739 ;
  assign n29741 = n29562 & n29740 ;
  assign n29742 = n28577 & ~n29741 ;
  assign n29743 = ~n29303 & ~n29742 ;
  assign n29744 = ~n28569 & ~n29743 ;
  assign n29842 = ~n8460 & n28572 ;
  assign n29841 = ~n12590 & ~n28572 ;
  assign n29843 = n28997 & ~n29841 ;
  assign n29844 = ~n29842 & n29843 ;
  assign n29779 = ~n8385 & ~n28634 ;
  assign n29746 = n12590 & n28619 ;
  assign n29778 = n8460 & n28630 ;
  assign n29845 = ~n29746 & ~n29778 ;
  assign n29846 = ~n29779 & n29845 ;
  assign n29732 = ~n8402 & ~n28624 ;
  assign n29745 = ~n8410 & ~n28556 ;
  assign n29847 = ~n29732 & ~n29745 ;
  assign n29848 = n29846 & n29847 ;
  assign n29748 = ~n17995 & n19792 ;
  assign n29758 = ~n18117 & ~n18918 ;
  assign n29756 = ~n17935 & ~n18914 ;
  assign n29757 = ~n18912 & ~n18991 ;
  assign n29762 = ~n29756 & ~n29757 ;
  assign n29763 = ~n29758 & n29762 ;
  assign n29753 = \core_c_dec_IRE_reg[11]/NET0131  & ~n8402 ;
  assign n29755 = ~n18189 & ~n18907 ;
  assign n29761 = ~n29753 & ~n29755 ;
  assign n29764 = n19874 & n29761 ;
  assign n29771 = n29763 & n29764 ;
  assign n29772 = ~n18085 & n19854 ;
  assign n29773 = n29771 & n29772 ;
  assign n29752 = n18099 & ~n19857 ;
  assign n29754 = n18162 & ~n18895 ;
  assign n29767 = ~n29752 & ~n29754 ;
  assign n29759 = n18740 & ~n18775 ;
  assign n29760 = ~n17998 & n18765 ;
  assign n29768 = ~n29759 & ~n29760 ;
  assign n29769 = n29767 & n29768 ;
  assign n29747 = n18745 & ~n18781 ;
  assign n29749 = ~n18102 & ~n18720 ;
  assign n29765 = ~n29747 & ~n29749 ;
  assign n29750 = n18088 & ~n18898 ;
  assign n29751 = n18124 & ~n19818 ;
  assign n29766 = ~n29750 & ~n29751 ;
  assign n29770 = n29765 & n29766 ;
  assign n29774 = n29769 & n29770 ;
  assign n29775 = n29773 & n29774 ;
  assign n29776 = n29748 & n29775 ;
  assign n29777 = n28636 & ~n29776 ;
  assign n29798 = n18790 & n19731 ;
  assign n29793 = n17945 & n18153 ;
  assign n29794 = n19996 & ~n29793 ;
  assign n29795 = n18076 & n29794 ;
  assign n29782 = n18162 & n18179 ;
  assign n29783 = n18124 & n18157 ;
  assign n29786 = ~n29782 & ~n29783 ;
  assign n29784 = n18107 & n18171 ;
  assign n29785 = n17915 & n18111 ;
  assign n29787 = ~n29784 & ~n29785 ;
  assign n29788 = n29786 & n29787 ;
  assign n29789 = ~n17931 & ~n29788 ;
  assign n29807 = ~n18108 & n18136 ;
  assign n29791 = ~n17935 & ~n18091 ;
  assign n29792 = n18147 & ~n18175 ;
  assign n29825 = ~n29791 & ~n29792 ;
  assign n29826 = ~n29807 & n29825 ;
  assign n29832 = n17984 & n29826 ;
  assign n29833 = ~n29789 & n29832 ;
  assign n29836 = n29795 & n29833 ;
  assign n29837 = n29798 & n29836 ;
  assign n29805 = n18088 & ~n19979 ;
  assign n29796 = n17945 & ~n18047 ;
  assign n29829 = n18041 & ~n29796 ;
  assign n29830 = ~n29805 & n29829 ;
  assign n29802 = ~n18167 & n18178 ;
  assign n29803 = n18103 & n18120 ;
  assign n29814 = ~n29802 & ~n29803 ;
  assign n29806 = n18132 & n18188 ;
  assign n29811 = n18106 & n18172 ;
  assign n29815 = ~n29806 & ~n29811 ;
  assign n29816 = n29814 & n29815 ;
  assign n29799 = \core_c_dec_IRE_reg[11]/NET0131  & ~n8410 ;
  assign n29812 = ~n18060 & ~n29799 ;
  assign n29780 = n17921 & ~n18117 ;
  assign n29800 = ~n18129 & n18158 ;
  assign n29813 = ~n29780 & ~n29800 ;
  assign n29817 = n29812 & n29813 ;
  assign n29823 = n29816 & n29817 ;
  assign n29781 = n18100 & ~n18121 ;
  assign n29790 = ~n18133 & n18184 ;
  assign n29824 = ~n29781 & ~n29790 ;
  assign n29827 = n29823 & n29824 ;
  assign n29810 = n18166 & n18179 ;
  assign n29808 = n18148 & ~n18175 ;
  assign n29809 = n17915 & n18116 ;
  assign n29820 = ~n29808 & ~n29809 ;
  assign n29821 = ~n29810 & n29820 ;
  assign n29797 = n18131 & n18188 ;
  assign n29818 = ~n18065 & ~n29797 ;
  assign n29801 = n18128 & n18157 ;
  assign n29804 = n18103 & n18119 ;
  assign n29819 = ~n29801 & ~n29804 ;
  assign n29822 = n29818 & n29819 ;
  assign n29828 = n29821 & n29822 ;
  assign n29831 = n29827 & n29828 ;
  assign n29834 = n29830 & n29831 ;
  assign n29835 = n19999 & n29834 ;
  assign n29838 = n18799 & n29835 ;
  assign n29839 = n29837 & n29838 ;
  assign n29840 = n28627 & ~n29839 ;
  assign n29849 = ~n29777 & ~n29840 ;
  assign n29850 = n29848 & n29849 ;
  assign n29851 = ~n29844 & n29850 ;
  assign n29852 = ~n29308 & n29851 ;
  assign n29853 = ~n29744 & n29852 ;
  assign n29854 = ~n29737 & n29853 ;
  assign n29855 = n28719 & ~n29854 ;
  assign n29858 = n8460 & n28725 ;
  assign n29859 = \core_eu_em_mac_em_reg_myopwe_DO_reg[11]/P0001  & n28544 ;
  assign n29861 = n8350 & ~n28652 ;
  assign n29860 = n8346 & n28652 ;
  assign n29862 = ~n28660 & ~n29860 ;
  assign n29863 = ~n29861 & n29862 ;
  assign n29864 = n28739 & n29863 ;
  assign n29873 = ~n29859 & ~n29864 ;
  assign n29865 = n8338 & n28705 ;
  assign n29866 = n8342 & ~n28705 ;
  assign n29867 = ~n29865 & ~n29866 ;
  assign n29868 = n28735 & n29867 ;
  assign n29869 = ~\core_c_psq_MSTAT_reg_DO_reg[0]/P0002  & ~\core_eu_em_mac_em_reg_mfrwe_DO_reg[11]/P0001  ;
  assign n29870 = \core_c_psq_MSTAT_reg_DO_reg[0]/P0002  & ~\core_eu_em_mac_em_reg_mfswe_DO_reg[11]/P0001  ;
  assign n29871 = ~n29869 & ~n29870 ;
  assign n29872 = n28741 & n29871 ;
  assign n29874 = ~n29868 & ~n29872 ;
  assign n29875 = n29873 & n29874 ;
  assign n29876 = ~n29707 & ~n29875 ;
  assign n29857 = n12590 & n28729 ;
  assign n29877 = ~n28543 & ~n29857 ;
  assign n29878 = ~n29876 & n29877 ;
  assign n29879 = ~n29858 & n29878 ;
  assign n29856 = ~\core_eu_em_mac_em_reg_myopwe_DO_reg[11]/P0001  & n28543 ;
  assign n29880 = ~n28719 & ~n29856 ;
  assign n29881 = ~n29879 & n29880 ;
  assign n29882 = ~n29855 & ~n29881 ;
  assign n29885 = ~n20053 & n28561 ;
  assign n29884 = \core_c_dec_MTAR_E_reg/P0001  & n19848 ;
  assign n29886 = ~n28564 & ~n29884 ;
  assign n29887 = ~n29885 & n29886 ;
  assign n29888 = n28559 & ~n29887 ;
  assign n29889 = ~n7753 & ~n28594 ;
  assign n29890 = ~n7737 & ~n28589 ;
  assign n29891 = ~n29889 & ~n29890 ;
  assign n29892 = n29562 & n29891 ;
  assign n29893 = n28577 & ~n29892 ;
  assign n29894 = ~n29303 & ~n29893 ;
  assign n29895 = ~n28569 & ~n29894 ;
  assign n29948 = ~n7859 & n28572 ;
  assign n29947 = ~n12556 & ~n28572 ;
  assign n29949 = n28997 & ~n29947 ;
  assign n29950 = ~n29948 & n29949 ;
  assign n29910 = ~n17980 & ~n19856 ;
  assign n29911 = n17945 & ~n29910 ;
  assign n29920 = n18158 & n18742 ;
  assign n29917 = n18089 & n18905 ;
  assign n29919 = \core_c_dec_IRE_reg[11]/NET0131  & ~n7809 ;
  assign n29922 = ~n29917 & ~n29919 ;
  assign n29923 = ~n29920 & n29922 ;
  assign n29924 = ~n18783 & n29923 ;
  assign n29930 = ~n29911 & n29924 ;
  assign n29916 = ~n17924 & ~n18149 ;
  assign n29918 = n18765 & ~n19979 ;
  assign n29931 = ~n29916 & ~n29918 ;
  assign n29932 = n29930 & n29931 ;
  assign n29921 = ~n18108 & ~n18915 ;
  assign n29908 = ~n17922 & ~n19864 ;
  assign n29909 = ~n18121 & n18752 ;
  assign n29927 = ~n29908 & ~n29909 ;
  assign n29928 = ~n29921 & n29927 ;
  assign n29898 = ~n18133 & ~n18919 ;
  assign n29905 = ~n18159 & n18741 ;
  assign n29925 = ~n29898 & ~n29905 ;
  assign n29906 = ~n18091 & n18749 ;
  assign n29907 = ~n18180 & n18746 ;
  assign n29926 = ~n29906 & ~n29907 ;
  assign n29929 = n29925 & n29926 ;
  assign n29933 = n29928 & n29929 ;
  assign n29936 = n29932 & n29933 ;
  assign n29912 = ~n17981 & ~n18719 ;
  assign n29913 = n17839 & ~n29912 ;
  assign n29914 = ~n18046 & ~n29913 ;
  assign n29915 = ~n17938 & ~n29914 ;
  assign n29937 = n19997 & ~n29915 ;
  assign n29938 = n29936 & n29937 ;
  assign n29899 = ~n18123 & ~n18180 ;
  assign n29900 = n18099 & n18157 ;
  assign n29901 = n18090 & n18111 ;
  assign n29902 = ~n29900 & ~n29901 ;
  assign n29903 = ~n29899 & n29902 ;
  assign n29904 = n17931 & ~n29903 ;
  assign n29934 = n18042 & n29579 ;
  assign n29935 = ~n29904 & n29934 ;
  assign n29939 = n19716 & n29935 ;
  assign n29940 = n29798 & n29939 ;
  assign n29941 = n29938 & n29940 ;
  assign n29942 = n18800 & n29941 ;
  assign n29943 = n28627 & ~n29942 ;
  assign n29946 = n12556 & n28619 ;
  assign n29883 = ~n7784 & ~n28634 ;
  assign n29896 = n7859 & n28630 ;
  assign n29951 = ~n29883 & ~n29896 ;
  assign n29952 = ~n29946 & n29951 ;
  assign n29945 = ~n7809 & ~n28556 ;
  assign n29897 = ~n19895 & n28636 ;
  assign n29944 = ~n7801 & ~n28624 ;
  assign n29953 = ~n29897 & ~n29944 ;
  assign n29954 = ~n29945 & n29953 ;
  assign n29955 = n29952 & n29954 ;
  assign n29956 = ~n29943 & n29955 ;
  assign n29957 = ~n29950 & n29956 ;
  assign n29958 = ~n29308 & n29957 ;
  assign n29959 = ~n29895 & n29958 ;
  assign n29960 = ~n29888 & n29959 ;
  assign n29961 = n28719 & ~n29960 ;
  assign n29963 = n12556 & ~n28728 ;
  assign n29964 = ~\core_c_psq_MSTAT_reg_DO_reg[0]/P0002  & ~\core_eu_em_mac_em_reg_mfrwe_DO_reg[10]/P0001  ;
  assign n29965 = \core_c_psq_MSTAT_reg_DO_reg[0]/P0002  & ~\core_eu_em_mac_em_reg_mfswe_DO_reg[10]/P0001  ;
  assign n29966 = ~n29964 & ~n29965 ;
  assign n29967 = n28741 & n29966 ;
  assign n29977 = \core_eu_em_mac_em_reg_myopwe_DO_reg[10]/P0001  & ~n28545 ;
  assign n29978 = ~n29967 & ~n29977 ;
  assign n29969 = n7741 & ~n28652 ;
  assign n29968 = n7757 & n28652 ;
  assign n29970 = ~n28660 & ~n29968 ;
  assign n29971 = ~n29969 & n29970 ;
  assign n29972 = n28739 & n29971 ;
  assign n29973 = n7745 & n28705 ;
  assign n29974 = n7749 & ~n28705 ;
  assign n29975 = ~n29973 & ~n29974 ;
  assign n29976 = n28735 & n29975 ;
  assign n29979 = ~n29972 & ~n29976 ;
  assign n29980 = n29978 & n29979 ;
  assign n29981 = ~n28725 & n29980 ;
  assign n29982 = ~n29963 & n29981 ;
  assign n29962 = ~n7859 & n29643 ;
  assign n29983 = ~\core_eu_em_mac_em_reg_myopwe_DO_reg[10]/P0001  & n28543 ;
  assign n29984 = ~n28719 & ~n29983 ;
  assign n29985 = ~n29962 & n29984 ;
  assign n29986 = ~n29982 & n29985 ;
  assign n29987 = ~n29961 & ~n29986 ;
  assign n29988 = n19504 & n28660 ;
  assign n29989 = ~n29653 & ~n29988 ;
  assign n29990 = ~n28649 & ~n29989 ;
  assign n29991 = \core_eu_em_mac_em_reg_mxopwe_DO_reg[9]/P0001  & n28649 ;
  assign n29992 = ~n29990 & ~n29991 ;
  assign n29993 = ~n28550 & ~n29992 ;
  assign n29994 = n28550 & ~n29641 ;
  assign n29995 = ~n29993 & ~n29994 ;
  assign n29996 = n17836 & n28660 ;
  assign n29997 = ~n29712 & ~n29996 ;
  assign n29998 = ~n28649 & ~n29997 ;
  assign n29999 = \core_eu_em_mac_em_reg_mxopwe_DO_reg[13]/P0001  & n28649 ;
  assign n30000 = ~n29998 & ~n29999 ;
  assign n30001 = ~n28550 & ~n30000 ;
  assign n30002 = n28550 & ~n29702 ;
  assign n30003 = ~n30001 & ~n30002 ;
  assign n30004 = n23757 & n28660 ;
  assign n30005 = ~n29863 & ~n30004 ;
  assign n30006 = ~n28649 & ~n30005 ;
  assign n30007 = \core_eu_em_mac_em_reg_mxopwe_DO_reg[11]/P0001  & n28649 ;
  assign n30008 = ~n30006 & ~n30007 ;
  assign n30009 = ~n28550 & ~n30008 ;
  assign n30010 = n28550 & ~n29854 ;
  assign n30011 = ~n30009 & ~n30010 ;
  assign n30012 = n19848 & n28660 ;
  assign n30013 = ~n29971 & ~n30012 ;
  assign n30014 = ~n28649 & ~n30013 ;
  assign n30015 = \core_eu_em_mac_em_reg_mxopwe_DO_reg[10]/P0001  & n28649 ;
  assign n30016 = ~n30014 & ~n30015 ;
  assign n30017 = ~n28550 & ~n30016 ;
  assign n30018 = n28550 & ~n29960 ;
  assign n30019 = ~n30017 & ~n30018 ;
  assign n30021 = n9178 & n28725 ;
  assign n30020 = n12624 & n28729 ;
  assign n30031 = ~\core_c_psq_MSTAT_reg_DO_reg[0]/P0002  & ~\core_eu_em_mac_em_reg_mfrwe_DO_reg[12]/P0001  ;
  assign n30032 = \core_c_psq_MSTAT_reg_DO_reg[0]/P0002  & ~\core_eu_em_mac_em_reg_mfswe_DO_reg[12]/P0001  ;
  assign n30033 = ~n30031 & ~n30032 ;
  assign n30034 = n28741 & n30033 ;
  assign n30022 = n9064 & n28705 ;
  assign n30023 = n9068 & ~n28705 ;
  assign n30024 = ~n30022 & ~n30023 ;
  assign n30025 = n28735 & n30024 ;
  assign n30027 = n9060 & ~n28652 ;
  assign n30026 = n9076 & n28652 ;
  assign n30028 = ~n28660 & ~n30026 ;
  assign n30029 = ~n30027 & n30028 ;
  assign n30030 = n28739 & n30029 ;
  assign n30035 = ~n30025 & ~n30030 ;
  assign n30036 = ~n30034 & n30035 ;
  assign n30037 = ~n30020 & n30036 ;
  assign n30038 = ~n30021 & n30037 ;
  assign n30039 = ~n28543 & ~n30038 ;
  assign n30040 = \core_eu_em_mac_em_reg_myopwe_DO_reg[12]/P0001  & ~n28545 ;
  assign n30041 = ~n28719 & ~n30040 ;
  assign n30042 = ~n30039 & n30041 ;
  assign n30092 = ~n14413 & n28561 ;
  assign n30091 = \core_c_dec_MTAR_E_reg/P0001  & n23920 ;
  assign n30093 = ~n28564 & ~n30091 ;
  assign n30094 = ~n30092 & n30093 ;
  assign n30095 = n28559 & ~n30094 ;
  assign n30096 = ~n9072 & ~n28594 ;
  assign n30097 = ~n9056 & ~n28589 ;
  assign n30098 = ~n30096 & ~n30097 ;
  assign n30099 = n29562 & n30098 ;
  assign n30100 = n28577 & ~n30099 ;
  assign n30101 = ~n29303 & ~n30100 ;
  assign n30102 = ~n28569 & ~n30101 ;
  assign n30104 = ~n9178 & n28572 ;
  assign n30103 = ~n12624 & ~n28572 ;
  assign n30105 = n28997 & ~n30103 ;
  assign n30106 = ~n30104 & n30105 ;
  assign n30109 = n9178 & n28630 ;
  assign n30107 = ~n9103 & ~n28634 ;
  assign n30108 = n12624 & n28619 ;
  assign n30144 = ~n30107 & ~n30108 ;
  assign n30145 = ~n30109 & n30144 ;
  assign n30110 = ~n9120 & ~n28624 ;
  assign n30111 = ~n9128 & ~n28556 ;
  assign n30146 = ~n30110 & ~n30111 ;
  assign n30147 = n30145 & n30146 ;
  assign n30055 = ~n17998 & n18088 ;
  assign n30056 = n18162 & ~n18781 ;
  assign n30081 = ~n30055 & ~n30056 ;
  assign n30061 = ~n18170 & n20996 ;
  assign n30062 = ~n18182 & n20104 ;
  assign n30082 = ~n30061 & ~n30062 ;
  assign n30083 = n30081 & n30082 ;
  assign n30043 = n18191 & n18905 ;
  assign n30059 = \core_c_dec_IRE_reg[11]/NET0131  & ~n9120 ;
  assign n30065 = ~n30043 & ~n30059 ;
  assign n30054 = n18055 & ~n20096 ;
  assign n30057 = n17986 & n18752 ;
  assign n30066 = ~n30054 & ~n30057 ;
  assign n30069 = n30065 & n30066 ;
  assign n30058 = n18039 & ~n19870 ;
  assign n30070 = ~n17969 & ~n30058 ;
  assign n30071 = n30069 & n30070 ;
  assign n30064 = n18153 & n18741 ;
  assign n30060 = n18191 & n18749 ;
  assign n30063 = n18056 & n18756 ;
  assign n30067 = ~n30060 & ~n30063 ;
  assign n30068 = ~n30064 & n30067 ;
  assign n30072 = n19812 & n30068 ;
  assign n30079 = n30071 & n30072 ;
  assign n30052 = ~n17924 & n19808 ;
  assign n30053 = n18099 & ~n18720 ;
  assign n30080 = ~n30052 & ~n30053 ;
  assign n30084 = n30079 & n30080 ;
  assign n30048 = n18071 & n18124 ;
  assign n30049 = n18187 & n18893 ;
  assign n30075 = ~n30048 & ~n30049 ;
  assign n30050 = n18070 & n18740 ;
  assign n30051 = n18043 & n18751 ;
  assign n30076 = ~n30050 & ~n30051 ;
  assign n30077 = n30075 & n30076 ;
  assign n30044 = n18766 & ~n18914 ;
  assign n30045 = ~n18912 & n19862 ;
  assign n30073 = ~n30044 & ~n30045 ;
  assign n30046 = n18759 & ~n18907 ;
  assign n30047 = n18139 & n18745 ;
  assign n30074 = ~n30046 & ~n30047 ;
  assign n30078 = n30073 & n30074 ;
  assign n30085 = n30077 & n30078 ;
  assign n30086 = n30084 & n30085 ;
  assign n30087 = n30083 & n30086 ;
  assign n30088 = n19791 & n30087 ;
  assign n30089 = n29748 & n30088 ;
  assign n30090 = n28636 & ~n30089 ;
  assign n30123 = ~n18121 & ~n18743 ;
  assign n30120 = ~n18159 & ~n20096 ;
  assign n30122 = ~n18091 & n18766 ;
  assign n30128 = ~n30120 & ~n30122 ;
  assign n30129 = ~n30123 & n30128 ;
  assign n30135 = ~n18085 & n30129 ;
  assign n30136 = n29579 & n30135 ;
  assign n30139 = n18064 & n30136 ;
  assign n30140 = n29795 & n30139 ;
  assign n30124 = ~n17924 & n18176 ;
  assign n30113 = n17945 & ~n18152 ;
  assign n30116 = ~n17938 & ~n18149 ;
  assign n30132 = ~n30113 & ~n30116 ;
  assign n30133 = ~n30124 & n30132 ;
  assign n30115 = ~n18180 & ~n18919 ;
  assign n30117 = ~n17922 & ~n19870 ;
  assign n30126 = ~n30115 & ~n30117 ;
  assign n30118 = ~n18096 & n18752 ;
  assign n30119 = ~n18108 & n19862 ;
  assign n30127 = ~n30118 & ~n30119 ;
  assign n30130 = n30126 & n30127 ;
  assign n30112 = ~n18170 & n19717 ;
  assign n30114 = ~n18133 & ~n18915 ;
  assign n30121 = \core_c_dec_IRE_reg[11]/NET0131  & ~n9128 ;
  assign n30125 = ~n30114 & ~n30121 ;
  assign n30131 = ~n30112 & n30125 ;
  assign n30134 = n30130 & n30131 ;
  assign n30137 = n30133 & n30134 ;
  assign n30138 = n17988 & n30137 ;
  assign n30141 = n20159 & n30138 ;
  assign n30142 = n30140 & n30141 ;
  assign n30143 = n28627 & ~n30142 ;
  assign n30148 = ~n30090 & ~n30143 ;
  assign n30149 = n30147 & n30148 ;
  assign n30150 = ~n30106 & n30149 ;
  assign n30151 = ~n29308 & n30150 ;
  assign n30152 = ~n30102 & n30151 ;
  assign n30153 = ~n30095 & n30152 ;
  assign n30154 = n28719 & n30153 ;
  assign n30155 = ~n30042 & ~n30154 ;
  assign n30156 = n23920 & n28660 ;
  assign n30157 = ~n30029 & ~n30156 ;
  assign n30158 = ~n28649 & ~n30157 ;
  assign n30159 = \core_eu_em_mac_em_reg_mxopwe_DO_reg[12]/P0001  & n28649 ;
  assign n30160 = ~n30158 & ~n30159 ;
  assign n30161 = ~n28550 & ~n30160 ;
  assign n30162 = n28550 & ~n30153 ;
  assign n30163 = ~n30161 & ~n30162 ;
  assign n30165 = n11265 & n28725 ;
  assign n30164 = n13006 & n28729 ;
  assign n30175 = ~\core_c_psq_MSTAT_reg_DO_reg[0]/P0002  & ~\core_eu_em_mac_em_reg_mfrwe_DO_reg[7]/P0001  ;
  assign n30176 = \core_c_psq_MSTAT_reg_DO_reg[0]/P0002  & ~\core_eu_em_mac_em_reg_mfswe_DO_reg[7]/P0001  ;
  assign n30177 = ~n30175 & ~n30176 ;
  assign n30178 = n28741 & n30177 ;
  assign n30166 = n11176 & n28705 ;
  assign n30167 = n11180 & ~n28705 ;
  assign n30168 = ~n30166 & ~n30167 ;
  assign n30169 = n28735 & n30168 ;
  assign n30171 = n11188 & ~n28652 ;
  assign n30170 = n11184 & n28652 ;
  assign n30172 = ~n28660 & ~n30170 ;
  assign n30173 = ~n30171 & n30172 ;
  assign n30174 = n28739 & n30173 ;
  assign n30179 = ~n30169 & ~n30174 ;
  assign n30180 = ~n30178 & n30179 ;
  assign n30181 = ~n30164 & n30180 ;
  assign n30182 = ~n30165 & n30181 ;
  assign n30183 = ~n28543 & ~n30182 ;
  assign n30184 = \core_eu_em_mac_em_reg_myopwe_DO_reg[7]/P0001  & ~n28545 ;
  assign n30185 = ~n28719 & ~n30184 ;
  assign n30186 = ~n30183 & n30185 ;
  assign n30189 = ~n23253 & n28561 ;
  assign n30188 = \core_c_dec_MTAR_E_reg/P0001  & n19972 ;
  assign n30190 = ~n28564 & ~n30188 ;
  assign n30191 = ~n30189 & n30190 ;
  assign n30192 = n28559 & ~n30191 ;
  assign n30193 = ~n11192 & ~n28594 ;
  assign n30194 = ~n11196 & ~n28589 ;
  assign n30195 = ~n30193 & ~n30194 ;
  assign n30196 = n29562 & n30195 ;
  assign n30197 = n28577 & ~n30196 ;
  assign n30198 = ~n29303 & ~n30197 ;
  assign n30199 = ~n28569 & ~n30198 ;
  assign n30201 = ~n13006 & ~n28572 ;
  assign n30200 = ~n11265 & n28572 ;
  assign n30202 = n28997 & ~n30200 ;
  assign n30203 = ~n30201 & n30202 ;
  assign n30249 = ~n11239 & ~n28556 ;
  assign n30204 = ~n11231 & ~n28624 ;
  assign n30212 = \core_c_dec_IRE_reg[11]/NET0131  & ~n11231 ;
  assign n30214 = n18001 & n18125 ;
  assign n30224 = ~n30212 & ~n30214 ;
  assign n30215 = n18188 & n18191 ;
  assign n30218 = n18056 & n18103 ;
  assign n30225 = ~n30215 & ~n30218 ;
  assign n30226 = n30224 & n30225 ;
  assign n30210 = n18039 & n18188 ;
  assign n30227 = ~n18018 & ~n30210 ;
  assign n30228 = n30226 & n30227 ;
  assign n30229 = n18902 & n19812 ;
  assign n30236 = n30228 & n30229 ;
  assign n30206 = n18111 & ~n18898 ;
  assign n30207 = ~n18165 & n20996 ;
  assign n30237 = ~n30206 & ~n30207 ;
  assign n30240 = n30236 & n30237 ;
  assign n30220 = n18163 & ~n18912 ;
  assign n30221 = n18184 & ~n18918 ;
  assign n30232 = ~n30220 & ~n30221 ;
  assign n30222 = n17980 & n18751 ;
  assign n30223 = ~n18909 & n19720 ;
  assign n30233 = ~n30222 & ~n30223 ;
  assign n30234 = n30232 & n30233 ;
  assign n30208 = ~n18914 & ~n18991 ;
  assign n30209 = ~n17935 & ~n18079 ;
  assign n30230 = ~n30208 & ~n30209 ;
  assign n30213 = n18124 & n19801 ;
  assign n30219 = n18128 & ~n18907 ;
  assign n30231 = ~n30213 & ~n30219 ;
  assign n30235 = n30230 & n30231 ;
  assign n30241 = n30234 & n30235 ;
  assign n30242 = n30240 & n30241 ;
  assign n30217 = ~n17998 & n18115 ;
  assign n30211 = ~n18175 & n18922 ;
  assign n30216 = n18099 & ~n18895 ;
  assign n30238 = ~n30211 & ~n30216 ;
  assign n30239 = ~n30217 & n30238 ;
  assign n30243 = n18790 & n30239 ;
  assign n30244 = n18892 & n30243 ;
  assign n30245 = n30242 & n30244 ;
  assign n30246 = n28636 & ~n30245 ;
  assign n30252 = ~n30204 & ~n30246 ;
  assign n30253 = ~n30249 & n30252 ;
  assign n30187 = ~n20030 & n28627 ;
  assign n30248 = ~n11062 & ~n28634 ;
  assign n30205 = n11265 & n28630 ;
  assign n30247 = n13006 & n28619 ;
  assign n30250 = ~n30205 & ~n30247 ;
  assign n30251 = ~n30248 & n30250 ;
  assign n30254 = ~n30187 & n30251 ;
  assign n30255 = n30253 & n30254 ;
  assign n30256 = ~n30203 & n30255 ;
  assign n30257 = ~n29308 & n30256 ;
  assign n30258 = ~n30199 & n30257 ;
  assign n30259 = ~n30192 & n30258 ;
  assign n30260 = n28719 & n30259 ;
  assign n30261 = ~n30186 & ~n30260 ;
  assign n30262 = \sport1_regs_FSDIVreg_DO_reg[14]/NET0131  & n28786 ;
  assign n30263 = ~\sport1_cfg_FSi_cnt_reg[14]/NET0131  & ~n28869 ;
  assign n30264 = n28855 & ~n28870 ;
  assign n30265 = ~n30263 & n30264 ;
  assign n30266 = ~n30262 & ~n30265 ;
  assign n30267 = n12715 & n28729 ;
  assign n30268 = n12688 & n28725 ;
  assign n30278 = ~\core_c_psq_MSTAT_reg_DO_reg[0]/P0002  & ~\core_eu_em_mac_em_reg_mfrwe_DO_reg[14]/P0001  ;
  assign n30279 = \core_c_psq_MSTAT_reg_DO_reg[0]/P0002  & ~\core_eu_em_mac_em_reg_mfswe_DO_reg[14]/P0001  ;
  assign n30280 = ~n30278 & ~n30279 ;
  assign n30281 = n28741 & n30280 ;
  assign n30269 = n11862 & n28705 ;
  assign n30270 = n11866 & ~n28705 ;
  assign n30271 = ~n30269 & ~n30270 ;
  assign n30272 = n28735 & n30271 ;
  assign n30274 = n11874 & ~n28652 ;
  assign n30273 = n11870 & n28652 ;
  assign n30275 = ~n28660 & ~n30273 ;
  assign n30276 = ~n30274 & n30275 ;
  assign n30277 = n28739 & n30276 ;
  assign n30282 = ~n30272 & ~n30277 ;
  assign n30283 = ~n30281 & n30282 ;
  assign n30284 = ~n30268 & n30283 ;
  assign n30285 = ~n30267 & n30284 ;
  assign n30286 = ~n28543 & ~n30285 ;
  assign n30287 = \core_eu_em_mac_em_reg_myopwe_DO_reg[14]/P0001  & ~n28545 ;
  assign n30288 = ~n28719 & ~n30287 ;
  assign n30289 = ~n30286 & n30288 ;
  assign n30292 = n14540 & n28561 ;
  assign n30291 = \core_c_dec_MTAR_E_reg/P0001  & n20150 ;
  assign n30293 = ~n28564 & ~n30291 ;
  assign n30294 = ~n30292 & n30293 ;
  assign n30295 = n28559 & ~n30294 ;
  assign n30296 = ~n11878 & ~n28594 ;
  assign n30297 = ~n11882 & ~n28589 ;
  assign n30298 = ~n30296 & ~n30297 ;
  assign n30299 = n29562 & n30298 ;
  assign n30300 = n28577 & ~n30299 ;
  assign n30301 = ~n29303 & ~n30300 ;
  assign n30302 = ~n28569 & ~n30301 ;
  assign n30310 = ~n12688 & n28572 ;
  assign n30309 = ~n12715 & ~n28572 ;
  assign n30311 = n28997 & ~n30309 ;
  assign n30312 = ~n30310 & n30311 ;
  assign n30308 = ~n21226 & n28636 ;
  assign n30290 = ~n20192 & n28627 ;
  assign n30305 = n12715 & n28619 ;
  assign n30303 = ~n11837 & ~n28634 ;
  assign n30304 = n12688 & n28630 ;
  assign n30313 = ~n30303 & ~n30304 ;
  assign n30314 = ~n30305 & n30313 ;
  assign n30306 = ~n11854 & ~n28556 ;
  assign n30307 = ~n11846 & ~n28624 ;
  assign n30315 = ~n30306 & ~n30307 ;
  assign n30316 = n30314 & n30315 ;
  assign n30317 = ~n30290 & n30316 ;
  assign n30318 = ~n30308 & n30317 ;
  assign n30319 = ~n30312 & n30318 ;
  assign n30320 = ~n29308 & n30319 ;
  assign n30321 = ~n30302 & n30320 ;
  assign n30322 = ~n30295 & n30321 ;
  assign n30323 = n28719 & n30322 ;
  assign n30324 = ~n30289 & ~n30323 ;
  assign n30325 = \sport0_regs_FSDIVreg_DO_reg[14]/NET0131  & n28876 ;
  assign n30326 = ~\sport0_cfg_FSi_cnt_reg[14]/NET0131  & ~n28959 ;
  assign n30327 = n28945 & ~n28960 ;
  assign n30328 = ~n30326 & n30327 ;
  assign n30329 = ~n30325 & ~n30328 ;
  assign n30330 = n19972 & n28660 ;
  assign n30331 = ~n30173 & ~n30330 ;
  assign n30332 = ~n28649 & ~n30331 ;
  assign n30333 = \core_eu_em_mac_em_reg_mxopwe_DO_reg[7]/P0001  & n28649 ;
  assign n30334 = ~n30332 & ~n30333 ;
  assign n30335 = ~n28550 & ~n30334 ;
  assign n30336 = n28550 & ~n30259 ;
  assign n30337 = ~n30335 & ~n30336 ;
  assign n30338 = n20150 & n28660 ;
  assign n30339 = ~n30276 & ~n30338 ;
  assign n30340 = ~n28649 & ~n30339 ;
  assign n30341 = \core_eu_em_mac_em_reg_mxopwe_DO_reg[14]/P0001  & n28649 ;
  assign n30342 = ~n30340 & ~n30341 ;
  assign n30343 = ~n28550 & ~n30342 ;
  assign n30344 = n28550 & ~n30322 ;
  assign n30345 = ~n30343 & ~n30344 ;
  assign n30395 = ~n14658 & n28561 ;
  assign n30394 = \core_c_dec_MTAR_E_reg/P0001  & n23860 ;
  assign n30396 = ~n28564 & ~n30394 ;
  assign n30397 = ~n30395 & n30396 ;
  assign n30398 = n28559 & ~n30397 ;
  assign n30399 = ~n10534 & ~n28594 ;
  assign n30400 = ~n10538 & ~n28589 ;
  assign n30401 = ~n30399 & ~n30400 ;
  assign n30402 = n29562 & n30401 ;
  assign n30403 = n28577 & ~n30402 ;
  assign n30404 = ~n29303 & ~n30403 ;
  assign n30405 = ~n28569 & ~n30404 ;
  assign n30407 = ~n10638 & n28572 ;
  assign n30406 = ~n13041 & ~n28572 ;
  assign n30408 = n28997 & ~n30406 ;
  assign n30409 = ~n30407 & n30408 ;
  assign n30355 = ~n18091 & n19862 ;
  assign n30356 = ~n18108 & n18756 ;
  assign n30373 = ~n30355 & ~n30356 ;
  assign n30359 = ~n18133 & ~n20096 ;
  assign n30360 = n18043 & n18748 ;
  assign n30374 = ~n30359 & ~n30360 ;
  assign n30377 = n30373 & n30374 ;
  assign n30347 = ~n18170 & n18732 ;
  assign n30371 = ~n18140 & ~n30347 ;
  assign n30353 = ~n18180 & ~n18743 ;
  assign n30354 = ~n18159 & n18752 ;
  assign n30372 = ~n30353 & ~n30354 ;
  assign n30378 = n30371 & n30372 ;
  assign n30385 = n30377 & n30378 ;
  assign n30363 = ~n17922 & ~n18915 ;
  assign n30361 = n18070 & n18765 ;
  assign n30362 = ~n18110 & n18147 ;
  assign n30375 = ~n30361 & ~n30362 ;
  assign n30376 = ~n30363 & n30375 ;
  assign n30386 = ~n18085 & n30376 ;
  assign n30387 = n30385 & n30386 ;
  assign n30346 = ~n18161 & n19717 ;
  assign n30381 = n29052 & ~n30346 ;
  assign n30350 = n17925 & ~n29063 ;
  assign n30351 = n18088 & ~n18775 ;
  assign n30382 = ~n30350 & ~n30351 ;
  assign n30383 = n30381 & n30382 ;
  assign n30352 = ~n17924 & n18719 ;
  assign n30348 = n18748 & n18761 ;
  assign n30368 = ~n18058 & ~n30348 ;
  assign n30369 = ~n30352 & n30368 ;
  assign n30349 = n18089 & n19863 ;
  assign n30358 = \core_c_dec_IRE_reg[11]/NET0131  & ~n10575 ;
  assign n30365 = ~n30349 & ~n30358 ;
  assign n30357 = n17986 & n18905 ;
  assign n30364 = n18153 & n18766 ;
  assign n30366 = ~n30357 & ~n30364 ;
  assign n30367 = n30365 & n30366 ;
  assign n30370 = ~n18069 & n30367 ;
  assign n30379 = n30369 & n30370 ;
  assign n30380 = n18041 & ~n19991 ;
  assign n30384 = n30379 & n30380 ;
  assign n30388 = n30383 & n30384 ;
  assign n30389 = n18726 & n30388 ;
  assign n30390 = n30387 & n30389 ;
  assign n30391 = n19977 & n30390 ;
  assign n30392 = n29047 & n30391 ;
  assign n30393 = n28627 & ~n30392 ;
  assign n30445 = ~n10461 & ~n28634 ;
  assign n30443 = n10638 & n28630 ;
  assign n30444 = n13041 & n28619 ;
  assign n30448 = ~n30443 & ~n30444 ;
  assign n30449 = ~n30445 & n30448 ;
  assign n30447 = ~n10567 & ~n28624 ;
  assign n30413 = ~n18098 & ~n18781 ;
  assign n30414 = n18751 & ~n19818 ;
  assign n30432 = ~n30413 & ~n30414 ;
  assign n30415 = ~n18170 & n19808 ;
  assign n30416 = ~n18182 & n19785 ;
  assign n30433 = ~n30415 & ~n30416 ;
  assign n30436 = n30432 & n30433 ;
  assign n30427 = n18763 & ~n18907 ;
  assign n30417 = ~n18912 & ~n18919 ;
  assign n30410 = n17952 & n18746 ;
  assign n30420 = \core_c_dec_IRE_reg[11]/NET0131  & ~n10567 ;
  assign n30428 = ~n30410 & ~n30420 ;
  assign n30429 = ~n30417 & n30428 ;
  assign n30430 = ~n30427 & n30429 ;
  assign n30411 = n18748 & ~n18898 ;
  assign n30412 = n18740 & ~n18895 ;
  assign n30431 = ~n30411 & ~n30412 ;
  assign n30437 = n30430 & n30431 ;
  assign n30438 = n30436 & n30437 ;
  assign n30421 = n18001 & n18745 ;
  assign n30422 = ~n18037 & ~n30421 ;
  assign n30423 = ~n29533 & n30422 ;
  assign n30424 = n29536 & n30423 ;
  assign n30425 = ~n17931 & ~n30424 ;
  assign n30426 = ~n17924 & n18080 ;
  assign n30418 = ~n17938 & n18922 ;
  assign n30419 = ~n17998 & n18111 ;
  assign n30434 = ~n30418 & ~n30419 ;
  assign n30435 = ~n30426 & n30434 ;
  assign n30439 = ~n30425 & n30435 ;
  assign n30440 = n30438 & n30439 ;
  assign n30441 = n29522 & n30440 ;
  assign n30442 = n28636 & ~n30441 ;
  assign n30446 = ~n10575 & ~n28556 ;
  assign n30450 = ~n30442 & ~n30446 ;
  assign n30451 = ~n30447 & n30450 ;
  assign n30452 = n30449 & n30451 ;
  assign n30453 = ~n30393 & n30452 ;
  assign n30454 = ~n30409 & n30453 ;
  assign n30455 = ~n29308 & n30454 ;
  assign n30456 = ~n30405 & n30455 ;
  assign n30457 = ~n30398 & n30456 ;
  assign n30458 = n28719 & ~n30457 ;
  assign n30461 = n10638 & n28725 ;
  assign n30462 = \core_eu_em_mac_em_reg_myopwe_DO_reg[8]/P0001  & n28544 ;
  assign n30464 = n10530 & ~n28652 ;
  assign n30463 = n10526 & n28652 ;
  assign n30465 = ~n28660 & ~n30463 ;
  assign n30466 = ~n30464 & n30465 ;
  assign n30467 = n28739 & n30466 ;
  assign n30476 = ~n30462 & ~n30467 ;
  assign n30468 = n10518 & n28705 ;
  assign n30469 = n10522 & ~n28705 ;
  assign n30470 = ~n30468 & ~n30469 ;
  assign n30471 = n28735 & n30470 ;
  assign n30472 = ~\core_c_psq_MSTAT_reg_DO_reg[0]/P0002  & ~\core_eu_em_mac_em_reg_mfrwe_DO_reg[8]/P0001  ;
  assign n30473 = \core_c_psq_MSTAT_reg_DO_reg[0]/P0002  & ~\core_eu_em_mac_em_reg_mfswe_DO_reg[8]/P0001  ;
  assign n30474 = ~n30472 & ~n30473 ;
  assign n30475 = n28741 & n30474 ;
  assign n30477 = ~n30471 & ~n30475 ;
  assign n30478 = n30476 & n30477 ;
  assign n30479 = ~n29707 & ~n30478 ;
  assign n30460 = n13041 & n28729 ;
  assign n30480 = ~n28543 & ~n30460 ;
  assign n30481 = ~n30479 & n30480 ;
  assign n30482 = ~n30461 & n30481 ;
  assign n30459 = ~\core_eu_em_mac_em_reg_myopwe_DO_reg[8]/P0001  & n28543 ;
  assign n30483 = ~n28719 & ~n30459 ;
  assign n30484 = ~n30482 & n30483 ;
  assign n30485 = ~n30458 & ~n30484 ;
  assign n30486 = n23860 & n28660 ;
  assign n30487 = ~n30466 & ~n30486 ;
  assign n30488 = ~n28649 & ~n30487 ;
  assign n30489 = \core_eu_em_mac_em_reg_mxopwe_DO_reg[8]/P0001  & n28649 ;
  assign n30490 = ~n30488 & ~n30489 ;
  assign n30491 = ~n28550 & ~n30490 ;
  assign n30492 = n28550 & ~n30457 ;
  assign n30493 = ~n30491 & ~n30492 ;
  assign n30494 = ~n14610 & n28561 ;
  assign n30495 = \core_c_dec_MTAR_E_reg/P0001  & n21663 ;
  assign n30496 = ~n28564 & ~n30495 ;
  assign n30497 = ~n30494 & n30496 ;
  assign n30498 = n28559 & ~n30497 ;
  assign n30505 = ~n8113 & n28577 ;
  assign n30504 = ~n12870 & ~n28577 ;
  assign n30506 = ~n28575 & ~n30504 ;
  assign n30507 = ~n30505 & n30506 ;
  assign n30508 = ~n28576 & ~n30507 ;
  assign n30509 = n28569 & ~n30508 ;
  assign n30515 = ~n7885 & ~n28589 ;
  assign n30513 = ~n7905 & ~n28598 ;
  assign n30514 = ~n7909 & ~n28594 ;
  assign n30516 = ~n30513 & ~n30514 ;
  assign n30517 = ~n30515 & n30516 ;
  assign n30518 = n28607 & n30517 ;
  assign n30519 = n28572 & n30518 ;
  assign n30512 = ~n8113 & ~n28572 ;
  assign n30520 = n28584 & ~n30512 ;
  assign n30521 = ~n30519 & n30520 ;
  assign n30501 = ~n21700 & n28627 ;
  assign n30499 = ~n21958 & n28636 ;
  assign n30500 = n8113 & n28630 ;
  assign n30522 = ~n30499 & ~n30500 ;
  assign n30510 = ~n7952 & ~n28634 ;
  assign n30511 = n12870 & n28619 ;
  assign n30523 = ~n30510 & ~n30511 ;
  assign n30524 = n30522 & n30523 ;
  assign n30502 = ~n7987 & ~n28624 ;
  assign n30503 = ~n7991 & ~n28556 ;
  assign n30525 = ~n30502 & ~n30503 ;
  assign n30526 = n30524 & n30525 ;
  assign n30527 = ~n30501 & n30526 ;
  assign n30528 = ~n30521 & n30527 ;
  assign n30529 = ~n30509 & n30528 ;
  assign n30530 = ~n30498 & n30529 ;
  assign n30531 = n28550 & ~n30530 ;
  assign n30537 = n21663 & n28660 ;
  assign n30534 = n7901 & ~n28652 ;
  assign n30533 = n7889 & n28652 ;
  assign n30535 = ~n28660 & ~n30533 ;
  assign n30536 = ~n30534 & n30535 ;
  assign n30538 = ~n28649 & ~n30536 ;
  assign n30539 = ~n30537 & n30538 ;
  assign n30532 = ~\core_eu_em_mac_em_reg_mxopwe_DO_reg[3]/P0001  & n28649 ;
  assign n30540 = ~n28550 & ~n30532 ;
  assign n30541 = ~n30539 & n30540 ;
  assign n30542 = ~n30531 & ~n30541 ;
  assign n30545 = ~n14564 & n28561 ;
  assign n30544 = \core_c_dec_MTAR_E_reg/P0001  & n19559 ;
  assign n30546 = ~n28564 & ~n30544 ;
  assign n30547 = ~n30545 & n30546 ;
  assign n30548 = n28559 & ~n30547 ;
  assign n30550 = ~n12520 & ~n28577 ;
  assign n30549 = ~n7607 & n28577 ;
  assign n30551 = ~n28575 & ~n30549 ;
  assign n30552 = ~n30550 & n30551 ;
  assign n30553 = ~n28576 & ~n30552 ;
  assign n30554 = n28569 & ~n30553 ;
  assign n30620 = ~n7449 & ~n28589 ;
  assign n30618 = ~n7473 & ~n28598 ;
  assign n30619 = ~n7469 & ~n28594 ;
  assign n30621 = ~n30618 & ~n30619 ;
  assign n30622 = ~n30620 & n30621 ;
  assign n30623 = n28607 & n30622 ;
  assign n30624 = n28572 & n30623 ;
  assign n30617 = ~n7607 & ~n28572 ;
  assign n30625 = n28584 & ~n30617 ;
  assign n30626 = ~n30624 & n30625 ;
  assign n30579 = n18766 & ~n18912 ;
  assign n30571 = n18124 & n18147 ;
  assign n30573 = ~n18918 & n20308 ;
  assign n30596 = ~n30571 & ~n30573 ;
  assign n30597 = ~n30579 & n30596 ;
  assign n30607 = n18724 & n30597 ;
  assign n30608 = n18796 & n30607 ;
  assign n30588 = ~n18018 & ~n29242 ;
  assign n30572 = n17952 & n18749 ;
  assign n30578 = ~n18123 & n18148 ;
  assign n30589 = ~n30572 & ~n30578 ;
  assign n30590 = n30588 & n30589 ;
  assign n30582 = n17921 & n18752 ;
  assign n30580 = n18055 & n18754 ;
  assign n30581 = n18055 & n18759 ;
  assign n30585 = ~n30580 & ~n30581 ;
  assign n30586 = ~n30582 & n30585 ;
  assign n30558 = n18056 & n19862 ;
  assign n30577 = \core_c_dec_IRE_reg[11]/NET0131  & ~n7377 ;
  assign n30583 = ~n30558 & ~n30577 ;
  assign n30567 = n18153 & ~n18919 ;
  assign n30569 = n18001 & n18749 ;
  assign n30584 = ~n30567 & ~n30569 ;
  assign n30587 = n30583 & n30584 ;
  assign n30591 = n30586 & n30587 ;
  assign n30600 = n30590 & n30591 ;
  assign n30601 = n29049 & n29239 ;
  assign n30605 = n30600 & n30601 ;
  assign n30562 = n18070 & n18187 ;
  assign n30563 = n18139 & n18758 ;
  assign n30594 = ~n30562 & ~n30563 ;
  assign n30568 = ~n18091 & ~n18743 ;
  assign n30570 = n18046 & n18162 ;
  assign n30595 = ~n30568 & ~n30570 ;
  assign n30598 = n30594 & n30595 ;
  assign n30559 = n18071 & n18183 ;
  assign n30592 = n18038 & ~n30559 ;
  assign n30560 = n18905 & ~n18907 ;
  assign n30561 = n18115 & n18893 ;
  assign n30593 = ~n30560 & ~n30561 ;
  assign n30599 = n30592 & n30593 ;
  assign n30606 = n30598 & n30599 ;
  assign n30609 = n30605 & n30606 ;
  assign n30564 = n18171 & ~n18781 ;
  assign n30565 = ~n17924 & n20996 ;
  assign n30602 = ~n30564 & ~n30565 ;
  assign n30566 = n18745 & ~n19804 ;
  assign n30574 = n17915 & n18751 ;
  assign n30575 = ~n18192 & ~n30574 ;
  assign n30576 = ~n17929 & ~n30575 ;
  assign n30603 = ~n30566 & ~n30576 ;
  assign n30604 = n30602 & n30603 ;
  assign n30610 = n29252 & n30604 ;
  assign n30611 = n30609 & n30610 ;
  assign n30612 = n30608 & n30611 ;
  assign n30613 = n20107 & n30612 ;
  assign n30614 = n28627 & ~n30613 ;
  assign n30543 = n7607 & n28630 ;
  assign n30557 = ~n7422 & ~n28634 ;
  assign n30627 = ~n30543 & ~n30557 ;
  assign n30615 = n12520 & n28619 ;
  assign n30616 = ~n20326 & n28636 ;
  assign n30628 = ~n30615 & ~n30616 ;
  assign n30629 = n30627 & n30628 ;
  assign n30555 = ~n7377 & ~n28556 ;
  assign n30556 = ~n7381 & ~n28624 ;
  assign n30630 = ~n30555 & ~n30556 ;
  assign n30631 = n30629 & n30630 ;
  assign n30632 = ~n30614 & n30631 ;
  assign n30633 = ~n30626 & n30632 ;
  assign n30634 = ~n30554 & n30633 ;
  assign n30635 = ~n30548 & n30634 ;
  assign n30636 = n28550 & ~n30635 ;
  assign n30642 = n19559 & n28660 ;
  assign n30639 = n7457 & ~n28652 ;
  assign n30638 = n7465 & n28652 ;
  assign n30640 = ~n28660 & ~n30638 ;
  assign n30641 = ~n30639 & n30640 ;
  assign n30643 = ~n28649 & ~n30641 ;
  assign n30644 = ~n30642 & n30643 ;
  assign n30637 = ~\core_eu_em_mac_em_reg_mxopwe_DO_reg[0]/P0001  & n28649 ;
  assign n30645 = ~n28550 & ~n30637 ;
  assign n30646 = ~n30644 & n30645 ;
  assign n30647 = ~n30636 & ~n30646 ;
  assign n30649 = n7607 & n28725 ;
  assign n30648 = n12520 & n28729 ;
  assign n30655 = ~\core_c_psq_MSTAT_reg_DO_reg[0]/P0002  & ~\core_eu_em_mac_em_reg_mfrwe_DO_reg[0]/P0001  ;
  assign n30656 = \core_c_psq_MSTAT_reg_DO_reg[0]/P0002  & ~\core_eu_em_mac_em_reg_mfswe_DO_reg[0]/P0001  ;
  assign n30657 = ~n30655 & ~n30656 ;
  assign n30658 = n28741 & n30657 ;
  assign n30650 = n7453 & n28705 ;
  assign n30651 = n7461 & ~n28705 ;
  assign n30652 = ~n30650 & ~n30651 ;
  assign n30653 = n28735 & n30652 ;
  assign n30654 = n28739 & n30641 ;
  assign n30659 = ~n30653 & ~n30654 ;
  assign n30660 = ~n30658 & n30659 ;
  assign n30661 = ~n30648 & n30660 ;
  assign n30662 = ~n30649 & n30661 ;
  assign n30663 = ~n28543 & ~n30662 ;
  assign n30664 = \core_eu_em_mac_em_reg_myopwe_DO_reg[0]/P0001  & ~n28545 ;
  assign n30665 = ~n30663 & ~n30664 ;
  assign n30666 = ~n28719 & ~n30665 ;
  assign n30667 = n28719 & ~n30635 ;
  assign n30668 = ~n30666 & ~n30667 ;
  assign n30670 = n8113 & n28725 ;
  assign n30669 = n12870 & n28729 ;
  assign n30676 = ~\core_c_psq_MSTAT_reg_DO_reg[0]/P0002  & ~\core_eu_em_mac_em_reg_mfrwe_DO_reg[3]/P0001  ;
  assign n30677 = \core_c_psq_MSTAT_reg_DO_reg[0]/P0002  & ~\core_eu_em_mac_em_reg_mfswe_DO_reg[3]/P0001  ;
  assign n30678 = ~n30676 & ~n30677 ;
  assign n30679 = n28741 & n30678 ;
  assign n30671 = n7897 & n28705 ;
  assign n30672 = n7893 & ~n28705 ;
  assign n30673 = ~n30671 & ~n30672 ;
  assign n30674 = n28735 & n30673 ;
  assign n30675 = n28739 & n30536 ;
  assign n30680 = ~n30674 & ~n30675 ;
  assign n30681 = ~n30679 & n30680 ;
  assign n30682 = ~n30669 & n30681 ;
  assign n30683 = ~n30670 & n30682 ;
  assign n30684 = ~n28543 & ~n30683 ;
  assign n30685 = \core_eu_em_mac_em_reg_myopwe_DO_reg[3]/P0001  & ~n28545 ;
  assign n30686 = ~n30684 & ~n30685 ;
  assign n30687 = ~n28719 & ~n30686 ;
  assign n30688 = n28719 & ~n30530 ;
  assign n30689 = ~n30687 & ~n30688 ;
  assign n30690 = n17805 & n28530 ;
  assign n30691 = n19972 & n30690 ;
  assign n30692 = ~n19385 & ~n30691 ;
  assign n30693 = n28532 & ~n30692 ;
  assign n30694 = ~n18268 & n28534 ;
  assign n30695 = \core_eu_em_mac_em_reg_mr2swe_DO_reg[7]/P0001  & ~n30694 ;
  assign n30696 = ~n30693 & ~n30695 ;
  assign n30697 = ~n18262 & ~n30696 ;
  assign n30698 = n18262 & ~n22883 ;
  assign n30699 = ~n30697 & ~n30698 ;
  assign n30700 = \tm_tcr_reg_DO_reg[1]/NET0131  & n20355 ;
  assign n30702 = ~\tm_TCR_TMP_reg[0]/NET0131  & n22411 ;
  assign n30704 = ~\tm_TCR_TMP_reg[1]/NET0131  & n30702 ;
  assign n30703 = \tm_TCR_TMP_reg[1]/NET0131  & ~n30702 ;
  assign n30705 = ~n22400 & ~n30703 ;
  assign n30706 = ~n30704 & n30705 ;
  assign n30701 = ~\tm_tpr_reg_DO_reg[1]/NET0131  & n22400 ;
  assign n30707 = ~n20355 & ~n30701 ;
  assign n30708 = ~n30706 & n30707 ;
  assign n30709 = ~n30700 & ~n30708 ;
  assign n30710 = \tm_tcr_reg_DO_reg[2]/NET0131  & n20355 ;
  assign n30713 = \tm_TCR_TMP_reg[2]/NET0131  & ~n30704 ;
  assign n30712 = ~\tm_TCR_TMP_reg[2]/NET0131  & n30704 ;
  assign n30714 = ~n22400 & ~n30712 ;
  assign n30715 = ~n30713 & n30714 ;
  assign n30711 = ~\tm_tpr_reg_DO_reg[2]/NET0131  & n22400 ;
  assign n30716 = ~n20355 & ~n30711 ;
  assign n30717 = ~n30715 & n30716 ;
  assign n30718 = ~n30710 & ~n30717 ;
  assign n30719 = ~\tm_tpr_reg_DO_reg[6]/NET0131  & n22400 ;
  assign n30720 = \tm_TCR_TMP_reg[6]/NET0131  & ~n27895 ;
  assign n30721 = ~n22400 & ~n27896 ;
  assign n30722 = ~n30720 & n30721 ;
  assign n30723 = ~n30719 & ~n30722 ;
  assign n30724 = ~n20355 & ~n30723 ;
  assign n30725 = ~\tm_tcr_reg_DO_reg[6]/NET0131  & n20355 ;
  assign n30726 = ~n30724 & ~n30725 ;
  assign n30727 = \tm_tcr_reg_DO_reg[5]/NET0131  & n20355 ;
  assign n30729 = \tm_TCR_TMP_reg[4]/NET0131  & n27890 ;
  assign n30733 = ~n27893 & ~n30729 ;
  assign n30734 = n22411 & ~n30733 ;
  assign n30735 = \tm_TCR_TMP_reg[5]/NET0131  & ~n30734 ;
  assign n30730 = \tm_TCR_TMP_reg[5]/NET0131  & n30729 ;
  assign n30731 = ~n27894 & ~n30730 ;
  assign n30732 = n22411 & ~n30731 ;
  assign n30736 = ~n22400 & ~n30732 ;
  assign n30737 = ~n30735 & n30736 ;
  assign n30728 = ~\tm_tpr_reg_DO_reg[5]/NET0131  & n22400 ;
  assign n30738 = ~n20355 & ~n30728 ;
  assign n30739 = ~n30737 & n30738 ;
  assign n30740 = ~n30727 & ~n30739 ;
  assign n30743 = ~n21382 & n22650 ;
  assign n30741 = ~\sport1_cfg_RFSg_d1_reg/NET0131  & \sport1_regs_SCTLreg_DO_reg[11]/NET0131  ;
  assign n30742 = ~\sport1_regs_SCTLreg_DO_reg[12]/NET0131  & n30741 ;
  assign n30745 = \sport1_cfg_RFSg_d3_reg/NET0131  & \sport1_regs_SCTLreg_DO_reg[11]/NET0131  ;
  assign n30744 = \sport1_cfg_RFSg_d2_reg/NET0131  & ~\sport1_regs_SCTLreg_DO_reg[11]/NET0131  ;
  assign n30746 = \sport1_regs_SCTLreg_DO_reg[12]/NET0131  & ~n30744 ;
  assign n30747 = ~n30745 & n30746 ;
  assign n30748 = ~n30742 & ~n30747 ;
  assign n30749 = ~n30743 & n30748 ;
  assign n30750 = \sport1_rxctl_RCS_reg[0]/NET0131  & ~n30749 ;
  assign n30751 = ~\sport1_rxctl_LMcnt_reg[0]/NET0131  & ~\sport1_rxctl_LMcnt_reg[1]/NET0131  ;
  assign n30752 = ~\sport1_rxctl_LMcnt_reg[2]/NET0131  & n30751 ;
  assign n30753 = ~\sport1_rxctl_LMcnt_reg[3]/NET0131  & n30752 ;
  assign n30754 = ~\sport1_rxctl_LMcnt_reg[4]/NET0131  & n30753 ;
  assign n30755 = ~n30750 & ~n30754 ;
  assign n30760 = \sport1_rxctl_RXSHT_reg[0]/P0001  & n30755 ;
  assign n30759 = ~\sport1_regs_SCTLreg_DO_reg[4]/NET0131  & ~\sport1_regs_SCTLreg_DO_reg[5]/NET0131  ;
  assign n30761 = \sport1_rxctl_sht2nd_reg/P0001  & ~n30759 ;
  assign n30762 = n30760 & n30761 ;
  assign n30756 = \sport1_rxctl_RXSHT_reg[15]/P0001  & ~n30755 ;
  assign n30757 = ~\sport1_rxctl_sht2nd_reg/P0001  & n30755 ;
  assign n30758 = \sport1_rxctl_RXSHT_reg[14]/P0001  & n30757 ;
  assign n30763 = ~n30756 & ~n30758 ;
  assign n30764 = ~n30762 & n30763 ;
  assign n30767 = n19933 & ~n21390 ;
  assign n30765 = ~\sport0_cfg_RFSg_d1_reg/NET0131  & \sport0_regs_SCTLreg_DO_reg[11]/NET0131  ;
  assign n30766 = ~\sport0_regs_SCTLreg_DO_reg[12]/NET0131  & n30765 ;
  assign n30769 = \sport0_cfg_RFSg_d3_reg/NET0131  & \sport0_regs_SCTLreg_DO_reg[11]/NET0131  ;
  assign n30768 = \sport0_cfg_RFSg_d2_reg/NET0131  & ~\sport0_regs_SCTLreg_DO_reg[11]/NET0131  ;
  assign n30770 = \sport0_regs_SCTLreg_DO_reg[12]/NET0131  & ~n30768 ;
  assign n30771 = ~n30769 & n30770 ;
  assign n30772 = ~n30766 & ~n30771 ;
  assign n30773 = ~n30767 & n30772 ;
  assign n30774 = \sport0_rxctl_RCS_reg[0]/NET0131  & ~n30773 ;
  assign n30775 = ~\sport0_rxctl_LMcnt_reg[0]/NET0131  & ~\sport0_rxctl_LMcnt_reg[1]/NET0131  ;
  assign n30776 = ~\sport0_rxctl_LMcnt_reg[2]/NET0131  & n30775 ;
  assign n30777 = ~\sport0_rxctl_LMcnt_reg[3]/NET0131  & n30776 ;
  assign n30778 = ~\sport0_rxctl_LMcnt_reg[4]/NET0131  & n30777 ;
  assign n30779 = ~n30774 & ~n30778 ;
  assign n30784 = \sport0_rxctl_RXSHT_reg[0]/P0001  & n30779 ;
  assign n30783 = ~\sport0_regs_SCTLreg_DO_reg[4]/NET0131  & ~\sport0_regs_SCTLreg_DO_reg[5]/NET0131  ;
  assign n30785 = \sport0_rxctl_sht2nd_reg/P0001  & ~n30783 ;
  assign n30786 = n30784 & n30785 ;
  assign n30780 = \sport0_rxctl_RXSHT_reg[10]/P0001  & ~n30779 ;
  assign n30781 = ~\sport0_rxctl_sht2nd_reg/P0001  & n30779 ;
  assign n30782 = \sport0_rxctl_RXSHT_reg[9]/P0001  & n30781 ;
  assign n30787 = ~n30780 & ~n30782 ;
  assign n30788 = ~n30786 & n30787 ;
  assign n30790 = \sport1_rxctl_RXSHT_reg[9]/P0001  & n30757 ;
  assign n30789 = \sport1_rxctl_RXSHT_reg[10]/P0001  & ~n30755 ;
  assign n30791 = ~n30762 & ~n30789 ;
  assign n30792 = ~n30790 & n30791 ;
  assign n30794 = \sport1_rxctl_RXSHT_reg[10]/P0001  & n30757 ;
  assign n30793 = \sport1_rxctl_RXSHT_reg[11]/P0001  & ~n30755 ;
  assign n30795 = ~n30762 & ~n30793 ;
  assign n30796 = ~n30794 & n30795 ;
  assign n30797 = n18262 & n22926 ;
  assign n30799 = n18276 & n30690 ;
  assign n30800 = ~n19385 & ~n30799 ;
  assign n30801 = n28532 & ~n30800 ;
  assign n30798 = \core_eu_em_mac_em_reg_mr2swe_DO_reg[6]/P0001  & ~n28534 ;
  assign n30802 = n28529 & ~n30798 ;
  assign n30803 = ~n30801 & n30802 ;
  assign n30804 = ~n30797 & ~n30803 ;
  assign n30806 = \sport1_rxctl_RXSHT_reg[11]/P0001  & n30757 ;
  assign n30805 = \sport1_rxctl_RXSHT_reg[12]/P0001  & ~n30755 ;
  assign n30807 = ~n30762 & ~n30805 ;
  assign n30808 = ~n30806 & n30807 ;
  assign n30810 = \sport1_rxctl_RXSHT_reg[12]/P0001  & n30757 ;
  assign n30809 = \sport1_rxctl_RXSHT_reg[13]/P0001  & ~n30755 ;
  assign n30811 = ~n30762 & ~n30809 ;
  assign n30812 = ~n30810 & n30811 ;
  assign n30814 = \sport1_rxctl_RXSHT_reg[13]/P0001  & n30757 ;
  assign n30813 = \sport1_rxctl_RXSHT_reg[14]/P0001  & ~n30755 ;
  assign n30815 = ~n30762 & ~n30813 ;
  assign n30816 = ~n30814 & n30815 ;
  assign n30818 = \sport1_rxctl_RXSHT_reg[1]/P0001  & n30757 ;
  assign n30817 = \sport1_rxctl_RXSHT_reg[2]/P0001  & ~n30755 ;
  assign n30819 = ~n30762 & ~n30817 ;
  assign n30820 = ~n30818 & n30819 ;
  assign n30822 = \sport1_rxctl_RXSHT_reg[2]/P0001  & n30757 ;
  assign n30821 = \sport1_rxctl_RXSHT_reg[3]/P0001  & ~n30755 ;
  assign n30823 = ~n30762 & ~n30821 ;
  assign n30824 = ~n30822 & n30823 ;
  assign n30826 = \sport1_rxctl_RXSHT_reg[3]/P0001  & n30757 ;
  assign n30825 = \sport1_rxctl_RXSHT_reg[4]/P0001  & ~n30755 ;
  assign n30827 = ~n30762 & ~n30825 ;
  assign n30828 = ~n30826 & n30827 ;
  assign n30830 = \sport1_rxctl_RXSHT_reg[4]/P0001  & n30757 ;
  assign n30829 = \sport1_rxctl_RXSHT_reg[5]/P0001  & ~n30755 ;
  assign n30831 = ~n30762 & ~n30829 ;
  assign n30832 = ~n30830 & n30831 ;
  assign n30834 = \sport1_rxctl_RXSHT_reg[5]/P0001  & n30757 ;
  assign n30833 = \sport1_rxctl_RXSHT_reg[6]/P0001  & ~n30755 ;
  assign n30835 = ~n30762 & ~n30833 ;
  assign n30836 = ~n30834 & n30835 ;
  assign n30838 = \sport1_rxctl_RXSHT_reg[7]/P0001  & n30757 ;
  assign n30837 = \sport1_rxctl_RXSHT_reg[8]/P0001  & ~n30755 ;
  assign n30839 = ~n30762 & ~n30837 ;
  assign n30840 = ~n30838 & n30839 ;
  assign n30842 = \sport1_rxctl_RXSHT_reg[8]/P0001  & n30757 ;
  assign n30841 = \sport1_rxctl_RXSHT_reg[9]/P0001  & ~n30755 ;
  assign n30843 = ~n30762 & ~n30841 ;
  assign n30844 = ~n30842 & n30843 ;
  assign n30846 = \sport0_rxctl_RXSHT_reg[10]/P0001  & n30781 ;
  assign n30845 = \sport0_rxctl_RXSHT_reg[11]/P0001  & ~n30779 ;
  assign n30847 = ~n30786 & ~n30845 ;
  assign n30848 = ~n30846 & n30847 ;
  assign n30850 = \sport0_rxctl_RXSHT_reg[13]/P0001  & n30781 ;
  assign n30849 = \sport0_rxctl_RXSHT_reg[14]/P0001  & ~n30779 ;
  assign n30851 = ~n30786 & ~n30849 ;
  assign n30852 = ~n30850 & n30851 ;
  assign n30854 = \sport0_rxctl_RXSHT_reg[14]/P0001  & n30781 ;
  assign n30853 = \sport0_rxctl_RXSHT_reg[15]/P0001  & ~n30779 ;
  assign n30855 = ~n30786 & ~n30853 ;
  assign n30856 = ~n30854 & n30855 ;
  assign n30858 = \sport0_rxctl_RXSHT_reg[1]/P0001  & n30781 ;
  assign n30857 = \sport0_rxctl_RXSHT_reg[2]/P0001  & ~n30779 ;
  assign n30859 = ~n30786 & ~n30857 ;
  assign n30860 = ~n30858 & n30859 ;
  assign n30862 = \sport0_rxctl_RXSHT_reg[2]/P0001  & n30781 ;
  assign n30861 = \sport0_rxctl_RXSHT_reg[3]/P0001  & ~n30779 ;
  assign n30863 = ~n30786 & ~n30861 ;
  assign n30864 = ~n30862 & n30863 ;
  assign n30866 = \sport0_rxctl_RXSHT_reg[3]/P0001  & n30781 ;
  assign n30865 = \sport0_rxctl_RXSHT_reg[4]/P0001  & ~n30779 ;
  assign n30867 = ~n30786 & ~n30865 ;
  assign n30868 = ~n30866 & n30867 ;
  assign n30870 = \sport0_rxctl_RXSHT_reg[4]/P0001  & n30781 ;
  assign n30869 = \sport0_rxctl_RXSHT_reg[5]/P0001  & ~n30779 ;
  assign n30871 = ~n30786 & ~n30869 ;
  assign n30872 = ~n30870 & n30871 ;
  assign n30874 = \sport0_rxctl_RXSHT_reg[5]/P0001  & n30781 ;
  assign n30873 = \sport0_rxctl_RXSHT_reg[6]/P0001  & ~n30779 ;
  assign n30875 = ~n30786 & ~n30873 ;
  assign n30876 = ~n30874 & n30875 ;
  assign n30878 = \sport0_rxctl_RXSHT_reg[6]/P0001  & n30781 ;
  assign n30877 = \sport0_rxctl_RXSHT_reg[7]/P0001  & ~n30779 ;
  assign n30879 = ~n30786 & ~n30877 ;
  assign n30880 = ~n30878 & n30879 ;
  assign n30882 = \sport0_rxctl_RXSHT_reg[7]/P0001  & n30781 ;
  assign n30881 = \sport0_rxctl_RXSHT_reg[8]/P0001  & ~n30779 ;
  assign n30883 = ~n30786 & ~n30881 ;
  assign n30884 = ~n30882 & n30883 ;
  assign n30886 = \sport0_rxctl_RXSHT_reg[8]/P0001  & n30781 ;
  assign n30885 = \sport0_rxctl_RXSHT_reg[9]/P0001  & ~n30779 ;
  assign n30887 = ~n30786 & ~n30885 ;
  assign n30888 = ~n30886 & n30887 ;
  assign n30890 = \sport1_rxctl_RXSHT_reg[6]/P0001  & n30757 ;
  assign n30889 = \sport1_rxctl_RXSHT_reg[7]/P0001  & ~n30755 ;
  assign n30891 = ~n30762 & ~n30889 ;
  assign n30892 = ~n30890 & n30891 ;
  assign n30894 = \sport0_rxctl_RXSHT_reg[12]/P0001  & n30781 ;
  assign n30893 = \sport0_rxctl_RXSHT_reg[13]/P0001  & ~n30779 ;
  assign n30895 = ~n30786 & ~n30893 ;
  assign n30896 = ~n30894 & n30895 ;
  assign n30898 = \sport0_rxctl_RXSHT_reg[11]/P0001  & n30781 ;
  assign n30897 = \sport0_rxctl_RXSHT_reg[12]/P0001  & ~n30779 ;
  assign n30899 = ~n30786 & ~n30897 ;
  assign n30900 = ~n30898 & n30899 ;
  assign n30902 = ~n19205 & n19243 ;
  assign n30901 = ~\core_eu_ec_cun_AN_reg/P0001  & n19205 ;
  assign n30903 = n4150 & ~n30901 ;
  assign n30904 = ~n30902 & n30903 ;
  assign n30905 = n17799 & n17805 ;
  assign n30906 = n19972 & n30905 ;
  assign n30907 = ~n17823 & ~n30906 ;
  assign n30908 = n17808 & ~n30907 ;
  assign n30909 = n17811 & ~n17827 ;
  assign n30910 = \core_eu_em_mac_em_reg_mr2rwe_DO_reg[7]/P0001  & ~n30909 ;
  assign n30911 = ~n30908 & ~n30910 ;
  assign n30912 = ~n14752 & ~n30911 ;
  assign n30913 = n14752 & ~n22883 ;
  assign n30914 = ~n30912 & ~n30913 ;
  assign n30915 = \tm_tcr_reg_DO_reg[13]/NET0131  & n20355 ;
  assign n30917 = \tm_TCR_TMP_reg[13]/NET0131  & ~n25840 ;
  assign n30918 = ~n22400 & ~n25841 ;
  assign n30919 = ~n30917 & n30918 ;
  assign n30916 = ~\tm_tpr_reg_DO_reg[13]/NET0131  & n22400 ;
  assign n30920 = ~n20355 & ~n30916 ;
  assign n30921 = ~n30919 & n30920 ;
  assign n30922 = ~n30915 & ~n30921 ;
  assign n30923 = n14752 & n22926 ;
  assign n30924 = ~\core_eu_em_mac_em_reg_mr2rwe_DO_reg[6]/P0001  & ~n17799 ;
  assign n30925 = ~n17809 & n18276 ;
  assign n30926 = n17811 & ~n30925 ;
  assign n30927 = ~n30924 & ~n30926 ;
  assign n30928 = ~n17823 & ~n30927 ;
  assign n30929 = ~\core_eu_em_mac_em_reg_mr2rwe_DO_reg[6]/P0001  & ~n17808 ;
  assign n30930 = ~n30928 & ~n30929 ;
  assign n30931 = n17829 & ~n30930 ;
  assign n30932 = ~n30923 & ~n30931 ;
  assign n30933 = \core_c_dec_pMFMAC_Ei_reg/NET0131  & n4117 ;
  assign n30934 = ~n4117 & ~n19701 ;
  assign n30953 = ~n6116 & n6956 ;
  assign n30935 = n6028 & n19696 ;
  assign n30954 = ~n26373 & n30935 ;
  assign n30955 = ~n30953 & ~n30954 ;
  assign n30937 = n6028 & n21248 ;
  assign n30940 = ~n18839 & ~n25469 ;
  assign n30941 = ~n24646 & n30940 ;
  assign n30942 = ~n30937 & n30941 ;
  assign n30936 = ~n24644 & ~n30935 ;
  assign n30938 = ~n6024 & n6119 ;
  assign n30939 = \core_c_dec_IR_reg[15]/NET0131  & n30938 ;
  assign n30943 = n30936 & ~n30939 ;
  assign n30944 = n30942 & n30943 ;
  assign n30945 = \core_c_dec_IR_reg[17]/NET0131  & n6028 ;
  assign n30946 = ~n6956 & ~n18839 ;
  assign n30947 = ~n25081 & n30946 ;
  assign n30948 = ~n30945 & n30947 ;
  assign n30949 = \core_c_dec_IR_reg[0]/NET0131  & ~n30948 ;
  assign n30950 = \core_c_dec_IR_reg[4]/NET0131  & n30948 ;
  assign n30951 = ~n30949 & ~n30950 ;
  assign n30973 = ~n30944 & n30951 ;
  assign n30974 = n30955 & n30973 ;
  assign n30964 = \core_c_dec_IR_reg[3]/NET0131  & ~n30948 ;
  assign n30965 = \core_c_dec_IR_reg[7]/NET0131  & n30948 ;
  assign n30966 = ~n30964 & ~n30965 ;
  assign n30956 = \core_c_dec_IR_reg[2]/NET0131  & ~n30948 ;
  assign n30957 = \core_c_dec_IR_reg[6]/NET0131  & n30948 ;
  assign n30958 = ~n30956 & ~n30957 ;
  assign n30959 = \core_c_dec_IR_reg[1]/NET0131  & ~n30948 ;
  assign n30960 = \core_c_dec_IR_reg[5]/NET0131  & n30948 ;
  assign n30961 = ~n30959 & ~n30960 ;
  assign n30977 = ~n30958 & n30961 ;
  assign n30978 = ~n30966 & n30977 ;
  assign n30982 = n30974 & n30978 ;
  assign n30952 = ~n30944 & ~n30951 ;
  assign n30970 = n30952 & n30955 ;
  assign n30979 = n30970 & n30978 ;
  assign n30962 = n30958 & ~n30961 ;
  assign n30963 = n30955 & n30962 ;
  assign n30980 = ~n30944 & n30966 ;
  assign n30981 = n30963 & n30980 ;
  assign n30983 = ~n30979 & ~n30981 ;
  assign n30984 = ~n30982 & n30983 ;
  assign n30969 = ~n30958 & ~n30961 ;
  assign n30975 = n30966 & n30974 ;
  assign n30976 = n30969 & n30975 ;
  assign n30967 = n30963 & ~n30966 ;
  assign n30968 = n30952 & n30967 ;
  assign n30971 = n30966 & n30970 ;
  assign n30972 = n30969 & n30971 ;
  assign n30985 = ~n30968 & ~n30972 ;
  assign n30986 = ~n30976 & n30985 ;
  assign n30987 = n30984 & n30986 ;
  assign n30988 = n30934 & ~n30987 ;
  assign n30989 = ~n30933 & ~n30988 ;
  assign n30990 = \core_c_dec_MFMAC_Ei_reg/NET0131  & n4117 ;
  assign n30991 = n25047 & ~n30987 ;
  assign n30992 = ~n30990 & ~n30991 ;
  assign n30993 = \sport1_regs_FSDIVreg_DO_reg[11]/NET0131  & n28786 ;
  assign n30994 = ~\sport1_cfg_FSi_cnt_reg[11]/NET0131  & ~n28866 ;
  assign n30995 = n28855 & ~n28867 ;
  assign n30996 = ~n30994 & n30995 ;
  assign n30997 = ~n30993 & ~n30996 ;
  assign n30998 = \sport0_regs_FSDIVreg_DO_reg[11]/NET0131  & n28876 ;
  assign n30999 = ~\sport0_cfg_FSi_cnt_reg[11]/NET0131  & ~n28956 ;
  assign n31000 = n28945 & ~n28957 ;
  assign n31001 = ~n30999 & n31000 ;
  assign n31002 = ~n30998 & ~n31001 ;
  assign n31003 = \tm_tcr_reg_DO_reg[0]/NET0131  & n20355 ;
  assign n31005 = \tm_TCR_TMP_reg[0]/NET0131  & ~n22411 ;
  assign n31006 = ~n22400 & ~n30702 ;
  assign n31007 = ~n31005 & n31006 ;
  assign n31004 = ~\tm_tpr_reg_DO_reg[0]/NET0131  & n22400 ;
  assign n31008 = ~n20355 & ~n31004 ;
  assign n31009 = ~n31007 & n31008 ;
  assign n31010 = ~n31003 & ~n31009 ;
  assign n31011 = \tm_tcr_reg_DO_reg[3]/NET0131  & n20355 ;
  assign n31014 = \tm_TCR_TMP_reg[3]/NET0131  & ~n30712 ;
  assign n31013 = n20359 & n30702 ;
  assign n31015 = ~n22400 & ~n31013 ;
  assign n31016 = ~n31014 & n31015 ;
  assign n31012 = ~\tm_tpr_reg_DO_reg[3]/NET0131  & n22400 ;
  assign n31017 = ~n20355 & ~n31012 ;
  assign n31018 = ~n31016 & n31017 ;
  assign n31019 = ~n31011 & ~n31018 ;
  assign n31020 = \tm_tcr_reg_DO_reg[4]/NET0131  & n20355 ;
  assign n31022 = \tm_TCR_TMP_reg[4]/NET0131  & ~n22411 ;
  assign n31023 = ~n22400 & ~n30734 ;
  assign n31024 = ~n31022 & n31023 ;
  assign n31021 = ~\tm_tpr_reg_DO_reg[4]/NET0131  & n22400 ;
  assign n31025 = ~n20355 & ~n31021 ;
  assign n31026 = ~n31024 & n31025 ;
  assign n31027 = ~n31020 & ~n31026 ;
  assign n31030 = n20957 & n20976 ;
  assign n31039 = ~n20882 & n20966 ;
  assign n31040 = ~n20974 & n31039 ;
  assign n31031 = ~n20966 & n20974 ;
  assign n31032 = ~\sport0_rxctl_RX_reg[4]/P0001  & ~n20914 ;
  assign n31033 = n20878 & ~n31032 ;
  assign n31034 = \sport0_rxctl_RX_reg[6]/P0001  & ~n31033 ;
  assign n31035 = ~\sport0_rxctl_RX_reg[6]/P0001  & n20884 ;
  assign n31036 = ~n20891 & ~n31035 ;
  assign n31037 = ~n31034 & n31036 ;
  assign n31038 = n20882 & n31037 ;
  assign n31041 = ~n31031 & ~n31038 ;
  assign n31042 = ~n31040 & n31041 ;
  assign n31043 = n31030 & n31042 ;
  assign n31045 = ~\sport0_rxctl_RX_reg[4]/P0001  & n20878 ;
  assign n31046 = ~\sport0_rxctl_RX_reg[6]/P0001  & n31045 ;
  assign n31049 = ~n31043 & ~n31046 ;
  assign n31050 = ~\sport0_regs_SCTLreg_DO_reg[4]/NET0131  & ~n31049 ;
  assign n31051 = ~\sport0_rxctl_RX_reg[7]/P0001  & ~n31050 ;
  assign n31044 = ~\sport0_rxctl_RX_reg[7]/P0001  & ~n31043 ;
  assign n31047 = ~\sport0_regs_SCTLreg_DO_reg[4]/NET0131  & n31046 ;
  assign n31048 = ~n31044 & n31047 ;
  assign n31052 = \sport0_regs_SCTLreg_DO_reg[5]/NET0131  & ~n31048 ;
  assign n31053 = ~n31051 & n31052 ;
  assign n31029 = ~\sport0_regs_SCTLreg_DO_reg[5]/NET0131  & ~\sport0_rxctl_RX_reg[12]/P0001  ;
  assign n31054 = \sport0_rxctl_ldRX_cmp_reg/P0001  & ~n31029 ;
  assign n31055 = ~n31053 & n31054 ;
  assign n31056 = ~\sport0_rxctl_ldRX_cmp_reg/P0001  & n20869 ;
  assign n31057 = n9178 & n31056 ;
  assign n31058 = ~n31055 & ~n31057 ;
  assign n31059 = ~n20868 & ~n31058 ;
  assign n31028 = \sport0_rxctl_RX_reg[12]/P0001  & n20871 ;
  assign n31060 = \sport0_rxctl_RXSHT_reg[12]/P0001  & n20868 ;
  assign n31061 = ~n31028 & ~n31060 ;
  assign n31062 = ~n31059 & n31061 ;
  assign n31063 = ~\core_c_dec_MTAR_E_reg/P0001  & ~\core_c_dec_updAR_E_reg/P0001  ;
  assign n31064 = n14666 & ~n31063 ;
  assign n31065 = ~n29291 & n31064 ;
  assign n31066 = \core_eu_ea_alu_ea_reg_arswe_DO_reg[15]/P0001  & ~n31064 ;
  assign n31067 = ~n31065 & ~n31066 ;
  assign n31069 = ~\core_c_dec_IR_reg[20]/NET0131  & ~\core_c_dec_IR_reg[21]/NET0131  ;
  assign n31070 = \core_c_dec_IR_reg[22]/NET0131  & ~\core_c_dec_IR_reg[23]/NET0131  ;
  assign n31071 = ~n31069 & n31070 ;
  assign n31072 = ~n25244 & ~n31071 ;
  assign n31073 = ~n25081 & n31072 ;
  assign n31074 = \core_c_dec_IR_reg[1]/NET0131  & ~n31073 ;
  assign n31075 = \core_c_dec_IR_reg[5]/NET0131  & n31073 ;
  assign n31076 = ~n31074 & ~n31075 ;
  assign n31077 = \core_c_dec_IR_reg[2]/NET0131  & ~n31073 ;
  assign n31078 = \core_c_dec_IR_reg[6]/NET0131  & n31073 ;
  assign n31079 = ~n31077 & ~n31078 ;
  assign n31080 = ~n31076 & ~n31079 ;
  assign n31081 = ~n25081 & ~n30938 ;
  assign n31082 = ~\core_c_dec_IR_reg[15]/NET0131  & ~n31081 ;
  assign n31084 = ~n18839 & ~n24441 ;
  assign n31085 = ~n13578 & n31084 ;
  assign n31086 = ~n11744 & n31085 ;
  assign n31083 = ~n11745 & ~n25244 ;
  assign n31087 = ~n30945 & n31083 ;
  assign n31088 = n31086 & n31087 ;
  assign n31089 = ~n31082 & n31088 ;
  assign n31091 = \core_c_dec_IR_reg[11]/NET0131  & n30935 ;
  assign n31090 = \core_c_dec_IR_reg[10]/NET0131  & n30935 ;
  assign n31092 = ~n25244 & ~n30953 ;
  assign n31093 = ~n31090 & n31092 ;
  assign n31094 = ~n31091 & n31093 ;
  assign n31095 = ~n31089 & n31094 ;
  assign n31096 = \core_c_dec_IR_reg[0]/NET0131  & ~n31073 ;
  assign n31097 = \core_c_dec_IR_reg[4]/NET0131  & n31073 ;
  assign n31098 = ~n31096 & ~n31097 ;
  assign n31099 = n31095 & ~n31098 ;
  assign n31100 = \core_c_dec_IR_reg[3]/NET0131  & ~n31073 ;
  assign n31101 = \core_c_dec_IR_reg[7]/NET0131  & n31073 ;
  assign n31102 = ~n31100 & ~n31101 ;
  assign n31103 = n31099 & n31102 ;
  assign n31104 = n31080 & n31103 ;
  assign n31105 = \core_c_dec_IR_reg[20]/NET0131  & n6023 ;
  assign n31106 = ~n4117 & ~n31105 ;
  assign n31107 = ~n31104 & n31106 ;
  assign n31068 = ~\core_c_dec_MTMY1_E_reg/P0001  & n4117 ;
  assign n31108 = n4116 & ~n31068 ;
  assign n31109 = ~n31107 & n31108 ;
  assign n31111 = n31095 & n31098 ;
  assign n31112 = n31102 & n31111 ;
  assign n31113 = n31080 & n31112 ;
  assign n31114 = ~\core_c_dec_IR_reg[20]/NET0131  & n6023 ;
  assign n31115 = ~n4117 & ~n31114 ;
  assign n31116 = ~n31113 & n31115 ;
  assign n31110 = ~\core_c_dec_MTMY0_E_reg/P0001  & n4117 ;
  assign n31117 = n4116 & ~n31110 ;
  assign n31118 = ~n31116 & n31117 ;
  assign n31119 = \core_c_dec_MTAY1_E_reg/P0001  & n4117 ;
  assign n31120 = ~n4117 & n31099 ;
  assign n31121 = n31076 & n31102 ;
  assign n31122 = ~n31079 & n31121 ;
  assign n31123 = n31120 & n31122 ;
  assign n31124 = ~n31119 & ~n31123 ;
  assign n31125 = n4116 & ~n31124 ;
  assign n31126 = \core_c_dec_MTAY0_E_reg/P0001  & n4117 ;
  assign n31127 = ~n4117 & n31111 ;
  assign n31128 = n31122 & n31127 ;
  assign n31129 = ~n31126 & ~n31128 ;
  assign n31130 = n4116 & ~n31129 ;
  assign n31131 = ~\sport0_cfg_SCLKi_cnt_reg[11]/NET0131  & ~n19548 ;
  assign n31132 = n19197 & ~n19549 ;
  assign n31133 = ~n31131 & n31132 ;
  assign n31134 = n13804 & ~n31063 ;
  assign n31135 = ~n29291 & n31134 ;
  assign n31136 = \core_eu_ea_alu_ea_reg_arrwe_DO_reg[15]/P0001  & ~n31134 ;
  assign n31137 = ~n31135 & ~n31136 ;
  assign n31140 = n18271 & ~n23757 ;
  assign n31139 = ~\core_eu_em_mac_em_reg_mr0swe_DO_reg[11]/P0001  & ~n18271 ;
  assign n31141 = n18273 & ~n31139 ;
  assign n31142 = ~n31140 & n31141 ;
  assign n31138 = \core_eu_em_mac_em_reg_mr0swe_DO_reg[11]/P0001  & ~n18266 ;
  assign n31143 = ~n18270 & ~n31138 ;
  assign n31144 = ~n31142 & n31143 ;
  assign n31145 = ~n18262 & ~n31144 ;
  assign n31146 = n18262 & ~n19618 ;
  assign n31147 = ~n31145 & ~n31146 ;
  assign n31148 = n14752 & n19618 ;
  assign n31149 = n18328 & n23757 ;
  assign n31150 = \core_eu_em_mac_em_reg_mr0rwe_DO_reg[11]/P0001  & ~n18330 ;
  assign n31151 = n18334 & ~n31150 ;
  assign n31152 = ~n31149 & n31151 ;
  assign n31153 = ~n31148 & ~n31152 ;
  assign n31154 = ~\sice_RCS_reg[1]/NET0131  & ~\sice_RST_req_reg/NET0131  ;
  assign n31155 = ~\sice_RCS_reg[0]/NET0131  & ~n31154 ;
  assign n31156 = IACKn_pad & \sice_RCS_reg[0]/NET0131  ;
  assign n31157 = ~\sice_RCS_reg[1]/NET0131  & n31156 ;
  assign n31158 = ~n31155 & ~n31157 ;
  assign n31160 = n19499 & ~n23757 ;
  assign n31159 = ~\core_eu_em_mac_em_reg_mr1swe_DO_reg[11]/P0001  & ~n19499 ;
  assign n31161 = n19501 & ~n31159 ;
  assign n31162 = ~n31160 & n31161 ;
  assign n31163 = \core_eu_em_mac_em_reg_mr1swe_DO_reg[11]/P0001  & ~n19383 ;
  assign n31164 = ~n19508 & ~n31163 ;
  assign n31165 = ~n31162 & n31164 ;
  assign n31166 = ~n18262 & ~n31165 ;
  assign n31167 = n18262 & ~n19436 ;
  assign n31168 = ~n31166 & ~n31167 ;
  assign n31169 = \core_eu_ea_alu_ea_reg_ay0swe_DO_reg[0]/P0001  & ~n21990 ;
  assign n31170 = ~n13806 & ~n24517 ;
  assign n31171 = \core_c_dec_DIVS_E_reg/P0001  & ~n14486 ;
  assign n31172 = ~\core_c_dec_DIVS_E_reg/P0001  & n19222 ;
  assign n31173 = ~n31171 & ~n31172 ;
  assign n31174 = n13837 & ~n31173 ;
  assign n31175 = ~n13837 & n31173 ;
  assign n31176 = ~n31174 & ~n31175 ;
  assign n31178 = ~\core_c_dec_DIVS_E_reg/P0001  & ~n31176 ;
  assign n31177 = \core_c_dec_DIVS_E_reg/P0001  & n31176 ;
  assign n31179 = n13806 & ~n31177 ;
  assign n31180 = ~n31178 & n31179 ;
  assign n31181 = ~n31170 & ~n31180 ;
  assign n31182 = n21990 & n31181 ;
  assign n31183 = ~n31169 & ~n31182 ;
  assign n31184 = \core_eu_ea_alu_ea_reg_ay0rwe_DO_reg[0]/P0001  & ~n22158 ;
  assign n31185 = n22158 & n31181 ;
  assign n31186 = ~n31184 & ~n31185 ;
  assign n31187 = ~\sport1_cfg_SCLKi_cnt_reg[11]/NET0131  & ~n20249 ;
  assign n31188 = n19130 & ~n20250 ;
  assign n31189 = ~n31187 & n31188 ;
  assign n31206 = n14564 & n19206 ;
  assign n31207 = ~n14573 & n31206 ;
  assign n31208 = n14586 & n31207 ;
  assign n31209 = n14610 & n31208 ;
  assign n31210 = n14600 & n31209 ;
  assign n31211 = n14634 & n31210 ;
  assign n31212 = n14623 & n31211 ;
  assign n31213 = n23253 & n31212 ;
  assign n31214 = n14658 & n31213 ;
  assign n31215 = n14649 & n31214 ;
  assign n31216 = n20053 & n31215 ;
  assign n31217 = n14424 & n31216 ;
  assign n31218 = n14413 & n31217 ;
  assign n31219 = n14551 & n31218 ;
  assign n31220 = ~n14540 & n31219 ;
  assign n31221 = n19222 & n31220 ;
  assign n31197 = \core_c_psq_ststk_sts7x23_STcell_reg[5][0]/P0001  & n14699 ;
  assign n31195 = \core_c_psq_ststk_sts7x23_STcell_reg[3][0]/P0001  & n14704 ;
  assign n31196 = \core_c_psq_ststk_sts7x23_STcell_reg[6][0]/P0001  & n14711 ;
  assign n31200 = ~n31195 & ~n31196 ;
  assign n31201 = ~n31197 & n31200 ;
  assign n31191 = \core_c_psq_ststk_sts7x23_STcell_reg[2][0]/P0001  & n14713 ;
  assign n31192 = \core_c_psq_ststk_sts7x23_STcell_reg[0][0]/P0001  & n14702 ;
  assign n31198 = ~n31191 & ~n31192 ;
  assign n31193 = \core_c_psq_ststk_sts7x23_STcell_reg[1][0]/P0001  & n14708 ;
  assign n31194 = \core_c_psq_ststk_sts7x23_STcell_reg[4][0]/P0001  & n14706 ;
  assign n31199 = ~n31193 & ~n31194 ;
  assign n31202 = n31198 & n31199 ;
  assign n31203 = n31201 & n31202 ;
  assign n31204 = n14697 & ~n31203 ;
  assign n31205 = \core_c_dec_MTASTAT_E_reg/P0001  & n7607 ;
  assign n31222 = ~n31204 & ~n31205 ;
  assign n31223 = ~n19205 & n31222 ;
  assign n31224 = ~n31221 & n31223 ;
  assign n31190 = ~\core_eu_ec_cun_AZ_reg/P0001  & n19205 ;
  assign n31225 = n4150 & ~n31190 ;
  assign n31226 = ~n31224 & n31225 ;
  assign n31227 = n14752 & n19436 ;
  assign n31228 = n19776 & n23757 ;
  assign n31229 = \core_eu_em_mac_em_reg_mr1rwe_DO_reg[11]/P0001  & ~n17809 ;
  assign n31230 = n19780 & ~n31229 ;
  assign n31231 = ~n31228 & n31230 ;
  assign n31232 = ~n31227 & ~n31231 ;
  assign n31251 = n13806 & n31176 ;
  assign n31233 = ~n5950 & n13806 ;
  assign n31234 = n19202 & ~n31233 ;
  assign n31236 = \core_c_dec_MTASTAT_E_reg/P0001  & n10911 ;
  assign n31243 = \core_c_psq_ststk_sts7x23_STcell_reg[6][5]/P0001  & n14711 ;
  assign n31241 = \core_c_psq_ststk_sts7x23_STcell_reg[3][5]/P0001  & n14704 ;
  assign n31242 = \core_c_psq_ststk_sts7x23_STcell_reg[5][5]/P0001  & n14699 ;
  assign n31246 = ~n31241 & ~n31242 ;
  assign n31247 = ~n31243 & n31246 ;
  assign n31237 = \core_c_psq_ststk_sts7x23_STcell_reg[2][5]/P0001  & n14713 ;
  assign n31238 = \core_c_psq_ststk_sts7x23_STcell_reg[0][5]/P0001  & n14702 ;
  assign n31244 = ~n31237 & ~n31238 ;
  assign n31239 = \core_c_psq_ststk_sts7x23_STcell_reg[4][5]/P0001  & n14706 ;
  assign n31240 = \core_c_psq_ststk_sts7x23_STcell_reg[1][5]/P0001  & n14708 ;
  assign n31245 = ~n31239 & ~n31240 ;
  assign n31248 = n31244 & n31245 ;
  assign n31249 = n31247 & n31248 ;
  assign n31250 = n14697 & ~n31249 ;
  assign n31252 = ~n31236 & ~n31250 ;
  assign n31253 = ~n31234 & n31252 ;
  assign n31254 = ~n31251 & n31253 ;
  assign n31235 = ~\core_eu_ec_cun_AQ_reg/P0001  & n31234 ;
  assign n31255 = n4150 & ~n31235 ;
  assign n31256 = ~n31254 & n31255 ;
  assign n31257 = \core_c_dec_pMFALU_Ei_reg/NET0131  & n4117 ;
  assign n31260 = n30967 & n30973 ;
  assign n31258 = n30955 & n30961 ;
  assign n31259 = n30980 & n31258 ;
  assign n31261 = \core_c_dec_IR_reg[8]/NET0131  & n30935 ;
  assign n31262 = \core_c_dec_IR_reg[18]/NET0131  & ~n30935 ;
  assign n31263 = ~n31261 & ~n31262 ;
  assign n31264 = ~n30936 & ~n31263 ;
  assign n31265 = ~\core_c_dec_IR_reg[1]/NET0131  & ~\core_c_dec_IR_reg[2]/NET0131  ;
  assign n31266 = n31264 & n31265 ;
  assign n31267 = \core_c_dec_IR_reg[9]/NET0131  & n30935 ;
  assign n31268 = \core_c_dec_IR_reg[19]/NET0131  & ~n30935 ;
  assign n31269 = ~n31267 & ~n31268 ;
  assign n31270 = ~\core_c_dec_IR_reg[0]/NET0131  & ~n31269 ;
  assign n31271 = ~\core_c_dec_IR_reg[3]/NET0131  & n31270 ;
  assign n31272 = n31266 & n31271 ;
  assign n31273 = ~n31259 & ~n31272 ;
  assign n31274 = ~n31260 & n31273 ;
  assign n31275 = n30934 & ~n31274 ;
  assign n31276 = ~n31257 & ~n31275 ;
  assign n31277 = \core_c_dec_MFALU_Ei_reg/NET0131  & n4117 ;
  assign n31278 = n25047 & ~n31274 ;
  assign n31279 = ~n31277 & ~n31278 ;
  assign n31280 = \sport1_txctl_TXSHT_reg[6]/P0001  & ~n22677 ;
  assign n31281 = \sport1_txctl_TX_reg[7]/P0001  & n22677 ;
  assign n31282 = ~n31280 & ~n31281 ;
  assign n31283 = \sport1_regs_FSDIVreg_DO_reg[10]/NET0131  & n28786 ;
  assign n31284 = ~\sport1_cfg_FSi_cnt_reg[10]/NET0131  & ~n28865 ;
  assign n31285 = n28855 & ~n28866 ;
  assign n31286 = ~n31284 & n31285 ;
  assign n31287 = ~n31283 & ~n31286 ;
  assign n31288 = \sport1_regs_FSDIVreg_DO_reg[12]/NET0131  & n28786 ;
  assign n31289 = ~\sport1_cfg_FSi_cnt_reg[12]/NET0131  & ~n28867 ;
  assign n31290 = n28855 & ~n28868 ;
  assign n31291 = ~n31289 & n31290 ;
  assign n31292 = ~n31288 & ~n31291 ;
  assign n31293 = \sport0_regs_FSDIVreg_DO_reg[10]/NET0131  & n28876 ;
  assign n31294 = ~\sport0_cfg_FSi_cnt_reg[10]/NET0131  & ~n28955 ;
  assign n31295 = n28945 & ~n28956 ;
  assign n31296 = ~n31294 & n31295 ;
  assign n31297 = ~n31293 & ~n31296 ;
  assign n31298 = \sport0_txctl_TXSHT_reg[6]/P0001  & ~n19960 ;
  assign n31299 = \sport0_txctl_TX_reg[7]/P0001  & n19960 ;
  assign n31300 = ~n31298 & ~n31299 ;
  assign n31301 = \sport0_regs_FSDIVreg_DO_reg[12]/NET0131  & n28876 ;
  assign n31302 = ~\sport0_cfg_FSi_cnt_reg[12]/NET0131  & ~n28957 ;
  assign n31303 = n28945 & ~n28958 ;
  assign n31304 = ~n31302 & n31303 ;
  assign n31305 = ~n31301 & ~n31304 ;
  assign n31306 = \core_dag_ilm2reg_M_E_reg[1]/NET0131  & ~n5692 ;
  assign n31307 = n4055 & ~n25690 ;
  assign n31309 = \sport1_regs_AUTOreg_DO_reg[3]/NET0131  & n5966 ;
  assign n31310 = \sport1_regs_AUTOreg_DO_reg[8]/NET0131  & n5968 ;
  assign n31308 = \sport0_regs_AUTOreg_DO_reg[3]/NET0131  & n5970 ;
  assign n31311 = \sport0_regs_AUTOreg_DO_reg[8]/NET0131  & n4050 ;
  assign n31312 = ~n31308 & ~n31311 ;
  assign n31313 = ~n31310 & n31312 ;
  assign n31314 = ~n31309 & n31313 ;
  assign n31315 = ~n31307 & n31314 ;
  assign n31316 = n5692 & ~n31315 ;
  assign n31317 = ~n31306 & ~n31316 ;
  assign n31318 = \core_dag_ilm2reg_M_E_reg[0]/NET0131  & ~n5692 ;
  assign n31319 = n4055 & ~n25696 ;
  assign n31321 = \sport1_regs_AUTOreg_DO_reg[2]/NET0131  & n5966 ;
  assign n31322 = \sport1_regs_AUTOreg_DO_reg[7]/NET0131  & n5968 ;
  assign n31320 = \sport0_regs_AUTOreg_DO_reg[7]/NET0131  & n4050 ;
  assign n31323 = \sport0_regs_AUTOreg_DO_reg[2]/NET0131  & n5970 ;
  assign n31324 = ~n31320 & ~n31323 ;
  assign n31325 = ~n31322 & n31324 ;
  assign n31326 = ~n31321 & n31325 ;
  assign n31327 = ~n31319 & n31326 ;
  assign n31328 = n5692 & ~n31327 ;
  assign n31329 = ~n31318 & ~n31328 ;
  assign n31332 = ~n26060 & ~n31329 ;
  assign n31333 = ~n26075 & n31329 ;
  assign n31334 = ~n31332 & ~n31333 ;
  assign n31335 = n31317 & ~n31334 ;
  assign n31330 = ~n31317 & n31329 ;
  assign n31331 = ~n26059 & n31330 ;
  assign n31336 = ~n31317 & ~n31329 ;
  assign n31337 = ~n26074 & n31336 ;
  assign n31338 = ~n31331 & ~n31337 ;
  assign n31339 = ~n31335 & n31338 ;
  assign n31340 = n10289 & n31339 ;
  assign n31343 = \core_dag_ilm2reg_M7_we_DO_reg[9]/NET0131  & n31337 ;
  assign n31346 = \core_dag_ilm2reg_M6_we_DO_reg[9]/NET0131  & n31331 ;
  assign n31347 = ~n31343 & ~n31346 ;
  assign n31348 = ~n21579 & n31347 ;
  assign n31341 = n31317 & n31332 ;
  assign n31342 = \core_dag_ilm2reg_M5_we_DO_reg[9]/NET0131  & n31341 ;
  assign n31344 = n31317 & n31333 ;
  assign n31345 = \core_dag_ilm2reg_M4_we_DO_reg[9]/NET0131  & n31344 ;
  assign n31349 = ~n31342 & ~n31345 ;
  assign n31350 = n31348 & n31349 ;
  assign n31351 = ~n31340 & n31350 ;
  assign n31352 = ~\core_dag_ilm2reg_M_reg[9]/NET0131  & n21579 ;
  assign n31353 = ~n31351 & ~n31352 ;
  assign n31354 = n9178 & n31339 ;
  assign n31356 = \core_dag_ilm2reg_M7_we_DO_reg[12]/NET0131  & n31337 ;
  assign n31358 = \core_dag_ilm2reg_M6_we_DO_reg[12]/NET0131  & n31331 ;
  assign n31359 = ~n31356 & ~n31358 ;
  assign n31360 = ~n21579 & n31359 ;
  assign n31355 = \core_dag_ilm2reg_M5_we_DO_reg[12]/NET0131  & n31341 ;
  assign n31357 = \core_dag_ilm2reg_M4_we_DO_reg[12]/NET0131  & n31344 ;
  assign n31361 = ~n31355 & ~n31357 ;
  assign n31362 = n31360 & n31361 ;
  assign n31363 = ~n31354 & n31362 ;
  assign n31364 = ~\core_dag_ilm2reg_M_reg[12]/NET0131  & n21579 ;
  assign n31365 = ~n31363 & ~n31364 ;
  assign n31366 = n8460 & n31339 ;
  assign n31368 = \core_dag_ilm2reg_M7_we_DO_reg[11]/NET0131  & n31337 ;
  assign n31370 = \core_dag_ilm2reg_M6_we_DO_reg[11]/NET0131  & n31331 ;
  assign n31371 = ~n31368 & ~n31370 ;
  assign n31372 = ~n21579 & n31371 ;
  assign n31367 = \core_dag_ilm2reg_M5_we_DO_reg[11]/NET0131  & n31341 ;
  assign n31369 = \core_dag_ilm2reg_M4_we_DO_reg[11]/NET0131  & n31344 ;
  assign n31373 = ~n31367 & ~n31369 ;
  assign n31374 = n31372 & n31373 ;
  assign n31375 = ~n31366 & n31374 ;
  assign n31376 = ~\core_dag_ilm2reg_M_reg[11]/NET0131  & n21579 ;
  assign n31377 = ~n31375 & ~n31376 ;
  assign n31378 = n7859 & n31339 ;
  assign n31380 = \core_dag_ilm2reg_M7_we_DO_reg[10]/NET0131  & n31337 ;
  assign n31382 = \core_dag_ilm2reg_M6_we_DO_reg[10]/NET0131  & n31331 ;
  assign n31383 = ~n31380 & ~n31382 ;
  assign n31384 = ~n21579 & n31383 ;
  assign n31379 = \core_dag_ilm2reg_M5_we_DO_reg[10]/NET0131  & n31341 ;
  assign n31381 = \core_dag_ilm2reg_M4_we_DO_reg[10]/NET0131  & n31344 ;
  assign n31385 = ~n31379 & ~n31381 ;
  assign n31386 = n31384 & n31385 ;
  assign n31387 = ~n31378 & n31386 ;
  assign n31388 = ~\core_dag_ilm2reg_M_reg[10]/NET0131  & n21579 ;
  assign n31389 = ~n31387 & ~n31388 ;
  assign n31390 = \core_c_dec_IRE_reg[1]/NET0131  & ~n5692 ;
  assign n31391 = \core_c_dec_IR_reg[1]/NET0131  & n4055 ;
  assign n31392 = n31314 & ~n31391 ;
  assign n31393 = n5692 & ~n31392 ;
  assign n31394 = ~n31390 & ~n31393 ;
  assign n31395 = \core_c_dec_IRE_reg[0]/NET0131  & ~n5692 ;
  assign n31396 = \core_c_dec_IR_reg[0]/NET0131  & n4055 ;
  assign n31397 = n31326 & ~n31396 ;
  assign n31398 = n5692 & ~n31397 ;
  assign n31399 = ~n31395 & ~n31398 ;
  assign n31402 = ~n26080 & n31399 ;
  assign n31403 = ~n26076 & ~n31399 ;
  assign n31404 = ~n31402 & ~n31403 ;
  assign n31405 = n31394 & ~n31404 ;
  assign n31400 = ~n31394 & n31399 ;
  assign n31401 = ~n26079 & n31400 ;
  assign n31406 = ~n31394 & ~n31399 ;
  assign n31407 = ~n26077 & n31406 ;
  assign n31408 = ~n31401 & ~n31407 ;
  assign n31409 = ~n31405 & n31408 ;
  assign n31410 = n10289 & n31409 ;
  assign n31413 = \core_dag_ilm1reg_M3_we_DO_reg[9]/NET0131  & n31407 ;
  assign n31416 = \core_dag_ilm1reg_M2_we_DO_reg[9]/NET0131  & n31401 ;
  assign n31417 = ~n31413 & ~n31416 ;
  assign n31418 = ~n21592 & n31417 ;
  assign n31411 = n31394 & n31402 ;
  assign n31412 = \core_dag_ilm1reg_M0_we_DO_reg[9]/NET0131  & n31411 ;
  assign n31414 = n31394 & n31403 ;
  assign n31415 = \core_dag_ilm1reg_M1_we_DO_reg[9]/NET0131  & n31414 ;
  assign n31419 = ~n31412 & ~n31415 ;
  assign n31420 = n31418 & n31419 ;
  assign n31421 = ~n31410 & n31420 ;
  assign n31422 = ~\core_dag_ilm1reg_M_reg[9]/NET0131  & n21592 ;
  assign n31423 = ~n31421 & ~n31422 ;
  assign n31424 = n10638 & n31409 ;
  assign n31426 = \core_dag_ilm1reg_M3_we_DO_reg[8]/NET0131  & n31407 ;
  assign n31428 = \core_dag_ilm1reg_M2_we_DO_reg[8]/NET0131  & n31401 ;
  assign n31429 = ~n31426 & ~n31428 ;
  assign n31430 = ~n21592 & n31429 ;
  assign n31425 = \core_dag_ilm1reg_M0_we_DO_reg[8]/NET0131  & n31411 ;
  assign n31427 = \core_dag_ilm1reg_M1_we_DO_reg[8]/NET0131  & n31414 ;
  assign n31431 = ~n31425 & ~n31427 ;
  assign n31432 = n31430 & n31431 ;
  assign n31433 = ~n31424 & n31432 ;
  assign n31434 = ~\core_dag_ilm1reg_M_reg[8]/NET0131  & n21592 ;
  assign n31435 = ~n31433 & ~n31434 ;
  assign n31436 = n7340 & n31409 ;
  assign n31438 = \core_dag_ilm1reg_M3_we_DO_reg[13]/NET0131  & n31407 ;
  assign n31440 = \core_dag_ilm1reg_M2_we_DO_reg[13]/NET0131  & n31401 ;
  assign n31441 = ~n31438 & ~n31440 ;
  assign n31442 = ~n21592 & n31441 ;
  assign n31437 = \core_dag_ilm1reg_M0_we_DO_reg[13]/NET0131  & n31411 ;
  assign n31439 = \core_dag_ilm1reg_M1_we_DO_reg[13]/NET0131  & n31414 ;
  assign n31443 = ~n31437 & ~n31439 ;
  assign n31444 = n31442 & n31443 ;
  assign n31445 = ~n31436 & n31444 ;
  assign n31446 = ~\core_dag_ilm1reg_M_reg[13]/NET0131  & n21592 ;
  assign n31447 = ~n31445 & ~n31446 ;
  assign n31448 = n8460 & n31409 ;
  assign n31450 = \core_dag_ilm1reg_M3_we_DO_reg[11]/NET0131  & n31407 ;
  assign n31452 = \core_dag_ilm1reg_M2_we_DO_reg[11]/NET0131  & n31401 ;
  assign n31453 = ~n31450 & ~n31452 ;
  assign n31454 = ~n21592 & n31453 ;
  assign n31449 = \core_dag_ilm1reg_M0_we_DO_reg[11]/NET0131  & n31411 ;
  assign n31451 = \core_dag_ilm1reg_M1_we_DO_reg[11]/NET0131  & n31414 ;
  assign n31455 = ~n31449 & ~n31451 ;
  assign n31456 = n31454 & n31455 ;
  assign n31457 = ~n31448 & n31456 ;
  assign n31458 = ~\core_dag_ilm1reg_M_reg[11]/NET0131  & n21592 ;
  assign n31459 = ~n31457 & ~n31458 ;
  assign n31460 = n7859 & n31409 ;
  assign n31462 = \core_dag_ilm1reg_M3_we_DO_reg[10]/NET0131  & n31407 ;
  assign n31464 = \core_dag_ilm1reg_M2_we_DO_reg[10]/NET0131  & n31401 ;
  assign n31465 = ~n31462 & ~n31464 ;
  assign n31466 = ~n21592 & n31465 ;
  assign n31461 = \core_dag_ilm1reg_M0_we_DO_reg[10]/NET0131  & n31411 ;
  assign n31463 = \core_dag_ilm1reg_M1_we_DO_reg[10]/NET0131  & n31414 ;
  assign n31467 = ~n31461 & ~n31463 ;
  assign n31468 = n31466 & n31467 ;
  assign n31469 = ~n31460 & n31468 ;
  assign n31470 = ~\core_dag_ilm1reg_M_reg[10]/NET0131  & n21592 ;
  assign n31471 = ~n31469 & ~n31470 ;
  assign n31473 = n19499 & ~n19848 ;
  assign n31472 = ~\core_eu_em_mac_em_reg_mr1swe_DO_reg[10]/P0001  & ~n19499 ;
  assign n31474 = n19501 & ~n31472 ;
  assign n31475 = ~n31473 & n31474 ;
  assign n31476 = \core_eu_em_mac_em_reg_mr1swe_DO_reg[10]/P0001  & ~n19383 ;
  assign n31477 = ~n19508 & ~n31476 ;
  assign n31478 = ~n31475 & n31477 ;
  assign n31479 = ~n18262 & ~n31478 ;
  assign n31480 = ~\core_c_psq_MSTAT_reg_DO_reg[4]/NET0131  & ~n19516 ;
  assign n31481 = \core_c_psq_MSTAT_reg_DO_reg[4]/NET0131  & n19434 ;
  assign n31482 = ~n31480 & ~n31481 ;
  assign n31483 = n18262 & ~n31482 ;
  assign n31484 = ~n31479 & ~n31483 ;
  assign n31485 = n14752 & n31482 ;
  assign n31486 = n19776 & n19848 ;
  assign n31487 = \core_eu_em_mac_em_reg_mr1rwe_DO_reg[10]/P0001  & ~n17809 ;
  assign n31488 = n19780 & ~n31487 ;
  assign n31489 = ~n31486 & n31488 ;
  assign n31490 = ~n31485 & ~n31489 ;
  assign n31522 = \clkc_STDcnt_reg[0]/NET0131  & \clkc_STDcnt_reg[1]/NET0131  ;
  assign n31523 = \clkc_STDcnt_reg[2]/NET0131  & n31522 ;
  assign n31524 = \clkc_STDcnt_reg[3]/NET0131  & n31523 ;
  assign n31525 = \clkc_STDcnt_reg[4]/NET0131  & n31524 ;
  assign n31526 = \clkc_STDcnt_reg[5]/NET0131  & n31525 ;
  assign n31527 = \clkc_STDcnt_reg[6]/NET0131  & n31526 ;
  assign n31528 = \clkc_STDcnt_reg[7]/NET0131  & n31527 ;
  assign n31529 = \clkc_STDcnt_reg[8]/NET0131  & n31528 ;
  assign n31530 = \clkc_STDcnt_reg[9]/NET0131  & n31529 ;
  assign n31532 = \clkc_STDcnt_reg[10]/NET0131  & n31530 ;
  assign n31491 = ~\clkc_STDcnt_reg[8]/NET0131  & \clkc_ckr_reg_DO_reg[5]/NET0131  ;
  assign n31495 = \clkc_STDcnt_reg[7]/NET0131  & ~\clkc_ckr_reg_DO_reg[4]/NET0131  ;
  assign n31509 = ~n31491 & ~n31495 ;
  assign n31496 = ~\clkc_STDcnt_reg[7]/NET0131  & \clkc_ckr_reg_DO_reg[4]/NET0131  ;
  assign n31500 = ~\clkc_STDcnt_reg[5]/NET0131  & \clkc_ckr_reg_DO_reg[2]/NET0131  ;
  assign n31510 = ~n31496 & ~n31500 ;
  assign n31517 = n31509 & n31510 ;
  assign n31492 = ~\clkc_STDcnt_reg[9]/NET0131  & ~\clkc_ckr_reg_DO_reg[6]/NET0131  ;
  assign n31493 = \clkc_STDcnt_reg[9]/NET0131  & \clkc_ckr_reg_DO_reg[6]/NET0131  ;
  assign n31494 = ~n31492 & ~n31493 ;
  assign n31497 = ~\clkc_STDcnt_reg[10]/NET0131  & ~\clkc_ckr_reg_DO_reg[7]/NET0131  ;
  assign n31498 = \clkc_STDcnt_reg[10]/NET0131  & \clkc_ckr_reg_DO_reg[7]/NET0131  ;
  assign n31499 = ~n31497 & ~n31498 ;
  assign n31518 = ~n31494 & ~n31499 ;
  assign n31519 = n31517 & n31518 ;
  assign n31505 = \clkc_STDcnt_reg[3]/NET0131  & ~\clkc_ckr_reg_DO_reg[0]/NET0131  ;
  assign n31506 = \clkc_STDcnt_reg[6]/NET0131  & ~\clkc_ckr_reg_DO_reg[3]/NET0131  ;
  assign n31513 = ~n31505 & ~n31506 ;
  assign n31507 = ~\clkc_STDcnt_reg[3]/NET0131  & \clkc_ckr_reg_DO_reg[0]/NET0131  ;
  assign n31508 = \clkc_STDcnt_reg[8]/NET0131  & ~\clkc_ckr_reg_DO_reg[5]/NET0131  ;
  assign n31514 = ~n31507 & ~n31508 ;
  assign n31515 = n31513 & n31514 ;
  assign n31501 = \clkc_STDcnt_reg[5]/NET0131  & ~\clkc_ckr_reg_DO_reg[2]/NET0131  ;
  assign n31502 = \clkc_STDcnt_reg[4]/NET0131  & ~\clkc_ckr_reg_DO_reg[1]/NET0131  ;
  assign n31511 = ~n31501 & ~n31502 ;
  assign n31503 = ~\clkc_STDcnt_reg[4]/NET0131  & \clkc_ckr_reg_DO_reg[1]/NET0131  ;
  assign n31504 = ~\clkc_STDcnt_reg[6]/NET0131  & \clkc_ckr_reg_DO_reg[3]/NET0131  ;
  assign n31512 = ~n31503 & ~n31504 ;
  assign n31516 = n31511 & n31512 ;
  assign n31520 = n31515 & n31516 ;
  assign n31521 = n31519 & n31520 ;
  assign n31531 = ~\clkc_STDcnt_reg[10]/NET0131  & ~n31530 ;
  assign n31533 = ~n31521 & ~n31531 ;
  assign n31534 = ~n31532 & n31533 ;
  assign n31535 = \core_c_psq_Iact_E_reg[6]/NET0131  & ~n4116 ;
  assign n31536 = ~\sport0_regs_AUTOreg_DO_reg[1]/NET0131  & \sport0_txctl_c_sync1_reg/P0001  ;
  assign n31537 = ~\sport0_txctl_c_sync2_reg/P0001  & n31536 ;
  assign n31538 = \core_dag_modulo1_T0wrap_reg/P0001  & \sport0_regs_AUTOreg_DO_reg[1]/NET0131  ;
  assign n31539 = ~\core_c_psq_IFC_reg[14]/NET0131  & ~\core_c_psq_Iflag_reg[6]/NET0131  ;
  assign n31540 = ~n31538 & n31539 ;
  assign n31541 = ~n31537 & n31540 ;
  assign n31542 = ~\core_c_psq_IFC_reg[6]/NET0131  & ~n31541 ;
  assign n31543 = ~n31535 & n31542 ;
  assign n31545 = ~n31076 & n31079 ;
  assign n31546 = n31103 & n31545 ;
  assign n31547 = n6023 & n6025 ;
  assign n31548 = ~n4117 & ~n31547 ;
  assign n31549 = ~n31546 & n31548 ;
  assign n31544 = ~\core_c_dec_MTMX1_E_reg/P0001  & n4117 ;
  assign n31550 = n4116 & ~n31544 ;
  assign n31551 = ~n31549 & n31550 ;
  assign n31553 = n31112 & n31545 ;
  assign n31554 = n6023 & n19697 ;
  assign n31555 = ~n4117 & ~n31554 ;
  assign n31556 = ~n31553 & n31555 ;
  assign n31552 = ~\core_c_dec_MTMX0_E_reg/P0001  & n4117 ;
  assign n31557 = n4116 & ~n31552 ;
  assign n31558 = ~n31556 & n31557 ;
  assign n31562 = n31094 & n31121 ;
  assign n31561 = n31079 & ~n31089 ;
  assign n31563 = ~n31098 & n31561 ;
  assign n31564 = n31562 & n31563 ;
  assign n31560 = n6023 & n20606 ;
  assign n31565 = ~n4117 & ~n31560 ;
  assign n31566 = ~n31564 & n31565 ;
  assign n31559 = ~\core_c_dec_MTAX1_E_reg/P0001  & n4117 ;
  assign n31567 = n4116 & ~n31559 ;
  assign n31568 = ~n31566 & n31567 ;
  assign n31569 = ~\sport0_cfg_SCLKi_cnt_reg[14]/NET0131  & ~n19552 ;
  assign n31570 = n19197 & ~n29228 ;
  assign n31571 = ~n31569 & n31570 ;
  assign n31572 = ~\core_c_psq_MSTAT_reg_DO_reg[4]/NET0131  & n17789 ;
  assign n31573 = \core_c_psq_MSTAT_reg_DO_reg[4]/NET0131  & n25067 ;
  assign n31574 = ~n31572 & ~n31573 ;
  assign n31575 = ~\sport1_cfg_SCLKi_cnt_reg[14]/NET0131  & ~n20253 ;
  assign n31576 = n19130 & ~n29407 ;
  assign n31577 = ~n31575 & n31576 ;
  assign n31580 = n31098 & n31561 ;
  assign n31581 = ~n4117 & n31580 ;
  assign n31582 = n31562 & n31581 ;
  assign n31578 = n6116 & n25725 ;
  assign n31579 = \core_c_dec_MTAX0_E_reg/P0001  & n4117 ;
  assign n31583 = ~n31578 & ~n31579 ;
  assign n31584 = ~n31582 & n31583 ;
  assign n31585 = n4116 & ~n31584 ;
  assign n31586 = ~\sport1_cfg_FSi_reg/NET0131  & ~n28854 ;
  assign n31598 = ~\sport1_cfg_FSi_cnt_reg[2]/NET0131  & \sport1_regs_SCTLreg_DO_reg[2]/NET0131  ;
  assign n31599 = \sport1_cfg_FSi_cnt_reg[0]/NET0131  & ~\sport1_regs_SCTLreg_DO_reg[0]/NET0131  ;
  assign n31605 = ~n31598 & ~n31599 ;
  assign n31600 = \sport1_cfg_FSi_cnt_reg[3]/NET0131  & ~\sport1_regs_SCTLreg_DO_reg[3]/NET0131  ;
  assign n31601 = ~\sport1_cfg_FSi_cnt_reg[3]/NET0131  & \sport1_regs_SCTLreg_DO_reg[3]/NET0131  ;
  assign n31606 = ~n31600 & ~n31601 ;
  assign n31607 = n31605 & n31606 ;
  assign n31592 = ~\sport1_cfg_FSi_cnt_reg[1]/NET0131  & \sport1_regs_SCTLreg_DO_reg[1]/NET0131  ;
  assign n31593 = \sport1_cfg_FSi_cnt_reg[4]/NET0131  & ~\sport1_regs_MWORDreg_DO_reg[10]/NET0131  ;
  assign n31602 = ~n31592 & ~n31593 ;
  assign n31594 = \sport1_cfg_FSi_cnt_reg[1]/NET0131  & ~\sport1_regs_SCTLreg_DO_reg[1]/NET0131  ;
  assign n31595 = ~\sport1_cfg_FSi_cnt_reg[4]/NET0131  & \sport1_regs_MWORDreg_DO_reg[10]/NET0131  ;
  assign n31603 = ~n31594 & ~n31595 ;
  assign n31596 = \sport1_cfg_FSi_cnt_reg[2]/NET0131  & ~\sport1_regs_SCTLreg_DO_reg[2]/NET0131  ;
  assign n31597 = ~\sport1_cfg_FSi_cnt_reg[0]/NET0131  & \sport1_regs_SCTLreg_DO_reg[0]/NET0131  ;
  assign n31604 = ~n31596 & ~n31597 ;
  assign n31608 = n31603 & n31604 ;
  assign n31609 = n31602 & n31608 ;
  assign n31610 = n31607 & n31609 ;
  assign n31587 = \sport1_cfg_FSi_cnt_reg[0]/NET0131  & \sport1_cfg_FSi_cnt_reg[1]/NET0131  ;
  assign n31588 = \sport1_cfg_FSi_cnt_reg[2]/NET0131  & \sport1_cfg_FSi_cnt_reg[3]/NET0131  ;
  assign n31589 = ~\sport1_cfg_FSi_cnt_reg[4]/NET0131  & \sport1_regs_MWORDreg_DO_reg[9]/NET0131  ;
  assign n31590 = n31588 & n31589 ;
  assign n31591 = n31587 & n31590 ;
  assign n31611 = \sport1_cfg_SP_ENg_reg/NET0131  & \sport1_regs_SCTLreg_DO_reg[10]/NET0131  ;
  assign n31612 = ~n31591 & n31611 ;
  assign n31613 = ~n31610 & n31612 ;
  assign n31614 = \sport1_cfg_FSi_reg/NET0131  & ~n31613 ;
  assign n31615 = ~n31586 & ~n31614 ;
  assign n31616 = ~\sport0_cfg_FSi_reg/NET0131  & ~n28944 ;
  assign n31628 = ~\sport0_cfg_FSi_cnt_reg[2]/NET0131  & \sport0_regs_SCTLreg_DO_reg[2]/NET0131  ;
  assign n31629 = \sport0_cfg_FSi_cnt_reg[0]/NET0131  & ~\sport0_regs_SCTLreg_DO_reg[0]/NET0131  ;
  assign n31635 = ~n31628 & ~n31629 ;
  assign n31630 = \sport0_cfg_FSi_cnt_reg[3]/NET0131  & ~\sport0_regs_SCTLreg_DO_reg[3]/NET0131  ;
  assign n31631 = ~\sport0_cfg_FSi_cnt_reg[3]/NET0131  & \sport0_regs_SCTLreg_DO_reg[3]/NET0131  ;
  assign n31636 = ~n31630 & ~n31631 ;
  assign n31637 = n31635 & n31636 ;
  assign n31622 = ~\sport0_cfg_FSi_cnt_reg[1]/NET0131  & \sport0_regs_SCTLreg_DO_reg[1]/NET0131  ;
  assign n31623 = \sport0_cfg_FSi_cnt_reg[4]/NET0131  & ~\sport0_regs_MWORDreg_DO_reg[10]/NET0131  ;
  assign n31632 = ~n31622 & ~n31623 ;
  assign n31624 = \sport0_cfg_FSi_cnt_reg[1]/NET0131  & ~\sport0_regs_SCTLreg_DO_reg[1]/NET0131  ;
  assign n31625 = ~\sport0_cfg_FSi_cnt_reg[4]/NET0131  & \sport0_regs_MWORDreg_DO_reg[10]/NET0131  ;
  assign n31633 = ~n31624 & ~n31625 ;
  assign n31626 = \sport0_cfg_FSi_cnt_reg[2]/NET0131  & ~\sport0_regs_SCTLreg_DO_reg[2]/NET0131  ;
  assign n31627 = ~\sport0_cfg_FSi_cnt_reg[0]/NET0131  & \sport0_regs_SCTLreg_DO_reg[0]/NET0131  ;
  assign n31634 = ~n31626 & ~n31627 ;
  assign n31638 = n31633 & n31634 ;
  assign n31639 = n31632 & n31638 ;
  assign n31640 = n31637 & n31639 ;
  assign n31617 = \sport0_cfg_FSi_cnt_reg[0]/NET0131  & \sport0_cfg_FSi_cnt_reg[1]/NET0131  ;
  assign n31618 = \sport0_cfg_FSi_cnt_reg[2]/NET0131  & \sport0_cfg_FSi_cnt_reg[3]/NET0131  ;
  assign n31619 = ~\sport0_cfg_FSi_cnt_reg[4]/NET0131  & \sport0_regs_MWORDreg_DO_reg[9]/NET0131  ;
  assign n31620 = n31618 & n31619 ;
  assign n31621 = n31617 & n31620 ;
  assign n31641 = \sport0_cfg_SP_ENg_reg/NET0131  & \sport0_regs_SCTLreg_DO_reg[10]/NET0131  ;
  assign n31642 = ~n31621 & n31641 ;
  assign n31643 = ~n31640 & n31642 ;
  assign n31644 = \sport0_cfg_FSi_reg/NET0131  & ~n31643 ;
  assign n31645 = ~n31616 & ~n31644 ;
  assign n31646 = \core_c_dec_pMFSHT_Ei_reg/NET0131  & n4117 ;
  assign n31647 = ~n30966 & n30969 ;
  assign n31648 = n30970 & n31647 ;
  assign n31653 = \core_c_dec_IR_reg[1]/NET0131  & \core_c_dec_IR_reg[2]/NET0131  ;
  assign n31654 = n31264 & n31653 ;
  assign n31655 = n31271 & n31654 ;
  assign n31657 = ~n31648 & ~n31655 ;
  assign n31650 = n30958 & n30961 ;
  assign n31651 = ~n30966 & n31650 ;
  assign n31656 = n30974 & n31651 ;
  assign n31649 = n30974 & n31647 ;
  assign n31652 = n30970 & n31651 ;
  assign n31658 = ~n31649 & ~n31652 ;
  assign n31659 = ~n31656 & n31658 ;
  assign n31660 = n31657 & n31659 ;
  assign n31661 = n30934 & ~n31660 ;
  assign n31662 = ~n31646 & ~n31661 ;
  assign n31663 = \core_c_dec_MFSHT_Ei_reg/NET0131  & n4117 ;
  assign n31664 = n25047 & ~n31660 ;
  assign n31665 = ~n31663 & ~n31664 ;
  assign n31666 = \tm_tsr_reg_DO_reg[4]/NET0131  & ~n25491 ;
  assign n31667 = \tm_TSR_TMP_reg[4]/NET0131  & ~n25493 ;
  assign n31668 = ~n25494 & ~n31667 ;
  assign n31669 = n25491 & ~n31668 ;
  assign n31670 = ~n31666 & ~n31669 ;
  assign n31671 = \sport0_regs_FSDIVreg_DO_reg[7]/NET0131  & n28876 ;
  assign n31672 = ~\sport0_cfg_FSi_cnt_reg[7]/NET0131  & ~n28952 ;
  assign n31673 = ~n28953 & ~n31672 ;
  assign n31674 = n28945 & n31673 ;
  assign n31675 = ~n31671 & ~n31674 ;
  assign n31676 = \sport1_regs_FSDIVreg_DO_reg[7]/NET0131  & n28786 ;
  assign n31677 = ~\sport1_cfg_FSi_cnt_reg[7]/NET0131  & ~n28862 ;
  assign n31678 = ~n28863 & ~n31677 ;
  assign n31679 = n28855 & n31678 ;
  assign n31680 = ~n31676 & ~n31679 ;
  assign n31681 = \sport1_regs_FSDIVreg_DO_reg[8]/NET0131  & n28786 ;
  assign n31682 = ~\sport1_cfg_FSi_cnt_reg[8]/NET0131  & ~n28863 ;
  assign n31683 = n28855 & ~n28864 ;
  assign n31684 = ~n31682 & n31683 ;
  assign n31685 = ~n31681 & ~n31684 ;
  assign n31686 = \sport0_regs_FSDIVreg_DO_reg[8]/NET0131  & n28876 ;
  assign n31687 = ~\sport0_cfg_FSi_cnt_reg[8]/NET0131  & ~n28953 ;
  assign n31688 = n28945 & ~n28954 ;
  assign n31689 = ~n31687 & n31688 ;
  assign n31690 = ~n31686 & ~n31689 ;
  assign n31696 = ~\sport1_rxctl_RCS_reg[0]/NET0131  & ~\sport1_rxctl_RCS_reg[2]/NET0131  ;
  assign n31697 = \sport1_rxctl_RCS_reg[1]/NET0131  & n31696 ;
  assign n31698 = \sport1_rxctl_RCS_reg[0]/NET0131  & \sport1_rxctl_RCS_reg[2]/NET0131  ;
  assign n31699 = ~\sport1_rxctl_RCS_reg[1]/NET0131  & ~n31696 ;
  assign n31700 = ~n31698 & n31699 ;
  assign n31701 = ~n30750 & n31700 ;
  assign n31702 = ~n31697 & ~n31701 ;
  assign n31691 = ~\sport1_rxctl_Bcnt_reg[0]/NET0131  & ~\sport1_rxctl_Bcnt_reg[1]/NET0131  ;
  assign n31692 = ~\sport1_rxctl_Bcnt_reg[2]/NET0131  & n31691 ;
  assign n31693 = ~\sport1_rxctl_Bcnt_reg[3]/NET0131  & n31692 ;
  assign n31703 = ~\sport1_rxctl_Bcnt_reg[4]/NET0131  & n31693 ;
  assign n31704 = ~n31701 & n31703 ;
  assign n31705 = ~n31702 & ~n31704 ;
  assign n31707 = \sport1_regs_SCTLreg_DO_reg[3]/NET0131  & ~n31705 ;
  assign n31694 = \sport1_rxctl_Bcnt_reg[3]/NET0131  & ~n31692 ;
  assign n31695 = ~n31693 & ~n31694 ;
  assign n31706 = ~n31695 & n31705 ;
  assign n31708 = ~\sport1_rxctl_TAG_SLOT_reg/P0001  & ~n31706 ;
  assign n31709 = ~n31707 & n31708 ;
  assign n31711 = \sport1_rxctl_Bcnt_reg[2]/NET0131  & ~n31691 ;
  assign n31712 = ~n31692 & ~n31711 ;
  assign n31713 = n31705 & ~n31712 ;
  assign n31710 = \sport1_regs_SCTLreg_DO_reg[2]/NET0131  & ~n31705 ;
  assign n31714 = ~\sport1_rxctl_TAG_SLOT_reg/P0001  & ~n31710 ;
  assign n31715 = ~n31713 & n31714 ;
  assign n31717 = \sport1_rxctl_Bcnt_reg[0]/NET0131  & \sport1_rxctl_Bcnt_reg[1]/NET0131  ;
  assign n31718 = ~n31691 & ~n31717 ;
  assign n31719 = n31705 & ~n31718 ;
  assign n31716 = \sport1_regs_SCTLreg_DO_reg[1]/NET0131  & ~n31705 ;
  assign n31720 = ~\sport1_rxctl_TAG_SLOT_reg/P0001  & ~n31716 ;
  assign n31721 = ~n31719 & n31720 ;
  assign n31723 = \sport1_regs_SCTLreg_DO_reg[0]/NET0131  & ~n31705 ;
  assign n31722 = ~\sport1_rxctl_Bcnt_reg[0]/NET0131  & n31705 ;
  assign n31724 = ~\sport1_rxctl_TAG_SLOT_reg/P0001  & ~n31722 ;
  assign n31725 = ~n31723 & n31724 ;
  assign n31726 = n11525 & n31339 ;
  assign n31729 = \core_dag_ilm2reg_M4_we_DO_reg[6]/NET0131  & n31344 ;
  assign n31727 = \core_dag_ilm2reg_M5_we_DO_reg[6]/NET0131  & n31341 ;
  assign n31728 = \core_dag_ilm2reg_M6_we_DO_reg[6]/NET0131  & n31331 ;
  assign n31730 = \core_dag_ilm2reg_M7_we_DO_reg[6]/NET0131  & n31337 ;
  assign n31731 = ~n31728 & ~n31730 ;
  assign n31732 = ~n31727 & n31731 ;
  assign n31733 = ~n31729 & n31732 ;
  assign n31734 = ~n31726 & n31733 ;
  assign n31735 = n10911 & n31339 ;
  assign n31738 = \core_dag_ilm2reg_M4_we_DO_reg[5]/NET0131  & n31344 ;
  assign n31736 = \core_dag_ilm2reg_M5_we_DO_reg[5]/NET0131  & n31341 ;
  assign n31737 = \core_dag_ilm2reg_M6_we_DO_reg[5]/NET0131  & n31331 ;
  assign n31739 = \core_dag_ilm2reg_M7_we_DO_reg[5]/NET0131  & n31337 ;
  assign n31740 = ~n31737 & ~n31739 ;
  assign n31741 = ~n31736 & n31740 ;
  assign n31742 = ~n31738 & n31741 ;
  assign n31743 = ~n31735 & n31742 ;
  assign n31744 = n10069 & n31339 ;
  assign n31747 = \core_dag_ilm2reg_M5_we_DO_reg[4]/NET0131  & n31341 ;
  assign n31745 = \core_dag_ilm2reg_M4_we_DO_reg[4]/NET0131  & n31344 ;
  assign n31746 = \core_dag_ilm2reg_M7_we_DO_reg[4]/NET0131  & n31337 ;
  assign n31748 = \core_dag_ilm2reg_M6_we_DO_reg[4]/NET0131  & n31331 ;
  assign n31749 = ~n31746 & ~n31748 ;
  assign n31750 = ~n31745 & n31749 ;
  assign n31751 = ~n31747 & n31750 ;
  assign n31752 = ~n31744 & n31751 ;
  assign n31753 = n8113 & n31339 ;
  assign n31756 = \core_dag_ilm2reg_M5_we_DO_reg[3]/NET0131  & n31341 ;
  assign n31754 = \core_dag_ilm2reg_M4_we_DO_reg[3]/NET0131  & n31344 ;
  assign n31755 = \core_dag_ilm2reg_M7_we_DO_reg[3]/NET0131  & n31337 ;
  assign n31757 = \core_dag_ilm2reg_M6_we_DO_reg[3]/NET0131  & n31331 ;
  assign n31758 = ~n31755 & ~n31757 ;
  assign n31759 = ~n31754 & n31758 ;
  assign n31760 = ~n31756 & n31759 ;
  assign n31761 = ~n31753 & n31760 ;
  assign n31762 = n8715 & n31339 ;
  assign n31765 = \core_dag_ilm2reg_M5_we_DO_reg[2]/NET0131  & n31341 ;
  assign n31763 = \core_dag_ilm2reg_M4_we_DO_reg[2]/NET0131  & n31344 ;
  assign n31764 = \core_dag_ilm2reg_M7_we_DO_reg[2]/NET0131  & n31337 ;
  assign n31766 = \core_dag_ilm2reg_M6_we_DO_reg[2]/NET0131  & n31331 ;
  assign n31767 = ~n31764 & ~n31766 ;
  assign n31768 = ~n31763 & n31767 ;
  assign n31769 = ~n31765 & n31768 ;
  assign n31770 = ~n31762 & n31769 ;
  assign n31771 = n9435 & n31339 ;
  assign n31774 = \core_dag_ilm2reg_M5_we_DO_reg[1]/NET0131  & n31341 ;
  assign n31772 = \core_dag_ilm2reg_M4_we_DO_reg[1]/NET0131  & n31344 ;
  assign n31773 = \core_dag_ilm2reg_M7_we_DO_reg[1]/NET0131  & n31337 ;
  assign n31775 = \core_dag_ilm2reg_M6_we_DO_reg[1]/NET0131  & n31331 ;
  assign n31776 = ~n31773 & ~n31775 ;
  assign n31777 = ~n31772 & n31776 ;
  assign n31778 = ~n31774 & n31777 ;
  assign n31779 = ~n31771 & n31778 ;
  assign n31780 = n8715 & n31409 ;
  assign n31783 = \core_dag_ilm1reg_M1_we_DO_reg[2]/NET0131  & n31414 ;
  assign n31781 = \core_dag_ilm1reg_M0_we_DO_reg[2]/NET0131  & n31411 ;
  assign n31782 = \core_dag_ilm1reg_M2_we_DO_reg[2]/NET0131  & n31401 ;
  assign n31784 = \core_dag_ilm1reg_M3_we_DO_reg[2]/NET0131  & n31407 ;
  assign n31785 = ~n31782 & ~n31784 ;
  assign n31786 = ~n31781 & n31785 ;
  assign n31787 = ~n31783 & n31786 ;
  assign n31788 = ~n31780 & n31787 ;
  assign n31789 = n9435 & n31409 ;
  assign n31792 = \core_dag_ilm1reg_M1_we_DO_reg[1]/NET0131  & n31414 ;
  assign n31790 = \core_dag_ilm1reg_M0_we_DO_reg[1]/NET0131  & n31411 ;
  assign n31791 = \core_dag_ilm1reg_M2_we_DO_reg[1]/NET0131  & n31401 ;
  assign n31793 = \core_dag_ilm1reg_M3_we_DO_reg[1]/NET0131  & n31407 ;
  assign n31794 = ~n31791 & ~n31793 ;
  assign n31795 = ~n31790 & n31794 ;
  assign n31796 = ~n31792 & n31795 ;
  assign n31797 = ~n31789 & n31796 ;
  assign n31798 = n7607 & n31409 ;
  assign n31801 = \core_dag_ilm1reg_M1_we_DO_reg[0]/NET0131  & n31414 ;
  assign n31799 = \core_dag_ilm1reg_M0_we_DO_reg[0]/NET0131  & n31411 ;
  assign n31800 = \core_dag_ilm1reg_M2_we_DO_reg[0]/NET0131  & n31401 ;
  assign n31802 = \core_dag_ilm1reg_M3_we_DO_reg[0]/NET0131  & n31407 ;
  assign n31803 = ~n31800 & ~n31802 ;
  assign n31804 = ~n31799 & n31803 ;
  assign n31805 = ~n31801 & n31804 ;
  assign n31806 = ~n31798 & n31805 ;
  assign n31807 = n11525 & n31409 ;
  assign n31810 = \core_dag_ilm1reg_M0_we_DO_reg[6]/NET0131  & n31411 ;
  assign n31808 = \core_dag_ilm1reg_M1_we_DO_reg[6]/NET0131  & n31414 ;
  assign n31809 = \core_dag_ilm1reg_M3_we_DO_reg[6]/NET0131  & n31407 ;
  assign n31811 = \core_dag_ilm1reg_M2_we_DO_reg[6]/NET0131  & n31401 ;
  assign n31812 = ~n31809 & ~n31811 ;
  assign n31813 = ~n31808 & n31812 ;
  assign n31814 = ~n31810 & n31813 ;
  assign n31815 = ~n31807 & n31814 ;
  assign n31816 = n10911 & n31409 ;
  assign n31819 = \core_dag_ilm1reg_M0_we_DO_reg[5]/NET0131  & n31411 ;
  assign n31817 = \core_dag_ilm1reg_M1_we_DO_reg[5]/NET0131  & n31414 ;
  assign n31818 = \core_dag_ilm1reg_M3_we_DO_reg[5]/NET0131  & n31407 ;
  assign n31820 = \core_dag_ilm1reg_M2_we_DO_reg[5]/NET0131  & n31401 ;
  assign n31821 = ~n31818 & ~n31820 ;
  assign n31822 = ~n31817 & n31821 ;
  assign n31823 = ~n31819 & n31822 ;
  assign n31824 = ~n31816 & n31823 ;
  assign n31825 = n10069 & n31409 ;
  assign n31828 = \core_dag_ilm1reg_M0_we_DO_reg[4]/NET0131  & n31411 ;
  assign n31826 = \core_dag_ilm1reg_M1_we_DO_reg[4]/NET0131  & n31414 ;
  assign n31827 = \core_dag_ilm1reg_M3_we_DO_reg[4]/NET0131  & n31407 ;
  assign n31829 = \core_dag_ilm1reg_M2_we_DO_reg[4]/NET0131  & n31401 ;
  assign n31830 = ~n31827 & ~n31829 ;
  assign n31831 = ~n31826 & n31830 ;
  assign n31832 = ~n31828 & n31831 ;
  assign n31833 = ~n31825 & n31832 ;
  assign n31834 = ~\sport0_cfg_SCLKi_cnt_reg[7]/NET0131  & ~n19544 ;
  assign n31835 = n19197 & ~n19545 ;
  assign n31836 = ~n31834 & n31835 ;
  assign n31837 = \core_eu_em_mac_em_reg_mfswe_DO_reg[10]/P0001  & ~n20864 ;
  assign n31838 = n20864 & ~n31482 ;
  assign n31839 = ~n31837 & ~n31838 ;
  assign n31840 = \core_c_dec_MACdep_Eg_reg/P0001  & n4117 ;
  assign n31841 = ~n26346 & ~n26371 ;
  assign n31842 = \core_c_dec_updMR_E_reg/P0001  & ~n31841 ;
  assign n31843 = \core_c_dec_updMF_E_reg/P0001  & n20470 ;
  assign n31844 = ~n26358 & n31843 ;
  assign n31845 = ~n31842 & ~n31844 ;
  assign n31846 = n18848 & ~n31845 ;
  assign n31847 = n13803 & n31846 ;
  assign n31848 = ~n31840 & ~n31847 ;
  assign n31849 = n4116 & ~n31848 ;
  assign n31851 = \sport1_rxctl_Bcnt_reg[4]/NET0131  & ~n31693 ;
  assign n31852 = ~n31703 & ~n31851 ;
  assign n31853 = n31705 & n31852 ;
  assign n31850 = ~\sport1_regs_MWORDreg_DO_reg[10]/NET0131  & ~n31705 ;
  assign n31854 = ~\sport1_rxctl_TAG_SLOT_reg/P0001  & ~n31850 ;
  assign n31855 = ~n31853 & n31854 ;
  assign n31856 = ~\sport0_rxctl_RCS_reg[0]/NET0131  & ~\sport0_rxctl_RCS_reg[2]/NET0131  ;
  assign n31857 = \sport0_rxctl_RCS_reg[1]/NET0131  & n31856 ;
  assign n31858 = \sport0_rxctl_RCS_reg[0]/NET0131  & \sport0_rxctl_RCS_reg[2]/NET0131  ;
  assign n31859 = ~\sport0_rxctl_RCS_reg[1]/NET0131  & ~n31856 ;
  assign n31860 = ~n31858 & n31859 ;
  assign n31861 = ~n30774 & n31860 ;
  assign n31862 = ~n31857 & ~n31861 ;
  assign n31863 = ~\sport0_rxctl_Bcnt_reg[0]/NET0131  & ~\sport0_rxctl_Bcnt_reg[1]/NET0131  ;
  assign n31864 = ~\sport0_rxctl_Bcnt_reg[2]/NET0131  & n31863 ;
  assign n31865 = ~\sport0_rxctl_Bcnt_reg[3]/NET0131  & n31864 ;
  assign n31866 = ~\sport0_rxctl_Bcnt_reg[4]/NET0131  & n31865 ;
  assign n31867 = ~n31861 & n31866 ;
  assign n31868 = ~n31862 & ~n31867 ;
  assign n31870 = \sport0_rxctl_Bcnt_reg[4]/NET0131  & ~n31865 ;
  assign n31871 = ~n31866 & ~n31870 ;
  assign n31872 = n31868 & n31871 ;
  assign n31869 = ~\sport0_regs_MWORDreg_DO_reg[10]/NET0131  & ~n31868 ;
  assign n31873 = ~\sport0_rxctl_TAG_SLOT_reg/P0001  & ~n31869 ;
  assign n31874 = ~n31872 & n31873 ;
  assign n31876 = \sport0_rxctl_Bcnt_reg[3]/NET0131  & ~n31864 ;
  assign n31877 = ~n31865 & ~n31876 ;
  assign n31878 = n31868 & ~n31877 ;
  assign n31875 = \sport0_regs_SCTLreg_DO_reg[3]/NET0131  & ~n31868 ;
  assign n31879 = ~\sport0_rxctl_TAG_SLOT_reg/P0001  & ~n31875 ;
  assign n31880 = ~n31878 & n31879 ;
  assign n31882 = \sport0_rxctl_Bcnt_reg[2]/NET0131  & ~n31863 ;
  assign n31883 = ~n31864 & ~n31882 ;
  assign n31884 = n31868 & ~n31883 ;
  assign n31881 = \sport0_regs_SCTLreg_DO_reg[2]/NET0131  & ~n31868 ;
  assign n31885 = ~\sport0_rxctl_TAG_SLOT_reg/P0001  & ~n31881 ;
  assign n31886 = ~n31884 & n31885 ;
  assign n31888 = \sport0_rxctl_Bcnt_reg[0]/NET0131  & \sport0_rxctl_Bcnt_reg[1]/NET0131  ;
  assign n31889 = ~n31863 & ~n31888 ;
  assign n31890 = n31868 & ~n31889 ;
  assign n31887 = \sport0_regs_SCTLreg_DO_reg[1]/NET0131  & ~n31868 ;
  assign n31891 = ~\sport0_rxctl_TAG_SLOT_reg/P0001  & ~n31887 ;
  assign n31892 = ~n31890 & n31891 ;
  assign n31894 = \sport0_regs_SCTLreg_DO_reg[0]/NET0131  & ~n31868 ;
  assign n31893 = ~\sport0_rxctl_Bcnt_reg[0]/NET0131  & n31868 ;
  assign n31895 = ~\sport0_rxctl_TAG_SLOT_reg/P0001  & ~n31893 ;
  assign n31896 = ~n31894 & n31895 ;
  assign n31897 = ~\sport1_cfg_SCLKi_cnt_reg[7]/NET0131  & ~n20236 ;
  assign n31898 = n19130 & ~n20237 ;
  assign n31899 = ~n31897 & n31898 ;
  assign n31900 = \core_c_psq_Iact_E_reg[5]/NET0131  & ~n4116 ;
  assign n31902 = \core_dag_modulo1_R0wrap_reg/P0001  & \sport0_regs_AUTOreg_DO_reg[0]/NET0131  ;
  assign n31901 = ~\sport0_regs_AUTOreg_DO_reg[0]/NET0131  & \sport0_rxctl_ISRa_reg/P0001  ;
  assign n31903 = ~\core_c_psq_IFC_reg[13]/NET0131  & ~\core_c_psq_Iflag_reg[5]/NET0131  ;
  assign n31904 = ~n31901 & n31903 ;
  assign n31905 = ~n31902 & n31904 ;
  assign n31906 = ~\core_c_psq_IFC_reg[5]/NET0131  & ~n31905 ;
  assign n31907 = ~n31900 & n31906 ;
  assign n31911 = ~\clkc_oscntr_reg_DO_reg[10]/NET0131  & ~\clkc_oscntr_reg_DO_reg[11]/NET0131  ;
  assign n31912 = ~\clkc_oscntr_reg_DO_reg[6]/NET0131  & ~\clkc_oscntr_reg_DO_reg[7]/NET0131  ;
  assign n31913 = n31911 & n31912 ;
  assign n31914 = \T_TMODE[0]_pad  & ~\clkc_oscntr_reg_DO_reg[5]/NET0131  ;
  assign n31915 = n31913 & n31914 ;
  assign n31916 = ~\T_TMODE[0]_pad  & \clkc_oscntr_reg_DO_reg[5]/NET0131  ;
  assign n31917 = \clkc_oscntr_reg_DO_reg[6]/NET0131  & n31916 ;
  assign n31918 = \clkc_oscntr_reg_DO_reg[11]/NET0131  & \clkc_oscntr_reg_DO_reg[8]/NET0131  ;
  assign n31919 = \clkc_oscntr_reg_DO_reg[9]/NET0131  & n31918 ;
  assign n31920 = n31917 & n31919 ;
  assign n31921 = ~n31915 & ~n31920 ;
  assign n31922 = ~\clkc_oscntr_reg_DO_reg[7]/NET0131  & \clkc_oscntr_reg_DO_reg[9]/NET0131  ;
  assign n31908 = \sport0_regs_AUTO_a_reg[14]/NET0131  & \sport0_regs_AUTO_a_reg[15]/NET0131  ;
  assign n31910 = ~\clkc_oscntr_reg_DO_reg[10]/NET0131  & \clkc_oscntr_reg_DO_reg[8]/NET0131  ;
  assign n31923 = n31908 & ~n31910 ;
  assign n31924 = ~n31922 & n31923 ;
  assign n31925 = n23418 & n31924 ;
  assign n31926 = ~n31921 & n31925 ;
  assign n31909 = \clkc_Cnt128_reg/NET0131  & ~n31908 ;
  assign n31927 = ~\clkc_Cnt4096_reg/NET0131  & ~n31909 ;
  assign n31928 = ~n31926 & n31927 ;
  assign n31929 = ~\clkc_Awake_reg/NET0131  & ~n31928 ;
  assign n31930 = n27915 & ~n28054 ;
  assign n31931 = \core_c_psq_CNTR_reg_DO_reg[13]/NET0131  & ~n27915 ;
  assign n31932 = ~n31930 & ~n31931 ;
  assign n31933 = \tm_tsr_reg_DO_reg[0]/NET0131  & ~n25491 ;
  assign n31934 = \core_c_psq_PCS_reg[3]/NET0131  & \tm_TSR_TMP_reg[0]/NET0131  ;
  assign n31935 = ~\core_c_psq_PCS_reg[3]/NET0131  & ~\tm_TSR_TMP_reg[0]/NET0131  ;
  assign n31936 = ~n31934 & ~n31935 ;
  assign n31937 = n25491 & ~n31936 ;
  assign n31938 = ~n31933 & ~n31937 ;
  assign n31941 = n18271 & ~n18974 ;
  assign n31940 = ~\core_eu_em_mac_em_reg_mr0swe_DO_reg[1]/P0001  & ~n18271 ;
  assign n31942 = n18273 & ~n31940 ;
  assign n31943 = ~n31941 & n31942 ;
  assign n31939 = \core_eu_em_mac_em_reg_mr0swe_DO_reg[1]/P0001  & ~n18266 ;
  assign n31944 = ~n18270 & ~n31939 ;
  assign n31945 = ~n31943 & n31944 ;
  assign n31946 = ~n18262 & ~n31945 ;
  assign n31947 = n18262 & n19667 ;
  assign n31948 = ~n31946 & ~n31947 ;
  assign n31949 = n14752 & ~n19667 ;
  assign n31950 = n18328 & n18974 ;
  assign n31951 = \core_eu_em_mac_em_reg_mr0rwe_DO_reg[1]/P0001  & ~n18330 ;
  assign n31952 = n18334 & ~n31951 ;
  assign n31953 = ~n31950 & n31952 ;
  assign n31954 = ~n31949 & ~n31953 ;
  assign n31955 = \core_eu_em_mac_em_reg_mfrwe_DO_reg[10]/P0001  & ~n20990 ;
  assign n31956 = n20990 & ~n31482 ;
  assign n31957 = ~n31955 & ~n31956 ;
  assign n31959 = \core_dag_modulo1_R1wrap_reg/P0001  & \sport1_regs_AUTOreg_DO_reg[0]/NET0131  ;
  assign n31958 = ~\sport1_regs_AUTOreg_DO_reg[0]/NET0131  & \sport1_rxctl_ISRa_reg/P0001  ;
  assign n31960 = ~\core_c_psq_IFC_reg[9]/NET0131  & ~n31958 ;
  assign n31961 = ~n31959 & n31960 ;
  assign n31962 = \memc_usysr_DO_reg[11]/NET0131  & ~n31961 ;
  assign n31963 = ~\core_c_psq_Iflag_reg[1]/NET0131  & ~n31962 ;
  assign n31964 = n21416 & ~n31963 ;
  assign n31965 = ~\core_c_dec_MFDAG1_Ei_reg/NET0131  & n4117 ;
  assign n31966 = ~n30936 & n31269 ;
  assign n31967 = ~\core_c_dec_IR_reg[2]/NET0131  & n31966 ;
  assign n31968 = \core_c_dec_IR_reg[3]/NET0131  & ~n31263 ;
  assign n31981 = n19301 & n31968 ;
  assign n31982 = n31967 & n31981 ;
  assign n31976 = n19267 & n31968 ;
  assign n31977 = n31967 & n31976 ;
  assign n31978 = ~\core_c_dec_IR_reg[3]/NET0131  & ~n31269 ;
  assign n31979 = \core_c_dec_IR_reg[0]/NET0131  & n31978 ;
  assign n31980 = n31654 & n31979 ;
  assign n31984 = ~n31977 & ~n31980 ;
  assign n31985 = ~n31982 & n31984 ;
  assign n31969 = n19270 & n31968 ;
  assign n31970 = n31967 & n31969 ;
  assign n31971 = ~n4117 & ~n31970 ;
  assign n31972 = ~\core_c_dec_IR_reg[3]/NET0131  & ~n31263 ;
  assign n31973 = n31966 & n31972 ;
  assign n31974 = n19298 & n31968 ;
  assign n31975 = n31967 & n31974 ;
  assign n31983 = ~n31973 & ~n31975 ;
  assign n31986 = n31971 & n31983 ;
  assign n31987 = n31985 & n31986 ;
  assign n31988 = ~n31965 & ~n31987 ;
  assign n31989 = \core_c_dec_Long_Eg_reg/P0001  & n4118 ;
  assign n32000 = ~n31090 & ~n31262 ;
  assign n32001 = ~n30935 & n31083 ;
  assign n32002 = ~n32000 & ~n32001 ;
  assign n32003 = ~n31091 & ~n31268 ;
  assign n32004 = n32002 & ~n32003 ;
  assign n32005 = \core_c_dec_IR_reg[0]/NET0131  & ~n30935 ;
  assign n32006 = \core_c_dec_IR_reg[4]/NET0131  & n30935 ;
  assign n32007 = ~n32005 & ~n32006 ;
  assign n32008 = n32004 & ~n32007 ;
  assign n31990 = \core_c_dec_IR_reg[3]/NET0131  & ~n30935 ;
  assign n31991 = \core_c_dec_IR_reg[7]/NET0131  & n30935 ;
  assign n31992 = ~n31990 & ~n31991 ;
  assign n31993 = \core_c_dec_IR_reg[2]/NET0131  & ~n30935 ;
  assign n31994 = \core_c_dec_IR_reg[6]/NET0131  & n30935 ;
  assign n31995 = ~n31993 & ~n31994 ;
  assign n31996 = \core_c_dec_IR_reg[1]/NET0131  & ~n30935 ;
  assign n31997 = \core_c_dec_IR_reg[5]/NET0131  & n30935 ;
  assign n31998 = ~n31996 & ~n31997 ;
  assign n31999 = ~n31995 & ~n31998 ;
  assign n32009 = ~n31992 & n31999 ;
  assign n32010 = n32008 & n32009 ;
  assign n32023 = \core_c_dec_IR_reg[3]/NET0131  & ~n31269 ;
  assign n32024 = \core_c_dec_IR_reg[0]/NET0131  & n32023 ;
  assign n32025 = n31654 & n32024 ;
  assign n32011 = ~\core_c_dec_IR_reg[13]/NET0131  & ~\core_c_dec_IR_reg[5]/NET0131  ;
  assign n32012 = ~\core_c_dec_IR_reg[7]/NET0131  & n32011 ;
  assign n32013 = n24815 & ~n32012 ;
  assign n32026 = ~n21250 & ~n25249 ;
  assign n32027 = ~n32013 & n32026 ;
  assign n32028 = ~n32025 & n32027 ;
  assign n32029 = ~n32010 & n32028 ;
  assign n32021 = n31992 & n31995 ;
  assign n32022 = n32008 & n32021 ;
  assign n32014 = n31995 & n31998 ;
  assign n32015 = n32007 & n32014 ;
  assign n32016 = n31992 & n32004 ;
  assign n32017 = n32015 & n32016 ;
  assign n32018 = ~n31992 & n32002 ;
  assign n32019 = n32003 & n32018 ;
  assign n32020 = n31999 & n32019 ;
  assign n32030 = ~n32017 & ~n32020 ;
  assign n32031 = ~n32022 & n32030 ;
  assign n32032 = n32029 & n32031 ;
  assign n32033 = n23231 & ~n32032 ;
  assign n32034 = ~n31989 & ~n32033 ;
  assign n32035 = \sice_ICYC_reg[23]/NET0131  & n20785 ;
  assign n32036 = ~\core_c_psq_PCS_reg[3]/NET0131  & ~n32035 ;
  assign n32037 = ~\core_c_dec_Dummy_E_reg/NET0131  & ~n4093 ;
  assign n32038 = n32036 & n32037 ;
  assign n32039 = n22584 & n32038 ;
  assign n32040 = \sice_IIRC_reg[18]/NET0131  & n32039 ;
  assign n32041 = \sice_IIRC_reg[19]/NET0131  & n32040 ;
  assign n32042 = \sice_IIRC_reg[20]/NET0131  & n32041 ;
  assign n32043 = ~\sice_IIRC_reg[20]/NET0131  & ~n32041 ;
  assign n32044 = ~n32042 & ~n32043 ;
  assign n32045 = n6111 & ~n6164 ;
  assign n32046 = ~n6121 & n32045 ;
  assign n32047 = ~n6047 & n32046 ;
  assign n32048 = ~n6112 & ~n32047 ;
  assign n32055 = n7622 & ~n32048 ;
  assign n32049 = n6546 & n32048 ;
  assign n32050 = ~n6101 & n6121 ;
  assign n32051 = ~n6111 & ~n32050 ;
  assign n32052 = ~n6047 & n6165 ;
  assign n32053 = n6111 & ~n32052 ;
  assign n32054 = ~n32051 & ~n32053 ;
  assign n32056 = ~n32049 & n32054 ;
  assign n32057 = ~n32055 & n32056 ;
  assign n32062 = n9497 & ~n32048 ;
  assign n32058 = n6047 & ~n6121 ;
  assign n32059 = ~n9452 & n32058 ;
  assign n32060 = ~n9445 & n32048 ;
  assign n32061 = ~n32059 & n32060 ;
  assign n32063 = ~n32054 & ~n32061 ;
  assign n32064 = ~n32062 & n32063 ;
  assign n32065 = ~n32057 & ~n32064 ;
  assign n32066 = ~n6106 & ~n6111 ;
  assign n32067 = ~n6101 & n32066 ;
  assign n32068 = ~n32053 & ~n32067 ;
  assign n32069 = ~n32065 & ~n32068 ;
  assign n32071 = ~n7340 & n32048 ;
  assign n32070 = ~n7607 & ~n32048 ;
  assign n32072 = n32054 & ~n32070 ;
  assign n32073 = ~n32071 & n32072 ;
  assign n32075 = n6951 & ~n32048 ;
  assign n32074 = n6158 & n32048 ;
  assign n32076 = ~n32054 & ~n32074 ;
  assign n32077 = ~n32075 & n32076 ;
  assign n32078 = ~n32073 & ~n32077 ;
  assign n32079 = n32068 & ~n32078 ;
  assign n32080 = ~n32069 & ~n32079 ;
  assign n32081 = \core_c_psq_DMOVL_reg_DO_reg[3]/NET0131  & ~n25009 ;
  assign n32082 = n32080 & n32081 ;
  assign n32083 = ~PM_bdry_sel_pad & n20698 ;
  assign n32084 = \core_c_psq_PMOVL_regh_DO_reg[3]/NET0131  & ~n19702 ;
  assign n32085 = ~n20687 & n32084 ;
  assign n32086 = ~n32083 & n32085 ;
  assign n32087 = ~n25081 & ~n32086 ;
  assign n32088 = ~n32082 & n32087 ;
  assign n32089 = n11741 & ~n32088 ;
  assign n32090 = ~\T_TMODE[1]_pad  & ~n4117 ;
  assign n32091 = ~n32089 & n32090 ;
  assign n32092 = n4068 & n4117 ;
  assign n32093 = ~n32091 & ~n32092 ;
  assign n32094 = n10638 & n31339 ;
  assign n32096 = \core_dag_ilm2reg_M6_we_DO_reg[8]/NET0131  & n31331 ;
  assign n32098 = \core_dag_ilm2reg_M7_we_DO_reg[8]/NET0131  & n31337 ;
  assign n32099 = ~n32096 & ~n32098 ;
  assign n32100 = ~n21579 & n32099 ;
  assign n32095 = \core_dag_ilm2reg_M5_we_DO_reg[8]/NET0131  & n31341 ;
  assign n32097 = \core_dag_ilm2reg_M4_we_DO_reg[8]/NET0131  & n31344 ;
  assign n32101 = ~n32095 & ~n32097 ;
  assign n32102 = n32100 & n32101 ;
  assign n32103 = ~n32094 & n32102 ;
  assign n32104 = ~\core_dag_ilm2reg_M_reg[8]/NET0131  & n21579 ;
  assign n32105 = ~n32103 & ~n32104 ;
  assign n32106 = n7340 & n31339 ;
  assign n32108 = \core_dag_ilm2reg_M7_we_DO_reg[13]/NET0131  & n31337 ;
  assign n32110 = \core_dag_ilm2reg_M6_we_DO_reg[13]/NET0131  & n31331 ;
  assign n32111 = ~n32108 & ~n32110 ;
  assign n32112 = ~n21579 & n32111 ;
  assign n32107 = \core_dag_ilm2reg_M4_we_DO_reg[13]/NET0131  & n31344 ;
  assign n32109 = \core_dag_ilm2reg_M5_we_DO_reg[13]/NET0131  & n31341 ;
  assign n32113 = ~n32107 & ~n32109 ;
  assign n32114 = n32112 & n32113 ;
  assign n32115 = ~n32106 & n32114 ;
  assign n32116 = ~\core_dag_ilm2reg_M_reg[13]/NET0131  & n21579 ;
  assign n32117 = ~n32115 & ~n32116 ;
  assign n32118 = n9178 & n31409 ;
  assign n32120 = \core_dag_ilm1reg_M3_we_DO_reg[12]/NET0131  & n31407 ;
  assign n32122 = \core_dag_ilm1reg_M2_we_DO_reg[12]/NET0131  & n31401 ;
  assign n32123 = ~n32120 & ~n32122 ;
  assign n32124 = ~n21592 & n32123 ;
  assign n32119 = \core_dag_ilm1reg_M1_we_DO_reg[12]/NET0131  & n31414 ;
  assign n32121 = \core_dag_ilm1reg_M0_we_DO_reg[12]/NET0131  & n31411 ;
  assign n32125 = ~n32119 & ~n32121 ;
  assign n32126 = n32124 & n32125 ;
  assign n32127 = ~n32118 & n32126 ;
  assign n32128 = ~\core_dag_ilm1reg_M_reg[12]/NET0131  & n21592 ;
  assign n32129 = ~n32127 & ~n32128 ;
  assign n32130 = n11265 & n31339 ;
  assign n32132 = \core_dag_ilm2reg_M7_we_DO_reg[7]/NET0131  & n31337 ;
  assign n32134 = \core_dag_ilm2reg_M6_we_DO_reg[7]/NET0131  & n31331 ;
  assign n32135 = ~n32132 & ~n32134 ;
  assign n32136 = ~n21579 & n32135 ;
  assign n32131 = \core_dag_ilm2reg_M4_we_DO_reg[7]/NET0131  & n31344 ;
  assign n32133 = \core_dag_ilm2reg_M5_we_DO_reg[7]/NET0131  & n31341 ;
  assign n32137 = ~n32131 & ~n32133 ;
  assign n32138 = n32136 & n32137 ;
  assign n32139 = ~n32130 & n32138 ;
  assign n32140 = ~\core_dag_ilm2reg_M_reg[7]/NET0131  & n21579 ;
  assign n32141 = ~n32139 & ~n32140 ;
  assign n32142 = n7607 & n31339 ;
  assign n32144 = \core_dag_ilm2reg_M7_we_DO_reg[0]/NET0131  & n31337 ;
  assign n32146 = \core_dag_ilm2reg_M6_we_DO_reg[0]/NET0131  & n31331 ;
  assign n32147 = ~n32144 & ~n32146 ;
  assign n32148 = ~n21579 & n32147 ;
  assign n32143 = \core_dag_ilm2reg_M4_we_DO_reg[0]/NET0131  & n31344 ;
  assign n32145 = \core_dag_ilm2reg_M5_we_DO_reg[0]/NET0131  & n31341 ;
  assign n32149 = ~n32143 & ~n32145 ;
  assign n32150 = n32148 & n32149 ;
  assign n32151 = ~n32142 & n32150 ;
  assign n32152 = ~\core_dag_ilm2reg_M_reg[0]/NET0131  & n21579 ;
  assign n32153 = ~n32151 & ~n32152 ;
  assign n32154 = n11265 & n31409 ;
  assign n32156 = \core_dag_ilm1reg_M3_we_DO_reg[7]/NET0131  & n31407 ;
  assign n32158 = \core_dag_ilm1reg_M2_we_DO_reg[7]/NET0131  & n31401 ;
  assign n32159 = ~n32156 & ~n32158 ;
  assign n32160 = ~n21592 & n32159 ;
  assign n32155 = \core_dag_ilm1reg_M1_we_DO_reg[7]/NET0131  & n31414 ;
  assign n32157 = \core_dag_ilm1reg_M0_we_DO_reg[7]/NET0131  & n31411 ;
  assign n32161 = ~n32155 & ~n32157 ;
  assign n32162 = n32160 & n32161 ;
  assign n32163 = ~n32154 & n32162 ;
  assign n32164 = ~\core_dag_ilm1reg_M_reg[7]/NET0131  & n21592 ;
  assign n32165 = ~n32163 & ~n32164 ;
  assign n32166 = n8113 & n31409 ;
  assign n32168 = \core_dag_ilm1reg_M2_we_DO_reg[3]/NET0131  & n31401 ;
  assign n32170 = \core_dag_ilm1reg_M3_we_DO_reg[3]/NET0131  & n31407 ;
  assign n32171 = ~n32168 & ~n32170 ;
  assign n32172 = ~n21592 & n32171 ;
  assign n32167 = \core_dag_ilm1reg_M0_we_DO_reg[3]/NET0131  & n31411 ;
  assign n32169 = \core_dag_ilm1reg_M1_we_DO_reg[3]/NET0131  & n31414 ;
  assign n32173 = ~n32167 & ~n32169 ;
  assign n32174 = n32172 & n32173 ;
  assign n32175 = ~n32166 & n32174 ;
  assign n32176 = ~\core_dag_ilm1reg_M_reg[3]/NET0131  & n21592 ;
  assign n32177 = ~n32175 & ~n32176 ;
  assign n32178 = \sport1_regs_FSDIVreg_DO_reg[4]/NET0131  & n28786 ;
  assign n32179 = ~\sport1_cfg_FSi_cnt_reg[4]/NET0131  & ~n28859 ;
  assign n32180 = ~n28860 & ~n32179 ;
  assign n32181 = n28855 & n32180 ;
  assign n32182 = ~n32178 & ~n32181 ;
  assign n32183 = \sport0_regs_FSDIVreg_DO_reg[4]/NET0131  & n28876 ;
  assign n32184 = ~\sport0_cfg_FSi_cnt_reg[4]/NET0131  & ~n28949 ;
  assign n32185 = ~n28950 & ~n32184 ;
  assign n32186 = n28945 & n32185 ;
  assign n32187 = ~n32183 & ~n32186 ;
  assign n32188 = \sport1_regs_FSDIVreg_DO_reg[6]/NET0131  & n28786 ;
  assign n32189 = ~\sport1_cfg_FSi_cnt_reg[6]/NET0131  & ~n28861 ;
  assign n32190 = ~n28862 & ~n32189 ;
  assign n32191 = n28855 & n32190 ;
  assign n32192 = ~n32188 & ~n32191 ;
  assign n32193 = \sport0_regs_FSDIVreg_DO_reg[6]/NET0131  & n28876 ;
  assign n32194 = ~\sport0_cfg_FSi_cnt_reg[6]/NET0131  & ~n28951 ;
  assign n32195 = ~n28952 & ~n32194 ;
  assign n32196 = n28945 & n32195 ;
  assign n32197 = ~n32193 & ~n32196 ;
  assign n32198 = \tm_tsr_reg_DO_reg[1]/NET0131  & ~n25491 ;
  assign n32199 = ~\tm_TSR_TMP_reg[1]/NET0131  & n31935 ;
  assign n32200 = \tm_TSR_TMP_reg[1]/NET0131  & ~n31935 ;
  assign n32201 = ~n32199 & ~n32200 ;
  assign n32202 = n25491 & ~n32201 ;
  assign n32203 = ~n32198 & ~n32202 ;
  assign n32204 = \tm_tsr_reg_DO_reg[2]/NET0131  & ~n25491 ;
  assign n32205 = \tm_TSR_TMP_reg[2]/NET0131  & ~n32199 ;
  assign n32206 = n22402 & n31935 ;
  assign n32207 = ~n32205 & ~n32206 ;
  assign n32208 = n25491 & ~n32207 ;
  assign n32209 = ~n32204 & ~n32208 ;
  assign n32210 = \tm_TSR_TMP_reg[3]/NET0131  & ~n32206 ;
  assign n32211 = ~\core_c_psq_PCS_reg[3]/NET0131  & n22404 ;
  assign n32212 = ~n32210 & ~n32211 ;
  assign n32213 = n25491 & ~n32212 ;
  assign n32214 = \tm_tsr_reg_DO_reg[3]/NET0131  & ~n25491 ;
  assign n32215 = ~n32213 & ~n32214 ;
  assign n32216 = ~\sport1_regs_AUTOreg_DO_reg[1]/NET0131  & \sport1_txctl_c_sync1_reg/P0001  ;
  assign n32217 = ~\sport1_txctl_c_sync2_reg/P0001  & n32216 ;
  assign n32218 = \core_dag_modulo1_T1wrap_reg/P0001  & \sport1_regs_AUTOreg_DO_reg[1]/NET0131  ;
  assign n32219 = ~\core_c_psq_IFC_reg[10]/NET0131  & ~n32218 ;
  assign n32220 = ~n32217 & n32219 ;
  assign n32221 = \memc_usysr_DO_reg[11]/NET0131  & ~n32220 ;
  assign n32222 = ~\core_c_psq_Iflag_reg[2]/NET0131  & ~n32221 ;
  assign n32223 = n21406 & ~n32222 ;
  assign n32224 = n19203 & n23586 ;
  assign n32225 = n19202 & ~n32224 ;
  assign n32234 = \core_c_psq_ststk_sts7x23_STcell_reg[2][7]/P0001  & n14713 ;
  assign n32232 = \core_c_psq_ststk_sts7x23_STcell_reg[4][7]/P0001  & n14706 ;
  assign n32233 = \core_c_psq_ststk_sts7x23_STcell_reg[0][7]/P0001  & n14702 ;
  assign n32237 = ~n32232 & ~n32233 ;
  assign n32238 = ~n32234 & n32237 ;
  assign n32228 = \core_c_psq_ststk_sts7x23_STcell_reg[1][7]/P0001  & n14708 ;
  assign n32229 = \core_c_psq_ststk_sts7x23_STcell_reg[5][7]/P0001  & n14699 ;
  assign n32235 = ~n32228 & ~n32229 ;
  assign n32230 = \core_c_psq_ststk_sts7x23_STcell_reg[6][7]/P0001  & n14711 ;
  assign n32231 = \core_c_psq_ststk_sts7x23_STcell_reg[3][7]/P0001  & n14704 ;
  assign n32236 = ~n32230 & ~n32231 ;
  assign n32239 = n32235 & n32236 ;
  assign n32240 = n32238 & n32239 ;
  assign n32241 = n14697 & ~n32240 ;
  assign n32227 = \core_c_dec_MTASTAT_E_reg/P0001  & n11265 ;
  assign n32243 = n17938 & ~n23664 ;
  assign n32242 = ~n17938 & n23664 ;
  assign n32244 = n23586 & ~n32242 ;
  assign n32245 = ~n32243 & n32244 ;
  assign n32246 = n13803 & n32245 ;
  assign n32247 = ~n32227 & ~n32246 ;
  assign n32248 = ~n32241 & n32247 ;
  assign n32249 = ~n32225 & n32248 ;
  assign n32226 = ~\core_eu_ec_cun_SS_reg/P0001  & n32225 ;
  assign n32250 = n4150 & ~n32226 ;
  assign n32251 = ~n32249 & n32250 ;
  assign n32253 = ~n19205 & n19263 ;
  assign n32252 = ~\core_eu_ec_cun_AV_reg/P0001  & n19205 ;
  assign n32254 = n4150 & ~n32252 ;
  assign n32255 = ~n32253 & n32254 ;
  assign n32256 = ~\sport0_cfg_SCLKi_cnt_reg[12]/NET0131  & ~n19549 ;
  assign n32257 = n19197 & ~n19550 ;
  assign n32258 = ~n32256 & n32257 ;
  assign n32259 = ~\sport0_cfg_SCLKi_cnt_reg[10]/NET0131  & ~n19547 ;
  assign n32260 = n19197 & ~n19548 ;
  assign n32261 = ~n32259 & n32260 ;
  assign n32262 = \sport1_rxctl_LMcnt_reg[2]/NET0131  & ~n30751 ;
  assign n32263 = ~n30752 & ~n32262 ;
  assign n32264 = ~n30754 & n31705 ;
  assign n32265 = ~n32263 & n32264 ;
  assign n32266 = \core_c_dec_MTSR1_E_reg/P0001  & n4117 ;
  assign n32267 = n31080 & ~n31102 ;
  assign n32268 = n31120 & n32267 ;
  assign n32269 = ~n32266 & ~n32268 ;
  assign n32270 = n4116 & ~n32269 ;
  assign n32271 = \core_c_dec_MTSR0_E_reg/P0001  & n4117 ;
  assign n32272 = n31127 & n32267 ;
  assign n32273 = ~n32271 & ~n32272 ;
  assign n32274 = n4116 & ~n32273 ;
  assign n32275 = \core_c_dec_MTSI_E_reg/P0001  & n4117 ;
  assign n32276 = n31076 & ~n31102 ;
  assign n32277 = n31079 & n32276 ;
  assign n32278 = n31127 & n32277 ;
  assign n32279 = ~n32275 & ~n32278 ;
  assign n32280 = n4116 & ~n32279 ;
  assign n32281 = \core_c_dec_MTSE_E_reg/P0001  & n4117 ;
  assign n32282 = n31120 & n32277 ;
  assign n32283 = ~n32281 & ~n32282 ;
  assign n32284 = n4116 & ~n32283 ;
  assign n32285 = \core_c_dec_MTMR2_E_reg/P0001  & n4117 ;
  assign n32286 = ~n31079 & n32276 ;
  assign n32287 = n31120 & n32286 ;
  assign n32288 = ~n32285 & ~n32287 ;
  assign n32289 = n4116 & ~n32288 ;
  assign n32290 = \core_c_dec_MTMR1_E_reg/P0001  & n4117 ;
  assign n32291 = n31127 & n32286 ;
  assign n32292 = ~n32290 & ~n32291 ;
  assign n32293 = n4116 & ~n32292 ;
  assign n32294 = \core_c_dec_MTMR0_E_reg/P0001  & n4117 ;
  assign n32295 = ~n31102 & n31545 ;
  assign n32296 = n31120 & n32295 ;
  assign n32297 = ~n32294 & ~n32296 ;
  assign n32298 = n4116 & ~n32297 ;
  assign n32299 = \core_c_dec_MTAR_E_reg/P0001  & n4117 ;
  assign n32300 = n31127 & n32295 ;
  assign n32301 = ~n32299 & ~n32300 ;
  assign n32302 = n4116 & ~n32301 ;
  assign n32303 = \sport1_rxctl_LMcnt_reg[3]/NET0131  & ~n30752 ;
  assign n32304 = ~n30753 & ~n32303 ;
  assign n32305 = n32264 & ~n32304 ;
  assign n32306 = \sport1_rxctl_LMcnt_reg[0]/NET0131  & \sport1_rxctl_LMcnt_reg[1]/NET0131  ;
  assign n32307 = ~n30751 & ~n32306 ;
  assign n32308 = n32264 & ~n32307 ;
  assign n32309 = ~n30778 & n31868 ;
  assign n32310 = \sport0_rxctl_LMcnt_reg[3]/NET0131  & ~n30776 ;
  assign n32311 = ~n30777 & ~n32310 ;
  assign n32312 = n32309 & ~n32311 ;
  assign n32313 = \sport0_rxctl_LMcnt_reg[2]/NET0131  & ~n30775 ;
  assign n32314 = ~n30776 & ~n32313 ;
  assign n32315 = n32309 & ~n32314 ;
  assign n32316 = \sport0_rxctl_LMcnt_reg[0]/NET0131  & \sport0_rxctl_LMcnt_reg[1]/NET0131  ;
  assign n32317 = ~n30775 & ~n32316 ;
  assign n32318 = n32309 & ~n32317 ;
  assign n32319 = ~\sport0_rxctl_LMcnt_reg[0]/NET0131  & n32309 ;
  assign n32320 = \clkc_oscntr_reg_DO_reg[4]/NET0131  & n31917 ;
  assign n32321 = ~\clkc_oscntr_reg_DO_reg[4]/NET0131  & ~\clkc_oscntr_reg_DO_reg[5]/NET0131  ;
  assign n32322 = \T_TMODE[0]_pad  & ~\clkc_oscntr_reg_DO_reg[6]/NET0131  ;
  assign n32323 = n32321 & n32322 ;
  assign n32324 = ~n32320 & ~n32323 ;
  assign n32325 = n23417 & ~n32324 ;
  assign n32326 = \sport0_regs_AUTO_a_reg[15]/NET0131  & ~n32325 ;
  assign n32329 = n20848 & n26045 ;
  assign n32330 = n32321 & n32329 ;
  assign n32327 = ~\clkc_oscntr_reg_DO_reg[8]/NET0131  & ~\clkc_oscntr_reg_DO_reg[9]/NET0131  ;
  assign n32328 = ~\sport0_regs_AUTO_a_reg[15]/NET0131  & n32327 ;
  assign n32331 = n31913 & n32328 ;
  assign n32332 = n32330 & n32331 ;
  assign n32333 = ~n32326 & ~n32332 ;
  assign n32334 = ~\clkc_Cnt128_reg/NET0131  & ~n32333 ;
  assign n32335 = ~\clkc_Awake_reg/NET0131  & ~n32334 ;
  assign n32336 = ~\sport1_cfg_SCLKi_cnt_reg[12]/NET0131  & ~n20250 ;
  assign n32337 = n19130 & ~n20251 ;
  assign n32338 = ~n32336 & n32337 ;
  assign n32339 = ~\sport1_cfg_SCLKi_cnt_reg[10]/NET0131  & ~n20240 ;
  assign n32340 = n19130 & ~n20249 ;
  assign n32341 = ~n32339 & n32340 ;
  assign n32342 = ~\sport1_rxctl_LMcnt_reg[0]/NET0131  & n32264 ;
  assign n32343 = \core_c_dec_MTSR1_E_reg/P0001  & ~n19504 ;
  assign n32344 = ~\core_c_dec_MTSR1_E_reg/P0001  & n29626 ;
  assign n32345 = ~n32343 & ~n32344 ;
  assign n32346 = n18717 & ~n32345 ;
  assign n32347 = ~\core_eu_es_sht_es_reg_sr1swe_DO_reg[9]/P0001  & ~n18717 ;
  assign n32348 = ~n32346 & ~n32347 ;
  assign n32351 = n4064 & n13757 ;
  assign n32350 = \core_c_psq_T_IRQE0_reg/P0001  & ~\core_c_psq_T_IRQE0_s1_reg/P0001  ;
  assign n32352 = ~\core_c_psq_IFC_reg[11]/NET0131  & ~\core_c_psq_Iflag_reg[3]/NET0131  ;
  assign n32353 = ~n32350 & n32352 ;
  assign n32354 = ~n32351 & n32353 ;
  assign n32349 = \core_c_psq_Iact_E_reg[3]/NET0131  & ~n4116 ;
  assign n32355 = ~\core_c_psq_IFC_reg[3]/NET0131  & ~n32349 ;
  assign n32356 = ~n32354 & n32355 ;
  assign n32357 = \core_c_psq_Iact_E_reg[0]/NET0131  & ~n4116 ;
  assign n32358 = ~\T_TMODE[0]_pad  & ~\tm_TINT_GEN1_reg/NET0131  ;
  assign n32359 = \tm_TINT_GEN2_reg/NET0131  & n32358 ;
  assign n32360 = ~\core_c_psq_IFC_reg[8]/NET0131  & ~\core_c_psq_Iflag_reg[0]/NET0131  ;
  assign n32361 = ~n32359 & n32360 ;
  assign n32362 = ~\core_c_psq_IFC_reg[0]/NET0131  & ~n32361 ;
  assign n32363 = ~n32357 & n32362 ;
  assign n32364 = ~\core_c_psq_PCS_reg[3]/NET0131  & ~n4112 ;
  assign n32365 = ~\core_c_dec_MTIMASK_Eg_reg/P0001  & ~n14697 ;
  assign n32366 = ~n5950 & ~n32365 ;
  assign n32367 = ~n32364 & n32366 ;
  assign n32368 = \core_c_dec_MTIMASK_Eg_reg/P0001  & ~n8113 ;
  assign n32372 = \core_c_psq_ststk_sts7x23_STcell_reg[5][18]/P0001  & n14699 ;
  assign n32373 = \core_c_psq_ststk_sts7x23_STcell_reg[3][18]/P0001  & n14704 ;
  assign n32378 = ~n32372 & ~n32373 ;
  assign n32374 = \core_c_psq_ststk_sts7x23_STcell_reg[0][18]/P0001  & n14702 ;
  assign n32375 = \core_c_psq_ststk_sts7x23_STcell_reg[4][18]/P0001  & n14706 ;
  assign n32379 = ~n32374 & ~n32375 ;
  assign n32380 = n32378 & n32379 ;
  assign n32369 = \core_c_psq_ststk_sts7x23_STcell_reg[1][18]/P0001  & n14708 ;
  assign n32376 = ~\core_c_dec_MTIMASK_Eg_reg/P0001  & ~n32369 ;
  assign n32370 = \core_c_psq_ststk_sts7x23_STcell_reg[2][18]/P0001  & n14713 ;
  assign n32371 = \core_c_psq_ststk_sts7x23_STcell_reg[6][18]/P0001  & n14711 ;
  assign n32377 = ~n32370 & ~n32371 ;
  assign n32381 = n32376 & n32377 ;
  assign n32382 = n32380 & n32381 ;
  assign n32383 = ~n32368 & ~n32382 ;
  assign n32384 = n32367 & n32383 ;
  assign n32385 = ~\core_c_psq_Iact_E_reg[2]/NET0131  & n5299 ;
  assign n32386 = \core_c_psq_ICNTL_reg_DO_reg[4]/NET0131  & ~n32385 ;
  assign n32387 = n32364 & ~n32386 ;
  assign n32388 = \core_c_psq_IMASK_reg[3]/NET0131  & ~n32387 ;
  assign n32389 = ~n32367 & n32388 ;
  assign n32390 = ~n32384 & ~n32389 ;
  assign n32391 = n17833 & ~n32345 ;
  assign n32392 = ~\core_eu_es_sht_es_reg_sr1rwe_DO_reg[9]/P0001  & ~n17833 ;
  assign n32393 = ~n32391 & ~n32392 ;
  assign n32401 = ~\sport0_rxctl_ldRX_cmp_reg/P0001  & n12688 ;
  assign n32395 = \sport0_rxctl_RX_reg[0]/P0001  & \sport0_rxctl_RX_reg[2]/P0001  ;
  assign n32396 = n20913 & n32395 ;
  assign n32397 = ~n20888 & n32396 ;
  assign n32398 = n20881 & n32397 ;
  assign n32399 = ~\sport0_rxctl_RX_reg[7]/P0001  & n20875 ;
  assign n32400 = ~n32398 & n32399 ;
  assign n32402 = \sport0_rxctl_RX_reg[14]/P0001  & n20873 ;
  assign n32403 = ~n20868 & ~n32402 ;
  assign n32404 = ~n32400 & n32403 ;
  assign n32405 = ~n32401 & n32404 ;
  assign n32394 = ~\sport0_rxctl_RXSHT_reg[14]/P0001  & n20868 ;
  assign n32406 = ~n20871 & ~n32394 ;
  assign n32407 = ~n32405 & n32406 ;
  assign n32408 = \sport0_rxctl_RX_reg[14]/P0001  & n20871 ;
  assign n32409 = ~n32407 & ~n32408 ;
  assign n32411 = ~\sport0_rxctl_ldRX_cmp_reg/P0001  & n12743 ;
  assign n32412 = \sport0_rxctl_RX_reg[15]/P0001  & n20873 ;
  assign n32413 = ~n20868 & ~n32412 ;
  assign n32414 = ~n32400 & n32413 ;
  assign n32415 = ~n32411 & n32414 ;
  assign n32410 = ~\sport0_rxctl_RXSHT_reg[15]/P0001  & n20868 ;
  assign n32416 = ~n20871 & ~n32410 ;
  assign n32417 = ~n32415 & n32416 ;
  assign n32418 = \sport0_rxctl_RX_reg[15]/P0001  & n20871 ;
  assign n32419 = ~n32417 & ~n32418 ;
  assign n32420 = ~n29560 & n31064 ;
  assign n32421 = \core_eu_ea_alu_ea_reg_arswe_DO_reg[9]/P0001  & ~n31064 ;
  assign n32422 = ~n32420 & ~n32421 ;
  assign n32423 = n27915 & ~n28023 ;
  assign n32424 = \core_c_psq_CNTR_reg_DO_reg[9]/NET0131  & ~n27915 ;
  assign n32425 = ~n32423 & ~n32424 ;
  assign n32426 = n27915 & ~n27978 ;
  assign n32427 = \core_c_psq_CNTR_reg_DO_reg[8]/NET0131  & ~n27915 ;
  assign n32428 = ~n32426 & ~n32427 ;
  assign n32429 = n27915 & ~n27993 ;
  assign n32430 = \core_c_psq_CNTR_reg_DO_reg[4]/NET0131  & ~n27915 ;
  assign n32431 = ~n32429 & ~n32430 ;
  assign n32432 = n27915 & ~n28038 ;
  assign n32433 = \core_c_psq_CNTR_reg_DO_reg[3]/NET0131  & ~n27915 ;
  assign n32434 = ~n32432 & ~n32433 ;
  assign n32435 = ~n30397 & n31064 ;
  assign n32436 = \core_eu_ea_alu_ea_reg_arswe_DO_reg[8]/P0001  & ~n31064 ;
  assign n32437 = ~n32435 & ~n32436 ;
  assign n32438 = n27915 & ~n28069 ;
  assign n32439 = \core_c_psq_CNTR_reg_DO_reg[2]/NET0131  & ~n27915 ;
  assign n32440 = ~n32438 & ~n32439 ;
  assign n32441 = n27915 & ~n27948 ;
  assign n32442 = \core_c_psq_CNTR_reg_DO_reg[12]/NET0131  & ~n27915 ;
  assign n32443 = ~n32441 & ~n32442 ;
  assign n32444 = n27915 & ~n28143 ;
  assign n32445 = \core_c_psq_CNTR_reg_DO_reg[11]/NET0131  & ~n27915 ;
  assign n32446 = ~n32444 & ~n32445 ;
  assign n32447 = n27915 & ~n27963 ;
  assign n32448 = \core_c_psq_CNTR_reg_DO_reg[10]/NET0131  & ~n27915 ;
  assign n32449 = ~n32447 & ~n32448 ;
  assign n32450 = ~n30191 & n31064 ;
  assign n32451 = \core_eu_ea_alu_ea_reg_arswe_DO_reg[7]/P0001  & ~n31064 ;
  assign n32452 = ~n32450 & ~n32451 ;
  assign n32453 = ~IACKn_pad & ~\idma_IAL_reg/P0001  ;
  assign n32454 = \memc_MMR_web_reg/NET0131  & n32453 ;
  assign n32455 = ~n20073 & ~n32454 ;
  assign n32456 = ~\idma_IAL_reg/P0001  & ~n10638 ;
  assign n32457 = ~\idma_IADi_reg[8]/P0001  & \idma_IAL_reg/P0001  ;
  assign n32458 = ~n32456 & ~n32457 ;
  assign n32459 = n32455 & n32458 ;
  assign n32460 = ~\idma_DCTL_reg[14]/NET0131  & \idma_PM_1st_reg/NET0131  ;
  assign n32461 = \auctl_DSack_reg/NET0131  & ~n32460 ;
  assign n32462 = n20382 & n32460 ;
  assign n32463 = ~n32461 & ~n32462 ;
  assign n32464 = \idma_WRcyc_reg/NET0131  & ~n32463 ;
  assign n32465 = ~n20394 & ~n32464 ;
  assign n32466 = ~n32454 & ~n32460 ;
  assign n32467 = ~n32465 & n32466 ;
  assign n32468 = \idma_DCTL_reg[0]/NET0131  & n32467 ;
  assign n32469 = \idma_DCTL_reg[1]/NET0131  & n32468 ;
  assign n32470 = \idma_DCTL_reg[2]/NET0131  & n32469 ;
  assign n32471 = \idma_DCTL_reg[3]/NET0131  & n32470 ;
  assign n32472 = \idma_DCTL_reg[4]/NET0131  & n32471 ;
  assign n32473 = \idma_DCTL_reg[5]/NET0131  & n32472 ;
  assign n32474 = \idma_DCTL_reg[6]/NET0131  & n32473 ;
  assign n32475 = \idma_DCTL_reg[7]/NET0131  & n32474 ;
  assign n32477 = \idma_DCTL_reg[8]/NET0131  & n32475 ;
  assign n32476 = ~\idma_DCTL_reg[8]/NET0131  & ~n32475 ;
  assign n32478 = ~n32455 & ~n32476 ;
  assign n32479 = ~n32477 & n32478 ;
  assign n32480 = ~n32459 & ~n32479 ;
  assign n32481 = ~\idma_IAL_reg/P0001  & ~n10289 ;
  assign n32482 = ~\idma_IADi_reg[9]/P0001  & \idma_IAL_reg/P0001  ;
  assign n32483 = ~n32481 & ~n32482 ;
  assign n32484 = n32455 & n32483 ;
  assign n32486 = \idma_DCTL_reg[9]/NET0131  & n32477 ;
  assign n32485 = ~\idma_DCTL_reg[9]/NET0131  & ~n32477 ;
  assign n32487 = ~n32455 & ~n32485 ;
  assign n32488 = ~n32486 & n32487 ;
  assign n32489 = ~n32484 & ~n32488 ;
  assign n32491 = ~\idma_IAL_reg/P0001  & ~n7340 ;
  assign n32490 = ~\idma_IADi_reg[13]/P0001  & \idma_IAL_reg/P0001  ;
  assign n32492 = n32455 & ~n32490 ;
  assign n32493 = ~n32491 & n32492 ;
  assign n32494 = \idma_DCTL_reg[10]/NET0131  & n32486 ;
  assign n32495 = \idma_DCTL_reg[11]/NET0131  & n32494 ;
  assign n32496 = \idma_DCTL_reg[12]/NET0131  & n32495 ;
  assign n32498 = \idma_DCTL_reg[13]/NET0131  & n32496 ;
  assign n32497 = ~\idma_DCTL_reg[13]/NET0131  & ~n32496 ;
  assign n32499 = ~n32455 & ~n32497 ;
  assign n32500 = ~n32498 & n32499 ;
  assign n32501 = ~n32493 & ~n32500 ;
  assign n32502 = ~\idma_DCTL_reg[12]/NET0131  & ~n32495 ;
  assign n32503 = ~n32496 & ~n32502 ;
  assign n32504 = ~n32455 & ~n32503 ;
  assign n32505 = ~\idma_IAL_reg/P0001  & n9178 ;
  assign n32506 = \idma_IADi_reg[12]/P0001  & \idma_IAL_reg/P0001  ;
  assign n32507 = n32455 & ~n32506 ;
  assign n32508 = ~n32505 & n32507 ;
  assign n32509 = ~n32504 & ~n32508 ;
  assign n32510 = ~\idma_IAL_reg/P0001  & ~n8460 ;
  assign n32511 = ~\idma_IADi_reg[11]/P0001  & \idma_IAL_reg/P0001  ;
  assign n32512 = ~n32510 & ~n32511 ;
  assign n32513 = n32455 & n32512 ;
  assign n32514 = ~\idma_DCTL_reg[11]/NET0131  & ~n32494 ;
  assign n32515 = ~n32455 & ~n32495 ;
  assign n32516 = ~n32514 & n32515 ;
  assign n32517 = ~n32513 & ~n32516 ;
  assign n32518 = ~\idma_IAL_reg/P0001  & ~n7859 ;
  assign n32519 = ~\idma_IADi_reg[10]/P0001  & \idma_IAL_reg/P0001  ;
  assign n32520 = ~n32518 & ~n32519 ;
  assign n32521 = n32455 & n32520 ;
  assign n32522 = ~\idma_DCTL_reg[10]/NET0131  & ~n32486 ;
  assign n32523 = ~n32455 & ~n32494 ;
  assign n32524 = ~n32522 & n32523 ;
  assign n32525 = ~n32521 & ~n32524 ;
  assign n32526 = ~n28990 & n31064 ;
  assign n32527 = \core_eu_ea_alu_ea_reg_arswe_DO_reg[6]/P0001  & ~n31064 ;
  assign n32528 = ~n32526 & ~n32527 ;
  assign n32530 = ~\sport0_rxctl_ldRX_cmp_reg/P0001  & n7340 ;
  assign n32531 = \sport0_rxctl_RX_reg[13]/P0001  & n20873 ;
  assign n32532 = ~n20868 & ~n32531 ;
  assign n32533 = ~n32400 & n32532 ;
  assign n32534 = ~n32530 & n32533 ;
  assign n32529 = ~\sport0_rxctl_RXSHT_reg[13]/P0001  & n20868 ;
  assign n32535 = ~n20871 & ~n32529 ;
  assign n32536 = ~n32534 & n32535 ;
  assign n32537 = \sport0_rxctl_RX_reg[13]/P0001  & n20871 ;
  assign n32538 = ~n32536 & ~n32537 ;
  assign n32539 = ~\idma_IAL_reg/P0001  & ~n11265 ;
  assign n32540 = ~\idma_IADi_reg[7]/P0001  & \idma_IAL_reg/P0001  ;
  assign n32541 = ~n32539 & ~n32540 ;
  assign n32542 = n32455 & n32541 ;
  assign n32543 = ~\idma_DCTL_reg[7]/NET0131  & ~n32474 ;
  assign n32544 = ~n32455 & ~n32475 ;
  assign n32545 = ~n32543 & n32544 ;
  assign n32546 = ~n32542 & ~n32545 ;
  assign n32547 = ~\idma_IAL_reg/P0001  & ~n10911 ;
  assign n32548 = ~\idma_IADi_reg[5]/P0001  & \idma_IAL_reg/P0001  ;
  assign n32549 = ~n32547 & ~n32548 ;
  assign n32550 = n32455 & n32549 ;
  assign n32551 = ~\idma_DCTL_reg[5]/NET0131  & ~n32472 ;
  assign n32552 = ~n32473 & ~n32551 ;
  assign n32553 = ~n32455 & n32552 ;
  assign n32554 = ~n32550 & ~n32553 ;
  assign n32555 = ~\idma_IAL_reg/P0001  & ~n11525 ;
  assign n32556 = ~\idma_IADi_reg[6]/P0001  & \idma_IAL_reg/P0001  ;
  assign n32557 = ~n32555 & ~n32556 ;
  assign n32558 = n32455 & n32557 ;
  assign n32559 = ~\idma_DCTL_reg[6]/NET0131  & ~n32473 ;
  assign n32560 = ~n32455 & ~n32474 ;
  assign n32561 = ~n32559 & n32560 ;
  assign n32562 = ~n32558 & ~n32561 ;
  assign n32563 = ~\idma_IAL_reg/P0001  & ~n10069 ;
  assign n32564 = ~\idma_IADi_reg[4]/P0001  & \idma_IAL_reg/P0001  ;
  assign n32565 = ~n32563 & ~n32564 ;
  assign n32566 = n32455 & n32565 ;
  assign n32567 = ~\idma_DCTL_reg[4]/NET0131  & ~n32471 ;
  assign n32568 = ~n32472 & ~n32567 ;
  assign n32569 = ~n32455 & n32568 ;
  assign n32570 = ~n32566 & ~n32569 ;
  assign n32571 = ~\idma_IAL_reg/P0001  & ~n8113 ;
  assign n32572 = ~\idma_IADi_reg[3]/P0001  & \idma_IAL_reg/P0001  ;
  assign n32573 = ~n32571 & ~n32572 ;
  assign n32574 = n32455 & n32573 ;
  assign n32575 = ~\idma_DCTL_reg[3]/NET0131  & ~n32470 ;
  assign n32576 = ~n32471 & ~n32575 ;
  assign n32577 = ~n32455 & n32576 ;
  assign n32578 = ~n32574 & ~n32577 ;
  assign n32579 = ~\idma_IAL_reg/P0001  & ~n8715 ;
  assign n32580 = ~\idma_IADi_reg[2]/P0001  & \idma_IAL_reg/P0001  ;
  assign n32581 = ~n32579 & ~n32580 ;
  assign n32582 = n32455 & n32581 ;
  assign n32583 = ~\idma_DCTL_reg[2]/NET0131  & ~n32469 ;
  assign n32584 = ~n32470 & ~n32583 ;
  assign n32585 = ~n32455 & n32584 ;
  assign n32586 = ~n32582 & ~n32585 ;
  assign n32587 = ~\idma_IAL_reg/P0001  & ~n7607 ;
  assign n32588 = ~\idma_IADi_reg[0]/P0001  & \idma_IAL_reg/P0001  ;
  assign n32589 = ~n32587 & ~n32588 ;
  assign n32590 = n32455 & n32589 ;
  assign n32591 = ~\idma_DCTL_reg[0]/NET0131  & ~n32467 ;
  assign n32592 = ~n32468 & ~n32591 ;
  assign n32593 = ~n32455 & n32592 ;
  assign n32594 = ~n32590 & ~n32593 ;
  assign n32595 = ~n29042 & n31064 ;
  assign n32596 = \core_eu_ea_alu_ea_reg_arswe_DO_reg[5]/P0001  & ~n31064 ;
  assign n32597 = ~n32595 & ~n32596 ;
  assign n32598 = n27915 & ~n28098 ;
  assign n32599 = \core_c_psq_CNTR_reg_DO_reg[7]/NET0131  & ~n27915 ;
  assign n32600 = ~n32598 & ~n32599 ;
  assign n32601 = n27915 & ~n28113 ;
  assign n32602 = \core_c_psq_CNTR_reg_DO_reg[6]/NET0131  & ~n27915 ;
  assign n32603 = ~n32601 & ~n32602 ;
  assign n32604 = \core_c_psq_CNTR_reg_DO_reg[0]/NET0131  & ~n27915 ;
  assign n32605 = ~n28083 & ~n32604 ;
  assign n32606 = n31697 & n31703 ;
  assign n32607 = ~\sport1_rxctl_Wcnt_reg[0]/NET0131  & ~\sport1_rxctl_Wcnt_reg[1]/NET0131  ;
  assign n32608 = ~\sport1_rxctl_Wcnt_reg[2]/NET0131  & ~\sport1_rxctl_Wcnt_reg[3]/NET0131  ;
  assign n32609 = n32607 & n32608 ;
  assign n32610 = n20408 & n32609 ;
  assign n32611 = n32606 & n32610 ;
  assign n32612 = ~n31702 & ~n32611 ;
  assign n32613 = n32606 & ~n32610 ;
  assign n32614 = n32607 & n32613 ;
  assign n32615 = ~\sport1_rxctl_Wcnt_reg[2]/NET0131  & n32614 ;
  assign n32616 = ~\sport1_rxctl_Wcnt_reg[3]/NET0131  & n32615 ;
  assign n32617 = \sport1_rxctl_Wcnt_reg[4]/NET0131  & ~n32616 ;
  assign n32618 = ~\sport1_rxctl_Wcnt_reg[4]/NET0131  & n32616 ;
  assign n32619 = ~n32617 & ~n32618 ;
  assign n32620 = n32612 & ~n32619 ;
  assign n32621 = \sport1_regs_MWORDreg_DO_reg[4]/NET0131  & ~n32612 ;
  assign n32622 = ~n32620 & ~n32621 ;
  assign n32623 = n27915 & ~n28128 ;
  assign n32624 = \core_c_psq_CNTR_reg_DO_reg[5]/NET0131  & ~n27915 ;
  assign n32625 = ~n32623 & ~n32624 ;
  assign n32626 = n27915 & ~n28008 ;
  assign n32627 = \core_c_psq_CNTR_reg_DO_reg[1]/NET0131  & ~n27915 ;
  assign n32628 = ~n32626 & ~n32627 ;
  assign n32629 = ~n29132 & n31064 ;
  assign n32630 = \core_eu_ea_alu_ea_reg_arswe_DO_reg[4]/P0001  & ~n31064 ;
  assign n32631 = ~n32629 & ~n32630 ;
  assign n32632 = \core_c_dec_MFMY1_E_reg/P0001  & n4117 ;
  assign n32633 = ~n4117 & n30972 ;
  assign n32634 = ~n32632 & ~n32633 ;
  assign n32635 = \core_c_dec_MFMY0_E_reg/P0001  & n4117 ;
  assign n32636 = ~n4117 & n30976 ;
  assign n32637 = ~n32635 & ~n32636 ;
  assign n32638 = \core_c_dec_MFMX0_E_reg/P0001  & n4117 ;
  assign n32639 = ~n4117 & n30975 ;
  assign n32640 = n30962 & n32639 ;
  assign n32641 = ~n32638 & ~n32640 ;
  assign n32642 = \core_c_dec_MFAY1_E_reg/P0001  & n4117 ;
  assign n32643 = ~n4117 & n30971 ;
  assign n32644 = n30977 & n32643 ;
  assign n32645 = ~n32642 & ~n32644 ;
  assign n32646 = \core_c_dec_MFAY0_E_reg/P0001  & n4117 ;
  assign n32647 = n30977 & n32639 ;
  assign n32648 = ~n32646 & ~n32647 ;
  assign n32649 = ~n30497 & n31064 ;
  assign n32650 = \core_eu_ea_alu_ea_reg_arswe_DO_reg[3]/P0001  & ~n31064 ;
  assign n32651 = ~n32649 & ~n32650 ;
  assign n32652 = n31857 & n31866 ;
  assign n32653 = ~\sport0_rxctl_Wcnt_reg[0]/NET0131  & ~\sport0_rxctl_Wcnt_reg[1]/NET0131  ;
  assign n32654 = ~\sport0_rxctl_Wcnt_reg[2]/NET0131  & ~\sport0_rxctl_Wcnt_reg[3]/NET0131  ;
  assign n32655 = n32653 & n32654 ;
  assign n32656 = n20430 & n32655 ;
  assign n32657 = n32652 & n32656 ;
  assign n32658 = ~n31862 & ~n32657 ;
  assign n32659 = n32652 & ~n32656 ;
  assign n32660 = n32653 & n32659 ;
  assign n32661 = ~\sport0_rxctl_Wcnt_reg[2]/NET0131  & n32660 ;
  assign n32662 = ~\sport0_rxctl_Wcnt_reg[3]/NET0131  & n32661 ;
  assign n32663 = \sport0_rxctl_Wcnt_reg[4]/NET0131  & ~n32662 ;
  assign n32664 = ~\sport0_rxctl_Wcnt_reg[4]/NET0131  & n32662 ;
  assign n32665 = ~n32663 & ~n32664 ;
  assign n32666 = n32658 & ~n32665 ;
  assign n32667 = \sport0_regs_MWORDreg_DO_reg[4]/NET0131  & ~n32658 ;
  assign n32668 = ~n32666 & ~n32667 ;
  assign n32669 = ~n28566 & n31064 ;
  assign n32670 = \core_eu_ea_alu_ea_reg_arswe_DO_reg[2]/P0001  & ~n31064 ;
  assign n32671 = ~n32669 & ~n32670 ;
  assign n32672 = ~n29183 & n31064 ;
  assign n32673 = \core_eu_ea_alu_ea_reg_arswe_DO_reg[1]/P0001  & ~n31064 ;
  assign n32674 = ~n32672 & ~n32673 ;
  assign n32675 = ~\idma_IAL_reg/P0001  & ~n9435 ;
  assign n32676 = ~\idma_IADi_reg[1]/P0001  & \idma_IAL_reg/P0001  ;
  assign n32677 = ~n32675 & ~n32676 ;
  assign n32678 = n32455 & n32677 ;
  assign n32679 = ~\idma_DCTL_reg[1]/NET0131  & ~n32468 ;
  assign n32680 = ~n32469 & ~n32679 ;
  assign n32681 = ~n32455 & n32680 ;
  assign n32682 = ~n32678 & ~n32681 ;
  assign n32683 = ~n30294 & n31064 ;
  assign n32684 = \core_eu_ea_alu_ea_reg_arswe_DO_reg[14]/P0001  & ~n31064 ;
  assign n32685 = ~n32683 & ~n32684 ;
  assign n32686 = ~n29674 & n31064 ;
  assign n32687 = \core_eu_ea_alu_ea_reg_arswe_DO_reg[13]/P0001  & ~n31064 ;
  assign n32688 = ~n32686 & ~n32687 ;
  assign n32689 = ~n30094 & n31064 ;
  assign n32690 = \core_eu_ea_alu_ea_reg_arswe_DO_reg[12]/P0001  & ~n31064 ;
  assign n32691 = ~n32689 & ~n32690 ;
  assign n32692 = ~n29736 & n31064 ;
  assign n32693 = \core_eu_ea_alu_ea_reg_arswe_DO_reg[11]/P0001  & ~n31064 ;
  assign n32694 = ~n32692 & ~n32693 ;
  assign n32695 = ~n29887 & n31064 ;
  assign n32696 = \core_eu_ea_alu_ea_reg_arswe_DO_reg[10]/P0001  & ~n31064 ;
  assign n32697 = ~n32695 & ~n32696 ;
  assign n32698 = ~n30547 & n31064 ;
  assign n32699 = \core_eu_ea_alu_ea_reg_arswe_DO_reg[0]/P0001  & ~n31064 ;
  assign n32700 = ~n32698 & ~n32699 ;
  assign n32701 = ~n29560 & n31134 ;
  assign n32702 = \core_eu_ea_alu_ea_reg_arrwe_DO_reg[9]/P0001  & ~n31134 ;
  assign n32703 = ~n32701 & ~n32702 ;
  assign n32704 = ~n30397 & n31134 ;
  assign n32705 = \core_eu_ea_alu_ea_reg_arrwe_DO_reg[8]/P0001  & ~n31134 ;
  assign n32706 = ~n32704 & ~n32705 ;
  assign n32707 = ~n30191 & n31134 ;
  assign n32708 = \core_eu_ea_alu_ea_reg_arrwe_DO_reg[7]/P0001  & ~n31134 ;
  assign n32709 = ~n32707 & ~n32708 ;
  assign n32710 = ~n28990 & n31134 ;
  assign n32711 = \core_eu_ea_alu_ea_reg_arrwe_DO_reg[6]/P0001  & ~n31134 ;
  assign n32712 = ~n32710 & ~n32711 ;
  assign n32713 = ~n29132 & n31134 ;
  assign n32714 = \core_eu_ea_alu_ea_reg_arrwe_DO_reg[4]/P0001  & ~n31134 ;
  assign n32715 = ~n32713 & ~n32714 ;
  assign n32716 = ~n30497 & n31134 ;
  assign n32717 = \core_eu_ea_alu_ea_reg_arrwe_DO_reg[3]/P0001  & ~n31134 ;
  assign n32718 = ~n32716 & ~n32717 ;
  assign n32719 = ~n29042 & n31134 ;
  assign n32720 = \core_eu_ea_alu_ea_reg_arrwe_DO_reg[5]/P0001  & ~n31134 ;
  assign n32721 = ~n32719 & ~n32720 ;
  assign n32722 = ~\clkc_STDcnt_reg[8]/NET0131  & ~n31528 ;
  assign n32723 = ~n31521 & ~n31529 ;
  assign n32724 = ~n32722 & n32723 ;
  assign n32725 = ~\clkc_STDcnt_reg[6]/NET0131  & ~n31526 ;
  assign n32726 = ~n31521 & ~n31527 ;
  assign n32727 = ~n32725 & n32726 ;
  assign n32728 = ~\sport0_cfg_SCLKi_cnt_reg[8]/NET0131  & ~n19545 ;
  assign n32729 = n19197 & ~n19546 ;
  assign n32730 = ~n32728 & n32729 ;
  assign n32731 = ~n28566 & n31134 ;
  assign n32732 = \core_eu_ea_alu_ea_reg_arrwe_DO_reg[2]/P0001  & ~n31134 ;
  assign n32733 = ~n32731 & ~n32732 ;
  assign n32734 = ~\sport1_cfg_SCLKi_cnt_reg[8]/NET0131  & ~n20237 ;
  assign n32735 = n19130 & ~n20238 ;
  assign n32736 = ~n32734 & n32735 ;
  assign n32737 = ~n29183 & n31134 ;
  assign n32738 = \core_eu_ea_alu_ea_reg_arrwe_DO_reg[1]/P0001  & ~n31134 ;
  assign n32739 = ~n32737 & ~n32738 ;
  assign n32740 = ~n30294 & n31134 ;
  assign n32741 = \core_eu_ea_alu_ea_reg_arrwe_DO_reg[14]/P0001  & ~n31134 ;
  assign n32742 = ~n32740 & ~n32741 ;
  assign n32743 = ~n29674 & n31134 ;
  assign n32744 = \core_eu_ea_alu_ea_reg_arrwe_DO_reg[13]/P0001  & ~n31134 ;
  assign n32745 = ~n32743 & ~n32744 ;
  assign n32746 = ~n30094 & n31134 ;
  assign n32747 = \core_eu_ea_alu_ea_reg_arrwe_DO_reg[12]/P0001  & ~n31134 ;
  assign n32748 = ~n32746 & ~n32747 ;
  assign n32749 = ~n29736 & n31134 ;
  assign n32750 = \core_eu_ea_alu_ea_reg_arrwe_DO_reg[11]/P0001  & ~n31134 ;
  assign n32751 = ~n32749 & ~n32750 ;
  assign n32752 = ~n29887 & n31134 ;
  assign n32753 = \core_eu_ea_alu_ea_reg_arrwe_DO_reg[10]/P0001  & ~n31134 ;
  assign n32754 = ~n32752 & ~n32753 ;
  assign n32755 = ~n30547 & n31134 ;
  assign n32756 = \core_eu_ea_alu_ea_reg_arrwe_DO_reg[0]/P0001  & ~n31134 ;
  assign n32757 = ~n32755 & ~n32756 ;
  assign n32758 = \bdma_BCTL_reg[3]/NET0131  & n13757 ;
  assign n32759 = ~\bdma_BRST_s2_reg/NET0131  & ~\sice_IRST_syn_reg/P0001  ;
  assign n32760 = ~n32758 & n32759 ;
  assign n32807 = n11525 & n32048 ;
  assign n32808 = n11265 & ~n32048 ;
  assign n32809 = n32068 & ~n32808 ;
  assign n32810 = ~n32807 & n32809 ;
  assign n32812 = ~n11280 & n32048 ;
  assign n32811 = ~n10954 & ~n32048 ;
  assign n32813 = ~n32068 & ~n32811 ;
  assign n32814 = ~n32812 & n32813 ;
  assign n32815 = ~n32810 & ~n32814 ;
  assign n32816 = n32054 & ~n32815 ;
  assign n32817 = ~n10930 & ~n32048 ;
  assign n32818 = ~n10967 & n32058 ;
  assign n32819 = ~n10978 & ~n32818 ;
  assign n32820 = n32048 & ~n32819 ;
  assign n32821 = ~n32068 & ~n32820 ;
  assign n32822 = ~n32817 & n32821 ;
  assign n32824 = ~n10994 & n32048 ;
  assign n32823 = ~n11023 & ~n32048 ;
  assign n32825 = n32068 & ~n32823 ;
  assign n32826 = ~n32824 & n32825 ;
  assign n32827 = ~n32822 & ~n32826 ;
  assign n32828 = ~n32054 & ~n32827 ;
  assign n32829 = ~n32816 & ~n32828 ;
  assign n32877 = n10911 & ~n32048 ;
  assign n32876 = n10638 & n32048 ;
  assign n32878 = n32068 & ~n32876 ;
  assign n32879 = ~n32877 & n32878 ;
  assign n32881 = ~n10663 & ~n32048 ;
  assign n32880 = ~n10343 & n32048 ;
  assign n32882 = ~n32068 & ~n32880 ;
  assign n32883 = ~n32881 & n32882 ;
  assign n32884 = ~n32879 & ~n32883 ;
  assign n32885 = n32054 & ~n32884 ;
  assign n32886 = ~n11654 & ~n32048 ;
  assign n32887 = ~n11609 & n32058 ;
  assign n32888 = ~n11620 & ~n32887 ;
  assign n32889 = n32048 & ~n32888 ;
  assign n32890 = ~n32068 & ~n32889 ;
  assign n32891 = ~n32886 & n32890 ;
  assign n32893 = ~n10414 & n32048 ;
  assign n32892 = ~n10384 & ~n32048 ;
  assign n32894 = n32068 & ~n32892 ;
  assign n32895 = ~n32893 & n32894 ;
  assign n32896 = ~n32891 & ~n32895 ;
  assign n32897 = ~n32054 & ~n32896 ;
  assign n32898 = ~n32885 & ~n32897 ;
  assign n32947 = n32829 & n32898 ;
  assign n32900 = n9435 & ~n32048 ;
  assign n32899 = n9178 & n32048 ;
  assign n32901 = n32068 & ~n32899 ;
  assign n32902 = ~n32900 & n32901 ;
  assign n32904 = ~n8962 & n32048 ;
  assign n32903 = ~n8926 & ~n32048 ;
  assign n32905 = ~n32068 & ~n32903 ;
  assign n32906 = ~n32904 & n32905 ;
  assign n32907 = ~n32902 & ~n32906 ;
  assign n32908 = n32054 & ~n32907 ;
  assign n32909 = ~n8945 & ~n32048 ;
  assign n32910 = ~n8845 & n32058 ;
  assign n32911 = ~n8856 & ~n32910 ;
  assign n32912 = n32048 & ~n32911 ;
  assign n32913 = ~n32068 & ~n32912 ;
  assign n32914 = ~n32909 & n32913 ;
  assign n32916 = ~n8873 & n32048 ;
  assign n32915 = ~n8903 & ~n32048 ;
  assign n32917 = n32068 & ~n32915 ;
  assign n32918 = ~n32916 & n32917 ;
  assign n32919 = ~n32914 & ~n32918 ;
  assign n32920 = ~n32054 & ~n32919 ;
  assign n32921 = ~n32908 & ~n32920 ;
  assign n32923 = n8715 & ~n32048 ;
  assign n32922 = n8460 & n32048 ;
  assign n32924 = n32068 & ~n32922 ;
  assign n32925 = ~n32923 & n32924 ;
  assign n32927 = ~n8246 & n32048 ;
  assign n32926 = ~n8794 & ~n32048 ;
  assign n32928 = ~n32068 & ~n32926 ;
  assign n32929 = ~n32927 & n32928 ;
  assign n32930 = ~n32925 & ~n32929 ;
  assign n32931 = n32054 & ~n32930 ;
  assign n32932 = ~n8813 & ~n32048 ;
  assign n32933 = ~n8723 & n32058 ;
  assign n32934 = ~n8819 & ~n32933 ;
  assign n32935 = n32048 & ~n32934 ;
  assign n32936 = ~n32068 & ~n32935 ;
  assign n32937 = ~n32932 & n32936 ;
  assign n32939 = ~n8750 & n32048 ;
  assign n32938 = ~n8773 & ~n32048 ;
  assign n32940 = n32068 & ~n32938 ;
  assign n32941 = ~n32939 & n32940 ;
  assign n32942 = ~n32937 & ~n32941 ;
  assign n32943 = ~n32054 & ~n32942 ;
  assign n32944 = ~n32931 & ~n32943 ;
  assign n32948 = n32921 & n32944 ;
  assign n32949 = n32947 & n32948 ;
  assign n32945 = ~n24649 & ~n32080 ;
  assign n32762 = n10638 & ~n32048 ;
  assign n32761 = n10911 & n32048 ;
  assign n32763 = n32068 & ~n32761 ;
  assign n32764 = ~n32762 & n32763 ;
  assign n32766 = ~n10343 & ~n32048 ;
  assign n32765 = ~n10663 & n32048 ;
  assign n32767 = ~n32068 & ~n32765 ;
  assign n32768 = ~n32766 & n32767 ;
  assign n32769 = ~n32764 & ~n32768 ;
  assign n32770 = n32054 & ~n32769 ;
  assign n32771 = ~n10324 & ~n32048 ;
  assign n32772 = ~n10356 & n32058 ;
  assign n32773 = ~n10367 & ~n32772 ;
  assign n32774 = n32048 & ~n32773 ;
  assign n32775 = ~n32068 & ~n32774 ;
  assign n32776 = ~n32771 & n32775 ;
  assign n32778 = ~n10384 & n32048 ;
  assign n32777 = ~n10414 & ~n32048 ;
  assign n32779 = n32068 & ~n32777 ;
  assign n32780 = ~n32778 & n32779 ;
  assign n32781 = ~n32776 & ~n32780 ;
  assign n32782 = ~n32054 & ~n32781 ;
  assign n32783 = ~n32770 & ~n32782 ;
  assign n32785 = n11525 & ~n32048 ;
  assign n32784 = n11265 & n32048 ;
  assign n32786 = n32068 & ~n32784 ;
  assign n32787 = ~n32785 & n32786 ;
  assign n32789 = ~n11280 & ~n32048 ;
  assign n32788 = ~n10954 & n32048 ;
  assign n32790 = ~n32068 & ~n32788 ;
  assign n32791 = ~n32789 & n32790 ;
  assign n32792 = ~n32787 & ~n32791 ;
  assign n32793 = n32054 & ~n32792 ;
  assign n32794 = ~n11579 & ~n32048 ;
  assign n32795 = ~n11540 & n32058 ;
  assign n32796 = ~n11551 & ~n32795 ;
  assign n32797 = n32048 & ~n32796 ;
  assign n32798 = ~n32068 & ~n32797 ;
  assign n32799 = ~n32794 & n32798 ;
  assign n32801 = ~n11023 & n32048 ;
  assign n32800 = ~n10994 & ~n32048 ;
  assign n32802 = n32068 & ~n32800 ;
  assign n32803 = ~n32801 & n32802 ;
  assign n32804 = ~n32799 & ~n32803 ;
  assign n32805 = ~n32054 & ~n32804 ;
  assign n32806 = ~n32793 & ~n32805 ;
  assign n32946 = n32783 & n32806 ;
  assign n32950 = n32945 & n32946 ;
  assign n32831 = n10069 & ~n32048 ;
  assign n32830 = n10289 & n32048 ;
  assign n32832 = n32068 & ~n32830 ;
  assign n32833 = ~n32831 & n32832 ;
  assign n32835 = ~n10302 & ~n32048 ;
  assign n32834 = ~n9752 & n32048 ;
  assign n32836 = ~n32068 & ~n32834 ;
  assign n32837 = ~n32835 & n32836 ;
  assign n32838 = ~n32833 & ~n32837 ;
  assign n32839 = n32054 & ~n32838 ;
  assign n32840 = ~n11720 & ~n32048 ;
  assign n32841 = ~n11668 & n32058 ;
  assign n32842 = ~n11692 & ~n32841 ;
  assign n32843 = n32048 & ~n32842 ;
  assign n32844 = ~n32068 & ~n32843 ;
  assign n32845 = ~n32840 & n32844 ;
  assign n32847 = ~n9733 & n32048 ;
  assign n32846 = ~n9786 & ~n32048 ;
  assign n32848 = n32068 & ~n32846 ;
  assign n32849 = ~n32847 & n32848 ;
  assign n32850 = ~n32845 & ~n32849 ;
  assign n32851 = ~n32054 & ~n32850 ;
  assign n32852 = ~n32839 & ~n32851 ;
  assign n32854 = n8113 & ~n32048 ;
  assign n32853 = n7859 & n32048 ;
  assign n32855 = n32068 & ~n32853 ;
  assign n32856 = ~n32854 & n32855 ;
  assign n32858 = ~n8224 & ~n32048 ;
  assign n32857 = ~n7644 & n32048 ;
  assign n32859 = ~n32068 & ~n32857 ;
  assign n32860 = ~n32858 & n32859 ;
  assign n32861 = ~n32856 & ~n32860 ;
  assign n32862 = n32054 & ~n32861 ;
  assign n32863 = ~n8211 & ~n32048 ;
  assign n32864 = ~n8121 & n32058 ;
  assign n32865 = ~n8162 & ~n32864 ;
  assign n32866 = n32048 & ~n32865 ;
  assign n32867 = ~n32068 & ~n32866 ;
  assign n32868 = ~n32863 & n32867 ;
  assign n32870 = ~n8149 & n32048 ;
  assign n32869 = ~n8190 & ~n32048 ;
  assign n32871 = n32068 & ~n32869 ;
  assign n32872 = ~n32870 & n32871 ;
  assign n32873 = ~n32868 & ~n32872 ;
  assign n32874 = ~n32054 & ~n32873 ;
  assign n32875 = ~n32862 & ~n32874 ;
  assign n32951 = n32852 & n32875 ;
  assign n32952 = n32950 & n32951 ;
  assign n32953 = n32949 & n32952 ;
  assign n32954 = n20386 & ~n32465 ;
  assign n32955 = ~\idma_DCTL_reg[14]/NET0131  & ~n32465 ;
  assign n32956 = \idma_PM_1st_reg/NET0131  & ~n32955 ;
  assign n32957 = ~n32954 & ~n32956 ;
  assign n32958 = n20074 & n32957 ;
  assign n32959 = n4150 & ~n25780 ;
  assign n32960 = \tm_tcr_reg_DO_reg[12]/NET0131  & n20355 ;
  assign n32962 = \tm_TCR_TMP_reg[12]/NET0131  & ~n25839 ;
  assign n32963 = ~n22400 & ~n25840 ;
  assign n32964 = ~n32962 & n32963 ;
  assign n32961 = ~\tm_tpr_reg_DO_reg[12]/NET0131  & n22400 ;
  assign n32965 = ~n20355 & ~n32961 ;
  assign n32966 = ~n32964 & n32965 ;
  assign n32967 = ~n32960 & ~n32966 ;
  assign n32968 = \sport1_rxctl_LMcnt_reg[4]/NET0131  & ~n30753 ;
  assign n32969 = n31705 & ~n32968 ;
  assign n32970 = \sport0_rxctl_LMcnt_reg[4]/NET0131  & ~n30777 ;
  assign n32971 = n31868 & ~n32970 ;
  assign n32972 = n4055 & ~n6033 ;
  assign n32973 = n5692 & n5974 ;
  assign n32974 = ~n32972 & n32973 ;
  assign n32975 = ~\core_dag_ilm2reg_IL_E_reg[1]/P0001  & ~n5692 ;
  assign n32976 = ~n32974 & ~n32975 ;
  assign n32977 = n4055 & ~n6036 ;
  assign n32978 = n5692 & n5989 ;
  assign n32979 = ~n32977 & n32978 ;
  assign n32980 = ~\core_dag_ilm2reg_IL_E_reg[0]/P0001  & ~n5692 ;
  assign n32981 = ~n32979 & ~n32980 ;
  assign n32982 = ~n32976 & n32981 ;
  assign n32983 = n25955 & n32982 ;
  assign n32984 = n32976 & ~n32981 ;
  assign n32985 = n25965 & n32984 ;
  assign n32990 = ~n32983 & ~n32985 ;
  assign n32986 = ~n32976 & ~n32981 ;
  assign n32987 = n25954 & n32986 ;
  assign n32988 = n32976 & n32981 ;
  assign n32989 = n25959 & n32988 ;
  assign n32991 = ~n32987 & ~n32989 ;
  assign n32992 = n32990 & n32991 ;
  assign n32993 = n11265 & ~n32992 ;
  assign n32994 = ~n25965 & n32984 ;
  assign n32995 = \core_dag_ilm2reg_L6_we_DO_reg[7]/NET0131  & n32994 ;
  assign n33002 = ~n21579 & ~n32995 ;
  assign n33000 = ~n25955 & n32982 ;
  assign n33001 = \core_dag_ilm2reg_L5_we_DO_reg[7]/NET0131  & n33000 ;
  assign n32996 = ~n25954 & n32986 ;
  assign n32997 = \core_dag_ilm2reg_L4_we_DO_reg[7]/NET0131  & n32996 ;
  assign n32998 = ~n25959 & n32988 ;
  assign n32999 = \core_dag_ilm2reg_L7_we_DO_reg[7]/NET0131  & n32998 ;
  assign n33003 = ~n32997 & ~n32999 ;
  assign n33004 = ~n33001 & n33003 ;
  assign n33005 = n33002 & n33004 ;
  assign n33006 = ~n32993 & n33005 ;
  assign n33007 = ~\core_dag_ilm2reg_L_reg[7]/NET0131  & n21579 ;
  assign n33008 = ~n33006 & ~n33007 ;
  assign n33009 = n11525 & ~n32992 ;
  assign n33010 = \core_dag_ilm2reg_L6_we_DO_reg[6]/NET0131  & n32994 ;
  assign n33014 = ~n21579 & ~n33010 ;
  assign n33013 = \core_dag_ilm2reg_L5_we_DO_reg[6]/NET0131  & n33000 ;
  assign n33011 = \core_dag_ilm2reg_L4_we_DO_reg[6]/NET0131  & n32996 ;
  assign n33012 = \core_dag_ilm2reg_L7_we_DO_reg[6]/NET0131  & n32998 ;
  assign n33015 = ~n33011 & ~n33012 ;
  assign n33016 = ~n33013 & n33015 ;
  assign n33017 = n33014 & n33016 ;
  assign n33018 = ~n33009 & n33017 ;
  assign n33019 = ~\core_dag_ilm2reg_L_reg[6]/NET0131  & n21579 ;
  assign n33020 = ~n33018 & ~n33019 ;
  assign n33021 = n10069 & ~n32992 ;
  assign n33022 = \core_dag_ilm2reg_L4_we_DO_reg[4]/NET0131  & n32996 ;
  assign n33026 = ~n21579 & ~n33022 ;
  assign n33025 = \core_dag_ilm2reg_L7_we_DO_reg[4]/NET0131  & n32998 ;
  assign n33023 = \core_dag_ilm2reg_L6_we_DO_reg[4]/NET0131  & n32994 ;
  assign n33024 = \core_dag_ilm2reg_L5_we_DO_reg[4]/NET0131  & n33000 ;
  assign n33027 = ~n33023 & ~n33024 ;
  assign n33028 = ~n33025 & n33027 ;
  assign n33029 = n33026 & n33028 ;
  assign n33030 = ~n33021 & n33029 ;
  assign n33031 = ~\core_dag_ilm2reg_L_reg[4]/NET0131  & n21579 ;
  assign n33032 = ~n33030 & ~n33031 ;
  assign n33033 = n8113 & ~n32992 ;
  assign n33034 = \core_dag_ilm2reg_L6_we_DO_reg[3]/NET0131  & n32994 ;
  assign n33038 = ~n21579 & ~n33034 ;
  assign n33037 = \core_dag_ilm2reg_L5_we_DO_reg[3]/NET0131  & n33000 ;
  assign n33035 = \core_dag_ilm2reg_L4_we_DO_reg[3]/NET0131  & n32996 ;
  assign n33036 = \core_dag_ilm2reg_L7_we_DO_reg[3]/NET0131  & n32998 ;
  assign n33039 = ~n33035 & ~n33036 ;
  assign n33040 = ~n33037 & n33039 ;
  assign n33041 = n33038 & n33040 ;
  assign n33042 = ~n33033 & n33041 ;
  assign n33043 = ~\core_dag_ilm2reg_L_reg[3]/NET0131  & n21579 ;
  assign n33044 = ~n33042 & ~n33043 ;
  assign n33045 = n8715 & ~n32992 ;
  assign n33046 = \core_dag_ilm2reg_L6_we_DO_reg[2]/NET0131  & n32994 ;
  assign n33050 = ~n21579 & ~n33046 ;
  assign n33049 = \core_dag_ilm2reg_L5_we_DO_reg[2]/NET0131  & n33000 ;
  assign n33047 = \core_dag_ilm2reg_L4_we_DO_reg[2]/NET0131  & n32996 ;
  assign n33048 = \core_dag_ilm2reg_L7_we_DO_reg[2]/NET0131  & n32998 ;
  assign n33051 = ~n33047 & ~n33048 ;
  assign n33052 = ~n33049 & n33051 ;
  assign n33053 = n33050 & n33052 ;
  assign n33054 = ~n33045 & n33053 ;
  assign n33055 = ~\core_dag_ilm2reg_L_reg[2]/NET0131  & n21579 ;
  assign n33056 = ~n33054 & ~n33055 ;
  assign n33057 = n9435 & ~n32992 ;
  assign n33058 = \core_dag_ilm2reg_L4_we_DO_reg[1]/NET0131  & n32996 ;
  assign n33062 = ~n21579 & ~n33058 ;
  assign n33061 = \core_dag_ilm2reg_L7_we_DO_reg[1]/NET0131  & n32998 ;
  assign n33059 = \core_dag_ilm2reg_L6_we_DO_reg[1]/NET0131  & n32994 ;
  assign n33060 = \core_dag_ilm2reg_L5_we_DO_reg[1]/NET0131  & n33000 ;
  assign n33063 = ~n33059 & ~n33060 ;
  assign n33064 = ~n33061 & n33063 ;
  assign n33065 = n33062 & n33064 ;
  assign n33066 = ~n33057 & n33065 ;
  assign n33067 = ~\core_dag_ilm2reg_L_reg[1]/NET0131  & n21579 ;
  assign n33068 = ~n33066 & ~n33067 ;
  assign n33069 = n7607 & ~n32992 ;
  assign n33070 = \core_dag_ilm2reg_L6_we_DO_reg[0]/NET0131  & n32994 ;
  assign n33074 = ~n21579 & ~n33070 ;
  assign n33073 = \core_dag_ilm2reg_L5_we_DO_reg[0]/NET0131  & n33000 ;
  assign n33071 = \core_dag_ilm2reg_L4_we_DO_reg[0]/NET0131  & n32996 ;
  assign n33072 = \core_dag_ilm2reg_L7_we_DO_reg[0]/NET0131  & n32998 ;
  assign n33075 = ~n33071 & ~n33072 ;
  assign n33076 = ~n33073 & n33075 ;
  assign n33077 = n33074 & n33076 ;
  assign n33078 = ~n33069 & n33077 ;
  assign n33079 = ~\core_dag_ilm2reg_L_reg[0]/NET0131  & n21579 ;
  assign n33080 = ~n33078 & ~n33079 ;
  assign n33081 = ~\core_c_dec_IRE_reg[3]/NET0131  & ~n5692 ;
  assign n33082 = \core_c_dec_IR_reg[3]/NET0131  & n4055 ;
  assign n33083 = n32973 & ~n33082 ;
  assign n33084 = ~n33081 & ~n33083 ;
  assign n33085 = ~\core_c_dec_IRE_reg[2]/NET0131  & ~n5692 ;
  assign n33086 = \core_c_dec_IR_reg[2]/NET0131  & n4055 ;
  assign n33087 = n32978 & ~n33086 ;
  assign n33088 = ~n33085 & ~n33087 ;
  assign n33089 = n33084 & n33088 ;
  assign n33090 = n25976 & n33089 ;
  assign n33091 = ~n33084 & ~n33088 ;
  assign n33092 = n25975 & n33091 ;
  assign n33097 = ~n33090 & ~n33092 ;
  assign n33093 = n33084 & ~n33088 ;
  assign n33094 = n25973 & n33093 ;
  assign n33095 = ~n33084 & n33088 ;
  assign n33096 = n25974 & n33095 ;
  assign n33098 = ~n33094 & ~n33096 ;
  assign n33099 = n33097 & n33098 ;
  assign n33100 = n11265 & ~n33099 ;
  assign n33101 = ~n25976 & n33089 ;
  assign n33102 = \core_dag_ilm1reg_L3_we_DO_reg[7]/NET0131  & n33101 ;
  assign n33103 = ~n25975 & n33091 ;
  assign n33104 = \core_dag_ilm1reg_L0_we_DO_reg[7]/NET0131  & n33103 ;
  assign n33109 = ~n33102 & ~n33104 ;
  assign n33105 = ~n25974 & n33095 ;
  assign n33106 = \core_dag_ilm1reg_L1_we_DO_reg[7]/NET0131  & n33105 ;
  assign n33107 = ~n25973 & n33093 ;
  assign n33108 = \core_dag_ilm1reg_L2_we_DO_reg[7]/NET0131  & n33107 ;
  assign n33110 = ~n33106 & ~n33108 ;
  assign n33111 = n33109 & n33110 ;
  assign n33112 = ~n21592 & n33111 ;
  assign n33113 = ~n33100 & n33112 ;
  assign n33114 = ~\core_dag_ilm1reg_L_reg[7]/NET0131  & n21592 ;
  assign n33115 = ~n33113 & ~n33114 ;
  assign n33116 = n11525 & ~n33099 ;
  assign n33117 = \core_dag_ilm1reg_L1_we_DO_reg[6]/NET0131  & n33105 ;
  assign n33118 = \core_dag_ilm1reg_L2_we_DO_reg[6]/NET0131  & n33107 ;
  assign n33121 = ~n33117 & ~n33118 ;
  assign n33119 = \core_dag_ilm1reg_L3_we_DO_reg[6]/NET0131  & n33101 ;
  assign n33120 = \core_dag_ilm1reg_L0_we_DO_reg[6]/NET0131  & n33103 ;
  assign n33122 = ~n33119 & ~n33120 ;
  assign n33123 = n33121 & n33122 ;
  assign n33124 = ~n21592 & n33123 ;
  assign n33125 = ~n33116 & n33124 ;
  assign n33126 = ~\core_dag_ilm1reg_L_reg[6]/NET0131  & n21592 ;
  assign n33127 = ~n33125 & ~n33126 ;
  assign n33128 = n10911 & ~n33099 ;
  assign n33129 = \core_dag_ilm1reg_L1_we_DO_reg[5]/NET0131  & n33105 ;
  assign n33130 = \core_dag_ilm1reg_L2_we_DO_reg[5]/NET0131  & n33107 ;
  assign n33133 = ~n33129 & ~n33130 ;
  assign n33131 = \core_dag_ilm1reg_L3_we_DO_reg[5]/NET0131  & n33101 ;
  assign n33132 = \core_dag_ilm1reg_L0_we_DO_reg[5]/NET0131  & n33103 ;
  assign n33134 = ~n33131 & ~n33132 ;
  assign n33135 = n33133 & n33134 ;
  assign n33136 = ~n21592 & n33135 ;
  assign n33137 = ~n33128 & n33136 ;
  assign n33138 = ~\core_dag_ilm1reg_L_reg[5]/NET0131  & n21592 ;
  assign n33139 = ~n33137 & ~n33138 ;
  assign n33140 = n10069 & ~n33099 ;
  assign n33141 = \core_dag_ilm1reg_L1_we_DO_reg[4]/NET0131  & n33105 ;
  assign n33142 = \core_dag_ilm1reg_L2_we_DO_reg[4]/NET0131  & n33107 ;
  assign n33145 = ~n33141 & ~n33142 ;
  assign n33143 = \core_dag_ilm1reg_L3_we_DO_reg[4]/NET0131  & n33101 ;
  assign n33144 = \core_dag_ilm1reg_L0_we_DO_reg[4]/NET0131  & n33103 ;
  assign n33146 = ~n33143 & ~n33144 ;
  assign n33147 = n33145 & n33146 ;
  assign n33148 = ~n21592 & n33147 ;
  assign n33149 = ~n33140 & n33148 ;
  assign n33150 = ~\core_dag_ilm1reg_L_reg[4]/NET0131  & n21592 ;
  assign n33151 = ~n33149 & ~n33150 ;
  assign n33152 = n8113 & ~n33099 ;
  assign n33153 = \core_dag_ilm1reg_L1_we_DO_reg[3]/NET0131  & n33105 ;
  assign n33154 = \core_dag_ilm1reg_L2_we_DO_reg[3]/NET0131  & n33107 ;
  assign n33157 = ~n33153 & ~n33154 ;
  assign n33155 = \core_dag_ilm1reg_L3_we_DO_reg[3]/NET0131  & n33101 ;
  assign n33156 = \core_dag_ilm1reg_L0_we_DO_reg[3]/NET0131  & n33103 ;
  assign n33158 = ~n33155 & ~n33156 ;
  assign n33159 = n33157 & n33158 ;
  assign n33160 = ~n21592 & n33159 ;
  assign n33161 = ~n33152 & n33160 ;
  assign n33162 = ~\core_dag_ilm1reg_L_reg[3]/NET0131  & n21592 ;
  assign n33163 = ~n33161 & ~n33162 ;
  assign n33164 = n8715 & ~n33099 ;
  assign n33165 = \core_dag_ilm1reg_L1_we_DO_reg[2]/NET0131  & n33105 ;
  assign n33166 = \core_dag_ilm1reg_L2_we_DO_reg[2]/NET0131  & n33107 ;
  assign n33169 = ~n33165 & ~n33166 ;
  assign n33167 = \core_dag_ilm1reg_L3_we_DO_reg[2]/NET0131  & n33101 ;
  assign n33168 = \core_dag_ilm1reg_L0_we_DO_reg[2]/NET0131  & n33103 ;
  assign n33170 = ~n33167 & ~n33168 ;
  assign n33171 = n33169 & n33170 ;
  assign n33172 = ~n21592 & n33171 ;
  assign n33173 = ~n33164 & n33172 ;
  assign n33174 = ~\core_dag_ilm1reg_L_reg[2]/NET0131  & n21592 ;
  assign n33175 = ~n33173 & ~n33174 ;
  assign n33176 = n9435 & ~n33099 ;
  assign n33177 = \core_dag_ilm1reg_L3_we_DO_reg[1]/NET0131  & n33101 ;
  assign n33178 = \core_dag_ilm1reg_L0_we_DO_reg[1]/NET0131  & n33103 ;
  assign n33181 = ~n33177 & ~n33178 ;
  assign n33179 = \core_dag_ilm1reg_L1_we_DO_reg[1]/NET0131  & n33105 ;
  assign n33180 = \core_dag_ilm1reg_L2_we_DO_reg[1]/NET0131  & n33107 ;
  assign n33182 = ~n33179 & ~n33180 ;
  assign n33183 = n33181 & n33182 ;
  assign n33184 = ~n21592 & n33183 ;
  assign n33185 = ~n33176 & n33184 ;
  assign n33186 = ~\core_dag_ilm1reg_L_reg[1]/NET0131  & n21592 ;
  assign n33187 = ~n33185 & ~n33186 ;
  assign n33188 = n7607 & ~n33099 ;
  assign n33189 = \core_dag_ilm1reg_L1_we_DO_reg[0]/NET0131  & n33105 ;
  assign n33190 = \core_dag_ilm1reg_L2_we_DO_reg[0]/NET0131  & n33107 ;
  assign n33193 = ~n33189 & ~n33190 ;
  assign n33191 = \core_dag_ilm1reg_L3_we_DO_reg[0]/NET0131  & n33101 ;
  assign n33192 = \core_dag_ilm1reg_L0_we_DO_reg[0]/NET0131  & n33103 ;
  assign n33194 = ~n33191 & ~n33192 ;
  assign n33195 = n33193 & n33194 ;
  assign n33196 = ~n21592 & n33195 ;
  assign n33197 = ~n33188 & n33196 ;
  assign n33198 = ~\core_dag_ilm1reg_L_reg[0]/NET0131  & n21592 ;
  assign n33199 = ~n33197 & ~n33198 ;
  assign n33200 = \core_c_psq_TRAP_Eg_reg/NET0131  & ~n19477 ;
  assign n33214 = ~n19480 & ~n19486 ;
  assign n33215 = n19495 & n33214 ;
  assign n33216 = ~n19483 & n33215 ;
  assign n33202 = ~\core_c_psq_Iflag_reg[2]/NET0131  & \memc_usysr_DO_reg[11]/NET0131  ;
  assign n33201 = ~\core_c_psq_Iflag_reg[12]/NET0131  & ~\memc_usysr_DO_reg[11]/NET0131  ;
  assign n33203 = \core_c_psq_IMASK_reg[2]/NET0131  & ~n33201 ;
  assign n33204 = ~n33202 & n33203 ;
  assign n33205 = ~\core_c_psq_PCS_reg[3]/NET0131  & n33204 ;
  assign n33207 = ~\core_c_psq_Iflag_reg[11]/NET0131  & ~\memc_usysr_DO_reg[11]/NET0131  ;
  assign n33206 = ~\core_c_psq_Iflag_reg[1]/NET0131  & \memc_usysr_DO_reg[11]/NET0131  ;
  assign n33208 = \core_c_psq_IMASK_reg[1]/NET0131  & ~\core_c_psq_PCS_reg[3]/NET0131  ;
  assign n33209 = ~n33206 & n33208 ;
  assign n33210 = ~n33207 & n33209 ;
  assign n33211 = ~n33205 & ~n33210 ;
  assign n33212 = \core_c_psq_IMASK_reg[3]/NET0131  & \core_c_psq_Iflag_reg[0]/NET0131  ;
  assign n33213 = ~\core_c_psq_PCS_reg[3]/NET0131  & n33212 ;
  assign n33217 = \core_c_psq_IMASK_reg[0]/NET0131  & \core_c_psq_Iflag_reg[3]/NET0131  ;
  assign n33218 = ~\core_c_psq_PCS_reg[3]/NET0131  & n33217 ;
  assign n33219 = ~n33213 & ~n33218 ;
  assign n33220 = n33211 & n33219 ;
  assign n33221 = n33216 & n33220 ;
  assign n33222 = ~\core_c_psq_PCS_reg[7]/NET0131  & n33221 ;
  assign n33223 = ~n26030 & ~n33222 ;
  assign n33224 = n19477 & n33223 ;
  assign n33225 = n11741 & n33224 ;
  assign n33226 = ~n33200 & ~n33225 ;
  assign n33227 = \core_c_dec_MTIMASK_Eg_reg/P0001  & ~n11525 ;
  assign n33231 = \core_c_psq_ststk_sts7x23_STcell_reg[3][21]/P0001  & n14704 ;
  assign n33232 = \core_c_psq_ststk_sts7x23_STcell_reg[1][21]/P0001  & n14708 ;
  assign n33237 = ~n33231 & ~n33232 ;
  assign n33233 = \core_c_psq_ststk_sts7x23_STcell_reg[2][21]/P0001  & n14713 ;
  assign n33234 = \core_c_psq_ststk_sts7x23_STcell_reg[0][21]/P0001  & n14702 ;
  assign n33238 = ~n33233 & ~n33234 ;
  assign n33239 = n33237 & n33238 ;
  assign n33228 = \core_c_psq_ststk_sts7x23_STcell_reg[6][21]/P0001  & n14711 ;
  assign n33235 = ~\core_c_dec_MTIMASK_Eg_reg/P0001  & ~n33228 ;
  assign n33229 = \core_c_psq_ststk_sts7x23_STcell_reg[4][21]/P0001  & n14706 ;
  assign n33230 = \core_c_psq_ststk_sts7x23_STcell_reg[5][21]/P0001  & n14699 ;
  assign n33236 = ~n33229 & ~n33230 ;
  assign n33240 = n33235 & n33236 ;
  assign n33241 = n33239 & n33240 ;
  assign n33242 = ~n33227 & ~n33241 ;
  assign n33243 = n32367 & n33242 ;
  assign n33244 = ~\core_c_psq_Iact_E_reg[3]/NET0131  & n32385 ;
  assign n33245 = ~\core_c_psq_Iact_E_reg[4]/NET0131  & n33244 ;
  assign n33246 = ~\core_c_psq_Iact_E_reg[5]/NET0131  & n33245 ;
  assign n33247 = \core_c_psq_ICNTL_reg_DO_reg[4]/NET0131  & ~n33246 ;
  assign n33248 = n32364 & ~n33247 ;
  assign n33249 = \core_c_psq_IMASK_reg[6]/NET0131  & ~n33248 ;
  assign n33250 = ~n32367 & n33249 ;
  assign n33251 = ~n33243 & ~n33250 ;
  assign n33252 = \core_c_dec_MTIMASK_Eg_reg/P0001  & ~n10911 ;
  assign n33256 = \core_c_psq_ststk_sts7x23_STcell_reg[3][20]/P0001  & n14704 ;
  assign n33257 = \core_c_psq_ststk_sts7x23_STcell_reg[5][20]/P0001  & n14699 ;
  assign n33262 = ~n33256 & ~n33257 ;
  assign n33258 = \core_c_psq_ststk_sts7x23_STcell_reg[6][20]/P0001  & n14711 ;
  assign n33259 = \core_c_psq_ststk_sts7x23_STcell_reg[0][20]/P0001  & n14702 ;
  assign n33263 = ~n33258 & ~n33259 ;
  assign n33264 = n33262 & n33263 ;
  assign n33253 = \core_c_psq_ststk_sts7x23_STcell_reg[2][20]/P0001  & n14713 ;
  assign n33260 = ~\core_c_dec_MTIMASK_Eg_reg/P0001  & ~n33253 ;
  assign n33254 = \core_c_psq_ststk_sts7x23_STcell_reg[4][20]/P0001  & n14706 ;
  assign n33255 = \core_c_psq_ststk_sts7x23_STcell_reg[1][20]/P0001  & n14708 ;
  assign n33261 = ~n33254 & ~n33255 ;
  assign n33265 = n33260 & n33261 ;
  assign n33266 = n33264 & n33265 ;
  assign n33267 = ~n33252 & ~n33266 ;
  assign n33268 = n32367 & n33267 ;
  assign n33269 = \core_c_psq_ICNTL_reg_DO_reg[4]/NET0131  & ~n33245 ;
  assign n33270 = n32364 & ~n33269 ;
  assign n33271 = \core_c_psq_IMASK_reg[5]/NET0131  & ~n33270 ;
  assign n33272 = ~n32367 & n33271 ;
  assign n33273 = ~n33268 & ~n33272 ;
  assign n33274 = ~\core_c_dec_MFPSQ_Ei_reg/NET0131  & n4117 ;
  assign n33280 = ~\core_c_dec_IR_reg[2]/NET0131  & n19270 ;
  assign n33281 = ~n31653 & ~n33280 ;
  assign n33282 = n31264 & n33281 ;
  assign n33283 = n31978 & n33282 ;
  assign n33275 = \core_c_dec_IR_reg[2]/NET0131  & n31966 ;
  assign n33278 = n31974 & n33275 ;
  assign n33279 = n31969 & n33275 ;
  assign n33286 = ~n33278 & ~n33279 ;
  assign n33287 = ~n33283 & n33286 ;
  assign n33276 = n31981 & n33275 ;
  assign n33277 = ~n4117 & ~n33276 ;
  assign n33284 = n24442 & ~n25244 ;
  assign n33285 = ~n32025 & n33284 ;
  assign n33288 = n33277 & n33285 ;
  assign n33289 = n33287 & n33288 ;
  assign n33290 = ~n33274 & ~n33289 ;
  assign n33291 = n13739 & n13764 ;
  assign n33292 = ~\bdma_BWCOUNT_reg[7]/NET0131  & n33291 ;
  assign n33293 = ~\bdma_BWCOUNT_reg[8]/NET0131  & n33292 ;
  assign n33294 = ~\bdma_BWCOUNT_reg[9]/NET0131  & n33293 ;
  assign n33295 = ~\bdma_BWCOUNT_reg[10]/NET0131  & n33294 ;
  assign n33296 = ~\bdma_BWCOUNT_reg[11]/NET0131  & n33295 ;
  assign n33297 = ~\bdma_BWCOUNT_reg[12]/NET0131  & n33296 ;
  assign n33298 = ~\bdma_BWCOUNT_reg[13]/NET0131  & ~n33297 ;
  assign n33299 = \bdma_BWCOUNT_reg[13]/NET0131  & n33297 ;
  assign n33300 = ~n33298 & ~n33299 ;
  assign n33301 = ~n13763 & ~n33300 ;
  assign n33302 = ~n7340 & n13763 ;
  assign n33303 = ~n33301 & ~n33302 ;
  assign n33304 = \bdma_BEAD_reg[2]/NET0131  & n20769 ;
  assign n33305 = \bdma_BEAD_reg[3]/NET0131  & n33304 ;
  assign n33306 = \bdma_BEAD_reg[4]/NET0131  & n33305 ;
  assign n33307 = \bdma_BEAD_reg[5]/NET0131  & n33306 ;
  assign n33308 = \bdma_BEAD_reg[6]/NET0131  & n33307 ;
  assign n33309 = \bdma_BEAD_reg[7]/NET0131  & n33308 ;
  assign n33310 = \bdma_BEAD_reg[8]/NET0131  & n33309 ;
  assign n33311 = \bdma_BEAD_reg[9]/NET0131  & n33310 ;
  assign n33312 = \bdma_BEAD_reg[10]/NET0131  & n33311 ;
  assign n33313 = \bdma_BEAD_reg[11]/NET0131  & n33312 ;
  assign n33315 = ~\bdma_BEAD_reg[12]/NET0131  & ~n33313 ;
  assign n33314 = \bdma_BEAD_reg[12]/NET0131  & n33313 ;
  assign n33316 = ~n20765 & ~n33314 ;
  assign n33317 = ~n33315 & n33316 ;
  assign n33318 = n9178 & n20765 ;
  assign n33319 = ~n33317 & ~n33318 ;
  assign n33322 = n18271 & ~n19559 ;
  assign n33321 = ~\core_eu_em_mac_em_reg_mr0swe_DO_reg[0]/P0001  & ~n18271 ;
  assign n33323 = n18273 & ~n33321 ;
  assign n33324 = ~n33322 & n33323 ;
  assign n33320 = \core_eu_em_mac_em_reg_mr0swe_DO_reg[0]/P0001  & ~n18266 ;
  assign n33325 = ~n18270 & ~n33320 ;
  assign n33326 = ~n33324 & n33325 ;
  assign n33327 = ~n18262 & ~n33326 ;
  assign n33328 = n18262 & ~n19653 ;
  assign n33329 = ~n33327 & ~n33328 ;
  assign n33330 = n14752 & n19653 ;
  assign n33331 = n18328 & n19559 ;
  assign n33332 = \core_eu_em_mac_em_reg_mr0rwe_DO_reg[0]/P0001  & ~n18330 ;
  assign n33333 = n18334 & ~n33332 ;
  assign n33334 = ~n33331 & n33333 ;
  assign n33335 = ~n33330 & ~n33334 ;
  assign n33336 = \core_c_psq_cntstk_ptr_reg[2]/NET0131  & ~n13778 ;
  assign n33341 = ~n5950 & ~n27920 ;
  assign n33338 = ~\core_c_psq_Eqend_Ed_reg/P0001  & ~n13777 ;
  assign n33339 = ~n27907 & n33338 ;
  assign n33340 = ~n27911 & n33339 ;
  assign n33342 = ~\core_c_psq_cntstk_ptr_reg[2]/NET0131  & ~n33340 ;
  assign n33343 = n33341 & n33342 ;
  assign n33344 = ~n13779 & ~n33343 ;
  assign n33345 = ~\core_c_psq_cntstk_ptr_reg[2]/NET0131  & n13778 ;
  assign n33337 = ~\core_c_psq_cntstk_ptr_reg[2]/NET0131  & ~n13784 ;
  assign n33346 = ~n13775 & ~n33337 ;
  assign n33347 = ~n33345 & n33346 ;
  assign n33348 = ~n33344 & n33347 ;
  assign n33349 = ~n33336 & ~n33348 ;
  assign n33350 = ~\core_c_psq_cntstk_ptr_reg[0]/NET0131  & ~n33344 ;
  assign n33351 = \core_c_psq_cntstk_ptr_reg[0]/NET0131  & n33344 ;
  assign n33352 = ~n33350 & ~n33351 ;
  assign n33356 = \core_c_psq_ststk_sts7x23_STcell_reg[0][14]/P0001  & n14702 ;
  assign n33357 = \core_c_psq_ststk_sts7x23_STcell_reg[5][14]/P0001  & n14699 ;
  assign n33362 = ~n33356 & ~n33357 ;
  assign n33358 = \core_c_psq_ststk_sts7x23_STcell_reg[4][14]/P0001  & n14706 ;
  assign n33359 = \core_c_psq_ststk_sts7x23_STcell_reg[2][14]/P0001  & n14713 ;
  assign n33363 = ~n33358 & ~n33359 ;
  assign n33364 = n33362 & n33363 ;
  assign n33353 = \core_c_psq_ststk_sts7x23_STcell_reg[6][14]/P0001  & n14711 ;
  assign n33360 = ~\core_c_dec_Modctl_Eg_reg/P0001  & ~n33353 ;
  assign n33354 = \core_c_psq_ststk_sts7x23_STcell_reg[3][14]/P0001  & n14704 ;
  assign n33355 = \core_c_psq_ststk_sts7x23_STcell_reg[1][14]/P0001  & n14708 ;
  assign n33361 = ~n33354 & ~n33355 ;
  assign n33365 = n33360 & n33361 ;
  assign n33366 = n33364 & n33365 ;
  assign n33367 = ~\core_c_dec_IRE_reg[3]/NET0131  & \core_c_psq_MSTAT_reg_DO_reg[6]/NET0131  ;
  assign n33368 = \core_c_dec_Modctl_Eg_reg/P0001  & ~n6071 ;
  assign n33369 = ~n33367 & n33368 ;
  assign n33370 = ~\core_c_dec_MTMSTAT_Eg_reg/P0001  & ~n33369 ;
  assign n33371 = ~n33366 & n33370 ;
  assign n33372 = \core_c_dec_MTMSTAT_Eg_reg/P0001  & n11525 ;
  assign n33373 = ~n33371 & ~n33372 ;
  assign n33374 = n23243 & ~n33373 ;
  assign n33375 = \core_c_psq_MSTAT_reg_DO_reg[6]/NET0131  & ~n23243 ;
  assign n33376 = ~n33374 & ~n33375 ;
  assign n33384 = \core_c_psq_ststk_sts7x23_STcell_reg[2][13]/P0001  & n14713 ;
  assign n33385 = \core_c_psq_ststk_sts7x23_STcell_reg[5][13]/P0001  & n14699 ;
  assign n33390 = ~n33384 & ~n33385 ;
  assign n33386 = \core_c_psq_ststk_sts7x23_STcell_reg[1][13]/P0001  & n14708 ;
  assign n33387 = \core_c_psq_ststk_sts7x23_STcell_reg[3][13]/P0001  & n14704 ;
  assign n33391 = ~n33386 & ~n33387 ;
  assign n33392 = n33390 & n33391 ;
  assign n33381 = \core_c_psq_ststk_sts7x23_STcell_reg[0][13]/P0001  & n14702 ;
  assign n33388 = ~\core_c_dec_Modctl_Eg_reg/P0001  & ~n33381 ;
  assign n33382 = \core_c_psq_ststk_sts7x23_STcell_reg[4][13]/P0001  & n14706 ;
  assign n33383 = \core_c_psq_ststk_sts7x23_STcell_reg[6][13]/P0001  & n14711 ;
  assign n33389 = ~n33382 & ~n33383 ;
  assign n33393 = n33388 & n33389 ;
  assign n33394 = n33392 & n33393 ;
  assign n33378 = \core_c_dec_IRE_reg[14]/NET0131  & \core_c_dec_IRE_reg[15]/NET0131  ;
  assign n33377 = ~\core_c_dec_IRE_reg[15]/NET0131  & \core_c_psq_MSTAT_reg_DO_reg[5]/NET0131  ;
  assign n33379 = \core_c_dec_Modctl_Eg_reg/P0001  & ~n33377 ;
  assign n33380 = ~n33378 & n33379 ;
  assign n33395 = ~\core_c_dec_MTMSTAT_Eg_reg/P0001  & ~n33380 ;
  assign n33396 = ~n33394 & n33395 ;
  assign n33397 = \core_c_dec_MTMSTAT_Eg_reg/P0001  & n10911 ;
  assign n33398 = ~n33396 & ~n33397 ;
  assign n33399 = n23243 & ~n33398 ;
  assign n33400 = \core_c_psq_MSTAT_reg_DO_reg[5]/NET0131  & ~n23243 ;
  assign n33401 = ~n33399 & ~n33400 ;
  assign n33409 = \core_c_psq_ststk_sts7x23_STcell_reg[6][11]/P0001  & n14711 ;
  assign n33410 = \core_c_psq_ststk_sts7x23_STcell_reg[1][11]/P0001  & n14708 ;
  assign n33415 = ~n33409 & ~n33410 ;
  assign n33411 = \core_c_psq_ststk_sts7x23_STcell_reg[5][11]/P0001  & n14699 ;
  assign n33412 = \core_c_psq_ststk_sts7x23_STcell_reg[3][11]/P0001  & n14704 ;
  assign n33416 = ~n33411 & ~n33412 ;
  assign n33417 = n33415 & n33416 ;
  assign n33406 = \core_c_psq_ststk_sts7x23_STcell_reg[0][11]/P0001  & n14702 ;
  assign n33413 = ~\core_c_dec_Modctl_Eg_reg/P0001  & ~n33406 ;
  assign n33407 = \core_c_psq_ststk_sts7x23_STcell_reg[4][11]/P0001  & n14706 ;
  assign n33408 = \core_c_psq_ststk_sts7x23_STcell_reg[2][11]/P0001  & n14713 ;
  assign n33414 = ~n33407 & ~n33408 ;
  assign n33418 = n33413 & n33414 ;
  assign n33419 = n33417 & n33418 ;
  assign n33403 = \core_c_dec_IRE_reg[10]/NET0131  & \core_c_dec_IRE_reg[13]/NET0131  ;
  assign n33402 = ~\core_c_dec_IRE_reg[13]/NET0131  & \core_c_psq_MSTAT_reg_DO_reg[3]/NET0131  ;
  assign n33404 = \core_c_dec_Modctl_Eg_reg/P0001  & ~n33402 ;
  assign n33405 = ~n33403 & n33404 ;
  assign n33420 = ~\core_c_dec_MTMSTAT_Eg_reg/P0001  & ~n33405 ;
  assign n33421 = ~n33419 & n33420 ;
  assign n33422 = \core_c_dec_MTMSTAT_Eg_reg/P0001  & n8113 ;
  assign n33423 = ~n33421 & ~n33422 ;
  assign n33424 = n23243 & ~n33423 ;
  assign n33425 = \core_c_psq_MSTAT_reg_DO_reg[3]/NET0131  & ~n23243 ;
  assign n33426 = ~n33424 & ~n33425 ;
  assign n33430 = \core_c_psq_ststk_sts7x23_STcell_reg[4][10]/P0001  & n14706 ;
  assign n33431 = \core_c_psq_ststk_sts7x23_STcell_reg[1][10]/P0001  & n14708 ;
  assign n33436 = ~n33430 & ~n33431 ;
  assign n33432 = \core_c_psq_ststk_sts7x23_STcell_reg[3][10]/P0001  & n14704 ;
  assign n33433 = \core_c_psq_ststk_sts7x23_STcell_reg[6][10]/P0001  & n14711 ;
  assign n33437 = ~n33432 & ~n33433 ;
  assign n33438 = n33436 & n33437 ;
  assign n33427 = \core_c_psq_ststk_sts7x23_STcell_reg[5][10]/P0001  & n14699 ;
  assign n33434 = ~\core_c_dec_Modctl_Eg_reg/P0001  & ~n33427 ;
  assign n33428 = \core_c_psq_ststk_sts7x23_STcell_reg[2][10]/P0001  & n14713 ;
  assign n33429 = \core_c_psq_ststk_sts7x23_STcell_reg[0][10]/P0001  & n14702 ;
  assign n33435 = ~n33428 & ~n33429 ;
  assign n33439 = n33434 & n33435 ;
  assign n33440 = n33438 & n33439 ;
  assign n33441 = ~\core_c_dec_IRE_reg[9]/NET0131  & \core_c_psq_MSTAT_reg_DO_reg[2]/NET0131  ;
  assign n33442 = \core_c_dec_Modctl_Eg_reg/P0001  & ~n13818 ;
  assign n33443 = ~n33441 & n33442 ;
  assign n33444 = ~\core_c_dec_MTMSTAT_Eg_reg/P0001  & ~n33443 ;
  assign n33445 = ~n33440 & n33444 ;
  assign n33446 = \core_c_dec_MTMSTAT_Eg_reg/P0001  & n8715 ;
  assign n33447 = ~n33445 & ~n33446 ;
  assign n33448 = n23243 & ~n33447 ;
  assign n33449 = \core_c_psq_MSTAT_reg_DO_reg[2]/NET0131  & ~n23243 ;
  assign n33450 = ~n33448 & ~n33449 ;
  assign n33458 = \core_c_psq_ststk_sts7x23_STcell_reg[2][9]/P0001  & n14713 ;
  assign n33459 = \core_c_psq_ststk_sts7x23_STcell_reg[5][9]/P0001  & n14699 ;
  assign n33464 = ~n33458 & ~n33459 ;
  assign n33460 = \core_c_psq_ststk_sts7x23_STcell_reg[1][9]/P0001  & n14708 ;
  assign n33461 = \core_c_psq_ststk_sts7x23_STcell_reg[3][9]/P0001  & n14704 ;
  assign n33465 = ~n33460 & ~n33461 ;
  assign n33466 = n33464 & n33465 ;
  assign n33455 = \core_c_psq_ststk_sts7x23_STcell_reg[0][9]/P0001  & n14702 ;
  assign n33462 = ~\core_c_dec_Modctl_Eg_reg/P0001  & ~n33455 ;
  assign n33456 = \core_c_psq_ststk_sts7x23_STcell_reg[4][9]/P0001  & n14706 ;
  assign n33457 = \core_c_psq_ststk_sts7x23_STcell_reg[6][9]/P0001  & n14711 ;
  assign n33463 = ~n33456 & ~n33457 ;
  assign n33467 = n33462 & n33463 ;
  assign n33468 = n33466 & n33467 ;
  assign n33452 = \core_c_dec_IRE_reg[5]/NET0131  & \core_c_dec_IRE_reg[6]/NET0131  ;
  assign n33451 = ~\core_c_dec_IRE_reg[5]/NET0131  & \core_c_psq_MSTAT_reg_DO_reg[1]/NET0131  ;
  assign n33453 = \core_c_dec_Modctl_Eg_reg/P0001  & ~n33451 ;
  assign n33454 = ~n33452 & n33453 ;
  assign n33469 = ~\core_c_dec_MTMSTAT_Eg_reg/P0001  & ~n33454 ;
  assign n33470 = ~n33468 & n33469 ;
  assign n33471 = \core_c_dec_MTMSTAT_Eg_reg/P0001  & n9435 ;
  assign n33472 = ~n33470 & ~n33471 ;
  assign n33473 = n23243 & ~n33472 ;
  assign n33474 = \core_c_psq_MSTAT_reg_DO_reg[1]/NET0131  & ~n23243 ;
  assign n33475 = ~n33473 & ~n33474 ;
  assign n33476 = \core_c_dec_MTIMASK_Eg_reg/P0001  & ~n10289 ;
  assign n33480 = \core_c_psq_ststk_sts7x23_STcell_reg[3][24]/P0001  & n14704 ;
  assign n33481 = \core_c_psq_ststk_sts7x23_STcell_reg[5][24]/P0001  & n14699 ;
  assign n33486 = ~n33480 & ~n33481 ;
  assign n33482 = \core_c_psq_ststk_sts7x23_STcell_reg[6][24]/P0001  & n14711 ;
  assign n33483 = \core_c_psq_ststk_sts7x23_STcell_reg[0][24]/P0001  & n14702 ;
  assign n33487 = ~n33482 & ~n33483 ;
  assign n33488 = n33486 & n33487 ;
  assign n33477 = \core_c_psq_ststk_sts7x23_STcell_reg[2][24]/P0001  & n14713 ;
  assign n33484 = ~\core_c_dec_MTIMASK_Eg_reg/P0001  & ~n33477 ;
  assign n33478 = \core_c_psq_ststk_sts7x23_STcell_reg[4][24]/P0001  & n14706 ;
  assign n33479 = \core_c_psq_ststk_sts7x23_STcell_reg[1][24]/P0001  & n14708 ;
  assign n33485 = ~n33478 & ~n33479 ;
  assign n33489 = n33484 & n33485 ;
  assign n33490 = n33488 & n33489 ;
  assign n33491 = ~n33476 & ~n33490 ;
  assign n33492 = n32367 & n33491 ;
  assign n33493 = ~\core_c_psq_Iact_E_reg[6]/NET0131  & n33246 ;
  assign n33494 = ~\core_c_psq_Iact_E_reg[7]/NET0131  & n33493 ;
  assign n33495 = ~\core_c_psq_Iact_E_reg[8]/NET0131  & n33494 ;
  assign n33496 = \core_c_psq_ICNTL_reg_DO_reg[4]/NET0131  & ~n33495 ;
  assign n33497 = n32364 & ~n33496 ;
  assign n33498 = \core_c_psq_IMASK_reg[9]/NET0131  & ~n33497 ;
  assign n33499 = ~n32367 & n33498 ;
  assign n33500 = ~n33492 & ~n33499 ;
  assign n33501 = \core_c_dec_MTIMASK_Eg_reg/P0001  & ~n9435 ;
  assign n33505 = \core_c_psq_ststk_sts7x23_STcell_reg[5][16]/P0001  & n14699 ;
  assign n33506 = \core_c_psq_ststk_sts7x23_STcell_reg[3][16]/P0001  & n14704 ;
  assign n33511 = ~n33505 & ~n33506 ;
  assign n33507 = \core_c_psq_ststk_sts7x23_STcell_reg[0][16]/P0001  & n14702 ;
  assign n33508 = \core_c_psq_ststk_sts7x23_STcell_reg[4][16]/P0001  & n14706 ;
  assign n33512 = ~n33507 & ~n33508 ;
  assign n33513 = n33511 & n33512 ;
  assign n33502 = \core_c_psq_ststk_sts7x23_STcell_reg[1][16]/P0001  & n14708 ;
  assign n33509 = ~\core_c_dec_MTIMASK_Eg_reg/P0001  & ~n33502 ;
  assign n33503 = \core_c_psq_ststk_sts7x23_STcell_reg[2][16]/P0001  & n14713 ;
  assign n33504 = \core_c_psq_ststk_sts7x23_STcell_reg[6][16]/P0001  & n14711 ;
  assign n33510 = ~n33503 & ~n33504 ;
  assign n33514 = n33509 & n33510 ;
  assign n33515 = n33513 & n33514 ;
  assign n33516 = ~n33501 & ~n33515 ;
  assign n33517 = n32367 & n33516 ;
  assign n33518 = \core_c_psq_ICNTL_reg_DO_reg[4]/NET0131  & \core_c_psq_Iact_E_reg[0]/NET0131  ;
  assign n33519 = n32364 & ~n33518 ;
  assign n33520 = \core_c_psq_IMASK_reg[1]/NET0131  & ~n33519 ;
  assign n33521 = ~n32367 & n33520 ;
  assign n33522 = ~n33517 & ~n33521 ;
  assign n33523 = ~n4117 & n31648 ;
  assign n33524 = \core_c_dec_MFSR1_E_reg/P0001  & n4117 ;
  assign n33525 = ~n33523 & ~n33524 ;
  assign n33526 = ~n4117 & n31649 ;
  assign n33527 = \core_c_dec_MFSR0_E_reg/P0001  & n4117 ;
  assign n33528 = ~n33526 & ~n33527 ;
  assign n33529 = ~n4117 & n31656 ;
  assign n33530 = \core_c_dec_MFSI_E_reg/P0001  & n4117 ;
  assign n33531 = ~n33529 & ~n33530 ;
  assign n33532 = ~n4117 & n31652 ;
  assign n33533 = \core_c_dec_MFSE_E_reg/P0001  & n4117 ;
  assign n33534 = ~n33532 & ~n33533 ;
  assign n33535 = \core_c_dec_MFMX1_E_reg/P0001  & n4117 ;
  assign n33536 = n30962 & n32643 ;
  assign n33537 = ~n33535 & ~n33536 ;
  assign n33538 = ~n4117 & n30979 ;
  assign n33539 = \core_c_dec_MFMR2_E_reg/P0001  & n4117 ;
  assign n33540 = ~n33538 & ~n33539 ;
  assign n33541 = ~n4117 & n30982 ;
  assign n33542 = \core_c_dec_MFMR1_E_reg/P0001  & n4117 ;
  assign n33543 = ~n33541 & ~n33542 ;
  assign n33544 = ~n4117 & n30968 ;
  assign n33545 = \core_c_dec_MFMR0_E_reg/P0001  & n4117 ;
  assign n33546 = ~n33544 & ~n33545 ;
  assign n33547 = \core_c_dec_MFAX1_E_reg/P0001  & n4117 ;
  assign n33548 = n31650 & n32643 ;
  assign n33549 = ~n33547 & ~n33548 ;
  assign n33550 = ~n4117 & n31260 ;
  assign n33551 = \core_c_dec_MFAR_E_reg/P0001  & n4117 ;
  assign n33552 = ~n33550 & ~n33551 ;
  assign n33553 = \sport1_regs_MWORDreg_DO_reg[7]/NET0131  & ~n32612 ;
  assign n33554 = n20407 & n32616 ;
  assign n33555 = \sport1_rxctl_Wcnt_reg[7]/NET0131  & ~n33554 ;
  assign n33556 = n32612 & n33555 ;
  assign n33557 = ~n33553 & ~n33556 ;
  assign n33558 = ~\sport1_rxctl_Wcnt_reg[5]/NET0131  & n32618 ;
  assign n33559 = \sport1_rxctl_Wcnt_reg[6]/NET0131  & ~n33558 ;
  assign n33560 = ~n33554 & ~n33559 ;
  assign n33561 = n32612 & ~n33560 ;
  assign n33562 = \sport1_regs_MWORDreg_DO_reg[6]/NET0131  & ~n32612 ;
  assign n33563 = ~n33561 & ~n33562 ;
  assign n33564 = ~\sport1_regs_MWORDreg_DO_reg[5]/NET0131  & ~n32612 ;
  assign n33565 = \sport1_rxctl_Wcnt_reg[5]/NET0131  & ~n32618 ;
  assign n33566 = ~n33558 & ~n33565 ;
  assign n33567 = n32612 & n33566 ;
  assign n33568 = ~n33564 & ~n33567 ;
  assign n33569 = \sport1_regs_MWORDreg_DO_reg[3]/NET0131  & ~n32612 ;
  assign n33570 = \sport1_rxctl_Wcnt_reg[3]/NET0131  & ~n32615 ;
  assign n33571 = ~n32616 & ~n33570 ;
  assign n33572 = n32612 & ~n33571 ;
  assign n33573 = ~n33569 & ~n33572 ;
  assign n33574 = ~\sport1_regs_MWORDreg_DO_reg[2]/NET0131  & ~n32612 ;
  assign n33575 = \sport1_rxctl_Wcnt_reg[2]/NET0131  & ~n32614 ;
  assign n33576 = ~n32615 & ~n33575 ;
  assign n33577 = n32612 & n33576 ;
  assign n33578 = ~n33574 & ~n33577 ;
  assign n33579 = ~\sport1_rxctl_Wcnt_reg[0]/NET0131  & n32613 ;
  assign n33580 = \sport1_rxctl_Wcnt_reg[1]/NET0131  & ~n33579 ;
  assign n33581 = ~n32614 & ~n33580 ;
  assign n33582 = n32612 & ~n33581 ;
  assign n33583 = \sport1_regs_MWORDreg_DO_reg[1]/NET0131  & ~n32612 ;
  assign n33584 = ~n33582 & ~n33583 ;
  assign n33585 = \sport1_rxctl_Wcnt_reg[0]/NET0131  & ~n32613 ;
  assign n33586 = ~n33579 & ~n33585 ;
  assign n33587 = n32612 & ~n33586 ;
  assign n33588 = \sport1_regs_MWORDreg_DO_reg[0]/NET0131  & ~n32612 ;
  assign n33589 = ~n33587 & ~n33588 ;
  assign n33590 = \sport0_regs_MWORDreg_DO_reg[7]/NET0131  & ~n32658 ;
  assign n33591 = n20429 & n32662 ;
  assign n33592 = \sport0_rxctl_Wcnt_reg[7]/NET0131  & ~n33591 ;
  assign n33593 = n32658 & n33592 ;
  assign n33594 = ~n33590 & ~n33593 ;
  assign n33595 = ~\sport0_regs_MWORDreg_DO_reg[5]/NET0131  & ~n32658 ;
  assign n33596 = \sport0_rxctl_Wcnt_reg[5]/NET0131  & ~n32664 ;
  assign n33597 = ~\sport0_rxctl_Wcnt_reg[5]/NET0131  & n32664 ;
  assign n33598 = ~n33596 & ~n33597 ;
  assign n33599 = n32658 & n33598 ;
  assign n33600 = ~n33595 & ~n33599 ;
  assign n33601 = \sport0_regs_MWORDreg_DO_reg[3]/NET0131  & ~n32658 ;
  assign n33602 = \sport0_rxctl_Wcnt_reg[3]/NET0131  & ~n32661 ;
  assign n33603 = ~n32662 & ~n33602 ;
  assign n33604 = n32658 & ~n33603 ;
  assign n33605 = ~n33601 & ~n33604 ;
  assign n33606 = ~\sport0_rxctl_Wcnt_reg[0]/NET0131  & n32659 ;
  assign n33607 = \sport0_rxctl_Wcnt_reg[1]/NET0131  & ~n33606 ;
  assign n33608 = ~n32660 & ~n33607 ;
  assign n33609 = n32658 & ~n33608 ;
  assign n33610 = \sport0_regs_MWORDreg_DO_reg[1]/NET0131  & ~n32658 ;
  assign n33611 = ~n33609 & ~n33610 ;
  assign n33612 = \sport0_rxctl_Wcnt_reg[0]/NET0131  & ~n32659 ;
  assign n33613 = ~n33606 & ~n33612 ;
  assign n33614 = n32658 & ~n33613 ;
  assign n33615 = \sport0_regs_MWORDreg_DO_reg[0]/NET0131  & ~n32658 ;
  assign n33616 = ~n33614 & ~n33615 ;
  assign n33617 = \clkc_oscntr_reg_DO_reg[10]/NET0131  & n23424 ;
  assign n33618 = \clkc_oscntr_reg_DO_reg[11]/NET0131  & ~n33617 ;
  assign n33619 = ~\clkc_oscntr_reg_DO_reg[11]/NET0131  & n33617 ;
  assign n33620 = ~n33618 & ~n33619 ;
  assign n33621 = ~\sport0_regs_MWORDreg_DO_reg[2]/NET0131  & ~n32658 ;
  assign n33622 = \sport0_rxctl_Wcnt_reg[2]/NET0131  & ~n32660 ;
  assign n33623 = ~n32661 & ~n33622 ;
  assign n33624 = n32658 & n33623 ;
  assign n33625 = ~n33621 & ~n33624 ;
  assign n33626 = \sport0_rxctl_Wcnt_reg[6]/NET0131  & ~n33597 ;
  assign n33627 = ~n33591 & ~n33626 ;
  assign n33628 = n32658 & ~n33627 ;
  assign n33629 = \sport0_regs_MWORDreg_DO_reg[6]/NET0131  & ~n32658 ;
  assign n33630 = ~n33628 & ~n33629 ;
  assign n33631 = ~\sice_IIRC_reg[16]/NET0131  & ~n22581 ;
  assign n33632 = ~n22582 & ~n33631 ;
  assign n33633 = \core_c_dec_MFAX0_E_reg/P0001  & n4117 ;
  assign n33634 = n31650 & n32639 ;
  assign n33635 = ~n33633 & ~n33634 ;
  assign n33636 = n10289 & ~n32992 ;
  assign n33637 = \core_dag_ilm2reg_L6_we_DO_reg[9]/NET0131  & n32994 ;
  assign n33641 = ~n21579 & ~n33637 ;
  assign n33640 = \core_dag_ilm2reg_L5_we_DO_reg[9]/NET0131  & n33000 ;
  assign n33638 = \core_dag_ilm2reg_L4_we_DO_reg[9]/NET0131  & n32996 ;
  assign n33639 = \core_dag_ilm2reg_L7_we_DO_reg[9]/NET0131  & n32998 ;
  assign n33642 = ~n33638 & ~n33639 ;
  assign n33643 = ~n33640 & n33642 ;
  assign n33644 = n33641 & n33643 ;
  assign n33645 = ~n33636 & n33644 ;
  assign n33646 = ~\core_dag_ilm2reg_L_reg[9]/NET0131  & n21579 ;
  assign n33647 = ~n33645 & ~n33646 ;
  assign n33648 = n10638 & ~n32992 ;
  assign n33649 = \core_dag_ilm2reg_L6_we_DO_reg[8]/NET0131  & n32994 ;
  assign n33653 = ~n21579 & ~n33649 ;
  assign n33652 = \core_dag_ilm2reg_L5_we_DO_reg[8]/NET0131  & n33000 ;
  assign n33650 = \core_dag_ilm2reg_L4_we_DO_reg[8]/NET0131  & n32996 ;
  assign n33651 = \core_dag_ilm2reg_L7_we_DO_reg[8]/NET0131  & n32998 ;
  assign n33654 = ~n33650 & ~n33651 ;
  assign n33655 = ~n33652 & n33654 ;
  assign n33656 = n33653 & n33655 ;
  assign n33657 = ~n33648 & n33656 ;
  assign n33658 = ~\core_dag_ilm2reg_L_reg[8]/NET0131  & n21579 ;
  assign n33659 = ~n33657 & ~n33658 ;
  assign n33660 = n9178 & ~n32992 ;
  assign n33661 = \core_dag_ilm2reg_L6_we_DO_reg[12]/NET0131  & n32994 ;
  assign n33665 = ~n21579 & ~n33661 ;
  assign n33664 = \core_dag_ilm2reg_L5_we_DO_reg[12]/NET0131  & n33000 ;
  assign n33662 = \core_dag_ilm2reg_L4_we_DO_reg[12]/NET0131  & n32996 ;
  assign n33663 = \core_dag_ilm2reg_L7_we_DO_reg[12]/NET0131  & n32998 ;
  assign n33666 = ~n33662 & ~n33663 ;
  assign n33667 = ~n33664 & n33666 ;
  assign n33668 = n33665 & n33667 ;
  assign n33669 = ~n33660 & n33668 ;
  assign n33670 = ~\core_dag_ilm2reg_L_reg[12]/NET0131  & n21579 ;
  assign n33671 = ~n33669 & ~n33670 ;
  assign n33672 = n8460 & ~n32992 ;
  assign n33673 = \core_dag_ilm2reg_L6_we_DO_reg[11]/NET0131  & n32994 ;
  assign n33677 = ~n21579 & ~n33673 ;
  assign n33676 = \core_dag_ilm2reg_L5_we_DO_reg[11]/NET0131  & n33000 ;
  assign n33674 = \core_dag_ilm2reg_L4_we_DO_reg[11]/NET0131  & n32996 ;
  assign n33675 = \core_dag_ilm2reg_L7_we_DO_reg[11]/NET0131  & n32998 ;
  assign n33678 = ~n33674 & ~n33675 ;
  assign n33679 = ~n33676 & n33678 ;
  assign n33680 = n33677 & n33679 ;
  assign n33681 = ~n33672 & n33680 ;
  assign n33682 = ~\core_dag_ilm2reg_L_reg[11]/NET0131  & n21579 ;
  assign n33683 = ~n33681 & ~n33682 ;
  assign n33692 = ~n6008 & n32984 ;
  assign n33693 = ~n5964 & n32986 ;
  assign n33696 = ~n33692 & ~n33693 ;
  assign n33694 = ~n6000 & n32988 ;
  assign n33695 = ~n6015 & n32982 ;
  assign n33697 = ~n33694 & ~n33695 ;
  assign n33698 = n33696 & n33697 ;
  assign n33699 = n20755 & ~n33698 ;
  assign n33684 = n6008 & n32984 ;
  assign n33685 = \core_dag_ilm2reg_I6_we_DO_reg[9]/NET0131  & n33684 ;
  assign n33700 = ~n21579 & ~n33685 ;
  assign n33690 = n5964 & n32986 ;
  assign n33691 = \core_dag_ilm2reg_I4_we_DO_reg[9]/NET0131  & n33690 ;
  assign n33686 = n6000 & n32988 ;
  assign n33687 = \core_dag_ilm2reg_I7_we_DO_reg[9]/NET0131  & n33686 ;
  assign n33688 = n6015 & n32982 ;
  assign n33689 = \core_dag_ilm2reg_I5_we_DO_reg[9]/NET0131  & n33688 ;
  assign n33701 = ~n33687 & ~n33689 ;
  assign n33702 = ~n33691 & n33701 ;
  assign n33703 = n33700 & n33702 ;
  assign n33704 = ~n33699 & n33703 ;
  assign n33705 = ~\core_dag_ilm2reg_I_reg[9]/NET0131  & n21579 ;
  assign n33706 = ~n33704 & ~n33705 ;
  assign n33711 = n20624 & ~n33698 ;
  assign n33707 = \core_dag_ilm2reg_I6_we_DO_reg[6]/NET0131  & n33684 ;
  assign n33712 = ~n21579 & ~n33707 ;
  assign n33710 = \core_dag_ilm2reg_I4_we_DO_reg[6]/NET0131  & n33690 ;
  assign n33708 = \core_dag_ilm2reg_I7_we_DO_reg[6]/NET0131  & n33686 ;
  assign n33709 = \core_dag_ilm2reg_I5_we_DO_reg[6]/NET0131  & n33688 ;
  assign n33713 = ~n33708 & ~n33709 ;
  assign n33714 = ~n33710 & n33713 ;
  assign n33715 = n33712 & n33714 ;
  assign n33716 = ~n33711 & n33715 ;
  assign n33717 = ~\core_dag_ilm2reg_I_reg[6]/NET0131  & n21579 ;
  assign n33718 = ~n33716 & ~n33717 ;
  assign n33723 = n20634 & ~n33698 ;
  assign n33719 = \core_dag_ilm2reg_I6_we_DO_reg[5]/NET0131  & n33684 ;
  assign n33724 = ~n21579 & ~n33719 ;
  assign n33722 = \core_dag_ilm2reg_I4_we_DO_reg[5]/NET0131  & n33690 ;
  assign n33720 = \core_dag_ilm2reg_I7_we_DO_reg[5]/NET0131  & n33686 ;
  assign n33721 = \core_dag_ilm2reg_I5_we_DO_reg[5]/NET0131  & n33688 ;
  assign n33725 = ~n33720 & ~n33721 ;
  assign n33726 = ~n33722 & n33725 ;
  assign n33727 = n33724 & n33726 ;
  assign n33728 = ~n33723 & n33727 ;
  assign n33729 = ~\core_dag_ilm2reg_I_reg[5]/NET0131  & n21579 ;
  assign n33730 = ~n33728 & ~n33729 ;
  assign n33735 = n20644 & ~n33698 ;
  assign n33731 = \core_dag_ilm2reg_I6_we_DO_reg[4]/NET0131  & n33684 ;
  assign n33736 = ~n21579 & ~n33731 ;
  assign n33734 = \core_dag_ilm2reg_I4_we_DO_reg[4]/NET0131  & n33690 ;
  assign n33732 = \core_dag_ilm2reg_I7_we_DO_reg[4]/NET0131  & n33686 ;
  assign n33733 = \core_dag_ilm2reg_I5_we_DO_reg[4]/NET0131  & n33688 ;
  assign n33737 = ~n33732 & ~n33733 ;
  assign n33738 = ~n33734 & n33737 ;
  assign n33739 = n33736 & n33738 ;
  assign n33740 = ~n33735 & n33739 ;
  assign n33741 = ~\core_dag_ilm2reg_I_reg[4]/NET0131  & n21579 ;
  assign n33742 = ~n33740 & ~n33741 ;
  assign n33747 = n13262 & ~n33698 ;
  assign n33743 = \core_dag_ilm2reg_I6_we_DO_reg[3]/NET0131  & n33684 ;
  assign n33748 = ~n21579 & ~n33743 ;
  assign n33746 = \core_dag_ilm2reg_I4_we_DO_reg[3]/NET0131  & n33690 ;
  assign n33744 = \core_dag_ilm2reg_I5_we_DO_reg[3]/NET0131  & n33688 ;
  assign n33745 = \core_dag_ilm2reg_I7_we_DO_reg[3]/NET0131  & n33686 ;
  assign n33749 = ~n33744 & ~n33745 ;
  assign n33750 = ~n33746 & n33749 ;
  assign n33751 = n33748 & n33750 ;
  assign n33752 = ~n33747 & n33751 ;
  assign n33753 = ~\core_dag_ilm2reg_I_reg[3]/NET0131  & n21579 ;
  assign n33754 = ~n33752 & ~n33753 ;
  assign n33759 = ~n20663 & ~n33698 ;
  assign n33755 = \core_dag_ilm2reg_I6_we_DO_reg[2]/NET0131  & n33684 ;
  assign n33760 = ~n21579 & ~n33755 ;
  assign n33758 = \core_dag_ilm2reg_I4_we_DO_reg[2]/NET0131  & n33690 ;
  assign n33756 = \core_dag_ilm2reg_I7_we_DO_reg[2]/NET0131  & n33686 ;
  assign n33757 = \core_dag_ilm2reg_I5_we_DO_reg[2]/NET0131  & n33688 ;
  assign n33761 = ~n33756 & ~n33757 ;
  assign n33762 = ~n33758 & n33761 ;
  assign n33763 = n33760 & n33762 ;
  assign n33764 = ~n33759 & n33763 ;
  assign n33765 = ~\core_dag_ilm2reg_I_reg[2]/NET0131  & n21579 ;
  assign n33766 = ~n33764 & ~n33765 ;
  assign n33771 = ~n20674 & ~n33698 ;
  assign n33767 = \core_dag_ilm2reg_I6_we_DO_reg[1]/NET0131  & n33684 ;
  assign n33772 = ~n21579 & ~n33767 ;
  assign n33770 = \core_dag_ilm2reg_I4_we_DO_reg[1]/NET0131  & n33690 ;
  assign n33768 = \core_dag_ilm2reg_I5_we_DO_reg[1]/NET0131  & n33688 ;
  assign n33769 = \core_dag_ilm2reg_I7_we_DO_reg[1]/NET0131  & n33686 ;
  assign n33773 = ~n33768 & ~n33769 ;
  assign n33774 = ~n33770 & n33773 ;
  assign n33775 = n33772 & n33774 ;
  assign n33776 = ~n33771 & n33775 ;
  assign n33777 = ~\core_dag_ilm2reg_I_reg[1]/NET0131  & n21579 ;
  assign n33778 = ~n33776 & ~n33777 ;
  assign n33783 = ~n20685 & ~n33698 ;
  assign n33779 = \core_dag_ilm2reg_I6_we_DO_reg[13]/NET0131  & n33684 ;
  assign n33784 = ~n21579 & ~n33779 ;
  assign n33782 = \core_dag_ilm2reg_I4_we_DO_reg[13]/NET0131  & n33690 ;
  assign n33780 = \core_dag_ilm2reg_I5_we_DO_reg[13]/NET0131  & n33688 ;
  assign n33781 = \core_dag_ilm2reg_I7_we_DO_reg[13]/NET0131  & n33686 ;
  assign n33785 = ~n33780 & ~n33781 ;
  assign n33786 = ~n33782 & n33785 ;
  assign n33787 = n33784 & n33786 ;
  assign n33788 = ~n33783 & n33787 ;
  assign n33789 = ~\core_dag_ilm2reg_I_reg[13]/NET0131  & n21579 ;
  assign n33790 = ~n33788 & ~n33789 ;
  assign n33795 = ~n20696 & ~n33698 ;
  assign n33791 = \core_dag_ilm2reg_I6_we_DO_reg[12]/NET0131  & n33684 ;
  assign n33796 = ~n21579 & ~n33791 ;
  assign n33794 = \core_dag_ilm2reg_I4_we_DO_reg[12]/NET0131  & n33690 ;
  assign n33792 = \core_dag_ilm2reg_I7_we_DO_reg[12]/NET0131  & n33686 ;
  assign n33793 = \core_dag_ilm2reg_I5_we_DO_reg[12]/NET0131  & n33688 ;
  assign n33797 = ~n33792 & ~n33793 ;
  assign n33798 = ~n33794 & n33797 ;
  assign n33799 = n33796 & n33798 ;
  assign n33800 = ~n33795 & n33799 ;
  assign n33801 = ~\core_dag_ilm2reg_I_reg[12]/NET0131  & n21579 ;
  assign n33802 = ~n33800 & ~n33801 ;
  assign n33807 = ~n20729 & ~n33698 ;
  assign n33803 = \core_dag_ilm2reg_I6_we_DO_reg[0]/NET0131  & n33684 ;
  assign n33808 = ~n21579 & ~n33803 ;
  assign n33806 = \core_dag_ilm2reg_I4_we_DO_reg[0]/NET0131  & n33690 ;
  assign n33804 = \core_dag_ilm2reg_I7_we_DO_reg[0]/NET0131  & n33686 ;
  assign n33805 = \core_dag_ilm2reg_I5_we_DO_reg[0]/NET0131  & n33688 ;
  assign n33809 = ~n33804 & ~n33805 ;
  assign n33810 = ~n33806 & n33809 ;
  assign n33811 = n33808 & n33810 ;
  assign n33812 = ~n33807 & n33811 ;
  assign n33813 = ~\core_dag_ilm2reg_I_reg[0]/NET0131  & n21579 ;
  assign n33814 = ~n33812 & ~n33813 ;
  assign n33815 = n10289 & ~n33099 ;
  assign n33816 = \core_dag_ilm1reg_L1_we_DO_reg[9]/NET0131  & n33105 ;
  assign n33817 = \core_dag_ilm1reg_L2_we_DO_reg[9]/NET0131  & n33107 ;
  assign n33820 = ~n33816 & ~n33817 ;
  assign n33818 = \core_dag_ilm1reg_L3_we_DO_reg[9]/NET0131  & n33101 ;
  assign n33819 = \core_dag_ilm1reg_L0_we_DO_reg[9]/NET0131  & n33103 ;
  assign n33821 = ~n33818 & ~n33819 ;
  assign n33822 = n33820 & n33821 ;
  assign n33823 = ~n21592 & n33822 ;
  assign n33824 = ~n33815 & n33823 ;
  assign n33825 = ~\core_dag_ilm1reg_L_reg[9]/NET0131  & n21592 ;
  assign n33826 = ~n33824 & ~n33825 ;
  assign n33827 = n10638 & ~n33099 ;
  assign n33828 = \core_dag_ilm1reg_L3_we_DO_reg[8]/NET0131  & n33101 ;
  assign n33829 = \core_dag_ilm1reg_L0_we_DO_reg[8]/NET0131  & n33103 ;
  assign n33832 = ~n33828 & ~n33829 ;
  assign n33830 = \core_dag_ilm1reg_L1_we_DO_reg[8]/NET0131  & n33105 ;
  assign n33831 = \core_dag_ilm1reg_L2_we_DO_reg[8]/NET0131  & n33107 ;
  assign n33833 = ~n33830 & ~n33831 ;
  assign n33834 = n33832 & n33833 ;
  assign n33835 = ~n21592 & n33834 ;
  assign n33836 = ~n33827 & n33835 ;
  assign n33837 = ~\core_dag_ilm1reg_L_reg[8]/NET0131  & n21592 ;
  assign n33838 = ~n33836 & ~n33837 ;
  assign n33839 = n7340 & ~n33099 ;
  assign n33840 = \core_dag_ilm1reg_L3_we_DO_reg[13]/NET0131  & n33101 ;
  assign n33841 = \core_dag_ilm1reg_L0_we_DO_reg[13]/NET0131  & n33103 ;
  assign n33844 = ~n33840 & ~n33841 ;
  assign n33842 = \core_dag_ilm1reg_L1_we_DO_reg[13]/NET0131  & n33105 ;
  assign n33843 = \core_dag_ilm1reg_L2_we_DO_reg[13]/NET0131  & n33107 ;
  assign n33845 = ~n33842 & ~n33843 ;
  assign n33846 = n33844 & n33845 ;
  assign n33847 = ~n21592 & n33846 ;
  assign n33848 = ~n33839 & n33847 ;
  assign n33849 = ~\core_dag_ilm1reg_L_reg[13]/NET0131  & n21592 ;
  assign n33850 = ~n33848 & ~n33849 ;
  assign n33851 = n9178 & ~n33099 ;
  assign n33852 = \core_dag_ilm1reg_L3_we_DO_reg[12]/NET0131  & n33101 ;
  assign n33853 = \core_dag_ilm1reg_L0_we_DO_reg[12]/NET0131  & n33103 ;
  assign n33856 = ~n33852 & ~n33853 ;
  assign n33854 = \core_dag_ilm1reg_L1_we_DO_reg[12]/NET0131  & n33105 ;
  assign n33855 = \core_dag_ilm1reg_L2_we_DO_reg[12]/NET0131  & n33107 ;
  assign n33857 = ~n33854 & ~n33855 ;
  assign n33858 = n33856 & n33857 ;
  assign n33859 = ~n21592 & n33858 ;
  assign n33860 = ~n33851 & n33859 ;
  assign n33861 = ~\core_dag_ilm1reg_L_reg[12]/NET0131  & n21592 ;
  assign n33862 = ~n33860 & ~n33861 ;
  assign n33863 = n8460 & ~n33099 ;
  assign n33864 = \core_dag_ilm1reg_L1_we_DO_reg[11]/NET0131  & n33105 ;
  assign n33865 = \core_dag_ilm1reg_L2_we_DO_reg[11]/NET0131  & n33107 ;
  assign n33868 = ~n33864 & ~n33865 ;
  assign n33866 = \core_dag_ilm1reg_L3_we_DO_reg[11]/NET0131  & n33101 ;
  assign n33867 = \core_dag_ilm1reg_L0_we_DO_reg[11]/NET0131  & n33103 ;
  assign n33869 = ~n33866 & ~n33867 ;
  assign n33870 = n33868 & n33869 ;
  assign n33871 = ~n21592 & n33870 ;
  assign n33872 = ~n33863 & n33871 ;
  assign n33873 = ~\core_dag_ilm1reg_L_reg[11]/NET0131  & n21592 ;
  assign n33874 = ~n33872 & ~n33873 ;
  assign n33875 = n7859 & ~n33099 ;
  assign n33876 = \core_dag_ilm1reg_L1_we_DO_reg[10]/NET0131  & n33105 ;
  assign n33877 = \core_dag_ilm1reg_L2_we_DO_reg[10]/NET0131  & n33107 ;
  assign n33880 = ~n33876 & ~n33877 ;
  assign n33878 = \core_dag_ilm1reg_L3_we_DO_reg[10]/NET0131  & n33101 ;
  assign n33879 = \core_dag_ilm1reg_L0_we_DO_reg[10]/NET0131  & n33103 ;
  assign n33881 = ~n33878 & ~n33879 ;
  assign n33882 = n33880 & n33881 ;
  assign n33883 = ~n21592 & n33882 ;
  assign n33884 = ~n33875 & n33883 ;
  assign n33885 = ~\core_dag_ilm1reg_L_reg[10]/NET0131  & n21592 ;
  assign n33886 = ~n33884 & ~n33885 ;
  assign n33890 = ~n6067 & n33095 ;
  assign n33891 = ~n6075 & n33089 ;
  assign n33894 = ~n33890 & ~n33891 ;
  assign n33892 = ~n6058 & n33091 ;
  assign n33893 = ~n6084 & n33093 ;
  assign n33895 = ~n33892 & ~n33893 ;
  assign n33896 = n33894 & n33895 ;
  assign n33897 = n24062 & ~n33896 ;
  assign n33887 = n24166 & n33091 ;
  assign n33899 = ~n21592 & ~n33887 ;
  assign n33898 = n10402 & n33095 ;
  assign n33888 = n24064 & n33089 ;
  assign n33889 = n10398 & n33093 ;
  assign n33900 = ~n33888 & ~n33889 ;
  assign n33901 = ~n33898 & n33900 ;
  assign n33902 = n33899 & n33901 ;
  assign n33903 = ~n33897 & n33902 ;
  assign n33904 = ~\core_dag_ilm1reg_I_reg[8]/NET0131  & n21592 ;
  assign n33905 = ~n33903 & ~n33904 ;
  assign n33907 = n24068 & ~n33896 ;
  assign n33906 = n10369 & n33091 ;
  assign n33913 = ~n21592 & ~n33906 ;
  assign n33912 = n24149 & n33095 ;
  assign n33908 = n6075 & n33089 ;
  assign n33909 = \core_dag_ilm1reg_I3_we_DO_reg[5]/NET0131  & n33908 ;
  assign n33910 = n6084 & n33093 ;
  assign n33911 = \core_dag_ilm1reg_I2_we_DO_reg[5]/NET0131  & n33910 ;
  assign n33914 = ~n33909 & ~n33911 ;
  assign n33915 = ~n33912 & n33914 ;
  assign n33916 = n33913 & n33915 ;
  assign n33917 = ~n33907 & n33916 ;
  assign n33918 = ~\core_dag_ilm1reg_I_reg[5]/NET0131  & n21592 ;
  assign n33919 = ~n33917 & ~n33918 ;
  assign n33920 = n24074 & ~n33896 ;
  assign n33921 = n8891 & n33095 ;
  assign n33926 = ~n21592 & ~n33921 ;
  assign n33925 = \core_dag_ilm1reg_I3_we_DO_reg[1]/NET0131  & n33908 ;
  assign n33922 = n6058 & n33091 ;
  assign n33923 = \core_dag_ilm1reg_I0_we_DO_reg[1]/NET0131  & n33922 ;
  assign n33924 = \core_dag_ilm1reg_I2_we_DO_reg[1]/NET0131  & n33910 ;
  assign n33927 = ~n33923 & ~n33924 ;
  assign n33928 = ~n33925 & n33927 ;
  assign n33929 = n33926 & n33928 ;
  assign n33930 = ~n33920 & n33929 ;
  assign n33931 = ~\core_dag_ilm1reg_I_reg[1]/NET0131  & n21592 ;
  assign n33932 = ~n33930 & ~n33931 ;
  assign n33936 = n24080 & ~n33896 ;
  assign n33933 = n6136 & n33091 ;
  assign n33939 = ~n21592 & ~n33933 ;
  assign n33937 = n6067 & n33095 ;
  assign n33938 = \core_dag_ilm1reg_I1_we_DO_reg[13]/NET0131  & n33937 ;
  assign n33934 = n24082 & n33089 ;
  assign n33935 = \core_dag_ilm1reg_I2_we_DO_reg[13]/NET0131  & n33910 ;
  assign n33940 = ~n33934 & ~n33935 ;
  assign n33941 = ~n33938 & n33940 ;
  assign n33942 = n33939 & n33941 ;
  assign n33943 = ~n33936 & n33942 ;
  assign n33944 = ~\core_dag_ilm1reg_I_reg[13]/NET0131  & n21592 ;
  assign n33945 = ~n33943 & ~n33944 ;
  assign n33947 = ~n24086 & ~n33896 ;
  assign n33946 = n24134 & n33093 ;
  assign n33951 = ~n21592 & ~n33946 ;
  assign n33950 = \core_dag_ilm1reg_I0_we_DO_reg[12]/NET0131  & n33922 ;
  assign n33948 = \core_dag_ilm1reg_I1_we_DO_reg[12]/NET0131  & n33937 ;
  assign n33949 = n8869 & n33089 ;
  assign n33952 = ~n33948 & ~n33949 ;
  assign n33953 = ~n33950 & n33952 ;
  assign n33954 = n33951 & n33953 ;
  assign n33955 = ~n33947 & n33954 ;
  assign n33956 = ~\core_dag_ilm1reg_I_reg[12]/NET0131  & n21592 ;
  assign n33957 = ~n33955 & ~n33956 ;
  assign n33961 = ~n24091 & ~n33896 ;
  assign n33958 = \core_dag_ilm1reg_I1_we_DO_reg[11]/NET0131  & n33937 ;
  assign n33963 = ~n21592 & ~n33958 ;
  assign n33962 = \core_dag_ilm1reg_I0_we_DO_reg[11]/NET0131  & n33922 ;
  assign n33959 = n8734 & n33093 ;
  assign n33960 = \core_dag_ilm1reg_I3_we_DO_reg[11]/NET0131  & n33908 ;
  assign n33964 = ~n33959 & ~n33960 ;
  assign n33965 = ~n33962 & n33964 ;
  assign n33966 = n33963 & n33965 ;
  assign n33967 = ~n33961 & n33966 ;
  assign n33968 = ~\core_dag_ilm1reg_I_reg[11]/NET0131  & n21592 ;
  assign n33969 = ~n33967 & ~n33968 ;
  assign n33973 = n23763 & ~n33896 ;
  assign n33970 = \core_dag_ilm1reg_I1_we_DO_reg[10]/NET0131  & n33937 ;
  assign n33975 = ~n21592 & ~n33970 ;
  assign n33974 = \core_dag_ilm1reg_I0_we_DO_reg[10]/NET0131  & n33922 ;
  assign n33971 = n8133 & n33093 ;
  assign n33972 = \core_dag_ilm1reg_I3_we_DO_reg[10]/NET0131  & n33908 ;
  assign n33976 = ~n33971 & ~n33972 ;
  assign n33977 = ~n33974 & n33976 ;
  assign n33978 = n33975 & n33977 ;
  assign n33979 = ~n33973 & n33978 ;
  assign n33980 = ~\core_dag_ilm1reg_I_reg[10]/NET0131  & n21592 ;
  assign n33981 = ~n33979 & ~n33980 ;
  assign n33982 = ~\sice_ICYC_reg[16]/NET0131  & ~n20745 ;
  assign n33983 = ~n20746 & ~n33982 ;
  assign n33984 = \core_c_dec_MTSR1_E_reg/P0001  & ~n23920 ;
  assign n33985 = ~\core_c_dec_MTSR1_E_reg/P0001  & n30142 ;
  assign n33986 = ~n33984 & ~n33985 ;
  assign n33987 = n18717 & ~n33986 ;
  assign n33988 = ~\core_eu_es_sht_es_reg_sr1swe_DO_reg[12]/P0001  & ~n18717 ;
  assign n33989 = ~n33987 & ~n33988 ;
  assign n33990 = n17833 & ~n33986 ;
  assign n33991 = ~\core_eu_es_sht_es_reg_sr1rwe_DO_reg[12]/P0001  & ~n17833 ;
  assign n33992 = ~n33990 & ~n33991 ;
  assign n33995 = n18271 & ~n19848 ;
  assign n33994 = ~\core_eu_em_mac_em_reg_mr0swe_DO_reg[10]/P0001  & ~n18271 ;
  assign n33996 = n18273 & ~n33994 ;
  assign n33997 = ~n33995 & n33996 ;
  assign n33993 = \core_eu_em_mac_em_reg_mr0swe_DO_reg[10]/P0001  & ~n18266 ;
  assign n33998 = ~n18270 & ~n33993 ;
  assign n33999 = ~n33997 & n33998 ;
  assign n34000 = ~n18262 & ~n33999 ;
  assign n34001 = n18262 & n19643 ;
  assign n34002 = ~n34000 & ~n34001 ;
  assign n34003 = \sport1_txctl_TXSHT_reg[10]/P0001  & ~n22677 ;
  assign n34004 = \sport1_txctl_TX_reg[11]/P0001  & n22677 ;
  assign n34005 = ~n34003 & ~n34004 ;
  assign n34006 = n14752 & ~n19643 ;
  assign n34007 = n18328 & n19848 ;
  assign n34008 = \core_eu_em_mac_em_reg_mr0rwe_DO_reg[10]/P0001  & ~n18330 ;
  assign n34009 = n18334 & ~n34008 ;
  assign n34010 = ~n34007 & n34009 ;
  assign n34011 = ~n34006 & ~n34010 ;
  assign n34012 = \sport1_rxctl_RCS_reg[1]/NET0131  & ~n31705 ;
  assign n34013 = \sport0_rxctl_RCS_reg[1]/NET0131  & ~n31868 ;
  assign n34014 = \sport0_txctl_TXSHT_reg[10]/P0001  & ~n19960 ;
  assign n34015 = \sport0_txctl_TX_reg[11]/P0001  & n19960 ;
  assign n34016 = ~n34014 & ~n34015 ;
  assign n34017 = ~\sport0_cfg_SCLKi_cnt_reg[6]/NET0131  & ~n19538 ;
  assign n34018 = ~n19544 & ~n34017 ;
  assign n34019 = n19197 & n34018 ;
  assign n34020 = ~\sport0_cfg_SCLKi_cnt_reg[4]/NET0131  & ~n19535 ;
  assign n34021 = ~n19536 & ~n34020 ;
  assign n34022 = n19197 & n34021 ;
  assign n34023 = ~\core_c_dec_MFDAG2_Ei_reg/NET0131  & n4117 ;
  assign n34024 = ~n30936 & n31263 ;
  assign n34027 = \core_c_dec_IR_reg[1]/NET0131  & n34024 ;
  assign n34028 = ~\core_c_dec_IR_reg[2]/NET0131  & n34027 ;
  assign n34029 = ~\core_c_dec_IR_reg[1]/NET0131  & \core_c_dec_IR_reg[2]/NET0131  ;
  assign n34030 = n34024 & n34029 ;
  assign n34031 = ~n34028 & ~n34030 ;
  assign n34032 = n31271 & ~n34031 ;
  assign n34041 = n6091 & ~n31269 ;
  assign n34042 = n34027 & n34041 ;
  assign n34025 = n31265 & n34024 ;
  assign n34026 = n31270 & n34025 ;
  assign n34035 = n32024 & n34025 ;
  assign n34043 = ~n34026 & ~n34035 ;
  assign n34044 = ~n34042 & n34043 ;
  assign n34045 = ~n34032 & n34044 ;
  assign n34033 = n32024 & n34028 ;
  assign n34034 = ~n4117 & ~n34033 ;
  assign n34036 = ~n31653 & n31979 ;
  assign n34037 = n6095 & n19298 ;
  assign n34038 = ~n31269 & n34037 ;
  assign n34039 = ~n34036 & ~n34038 ;
  assign n34040 = n34024 & ~n34039 ;
  assign n34046 = n34034 & ~n34040 ;
  assign n34047 = n34045 & n34046 ;
  assign n34048 = ~n34023 & ~n34047 ;
  assign n34049 = ~\sport1_cfg_SCLKi_cnt_reg[6]/NET0131  & ~n20235 ;
  assign n34050 = ~n20236 & ~n34049 ;
  assign n34051 = n19130 & n34050 ;
  assign n34052 = ~\sport1_cfg_SCLKi_cnt_reg[4]/NET0131  & ~n20233 ;
  assign n34053 = ~n20234 & ~n34052 ;
  assign n34054 = n19130 & n34053 ;
  assign n34055 = \core_c_psq_SSTAT_reg[2]/NET0131  & ~n13778 ;
  assign n34056 = ~n33341 & ~n34055 ;
  assign n34057 = n33337 & n33341 ;
  assign n34058 = ~n34056 & ~n34057 ;
  assign n34059 = \bdma_BCTL_reg[0]/NET0131  & ~n6914 ;
  assign n34060 = ~n5733 & ~n34059 ;
  assign n34061 = n19923 & ~n34060 ;
  assign n34062 = ~\bdma_BCTL_reg[0]/NET0131  & \bdma_BCTL_reg[1]/NET0131  ;
  assign n34063 = ~n34061 & ~n34062 ;
  assign n34064 = ~n5729 & ~n34059 ;
  assign n34065 = ~n13146 & ~n34064 ;
  assign n34066 = n19923 & ~n34065 ;
  assign n34067 = ~n25024 & ~n34066 ;
  assign n34068 = ~n34063 & n34067 ;
  assign n34069 = \bdma_BRdataBUF_reg[0]/P0001  & ~n34068 ;
  assign n34070 = \T_ED[0]_pad  & n34061 ;
  assign n34071 = n34067 & n34070 ;
  assign n34072 = ~n34069 & ~n34071 ;
  assign n34073 = \bdma_BWCOUNT_reg[11]/NET0131  & ~n33295 ;
  assign n34074 = ~n13763 & ~n33296 ;
  assign n34075 = ~n34073 & n34074 ;
  assign n34076 = ~n8460 & n13763 ;
  assign n34077 = ~n34075 & ~n34076 ;
  assign n34079 = \bdma_BIAD_reg[0]/NET0131  & ~n13755 ;
  assign n34080 = \bdma_BIAD_reg[1]/NET0131  & n34079 ;
  assign n34081 = \bdma_BIAD_reg[2]/NET0131  & n34080 ;
  assign n34082 = \bdma_BIAD_reg[3]/NET0131  & n34081 ;
  assign n34083 = \bdma_BIAD_reg[4]/NET0131  & n34082 ;
  assign n34084 = \bdma_BIAD_reg[5]/NET0131  & n34083 ;
  assign n34085 = \bdma_BIAD_reg[6]/NET0131  & n34084 ;
  assign n34086 = \bdma_BIAD_reg[7]/NET0131  & n34085 ;
  assign n34087 = \bdma_BIAD_reg[8]/NET0131  & n34086 ;
  assign n34088 = \bdma_BIAD_reg[9]/NET0131  & n34087 ;
  assign n34089 = \bdma_BIAD_reg[10]/NET0131  & n34088 ;
  assign n34090 = \bdma_BIAD_reg[11]/NET0131  & n34089 ;
  assign n34092 = \bdma_BIAD_reg[12]/NET0131  & n34090 ;
  assign n34078 = n7232 & n20764 ;
  assign n34091 = ~\bdma_BIAD_reg[12]/NET0131  & ~n34090 ;
  assign n34093 = ~n34078 & ~n34091 ;
  assign n34094 = ~n34092 & n34093 ;
  assign n34095 = n9178 & n34078 ;
  assign n34096 = ~n34094 & ~n34095 ;
  assign n34097 = ~\bdma_BIAD_reg[11]/NET0131  & ~n34089 ;
  assign n34098 = ~n34078 & ~n34090 ;
  assign n34099 = ~n34097 & n34098 ;
  assign n34100 = n8460 & n34078 ;
  assign n34101 = ~n34099 & ~n34100 ;
  assign n34102 = \bdma_BEAD_reg[13]/NET0131  & ~n33314 ;
  assign n34103 = ~\bdma_BEAD_reg[13]/NET0131  & n33314 ;
  assign n34104 = ~n34102 & ~n34103 ;
  assign n34105 = ~n20765 & ~n34104 ;
  assign n34106 = n7340 & n20765 ;
  assign n34107 = ~n34105 & ~n34106 ;
  assign n34108 = ~\bdma_BEAD_reg[11]/NET0131  & ~n33312 ;
  assign n34109 = ~n20765 & ~n33313 ;
  assign n34110 = ~n34108 & n34109 ;
  assign n34111 = n8460 & n20765 ;
  assign n34112 = ~n34110 & ~n34111 ;
  assign n34113 = \core_c_dec_MTIMASK_Eg_reg/P0001  & ~n10638 ;
  assign n34117 = \core_c_psq_ststk_sts7x23_STcell_reg[6][23]/P0001  & n14711 ;
  assign n34118 = \core_c_psq_ststk_sts7x23_STcell_reg[2][23]/P0001  & n14713 ;
  assign n34123 = ~n34117 & ~n34118 ;
  assign n34119 = \core_c_psq_ststk_sts7x23_STcell_reg[0][23]/P0001  & n14702 ;
  assign n34120 = \core_c_psq_ststk_sts7x23_STcell_reg[1][23]/P0001  & n14708 ;
  assign n34124 = ~n34119 & ~n34120 ;
  assign n34125 = n34123 & n34124 ;
  assign n34114 = \core_c_psq_ststk_sts7x23_STcell_reg[3][23]/P0001  & n14704 ;
  assign n34121 = ~\core_c_dec_MTIMASK_Eg_reg/P0001  & ~n34114 ;
  assign n34115 = \core_c_psq_ststk_sts7x23_STcell_reg[5][23]/P0001  & n14699 ;
  assign n34116 = \core_c_psq_ststk_sts7x23_STcell_reg[4][23]/P0001  & n14706 ;
  assign n34122 = ~n34115 & ~n34116 ;
  assign n34126 = n34121 & n34122 ;
  assign n34127 = n34125 & n34126 ;
  assign n34128 = ~n34113 & ~n34127 ;
  assign n34129 = n32367 & n34128 ;
  assign n34130 = \core_c_psq_ICNTL_reg_DO_reg[4]/NET0131  & ~n33494 ;
  assign n34131 = n32364 & ~n34130 ;
  assign n34132 = \core_c_psq_IMASK_reg[8]/NET0131  & ~n34131 ;
  assign n34133 = ~n32367 & n34132 ;
  assign n34134 = ~n34129 & ~n34133 ;
  assign n34135 = \bdma_BRdataBUF_reg[5]/P0001  & ~n34068 ;
  assign n34136 = \T_ED[5]_pad  & ~n25024 ;
  assign n34137 = n34061 & n34136 ;
  assign n34138 = ~n34135 & ~n34137 ;
  assign n34139 = \bdma_BRdataBUF_reg[7]/P0001  & ~n34068 ;
  assign n34140 = \T_ED[7]_pad  & ~n25024 ;
  assign n34141 = n34061 & n34140 ;
  assign n34142 = ~n34139 & ~n34141 ;
  assign n34143 = \bdma_BRdataBUF_reg[4]/P0001  & ~n34068 ;
  assign n34144 = \T_ED[4]_pad  & ~n25024 ;
  assign n34145 = n34061 & n34144 ;
  assign n34146 = ~n34143 & ~n34145 ;
  assign n34147 = \bdma_BRdataBUF_reg[6]/P0001  & ~n34068 ;
  assign n34148 = \T_ED[6]_pad  & ~n25024 ;
  assign n34149 = n34061 & n34148 ;
  assign n34150 = ~n34147 & ~n34149 ;
  assign n34151 = \bdma_BRdataBUF_reg[3]/P0001  & ~n34068 ;
  assign n34152 = \T_ED[3]_pad  & ~n25024 ;
  assign n34153 = n34061 & n34152 ;
  assign n34154 = ~n34151 & ~n34153 ;
  assign n34155 = \bdma_BRdataBUF_reg[2]/P0001  & ~n34068 ;
  assign n34156 = \T_ED[2]_pad  & ~n25024 ;
  assign n34157 = n34061 & n34156 ;
  assign n34158 = ~n34155 & ~n34157 ;
  assign n34159 = \bdma_BRdataBUF_reg[1]/P0001  & ~n34068 ;
  assign n34160 = \T_ED[1]_pad  & ~n25024 ;
  assign n34161 = n34061 & n34160 ;
  assign n34162 = ~n34159 & ~n34161 ;
  assign n34163 = ~\sice_ICYC_reg[20]/NET0131  & ~n20749 ;
  assign n34164 = ~n20750 & ~n34163 ;
  assign n34165 = \sice_IIRC_reg[21]/NET0131  & n32042 ;
  assign n34166 = \sice_IIRC_reg[22]/NET0131  & n34165 ;
  assign n34167 = ~\sice_IIRC_reg[23]/NET0131  & ~n34166 ;
  assign n34168 = \sice_IIRC_reg[23]/NET0131  & n34166 ;
  assign n34169 = ~n34167 & ~n34168 ;
  assign n34170 = ~\clkc_oscntr_reg_DO_reg[10]/NET0131  & ~n23424 ;
  assign n34171 = ~n33617 & ~n34170 ;
  assign n34172 = \core_c_dec_MTIMASK_Eg_reg/P0001  & ~n11265 ;
  assign n34176 = \core_c_psq_ststk_sts7x23_STcell_reg[2][22]/P0001  & n14713 ;
  assign n34177 = \core_c_psq_ststk_sts7x23_STcell_reg[6][22]/P0001  & n14711 ;
  assign n34182 = ~n34176 & ~n34177 ;
  assign n34178 = \core_c_psq_ststk_sts7x23_STcell_reg[1][22]/P0001  & n14708 ;
  assign n34179 = \core_c_psq_ststk_sts7x23_STcell_reg[5][22]/P0001  & n14699 ;
  assign n34183 = ~n34178 & ~n34179 ;
  assign n34184 = n34182 & n34183 ;
  assign n34173 = \core_c_psq_ststk_sts7x23_STcell_reg[4][22]/P0001  & n14706 ;
  assign n34180 = ~\core_c_dec_MTIMASK_Eg_reg/P0001  & ~n34173 ;
  assign n34174 = \core_c_psq_ststk_sts7x23_STcell_reg[3][22]/P0001  & n14704 ;
  assign n34175 = \core_c_psq_ststk_sts7x23_STcell_reg[0][22]/P0001  & n14702 ;
  assign n34181 = ~n34174 & ~n34175 ;
  assign n34185 = n34180 & n34181 ;
  assign n34186 = n34184 & n34185 ;
  assign n34187 = ~n34172 & ~n34186 ;
  assign n34188 = n32367 & n34187 ;
  assign n34189 = \core_c_psq_ICNTL_reg_DO_reg[4]/NET0131  & ~n33493 ;
  assign n34190 = n32364 & ~n34189 ;
  assign n34191 = \core_c_psq_IMASK_reg[7]/NET0131  & ~n34190 ;
  assign n34192 = ~n32367 & n34191 ;
  assign n34193 = ~n34188 & ~n34192 ;
  assign n34194 = \core_c_dec_MTIMASK_Eg_reg/P0001  & ~n8715 ;
  assign n34198 = \core_c_psq_ststk_sts7x23_STcell_reg[2][17]/P0001  & n14713 ;
  assign n34199 = \core_c_psq_ststk_sts7x23_STcell_reg[6][17]/P0001  & n14711 ;
  assign n34204 = ~n34198 & ~n34199 ;
  assign n34200 = \core_c_psq_ststk_sts7x23_STcell_reg[1][17]/P0001  & n14708 ;
  assign n34201 = \core_c_psq_ststk_sts7x23_STcell_reg[5][17]/P0001  & n14699 ;
  assign n34205 = ~n34200 & ~n34201 ;
  assign n34206 = n34204 & n34205 ;
  assign n34195 = \core_c_psq_ststk_sts7x23_STcell_reg[4][17]/P0001  & n14706 ;
  assign n34202 = ~\core_c_dec_MTIMASK_Eg_reg/P0001  & ~n34195 ;
  assign n34196 = \core_c_psq_ststk_sts7x23_STcell_reg[3][17]/P0001  & n14704 ;
  assign n34197 = \core_c_psq_ststk_sts7x23_STcell_reg[0][17]/P0001  & n14702 ;
  assign n34203 = ~n34196 & ~n34197 ;
  assign n34207 = n34202 & n34203 ;
  assign n34208 = n34206 & n34207 ;
  assign n34209 = ~n34194 & ~n34208 ;
  assign n34210 = n32367 & n34209 ;
  assign n34211 = \core_c_psq_ICNTL_reg_DO_reg[4]/NET0131  & ~n5299 ;
  assign n34212 = n32364 & ~n34211 ;
  assign n34213 = \core_c_psq_IMASK_reg[2]/NET0131  & ~n34212 ;
  assign n34214 = ~n32367 & n34213 ;
  assign n34215 = ~n34210 & ~n34214 ;
  assign n34216 = ~\clkc_oscntr_reg_DO_reg[8]/NET0131  & ~n23421 ;
  assign n34217 = ~n23422 & ~n34216 ;
  assign n34218 = \core_c_dec_MTIMASK_Eg_reg/P0001  & ~n10069 ;
  assign n34222 = \core_c_psq_ststk_sts7x23_STcell_reg[2][19]/P0001  & n14713 ;
  assign n34223 = \core_c_psq_ststk_sts7x23_STcell_reg[6][19]/P0001  & n14711 ;
  assign n34228 = ~n34222 & ~n34223 ;
  assign n34224 = \core_c_psq_ststk_sts7x23_STcell_reg[1][19]/P0001  & n14708 ;
  assign n34225 = \core_c_psq_ststk_sts7x23_STcell_reg[5][19]/P0001  & n14699 ;
  assign n34229 = ~n34224 & ~n34225 ;
  assign n34230 = n34228 & n34229 ;
  assign n34219 = \core_c_psq_ststk_sts7x23_STcell_reg[4][19]/P0001  & n14706 ;
  assign n34226 = ~\core_c_dec_MTIMASK_Eg_reg/P0001  & ~n34219 ;
  assign n34220 = \core_c_psq_ststk_sts7x23_STcell_reg[3][19]/P0001  & n14704 ;
  assign n34221 = \core_c_psq_ststk_sts7x23_STcell_reg[0][19]/P0001  & n14702 ;
  assign n34227 = ~n34220 & ~n34221 ;
  assign n34231 = n34226 & n34227 ;
  assign n34232 = n34230 & n34231 ;
  assign n34233 = ~n34218 & ~n34232 ;
  assign n34234 = n32367 & n34233 ;
  assign n34235 = \core_c_psq_ICNTL_reg_DO_reg[4]/NET0131  & ~n33244 ;
  assign n34236 = n32364 & ~n34235 ;
  assign n34237 = \core_c_psq_IMASK_reg[4]/NET0131  & ~n34236 ;
  assign n34238 = ~n32367 & n34237 ;
  assign n34239 = ~n34234 & ~n34238 ;
  assign n34240 = \sport0_regs_FSDIVreg_DO_reg[3]/NET0131  & n28876 ;
  assign n34241 = ~\sport0_cfg_FSi_cnt_reg[3]/NET0131  & ~n28948 ;
  assign n34242 = ~n28949 & ~n34241 ;
  assign n34243 = n28945 & n34242 ;
  assign n34244 = ~n34240 & ~n34243 ;
  assign n34245 = ~\sice_ICYC_reg[12]/NET0131  & ~n20741 ;
  assign n34246 = ~n20742 & ~n34245 ;
  assign n34247 = \sport1_regs_FSDIVreg_DO_reg[3]/NET0131  & n28786 ;
  assign n34248 = ~\sport1_cfg_FSi_cnt_reg[3]/NET0131  & ~n28858 ;
  assign n34249 = ~n28859 & ~n34248 ;
  assign n34250 = n28855 & n34249 ;
  assign n34251 = ~n34247 & ~n34250 ;
  assign n34252 = ~\sice_IIRC_reg[12]/NET0131  & ~n20856 ;
  assign n34253 = ~n20857 & ~n34252 ;
  assign n34254 = ~\core_c_dec_Dummy_E_reg/NET0131  & \core_c_dec_MTSB_E_reg/P0001  ;
  assign n34260 = ~n9268 & ~n26276 ;
  assign n34261 = n7365 & ~n34260 ;
  assign n34262 = ~n23671 & n34261 ;
  assign n34259 = n9268 & n26276 ;
  assign n34263 = n8489 & n27488 ;
  assign n34264 = ~n34259 & ~n34263 ;
  assign n34265 = ~n34262 & n34264 ;
  assign n34266 = ~n7983 & ~n29493 ;
  assign n34267 = ~n8489 & ~n27488 ;
  assign n34268 = ~n34266 & ~n34267 ;
  assign n34269 = ~n34265 & n34268 ;
  assign n34257 = ~n7168 & n29480 ;
  assign n34258 = n7983 & n29493 ;
  assign n34270 = ~n34257 & ~n34258 ;
  assign n34271 = ~n34269 & n34270 ;
  assign n34256 = n7168 & ~n29480 ;
  assign n34255 = \core_c_dec_IRE_reg[11]/NET0131  & \core_c_dec_IRE_reg[12]/NET0131  ;
  assign n34272 = n23585 & n34255 ;
  assign n34273 = n13803 & n34272 ;
  assign n34274 = ~n34256 & n34273 ;
  assign n34275 = ~n34271 & n34274 ;
  assign n34276 = ~n34254 & ~n34275 ;
  assign n34277 = n14664 & ~n34276 ;
  assign n34278 = \core_c_dec_MTSB_E_reg/P0001  & ~n9435 ;
  assign n34279 = ~\core_c_dec_MTSB_E_reg/P0001  & ~n26276 ;
  assign n34280 = ~n34278 & ~n34279 ;
  assign n34281 = n34277 & ~n34280 ;
  assign n34282 = ~\core_eu_es_sht_es_reg_SBs_reg[1]/P0001  & ~n34277 ;
  assign n34283 = ~n34281 & ~n34282 ;
  assign n34284 = \core_c_dec_MTSB_E_reg/P0001  & ~n7607 ;
  assign n34285 = ~\core_c_dec_MTSB_E_reg/P0001  & n23671 ;
  assign n34286 = ~n34284 & ~n34285 ;
  assign n34287 = n34277 & ~n34286 ;
  assign n34288 = ~\core_eu_es_sht_es_reg_SBs_reg[0]/P0001  & ~n34277 ;
  assign n34289 = ~n34287 & ~n34288 ;
  assign n34290 = \core_c_dec_MTSB_E_reg/P0001  & ~n8113 ;
  assign n34291 = ~\core_c_dec_MTSB_E_reg/P0001  & ~n29493 ;
  assign n34292 = ~n34290 & ~n34291 ;
  assign n34293 = n34277 & ~n34292 ;
  assign n34294 = ~\core_eu_es_sht_es_reg_SBs_reg[3]/P0001  & ~n34277 ;
  assign n34295 = ~n34293 & ~n34294 ;
  assign n34296 = n13801 & ~n34276 ;
  assign n34297 = ~n34292 & n34296 ;
  assign n34298 = ~\core_eu_es_sht_es_reg_SBr_reg[3]/P0001  & ~n34296 ;
  assign n34299 = ~n34297 & ~n34298 ;
  assign n34300 = \core_c_dec_MTSB_E_reg/P0001  & ~n8715 ;
  assign n34301 = ~\core_c_dec_MTSB_E_reg/P0001  & ~n27488 ;
  assign n34302 = ~n34300 & ~n34301 ;
  assign n34303 = n34277 & ~n34302 ;
  assign n34304 = ~\core_eu_es_sht_es_reg_SBs_reg[2]/P0001  & ~n34277 ;
  assign n34305 = ~n34303 & ~n34304 ;
  assign n34306 = n34296 & ~n34302 ;
  assign n34307 = ~\core_eu_es_sht_es_reg_SBr_reg[2]/P0001  & ~n34296 ;
  assign n34308 = ~n34306 & ~n34307 ;
  assign n34309 = \core_c_dec_MTSB_E_reg/P0001  & ~n10069 ;
  assign n34310 = ~\core_c_dec_MTSB_E_reg/P0001  & n29480 ;
  assign n34311 = ~n34309 & ~n34310 ;
  assign n34312 = n34296 & ~n34311 ;
  assign n34313 = ~\core_eu_es_sht_es_reg_SBr_reg[4]/P0001  & ~n34296 ;
  assign n34314 = ~n34312 & ~n34313 ;
  assign n34315 = ~n34280 & n34296 ;
  assign n34316 = ~\core_eu_es_sht_es_reg_SBr_reg[1]/P0001  & ~n34296 ;
  assign n34317 = ~n34315 & ~n34316 ;
  assign n34318 = n34277 & ~n34311 ;
  assign n34319 = ~\core_eu_es_sht_es_reg_SBs_reg[4]/P0001  & ~n34277 ;
  assign n34320 = ~n34318 & ~n34319 ;
  assign n34321 = ~n34286 & n34296 ;
  assign n34322 = ~\core_eu_es_sht_es_reg_SBr_reg[0]/P0001  & ~n34296 ;
  assign n34323 = ~n34321 & ~n34322 ;
  assign n34326 = n18271 & ~n19504 ;
  assign n34325 = ~\core_eu_em_mac_em_reg_mr0swe_DO_reg[9]/P0001  & ~n18271 ;
  assign n34327 = n18273 & ~n34325 ;
  assign n34328 = ~n34326 & n34327 ;
  assign n34324 = \core_eu_em_mac_em_reg_mr0swe_DO_reg[9]/P0001  & ~n18266 ;
  assign n34329 = ~n18270 & ~n34324 ;
  assign n34330 = ~n34328 & n34329 ;
  assign n34331 = ~n18262 & ~n34330 ;
  assign n34332 = n18262 & ~n19646 ;
  assign n34333 = ~n34331 & ~n34332 ;
  assign n34334 = n14752 & n19646 ;
  assign n34335 = n18328 & n19504 ;
  assign n34336 = \core_eu_em_mac_em_reg_mr0rwe_DO_reg[9]/P0001  & ~n18330 ;
  assign n34337 = n18334 & ~n34336 ;
  assign n34338 = ~n34335 & n34337 ;
  assign n34339 = ~n34334 & ~n34338 ;
  assign n34342 = \sport0_rxctl_RX_reg[4]/P0001  & ~n20914 ;
  assign n34343 = \sport0_rxctl_RX_reg[2]/P0001  & ~\sport0_rxctl_RX_reg[4]/P0001  ;
  assign n34344 = ~n20878 & ~n34343 ;
  assign n34345 = ~n34342 & n34344 ;
  assign n34346 = ~n20905 & ~n34345 ;
  assign n34347 = ~\sport0_rxctl_RX_reg[6]/P0001  & ~n34346 ;
  assign n34348 = \sport0_rxctl_RX_reg[0]/P0001  & ~\sport0_rxctl_RX_reg[6]/P0001  ;
  assign n34349 = n31045 & ~n34348 ;
  assign n34350 = ~n34347 & ~n34349 ;
  assign n34351 = n20882 & ~n34350 ;
  assign n34352 = ~n20882 & n31037 ;
  assign n34353 = ~n34351 & ~n34352 ;
  assign n34354 = n31031 & n34353 ;
  assign n34355 = ~n20925 & ~n20926 ;
  assign n34356 = ~\sport0_rxctl_RX_reg[4]/P0001  & ~n34355 ;
  assign n34357 = ~\sport0_rxctl_RX_reg[6]/P0001  & ~n20931 ;
  assign n34358 = ~n34356 & n34357 ;
  assign n34359 = n20882 & ~n34358 ;
  assign n34360 = ~n20882 & n34350 ;
  assign n34361 = ~n34359 & ~n34360 ;
  assign n34362 = ~n34354 & n34361 ;
  assign n34363 = n34354 & ~n34361 ;
  assign n34364 = ~n34362 & ~n34363 ;
  assign n34365 = n31043 & n34353 ;
  assign n34366 = ~\sport0_rxctl_RX_reg[7]/P0001  & ~n34365 ;
  assign n34368 = n34364 & ~n34366 ;
  assign n34367 = ~n34364 & n34366 ;
  assign n34369 = n20875 & ~n34367 ;
  assign n34370 = ~n34368 & n34369 ;
  assign n34371 = ~\sport0_rxctl_ldRX_cmp_reg/P0001  & n10638 ;
  assign n34341 = \sport0_rxctl_RX_reg[8]/P0001  & n20873 ;
  assign n34372 = ~n20868 & ~n34341 ;
  assign n34373 = ~n34371 & n34372 ;
  assign n34374 = ~n34370 & n34373 ;
  assign n34340 = ~\sport0_rxctl_RXSHT_reg[8]/P0001  & n20868 ;
  assign n34375 = ~n20871 & ~n34340 ;
  assign n34376 = ~n34374 & n34375 ;
  assign n34377 = \sport0_rxctl_RX_reg[8]/P0001  & n20871 ;
  assign n34378 = ~n34376 & ~n34377 ;
  assign n34379 = ~n17796 & n18262 ;
  assign n34380 = ~\core_eu_em_mac_em_reg_mr2swe_DO_reg[2]/P0001  & ~n28530 ;
  assign n34381 = n17814 & ~n19381 ;
  assign n34382 = n28534 & ~n34381 ;
  assign n34383 = ~n34380 & ~n34382 ;
  assign n34384 = ~n19385 & ~n34383 ;
  assign n34385 = ~\core_eu_em_mac_em_reg_mr2swe_DO_reg[2]/P0001  & ~n28532 ;
  assign n34386 = ~n34384 & ~n34385 ;
  assign n34387 = n28529 & ~n34386 ;
  assign n34388 = ~n34379 & ~n34387 ;
  assign n34391 = ~n20882 & n34358 ;
  assign n34392 = \sport0_rxctl_RX_reg[2]/P0001  & n31045 ;
  assign n34393 = ~\sport0_rxctl_RX_reg[6]/P0001  & ~n20961 ;
  assign n34394 = ~n34392 & n34393 ;
  assign n34395 = n20882 & n34394 ;
  assign n34396 = ~n34391 & ~n34395 ;
  assign n34397 = n34363 & n34396 ;
  assign n34398 = n34364 & n34365 ;
  assign n34399 = ~\sport0_rxctl_RX_reg[7]/P0001  & ~n34398 ;
  assign n34400 = ~n20882 & n34394 ;
  assign n34401 = ~\sport0_rxctl_RX_reg[6]/P0001  & n31033 ;
  assign n34402 = \sport0_regs_SCTLreg_DO_reg[4]/NET0131  & n34401 ;
  assign n34403 = ~n34400 & ~n34402 ;
  assign n34404 = n34399 & ~n34403 ;
  assign n34405 = ~n34399 & n34403 ;
  assign n34406 = ~n34404 & ~n34405 ;
  assign n34408 = ~n34397 & ~n34406 ;
  assign n34407 = n34397 & n34406 ;
  assign n34409 = n20875 & ~n34407 ;
  assign n34410 = ~n34408 & n34409 ;
  assign n34411 = ~\sport0_rxctl_ldRX_cmp_reg/P0001  & n7859 ;
  assign n34390 = \sport0_rxctl_RX_reg[10]/P0001  & n20873 ;
  assign n34412 = ~n20868 & ~n34390 ;
  assign n34413 = ~n34411 & n34412 ;
  assign n34414 = ~n34410 & n34413 ;
  assign n34389 = ~\sport0_rxctl_RXSHT_reg[10]/P0001  & n20868 ;
  assign n34415 = ~n20871 & ~n34389 ;
  assign n34416 = ~n34414 & n34415 ;
  assign n34417 = \sport0_rxctl_RX_reg[10]/P0001  & n20871 ;
  assign n34418 = ~n34416 & ~n34417 ;
  assign n34420 = ~\idma_DCTL_reg[11]/NET0131  & ~\idma_DCTL_reg[12]/NET0131  ;
  assign n34421 = ~\idma_DCTL_reg[13]/NET0131  & ~\idma_DCTL_reg[1]/NET0131  ;
  assign n34428 = n34420 & n34421 ;
  assign n34419 = ~\idma_DCTL_reg[0]/NET0131  & ~\idma_DCTL_reg[10]/NET0131  ;
  assign n34429 = n20386 & n34419 ;
  assign n34430 = n34428 & n34429 ;
  assign n34424 = ~\idma_DCTL_reg[6]/NET0131  & ~\idma_DCTL_reg[7]/NET0131  ;
  assign n34425 = ~\idma_DCTL_reg[8]/NET0131  & ~\idma_DCTL_reg[9]/NET0131  ;
  assign n34426 = n34424 & n34425 ;
  assign n34422 = ~\idma_DCTL_reg[2]/NET0131  & ~\idma_DCTL_reg[3]/NET0131  ;
  assign n34423 = ~\idma_DCTL_reg[4]/NET0131  & ~\idma_DCTL_reg[5]/NET0131  ;
  assign n34427 = n34422 & n34423 ;
  assign n34431 = n34426 & n34427 ;
  assign n34432 = n34430 & n34431 ;
  assign n34433 = n32464 & n34432 ;
  assign n34434 = ~n4060 & ~n34433 ;
  assign n34435 = ~\clkc_OUTcnt_reg[4]/NET0131  & ~n19470 ;
  assign n34436 = ~n19471 & ~n34435 ;
  assign n34437 = ~n19467 & n34436 ;
  assign n34438 = ~\clkc_STDcnt_reg[4]/NET0131  & ~n31524 ;
  assign n34439 = ~n31525 & ~n34438 ;
  assign n34440 = ~n31521 & n34439 ;
  assign n34458 = ~\core_c_psq_IMASK_reg[0]/NET0131  & ~n32366 ;
  assign n34441 = \core_c_dec_MTIMASK_Eg_reg/P0001  & ~n7607 ;
  assign n34445 = \core_c_psq_ststk_sts7x23_STcell_reg[6][15]/P0001  & n14711 ;
  assign n34446 = \core_c_psq_ststk_sts7x23_STcell_reg[2][15]/P0001  & n14713 ;
  assign n34451 = ~n34445 & ~n34446 ;
  assign n34447 = \core_c_psq_ststk_sts7x23_STcell_reg[0][15]/P0001  & n14702 ;
  assign n34448 = \core_c_psq_ststk_sts7x23_STcell_reg[1][15]/P0001  & n14708 ;
  assign n34452 = ~n34447 & ~n34448 ;
  assign n34453 = n34451 & n34452 ;
  assign n34442 = \core_c_psq_ststk_sts7x23_STcell_reg[3][15]/P0001  & n14704 ;
  assign n34449 = ~\core_c_dec_MTIMASK_Eg_reg/P0001  & ~n34442 ;
  assign n34443 = \core_c_psq_ststk_sts7x23_STcell_reg[5][15]/P0001  & n14699 ;
  assign n34444 = \core_c_psq_ststk_sts7x23_STcell_reg[4][15]/P0001  & n14706 ;
  assign n34450 = ~n34443 & ~n34444 ;
  assign n34454 = n34449 & n34450 ;
  assign n34455 = n34453 & n34454 ;
  assign n34456 = ~n34441 & ~n34455 ;
  assign n34457 = n32366 & ~n34456 ;
  assign n34459 = ~n32364 & ~n34457 ;
  assign n34460 = ~n34458 & n34459 ;
  assign n34461 = \core_c_dec_MTTX1_E_reg/P0001  & n4117 ;
  assign n34462 = n31995 & ~n31998 ;
  assign n34463 = ~n4117 & ~n32007 ;
  assign n34464 = ~n32003 & n34463 ;
  assign n34465 = n34462 & n34464 ;
  assign n34466 = n32018 & n34465 ;
  assign n34467 = ~n34461 & ~n34466 ;
  assign n34468 = n4116 & ~n34467 ;
  assign n34469 = \core_c_dec_MTTX0_E_reg/P0001  & n4117 ;
  assign n34470 = n32014 & n34464 ;
  assign n34471 = n32018 & n34470 ;
  assign n34472 = ~n34469 & ~n34471 ;
  assign n34473 = n4116 & ~n34472 ;
  assign n34474 = \core_c_dec_MTMreg_E_reg[1]/P0001  & n4117 ;
  assign n34475 = n31992 & ~n32000 ;
  assign n34476 = ~n31995 & n34475 ;
  assign n34477 = n31998 & ~n32007 ;
  assign n34478 = ~n32001 & n32003 ;
  assign n34479 = ~n4117 & n34478 ;
  assign n34480 = n34477 & n34479 ;
  assign n34481 = n34476 & n34480 ;
  assign n34482 = ~n34474 & ~n34481 ;
  assign n34483 = n4116 & ~n34482 ;
  assign n34485 = \sport1_txctl_Bcnt_reg[4]/NET0131  & ~n22674 ;
  assign n34486 = ~n22675 & ~n34485 ;
  assign n34487 = n23265 & n34486 ;
  assign n34484 = ~\sport1_regs_MWORDreg_DO_reg[10]/NET0131  & ~n23265 ;
  assign n34488 = ~\sport1_rxctl_TAG_SLOT_reg/P0001  & ~n34484 ;
  assign n34489 = ~n34487 & n34488 ;
  assign n34491 = \sport0_txctl_Bcnt_reg[4]/NET0131  & ~n19957 ;
  assign n34492 = ~n19958 & ~n34491 ;
  assign n34493 = n23277 & n34492 ;
  assign n34490 = ~\sport0_regs_MWORDreg_DO_reg[10]/NET0131  & ~n23277 ;
  assign n34494 = ~\sport0_rxctl_TAG_SLOT_reg/P0001  & ~n34490 ;
  assign n34495 = ~n34493 & n34494 ;
  assign n34496 = ~n10289 & n13763 ;
  assign n34497 = \bdma_BWCOUNT_reg[9]/NET0131  & ~n33293 ;
  assign n34498 = ~n13763 & ~n33294 ;
  assign n34499 = ~n34497 & n34498 ;
  assign n34500 = ~n34496 & ~n34499 ;
  assign n34501 = ~n10638 & n13763 ;
  assign n34502 = \bdma_BWCOUNT_reg[8]/NET0131  & ~n33292 ;
  assign n34503 = ~n13763 & ~n33293 ;
  assign n34504 = ~n34502 & n34503 ;
  assign n34505 = ~n34501 & ~n34504 ;
  assign n34506 = \bdma_BWCOUNT_reg[12]/NET0131  & ~n33296 ;
  assign n34507 = ~n13763 & ~n33297 ;
  assign n34508 = ~n34506 & n34507 ;
  assign n34509 = ~n9178 & n13763 ;
  assign n34510 = ~n34508 & ~n34509 ;
  assign n34511 = \bdma_BWCOUNT_reg[10]/NET0131  & ~n33294 ;
  assign n34512 = ~n13763 & ~n33295 ;
  assign n34513 = ~n34511 & n34512 ;
  assign n34514 = ~n7859 & n13763 ;
  assign n34515 = ~n34513 & ~n34514 ;
  assign n34516 = ~\bdma_BIAD_reg[9]/NET0131  & ~n34087 ;
  assign n34517 = ~n34078 & ~n34088 ;
  assign n34518 = ~n34516 & n34517 ;
  assign n34519 = n10289 & n34078 ;
  assign n34520 = ~n34518 & ~n34519 ;
  assign n34521 = ~\bdma_BIAD_reg[8]/NET0131  & ~n34086 ;
  assign n34522 = ~n34078 & ~n34087 ;
  assign n34523 = ~n34521 & n34522 ;
  assign n34524 = n10638 & n34078 ;
  assign n34525 = ~n34523 & ~n34524 ;
  assign n34526 = \bdma_BIAD_reg[13]/NET0131  & ~n34092 ;
  assign n34527 = ~\bdma_BIAD_reg[13]/NET0131  & n34092 ;
  assign n34528 = ~n34526 & ~n34527 ;
  assign n34529 = ~n34078 & ~n34528 ;
  assign n34530 = n7340 & n34078 ;
  assign n34531 = ~n34529 & ~n34530 ;
  assign n34532 = ~\bdma_BIAD_reg[10]/NET0131  & ~n34088 ;
  assign n34533 = ~n34078 & ~n34089 ;
  assign n34534 = ~n34532 & n34533 ;
  assign n34535 = n7859 & n34078 ;
  assign n34536 = ~n34534 & ~n34535 ;
  assign n34537 = ~\bdma_BEAD_reg[9]/NET0131  & ~n33310 ;
  assign n34538 = ~n20765 & ~n33311 ;
  assign n34539 = ~n34537 & n34538 ;
  assign n34540 = n10289 & n20765 ;
  assign n34541 = ~n34539 & ~n34540 ;
  assign n34542 = ~\bdma_BEAD_reg[8]/NET0131  & ~n33309 ;
  assign n34543 = ~n20765 & ~n33310 ;
  assign n34544 = ~n34542 & n34543 ;
  assign n34545 = n10638 & n20765 ;
  assign n34546 = ~n34544 & ~n34545 ;
  assign n34547 = ~\bdma_BEAD_reg[10]/NET0131  & ~n33311 ;
  assign n34548 = ~n20765 & ~n33312 ;
  assign n34549 = ~n34547 & n34548 ;
  assign n34550 = n7859 & n20765 ;
  assign n34551 = ~n34549 & ~n34550 ;
  assign n34552 = \sport1_txctl_TXSHT_reg[3]/P0001  & ~n22677 ;
  assign n34553 = \sport1_txctl_TX_reg[4]/P0001  & n22677 ;
  assign n34554 = ~n34552 & ~n34553 ;
  assign n34555 = \core_c_dec_MFSPT_Ei_reg/NET0131  & n4117 ;
  assign n34556 = ~\core_c_dec_IR_reg[2]/NET0131  & n31264 ;
  assign n34557 = ~n31269 & n34556 ;
  assign n34558 = n25864 & n34557 ;
  assign n34559 = ~n34555 & ~n34558 ;
  assign n34560 = \bdma_BWCOUNT_reg[7]/NET0131  & ~n33291 ;
  assign n34561 = ~n13763 & ~n33292 ;
  assign n34562 = ~n34560 & n34561 ;
  assign n34563 = ~n11265 & n13763 ;
  assign n34564 = ~n34562 & ~n34563 ;
  assign n34565 = ~n11525 & n13763 ;
  assign n34566 = \bdma_BWCOUNT_reg[6]/NET0131  & ~n13769 ;
  assign n34567 = ~n13763 & ~n33291 ;
  assign n34568 = ~n34566 & n34567 ;
  assign n34569 = ~n34565 & ~n34568 ;
  assign n34570 = \sport0_txctl_TXSHT_reg[3]/P0001  & ~n19960 ;
  assign n34571 = \sport0_txctl_TX_reg[4]/P0001  & n19960 ;
  assign n34572 = ~n34570 & ~n34571 ;
  assign n34573 = ~\bdma_BWCOUNT_reg[3]/NET0131  & n13766 ;
  assign n34574 = \bdma_BWCOUNT_reg[4]/NET0131  & ~n34573 ;
  assign n34575 = ~n13763 & ~n13767 ;
  assign n34576 = ~n34574 & n34575 ;
  assign n34577 = ~n10069 & n13763 ;
  assign n34578 = ~n34576 & ~n34577 ;
  assign n34579 = \bdma_BWCOUNT_reg[3]/NET0131  & ~n13766 ;
  assign n34580 = ~n13763 & ~n34573 ;
  assign n34581 = ~n34579 & n34580 ;
  assign n34582 = ~n8113 & n13763 ;
  assign n34583 = ~n34581 & ~n34582 ;
  assign n34584 = \bdma_BWCOUNT_reg[2]/NET0131  & ~n13765 ;
  assign n34585 = ~n13763 & ~n13766 ;
  assign n34586 = ~n34584 & n34585 ;
  assign n34587 = ~n8715 & n13763 ;
  assign n34588 = ~n34586 & ~n34587 ;
  assign n34589 = \bdma_BWCOUNT_reg[0]/NET0131  & n13755 ;
  assign n34590 = ~n13763 & ~n13764 ;
  assign n34591 = ~n34589 & n34590 ;
  assign n34592 = ~n7607 & n13763 ;
  assign n34593 = ~n34591 & ~n34592 ;
  assign n34594 = ~\bdma_BIAD_reg[6]/NET0131  & ~n34084 ;
  assign n34595 = ~n34078 & ~n34085 ;
  assign n34596 = ~n34594 & n34595 ;
  assign n34597 = n11525 & n34078 ;
  assign n34598 = ~n34596 & ~n34597 ;
  assign n34599 = ~\bdma_BIAD_reg[7]/NET0131  & ~n34085 ;
  assign n34600 = ~n34078 & ~n34086 ;
  assign n34601 = ~n34599 & n34600 ;
  assign n34602 = n11265 & n34078 ;
  assign n34603 = ~n34601 & ~n34602 ;
  assign n34604 = ~\bdma_BIAD_reg[5]/NET0131  & ~n34083 ;
  assign n34605 = ~n34078 & ~n34084 ;
  assign n34606 = ~n34604 & n34605 ;
  assign n34607 = n10911 & n34078 ;
  assign n34608 = ~n34606 & ~n34607 ;
  assign n34609 = ~\bdma_BIAD_reg[4]/NET0131  & ~n34082 ;
  assign n34610 = ~n34078 & ~n34083 ;
  assign n34611 = ~n34609 & n34610 ;
  assign n34612 = n10069 & n34078 ;
  assign n34613 = ~n34611 & ~n34612 ;
  assign n34614 = ~\bdma_BIAD_reg[3]/NET0131  & ~n34081 ;
  assign n34615 = ~n34078 & ~n34082 ;
  assign n34616 = ~n34614 & n34615 ;
  assign n34617 = n8113 & n34078 ;
  assign n34618 = ~n34616 & ~n34617 ;
  assign n34619 = ~\bdma_BIAD_reg[2]/NET0131  & ~n34080 ;
  assign n34620 = ~n34078 & ~n34081 ;
  assign n34621 = ~n34619 & n34620 ;
  assign n34622 = n8715 & n34078 ;
  assign n34623 = ~n34621 & ~n34622 ;
  assign n34624 = ~\bdma_BIAD_reg[1]/NET0131  & ~n34079 ;
  assign n34625 = ~n34078 & ~n34080 ;
  assign n34626 = ~n34624 & n34625 ;
  assign n34627 = n9435 & n34078 ;
  assign n34628 = ~n34626 & ~n34627 ;
  assign n34629 = ~\bdma_BIAD_reg[0]/NET0131  & n13755 ;
  assign n34630 = ~n34078 & ~n34079 ;
  assign n34631 = ~n34629 & n34630 ;
  assign n34632 = n7607 & n34078 ;
  assign n34633 = ~n34631 & ~n34632 ;
  assign n34634 = n18868 & n32038 ;
  assign n34635 = ~\sice_IIRC_reg[5]/NET0131  & ~n34634 ;
  assign n34636 = n18869 & n32038 ;
  assign n34637 = ~n34635 & ~n34636 ;
  assign n34638 = \sice_IIRC_reg[0]/NET0131  & ~n32038 ;
  assign n34639 = ~\sice_IIRC_reg[0]/NET0131  & n32038 ;
  assign n34640 = ~n34638 & ~n34639 ;
  assign n34641 = ~\sice_IIRC_reg[18]/NET0131  & ~n32039 ;
  assign n34642 = ~n32040 & ~n34641 ;
  assign n34643 = ~\sice_IIRC_reg[19]/NET0131  & ~n32040 ;
  assign n34644 = ~n32041 & ~n34643 ;
  assign n34645 = ~\sice_IIRC_reg[21]/NET0131  & ~n32042 ;
  assign n34646 = ~n34165 & ~n34645 ;
  assign n34647 = ~\sice_IIRC_reg[22]/NET0131  & ~n34165 ;
  assign n34648 = ~n34166 & ~n34647 ;
  assign n34649 = ~\clkc_oscntr_reg_DO_reg[7]/NET0131  & ~n23420 ;
  assign n34650 = ~n23421 & ~n34649 ;
  assign n34651 = n7340 & ~n32992 ;
  assign n34652 = \core_dag_ilm2reg_L5_we_DO_reg[13]/NET0131  & n33000 ;
  assign n34656 = ~n21579 & ~n34652 ;
  assign n34655 = \core_dag_ilm2reg_L7_we_DO_reg[13]/NET0131  & n32998 ;
  assign n34653 = \core_dag_ilm2reg_L6_we_DO_reg[13]/NET0131  & n32994 ;
  assign n34654 = \core_dag_ilm2reg_L4_we_DO_reg[13]/NET0131  & n32996 ;
  assign n34657 = ~n34653 & ~n34654 ;
  assign n34658 = ~n34655 & n34657 ;
  assign n34659 = n34656 & n34658 ;
  assign n34660 = ~n34651 & n34659 ;
  assign n34661 = ~\core_dag_ilm2reg_L_reg[13]/NET0131  & n21579 ;
  assign n34662 = ~n34660 & ~n34661 ;
  assign n34663 = n7859 & ~n32992 ;
  assign n34664 = \core_dag_ilm2reg_L5_we_DO_reg[10]/NET0131  & n33000 ;
  assign n34668 = ~n21579 & ~n34664 ;
  assign n34667 = \core_dag_ilm2reg_L7_we_DO_reg[10]/NET0131  & n32998 ;
  assign n34665 = \core_dag_ilm2reg_L6_we_DO_reg[10]/NET0131  & n32994 ;
  assign n34666 = \core_dag_ilm2reg_L4_we_DO_reg[10]/NET0131  & n32996 ;
  assign n34669 = ~n34665 & ~n34666 ;
  assign n34670 = ~n34667 & n34669 ;
  assign n34671 = n34668 & n34670 ;
  assign n34672 = ~n34663 & n34671 ;
  assign n34673 = ~\core_dag_ilm2reg_L_reg[10]/NET0131  & n21579 ;
  assign n34674 = ~n34672 & ~n34673 ;
  assign n34679 = n20602 & ~n33698 ;
  assign n34675 = \core_dag_ilm2reg_I6_we_DO_reg[8]/NET0131  & n33684 ;
  assign n34680 = ~n21579 & ~n34675 ;
  assign n34678 = \core_dag_ilm2reg_I5_we_DO_reg[8]/NET0131  & n33688 ;
  assign n34676 = \core_dag_ilm2reg_I7_we_DO_reg[8]/NET0131  & n33686 ;
  assign n34677 = \core_dag_ilm2reg_I4_we_DO_reg[8]/NET0131  & n33690 ;
  assign n34681 = ~n34676 & ~n34677 ;
  assign n34682 = ~n34678 & n34681 ;
  assign n34683 = n34680 & n34682 ;
  assign n34684 = ~n34679 & n34683 ;
  assign n34685 = ~\core_dag_ilm2reg_I_reg[8]/NET0131  & n21579 ;
  assign n34686 = ~n34684 & ~n34685 ;
  assign n34691 = ~n20707 & ~n33698 ;
  assign n34687 = \core_dag_ilm2reg_I6_we_DO_reg[11]/NET0131  & n33684 ;
  assign n34692 = ~n21579 & ~n34687 ;
  assign n34690 = \core_dag_ilm2reg_I5_we_DO_reg[11]/NET0131  & n33688 ;
  assign n34688 = \core_dag_ilm2reg_I7_we_DO_reg[11]/NET0131  & n33686 ;
  assign n34689 = \core_dag_ilm2reg_I4_we_DO_reg[11]/NET0131  & n33690 ;
  assign n34693 = ~n34688 & ~n34689 ;
  assign n34694 = ~n34690 & n34693 ;
  assign n34695 = n34692 & n34694 ;
  assign n34696 = ~n34691 & n34695 ;
  assign n34697 = ~\core_dag_ilm2reg_I_reg[11]/NET0131  & n21579 ;
  assign n34698 = ~n34696 & ~n34697 ;
  assign n34703 = n20718 & ~n33698 ;
  assign n34699 = \core_dag_ilm2reg_I6_we_DO_reg[10]/NET0131  & n33684 ;
  assign n34704 = ~n21579 & ~n34699 ;
  assign n34702 = \core_dag_ilm2reg_I5_we_DO_reg[10]/NET0131  & n33688 ;
  assign n34700 = \core_dag_ilm2reg_I7_we_DO_reg[10]/NET0131  & n33686 ;
  assign n34701 = \core_dag_ilm2reg_I4_we_DO_reg[10]/NET0131  & n33690 ;
  assign n34705 = ~n34700 & ~n34701 ;
  assign n34706 = ~n34702 & n34705 ;
  assign n34707 = n34704 & n34706 ;
  assign n34708 = ~n34703 & n34707 ;
  assign n34709 = ~\core_dag_ilm2reg_I_reg[10]/NET0131  & n21579 ;
  assign n34710 = ~n34708 & ~n34709 ;
  assign n34715 = ~n24098 & ~n33896 ;
  assign n34711 = \core_dag_ilm1reg_I2_we_DO_reg[9]/NET0131  & n33910 ;
  assign n34716 = ~n21592 & ~n34711 ;
  assign n34714 = \core_dag_ilm1reg_I3_we_DO_reg[9]/NET0131  & n33908 ;
  assign n34712 = \core_dag_ilm1reg_I1_we_DO_reg[9]/NET0131  & n33937 ;
  assign n34713 = \core_dag_ilm1reg_I0_we_DO_reg[9]/NET0131  & n33922 ;
  assign n34717 = ~n34712 & ~n34713 ;
  assign n34718 = ~n34714 & n34717 ;
  assign n34719 = n34716 & n34718 ;
  assign n34720 = ~n34715 & n34719 ;
  assign n34721 = ~\core_dag_ilm1reg_I_reg[9]/NET0131  & n21592 ;
  assign n34722 = ~n34720 & ~n34721 ;
  assign n34723 = n10911 & ~n32992 ;
  assign n34724 = \core_dag_ilm2reg_L7_we_DO_reg[5]/NET0131  & n32998 ;
  assign n34728 = ~n21579 & ~n34724 ;
  assign n34727 = \core_dag_ilm2reg_L5_we_DO_reg[5]/NET0131  & n33000 ;
  assign n34725 = \core_dag_ilm2reg_L4_we_DO_reg[5]/NET0131  & n32996 ;
  assign n34726 = \core_dag_ilm2reg_L6_we_DO_reg[5]/NET0131  & n32994 ;
  assign n34729 = ~n34725 & ~n34726 ;
  assign n34730 = ~n34727 & n34729 ;
  assign n34731 = n34728 & n34730 ;
  assign n34732 = ~n34723 & n34731 ;
  assign n34733 = ~\core_dag_ilm2reg_L_reg[5]/NET0131  & n21579 ;
  assign n34734 = ~n34732 & ~n34733 ;
  assign n34739 = n20614 & ~n33698 ;
  assign n34735 = \core_dag_ilm2reg_I6_we_DO_reg[7]/NET0131  & n33684 ;
  assign n34740 = ~n21579 & ~n34735 ;
  assign n34738 = \core_dag_ilm2reg_I4_we_DO_reg[7]/NET0131  & n33690 ;
  assign n34736 = \core_dag_ilm2reg_I5_we_DO_reg[7]/NET0131  & n33688 ;
  assign n34737 = \core_dag_ilm2reg_I7_we_DO_reg[7]/NET0131  & n33686 ;
  assign n34741 = ~n34736 & ~n34737 ;
  assign n34742 = ~n34738 & n34741 ;
  assign n34743 = n34740 & n34742 ;
  assign n34744 = ~n34739 & n34743 ;
  assign n34745 = ~\core_dag_ilm2reg_I_reg[7]/NET0131  & n21579 ;
  assign n34746 = ~n34744 & ~n34745 ;
  assign n34751 = ~n24106 & ~n33896 ;
  assign n34747 = n24170 & n33091 ;
  assign n34752 = ~n21592 & ~n34747 ;
  assign n34750 = \core_dag_ilm1reg_I1_we_DO_reg[7]/NET0131  & n33937 ;
  assign n34748 = \core_dag_ilm1reg_I3_we_DO_reg[7]/NET0131  & n33908 ;
  assign n34749 = \core_dag_ilm1reg_I2_we_DO_reg[7]/NET0131  & n33910 ;
  assign n34753 = ~n34748 & ~n34749 ;
  assign n34754 = ~n34750 & n34753 ;
  assign n34755 = n34752 & n34754 ;
  assign n34756 = ~n34751 & n34755 ;
  assign n34757 = ~\core_dag_ilm1reg_I_reg[7]/NET0131  & n21592 ;
  assign n34758 = ~n34756 & ~n34757 ;
  assign n34763 = ~n24111 & ~n33896 ;
  assign n34759 = n24173 & n33091 ;
  assign n34764 = ~n21592 & ~n34759 ;
  assign n34762 = \core_dag_ilm1reg_I1_we_DO_reg[6]/NET0131  & n33937 ;
  assign n34760 = \core_dag_ilm1reg_I3_we_DO_reg[6]/NET0131  & n33908 ;
  assign n34761 = \core_dag_ilm1reg_I2_we_DO_reg[6]/NET0131  & n33910 ;
  assign n34765 = ~n34760 & ~n34761 ;
  assign n34766 = ~n34762 & n34765 ;
  assign n34767 = n34764 & n34766 ;
  assign n34768 = ~n34763 & n34767 ;
  assign n34769 = ~\core_dag_ilm1reg_I_reg[6]/NET0131  & n21592 ;
  assign n34770 = ~n34768 & ~n34769 ;
  assign n34775 = ~n24118 & ~n33896 ;
  assign n34771 = \core_dag_ilm1reg_I2_we_DO_reg[4]/NET0131  & n33910 ;
  assign n34776 = ~n21592 & ~n34771 ;
  assign n34774 = \core_dag_ilm1reg_I3_we_DO_reg[4]/NET0131  & n33908 ;
  assign n34772 = \core_dag_ilm1reg_I1_we_DO_reg[4]/NET0131  & n33937 ;
  assign n34773 = \core_dag_ilm1reg_I0_we_DO_reg[4]/NET0131  & n33922 ;
  assign n34777 = ~n34772 & ~n34773 ;
  assign n34778 = ~n34774 & n34777 ;
  assign n34779 = n34776 & n34778 ;
  assign n34780 = ~n34775 & n34779 ;
  assign n34781 = ~\core_dag_ilm1reg_I_reg[4]/NET0131  & n21592 ;
  assign n34782 = ~n34780 & ~n34781 ;
  assign n34786 = n23886 & ~n33896 ;
  assign n34783 = \core_dag_ilm1reg_I2_we_DO_reg[3]/NET0131  & n33910 ;
  assign n34788 = ~n21592 & ~n34783 ;
  assign n34787 = \core_dag_ilm1reg_I0_we_DO_reg[3]/NET0131  & n33922 ;
  assign n34784 = \core_dag_ilm1reg_I1_we_DO_reg[3]/NET0131  & n33937 ;
  assign n34785 = \core_dag_ilm1reg_I3_we_DO_reg[3]/NET0131  & n33908 ;
  assign n34789 = ~n34784 & ~n34785 ;
  assign n34790 = ~n34787 & n34789 ;
  assign n34791 = n34788 & n34790 ;
  assign n34792 = ~n34786 & n34791 ;
  assign n34793 = ~\core_dag_ilm1reg_I_reg[3]/NET0131  & n21592 ;
  assign n34794 = ~n34792 & ~n34793 ;
  assign n34799 = ~n24124 & ~n33896 ;
  assign n34795 = \core_dag_ilm1reg_I0_we_DO_reg[2]/NET0131  & n33922 ;
  assign n34800 = ~n21592 & ~n34795 ;
  assign n34798 = \core_dag_ilm1reg_I3_we_DO_reg[2]/NET0131  & n33908 ;
  assign n34796 = \core_dag_ilm1reg_I1_we_DO_reg[2]/NET0131  & n33937 ;
  assign n34797 = \core_dag_ilm1reg_I2_we_DO_reg[2]/NET0131  & n33910 ;
  assign n34801 = ~n34796 & ~n34797 ;
  assign n34802 = ~n34798 & n34801 ;
  assign n34803 = n34800 & n34802 ;
  assign n34804 = ~n34799 & n34803 ;
  assign n34805 = ~\core_dag_ilm1reg_I_reg[2]/NET0131  & n21592 ;
  assign n34806 = ~n34804 & ~n34805 ;
  assign n34811 = ~n24143 & ~n33896 ;
  assign n34807 = \core_dag_ilm1reg_I2_we_DO_reg[0]/NET0131  & n33910 ;
  assign n34812 = ~n21592 & ~n34807 ;
  assign n34810 = \core_dag_ilm1reg_I1_we_DO_reg[0]/NET0131  & n33937 ;
  assign n34808 = \core_dag_ilm1reg_I3_we_DO_reg[0]/NET0131  & n33908 ;
  assign n34809 = \core_dag_ilm1reg_I0_we_DO_reg[0]/NET0131  & n33922 ;
  assign n34813 = ~n34808 & ~n34809 ;
  assign n34814 = ~n34810 & n34813 ;
  assign n34815 = n34812 & n34814 ;
  assign n34816 = ~n34811 & n34815 ;
  assign n34817 = ~\core_dag_ilm1reg_I_reg[0]/NET0131  & n21592 ;
  assign n34818 = ~n34816 & ~n34817 ;
  assign n34819 = ~n5950 & ~n27908 ;
  assign n34820 = \core_c_psq_cntstk_ptr_reg[2]/NET0131  & n33341 ;
  assign n34821 = \core_c_psq_CNTRval_reg/NET0131  & ~n34820 ;
  assign n34822 = ~n34819 & ~n34821 ;
  assign n34823 = ~\sice_IIRC_reg[8]/NET0131  & ~n18871 ;
  assign n34824 = ~n20853 & ~n34823 ;
  assign n34827 = ~n26336 & n28982 ;
  assign n34825 = \sice_ICS_reg[2]/NET0131  & n26064 ;
  assign n34826 = \sice_SPC_reg[20]/P0001  & n34825 ;
  assign n34828 = \sice_SPC_reg[22]/P0001  & ~n34825 ;
  assign n34829 = ~n34826 & ~n34828 ;
  assign n34830 = ~n34827 & n34829 ;
  assign n34835 = \sice_IIRC_reg[21]/NET0131  & n24267 ;
  assign n34836 = \sice_DMR2_reg[15]/NET0131  & n25025 ;
  assign n34850 = ~n34835 & ~n34836 ;
  assign n34837 = \sice_CLR_I_reg/NET0131  & n23029 ;
  assign n34838 = \sice_idr1_reg_DO_reg[9]/P0001  & n26968 ;
  assign n34851 = ~n34837 & ~n34838 ;
  assign n34857 = n34850 & n34851 ;
  assign n34831 = n23028 & n25053 ;
  assign n34832 = \sice_IBR1_reg[15]/P0001  & n34831 ;
  assign n34848 = ~n25084 & ~n34832 ;
  assign n34833 = \sice_IMR2_reg[15]/NET0131  & n25034 ;
  assign n34834 = \sice_DBR1_reg[16]/P0001  & n25054 ;
  assign n34849 = ~n34833 & ~n34834 ;
  assign n34858 = n34848 & n34849 ;
  assign n34859 = n34857 & n34858 ;
  assign n34846 = n25033 & n25053 ;
  assign n34847 = \sice_IMR1_reg[15]/NET0131  & n34846 ;
  assign n34844 = \core_c_dec_IR_reg[21]/NET0131  & n28203 ;
  assign n34845 = \sice_IBR2_reg[15]/P0001  & n25074 ;
  assign n34854 = ~n34844 & ~n34845 ;
  assign n34855 = ~n34847 & n34854 ;
  assign n34839 = \sice_DMR1_reg[15]/NET0131  & n27903 ;
  assign n34840 = \sice_ICYC_reg[21]/NET0131  & n23409 ;
  assign n34852 = ~n34839 & ~n34840 ;
  assign n34841 = n23027 & n25010 ;
  assign n34842 = \sice_IRR_reg[11]/P0001  & n34841 ;
  assign n34843 = \sice_DBR2_reg[16]/P0001  & n25012 ;
  assign n34853 = ~n34842 & ~n34843 ;
  assign n34856 = n34852 & n34853 ;
  assign n34860 = n34855 & n34856 ;
  assign n34861 = n34859 & n34860 ;
  assign n34862 = n34827 & n34861 ;
  assign n34863 = ~n34830 & ~n34862 ;
  assign n34864 = n18262 & ~n24721 ;
  assign n34865 = ~\core_eu_em_mac_em_reg_mr2swe_DO_reg[5]/P0001  & ~n28530 ;
  assign n34866 = ~n19381 & n20259 ;
  assign n34867 = n28534 & ~n34866 ;
  assign n34868 = ~n34865 & ~n34867 ;
  assign n34869 = ~n19385 & ~n34868 ;
  assign n34870 = ~\core_eu_em_mac_em_reg_mr2swe_DO_reg[5]/P0001  & ~n28532 ;
  assign n34871 = ~n34869 & ~n34870 ;
  assign n34872 = n28529 & ~n34871 ;
  assign n34873 = ~n34864 & ~n34872 ;
  assign n34874 = \core_c_dec_MTMSTAT_Eg_reg/P0001  & ~n10069 ;
  assign n34878 = \core_c_psq_ststk_sts7x23_STcell_reg[1][12]/P0001  & n14708 ;
  assign n34879 = \core_c_psq_ststk_sts7x23_STcell_reg[6][12]/P0001  & n14711 ;
  assign n34884 = ~n34878 & ~n34879 ;
  assign n34880 = \core_c_psq_ststk_sts7x23_STcell_reg[5][12]/P0001  & n14699 ;
  assign n34881 = \core_c_psq_ststk_sts7x23_STcell_reg[4][12]/P0001  & n14706 ;
  assign n34885 = ~n34880 & ~n34881 ;
  assign n34886 = n34884 & n34885 ;
  assign n34875 = \core_c_psq_ststk_sts7x23_STcell_reg[0][12]/P0001  & n14702 ;
  assign n34882 = ~\core_c_dec_Modctl_Eg_reg/P0001  & ~n34875 ;
  assign n34876 = \core_c_psq_ststk_sts7x23_STcell_reg[2][12]/P0001  & n14713 ;
  assign n34877 = \core_c_psq_ststk_sts7x23_STcell_reg[3][12]/P0001  & n14704 ;
  assign n34883 = ~n34876 & ~n34877 ;
  assign n34887 = n34882 & n34883 ;
  assign n34888 = n34886 & n34887 ;
  assign n34889 = ~\core_c_dec_IRE_reg[11]/NET0131  & \core_c_psq_MSTAT_reg_DO_reg[4]/NET0131  ;
  assign n34890 = \core_c_dec_Modctl_Eg_reg/P0001  & ~n34255 ;
  assign n34891 = ~n34889 & n34890 ;
  assign n34892 = ~n34888 & ~n34891 ;
  assign n34893 = ~\core_c_dec_MTMSTAT_Eg_reg/P0001  & ~n34892 ;
  assign n34894 = ~n34874 & ~n34893 ;
  assign n34895 = \core_c_dec_MTMSTAT_Eg_reg/P0001  & ~n7607 ;
  assign n34897 = \core_c_dec_IRE_reg[4]/NET0131  & \core_c_dec_IRE_reg[7]/NET0131  ;
  assign n34896 = ~\core_c_dec_IRE_reg[7]/NET0131  & \core_c_psq_MSTAT_reg_DO_reg[0]/P0002  ;
  assign n34898 = \core_c_dec_Modctl_Eg_reg/P0001  & ~n34896 ;
  assign n34899 = ~n34897 & n34898 ;
  assign n34903 = \core_c_psq_ststk_sts7x23_STcell_reg[3][8]/P0001  & n14704 ;
  assign n34904 = \core_c_psq_ststk_sts7x23_STcell_reg[4][8]/P0001  & n14706 ;
  assign n34909 = ~n34903 & ~n34904 ;
  assign n34905 = \core_c_psq_ststk_sts7x23_STcell_reg[5][8]/P0001  & n14699 ;
  assign n34906 = \core_c_psq_ststk_sts7x23_STcell_reg[0][8]/P0001  & n14702 ;
  assign n34910 = ~n34905 & ~n34906 ;
  assign n34911 = n34909 & n34910 ;
  assign n34900 = \core_c_psq_ststk_sts7x23_STcell_reg[6][8]/P0001  & n14711 ;
  assign n34907 = ~\core_c_dec_Modctl_Eg_reg/P0001  & ~n34900 ;
  assign n34901 = \core_c_psq_ststk_sts7x23_STcell_reg[1][8]/P0001  & n14708 ;
  assign n34902 = \core_c_psq_ststk_sts7x23_STcell_reg[2][8]/P0001  & n14713 ;
  assign n34908 = ~n34901 & ~n34902 ;
  assign n34912 = n34907 & n34908 ;
  assign n34913 = n34911 & n34912 ;
  assign n34914 = ~n34899 & ~n34913 ;
  assign n34915 = ~\core_c_dec_MTMSTAT_Eg_reg/P0001  & ~n34914 ;
  assign n34916 = ~n34895 & ~n34915 ;
  assign n34917 = \bdma_WRlat_reg/P0001  & n13150 ;
  assign n34918 = \bdma_WRlat_reg/P0001  & ~n34065 ;
  assign n34919 = \bdma_WRlat_reg/P0001  & ~n34060 ;
  assign n34920 = \bdma_BWdataBUF_reg[6]/P0001  & ~n34919 ;
  assign n34921 = \bdma_BWdataBUF_h_reg[6]/P0001  & n34919 ;
  assign n34922 = ~n34920 & ~n34921 ;
  assign n34923 = ~n34918 & ~n34922 ;
  assign n34924 = \bdma_BWdataBUF_h_reg[14]/P0001  & n34918 ;
  assign n34925 = ~n34923 & ~n34924 ;
  assign n34926 = ~n34917 & ~n34925 ;
  assign n34927 = \bdma_BWdataBUF_h_reg[22]/P0001  & n34917 ;
  assign n34928 = ~n34926 & ~n34927 ;
  assign n34929 = \bdma_BWdataBUF_reg[5]/P0001  & ~n34919 ;
  assign n34930 = \bdma_BWdataBUF_h_reg[5]/P0001  & n34919 ;
  assign n34931 = ~n34929 & ~n34930 ;
  assign n34932 = ~n34918 & ~n34931 ;
  assign n34933 = \bdma_BWdataBUF_h_reg[13]/P0001  & n34918 ;
  assign n34934 = ~n34932 & ~n34933 ;
  assign n34935 = ~n34917 & ~n34934 ;
  assign n34936 = \bdma_BWdataBUF_h_reg[21]/P0001  & n34917 ;
  assign n34937 = ~n34935 & ~n34936 ;
  assign n34938 = \bdma_BWdataBUF_reg[7]/P0001  & ~n34919 ;
  assign n34939 = \bdma_BWdataBUF_h_reg[7]/P0001  & n34919 ;
  assign n34940 = ~n34938 & ~n34939 ;
  assign n34941 = ~n34918 & ~n34940 ;
  assign n34942 = \bdma_BWdataBUF_h_reg[15]/P0001  & n34918 ;
  assign n34943 = ~n34941 & ~n34942 ;
  assign n34944 = ~n34917 & ~n34943 ;
  assign n34945 = \bdma_BWdataBUF_h_reg[23]/P0001  & n34917 ;
  assign n34946 = ~n34944 & ~n34945 ;
  assign n34947 = \bdma_BWdataBUF_reg[4]/P0001  & ~n34919 ;
  assign n34948 = \bdma_BWdataBUF_h_reg[4]/P0001  & n34919 ;
  assign n34949 = ~n34947 & ~n34948 ;
  assign n34950 = ~n34918 & ~n34949 ;
  assign n34951 = \bdma_BWdataBUF_h_reg[12]/P0001  & n34918 ;
  assign n34952 = ~n34950 & ~n34951 ;
  assign n34953 = ~n34917 & ~n34952 ;
  assign n34954 = \bdma_BWdataBUF_h_reg[20]/P0001  & n34917 ;
  assign n34955 = ~n34953 & ~n34954 ;
  assign n34956 = \bdma_BWdataBUF_reg[3]/P0001  & ~n34919 ;
  assign n34957 = \bdma_BWdataBUF_h_reg[3]/P0001  & n34919 ;
  assign n34958 = ~n34956 & ~n34957 ;
  assign n34959 = ~n34918 & ~n34958 ;
  assign n34960 = \bdma_BWdataBUF_h_reg[11]/P0001  & n34918 ;
  assign n34961 = ~n34959 & ~n34960 ;
  assign n34962 = ~n34917 & ~n34961 ;
  assign n34963 = \bdma_BWdataBUF_h_reg[19]/P0001  & n34917 ;
  assign n34964 = ~n34962 & ~n34963 ;
  assign n34965 = \bdma_BWdataBUF_reg[2]/P0001  & ~n34919 ;
  assign n34966 = \bdma_BWdataBUF_h_reg[2]/P0001  & n34919 ;
  assign n34967 = ~n34965 & ~n34966 ;
  assign n34968 = ~n34918 & ~n34967 ;
  assign n34969 = \bdma_BWdataBUF_h_reg[10]/P0001  & n34918 ;
  assign n34970 = ~n34968 & ~n34969 ;
  assign n34971 = ~n34917 & ~n34970 ;
  assign n34972 = \bdma_BWdataBUF_h_reg[18]/P0001  & n34917 ;
  assign n34973 = ~n34971 & ~n34972 ;
  assign n34974 = \bdma_BWdataBUF_reg[1]/P0001  & ~n34919 ;
  assign n34975 = \bdma_BWdataBUF_h_reg[1]/P0001  & n34919 ;
  assign n34976 = ~n34974 & ~n34975 ;
  assign n34977 = ~n34918 & ~n34976 ;
  assign n34978 = \bdma_BWdataBUF_h_reg[9]/P0001  & n34918 ;
  assign n34979 = ~n34977 & ~n34978 ;
  assign n34980 = ~n34917 & ~n34979 ;
  assign n34981 = \bdma_BWdataBUF_h_reg[17]/P0001  & n34917 ;
  assign n34982 = ~n34980 & ~n34981 ;
  assign n34983 = \bdma_BWdataBUF_reg[0]/P0001  & ~n34919 ;
  assign n34984 = \bdma_BWdataBUF_h_reg[0]/P0001  & n34919 ;
  assign n34985 = ~n34983 & ~n34984 ;
  assign n34986 = ~n34918 & ~n34985 ;
  assign n34987 = \bdma_BWdataBUF_h_reg[8]/P0001  & n34918 ;
  assign n34988 = ~n34986 & ~n34987 ;
  assign n34989 = ~n34917 & ~n34988 ;
  assign n34990 = \bdma_BWdataBUF_h_reg[16]/P0001  & n34917 ;
  assign n34991 = ~n34989 & ~n34990 ;
  assign n34992 = \sice_SPC_reg[11]/P0001  & n34825 ;
  assign n34993 = \sice_SPC_reg[13]/P0001  & ~n34825 ;
  assign n34994 = ~n34992 & ~n34993 ;
  assign n34995 = ~n34827 & n34994 ;
  assign n34999 = \sice_IMR1_reg[6]/NET0131  & n34846 ;
  assign n35000 = \sice_idr1_reg_DO_reg[0]/P0001  & n26968 ;
  assign n35012 = ~n34999 & ~n35000 ;
  assign n35001 = \sice_DMR1_reg[6]/NET0131  & n27903 ;
  assign n35002 = \sice_IIRC_reg[12]/NET0131  & n24267 ;
  assign n35013 = ~n35001 & ~n35002 ;
  assign n35020 = n35012 & n35013 ;
  assign n34998 = \sice_ITR_reg[2]/NET0131  & n25084 ;
  assign n34996 = \sice_DMR2_reg[6]/NET0131  & n25025 ;
  assign n34997 = \sice_DBR1_reg[7]/P0001  & n25054 ;
  assign n35011 = ~n34996 & ~n34997 ;
  assign n35021 = ~n34998 & n35011 ;
  assign n35022 = n35020 & n35021 ;
  assign n35007 = \sice_ICYC_reg[12]/NET0131  & n23409 ;
  assign n35008 = ~\sice_IAR_reg[2]/NET0131  & n25083 ;
  assign n35016 = ~n35007 & ~n35008 ;
  assign n35009 = \sice_IBR2_reg[6]/P0001  & n25074 ;
  assign n35010 = \core_c_dec_IR_reg[12]/NET0131  & n28203 ;
  assign n35017 = ~n35009 & ~n35010 ;
  assign n35018 = n35016 & n35017 ;
  assign n35003 = \sice_IMR2_reg[6]/NET0131  & n25034 ;
  assign n35004 = \sice_IBR1_reg[6]/P0001  & n34831 ;
  assign n35014 = ~n35003 & ~n35004 ;
  assign n35005 = \sice_DBR2_reg[7]/P0001  & n25012 ;
  assign n35006 = \sice_IRR_reg[2]/P0001  & n34841 ;
  assign n35015 = ~n35005 & ~n35006 ;
  assign n35019 = n35014 & n35015 ;
  assign n35023 = n35018 & n35019 ;
  assign n35024 = n35022 & n35023 ;
  assign n35025 = n34827 & n35024 ;
  assign n35026 = ~n34995 & ~n35025 ;
  assign n35027 = \sice_SPC_reg[10]/P0001  & n34825 ;
  assign n35028 = \sice_SPC_reg[12]/P0001  & ~n34825 ;
  assign n35029 = ~n35027 & ~n35028 ;
  assign n35030 = ~n34827 & n35029 ;
  assign n35032 = \sice_IMR2_reg[5]/NET0131  & n25034 ;
  assign n35033 = \sice_ICYC_reg[11]/NET0131  & n23409 ;
  assign n35046 = ~n35032 & ~n35033 ;
  assign n35035 = \sice_DBR1_reg[6]/P0001  & n25054 ;
  assign n35036 = \core_c_dec_IR_reg[11]/NET0131  & n28203 ;
  assign n35047 = ~n35035 & ~n35036 ;
  assign n35054 = n35046 & n35047 ;
  assign n35034 = \sice_ITR_reg[1]/NET0131  & n25084 ;
  assign n35031 = \sice_IBR2_reg[5]/P0001  & n25074 ;
  assign n35045 = ~n35008 & ~n35031 ;
  assign n35055 = ~n35034 & n35045 ;
  assign n35056 = n35054 & n35055 ;
  assign n35041 = \sice_DBR2_reg[6]/P0001  & n25012 ;
  assign n35042 = \sice_IIRC_reg[11]/NET0131  & n24267 ;
  assign n35050 = ~n35041 & ~n35042 ;
  assign n35043 = \sice_DMR1_reg[5]/NET0131  & n27903 ;
  assign n35044 = \sice_IRR_reg[1]/P0001  & n34841 ;
  assign n35051 = ~n35043 & ~n35044 ;
  assign n35052 = n35050 & n35051 ;
  assign n35037 = \sice_IMR1_reg[5]/NET0131  & n34846 ;
  assign n35038 = \sice_DMR2_reg[5]/NET0131  & n25025 ;
  assign n35048 = ~n35037 & ~n35038 ;
  assign n35039 = \sice_IBR1_reg[5]/P0001  & n34831 ;
  assign n35040 = \sice_idr0_reg_DO_reg[11]/P0001  & n26968 ;
  assign n35049 = ~n35039 & ~n35040 ;
  assign n35053 = n35048 & n35049 ;
  assign n35057 = n35052 & n35053 ;
  assign n35058 = n35056 & n35057 ;
  assign n35059 = n34827 & n35058 ;
  assign n35060 = ~n35030 & ~n35059 ;
  assign n35061 = \sice_SPC_reg[9]/P0001  & n34825 ;
  assign n35062 = \sice_SPC_reg[11]/P0001  & ~n34825 ;
  assign n35063 = ~n35061 & ~n35062 ;
  assign n35064 = ~n34827 & n35063 ;
  assign n35066 = \sice_IMR2_reg[4]/NET0131  & n25034 ;
  assign n35067 = \sice_IIRC_reg[10]/NET0131  & n24267 ;
  assign n35080 = ~n35066 & ~n35067 ;
  assign n35069 = \sice_DBR1_reg[5]/P0001  & n25054 ;
  assign n35070 = \core_c_dec_IR_reg[10]/NET0131  & n28203 ;
  assign n35081 = ~n35069 & ~n35070 ;
  assign n35088 = n35080 & n35081 ;
  assign n35068 = \sice_ITR_reg[0]/NET0131  & n25084 ;
  assign n35065 = \sice_IBR2_reg[4]/P0001  & n25074 ;
  assign n35079 = ~n35008 & ~n35065 ;
  assign n35089 = ~n35068 & n35079 ;
  assign n35090 = n35088 & n35089 ;
  assign n35075 = \sice_DMR2_reg[4]/NET0131  & n25025 ;
  assign n35076 = \sice_DBR2_reg[5]/P0001  & n25012 ;
  assign n35084 = ~n35075 & ~n35076 ;
  assign n35077 = \sice_DMR1_reg[4]/NET0131  & n27903 ;
  assign n35078 = \sice_IRR_reg[0]/P0001  & n34841 ;
  assign n35085 = ~n35077 & ~n35078 ;
  assign n35086 = n35084 & n35085 ;
  assign n35071 = \sice_IMR1_reg[4]/NET0131  & n34846 ;
  assign n35072 = \sice_ICYC_reg[10]/NET0131  & n23409 ;
  assign n35082 = ~n35071 & ~n35072 ;
  assign n35073 = \sice_IBR1_reg[4]/P0001  & n34831 ;
  assign n35074 = \sice_idr0_reg_DO_reg[10]/P0001  & n26968 ;
  assign n35083 = ~n35073 & ~n35074 ;
  assign n35087 = n35082 & n35083 ;
  assign n35091 = n35086 & n35087 ;
  assign n35092 = n35090 & n35091 ;
  assign n35093 = n34827 & n35092 ;
  assign n35094 = ~n35064 & ~n35093 ;
  assign n35095 = ~\sice_ICYC_reg[8]/NET0131  & ~n18863 ;
  assign n35096 = ~n20738 & ~n35095 ;
  assign n35097 = ~\clkc_oscntr_reg_DO_reg[6]/NET0131  & ~n23419 ;
  assign n35098 = ~n23420 & ~n35097 ;
  assign n35099 = n18262 & n25069 ;
  assign n35100 = ~\core_eu_em_mac_em_reg_mr2swe_DO_reg[4]/P0001  & ~n28530 ;
  assign n35101 = ~n19381 & n20080 ;
  assign n35102 = n28534 & ~n35101 ;
  assign n35103 = ~n35100 & ~n35102 ;
  assign n35104 = ~n19385 & ~n35103 ;
  assign n35105 = ~\core_eu_em_mac_em_reg_mr2swe_DO_reg[4]/P0001  & ~n28532 ;
  assign n35106 = ~n35104 & ~n35105 ;
  assign n35107 = n28529 & ~n35106 ;
  assign n35108 = ~n35099 & ~n35107 ;
  assign n35109 = n18262 & ~n25088 ;
  assign n35110 = ~\core_eu_em_mac_em_reg_mr2swe_DO_reg[0]/P0001  & ~n28530 ;
  assign n35111 = ~n19381 & n19559 ;
  assign n35112 = n28534 & ~n35111 ;
  assign n35113 = ~n35110 & ~n35112 ;
  assign n35114 = ~n19385 & ~n35113 ;
  assign n35115 = ~\core_eu_em_mac_em_reg_mr2swe_DO_reg[0]/P0001  & ~n28532 ;
  assign n35116 = ~n35114 & ~n35115 ;
  assign n35117 = n28529 & ~n35116 ;
  assign n35118 = ~n35109 & ~n35117 ;
  assign n35119 = n6560 & n6599 ;
  assign n35120 = n8198 & ~n35119 ;
  assign n35121 = \core_dag_ilm1reg_STEALI_E_reg[2]/P0001  & ~n35120 ;
  assign n35122 = n6221 & n6315 ;
  assign n35123 = ~n7631 & ~n35122 ;
  assign n35124 = ~\core_dag_ilm1reg_STEALI_E_reg[2]/P0001  & ~n35123 ;
  assign n35125 = ~n35121 & ~n35124 ;
  assign n35126 = \auctl_T0Sack_reg/NET0131  & n35125 ;
  assign n35127 = \auctl_R0Sack_reg/NET0131  & n35125 ;
  assign n35128 = \auctl_T1Sack_reg/NET0131  & n35125 ;
  assign n35129 = \auctl_R1Sack_reg/NET0131  & n35125 ;
  assign n35130 = \core_c_dec_MTIreg_E_reg[4]/P0001  & n4117 ;
  assign n35131 = n32000 & ~n32001 ;
  assign n35132 = n31992 & n35131 ;
  assign n35133 = ~n4117 & n32007 ;
  assign n35134 = ~n32003 & n35133 ;
  assign n35135 = n32014 & n35134 ;
  assign n35136 = n35132 & n35135 ;
  assign n35137 = ~n35130 & ~n35136 ;
  assign n35138 = n4116 & ~n35137 ;
  assign n35139 = ~\core_c_dec_IRE_reg[0]/NET0131  & ~\core_c_dec_IRE_reg[1]/NET0131  ;
  assign n35140 = ~\core_c_dec_IRE_reg[2]/NET0131  & n35139 ;
  assign n35141 = \clkc_SIDLE_s1_reg/NET0131  & ~\clkc_SIDLE_s2_reg/NET0131  ;
  assign n35142 = ~n35140 & n35141 ;
  assign n35144 = ~\clkc_SlowDn_reg/NET0131  & ~n35142 ;
  assign n35143 = ~\clkc_STBY_reg/NET0131  & n35142 ;
  assign n35145 = n23018 & ~n35143 ;
  assign n35146 = ~n35144 & n35145 ;
  assign n35147 = n33221 & n35146 ;
  assign n35148 = ~\clkc_STDcnt_reg[7]/NET0131  & ~n31527 ;
  assign n35149 = ~n31521 & ~n31528 ;
  assign n35150 = ~n35148 & n35149 ;
  assign n35151 = \core_c_dec_MTIreg_E_reg[7]/P0001  & n4117 ;
  assign n35152 = n34465 & n35132 ;
  assign n35153 = ~n35151 & ~n35152 ;
  assign n35154 = n4116 & ~n35153 ;
  assign n35155 = \core_c_dec_MTDMOVL_E_reg/P0001  & n4117 ;
  assign n35156 = n32020 & n34463 ;
  assign n35157 = ~n35155 & ~n35156 ;
  assign n35158 = n4116 & ~n35157 ;
  assign n35160 = ~n4117 & ~n32017 ;
  assign n35159 = ~\core_c_dec_MTASTAT_E_reg/P0001  & n4117 ;
  assign n35161 = n4116 & ~n35159 ;
  assign n35162 = ~n35160 & n35161 ;
  assign n35163 = \core_c_dec_MTSB_E_reg/P0001  & n4117 ;
  assign n35164 = n32004 & n35133 ;
  assign n35165 = n31992 & n31999 ;
  assign n35166 = n35164 & n35165 ;
  assign n35167 = ~n35163 & ~n35166 ;
  assign n35168 = n4116 & ~n35167 ;
  assign n35169 = \core_c_dec_MTRX1_E_reg/P0001  & n4117 ;
  assign n35170 = n34462 & n35134 ;
  assign n35171 = n32018 & n35170 ;
  assign n35172 = ~n35169 & ~n35171 ;
  assign n35173 = n4116 & ~n35172 ;
  assign n35174 = \core_c_dec_MTRX0_E_reg/P0001  & n4117 ;
  assign n35175 = n32018 & n35135 ;
  assign n35176 = ~n35174 & ~n35175 ;
  assign n35177 = n4116 & ~n35176 ;
  assign n35178 = \core_c_dec_MTPMOVL_E_reg/P0001  & n4117 ;
  assign n35179 = n32020 & n35133 ;
  assign n35180 = ~n35178 & ~n35179 ;
  assign n35181 = n4116 & ~n35180 ;
  assign n35182 = \core_c_dec_MTOWRCNTR_Eg_reg/P0001  & n4117 ;
  assign n35183 = ~n31995 & n31998 ;
  assign n35184 = n11741 & n35183 ;
  assign n35185 = ~n31992 & n35184 ;
  assign n35186 = n32004 & n34463 ;
  assign n35187 = n35185 & n35186 ;
  assign n35188 = ~n35182 & ~n35187 ;
  assign n35189 = n4116 & ~n35188 ;
  assign n35190 = \core_c_dec_MTMreg_E_reg[7]/P0001  & n4117 ;
  assign n35191 = n34464 & n35132 ;
  assign n35192 = n31999 & n35191 ;
  assign n35193 = ~n35190 & ~n35192 ;
  assign n35194 = n4116 & ~n35193 ;
  assign n35195 = \core_c_dec_MTMreg_E_reg[6]/P0001  & n4117 ;
  assign n35196 = n35132 & n35134 ;
  assign n35197 = n31999 & n35196 ;
  assign n35198 = ~n35195 & ~n35197 ;
  assign n35199 = n4116 & ~n35198 ;
  assign n35200 = \core_c_dec_MTMreg_E_reg[5]/P0001  & n4117 ;
  assign n35201 = n35183 & n35191 ;
  assign n35202 = ~n35200 & ~n35201 ;
  assign n35203 = n4116 & ~n35202 ;
  assign n35204 = \core_c_dec_MTMreg_E_reg[4]/P0001  & n4117 ;
  assign n35205 = n35183 & n35196 ;
  assign n35206 = ~n35204 & ~n35205 ;
  assign n35207 = n4116 & ~n35206 ;
  assign n35208 = ~n31998 & ~n32007 ;
  assign n35209 = n34479 & n35208 ;
  assign n35210 = n34476 & n35209 ;
  assign n35211 = \core_c_dec_MTMreg_E_reg[3]/P0001  & n4117 ;
  assign n35212 = ~n35210 & ~n35211 ;
  assign n35213 = n4116 & ~n35212 ;
  assign n35214 = ~n31998 & n32007 ;
  assign n35215 = n34479 & n35214 ;
  assign n35216 = n34476 & n35215 ;
  assign n35217 = \core_c_dec_MTMreg_E_reg[2]/P0001  & n4117 ;
  assign n35218 = ~n35216 & ~n35217 ;
  assign n35219 = n4116 & ~n35218 ;
  assign n35220 = \core_c_dec_MTMreg_E_reg[0]/P0001  & n4117 ;
  assign n35221 = n34475 & n34479 ;
  assign n35222 = n32007 & n35183 ;
  assign n35223 = n35221 & n35222 ;
  assign n35224 = ~n35220 & ~n35223 ;
  assign n35225 = n4116 & ~n35224 ;
  assign n35226 = ~n31992 & n35131 ;
  assign n35227 = n34465 & n35226 ;
  assign n35228 = \core_c_dec_MTLreg_E_reg[7]/P0001  & n4117 ;
  assign n35229 = ~n35227 & ~n35228 ;
  assign n35230 = n4116 & ~n35229 ;
  assign n35231 = n35170 & n35226 ;
  assign n35232 = \core_c_dec_MTLreg_E_reg[6]/P0001  & n4117 ;
  assign n35233 = ~n35231 & ~n35232 ;
  assign n35234 = n4116 & ~n35233 ;
  assign n35235 = n34470 & n35226 ;
  assign n35236 = \core_c_dec_MTLreg_E_reg[5]/P0001  & n4117 ;
  assign n35237 = ~n35235 & ~n35236 ;
  assign n35238 = n4116 & ~n35237 ;
  assign n35239 = \core_c_dec_MTLreg_E_reg[4]/P0001  & n4117 ;
  assign n35240 = n35135 & n35226 ;
  assign n35241 = ~n35239 & ~n35240 ;
  assign n35242 = n4116 & ~n35241 ;
  assign n35243 = \core_c_dec_MTLreg_E_reg[3]/P0001  & n4117 ;
  assign n35244 = ~n4117 & n32019 ;
  assign n35245 = n31995 & n35244 ;
  assign n35246 = n35208 & n35245 ;
  assign n35247 = ~n35243 & ~n35246 ;
  assign n35248 = n4116 & ~n35247 ;
  assign n35249 = \core_c_dec_MTLreg_E_reg[2]/P0001  & n4117 ;
  assign n35250 = n35214 & n35245 ;
  assign n35251 = ~n35249 & ~n35250 ;
  assign n35252 = n4116 & ~n35251 ;
  assign n35253 = \core_c_dec_MTLreg_E_reg[1]/P0001  & n4117 ;
  assign n35254 = n34477 & n35245 ;
  assign n35255 = ~n35253 & ~n35254 ;
  assign n35256 = n4116 & ~n35255 ;
  assign n35257 = \core_c_dec_MTLreg_E_reg[0]/P0001  & n4117 ;
  assign n35258 = n32015 & n35244 ;
  assign n35259 = ~n35257 & ~n35258 ;
  assign n35260 = n4116 & ~n35259 ;
  assign n35261 = \core_c_dec_MTIreg_E_reg[6]/P0001  & n4117 ;
  assign n35262 = n35132 & n35170 ;
  assign n35263 = ~n35261 & ~n35262 ;
  assign n35264 = n4116 & ~n35263 ;
  assign n35265 = \core_c_dec_MTIreg_E_reg[5]/P0001  & n4117 ;
  assign n35266 = n34470 & n35132 ;
  assign n35267 = ~n35265 & ~n35266 ;
  assign n35268 = n4116 & ~n35267 ;
  assign n35269 = n31995 & n34475 ;
  assign n35270 = n35209 & n35269 ;
  assign n35271 = \core_c_dec_MTIreg_E_reg[3]/P0001  & n4117 ;
  assign n35272 = ~n35270 & ~n35271 ;
  assign n35273 = n4116 & ~n35272 ;
  assign n35274 = n35215 & n35269 ;
  assign n35275 = \core_c_dec_MTIreg_E_reg[2]/P0001  & n4117 ;
  assign n35276 = ~n35274 & ~n35275 ;
  assign n35277 = n4116 & ~n35276 ;
  assign n35278 = \core_c_dec_MTIreg_E_reg[1]/P0001  & n4117 ;
  assign n35279 = n34480 & n35269 ;
  assign n35280 = ~n35278 & ~n35279 ;
  assign n35281 = n4116 & ~n35280 ;
  assign n35282 = n14752 & n25069 ;
  assign n35283 = ~\core_eu_em_mac_em_reg_mr2rwe_DO_reg[4]/P0001  & ~n17799 ;
  assign n35284 = ~n17809 & n20080 ;
  assign n35285 = n17811 & ~n35284 ;
  assign n35286 = ~n35283 & ~n35285 ;
  assign n35287 = ~n17823 & ~n35286 ;
  assign n35288 = ~\core_eu_em_mac_em_reg_mr2rwe_DO_reg[4]/P0001  & ~n17808 ;
  assign n35289 = ~n35287 & ~n35288 ;
  assign n35290 = n17829 & ~n35289 ;
  assign n35291 = ~n35282 & ~n35290 ;
  assign n35292 = \core_c_dec_MTIreg_E_reg[0]/P0001  & n4117 ;
  assign n35293 = n32015 & n35221 ;
  assign n35294 = ~n35292 & ~n35293 ;
  assign n35295 = n4116 & ~n35294 ;
  assign n35296 = \core_c_dec_MTIFC_Eg_reg/P0001  & n4117 ;
  assign n35297 = n35164 & n35185 ;
  assign n35298 = ~n35296 & ~n35297 ;
  assign n35299 = n4116 & ~n35298 ;
  assign n35300 = \core_c_dec_MTIDR_E_reg/P0001  & n4117 ;
  assign n35301 = n35222 & n35244 ;
  assign n35302 = ~n35300 & ~n35301 ;
  assign n35303 = n4116 & ~n35302 ;
  assign n35304 = \core_c_dec_MTICNTL_Eg_reg/P0001  & n4117 ;
  assign n35305 = n31992 & n35184 ;
  assign n35306 = n35164 & n35305 ;
  assign n35307 = ~n35304 & ~n35306 ;
  assign n35308 = n4116 & ~n35307 ;
  assign n35309 = \core_c_dec_MTCNTR_Eg_reg/P0001  & n4117 ;
  assign n35310 = n35186 & n35305 ;
  assign n35311 = ~n35309 & ~n35310 ;
  assign n35312 = n4116 & ~n35311 ;
  assign n35313 = \bdma_BWCOUNT_reg[1]/NET0131  & ~n13764 ;
  assign n35314 = ~n13763 & ~n13765 ;
  assign n35315 = ~n35313 & n35314 ;
  assign n35316 = ~n9435 & n13763 ;
  assign n35317 = ~n35315 & ~n35316 ;
  assign n35318 = n13746 & ~n34589 ;
  assign n35320 = ~n19205 & n19296 ;
  assign n35319 = ~\core_eu_ec_cun_AC_reg/P0001  & n19205 ;
  assign n35321 = n4150 & ~n35319 ;
  assign n35322 = ~n35320 & n35321 ;
  assign n35323 = \core_c_dec_MTSR1_E_reg/P0001  & ~n19848 ;
  assign n35324 = ~\core_c_dec_MTSR1_E_reg/P0001  & n29942 ;
  assign n35325 = ~n35323 & ~n35324 ;
  assign n35326 = n18717 & ~n35325 ;
  assign n35327 = ~\core_eu_es_sht_es_reg_sr1swe_DO_reg[10]/P0001  & ~n18717 ;
  assign n35328 = ~n35326 & ~n35327 ;
  assign n35329 = n17833 & ~n35325 ;
  assign n35330 = ~\core_eu_es_sht_es_reg_sr1rwe_DO_reg[10]/P0001  & ~n17833 ;
  assign n35331 = ~n35329 & ~n35330 ;
  assign n35332 = \core_c_dec_MTSR0_E_reg/P0001  & ~n23860 ;
  assign n35333 = ~\core_c_dec_MTSR0_E_reg/P0001  & n30441 ;
  assign n35334 = ~n35332 & ~n35333 ;
  assign n35335 = n18886 & ~n35334 ;
  assign n35336 = ~\core_eu_es_sht_es_reg_sr0swe_DO_reg[8]/P0001  & ~n18886 ;
  assign n35337 = ~n35335 & ~n35336 ;
  assign n35338 = n19034 & ~n35334 ;
  assign n35339 = ~\core_eu_es_sht_es_reg_sr0rwe_DO_reg[8]/P0001  & ~n19034 ;
  assign n35340 = ~n35338 & ~n35339 ;
  assign n35341 = n14752 & ~n24721 ;
  assign n35342 = ~\core_eu_em_mac_em_reg_mr2rwe_DO_reg[5]/P0001  & ~n17799 ;
  assign n35343 = ~n17809 & n20259 ;
  assign n35344 = n17811 & ~n35343 ;
  assign n35345 = ~n35342 & ~n35344 ;
  assign n35346 = ~n17823 & ~n35345 ;
  assign n35347 = ~\core_eu_em_mac_em_reg_mr2rwe_DO_reg[5]/P0001  & ~n17808 ;
  assign n35348 = ~n35346 & ~n35347 ;
  assign n35349 = n17829 & ~n35348 ;
  assign n35350 = ~n35341 & ~n35349 ;
  assign n35353 = n18271 & ~n23860 ;
  assign n35352 = ~\core_eu_em_mac_em_reg_mr0swe_DO_reg[8]/P0001  & ~n18271 ;
  assign n35354 = n18273 & ~n35352 ;
  assign n35355 = ~n35353 & n35354 ;
  assign n35351 = \core_eu_em_mac_em_reg_mr0swe_DO_reg[8]/P0001  & ~n18266 ;
  assign n35356 = ~n18270 & ~n35351 ;
  assign n35357 = ~n35355 & n35356 ;
  assign n35358 = ~n18262 & ~n35357 ;
  assign n35359 = n18262 & n19633 ;
  assign n35360 = ~n35358 & ~n35359 ;
  assign n35361 = n14752 & ~n19633 ;
  assign n35362 = n18328 & n23860 ;
  assign n35363 = \core_eu_em_mac_em_reg_mr0rwe_DO_reg[8]/P0001  & ~n18330 ;
  assign n35364 = n18334 & ~n35363 ;
  assign n35365 = ~n35362 & n35364 ;
  assign n35366 = ~n35361 & ~n35365 ;
  assign n35367 = \bdma_BWRn_reg/NET0131  & ~\bdma_WRlat_reg/P0001  ;
  assign n35368 = ~\bdma_BCTL_reg[4]/NET0131  & ~\bdma_BCTL_reg[5]/NET0131  ;
  assign n35369 = \bdma_BCTL_reg[6]/NET0131  & ~n35368 ;
  assign n35370 = \bdma_BCTL_reg[7]/NET0131  & n35369 ;
  assign n35371 = \bdma_BWcnt_reg[4]/NET0131  & ~n35370 ;
  assign n35372 = ~\bdma_BWcnt_reg[4]/NET0131  & n35370 ;
  assign n35391 = ~n35371 & ~n35372 ;
  assign n35373 = ~\bdma_BCTL_reg[6]/NET0131  & n35368 ;
  assign n35374 = ~n35369 & ~n35373 ;
  assign n35375 = \bdma_BWcnt_reg[2]/NET0131  & ~n35374 ;
  assign n35376 = ~\bdma_BWcnt_reg[2]/NET0131  & n35374 ;
  assign n35392 = ~n35375 & ~n35376 ;
  assign n35393 = n35391 & n35392 ;
  assign n35377 = ~\bdma_BCTL_reg[7]/NET0131  & ~n35369 ;
  assign n35378 = ~\bdma_BWcnt_reg[4]/NET0131  & ~n35377 ;
  assign n35380 = ~\bdma_BWcnt_reg[3]/NET0131  & n35378 ;
  assign n35379 = \bdma_BWcnt_reg[3]/NET0131  & ~n35378 ;
  assign n35381 = \bdma_BCTL_reg[4]/NET0131  & \bdma_BCTL_reg[5]/NET0131  ;
  assign n35382 = ~n35368 & ~n35381 ;
  assign n35384 = ~\bdma_BWcnt_reg[1]/NET0131  & ~n35382 ;
  assign n35383 = \bdma_BWcnt_reg[1]/NET0131  & n35382 ;
  assign n35386 = \bdma_BCTL_reg[4]/NET0131  & \bdma_BWcnt_reg[0]/NET0131  ;
  assign n35385 = ~\bdma_BCTL_reg[4]/NET0131  & ~\bdma_BWcnt_reg[0]/NET0131  ;
  assign n35387 = \bdma_BCTL_reg[2]/NET0131  & ~n35385 ;
  assign n35388 = ~n35386 & n35387 ;
  assign n35389 = ~n35383 & n35388 ;
  assign n35390 = ~n35384 & n35389 ;
  assign n35394 = ~n35379 & n35390 ;
  assign n35395 = ~n35380 & n35394 ;
  assign n35396 = n35393 & n35395 ;
  assign n35397 = ~n35367 & ~n35396 ;
  assign n35400 = ~\sport0_regs_SCTLreg_DO_reg[4]/NET0131  & ~n34401 ;
  assign n35401 = \sport0_regs_SCTLreg_DO_reg[4]/NET0131  & ~n31046 ;
  assign n35402 = ~n35400 & ~n35401 ;
  assign n35404 = ~n31044 & ~n35402 ;
  assign n35403 = n31044 & n35402 ;
  assign n35405 = n20875 & ~n35403 ;
  assign n35406 = ~n35404 & n35405 ;
  assign n35407 = ~\sport0_rxctl_ldRX_cmp_reg/P0001  & n8460 ;
  assign n35399 = \sport0_rxctl_RX_reg[11]/P0001  & n20873 ;
  assign n35408 = ~n20868 & ~n35399 ;
  assign n35409 = ~n35407 & n35408 ;
  assign n35410 = ~n35406 & n35409 ;
  assign n35398 = ~\sport0_rxctl_RXSHT_reg[11]/P0001  & n20868 ;
  assign n35411 = ~n20871 & ~n35398 ;
  assign n35412 = ~n35410 & n35411 ;
  assign n35413 = \sport0_rxctl_RX_reg[11]/P0001  & n20871 ;
  assign n35414 = ~n35412 & ~n35413 ;
  assign n35415 = ~IACKn_pad & ~n20384 ;
  assign n35416 = ~n20821 & n35415 ;
  assign n35417 = n32465 & ~n35416 ;
  assign n35418 = ~n4117 & ~n25009 ;
  assign n35419 = ~n32852 & n35418 ;
  assign n35420 = ~\core_dag_ilm1reg_DMA_pi_DO_reg[9]/NET0131  & ~n35418 ;
  assign n35421 = ~n35419 & ~n35420 ;
  assign n35422 = ~n32898 & n35418 ;
  assign n35423 = ~\core_dag_ilm1reg_DMA_pi_DO_reg[8]/NET0131  & ~n35418 ;
  assign n35424 = ~n35422 & ~n35423 ;
  assign n35425 = ~n32806 & n35418 ;
  assign n35426 = ~\core_dag_ilm1reg_DMA_pi_DO_reg[7]/NET0131  & ~n35418 ;
  assign n35427 = ~n35425 & ~n35426 ;
  assign n35428 = ~n32829 & n35418 ;
  assign n35429 = ~\core_dag_ilm1reg_DMA_pi_DO_reg[6]/NET0131  & ~n35418 ;
  assign n35430 = ~n35428 & ~n35429 ;
  assign n35431 = ~n32783 & n35418 ;
  assign n35432 = ~\core_dag_ilm1reg_DMA_pi_DO_reg[5]/NET0131  & ~n35418 ;
  assign n35433 = ~n35431 & ~n35432 ;
  assign n35435 = ~n9752 & ~n32048 ;
  assign n35434 = ~n10302 & n32048 ;
  assign n35436 = n32054 & ~n35434 ;
  assign n35437 = ~n35435 & n35436 ;
  assign n35439 = ~n9767 & ~n32048 ;
  assign n35438 = ~n9805 & n32058 ;
  assign n35440 = ~n9790 & ~n35438 ;
  assign n35441 = ~n32054 & n35440 ;
  assign n35442 = ~n35439 & n35441 ;
  assign n35443 = ~n35437 & ~n35442 ;
  assign n35444 = ~n32068 & ~n35443 ;
  assign n35446 = ~n9786 & n32048 ;
  assign n35445 = ~n9733 & ~n32048 ;
  assign n35447 = ~n32054 & ~n35445 ;
  assign n35448 = ~n35446 & n35447 ;
  assign n35450 = n10069 & n32048 ;
  assign n35449 = n10289 & ~n32048 ;
  assign n35451 = n32054 & ~n35449 ;
  assign n35452 = ~n35450 & n35451 ;
  assign n35453 = ~n35448 & ~n35452 ;
  assign n35454 = n32068 & ~n35453 ;
  assign n35455 = ~n35444 & ~n35454 ;
  assign n35456 = n35418 & ~n35455 ;
  assign n35457 = ~\core_dag_ilm1reg_DMA_pi_DO_reg[4]/NET0131  & ~n35418 ;
  assign n35458 = ~n35456 & ~n35457 ;
  assign n35460 = ~n8224 & n32048 ;
  assign n35459 = ~n7644 & ~n32048 ;
  assign n35461 = n32054 & ~n35459 ;
  assign n35462 = ~n35460 & n35461 ;
  assign n35464 = ~n9695 & ~n32048 ;
  assign n35463 = ~n9666 & n32058 ;
  assign n35465 = ~n9700 & ~n35463 ;
  assign n35466 = ~n32054 & n35465 ;
  assign n35467 = ~n35464 & n35466 ;
  assign n35468 = ~n35462 & ~n35467 ;
  assign n35469 = ~n32068 & ~n35468 ;
  assign n35471 = ~n8190 & n32048 ;
  assign n35470 = ~n8149 & ~n32048 ;
  assign n35472 = ~n32054 & ~n35470 ;
  assign n35473 = ~n35471 & n35472 ;
  assign n35475 = n8113 & n32048 ;
  assign n35474 = n7859 & ~n32048 ;
  assign n35476 = n32054 & ~n35474 ;
  assign n35477 = ~n35475 & n35476 ;
  assign n35478 = ~n35473 & ~n35477 ;
  assign n35479 = n32068 & ~n35478 ;
  assign n35480 = ~n35469 & ~n35479 ;
  assign n35481 = n35418 & ~n35480 ;
  assign n35482 = ~\core_dag_ilm1reg_DMA_pi_DO_reg[3]/NET0131  & ~n35418 ;
  assign n35483 = ~n35481 & ~n35482 ;
  assign n35485 = ~n8246 & ~n32048 ;
  assign n35484 = ~n8794 & n32048 ;
  assign n35486 = n32054 & ~n35484 ;
  assign n35487 = ~n35485 & n35486 ;
  assign n35489 = ~n9625 & ~n32048 ;
  assign n35488 = ~n9600 & n32058 ;
  assign n35490 = ~n9633 & ~n35488 ;
  assign n35491 = ~n32054 & n35490 ;
  assign n35492 = ~n35489 & n35491 ;
  assign n35493 = ~n35487 & ~n35492 ;
  assign n35494 = ~n32068 & ~n35493 ;
  assign n35496 = ~n8773 & n32048 ;
  assign n35495 = ~n8750 & ~n32048 ;
  assign n35497 = ~n32054 & ~n35495 ;
  assign n35498 = ~n35496 & n35497 ;
  assign n35500 = n8715 & n32048 ;
  assign n35499 = n8460 & ~n32048 ;
  assign n35501 = n32054 & ~n35499 ;
  assign n35502 = ~n35500 & n35501 ;
  assign n35503 = ~n35498 & ~n35502 ;
  assign n35504 = n32068 & ~n35503 ;
  assign n35505 = ~n35494 & ~n35504 ;
  assign n35506 = n35418 & ~n35505 ;
  assign n35507 = ~\core_dag_ilm1reg_DMA_pi_DO_reg[2]/NET0131  & ~n35418 ;
  assign n35508 = ~n35506 & ~n35507 ;
  assign n35510 = ~n8962 & ~n32048 ;
  assign n35509 = ~n8926 & n32048 ;
  assign n35511 = n32054 & ~n35509 ;
  assign n35512 = ~n35510 & n35511 ;
  assign n35514 = ~n9559 & ~n32048 ;
  assign n35513 = ~n9528 & n32058 ;
  assign n35515 = ~n9567 & ~n35513 ;
  assign n35516 = ~n32054 & n35515 ;
  assign n35517 = ~n35514 & n35516 ;
  assign n35518 = ~n35512 & ~n35517 ;
  assign n35519 = ~n32068 & ~n35518 ;
  assign n35521 = ~n8903 & n32048 ;
  assign n35520 = ~n8873 & ~n32048 ;
  assign n35522 = ~n32054 & ~n35520 ;
  assign n35523 = ~n35521 & n35522 ;
  assign n35525 = n9435 & n32048 ;
  assign n35524 = n9178 & ~n32048 ;
  assign n35526 = n32054 & ~n35524 ;
  assign n35527 = ~n35525 & n35526 ;
  assign n35528 = ~n35523 & ~n35527 ;
  assign n35529 = n32068 & ~n35528 ;
  assign n35530 = ~n35519 & ~n35529 ;
  assign n35531 = n35418 & ~n35530 ;
  assign n35532 = ~\core_dag_ilm1reg_DMA_pi_DO_reg[1]/NET0131  & ~n35418 ;
  assign n35533 = ~n35531 & ~n35532 ;
  assign n35534 = \core_dag_ilm1reg_DMA_pi_DO_reg[13]/NET0131  & ~n35418 ;
  assign n35535 = ~n32080 & n35418 ;
  assign n35536 = ~n35534 & ~n35535 ;
  assign n35537 = ~n32921 & n35418 ;
  assign n35538 = ~\core_dag_ilm1reg_DMA_pi_DO_reg[12]/NET0131  & ~n35418 ;
  assign n35539 = ~n35537 & ~n35538 ;
  assign n35540 = ~n32944 & n35418 ;
  assign n35541 = ~\core_dag_ilm1reg_DMA_pi_DO_reg[11]/NET0131  & ~n35418 ;
  assign n35542 = ~n35540 & ~n35541 ;
  assign n35543 = ~n32875 & n35418 ;
  assign n35544 = ~\core_dag_ilm1reg_DMA_pi_DO_reg[10]/NET0131  & ~n35418 ;
  assign n35545 = ~n35543 & ~n35544 ;
  assign n35547 = ~n7622 & n32048 ;
  assign n35546 = ~n6546 & ~n32048 ;
  assign n35548 = n32054 & ~n35546 ;
  assign n35549 = ~n35547 & n35548 ;
  assign n35550 = ~n6911 & ~n32048 ;
  assign n35551 = ~n6980 & n32058 ;
  assign n35552 = ~n6957 & ~n35551 ;
  assign n35553 = ~n32054 & n35552 ;
  assign n35554 = ~n35550 & n35553 ;
  assign n35555 = ~n35549 & ~n35554 ;
  assign n35556 = ~n32068 & ~n35555 ;
  assign n35558 = ~n6951 & n32048 ;
  assign n35557 = ~n6158 & ~n32048 ;
  assign n35559 = ~n32054 & ~n35557 ;
  assign n35560 = ~n35558 & n35559 ;
  assign n35562 = n7607 & n32048 ;
  assign n35561 = n7340 & ~n32048 ;
  assign n35563 = n32054 & ~n35561 ;
  assign n35564 = ~n35562 & n35563 ;
  assign n35565 = ~n35560 & ~n35564 ;
  assign n35566 = n32068 & ~n35565 ;
  assign n35567 = ~n35556 & ~n35566 ;
  assign n35568 = n35418 & ~n35567 ;
  assign n35569 = ~\core_dag_ilm1reg_DMA_pi_DO_reg[0]/NET0131  & ~n35418 ;
  assign n35570 = ~n35568 & ~n35569 ;
  assign n35571 = \core_c_dec_MTMSTAT_Eg_reg/P0001  & n4118 ;
  assign n35572 = n23231 & n32022 ;
  assign n35573 = n31998 & n35572 ;
  assign n35574 = ~n35571 & ~n35573 ;
  assign n35575 = ~\bdma_BEAD_reg[7]/NET0131  & ~n33308 ;
  assign n35576 = ~n20765 & ~n33309 ;
  assign n35577 = ~n35575 & n35576 ;
  assign n35578 = n11265 & n20765 ;
  assign n35579 = ~n35577 & ~n35578 ;
  assign n35580 = ~\bdma_BEAD_reg[6]/NET0131  & ~n33307 ;
  assign n35581 = ~n20765 & ~n33308 ;
  assign n35582 = ~n35580 & n35581 ;
  assign n35583 = n11525 & n20765 ;
  assign n35584 = ~n35582 & ~n35583 ;
  assign n35585 = ~\bdma_BEAD_reg[5]/NET0131  & ~n33306 ;
  assign n35586 = ~n20765 & ~n33307 ;
  assign n35587 = ~n35585 & n35586 ;
  assign n35588 = n10911 & n20765 ;
  assign n35589 = ~n35587 & ~n35588 ;
  assign n35590 = \sport1_regs_FSDIVreg_DO_reg[0]/NET0131  & n28786 ;
  assign n35591 = ~\sport1_cfg_FSi_cnt_reg[0]/NET0131  & ~\sport1_cfg_SP_ENg_reg/NET0131  ;
  assign n35592 = ~n28856 & ~n35591 ;
  assign n35593 = n28855 & n35592 ;
  assign n35594 = ~n35590 & ~n35593 ;
  assign n35595 = \sport0_regs_FSDIVreg_DO_reg[0]/NET0131  & n28876 ;
  assign n35596 = ~\sport0_cfg_FSi_cnt_reg[0]/NET0131  & ~\sport0_cfg_SP_ENg_reg/NET0131  ;
  assign n35597 = ~n28946 & ~n35596 ;
  assign n35598 = n28945 & n35597 ;
  assign n35599 = ~n35595 & ~n35598 ;
  assign n35600 = n14752 & ~n25088 ;
  assign n35601 = ~\core_eu_em_mac_em_reg_mr2rwe_DO_reg[0]/P0001  & ~n17799 ;
  assign n35602 = ~n17809 & n19559 ;
  assign n35603 = n17811 & ~n35602 ;
  assign n35604 = ~n35601 & ~n35603 ;
  assign n35605 = ~n17823 & ~n35604 ;
  assign n35606 = ~\core_eu_em_mac_em_reg_mr2rwe_DO_reg[0]/P0001  & ~n17808 ;
  assign n35607 = ~n35605 & ~n35606 ;
  assign n35608 = n17829 & ~n35607 ;
  assign n35609 = ~n35600 & ~n35608 ;
  assign n35610 = ~\sice_ICYC_reg[23]/NET0131  & ~n20785 ;
  assign n35611 = ~n32035 & ~n35610 ;
  assign n35612 = \core_c_dec_MTtoppcs_Eg_reg/P0001  & n4118 ;
  assign n35613 = n23231 & n32010 ;
  assign n35614 = ~n35612 & ~n35613 ;
  assign n35615 = \sport0_regs_FSDIVreg_DO_reg[1]/NET0131  & n28876 ;
  assign n35616 = ~\sport0_cfg_FSi_cnt_reg[1]/NET0131  & ~n28946 ;
  assign n35617 = ~n28947 & ~n35616 ;
  assign n35618 = n28945 & n35617 ;
  assign n35619 = ~n35615 & ~n35618 ;
  assign n35620 = \sport1_regs_FSDIVreg_DO_reg[1]/NET0131  & n28786 ;
  assign n35621 = ~\sport1_cfg_FSi_cnt_reg[1]/NET0131  & ~n28856 ;
  assign n35622 = ~n28857 & ~n35621 ;
  assign n35623 = n28855 & n35622 ;
  assign n35624 = ~n35620 & ~n35623 ;
  assign n35625 = \sport1_regs_FSDIVreg_DO_reg[2]/NET0131  & n28786 ;
  assign n35626 = ~\sport1_cfg_FSi_cnt_reg[2]/NET0131  & ~n28857 ;
  assign n35627 = ~n28858 & ~n35626 ;
  assign n35628 = n28855 & n35627 ;
  assign n35629 = ~n35625 & ~n35628 ;
  assign n35630 = \sport1_regs_FSDIVreg_DO_reg[5]/NET0131  & n28786 ;
  assign n35631 = ~\sport1_cfg_FSi_cnt_reg[5]/NET0131  & ~n28860 ;
  assign n35632 = ~n28861 & ~n35631 ;
  assign n35633 = n28855 & n35632 ;
  assign n35634 = ~n35630 & ~n35633 ;
  assign n35635 = \sport1_regs_FSDIVreg_DO_reg[9]/NET0131  & n28786 ;
  assign n35636 = ~\sport1_cfg_FSi_cnt_reg[9]/NET0131  & ~n28864 ;
  assign n35637 = n28855 & ~n28865 ;
  assign n35638 = ~n35636 & n35637 ;
  assign n35639 = ~n35635 & ~n35638 ;
  assign n35640 = \sport0_regs_FSDIVreg_DO_reg[13]/NET0131  & n28876 ;
  assign n35641 = ~\sport0_cfg_FSi_cnt_reg[13]/NET0131  & ~n28958 ;
  assign n35642 = n28945 & ~n28959 ;
  assign n35643 = ~n35641 & n35642 ;
  assign n35644 = ~n35640 & ~n35643 ;
  assign n35645 = \sport0_regs_FSDIVreg_DO_reg[2]/NET0131  & n28876 ;
  assign n35646 = ~\sport0_cfg_FSi_cnt_reg[2]/NET0131  & ~n28947 ;
  assign n35647 = ~n28948 & ~n35646 ;
  assign n35648 = n28945 & n35647 ;
  assign n35649 = ~n35645 & ~n35648 ;
  assign n35650 = \sport0_regs_FSDIVreg_DO_reg[5]/NET0131  & n28876 ;
  assign n35651 = ~\sport0_cfg_FSi_cnt_reg[5]/NET0131  & ~n28950 ;
  assign n35652 = ~n28951 & ~n35651 ;
  assign n35653 = n28945 & n35652 ;
  assign n35654 = ~n35650 & ~n35653 ;
  assign n35655 = ~\sice_ICYC_reg[4]/NET0131  & ~n18858 ;
  assign n35656 = ~n18859 & ~n35655 ;
  assign n35657 = \sport0_regs_FSDIVreg_DO_reg[9]/NET0131  & n28876 ;
  assign n35658 = ~\sport0_cfg_FSi_cnt_reg[9]/NET0131  & ~n28954 ;
  assign n35659 = n28945 & ~n28955 ;
  assign n35660 = ~n35658 & n35659 ;
  assign n35661 = ~n35657 & ~n35660 ;
  assign n35662 = ~\clkc_oscntr_reg_DO_reg[4]/NET0131  & ~n23417 ;
  assign n35663 = ~n23418 & ~n35662 ;
  assign n35664 = ~\sice_IIRC_reg[4]/NET0131  & ~n18867 ;
  assign n35665 = ~n18868 & ~n35664 ;
  assign n35666 = \sport1_regs_FSDIVreg_DO_reg[13]/NET0131  & n28786 ;
  assign n35667 = ~\sport1_cfg_FSi_cnt_reg[13]/NET0131  & ~n28868 ;
  assign n35668 = n28855 & ~n28869 ;
  assign n35669 = ~n35667 & n35668 ;
  assign n35670 = ~n35666 & ~n35669 ;
  assign n35671 = n26967 & n34841 ;
  assign n35672 = \sice_IRR_reg[4]/P0001  & ~n35671 ;
  assign n35673 = \sice_SPC_reg[14]/P0001  & n35671 ;
  assign n35674 = ~n35672 & ~n35673 ;
  assign n35675 = n4093 & ~n35674 ;
  assign n35676 = \core_c_psq_EXA_reg[4]/P0001  & ~n4093 ;
  assign n35677 = ~n35675 & ~n35676 ;
  assign n35678 = \sice_IRR_reg[9]/P0001  & ~n35671 ;
  assign n35679 = \sice_SPC_reg[19]/P0001  & n35671 ;
  assign n35680 = ~n35678 & ~n35679 ;
  assign n35681 = n4093 & ~n35680 ;
  assign n35682 = \core_c_psq_EXA_reg[9]/P0001  & ~n4093 ;
  assign n35683 = ~n35681 & ~n35682 ;
  assign n35684 = \sice_IRR_reg[8]/P0001  & ~n35671 ;
  assign n35685 = \sice_SPC_reg[18]/P0001  & n35671 ;
  assign n35686 = ~n35684 & ~n35685 ;
  assign n35687 = n4093 & ~n35686 ;
  assign n35688 = \core_c_psq_EXA_reg[8]/P0001  & ~n4093 ;
  assign n35689 = ~n35687 & ~n35688 ;
  assign n35690 = \sice_IRR_reg[7]/P0001  & ~n35671 ;
  assign n35691 = \sice_SPC_reg[17]/P0001  & n35671 ;
  assign n35692 = ~n35690 & ~n35691 ;
  assign n35693 = n4093 & ~n35692 ;
  assign n35694 = \core_c_psq_EXA_reg[7]/P0001  & ~n4093 ;
  assign n35695 = ~n35693 & ~n35694 ;
  assign n35696 = \sice_IRR_reg[6]/P0001  & ~n35671 ;
  assign n35697 = \sice_SPC_reg[16]/P0001  & n35671 ;
  assign n35698 = ~n35696 & ~n35697 ;
  assign n35699 = n4093 & ~n35698 ;
  assign n35700 = \core_c_psq_EXA_reg[6]/P0001  & ~n4093 ;
  assign n35701 = ~n35699 & ~n35700 ;
  assign n35702 = \sice_IRR_reg[5]/P0001  & ~n35671 ;
  assign n35703 = \sice_SPC_reg[15]/P0001  & n35671 ;
  assign n35704 = ~n35702 & ~n35703 ;
  assign n35705 = n4093 & ~n35704 ;
  assign n35706 = \core_c_psq_EXA_reg[5]/P0001  & ~n4093 ;
  assign n35707 = ~n35705 & ~n35706 ;
  assign n35708 = \sice_IRR_reg[3]/P0001  & ~n35671 ;
  assign n35709 = \sice_SPC_reg[13]/P0001  & n35671 ;
  assign n35710 = ~n35708 & ~n35709 ;
  assign n35711 = n4093 & ~n35710 ;
  assign n35712 = \core_c_psq_EXA_reg[3]/P0001  & ~n4093 ;
  assign n35713 = ~n35711 & ~n35712 ;
  assign n35714 = \sice_IRR_reg[2]/P0001  & ~n35671 ;
  assign n35715 = \sice_SPC_reg[12]/P0001  & n35671 ;
  assign n35716 = ~n35714 & ~n35715 ;
  assign n35717 = n4093 & ~n35716 ;
  assign n35718 = \core_c_psq_EXA_reg[2]/P0001  & ~n4093 ;
  assign n35719 = ~n35717 & ~n35718 ;
  assign n35720 = \sice_IRR_reg[13]/P0001  & ~n35671 ;
  assign n35721 = \sice_SPC_reg[23]/P0001  & n35671 ;
  assign n35722 = ~n35720 & ~n35721 ;
  assign n35723 = n4093 & ~n35722 ;
  assign n35724 = \core_c_psq_EXA_reg[13]/P0001  & ~n4093 ;
  assign n35725 = ~n35723 & ~n35724 ;
  assign n35726 = \sice_IRR_reg[1]/P0001  & ~n35671 ;
  assign n35727 = \sice_SPC_reg[11]/P0001  & n35671 ;
  assign n35728 = ~n35726 & ~n35727 ;
  assign n35729 = n4093 & ~n35728 ;
  assign n35730 = \core_c_psq_EXA_reg[1]/P0001  & ~n4093 ;
  assign n35731 = ~n35729 & ~n35730 ;
  assign n35732 = \sice_IRR_reg[12]/P0001  & ~n35671 ;
  assign n35733 = \sice_SPC_reg[22]/P0001  & n35671 ;
  assign n35734 = ~n35732 & ~n35733 ;
  assign n35735 = n4093 & ~n35734 ;
  assign n35736 = \core_c_psq_EXA_reg[12]/P0001  & ~n4093 ;
  assign n35737 = ~n35735 & ~n35736 ;
  assign n35738 = \sice_IRR_reg[11]/P0001  & ~n35671 ;
  assign n35739 = \sice_SPC_reg[21]/P0001  & n35671 ;
  assign n35740 = ~n35738 & ~n35739 ;
  assign n35741 = n4093 & ~n35740 ;
  assign n35742 = \core_c_psq_EXA_reg[11]/P0001  & ~n4093 ;
  assign n35743 = ~n35741 & ~n35742 ;
  assign n35744 = \sice_IRR_reg[10]/P0001  & ~n35671 ;
  assign n35745 = \sice_SPC_reg[20]/P0001  & n35671 ;
  assign n35746 = ~n35744 & ~n35745 ;
  assign n35747 = n4093 & ~n35746 ;
  assign n35748 = \core_c_psq_EXA_reg[10]/P0001  & ~n4093 ;
  assign n35749 = ~n35747 & ~n35748 ;
  assign n35750 = \sice_IRR_reg[0]/P0001  & ~n35671 ;
  assign n35751 = \sice_SPC_reg[10]/P0001  & n35671 ;
  assign n35752 = ~n35750 & ~n35751 ;
  assign n35753 = n4093 & ~n35752 ;
  assign n35754 = \core_c_psq_EXA_reg[0]/P0001  & ~n4093 ;
  assign n35755 = ~n35753 & ~n35754 ;
  assign n35756 = n31264 & n34029 ;
  assign n35757 = ~n4117 & n31271 ;
  assign n35758 = n35756 & n35757 ;
  assign n35759 = \core_c_dec_MFICNTL_E_reg/P0001  & n4117 ;
  assign n35760 = ~n35758 & ~n35759 ;
  assign n35761 = \sport0_txctl_TXSHT_reg[13]/P0001  & ~n19960 ;
  assign n35762 = \sport0_txctl_TX_reg[14]/P0001  & n19960 ;
  assign n35763 = ~n35761 & ~n35762 ;
  assign n35764 = \sport0_txctl_TXSHT_reg[9]/P0001  & ~n19960 ;
  assign n35765 = \sport0_txctl_TX_reg[10]/P0001  & n19960 ;
  assign n35766 = ~n35764 & ~n35765 ;
  assign n35767 = \sport0_txctl_TXSHT_reg[8]/P0001  & ~n19960 ;
  assign n35768 = \sport0_txctl_TX_reg[9]/P0001  & n19960 ;
  assign n35769 = ~n35767 & ~n35768 ;
  assign n35770 = \sport0_txctl_TXSHT_reg[7]/P0001  & ~n19960 ;
  assign n35771 = \sport0_txctl_TX_reg[8]/P0001  & n19960 ;
  assign n35772 = ~n35770 & ~n35771 ;
  assign n35773 = \sport1_txctl_TXSHT_reg[8]/P0001  & ~n22677 ;
  assign n35774 = \sport1_txctl_TX_reg[9]/P0001  & n22677 ;
  assign n35775 = ~n35773 & ~n35774 ;
  assign n35776 = \sport0_txctl_TXSHT_reg[5]/P0001  & ~n19960 ;
  assign n35777 = \sport0_txctl_TX_reg[6]/P0001  & n19960 ;
  assign n35778 = ~n35776 & ~n35777 ;
  assign n35779 = \sport1_txctl_TXSHT_reg[7]/P0001  & ~n22677 ;
  assign n35780 = \sport1_txctl_TX_reg[8]/P0001  & n22677 ;
  assign n35781 = ~n35779 & ~n35780 ;
  assign n35782 = ~\sice_ICYC_reg[15]/NET0131  & ~n20744 ;
  assign n35783 = ~n20745 & ~n35782 ;
  assign n35784 = \sport0_txctl_TXSHT_reg[4]/P0001  & ~n19960 ;
  assign n35785 = \sport0_txctl_TX_reg[5]/P0001  & n19960 ;
  assign n35786 = ~n35784 & ~n35785 ;
  assign n35787 = ~\sice_IIRC_reg[15]/NET0131  & ~n20859 ;
  assign n35788 = ~n22581 & ~n35787 ;
  assign n35789 = \sport1_txctl_TXSHT_reg[5]/P0001  & ~n22677 ;
  assign n35790 = \sport1_txctl_TX_reg[6]/P0001  & n22677 ;
  assign n35791 = ~n35789 & ~n35790 ;
  assign n35792 = \sport1_txctl_TXSHT_reg[4]/P0001  & ~n22677 ;
  assign n35793 = \sport1_txctl_TX_reg[5]/P0001  & n22677 ;
  assign n35794 = ~n35792 & ~n35793 ;
  assign n35795 = \sport0_txctl_TXSHT_reg[2]/P0001  & ~n19960 ;
  assign n35796 = \sport0_txctl_TX_reg[3]/P0001  & n19960 ;
  assign n35797 = ~n35795 & ~n35796 ;
  assign n35798 = \sice_ICYC_reg[0]/NET0131  & ~n32036 ;
  assign n35799 = ~\sice_ICYC_reg[0]/NET0131  & n32036 ;
  assign n35800 = ~n35798 & ~n35799 ;
  assign n35801 = \sice_SPC_reg[5]/P0001  & ~n26297 ;
  assign n35806 = \core_c_dec_IR_reg[5]/NET0131  & n28203 ;
  assign n35807 = \sice_DBR2_reg[0]/P0001  & n25012 ;
  assign n35812 = ~n35806 & ~n35807 ;
  assign n35808 = \sice_ICYC_reg[5]/NET0131  & n23409 ;
  assign n35809 = \sice_idr0_reg_DO_reg[5]/P0001  & n26968 ;
  assign n35813 = ~n35808 & ~n35809 ;
  assign n35810 = \sice_IIRC_reg[5]/NET0131  & n24267 ;
  assign n35811 = \sice_DBR1_reg[0]/P0001  & n25054 ;
  assign n35814 = ~n35810 & ~n35811 ;
  assign n35815 = n35813 & n35814 ;
  assign n35816 = n35812 & n35815 ;
  assign n35817 = n34827 & n35816 ;
  assign n35802 = \sice_SPC_reg[4]/P0001  & n34825 ;
  assign n35803 = \sice_SPC_reg[6]/P0001  & ~n34825 ;
  assign n35804 = ~n35802 & ~n35803 ;
  assign n35805 = ~n34827 & n35804 ;
  assign n35818 = n26297 & ~n35805 ;
  assign n35819 = ~n35817 & n35818 ;
  assign n35820 = ~n35801 & ~n35819 ;
  assign n35821 = \sice_SPC_reg[8]/P0001  & n34825 ;
  assign n35822 = \sice_SPC_reg[10]/P0001  & ~n34825 ;
  assign n35823 = ~n35821 & ~n35822 ;
  assign n35824 = ~n34827 & n35823 ;
  assign n35833 = \sice_DBR1_reg[4]/P0001  & n25054 ;
  assign n35834 = \sice_idr0_reg_DO_reg[9]/P0001  & n26968 ;
  assign n35841 = ~n35833 & ~n35834 ;
  assign n35835 = \sice_DMR1_reg[3]/NET0131  & n27903 ;
  assign n35836 = \sice_ICYC_reg[9]/NET0131  & n23409 ;
  assign n35842 = ~n35835 & ~n35836 ;
  assign n35843 = n35841 & n35842 ;
  assign n35829 = \sice_DMR2_reg[3]/NET0131  & n25025 ;
  assign n35830 = \sice_IBR1_reg[3]/P0001  & n34831 ;
  assign n35839 = ~n35829 & ~n35830 ;
  assign n35831 = \sice_IIRC_reg[9]/NET0131  & n24267 ;
  assign n35832 = \sice_IMR2_reg[3]/NET0131  & n25034 ;
  assign n35840 = ~n35831 & ~n35832 ;
  assign n35844 = n35839 & n35840 ;
  assign n35825 = \core_c_dec_IR_reg[9]/NET0131  & n28203 ;
  assign n35826 = \sice_DBR2_reg[4]/P0001  & n25012 ;
  assign n35837 = ~n35825 & ~n35826 ;
  assign n35827 = \sice_IBR2_reg[3]/P0001  & n25074 ;
  assign n35828 = \sice_IMR1_reg[3]/NET0131  & n34846 ;
  assign n35838 = ~n35827 & ~n35828 ;
  assign n35845 = n35837 & n35838 ;
  assign n35846 = n35844 & n35845 ;
  assign n35847 = n35843 & n35846 ;
  assign n35848 = n34827 & n35847 ;
  assign n35849 = ~n35824 & ~n35848 ;
  assign n35850 = \sport0_txctl_TXSHT_reg[1]/P0001  & ~n19960 ;
  assign n35851 = \sport0_txctl_TX_reg[2]/P0001  & n19960 ;
  assign n35852 = ~n35850 & ~n35851 ;
  assign n35853 = \sice_SPC_reg[5]/P0001  & n34825 ;
  assign n35854 = \sice_SPC_reg[7]/P0001  & ~n34825 ;
  assign n35855 = ~n35853 & ~n35854 ;
  assign n35856 = ~n34827 & n35855 ;
  assign n35865 = \sice_IBR2_reg[0]/P0001  & n25074 ;
  assign n35866 = \sice_idr0_reg_DO_reg[6]/P0001  & n26968 ;
  assign n35873 = ~n35865 & ~n35866 ;
  assign n35867 = \sice_DBR2_reg[1]/P0001  & n25012 ;
  assign n35868 = \sice_ICYC_reg[6]/NET0131  & n23409 ;
  assign n35874 = ~n35867 & ~n35868 ;
  assign n35875 = n35873 & n35874 ;
  assign n35861 = \sice_IMR2_reg[0]/NET0131  & n25034 ;
  assign n35862 = \sice_IBR1_reg[0]/P0001  & n34831 ;
  assign n35871 = ~n35861 & ~n35862 ;
  assign n35863 = \sice_IIRC_reg[6]/NET0131  & n24267 ;
  assign n35864 = \sice_IMR1_reg[0]/NET0131  & n34846 ;
  assign n35872 = ~n35863 & ~n35864 ;
  assign n35876 = n35871 & n35872 ;
  assign n35857 = \core_c_dec_IR_reg[6]/NET0131  & n28203 ;
  assign n35858 = \sice_DMR1_reg[0]/NET0131  & n27903 ;
  assign n35869 = ~n35857 & ~n35858 ;
  assign n35859 = \sice_DMR2_reg[0]/NET0131  & n25025 ;
  assign n35860 = \sice_DBR1_reg[1]/P0001  & n25054 ;
  assign n35870 = ~n35859 & ~n35860 ;
  assign n35877 = n35869 & n35870 ;
  assign n35878 = n35876 & n35877 ;
  assign n35879 = n35875 & n35878 ;
  assign n35880 = n34827 & n35879 ;
  assign n35881 = ~n35856 & ~n35880 ;
  assign n35882 = \sport0_txctl_TXSHT_reg[0]/P0001  & ~n19960 ;
  assign n35883 = \sport0_txctl_TX_reg[1]/P0001  & n19960 ;
  assign n35884 = ~n35882 & ~n35883 ;
  assign n35885 = \sport1_txctl_TXSHT_reg[2]/P0001  & ~n22677 ;
  assign n35886 = \sport1_txctl_TX_reg[3]/P0001  & n22677 ;
  assign n35887 = ~n35885 & ~n35886 ;
  assign n35888 = \sport1_txctl_TXSHT_reg[1]/P0001  & ~n22677 ;
  assign n35889 = \sport1_txctl_TX_reg[2]/P0001  & n22677 ;
  assign n35890 = ~n35888 & ~n35889 ;
  assign n35891 = n18262 & n31574 ;
  assign n35892 = ~\core_eu_em_mac_em_reg_mr2swe_DO_reg[3]/P0001  & ~n28530 ;
  assign n35893 = ~n19381 & n21663 ;
  assign n35894 = n28534 & ~n35893 ;
  assign n35895 = ~n35892 & ~n35894 ;
  assign n35896 = ~n19385 & ~n35895 ;
  assign n35897 = ~\core_eu_em_mac_em_reg_mr2swe_DO_reg[3]/P0001  & ~n28532 ;
  assign n35898 = ~n35896 & ~n35897 ;
  assign n35899 = n28529 & ~n35898 ;
  assign n35900 = ~n35891 & ~n35899 ;
  assign n35901 = \sport0_txctl_TX_reg[0]/P0001  & n19960 ;
  assign n35902 = \sport1_txctl_TXSHT_reg[0]/P0001  & ~n22677 ;
  assign n35903 = \sport1_txctl_TX_reg[1]/P0001  & n22677 ;
  assign n35904 = ~n35902 & ~n35903 ;
  assign n35906 = ~n5582 & ~n20208 ;
  assign n35907 = n12442 & ~n35906 ;
  assign n35905 = \memc_Pwrite_E_reg/NET0131  & ~n5607 ;
  assign n35908 = \memc_Dwrite_E_reg/NET0131  & ~n5600 ;
  assign n35909 = ~n35905 & ~n35908 ;
  assign n35910 = ~n35907 & n35909 ;
  assign n35911 = ~n5581 & ~n5597 ;
  assign n35912 = n5560 & n35911 ;
  assign n35913 = n5586 & n35912 ;
  assign n35914 = \bdma_BCTL_reg[2]/NET0131  & n35913 ;
  assign n35916 = ~n12442 & n20208 ;
  assign n35917 = \memc_Pread_E_reg/NET0131  & n5606 ;
  assign n35915 = n5599 & ~n14732 ;
  assign n35918 = ~n35913 & ~n35915 ;
  assign n35919 = ~n35917 & n35918 ;
  assign n35920 = ~n35916 & n35919 ;
  assign n35921 = ~n35914 & ~n35920 ;
  assign n35922 = n12442 & n20208 ;
  assign n35923 = \memc_Pwrite_E_reg/NET0131  & n5606 ;
  assign n35924 = \memc_Dwrite_E_reg/NET0131  & n5599 ;
  assign n35925 = ~n35923 & ~n35924 ;
  assign n35926 = ~n35922 & n35925 ;
  assign n35927 = \sport1_txctl_TX_reg[0]/P0001  & n22677 ;
  assign n35928 = ~n5556 & ~n35912 ;
  assign n35929 = \core_c_psq_PCS_reg[12]/NET0131  & ~\emc_eRDY_reg/NET0131  ;
  assign n35930 = \core_c_psq_PCS_reg[1]/NET0131  & ~n4068 ;
  assign n35931 = ~n35929 & ~n35930 ;
  assign n35932 = n5700 & n35931 ;
  assign n35933 = ~\core_c_psq_PCS_reg[3]/NET0131  & ~n35932 ;
  assign n35934 = n19047 & ~n35933 ;
  assign n35935 = n4118 & ~n35934 ;
  assign n35936 = \core_c_dec_MTSR0_E_reg/P0001  & ~n19504 ;
  assign n35937 = ~\core_c_dec_MTSR0_E_reg/P0001  & n29555 ;
  assign n35938 = ~n35936 & ~n35937 ;
  assign n35939 = n18886 & ~n35938 ;
  assign n35940 = ~\core_eu_es_sht_es_reg_sr0swe_DO_reg[9]/P0001  & ~n18886 ;
  assign n35941 = ~n35939 & ~n35940 ;
  assign n35942 = n19034 & ~n35938 ;
  assign n35943 = ~\core_eu_es_sht_es_reg_sr0rwe_DO_reg[9]/P0001  & ~n19034 ;
  assign n35944 = ~n35942 & ~n35943 ;
  assign n35945 = n18513 & ~n23044 ;
  assign n35946 = n18471 & ~n35945 ;
  assign n35948 = \sport0_regs_SCTLreg_DO_reg[4]/NET0131  & n35946 ;
  assign n35947 = ~\sport0_regs_SCTLreg_DO_reg[4]/NET0131  & ~n35946 ;
  assign n35949 = \sport0_txctl_ldTX_cmp_reg/P0001  & ~n35947 ;
  assign n35950 = ~n35948 & n35949 ;
  assign n35952 = ~n10911 & ~n18519 ;
  assign n35951 = ~\sport0_txctl_TX_reg[5]/P0001  & n18519 ;
  assign n35953 = ~\sport0_txctl_ldTX_cmp_reg/P0001  & ~n35951 ;
  assign n35954 = ~n35952 & n35953 ;
  assign n35955 = ~n35950 & ~n35954 ;
  assign n35956 = \ISCLK0_pad  & \sport0_cfg_SCLKi_h_reg/NET0131  ;
  assign n35958 = \T_SCLK0_pad  & \sport0_regs_SCTLreg_DO_reg[13]/NET0131  ;
  assign n35957 = ~\T_SCLK0_pad  & ~\sport0_regs_SCTLreg_DO_reg[13]/NET0131  ;
  assign n35959 = ~\ISCLK0_pad  & ~n35957 ;
  assign n35960 = ~n35958 & n35959 ;
  assign n35961 = ~n35956 & ~n35960 ;
  assign n35962 = \ISCLK1_pad  & \sport1_cfg_SCLKi_h_reg/NET0131  ;
  assign n35964 = \T_SCLK1_pad  & \sport1_regs_SCTLreg_DO_reg[13]/NET0131  ;
  assign n35963 = ~\T_SCLK1_pad  & ~\sport1_regs_SCTLreg_DO_reg[13]/NET0131  ;
  assign n35965 = ~\ISCLK1_pad  & ~n35963 ;
  assign n35966 = ~n35964 & n35965 ;
  assign n35967 = ~n35962 & ~n35966 ;
  assign n35968 = \core_c_dec_MTSR1_E_reg/P0001  & ~n23860 ;
  assign n35969 = ~\core_c_dec_MTSR1_E_reg/P0001  & n30392 ;
  assign n35970 = ~n35968 & ~n35969 ;
  assign n35971 = n18717 & ~n35970 ;
  assign n35972 = ~\core_eu_es_sht_es_reg_sr1swe_DO_reg[8]/P0001  & ~n18717 ;
  assign n35973 = ~n35971 & ~n35972 ;
  assign n35974 = ~n13806 & ~n19222 ;
  assign n35975 = n13806 & n14540 ;
  assign n35976 = ~n35974 & ~n35975 ;
  assign n35977 = n14667 & ~n35976 ;
  assign n35978 = \core_eu_ea_alu_ea_reg_afswe_DO_reg[15]/P0001  & ~n14667 ;
  assign n35979 = ~n35977 & ~n35978 ;
  assign n35980 = n13805 & ~n35976 ;
  assign n35981 = \core_eu_ea_alu_ea_reg_afrwe_DO_reg[15]/P0001  & ~n13805 ;
  assign n35982 = ~n35980 & ~n35981 ;
  assign n35983 = \core_c_dec_MTSR1_E_reg/P0001  & ~n23757 ;
  assign n35984 = ~\core_c_dec_MTSR1_E_reg/P0001  & n29839 ;
  assign n35985 = ~n35983 & ~n35984 ;
  assign n35986 = n18717 & ~n35985 ;
  assign n35987 = ~\core_eu_es_sht_es_reg_sr1swe_DO_reg[11]/P0001  & ~n18717 ;
  assign n35988 = ~n35986 & ~n35987 ;
  assign n35989 = n17833 & ~n35970 ;
  assign n35990 = ~\core_eu_es_sht_es_reg_sr1rwe_DO_reg[8]/P0001  & ~n17833 ;
  assign n35991 = ~n35989 & ~n35990 ;
  assign n35992 = n17833 & ~n35985 ;
  assign n35993 = ~\core_eu_es_sht_es_reg_sr1rwe_DO_reg[11]/P0001  & ~n17833 ;
  assign n35994 = ~n35992 & ~n35993 ;
  assign n35995 = \core_c_dec_MTSR0_E_reg/P0001  & ~n17820 ;
  assign n35996 = ~\core_c_dec_MTSR0_E_reg/P0001  & n29285 ;
  assign n35997 = ~n35995 & ~n35996 ;
  assign n35998 = n18886 & ~n35997 ;
  assign n35999 = ~\core_eu_es_sht_es_reg_sr0swe_DO_reg[15]/P0001  & ~n18886 ;
  assign n36000 = ~n35998 & ~n35999 ;
  assign n36002 = \sport0_txctl_Bcnt_reg[3]/NET0131  & ~n19956 ;
  assign n36003 = ~n19957 & ~n36002 ;
  assign n36004 = n23277 & ~n36003 ;
  assign n36001 = \sport0_regs_SCTLreg_DO_reg[3]/NET0131  & ~n23277 ;
  assign n36005 = ~\sport0_rxctl_TAG_SLOT_reg/P0001  & ~n36001 ;
  assign n36006 = ~n36004 & n36005 ;
  assign n36008 = \sport1_txctl_Bcnt_reg[3]/NET0131  & ~n22673 ;
  assign n36009 = ~n22674 & ~n36008 ;
  assign n36010 = n23265 & ~n36009 ;
  assign n36007 = \sport1_regs_SCTLreg_DO_reg[3]/NET0131  & ~n23265 ;
  assign n36011 = ~\sport1_rxctl_TAG_SLOT_reg/P0001  & ~n36007 ;
  assign n36012 = ~n36010 & n36011 ;
  assign n36014 = \sport1_txctl_Bcnt_reg[2]/NET0131  & ~n22672 ;
  assign n36015 = ~n22673 & ~n36014 ;
  assign n36016 = n23265 & ~n36015 ;
  assign n36013 = \sport1_regs_SCTLreg_DO_reg[2]/NET0131  & ~n23265 ;
  assign n36017 = ~\sport1_rxctl_TAG_SLOT_reg/P0001  & ~n36013 ;
  assign n36018 = ~n36016 & n36017 ;
  assign n36019 = n19034 & ~n35997 ;
  assign n36020 = ~\core_eu_es_sht_es_reg_sr0rwe_DO_reg[15]/P0001  & ~n19034 ;
  assign n36021 = ~n36019 & ~n36020 ;
  assign n36023 = \sport1_txctl_Bcnt_reg[0]/NET0131  & \sport1_txctl_Bcnt_reg[1]/NET0131  ;
  assign n36024 = ~n22672 & ~n36023 ;
  assign n36025 = n23265 & ~n36024 ;
  assign n36022 = \sport1_regs_SCTLreg_DO_reg[1]/NET0131  & ~n23265 ;
  assign n36026 = ~\sport1_rxctl_TAG_SLOT_reg/P0001  & ~n36022 ;
  assign n36027 = ~n36025 & n36026 ;
  assign n36028 = ~T_IRDn_pad & ~T_ISn_pad ;
  assign n36030 = \sport1_regs_SCTLreg_DO_reg[0]/NET0131  & ~n23265 ;
  assign n36029 = ~\sport1_txctl_Bcnt_reg[0]/NET0131  & n23265 ;
  assign n36031 = ~\sport1_rxctl_TAG_SLOT_reg/P0001  & ~n36029 ;
  assign n36032 = ~n36030 & n36031 ;
  assign n36034 = \sport0_txctl_Bcnt_reg[0]/NET0131  & \sport0_txctl_Bcnt_reg[1]/NET0131  ;
  assign n36035 = ~n19955 & ~n36034 ;
  assign n36036 = n23277 & ~n36035 ;
  assign n36033 = \sport0_regs_SCTLreg_DO_reg[1]/NET0131  & ~n23277 ;
  assign n36037 = ~\sport0_rxctl_TAG_SLOT_reg/P0001  & ~n36033 ;
  assign n36038 = ~n36036 & n36037 ;
  assign n36040 = \sport0_regs_SCTLreg_DO_reg[0]/NET0131  & ~n23277 ;
  assign n36039 = ~\sport0_txctl_Bcnt_reg[0]/NET0131  & n23277 ;
  assign n36041 = ~\sport0_rxctl_TAG_SLOT_reg/P0001  & ~n36039 ;
  assign n36042 = ~n36040 & n36041 ;
  assign n36044 = \sport0_txctl_Bcnt_reg[2]/NET0131  & ~n19955 ;
  assign n36045 = ~n19956 & ~n36044 ;
  assign n36046 = n23277 & ~n36045 ;
  assign n36043 = \sport0_regs_SCTLreg_DO_reg[2]/NET0131  & ~n23277 ;
  assign n36047 = ~\sport0_rxctl_TAG_SLOT_reg/P0001  & ~n36043 ;
  assign n36048 = ~n36046 & n36047 ;
  assign n36049 = n23715 & ~n33221 ;
  assign n36050 = ~\clkc_OUTcnt_reg[3]/NET0131  & ~n19469 ;
  assign n36051 = ~n19470 & ~n36050 ;
  assign n36052 = ~n19467 & n36051 ;
  assign n36053 = ~\clkc_STDcnt_reg[3]/NET0131  & ~n31523 ;
  assign n36054 = ~n31524 & ~n36053 ;
  assign n36055 = ~n31521 & n36054 ;
  assign n36057 = n6115 & n21249 ;
  assign n36059 = n21256 & ~n36057 ;
  assign n36058 = ~\core_c_dec_IR_reg[17]/NET0131  & n19529 ;
  assign n36060 = ~n21428 & ~n36058 ;
  assign n36061 = n36059 & n36060 ;
  assign n36062 = n14729 & n36061 ;
  assign n36056 = ~\core_c_dec_Usecond_E_reg/P0001  & n4117 ;
  assign n36063 = n4116 & ~n36056 ;
  assign n36064 = ~n36062 & n36063 ;
  assign n36065 = ~\sport0_cfg_SCLKi_cnt_reg[3]/NET0131  & ~n19534 ;
  assign n36066 = ~n19535 & ~n36065 ;
  assign n36067 = n19197 & n36066 ;
  assign n36068 = \idma_WRcyc_reg/NET0131  & ~n32460 ;
  assign n36069 = n20382 & n36068 ;
  assign n36070 = ~n20386 & n20821 ;
  assign n36071 = ~\idma_DSreq_reg/NET0131  & ~n36070 ;
  assign n36072 = ~n36069 & n36071 ;
  assign n36073 = n20070 & n22457 ;
  assign n36074 = n10638 & n36073 ;
  assign n36075 = n12688 & n18946 ;
  assign n36076 = \IRFS1_pad  & ~n36073 ;
  assign n36077 = ~n36075 & ~n36076 ;
  assign n36078 = ~n36074 & n36077 ;
  assign n36079 = n10289 & n36073 ;
  assign n36080 = \ITFS1_pad  & ~n36073 ;
  assign n36081 = ~n36075 & ~n36080 ;
  assign n36082 = ~n36079 & n36081 ;
  assign n36083 = n9435 & n36073 ;
  assign n36084 = \sport1_regs_SCTLreg_DO_reg[1]/NET0131  & ~n36073 ;
  assign n36085 = ~n36075 & ~n36084 ;
  assign n36086 = ~n36083 & n36085 ;
  assign n36087 = n8460 & n36073 ;
  assign n36088 = \sport1_regs_SCTLreg_DO_reg[11]/NET0131  & ~n36073 ;
  assign n36089 = ~n36075 & ~n36088 ;
  assign n36090 = ~n36087 & n36089 ;
  assign n36091 = n7859 & n36073 ;
  assign n36092 = \sport1_regs_SCTLreg_DO_reg[10]/NET0131  & ~n36073 ;
  assign n36093 = ~n36075 & ~n36092 ;
  assign n36094 = ~n36091 & n36093 ;
  assign n36095 = n7607 & n36073 ;
  assign n36096 = \sport1_regs_SCTLreg_DO_reg[0]/NET0131  & ~n36073 ;
  assign n36097 = ~n36075 & ~n36096 ;
  assign n36098 = ~n36095 & n36097 ;
  assign n36099 = ~\sport1_regs_MWORDreg_DO_reg[2]/NET0131  & ~n18946 ;
  assign n36100 = ~n8715 & n18948 ;
  assign n36101 = ~n36099 & ~n36100 ;
  assign n36102 = ~\sport1_regs_MWORDreg_DO_reg[3]/NET0131  & ~n18946 ;
  assign n36103 = ~n8113 & n18948 ;
  assign n36104 = ~n36102 & ~n36103 ;
  assign n36105 = ~\sport1_regs_MWORDreg_DO_reg[10]/NET0131  & ~n18946 ;
  assign n36106 = ~n12743 & n18948 ;
  assign n36107 = ~n36105 & ~n36106 ;
  assign n36108 = n18227 & n20071 ;
  assign n36109 = n11265 & n36108 ;
  assign n36110 = \sport1_regs_FSDIVreg_DO_reg[7]/NET0131  & ~n36108 ;
  assign n36111 = ~n36075 & ~n36110 ;
  assign n36112 = ~n36109 & n36111 ;
  assign n36113 = n11525 & n36108 ;
  assign n36114 = \sport1_regs_FSDIVreg_DO_reg[6]/NET0131  & ~n36108 ;
  assign n36115 = ~n36075 & ~n36114 ;
  assign n36116 = ~n36113 & n36115 ;
  assign n36117 = n10911 & n36108 ;
  assign n36118 = \sport1_regs_FSDIVreg_DO_reg[5]/NET0131  & ~n36108 ;
  assign n36119 = ~n36075 & ~n36118 ;
  assign n36120 = ~n36117 & n36119 ;
  assign n36121 = n10069 & n36108 ;
  assign n36122 = \sport1_regs_FSDIVreg_DO_reg[4]/NET0131  & ~n36108 ;
  assign n36123 = ~n36075 & ~n36122 ;
  assign n36124 = ~n36121 & n36123 ;
  assign n36125 = n8113 & n36108 ;
  assign n36126 = \sport1_regs_FSDIVreg_DO_reg[3]/NET0131  & ~n36108 ;
  assign n36127 = ~n36075 & ~n36126 ;
  assign n36128 = ~n36125 & n36127 ;
  assign n36129 = n8715 & n36108 ;
  assign n36130 = \sport1_regs_FSDIVreg_DO_reg[2]/NET0131  & ~n36108 ;
  assign n36131 = ~n36075 & ~n36130 ;
  assign n36132 = ~n36129 & n36131 ;
  assign n36133 = n9435 & n36108 ;
  assign n36134 = \sport1_regs_FSDIVreg_DO_reg[1]/NET0131  & ~n36108 ;
  assign n36135 = ~n36075 & ~n36134 ;
  assign n36136 = ~n36133 & n36135 ;
  assign n36137 = n7607 & n36108 ;
  assign n36138 = \sport1_regs_FSDIVreg_DO_reg[0]/NET0131  & ~n36108 ;
  assign n36139 = ~n36075 & ~n36138 ;
  assign n36140 = ~n36137 & n36139 ;
  assign n36141 = ~\sport1_cfg_SCLKi_cnt_reg[3]/NET0131  & ~n20232 ;
  assign n36142 = ~n20233 & ~n36141 ;
  assign n36143 = n19130 & n36142 ;
  assign n36144 = n10289 & n18229 ;
  assign n36145 = \ITFS0_pad  & ~n18229 ;
  assign n36146 = ~n18232 & ~n36145 ;
  assign n36147 = ~n36144 & n36146 ;
  assign n36148 = n10638 & n18229 ;
  assign n36149 = \IRFS0_pad  & ~n18229 ;
  assign n36150 = ~n18232 & ~n36149 ;
  assign n36151 = ~n36148 & n36150 ;
  assign n36152 = n9435 & n18229 ;
  assign n36153 = \sport0_regs_SCTLreg_DO_reg[1]/NET0131  & ~n18229 ;
  assign n36154 = ~n18232 & ~n36153 ;
  assign n36155 = ~n36152 & n36154 ;
  assign n36156 = n8460 & n18229 ;
  assign n36157 = \sport0_regs_SCTLreg_DO_reg[11]/NET0131  & ~n18229 ;
  assign n36158 = ~n18232 & ~n36157 ;
  assign n36159 = ~n36156 & n36158 ;
  assign n36160 = n7859 & n18229 ;
  assign n36161 = \sport0_regs_SCTLreg_DO_reg[10]/NET0131  & ~n18229 ;
  assign n36162 = ~n18232 & ~n36161 ;
  assign n36163 = ~n36160 & n36162 ;
  assign n36164 = n7607 & n18229 ;
  assign n36165 = \sport0_regs_SCTLreg_DO_reg[0]/NET0131  & ~n18229 ;
  assign n36166 = ~n18232 & ~n36165 ;
  assign n36167 = ~n36164 & n36166 ;
  assign n36168 = ~\sport0_regs_MWORDreg_DO_reg[3]/NET0131  & ~n18231 ;
  assign n36169 = ~n8113 & n19015 ;
  assign n36170 = ~n36168 & ~n36169 ;
  assign n36171 = ~\sport0_regs_MWORDreg_DO_reg[2]/NET0131  & ~n18231 ;
  assign n36172 = ~n8715 & n19015 ;
  assign n36173 = ~n36171 & ~n36172 ;
  assign n36174 = ~\sport0_regs_MWORDreg_DO_reg[10]/NET0131  & ~n18231 ;
  assign n36175 = ~n12743 & n19015 ;
  assign n36176 = ~n36174 & ~n36175 ;
  assign n36177 = n11265 & n18652 ;
  assign n36178 = \sport0_regs_FSDIVreg_DO_reg[7]/NET0131  & ~n18652 ;
  assign n36179 = ~n18232 & ~n36178 ;
  assign n36180 = ~n36177 & n36179 ;
  assign n36181 = n11525 & n18652 ;
  assign n36182 = \sport0_regs_FSDIVreg_DO_reg[6]/NET0131  & ~n18652 ;
  assign n36183 = ~n18232 & ~n36182 ;
  assign n36184 = ~n36181 & n36183 ;
  assign n36185 = n10911 & n18652 ;
  assign n36186 = \sport0_regs_FSDIVreg_DO_reg[5]/NET0131  & ~n18652 ;
  assign n36187 = ~n18232 & ~n36186 ;
  assign n36188 = ~n36185 & n36187 ;
  assign n36189 = n10069 & n18652 ;
  assign n36190 = \sport0_regs_FSDIVreg_DO_reg[4]/NET0131  & ~n18652 ;
  assign n36191 = ~n18232 & ~n36190 ;
  assign n36192 = ~n36189 & n36191 ;
  assign n36193 = n8113 & n18652 ;
  assign n36194 = \sport0_regs_FSDIVreg_DO_reg[3]/NET0131  & ~n18652 ;
  assign n36195 = ~n18232 & ~n36194 ;
  assign n36196 = ~n36193 & n36195 ;
  assign n36197 = n8715 & n18652 ;
  assign n36198 = \sport0_regs_FSDIVreg_DO_reg[2]/NET0131  & ~n18652 ;
  assign n36199 = ~n18232 & ~n36198 ;
  assign n36200 = ~n36197 & n36199 ;
  assign n36201 = n9435 & n18652 ;
  assign n36202 = \sport0_regs_FSDIVreg_DO_reg[1]/NET0131  & ~n18652 ;
  assign n36203 = ~n18232 & ~n36202 ;
  assign n36204 = ~n36201 & n36203 ;
  assign n36205 = n7607 & n18652 ;
  assign n36206 = \sport0_regs_FSDIVreg_DO_reg[0]/NET0131  & ~n18652 ;
  assign n36207 = ~n18232 & ~n36206 ;
  assign n36208 = ~n36205 & n36207 ;
  assign n36209 = n7232 & n7283 ;
  assign n36210 = n13762 & n36209 ;
  assign n36211 = ~n25671 & n36210 ;
  assign n36212 = \PIO_out[6]_pad  & ~n36211 ;
  assign n36213 = n11525 & n36211 ;
  assign n36214 = ~n36212 & ~n36213 ;
  assign n36215 = \PIO_oe[6]_pad  & ~n36214 ;
  assign n36216 = ~\PIO_oe[6]_pad  & \pio_PIO_RES_reg[6]/NET0131  ;
  assign n36217 = ~n36215 & ~n36216 ;
  assign n36218 = ~n25679 & n36210 ;
  assign n36219 = \PIO_out[4]_pad  & ~n36218 ;
  assign n36220 = n10069 & n36218 ;
  assign n36221 = ~n36219 & ~n36220 ;
  assign n36222 = \PIO_oe[4]_pad  & ~n36221 ;
  assign n36223 = ~\PIO_oe[4]_pad  & \pio_PIO_RES_reg[4]/NET0131  ;
  assign n36224 = ~n36222 & ~n36223 ;
  assign n36225 = ~n25666 & n36210 ;
  assign n36226 = \PIO_out[2]_pad  & ~n36225 ;
  assign n36227 = n8715 & n36225 ;
  assign n36228 = ~n36226 & ~n36227 ;
  assign n36229 = \PIO_oe[2]_pad  & ~n36228 ;
  assign n36230 = ~\PIO_oe[2]_pad  & \pio_PIO_RES_reg[2]/NET0131  ;
  assign n36231 = ~n36229 & ~n36230 ;
  assign n36232 = ~n25661 & n36210 ;
  assign n36233 = \PIO_out[10]_pad  & ~n36232 ;
  assign n36234 = n12688 & n36232 ;
  assign n36235 = ~n36233 & ~n36234 ;
  assign n36236 = \PIO_oe[10]_pad  & ~n36235 ;
  assign n36237 = ~\PIO_oe[10]_pad  & \pio_PIO_RES_reg[10]/NET0131  ;
  assign n36238 = ~n36236 & ~n36237 ;
  assign n36239 = ~n25656 & n36210 ;
  assign n36240 = \PIO_out[0]_pad  & ~n36239 ;
  assign n36241 = n7607 & n36239 ;
  assign n36242 = ~n36240 & ~n36241 ;
  assign n36243 = \PIO_oe[0]_pad  & ~n36242 ;
  assign n36244 = ~\PIO_oe[0]_pad  & \pio_PIO_RES_reg[0]/NET0131  ;
  assign n36245 = ~n36243 & ~n36244 ;
  assign n36246 = \sice_DMR1_reg[8]/NET0131  & ~n27904 ;
  assign n36247 = \sice_SPC_reg[14]/P0001  & n27904 ;
  assign n36248 = ~n36246 & ~n36247 ;
  assign n36249 = \core_c_psq_T_IRQL0p_reg/P0001  & \core_c_psq_irql0_de_OUT_reg/P0001  ;
  assign n36250 = ~\core_c_psq_T_IRQL0p_reg/P0001  & ~\core_c_psq_irql0_de_OUT_reg/P0001  ;
  assign n36251 = \core_c_psq_irql0_de_IN_syn_reg/P0001  & ~n36250 ;
  assign n36252 = ~n36249 & ~n36251 ;
  assign n36253 = ~n25651 & n36210 ;
  assign n36254 = \PIO_out[9]_pad  & ~n36253 ;
  assign n36255 = n7340 & n36253 ;
  assign n36256 = ~n36254 & ~n36255 ;
  assign n36257 = \PIO_oe[9]_pad  & ~n36256 ;
  assign n36258 = ~\PIO_oe[9]_pad  & \pio_PIO_RES_reg[9]/NET0131  ;
  assign n36259 = ~n36257 & ~n36258 ;
  assign n36260 = \PIO_out[8]_pad  & ~n36253 ;
  assign n36261 = n9178 & n36253 ;
  assign n36262 = ~n36260 & ~n36261 ;
  assign n36263 = \PIO_oe[8]_pad  & ~n36262 ;
  assign n36264 = ~\PIO_oe[8]_pad  & \pio_PIO_RES_reg[8]/NET0131  ;
  assign n36265 = ~n36263 & ~n36264 ;
  assign n36266 = \PIO_out[5]_pad  & ~n36218 ;
  assign n36267 = n10911 & n36218 ;
  assign n36268 = ~n36266 & ~n36267 ;
  assign n36269 = \PIO_oe[5]_pad  & ~n36268 ;
  assign n36270 = ~\PIO_oe[5]_pad  & \pio_PIO_RES_reg[5]/NET0131  ;
  assign n36271 = ~n36269 & ~n36270 ;
  assign n36272 = \PIO_out[7]_pad  & ~n36211 ;
  assign n36273 = n11265 & n36211 ;
  assign n36274 = ~n36272 & ~n36273 ;
  assign n36275 = \PIO_oe[7]_pad  & ~n36274 ;
  assign n36276 = ~\PIO_oe[7]_pad  & \pio_PIO_RES_reg[7]/NET0131  ;
  assign n36277 = ~n36275 & ~n36276 ;
  assign n36278 = \PIO_out[3]_pad  & ~n36225 ;
  assign n36279 = n8113 & n36225 ;
  assign n36280 = ~n36278 & ~n36279 ;
  assign n36281 = \PIO_oe[3]_pad  & ~n36280 ;
  assign n36282 = ~\PIO_oe[3]_pad  & \pio_PIO_RES_reg[3]/NET0131  ;
  assign n36283 = ~n36281 & ~n36282 ;
  assign n36284 = \PIO_out[1]_pad  & ~n36239 ;
  assign n36285 = n9435 & n36239 ;
  assign n36286 = ~n36284 & ~n36285 ;
  assign n36287 = \PIO_oe[1]_pad  & ~n36286 ;
  assign n36288 = ~\PIO_oe[1]_pad  & \pio_PIO_RES_reg[1]/NET0131  ;
  assign n36289 = ~n36287 & ~n36288 ;
  assign n36290 = \sice_SPC_reg[7]/P0001  & ~n26297 ;
  assign n36303 = \sice_DBR1_reg[2]/P0001  & n25054 ;
  assign n36304 = \sice_IMR1_reg[1]/NET0131  & n34846 ;
  assign n36311 = ~n36303 & ~n36304 ;
  assign n36305 = \sice_IIRC_reg[7]/NET0131  & n24267 ;
  assign n36306 = \sice_ICYC_reg[7]/NET0131  & n23409 ;
  assign n36312 = ~n36305 & ~n36306 ;
  assign n36313 = n36311 & n36312 ;
  assign n36299 = \sice_DMR2_reg[1]/NET0131  & n25025 ;
  assign n36300 = \sice_DBR2_reg[2]/P0001  & n25012 ;
  assign n36309 = ~n36299 & ~n36300 ;
  assign n36301 = \sice_idr0_reg_DO_reg[7]/P0001  & n26968 ;
  assign n36302 = \sice_IBR2_reg[1]/P0001  & n25074 ;
  assign n36310 = ~n36301 & ~n36302 ;
  assign n36314 = n36309 & n36310 ;
  assign n36295 = \sice_DMR1_reg[1]/NET0131  & n27903 ;
  assign n36296 = \sice_IMR2_reg[1]/NET0131  & n25034 ;
  assign n36307 = ~n36295 & ~n36296 ;
  assign n36297 = \sice_IBR1_reg[1]/P0001  & n34831 ;
  assign n36298 = \core_c_dec_IR_reg[7]/NET0131  & n28203 ;
  assign n36308 = ~n36297 & ~n36298 ;
  assign n36315 = n36307 & n36308 ;
  assign n36316 = n36314 & n36315 ;
  assign n36317 = n36313 & n36316 ;
  assign n36318 = n34827 & n36317 ;
  assign n36291 = \sice_SPC_reg[6]/P0001  & n34825 ;
  assign n36292 = \sice_SPC_reg[8]/P0001  & ~n34825 ;
  assign n36293 = ~n36291 & ~n36292 ;
  assign n36294 = ~n34827 & n36293 ;
  assign n36319 = n26297 & ~n36294 ;
  assign n36320 = ~n36318 & n36319 ;
  assign n36321 = ~n36290 & ~n36320 ;
  assign n36322 = \sice_SPC_reg[8]/P0001  & ~n26297 ;
  assign n36335 = \sice_DBR1_reg[3]/P0001  & n25054 ;
  assign n36336 = \sice_IMR1_reg[2]/NET0131  & n34846 ;
  assign n36343 = ~n36335 & ~n36336 ;
  assign n36337 = \sice_IIRC_reg[8]/NET0131  & n24267 ;
  assign n36338 = \sice_ICYC_reg[8]/NET0131  & n23409 ;
  assign n36344 = ~n36337 & ~n36338 ;
  assign n36345 = n36343 & n36344 ;
  assign n36331 = \sice_DMR2_reg[2]/NET0131  & n25025 ;
  assign n36332 = \sice_DBR2_reg[3]/P0001  & n25012 ;
  assign n36341 = ~n36331 & ~n36332 ;
  assign n36333 = \sice_idr0_reg_DO_reg[8]/P0001  & n26968 ;
  assign n36334 = \sice_IBR2_reg[2]/P0001  & n25074 ;
  assign n36342 = ~n36333 & ~n36334 ;
  assign n36346 = n36341 & n36342 ;
  assign n36327 = \sice_DMR1_reg[2]/NET0131  & n27903 ;
  assign n36328 = \sice_IMR2_reg[2]/NET0131  & n25034 ;
  assign n36339 = ~n36327 & ~n36328 ;
  assign n36329 = \sice_IBR1_reg[2]/P0001  & n34831 ;
  assign n36330 = \core_c_dec_IR_reg[8]/NET0131  & n28203 ;
  assign n36340 = ~n36329 & ~n36330 ;
  assign n36347 = n36339 & n36340 ;
  assign n36348 = n36346 & n36347 ;
  assign n36349 = n36345 & n36348 ;
  assign n36350 = n34827 & n36349 ;
  assign n36323 = \sice_SPC_reg[7]/P0001  & n34825 ;
  assign n36324 = \sice_SPC_reg[9]/P0001  & ~n34825 ;
  assign n36325 = ~n36323 & ~n36324 ;
  assign n36326 = ~n34827 & n36325 ;
  assign n36351 = n26297 & ~n36326 ;
  assign n36352 = ~n36350 & n36351 ;
  assign n36353 = ~n36322 & ~n36352 ;
  assign n36354 = \idma_WRcyc_reg/NET0131  & n32463 ;
  assign n36355 = ~n20384 & ~n36354 ;
  assign n36356 = \PIO_out[11]_pad  & ~n36232 ;
  assign n36357 = n12743 & n36232 ;
  assign n36358 = ~n36356 & ~n36357 ;
  assign n36359 = \PIO_oe[11]_pad  & ~n36358 ;
  assign n36360 = ~\PIO_oe[11]_pad  & \pio_PIO_RES_reg[11]/NET0131  ;
  assign n36361 = ~n36359 & ~n36360 ;
  assign n36363 = n20398 & n21422 ;
  assign n36362 = \core_eu_em_mac_em_dec_emcorepi_DO_reg[10]/P0001  & ~n18848 ;
  assign n36364 = \core_c_dec_IR_reg[16]/NET0131  & n18847 ;
  assign n36365 = n5123 & n36364 ;
  assign n36366 = ~n36362 & ~n36365 ;
  assign n36367 = ~n36363 & n36366 ;
  assign n36368 = ~n5951 & ~n6988 ;
  assign n36369 = ~n11738 & ~n36368 ;
  assign n36370 = n11764 & ~n36369 ;
  assign n36371 = n9513 & n12197 ;
  assign n36372 = ~n11735 & ~n36371 ;
  assign n36373 = ~n36370 & ~n36372 ;
  assign n36374 = n23032 & n34846 ;
  assign n36375 = \core_eu_em_mac_em_dec_emcorepi_DO_reg[1]/P0001  & ~n18848 ;
  assign n36376 = \core_c_dec_IR_reg[14]/NET0131  & ~\core_c_dec_IR_reg[15]/NET0131  ;
  assign n36377 = ~\core_c_dec_IR_reg[16]/NET0131  & ~n36376 ;
  assign n36378 = n18848 & n36377 ;
  assign n36379 = ~n36375 & ~n36378 ;
  assign n36380 = \core_c_psq_Iact_E_reg[2]/NET0131  & ~n19477 ;
  assign n36381 = n19477 & ~n33213 ;
  assign n36382 = n33205 & n33216 ;
  assign n36383 = n36381 & n36382 ;
  assign n36384 = ~n36380 & ~n36383 ;
  assign n36385 = \clkc_ckSTDCLK_STDCLK_reg_Q_reg/NET0131  & ~n31521 ;
  assign n36386 = ~\clkc_ckSTDCLK_STDCLK_reg_Q_reg/NET0131  & n31521 ;
  assign n36387 = ~n36385 & ~n36386 ;
  assign n36388 = n23032 & n34831 ;
  assign n36389 = \sport1_regs_MWORDreg_DO_reg[7]/NET0131  & n23274 ;
  assign n36390 = ~\sport1_txctl_Wcnt_reg[0]/NET0131  & n23726 ;
  assign n36391 = ~\sport1_txctl_Wcnt_reg[1]/NET0131  & n36390 ;
  assign n36392 = ~\sport1_txctl_Wcnt_reg[2]/NET0131  & n36391 ;
  assign n36393 = ~\sport1_txctl_Wcnt_reg[3]/NET0131  & n36392 ;
  assign n36394 = ~\sport1_txctl_Wcnt_reg[4]/NET0131  & n36393 ;
  assign n36395 = ~\sport1_txctl_Wcnt_reg[5]/NET0131  & n36394 ;
  assign n36396 = ~\sport1_txctl_Wcnt_reg[6]/NET0131  & n36395 ;
  assign n36397 = ~n23274 & ~n36396 ;
  assign n36398 = \sport1_txctl_Wcnt_reg[7]/NET0131  & n36397 ;
  assign n36399 = ~n36389 & ~n36398 ;
  assign n36400 = \sport1_txctl_Wcnt_reg[5]/NET0131  & ~n36394 ;
  assign n36401 = ~n36395 & ~n36400 ;
  assign n36402 = ~n23274 & n36401 ;
  assign n36403 = ~\sport1_regs_MWORDreg_DO_reg[5]/NET0131  & n23274 ;
  assign n36404 = ~n36402 & ~n36403 ;
  assign n36405 = \sport0_regs_MWORDreg_DO_reg[7]/NET0131  & n23286 ;
  assign n36406 = ~\sport0_txctl_Wcnt_reg[0]/NET0131  & n23744 ;
  assign n36407 = ~\sport0_txctl_Wcnt_reg[1]/NET0131  & n36406 ;
  assign n36408 = ~\sport0_txctl_Wcnt_reg[2]/NET0131  & n36407 ;
  assign n36409 = ~\sport0_txctl_Wcnt_reg[3]/NET0131  & n36408 ;
  assign n36410 = ~\sport0_txctl_Wcnt_reg[4]/NET0131  & n36409 ;
  assign n36411 = ~\sport0_txctl_Wcnt_reg[5]/NET0131  & n36410 ;
  assign n36412 = ~\sport0_txctl_Wcnt_reg[6]/NET0131  & n36411 ;
  assign n36413 = ~n23286 & ~n36412 ;
  assign n36414 = \sport0_txctl_Wcnt_reg[7]/NET0131  & n36413 ;
  assign n36415 = ~n36405 & ~n36414 ;
  assign n36416 = \sport0_txctl_Wcnt_reg[5]/NET0131  & ~n36410 ;
  assign n36417 = ~n36411 & ~n36416 ;
  assign n36418 = ~n23286 & n36417 ;
  assign n36419 = ~\sport0_regs_MWORDreg_DO_reg[5]/NET0131  & n23286 ;
  assign n36420 = ~n36418 & ~n36419 ;
  assign n36421 = ~\idma_WRcnt_reg[2]/NET0131  & ~n20459 ;
  assign n36422 = \idma_WRcnt_reg[2]/NET0131  & n20459 ;
  assign n36423 = ~n36421 & ~n36422 ;
  assign n36424 = ~n20455 & ~n36423 ;
  assign n36425 = ~\memc_usysr_DO_reg[9]/NET0131  & n20455 ;
  assign n36426 = ~n36424 & ~n36425 ;
  assign n36427 = ~n21137 & ~n21138 ;
  assign n36429 = \core_c_dec_IRE_reg[4]/NET0131  & \core_c_dec_Stkctl_Eg_reg/P0001  ;
  assign n36430 = ~\core_c_dec_MFtoppcs_Eg_reg/P0001  & ~n36429 ;
  assign n36431 = \core_c_dec_RET_Ed_reg/P0001  & ~n4184 ;
  assign n36432 = n36430 & ~n36431 ;
  assign n36433 = ~n4842 & n36432 ;
  assign n36434 = ~n5950 & ~n36433 ;
  assign n36435 = ~\core_c_psq_pcstk_ptr_reg[4]/NET0131  & n36434 ;
  assign n36436 = ~\core_c_dec_Call_Ed_reg/P0001  & ~\core_c_dec_RET_Ed_reg/P0001  ;
  assign n36437 = ~\core_c_psq_Eqend_Ed_reg/P0001  & ~\core_c_psq_TRAP_Eg_reg/NET0131  ;
  assign n36438 = n36436 & n36437 ;
  assign n36439 = n21134 & n36438 ;
  assign n36440 = n36430 & n36439 ;
  assign n36441 = n36435 & ~n36440 ;
  assign n36442 = ~n36427 & ~n36441 ;
  assign n36428 = ~n4217 & ~n36427 ;
  assign n36443 = ~n4208 & ~n21137 ;
  assign n36444 = ~n36428 & ~n36443 ;
  assign n36445 = ~n36442 & n36444 ;
  assign n36446 = \core_c_psq_pcstk_ptr_reg[3]/NET0131  & ~n36445 ;
  assign n36447 = ~\core_c_psq_pcstk_ptr_reg[3]/NET0131  & n36445 ;
  assign n36448 = ~n36446 & ~n36447 ;
  assign n36449 = ~\core_c_psq_pcstk_ptr_reg[0]/NET0131  & ~n36442 ;
  assign n36450 = \core_c_psq_pcstk_ptr_reg[1]/NET0131  & n36427 ;
  assign n36451 = ~n36449 & ~n36450 ;
  assign n36452 = ~\core_c_psq_pcstk_ptr_reg[1]/NET0131  & ~n36427 ;
  assign n36453 = ~\core_c_psq_pcstk_ptr_reg[0]/NET0131  & ~n36452 ;
  assign n36454 = ~n36451 & ~n36453 ;
  assign n36455 = \core_c_psq_pcstk_ptr_reg[2]/NET0131  & ~n36454 ;
  assign n36456 = ~\core_c_psq_pcstk_ptr_reg[2]/NET0131  & n36454 ;
  assign n36457 = ~n36455 & ~n36456 ;
  assign n36458 = ~n36450 & ~n36452 ;
  assign n36459 = n36449 & ~n36458 ;
  assign n36460 = ~n36449 & n36458 ;
  assign n36461 = ~n36459 & ~n36460 ;
  assign n36462 = \core_c_psq_pcstk_ptr_reg[0]/NET0131  & n36442 ;
  assign n36463 = ~n36449 & ~n36462 ;
  assign n36464 = \core_c_psq_Iact_E_reg[1]/NET0131  & ~n19477 ;
  assign n36465 = ~n33204 & n33210 ;
  assign n36466 = n33216 & n36465 ;
  assign n36467 = n36381 & n36466 ;
  assign n36468 = ~n36464 & ~n36467 ;
  assign n36469 = \core_c_psq_Iact_E_reg[0]/NET0131  & ~n19477 ;
  assign n36470 = ~n19488 & ~n33212 ;
  assign n36471 = ~n19480 & n36470 ;
  assign n36472 = n33218 & n36471 ;
  assign n36473 = n19494 & n36472 ;
  assign n36474 = n33211 & n36473 ;
  assign n36475 = n19487 & n36474 ;
  assign n36476 = ~n36469 & ~n36475 ;
  assign n36477 = \core_c_dec_MTIMASK_Eg_reg/P0001  & n4118 ;
  assign n36478 = ~n31998 & n35572 ;
  assign n36479 = ~n36477 & ~n36478 ;
  assign n36480 = \core_c_dec_MFTX1_E_reg/P0001  & n4117 ;
  assign n36481 = n25734 & n34556 ;
  assign n36482 = n32024 & n36481 ;
  assign n36483 = ~n36480 & ~n36482 ;
  assign n36484 = \core_c_dec_MFTX0_E_reg/P0001  & n4117 ;
  assign n36485 = n31266 & n32023 ;
  assign n36486 = n26100 & n36485 ;
  assign n36487 = ~n36484 & ~n36486 ;
  assign n36488 = \core_c_dec_MFSSTAT_E_reg/P0001  & n4117 ;
  assign n36489 = n31271 & n36481 ;
  assign n36490 = ~n36488 & ~n36489 ;
  assign n36491 = \core_c_dec_MFRX1_E_reg/P0001  & n4117 ;
  assign n36492 = ~n4117 & n34038 ;
  assign n36493 = n31264 & n36492 ;
  assign n36494 = ~n36491 & ~n36493 ;
  assign n36495 = \core_c_dec_MFRX0_E_reg/P0001  & n4117 ;
  assign n36496 = n25729 & n36485 ;
  assign n36497 = ~n36495 & ~n36496 ;
  assign n36498 = ~n4117 & ~n33278 ;
  assign n36499 = ~\core_c_dec_MFPMOVL_E_reg/P0001  & n4117 ;
  assign n36500 = ~n36498 & ~n36499 ;
  assign n36501 = \core_c_dec_MFMreg_E_reg[7]/P0001  & n4117 ;
  assign n36502 = n26100 & n34042 ;
  assign n36503 = ~n36501 & ~n36502 ;
  assign n36504 = \core_c_dec_MFMreg_E_reg[6]/P0001  & n4117 ;
  assign n36505 = n25729 & n34042 ;
  assign n36506 = ~n36504 & ~n36505 ;
  assign n36507 = n26100 & n31978 ;
  assign n36508 = n34030 & n36507 ;
  assign n36509 = \core_c_dec_MFMreg_E_reg[5]/P0001  & n4117 ;
  assign n36510 = ~n36508 & ~n36509 ;
  assign n36511 = \core_c_dec_MFMreg_E_reg[4]/P0001  & n4117 ;
  assign n36512 = n34030 & n35757 ;
  assign n36513 = ~n36511 & ~n36512 ;
  assign n36514 = \core_c_dec_MFMreg_E_reg[3]/P0001  & n4117 ;
  assign n36515 = n6091 & ~n31263 ;
  assign n36516 = n19301 & n31966 ;
  assign n36517 = ~n4117 & n36516 ;
  assign n36518 = n36515 & n36517 ;
  assign n36519 = ~n36514 & ~n36518 ;
  assign n36520 = \core_c_dec_MFMreg_E_reg[2]/P0001  & n4117 ;
  assign n36521 = n19298 & n31966 ;
  assign n36522 = ~n4117 & n36521 ;
  assign n36523 = n36515 & n36522 ;
  assign n36524 = ~n36520 & ~n36523 ;
  assign n36525 = \core_c_dec_MFMreg_E_reg[1]/P0001  & n4117 ;
  assign n36526 = n19267 & n31966 ;
  assign n36527 = ~n4117 & n36526 ;
  assign n36528 = n36515 & n36527 ;
  assign n36529 = ~n36525 & ~n36528 ;
  assign n36530 = \core_c_dec_MFMreg_E_reg[0]/P0001  & n4117 ;
  assign n36531 = n19270 & n31973 ;
  assign n36532 = n25852 & n36531 ;
  assign n36533 = ~n36530 & ~n36532 ;
  assign n36534 = \core_c_dec_MFMSTAT_E_reg/P0001  & n4117 ;
  assign n36535 = n31266 & n36507 ;
  assign n36536 = ~n36534 & ~n36535 ;
  assign n36537 = ~\core_c_dec_MFLreg_E_reg[7]/P0001  & n4117 ;
  assign n36538 = ~n34034 & ~n36537 ;
  assign n36539 = \core_c_dec_MFLreg_E_reg[6]/P0001  & n4117 ;
  assign n36540 = n34024 & n36492 ;
  assign n36541 = ~n36539 & ~n36540 ;
  assign n36542 = ~n4117 & ~n34035 ;
  assign n36543 = ~\core_c_dec_MFLreg_E_reg[5]/P0001  & n4117 ;
  assign n36544 = ~n36542 & ~n36543 ;
  assign n36545 = \core_c_dec_MFLreg_E_reg[4]/P0001  & n4117 ;
  assign n36546 = n25864 & n34026 ;
  assign n36547 = ~n36545 & ~n36546 ;
  assign n36548 = ~n4117 & n31982 ;
  assign n36549 = \core_c_dec_MFLreg_E_reg[3]/P0001  & n4117 ;
  assign n36550 = ~n36548 & ~n36549 ;
  assign n36551 = ~n4117 & n31975 ;
  assign n36552 = \core_c_dec_MFLreg_E_reg[2]/P0001  & n4117 ;
  assign n36553 = ~n36551 & ~n36552 ;
  assign n36554 = ~\core_c_dec_MFLreg_E_reg[0]/P0001  & n4117 ;
  assign n36555 = ~n31971 & ~n36554 ;
  assign n36556 = \core_c_dec_MFIreg_E_reg[7]/P0001  & n4117 ;
  assign n36557 = n34028 & n36507 ;
  assign n36558 = ~n36556 & ~n36557 ;
  assign n36559 = \core_c_dec_MFIreg_E_reg[6]/P0001  & n4117 ;
  assign n36560 = n34028 & n35757 ;
  assign n36561 = ~n36559 & ~n36560 ;
  assign n36562 = \core_c_dec_MFIreg_E_reg[5]/P0001  & n4117 ;
  assign n36563 = n34025 & n36507 ;
  assign n36564 = ~n36562 & ~n36563 ;
  assign n36565 = \core_c_dec_MFIreg_E_reg[4]/P0001  & n4117 ;
  assign n36566 = n34025 & n35757 ;
  assign n36567 = ~n36565 & ~n36566 ;
  assign n36568 = \core_c_dec_MFIreg_E_reg[3]/P0001  & n4117 ;
  assign n36569 = n6093 & ~n31263 ;
  assign n36570 = n36517 & n36569 ;
  assign n36571 = ~n36568 & ~n36570 ;
  assign n36572 = \core_c_dec_MFIreg_E_reg[1]/P0001  & n4117 ;
  assign n36573 = n36527 & n36569 ;
  assign n36574 = ~n36572 & ~n36573 ;
  assign n36575 = \core_c_dec_MFIreg_E_reg[0]/P0001  & n4117 ;
  assign n36576 = n31265 & n31973 ;
  assign n36577 = n25729 & n36576 ;
  assign n36578 = ~n36575 & ~n36577 ;
  assign n36579 = \core_c_dec_MFIMASK_E_reg/P0001  & n4117 ;
  assign n36580 = n31979 & n36481 ;
  assign n36581 = ~n36579 & ~n36580 ;
  assign n36582 = ~n4117 & n33279 ;
  assign n36583 = \core_c_dec_MFIDR_E_reg/P0001  & n4117 ;
  assign n36584 = ~n36582 & ~n36583 ;
  assign n36585 = ~\core_c_dec_MFDMOVL_E_reg/P0001  & n4117 ;
  assign n36586 = ~n33277 & ~n36585 ;
  assign n36587 = \core_c_dec_MFASTAT_E_reg/P0001  & n4117 ;
  assign n36588 = n31266 & n35757 ;
  assign n36589 = ~n36587 & ~n36588 ;
  assign n36590 = ~\bdma_BEAD_reg[4]/NET0131  & ~n33305 ;
  assign n36591 = ~n20765 & ~n33306 ;
  assign n36592 = ~n36590 & n36591 ;
  assign n36593 = n10069 & n20765 ;
  assign n36594 = ~n36592 & ~n36593 ;
  assign n36595 = ~\bdma_BEAD_reg[3]/NET0131  & ~n33304 ;
  assign n36596 = ~n20765 & ~n33305 ;
  assign n36597 = ~n36595 & n36596 ;
  assign n36598 = n8113 & n20765 ;
  assign n36599 = ~n36597 & ~n36598 ;
  assign n36600 = \core_c_dec_MFIreg_E_reg[2]/P0001  & n4117 ;
  assign n36601 = n36522 & n36569 ;
  assign n36602 = ~n36600 & ~n36601 ;
  assign n36603 = n4215 & n36427 ;
  assign n36604 = n4218 & ~n36427 ;
  assign n36605 = n36441 & n36604 ;
  assign n36606 = ~\core_c_psq_pcstk_ptr_reg[4]/NET0131  & ~n36605 ;
  assign n36607 = ~n36603 & ~n36606 ;
  assign n36608 = ~\sice_ICYC_reg[19]/NET0131  & ~n20748 ;
  assign n36609 = ~n20749 & ~n36608 ;
  assign n36610 = \core_c_dec_MFtoppcs_Eg_reg/P0001  & n4118 ;
  assign n36611 = n23231 & n32025 ;
  assign n36612 = ~n36610 & ~n36611 ;
  assign n36613 = \sice_SPC_reg[22]/P0001  & n34825 ;
  assign n36614 = T_ID_pad & ~n34825 ;
  assign n36615 = ~n36613 & ~n36614 ;
  assign n36616 = ~n34827 & n36615 ;
  assign n36624 = \emc_eRDY_reg/NET0131  & n35008 ;
  assign n36617 = \sice_IMR1_reg[17]/NET0131  & n34846 ;
  assign n36632 = ~n25084 & ~n36617 ;
  assign n36618 = \sice_CMRW_reg/NET0131  & n23029 ;
  assign n36619 = \sice_DMR1_reg[17]/NET0131  & n27903 ;
  assign n36633 = ~n36618 & ~n36619 ;
  assign n36642 = n36632 & n36633 ;
  assign n36643 = ~n36624 & n36642 ;
  assign n36631 = \sice_DMR2_reg[17]/NET0131  & n25025 ;
  assign n36629 = \sice_ICYC_reg[23]/NET0131  & n23409 ;
  assign n36630 = \sice_IBR1_reg[17]/P0001  & n34831 ;
  assign n36638 = ~n36629 & ~n36630 ;
  assign n36639 = ~n36631 & n36638 ;
  assign n36625 = \core_c_dec_IR_reg[23]/NET0131  & n28203 ;
  assign n36626 = \sice_IRR_reg[13]/P0001  & n34841 ;
  assign n36636 = ~n36625 & ~n36626 ;
  assign n36627 = \sice_IIRC_reg[23]/NET0131  & n24267 ;
  assign n36628 = \sice_IMR2_reg[17]/NET0131  & n25034 ;
  assign n36637 = ~n36627 & ~n36628 ;
  assign n36640 = n36636 & n36637 ;
  assign n36620 = \sice_DBR1_reg[18]/P0001  & n25054 ;
  assign n36621 = \sice_DBR2_reg[18]/P0001  & n25012 ;
  assign n36634 = ~n36620 & ~n36621 ;
  assign n36622 = \sice_IBR2_reg[17]/P0001  & n25074 ;
  assign n36623 = \sice_idr1_reg_DO_reg[11]/P0001  & n26968 ;
  assign n36635 = ~n36622 & ~n36623 ;
  assign n36641 = n36634 & n36635 ;
  assign n36644 = n36640 & n36641 ;
  assign n36645 = n36639 & n36644 ;
  assign n36646 = n36643 & n36645 ;
  assign n36647 = n34827 & n36646 ;
  assign n36648 = ~n36616 & ~n36647 ;
  assign n36649 = \sice_SPC_reg[21]/P0001  & n34825 ;
  assign n36650 = \sice_SPC_reg[23]/P0001  & ~n34825 ;
  assign n36651 = ~n36649 & ~n36650 ;
  assign n36652 = ~n34827 & n36651 ;
  assign n36660 = \sice_IDONE_reg/NET0131  & n35008 ;
  assign n36653 = \sice_IMR1_reg[16]/NET0131  & n34846 ;
  assign n36668 = ~n25084 & ~n36653 ;
  assign n36654 = \sice_IIRC_reg[22]/NET0131  & n24267 ;
  assign n36655 = \sice_DMR1_reg[16]/NET0131  & n27903 ;
  assign n36669 = ~n36654 & ~n36655 ;
  assign n36678 = n36668 & n36669 ;
  assign n36679 = ~n36660 & n36678 ;
  assign n36667 = \sice_DMR2_reg[16]/NET0131  & n25025 ;
  assign n36665 = \sice_IBR2_reg[16]/P0001  & n25074 ;
  assign n36666 = \sice_IBR1_reg[16]/P0001  & n34831 ;
  assign n36674 = ~n36665 & ~n36666 ;
  assign n36675 = ~n36667 & n36674 ;
  assign n36661 = \core_c_dec_IR_reg[22]/NET0131  & n28203 ;
  assign n36662 = \sice_IRR_reg[12]/P0001  & n34841 ;
  assign n36672 = ~n36661 & ~n36662 ;
  assign n36663 = \sice_ICYC_reg[22]/NET0131  & n23409 ;
  assign n36664 = \sice_IMR2_reg[16]/NET0131  & n25034 ;
  assign n36673 = ~n36663 & ~n36664 ;
  assign n36676 = n36672 & n36673 ;
  assign n36656 = \sice_DBR1_reg[17]/P0001  & n25054 ;
  assign n36657 = \sice_DBR2_reg[17]/P0001  & n25012 ;
  assign n36670 = ~n36656 & ~n36657 ;
  assign n36658 = \sice_CLR_M_reg/NET0131  & n23029 ;
  assign n36659 = \sice_idr1_reg_DO_reg[10]/P0001  & n26968 ;
  assign n36671 = ~n36658 & ~n36659 ;
  assign n36677 = n36670 & n36671 ;
  assign n36680 = n36676 & n36677 ;
  assign n36681 = n36675 & n36680 ;
  assign n36682 = n36679 & n36681 ;
  assign n36683 = n34827 & n36682 ;
  assign n36684 = ~n36652 & ~n36683 ;
  assign n36685 = \sice_SPC_reg[19]/P0001  & n34825 ;
  assign n36686 = \sice_SPC_reg[21]/P0001  & ~n34825 ;
  assign n36687 = ~n36685 & ~n36686 ;
  assign n36688 = ~n34827 & n36687 ;
  assign n36696 = ~n4068 & n35008 ;
  assign n36689 = \sice_IMR1_reg[14]/NET0131  & n34846 ;
  assign n36704 = ~n25084 & ~n36689 ;
  assign n36690 = \sice_IIRC_reg[20]/NET0131  & n24267 ;
  assign n36691 = \sice_DMR1_reg[14]/NET0131  & n27903 ;
  assign n36705 = ~n36690 & ~n36691 ;
  assign n36714 = n36704 & n36705 ;
  assign n36715 = ~n36696 & n36714 ;
  assign n36703 = \sice_DMR2_reg[14]/NET0131  & n25025 ;
  assign n36701 = \sice_IBR2_reg[14]/P0001  & n25074 ;
  assign n36702 = \sice_IBR1_reg[14]/P0001  & n34831 ;
  assign n36710 = ~n36701 & ~n36702 ;
  assign n36711 = ~n36703 & n36710 ;
  assign n36697 = \core_c_dec_IR_reg[20]/NET0131  & n28203 ;
  assign n36698 = \sice_IRR_reg[10]/P0001  & n34841 ;
  assign n36708 = ~n36697 & ~n36698 ;
  assign n36699 = \sice_ICYC_reg[20]/NET0131  & n23409 ;
  assign n36700 = \sice_IMR2_reg[14]/NET0131  & n25034 ;
  assign n36709 = ~n36699 & ~n36700 ;
  assign n36712 = n36708 & n36709 ;
  assign n36692 = \sice_DBR1_reg[15]/P0001  & n25054 ;
  assign n36693 = \sice_DBR2_reg[15]/P0001  & n25012 ;
  assign n36706 = ~n36692 & ~n36693 ;
  assign n36694 = \sice_GO_NX_reg/NET0131  & n23029 ;
  assign n36695 = \sice_idr1_reg_DO_reg[8]/P0001  & n26968 ;
  assign n36707 = ~n36694 & ~n36695 ;
  assign n36713 = n36706 & n36707 ;
  assign n36716 = n36712 & n36713 ;
  assign n36717 = n36711 & n36716 ;
  assign n36718 = n36715 & n36717 ;
  assign n36719 = n34827 & n36718 ;
  assign n36720 = ~n36688 & ~n36719 ;
  assign n36721 = \sice_SPC_reg[18]/P0001  & n34825 ;
  assign n36722 = \sice_SPC_reg[20]/P0001  & ~n34825 ;
  assign n36723 = ~n36721 & ~n36722 ;
  assign n36724 = ~n34827 & n36723 ;
  assign n36732 = \core_c_psq_MGNT_reg/NET0131  & n35008 ;
  assign n36725 = \sice_IMR1_reg[13]/NET0131  & n34846 ;
  assign n36740 = ~n25084 & ~n36725 ;
  assign n36726 = \sice_IIRC_reg[19]/NET0131  & n24267 ;
  assign n36727 = \sice_DMR1_reg[13]/NET0131  & n27903 ;
  assign n36741 = ~n36726 & ~n36727 ;
  assign n36750 = n36740 & n36741 ;
  assign n36751 = ~n36732 & n36750 ;
  assign n36739 = \sice_DMR2_reg[13]/NET0131  & n25025 ;
  assign n36737 = \sice_IBR2_reg[13]/P0001  & n25074 ;
  assign n36738 = \sice_IBR1_reg[13]/P0001  & n34831 ;
  assign n36746 = ~n36737 & ~n36738 ;
  assign n36747 = ~n36739 & n36746 ;
  assign n36733 = \core_c_dec_IR_reg[19]/NET0131  & n28203 ;
  assign n36734 = \sice_IRR_reg[9]/P0001  & n34841 ;
  assign n36744 = ~n36733 & ~n36734 ;
  assign n36735 = \sice_ICYC_reg[19]/NET0131  & n23409 ;
  assign n36736 = \sice_IMR2_reg[13]/NET0131  & n25034 ;
  assign n36745 = ~n36735 & ~n36736 ;
  assign n36748 = n36744 & n36745 ;
  assign n36728 = \sice_DBR1_reg[14]/P0001  & n25054 ;
  assign n36729 = \sice_DBR2_reg[14]/P0001  & n25012 ;
  assign n36742 = ~n36728 & ~n36729 ;
  assign n36730 = ~n23018 & n23029 ;
  assign n36731 = \sice_idr1_reg_DO_reg[7]/P0001  & n26968 ;
  assign n36743 = ~n36730 & ~n36731 ;
  assign n36749 = n36742 & n36743 ;
  assign n36752 = n36748 & n36749 ;
  assign n36753 = n36747 & n36752 ;
  assign n36754 = n36751 & n36753 ;
  assign n36755 = n34827 & n36754 ;
  assign n36756 = ~n36724 & ~n36755 ;
  assign n36757 = \sice_SPC_reg[17]/P0001  & n34825 ;
  assign n36758 = \sice_SPC_reg[19]/P0001  & ~n34825 ;
  assign n36759 = ~n36757 & ~n36758 ;
  assign n36760 = ~n34827 & n36759 ;
  assign n36768 = \core_c_psq_PCS_reg[3]/NET0131  & n35008 ;
  assign n36761 = \sice_IMR1_reg[12]/NET0131  & n34846 ;
  assign n36776 = ~n25084 & ~n36761 ;
  assign n36762 = \sice_IIRC_reg[18]/NET0131  & n24267 ;
  assign n36763 = \sice_DMR1_reg[12]/NET0131  & n27903 ;
  assign n36777 = ~n36762 & ~n36763 ;
  assign n36786 = n36776 & n36777 ;
  assign n36787 = ~n36768 & n36786 ;
  assign n36775 = \sice_DMR2_reg[12]/NET0131  & n25025 ;
  assign n36773 = \sice_IBR2_reg[12]/P0001  & n25074 ;
  assign n36774 = \sice_IBR1_reg[12]/P0001  & n34831 ;
  assign n36782 = ~n36773 & ~n36774 ;
  assign n36783 = ~n36775 & n36782 ;
  assign n36769 = \core_c_dec_IR_reg[18]/NET0131  & n28203 ;
  assign n36770 = \sice_IRR_reg[8]/P0001  & n34841 ;
  assign n36780 = ~n36769 & ~n36770 ;
  assign n36771 = \sice_ICYC_reg[18]/NET0131  & n23409 ;
  assign n36772 = \sice_IMR2_reg[12]/NET0131  & n25034 ;
  assign n36781 = ~n36771 & ~n36772 ;
  assign n36784 = n36780 & n36781 ;
  assign n36764 = \sice_DBR1_reg[13]/P0001  & n25054 ;
  assign n36765 = \sice_DBR2_reg[13]/P0001  & n25012 ;
  assign n36778 = ~n36764 & ~n36765 ;
  assign n36766 = \sice_IRST_reg/NET0131  & n23029 ;
  assign n36767 = \sice_idr1_reg_DO_reg[6]/P0001  & n26968 ;
  assign n36779 = ~n36766 & ~n36767 ;
  assign n36785 = n36778 & n36779 ;
  assign n36788 = n36784 & n36785 ;
  assign n36789 = n36783 & n36788 ;
  assign n36790 = n36787 & n36789 ;
  assign n36791 = n34827 & n36790 ;
  assign n36792 = ~n36760 & ~n36791 ;
  assign n36793 = \core_c_dec_MFSB_E_reg/P0001  & n4117 ;
  assign n36794 = n31654 & n35757 ;
  assign n36795 = ~n36793 & ~n36794 ;
  assign n36796 = ~n4117 & n31977 ;
  assign n36797 = \core_c_dec_MFLreg_E_reg[1]/P0001  & n4117 ;
  assign n36798 = ~n36796 & ~n36797 ;
  assign n36799 = \core_c_dec_MFCNTR_E_reg/P0001  & n4117 ;
  assign n36800 = n35756 & n36507 ;
  assign n36801 = ~n36799 & ~n36800 ;
  assign n36802 = \sice_SPC_reg[12]/P0001  & n34825 ;
  assign n36803 = \sice_SPC_reg[14]/P0001  & ~n34825 ;
  assign n36804 = ~n36802 & ~n36803 ;
  assign n36805 = ~n34827 & n36804 ;
  assign n36806 = \sice_IMR2_reg[7]/NET0131  & n25034 ;
  assign n36819 = ~n25083 & ~n36806 ;
  assign n36807 = \sice_IRR_reg[3]/P0001  & n34841 ;
  assign n36808 = \sice_IBR1_reg[7]/P0001  & n34831 ;
  assign n36820 = ~n36807 & ~n36808 ;
  assign n36809 = \sice_IBR2_reg[7]/P0001  & n25074 ;
  assign n36810 = \core_c_dec_IR_reg[13]/NET0131  & n28203 ;
  assign n36821 = ~n36809 & ~n36810 ;
  assign n36828 = n36820 & n36821 ;
  assign n36829 = n36819 & n36828 ;
  assign n36815 = \sice_DBR2_reg[8]/P0001  & n25012 ;
  assign n36816 = \sice_DBR1_reg[8]/P0001  & n25054 ;
  assign n36824 = ~n36815 & ~n36816 ;
  assign n36817 = \sice_IIRC_reg[13]/NET0131  & n24267 ;
  assign n36818 = \sice_idr1_reg_DO_reg[1]/P0001  & n26968 ;
  assign n36825 = ~n36817 & ~n36818 ;
  assign n36826 = n36824 & n36825 ;
  assign n36811 = \sice_DMR2_reg[7]/NET0131  & n25025 ;
  assign n36812 = \sice_ICYC_reg[13]/NET0131  & n23409 ;
  assign n36822 = ~n36811 & ~n36812 ;
  assign n36813 = \sice_IMR1_reg[7]/NET0131  & n34846 ;
  assign n36814 = \sice_DMR1_reg[7]/NET0131  & n27903 ;
  assign n36823 = ~n36813 & ~n36814 ;
  assign n36827 = n36822 & n36823 ;
  assign n36830 = n36826 & n36827 ;
  assign n36831 = n36829 & n36830 ;
  assign n36832 = n34827 & n36831 ;
  assign n36833 = ~n36805 & ~n36832 ;
  assign n36834 = \sice_SPC_reg[13]/P0001  & n34825 ;
  assign n36835 = \sice_SPC_reg[15]/P0001  & ~n34825 ;
  assign n36836 = ~n36834 & ~n36835 ;
  assign n36837 = ~n34827 & n36836 ;
  assign n36838 = \sice_DBR1_reg[9]/P0001  & n25054 ;
  assign n36851 = ~n25083 & ~n36838 ;
  assign n36839 = \sice_IRR_reg[4]/P0001  & n34841 ;
  assign n36840 = \sice_IMR2_reg[8]/NET0131  & n25034 ;
  assign n36852 = ~n36839 & ~n36840 ;
  assign n36841 = \sice_IBR2_reg[8]/P0001  & n25074 ;
  assign n36842 = \core_c_dec_IR_reg[14]/NET0131  & n28203 ;
  assign n36853 = ~n36841 & ~n36842 ;
  assign n36860 = n36852 & n36853 ;
  assign n36861 = n36851 & n36860 ;
  assign n36847 = \sice_IIRC_reg[14]/NET0131  & n24267 ;
  assign n36848 = \sice_DBR2_reg[9]/P0001  & n25012 ;
  assign n36856 = ~n36847 & ~n36848 ;
  assign n36849 = \sice_DMR1_reg[8]/NET0131  & n27903 ;
  assign n36850 = \sice_idr1_reg_DO_reg[2]/P0001  & n26968 ;
  assign n36857 = ~n36849 & ~n36850 ;
  assign n36858 = n36856 & n36857 ;
  assign n36843 = \sice_DMR2_reg[8]/NET0131  & n25025 ;
  assign n36844 = \sice_ICYC_reg[14]/NET0131  & n23409 ;
  assign n36854 = ~n36843 & ~n36844 ;
  assign n36845 = \sice_IMR1_reg[8]/NET0131  & n34846 ;
  assign n36846 = \sice_IBR1_reg[8]/P0001  & n34831 ;
  assign n36855 = ~n36845 & ~n36846 ;
  assign n36859 = n36854 & n36855 ;
  assign n36862 = n36858 & n36859 ;
  assign n36863 = n36861 & n36862 ;
  assign n36864 = n34827 & n36863 ;
  assign n36865 = ~n36837 & ~n36864 ;
  assign n36866 = \sice_SPC_reg[14]/P0001  & n34825 ;
  assign n36867 = \sice_SPC_reg[16]/P0001  & ~n34825 ;
  assign n36868 = ~n36866 & ~n36867 ;
  assign n36869 = ~n34827 & n36868 ;
  assign n36870 = \sice_DBR1_reg[10]/P0001  & n25054 ;
  assign n36883 = ~n25083 & ~n36870 ;
  assign n36871 = \sice_IRR_reg[5]/P0001  & n34841 ;
  assign n36872 = \sice_IMR2_reg[9]/NET0131  & n25034 ;
  assign n36884 = ~n36871 & ~n36872 ;
  assign n36873 = \sice_IBR2_reg[9]/P0001  & n25074 ;
  assign n36874 = \core_c_dec_IR_reg[15]/NET0131  & n28203 ;
  assign n36885 = ~n36873 & ~n36874 ;
  assign n36892 = n36884 & n36885 ;
  assign n36893 = n36883 & n36892 ;
  assign n36879 = \sice_IIRC_reg[15]/NET0131  & n24267 ;
  assign n36880 = \sice_DBR2_reg[10]/P0001  & n25012 ;
  assign n36888 = ~n36879 & ~n36880 ;
  assign n36881 = \sice_DMR1_reg[9]/NET0131  & n27903 ;
  assign n36882 = \sice_idr1_reg_DO_reg[3]/P0001  & n26968 ;
  assign n36889 = ~n36881 & ~n36882 ;
  assign n36890 = n36888 & n36889 ;
  assign n36875 = \sice_DMR2_reg[9]/NET0131  & n25025 ;
  assign n36876 = \sice_ICYC_reg[15]/NET0131  & n23409 ;
  assign n36886 = ~n36875 & ~n36876 ;
  assign n36877 = \sice_IMR1_reg[9]/NET0131  & n34846 ;
  assign n36878 = \sice_IBR1_reg[9]/P0001  & n34831 ;
  assign n36887 = ~n36877 & ~n36878 ;
  assign n36891 = n36886 & n36887 ;
  assign n36894 = n36890 & n36891 ;
  assign n36895 = n36893 & n36894 ;
  assign n36896 = n34827 & n36895 ;
  assign n36897 = ~n36869 & ~n36896 ;
  assign n36898 = ~\sice_ICYC_reg[11]/NET0131  & ~n20740 ;
  assign n36899 = ~n20741 & ~n36898 ;
  assign n36900 = ~\sice_IIRC_reg[11]/NET0131  & ~n20855 ;
  assign n36901 = ~n20856 & ~n36900 ;
  assign n36902 = \sice_SPC_reg[16]/P0001  & n34825 ;
  assign n36903 = \sice_SPC_reg[18]/P0001  & ~n34825 ;
  assign n36904 = ~n36902 & ~n36903 ;
  assign n36905 = ~n34827 & n36904 ;
  assign n36906 = \sice_DBR1_reg[12]/P0001  & n25054 ;
  assign n36919 = ~n25083 & ~n36906 ;
  assign n36907 = \sice_IRR_reg[7]/P0001  & n34841 ;
  assign n36908 = \sice_IMR2_reg[11]/NET0131  & n25034 ;
  assign n36920 = ~n36907 & ~n36908 ;
  assign n36909 = \sice_IBR2_reg[11]/P0001  & n25074 ;
  assign n36910 = \sice_idr1_reg_DO_reg[5]/P0001  & n26968 ;
  assign n36921 = ~n36909 & ~n36910 ;
  assign n36928 = n36920 & n36921 ;
  assign n36929 = n36919 & n36928 ;
  assign n36915 = \sice_IIRC_reg[17]/NET0131  & n24267 ;
  assign n36916 = \sice_DBR2_reg[12]/P0001  & n25012 ;
  assign n36924 = ~n36915 & ~n36916 ;
  assign n36917 = \sice_DMR1_reg[11]/NET0131  & n27903 ;
  assign n36918 = \core_c_dec_IR_reg[17]/NET0131  & n28203 ;
  assign n36925 = ~n36917 & ~n36918 ;
  assign n36926 = n36924 & n36925 ;
  assign n36911 = \sice_DMR2_reg[11]/NET0131  & n25025 ;
  assign n36912 = \sice_ICYC_reg[17]/NET0131  & n23409 ;
  assign n36922 = ~n36911 & ~n36912 ;
  assign n36913 = \sice_IMR1_reg[11]/NET0131  & n34846 ;
  assign n36914 = \sice_IBR1_reg[11]/P0001  & n34831 ;
  assign n36923 = ~n36913 & ~n36914 ;
  assign n36927 = n36922 & n36923 ;
  assign n36930 = n36926 & n36927 ;
  assign n36931 = n36929 & n36930 ;
  assign n36932 = n34827 & n36931 ;
  assign n36933 = ~n36905 & ~n36932 ;
  assign n36934 = ~\memc_Dread_E_reg/NET0131  & ~\memc_Dwrite_E_reg/NET0131  ;
  assign n36935 = n5435 & ~n36934 ;
  assign n36936 = ~n4068 & n36935 ;
  assign n36937 = ~n19054 & n36936 ;
  assign n36938 = \emc_DMcst_reg/NET0131  & ~n23398 ;
  assign n36939 = n19054 & n36938 ;
  assign n36940 = ~n36937 & ~n36939 ;
  assign n36941 = \sice_SPC_reg[15]/P0001  & n34825 ;
  assign n36942 = \sice_SPC_reg[17]/P0001  & ~n34825 ;
  assign n36943 = ~n36941 & ~n36942 ;
  assign n36944 = ~n34827 & n36943 ;
  assign n36945 = \sice_DBR1_reg[11]/P0001  & n25054 ;
  assign n36958 = ~n25083 & ~n36945 ;
  assign n36946 = \sice_IRR_reg[6]/P0001  & n34841 ;
  assign n36947 = \sice_IMR2_reg[10]/NET0131  & n25034 ;
  assign n36959 = ~n36946 & ~n36947 ;
  assign n36948 = \sice_IBR2_reg[10]/P0001  & n25074 ;
  assign n36949 = \sice_idr1_reg_DO_reg[4]/P0001  & n26968 ;
  assign n36960 = ~n36948 & ~n36949 ;
  assign n36967 = n36959 & n36960 ;
  assign n36968 = n36958 & n36967 ;
  assign n36954 = \sice_IIRC_reg[16]/NET0131  & n24267 ;
  assign n36955 = \sice_DBR2_reg[11]/P0001  & n25012 ;
  assign n36963 = ~n36954 & ~n36955 ;
  assign n36956 = \sice_DMR1_reg[10]/NET0131  & n27903 ;
  assign n36957 = \core_c_dec_IR_reg[16]/NET0131  & n28203 ;
  assign n36964 = ~n36956 & ~n36957 ;
  assign n36965 = n36963 & n36964 ;
  assign n36950 = \sice_DMR2_reg[10]/NET0131  & n25025 ;
  assign n36951 = \sice_ICYC_reg[16]/NET0131  & n23409 ;
  assign n36961 = ~n36950 & ~n36951 ;
  assign n36952 = \sice_IMR1_reg[10]/NET0131  & n34846 ;
  assign n36953 = \sice_IBR1_reg[10]/P0001  & n34831 ;
  assign n36962 = ~n36952 & ~n36953 ;
  assign n36966 = n36961 & n36962 ;
  assign n36969 = n36965 & n36966 ;
  assign n36970 = n36968 & n36969 ;
  assign n36971 = n34827 & n36970 ;
  assign n36972 = ~n36944 & ~n36971 ;
  assign n36973 = \sice_SPC_reg[4]/P0001  & ~n26297 ;
  assign n36978 = \sice_idr0_reg_DO_reg[4]/P0001  & n26968 ;
  assign n36979 = \core_c_dec_IR_reg[4]/NET0131  & n28203 ;
  assign n36982 = ~n36978 & ~n36979 ;
  assign n36980 = \sice_ICYC_reg[4]/NET0131  & n23409 ;
  assign n36981 = \sice_IIRC_reg[4]/NET0131  & n24267 ;
  assign n36983 = ~n36980 & ~n36981 ;
  assign n36984 = n36982 & n36983 ;
  assign n36985 = n34827 & n36984 ;
  assign n36974 = \sice_SPC_reg[3]/P0001  & n34825 ;
  assign n36975 = \sice_SPC_reg[5]/P0001  & ~n34825 ;
  assign n36976 = ~n36974 & ~n36975 ;
  assign n36977 = ~n34827 & n36976 ;
  assign n36986 = n26297 & ~n36977 ;
  assign n36987 = ~n36985 & n36986 ;
  assign n36988 = ~n36973 & ~n36987 ;
  assign n36989 = \sice_SPC_reg[3]/P0001  & ~n26297 ;
  assign n36994 = \sice_idr0_reg_DO_reg[3]/P0001  & n26968 ;
  assign n36995 = \core_c_dec_IR_reg[3]/NET0131  & n28203 ;
  assign n36998 = ~n36994 & ~n36995 ;
  assign n36996 = \sice_ICYC_reg[3]/NET0131  & n23409 ;
  assign n36997 = \sice_IIRC_reg[3]/NET0131  & n24267 ;
  assign n36999 = ~n36996 & ~n36997 ;
  assign n37000 = n36998 & n36999 ;
  assign n37001 = n34827 & n37000 ;
  assign n36990 = \sice_SPC_reg[2]/P0001  & n34825 ;
  assign n36991 = \sice_SPC_reg[4]/P0001  & ~n34825 ;
  assign n36992 = ~n36990 & ~n36991 ;
  assign n36993 = ~n34827 & n36992 ;
  assign n37002 = n26297 & ~n36993 ;
  assign n37003 = ~n37001 & n37002 ;
  assign n37004 = ~n36989 & ~n37003 ;
  assign n37005 = \sice_SPC_reg[2]/P0001  & ~n26297 ;
  assign n37010 = \sice_idr0_reg_DO_reg[2]/P0001  & n26968 ;
  assign n37011 = \core_c_dec_IR_reg[2]/NET0131  & n28203 ;
  assign n37014 = ~n37010 & ~n37011 ;
  assign n37012 = \sice_ICYC_reg[2]/NET0131  & n23409 ;
  assign n37013 = \sice_IIRC_reg[2]/NET0131  & n24267 ;
  assign n37015 = ~n37012 & ~n37013 ;
  assign n37016 = n37014 & n37015 ;
  assign n37017 = n34827 & n37016 ;
  assign n37006 = \sice_SPC_reg[1]/P0001  & n34825 ;
  assign n37007 = \sice_SPC_reg[3]/P0001  & ~n34825 ;
  assign n37008 = ~n37006 & ~n37007 ;
  assign n37009 = ~n34827 & n37008 ;
  assign n37018 = n26297 & ~n37009 ;
  assign n37019 = ~n37017 & n37018 ;
  assign n37020 = ~n37005 & ~n37019 ;
  assign n37021 = \sice_SPC_reg[1]/P0001  & ~n26297 ;
  assign n37026 = \sice_idr0_reg_DO_reg[1]/P0001  & n26968 ;
  assign n37027 = \core_c_dec_IR_reg[1]/NET0131  & n28203 ;
  assign n37030 = ~n37026 & ~n37027 ;
  assign n37028 = \sice_ICYC_reg[1]/NET0131  & n23409 ;
  assign n37029 = \sice_IIRC_reg[1]/NET0131  & n24267 ;
  assign n37031 = ~n37028 & ~n37029 ;
  assign n37032 = n37030 & n37031 ;
  assign n37033 = n34827 & n37032 ;
  assign n37022 = \sice_SPC_reg[0]/P0001  & n34825 ;
  assign n37023 = \sice_SPC_reg[2]/P0001  & ~n34825 ;
  assign n37024 = ~n37022 & ~n37023 ;
  assign n37025 = ~n34827 & n37024 ;
  assign n37034 = n26297 & ~n37025 ;
  assign n37035 = ~n37033 & n37034 ;
  assign n37036 = ~n37021 & ~n37035 ;
  assign n37037 = n14752 & n31574 ;
  assign n37038 = ~\core_eu_em_mac_em_reg_mr2rwe_DO_reg[3]/P0001  & ~n17799 ;
  assign n37039 = ~n17809 & n21663 ;
  assign n37040 = n17811 & ~n37039 ;
  assign n37041 = ~n37038 & ~n37040 ;
  assign n37042 = ~n17823 & ~n37041 ;
  assign n37043 = ~\core_eu_em_mac_em_reg_mr2rwe_DO_reg[3]/P0001  & ~n17808 ;
  assign n37044 = ~n37042 & ~n37043 ;
  assign n37045 = n17829 & ~n37044 ;
  assign n37046 = ~n37037 & ~n37045 ;
  assign n37047 = ~\clkc_STDcnt_reg[0]/NET0131  & ~n31521 ;
  assign n37048 = ~\clkc_STDcnt_reg[9]/NET0131  & ~n31529 ;
  assign n37049 = ~n31521 & ~n31530 ;
  assign n37050 = ~n37048 & n37049 ;
  assign n37053 = ~n31031 & ~n34353 ;
  assign n37054 = ~n34354 & ~n37053 ;
  assign n37056 = ~n31044 & n37054 ;
  assign n37055 = n31044 & ~n37054 ;
  assign n37057 = n20875 & ~n37055 ;
  assign n37058 = ~n37056 & n37057 ;
  assign n37059 = ~\sport0_rxctl_ldRX_cmp_reg/P0001  & n11265 ;
  assign n37052 = \sport0_rxctl_RX_reg[7]/P0001  & n20873 ;
  assign n37060 = ~n20868 & ~n37052 ;
  assign n37061 = ~n37059 & n37060 ;
  assign n37062 = ~n37058 & n37061 ;
  assign n37051 = ~\sport0_rxctl_RXSHT_reg[7]/P0001  & n20868 ;
  assign n37063 = ~n20871 & ~n37051 ;
  assign n37064 = ~n37062 & n37063 ;
  assign n37065 = \sport0_rxctl_RX_reg[7]/P0001  & n20871 ;
  assign n37066 = ~n37064 & ~n37065 ;
  assign n37067 = \core_c_dec_MTSR1_E_reg/P0001  & ~n20259 ;
  assign n37068 = ~\core_c_dec_MTSR1_E_reg/P0001  & n29085 ;
  assign n37069 = ~n37067 & ~n37068 ;
  assign n37070 = n18717 & ~n37069 ;
  assign n37071 = ~\core_eu_es_sht_es_reg_sr1swe_DO_reg[5]/P0001  & ~n18717 ;
  assign n37072 = ~n37070 & ~n37071 ;
  assign n37073 = \core_c_dec_MTSR1_E_reg/P0001  & ~n19559 ;
  assign n37074 = ~\core_c_dec_MTSR1_E_reg/P0001  & n30613 ;
  assign n37075 = ~n37073 & ~n37074 ;
  assign n37076 = n18717 & ~n37075 ;
  assign n37077 = ~\core_eu_es_sht_es_reg_sr1swe_DO_reg[0]/P0001  & ~n18717 ;
  assign n37078 = ~n37076 & ~n37077 ;
  assign n37079 = n17833 & ~n37075 ;
  assign n37080 = ~\core_eu_es_sht_es_reg_sr1rwe_DO_reg[0]/P0001  & ~n17833 ;
  assign n37081 = ~n37079 & ~n37080 ;
  assign n37082 = \core_c_dec_MTSR0_E_reg/P0001  & ~n23920 ;
  assign n37083 = ~\core_c_dec_MTSR0_E_reg/P0001  & n30089 ;
  assign n37084 = ~n37082 & ~n37083 ;
  assign n37085 = n18886 & ~n37084 ;
  assign n37086 = ~\core_eu_es_sht_es_reg_sr0swe_DO_reg[12]/P0001  & ~n18886 ;
  assign n37087 = ~n37085 & ~n37086 ;
  assign n37088 = n19034 & ~n37084 ;
  assign n37089 = ~\core_eu_es_sht_es_reg_sr0rwe_DO_reg[12]/P0001  & ~n19034 ;
  assign n37090 = ~n37088 & ~n37089 ;
  assign n37093 = n18271 & ~n19972 ;
  assign n37092 = ~\core_eu_em_mac_em_reg_mr0swe_DO_reg[7]/P0001  & ~n18271 ;
  assign n37094 = n18273 & ~n37092 ;
  assign n37095 = ~n37093 & n37094 ;
  assign n37091 = \core_eu_em_mac_em_reg_mr0swe_DO_reg[7]/P0001  & ~n18266 ;
  assign n37096 = ~n18270 & ~n37091 ;
  assign n37097 = ~n37095 & n37096 ;
  assign n37098 = ~n18262 & ~n37097 ;
  assign n37099 = n18262 & ~n19623 ;
  assign n37100 = ~n37098 & ~n37099 ;
  assign n37101 = n14752 & n19623 ;
  assign n37102 = n18328 & n19972 ;
  assign n37103 = \core_eu_em_mac_em_reg_mr0rwe_DO_reg[7]/P0001  & ~n18330 ;
  assign n37104 = n18334 & ~n37103 ;
  assign n37105 = ~n37102 & n37104 ;
  assign n37106 = ~n37101 & ~n37105 ;
  assign n37109 = ~n34363 & ~n34396 ;
  assign n37110 = ~n34397 & ~n37109 ;
  assign n37112 = ~n34399 & n37110 ;
  assign n37111 = n34399 & ~n37110 ;
  assign n37113 = n20875 & ~n37111 ;
  assign n37114 = ~n37112 & n37113 ;
  assign n37115 = ~\sport0_rxctl_ldRX_cmp_reg/P0001  & n10289 ;
  assign n37108 = \sport0_rxctl_RX_reg[9]/P0001  & n20873 ;
  assign n37116 = ~n20868 & ~n37108 ;
  assign n37117 = ~n37115 & n37116 ;
  assign n37118 = ~n37114 & n37117 ;
  assign n37107 = ~\sport0_rxctl_RXSHT_reg[9]/P0001  & n20868 ;
  assign n37119 = ~n20871 & ~n37107 ;
  assign n37120 = ~n37118 & n37119 ;
  assign n37121 = \sport0_rxctl_RX_reg[9]/P0001  & n20871 ;
  assign n37122 = ~n37120 & ~n37121 ;
  assign n37123 = n17833 & ~n37069 ;
  assign n37124 = ~\core_eu_es_sht_es_reg_sr1rwe_DO_reg[5]/P0001  & ~n17833 ;
  assign n37125 = ~n37123 & ~n37124 ;
  assign n37126 = \core_c_dec_MTSR0_E_reg/P0001  & ~n19972 ;
  assign n37127 = ~\core_c_dec_MTSR0_E_reg/P0001  & n30245 ;
  assign n37128 = ~n37126 & ~n37127 ;
  assign n37129 = n18886 & ~n37128 ;
  assign n37130 = ~\core_eu_es_sht_es_reg_sr0swe_DO_reg[7]/P0001  & ~n18886 ;
  assign n37131 = ~n37129 & ~n37130 ;
  assign n37132 = \core_c_dec_MTSR0_E_reg/P0001  & ~n23757 ;
  assign n37133 = ~\core_c_dec_MTSR0_E_reg/P0001  & n29776 ;
  assign n37134 = ~n37132 & ~n37133 ;
  assign n37135 = n18886 & ~n37134 ;
  assign n37136 = ~\core_eu_es_sht_es_reg_sr0swe_DO_reg[11]/P0001  & ~n18886 ;
  assign n37137 = ~n37135 & ~n37136 ;
  assign n37138 = n19034 & ~n37128 ;
  assign n37139 = ~\core_eu_es_sht_es_reg_sr0rwe_DO_reg[7]/P0001  & ~n19034 ;
  assign n37140 = ~n37138 & ~n37139 ;
  assign n37141 = n19034 & ~n37134 ;
  assign n37142 = ~\core_eu_es_sht_es_reg_sr0rwe_DO_reg[11]/P0001  & ~n19034 ;
  assign n37143 = ~n37141 & ~n37142 ;
  assign n37144 = ~\clkc_STDcnt_reg[5]/NET0131  & ~n31525 ;
  assign n37145 = ~n31521 & ~n31526 ;
  assign n37146 = ~n37144 & n37145 ;
  assign n37147 = ~\clkc_STDcnt_reg[2]/NET0131  & ~n31522 ;
  assign n37148 = ~n31523 & ~n37147 ;
  assign n37149 = ~n31521 & n37148 ;
  assign n37150 = ~n25833 & ~n25835 ;
  assign n37151 = ~n22424 & n37150 ;
  assign n37152 = n22424 & ~n37150 ;
  assign n37153 = ~n37151 & ~n37152 ;
  assign n37154 = n22411 & ~n37153 ;
  assign n37155 = \tm_TCR_TMP_reg[11]/NET0131  & ~n22411 ;
  assign n37156 = ~n37154 & ~n37155 ;
  assign n37157 = ~n22400 & ~n37156 ;
  assign n37158 = \tm_tpr_reg_DO_reg[11]/NET0131  & n22400 ;
  assign n37159 = ~n37157 & ~n37158 ;
  assign n37160 = ~n20355 & ~n37159 ;
  assign n37161 = \tm_tcr_reg_DO_reg[11]/NET0131  & n20355 ;
  assign n37162 = ~n37160 & ~n37161 ;
  assign n37163 = \T_ED[1]_pad  & n34066 ;
  assign n37164 = \bdma_BCTL_reg[0]/NET0131  & \bdma_BCTL_reg[1]/NET0131  ;
  assign n37165 = ~n34061 & n37164 ;
  assign n37166 = ~n34066 & ~n37165 ;
  assign n37167 = \bdma_BRdataBUF_reg[9]/P0001  & n37166 ;
  assign n37168 = ~n37163 & ~n37167 ;
  assign n37169 = \T_ED[0]_pad  & n34066 ;
  assign n37170 = \bdma_BRdataBUF_reg[8]/P0001  & n37166 ;
  assign n37171 = ~n37169 & ~n37170 ;
  assign n37172 = \T_ED[7]_pad  & n34066 ;
  assign n37173 = \bdma_BRdataBUF_reg[15]/P0001  & n37166 ;
  assign n37174 = ~n37172 & ~n37173 ;
  assign n37175 = \T_ED[6]_pad  & n34066 ;
  assign n37176 = \bdma_BRdataBUF_reg[14]/P0001  & n37166 ;
  assign n37177 = ~n37175 & ~n37176 ;
  assign n37178 = \T_ED[5]_pad  & n34066 ;
  assign n37179 = \bdma_BRdataBUF_reg[13]/P0001  & n37166 ;
  assign n37180 = ~n37178 & ~n37179 ;
  assign n37181 = \T_ED[4]_pad  & n34066 ;
  assign n37182 = \bdma_BRdataBUF_reg[12]/P0001  & n37166 ;
  assign n37183 = ~n37181 & ~n37182 ;
  assign n37184 = \T_ED[3]_pad  & n34066 ;
  assign n37185 = \bdma_BRdataBUF_reg[11]/P0001  & n37166 ;
  assign n37186 = ~n37184 & ~n37185 ;
  assign n37187 = \T_ED[2]_pad  & n34066 ;
  assign n37188 = \bdma_BRdataBUF_reg[10]/P0001  & n37166 ;
  assign n37189 = ~n37187 & ~n37188 ;
  assign n37190 = \sice_SPC_reg[0]/P0001  & ~n26297 ;
  assign n37191 = \sice_idr0_reg_DO_reg[0]/P0001  & n26968 ;
  assign n37192 = \sice_ICYC_reg[0]/NET0131  & n23409 ;
  assign n37195 = ~n37191 & ~n37192 ;
  assign n37193 = \sice_IIRC_reg[0]/NET0131  & n24267 ;
  assign n37194 = \core_c_dec_IR_reg[0]/NET0131  & n28203 ;
  assign n37196 = ~n37193 & ~n37194 ;
  assign n37197 = n37195 & n37196 ;
  assign n37198 = n34827 & ~n37197 ;
  assign n37199 = \sice_SPC_reg[1]/P0001  & ~n28982 ;
  assign n37200 = ~n37198 & ~n37199 ;
  assign n37201 = n26297 & ~n37200 ;
  assign n37202 = ~n37190 & ~n37201 ;
  assign n37203 = ~\clkc_STDcnt_reg[0]/NET0131  & ~\clkc_STDcnt_reg[1]/NET0131  ;
  assign n37204 = ~n31522 & ~n37203 ;
  assign n37205 = ~n31521 & n37204 ;
  assign n37206 = \sport0_regs_MWORDreg_DO_reg[9]/NET0131  & n28944 ;
  assign n37207 = \sport1_regs_MWORDreg_DO_reg[9]/NET0131  & n28854 ;
  assign n37208 = \core_c_dec_updMF_E_reg/P0001  & n4118 ;
  assign n37209 = n18848 & n20378 ;
  assign n37210 = ~n37208 & ~n37209 ;
  assign n37211 = \core_c_psq_SSTAT_reg[0]/NET0131  & n21137 ;
  assign n37212 = ~n36434 & ~n37211 ;
  assign n37213 = ~n4218 & n36435 ;
  assign n37214 = ~n37212 & ~n37213 ;
  assign n37215 = ~n36073 & ~n36075 ;
  assign n37216 = \sport1_regs_SCTLreg_DO_reg[3]/NET0131  & n37215 ;
  assign n37217 = n7270 & n18235 ;
  assign n37218 = n36073 & ~n37217 ;
  assign n37219 = n8113 & n37218 ;
  assign n37220 = ~n37216 & ~n37219 ;
  assign n37221 = \sport1_regs_SCTLreg_DO_reg[2]/NET0131  & n37215 ;
  assign n37222 = n8715 & n37218 ;
  assign n37223 = ~n37221 & ~n37222 ;
  assign n37224 = \sport0_regs_SCTLreg_DO_reg[3]/NET0131  & n18233 ;
  assign n37225 = n8113 & n18237 ;
  assign n37226 = ~n37224 & ~n37225 ;
  assign n37227 = \sport0_regs_SCTLreg_DO_reg[2]/NET0131  & n18233 ;
  assign n37228 = n8715 & n18237 ;
  assign n37229 = ~n37227 & ~n37228 ;
  assign n37230 = ~\idma_IAL_reg/P0001  & n12688 ;
  assign n37231 = \idma_IADi_reg[14]/P0001  & \idma_IAL_reg/P0001  ;
  assign n37232 = ~n37230 & ~n37231 ;
  assign n37233 = n32455 & ~n37232 ;
  assign n37234 = \idma_DCTL_reg[14]/NET0131  & ~n32455 ;
  assign n37235 = ~n37233 & ~n37234 ;
  assign n37236 = \core_c_psq_Iact_E_reg[6]/NET0131  & ~n19477 ;
  assign n37237 = ~n19488 & n19493 ;
  assign n37238 = n19487 & n37237 ;
  assign n37239 = ~n37236 & ~n37238 ;
  assign n37240 = \bdma_BEAD_reg[11]/NET0131  & \bdma_BM_cyc_reg/P0001  ;
  assign n37243 = \core_dag_ilm2reg_PMA_pi_DO_reg[11]/NET0131  & ~n5608 ;
  assign n37241 = \core_dag_ilm1reg_DMA_pi_DO_reg[11]/NET0131  & n5602 ;
  assign n37242 = \emc_ECMA_reg[11]/P0001  & \emc_ECMcs_reg/NET0131  ;
  assign n37244 = ~n37241 & ~n37242 ;
  assign n37245 = ~n37243 & n37244 ;
  assign n37246 = ~\bdma_BM_cyc_reg/P0001  & ~n37245 ;
  assign n37247 = ~n37240 & ~n37246 ;
  assign n37248 = n36427 & ~n36440 ;
  assign n37249 = n4190 & n37248 ;
  assign n37250 = \core_c_psq_pcstk_cnts16x14_PCcell_reg[2][7]/P0001  & ~n37249 ;
  assign n37251 = ~\core_c_dec_MTtoppcs_Eg_reg/P0001  & n5355 ;
  assign n37252 = \core_c_dec_MTtoppcs_Eg_reg/P0001  & n11265 ;
  assign n37253 = ~n37251 & ~n37252 ;
  assign n37254 = ~\core_c_psq_TRAP_Eg_reg/NET0131  & ~n37253 ;
  assign n37255 = \core_c_psq_EXA_reg[7]/P0001  & \core_c_psq_TRAP_Eg_reg/NET0131  ;
  assign n37256 = ~n37254 & ~n37255 ;
  assign n37257 = n37249 & ~n37256 ;
  assign n37258 = ~n37250 & ~n37257 ;
  assign n37259 = \core_c_psq_pcstk_cnts16x14_PCcell_reg[2][5]/P0001  & ~n37249 ;
  assign n37260 = ~\core_c_dec_MTtoppcs_Eg_reg/P0001  & n5304 ;
  assign n37261 = \core_c_dec_MTtoppcs_Eg_reg/P0001  & n10911 ;
  assign n37262 = ~n37260 & ~n37261 ;
  assign n37263 = ~\core_c_psq_TRAP_Eg_reg/NET0131  & ~n37262 ;
  assign n37264 = \core_c_psq_EXA_reg[5]/P0001  & \core_c_psq_TRAP_Eg_reg/NET0131  ;
  assign n37265 = ~n37263 & ~n37264 ;
  assign n37266 = n37249 & ~n37265 ;
  assign n37267 = ~n37259 & ~n37266 ;
  assign n37268 = \core_c_psq_pcstk_cnts16x14_PCcell_reg[2][4]/P0001  & ~n37249 ;
  assign n37269 = ~\core_c_dec_MTtoppcs_Eg_reg/P0001  & n5270 ;
  assign n37270 = \core_c_dec_MTtoppcs_Eg_reg/P0001  & n10069 ;
  assign n37271 = ~n37269 & ~n37270 ;
  assign n37272 = ~\core_c_psq_TRAP_Eg_reg/NET0131  & ~n37271 ;
  assign n37273 = \core_c_psq_EXA_reg[4]/P0001  & \core_c_psq_TRAP_Eg_reg/NET0131  ;
  assign n37274 = ~n37272 & ~n37273 ;
  assign n37275 = n37249 & ~n37274 ;
  assign n37276 = ~n37268 & ~n37275 ;
  assign n37277 = \core_c_psq_pcstk_cnts16x14_PCcell_reg[2][3]/P0001  & ~n37249 ;
  assign n37278 = ~\core_c_dec_MTtoppcs_Eg_reg/P0001  & n5233 ;
  assign n37279 = \core_c_dec_MTtoppcs_Eg_reg/P0001  & n8113 ;
  assign n37280 = ~n37278 & ~n37279 ;
  assign n37281 = ~\core_c_psq_TRAP_Eg_reg/NET0131  & ~n37280 ;
  assign n37282 = \core_c_psq_EXA_reg[3]/P0001  & \core_c_psq_TRAP_Eg_reg/NET0131  ;
  assign n37283 = ~n37281 & ~n37282 ;
  assign n37284 = n37249 & ~n37283 ;
  assign n37285 = ~n37277 & ~n37284 ;
  assign n37286 = \core_c_psq_pcstk_cnts16x14_PCcell_reg[2][1]/P0001  & ~n37249 ;
  assign n37287 = ~\core_c_dec_MTtoppcs_Eg_reg/P0001  & n5158 ;
  assign n37288 = \core_c_dec_MTtoppcs_Eg_reg/P0001  & n9435 ;
  assign n37289 = ~n37287 & ~n37288 ;
  assign n37290 = ~\core_c_psq_TRAP_Eg_reg/NET0131  & ~n37289 ;
  assign n37291 = \core_c_psq_EXA_reg[1]/P0001  & \core_c_psq_TRAP_Eg_reg/NET0131  ;
  assign n37292 = ~n37290 & ~n37291 ;
  assign n37293 = n37249 & ~n37292 ;
  assign n37294 = ~n37286 & ~n37293 ;
  assign n37295 = \core_c_psq_pcstk_cnts16x14_PCcell_reg[2][11]/P0001  & ~n37249 ;
  assign n37296 = ~\core_c_dec_MTtoppcs_Eg_reg/P0001  & n5131 ;
  assign n37297 = \core_c_dec_MTtoppcs_Eg_reg/P0001  & n8460 ;
  assign n37298 = ~n37296 & ~n37297 ;
  assign n37299 = ~\core_c_psq_TRAP_Eg_reg/NET0131  & ~n37298 ;
  assign n37300 = \core_c_psq_EXA_reg[11]/P0001  & \core_c_psq_TRAP_Eg_reg/NET0131  ;
  assign n37301 = ~n37299 & ~n37300 ;
  assign n37302 = n37249 & ~n37301 ;
  assign n37303 = ~n37295 & ~n37302 ;
  assign n37304 = \core_c_psq_pcstk_cnts16x14_PCcell_reg[2][10]/P0001  & ~n37249 ;
  assign n37305 = ~\core_c_dec_MTtoppcs_Eg_reg/P0001  & n5093 ;
  assign n37306 = \core_c_dec_MTtoppcs_Eg_reg/P0001  & n7859 ;
  assign n37307 = ~n37305 & ~n37306 ;
  assign n37308 = ~\core_c_psq_TRAP_Eg_reg/NET0131  & ~n37307 ;
  assign n37309 = \core_c_psq_EXA_reg[10]/P0001  & \core_c_psq_TRAP_Eg_reg/NET0131  ;
  assign n37310 = ~n37308 & ~n37309 ;
  assign n37311 = n37249 & ~n37310 ;
  assign n37312 = ~n37304 & ~n37311 ;
  assign n37313 = ~\core_c_dec_MTtoppcs_Eg_reg/P0001  & ~\core_c_psq_EXA_reg[0]/P0001  ;
  assign n37314 = \core_c_dec_MTtoppcs_Eg_reg/P0001  & n7607 ;
  assign n37315 = ~n37313 & ~n37314 ;
  assign n37316 = ~\core_c_psq_TRAP_Eg_reg/NET0131  & ~n37315 ;
  assign n37317 = \core_c_psq_EXA_reg[0]/P0001  & \core_c_psq_TRAP_Eg_reg/NET0131  ;
  assign n37318 = ~n37316 & ~n37317 ;
  assign n37319 = n37249 & ~n37318 ;
  assign n37320 = \core_c_psq_pcstk_cnts16x14_PCcell_reg[2][0]/P0001  & ~n37249 ;
  assign n37321 = ~n37319 & ~n37320 ;
  assign n37322 = n4218 & n37248 ;
  assign n37323 = \core_c_psq_pcstk_cnts16x14_PCcell_reg[1][9]/P0001  & ~n37322 ;
  assign n37324 = ~\core_c_dec_MTtoppcs_Eg_reg/P0001  & n5409 ;
  assign n37325 = \core_c_dec_MTtoppcs_Eg_reg/P0001  & n10289 ;
  assign n37326 = ~n37324 & ~n37325 ;
  assign n37327 = ~\core_c_psq_TRAP_Eg_reg/NET0131  & ~n37326 ;
  assign n37328 = \core_c_psq_EXA_reg[9]/P0001  & \core_c_psq_TRAP_Eg_reg/NET0131  ;
  assign n37329 = ~n37327 & ~n37328 ;
  assign n37330 = n37322 & ~n37329 ;
  assign n37331 = ~n37323 & ~n37330 ;
  assign n37332 = \core_c_psq_pcstk_cnts16x14_PCcell_reg[1][8]/P0001  & ~n37322 ;
  assign n37333 = ~\core_c_dec_MTtoppcs_Eg_reg/P0001  & n5382 ;
  assign n37334 = \core_c_dec_MTtoppcs_Eg_reg/P0001  & n10638 ;
  assign n37335 = ~n37333 & ~n37334 ;
  assign n37336 = ~\core_c_psq_TRAP_Eg_reg/NET0131  & ~n37335 ;
  assign n37337 = \core_c_psq_EXA_reg[8]/P0001  & \core_c_psq_TRAP_Eg_reg/NET0131  ;
  assign n37338 = ~n37336 & ~n37337 ;
  assign n37339 = n37322 & ~n37338 ;
  assign n37340 = ~n37332 & ~n37339 ;
  assign n37341 = \core_c_psq_pcstk_cnts16x14_PCcell_reg[1][7]/P0001  & ~n37322 ;
  assign n37342 = ~n37256 & n37322 ;
  assign n37343 = ~n37341 & ~n37342 ;
  assign n37344 = \core_c_psq_pcstk_cnts16x14_PCcell_reg[1][6]/P0001  & ~n37322 ;
  assign n37345 = ~\core_c_dec_MTtoppcs_Eg_reg/P0001  & n5328 ;
  assign n37346 = \core_c_dec_MTtoppcs_Eg_reg/P0001  & n11525 ;
  assign n37347 = ~n37345 & ~n37346 ;
  assign n37348 = ~\core_c_psq_TRAP_Eg_reg/NET0131  & ~n37347 ;
  assign n37349 = \core_c_psq_EXA_reg[6]/P0001  & \core_c_psq_TRAP_Eg_reg/NET0131  ;
  assign n37350 = ~n37348 & ~n37349 ;
  assign n37351 = n37322 & ~n37350 ;
  assign n37352 = ~n37344 & ~n37351 ;
  assign n37353 = \core_c_psq_pcstk_cnts16x14_PCcell_reg[1][3]/P0001  & ~n37322 ;
  assign n37354 = ~n37283 & n37322 ;
  assign n37355 = ~n37353 & ~n37354 ;
  assign n37356 = \core_c_psq_pcstk_cnts16x14_PCcell_reg[1][2]/P0001  & ~n37322 ;
  assign n37357 = ~\core_c_dec_MTtoppcs_Eg_reg/P0001  & n5195 ;
  assign n37358 = \core_c_dec_MTtoppcs_Eg_reg/P0001  & n8715 ;
  assign n37359 = ~n37357 & ~n37358 ;
  assign n37360 = ~\core_c_psq_TRAP_Eg_reg/NET0131  & ~n37359 ;
  assign n37361 = \core_c_psq_EXA_reg[2]/P0001  & \core_c_psq_TRAP_Eg_reg/NET0131  ;
  assign n37362 = ~n37360 & ~n37361 ;
  assign n37363 = n37322 & ~n37362 ;
  assign n37364 = ~n37356 & ~n37363 ;
  assign n37365 = \core_c_psq_pcstk_cnts16x14_PCcell_reg[1][1]/P0001  & ~n37322 ;
  assign n37366 = ~n37292 & n37322 ;
  assign n37367 = ~n37365 & ~n37366 ;
  assign n37368 = \core_c_psq_pcstk_cnts16x14_PCcell_reg[1][13]/P0001  & ~n37322 ;
  assign n37369 = ~\core_c_dec_MTtoppcs_Eg_reg/P0001  & n5649 ;
  assign n37370 = \core_c_dec_MTtoppcs_Eg_reg/P0001  & n7340 ;
  assign n37371 = ~n37369 & ~n37370 ;
  assign n37372 = ~\core_c_psq_TRAP_Eg_reg/NET0131  & ~n37371 ;
  assign n37373 = \core_c_psq_EXA_reg[13]/P0001  & \core_c_psq_TRAP_Eg_reg/NET0131  ;
  assign n37374 = ~n37372 & ~n37373 ;
  assign n37375 = n37322 & ~n37374 ;
  assign n37376 = ~n37368 & ~n37375 ;
  assign n37377 = \core_c_psq_pcstk_cnts16x14_PCcell_reg[1][12]/P0001  & ~n37322 ;
  assign n37378 = ~\core_c_dec_MTtoppcs_Eg_reg/P0001  & n5624 ;
  assign n37379 = \core_c_dec_MTtoppcs_Eg_reg/P0001  & n9178 ;
  assign n37380 = ~n37378 & ~n37379 ;
  assign n37381 = ~\core_c_psq_TRAP_Eg_reg/NET0131  & ~n37380 ;
  assign n37382 = \core_c_psq_EXA_reg[12]/P0001  & \core_c_psq_TRAP_Eg_reg/NET0131  ;
  assign n37383 = ~n37381 & ~n37382 ;
  assign n37384 = n37322 & ~n37383 ;
  assign n37385 = ~n37377 & ~n37384 ;
  assign n37386 = \core_c_psq_pcstk_cnts16x14_PCcell_reg[1][11]/P0001  & ~n37322 ;
  assign n37387 = ~n37301 & n37322 ;
  assign n37388 = ~n37386 & ~n37387 ;
  assign n37389 = \core_c_psq_pcstk_cnts16x14_PCcell_reg[1][10]/P0001  & ~n37322 ;
  assign n37390 = ~n37310 & n37322 ;
  assign n37391 = ~n37389 & ~n37390 ;
  assign n37392 = ~n37318 & n37322 ;
  assign n37393 = \core_c_psq_pcstk_cnts16x14_PCcell_reg[1][0]/P0001  & ~n37322 ;
  assign n37394 = ~n37392 & ~n37393 ;
  assign n37395 = n4222 & n37248 ;
  assign n37396 = \core_c_psq_pcstk_cnts16x14_PCcell_reg[15][9]/P0001  & ~n37395 ;
  assign n37397 = ~n37329 & n37395 ;
  assign n37398 = ~n37396 & ~n37397 ;
  assign n37399 = \core_c_psq_pcstk_cnts16x14_PCcell_reg[15][8]/P0001  & ~n37395 ;
  assign n37400 = ~n37338 & n37395 ;
  assign n37401 = ~n37399 & ~n37400 ;
  assign n37402 = \core_c_psq_pcstk_cnts16x14_PCcell_reg[15][7]/P0001  & ~n37395 ;
  assign n37403 = ~n37256 & n37395 ;
  assign n37404 = ~n37402 & ~n37403 ;
  assign n37405 = \core_c_psq_pcstk_cnts16x14_PCcell_reg[15][6]/P0001  & ~n37395 ;
  assign n37406 = ~n37350 & n37395 ;
  assign n37407 = ~n37405 & ~n37406 ;
  assign n37408 = \core_c_psq_pcstk_cnts16x14_PCcell_reg[15][5]/P0001  & ~n37395 ;
  assign n37409 = ~n37265 & n37395 ;
  assign n37410 = ~n37408 & ~n37409 ;
  assign n37411 = \core_c_psq_pcstk_cnts16x14_PCcell_reg[15][4]/P0001  & ~n37395 ;
  assign n37412 = ~n37274 & n37395 ;
  assign n37413 = ~n37411 & ~n37412 ;
  assign n37414 = \core_c_psq_pcstk_cnts16x14_PCcell_reg[15][3]/P0001  & ~n37395 ;
  assign n37415 = ~n37283 & n37395 ;
  assign n37416 = ~n37414 & ~n37415 ;
  assign n37417 = \core_c_psq_pcstk_cnts16x14_PCcell_reg[15][2]/P0001  & ~n37395 ;
  assign n37418 = ~n37362 & n37395 ;
  assign n37419 = ~n37417 & ~n37418 ;
  assign n37420 = \core_c_psq_pcstk_cnts16x14_PCcell_reg[15][1]/P0001  & ~n37395 ;
  assign n37421 = ~n37292 & n37395 ;
  assign n37422 = ~n37420 & ~n37421 ;
  assign n37423 = \core_c_psq_pcstk_cnts16x14_PCcell_reg[15][13]/P0001  & ~n37395 ;
  assign n37424 = ~n37374 & n37395 ;
  assign n37425 = ~n37423 & ~n37424 ;
  assign n37426 = \core_c_psq_pcstk_cnts16x14_PCcell_reg[15][12]/P0001  & ~n37395 ;
  assign n37427 = ~n37383 & n37395 ;
  assign n37428 = ~n37426 & ~n37427 ;
  assign n37429 = \core_c_psq_pcstk_cnts16x14_PCcell_reg[15][11]/P0001  & ~n37395 ;
  assign n37430 = ~n37301 & n37395 ;
  assign n37431 = ~n37429 & ~n37430 ;
  assign n37432 = \core_c_psq_pcstk_cnts16x14_PCcell_reg[15][10]/P0001  & ~n37395 ;
  assign n37433 = ~n37310 & n37395 ;
  assign n37434 = ~n37432 & ~n37433 ;
  assign n37435 = ~n37318 & n37395 ;
  assign n37436 = \core_c_psq_pcstk_cnts16x14_PCcell_reg[15][0]/P0001  & ~n37395 ;
  assign n37437 = ~n37435 & ~n37436 ;
  assign n37438 = n4224 & n37248 ;
  assign n37439 = \core_c_psq_pcstk_cnts16x14_PCcell_reg[14][9]/P0001  & ~n37438 ;
  assign n37440 = ~n37329 & n37438 ;
  assign n37441 = ~n37439 & ~n37440 ;
  assign n37442 = \core_c_psq_pcstk_cnts16x14_PCcell_reg[14][8]/P0001  & ~n37438 ;
  assign n37443 = ~n37338 & n37438 ;
  assign n37444 = ~n37442 & ~n37443 ;
  assign n37445 = \core_c_psq_pcstk_cnts16x14_PCcell_reg[14][7]/P0001  & ~n37438 ;
  assign n37446 = ~n37256 & n37438 ;
  assign n37447 = ~n37445 & ~n37446 ;
  assign n37448 = \core_c_psq_pcstk_cnts16x14_PCcell_reg[14][6]/P0001  & ~n37438 ;
  assign n37449 = ~n37350 & n37438 ;
  assign n37450 = ~n37448 & ~n37449 ;
  assign n37451 = \core_c_psq_pcstk_cnts16x14_PCcell_reg[14][5]/P0001  & ~n37438 ;
  assign n37452 = ~n37265 & n37438 ;
  assign n37453 = ~n37451 & ~n37452 ;
  assign n37454 = \core_c_psq_pcstk_cnts16x14_PCcell_reg[14][4]/P0001  & ~n37438 ;
  assign n37455 = ~n37274 & n37438 ;
  assign n37456 = ~n37454 & ~n37455 ;
  assign n37457 = \core_c_psq_pcstk_cnts16x14_PCcell_reg[14][3]/P0001  & ~n37438 ;
  assign n37458 = ~n37283 & n37438 ;
  assign n37459 = ~n37457 & ~n37458 ;
  assign n37460 = \core_c_psq_pcstk_cnts16x14_PCcell_reg[14][2]/P0001  & ~n37438 ;
  assign n37461 = ~n37362 & n37438 ;
  assign n37462 = ~n37460 & ~n37461 ;
  assign n37463 = \core_c_psq_pcstk_cnts16x14_PCcell_reg[14][1]/P0001  & ~n37438 ;
  assign n37464 = ~n37292 & n37438 ;
  assign n37465 = ~n37463 & ~n37464 ;
  assign n37466 = \core_c_psq_pcstk_cnts16x14_PCcell_reg[14][13]/P0001  & ~n37438 ;
  assign n37467 = ~n37374 & n37438 ;
  assign n37468 = ~n37466 & ~n37467 ;
  assign n37469 = \core_c_psq_pcstk_cnts16x14_PCcell_reg[14][12]/P0001  & ~n37438 ;
  assign n37470 = ~n37383 & n37438 ;
  assign n37471 = ~n37469 & ~n37470 ;
  assign n37472 = \core_c_psq_pcstk_cnts16x14_PCcell_reg[14][11]/P0001  & ~n37438 ;
  assign n37473 = ~n37301 & n37438 ;
  assign n37474 = ~n37472 & ~n37473 ;
  assign n37475 = \core_c_psq_pcstk_cnts16x14_PCcell_reg[14][10]/P0001  & ~n37438 ;
  assign n37476 = ~n37310 & n37438 ;
  assign n37477 = ~n37475 & ~n37476 ;
  assign n37478 = ~n37318 & n37438 ;
  assign n37479 = \core_c_psq_pcstk_cnts16x14_PCcell_reg[14][0]/P0001  & ~n37438 ;
  assign n37480 = ~n37478 & ~n37479 ;
  assign n37481 = n4194 & n37248 ;
  assign n37482 = \core_c_psq_pcstk_cnts16x14_PCcell_reg[13][9]/P0001  & ~n37481 ;
  assign n37483 = ~n37329 & n37481 ;
  assign n37484 = ~n37482 & ~n37483 ;
  assign n37485 = \core_c_psq_pcstk_cnts16x14_PCcell_reg[13][8]/P0001  & ~n37481 ;
  assign n37486 = ~n37338 & n37481 ;
  assign n37487 = ~n37485 & ~n37486 ;
  assign n37488 = \core_c_psq_pcstk_cnts16x14_PCcell_reg[13][7]/P0001  & ~n37481 ;
  assign n37489 = ~n37256 & n37481 ;
  assign n37490 = ~n37488 & ~n37489 ;
  assign n37491 = \core_c_psq_pcstk_cnts16x14_PCcell_reg[13][6]/P0001  & ~n37481 ;
  assign n37492 = ~n37350 & n37481 ;
  assign n37493 = ~n37491 & ~n37492 ;
  assign n37494 = \core_c_psq_pcstk_cnts16x14_PCcell_reg[13][5]/P0001  & ~n37481 ;
  assign n37495 = ~n37265 & n37481 ;
  assign n37496 = ~n37494 & ~n37495 ;
  assign n37497 = \core_c_psq_pcstk_cnts16x14_PCcell_reg[13][4]/P0001  & ~n37481 ;
  assign n37498 = ~n37274 & n37481 ;
  assign n37499 = ~n37497 & ~n37498 ;
  assign n37500 = \core_c_psq_pcstk_cnts16x14_PCcell_reg[13][3]/P0001  & ~n37481 ;
  assign n37501 = ~n37283 & n37481 ;
  assign n37502 = ~n37500 & ~n37501 ;
  assign n37503 = \core_c_psq_pcstk_cnts16x14_PCcell_reg[13][2]/P0001  & ~n37481 ;
  assign n37504 = ~n37362 & n37481 ;
  assign n37505 = ~n37503 & ~n37504 ;
  assign n37506 = \core_c_psq_pcstk_cnts16x14_PCcell_reg[13][1]/P0001  & ~n37481 ;
  assign n37507 = ~n37292 & n37481 ;
  assign n37508 = ~n37506 & ~n37507 ;
  assign n37509 = \core_c_psq_pcstk_cnts16x14_PCcell_reg[13][13]/P0001  & ~n37481 ;
  assign n37510 = ~n37374 & n37481 ;
  assign n37511 = ~n37509 & ~n37510 ;
  assign n37512 = \core_c_psq_pcstk_cnts16x14_PCcell_reg[13][12]/P0001  & ~n37481 ;
  assign n37513 = ~n37383 & n37481 ;
  assign n37514 = ~n37512 & ~n37513 ;
  assign n37515 = \core_c_psq_pcstk_cnts16x14_PCcell_reg[13][11]/P0001  & ~n37481 ;
  assign n37516 = ~n37301 & n37481 ;
  assign n37517 = ~n37515 & ~n37516 ;
  assign n37518 = \core_c_psq_pcstk_cnts16x14_PCcell_reg[13][10]/P0001  & ~n37481 ;
  assign n37519 = ~n37310 & n37481 ;
  assign n37520 = ~n37518 & ~n37519 ;
  assign n37521 = ~n37318 & n37481 ;
  assign n37522 = \core_c_psq_pcstk_cnts16x14_PCcell_reg[13][0]/P0001  & ~n37481 ;
  assign n37523 = ~n37521 & ~n37522 ;
  assign n37524 = n4205 & n37248 ;
  assign n37525 = \core_c_psq_pcstk_cnts16x14_PCcell_reg[12][9]/P0001  & ~n37524 ;
  assign n37526 = ~n37329 & n37524 ;
  assign n37527 = ~n37525 & ~n37526 ;
  assign n37528 = \core_c_psq_pcstk_cnts16x14_PCcell_reg[12][8]/P0001  & ~n37524 ;
  assign n37529 = ~n37338 & n37524 ;
  assign n37530 = ~n37528 & ~n37529 ;
  assign n37531 = \core_c_psq_pcstk_cnts16x14_PCcell_reg[12][7]/P0001  & ~n37524 ;
  assign n37532 = ~n37256 & n37524 ;
  assign n37533 = ~n37531 & ~n37532 ;
  assign n37534 = \core_c_psq_pcstk_cnts16x14_PCcell_reg[12][6]/P0001  & ~n37524 ;
  assign n37535 = ~n37350 & n37524 ;
  assign n37536 = ~n37534 & ~n37535 ;
  assign n37537 = \core_c_psq_pcstk_cnts16x14_PCcell_reg[12][5]/P0001  & ~n37524 ;
  assign n37538 = ~n37265 & n37524 ;
  assign n37539 = ~n37537 & ~n37538 ;
  assign n37540 = \core_c_psq_pcstk_cnts16x14_PCcell_reg[12][4]/P0001  & ~n37524 ;
  assign n37541 = ~n37274 & n37524 ;
  assign n37542 = ~n37540 & ~n37541 ;
  assign n37543 = \core_c_psq_pcstk_cnts16x14_PCcell_reg[12][3]/P0001  & ~n37524 ;
  assign n37544 = ~n37283 & n37524 ;
  assign n37545 = ~n37543 & ~n37544 ;
  assign n37546 = \core_c_psq_pcstk_cnts16x14_PCcell_reg[12][2]/P0001  & ~n37524 ;
  assign n37547 = ~n37362 & n37524 ;
  assign n37548 = ~n37546 & ~n37547 ;
  assign n37549 = \core_c_psq_pcstk_cnts16x14_PCcell_reg[12][1]/P0001  & ~n37524 ;
  assign n37550 = ~n37292 & n37524 ;
  assign n37551 = ~n37549 & ~n37550 ;
  assign n37552 = \core_c_psq_pcstk_cnts16x14_PCcell_reg[12][13]/P0001  & ~n37524 ;
  assign n37553 = ~n37374 & n37524 ;
  assign n37554 = ~n37552 & ~n37553 ;
  assign n37555 = \core_c_psq_pcstk_cnts16x14_PCcell_reg[12][12]/P0001  & ~n37524 ;
  assign n37556 = ~n37383 & n37524 ;
  assign n37557 = ~n37555 & ~n37556 ;
  assign n37558 = \core_c_psq_pcstk_cnts16x14_PCcell_reg[12][11]/P0001  & ~n37524 ;
  assign n37559 = ~n37301 & n37524 ;
  assign n37560 = ~n37558 & ~n37559 ;
  assign n37561 = \core_c_psq_pcstk_cnts16x14_PCcell_reg[12][10]/P0001  & ~n37524 ;
  assign n37562 = ~n37310 & n37524 ;
  assign n37563 = ~n37561 & ~n37562 ;
  assign n37564 = ~n37318 & n37524 ;
  assign n37565 = \core_c_psq_pcstk_cnts16x14_PCcell_reg[12][0]/P0001  & ~n37524 ;
  assign n37566 = ~n37564 & ~n37565 ;
  assign n37567 = n4202 & n37248 ;
  assign n37568 = \core_c_psq_pcstk_cnts16x14_PCcell_reg[11][9]/P0001  & ~n37567 ;
  assign n37569 = ~n37329 & n37567 ;
  assign n37570 = ~n37568 & ~n37569 ;
  assign n37571 = \core_c_psq_pcstk_cnts16x14_PCcell_reg[11][8]/P0001  & ~n37567 ;
  assign n37572 = ~n37338 & n37567 ;
  assign n37573 = ~n37571 & ~n37572 ;
  assign n37574 = \core_c_psq_pcstk_cnts16x14_PCcell_reg[11][7]/P0001  & ~n37567 ;
  assign n37575 = ~n37256 & n37567 ;
  assign n37576 = ~n37574 & ~n37575 ;
  assign n37577 = \core_c_psq_pcstk_cnts16x14_PCcell_reg[11][6]/P0001  & ~n37567 ;
  assign n37578 = ~n37350 & n37567 ;
  assign n37579 = ~n37577 & ~n37578 ;
  assign n37580 = \core_c_psq_pcstk_cnts16x14_PCcell_reg[11][5]/P0001  & ~n37567 ;
  assign n37581 = ~n37265 & n37567 ;
  assign n37582 = ~n37580 & ~n37581 ;
  assign n37583 = \core_c_psq_pcstk_cnts16x14_PCcell_reg[11][4]/P0001  & ~n37567 ;
  assign n37584 = ~n37274 & n37567 ;
  assign n37585 = ~n37583 & ~n37584 ;
  assign n37586 = \core_c_psq_pcstk_cnts16x14_PCcell_reg[11][3]/P0001  & ~n37567 ;
  assign n37587 = ~n37283 & n37567 ;
  assign n37588 = ~n37586 & ~n37587 ;
  assign n37589 = \core_c_psq_pcstk_cnts16x14_PCcell_reg[11][2]/P0001  & ~n37567 ;
  assign n37590 = ~n37362 & n37567 ;
  assign n37591 = ~n37589 & ~n37590 ;
  assign n37592 = \core_c_psq_pcstk_cnts16x14_PCcell_reg[11][1]/P0001  & ~n37567 ;
  assign n37593 = ~n37292 & n37567 ;
  assign n37594 = ~n37592 & ~n37593 ;
  assign n37595 = \core_c_psq_pcstk_cnts16x14_PCcell_reg[11][13]/P0001  & ~n37567 ;
  assign n37596 = ~n37374 & n37567 ;
  assign n37597 = ~n37595 & ~n37596 ;
  assign n37598 = \core_c_psq_pcstk_cnts16x14_PCcell_reg[11][12]/P0001  & ~n37567 ;
  assign n37599 = ~n37383 & n37567 ;
  assign n37600 = ~n37598 & ~n37599 ;
  assign n37601 = \core_c_psq_pcstk_cnts16x14_PCcell_reg[11][11]/P0001  & ~n37567 ;
  assign n37602 = ~n37301 & n37567 ;
  assign n37603 = ~n37601 & ~n37602 ;
  assign n37604 = \core_c_psq_pcstk_cnts16x14_PCcell_reg[11][10]/P0001  & ~n37567 ;
  assign n37605 = ~n37310 & n37567 ;
  assign n37606 = ~n37604 & ~n37605 ;
  assign n37607 = ~n37318 & n37567 ;
  assign n37608 = \core_c_psq_pcstk_cnts16x14_PCcell_reg[11][0]/P0001  & ~n37567 ;
  assign n37609 = ~n37607 & ~n37608 ;
  assign n37610 = n4228 & n37248 ;
  assign n37611 = \core_c_psq_pcstk_cnts16x14_PCcell_reg[10][9]/P0001  & ~n37610 ;
  assign n37612 = ~n37329 & n37610 ;
  assign n37613 = ~n37611 & ~n37612 ;
  assign n37614 = \core_c_psq_pcstk_cnts16x14_PCcell_reg[10][8]/P0001  & ~n37610 ;
  assign n37615 = ~n37338 & n37610 ;
  assign n37616 = ~n37614 & ~n37615 ;
  assign n37617 = \core_c_psq_pcstk_cnts16x14_PCcell_reg[10][7]/P0001  & ~n37610 ;
  assign n37618 = ~n37256 & n37610 ;
  assign n37619 = ~n37617 & ~n37618 ;
  assign n37620 = \core_c_psq_pcstk_cnts16x14_PCcell_reg[10][6]/P0001  & ~n37610 ;
  assign n37621 = ~n37350 & n37610 ;
  assign n37622 = ~n37620 & ~n37621 ;
  assign n37623 = \core_c_psq_pcstk_cnts16x14_PCcell_reg[10][5]/P0001  & ~n37610 ;
  assign n37624 = ~n37265 & n37610 ;
  assign n37625 = ~n37623 & ~n37624 ;
  assign n37626 = \core_c_psq_pcstk_cnts16x14_PCcell_reg[10][4]/P0001  & ~n37610 ;
  assign n37627 = ~n37274 & n37610 ;
  assign n37628 = ~n37626 & ~n37627 ;
  assign n37629 = \core_c_psq_pcstk_cnts16x14_PCcell_reg[10][3]/P0001  & ~n37610 ;
  assign n37630 = ~n37283 & n37610 ;
  assign n37631 = ~n37629 & ~n37630 ;
  assign n37632 = \core_c_psq_pcstk_cnts16x14_PCcell_reg[10][2]/P0001  & ~n37610 ;
  assign n37633 = ~n37362 & n37610 ;
  assign n37634 = ~n37632 & ~n37633 ;
  assign n37635 = \core_c_psq_pcstk_cnts16x14_PCcell_reg[10][1]/P0001  & ~n37610 ;
  assign n37636 = ~n37292 & n37610 ;
  assign n37637 = ~n37635 & ~n37636 ;
  assign n37638 = \core_c_psq_pcstk_cnts16x14_PCcell_reg[10][13]/P0001  & ~n37610 ;
  assign n37639 = ~n37374 & n37610 ;
  assign n37640 = ~n37638 & ~n37639 ;
  assign n37641 = \core_c_psq_pcstk_cnts16x14_PCcell_reg[10][12]/P0001  & ~n37610 ;
  assign n37642 = ~n37383 & n37610 ;
  assign n37643 = ~n37641 & ~n37642 ;
  assign n37644 = \core_c_psq_pcstk_cnts16x14_PCcell_reg[10][11]/P0001  & ~n37610 ;
  assign n37645 = ~n37301 & n37610 ;
  assign n37646 = ~n37644 & ~n37645 ;
  assign n37647 = \core_c_psq_pcstk_cnts16x14_PCcell_reg[10][10]/P0001  & ~n37610 ;
  assign n37648 = ~n37310 & n37610 ;
  assign n37649 = ~n37647 & ~n37648 ;
  assign n37650 = ~n37318 & n37610 ;
  assign n37651 = \core_c_psq_pcstk_cnts16x14_PCcell_reg[10][0]/P0001  & ~n37610 ;
  assign n37652 = ~n37650 & ~n37651 ;
  assign n37653 = ~n36440 & n36603 ;
  assign n37654 = \core_c_psq_pcstk_cnts16x14_PCcell_reg[0][9]/P0001  & ~n37653 ;
  assign n37655 = ~n37329 & n37653 ;
  assign n37656 = ~n37654 & ~n37655 ;
  assign n37657 = \core_c_psq_pcstk_cnts16x14_PCcell_reg[0][8]/P0001  & ~n37653 ;
  assign n37658 = ~n37338 & n37653 ;
  assign n37659 = ~n37657 & ~n37658 ;
  assign n37660 = \core_c_psq_pcstk_cnts16x14_PCcell_reg[0][7]/P0001  & ~n37653 ;
  assign n37661 = ~n37256 & n37653 ;
  assign n37662 = ~n37660 & ~n37661 ;
  assign n37663 = \core_c_psq_pcstk_cnts16x14_PCcell_reg[0][6]/P0001  & ~n37653 ;
  assign n37664 = ~n37350 & n37653 ;
  assign n37665 = ~n37663 & ~n37664 ;
  assign n37666 = \core_c_psq_pcstk_cnts16x14_PCcell_reg[0][5]/P0001  & ~n37653 ;
  assign n37667 = ~n37265 & n37653 ;
  assign n37668 = ~n37666 & ~n37667 ;
  assign n37669 = \core_c_psq_pcstk_cnts16x14_PCcell_reg[0][4]/P0001  & ~n37653 ;
  assign n37670 = ~n37274 & n37653 ;
  assign n37671 = ~n37669 & ~n37670 ;
  assign n37672 = \core_c_psq_pcstk_cnts16x14_PCcell_reg[0][3]/P0001  & ~n37653 ;
  assign n37673 = ~n37283 & n37653 ;
  assign n37674 = ~n37672 & ~n37673 ;
  assign n37675 = \core_c_psq_pcstk_cnts16x14_PCcell_reg[0][2]/P0001  & ~n37653 ;
  assign n37676 = ~n37362 & n37653 ;
  assign n37677 = ~n37675 & ~n37676 ;
  assign n37678 = \core_c_psq_pcstk_cnts16x14_PCcell_reg[0][1]/P0001  & ~n37653 ;
  assign n37679 = ~n37292 & n37653 ;
  assign n37680 = ~n37678 & ~n37679 ;
  assign n37681 = \core_c_psq_pcstk_cnts16x14_PCcell_reg[0][13]/P0001  & ~n37653 ;
  assign n37682 = ~n37374 & n37653 ;
  assign n37683 = ~n37681 & ~n37682 ;
  assign n37684 = \core_c_psq_pcstk_cnts16x14_PCcell_reg[0][12]/P0001  & ~n37653 ;
  assign n37685 = ~n37383 & n37653 ;
  assign n37686 = ~n37684 & ~n37685 ;
  assign n37687 = \core_c_psq_pcstk_cnts16x14_PCcell_reg[0][11]/P0001  & ~n37653 ;
  assign n37688 = ~n37301 & n37653 ;
  assign n37689 = ~n37687 & ~n37688 ;
  assign n37690 = \core_c_psq_pcstk_cnts16x14_PCcell_reg[0][10]/P0001  & ~n37653 ;
  assign n37691 = ~n37310 & n37653 ;
  assign n37692 = ~n37690 & ~n37691 ;
  assign n37693 = ~n37318 & n37653 ;
  assign n37694 = \core_c_psq_pcstk_cnts16x14_PCcell_reg[0][0]/P0001  & ~n37653 ;
  assign n37695 = ~n37693 & ~n37694 ;
  assign n37696 = \core_c_psq_Iact_E_reg[3]/NET0131  & ~n19477 ;
  assign n37697 = n19482 & n33213 ;
  assign n37698 = n33215 & n37697 ;
  assign n37699 = n19477 & n37698 ;
  assign n37700 = ~n37696 & ~n37699 ;
  assign n37701 = \core_c_psq_pcstk_cnts16x14_PCcell_reg[2][6]/P0001  & ~n37249 ;
  assign n37702 = n37249 & ~n37350 ;
  assign n37703 = ~n37701 & ~n37702 ;
  assign n37704 = ~\sport1_regs_MWORDreg_DO_reg[0]/NET0131  & n23274 ;
  assign n37705 = \sport1_txctl_Wcnt_reg[0]/NET0131  & ~n23264 ;
  assign n37706 = ~n36390 & ~n37705 ;
  assign n37707 = ~n23274 & n37706 ;
  assign n37708 = ~n37704 & ~n37707 ;
  assign n37709 = ~\sport1_regs_MWORDreg_DO_reg[6]/NET0131  & n23274 ;
  assign n37710 = \sport1_txctl_Wcnt_reg[6]/NET0131  & ~n36395 ;
  assign n37711 = n36397 & ~n37710 ;
  assign n37712 = ~n37709 & ~n37711 ;
  assign n37713 = \sport1_txctl_Wcnt_reg[3]/NET0131  & ~n36392 ;
  assign n37714 = ~n36393 & ~n37713 ;
  assign n37715 = ~n23274 & n37714 ;
  assign n37716 = ~\sport1_regs_MWORDreg_DO_reg[3]/NET0131  & n23274 ;
  assign n37717 = ~n37715 & ~n37716 ;
  assign n37718 = \sport1_txctl_Wcnt_reg[2]/NET0131  & ~n36391 ;
  assign n37719 = ~n36392 & ~n37718 ;
  assign n37720 = ~n23274 & n37719 ;
  assign n37721 = ~\sport1_regs_MWORDreg_DO_reg[2]/NET0131  & n23274 ;
  assign n37722 = ~n37720 & ~n37721 ;
  assign n37723 = ~\sport0_regs_MWORDreg_DO_reg[6]/NET0131  & n23286 ;
  assign n37724 = \sport0_txctl_Wcnt_reg[6]/NET0131  & ~n36411 ;
  assign n37725 = n36413 & ~n37724 ;
  assign n37726 = ~n37723 & ~n37725 ;
  assign n37727 = \sport0_txctl_Wcnt_reg[3]/NET0131  & ~n36408 ;
  assign n37728 = ~n36409 & ~n37727 ;
  assign n37729 = ~n23286 & n37728 ;
  assign n37730 = ~\sport0_regs_MWORDreg_DO_reg[3]/NET0131  & n23286 ;
  assign n37731 = ~n37729 & ~n37730 ;
  assign n37732 = \sport0_txctl_Wcnt_reg[2]/NET0131  & ~n36407 ;
  assign n37733 = ~n36408 & ~n37732 ;
  assign n37734 = ~n23286 & n37733 ;
  assign n37735 = ~\sport0_regs_MWORDreg_DO_reg[2]/NET0131  & n23286 ;
  assign n37736 = ~n37734 & ~n37735 ;
  assign n37737 = ~\sport0_regs_MWORDreg_DO_reg[0]/NET0131  & n23286 ;
  assign n37738 = \sport0_txctl_Wcnt_reg[0]/NET0131  & ~n23276 ;
  assign n37739 = ~n36406 & ~n37738 ;
  assign n37740 = ~n23286 & n37739 ;
  assign n37741 = ~n37737 & ~n37740 ;
  assign n37742 = ~n20068 & ~n32454 ;
  assign n37743 = ~n32483 & n37742 ;
  assign n37744 = ~\idma_DOVL_reg[9]/NET0131  & ~n37742 ;
  assign n37745 = ~n37743 & ~n37744 ;
  assign n37746 = ~n32458 & n37742 ;
  assign n37747 = ~\idma_DOVL_reg[8]/NET0131  & ~n37742 ;
  assign n37748 = ~n37746 & ~n37747 ;
  assign n37749 = ~n32520 & n37742 ;
  assign n37750 = ~\idma_DOVL_reg[10]/NET0131  & ~n37742 ;
  assign n37751 = ~n37749 & ~n37750 ;
  assign n37752 = ~n32512 & n37742 ;
  assign n37753 = ~\idma_DOVL_reg[11]/NET0131  & ~n37742 ;
  assign n37754 = ~n37752 & ~n37753 ;
  assign n37755 = \core_c_psq_pcstk_cnts16x14_PCcell_reg[2][12]/P0001  & ~n37249 ;
  assign n37756 = n37249 & ~n37383 ;
  assign n37757 = ~n37755 & ~n37756 ;
  assign n37758 = \core_c_psq_pcstk_cnts16x14_PCcell_reg[2][13]/P0001  & ~n37249 ;
  assign n37759 = n37249 & ~n37374 ;
  assign n37760 = ~n37758 & ~n37759 ;
  assign n37761 = \core_c_psq_pcstk_cnts16x14_PCcell_reg[1][5]/P0001  & ~n37322 ;
  assign n37762 = ~n37265 & n37322 ;
  assign n37763 = ~n37761 & ~n37762 ;
  assign n37764 = \core_c_psq_pcstk_cnts16x14_PCcell_reg[2][2]/P0001  & ~n37249 ;
  assign n37765 = n37249 & ~n37362 ;
  assign n37766 = ~n37764 & ~n37765 ;
  assign n37767 = n4220 & n37248 ;
  assign n37768 = \core_c_psq_pcstk_cnts16x14_PCcell_reg[9][9]/P0001  & ~n37767 ;
  assign n37769 = ~n37329 & n37767 ;
  assign n37770 = ~n37768 & ~n37769 ;
  assign n37771 = \core_c_psq_pcstk_cnts16x14_PCcell_reg[9][8]/P0001  & ~n37767 ;
  assign n37772 = ~n37338 & n37767 ;
  assign n37773 = ~n37771 & ~n37772 ;
  assign n37774 = \core_c_psq_pcstk_cnts16x14_PCcell_reg[9][7]/P0001  & ~n37767 ;
  assign n37775 = ~n37256 & n37767 ;
  assign n37776 = ~n37774 & ~n37775 ;
  assign n37777 = \core_c_psq_pcstk_cnts16x14_PCcell_reg[9][6]/P0001  & ~n37767 ;
  assign n37778 = ~n37350 & n37767 ;
  assign n37779 = ~n37777 & ~n37778 ;
  assign n37780 = \core_c_psq_pcstk_cnts16x14_PCcell_reg[9][5]/P0001  & ~n37767 ;
  assign n37781 = ~n37265 & n37767 ;
  assign n37782 = ~n37780 & ~n37781 ;
  assign n37783 = \core_c_psq_pcstk_cnts16x14_PCcell_reg[9][4]/P0001  & ~n37767 ;
  assign n37784 = ~n37274 & n37767 ;
  assign n37785 = ~n37783 & ~n37784 ;
  assign n37786 = \core_c_psq_pcstk_cnts16x14_PCcell_reg[9][3]/P0001  & ~n37767 ;
  assign n37787 = ~n37283 & n37767 ;
  assign n37788 = ~n37786 & ~n37787 ;
  assign n37789 = \core_c_psq_pcstk_cnts16x14_PCcell_reg[9][2]/P0001  & ~n37767 ;
  assign n37790 = ~n37362 & n37767 ;
  assign n37791 = ~n37789 & ~n37790 ;
  assign n37792 = \core_c_psq_pcstk_cnts16x14_PCcell_reg[9][1]/P0001  & ~n37767 ;
  assign n37793 = ~n37292 & n37767 ;
  assign n37794 = ~n37792 & ~n37793 ;
  assign n37795 = \core_c_psq_pcstk_cnts16x14_PCcell_reg[9][13]/P0001  & ~n37767 ;
  assign n37796 = ~n37374 & n37767 ;
  assign n37797 = ~n37795 & ~n37796 ;
  assign n37798 = \core_c_psq_pcstk_cnts16x14_PCcell_reg[9][12]/P0001  & ~n37767 ;
  assign n37799 = ~n37383 & n37767 ;
  assign n37800 = ~n37798 & ~n37799 ;
  assign n37801 = \core_c_psq_pcstk_cnts16x14_PCcell_reg[9][11]/P0001  & ~n37767 ;
  assign n37802 = ~n37301 & n37767 ;
  assign n37803 = ~n37801 & ~n37802 ;
  assign n37804 = \core_c_psq_pcstk_cnts16x14_PCcell_reg[9][10]/P0001  & ~n37767 ;
  assign n37805 = ~n37310 & n37767 ;
  assign n37806 = ~n37804 & ~n37805 ;
  assign n37807 = ~n37318 & n37767 ;
  assign n37808 = \core_c_psq_pcstk_cnts16x14_PCcell_reg[9][0]/P0001  & ~n37767 ;
  assign n37809 = ~n37807 & ~n37808 ;
  assign n37810 = n4209 & n37248 ;
  assign n37811 = \core_c_psq_pcstk_cnts16x14_PCcell_reg[8][9]/P0001  & ~n37810 ;
  assign n37812 = ~n37329 & n37810 ;
  assign n37813 = ~n37811 & ~n37812 ;
  assign n37814 = \core_c_psq_pcstk_cnts16x14_PCcell_reg[8][8]/P0001  & ~n37810 ;
  assign n37815 = ~n37338 & n37810 ;
  assign n37816 = ~n37814 & ~n37815 ;
  assign n37817 = \core_c_psq_pcstk_cnts16x14_PCcell_reg[8][7]/P0001  & ~n37810 ;
  assign n37818 = ~n37256 & n37810 ;
  assign n37819 = ~n37817 & ~n37818 ;
  assign n37820 = \core_c_psq_pcstk_cnts16x14_PCcell_reg[8][6]/P0001  & ~n37810 ;
  assign n37821 = ~n37350 & n37810 ;
  assign n37822 = ~n37820 & ~n37821 ;
  assign n37823 = \core_c_psq_pcstk_cnts16x14_PCcell_reg[8][5]/P0001  & ~n37810 ;
  assign n37824 = ~n37265 & n37810 ;
  assign n37825 = ~n37823 & ~n37824 ;
  assign n37826 = \core_c_psq_pcstk_cnts16x14_PCcell_reg[8][4]/P0001  & ~n37810 ;
  assign n37827 = ~n37274 & n37810 ;
  assign n37828 = ~n37826 & ~n37827 ;
  assign n37829 = \core_c_psq_pcstk_cnts16x14_PCcell_reg[8][3]/P0001  & ~n37810 ;
  assign n37830 = ~n37283 & n37810 ;
  assign n37831 = ~n37829 & ~n37830 ;
  assign n37832 = \core_c_psq_pcstk_cnts16x14_PCcell_reg[8][2]/P0001  & ~n37810 ;
  assign n37833 = ~n37362 & n37810 ;
  assign n37834 = ~n37832 & ~n37833 ;
  assign n37835 = \core_c_psq_pcstk_cnts16x14_PCcell_reg[8][1]/P0001  & ~n37810 ;
  assign n37836 = ~n37292 & n37810 ;
  assign n37837 = ~n37835 & ~n37836 ;
  assign n37838 = \core_c_psq_pcstk_cnts16x14_PCcell_reg[8][13]/P0001  & ~n37810 ;
  assign n37839 = ~n37374 & n37810 ;
  assign n37840 = ~n37838 & ~n37839 ;
  assign n37841 = \core_c_psq_pcstk_cnts16x14_PCcell_reg[8][12]/P0001  & ~n37810 ;
  assign n37842 = ~n37383 & n37810 ;
  assign n37843 = ~n37841 & ~n37842 ;
  assign n37844 = \core_c_psq_pcstk_cnts16x14_PCcell_reg[8][11]/P0001  & ~n37810 ;
  assign n37845 = ~n37301 & n37810 ;
  assign n37846 = ~n37844 & ~n37845 ;
  assign n37847 = \core_c_psq_pcstk_cnts16x14_PCcell_reg[8][10]/P0001  & ~n37810 ;
  assign n37848 = ~n37310 & n37810 ;
  assign n37849 = ~n37847 & ~n37848 ;
  assign n37850 = ~n37318 & n37810 ;
  assign n37851 = \core_c_psq_pcstk_cnts16x14_PCcell_reg[8][0]/P0001  & ~n37810 ;
  assign n37852 = ~n37850 & ~n37851 ;
  assign n37853 = n4226 & n37248 ;
  assign n37854 = \core_c_psq_pcstk_cnts16x14_PCcell_reg[7][9]/P0001  & ~n37853 ;
  assign n37855 = ~n37329 & n37853 ;
  assign n37856 = ~n37854 & ~n37855 ;
  assign n37857 = \core_c_psq_pcstk_cnts16x14_PCcell_reg[7][8]/P0001  & ~n37853 ;
  assign n37858 = ~n37338 & n37853 ;
  assign n37859 = ~n37857 & ~n37858 ;
  assign n37860 = \core_c_psq_pcstk_cnts16x14_PCcell_reg[7][7]/P0001  & ~n37853 ;
  assign n37861 = ~n37256 & n37853 ;
  assign n37862 = ~n37860 & ~n37861 ;
  assign n37863 = \core_c_psq_pcstk_cnts16x14_PCcell_reg[7][6]/P0001  & ~n37853 ;
  assign n37864 = ~n37350 & n37853 ;
  assign n37865 = ~n37863 & ~n37864 ;
  assign n37866 = \core_c_psq_pcstk_cnts16x14_PCcell_reg[7][5]/P0001  & ~n37853 ;
  assign n37867 = ~n37265 & n37853 ;
  assign n37868 = ~n37866 & ~n37867 ;
  assign n37869 = \core_c_psq_pcstk_cnts16x14_PCcell_reg[7][4]/P0001  & ~n37853 ;
  assign n37870 = ~n37274 & n37853 ;
  assign n37871 = ~n37869 & ~n37870 ;
  assign n37872 = \core_c_psq_pcstk_cnts16x14_PCcell_reg[7][3]/P0001  & ~n37853 ;
  assign n37873 = ~n37283 & n37853 ;
  assign n37874 = ~n37872 & ~n37873 ;
  assign n37875 = \core_c_psq_pcstk_cnts16x14_PCcell_reg[7][2]/P0001  & ~n37853 ;
  assign n37876 = ~n37362 & n37853 ;
  assign n37877 = ~n37875 & ~n37876 ;
  assign n37878 = \core_c_psq_pcstk_cnts16x14_PCcell_reg[7][1]/P0001  & ~n37853 ;
  assign n37879 = ~n37292 & n37853 ;
  assign n37880 = ~n37878 & ~n37879 ;
  assign n37881 = \core_c_psq_pcstk_cnts16x14_PCcell_reg[7][13]/P0001  & ~n37853 ;
  assign n37882 = ~n37374 & n37853 ;
  assign n37883 = ~n37881 & ~n37882 ;
  assign n37884 = \core_c_psq_pcstk_cnts16x14_PCcell_reg[7][12]/P0001  & ~n37853 ;
  assign n37885 = ~n37383 & n37853 ;
  assign n37886 = ~n37884 & ~n37885 ;
  assign n37887 = \core_c_psq_pcstk_cnts16x14_PCcell_reg[7][11]/P0001  & ~n37853 ;
  assign n37888 = ~n37301 & n37853 ;
  assign n37889 = ~n37887 & ~n37888 ;
  assign n37890 = \core_c_psq_pcstk_cnts16x14_PCcell_reg[7][10]/P0001  & ~n37853 ;
  assign n37891 = ~n37310 & n37853 ;
  assign n37892 = ~n37890 & ~n37891 ;
  assign n37893 = ~n37318 & n37853 ;
  assign n37894 = \core_c_psq_pcstk_cnts16x14_PCcell_reg[7][0]/P0001  & ~n37853 ;
  assign n37895 = ~n37893 & ~n37894 ;
  assign n37896 = n4213 & n37248 ;
  assign n37897 = \core_c_psq_pcstk_cnts16x14_PCcell_reg[6][9]/P0001  & ~n37896 ;
  assign n37898 = ~n37329 & n37896 ;
  assign n37899 = ~n37897 & ~n37898 ;
  assign n37900 = \core_c_psq_pcstk_cnts16x14_PCcell_reg[6][8]/P0001  & ~n37896 ;
  assign n37901 = ~n37338 & n37896 ;
  assign n37902 = ~n37900 & ~n37901 ;
  assign n37903 = \core_c_psq_pcstk_cnts16x14_PCcell_reg[6][7]/P0001  & ~n37896 ;
  assign n37904 = ~n37256 & n37896 ;
  assign n37905 = ~n37903 & ~n37904 ;
  assign n37906 = \core_c_psq_pcstk_cnts16x14_PCcell_reg[6][6]/P0001  & ~n37896 ;
  assign n37907 = ~n37350 & n37896 ;
  assign n37908 = ~n37906 & ~n37907 ;
  assign n37909 = \core_c_psq_pcstk_cnts16x14_PCcell_reg[6][4]/P0001  & ~n37896 ;
  assign n37910 = ~n37274 & n37896 ;
  assign n37911 = ~n37909 & ~n37910 ;
  assign n37912 = \core_c_psq_pcstk_cnts16x14_PCcell_reg[6][3]/P0001  & ~n37896 ;
  assign n37913 = ~n37283 & n37896 ;
  assign n37914 = ~n37912 & ~n37913 ;
  assign n37915 = \core_c_psq_pcstk_cnts16x14_PCcell_reg[6][5]/P0001  & ~n37896 ;
  assign n37916 = ~n37265 & n37896 ;
  assign n37917 = ~n37915 & ~n37916 ;
  assign n37918 = \core_c_psq_pcstk_cnts16x14_PCcell_reg[6][2]/P0001  & ~n37896 ;
  assign n37919 = ~n37362 & n37896 ;
  assign n37920 = ~n37918 & ~n37919 ;
  assign n37921 = \core_c_psq_pcstk_cnts16x14_PCcell_reg[6][13]/P0001  & ~n37896 ;
  assign n37922 = ~n37374 & n37896 ;
  assign n37923 = ~n37921 & ~n37922 ;
  assign n37924 = \core_c_psq_pcstk_cnts16x14_PCcell_reg[6][1]/P0001  & ~n37896 ;
  assign n37925 = ~n37292 & n37896 ;
  assign n37926 = ~n37924 & ~n37925 ;
  assign n37927 = \core_c_psq_pcstk_cnts16x14_PCcell_reg[6][12]/P0001  & ~n37896 ;
  assign n37928 = ~n37383 & n37896 ;
  assign n37929 = ~n37927 & ~n37928 ;
  assign n37930 = \core_c_psq_pcstk_cnts16x14_PCcell_reg[6][11]/P0001  & ~n37896 ;
  assign n37931 = ~n37301 & n37896 ;
  assign n37932 = ~n37930 & ~n37931 ;
  assign n37933 = \core_c_psq_pcstk_cnts16x14_PCcell_reg[6][10]/P0001  & ~n37896 ;
  assign n37934 = ~n37310 & n37896 ;
  assign n37935 = ~n37933 & ~n37934 ;
  assign n37936 = ~n37318 & n37896 ;
  assign n37937 = \core_c_psq_pcstk_cnts16x14_PCcell_reg[6][0]/P0001  & ~n37896 ;
  assign n37938 = ~n37936 & ~n37937 ;
  assign n37939 = n4197 & n37248 ;
  assign n37940 = \core_c_psq_pcstk_cnts16x14_PCcell_reg[5][9]/P0001  & ~n37939 ;
  assign n37941 = ~n37329 & n37939 ;
  assign n37942 = ~n37940 & ~n37941 ;
  assign n37943 = \core_c_psq_pcstk_cnts16x14_PCcell_reg[5][8]/P0001  & ~n37939 ;
  assign n37944 = ~n37338 & n37939 ;
  assign n37945 = ~n37943 & ~n37944 ;
  assign n37946 = \core_c_psq_pcstk_cnts16x14_PCcell_reg[5][7]/P0001  & ~n37939 ;
  assign n37947 = ~n37256 & n37939 ;
  assign n37948 = ~n37946 & ~n37947 ;
  assign n37949 = \core_c_psq_pcstk_cnts16x14_PCcell_reg[5][6]/P0001  & ~n37939 ;
  assign n37950 = ~n37350 & n37939 ;
  assign n37951 = ~n37949 & ~n37950 ;
  assign n37952 = \core_c_psq_pcstk_cnts16x14_PCcell_reg[5][5]/P0001  & ~n37939 ;
  assign n37953 = ~n37265 & n37939 ;
  assign n37954 = ~n37952 & ~n37953 ;
  assign n37955 = \core_c_psq_pcstk_cnts16x14_PCcell_reg[5][4]/P0001  & ~n37939 ;
  assign n37956 = ~n37274 & n37939 ;
  assign n37957 = ~n37955 & ~n37956 ;
  assign n37958 = \core_c_psq_pcstk_cnts16x14_PCcell_reg[5][3]/P0001  & ~n37939 ;
  assign n37959 = ~n37283 & n37939 ;
  assign n37960 = ~n37958 & ~n37959 ;
  assign n37961 = \core_c_psq_pcstk_cnts16x14_PCcell_reg[5][2]/P0001  & ~n37939 ;
  assign n37962 = ~n37362 & n37939 ;
  assign n37963 = ~n37961 & ~n37962 ;
  assign n37964 = \core_c_psq_pcstk_cnts16x14_PCcell_reg[5][1]/P0001  & ~n37939 ;
  assign n37965 = ~n37292 & n37939 ;
  assign n37966 = ~n37964 & ~n37965 ;
  assign n37967 = \core_c_psq_pcstk_cnts16x14_PCcell_reg[5][13]/P0001  & ~n37939 ;
  assign n37968 = ~n37374 & n37939 ;
  assign n37969 = ~n37967 & ~n37968 ;
  assign n37970 = \core_c_psq_pcstk_cnts16x14_PCcell_reg[5][12]/P0001  & ~n37939 ;
  assign n37971 = ~n37383 & n37939 ;
  assign n37972 = ~n37970 & ~n37971 ;
  assign n37973 = \core_c_psq_pcstk_cnts16x14_PCcell_reg[5][11]/P0001  & ~n37939 ;
  assign n37974 = ~n37301 & n37939 ;
  assign n37975 = ~n37973 & ~n37974 ;
  assign n37976 = ~n37318 & n37939 ;
  assign n37977 = \core_c_psq_pcstk_cnts16x14_PCcell_reg[5][0]/P0001  & ~n37939 ;
  assign n37978 = ~n37976 & ~n37977 ;
  assign n37979 = \core_c_psq_pcstk_cnts16x14_PCcell_reg[5][10]/P0001  & ~n37939 ;
  assign n37980 = ~n37310 & n37939 ;
  assign n37981 = ~n37979 & ~n37980 ;
  assign n37982 = n4200 & n37248 ;
  assign n37983 = \core_c_psq_pcstk_cnts16x14_PCcell_reg[4][9]/P0001  & ~n37982 ;
  assign n37984 = ~n37329 & n37982 ;
  assign n37985 = ~n37983 & ~n37984 ;
  assign n37986 = \core_c_psq_pcstk_cnts16x14_PCcell_reg[4][8]/P0001  & ~n37982 ;
  assign n37987 = ~n37338 & n37982 ;
  assign n37988 = ~n37986 & ~n37987 ;
  assign n37989 = \core_c_psq_pcstk_cnts16x14_PCcell_reg[4][7]/P0001  & ~n37982 ;
  assign n37990 = ~n37256 & n37982 ;
  assign n37991 = ~n37989 & ~n37990 ;
  assign n37992 = \core_c_psq_pcstk_cnts16x14_PCcell_reg[4][6]/P0001  & ~n37982 ;
  assign n37993 = ~n37350 & n37982 ;
  assign n37994 = ~n37992 & ~n37993 ;
  assign n37995 = \core_c_psq_pcstk_cnts16x14_PCcell_reg[4][5]/P0001  & ~n37982 ;
  assign n37996 = ~n37265 & n37982 ;
  assign n37997 = ~n37995 & ~n37996 ;
  assign n37998 = \core_c_psq_pcstk_cnts16x14_PCcell_reg[4][4]/P0001  & ~n37982 ;
  assign n37999 = ~n37274 & n37982 ;
  assign n38000 = ~n37998 & ~n37999 ;
  assign n38001 = \core_c_psq_pcstk_cnts16x14_PCcell_reg[4][3]/P0001  & ~n37982 ;
  assign n38002 = ~n37283 & n37982 ;
  assign n38003 = ~n38001 & ~n38002 ;
  assign n38004 = \core_c_psq_pcstk_cnts16x14_PCcell_reg[4][2]/P0001  & ~n37982 ;
  assign n38005 = ~n37362 & n37982 ;
  assign n38006 = ~n38004 & ~n38005 ;
  assign n38007 = \core_c_psq_pcstk_cnts16x14_PCcell_reg[4][1]/P0001  & ~n37982 ;
  assign n38008 = ~n37292 & n37982 ;
  assign n38009 = ~n38007 & ~n38008 ;
  assign n38010 = \core_c_psq_pcstk_cnts16x14_PCcell_reg[4][13]/P0001  & ~n37982 ;
  assign n38011 = ~n37374 & n37982 ;
  assign n38012 = ~n38010 & ~n38011 ;
  assign n38013 = \core_c_psq_pcstk_cnts16x14_PCcell_reg[4][12]/P0001  & ~n37982 ;
  assign n38014 = ~n37383 & n37982 ;
  assign n38015 = ~n38013 & ~n38014 ;
  assign n38016 = \core_c_psq_pcstk_cnts16x14_PCcell_reg[4][11]/P0001  & ~n37982 ;
  assign n38017 = ~n37301 & n37982 ;
  assign n38018 = ~n38016 & ~n38017 ;
  assign n38019 = \core_c_psq_pcstk_cnts16x14_PCcell_reg[4][10]/P0001  & ~n37982 ;
  assign n38020 = ~n37310 & n37982 ;
  assign n38021 = ~n38019 & ~n38020 ;
  assign n38022 = ~n37318 & n37982 ;
  assign n38023 = \core_c_psq_pcstk_cnts16x14_PCcell_reg[4][0]/P0001  & ~n37982 ;
  assign n38024 = ~n38022 & ~n38023 ;
  assign n38025 = n4211 & n37248 ;
  assign n38026 = \core_c_psq_pcstk_cnts16x14_PCcell_reg[3][9]/P0001  & ~n38025 ;
  assign n38027 = ~n37329 & n38025 ;
  assign n38028 = ~n38026 & ~n38027 ;
  assign n38029 = \core_c_psq_pcstk_cnts16x14_PCcell_reg[3][8]/P0001  & ~n38025 ;
  assign n38030 = ~n37338 & n38025 ;
  assign n38031 = ~n38029 & ~n38030 ;
  assign n38032 = \core_c_psq_pcstk_cnts16x14_PCcell_reg[3][7]/P0001  & ~n38025 ;
  assign n38033 = ~n37256 & n38025 ;
  assign n38034 = ~n38032 & ~n38033 ;
  assign n38035 = \core_c_psq_pcstk_cnts16x14_PCcell_reg[1][4]/P0001  & ~n37322 ;
  assign n38036 = ~n37274 & n37322 ;
  assign n38037 = ~n38035 & ~n38036 ;
  assign n38038 = \core_c_psq_pcstk_cnts16x14_PCcell_reg[3][6]/P0001  & ~n38025 ;
  assign n38039 = ~n37350 & n38025 ;
  assign n38040 = ~n38038 & ~n38039 ;
  assign n38041 = \core_c_psq_pcstk_cnts16x14_PCcell_reg[3][5]/P0001  & ~n38025 ;
  assign n38042 = ~n37265 & n38025 ;
  assign n38043 = ~n38041 & ~n38042 ;
  assign n38044 = \core_c_psq_pcstk_cnts16x14_PCcell_reg[3][4]/P0001  & ~n38025 ;
  assign n38045 = ~n37274 & n38025 ;
  assign n38046 = ~n38044 & ~n38045 ;
  assign n38047 = \core_c_psq_pcstk_cnts16x14_PCcell_reg[3][3]/P0001  & ~n38025 ;
  assign n38048 = ~n37283 & n38025 ;
  assign n38049 = ~n38047 & ~n38048 ;
  assign n38050 = \core_c_psq_pcstk_cnts16x14_PCcell_reg[3][2]/P0001  & ~n38025 ;
  assign n38051 = ~n37362 & n38025 ;
  assign n38052 = ~n38050 & ~n38051 ;
  assign n38053 = \core_c_psq_pcstk_cnts16x14_PCcell_reg[3][1]/P0001  & ~n38025 ;
  assign n38054 = ~n37292 & n38025 ;
  assign n38055 = ~n38053 & ~n38054 ;
  assign n38056 = \core_c_psq_pcstk_cnts16x14_PCcell_reg[3][13]/P0001  & ~n38025 ;
  assign n38057 = ~n37374 & n38025 ;
  assign n38058 = ~n38056 & ~n38057 ;
  assign n38059 = \core_c_psq_pcstk_cnts16x14_PCcell_reg[3][12]/P0001  & ~n38025 ;
  assign n38060 = ~n37383 & n38025 ;
  assign n38061 = ~n38059 & ~n38060 ;
  assign n38062 = \core_c_psq_pcstk_cnts16x14_PCcell_reg[3][11]/P0001  & ~n38025 ;
  assign n38063 = ~n37301 & n38025 ;
  assign n38064 = ~n38062 & ~n38063 ;
  assign n38065 = \core_c_psq_pcstk_cnts16x14_PCcell_reg[3][10]/P0001  & ~n38025 ;
  assign n38066 = ~n37310 & n38025 ;
  assign n38067 = ~n38065 & ~n38066 ;
  assign n38068 = ~n37318 & n38025 ;
  assign n38069 = \core_c_psq_pcstk_cnts16x14_PCcell_reg[3][0]/P0001  & ~n38025 ;
  assign n38070 = ~n38068 & ~n38069 ;
  assign n38071 = \core_c_psq_pcstk_cnts16x14_PCcell_reg[2][9]/P0001  & ~n37249 ;
  assign n38072 = n37249 & ~n37329 ;
  assign n38073 = ~n38071 & ~n38072 ;
  assign n38074 = \core_c_psq_pcstk_cnts16x14_PCcell_reg[2][8]/P0001  & ~n37249 ;
  assign n38075 = n37249 & ~n37338 ;
  assign n38076 = ~n38074 & ~n38075 ;
  assign n38077 = ~n32541 & n37742 ;
  assign n38078 = ~\idma_DOVL_reg[7]/NET0131  & ~n37742 ;
  assign n38079 = ~n38077 & ~n38078 ;
  assign n38080 = ~n32557 & n37742 ;
  assign n38081 = ~\idma_DOVL_reg[6]/NET0131  & ~n37742 ;
  assign n38082 = ~n38080 & ~n38081 ;
  assign n38083 = ~n32549 & n37742 ;
  assign n38084 = ~\idma_DOVL_reg[5]/NET0131  & ~n37742 ;
  assign n38085 = ~n38083 & ~n38084 ;
  assign n38086 = ~n32573 & n37742 ;
  assign n38087 = ~\idma_DOVL_reg[3]/NET0131  & ~n37742 ;
  assign n38088 = ~n38086 & ~n38087 ;
  assign n38089 = ~n32565 & n37742 ;
  assign n38090 = ~\idma_DOVL_reg[4]/NET0131  & ~n37742 ;
  assign n38091 = ~n38089 & ~n38090 ;
  assign n38092 = ~n32581 & n37742 ;
  assign n38093 = ~\idma_DOVL_reg[2]/NET0131  & ~n37742 ;
  assign n38094 = ~n38092 & ~n38093 ;
  assign n38095 = ~n32677 & n37742 ;
  assign n38096 = ~\idma_DOVL_reg[1]/NET0131  & ~n37742 ;
  assign n38097 = ~n38095 & ~n38096 ;
  assign n38098 = ~n32589 & n37742 ;
  assign n38099 = ~\idma_DOVL_reg[0]/NET0131  & ~n37742 ;
  assign n38100 = ~n38098 & ~n38099 ;
  assign n38101 = \sport0_regs_SCTLreg_DO_reg[7]/NET0131  & n18233 ;
  assign n38102 = n11265 & n18237 ;
  assign n38103 = ~n38101 & ~n38102 ;
  assign n38104 = \sport0_regs_SCTLreg_DO_reg[6]/NET0131  & n18233 ;
  assign n38105 = n11525 & n18237 ;
  assign n38106 = ~n38104 & ~n38105 ;
  assign n38107 = \sport0_regs_SCTLreg_DO_reg[5]/NET0131  & n18233 ;
  assign n38108 = n10911 & n18237 ;
  assign n38109 = ~n38107 & ~n38108 ;
  assign n38110 = \sport0_regs_SCTLreg_DO_reg[15]/NET0131  & n18233 ;
  assign n38111 = n12743 & n18237 ;
  assign n38112 = ~n38110 & ~n38111 ;
  assign n38113 = \ISCLK0_pad  & n18233 ;
  assign n38114 = n12688 & n18237 ;
  assign n38115 = ~n38113 & ~n38114 ;
  assign n38116 = \sport0_txctl_Wcnt_reg[4]/NET0131  & ~n36409 ;
  assign n38117 = ~n36410 & ~n38116 ;
  assign n38118 = ~n23286 & n38117 ;
  assign n38119 = ~\sport0_regs_MWORDreg_DO_reg[4]/NET0131  & n23286 ;
  assign n38120 = ~n38118 & ~n38119 ;
  assign n38121 = \sport1_txctl_Wcnt_reg[4]/NET0131  & ~n36393 ;
  assign n38122 = ~n36394 & ~n38121 ;
  assign n38123 = ~n23274 & n38122 ;
  assign n38124 = ~\sport1_regs_MWORDreg_DO_reg[4]/NET0131  & n23274 ;
  assign n38125 = ~n38123 & ~n38124 ;
  assign n38126 = ~\bdma_BEAD_reg[2]/NET0131  & ~n20769 ;
  assign n38127 = ~n20765 & ~n33304 ;
  assign n38128 = ~n38126 & n38127 ;
  assign n38129 = n8715 & n20765 ;
  assign n38130 = ~n38128 & ~n38129 ;
  assign n38131 = \sport1_txctl_Wcnt_reg[1]/NET0131  & ~n36390 ;
  assign n38132 = ~n36391 & ~n38131 ;
  assign n38133 = ~n23274 & n38132 ;
  assign n38134 = ~\sport1_regs_MWORDreg_DO_reg[1]/NET0131  & n23274 ;
  assign n38135 = ~n38133 & ~n38134 ;
  assign n38136 = \sport0_txctl_Wcnt_reg[1]/NET0131  & ~n36406 ;
  assign n38137 = ~n36407 & ~n38136 ;
  assign n38138 = ~n23286 & n38137 ;
  assign n38139 = ~\sport0_regs_MWORDreg_DO_reg[1]/NET0131  & n23286 ;
  assign n38140 = ~n38138 & ~n38139 ;
  assign n38141 = ~\idma_RDcnt_reg[2]/NET0131  & ~n20828 ;
  assign n38142 = \idma_RDcnt_reg[2]/NET0131  & n20828 ;
  assign n38143 = ~n38141 & ~n38142 ;
  assign n38144 = ~n20824 & ~n38143 ;
  assign n38145 = ~\memc_usysr_DO_reg[6]/NET0131  & n20824 ;
  assign n38146 = ~n38144 & ~n38145 ;
  assign n38147 = \sport1_regs_SCTLreg_DO_reg[7]/NET0131  & n37215 ;
  assign n38148 = n11265 & n37218 ;
  assign n38149 = ~n38147 & ~n38148 ;
  assign n38150 = \sport1_regs_SCTLreg_DO_reg[6]/NET0131  & n37215 ;
  assign n38151 = n11525 & n37218 ;
  assign n38152 = ~n38150 & ~n38151 ;
  assign n38153 = \sport1_regs_SCTLreg_DO_reg[5]/NET0131  & n37215 ;
  assign n38154 = n10911 & n37218 ;
  assign n38155 = ~n38153 & ~n38154 ;
  assign n38156 = \sport1_regs_SCTLreg_DO_reg[4]/NET0131  & n37215 ;
  assign n38157 = n10069 & n37218 ;
  assign n38158 = ~n38156 & ~n38157 ;
  assign n38159 = \sport1_regs_SCTLreg_DO_reg[15]/NET0131  & n37215 ;
  assign n38160 = n12743 & ~n37217 ;
  assign n38161 = n36073 & n38160 ;
  assign n38162 = ~n38159 & ~n38161 ;
  assign n38163 = \ISCLK1_pad  & n37215 ;
  assign n38164 = n12688 & ~n37217 ;
  assign n38165 = n36073 & n38164 ;
  assign n38166 = ~n38163 & ~n38165 ;
  assign n38167 = \sport1_regs_SCTLreg_DO_reg[13]/NET0131  & n37215 ;
  assign n38168 = n7340 & ~n37217 ;
  assign n38169 = n36073 & n38168 ;
  assign n38170 = ~n38167 & ~n38169 ;
  assign n38171 = \sport1_regs_SCTLreg_DO_reg[12]/NET0131  & n37215 ;
  assign n38172 = n9178 & ~n37217 ;
  assign n38173 = n36073 & n38172 ;
  assign n38174 = ~n38171 & ~n38173 ;
  assign n38175 = ~n36075 & ~n36108 ;
  assign n38176 = \sport1_regs_FSDIVreg_DO_reg[9]/NET0131  & n38175 ;
  assign n38177 = n36108 & ~n37217 ;
  assign n38178 = n10289 & n38177 ;
  assign n38179 = ~n38176 & ~n38178 ;
  assign n38180 = \sport1_regs_FSDIVreg_DO_reg[8]/NET0131  & n38175 ;
  assign n38181 = n10638 & n38177 ;
  assign n38182 = ~n38180 & ~n38181 ;
  assign n38183 = \sport1_regs_FSDIVreg_DO_reg[15]/NET0131  & n38175 ;
  assign n38184 = n36108 & n38160 ;
  assign n38185 = ~n38183 & ~n38184 ;
  assign n38186 = \sport1_regs_FSDIVreg_DO_reg[14]/NET0131  & n38175 ;
  assign n38187 = n36108 & n38164 ;
  assign n38188 = ~n38186 & ~n38187 ;
  assign n38189 = \sport1_regs_FSDIVreg_DO_reg[13]/NET0131  & n38175 ;
  assign n38190 = n36108 & n38168 ;
  assign n38191 = ~n38189 & ~n38190 ;
  assign n38192 = \sport1_regs_FSDIVreg_DO_reg[12]/NET0131  & n38175 ;
  assign n38193 = n36108 & n38172 ;
  assign n38194 = ~n38192 & ~n38193 ;
  assign n38195 = \sport1_regs_FSDIVreg_DO_reg[10]/NET0131  & n38175 ;
  assign n38196 = n7859 & n38177 ;
  assign n38197 = ~n38195 & ~n38196 ;
  assign n38198 = \sport1_regs_FSDIVreg_DO_reg[11]/NET0131  & n38175 ;
  assign n38199 = n8460 & n38177 ;
  assign n38200 = ~n38198 & ~n38199 ;
  assign n38201 = n14699 & ~n18220 ;
  assign n38202 = \core_c_psq_ststk_sts7x23_STcell_reg[6][9]/P0001  & ~n38201 ;
  assign n38203 = \core_c_psq_MSTAT_reg_DO_reg[1]/NET0131  & n38201 ;
  assign n38204 = ~n38202 & ~n38203 ;
  assign n38205 = \core_c_psq_ststk_sts7x23_STcell_reg[6][8]/P0001  & ~n38201 ;
  assign n38206 = \core_c_psq_MSTAT_reg_DO_reg[0]/P0002  & n38201 ;
  assign n38207 = ~n38205 & ~n38206 ;
  assign n38208 = \core_c_psq_ststk_sts7x23_STcell_reg[6][7]/P0001  & ~n38201 ;
  assign n38209 = \core_eu_ec_cun_SS_reg/P0001  & n38201 ;
  assign n38210 = ~n38208 & ~n38209 ;
  assign n38211 = \core_c_psq_ststk_sts7x23_STcell_reg[6][6]/P0001  & ~n38201 ;
  assign n38212 = ~n4174 & n38201 ;
  assign n38213 = ~n38211 & ~n38212 ;
  assign n38214 = \core_c_psq_ststk_sts7x23_STcell_reg[6][5]/P0001  & ~n38201 ;
  assign n38215 = \core_eu_ec_cun_AQ_reg/P0001  & n38201 ;
  assign n38216 = ~n38214 & ~n38215 ;
  assign n38217 = \core_c_psq_ststk_sts7x23_STcell_reg[6][4]/P0001  & ~n38201 ;
  assign n38218 = \core_eu_ec_cun_AS_reg/P0001  & n38201 ;
  assign n38219 = ~n38217 & ~n38218 ;
  assign n38220 = \core_c_psq_ststk_sts7x23_STcell_reg[6][3]/P0001  & ~n38201 ;
  assign n38221 = \core_eu_ec_cun_AC_reg/P0001  & n38201 ;
  assign n38222 = ~n38220 & ~n38221 ;
  assign n38223 = \core_c_psq_ststk_sts7x23_STcell_reg[6][2]/P0001  & ~n38201 ;
  assign n38224 = \core_eu_ec_cun_AV_reg/P0001  & n38201 ;
  assign n38225 = ~n38223 & ~n38224 ;
  assign n38226 = \core_c_psq_ststk_sts7x23_STcell_reg[6][24]/P0001  & ~n38201 ;
  assign n38227 = \core_c_psq_IMASK_reg[9]/NET0131  & n38201 ;
  assign n38228 = ~n38226 & ~n38227 ;
  assign n38229 = \core_c_psq_ststk_sts7x23_STcell_reg[6][23]/P0001  & ~n38201 ;
  assign n38230 = \core_c_psq_IMASK_reg[8]/NET0131  & n38201 ;
  assign n38231 = ~n38229 & ~n38230 ;
  assign n38232 = \core_c_psq_ststk_sts7x23_STcell_reg[6][22]/P0001  & ~n38201 ;
  assign n38233 = \core_c_psq_IMASK_reg[7]/NET0131  & n38201 ;
  assign n38234 = ~n38232 & ~n38233 ;
  assign n38235 = \core_c_psq_ststk_sts7x23_STcell_reg[6][21]/P0001  & ~n38201 ;
  assign n38236 = \core_c_psq_IMASK_reg[6]/NET0131  & n38201 ;
  assign n38237 = ~n38235 & ~n38236 ;
  assign n38238 = \core_c_psq_ststk_sts7x23_STcell_reg[6][20]/P0001  & ~n38201 ;
  assign n38239 = \core_c_psq_IMASK_reg[5]/NET0131  & n38201 ;
  assign n38240 = ~n38238 & ~n38239 ;
  assign n38241 = \core_c_psq_ststk_sts7x23_STcell_reg[6][1]/P0001  & ~n38201 ;
  assign n38242 = \core_eu_ec_cun_AN_reg/P0001  & n38201 ;
  assign n38243 = ~n38241 & ~n38242 ;
  assign n38244 = \core_c_psq_ststk_sts7x23_STcell_reg[6][19]/P0001  & ~n38201 ;
  assign n38245 = \core_c_psq_IMASK_reg[4]/NET0131  & n38201 ;
  assign n38246 = ~n38244 & ~n38245 ;
  assign n38247 = \core_c_psq_ststk_sts7x23_STcell_reg[6][18]/P0001  & ~n38201 ;
  assign n38248 = \core_c_psq_IMASK_reg[3]/NET0131  & n38201 ;
  assign n38249 = ~n38247 & ~n38248 ;
  assign n38250 = \core_c_psq_ststk_sts7x23_STcell_reg[6][17]/P0001  & ~n38201 ;
  assign n38251 = \core_c_psq_IMASK_reg[2]/NET0131  & n38201 ;
  assign n38252 = ~n38250 & ~n38251 ;
  assign n38253 = \core_c_psq_ststk_sts7x23_STcell_reg[6][16]/P0001  & ~n38201 ;
  assign n38254 = \core_c_psq_IMASK_reg[1]/NET0131  & n38201 ;
  assign n38255 = ~n38253 & ~n38254 ;
  assign n38256 = \core_c_psq_ststk_sts7x23_STcell_reg[6][15]/P0001  & ~n38201 ;
  assign n38257 = \core_c_psq_IMASK_reg[0]/NET0131  & n38201 ;
  assign n38258 = ~n38256 & ~n38257 ;
  assign n38259 = \core_c_psq_ststk_sts7x23_STcell_reg[6][14]/P0001  & ~n38201 ;
  assign n38260 = \core_c_psq_MSTAT_reg_DO_reg[6]/NET0131  & n38201 ;
  assign n38261 = ~n38259 & ~n38260 ;
  assign n38262 = \core_c_psq_ststk_sts7x23_STcell_reg[6][13]/P0001  & ~n38201 ;
  assign n38263 = \core_c_psq_MSTAT_reg_DO_reg[5]/NET0131  & n38201 ;
  assign n38264 = ~n38262 & ~n38263 ;
  assign n38267 = ~\sport0_rxctl_RX_reg[7]/P0001  & ~n31030 ;
  assign n38269 = n31042 & ~n38267 ;
  assign n38268 = ~n31042 & n38267 ;
  assign n38270 = n20875 & ~n38268 ;
  assign n38271 = ~n38269 & n38270 ;
  assign n38272 = ~\sport0_rxctl_ldRX_cmp_reg/P0001  & n11525 ;
  assign n38266 = \sport0_rxctl_RX_reg[6]/P0001  & n20873 ;
  assign n38273 = ~n20868 & ~n38266 ;
  assign n38274 = ~n38272 & n38273 ;
  assign n38275 = ~n38271 & n38274 ;
  assign n38265 = ~\sport0_rxctl_RXSHT_reg[6]/P0001  & n20868 ;
  assign n38276 = ~n20871 & ~n38265 ;
  assign n38277 = ~n38275 & n38276 ;
  assign n38278 = \sport0_rxctl_RX_reg[6]/P0001  & n20871 ;
  assign n38279 = ~n38277 & ~n38278 ;
  assign n38280 = \core_c_psq_ststk_sts7x23_STcell_reg[6][12]/P0001  & ~n38201 ;
  assign n38281 = \core_c_psq_MSTAT_reg_DO_reg[4]/NET0131  & n38201 ;
  assign n38282 = ~n38280 & ~n38281 ;
  assign n38283 = \core_c_psq_ststk_sts7x23_STcell_reg[6][11]/P0001  & ~n38201 ;
  assign n38284 = \core_c_psq_MSTAT_reg_DO_reg[3]/NET0131  & n38201 ;
  assign n38285 = ~n38283 & ~n38284 ;
  assign n38286 = \core_c_psq_ststk_sts7x23_STcell_reg[6][10]/P0001  & ~n38201 ;
  assign n38287 = \core_c_psq_MSTAT_reg_DO_reg[2]/NET0131  & n38201 ;
  assign n38288 = ~n38286 & ~n38287 ;
  assign n38289 = \core_c_psq_ststk_sts7x23_STcell_reg[6][0]/P0001  & ~n38201 ;
  assign n38290 = \core_eu_ec_cun_AZ_reg/P0001  & n38201 ;
  assign n38291 = ~n38289 & ~n38290 ;
  assign n38292 = n14706 & ~n18220 ;
  assign n38293 = \core_c_psq_ststk_sts7x23_STcell_reg[5][9]/P0001  & ~n38292 ;
  assign n38294 = \core_c_psq_MSTAT_reg_DO_reg[1]/NET0131  & n38292 ;
  assign n38295 = ~n38293 & ~n38294 ;
  assign n38296 = \core_c_psq_ststk_sts7x23_STcell_reg[5][8]/P0001  & ~n38292 ;
  assign n38297 = \core_c_psq_MSTAT_reg_DO_reg[0]/P0002  & n38292 ;
  assign n38298 = ~n38296 & ~n38297 ;
  assign n38299 = \core_c_psq_ststk_sts7x23_STcell_reg[5][7]/P0001  & ~n38292 ;
  assign n38300 = \core_eu_ec_cun_SS_reg/P0001  & n38292 ;
  assign n38301 = ~n38299 & ~n38300 ;
  assign n38302 = \core_c_psq_ststk_sts7x23_STcell_reg[5][6]/P0001  & ~n38292 ;
  assign n38303 = ~n4174 & n38292 ;
  assign n38304 = ~n38302 & ~n38303 ;
  assign n38305 = \core_c_psq_ststk_sts7x23_STcell_reg[5][5]/P0001  & ~n38292 ;
  assign n38306 = \core_eu_ec_cun_AQ_reg/P0001  & n38292 ;
  assign n38307 = ~n38305 & ~n38306 ;
  assign n38308 = \core_c_psq_ststk_sts7x23_STcell_reg[5][4]/P0001  & ~n38292 ;
  assign n38309 = \core_eu_ec_cun_AS_reg/P0001  & n38292 ;
  assign n38310 = ~n38308 & ~n38309 ;
  assign n38311 = \core_c_psq_ststk_sts7x23_STcell_reg[5][3]/P0001  & ~n38292 ;
  assign n38312 = \core_eu_ec_cun_AC_reg/P0001  & n38292 ;
  assign n38313 = ~n38311 & ~n38312 ;
  assign n38314 = \core_c_psq_ststk_sts7x23_STcell_reg[5][2]/P0001  & ~n38292 ;
  assign n38315 = \core_eu_ec_cun_AV_reg/P0001  & n38292 ;
  assign n38316 = ~n38314 & ~n38315 ;
  assign n38317 = \core_c_psq_ststk_sts7x23_STcell_reg[5][24]/P0001  & ~n38292 ;
  assign n38318 = \core_c_psq_IMASK_reg[9]/NET0131  & n38292 ;
  assign n38319 = ~n38317 & ~n38318 ;
  assign n38320 = \core_c_psq_ststk_sts7x23_STcell_reg[5][23]/P0001  & ~n38292 ;
  assign n38321 = \core_c_psq_IMASK_reg[8]/NET0131  & n38292 ;
  assign n38322 = ~n38320 & ~n38321 ;
  assign n38323 = \core_c_psq_ststk_sts7x23_STcell_reg[5][22]/P0001  & ~n38292 ;
  assign n38324 = \core_c_psq_IMASK_reg[7]/NET0131  & n38292 ;
  assign n38325 = ~n38323 & ~n38324 ;
  assign n38326 = \core_c_psq_ststk_sts7x23_STcell_reg[5][21]/P0001  & ~n38292 ;
  assign n38327 = \core_c_psq_IMASK_reg[6]/NET0131  & n38292 ;
  assign n38328 = ~n38326 & ~n38327 ;
  assign n38329 = \core_c_psq_ststk_sts7x23_STcell_reg[5][20]/P0001  & ~n38292 ;
  assign n38330 = \core_c_psq_IMASK_reg[5]/NET0131  & n38292 ;
  assign n38331 = ~n38329 & ~n38330 ;
  assign n38332 = \core_c_psq_ststk_sts7x23_STcell_reg[5][1]/P0001  & ~n38292 ;
  assign n38333 = \core_eu_ec_cun_AN_reg/P0001  & n38292 ;
  assign n38334 = ~n38332 & ~n38333 ;
  assign n38335 = \core_c_psq_ststk_sts7x23_STcell_reg[5][19]/P0001  & ~n38292 ;
  assign n38336 = \core_c_psq_IMASK_reg[4]/NET0131  & n38292 ;
  assign n38337 = ~n38335 & ~n38336 ;
  assign n38338 = \core_c_psq_ststk_sts7x23_STcell_reg[5][18]/P0001  & ~n38292 ;
  assign n38339 = \core_c_psq_IMASK_reg[3]/NET0131  & n38292 ;
  assign n38340 = ~n38338 & ~n38339 ;
  assign n38341 = \core_c_psq_ststk_sts7x23_STcell_reg[5][17]/P0001  & ~n38292 ;
  assign n38342 = \core_c_psq_IMASK_reg[2]/NET0131  & n38292 ;
  assign n38343 = ~n38341 & ~n38342 ;
  assign n38344 = \core_c_psq_ststk_sts7x23_STcell_reg[5][16]/P0001  & ~n38292 ;
  assign n38345 = \core_c_psq_IMASK_reg[1]/NET0131  & n38292 ;
  assign n38346 = ~n38344 & ~n38345 ;
  assign n38347 = \core_c_psq_ststk_sts7x23_STcell_reg[5][15]/P0001  & ~n38292 ;
  assign n38348 = \core_c_psq_IMASK_reg[0]/NET0131  & n38292 ;
  assign n38349 = ~n38347 & ~n38348 ;
  assign n38350 = \core_c_psq_ststk_sts7x23_STcell_reg[5][14]/P0001  & ~n38292 ;
  assign n38351 = \core_c_psq_MSTAT_reg_DO_reg[6]/NET0131  & n38292 ;
  assign n38352 = ~n38350 & ~n38351 ;
  assign n38353 = \core_c_psq_ststk_sts7x23_STcell_reg[5][13]/P0001  & ~n38292 ;
  assign n38354 = \core_c_psq_MSTAT_reg_DO_reg[5]/NET0131  & n38292 ;
  assign n38355 = ~n38353 & ~n38354 ;
  assign n38356 = \core_c_psq_ststk_sts7x23_STcell_reg[5][12]/P0001  & ~n38292 ;
  assign n38357 = \core_c_psq_MSTAT_reg_DO_reg[4]/NET0131  & n38292 ;
  assign n38358 = ~n38356 & ~n38357 ;
  assign n38359 = \core_c_psq_ststk_sts7x23_STcell_reg[5][11]/P0001  & ~n38292 ;
  assign n38360 = \core_c_psq_MSTAT_reg_DO_reg[3]/NET0131  & n38292 ;
  assign n38361 = ~n38359 & ~n38360 ;
  assign n38362 = \core_c_psq_ststk_sts7x23_STcell_reg[5][10]/P0001  & ~n38292 ;
  assign n38363 = \core_c_psq_MSTAT_reg_DO_reg[2]/NET0131  & n38292 ;
  assign n38364 = ~n38362 & ~n38363 ;
  assign n38365 = \core_c_psq_ststk_sts7x23_STcell_reg[5][0]/P0001  & ~n38292 ;
  assign n38366 = \core_eu_ec_cun_AZ_reg/P0001  & n38292 ;
  assign n38367 = ~n38365 & ~n38366 ;
  assign n38368 = ~\core_c_psq_ststk_ptr_reg[2]/NET0131  & n18679 ;
  assign n38369 = \core_c_psq_ststk_sts7x23_STcell_reg[4][9]/P0001  & ~n38368 ;
  assign n38370 = \core_c_psq_MSTAT_reg_DO_reg[1]/NET0131  & n38368 ;
  assign n38371 = ~n38369 & ~n38370 ;
  assign n38372 = \core_c_psq_ststk_sts7x23_STcell_reg[4][8]/P0001  & ~n38368 ;
  assign n38373 = \core_c_psq_MSTAT_reg_DO_reg[0]/P0002  & n38368 ;
  assign n38374 = ~n38372 & ~n38373 ;
  assign n38375 = \core_c_psq_ststk_sts7x23_STcell_reg[4][7]/P0001  & ~n38368 ;
  assign n38376 = \core_eu_ec_cun_SS_reg/P0001  & n38368 ;
  assign n38377 = ~n38375 & ~n38376 ;
  assign n38378 = \core_c_psq_ststk_sts7x23_STcell_reg[4][6]/P0001  & ~n38368 ;
  assign n38379 = ~n4174 & n38368 ;
  assign n38380 = ~n38378 & ~n38379 ;
  assign n38381 = \core_c_psq_ststk_sts7x23_STcell_reg[4][5]/P0001  & ~n38368 ;
  assign n38382 = \core_eu_ec_cun_AQ_reg/P0001  & n38368 ;
  assign n38383 = ~n38381 & ~n38382 ;
  assign n38384 = \core_c_psq_ststk_sts7x23_STcell_reg[4][4]/P0001  & ~n38368 ;
  assign n38385 = \core_eu_ec_cun_AS_reg/P0001  & n38368 ;
  assign n38386 = ~n38384 & ~n38385 ;
  assign n38387 = \core_c_psq_ststk_sts7x23_STcell_reg[4][3]/P0001  & ~n38368 ;
  assign n38388 = \core_eu_ec_cun_AC_reg/P0001  & n38368 ;
  assign n38389 = ~n38387 & ~n38388 ;
  assign n38390 = \core_c_psq_ststk_sts7x23_STcell_reg[4][2]/P0001  & ~n38368 ;
  assign n38391 = \core_eu_ec_cun_AV_reg/P0001  & n38368 ;
  assign n38392 = ~n38390 & ~n38391 ;
  assign n38393 = \core_c_psq_ststk_sts7x23_STcell_reg[4][24]/P0001  & ~n38368 ;
  assign n38394 = \core_c_psq_IMASK_reg[9]/NET0131  & n38368 ;
  assign n38395 = ~n38393 & ~n38394 ;
  assign n38396 = \core_c_psq_ststk_sts7x23_STcell_reg[4][23]/P0001  & ~n38368 ;
  assign n38397 = \core_c_psq_IMASK_reg[8]/NET0131  & n38368 ;
  assign n38398 = ~n38396 & ~n38397 ;
  assign n38399 = \core_c_psq_ststk_sts7x23_STcell_reg[4][22]/P0001  & ~n38368 ;
  assign n38400 = \core_c_psq_IMASK_reg[7]/NET0131  & n38368 ;
  assign n38401 = ~n38399 & ~n38400 ;
  assign n38402 = \core_c_psq_ststk_sts7x23_STcell_reg[4][21]/P0001  & ~n38368 ;
  assign n38403 = \core_c_psq_IMASK_reg[6]/NET0131  & n38368 ;
  assign n38404 = ~n38402 & ~n38403 ;
  assign n38405 = \core_c_psq_ststk_sts7x23_STcell_reg[4][20]/P0001  & ~n38368 ;
  assign n38406 = \core_c_psq_IMASK_reg[5]/NET0131  & n38368 ;
  assign n38407 = ~n38405 & ~n38406 ;
  assign n38408 = \core_c_psq_ststk_sts7x23_STcell_reg[4][1]/P0001  & ~n38368 ;
  assign n38409 = \core_eu_ec_cun_AN_reg/P0001  & n38368 ;
  assign n38410 = ~n38408 & ~n38409 ;
  assign n38411 = \core_c_psq_ststk_sts7x23_STcell_reg[4][19]/P0001  & ~n38368 ;
  assign n38412 = \core_c_psq_IMASK_reg[4]/NET0131  & n38368 ;
  assign n38413 = ~n38411 & ~n38412 ;
  assign n38414 = \core_c_psq_ststk_sts7x23_STcell_reg[4][18]/P0001  & ~n38368 ;
  assign n38415 = \core_c_psq_IMASK_reg[3]/NET0131  & n38368 ;
  assign n38416 = ~n38414 & ~n38415 ;
  assign n38417 = \core_c_psq_ststk_sts7x23_STcell_reg[4][17]/P0001  & ~n38368 ;
  assign n38418 = \core_c_psq_IMASK_reg[2]/NET0131  & n38368 ;
  assign n38419 = ~n38417 & ~n38418 ;
  assign n38420 = \core_c_psq_ststk_sts7x23_STcell_reg[4][16]/P0001  & ~n38368 ;
  assign n38421 = \core_c_psq_IMASK_reg[1]/NET0131  & n38368 ;
  assign n38422 = ~n38420 & ~n38421 ;
  assign n38423 = \core_c_psq_ststk_sts7x23_STcell_reg[4][15]/P0001  & ~n38368 ;
  assign n38424 = \core_c_psq_IMASK_reg[0]/NET0131  & n38368 ;
  assign n38425 = ~n38423 & ~n38424 ;
  assign n38426 = \core_c_psq_ststk_sts7x23_STcell_reg[4][14]/P0001  & ~n38368 ;
  assign n38427 = \core_c_psq_MSTAT_reg_DO_reg[6]/NET0131  & n38368 ;
  assign n38428 = ~n38426 & ~n38427 ;
  assign n38429 = \core_c_psq_ststk_sts7x23_STcell_reg[4][13]/P0001  & ~n38368 ;
  assign n38430 = \core_c_psq_MSTAT_reg_DO_reg[5]/NET0131  & n38368 ;
  assign n38431 = ~n38429 & ~n38430 ;
  assign n38432 = \core_c_psq_ststk_sts7x23_STcell_reg[4][12]/P0001  & ~n38368 ;
  assign n38433 = \core_c_psq_MSTAT_reg_DO_reg[4]/NET0131  & n38368 ;
  assign n38434 = ~n38432 & ~n38433 ;
  assign n38435 = \core_c_psq_ststk_sts7x23_STcell_reg[4][11]/P0001  & ~n38368 ;
  assign n38436 = \core_c_psq_MSTAT_reg_DO_reg[3]/NET0131  & n38368 ;
  assign n38437 = ~n38435 & ~n38436 ;
  assign n38438 = \core_c_psq_ststk_sts7x23_STcell_reg[4][10]/P0001  & ~n38368 ;
  assign n38439 = \core_c_psq_MSTAT_reg_DO_reg[2]/NET0131  & n38368 ;
  assign n38440 = ~n38438 & ~n38439 ;
  assign n38441 = \core_c_psq_ststk_sts7x23_STcell_reg[4][0]/P0001  & ~n38368 ;
  assign n38442 = \core_eu_ec_cun_AZ_reg/P0001  & n38368 ;
  assign n38443 = ~n38441 & ~n38442 ;
  assign n38444 = \core_c_psq_ststk_sts7x23_STcell_reg[3][9]/P0001  & ~n18221 ;
  assign n38445 = \core_c_psq_MSTAT_reg_DO_reg[1]/NET0131  & n18221 ;
  assign n38446 = ~n38444 & ~n38445 ;
  assign n38447 = \core_c_psq_ststk_sts7x23_STcell_reg[3][8]/P0001  & ~n18221 ;
  assign n38448 = \core_c_psq_MSTAT_reg_DO_reg[0]/P0002  & n18221 ;
  assign n38449 = ~n38447 & ~n38448 ;
  assign n38450 = \core_c_psq_ststk_sts7x23_STcell_reg[3][7]/P0001  & ~n18221 ;
  assign n38451 = \core_eu_ec_cun_SS_reg/P0001  & n18221 ;
  assign n38452 = ~n38450 & ~n38451 ;
  assign n38453 = \core_c_psq_ststk_sts7x23_STcell_reg[3][6]/P0001  & ~n18221 ;
  assign n38454 = ~n4174 & n18221 ;
  assign n38455 = ~n38453 & ~n38454 ;
  assign n38456 = \core_c_psq_ststk_sts7x23_STcell_reg[3][5]/P0001  & ~n18221 ;
  assign n38457 = \core_eu_ec_cun_AQ_reg/P0001  & n18221 ;
  assign n38458 = ~n38456 & ~n38457 ;
  assign n38459 = \core_c_psq_ststk_sts7x23_STcell_reg[3][4]/P0001  & ~n18221 ;
  assign n38460 = \core_eu_ec_cun_AS_reg/P0001  & n18221 ;
  assign n38461 = ~n38459 & ~n38460 ;
  assign n38462 = \core_c_psq_ststk_sts7x23_STcell_reg[3][3]/P0001  & ~n18221 ;
  assign n38463 = \core_eu_ec_cun_AC_reg/P0001  & n18221 ;
  assign n38464 = ~n38462 & ~n38463 ;
  assign n38465 = \core_c_psq_ststk_sts7x23_STcell_reg[3][2]/P0001  & ~n18221 ;
  assign n38466 = \core_eu_ec_cun_AV_reg/P0001  & n18221 ;
  assign n38467 = ~n38465 & ~n38466 ;
  assign n38468 = \core_c_psq_ststk_sts7x23_STcell_reg[3][24]/P0001  & ~n18221 ;
  assign n38469 = \core_c_psq_IMASK_reg[9]/NET0131  & n18221 ;
  assign n38470 = ~n38468 & ~n38469 ;
  assign n38471 = \core_c_psq_ststk_sts7x23_STcell_reg[3][23]/P0001  & ~n18221 ;
  assign n38472 = \core_c_psq_IMASK_reg[8]/NET0131  & n18221 ;
  assign n38473 = ~n38471 & ~n38472 ;
  assign n38474 = \core_c_psq_ststk_sts7x23_STcell_reg[3][22]/P0001  & ~n18221 ;
  assign n38475 = \core_c_psq_IMASK_reg[7]/NET0131  & n18221 ;
  assign n38476 = ~n38474 & ~n38475 ;
  assign n38477 = \core_c_psq_ststk_sts7x23_STcell_reg[3][21]/P0001  & ~n18221 ;
  assign n38478 = \core_c_psq_IMASK_reg[6]/NET0131  & n18221 ;
  assign n38479 = ~n38477 & ~n38478 ;
  assign n38480 = \core_c_psq_ststk_sts7x23_STcell_reg[3][20]/P0001  & ~n18221 ;
  assign n38481 = \core_c_psq_IMASK_reg[5]/NET0131  & n18221 ;
  assign n38482 = ~n38480 & ~n38481 ;
  assign n38483 = \core_c_psq_ststk_sts7x23_STcell_reg[3][1]/P0001  & ~n18221 ;
  assign n38484 = \core_eu_ec_cun_AN_reg/P0001  & n18221 ;
  assign n38485 = ~n38483 & ~n38484 ;
  assign n38486 = \core_c_psq_ststk_sts7x23_STcell_reg[3][19]/P0001  & ~n18221 ;
  assign n38487 = \core_c_psq_IMASK_reg[4]/NET0131  & n18221 ;
  assign n38488 = ~n38486 & ~n38487 ;
  assign n38489 = ~n18213 & n18717 ;
  assign n38490 = ~\core_eu_es_sht_es_reg_sr1swe_DO_reg[13]/P0001  & ~n18717 ;
  assign n38491 = ~n38489 & ~n38490 ;
  assign n38492 = \core_c_psq_ststk_sts7x23_STcell_reg[3][18]/P0001  & ~n18221 ;
  assign n38493 = \core_c_psq_IMASK_reg[3]/NET0131  & n18221 ;
  assign n38494 = ~n38492 & ~n38493 ;
  assign n38495 = \core_c_psq_ststk_sts7x23_STcell_reg[3][17]/P0001  & ~n18221 ;
  assign n38496 = \core_c_psq_IMASK_reg[2]/NET0131  & n18221 ;
  assign n38497 = ~n38495 & ~n38496 ;
  assign n38498 = \sport0_regs_SCTLreg_DO_reg[13]/NET0131  & n18233 ;
  assign n38499 = n7340 & n18237 ;
  assign n38500 = ~n38498 & ~n38499 ;
  assign n38501 = \core_c_psq_ststk_sts7x23_STcell_reg[3][16]/P0001  & ~n18221 ;
  assign n38502 = \core_c_psq_IMASK_reg[1]/NET0131  & n18221 ;
  assign n38503 = ~n38501 & ~n38502 ;
  assign n38504 = \core_c_psq_ststk_sts7x23_STcell_reg[3][15]/P0001  & ~n18221 ;
  assign n38505 = \core_c_psq_IMASK_reg[0]/NET0131  & n18221 ;
  assign n38506 = ~n38504 & ~n38505 ;
  assign n38507 = \core_c_psq_ststk_sts7x23_STcell_reg[3][14]/P0001  & ~n18221 ;
  assign n38508 = \core_c_psq_MSTAT_reg_DO_reg[6]/NET0131  & n18221 ;
  assign n38509 = ~n38507 & ~n38508 ;
  assign n38510 = \core_c_psq_ststk_sts7x23_STcell_reg[3][13]/P0001  & ~n18221 ;
  assign n38511 = \core_c_psq_MSTAT_reg_DO_reg[5]/NET0131  & n18221 ;
  assign n38512 = ~n38510 & ~n38511 ;
  assign n38513 = \core_c_psq_ststk_sts7x23_STcell_reg[3][12]/P0001  & ~n18221 ;
  assign n38514 = \core_c_psq_MSTAT_reg_DO_reg[4]/NET0131  & n18221 ;
  assign n38515 = ~n38513 & ~n38514 ;
  assign n38516 = \core_c_psq_ststk_sts7x23_STcell_reg[3][11]/P0001  & ~n18221 ;
  assign n38517 = \core_c_psq_MSTAT_reg_DO_reg[3]/NET0131  & n18221 ;
  assign n38518 = ~n38516 & ~n38517 ;
  assign n38519 = \core_c_psq_ststk_sts7x23_STcell_reg[3][10]/P0001  & ~n18221 ;
  assign n38520 = \core_c_psq_MSTAT_reg_DO_reg[2]/NET0131  & n18221 ;
  assign n38521 = ~n38519 & ~n38520 ;
  assign n38522 = ~n26090 & ~n34434 ;
  assign n38523 = \T_TMODE[1]_pad  & \core_c_dec_PPclr_reg/P0001  ;
  assign n38524 = ~n32093 & ~n38523 ;
  assign n38525 = \T_PIOin[0]_pad  & ~n25656 ;
  assign n38526 = \pio_PIO_IN_P_reg[0]/P0001  & n25656 ;
  assign n38527 = ~n38525 & ~n38526 ;
  assign n38528 = \T_PIOin[10]_pad  & ~n25661 ;
  assign n38529 = \pio_PIO_IN_P_reg[10]/P0001  & n25661 ;
  assign n38530 = ~n38528 & ~n38529 ;
  assign n38531 = \T_PIOin[11]_pad  & ~n25661 ;
  assign n38532 = \pio_PIO_IN_P_reg[11]/P0001  & n25661 ;
  assign n38533 = ~n38531 & ~n38532 ;
  assign n38534 = \T_PIOin[1]_pad  & ~n25656 ;
  assign n38535 = \pio_PIO_IN_P_reg[1]/P0001  & n25656 ;
  assign n38536 = ~n38534 & ~n38535 ;
  assign n38537 = \T_PIOin[2]_pad  & ~n25666 ;
  assign n38538 = \pio_PIO_IN_P_reg[2]/P0001  & n25666 ;
  assign n38539 = ~n38537 & ~n38538 ;
  assign n38540 = \T_PIOin[3]_pad  & ~n25666 ;
  assign n38541 = \pio_PIO_IN_P_reg[3]/P0001  & n25666 ;
  assign n38542 = ~n38540 & ~n38541 ;
  assign n38543 = \T_PIOin[4]_pad  & ~n25679 ;
  assign n38544 = \pio_PIO_IN_P_reg[4]/P0001  & n25679 ;
  assign n38545 = ~n38543 & ~n38544 ;
  assign n38546 = \T_PIOin[5]_pad  & ~n25679 ;
  assign n38547 = \pio_PIO_IN_P_reg[5]/P0001  & n25679 ;
  assign n38548 = ~n38546 & ~n38547 ;
  assign n38549 = \T_PIOin[6]_pad  & ~n25671 ;
  assign n38550 = \pio_PIO_IN_P_reg[6]/P0001  & n25671 ;
  assign n38551 = ~n38549 & ~n38550 ;
  assign n38552 = \T_PIOin[7]_pad  & ~n25671 ;
  assign n38553 = \pio_PIO_IN_P_reg[7]/P0001  & n25671 ;
  assign n38554 = ~n38552 & ~n38553 ;
  assign n38555 = \T_PIOin[8]_pad  & ~n25651 ;
  assign n38556 = \pio_PIO_IN_P_reg[8]/P0001  & n25651 ;
  assign n38557 = ~n38555 & ~n38556 ;
  assign n38558 = \T_PIOin[9]_pad  & ~n25651 ;
  assign n38559 = \pio_PIO_IN_P_reg[9]/P0001  & n25651 ;
  assign n38560 = ~n38558 & ~n38559 ;
  assign n38561 = \pio_PIO_RES_reg[0]/NET0131  & ~n25656 ;
  assign n38562 = \pio_PIO_RES_OUT_reg[0]/P0001  & n25656 ;
  assign n38563 = ~n38561 & ~n38562 ;
  assign n38564 = \pio_PIO_RES_reg[10]/NET0131  & ~n25661 ;
  assign n38565 = \pio_PIO_RES_OUT_reg[10]/P0001  & n25661 ;
  assign n38566 = ~n38564 & ~n38565 ;
  assign n38567 = \pio_PIO_RES_reg[2]/NET0131  & ~n25666 ;
  assign n38568 = \pio_PIO_RES_OUT_reg[2]/P0001  & n25666 ;
  assign n38569 = ~n38567 & ~n38568 ;
  assign n38570 = \pio_PIO_RES_reg[4]/NET0131  & ~n25679 ;
  assign n38571 = \pio_PIO_RES_OUT_reg[4]/P0001  & n25679 ;
  assign n38572 = ~n38570 & ~n38571 ;
  assign n38573 = \pio_PIO_RES_reg[6]/NET0131  & ~n25671 ;
  assign n38574 = \pio_PIO_RES_OUT_reg[6]/P0001  & n25671 ;
  assign n38575 = ~n38573 & ~n38574 ;
  assign n38576 = \sice_GO_NXi_reg/NET0131  & ~n23033 ;
  assign n38577 = \sice_SPC_reg[20]/P0001  & n23033 ;
  assign n38578 = ~n38576 & ~n38577 ;
  assign n38579 = ~n20442 & n30779 ;
  assign n38580 = ~\sport0_rxctl_RXSHT_reg[0]/P0001  & ~n30779 ;
  assign n38581 = ~n38579 & ~n38580 ;
  assign n38582 = \sport0_rxctl_RXSHT_reg[1]/P0001  & ~n30779 ;
  assign n38583 = ~n30784 & ~n38582 ;
  assign n38584 = ~n20420 & n30755 ;
  assign n38585 = ~\sport1_rxctl_RXSHT_reg[0]/P0001  & ~n30755 ;
  assign n38586 = ~n38584 & ~n38585 ;
  assign n38587 = \sport1_rxctl_RXSHT_reg[1]/P0001  & ~n30755 ;
  assign n38588 = ~n30760 & ~n38587 ;
  assign CLKO_pad = n4047 ;
  assign \CMAinx[0]_pad  = ~n5073 ;
  assign \CMAinx[10]_pad  = ~n5120 ;
  assign \CMAinx[11]_pad  = ~n5149 ;
  assign \CMAinx[1]_pad  = ~n5176 ;
  assign \CMAinx[2]_pad  = ~n5215 ;
  assign \CMAinx[3]_pad  = ~n5252 ;
  assign \CMAinx[4]_pad  = ~n5286 ;
  assign \CMAinx[5]_pad  = ~n5318 ;
  assign \CMAinx[6]_pad  = ~n5345 ;
  assign \CMAinx[7]_pad  = ~n5372 ;
  assign \CMAinx[8]_pad  = ~n5399 ;
  assign \CMAinx[9]_pad  = ~n5426 ;
  assign CMSn_pad = n5613 ;
  assign CM_cs_pad = n5725 ;
  assign \CM_wd[0]_pad  = ~n5741 ;
  assign \CM_wd[10]_pad  = ~n5747 ;
  assign \CM_wd[11]_pad  = ~n5753 ;
  assign \CM_wd[12]_pad  = ~n5759 ;
  assign \CM_wd[13]_pad  = ~n5765 ;
  assign \CM_wd[14]_pad  = ~n5771 ;
  assign \CM_wd[15]_pad  = ~n5777 ;
  assign \CM_wd[16]_pad  = ~n5783 ;
  assign \CM_wd[17]_pad  = ~n5789 ;
  assign \CM_wd[18]_pad  = ~n5795 ;
  assign \CM_wd[19]_pad  = ~n5801 ;
  assign \CM_wd[1]_pad  = ~n5807 ;
  assign \CM_wd[20]_pad  = ~n5813 ;
  assign \CM_wd[21]_pad  = ~n5819 ;
  assign \CM_wd[22]_pad  = ~n5825 ;
  assign \CM_wd[23]_pad  = ~n5831 ;
  assign \CM_wd[2]_pad  = ~n5837 ;
  assign \CM_wd[3]_pad  = ~n5843 ;
  assign \CM_wd[4]_pad  = ~n5849 ;
  assign \CM_wd[5]_pad  = ~n5855 ;
  assign \CM_wd[6]_pad  = ~n5861 ;
  assign \CM_wd[7]_pad  = ~n5867 ;
  assign \CM_wd[8]_pad  = ~n5873 ;
  assign \CM_wd[9]_pad  = ~n5879 ;
  assign CM_web_pad = n5891 ;
  assign \CMo_cs0_pad  = n5924 ;
  assign \CMo_cs1_pad  = n5925 ;
  assign \CMo_cs2_pad  = n5927 ;
  assign \CMo_cs3_pad  = n5928 ;
  assign \CMo_cs4_pad  = n5931 ;
  assign \CMo_cs5_pad  = n5932 ;
  assign \CMo_cs6_pad  = n5934 ;
  assign \CMo_cs7_pad  = n5935 ;
  assign \DMAinx[0]_pad  = n7628 ;
  assign \DMAinx[10]_pad  = ~n8230 ;
  assign \DMAinx[11]_pad  = ~n8835 ;
  assign \DMAinx[12]_pad  = ~n9440 ;
  assign \DMAinx[13]_pad  = ~n9513 ;
  assign \DMAinx[1]_pad  = ~n9585 ;
  assign \DMAinx[2]_pad  = ~n9651 ;
  assign \DMAinx[3]_pad  = n9717 ;
  assign \DMAinx[4]_pad  = n10308 ;
  assign \DMAinx[5]_pad  = ~n10916 ;
  assign \DMAinx[6]_pad  = ~n11530 ;
  assign \DMAinx[7]_pad  = ~n11596 ;
  assign \DMAinx[8]_pad  = n11660 ;
  assign \DMAinx[9]_pad  = ~n11726 ;
  assign DMSn_pad = ~n5602 ;
  assign DM_cs_pad = n11767 ;
  assign \DM_wd[0]_pad  = ~n11780 ;
  assign \DM_wd[10]_pad  = ~n11789 ;
  assign \DM_wd[11]_pad  = ~n11798 ;
  assign \DM_wd[12]_pad  = ~n11807 ;
  assign \DM_wd[13]_pad  = ~n11816 ;
  assign \DM_wd[14]_pad  = ~n11962 ;
  assign \DM_wd[15]_pad  = ~n12104 ;
  assign \DM_wd[1]_pad  = ~n12113 ;
  assign \DM_wd[2]_pad  = ~n12122 ;
  assign \DM_wd[3]_pad  = ~n12131 ;
  assign \DM_wd[4]_pad  = ~n12140 ;
  assign \DM_wd[5]_pad  = ~n12149 ;
  assign \DM_wd[6]_pad  = ~n12158 ;
  assign \DM_wd[7]_pad  = ~n12167 ;
  assign \DM_wd[8]_pad  = ~n12176 ;
  assign \DM_wd[9]_pad  = ~n12185 ;
  assign \DMo_cs0_pad  = n12214 ;
  assign \DMo_cs1_pad  = n12217 ;
  assign \DMo_cs2_pad  = n12220 ;
  assign \DMo_cs3_pad  = n12222 ;
  assign \DMo_cs4_pad  = n12226 ;
  assign \DMo_cs5_pad  = n12229 ;
  assign \DMo_cs6_pad  = n12231 ;
  assign \DMo_cs7_pad  = n12233 ;
  assign \DSPCLK_cm1_pad  = ~n12245 ;
  assign \EA_do[0]_pad  = ~n12260 ;
  assign \EA_do[10]_pad  = ~n12270 ;
  assign \EA_do[12]_pad  = ~n12296 ;
  assign \EA_do[13]_pad  = ~n12316 ;
  assign \EA_do[14]_pad  = ~n12336 ;
  assign \EA_do[1]_pad  = ~n12348 ;
  assign \EA_do[2]_pad  = ~n12360 ;
  assign \EA_do[3]_pad  = ~n12372 ;
  assign \EA_do[4]_pad  = ~n12384 ;
  assign \EA_do[5]_pad  = ~n12396 ;
  assign \EA_do[6]_pad  = ~n12408 ;
  assign \EA_do[7]_pad  = ~n12420 ;
  assign \EA_do[8]_pad  = ~n12430 ;
  assign \EA_do[9]_pad  = ~n12440 ;
  assign EA_oe_pad = n12450 ;
  assign \ED_do[0]_pad  = ~n12527 ;
  assign \ED_do[10]_pad  = ~n12561 ;
  assign \ED_do[11]_pad  = ~n12595 ;
  assign \ED_do[12]_pad  = ~n12629 ;
  assign \ED_do[13]_pad  = ~n12663 ;
  assign \ED_do[14]_pad  = ~n12720 ;
  assign \ED_do[15]_pad  = ~n12774 ;
  assign \ED_do[1]_pad  = ~n12808 ;
  assign \ED_do[2]_pad  = ~n12842 ;
  assign \ED_do[3]_pad  = ~n12876 ;
  assign \ED_do[4]_pad  = ~n12910 ;
  assign \ED_do[5]_pad  = ~n12944 ;
  assign \ED_do[6]_pad  = ~n12978 ;
  assign \ED_do[7]_pad  = ~n13012 ;
  assign \ED_do[8]_pad  = ~n13046 ;
  assign \ED_do[9]_pad  = ~n13080 ;
  assign \ED_oe_14_8_pad  = ~n13081 ;
  assign \ED_oe_7_0_pad  = ~n13082 ;
  assign \IAD_do[0]_pad  = n13087 ;
  assign \IAD_do[10]_pad  = ~n13089 ;
  assign \IAD_do[11]_pad  = n13091 ;
  assign \IAD_do[12]_pad  = n13092 ;
  assign \IAD_do[13]_pad  = ~n13094 ;
  assign \IAD_do[14]_pad  = n13095 ;
  assign \IAD_do[15]_pad  = ~n13097 ;
  assign \IAD_do[1]_pad  = n13101 ;
  assign \IAD_do[2]_pad  = ~n13105 ;
  assign \IAD_do[3]_pad  = n13109 ;
  assign \IAD_do[4]_pad  = n13113 ;
  assign \IAD_do[5]_pad  = ~n13117 ;
  assign \IAD_do[6]_pad  = n13121 ;
  assign \IAD_do[7]_pad  = ~n13125 ;
  assign \IAD_do[8]_pad  = n13126 ;
  assign \IAD_do[9]_pad  = n13127 ;
  assign IAD_oe_pad = ~n13128 ;
  assign IDoe_pad = n13129 ;
  assign IOSn_pad = ~n5610 ;
  assign \PMAinx[0]_pad  = ~n13173 ;
  assign \PMAinx[10]_pad  = ~n13192 ;
  assign \PMAinx[11]_pad  = ~n13211 ;
  assign \PMAinx[1]_pad  = ~n13230 ;
  assign \PMAinx[2]_pad  = ~n13249 ;
  assign \PMAinx[3]_pad  = n13268 ;
  assign \PMAinx[4]_pad  = n13287 ;
  assign \PMAinx[5]_pad  = n13306 ;
  assign \PMAinx[6]_pad  = n13325 ;
  assign \PMAinx[7]_pad  = n13344 ;
  assign \PMAinx[8]_pad  = n13363 ;
  assign \PMAinx[9]_pad  = n13382 ;
  assign \PM_wd[0]_pad  = n13392 ;
  assign \PM_wd[10]_pad  = n13399 ;
  assign \PM_wd[11]_pad  = n13406 ;
  assign \PM_wd[12]_pad  = n13413 ;
  assign \PM_wd[13]_pad  = n13420 ;
  assign \PM_wd[14]_pad  = n13427 ;
  assign \PM_wd[15]_pad  = n13434 ;
  assign \PM_wd[1]_pad  = n13441 ;
  assign \PM_wd[2]_pad  = n13448 ;
  assign \PM_wd[3]_pad  = n13455 ;
  assign \PM_wd[4]_pad  = n13462 ;
  assign \PM_wd[5]_pad  = n13469 ;
  assign \PM_wd[6]_pad  = n13476 ;
  assign \PM_wd[7]_pad  = n13483 ;
  assign \PM_wd[8]_pad  = n13490 ;
  assign \PM_wd[9]_pad  = n13497 ;
  assign \PMo_cs0_pad  = n13588 ;
  assign \PMo_cs1_pad  = n13591 ;
  assign \PMo_cs2_pad  = n13594 ;
  assign \PMo_cs3_pad  = n13596 ;
  assign \PMo_cs4_pad  = n13601 ;
  assign \PMo_cs5_pad  = n13604 ;
  assign \PMo_cs6_pad  = n13606 ;
  assign \PMo_cs7_pad  = n13608 ;
  assign \PMo_oe0_pad  = ~1'b0 ;
  assign \RFS0_pad  = ~n13613 ;
  assign \RFS1_pad  = ~n13618 ;
  assign \SCLK0_pad  = ~n13621 ;
  assign \SCLK1_pad  = ~n13624 ;
  assign \TD0_pad  = n13672 ;
  assign \TD1_pad  = n13721 ;
  assign \TFS0_pad  = ~n13725 ;
  assign \TFS1_pad  = ~n13729 ;
  assign \T_ISn_syn_2  = ~T_ISn_pad ;
  assign WRn_pad = ~n13732 ;
  assign XTALoffn_pad = ~n12239 ;
  assign \_al_n0  = 1'b0 ;
  assign \bdma_BDMA_boot_reg/NET0131_reg_syn_3  = ~n13759 ;
  assign \bdma_BDMA_boot_reg/n0  = n13734 ;
  assign \bdma_BM_cyc_reg/P0000  = ~\bdma_BM_cyc_reg/P0001  ;
  assign \bdma_BWCOUNT_reg[5]/NET0131_reg_syn_3  = ~n13774 ;
  assign \core_c_psq_MGNT_reg/P0001  = ~\core_c_psq_MGNT_reg/NET0131  ;
  assign \core_c_psq_cntstk_cnts4x14_CNTcell_reg[0][5]/P0001_reg_syn_3  = ~n13783 ;
  assign \core_c_psq_cntstk_cnts4x14_CNTcell_reg[1][5]/P0001_reg_syn_3  = ~n13788 ;
  assign \core_c_psq_cntstk_cnts4x14_CNTcell_reg[2][5]/P0001_reg_syn_3  = ~n13793 ;
  assign \core_c_psq_cntstk_cnts4x14_CNTcell_reg[3][5]/P0001_reg_syn_3  = ~n13798 ;
  assign \core_eu_ea_alu_ea_reg_afrwe_DO_reg[12]/P0001_reg_syn_3  = n14429 ;
  assign \core_eu_ea_alu_ea_reg_afrwe_DO_reg[14]/P0001_reg_syn_3  = n14556 ;
  assign \core_eu_ea_alu_ea_reg_afrwe_DO_reg[1]/P0001_reg_syn_3  = ~n14578 ;
  assign \core_eu_ea_alu_ea_reg_afrwe_DO_reg[2]/P0001_reg_syn_3  = ~n14592 ;
  assign \core_eu_ea_alu_ea_reg_afrwe_DO_reg[4]/P0001_reg_syn_3  = ~n14615 ;
  assign \core_eu_ea_alu_ea_reg_afrwe_DO_reg[6]/P0001_reg_syn_3  = ~n14639 ;
  assign \core_eu_ea_alu_ea_reg_afrwe_DO_reg[9]/P0001_reg_syn_3  = ~n14663 ;
  assign \core_eu_ea_alu_ea_reg_afswe_DO_reg[12]/P0001_reg_syn_3  = n14670 ;
  assign \core_eu_ea_alu_ea_reg_afswe_DO_reg[14]/P0001_reg_syn_3  = n14673 ;
  assign \core_eu_ea_alu_ea_reg_afswe_DO_reg[1]/P0001_reg_syn_3  = ~n14676 ;
  assign \core_eu_ea_alu_ea_reg_afswe_DO_reg[2]/P0001_reg_syn_3  = ~n14679 ;
  assign \core_eu_ea_alu_ea_reg_afswe_DO_reg[4]/P0001_reg_syn_3  = ~n14682 ;
  assign \core_eu_ea_alu_ea_reg_afswe_DO_reg[6]/P0001_reg_syn_3  = ~n14685 ;
  assign \core_eu_ea_alu_ea_reg_afswe_DO_reg[9]/P0001_reg_syn_3  = ~n14688 ;
  assign \core_eu_ec_cun_MVi_pre_C_reg/P0001_reg_syn_3  = ~n14725 ;
  assign \core_eu_em_mac_em_reg_Sq_E_reg/P0001_reg_syn_3  = n14731 ;
  assign \emc_DMDreg_reg[8]/P0001_reg_syn_3  = ~n14740 ;
  assign \emc_DMDreg_reg[9]/P0001_reg_syn_3  = ~n14743 ;
  assign \emc_ECMcs_reg/P0001  = ~\emc_ECMcs_reg/NET0131  ;
  assign \emc_PMDreg_reg[8]/P0001_reg_syn_3  = ~n14748 ;
  assign \emc_PMDreg_reg[9]/P0001_reg_syn_3  = ~n14751 ;
  assign \g10/_0_  = n17831 ;
  assign \g1000/_0_  = n18216 ;
  assign \g10000/_0_  = ~n18224 ;
  assign \g10001/_0_  = ~n18239 ;
  assign \g10002/_0_  = ~n18243 ;
  assign \g10003/_0_  = ~n18246 ;
  assign \g10004/_0_  = ~n18249 ;
  assign \g10005/_0_  = ~n18252 ;
  assign \g10007/_0_  = ~n18255 ;
  assign \g10008/_0_  = ~n18258 ;
  assign \g10009/_0_  = ~n18261 ;
  assign \g1001/_3_  = ~n18293 ;
  assign \g10010/_0_  = ~n18296 ;
  assign \g10011/_0_  = ~n18299 ;
  assign \g10012/_0_  = ~n18302 ;
  assign \g10013/_0_  = ~n18305 ;
  assign \g10014/_0_  = ~n18308 ;
  assign \g10015/_0_  = ~n18311 ;
  assign \g10016/_0_  = ~n18314 ;
  assign \g10017/_0_  = ~n18317 ;
  assign \g10018/_0_  = ~n18320 ;
  assign \g10019/_0_  = ~n18323 ;
  assign \g1002/_3_  = n18337 ;
  assign \g10020/_0_  = ~n18340 ;
  assign \g10021/_0_  = ~n18343 ;
  assign \g10022/_0_  = ~n18346 ;
  assign \g10023/_0_  = ~n18349 ;
  assign \g10024/_0_  = ~n18352 ;
  assign \g10025/_0_  = ~n18355 ;
  assign \g10026/_0_  = ~n18358 ;
  assign \g10027/_0_  = ~n18361 ;
  assign \g10028/_0_  = ~n18365 ;
  assign \g10029/_0_  = ~n18368 ;
  assign \g1003/_0_  = n18524 ;
  assign \g10030/_0_  = ~n18527 ;
  assign \g10031/_0_  = ~n18530 ;
  assign \g10032/_0_  = ~n18533 ;
  assign \g10033/_0_  = ~n18536 ;
  assign \g10034/_0_  = ~n18539 ;
  assign \g10035/_0_  = ~n18542 ;
  assign \g10036/_0_  = ~n18545 ;
  assign \g10037/_0_  = ~n18548 ;
  assign \g10038/_0_  = ~n18551 ;
  assign \g10039/_0_  = ~n18554 ;
  assign \g10040/_0_  = ~n18557 ;
  assign \g10041/_0_  = ~n18560 ;
  assign \g10042/_0_  = ~n18563 ;
  assign \g10043/_0_  = ~n18566 ;
  assign \g10044/_0_  = ~n18569 ;
  assign \g10045/_0_  = ~n18572 ;
  assign \g10046/_0_  = ~n18575 ;
  assign \g10047/_0_  = ~n18578 ;
  assign \g10048/_0_  = ~n18581 ;
  assign \g10049/_0_  = ~n18584 ;
  assign \g10050/_0_  = ~n18587 ;
  assign \g10051/_0_  = ~n18590 ;
  assign \g10052/_0_  = ~n18593 ;
  assign \g10053/_0_  = ~n18597 ;
  assign \g10054/_0_  = ~n18600 ;
  assign \g10055/_0_  = ~n18603 ;
  assign \g10056/_0_  = ~n18606 ;
  assign \g10057/_0_  = ~n18609 ;
  assign \g10058/_0_  = ~n18612 ;
  assign \g10059/_0_  = ~n18615 ;
  assign \g10060/_0_  = ~n18618 ;
  assign \g10061/_0_  = ~n18621 ;
  assign \g10062/_0_  = ~n18624 ;
  assign \g10063/_0_  = ~n18627 ;
  assign \g10064/_0_  = ~n18630 ;
  assign \g10065/_0_  = ~n18633 ;
  assign \g10066/_0_  = ~n18636 ;
  assign \g10067/_0_  = ~n18639 ;
  assign \g10068/_0_  = ~n18642 ;
  assign \g10069/_0_  = ~n18645 ;
  assign \g10070/_0_  = ~n18648 ;
  assign \g10071/_0_  = ~n18651 ;
  assign \g10072/_0_  = ~n18657 ;
  assign \g10073/_0_  = ~n18660 ;
  assign \g10074/_0_  = ~n18663 ;
  assign \g10075/_0_  = ~n18666 ;
  assign \g10076/_0_  = ~n18669 ;
  assign \g10077/_0_  = ~n18672 ;
  assign \g10078/_0_  = ~n18675 ;
  assign \g10080/_0_  = ~n18678 ;
  assign \g10081/_0_  = ~n18687 ;
  assign \g10083/_0_  = ~n18692 ;
  assign \g10089/_0_  = ~n18695 ;
  assign \g1009/_0_  = ~n18701 ;
  assign \g10090/_0_  = ~n18704 ;
  assign \g10091/_0_  = ~n18707 ;
  assign \g10092/_0_  = ~n18710 ;
  assign \g10093/_0_  = ~n18713 ;
  assign \g10094/_0_  = ~n18716 ;
  assign \g1010/_0_  = n18836 ;
  assign \g10108/_3_  = ~n18852 ;
  assign \g1011/_0_  = ~n18855 ;
  assign \g10110/_0_  = n18864 ;
  assign \g10111/_0_  = n18873 ;
  assign \g10113/_3_  = ~n18877 ;
  assign \g10115/_3_  = ~n18881 ;
  assign \g1013/_0_  = n18884 ;
  assign \g1014/_0_  = n18945 ;
  assign \g10152/_0_  = ~n18950 ;
  assign \g10153/_0_  = ~n18953 ;
  assign \g10154/_0_  = ~n18956 ;
  assign \g10155/_0_  = n18959 ;
  assign \g10156/_0_  = ~n18962 ;
  assign \g10157/_0_  = ~n18965 ;
  assign \g10158/_0_  = ~n18968 ;
  assign \g10159/_0_  = n18971 ;
  assign \g1016/_0_  = n19013 ;
  assign \g10160/_0_  = ~n19017 ;
  assign \g10161/_0_  = ~n19020 ;
  assign \g10162/_0_  = ~n19023 ;
  assign \g10163/_0_  = n19027 ;
  assign \g10164/_0_  = ~n19030 ;
  assign \g10165/_0_  = ~n19033 ;
  assign \g1017/_0_  = n19037 ;
  assign \g10170/_3_  = ~n19059 ;
  assign \g1018/_0_  = n19062 ;
  assign \g10190/_3_  = n19064 ;
  assign \g10194/_3_  = ~n19066 ;
  assign \g10198/_0_  = ~n19133 ;
  assign \g10199/_0_  = ~n19200 ;
  assign \g102/_0_  = n19363 ;
  assign \g103/_0_  = ~n19392 ;
  assign \g104/_0_  = ~n19402 ;
  assign \g105/_0_  = ~n19409 ;
  assign \g10598/_0_  = n19413 ;
  assign \g106/_0_  = ~n19436 ;
  assign \g10667/_0_  = n19440 ;
  assign \g10683/_0_  = n19476 ;
  assign \g10685/_0_  = ~n19498 ;
  assign \g107/_0_  = ~n19527 ;
  assign \g10721/_0_  = n19533 ;
  assign \g10758/_0_  = n19540 ;
  assign \g10765/_0_  = n19543 ;
  assign \g10778/_0_  = n19554 ;
  assign \g10791/_0_  = n19555 ;
  assign \g108/_0_  = ~n19694 ;
  assign \g10887/_0_  = n19707 ;
  assign \g1089/_0_  = n19774 ;
  assign \g109/_0_  = n19783 ;
  assign \g1090/_0_  = n19845 ;
  assign \g1091/_0_  = n19900 ;
  assign \g1092/_0_  = n19903 ;
  assign \g10923/_0_  = n19906 ;
  assign \g1093/_0_  = n19909 ;
  assign \g10930/_0_  = n19915 ;
  assign \g10931/_0_  = n19918 ;
  assign \g10936/_0_  = ~n19926 ;
  assign \g1097/_0_  = n19929 ;
  assign \g11/_0_  = ~n19963 ;
  assign \g110/_0_  = n19969 ;
  assign \g1101/_0_  = n20035 ;
  assign \g11013/_0_  = n20044 ;
  assign \g1102/_0_  = ~n20058 ;
  assign \g1103/_0_  = ~n20061 ;
  assign \g11032/_0_  = ~n20077 ;
  assign \g1104/_0_  = n20147 ;
  assign \g1105/_0_  = n20197 ;
  assign \g1107/_0_  = n20200 ;
  assign \g11074/_0_  = n20222 ;
  assign \g11077/_0_  = n20225 ;
  assign \g1108/_0_  = n20228 ;
  assign \g1109/_0_  = n20231 ;
  assign \g11112/_0_  = n20242 ;
  assign \g11115/_0_  = n20245 ;
  assign \g11116/_0_  = n20248 ;
  assign \g11119/_0_  = n20255 ;
  assign \g11120/_0_  = n20256 ;
  assign \g1113/_0_  = n20293 ;
  assign \g1115/_0_  = n20331 ;
  assign \g1116/_0_  = n20334 ;
  assign \g1117/_0_  = n20337 ;
  assign \g11267/_0_  = n20340 ;
  assign \g11281/_0_  = ~n20353 ;
  assign \g11287/_0_  = n20375 ;
  assign \g11300/_0_  = ~n20380 ;
  assign \g11323/_0_  = ~n20385 ;
  assign \g11325/_2__syn_2  = n20396 ;
  assign \g11345/_2_  = ~n20399 ;
  assign \g11470/_0_  = n20405 ;
  assign \g11471/_0_  = n20423 ;
  assign \g11472/_0_  = n20427 ;
  assign \g11473/_0_  = n20445 ;
  assign \g11474/_0_  = n20449 ;
  assign \g11476/_0_  = n20452 ;
  assign \g11477/_0_  = n20463 ;
  assign \g11496/_0_  = ~n20482 ;
  assign \g11497/_0_  = ~n20491 ;
  assign \g11498/_0_  = ~n20500 ;
  assign \g11499/_0_  = ~n20506 ;
  assign \g11500/_0_  = ~n20515 ;
  assign \g11501/_0_  = ~n20521 ;
  assign \g11502/_0_  = ~n20530 ;
  assign \g11503/_0_  = ~n20536 ;
  assign \g11504/_0_  = ~n20544 ;
  assign \g11505/_0_  = ~n20552 ;
  assign \g11506/_0_  = ~n20558 ;
  assign \g11507/_0_  = ~n20564 ;
  assign \g11509/_0_  = n20567 ;
  assign \g11510/_0_  = n20570 ;
  assign \g11515/_0_  = ~n20588 ;
  assign \g11516/_0_  = n20591 ;
  assign \g11520/_0_  = ~n20594 ;
  assign \g11521/_0_  = ~n20600 ;
  assign \g11576/_0_  = n20612 ;
  assign \g11577/_0_  = n20622 ;
  assign \g11578/_0_  = n20632 ;
  assign \g11579/_0_  = n20642 ;
  assign \g11580/_0_  = n20652 ;
  assign \g11581/_0_  = n20660 ;
  assign \g11582/_0_  = n20671 ;
  assign \g11583/_0_  = n20682 ;
  assign \g11584/_0_  = n20693 ;
  assign \g11585/_0_  = n20704 ;
  assign \g11586/_0_  = n20715 ;
  assign \g11587/_0_  = n20726 ;
  assign \g11588/_0_  = n20737 ;
  assign \g11589/_0_  = n20753 ;
  assign \g11591/_0_  = n20763 ;
  assign \g11593/_0_  = ~n20773 ;
  assign \g11595/_0_  = ~n20780 ;
  assign \g11596/_0_  = ~n20783 ;
  assign \g11597/_0_  = n20786 ;
  assign \g11605/_0_  = n20791 ;
  assign \g11606/_0_  = n20794 ;
  assign \g11607/_0_  = n20797 ;
  assign \g11608/_0_  = n20800 ;
  assign \g11609/_0_  = n20803 ;
  assign \g11610/_0_  = n20806 ;
  assign \g11611/_0_  = n20809 ;
  assign \g11612/_0_  = n20812 ;
  assign \g11613/_0_  = n20815 ;
  assign \g11615/_0_  = n20820 ;
  assign \g11616/_0_  = n20832 ;
  assign \g11617/_0_  = n20837 ;
  assign \g11651/_3_  = ~n20840 ;
  assign \g11704/_0_  = n20842 ;
  assign \g11705/_0_  = n20844 ;
  assign \g11709/_0_  = n20852 ;
  assign \g11722/_0_  = n20861 ;
  assign \g11723/_0_  = n20863 ;
  assign \g119/_0_  = ~n20867 ;
  assign \g1192/_0_  = ~n20988 ;
  assign \g11994/_0_  = n20989 ;
  assign \g120/_0_  = ~n20993 ;
  assign \g1200/_0_  = n21051 ;
  assign \g12003/_0_  = n21054 ;
  assign \g1201/_0_  = n21057 ;
  assign \g12019/_0_  = n21060 ;
  assign \g1203/_3_  = ~n21070 ;
  assign \g1204/_3_  = n21076 ;
  assign \g1207/_0_  = n21129 ;
  assign \g1208/_0_  = n21132 ;
  assign \g12092/_0_  = ~n21140 ;
  assign \g1210/_0_  = n21179 ;
  assign \g1211/_0_  = n21231 ;
  assign \g1212/_0_  = n21234 ;
  assign \g1213/_0_  = n21237 ;
  assign \g12145/_0_  = n21246 ;
  assign \g12155/_0_  = n21254 ;
  assign \g12186/_0_  = n21261 ;
  assign \g12187/_0_  = n21264 ;
  assign \g12192/_0_  = n21267 ;
  assign \g12201/_0_  = ~n21276 ;
  assign \g12202/_0_  = ~n21280 ;
  assign \g12203/_0_  = ~n21284 ;
  assign \g12204/_0_  = ~n21287 ;
  assign \g12207/_0_  = n21290 ;
  assign \g12229/_3_  = n21300 ;
  assign \g12267/_0_  = ~n21301 ;
  assign \g12276/_0_  = n21304 ;
  assign \g12278/_0_  = n21307 ;
  assign \g12279/_0_  = n21310 ;
  assign \g12280/_0_  = n21313 ;
  assign \g12302/_0_  = ~n21315 ;
  assign \g12316/_0_  = ~n21322 ;
  assign \g12317/_0_  = ~n21326 ;
  assign \g12319/_0_  = ~n21330 ;
  assign \g12328/_3_  = n21339 ;
  assign \g1233/_0_  = n10069 ;
  assign \g12348/_0_  = ~n21343 ;
  assign \g12351/_0_  = ~n21347 ;
  assign \g12352/_0_  = ~n21351 ;
  assign \g12353/_0_  = ~n21355 ;
  assign \g12354/_0_  = ~n21359 ;
  assign \g12355/_0_  = ~n21363 ;
  assign \g1237/_0_  = n8113 ;
  assign \g124/_0_  = ~n21366 ;
  assign \g12444/_0_  = ~n21371 ;
  assign \g125/_0_  = ~n21374 ;
  assign \g12637/_0_  = n21382 ;
  assign \g12639/_0_  = n21390 ;
  assign \g12658/_0_  = n21399 ;
  assign \g12659/_0_  = ~n21409 ;
  assign \g12660/_0_  = ~n21419 ;
  assign \g12663/_0_  = ~n21425 ;
  assign \g12664/_0_  = n21432 ;
  assign \g12665/_0_  = n21437 ;
  assign \g12672/_3_  = n21446 ;
  assign \g12673/_3_  = n21455 ;
  assign \g12674/_3_  = n21464 ;
  assign \g12675/_3_  = n21473 ;
  assign \g12676/_3_  = n21482 ;
  assign \g12677/_3_  = n21491 ;
  assign \g12678/_0_  = ~n21496 ;
  assign \g12679/_3_  = n21505 ;
  assign \g12697/_3_  = n21514 ;
  assign \g12701/_3_  = n21523 ;
  assign \g12711/_2_  = ~n21535 ;
  assign \g12713/_2_  = ~n21541 ;
  assign \g12715/_2_  = ~n21549 ;
  assign \g12717/_2_  = ~n21555 ;
  assign \g12718/_2__syn_2  = ~n21562 ;
  assign \g1272/_0_  = ~n21577 ;
  assign \g12728/_1__syn_2  = ~n21579 ;
  assign \g12730/_3_  = n21588 ;
  assign \g12741/_1__syn_2  = ~n21592 ;
  assign \g12746/_0__syn_2  = ~n18689 ;
  assign \g12748/_0_  = ~n21598 ;
  assign \g12749/_0_  = ~n21601 ;
  assign \g12759/_1__syn_2  = ~n18233 ;
  assign \g12760/_0_  = n21605 ;
  assign \g12762/_0_  = ~n21609 ;
  assign \g12763/_0_  = ~n21612 ;
  assign \g12764/_0_  = ~n21615 ;
  assign \g12765/_0_  = ~n21618 ;
  assign \g12766/_0_  = ~n21621 ;
  assign \g12767/_0_  = ~n21624 ;
  assign \g12768/_0_  = ~n21627 ;
  assign \g12769/_0_  = ~n21630 ;
  assign \g12770/_0_  = ~n21633 ;
  assign \g12771/_0_  = ~n21636 ;
  assign \g12772/_0_  = ~n21639 ;
  assign \g12773/_0_  = ~n21642 ;
  assign \g12774/_0_  = ~n21645 ;
  assign \g12775/_0_  = ~n21648 ;
  assign \g12776/_0_  = ~n21651 ;
  assign \g12777/_0_  = ~n21654 ;
  assign \g12778/_0_  = ~n21657 ;
  assign \g12779/_0_  = ~n21660 ;
  assign \g1278/_0_  = n21705 ;
  assign \g12780/_0_  = ~n21709 ;
  assign \g12781/_0_  = ~n21712 ;
  assign \g12782/_0_  = ~n21715 ;
  assign \g12783/_0_  = ~n21718 ;
  assign \g12784/_0_  = ~n21721 ;
  assign \g12785/_0_  = ~n21724 ;
  assign \g12786/_0_  = ~n21727 ;
  assign \g12787/_0_  = ~n21730 ;
  assign \g12788/_0_  = ~n21733 ;
  assign \g12789/_0_  = ~n21736 ;
  assign \g12790/_0_  = ~n21739 ;
  assign \g12791/_0_  = ~n21742 ;
  assign \g12792/_0_  = ~n21745 ;
  assign \g12793/_0_  = ~n21748 ;
  assign \g12794/_0_  = ~n21751 ;
  assign \g12795/_0_  = ~n21754 ;
  assign \g12796/_0_  = ~n21757 ;
  assign \g12797/_0_  = ~n21760 ;
  assign \g12798/_0_  = ~n21764 ;
  assign \g12799/_0_  = ~n21767 ;
  assign \g12800/_0_  = ~n21770 ;
  assign \g12801/_0_  = ~n21773 ;
  assign \g12802/_0_  = ~n21776 ;
  assign \g12803/_0_  = ~n21779 ;
  assign \g12804/_0_  = ~n21782 ;
  assign \g12805/_0_  = ~n21785 ;
  assign \g12806/_0_  = ~n21788 ;
  assign \g12807/_0_  = ~n21791 ;
  assign \g12808/_0_  = ~n21794 ;
  assign \g12809/_0_  = ~n21797 ;
  assign \g1281/_0_  = ~n21803 ;
  assign \g12810/_0_  = ~n21806 ;
  assign \g12811/_0_  = ~n21809 ;
  assign \g12812/_0_  = ~n21812 ;
  assign \g12813/_0_  = ~n21815 ;
  assign \g12814/_0_  = ~n21818 ;
  assign \g12815/_0_  = ~n21821 ;
  assign \g12816/_0_  = ~n21824 ;
  assign \g12817/_0_  = ~n21827 ;
  assign \g12818/_0_  = ~n21830 ;
  assign \g12819/_0_  = ~n21833 ;
  assign \g1282/_0_  = ~n21836 ;
  assign \g12820/_0_  = ~n21839 ;
  assign \g12821/_0_  = ~n21842 ;
  assign \g12822/_0_  = ~n21845 ;
  assign \g12823/_0_  = ~n21848 ;
  assign \g12824/_0_  = ~n21851 ;
  assign \g12825/_0_  = ~n21854 ;
  assign \g12826/_0_  = ~n21857 ;
  assign \g12827/_0_  = ~n21860 ;
  assign \g12828/_0_  = ~n21863 ;
  assign \g12829/_0_  = ~n21866 ;
  assign \g12830/_0_  = ~n21869 ;
  assign \g12831/_0_  = n21873 ;
  assign \g12832/_0_  = n21879 ;
  assign \g12833/_0_  = ~n21881 ;
  assign \g12835/_0_  = ~n21884 ;
  assign \g12836/_0_  = ~n21887 ;
  assign \g12838/_0_  = ~n21890 ;
  assign \g12848/_0_  = n21895 ;
  assign \g12849/_0_  = n21899 ;
  assign \g1285/_0_  = n21902 ;
  assign \g12850/_0_  = ~n21905 ;
  assign \g12857/_0_  = n21909 ;
  assign \g12858/_0_  = n21912 ;
  assign \g12859/_0_  = n21915 ;
  assign \g12861/_0_  = n21918 ;
  assign \g12862/_0_  = n21921 ;
  assign \g12868/_0_  = n21926 ;
  assign \g12869/_0_  = n21929 ;
  assign \g1287/_0_  = n21963 ;
  assign \g12870/_0_  = n21966 ;
  assign \g12871/_0_  = n21969 ;
  assign \g12872/_0_  = n21972 ;
  assign \g12873/_0_  = n21975 ;
  assign \g12874/_0_  = n21979 ;
  assign \g12875/_0_  = n21982 ;
  assign \g12876/_0_  = n21985 ;
  assign \g12877/_0_  = n21988 ;
  assign \g12878/_0_  = n22000 ;
  assign \g12879/_0_  = n22009 ;
  assign \g12880/_0_  = n22018 ;
  assign \g12881/_0_  = n22027 ;
  assign \g12882/_0_  = n22036 ;
  assign \g12883/_0_  = n22045 ;
  assign \g12884/_0_  = n22054 ;
  assign \g12885/_0_  = n22063 ;
  assign \g12886/_0_  = n22072 ;
  assign \g12887/_0_  = n22081 ;
  assign \g12888/_0_  = n22090 ;
  assign \g12889/_0_  = n22099 ;
  assign \g1289/_0_  = n22102 ;
  assign \g12890/_0_  = n22111 ;
  assign \g12891/_0_  = n22120 ;
  assign \g12894/_0_  = n22123 ;
  assign \g12898/_0_  = n22127 ;
  assign \g12899/_0_  = n22130 ;
  assign \g12900/_0_  = n22133 ;
  assign \g12901/_0_  = n22136 ;
  assign \g12902/_0_  = n22139 ;
  assign \g12903/_0_  = n22142 ;
  assign \g12906/_0_  = n22145 ;
  assign \g12907/_0_  = n22148 ;
  assign \g12908/_0_  = ~n22157 ;
  assign \g12912/_0_  = n22161 ;
  assign \g12913/_0_  = n22164 ;
  assign \g12914/_0_  = n22167 ;
  assign \g12915/_0_  = n22170 ;
  assign \g12916/_0_  = n22173 ;
  assign \g12917/_0_  = n22176 ;
  assign \g12918/_0_  = n22179 ;
  assign \g12919/_0_  = n22182 ;
  assign \g12920/_0_  = ~n22185 ;
  assign \g12921/_0_  = n22188 ;
  assign \g12922/_0_  = n22191 ;
  assign \g12923/_0_  = n22194 ;
  assign \g12924/_0_  = n22197 ;
  assign \g12925/_0_  = n22200 ;
  assign \g12926/_0_  = n22203 ;
  assign \g12932/_0_  = n22206 ;
  assign \g12933/_0_  = n22209 ;
  assign \g12936/_0_  = n22212 ;
  assign \g12955/_0_  = n22215 ;
  assign \g13015/_0_  = n22218 ;
  assign \g13016/_0_  = n22221 ;
  assign \g13017/_0_  = n22224 ;
  assign \g13018/_0_  = n22227 ;
  assign \g13019/_0_  = n22229 ;
  assign \g13020/_0_  = n22232 ;
  assign \g13021/_0_  = n22235 ;
  assign \g13024/_0_  = n22238 ;
  assign \g13025/_0_  = n22241 ;
  assign \g13027/_0_  = n22244 ;
  assign \g13028/_0_  = n22247 ;
  assign \g13030/_0_  = n22250 ;
  assign \g13031/_0_  = n22253 ;
  assign \g13033/_0_  = n22256 ;
  assign \g13047/_0_  = n22259 ;
  assign \g13060/_0_  = n22262 ;
  assign \g13062/_0_  = n22265 ;
  assign \g13063/_0_  = n22268 ;
  assign \g13064/_0_  = n22271 ;
  assign \g13067/_0_  = n22274 ;
  assign \g13068/_0_  = n22277 ;
  assign \g13069/_0_  = n22280 ;
  assign \g13070/_0_  = n22283 ;
  assign \g13072/_0_  = n22286 ;
  assign \g13094/_0_  = ~n22288 ;
  assign \g13104/_0_  = n22294 ;
  assign \g13110/_0_  = n22297 ;
  assign \g13114/_0_  = n22301 ;
  assign \g13115/_0_  = n22304 ;
  assign \g13116/_0_  = n22307 ;
  assign \g13117/_0_  = n22310 ;
  assign \g13118/_0_  = n22313 ;
  assign \g13119/_0_  = n22316 ;
  assign \g13120/_0_  = n22319 ;
  assign \g13121/_0_  = n22322 ;
  assign \g13124/_0_  = n22325 ;
  assign \g13125/_0_  = n22328 ;
  assign \g13127/_0_  = n22331 ;
  assign \g13128/_0_  = n22334 ;
  assign \g13129/_0_  = n22337 ;
  assign \g13130/_0_  = n22340 ;
  assign \g13131/_0_  = n22343 ;
  assign \g13132/_0_  = n22346 ;
  assign \g13133/_0_  = n22349 ;
  assign \g13134/_0_  = n22352 ;
  assign \g13138/_0_  = n22355 ;
  assign \g13139/_0_  = n22358 ;
  assign \g13140/_0_  = n22361 ;
  assign \g13141/_0_  = n22364 ;
  assign \g13142/_0_  = n22367 ;
  assign \g13143/_0_  = n22370 ;
  assign \g13144/_0_  = n22373 ;
  assign \g13146/_0_  = n22376 ;
  assign \g13150/_0_  = n22379 ;
  assign \g13152/_0_  = n22382 ;
  assign \g13154/_0_  = n22385 ;
  assign \g13155/_0_  = ~n22388 ;
  assign \g13156/_0_  = n22391 ;
  assign \g13157/_0_  = n22394 ;
  assign \g13158/_0_  = n22397 ;
  assign \g1320/_3_  = ~n22432 ;
  assign \g13266/_0_  = n22435 ;
  assign \g13269/_0_  = n22438 ;
  assign \g13274/_0_  = n22441 ;
  assign \g13277/_0_  = n22444 ;
  assign \g13280/_0_  = n22447 ;
  assign \g13283/_0_  = n22450 ;
  assign \g13294/_0_  = n22453 ;
  assign \g13330/_0_  = ~n22456 ;
  assign \g13333/_0_  = n22461 ;
  assign \g13334/_0_  = n22464 ;
  assign \g13335/_0_  = n22467 ;
  assign \g13336/_0_  = n22470 ;
  assign \g13337/_0_  = n22473 ;
  assign \g13338/_0_  = n22476 ;
  assign \g13345/_0_  = n22480 ;
  assign \g13346/_0_  = n22483 ;
  assign \g13347/_0_  = n22487 ;
  assign \g13348/_0_  = n22490 ;
  assign \g13349/_0_  = n22493 ;
  assign \g13350/_0_  = n22496 ;
  assign \g13351/_0_  = n22499 ;
  assign \g13352/_0_  = n22502 ;
  assign \g13486/_0_  = n22504 ;
  assign \g13488/_0_  = n22506 ;
  assign \g13508/_0_  = ~n22509 ;
  assign \g13509/_0_  = ~n22512 ;
  assign \g13510/_0_  = ~n22515 ;
  assign \g13511/_0_  = ~n22518 ;
  assign \g13512/_0_  = ~n22521 ;
  assign \g13513/_0_  = ~n22524 ;
  assign \g13514/_0_  = ~n22527 ;
  assign \g13515/_0_  = ~n22530 ;
  assign \g13516/_0_  = ~n22533 ;
  assign \g13517/_0_  = ~n22536 ;
  assign \g13518/_0_  = ~n22539 ;
  assign \g13519/_0_  = ~n22542 ;
  assign \g13520/_0_  = ~n22545 ;
  assign \g13521/_0_  = ~n22548 ;
  assign \g13540/_0_  = n22551 ;
  assign \g13541/_0_  = n22554 ;
  assign \g13542/_0_  = n22557 ;
  assign \g13543/_0_  = n22560 ;
  assign \g13544/_0_  = n22563 ;
  assign \g13545/_0_  = n22566 ;
  assign \g13546/_0_  = n22569 ;
  assign \g13547/_0_  = n22572 ;
  assign \g13548/_0_  = n22575 ;
  assign \g13549/_0_  = n22578 ;
  assign \g13550/_0_  = n22580 ;
  assign \g13551/_0_  = n22585 ;
  assign \g13552/_0_  = n22587 ;
  assign \g13553/_0_  = n22589 ;
  assign \g13554/_0_  = n22592 ;
  assign \g13555/_0_  = n22595 ;
  assign \g13556/_0_  = n22598 ;
  assign \g13557/_0_  = n22601 ;
  assign \g13558/_0_  = n22604 ;
  assign \g13559/_0_  = n22607 ;
  assign \g13560/_0_  = n22610 ;
  assign \g13561/_0_  = n22613 ;
  assign \g13562/_0_  = n22616 ;
  assign \g13563/_0_  = n22619 ;
  assign \g13564/_0_  = n22622 ;
  assign \g13565/_0_  = n22625 ;
  assign \g13566/_0_  = n22628 ;
  assign \g13567/_0_  = n22631 ;
  assign \g13568/_0_  = n22634 ;
  assign \g13569/_0_  = n22637 ;
  assign \g13570/_0_  = n22640 ;
  assign \g13571/_0_  = n22643 ;
  assign \g13572/_0_  = n22646 ;
  assign \g137/_3_  = ~n22680 ;
  assign \g1387/_3_  = ~n22690 ;
  assign \g1388/_3_  = n22696 ;
  assign \g1389/_0_  = ~n22701 ;
  assign \g139/_0_  = ~n22883 ;
  assign \g1390/_0_  = n22916 ;
  assign \g1393/_0_  = n22919 ;
  assign \g140/_0_  = ~n22926 ;
  assign \g141/_0_  = ~n22929 ;
  assign \g14173/_0_  = n22933 ;
  assign \g14176/_0_  = n22936 ;
  assign \g142/_3_  = ~n22961 ;
  assign \g14273/_1__syn_2  = n20402 ;
  assign \g14274/_0_  = n22962 ;
  assign \g14280/_0_  = n22973 ;
  assign \g14281/_0_  = n22984 ;
  assign \g143/_3_  = ~n23001 ;
  assign \g14354/_3__syn_2  = n13779 ;
  assign \g14370/_0_  = n23004 ;
  assign \g14385/_0_  = n23008 ;
  assign \g14386/_0_  = n23011 ;
  assign \g144/_3_  = n23017 ;
  assign \g14407/_0_  = n23023 ;
  assign \g14412/_0_  = n23026 ;
  assign \g14435/_0_  = n23035 ;
  assign \g14439/_0_  = n23037 ;
  assign \g145/_0_  = ~n23089 ;
  assign \g14522/_0_  = n23091 ;
  assign \g14528/_0_  = ~n23093 ;
  assign \g14533/_0_  = ~n23116 ;
  assign \g14581/_1_  = ~n23117 ;
  assign \g14582/_0_  = ~n23118 ;
  assign \g146/_3_  = n23124 ;
  assign \g14671/_0_  = n23135 ;
  assign \g14672/_0_  = n23146 ;
  assign \g147/_0_  = ~n23188 ;
  assign \g1473/_0_  = ~n23205 ;
  assign \g148/_0_  = ~n23222 ;
  assign \g14826/_0_  = n19024 ;
  assign \g149/_0_  = n23228 ;
  assign \g14908/_0_  = ~n23234 ;
  assign \g14911/_0_  = ~n23240 ;
  assign \g14936/_2_  = n23243 ;
  assign \g1494/_0_  = ~n23259 ;
  assign \g1495/_0_  = ~n23262 ;
  assign \g14950/_2_  = n23274 ;
  assign \g14953/_2_  = n23286 ;
  assign \g15003/_0_  = n23290 ;
  assign \g15004/_0_  = ~n23293 ;
  assign \g15006/_0_  = ~n23296 ;
  assign \g15007/_0_  = ~n23299 ;
  assign \g15008/_0_  = ~n23302 ;
  assign \g15009/_0_  = ~n23305 ;
  assign \g15010/_0_  = ~n23308 ;
  assign \g15011/_0_  = ~n23311 ;
  assign \g15012/_0_  = ~n23314 ;
  assign \g15013/_0_  = ~n23317 ;
  assign \g15014/_0_  = ~n23320 ;
  assign \g15015/_0_  = ~n23323 ;
  assign \g15016/_0_  = ~n23326 ;
  assign \g15017/_0_  = ~n23329 ;
  assign \g15018/_0_  = ~n23332 ;
  assign \g15019/_0_  = ~n23335 ;
  assign \g15035/_0_  = ~n23339 ;
  assign \g15036/_0_  = ~n23342 ;
  assign \g15038/_0_  = ~n23349 ;
  assign \g15039/_0_  = ~n23355 ;
  assign \g15040/_0_  = ~n23361 ;
  assign \g15041/_0_  = ~n23367 ;
  assign \g15042/_0_  = ~n23373 ;
  assign \g15043/_0_  = ~n23379 ;
  assign \g15044/_0_  = ~n23385 ;
  assign \g15045/_0_  = ~n23391 ;
  assign \g15046/_0_  = ~n23397 ;
  assign \g15056/_00_  = ~n23403 ;
  assign \g151/_0_  = ~n23406 ;
  assign \g15193/_0_  = ~n23413 ;
  assign \g152/_0_  = ~n23416 ;
  assign \g15256/_0_  = n23425 ;
  assign \g153/_0_  = ~n23428 ;
  assign \g15393/_0_  = ~n23436 ;
  assign \g15394/_0_  = ~n23442 ;
  assign \g15395/_0_  = ~n23448 ;
  assign \g15396/_0_  = ~n23454 ;
  assign \g15397/_0_  = ~n23460 ;
  assign \g15398/_0_  = ~n23466 ;
  assign \g15399/_0_  = ~n23472 ;
  assign \g154/_0_  = ~n23475 ;
  assign \g15400/_0_  = ~n23481 ;
  assign \g15401/_0_  = ~n23487 ;
  assign \g15402/_0_  = ~n23493 ;
  assign \g15403/_0_  = ~n23499 ;
  assign \g15404/_0_  = ~n23505 ;
  assign \g15405/_0_  = ~n23511 ;
  assign \g15406/_0_  = ~n23517 ;
  assign \g15407/_0_  = ~n23523 ;
  assign \g15408/_0_  = ~n23529 ;
  assign \g15473/_0_  = n23534 ;
  assign \g15650/_0_  = n23536 ;
  assign \g15651/_0_  = n23538 ;
  assign \g15652/_0_  = n23540 ;
  assign \g15653/_0_  = n23542 ;
  assign \g15662/_0_  = ~n23545 ;
  assign \g15663/_0_  = ~n23548 ;
  assign \g15664/_0_  = ~n23551 ;
  assign \g15665/_0_  = ~n23554 ;
  assign \g15666/_0_  = ~n23557 ;
  assign \g15667/_0_  = ~n23560 ;
  assign \g15668/_0_  = ~n23563 ;
  assign \g15669/_0_  = ~n23566 ;
  assign \g15670/_0_  = ~n23569 ;
  assign \g15671/_0_  = ~n23572 ;
  assign \g15672/_0_  = ~n23575 ;
  assign \g15673/_0_  = ~n23578 ;
  assign \g15674/_0_  = ~n23581 ;
  assign \g15675/_0_  = ~n23584 ;
  assign \g1569/_0_  = n23676 ;
  assign \g1570/_0_  = n23680 ;
  assign \g1575/_0_  = n23686 ;
  assign \g1576/_0_  = n23689 ;
  assign \g15922/_1_  = ~n23690 ;
  assign \g15970/_0_  = n23691 ;
  assign \g16059/_0_  = n23694 ;
  assign \g1606/_3_  = ~n23704 ;
  assign \g16124/_0_  = n20576 ;
  assign \g16144/_0_  = ~n23706 ;
  assign \g16202/_0_  = n23709 ;
  assign \g16214/_0_  = n23713 ;
  assign \g16247/_0_  = n23719 ;
  assign \g16257/_0_  = n23725 ;
  assign \g16274/_1_  = n23726 ;
  assign \g16324/_0_  = n20787 ;
  assign \g16343/_1__syn_2  = n22291 ;
  assign \g16381/_0_  = ~n23730 ;
  assign \g16383/_0_  = ~n23739 ;
  assign \g16386/_0_  = n23742 ;
  assign \g16414/_1__syn_2  = n21906 ;
  assign \g16416/_0__syn_2  = n20864 ;
  assign \g16448/_0_  = n23743 ;
  assign \g16460/_1_  = n23744 ;
  assign \g16625/_3_  = n23033 ;
  assign \g16662/_0_  = ~n23751 ;
  assign \g16668/_1__syn_2  = n22477 ;
  assign \g16692/_0_  = ~n23753 ;
  assign \g16721/_0_  = n23760 ;
  assign \g16723/_0_  = ~n23765 ;
  assign \g16725/_0_  = n23769 ;
  assign \g16726/_0_  = ~n23772 ;
  assign \g16727/_0_  = n23775 ;
  assign \g16728/_0_  = ~n23778 ;
  assign \g16729/_0_  = ~n23781 ;
  assign \g16730/_0_  = n23785 ;
  assign \g16731/_0_  = n23788 ;
  assign \g16732/_0_  = ~n23791 ;
  assign \g16733/_0_  = ~n23794 ;
  assign \g16734/_0_  = n23797 ;
  assign \g16735/_0_  = n23801 ;
  assign \g16736/_0_  = ~n23804 ;
  assign \g16737/_0_  = ~n23807 ;
  assign \g16738/_0_  = ~n23810 ;
  assign \g16739/_0_  = n23813 ;
  assign \g16740/_0_  = n23817 ;
  assign \g16741/_0_  = ~n23820 ;
  assign \g16742/_0_  = ~n23823 ;
  assign \g16743/_0_  = n23826 ;
  assign \g16747/_0_  = n23830 ;
  assign \g16748/_0_  = n23833 ;
  assign \g16749/_0_  = n23836 ;
  assign \g16750/_0_  = n23839 ;
  assign \g16753/_0_  = n23842 ;
  assign \g16754/_0_  = n23845 ;
  assign \g16755/_0_  = n23848 ;
  assign \g16756/_0_  = n23851 ;
  assign \g16757/_0_  = n23854 ;
  assign \g16758/_0_  = n23857 ;
  assign \g16761/_0_  = n23863 ;
  assign \g16765/_0_  = ~n23868 ;
  assign \g16766/_0_  = ~n23871 ;
  assign \g16767/_0_  = ~n23874 ;
  assign \g16768/_0_  = ~n23877 ;
  assign \g16769/_0_  = ~n23880 ;
  assign \g16772/_0_  = ~n23883 ;
  assign \g16785/_0_  = ~n23888 ;
  assign \g16786/_0_  = n23892 ;
  assign \g16787/_0_  = ~n23895 ;
  assign \g16788/_0_  = n23898 ;
  assign \g16789/_0_  = ~n23901 ;
  assign \g16790/_0_  = ~n23904 ;
  assign \g16791/_0_  = n23907 ;
  assign \g16804/_0_  = n23911 ;
  assign \g16805/_0_  = n23914 ;
  assign \g16806/_0_  = n23917 ;
  assign \g16807/_0_  = n23923 ;
  assign \g16808/_0_  = n23926 ;
  assign \g16809/_0_  = n23929 ;
  assign \g16810/_0_  = n23933 ;
  assign \g16811/_0_  = n23936 ;
  assign \g16812/_0_  = n23939 ;
  assign \g16813/_0_  = n23942 ;
  assign \g16814/_0_  = n23945 ;
  assign \g16815/_0_  = n23948 ;
  assign \g16816/_0_  = ~n23951 ;
  assign \g16817/_0_  = n23954 ;
  assign \g16819/_0_  = ~n23961 ;
  assign \g16822/_0_  = ~n23964 ;
  assign \g16823/_0_  = ~n23967 ;
  assign \g16824/_0_  = ~n23970 ;
  assign \g16825/_0_  = ~n23973 ;
  assign \g16828/_0_  = ~n23976 ;
  assign \g16829/_0_  = ~n23979 ;
  assign \g16830/_0_  = ~n23982 ;
  assign \g16831/_0_  = ~n23985 ;
  assign \g16832/_0_  = ~n23988 ;
  assign \g16833/_0_  = ~n23991 ;
  assign \g16834/_0_  = ~n23994 ;
  assign \g16835/_0_  = ~n23997 ;
  assign \g16836/_0_  = ~n24000 ;
  assign \g16837/_0_  = ~n24007 ;
  assign \g16840/_0_  = ~n24010 ;
  assign \g16841/_0_  = ~n24013 ;
  assign \g16842/_0_  = ~n24016 ;
  assign \g16843/_0_  = ~n24019 ;
  assign \g16846/_0_  = ~n24026 ;
  assign \g16847/_0_  = ~n24029 ;
  assign \g16848/_0_  = ~n24032 ;
  assign \g16849/_0_  = ~n24035 ;
  assign \g16850/_0_  = ~n24038 ;
  assign \g16851/_0_  = ~n24041 ;
  assign \g16852/_0_  = ~n24044 ;
  assign \g16853/_0_  = ~n24047 ;
  assign \g16854/_0_  = n24050 ;
  assign \g16855/_0_  = n24053 ;
  assign \g16856/_0_  = n24056 ;
  assign \g16857/_0_  = n24059 ;
  assign \g16859/_0_  = ~n24065 ;
  assign \g16862/_0_  = n24071 ;
  assign \g16865/_0_  = n24077 ;
  assign \g16866/_0_  = ~n24083 ;
  assign \g16867/_0_  = ~n24088 ;
  assign \g16868/_0_  = ~n24093 ;
  assign \g16869/_0_  = ~n24095 ;
  assign \g16870/_0_  = ~n24101 ;
  assign \g16871/_0_  = ~n24103 ;
  assign \g16872/_0_  = ~n24108 ;
  assign \g16873/_0_  = ~n24113 ;
  assign \g16874/_0_  = ~n24115 ;
  assign \g16875/_0_  = ~n24121 ;
  assign \g16876/_0_  = ~n24126 ;
  assign \g16877/_0_  = n24129 ;
  assign \g16878/_0_  = ~n24132 ;
  assign \g16879/_0_  = ~n24135 ;
  assign \g16880/_0_  = ~n24137 ;
  assign \g16881/_0_  = ~n24140 ;
  assign \g16882/_0_  = ~n24146 ;
  assign \g16884/_0_  = ~n24148 ;
  assign \g16887/_0_  = ~n24151 ;
  assign \g16891/_0_  = ~n24153 ;
  assign \g16892/_0_  = ~n24156 ;
  assign \g16893/_0_  = n24159 ;
  assign \g16894/_0_  = ~n24161 ;
  assign \g16895/_0_  = ~n24163 ;
  assign \g16897/_0_  = ~n24165 ;
  assign \g16898/_0_  = ~n24168 ;
  assign \g16899/_0_  = ~n24171 ;
  assign \g16900/_0_  = ~n24174 ;
  assign \g16901/_0_  = ~n24176 ;
  assign \g16902/_0_  = ~n24178 ;
  assign \g16903/_0_  = ~n24180 ;
  assign \g16904/_0_  = ~n24183 ;
  assign \g16905/_0_  = ~n24185 ;
  assign \g16906/_0_  = ~n24187 ;
  assign \g16907/_0_  = ~n24189 ;
  assign \g16908/_0_  = ~n24192 ;
  assign \g16909/_0_  = ~n24195 ;
  assign \g16910/_0_  = ~n24197 ;
  assign \g16912/_0_  = n24200 ;
  assign \g16914/_0_  = n24203 ;
  assign \g16915/_0_  = n24206 ;
  assign \g16950/_0_  = ~n24209 ;
  assign \g16951/_0_  = ~n24212 ;
  assign \g16952/_0_  = ~n24215 ;
  assign \g16953/_0_  = ~n24218 ;
  assign \g16954/_0_  = ~n24221 ;
  assign \g16955/_0_  = ~n24224 ;
  assign \g16956/_0_  = ~n24227 ;
  assign \g16957/_0_  = ~n24230 ;
  assign \g16958/_0_  = ~n24233 ;
  assign \g16959/_0_  = ~n24236 ;
  assign \g16960/_0_  = ~n24239 ;
  assign \g16961/_0_  = ~n24242 ;
  assign \g16962/_0_  = ~n24245 ;
  assign \g16963/_0_  = ~n24248 ;
  assign \g16964/_0_  = ~n24251 ;
  assign \g16965/_0_  = ~n24254 ;
  assign \g16966/_0_  = ~n24257 ;
  assign \g16967/_0_  = ~n24260 ;
  assign \g16968/_0_  = ~n24263 ;
  assign \g16970/_0_  = ~n24266 ;
  assign \g17102/_3_  = n24270 ;
  assign \g17106/_0_  = ~n24275 ;
  assign \g17107/_0_  = n24278 ;
  assign \g17109/_0_  = ~n24281 ;
  assign \g17110/_0_  = ~n24284 ;
  assign \g17111/_0_  = ~n24287 ;
  assign \g17112/_0_  = ~n24290 ;
  assign \g17115/_0_  = ~n24293 ;
  assign \g17116/_0_  = ~n24296 ;
  assign \g17119/_0_  = ~n24299 ;
  assign \g17120/_0_  = ~n24302 ;
  assign \g17122/_0_  = ~n24305 ;
  assign \g17123/_0_  = ~n24308 ;
  assign \g17124/_0_  = ~n24311 ;
  assign \g17125/_0_  = ~n24314 ;
  assign \g17126/_0_  = ~n24317 ;
  assign \g17127/_0_  = ~n24320 ;
  assign \g17128/_0_  = ~n24323 ;
  assign \g17130/_0_  = ~n24326 ;
  assign \g17131/_0_  = ~n24329 ;
  assign \g17132/_0_  = ~n24332 ;
  assign \g17133/_0_  = ~n24335 ;
  assign \g17134/_0_  = ~n24338 ;
  assign \g17135/_0_  = ~n24341 ;
  assign \g17136/_0_  = ~n24344 ;
  assign \g17137/_0_  = ~n24347 ;
  assign \g17138/_0_  = ~n24350 ;
  assign \g17140/_0_  = ~n24353 ;
  assign \g17141/_0_  = ~n24356 ;
  assign \g17142/_0_  = ~n24359 ;
  assign \g17143/_0_  = ~n24362 ;
  assign \g17144/_0_  = ~n24365 ;
  assign \g17145/_0_  = ~n24368 ;
  assign \g17146/_0_  = ~n24371 ;
  assign \g17147/_0_  = ~n24374 ;
  assign \g17148/_0_  = ~n24377 ;
  assign \g17149/_0_  = ~n24380 ;
  assign \g17150/_0_  = ~n24383 ;
  assign \g17151/_0_  = ~n24386 ;
  assign \g17152/_0_  = ~n24389 ;
  assign \g17153/_0_  = ~n24392 ;
  assign \g17154/_0_  = ~n24395 ;
  assign \g17155/_0_  = n24398 ;
  assign \g17157/_0_  = n24401 ;
  assign \g17159/_0_  = n24409 ;
  assign \g17160/_0_  = n24412 ;
  assign \g17161/_0_  = n24415 ;
  assign \g17162/_0_  = n24418 ;
  assign \g17163/_0_  = n24425 ;
  assign \g17164/_0_  = n24428 ;
  assign \g17165/_0_  = n24431 ;
  assign \g17166/_0_  = n24434 ;
  assign \g17168/_0_  = ~n24437 ;
  assign \g17171/_0_  = ~n24440 ;
  assign \g17173/_0_  = n24445 ;
  assign \g17177/_0_  = n24448 ;
  assign \g17178/_0_  = ~n24451 ;
  assign \g17179/_0_  = ~n24454 ;
  assign \g17180/_0_  = ~n24457 ;
  assign \g17182/_0_  = n24460 ;
  assign \g17183/_0_  = n24463 ;
  assign \g17184/_0_  = n24466 ;
  assign \g17185/_0_  = n24469 ;
  assign \g17186/_0_  = n24472 ;
  assign \g17188/_0_  = n24475 ;
  assign \g17189/_0_  = n24478 ;
  assign \g17190/_0_  = n24481 ;
  assign \g17191/_0_  = n24484 ;
  assign \g17193/_0_  = n24487 ;
  assign \g17194/_0_  = n24490 ;
  assign \g17195/_0_  = n24493 ;
  assign \g17196/_0_  = n24496 ;
  assign \g17197/_0_  = n24499 ;
  assign \g17198/_0_  = n24502 ;
  assign \g17199/_0_  = n24505 ;
  assign \g17200/_0_  = n24508 ;
  assign \g17201/_0_  = n24511 ;
  assign \g17202/_0_  = n24514 ;
  assign \g17203/_0_  = n24520 ;
  assign \g17204/_0_  = n24523 ;
  assign \g17205/_0_  = n24526 ;
  assign \g17206/_0_  = n24529 ;
  assign \g17207/_0_  = n24532 ;
  assign \g17208/_0_  = ~n24535 ;
  assign \g17209/_0_  = n24538 ;
  assign \g17210/_0_  = n24541 ;
  assign \g17211/_0_  = ~n24544 ;
  assign \g17212/_0_  = n24547 ;
  assign \g17213/_0_  = n24550 ;
  assign \g17214/_0_  = n24553 ;
  assign \g17215/_0_  = n24556 ;
  assign \g17216/_0_  = n24559 ;
  assign \g17217/_0_  = n24562 ;
  assign \g17218/_0_  = n24565 ;
  assign \g17219/_0_  = n24568 ;
  assign \g17223/_0_  = n24571 ;
  assign \g17224/_0_  = n24574 ;
  assign \g17225/_0_  = n24577 ;
  assign \g17226/_0_  = n24580 ;
  assign \g17227/_0_  = n24583 ;
  assign \g17228/_0_  = n24586 ;
  assign \g17229/_0_  = ~n24589 ;
  assign \g17231/_0_  = ~n24592 ;
  assign \g17232/_0_  = ~n24595 ;
  assign \g17233/_0_  = n24597 ;
  assign \g17234/_0_  = ~n24600 ;
  assign \g17237/_0_  = ~n24603 ;
  assign \g17239/_0_  = ~n24606 ;
  assign \g17240/_0_  = n24609 ;
  assign \g17243/_0_  = ~n24612 ;
  assign \g17246/_0_  = ~n24615 ;
  assign \g17247/_0_  = ~n24618 ;
  assign \g17248/_0_  = ~n24621 ;
  assign \g17249/_0_  = ~n24624 ;
  assign \g17250/_0_  = ~n24627 ;
  assign \g17251/_0_  = n24630 ;
  assign \g17252/_0_  = n24633 ;
  assign \g17253/_0_  = ~n24636 ;
  assign \g17254/_0_  = n24639 ;
  assign \g17258/_0_  = ~n24642 ;
  assign \g17261/_0_  = ~n24651 ;
  assign \g17262/_0_  = ~n24654 ;
  assign \g17269/_0_  = n24657 ;
  assign \g17271/_0_  = ~n24660 ;
  assign \g17274/_0_  = ~n24663 ;
  assign \g17275/_0_  = ~n24666 ;
  assign \g17276/_0_  = ~n24669 ;
  assign \g17277/_0_  = ~n24672 ;
  assign \g17278/_0_  = ~n24675 ;
  assign \g17279/_0_  = ~n24678 ;
  assign \g17280/_0_  = ~n24681 ;
  assign \g17281/_0_  = ~n24684 ;
  assign \g17282/_0_  = ~n24687 ;
  assign \g17283/_0_  = ~n24690 ;
  assign \g17285/_0_  = ~n24693 ;
  assign \g17290/_0_  = n24696 ;
  assign \g17292/_0_  = ~n24699 ;
  assign \g17293/_0_  = ~n24702 ;
  assign \g17296/_0_  = n24705 ;
  assign \g17297/_0_  = n24708 ;
  assign \g17298/_0_  = ~n24710 ;
  assign \g173/_0_  = n24721 ;
  assign \g17303/_0_  = n24724 ;
  assign \g17304/_0_  = n24727 ;
  assign \g17305/_0_  = n24730 ;
  assign \g17306/_0_  = n24733 ;
  assign \g17307/_0_  = n24736 ;
  assign \g17308/_0_  = n24739 ;
  assign \g17309/_0_  = n24742 ;
  assign \g17310/_0_  = n24745 ;
  assign \g17311/_0_  = n24748 ;
  assign \g17312/_0_  = n24751 ;
  assign \g17314/_0_  = n24754 ;
  assign \g17315/_0_  = n24757 ;
  assign \g17316/_0_  = n24760 ;
  assign \g17317/_0_  = n24763 ;
  assign \g17318/_0_  = n24766 ;
  assign \g17319/_0_  = n24769 ;
  assign \g17320/_0_  = n24772 ;
  assign \g17321/_0_  = n24775 ;
  assign \g17322/_0_  = n24778 ;
  assign \g17323/_0_  = n24781 ;
  assign \g17324/_0_  = n24784 ;
  assign \g17325/_0_  = n24787 ;
  assign \g17326/_0_  = n24790 ;
  assign \g17327/_0_  = n24793 ;
  assign \g17328/_0_  = n24796 ;
  assign \g17329/_0_  = n24799 ;
  assign \g17330/_0_  = n24802 ;
  assign \g17331/_0_  = n24805 ;
  assign \g17332/_0_  = n24808 ;
  assign \g17333/_0_  = n24811 ;
  assign \g17335/_0_  = n24814 ;
  assign \g17336/_0_  = ~n24818 ;
  assign \g17337/_0_  = n24821 ;
  assign \g17338/_0_  = ~n24824 ;
  assign \g17339/_0_  = n24827 ;
  assign \g17340/_0_  = ~n24830 ;
  assign \g17342/_0_  = n24833 ;
  assign \g17343/_0_  = ~n24836 ;
  assign \g17347/_0_  = n24839 ;
  assign \g17350/_0_  = n24842 ;
  assign \g17354/_0_  = n24845 ;
  assign \g17356/_0_  = n24848 ;
  assign \g17357/_0_  = n24851 ;
  assign \g17358/_0_  = n24854 ;
  assign \g17359/_0_  = n24857 ;
  assign \g17360/_0_  = n24860 ;
  assign \g17415/_0_  = ~n24863 ;
  assign \g17441/_0_  = n24865 ;
  assign \g17442/_0_  = ~n24867 ;
  assign \g17451/_0_  = n24869 ;
  assign \g17457/_0_  = n24873 ;
  assign \g17458/_0_  = ~n24876 ;
  assign \g17459/_0_  = n24879 ;
  assign \g17460/_0_  = n24882 ;
  assign \g17461/_0_  = n24885 ;
  assign \g17462/_0_  = n24888 ;
  assign \g17463/_0_  = n24891 ;
  assign \g17464/_0_  = n24894 ;
  assign \g17465/_0_  = n24897 ;
  assign \g17466/_0_  = n24900 ;
  assign \g17467/_0_  = n24903 ;
  assign \g17468/_0_  = n24906 ;
  assign \g17469/_0_  = ~n24909 ;
  assign \g17470/_0_  = ~n24912 ;
  assign \g17471/_0_  = n24915 ;
  assign \g17472/_0_  = n24918 ;
  assign \g175/_3_  = ~n24931 ;
  assign \g1750/_0_  = ~n24946 ;
  assign \g176/_3_  = ~n24965 ;
  assign \g17619/_0_  = n24967 ;
  assign \g17620/_0_  = ~n24968 ;
  assign \g1763/_3_  = ~n24978 ;
  assign \g1764/_3_  = n24984 ;
  assign \g1768/_0_  = ~n24990 ;
  assign \g1769/_0_  = ~n24993 ;
  assign \g177/_3_  = ~n25006 ;
  assign \g17737/_0_  = ~n25009 ;
  assign \g17747/_0_  = n25013 ;
  assign \g178/_3_  = n25019 ;
  assign \g17814/_1_  = n21314 ;
  assign \g17815/_0_  = ~n25023 ;
  assign \g17821/_1_  = ~n25024 ;
  assign \g17821/_1__syn_2  = n25024 ;
  assign \g17872/_0_  = n25026 ;
  assign \g179/_3_  = n25032 ;
  assign \g17902/_0_  = n25035 ;
  assign \g180/_3_  = n25041 ;
  assign \g18020/_1_  = ~n25043 ;
  assign \g18057/_0_  = ~n25045 ;
  assign \g18096/_0_  = n25049 ;
  assign \g18099/_0_  = n25052 ;
  assign \g18107/_0_  = n25055 ;
  assign \g18133/_0_  = ~n25059 ;
  assign \g18140/_1_  = ~n23021 ;
  assign \g18153/_0_  = n25062 ;
  assign \g182/_0_  = ~n25069 ;
  assign \g18218/_0_  = ~n25073 ;
  assign \g18244/_0_  = n25075 ;
  assign \g18262/_0_  = n25079 ;
  assign \g18267/_0_  = n25082 ;
  assign \g18387/_1__syn_2  = n25085 ;
  assign \g184/_0_  = n25088 ;
  assign \g18478/_1_  = n23343 ;
  assign \g18585/_3_  = n22290 ;
  assign \g18608/_0_  = ~n25092 ;
  assign \g18609/_0_  = ~n25096 ;
  assign \g18613/_0_  = ~n25101 ;
  assign \g18618/_0_  = ~n25105 ;
  assign \g18647/_0_  = ~n25109 ;
  assign \g18687/_2_  = n20990 ;
  assign \g18707/_0_  = ~n25113 ;
  assign \g18748/_0_  = n25117 ;
  assign \g18753/_0_  = n25121 ;
  assign \g18758/_0_  = n25124 ;
  assign \g18759/_0_  = n25128 ;
  assign \g18760/_0_  = n25131 ;
  assign \g18761/_0_  = n25135 ;
  assign \g18762/_0_  = n25138 ;
  assign \g18763/_0_  = n25141 ;
  assign \g18764/_0_  = n25144 ;
  assign \g18765/_0_  = n25147 ;
  assign \g18766/_0_  = n25150 ;
  assign \g18767/_0_  = n25153 ;
  assign \g18768/_0_  = n25156 ;
  assign \g18770/_0_  = n25159 ;
  assign \g18771/_0_  = n25162 ;
  assign \g18788/_0_  = n25165 ;
  assign \g18796/_0_  = n25168 ;
  assign \g18800/_0_  = n25171 ;
  assign \g18801/_0_  = n25174 ;
  assign \g18802/_0_  = n25177 ;
  assign \g18803/_0_  = n25180 ;
  assign \g18804/_0_  = n25183 ;
  assign \g18805/_0_  = n25186 ;
  assign \g18807/_0_  = n25189 ;
  assign \g18840/_0_  = ~n25196 ;
  assign \g18843/_0_  = n25199 ;
  assign \g18844/_0_  = ~n25205 ;
  assign \g18846/_0_  = ~n25210 ;
  assign \g18847/_0_  = ~n25216 ;
  assign \g18848/_0_  = ~n25220 ;
  assign \g18849/_0_  = ~n25224 ;
  assign \g18850/_0_  = n25228 ;
  assign \g18851/_0_  = n25231 ;
  assign \g18852/_0_  = n25234 ;
  assign \g18853/_0_  = n25237 ;
  assign \g18854/_0_  = ~n25243 ;
  assign \g18855/_0_  = ~n25247 ;
  assign \g18856/_0_  = ~n20720 ;
  assign \g18858/_0_  = ~n20709 ;
  assign \g18860/_0_  = ~n25251 ;
  assign \g18861/_0_  = n25254 ;
  assign \g18863/_0_  = n25257 ;
  assign \g18864/_0_  = n25260 ;
  assign \g18866/_0_  = n25263 ;
  assign \g18867/_0_  = n25266 ;
  assign \g18868/_0_  = n25269 ;
  assign \g18869/_0_  = n25272 ;
  assign \g18870/_0_  = n25275 ;
  assign \g18871/_0_  = n25278 ;
  assign \g18872/_0_  = n25281 ;
  assign \g18873/_0_  = n25284 ;
  assign \g18874/_0_  = n25287 ;
  assign \g18875/_0_  = n25290 ;
  assign \g18876/_0_  = n25293 ;
  assign \g18877/_0_  = n25296 ;
  assign \g18878/_0_  = n25299 ;
  assign \g18879/_0_  = n25302 ;
  assign \g18880/_0_  = n25305 ;
  assign \g18881/_0_  = n25308 ;
  assign \g18882/_0_  = n25311 ;
  assign \g18883/_0_  = n25314 ;
  assign \g18888/_0_  = ~n25318 ;
  assign \g18892/_0_  = ~n25324 ;
  assign \g18895/_0_  = ~n25330 ;
  assign \g18896/_0_  = ~n25336 ;
  assign \g18897/_0_  = n25339 ;
  assign \g18905/_0_  = ~n25343 ;
  assign \g18908/_0_  = n25346 ;
  assign \g18909/_0_  = n25349 ;
  assign \g18912/_0_  = n25352 ;
  assign \g18918/_0_  = ~n25356 ;
  assign \g18919/_0_  = ~n25360 ;
  assign \g18920/_0_  = n25363 ;
  assign \g18921/_0_  = ~n25369 ;
  assign \g18922/_0_  = n25372 ;
  assign \g18924/_0_  = ~n25378 ;
  assign \g18925/_0_  = n25381 ;
  assign \g18927/_0_  = n25384 ;
  assign \g18930/_0_  = n25387 ;
  assign \g18966/_0_  = ~n25393 ;
  assign \g18968/_0_  = ~n25399 ;
  assign \g18970/_0_  = n25402 ;
  assign \g18974/_0_  = n25405 ;
  assign \g18975/_0_  = ~n25411 ;
  assign \g18977/_0_  = ~n25417 ;
  assign \g18981/_0_  = ~n20757 ;
  assign \g18983/_0_  = ~n20604 ;
  assign \g18985/_0_  = ~n20616 ;
  assign \g18987/_0_  = ~n20626 ;
  assign \g18989/_0_  = ~n20636 ;
  assign \g18991/_0_  = ~n25421 ;
  assign \g18992/_0_  = ~n25427 ;
  assign \g18993/_0_  = ~n25433 ;
  assign \g18994/_0_  = n25436 ;
  assign \g18995/_0_  = ~n25442 ;
  assign \g18996/_0_  = n25445 ;
  assign \g18997/_0_  = ~n25451 ;
  assign \g18998/_0_  = n25454 ;
  assign \g18999/_0_  = n25457 ;
  assign \g19001/_0_  = n25460 ;
  assign \g19003/_0_  = n25463 ;
  assign \g19005/_0_  = n25466 ;
  assign \g19006/_0_  = ~n25472 ;
  assign \g19014/_0_  = ~n20646 ;
  assign \g19016/_0_  = ~n20654 ;
  assign \g19018/_0_  = ~n20665 ;
  assign \g19020/_0_  = ~n20676 ;
  assign \g19022/_0_  = ~n20731 ;
  assign \g19056/_3_  = ~n25476 ;
  assign \g19058/_3_  = ~n25480 ;
  assign \g19060/_3_  = ~n25484 ;
  assign \g19062/_3_  = ~n25488 ;
  assign \g1910/_0_  = ~n25502 ;
  assign \g19186/_0_  = n21380 ;
  assign \g19188/_0_  = n21388 ;
  assign \g19235/_0_  = n25506 ;
  assign \g19239/_0_  = n25509 ;
  assign \g19244/_0_  = n25512 ;
  assign \g19253/_0_  = n25515 ;
  assign \g19254/_0_  = n25518 ;
  assign \g19259/_0_  = n25521 ;
  assign \g19261/_0_  = n25524 ;
  assign \g19267/_0_  = n25527 ;
  assign \g19277/_0_  = n25531 ;
  assign \g19278/_0_  = n25534 ;
  assign \g19280/_0_  = n25538 ;
  assign \g19281/_0_  = n25541 ;
  assign \g19282/_0_  = n25544 ;
  assign \g19283/_0_  = n25547 ;
  assign \g19284/_0_  = n25550 ;
  assign \g19285/_0_  = n25553 ;
  assign \g19286/_0_  = n25556 ;
  assign \g19287/_0_  = n25559 ;
  assign \g19288/_0_  = n25562 ;
  assign \g19289/_0_  = n25565 ;
  assign \g19290/_0_  = n25568 ;
  assign \g19291/_0_  = n25571 ;
  assign \g19292/_0_  = n25574 ;
  assign \g19293/_0_  = n25577 ;
  assign \g19294/_0_  = n25580 ;
  assign \g19295/_0_  = n25583 ;
  assign \g19296/_0_  = n25586 ;
  assign \g19297/_0_  = n25589 ;
  assign \g19298/_0_  = n25592 ;
  assign \g19299/_0_  = n25595 ;
  assign \g19300/_0_  = n25598 ;
  assign \g19301/_0_  = n25601 ;
  assign \g19302/_0_  = n25604 ;
  assign \g19303/_0_  = n25607 ;
  assign \g19304/_0_  = n25610 ;
  assign \g19305/_0_  = n25613 ;
  assign \g19306/_0_  = n25616 ;
  assign \g19307/_0_  = n25619 ;
  assign \g19308/_0_  = n25622 ;
  assign \g19315/_0_  = n25625 ;
  assign \g19316/_0_  = n25628 ;
  assign \g19317/_0_  = n25631 ;
  assign \g19318/_0_  = n25634 ;
  assign \g19319/_0_  = n25637 ;
  assign \g19320/_0_  = n25640 ;
  assign \g19321/_0_  = n25643 ;
  assign \g19322/_0_  = n25646 ;
  assign \g19323/_0_  = n25649 ;
  assign \g19325/_3_  = ~n25654 ;
  assign \g19326/_3_  = ~n25659 ;
  assign \g19333/_3_  = ~n25664 ;
  assign \g19341/_3_  = ~n25669 ;
  assign \g19347/_3_  = ~n25674 ;
  assign \g19377/_3_  = ~n25677 ;
  assign \g19381/_3_  = ~n25682 ;
  assign \g19393/_0_  = ~n25687 ;
  assign \g19401/_0_  = ~n25693 ;
  assign \g19402/_0_  = ~n25699 ;
  assign \g195/_2_  = ~n13516 ;
  assign \g19513/_0_  = n25700 ;
  assign \g19514/_0_  = n25701 ;
  assign \g19515/_0_  = n25702 ;
  assign \g19516/_0_  = n25703 ;
  assign \g1952/_3_  = ~n25711 ;
  assign \g19529/_0_  = n25712 ;
  assign \g19530/_0_  = n25713 ;
  assign \g19531/_0_  = n25714 ;
  assign \g19532/_0_  = n25715 ;
  assign \g19533/_0_  = n25716 ;
  assign \g19534/_0_  = n25717 ;
  assign \g19535/_0_  = n25718 ;
  assign \g19536/_0_  = n25719 ;
  assign \g19537/_0_  = n25720 ;
  assign \g19539/_0_  = n25721 ;
  assign \g19546/_0_  = n25722 ;
  assign \g19552/_0_  = n25723 ;
  assign \g19553/_0_  = n25724 ;
  assign \g19562/_0_  = n25728 ;
  assign \g19563/_0_  = n25732 ;
  assign \g19564/_0_  = n25736 ;
  assign \g19572/_0_  = ~n19702 ;
  assign \g19575/_0_  = n25737 ;
  assign \g19615/_0_  = n25738 ;
  assign \g19686/_0_  = ~n25739 ;
  assign \g19688/_0_  = ~n25740 ;
  assign \g197/_0_  = n25792 ;
  assign \g19729/_0_  = n25796 ;
  assign \g19774/_0_  = n25800 ;
  assign \g19777/_0_  = n25804 ;
  assign \g19791/_0_  = n25808 ;
  assign \g19818/_0_  = n25810 ;
  assign \g19819/_0_  = n25811 ;
  assign \g19828/_0_  = n25815 ;
  assign \g19852/_1_  = ~n6067 ;
  assign \g19860/_0_  = n25819 ;
  assign \g19861/_0_  = n25823 ;
  assign \g19864/_0_  = n25827 ;
  assign \g19886/_0_  = n25828 ;
  assign \g19887/_0_  = n25830 ;
  assign \g199/_0_  = ~n25849 ;
  assign \g19908/_0_  = ~n25850 ;
  assign \g19918/_0_  = n25854 ;
  assign \g19927/_0_  = n25858 ;
  assign \g19933/_0_  = n25862 ;
  assign \g200/_0_  = n22959 ;
  assign \g20019/_0_  = n25866 ;
  assign \g20046/_0_  = n25870 ;
  assign \g20068/_1_  = n23958 ;
  assign \g20080/_1_  = n24004 ;
  assign \g201/_0_  = ~n25900 ;
  assign \g20137/_0_  = n25904 ;
  assign \g20139/_0_  = ~n25909 ;
  assign \g20141/_0_  = n25913 ;
  assign \g20152/_1_  = ~n6075 ;
  assign \g20154/_00_  = n25918 ;
  assign \g202/_0_  = ~n25948 ;
  assign \g20206/_0_  = ~n25953 ;
  assign \g20211/_2_  = n25954 ;
  assign \g20217/_2_  = n25955 ;
  assign \g20239/_0_  = ~n25958 ;
  assign \g20265/_2_  = n25959 ;
  assign \g20266/_0_  = ~n25961 ;
  assign \g20272/_2_  = ~n25964 ;
  assign \g20278/_2_  = n25965 ;
  assign \g20283/_0_  = ~n18519 ;
  assign \g20285/_2_  = ~n25968 ;
  assign \g20288/_2__syn_2  = n23336 ;
  assign \g20293/_0_  = ~n25972 ;
  assign \g20295/_2_  = ~n20870 ;
  assign \g203/_0_  = ~n22999 ;
  assign \g20302/_2_  = n25973 ;
  assign \g20303/_2_  = n25974 ;
  assign \g20304/_2_  = n25975 ;
  assign \g20311/_2_  = n25976 ;
  assign \g20326/_0_  = ~n25980 ;
  assign \g20330/_0_  = ~n25982 ;
  assign \g2034/_0_  = ~n25988 ;
  assign \g20345/_0_  = n25992 ;
  assign \g20346/_0_  = n25995 ;
  assign \g2035/_0_  = ~n25998 ;
  assign \g20363/_0_  = ~n21241 ;
  assign \g20364/_0_  = ~n26002 ;
  assign \g204/_0_  = ~n26021 ;
  assign \g2047/_0_  = ~n26026 ;
  assign \g20483/_0_  = ~n26029 ;
  assign \g20493/_00_  = ~n26034 ;
  assign \g205/_0_  = n26040 ;
  assign \g20569/_0_  = n26042 ;
  assign \g20570/_0_  = n26044 ;
  assign \g20571/_0_  = n26046 ;
  assign \g206/_0_  = ~n26049 ;
  assign \g20613/_0_  = n26050 ;
  assign \g20615/_0_  = n26051 ;
  assign \g20657/_1__syn_2  = n26052 ;
  assign \g20660/_0_  = n26053 ;
  assign \g20685/_0_  = n26055 ;
  assign \g207/_0_  = ~n26058 ;
  assign \g20713/_1_  = n26059 ;
  assign \g20747/_1_  = n26060 ;
  assign \g20784/_0_  = ~n23018 ;
  assign \g20820/_1_  = n25042 ;
  assign \g20859/_0_  = n26063 ;
  assign \g20873/_2_  = n26065 ;
  assign \g20886/_0_  = n26066 ;
  assign \g20887/_0_  = n26067 ;
  assign \g20891/_2__syn_2  = ~n25666 ;
  assign \g20907/_2_  = n25071 ;
  assign \g20936/_2__syn_2  = ~n25661 ;
  assign \g20937/_1_  = ~n26068 ;
  assign \g20955/_0_  = n26070 ;
  assign \g20959/_2__syn_2  = ~n25656 ;
  assign \g20967/_0_  = n26071 ;
  assign \g20971/_2__syn_2  = ~n25679 ;
  assign \g20974/_1__syn_2  = n25684 ;
  assign \g21015/_1_  = ~n26073 ;
  assign \g21051/_2_  = n25057 ;
  assign \g21079/_1_  = n26074 ;
  assign \g21081/_1_  = n26075 ;
  assign \g21087/_2__syn_2  = ~n25671 ;
  assign \g21114/_1_  = n26076 ;
  assign \g21116/_1_  = n26077 ;
  assign \g21120/_2__syn_2  = ~n25651 ;
  assign \g21147/_0_  = n26078 ;
  assign \g21179/_1_  = n26079 ;
  assign \g21185/_1_  = n26080 ;
  assign \g21223/_0_  = n26082 ;
  assign \g21242/_0_  = n26084 ;
  assign \g21253/_0_  = ~n26085 ;
  assign \g21257/_0_  = ~n26087 ;
  assign \g21323/_1_  = n26089 ;
  assign \g21324/_1_  = n26090 ;
  assign \g21366/_0_  = ~n26092 ;
  assign \g21385/_2_  = ~n26094 ;
  assign \g21464/_0_  = n26096 ;
  assign \g21475/_3_  = ~n26099 ;
  assign \g21481/_0_  = ~n26102 ;
  assign \g21482/_0_  = ~n26104 ;
  assign \g21494/_3_  = ~n26107 ;
  assign \g21500/_3_  = ~n26110 ;
  assign \g21507/_3_  = ~n26113 ;
  assign \g21511/_3_  = ~n26116 ;
  assign \g21537/_1_  = n26119 ;
  assign \g21568/_0_  = ~n26122 ;
  assign \g21591/_0_  = ~n26125 ;
  assign \g21604/_0_  = ~n26129 ;
  assign \g21605/_3_  = n20602 ;
  assign \g21606/_0_  = ~n26132 ;
  assign \g21607/_0_  = ~n26135 ;
  assign \g21608/_0_  = ~n26138 ;
  assign \g21609/_0_  = ~n26141 ;
  assign \g21610/_0_  = ~n26144 ;
  assign \g21611/_0_  = ~n26147 ;
  assign \g21612/_0_  = ~n26150 ;
  assign \g21613/_0_  = ~n26153 ;
  assign \g21614/_0_  = ~n26156 ;
  assign \g21615/_0_  = ~n26159 ;
  assign \g21616/_0_  = ~n26162 ;
  assign \g21617/_0_  = ~n26165 ;
  assign \g21618/_0_  = ~n26168 ;
  assign \g21621/_0_  = ~n26170 ;
  assign \g21640/_0_  = ~n26173 ;
  assign \g21678/_0_  = ~n26176 ;
  assign \g21679/_0_  = ~n26179 ;
  assign \g21686/_0_  = ~n26182 ;
  assign \g21692/_3_  = ~n24098 ;
  assign \g21696/_0_  = ~n26185 ;
  assign \g21698/_0_  = ~n26188 ;
  assign \g21702/_3_  = n20718 ;
  assign \g21707/_0_  = ~n26191 ;
  assign \g21709/_0_  = ~n26194 ;
  assign \g21728/_0_  = ~n26197 ;
  assign \g21729/_0_  = ~n26200 ;
  assign \g21731/_0_  = ~n26203 ;
  assign \g21732/_0_  = ~n26206 ;
  assign \g21733/_0_  = ~n26209 ;
  assign \g21736/_0_  = ~n26212 ;
  assign \g21744/_3_  = ~n20707 ;
  assign \g21753/_0_  = ~n26215 ;
  assign \g21754/_0_  = ~n26218 ;
  assign \g21755/_0_  = ~n26221 ;
  assign \g21756/_0_  = ~n26224 ;
  assign \g21757/_0_  = ~n26227 ;
  assign \g21759/_0_  = ~n26230 ;
  assign \g21761/_0_  = ~n26233 ;
  assign \g21763/_0_  = ~n26236 ;
  assign \g21764/_0_  = ~n26239 ;
  assign \g21766/_0_  = ~n26242 ;
  assign \g2180/_0_  = ~n26259 ;
  assign \g21853/_3_  = n23886 ;
  assign \g21861/_3_  = ~n24111 ;
  assign \g21863/_3_  = ~n24118 ;
  assign \g21869/_3_  = n20614 ;
  assign \g2187/_0_  = n26281 ;
  assign \g21875/_3_  = ~n24124 ;
  assign \g21877/_3_  = ~n24143 ;
  assign \g21879/_3_  = ~n24106 ;
  assign \g2188/_0_  = n26284 ;
  assign \g21900/_0_  = ~n26286 ;
  assign \g22080/_0_  = n26287 ;
  assign \g22082/_0_  = n26288 ;
  assign \g22135/_0_  = n26289 ;
  assign \g22145/_1_  = n26290 ;
  assign \g22225/_0_  = n26291 ;
  assign \g223/_0_  = n25004 ;
  assign \g22354/_0_  = ~n26292 ;
  assign \g224/_0_  = ~n24929 ;
  assign \g22412/_0_  = n26302 ;
  assign \g22415/_1__syn_2  = ~n23020 ;
  assign \g225/_0_  = ~n24963 ;
  assign \g2257/_0_  = ~n5560 ;
  assign \g226/_3_  = ~n26319 ;
  assign \g22624/_0_  = ~n26320 ;
  assign \g227/_3_  = n26326 ;
  assign \g22702/_0_  = n26327 ;
  assign \g22919/_1__syn_2  = n25989 ;
  assign \g22933/_0_  = n26334 ;
  assign \g22954/_0_  = n26337 ;
  assign \g22989/_1_  = ~n26338 ;
  assign \g23529/_0_  = ~\T_IRQE1n_pad  ;
  assign \g23539/_0_  = ~\T_IRQ2n_pad  ;
  assign \g2362/_2_  = n26396 ;
  assign \g23766/_0_  = ~T_PWDn_pad ;
  assign \g24/_3_  = ~n26399 ;
  assign \g24018/_0_  = ~\T_IRQ0n_pad  ;
  assign \g2416/_0_  = n26962 ;
  assign \g2420/_0_  = ~n26966 ;
  assign \g24213/_0_  = ~\T_IRQL1n_pad  ;
  assign \g24301/_0_  = ~\T_IRQ1n_pad  ;
  assign \g2479/_0_  = ~n27036 ;
  assign \g248/_3_  = ~n27055 ;
  assign \g2480/_0_  = ~n27083 ;
  assign \g2481/_0_  = ~n27111 ;
  assign \g2482/_0_  = ~n27139 ;
  assign \g2483/_0_  = ~n27167 ;
  assign \g2484/_0_  = ~n27195 ;
  assign \g2485/_0_  = ~n27223 ;
  assign \g2486/_0_  = ~n27251 ;
  assign \g2487/_0_  = ~n27279 ;
  assign \g2488/_0_  = ~n27307 ;
  assign \g249/_3_  = n27313 ;
  assign \g2490/_0_  = ~n27341 ;
  assign \g2491/_0_  = ~n27369 ;
  assign \g2492/_0_  = ~n27397 ;
  assign \g2493/_0_  = ~n27425 ;
  assign \g2494/_0_  = ~n27453 ;
  assign \g2495/_0_  = ~n27481 ;
  assign \g2496/_0_  = n27493 ;
  assign \g2497/_0_  = n27496 ;
  assign \g2507/_0_  = ~n27506 ;
  assign \g2508/_0_  = ~n27515 ;
  assign \g2509/_0_  = ~n27524 ;
  assign \g2510/_0_  = ~n27533 ;
  assign \g2511/_0_  = ~n27542 ;
  assign \g2512/_0_  = ~n27551 ;
  assign \g2513/_0_  = ~n27560 ;
  assign \g2514/_0_  = ~n27586 ;
  assign \g2515/_0_  = ~n27612 ;
  assign \g2516/_0_  = ~n27621 ;
  assign \g25237/_0_  = ~\T_IRQE0n_pad  ;
  assign \g2558/_0_  = ~n27626 ;
  assign \g2562/_0_  = ~n27652 ;
  assign \g2563/_0_  = ~n27678 ;
  assign \g2564/_0_  = ~n27704 ;
  assign \g2565/_0_  = ~n27730 ;
  assign \g2566/_0_  = ~n27756 ;
  assign \g2567/_0_  = ~n27782 ;
  assign \g2699/_0_  = ~n26394 ;
  assign \g27/_2_  = ~n27786 ;
  assign \g271/_0_  = ~n26317 ;
  assign \g272/_3_  = ~n27805 ;
  assign \g273/_3_  = ~n27818 ;
  assign \g274/_3_  = n27824 ;
  assign \g275/_3_  = n27830 ;
  assign \g276/_3_  = ~n27840 ;
  assign \g277/_3_  = n27846 ;
  assign \g2787/_3_  = ~n27856 ;
  assign \g2788/_3_  = n27862 ;
  assign \g279/_0_  = ~n27872 ;
  assign \g2795/_0_  = n27878 ;
  assign \g2796/_0_  = n27881 ;
  assign \g280/_0_  = n27887 ;
  assign \g2842/_3_  = ~n27902 ;
  assign \g29/_1_  = n27904 ;
  assign \g2927/_0_  = ~n28157 ;
  assign \g2978/_0_  = ~n28167 ;
  assign \g2979/_0_  = ~n28172 ;
  assign \g2980/_0_  = ~n28177 ;
  assign \g2981/_0_  = ~n28182 ;
  assign \g2982/_0_  = ~n28187 ;
  assign \g2983/_0_  = ~n28192 ;
  assign \g2984/_0_  = ~n28197 ;
  assign \g2985/_0_  = ~n28202 ;
  assign \g3021/_3_  = n28210 ;
  assign \g3022/_3_  = n28216 ;
  assign \g3023/_3_  = n28222 ;
  assign \g3024/_3_  = n28228 ;
  assign \g3025/_3_  = n28234 ;
  assign \g3026/_3_  = n28240 ;
  assign \g3027/_3_  = n28246 ;
  assign \g3028/_3_  = n28252 ;
  assign \g3029/_3_  = n28261 ;
  assign \g3030/_3_  = n28270 ;
  assign \g3031/_3_  = n28279 ;
  assign \g3032/_3_  = n28288 ;
  assign \g3033/_3_  = n28297 ;
  assign \g3034/_3_  = n28306 ;
  assign \g3035/_3_  = n28315 ;
  assign \g3036/_3_  = n28324 ;
  assign \g3037/_3_  = n28330 ;
  assign \g3038/_3_  = n28336 ;
  assign \g3039/_3_  = n28342 ;
  assign \g3040/_3_  = n28348 ;
  assign \g3041/_3_  = n28354 ;
  assign \g3042/_3_  = n28360 ;
  assign \g3049/_0_  = ~n28363 ;
  assign \g3050/_0_  = ~n28366 ;
  assign \g3051/_0_  = ~n28369 ;
  assign \g3052/_0_  = ~n28372 ;
  assign \g3053/_0_  = ~n28375 ;
  assign \g3054/_0_  = ~n28378 ;
  assign \g3058/_0_  = ~n28381 ;
  assign \g3059/_0_  = ~n28384 ;
  assign \g3088/_0_  = ~n28393 ;
  assign \g3089/_0_  = ~n28401 ;
  assign \g3090/_0_  = ~n28409 ;
  assign \g3091/_0_  = ~n28417 ;
  assign \g3092/_0_  = ~n28425 ;
  assign \g3093/_0_  = ~n28433 ;
  assign \g3094/_0_  = ~n28441 ;
  assign \g3095/_0_  = ~n28449 ;
  assign \g314/_0_  = ~n27053 ;
  assign \g3147/_3_  = n28455 ;
  assign \g3148/_3_  = n28461 ;
  assign \g3189/_0_  = ~n28467 ;
  assign \g3190/_0_  = ~n28473 ;
  assign \g3191/_0_  = ~n28479 ;
  assign \g3192/_0_  = ~n28485 ;
  assign \g3193/_0_  = ~n28491 ;
  assign \g3194/_0_  = ~n28497 ;
  assign \g3195/_0_  = ~n28503 ;
  assign \g3196/_0_  = ~n28509 ;
  assign \g3197/_0_  = ~n28515 ;
  assign \g3198/_0_  = ~n28521 ;
  assign \g3199/_0_  = ~n28527 ;
  assign \g32/_0_  = n28542 ;
  assign \g320/_3_  = ~n28669 ;
  assign \g3200/_0_  = ~n28675 ;
  assign \g3201/_0_  = ~n28681 ;
  assign \g3202/_0_  = ~n28687 ;
  assign \g3203/_0_  = ~n28693 ;
  assign \g3204/_0_  = ~n28699 ;
  assign \g321/_3_  = ~n28755 ;
  assign \g325/_3_  = ~n28763 ;
  assign \g3271/_2_  = n26388 ;
  assign \g33/_0_  = n28773 ;
  assign \g3363/_0_  = n28785 ;
  assign \g3413/_0_  = ~n28875 ;
  assign \g3414/_0_  = ~n28965 ;
  assign \g352/_0_  = n27803 ;
  assign \g355/_0_  = ~n27816 ;
  assign \g356/_3_  = ~n28975 ;
  assign \g357/_3_  = n28981 ;
  assign \g35_dup/_1_  = n28982 ;
  assign \g36/_3_  = ~n28985 ;
  assign \g365/_3_  = ~n29038 ;
  assign \g366/_3_  = ~n29127 ;
  assign \g367/_3_  = ~n29178 ;
  assign \g368/_3_  = ~n29227 ;
  assign \g3687/_0_  = n29232 ;
  assign \g369/_3_  = ~n29340 ;
  assign \g37/_3_  = ~n29343 ;
  assign \g370/_3_  = ~n29364 ;
  assign \g372/_3_  = ~n29385 ;
  assign \g374/_3_  = ~n29406 ;
  assign \g3740/_0_  = n29411 ;
  assign \g375/_3_  = ~n29432 ;
  assign \g376/_3_  = ~n29453 ;
  assign \g3878/_0_  = ~n29461 ;
  assign \g3879/_0_  = ~n29466 ;
  assign \g388/_3_  = ~n29476 ;
  assign \g3880/_0_  = n29485 ;
  assign \g3881/_0_  = ~n29490 ;
  assign \g3882/_0_  = n29498 ;
  assign \g389/_3_  = n29504 ;
  assign \g3894/_0_  = ~n29507 ;
  assign \g3895/_0_  = ~n29510 ;
  assign \g3896/_0_  = ~n29513 ;
  assign \g3897/_0_  = n29516 ;
  assign \g3898/_0_  = n29519 ;
  assign \g392/_3_  = ~n29669 ;
  assign \g393/_3_  = ~n29731 ;
  assign \g394/_3_  = ~n29882 ;
  assign \g395/_3_  = ~n29987 ;
  assign \g396/_3_  = ~n29995 ;
  assign \g397/_3_  = ~n30003 ;
  assign \g398/_3_  = ~n30011 ;
  assign \g399/_3_  = ~n30019 ;
  assign \g401/_3_  = n30155 ;
  assign \g402/_3_  = ~n30163 ;
  assign \g404/_3_  = n30261 ;
  assign \g4048/_0_  = ~n30266 ;
  assign \g405/_3_  = n30324 ;
  assign \g4050/_0_  = ~n30329 ;
  assign \g406/_3_  = ~n30337 ;
  assign \g407/_3_  = ~n30345 ;
  assign \g410/_3_  = ~n30485 ;
  assign \g411/_3_  = ~n30493 ;
  assign \g412/_3_  = ~n30542 ;
  assign \g413/_3_  = ~n30647 ;
  assign \g415/_3_  = ~n30668 ;
  assign \g416/_3_  = ~n30689 ;
  assign \g42/_0_  = ~n30699 ;
  assign \g4216/_3_  = ~n30709 ;
  assign \g4217/_3_  = ~n30718 ;
  assign \g4218/_3_  = n30726 ;
  assign \g4219/_3_  = ~n30740 ;
  assign \g4296/_0_  = ~n30764 ;
  assign \g4297/_0_  = ~n30788 ;
  assign \g4298/_0_  = ~n30792 ;
  assign \g4299/_0_  = ~n30796 ;
  assign \g43/_0_  = n30804 ;
  assign \g4300/_0_  = ~n30808 ;
  assign \g4301/_0_  = ~n30812 ;
  assign \g4302/_0_  = ~n30816 ;
  assign \g4303/_0_  = ~n30820 ;
  assign \g4304/_0_  = ~n30824 ;
  assign \g4305/_0_  = ~n30828 ;
  assign \g4306/_0_  = ~n30832 ;
  assign \g4307/_0_  = ~n30836 ;
  assign \g4308/_0_  = ~n30840 ;
  assign \g4309/_0_  = ~n30844 ;
  assign \g4310/_0_  = ~n30848 ;
  assign \g4311/_0_  = ~n30852 ;
  assign \g4312/_0_  = ~n30856 ;
  assign \g4313/_0_  = ~n30860 ;
  assign \g4314/_0_  = ~n30864 ;
  assign \g4315/_0_  = ~n30868 ;
  assign \g4316/_0_  = ~n30872 ;
  assign \g4317/_0_  = ~n30876 ;
  assign \g4318/_0_  = ~n30880 ;
  assign \g4319/_0_  = ~n30884 ;
  assign \g4320/_0_  = ~n30888 ;
  assign \g4321/_0_  = ~n30892 ;
  assign \g4322/_0_  = ~n30896 ;
  assign \g4323/_0_  = ~n30900 ;
  assign \g436/_0_  = n30904 ;
  assign \g44/_0_  = ~n30914 ;
  assign \g448/_3_  = ~n30922 ;
  assign \g45/_0_  = n30932 ;
  assign \g4587/_0_  = ~n30989 ;
  assign \g4588/_0_  = ~n30992 ;
  assign \g46/_0_  = n17796 ;
  assign \g4601/_0_  = ~n30997 ;
  assign \g4602/_0_  = ~n31002 ;
  assign \g4613/_3_  = ~n31010 ;
  assign \g4614/_3_  = ~n31019 ;
  assign \g4615/_3_  = ~n31027 ;
  assign \g463/_0_  = ~n31062 ;
  assign \g465/_0_  = ~n31067 ;
  assign \g4653/_0_  = n31109 ;
  assign \g4654/_0_  = n31118 ;
  assign \g4655/_0_  = n31125 ;
  assign \g4656/_0_  = n31130 ;
  assign \g4659/_0_  = n31133 ;
  assign \g466/_0_  = ~n31137 ;
  assign \g468/_3_  = ~n31147 ;
  assign \g469/_3_  = n31153 ;
  assign \g4697/_0_  = ~n31158 ;
  assign \g47/_3_  = ~n31168 ;
  assign \g470/_0_  = ~n31183 ;
  assign \g471/_0_  = ~n31186 ;
  assign \g4755/_0_  = n31189 ;
  assign \g476/_0_  = n31226 ;
  assign \g48/_3_  = n31232 ;
  assign \g480/_00_  = n31256 ;
  assign \g4839/_0_  = ~n31276 ;
  assign \g4840/_0_  = ~n31279 ;
  assign \g485/_3_  = ~n31282 ;
  assign \g4854/_0_  = ~n31287 ;
  assign \g4855/_0_  = ~n31292 ;
  assign \g4859/_0_  = ~n31297 ;
  assign \g486/_3_  = ~n31300 ;
  assign \g4860/_0_  = ~n31305 ;
  assign \g4880/_0_  = n31353 ;
  assign \g4881/_0_  = n31365 ;
  assign \g4882/_0_  = n31377 ;
  assign \g4883/_0_  = n31389 ;
  assign \g4884/_0_  = n31423 ;
  assign \g4885/_0_  = n31435 ;
  assign \g4886/_0_  = n31447 ;
  assign \g4887/_0_  = n31459 ;
  assign \g4888/_0_  = n31471 ;
  assign \g49/_0_  = ~n31484 ;
  assign \g494/_0_  = ~n5673 ;
  assign \g499/_1_  = ~n5642 ;
  assign \g50/_0_  = n31490 ;
  assign \g5002/_0_  = n31534 ;
  assign \g5003/_0_  = n31543 ;
  assign \g5009/_0_  = n31551 ;
  assign \g5010/_0_  = n31558 ;
  assign \g5011/_0_  = n31568 ;
  assign \g5014/_0_  = n31571 ;
  assign \g51/_0_  = ~n31574 ;
  assign \g5105/_0_  = n31577 ;
  assign \g5129/_2_  = n31585 ;
  assign \g5132/_0_  = n31615 ;
  assign \g5135/_0_  = n31645 ;
  assign \g5168/_0_  = ~n31662 ;
  assign \g5169/_0_  = ~n31665 ;
  assign \g5173/_0_  = ~n31670 ;
  assign \g5224/_0_  = ~n31675 ;
  assign \g5225/_0_  = ~n31680 ;
  assign \g5226/_0_  = ~n31685 ;
  assign \g5227/_0_  = ~n31690 ;
  assign \g5334/_0_  = ~n31709 ;
  assign \g5335/_0_  = ~n31715 ;
  assign \g5336/_0_  = ~n31721 ;
  assign \g5337/_0_  = ~n31725 ;
  assign \g5338/_0_  = ~n31734 ;
  assign \g5339/_0_  = ~n31743 ;
  assign \g5340/_0_  = ~n31752 ;
  assign \g5341/_0_  = ~n31761 ;
  assign \g5342/_0_  = ~n31770 ;
  assign \g5343/_0_  = ~n31779 ;
  assign \g5344/_0_  = ~n31788 ;
  assign \g5345/_0_  = ~n31797 ;
  assign \g5346/_0_  = ~n31806 ;
  assign \g5347/_0_  = ~n31815 ;
  assign \g5348/_0_  = ~n31824 ;
  assign \g5349/_0_  = ~n31833 ;
  assign \g5395/_0_  = n31836 ;
  assign \g54/_0_  = ~n31839 ;
  assign \g5434/_0_  = n31849 ;
  assign \g5447/_0_  = n31855 ;
  assign \g5450/_0_  = n31874 ;
  assign \g5451/_0_  = ~n31880 ;
  assign \g5452/_0_  = ~n31886 ;
  assign \g5453/_0_  = ~n31892 ;
  assign \g5454/_0_  = ~n31896 ;
  assign \g5461/_0_  = n31899 ;
  assign \g5483/_0_  = n31907 ;
  assign \g5484/_0_  = n31929 ;
  assign \g5492/_0_  = ~n31932 ;
  assign \g5493/_0_  = ~n31938 ;
  assign \g5496/_3_  = ~n31948 ;
  assign \g5497/_3_  = n31954 ;
  assign \g55/_0_  = ~n31957 ;
  assign \g5500/_0_  = n31964 ;
  assign \g5502/_0_  = n31988 ;
  assign \g5503/_0_  = ~n32034 ;
  assign \g5506/_0_  = n32044 ;
  assign \g5511/_0_  = n32093 ;
  assign \g5518/_0_  = n32105 ;
  assign \g5519/_0_  = n32117 ;
  assign \g5520/_0_  = n32129 ;
  assign \g5522/_0_  = n32141 ;
  assign \g5523/_0_  = n32153 ;
  assign \g5524/_0_  = n32165 ;
  assign \g5525/_0_  = n32177 ;
  assign \g5532/_0_  = ~n32182 ;
  assign \g5533/_0_  = ~n32187 ;
  assign \g5534/_0_  = ~n32192 ;
  assign \g5535/_0_  = ~n32197 ;
  assign \g5536/_0_  = ~n32203 ;
  assign \g5537/_0_  = ~n32209 ;
  assign \g5538/_0_  = ~n32215 ;
  assign \g5546/_0_  = n32223 ;
  assign \g5555/_00_  = n32251 ;
  assign \g5593/_0_  = n4148 ;
  assign \g5614/_2_  = ~n6929 ;
  assign \g567/_0_  = n32255 ;
  assign \g5677/_0_  = n32258 ;
  assign \g5678/_0_  = n32261 ;
  assign \g5682/_0_  = n32265 ;
  assign \g5683/_0_  = n32270 ;
  assign \g5684/_0_  = n32274 ;
  assign \g5686/_0_  = n32280 ;
  assign \g5687/_0_  = n32284 ;
  assign \g5689/_0_  = n32289 ;
  assign \g5690/_0_  = n32293 ;
  assign \g5691/_0_  = n32298 ;
  assign \g5692/_0_  = n32302 ;
  assign \g5698/_0_  = n32305 ;
  assign \g5699/_0_  = n32308 ;
  assign \g5700/_0_  = n32312 ;
  assign \g5701/_0_  = n32315 ;
  assign \g5702/_0_  = n32318 ;
  assign \g5703/_0_  = n32319 ;
  assign \g5704/_0_  = n32335 ;
  assign \g5709/_0_  = n32338 ;
  assign \g5711/_0_  = n32341 ;
  assign \g5714/_0_  = n32342 ;
  assign \g572/_0_  = n32348 ;
  assign \g5723/_0_  = n32356 ;
  assign \g5724/_0_  = n32363 ;
  assign \g5725/_0_  = ~n32390 ;
  assign \g573/_0_  = n32393 ;
  assign \g5739/_0_  = ~n32409 ;
  assign \g5740/_0_  = ~n32419 ;
  assign \g575/_0_  = ~n32422 ;
  assign \g5756/_0_  = ~n32425 ;
  assign \g5757/_0_  = ~n32428 ;
  assign \g5758/_0_  = ~n32431 ;
  assign \g5759/_0_  = ~n32434 ;
  assign \g576/_0_  = ~n32437 ;
  assign \g5760/_0_  = ~n32440 ;
  assign \g5761/_0_  = ~n32443 ;
  assign \g5762/_0_  = ~n32446 ;
  assign \g5763/_0_  = ~n32449 ;
  assign \g577/_0_  = ~n32452 ;
  assign \g5772/_0_  = ~n32480 ;
  assign \g5773/_0_  = ~n32489 ;
  assign \g5774/_0_  = ~n32501 ;
  assign \g5775/_0_  = n32509 ;
  assign \g5776/_0_  = ~n32517 ;
  assign \g5777/_0_  = ~n32525 ;
  assign \g578/_0_  = ~n32528 ;
  assign \g5781/_0_  = ~n32538 ;
  assign \g5783/_0_  = ~n32546 ;
  assign \g5784/_0_  = ~n32554 ;
  assign \g5785/_0_  = ~n32562 ;
  assign \g5786/_0_  = ~n32570 ;
  assign \g5787/_0_  = ~n32578 ;
  assign \g5788/_0_  = ~n32586 ;
  assign \g5789/_0_  = ~n32594 ;
  assign \g579/_0_  = ~n32597 ;
  assign \g5790/_0_  = ~n32600 ;
  assign \g5791/_0_  = ~n32603 ;
  assign \g5792/_0_  = ~n32605 ;
  assign \g5794/_0_  = ~n32622 ;
  assign \g5795/_0_  = ~n32625 ;
  assign \g5796/_0_  = ~n32628 ;
  assign \g580/_0_  = ~n32631 ;
  assign \g5801/_0_  = ~n32634 ;
  assign \g5802/_0_  = ~n32637 ;
  assign \g5803/_0_  = ~n32641 ;
  assign \g5804/_0_  = ~n32645 ;
  assign \g5805/_0_  = ~n32648 ;
  assign \g581/_0_  = ~n32651 ;
  assign \g5814/_0_  = ~n32668 ;
  assign \g582/_0_  = ~n32671 ;
  assign \g583/_0_  = ~n32674 ;
  assign \g5849/_3_  = ~n32682 ;
  assign \g585/_0_  = ~n32685 ;
  assign \g586/_0_  = ~n32688 ;
  assign \g587/_0_  = ~n32691 ;
  assign \g588/_0_  = ~n32694 ;
  assign \g589/_0_  = ~n32697 ;
  assign \g590/_0_  = ~n32700 ;
  assign \g591/_0_  = ~n32703 ;
  assign \g592/_0_  = ~n32706 ;
  assign \g593/_0_  = ~n32709 ;
  assign \g594/_0_  = ~n32712 ;
  assign \g595/_0_  = ~n32715 ;
  assign \g596/_0_  = ~n32718 ;
  assign \g597/_0_  = ~n32721 ;
  assign \g5971/_0_  = n32724 ;
  assign \g5972/_0_  = n32727 ;
  assign \g5976/_0_  = n32730 ;
  assign \g598/_0_  = ~n32733 ;
  assign \g5989/_0_  = n32736 ;
  assign \g599/_0_  = ~n32739 ;
  assign \g600/_0_  = ~n32742 ;
  assign \g601/_0_  = ~n32745 ;
  assign \g602/_0_  = ~n32748 ;
  assign \g603/_0_  = ~n32751 ;
  assign \g604/_0_  = ~n32754 ;
  assign \g605/_0_  = ~n32757 ;
  assign \g6092/_0_  = ~n32760 ;
  assign \g6093/_2_  = ~n32953 ;
  assign \g6094/_0_  = ~n32958 ;
  assign \g6114/_0_  = n32959 ;
  assign \g614/_3_  = ~n32967 ;
  assign \g6148/_0_  = ~n32969 ;
  assign \g6149/_0_  = ~n32971 ;
  assign \g6171/_0_  = n33008 ;
  assign \g6172/_0_  = n33020 ;
  assign \g6173/_0_  = n33032 ;
  assign \g6174/_0_  = n33044 ;
  assign \g6175/_0_  = n33056 ;
  assign \g6176/_0_  = n33068 ;
  assign \g6177/_0_  = n33080 ;
  assign \g6178/_0_  = n33115 ;
  assign \g6179/_0_  = n33127 ;
  assign \g6180/_0_  = n33139 ;
  assign \g6181/_0_  = n33151 ;
  assign \g6182/_0_  = n33163 ;
  assign \g6183/_0_  = n33175 ;
  assign \g6184/_0_  = n33187 ;
  assign \g6185/_0_  = n33199 ;
  assign \g6186/_0_  = ~n33226 ;
  assign \g6187/_0_  = ~n33251 ;
  assign \g6193/_0_  = ~n33273 ;
  assign \g6196/_0_  = n33290 ;
  assign \g6197/_0_  = n33303 ;
  assign \g6198/_3_  = ~n33319 ;
  assign \g6200/_2_  = n31701 ;
  assign \g6202/_2_  = n31861 ;
  assign \g6203/_3_  = ~n33329 ;
  assign \g6204/_3_  = n33335 ;
  assign \g6209/_0_  = ~n33349 ;
  assign \g6211/_0_  = ~n33352 ;
  assign \g6215/_0_  = ~n33376 ;
  assign \g6217/_0_  = ~n33401 ;
  assign \g6219/_0_  = ~n33426 ;
  assign \g6220/_0_  = ~n33450 ;
  assign \g6222/_0_  = ~n33475 ;
  assign \g6224/_0_  = ~n33500 ;
  assign \g6228/_0_  = ~n33522 ;
  assign \g6238/_0_  = ~n33525 ;
  assign \g6239/_0_  = ~n33528 ;
  assign \g6240/_0_  = ~n33531 ;
  assign \g6242/_0_  = ~n33534 ;
  assign \g6243/_0_  = ~n33537 ;
  assign \g6244/_0_  = ~n33540 ;
  assign \g6245/_0_  = ~n33543 ;
  assign \g6246/_0_  = ~n33546 ;
  assign \g6248/_0_  = ~n33549 ;
  assign \g6249/_0_  = ~n33552 ;
  assign \g6259/_0_  = ~n33557 ;
  assign \g6260/_0_  = ~n33563 ;
  assign \g6261/_0_  = n33568 ;
  assign \g6262/_0_  = ~n33573 ;
  assign \g6263/_0_  = n33578 ;
  assign \g6264/_0_  = ~n33584 ;
  assign \g6265/_0_  = ~n33589 ;
  assign \g6266/_0_  = ~n33594 ;
  assign \g6267/_0_  = n33600 ;
  assign \g6268/_0_  = ~n33605 ;
  assign \g6269/_0_  = ~n33611 ;
  assign \g6270/_0_  = ~n33616 ;
  assign \g6271/_0_  = ~n33620 ;
  assign \g6272/_0_  = n33625 ;
  assign \g6277/_0_  = ~n33630 ;
  assign \g6318/_0_  = n33632 ;
  assign \g6326/_0_  = ~n33635 ;
  assign \g6329/_0_  = n33647 ;
  assign \g6330/_0_  = n33659 ;
  assign \g6331/_0_  = n33671 ;
  assign \g6332/_0_  = n33683 ;
  assign \g6333/_0_  = n33706 ;
  assign \g6334/_0_  = n33718 ;
  assign \g6335/_0_  = n33730 ;
  assign \g6336/_0_  = n33742 ;
  assign \g6337/_0_  = n33754 ;
  assign \g6338/_0_  = n33766 ;
  assign \g6339/_0_  = n33778 ;
  assign \g6340/_0_  = n33790 ;
  assign \g6341/_0_  = n33802 ;
  assign \g6342/_0_  = n33814 ;
  assign \g6343/_0_  = n33826 ;
  assign \g6344/_0_  = n33838 ;
  assign \g6345/_0_  = n33850 ;
  assign \g6346/_0_  = n33862 ;
  assign \g6347/_0_  = n33874 ;
  assign \g6348/_0_  = n33886 ;
  assign \g6349/_0_  = n33905 ;
  assign \g6350/_0_  = n33919 ;
  assign \g6351/_0_  = n33932 ;
  assign \g6352/_0_  = n33945 ;
  assign \g6353/_0_  = n33957 ;
  assign \g6354/_0_  = n33969 ;
  assign \g6355/_0_  = n33981 ;
  assign \g6361/_0_  = n33983 ;
  assign \g637/_0_  = n33989 ;
  assign \g638/_0_  = n33992 ;
  assign \g639/_3_  = ~n34002 ;
  assign \g64/_3_  = ~n34005 ;
  assign \g640/_3_  = n34011 ;
  assign \g6419/_0_  = n5681 ;
  assign \g6442/_0_  = ~n12234 ;
  assign \g6442/_1_  = n12234 ;
  assign \g6489/_0_  = n34012 ;
  assign \g6490/_0_  = n34013 ;
  assign \g65/_3_  = ~n34016 ;
  assign \g6513/_0_  = n34019 ;
  assign \g6515/_0_  = n34022 ;
  assign \g6571/_0_  = n34048 ;
  assign \g6588/_0_  = n34051 ;
  assign \g6589/_0_  = n34054 ;
  assign \g6638/_0_  = n34058 ;
  assign \g6639/_0_  = ~n34072 ;
  assign \g6653/_0_  = n34077 ;
  assign \g6654/_3_  = ~n34096 ;
  assign \g6655/_0_  = ~n34101 ;
  assign \g6656/_0_  = ~n34107 ;
  assign \g6657/_0_  = ~n34112 ;
  assign \g6687/_0_  = ~n34134 ;
  assign \g6688/_0_  = ~n34138 ;
  assign \g6689/_0_  = ~n34142 ;
  assign \g6690/_0_  = ~n34146 ;
  assign \g6691/_0_  = ~n34150 ;
  assign \g6692/_0_  = ~n34154 ;
  assign \g6693/_0_  = ~n34158 ;
  assign \g6694/_0_  = ~n34162 ;
  assign \g6701/_0_  = n34164 ;
  assign \g6706/_0_  = n34169 ;
  assign \g6711/_0_  = n34171 ;
  assign \g6727/_0_  = ~n34193 ;
  assign \g6728/_0_  = ~n34215 ;
  assign \g6736/_0_  = n34217 ;
  assign \g6739/_0_  = ~n34239 ;
  assign \g6742/_0_  = ~n34244 ;
  assign \g6746/_0_  = n34246 ;
  assign \g6752/_0_  = ~n34251 ;
  assign \g6771/_0_  = n34253 ;
  assign \g684/_0_  = n34283 ;
  assign \g685/_0_  = n34289 ;
  assign \g686/_0_  = n34295 ;
  assign \g687/_0_  = n34299 ;
  assign \g688/_0_  = n34305 ;
  assign \g689/_0_  = n34308 ;
  assign \g690/_0_  = n34314 ;
  assign \g691/_0_  = n34317 ;
  assign \g692/_0_  = n34320 ;
  assign \g693/_0_  = n34323 ;
  assign \g696/_3_  = ~n34333 ;
  assign \g697/_3_  = n34339 ;
  assign \g699/_0_  = ~n34378 ;
  assign \g7/_0_  = n34388 ;
  assign \g700/_0_  = ~n34418 ;
  assign \g7005/_0_  = n34434 ;
  assign \g7056/_0_  = n34437 ;
  assign \g7057/_0_  = n31705 ;
  assign \g7058/_0_  = n31868 ;
  assign \g7060/_0_  = n34440 ;
  assign \g7075/_0_  = n34460 ;
  assign \g7086/_0_  = n34468 ;
  assign \g7087/_0_  = n34473 ;
  assign \g7089/_0_  = n34483 ;
  assign \g7108/_0_  = n34489 ;
  assign \g7109/_0_  = n34495 ;
  assign \g7112/_0_  = ~n32088 ;
  assign \g7172/_2_  = ~n33344 ;
  assign \g7210/_2_  = ~n32658 ;
  assign \g7211/_0_  = n34500 ;
  assign \g7212/_0_  = n34505 ;
  assign \g7213/_0_  = n34510 ;
  assign \g7214/_0_  = n34515 ;
  assign \g7215/_0_  = ~n34520 ;
  assign \g7216/_0_  = ~n34525 ;
  assign \g7217/_3_  = ~n34531 ;
  assign \g7218/_0_  = ~n34536 ;
  assign \g7219/_0_  = ~n34541 ;
  assign \g7220/_0_  = ~n34546 ;
  assign \g7222/_0_  = ~n34551 ;
  assign \g7227/_2_  = ~n32612 ;
  assign \g723/_3_  = ~n34554 ;
  assign \g7234/_0_  = ~n34559 ;
  assign \g7237/_3_  = n34564 ;
  assign \g7238/_3_  = n34569 ;
  assign \g7239/_3_  = n13773 ;
  assign \g724/_3_  = ~n34572 ;
  assign \g7240/_3_  = n34578 ;
  assign \g7241/_3_  = n34583 ;
  assign \g7242/_3_  = n34588 ;
  assign \g7243/_3_  = n34593 ;
  assign \g7244/_0_  = ~n34598 ;
  assign \g7245/_0_  = ~n34603 ;
  assign \g7246/_0_  = ~n34608 ;
  assign \g7247/_0_  = ~n34613 ;
  assign \g7248/_0_  = ~n34618 ;
  assign \g7249/_0_  = ~n34623 ;
  assign \g7250/_0_  = ~n34628 ;
  assign \g7251/_0_  = ~n34633 ;
  assign \g7253/_0_  = n34637 ;
  assign \g7254/_0_  = ~n34640 ;
  assign \g7255/_0_  = n34642 ;
  assign \g7256/_0_  = n34644 ;
  assign \g7257/_0_  = n34646 ;
  assign \g7258/_0_  = n34648 ;
  assign \g7261/_0_  = n34650 ;
  assign \g7264/_0_  = n34662 ;
  assign \g7265/_0_  = n34674 ;
  assign \g7266/_0_  = n34686 ;
  assign \g7267/_0_  = n34698 ;
  assign \g7268/_0_  = n34710 ;
  assign \g7269/_0_  = n34722 ;
  assign \g7278/_0_  = n34734 ;
  assign \g7279/_0_  = n34746 ;
  assign \g7280/_0_  = n34758 ;
  assign \g7281/_0_  = n34770 ;
  assign \g7282/_0_  = n34782 ;
  assign \g7283/_0_  = n34794 ;
  assign \g7284/_0_  = n34806 ;
  assign \g7285/_0_  = n34818 ;
  assign \g7286/_3_  = ~n26973 ;
  assign \g7288/_3_  = ~n34822 ;
  assign \g7291/_0_  = n34824 ;
  assign \g7296/_3_  = n34863 ;
  assign \g73/_0_  = n34873 ;
  assign \g7302/_3_  = n34894 ;
  assign \g7306/_3_  = n34916 ;
  assign \g7310/_3_  = ~n34928 ;
  assign \g7311/_3_  = ~n34937 ;
  assign \g7312/_3_  = ~n34946 ;
  assign \g7313/_3_  = ~n34955 ;
  assign \g7314/_3_  = ~n34964 ;
  assign \g7315/_3_  = ~n34973 ;
  assign \g7316/_3_  = ~n34982 ;
  assign \g7317/_3_  = ~n34991 ;
  assign \g7323/_3_  = n35026 ;
  assign \g7324/_3_  = n35060 ;
  assign \g7325/_3_  = n35094 ;
  assign \g7327/_0_  = n35096 ;
  assign \g7362/_0_  = n35098 ;
  assign \g74/_0_  = n35108 ;
  assign \g75/_0_  = n35118 ;
  assign \g7512/_0_  = n13758 ;
  assign \g7513/_0_  = n35126 ;
  assign \g7514/_0_  = n35127 ;
  assign \g7515/_0_  = n35128 ;
  assign \g7516/_0_  = n35129 ;
  assign \g7518/_0_  = n35138 ;
  assign \g7528/_0_  = n35147 ;
  assign \g7529/_0_  = n35150 ;
  assign \g7548/_0_  = n35154 ;
  assign \g7549/_0_  = n35158 ;
  assign \g7550/_0_  = n35162 ;
  assign \g7575/_0_  = n35168 ;
  assign \g7576/_0_  = n35173 ;
  assign \g7577/_0_  = n35177 ;
  assign \g7578/_0_  = n35181 ;
  assign \g7579/_0_  = n35189 ;
  assign \g7580/_0_  = n35194 ;
  assign \g7581/_0_  = n35199 ;
  assign \g7582/_0_  = n35203 ;
  assign \g7583/_0_  = n35207 ;
  assign \g7584/_0_  = n35213 ;
  assign \g7585/_0_  = n35219 ;
  assign \g7586/_0_  = n35225 ;
  assign \g7587/_0_  = n35230 ;
  assign \g7588/_0_  = n35234 ;
  assign \g7589/_0_  = n35238 ;
  assign \g7590/_0_  = n35242 ;
  assign \g7591/_0_  = n35248 ;
  assign \g7592/_0_  = n35252 ;
  assign \g7593/_0_  = n35256 ;
  assign \g7594/_0_  = n35260 ;
  assign \g7595/_0_  = n35264 ;
  assign \g7596/_0_  = n35268 ;
  assign \g7597/_0_  = n35273 ;
  assign \g7598/_0_  = n35277 ;
  assign \g7599/_0_  = n35281 ;
  assign \g76/_0_  = n35291 ;
  assign \g7600/_0_  = n35295 ;
  assign \g7601/_0_  = n35299 ;
  assign \g7602/_0_  = n35303 ;
  assign \g7603/_0_  = n35308 ;
  assign \g7604/_0_  = n35312 ;
  assign \g7614/_0_  = n35317 ;
  assign \g7618/_0_  = ~n35318 ;
  assign \g762/_0_  = n35322 ;
  assign \g7634/_0_  = n32758 ;
  assign \g766/_0_  = n35328 ;
  assign \g767/_0_  = n35331 ;
  assign \g768/_0_  = n35337 ;
  assign \g769/_0_  = n35340 ;
  assign \g77/_0_  = n35350 ;
  assign \g770/_3_  = ~n35360 ;
  assign \g771/_3_  = n35366 ;
  assign \g7715/_0_  = ~n35397 ;
  assign \g774/_0_  = ~n35414 ;
  assign \g7746/_0_  = n35417 ;
  assign \g7753/_0_  = n35421 ;
  assign \g7754/_0_  = n35424 ;
  assign \g7755/_0_  = n35427 ;
  assign \g7756/_0_  = n35430 ;
  assign \g7757/_0_  = n35433 ;
  assign \g7758/_0_  = n35458 ;
  assign \g7759/_0_  = n35483 ;
  assign \g7760/_0_  = n35508 ;
  assign \g7761/_0_  = n35533 ;
  assign \g7762/_0_  = ~n35536 ;
  assign \g7763/_0_  = n35539 ;
  assign \g7764/_0_  = n35542 ;
  assign \g7765/_0_  = n35545 ;
  assign \g7766/_0_  = n35570 ;
  assign \g7778/_0_  = ~n35574 ;
  assign \g7779/_0_  = ~n35579 ;
  assign \g7780/_0_  = ~n35584 ;
  assign \g7781/_0_  = ~n35589 ;
  assign \g7782/_0_  = ~n35594 ;
  assign \g7784/_0_  = ~n35599 ;
  assign \g78/_0_  = n35609 ;
  assign \g7800/_0_  = n35611 ;
  assign \g7823/_3_  = ~n35614 ;
  assign \g7837/_0_  = ~n35619 ;
  assign \g7841/_0_  = ~n35624 ;
  assign \g7842/_0_  = ~n35629 ;
  assign \g7843/_0_  = ~n35634 ;
  assign \g7844/_0_  = ~n35639 ;
  assign \g7845/_0_  = ~n35644 ;
  assign \g7846/_0_  = ~n35649 ;
  assign \g7847/_0_  = ~n35654 ;
  assign \g7849/_0_  = n35656 ;
  assign \g7850/_0_  = ~n35661 ;
  assign \g7852/_0_  = n35663 ;
  assign \g7854/_0_  = n35665 ;
  assign \g7855/_0_  = ~n35670 ;
  assign \g7857/_0_  = ~n35677 ;
  assign \g7858/_0_  = ~n35683 ;
  assign \g7859/_0_  = ~n35689 ;
  assign \g7860/_0_  = ~n35695 ;
  assign \g7861/_0_  = ~n35701 ;
  assign \g7862/_0_  = ~n35707 ;
  assign \g7863/_0_  = ~n35713 ;
  assign \g7864/_0_  = ~n35719 ;
  assign \g7865/_0_  = ~n35725 ;
  assign \g7866/_0_  = ~n35731 ;
  assign \g7867/_0_  = ~n35737 ;
  assign \g7868/_0_  = ~n35743 ;
  assign \g7869/_0_  = ~n35749 ;
  assign \g7870/_0_  = ~n35755 ;
  assign \g7871/_0_  = ~n35760 ;
  assign \g79211/_3_  = ~n35763 ;
  assign \g79258/_3_  = ~n35766 ;
  assign \g79299/_3_  = ~n35769 ;
  assign \g79316/_2_  = ~n13534 ;
  assign \g79342/_3_  = ~n35772 ;
  assign \g79401/_3_  = ~n35775 ;
  assign \g79452/_3_  = ~n35778 ;
  assign \g79457/_3_  = ~n35781 ;
  assign \g7951/_0_  = n35783 ;
  assign \g79541/_3_  = ~n35786 ;
  assign \g7958/_0_  = n35788 ;
  assign \g79598/_3_  = ~n35791 ;
  assign \g79654/_3_  = ~n35794 ;
  assign \g79675/_3_  = ~n35797 ;
  assign \g7971/_0_  = ~n35800 ;
  assign \g7972/_0_  = ~n35820 ;
  assign \g7973/_3_  = n35849 ;
  assign \g79753/_3_  = ~n35852 ;
  assign \g7976/_3_  = n35881 ;
  assign \g79855/_3_  = ~n35884 ;
  assign \g79858/_3_  = ~n35887 ;
  assign \g79997/_3_  = ~n35890 ;
  assign \g8/_0_  = n35900 ;
  assign \g80008/_3_  = n11525 ;
  assign \g80011/_0_  = n35901 ;
  assign \g80104/_0_  = ~n19960 ;
  assign \g80172/_1_  = n12451 ;
  assign \g80195/_3_  = n8715 ;
  assign \g80238/_3_  = ~n35904 ;
  assign \g80290/_2_  = n7340 ;
  assign \g80294/_0_  = n10911 ;
  assign \g80302/_0_  = n11265 ;
  assign \g80327/_0_  = ~n35910 ;
  assign \g80360/_3_  = n10289 ;
  assign \g80373/_0_  = ~n35921 ;
  assign \g80401/_0_  = n7607 ;
  assign \g80410/_0_  = n8460 ;
  assign \g80475/_0_  = n7859 ;
  assign \g80476/_0_  = n10638 ;
  assign \g80516/_3_  = n35926 ;
  assign \g80536/_0_  = n35927 ;
  assign \g80537/_0_  = n9178 ;
  assign \g80572/_0_  = n35908 ;
  assign \g80573/_0_  = n35905 ;
  assign \g80609/_2_  = n12688 ;
  assign \g80610/_2_  = n12743 ;
  assign \g80676/_0_  = ~n22677 ;
  assign \g80798/_0_  = ~n35928 ;
  assign \g80807/_0_  = n25905 ;
  assign \g80890/_2_  = n5608 ;
  assign \g80904/_0_  = ~n25905 ;
  assign \g81719/_2_  = n19941 ;
  assign \g81746/_0_  = ~n5586 ;
  assign \g81775/_0_  = ~n5708 ;
  assign \g81872/_0_  = n35935 ;
  assign \g81961/_0_  = ~n4151 ;
  assign \g81968/_0_  = n4172 ;
  assign \g82096/_0_  = ~n4150 ;
  assign \g82123/_0_  = ~n4117 ;
  assign \g82147/_0_  = ~n4149 ;
  assign \g82147/_1_  = n4149 ;
  assign \g82335/_0_  = ~n5581 ;
  assign \g82338/_2_  = ~n5597 ;
  assign \g82368/_0_  = ~n4094 ;
  assign \g82460/_2_  = n22658 ;
  assign \g82469/_0_  = ~n19045 ;
  assign \g82481/_0_  = ~n4093 ;
  assign \g82625/_1_  = n12245 ;
  assign \g82711/_0_  = n5689 ;
  assign \g82772/_0_  = ~n4116 ;
  assign \g82946/_0_  = n22656 ;
  assign \g82947/_0_  = n19939 ;
  assign \g82956/_0_  = ~n5679 ;
  assign \g83003/_0_  = ~n4112 ;
  assign \g83006/_1_  = n12244 ;
  assign \g83415/_0_  = ~n5700 ;
  assign \g83498/_0_  = n4115 ;
  assign \g837/_0_  = n35941 ;
  assign \g838/_0_  = n35944 ;
  assign \g83863/_0_  = n12241 ;
  assign \g839/_0_  = ~n35955 ;
  assign \g84049/_3_  = ~n35961 ;
  assign \g84050/_3_  = ~n35967 ;
  assign \g84077/_2_  = ~n5692 ;
  assign \g842/_0_  = n35973 ;
  assign \g84245/_0_  = ~n4071 ;
  assign \g843/_0_  = ~n35979 ;
  assign \g844/_0_  = ~n35982 ;
  assign \g84448/_0_  = n6988 ;
  assign \g84478/_3_  = ~n35931 ;
  assign \g845/_0_  = n35988 ;
  assign \g846/_0_  = n35991 ;
  assign \g847/_0_  = n35994 ;
  assign \g848/_0_  = n36000 ;
  assign \g8487/_0_  = ~n36006 ;
  assign \g8488/_0_  = ~n36012 ;
  assign \g8489/_0_  = ~n36018 ;
  assign \g849/_0_  = n36021 ;
  assign \g8490/_0_  = ~n36027 ;
  assign \g84904/_0_  = n36028 ;
  assign \g8491/_0_  = ~n36032 ;
  assign \g8492/_0_  = ~n36038 ;
  assign \g8493/_0_  = ~n36042 ;
  assign \g8494/_0_  = ~n36048 ;
  assign \g8496/_0_  = n36049 ;
  assign \g8517/_0_  = n36052 ;
  assign \g8534/_0_  = n36055 ;
  assign \g8538/_0_  = n36064 ;
  assign \g8540/_0_  = n36067 ;
  assign \g8576/_2_  = n32038 ;
  assign \g8597/_0_  = ~n36072 ;
  assign \g8598/_0_  = ~n36078 ;
  assign \g8599/_0_  = ~n36082 ;
  assign \g8600/_0_  = ~n36086 ;
  assign \g8601/_0_  = ~n36090 ;
  assign \g8602/_0_  = ~n36094 ;
  assign \g8603/_0_  = ~n36098 ;
  assign \g8605/_0_  = n36101 ;
  assign \g8606/_0_  = n36104 ;
  assign \g8607/_0_  = n36107 ;
  assign \g8608/_0_  = ~n36112 ;
  assign \g8609/_0_  = ~n36116 ;
  assign \g8610/_0_  = ~n36120 ;
  assign \g8611/_0_  = ~n36124 ;
  assign \g8612/_0_  = ~n36128 ;
  assign \g8613/_0_  = ~n36132 ;
  assign \g8614/_0_  = ~n36136 ;
  assign \g8615/_0_  = ~n36140 ;
  assign \g8617/_0_  = n36143 ;
  assign \g8643/_0_  = ~n36147 ;
  assign \g8644/_0_  = ~n36151 ;
  assign \g8645/_0_  = ~n36155 ;
  assign \g8646/_0_  = ~n36159 ;
  assign \g8647/_0_  = ~n36163 ;
  assign \g8648/_0_  = ~n36167 ;
  assign \g8650/_0_  = n36170 ;
  assign \g8651/_0_  = n36173 ;
  assign \g8652/_0_  = n36176 ;
  assign \g8653/_0_  = ~n36180 ;
  assign \g8654/_0_  = ~n36184 ;
  assign \g8655/_0_  = ~n36188 ;
  assign \g8656/_0_  = ~n36192 ;
  assign \g8657/_0_  = ~n36196 ;
  assign \g8658/_0_  = ~n36200 ;
  assign \g8659/_0_  = ~n36204 ;
  assign \g8660/_0_  = ~n36208 ;
  assign \g8665/_00_  = ~n36217 ;
  assign \g8666/_00_  = ~n36224 ;
  assign \g8667/_00_  = ~n36231 ;
  assign \g8668/_00_  = ~n36238 ;
  assign \g8669/_00_  = ~n36245 ;
  assign \g86715/_0_  = ~n36248 ;
  assign \g86745/_3_  = n9435 ;
  assign \g8691/_0_  = ~n36252 ;
  assign \g8700/_0_  = ~n36259 ;
  assign \g8701/_0_  = ~n36265 ;
  assign \g8702/_0_  = ~n36271 ;
  assign \g8703/_0_  = ~n36277 ;
  assign \g8704/_0_  = ~n36283 ;
  assign \g8705/_0_  = ~n36289 ;
  assign \g87063/_0_  = ~n36321 ;
  assign \g87114/_0_  = ~n36353 ;
  assign \g8712/_0_  = ~n36355 ;
  assign \g8713/_0_  = ~n36361 ;
  assign \g8714/_0_  = ~n36367 ;
  assign \g87171/_1_  = ~n36373 ;
  assign \g87252/_1_  = n4099 ;
  assign \g87298/_0_  = n36374 ;
  assign \g8730/_0_  = ~n36379 ;
  assign \g8741/_0_  = ~n36384 ;
  assign \g8747/_0_  = ~n36387 ;
  assign \g87480/_0_  = n36388 ;
  assign \g87484/_2_  = n23032 ;
  assign \g87488/_1__syn_2  = n26297 ;
  assign \g8761/_0_  = ~n36399 ;
  assign \g8762/_0_  = n36404 ;
  assign \g8763/_0_  = ~n36415 ;
  assign \g8764/_0_  = n36420 ;
  assign \g8765/_0_  = n36426 ;
  assign \g8775/_0_  = ~n36448 ;
  assign \g8776/_0_  = ~n36457 ;
  assign \g8777/_0_  = ~n36461 ;
  assign \g8778/_0_  = ~n36463 ;
  assign \g8784/_0_  = ~n36468 ;
  assign \g8804/_0_  = ~n36476 ;
  assign \g8807/_0_  = ~n36479 ;
  assign \g8808/_0_  = ~n36483 ;
  assign \g8809/_0_  = ~n36487 ;
  assign \g8810/_0_  = ~n36490 ;
  assign \g8811/_0_  = ~n36494 ;
  assign \g8812/_0_  = ~n36497 ;
  assign \g8813/_0_  = n36500 ;
  assign \g8814/_0_  = ~n36503 ;
  assign \g8815/_0_  = ~n36506 ;
  assign \g8816/_0_  = ~n36510 ;
  assign \g8817/_0_  = ~n36513 ;
  assign \g8818/_0_  = ~n36519 ;
  assign \g8819/_0_  = ~n36524 ;
  assign \g8820/_0_  = ~n36529 ;
  assign \g8821/_0_  = ~n36533 ;
  assign \g8822/_0_  = ~n36536 ;
  assign \g8823/_0_  = n36538 ;
  assign \g8824/_0_  = ~n36541 ;
  assign \g8825/_0_  = n36544 ;
  assign \g8826/_0_  = ~n36547 ;
  assign \g8827/_0_  = ~n36550 ;
  assign \g8828/_0_  = ~n36553 ;
  assign \g8829/_0_  = n36555 ;
  assign \g8830/_0_  = ~n36558 ;
  assign \g8831/_0_  = ~n36561 ;
  assign \g8832/_0_  = ~n36564 ;
  assign \g8833/_0_  = ~n36567 ;
  assign \g8834/_0_  = ~n36571 ;
  assign \g8835/_0_  = ~n36574 ;
  assign \g8836/_0_  = ~n36578 ;
  assign \g8837/_0_  = ~n36581 ;
  assign \g8838/_0_  = ~n36584 ;
  assign \g8839/_0_  = n36586 ;
  assign \g8840/_0_  = ~n36589 ;
  assign \g8842/_0_  = ~n36594 ;
  assign \g8843/_0_  = ~n36599 ;
  assign \g8846/_0_  = ~n36602 ;
  assign \g8848/_0_  = n36607 ;
  assign \g8857/_0_  = n36609 ;
  assign \g8895/_0_  = ~n36612 ;
  assign \g8902/_3_  = n36648 ;
  assign \g8903/_3_  = n36684 ;
  assign \g8904/_3_  = n36720 ;
  assign \g8905/_3_  = n36756 ;
  assign \g8906/_3_  = n36792 ;
  assign \g8909/_0_  = ~n36795 ;
  assign \g8910/_0_  = ~n36798 ;
  assign \g8911/_0_  = ~n36801 ;
  assign \g8924/_3_  = n36833 ;
  assign \g8926/_3_  = n36865 ;
  assign \g8927/_3_  = n36897 ;
  assign \g8943/_0_  = n36899 ;
  assign \g8944/_0_  = n36901 ;
  assign \g8958/_3_  = n36933 ;
  assign \g8960/_00_  = ~n36940 ;
  assign \g8961/_3_  = n36972 ;
  assign \g8965/_0_  = ~n36988 ;
  assign \g8966/_0_  = ~n37004 ;
  assign \g8967/_0_  = ~n37020 ;
  assign \g8968/_0_  = ~n37036 ;
  assign \g9/_0_  = n37046 ;
  assign \g9123/_0_  = n32036 ;
  assign \g9125/_0_  = n37047 ;
  assign \g9126/_0_  = n37050 ;
  assign \g913/_0_  = ~n37066 ;
  assign \g915/_0_  = n37072 ;
  assign \g916/_0_  = n37078 ;
  assign \g917/_0_  = n37081 ;
  assign \g918/_0_  = n37087 ;
  assign \g919/_0_  = n37090 ;
  assign \g920/_3_  = ~n37100 ;
  assign \g921/_3_  = n37106 ;
  assign \g925/_0_  = ~n37122 ;
  assign \g926/_0_  = n37125 ;
  assign \g927/_0_  = n37131 ;
  assign \g928/_0_  = n37137 ;
  assign \g929/_0_  = n37140 ;
  assign \g930/_0_  = n37143 ;
  assign \g9336/_0_  = n37146 ;
  assign \g9337/_0_  = n37149 ;
  assign \g939/_3_  = ~n37162 ;
  assign \g9396/_0_  = ~n37168 ;
  assign \g9397/_0_  = ~n37171 ;
  assign \g9399/_0_  = ~n37174 ;
  assign \g9400/_0_  = ~n37177 ;
  assign \g9401/_0_  = ~n37180 ;
  assign \g9402/_0_  = ~n37183 ;
  assign \g9403/_0_  = ~n37186 ;
  assign \g9404/_0_  = ~n37189 ;
  assign \g9415/_0_  = n32613 ;
  assign \g9418/_0_  = n32659 ;
  assign \g9419/_0_  = ~n37202 ;
  assign \g9420/_0_  = n37205 ;
  assign \g9446/_0_  = n37206 ;
  assign \g9465/_0_  = n37207 ;
  assign \g9493/_0_  = ~n37210 ;
  assign \g9536/_0_  = n37214 ;
  assign \g9537/_0_  = ~n37220 ;
  assign \g9538/_0_  = ~n37223 ;
  assign \g9539/_0_  = ~n37226 ;
  assign \g9540/_0_  = ~n37229 ;
  assign \g9541/_0_  = ~n37235 ;
  assign \g9542/_0_  = ~n37239 ;
  assign \g955/_2_  = ~n37247 ;
  assign \g9561/_0_  = ~n37258 ;
  assign \g9562/_0_  = ~n37267 ;
  assign \g9563/_0_  = ~n37276 ;
  assign \g9564/_0_  = ~n37285 ;
  assign \g9565/_0_  = ~n37294 ;
  assign \g9566/_0_  = ~n37303 ;
  assign \g9567/_0_  = ~n37312 ;
  assign \g9568/_0_  = ~n37321 ;
  assign \g9569/_0_  = ~n37331 ;
  assign \g9570/_0_  = ~n37340 ;
  assign \g9571/_0_  = ~n37343 ;
  assign \g9572/_0_  = ~n37352 ;
  assign \g9573/_0_  = ~n37355 ;
  assign \g9574/_0_  = ~n37364 ;
  assign \g9575/_0_  = ~n37367 ;
  assign \g9576/_0_  = ~n37376 ;
  assign \g9577/_0_  = ~n37385 ;
  assign \g9578/_0_  = ~n37388 ;
  assign \g9579/_0_  = ~n37391 ;
  assign \g9580/_0_  = ~n37394 ;
  assign \g9581/_0_  = ~n37398 ;
  assign \g9582/_0_  = ~n37401 ;
  assign \g9583/_0_  = ~n37404 ;
  assign \g9584/_0_  = ~n37407 ;
  assign \g9585/_0_  = ~n37410 ;
  assign \g9586/_0_  = ~n37413 ;
  assign \g9587/_0_  = ~n37416 ;
  assign \g9588/_0_  = ~n37419 ;
  assign \g9589/_0_  = ~n37422 ;
  assign \g9590/_0_  = ~n37425 ;
  assign \g9591/_0_  = ~n37428 ;
  assign \g9592/_0_  = ~n37431 ;
  assign \g9593/_0_  = ~n37434 ;
  assign \g9594/_0_  = ~n37437 ;
  assign \g9595/_0_  = ~n37441 ;
  assign \g9596/_0_  = ~n37444 ;
  assign \g9597/_0_  = ~n37447 ;
  assign \g9598/_0_  = ~n37450 ;
  assign \g9599/_0_  = ~n37453 ;
  assign \g9600/_0_  = ~n37456 ;
  assign \g9601/_0_  = ~n37459 ;
  assign \g9602/_0_  = ~n37462 ;
  assign \g9603/_0_  = ~n37465 ;
  assign \g9604/_0_  = ~n37468 ;
  assign \g9605/_0_  = ~n37471 ;
  assign \g9606/_0_  = ~n37474 ;
  assign \g9607/_0_  = ~n37477 ;
  assign \g9608/_0_  = ~n37480 ;
  assign \g9609/_0_  = ~n37484 ;
  assign \g9610/_0_  = ~n37487 ;
  assign \g9611/_0_  = ~n37490 ;
  assign \g9612/_0_  = ~n37493 ;
  assign \g9613/_0_  = ~n37496 ;
  assign \g9614/_0_  = ~n37499 ;
  assign \g9615/_0_  = ~n37502 ;
  assign \g9616/_0_  = ~n37505 ;
  assign \g9617/_0_  = ~n37508 ;
  assign \g9618/_0_  = ~n37511 ;
  assign \g9619/_0_  = ~n37514 ;
  assign \g9620/_0_  = ~n37517 ;
  assign \g9621/_0_  = ~n37520 ;
  assign \g9622/_0_  = ~n37523 ;
  assign \g9623/_0_  = ~n37527 ;
  assign \g9624/_0_  = ~n37530 ;
  assign \g9625/_0_  = ~n37533 ;
  assign \g9626/_0_  = ~n37536 ;
  assign \g9627/_0_  = ~n37539 ;
  assign \g9628/_0_  = ~n37542 ;
  assign \g9629/_0_  = ~n37545 ;
  assign \g9630/_0_  = ~n37548 ;
  assign \g9631/_0_  = ~n37551 ;
  assign \g9632/_0_  = ~n37554 ;
  assign \g9633/_0_  = ~n37557 ;
  assign \g9634/_0_  = ~n37560 ;
  assign \g9635/_0_  = ~n37563 ;
  assign \g9636/_0_  = ~n37566 ;
  assign \g9637/_0_  = ~n37570 ;
  assign \g9638/_0_  = ~n37573 ;
  assign \g9639/_0_  = ~n37576 ;
  assign \g9640/_0_  = ~n37579 ;
  assign \g9641/_0_  = ~n37582 ;
  assign \g9642/_0_  = ~n37585 ;
  assign \g9643/_0_  = ~n37588 ;
  assign \g9644/_0_  = ~n37591 ;
  assign \g9645/_0_  = ~n37594 ;
  assign \g9646/_0_  = ~n37597 ;
  assign \g9647/_0_  = ~n37600 ;
  assign \g9648/_0_  = ~n37603 ;
  assign \g9649/_0_  = ~n37606 ;
  assign \g9650/_0_  = ~n37609 ;
  assign \g9651/_0_  = ~n37613 ;
  assign \g9652/_0_  = ~n37616 ;
  assign \g9653/_0_  = ~n37619 ;
  assign \g9654/_0_  = ~n37622 ;
  assign \g9655/_0_  = ~n37625 ;
  assign \g9656/_0_  = ~n37628 ;
  assign \g9657/_0_  = ~n37631 ;
  assign \g9658/_0_  = ~n37634 ;
  assign \g9659/_0_  = ~n37637 ;
  assign \g9660/_0_  = ~n37640 ;
  assign \g9661/_0_  = ~n37643 ;
  assign \g9662/_0_  = ~n37646 ;
  assign \g9663/_0_  = ~n37649 ;
  assign \g9664/_0_  = ~n37652 ;
  assign \g9665/_0_  = ~n37656 ;
  assign \g9666/_0_  = ~n37659 ;
  assign \g9667/_0_  = ~n37662 ;
  assign \g9668/_0_  = ~n37665 ;
  assign \g9669/_0_  = ~n37668 ;
  assign \g9670/_0_  = ~n37671 ;
  assign \g9671/_0_  = ~n37674 ;
  assign \g9672/_0_  = ~n37677 ;
  assign \g9673/_0_  = ~n37680 ;
  assign \g9674/_0_  = ~n37683 ;
  assign \g9675/_0_  = ~n37686 ;
  assign \g9676/_0_  = ~n37689 ;
  assign \g9677/_0_  = ~n37692 ;
  assign \g9678/_0_  = ~n37695 ;
  assign \g9681/_0_  = ~n37700 ;
  assign \g9683/_0_  = ~n37703 ;
  assign \g9689/_0_  = n37708 ;
  assign \g9692/_0_  = n37712 ;
  assign \g9694/_0_  = n37717 ;
  assign \g9695/_0_  = n37722 ;
  assign \g9701/_0_  = n37726 ;
  assign \g9702/_0_  = n37731 ;
  assign \g9703/_0_  = n37736 ;
  assign \g9704/_0_  = n37741 ;
  assign \g9709/_0_  = n37745 ;
  assign \g9710/_0_  = n37748 ;
  assign \g9711/_0_  = n37751 ;
  assign \g9712/_0_  = n37754 ;
  assign \g9720/_0_  = ~n37757 ;
  assign \g9721/_0_  = ~n37760 ;
  assign \g9722/_0_  = ~n37763 ;
  assign \g9726/_0_  = ~n37766 ;
  assign \g9733/_0_  = ~n37770 ;
  assign \g9734/_0_  = ~n37773 ;
  assign \g9735/_0_  = ~n37776 ;
  assign \g9736/_0_  = ~n37779 ;
  assign \g9737/_0_  = ~n37782 ;
  assign \g9738/_0_  = ~n37785 ;
  assign \g9739/_0_  = ~n37788 ;
  assign \g9740/_0_  = ~n37791 ;
  assign \g9741/_0_  = ~n37794 ;
  assign \g9742/_0_  = ~n37797 ;
  assign \g9743/_0_  = ~n37800 ;
  assign \g9744/_0_  = ~n37803 ;
  assign \g9745/_0_  = ~n37806 ;
  assign \g9746/_0_  = ~n37809 ;
  assign \g9747/_0_  = ~n37813 ;
  assign \g9748/_0_  = ~n37816 ;
  assign \g9749/_0_  = ~n37819 ;
  assign \g9750/_0_  = ~n37822 ;
  assign \g9751/_0_  = ~n37825 ;
  assign \g9752/_0_  = ~n37828 ;
  assign \g9753/_0_  = ~n37831 ;
  assign \g9754/_0_  = ~n37834 ;
  assign \g9755/_0_  = ~n37837 ;
  assign \g9756/_0_  = ~n37840 ;
  assign \g9757/_0_  = ~n37843 ;
  assign \g9758/_0_  = ~n37846 ;
  assign \g9759/_0_  = ~n37849 ;
  assign \g9760/_0_  = ~n37852 ;
  assign \g9761/_0_  = ~n37856 ;
  assign \g9762/_0_  = ~n37859 ;
  assign \g9763/_0_  = ~n37862 ;
  assign \g9764/_0_  = ~n37865 ;
  assign \g9765/_0_  = ~n37868 ;
  assign \g9766/_0_  = ~n37871 ;
  assign \g9767/_0_  = ~n37874 ;
  assign \g9768/_0_  = ~n37877 ;
  assign \g9769/_0_  = ~n37880 ;
  assign \g9770/_0_  = ~n37883 ;
  assign \g9771/_0_  = ~n37886 ;
  assign \g9772/_0_  = ~n37889 ;
  assign \g9773/_0_  = ~n37892 ;
  assign \g9774/_0_  = ~n37895 ;
  assign \g9775/_0_  = ~n37899 ;
  assign \g9776/_0_  = ~n37902 ;
  assign \g9777/_0_  = ~n37905 ;
  assign \g9778/_0_  = ~n37908 ;
  assign \g9779/_0_  = ~n37911 ;
  assign \g9780/_0_  = ~n37914 ;
  assign \g9781/_0_  = ~n37917 ;
  assign \g9782/_0_  = ~n37920 ;
  assign \g9783/_0_  = ~n37923 ;
  assign \g9784/_0_  = ~n37926 ;
  assign \g9785/_0_  = ~n37929 ;
  assign \g9786/_0_  = ~n37932 ;
  assign \g9787/_0_  = ~n37935 ;
  assign \g9788/_0_  = ~n37938 ;
  assign \g9789/_0_  = ~n37942 ;
  assign \g9790/_0_  = ~n37945 ;
  assign \g9791/_0_  = ~n37948 ;
  assign \g9792/_0_  = ~n37951 ;
  assign \g9793/_0_  = ~n37954 ;
  assign \g9794/_0_  = ~n37957 ;
  assign \g9795/_0_  = ~n37960 ;
  assign \g9796/_0_  = ~n37963 ;
  assign \g9797/_0_  = ~n37966 ;
  assign \g9798/_0_  = ~n37969 ;
  assign \g9799/_0_  = ~n37972 ;
  assign \g9800/_0_  = ~n37975 ;
  assign \g9801/_0_  = ~n37978 ;
  assign \g9802/_0_  = ~n37981 ;
  assign \g9803/_0_  = ~n37985 ;
  assign \g9804/_0_  = ~n37988 ;
  assign \g9805/_0_  = ~n37991 ;
  assign \g9806/_0_  = ~n37994 ;
  assign \g9807/_0_  = ~n37997 ;
  assign \g9808/_0_  = ~n38000 ;
  assign \g9809/_0_  = ~n38003 ;
  assign \g9810/_0_  = ~n38006 ;
  assign \g9811/_0_  = ~n38009 ;
  assign \g9812/_0_  = ~n38012 ;
  assign \g9813/_0_  = ~n38015 ;
  assign \g9814/_0_  = ~n38018 ;
  assign \g9815/_0_  = ~n38021 ;
  assign \g9816/_0_  = ~n38024 ;
  assign \g9817/_0_  = ~n38028 ;
  assign \g9818/_0_  = ~n38031 ;
  assign \g9819/_0_  = ~n38034 ;
  assign \g9820/_0_  = ~n38037 ;
  assign \g9821/_0_  = ~n38040 ;
  assign \g9822/_0_  = ~n38043 ;
  assign \g9823/_0_  = ~n38046 ;
  assign \g9824/_0_  = ~n38049 ;
  assign \g9825/_0_  = ~n38052 ;
  assign \g9826/_0_  = ~n38055 ;
  assign \g9827/_0_  = ~n38058 ;
  assign \g9828/_0_  = ~n38061 ;
  assign \g9829/_0_  = ~n38064 ;
  assign \g9830/_0_  = ~n38067 ;
  assign \g9831/_0_  = ~n38070 ;
  assign \g9832/_0_  = ~n38073 ;
  assign \g9833/_0_  = ~n38076 ;
  assign \g9835/_0_  = n38079 ;
  assign \g9836/_0_  = n38082 ;
  assign \g9837/_0_  = n38085 ;
  assign \g9838/_0_  = n38088 ;
  assign \g9839/_0_  = n38091 ;
  assign \g9840/_0_  = n38094 ;
  assign \g9841/_0_  = n38097 ;
  assign \g9842/_0_  = n38100 ;
  assign \g9844/_0_  = ~n38103 ;
  assign \g9845/_0_  = ~n38106 ;
  assign \g9846/_0_  = ~n38109 ;
  assign \g9848/_0_  = ~n38112 ;
  assign \g9849/_0_  = ~n38115 ;
  assign \g9850/_0_  = n38120 ;
  assign \g9851/_0_  = n38125 ;
  assign \g9853/_0_  = ~n38130 ;
  assign \g9854/_0_  = n38135 ;
  assign \g9855/_0_  = n38140 ;
  assign \g9856/_0_  = n38146 ;
  assign \g9857/_0_  = ~n38149 ;
  assign \g9858/_0_  = ~n38152 ;
  assign \g9859/_0_  = ~n38155 ;
  assign \g9860/_0_  = ~n38158 ;
  assign \g9862/_0_  = ~n38162 ;
  assign \g9863/_0_  = ~n38166 ;
  assign \g9864/_0_  = ~n38170 ;
  assign \g9865/_0_  = ~n38174 ;
  assign \g9867/_0_  = ~n38179 ;
  assign \g9868/_0_  = ~n38182 ;
  assign \g9876/_0_  = ~n38185 ;
  assign \g9877/_0_  = ~n38188 ;
  assign \g9878/_0_  = ~n38191 ;
  assign \g9879/_0_  = ~n38194 ;
  assign \g9880/_0_  = ~n38197 ;
  assign \g9881/_0_  = ~n38200 ;
  assign \g9898/_0_  = ~n38204 ;
  assign \g9900/_0_  = ~n38207 ;
  assign \g9901/_0_  = ~n38210 ;
  assign \g9902/_0_  = ~n38213 ;
  assign \g9903/_0_  = ~n38216 ;
  assign \g9904/_0_  = ~n38219 ;
  assign \g9905/_0_  = ~n38222 ;
  assign \g9906/_0_  = ~n38225 ;
  assign \g9907/_0_  = ~n38228 ;
  assign \g9908/_0_  = ~n38231 ;
  assign \g9909/_0_  = ~n38234 ;
  assign \g9910/_0_  = ~n38237 ;
  assign \g9911/_0_  = ~n38240 ;
  assign \g9912/_0_  = ~n38243 ;
  assign \g9913/_0_  = ~n38246 ;
  assign \g9914/_0_  = ~n38249 ;
  assign \g9915/_0_  = ~n38252 ;
  assign \g9916/_0_  = ~n38255 ;
  assign \g9917/_0_  = ~n38258 ;
  assign \g9918/_0_  = ~n38261 ;
  assign \g9919/_0_  = ~n38264 ;
  assign \g992/_0_  = ~n38279 ;
  assign \g9920/_0_  = ~n38282 ;
  assign \g9921/_0_  = ~n38285 ;
  assign \g9922/_0_  = ~n38288 ;
  assign \g9923/_0_  = ~n38291 ;
  assign \g9924/_0_  = ~n38295 ;
  assign \g9925/_0_  = ~n38298 ;
  assign \g9926/_0_  = ~n38301 ;
  assign \g9927/_0_  = ~n38304 ;
  assign \g9928/_0_  = ~n38307 ;
  assign \g9929/_0_  = ~n38310 ;
  assign \g9930/_0_  = ~n38313 ;
  assign \g9931/_0_  = ~n38316 ;
  assign \g9932/_0_  = ~n38319 ;
  assign \g9933/_0_  = ~n38322 ;
  assign \g9934/_0_  = ~n38325 ;
  assign \g9935/_0_  = ~n38328 ;
  assign \g9936/_0_  = ~n38331 ;
  assign \g9937/_0_  = ~n38334 ;
  assign \g9938/_0_  = ~n38337 ;
  assign \g9939/_0_  = ~n38340 ;
  assign \g9940/_0_  = ~n38343 ;
  assign \g9941/_0_  = ~n38346 ;
  assign \g9942/_0_  = ~n38349 ;
  assign \g9943/_0_  = ~n38352 ;
  assign \g9944/_0_  = ~n38355 ;
  assign \g9945/_0_  = ~n38358 ;
  assign \g9946/_0_  = ~n38361 ;
  assign \g9947/_0_  = ~n38364 ;
  assign \g9948/_0_  = ~n38367 ;
  assign \g9949/_0_  = ~n38371 ;
  assign \g9950/_0_  = ~n38374 ;
  assign \g9951/_0_  = ~n38377 ;
  assign \g9952/_0_  = ~n38380 ;
  assign \g9953/_0_  = ~n38383 ;
  assign \g9954/_0_  = ~n38386 ;
  assign \g9955/_0_  = ~n38389 ;
  assign \g9956/_0_  = ~n38392 ;
  assign \g9957/_0_  = ~n38395 ;
  assign \g9958/_0_  = ~n38398 ;
  assign \g9959/_0_  = ~n38401 ;
  assign \g9960/_0_  = ~n38404 ;
  assign \g9961/_0_  = ~n38407 ;
  assign \g9962/_0_  = ~n38410 ;
  assign \g9963/_0_  = ~n38413 ;
  assign \g9964/_0_  = ~n38416 ;
  assign \g9965/_0_  = ~n38419 ;
  assign \g9966/_0_  = ~n38422 ;
  assign \g9967/_0_  = ~n38425 ;
  assign \g9968/_0_  = ~n38428 ;
  assign \g9969/_0_  = ~n38431 ;
  assign \g9970/_0_  = ~n38434 ;
  assign \g9971/_0_  = ~n38437 ;
  assign \g9972/_0_  = ~n38440 ;
  assign \g9973/_0_  = ~n38443 ;
  assign \g9974/_0_  = ~n38446 ;
  assign \g9975/_0_  = ~n38449 ;
  assign \g9976/_0_  = ~n38452 ;
  assign \g9977/_0_  = ~n38455 ;
  assign \g9978/_0_  = ~n38458 ;
  assign \g9979/_0_  = ~n38461 ;
  assign \g9980/_0_  = ~n38464 ;
  assign \g9981/_0_  = ~n38467 ;
  assign \g9982/_0_  = ~n38470 ;
  assign \g9983/_0_  = ~n38473 ;
  assign \g9984/_0_  = ~n38476 ;
  assign \g9985/_0_  = ~n38479 ;
  assign \g9987/_0_  = ~n38482 ;
  assign \g9988/_0_  = ~n38485 ;
  assign \g9989/_0_  = ~n38488 ;
  assign \g999/_0_  = n38491 ;
  assign \g9990/_0_  = ~n38494 ;
  assign \g9991/_0_  = ~n38497 ;
  assign \g9992/_0_  = ~n38500 ;
  assign \g9993/_0_  = ~n38503 ;
  assign \g9994/_0_  = ~n38506 ;
  assign \g9995/_0_  = ~n38509 ;
  assign \g9996/_0_  = ~n38512 ;
  assign \g9997/_0_  = ~n38515 ;
  assign \g9998/_0_  = ~n38518 ;
  assign \g9999/_0_  = ~n38521 ;
  assign \idma_IDMA_boot_reg/NET0131_reg_syn_3  = ~n38522 ;
  assign \memc_EXTC_Eg_reg/NET0131  = ~n4068 ;
  assign \memc_EXTC_Eg_reg/NET0131_reg_syn_3  = ~n38524 ;
  assign \memc_EXTC_Eg_reg/n0  = n38523 ;
  assign \pio_PIO_IN_P_reg[0]/P0001_reg_syn_3  = ~n38527 ;
  assign \pio_PIO_IN_P_reg[10]/P0001_reg_syn_3  = ~n38530 ;
  assign \pio_PIO_IN_P_reg[11]/P0001_reg_syn_3  = ~n38533 ;
  assign \pio_PIO_IN_P_reg[1]/P0001_reg_syn_3  = ~n38536 ;
  assign \pio_PIO_IN_P_reg[2]/P0001_reg_syn_3  = ~n38539 ;
  assign \pio_PIO_IN_P_reg[3]/P0001_reg_syn_3  = ~n38542 ;
  assign \pio_PIO_IN_P_reg[4]/P0001_reg_syn_3  = ~n38545 ;
  assign \pio_PIO_IN_P_reg[5]/P0001_reg_syn_3  = ~n38548 ;
  assign \pio_PIO_IN_P_reg[6]/P0001_reg_syn_3  = ~n38551 ;
  assign \pio_PIO_IN_P_reg[7]/P0001_reg_syn_3  = ~n38554 ;
  assign \pio_PIO_IN_P_reg[8]/P0001_reg_syn_3  = ~n38557 ;
  assign \pio_PIO_IN_P_reg[9]/P0001_reg_syn_3  = ~n38560 ;
  assign \pio_PIO_RES_OUT_reg[0]/P0001_reg_syn_3  = ~n38563 ;
  assign \pio_PIO_RES_OUT_reg[10]/P0001_reg_syn_3  = ~n38566 ;
  assign \pio_PIO_RES_OUT_reg[2]/P0001_reg_syn_3  = ~n38569 ;
  assign \pio_PIO_RES_OUT_reg[4]/P0001_reg_syn_3  = ~n38572 ;
  assign \pio_PIO_RES_OUT_reg[6]/P0001_reg_syn_3  = ~n38575 ;
  assign \sice_GO_NXi_reg/NET0131_reg_syn_3  = ~n38578 ;
  assign \sport0_rxctl_RXSHT_reg[0]/P0001_reg_syn_3  = n38581 ;
  assign \sport0_rxctl_RXSHT_reg[1]/P0001_reg_syn_3  = ~n38583 ;
  assign \sport1_rxctl_RXSHT_reg[0]/P0001_reg_syn_3  = n38586 ;
  assign \sport1_rxctl_RXSHT_reg[1]/P0001_reg_syn_3  = ~n38588 ;
endmodule
