module top (dma_ack_o_pad, dma_nd_i_pad, dma_req_i_pad, \u0_csr_r_reg[0]/NET0131 , \u0_int_maska_r_reg[0]/NET0131 , \u0_int_maska_r_reg[10]/NET0131 , \u0_int_maska_r_reg[11]/NET0131 , \u0_int_maska_r_reg[12]/NET0131 , \u0_int_maska_r_reg[13]/NET0131 , \u0_int_maska_r_reg[14]/NET0131 , \u0_int_maska_r_reg[15]/NET0131 , \u0_int_maska_r_reg[16]/NET0131 , \u0_int_maska_r_reg[17]/NET0131 , \u0_int_maska_r_reg[18]/NET0131 , \u0_int_maska_r_reg[19]/NET0131 , \u0_int_maska_r_reg[1]/NET0131 , \u0_int_maska_r_reg[20]/NET0131 , \u0_int_maska_r_reg[21]/NET0131 , \u0_int_maska_r_reg[22]/NET0131 , \u0_int_maska_r_reg[23]/NET0131 , \u0_int_maska_r_reg[24]/NET0131 , \u0_int_maska_r_reg[25]/NET0131 , \u0_int_maska_r_reg[26]/NET0131 , \u0_int_maska_r_reg[27]/NET0131 , \u0_int_maska_r_reg[28]/NET0131 , \u0_int_maska_r_reg[29]/NET0131 , \u0_int_maska_r_reg[2]/NET0131 , \u0_int_maska_r_reg[30]/NET0131 , \u0_int_maska_r_reg[3]/NET0131 , \u0_int_maska_r_reg[4]/NET0131 , \u0_int_maska_r_reg[5]/NET0131 , \u0_int_maska_r_reg[6]/NET0131 , \u0_int_maska_r_reg[7]/NET0131 , \u0_int_maska_r_reg[8]/NET0131 , \u0_int_maska_r_reg[9]/NET0131 , \u0_int_maskb_r_reg[0]/NET0131 , \u0_int_maskb_r_reg[10]/NET0131 , \u0_int_maskb_r_reg[11]/NET0131 , \u0_int_maskb_r_reg[12]/NET0131 , \u0_int_maskb_r_reg[13]/NET0131 , \u0_int_maskb_r_reg[14]/NET0131 , \u0_int_maskb_r_reg[15]/NET0131 , \u0_int_maskb_r_reg[16]/NET0131 , \u0_int_maskb_r_reg[17]/NET0131 , \u0_int_maskb_r_reg[18]/NET0131 , \u0_int_maskb_r_reg[19]/NET0131 , \u0_int_maskb_r_reg[1]/NET0131 , \u0_int_maskb_r_reg[20]/NET0131 , \u0_int_maskb_r_reg[21]/NET0131 , \u0_int_maskb_r_reg[22]/NET0131 , \u0_int_maskb_r_reg[23]/NET0131 , \u0_int_maskb_r_reg[24]/NET0131 , \u0_int_maskb_r_reg[25]/NET0131 , \u0_int_maskb_r_reg[26]/NET0131 , \u0_int_maskb_r_reg[27]/NET0131 , \u0_int_maskb_r_reg[28]/NET0131 , \u0_int_maskb_r_reg[29]/NET0131 , \u0_int_maskb_r_reg[2]/NET0131 , \u0_int_maskb_r_reg[30]/NET0131 , \u0_int_maskb_r_reg[3]/NET0131 , \u0_int_maskb_r_reg[4]/NET0131 , \u0_int_maskb_r_reg[5]/NET0131 , \u0_int_maskb_r_reg[6]/NET0131 , \u0_int_maskb_r_reg[7]/NET0131 , \u0_int_maskb_r_reg[8]/NET0131 , \u0_int_maskb_r_reg[9]/NET0131 , \u0_u0_ch_adr0_r_reg[0]/P0001 , \u0_u0_ch_adr0_r_reg[10]/P0001 , \u0_u0_ch_adr0_r_reg[11]/P0001 , \u0_u0_ch_adr0_r_reg[12]/P0001 , \u0_u0_ch_adr0_r_reg[13]/P0001 , \u0_u0_ch_adr0_r_reg[14]/P0001 , \u0_u0_ch_adr0_r_reg[15]/P0001 , \u0_u0_ch_adr0_r_reg[16]/P0001 , \u0_u0_ch_adr0_r_reg[17]/P0001 , \u0_u0_ch_adr0_r_reg[18]/P0001 , \u0_u0_ch_adr0_r_reg[19]/P0001 , \u0_u0_ch_adr0_r_reg[1]/P0001 , \u0_u0_ch_adr0_r_reg[20]/P0001 , \u0_u0_ch_adr0_r_reg[21]/P0001 , \u0_u0_ch_adr0_r_reg[22]/P0001 , \u0_u0_ch_adr0_r_reg[23]/P0001 , \u0_u0_ch_adr0_r_reg[24]/P0001 , \u0_u0_ch_adr0_r_reg[25]/P0001 , \u0_u0_ch_adr0_r_reg[26]/P0001 , \u0_u0_ch_adr0_r_reg[27]/P0001 , \u0_u0_ch_adr0_r_reg[28]/P0001 , \u0_u0_ch_adr0_r_reg[29]/P0001 , \u0_u0_ch_adr0_r_reg[2]/P0001 , \u0_u0_ch_adr0_r_reg[3]/P0001 , \u0_u0_ch_adr0_r_reg[4]/P0001 , \u0_u0_ch_adr0_r_reg[5]/P0001 , \u0_u0_ch_adr0_r_reg[6]/P0001 , \u0_u0_ch_adr0_r_reg[7]/P0001 , \u0_u0_ch_adr0_r_reg[8]/P0001 , \u0_u0_ch_adr0_r_reg[9]/P0001 , \u0_u0_ch_adr1_r_reg[0]/P0001 , \u0_u0_ch_adr1_r_reg[10]/P0001 , \u0_u0_ch_adr1_r_reg[11]/P0001 , \u0_u0_ch_adr1_r_reg[12]/P0001 , \u0_u0_ch_adr1_r_reg[13]/P0001 , \u0_u0_ch_adr1_r_reg[14]/P0001 , \u0_u0_ch_adr1_r_reg[15]/P0001 , \u0_u0_ch_adr1_r_reg[16]/P0001 , \u0_u0_ch_adr1_r_reg[17]/P0001 , \u0_u0_ch_adr1_r_reg[18]/P0001 , \u0_u0_ch_adr1_r_reg[19]/P0001 , \u0_u0_ch_adr1_r_reg[1]/P0001 , \u0_u0_ch_adr1_r_reg[20]/P0001 , \u0_u0_ch_adr1_r_reg[21]/P0001 , \u0_u0_ch_adr1_r_reg[22]/P0001 , \u0_u0_ch_adr1_r_reg[23]/P0001 , \u0_u0_ch_adr1_r_reg[24]/P0001 , \u0_u0_ch_adr1_r_reg[25]/P0001 , \u0_u0_ch_adr1_r_reg[26]/P0001 , \u0_u0_ch_adr1_r_reg[27]/P0001 , \u0_u0_ch_adr1_r_reg[28]/P0001 , \u0_u0_ch_adr1_r_reg[29]/P0001 , \u0_u0_ch_adr1_r_reg[2]/P0001 , \u0_u0_ch_adr1_r_reg[3]/P0001 , \u0_u0_ch_adr1_r_reg[4]/P0001 , \u0_u0_ch_adr1_r_reg[5]/P0001 , \u0_u0_ch_adr1_r_reg[6]/P0001 , \u0_u0_ch_adr1_r_reg[7]/P0001 , \u0_u0_ch_adr1_r_reg[8]/P0001 , \u0_u0_ch_adr1_r_reg[9]/P0001 , \u0_u0_ch_busy_reg/P0001 , \u0_u0_ch_chk_sz_r_reg[0]/P0001 , \u0_u0_ch_chk_sz_r_reg[10]/P0001 , \u0_u0_ch_chk_sz_r_reg[1]/P0001 , \u0_u0_ch_chk_sz_r_reg[2]/P0001 , \u0_u0_ch_chk_sz_r_reg[3]/P0001 , \u0_u0_ch_chk_sz_r_reg[4]/P0001 , \u0_u0_ch_chk_sz_r_reg[5]/P0001 , \u0_u0_ch_chk_sz_r_reg[6]/P0001 , \u0_u0_ch_chk_sz_r_reg[7]/P0001 , \u0_u0_ch_chk_sz_r_reg[8]/P0001 , \u0_u0_ch_chk_sz_r_reg[9]/P0001 , \u0_u0_ch_csr_r2_reg[0]/NET0131 , \u0_u0_ch_csr_r2_reg[1]/NET0131 , \u0_u0_ch_csr_r2_reg[2]/NET0131 , \u0_u0_ch_csr_r3_reg[0]/NET0131 , \u0_u0_ch_csr_r3_reg[1]/NET0131 , \u0_u0_ch_csr_r3_reg[2]/NET0131 , \u0_u0_ch_csr_r_reg[0]/NET0131 , \u0_u0_ch_csr_r_reg[1]/NET0131 , \u0_u0_ch_csr_r_reg[2]/NET0131 , \u0_u0_ch_csr_r_reg[3]/NET0131 , \u0_u0_ch_csr_r_reg[4]/NET0131 , \u0_u0_ch_csr_r_reg[5]/NET0131 , \u0_u0_ch_csr_r_reg[6]/NET0131 , \u0_u0_ch_csr_r_reg[7]/NET0131 , \u0_u0_ch_csr_r_reg[8]/NET0131 , \u0_u0_ch_done_reg/P0002 , \u0_u0_ch_err_reg/NET0131 , \u0_u0_ch_stop_reg/P0001 , \u0_u0_ch_sz_inf_reg/NET0131 , \u0_u0_ch_tot_sz_r_reg[0]/P0001 , \u0_u0_ch_tot_sz_r_reg[10]/P0001 , \u0_u0_ch_tot_sz_r_reg[11]/P0001 , \u0_u0_ch_tot_sz_r_reg[1]/P0001 , \u0_u0_ch_tot_sz_r_reg[2]/P0001 , \u0_u0_ch_tot_sz_r_reg[3]/P0001 , \u0_u0_ch_tot_sz_r_reg[4]/P0001 , \u0_u0_ch_tot_sz_r_reg[5]/P0001 , \u0_u0_ch_tot_sz_r_reg[6]/P0001 , \u0_u0_ch_tot_sz_r_reg[7]/P0001 , \u0_u0_ch_tot_sz_r_reg[8]/P0001 , \u0_u0_ch_tot_sz_r_reg[9]/P0001 , \u0_u0_int_src_r_reg[1]/NET0131 , \u0_u0_int_src_r_reg[2]/NET0131 , \u0_u0_rest_en_reg/NET0131 , \u0_wb_rf_dout_reg[0]/P0001 , \u0_wb_rf_dout_reg[10]/P0001 , \u0_wb_rf_dout_reg[11]/P0001 , \u0_wb_rf_dout_reg[12]/P0001 , \u0_wb_rf_dout_reg[13]/P0001 , \u0_wb_rf_dout_reg[14]/P0001 , \u0_wb_rf_dout_reg[15]/P0001 , \u0_wb_rf_dout_reg[16]/P0001 , \u0_wb_rf_dout_reg[17]/P0001 , \u0_wb_rf_dout_reg[18]/P0001 , \u0_wb_rf_dout_reg[19]/P0001 , \u0_wb_rf_dout_reg[1]/P0001 , \u0_wb_rf_dout_reg[20]/P0001 , \u0_wb_rf_dout_reg[21]/P0001 , \u0_wb_rf_dout_reg[22]/P0001 , \u0_wb_rf_dout_reg[23]/P0001 , \u0_wb_rf_dout_reg[24]/P0001 , \u0_wb_rf_dout_reg[25]/P0001 , \u0_wb_rf_dout_reg[26]/P0001 , \u0_wb_rf_dout_reg[27]/P0001 , \u0_wb_rf_dout_reg[28]/P0001 , \u0_wb_rf_dout_reg[29]/P0001 , \u0_wb_rf_dout_reg[2]/P0001 , \u0_wb_rf_dout_reg[30]/P0001 , \u0_wb_rf_dout_reg[31]/P0001 , \u0_wb_rf_dout_reg[3]/P0001 , \u0_wb_rf_dout_reg[4]/P0001 , \u0_wb_rf_dout_reg[5]/P0001 , \u0_wb_rf_dout_reg[6]/P0001 , \u0_wb_rf_dout_reg[7]/P0001 , \u0_wb_rf_dout_reg[8]/P0001 , \u0_wb_rf_dout_reg[9]/P0001 , \u1_de_start_r_reg/P0001 , \u1_ndnr_reg[0]/P0001 , \u1_ndr_r_reg[0]/NET0131 , \u1_next_start_reg/P0001 , \u1_req_r_reg[0]/P0001 , \u2_adr0_cnt_reg[0]/P0001 , \u2_adr0_cnt_reg[10]/P0001 , \u2_adr0_cnt_reg[11]/P0001 , \u2_adr0_cnt_reg[12]/P0001 , \u2_adr0_cnt_reg[13]/P0001 , \u2_adr0_cnt_reg[14]/P0001 , \u2_adr0_cnt_reg[15]/P0001 , \u2_adr0_cnt_reg[16]/NET0131 , \u2_adr0_cnt_reg[17]/P0001 , \u2_adr0_cnt_reg[18]/P0001 , \u2_adr0_cnt_reg[19]/P0001 , \u2_adr0_cnt_reg[1]/P0001 , \u2_adr0_cnt_reg[20]/P0001 , \u2_adr0_cnt_reg[21]/P0001 , \u2_adr0_cnt_reg[22]/P0001 , \u2_adr0_cnt_reg[23]/P0001 , \u2_adr0_cnt_reg[24]/P0001 , \u2_adr0_cnt_reg[25]/P0001 , \u2_adr0_cnt_reg[26]/P0001 , \u2_adr0_cnt_reg[27]/P0001 , \u2_adr0_cnt_reg[28]/P0001 , \u2_adr0_cnt_reg[29]/P0001 , \u2_adr0_cnt_reg[2]/P0001 , \u2_adr0_cnt_reg[3]/P0001 , \u2_adr0_cnt_reg[4]/P0001 , \u2_adr0_cnt_reg[5]/P0001 , \u2_adr0_cnt_reg[6]/P0001 , \u2_adr0_cnt_reg[7]/P0001 , \u2_adr0_cnt_reg[8]/P0001 , \u2_adr0_cnt_reg[9]/P0001 , \u2_adr1_cnt_reg[0]/P0001 , \u2_adr1_cnt_reg[10]/P0001 , \u2_adr1_cnt_reg[11]/P0001 , \u2_adr1_cnt_reg[12]/P0001 , \u2_adr1_cnt_reg[13]/P0001 , \u2_adr1_cnt_reg[14]/P0001 , \u2_adr1_cnt_reg[15]/P0001 , \u2_adr1_cnt_reg[16]/NET0131 , \u2_adr1_cnt_reg[17]/P0001 , \u2_adr1_cnt_reg[18]/P0001 , \u2_adr1_cnt_reg[19]/P0001 , \u2_adr1_cnt_reg[1]/P0001 , \u2_adr1_cnt_reg[20]/P0001 , \u2_adr1_cnt_reg[21]/P0001 , \u2_adr1_cnt_reg[22]/P0001 , \u2_adr1_cnt_reg[23]/P0001 , \u2_adr1_cnt_reg[24]/P0001 , \u2_adr1_cnt_reg[25]/P0001 , \u2_adr1_cnt_reg[26]/P0001 , \u2_adr1_cnt_reg[27]/P0001 , \u2_adr1_cnt_reg[28]/P0001 , \u2_adr1_cnt_reg[29]/P0001 , \u2_adr1_cnt_reg[2]/P0001 , \u2_adr1_cnt_reg[3]/P0001 , \u2_adr1_cnt_reg[4]/P0001 , \u2_adr1_cnt_reg[5]/P0001 , \u2_adr1_cnt_reg[6]/P0001 , \u2_adr1_cnt_reg[7]/P0001 , \u2_adr1_cnt_reg[8]/P0001 , \u2_adr1_cnt_reg[9]/P0001 , \u2_chunk_0_reg/P0001 , \u2_chunk_cnt_is_0_r_reg/P0001 , \u2_chunk_cnt_reg[0]/NET0131 , \u2_chunk_cnt_reg[1]/NET0131 , \u2_chunk_cnt_reg[2]/NET0131 , \u2_chunk_cnt_reg[3]/NET0131 , \u2_chunk_cnt_reg[4]/NET0131 , \u2_chunk_cnt_reg[5]/NET0131 , \u2_chunk_cnt_reg[6]/NET0131 , \u2_chunk_cnt_reg[7]/NET0131 , \u2_chunk_cnt_reg[8]/NET0131 , \u2_chunk_dec_reg/P0001 , \u2_dma_abort_r_reg/NET0131 , \u2_mast0_adr_reg[10]/P0001 , \u2_mast0_adr_reg[11]/P0001 , \u2_mast0_adr_reg[12]/P0001 , \u2_mast0_adr_reg[13]/P0001 , \u2_mast0_adr_reg[14]/P0001 , \u2_mast0_adr_reg[15]/P0001 , \u2_mast0_adr_reg[16]/P0001 , \u2_mast0_adr_reg[17]/P0001 , \u2_mast0_adr_reg[18]/P0001 , \u2_mast0_adr_reg[19]/P0001 , \u2_mast0_adr_reg[20]/P0001 , \u2_mast0_adr_reg[21]/P0001 , \u2_mast0_adr_reg[22]/P0001 , \u2_mast0_adr_reg[23]/P0001 , \u2_mast0_adr_reg[24]/P0001 , \u2_mast0_adr_reg[25]/P0001 , \u2_mast0_adr_reg[26]/P0001 , \u2_mast0_adr_reg[27]/P0001 , \u2_mast0_adr_reg[28]/P0001 , \u2_mast0_adr_reg[29]/P0001 , \u2_mast0_adr_reg[2]/P0001 , \u2_mast0_adr_reg[30]/P0001 , \u2_mast0_adr_reg[31]/P0001 , \u2_mast0_adr_reg[3]/NET0131 , \u2_mast0_adr_reg[4]/P0001 , \u2_mast0_adr_reg[5]/P0001 , \u2_mast0_adr_reg[6]/P0001 , \u2_mast0_adr_reg[7]/P0001 , \u2_mast0_adr_reg[8]/P0001 , \u2_mast0_adr_reg[9]/P0001 , \u2_mast0_drdy_r_reg/P0001 , \u2_mast1_adr_reg[10]/P0001 , \u2_mast1_adr_reg[11]/P0001 , \u2_mast1_adr_reg[12]/P0001 , \u2_mast1_adr_reg[13]/P0001 , \u2_mast1_adr_reg[14]/P0001 , \u2_mast1_adr_reg[15]/P0001 , \u2_mast1_adr_reg[16]/P0001 , \u2_mast1_adr_reg[17]/P0001 , \u2_mast1_adr_reg[18]/P0001 , \u2_mast1_adr_reg[19]/P0001 , \u2_mast1_adr_reg[20]/P0001 , \u2_mast1_adr_reg[21]/P0001 , \u2_mast1_adr_reg[22]/P0001 , \u2_mast1_adr_reg[23]/P0001 , \u2_mast1_adr_reg[24]/P0001 , \u2_mast1_adr_reg[25]/P0001 , \u2_mast1_adr_reg[26]/P0001 , \u2_mast1_adr_reg[27]/P0001 , \u2_mast1_adr_reg[28]/P0001 , \u2_mast1_adr_reg[29]/P0001 , \u2_mast1_adr_reg[2]/P0001 , \u2_mast1_adr_reg[30]/P0001 , \u2_mast1_adr_reg[31]/P0001 , \u2_mast1_adr_reg[3]/P0001 , \u2_mast1_adr_reg[4]/P0001 , \u2_mast1_adr_reg[5]/P0001 , \u2_mast1_adr_reg[6]/P0001 , \u2_mast1_adr_reg[7]/P0001 , \u2_mast1_adr_reg[8]/P0001 , \u2_mast1_adr_reg[9]/P0001 , \u2_next_ch_reg/P0001 , \u2_read_r_reg/P0001 , \u2_state_reg[0]/NET0131 , \u2_state_reg[10]/NET0131 , \u2_state_reg[1]/NET0131 , \u2_state_reg[2]/NET0131 , \u2_state_reg[3]/NET0131 , \u2_state_reg[4]/NET0131 , \u2_state_reg[5]/NET0131 , \u2_state_reg[6]/NET0131 , \u2_state_reg[7]/NET0131 , \u2_state_reg[8]/NET0131 , \u2_state_reg[9]/NET0131 , \u2_tsz_cnt_is_0_r_reg/P0001 , \u2_tsz_cnt_reg[0]/NET0131 , \u2_tsz_cnt_reg[10]/NET0131 , \u2_tsz_cnt_reg[11]/NET0131 , \u2_tsz_cnt_reg[1]/NET0131 , \u2_tsz_cnt_reg[2]/NET0131 , \u2_tsz_cnt_reg[3]/NET0131 , \u2_tsz_cnt_reg[4]/NET0131 , \u2_tsz_cnt_reg[5]/NET0131 , \u2_tsz_cnt_reg[6]/NET0131 , \u2_tsz_cnt_reg[7]/NET0131 , \u2_tsz_cnt_reg[8]/NET0131 , \u2_tsz_cnt_reg[9]/NET0131 , \u2_u0_out_r_reg[0]/P0001 , \u2_u0_out_r_reg[10]/P0001 , \u2_u0_out_r_reg[11]/P0001 , \u2_u0_out_r_reg[12]/P0001 , \u2_u0_out_r_reg[13]/P0001 , \u2_u0_out_r_reg[14]/P0001 , \u2_u0_out_r_reg[15]/P0001 , \u2_u0_out_r_reg[16]/P0001 , \u2_u0_out_r_reg[1]/P0001 , \u2_u0_out_r_reg[2]/P0001 , \u2_u0_out_r_reg[3]/P0001 , \u2_u0_out_r_reg[4]/P0001 , \u2_u0_out_r_reg[5]/P0001 , \u2_u0_out_r_reg[6]/P0001 , \u2_u0_out_r_reg[7]/P0001 , \u2_u0_out_r_reg[8]/P0001 , \u2_u0_out_r_reg[9]/P0001 , \u2_u1_out_r_reg[0]/P0001 , \u2_u1_out_r_reg[10]/P0001 , \u2_u1_out_r_reg[11]/P0001 , \u2_u1_out_r_reg[12]/P0001 , \u2_u1_out_r_reg[13]/P0001 , \u2_u1_out_r_reg[14]/P0001 , \u2_u1_out_r_reg[15]/P0001 , \u2_u1_out_r_reg[16]/P0001 , \u2_u1_out_r_reg[1]/P0001 , \u2_u1_out_r_reg[2]/P0001 , \u2_u1_out_r_reg[3]/P0001 , \u2_u1_out_r_reg[4]/P0001 , \u2_u1_out_r_reg[5]/P0001 , \u2_u1_out_r_reg[6]/P0001 , \u2_u1_out_r_reg[7]/P0001 , \u2_u1_out_r_reg[8]/P0001 , \u2_u1_out_r_reg[9]/P0001 , \u2_write_hold_r_reg/P0001 , \u2_write_r_reg/P0001 , \u3_u0_mast_cyc_reg/P0001 , \u3_u0_mast_dout_reg[0]/P0001 , \u3_u0_mast_dout_reg[10]/P0001 , \u3_u0_mast_dout_reg[11]/P0001 , \u3_u0_mast_dout_reg[12]/P0001 , \u3_u0_mast_dout_reg[13]/P0001 , \u3_u0_mast_dout_reg[14]/P0001 , \u3_u0_mast_dout_reg[15]/P0001 , \u3_u0_mast_dout_reg[16]/P0001 , \u3_u0_mast_dout_reg[17]/P0001 , \u3_u0_mast_dout_reg[18]/P0001 , \u3_u0_mast_dout_reg[19]/P0001 , \u3_u0_mast_dout_reg[1]/P0001 , \u3_u0_mast_dout_reg[20]/P0001 , \u3_u0_mast_dout_reg[21]/P0001 , \u3_u0_mast_dout_reg[22]/P0001 , \u3_u0_mast_dout_reg[23]/P0001 , \u3_u0_mast_dout_reg[24]/P0001 , \u3_u0_mast_dout_reg[25]/P0001 , \u3_u0_mast_dout_reg[26]/P0001 , \u3_u0_mast_dout_reg[27]/P0001 , \u3_u0_mast_dout_reg[28]/P0001 , \u3_u0_mast_dout_reg[29]/P0001 , \u3_u0_mast_dout_reg[2]/P0001 , \u3_u0_mast_dout_reg[30]/P0001 , \u3_u0_mast_dout_reg[31]/P0001 , \u3_u0_mast_dout_reg[3]/P0001 , \u3_u0_mast_dout_reg[4]/P0001 , \u3_u0_mast_dout_reg[5]/P0001 , \u3_u0_mast_dout_reg[6]/P0001 , \u3_u0_mast_dout_reg[7]/P0001 , \u3_u0_mast_dout_reg[8]/P0001 , \u3_u0_mast_dout_reg[9]/P0001 , \u3_u0_mast_stb_reg/P0001 , \u3_u0_mast_we_r_reg/P0002 , \u3_u1_rf_ack_reg/P0001 , \u3_u1_slv_adr_reg[2]/NET0131 , \u3_u1_slv_adr_reg[3]/P0001 , \u3_u1_slv_adr_reg[4]/NET0131 , \u3_u1_slv_adr_reg[5]/P0001 , \u3_u1_slv_adr_reg[6]/NET0131 , \u3_u1_slv_adr_reg[7]/NET0131 , \u3_u1_slv_adr_reg[8]/NET0131 , \u3_u1_slv_adr_reg[9]/NET0131 , \u3_u1_slv_dout_reg[0]/P0001 , \u3_u1_slv_dout_reg[10]/P0001 , \u3_u1_slv_dout_reg[11]/P0001 , \u3_u1_slv_dout_reg[12]/P0001 , \u3_u1_slv_dout_reg[13]/P0001 , \u3_u1_slv_dout_reg[14]/P0001 , \u3_u1_slv_dout_reg[15]/P0001 , \u3_u1_slv_dout_reg[16]/P0001 , \u3_u1_slv_dout_reg[17]/P0001 , \u3_u1_slv_dout_reg[18]/P0001 , \u3_u1_slv_dout_reg[19]/P0001 , \u3_u1_slv_dout_reg[1]/P0001 , \u3_u1_slv_dout_reg[20]/P0001 , \u3_u1_slv_dout_reg[21]/P0001 , \u3_u1_slv_dout_reg[22]/P0001 , \u3_u1_slv_dout_reg[23]/P0001 , \u3_u1_slv_dout_reg[24]/P0001 , \u3_u1_slv_dout_reg[25]/P0001 , \u3_u1_slv_dout_reg[26]/P0001 , \u3_u1_slv_dout_reg[27]/P0001 , \u3_u1_slv_dout_reg[28]/P0001 , \u3_u1_slv_dout_reg[29]/P0001 , \u3_u1_slv_dout_reg[2]/P0001 , \u3_u1_slv_dout_reg[30]/P0001 , \u3_u1_slv_dout_reg[31]/P0001 , \u3_u1_slv_dout_reg[3]/P0001 , \u3_u1_slv_dout_reg[4]/P0001 , \u3_u1_slv_dout_reg[5]/P0001 , \u3_u1_slv_dout_reg[6]/P0001 , \u3_u1_slv_dout_reg[7]/P0001 , \u3_u1_slv_dout_reg[8]/P0001 , \u3_u1_slv_dout_reg[9]/P0001 , \u3_u1_slv_re_reg/P0001 , \u3_u1_slv_we_reg/P0001 , \u4_u0_mast_cyc_reg/P0001 , \u4_u0_mast_dout_reg[0]/P0001 , \u4_u0_mast_dout_reg[10]/P0001 , \u4_u0_mast_dout_reg[11]/P0001 , \u4_u0_mast_dout_reg[12]/P0001 , \u4_u0_mast_dout_reg[13]/P0001 , \u4_u0_mast_dout_reg[14]/P0001 , \u4_u0_mast_dout_reg[15]/P0001 , \u4_u0_mast_dout_reg[16]/P0001 , \u4_u0_mast_dout_reg[17]/P0001 , \u4_u0_mast_dout_reg[18]/P0001 , \u4_u0_mast_dout_reg[19]/P0001 , \u4_u0_mast_dout_reg[1]/P0001 , \u4_u0_mast_dout_reg[20]/P0001 , \u4_u0_mast_dout_reg[21]/P0001 , \u4_u0_mast_dout_reg[22]/P0001 , \u4_u0_mast_dout_reg[23]/P0001 , \u4_u0_mast_dout_reg[24]/P0001 , \u4_u0_mast_dout_reg[25]/P0001 , \u4_u0_mast_dout_reg[26]/P0001 , \u4_u0_mast_dout_reg[27]/P0001 , \u4_u0_mast_dout_reg[28]/P0001 , \u4_u0_mast_dout_reg[29]/P0001 , \u4_u0_mast_dout_reg[2]/P0001 , \u4_u0_mast_dout_reg[30]/P0001 , \u4_u0_mast_dout_reg[31]/P0001 , \u4_u0_mast_dout_reg[3]/P0001 , \u4_u0_mast_dout_reg[4]/P0001 , \u4_u0_mast_dout_reg[5]/P0001 , \u4_u0_mast_dout_reg[6]/P0001 , \u4_u0_mast_dout_reg[7]/P0001 , \u4_u0_mast_dout_reg[8]/P0001 , \u4_u0_mast_dout_reg[9]/P0001 , \u4_u0_mast_stb_reg/P0001 , \u4_u0_mast_we_r_reg/P0001 , \u4_u1_rf_ack_reg/P0001 , \u4_u1_slv_re_reg/P0001 , \u4_u1_slv_we_reg/P0001 , \wb0_ack_i_pad , \wb0_addr_i[0]_pad , \wb0_addr_i[10]_pad , \wb0_addr_i[11]_pad , \wb0_addr_i[12]_pad , \wb0_addr_i[13]_pad , \wb0_addr_i[14]_pad , \wb0_addr_i[15]_pad , \wb0_addr_i[16]_pad , \wb0_addr_i[17]_pad , \wb0_addr_i[18]_pad , \wb0_addr_i[19]_pad , \wb0_addr_i[1]_pad , \wb0_addr_i[20]_pad , \wb0_addr_i[21]_pad , \wb0_addr_i[22]_pad , \wb0_addr_i[23]_pad , \wb0_addr_i[24]_pad , \wb0_addr_i[25]_pad , \wb0_addr_i[26]_pad , \wb0_addr_i[27]_pad , \wb0_addr_i[28]_pad , \wb0_addr_i[29]_pad , \wb0_addr_i[2]_pad , \wb0_addr_i[30]_pad , \wb0_addr_i[31]_pad , \wb0_addr_i[3]_pad , \wb0_addr_i[4]_pad , \wb0_addr_i[5]_pad , \wb0_addr_i[6]_pad , \wb0_addr_i[7]_pad , \wb0_addr_i[8]_pad , \wb0_addr_i[9]_pad , \wb0_cyc_i_pad , \wb0_err_i_pad , \wb0_rty_i_pad , \wb0_sel_i[0]_pad , \wb0_sel_i[1]_pad , \wb0_sel_i[2]_pad , \wb0_sel_i[3]_pad , \wb0_stb_i_pad , \wb0_we_i_pad , \wb0m_data_i[0]_pad , \wb0m_data_i[10]_pad , \wb0m_data_i[11]_pad , \wb0m_data_i[12]_pad , \wb0m_data_i[13]_pad , \wb0m_data_i[14]_pad , \wb0m_data_i[15]_pad , \wb0m_data_i[16]_pad , \wb0m_data_i[17]_pad , \wb0m_data_i[18]_pad , \wb0m_data_i[19]_pad , \wb0m_data_i[1]_pad , \wb0m_data_i[20]_pad , \wb0m_data_i[21]_pad , \wb0m_data_i[22]_pad , \wb0m_data_i[23]_pad , \wb0m_data_i[24]_pad , \wb0m_data_i[25]_pad , \wb0m_data_i[26]_pad , \wb0m_data_i[27]_pad , \wb0m_data_i[28]_pad , \wb0m_data_i[29]_pad , \wb0m_data_i[2]_pad , \wb0m_data_i[30]_pad , \wb0m_data_i[31]_pad , \wb0m_data_i[3]_pad , \wb0m_data_i[4]_pad , \wb0m_data_i[5]_pad , \wb0m_data_i[6]_pad , \wb0m_data_i[7]_pad , \wb0m_data_i[8]_pad , \wb0m_data_i[9]_pad , \wb0s_data_i[0]_pad , \wb0s_data_i[10]_pad , \wb0s_data_i[11]_pad , \wb0s_data_i[12]_pad , \wb0s_data_i[13]_pad , \wb0s_data_i[14]_pad , \wb0s_data_i[15]_pad , \wb0s_data_i[16]_pad , \wb0s_data_i[17]_pad , \wb0s_data_i[18]_pad , \wb0s_data_i[19]_pad , \wb0s_data_i[1]_pad , \wb0s_data_i[20]_pad , \wb0s_data_i[21]_pad , \wb0s_data_i[22]_pad , \wb0s_data_i[23]_pad , \wb0s_data_i[24]_pad , \wb0s_data_i[25]_pad , \wb0s_data_i[26]_pad , \wb0s_data_i[27]_pad , \wb0s_data_i[28]_pad , \wb0s_data_i[29]_pad , \wb0s_data_i[2]_pad , \wb0s_data_i[30]_pad , \wb0s_data_i[31]_pad , \wb0s_data_i[3]_pad , \wb0s_data_i[4]_pad , \wb0s_data_i[5]_pad , \wb0s_data_i[6]_pad , \wb0s_data_i[7]_pad , \wb0s_data_i[8]_pad , \wb0s_data_i[9]_pad , \wb1_ack_i_pad , \wb1_addr_i[0]_pad , \wb1_addr_i[10]_pad , \wb1_addr_i[11]_pad , \wb1_addr_i[12]_pad , \wb1_addr_i[13]_pad , \wb1_addr_i[14]_pad , \wb1_addr_i[15]_pad , \wb1_addr_i[16]_pad , \wb1_addr_i[17]_pad , \wb1_addr_i[18]_pad , \wb1_addr_i[19]_pad , \wb1_addr_i[1]_pad , \wb1_addr_i[20]_pad , \wb1_addr_i[21]_pad , \wb1_addr_i[22]_pad , \wb1_addr_i[23]_pad , \wb1_addr_i[24]_pad , \wb1_addr_i[25]_pad , \wb1_addr_i[26]_pad , \wb1_addr_i[27]_pad , \wb1_addr_i[28]_pad , \wb1_addr_i[29]_pad , \wb1_addr_i[2]_pad , \wb1_addr_i[30]_pad , \wb1_addr_i[31]_pad , \wb1_addr_i[3]_pad , \wb1_addr_i[4]_pad , \wb1_addr_i[5]_pad , \wb1_addr_i[6]_pad , \wb1_addr_i[7]_pad , \wb1_addr_i[8]_pad , \wb1_addr_i[9]_pad , \wb1_cyc_i_pad , \wb1_err_i_pad , \wb1_rty_i_pad , \wb1_sel_i[0]_pad , \wb1_sel_i[1]_pad , \wb1_sel_i[2]_pad , \wb1_sel_i[3]_pad , \wb1_stb_i_pad , \wb1_we_i_pad , \wb1m_data_i[0]_pad , \wb1m_data_i[10]_pad , \wb1m_data_i[11]_pad , \wb1m_data_i[12]_pad , \wb1m_data_i[13]_pad , \wb1m_data_i[14]_pad , \wb1m_data_i[15]_pad , \wb1m_data_i[16]_pad , \wb1m_data_i[17]_pad , \wb1m_data_i[18]_pad , \wb1m_data_i[19]_pad , \wb1m_data_i[1]_pad , \wb1m_data_i[20]_pad , \wb1m_data_i[21]_pad , \wb1m_data_i[22]_pad , \wb1m_data_i[23]_pad , \wb1m_data_i[24]_pad , \wb1m_data_i[25]_pad , \wb1m_data_i[26]_pad , \wb1m_data_i[27]_pad , \wb1m_data_i[28]_pad , \wb1m_data_i[29]_pad , \wb1m_data_i[2]_pad , \wb1m_data_i[30]_pad , \wb1m_data_i[31]_pad , \wb1m_data_i[3]_pad , \wb1m_data_i[4]_pad , \wb1m_data_i[5]_pad , \wb1m_data_i[6]_pad , \wb1m_data_i[7]_pad , \wb1m_data_i[8]_pad , \wb1m_data_i[9]_pad , \wb1s_data_i[0]_pad , \wb1s_data_i[10]_pad , \wb1s_data_i[11]_pad , \wb1s_data_i[12]_pad , \wb1s_data_i[13]_pad , \wb1s_data_i[14]_pad , \wb1s_data_i[15]_pad , \wb1s_data_i[16]_pad , \wb1s_data_i[17]_pad , \wb1s_data_i[18]_pad , \wb1s_data_i[19]_pad , \wb1s_data_i[1]_pad , \wb1s_data_i[20]_pad , \wb1s_data_i[21]_pad , \wb1s_data_i[22]_pad , \wb1s_data_i[23]_pad , \wb1s_data_i[24]_pad , \wb1s_data_i[25]_pad , \wb1s_data_i[26]_pad , \wb1s_data_i[27]_pad , \wb1s_data_i[28]_pad , \wb1s_data_i[29]_pad , \wb1s_data_i[2]_pad , \wb1s_data_i[30]_pad , \wb1s_data_i[31]_pad , \wb1s_data_i[3]_pad , \wb1s_data_i[4]_pad , \wb1s_data_i[5]_pad , \wb1s_data_i[6]_pad , \wb1s_data_i[7]_pad , \wb1s_data_i[8]_pad , \wb1s_data_i[9]_pad , \_al_n0 , \_al_n1 , \g22594/_0_ , \g22595/_0_ , \g22599/_0_ , \g22600/_0_ , \g22606/_0_ , \g22607/_0_ , \g22610/_0_ , \g22614/_0_ , \g22615/_0_ , \g22616/_0_ , \g22619/_0_ , \g22620/_0_ , \g22626/_0_ , \g22635/_0_ , \g22650/_0_ , \g22651/_0_ , \g22692/_0_ , \g22727/_0_ , \g22729/_3_ , \g22774/_0_ , \g22775/_0_ , \g22776/_0_ , \g22777/_0_ , \g22779/_3_ , \g22780/_0_ , \g22781/_0_ , \g22782/_0_ , \g22784/_0_ , \g22785/_0_ , \g22786/_0_ , \g22787/_0_ , \g22789/_3_ , \g22790/_0_ , \g22791/_0_ , \g22792/_0_ , \g22793/_0_ , \g22794/_0_ , \g22795/_0_ , \g22796/_0_ , \g22797/_0_ , \g22798/_0_ , \g22799/_0_ , \g22838/_0_ , \g22839/_0_ , \g22841/_0_ , \g22842/_0_ , \g22847/_0_ , \g22848/_0_ , \g22849/_0_ , \g22850/_0_ , \g22851/_0_ , \g22852/_0_ , \g22853/_0_ , \g22854/_0_ , \g22855/_0_ , \g22856/_0_ , \g22857/_0_ , \g22858/_0_ , \g22859/_0_ , \g22860/_0_ , \g22861/_0_ , \g22862/_0_ , \g22863/_0_ , \g22864/_0_ , \g22865/_0_ , \g22867/_0_ , \g22868/_0_ , \g22869/_0_ , \g22871/_0_ , \g22872/_0_ , \g22873/_0_ , \g22874/_0_ , \g22875/_0_ , \g22876/_0_ , \g22878/_0_ , \g22882/_2_ , \g22995/_0_ , \g23030/_0_ , \g23046/_0_ , \g23077/_0_ , \g23111/_0_ , \g23115/_1_ , \g23124/_2_ , \g23126/_2_ , \g23128/_2_ , \g23130/_2_ , \g23132/_2_ , \g23134/_2_ , \g23136/_2_ , \g23137/_0_ , \g23140/_2_ , \g23142/_2_ , \g23144/_2_ , \g23146/_2_ , \g23148/_2_ , \g23150/_2_ , \g23152/_2_ , \g23154/_2_ , \g23156/_2_ , \g23158/_2_ , \g23160/_2_ , \g23162/_2_ , \g23163/_3_ , \g23164/_0_ , \g23166/_0_ , \g23168/_0_ , \g23170/_2_ , \g23172/_2_ , \g23174/_2_ , \g23175/_0_ , \g23177/_0_ , \g23180/_2_ , \g23220/_0_ , \g23238/_0_ , \g23239/_0_ , \g23240/_0_ , \g23241/_0_ , \g23242/_0_ , \g23243/_0_ , \g23244/_0_ , \g23245/_0_ , \g23247/_3_ , \g23248/_0_ , \g23249/_0_ , \g23250/_0_ , \g23251/_0_ , \g23252/_0_ , \g23253/_0_ , \g23255/_3_ , \g23260/_0_ , \g23284/_3_ , \g23285/_0_ , \g23334/_0_ , \g23343/_0_ , \g23366/_0_ , \g23402/_0_ , \g23403/_0_ , \g23404/_0_ , \g23405/_0_ , \g23407/_0_ , \g23408/_0_ , \g23409/_0_ , \g23410/_0_ , \g23411/_0_ , \g23413/_2_ , \g23415/_2_ , \g23417/_2_ , \g23542/_0_ , \g23607/_0_ , \g23608/_0_ , \g23609/_3_ , \g23707/_0_ , \g23708/_0_ , \g23709/_0_ , \g23710/_0_ , \g23711/_0_ , \g23712/_0_ , \g23713/_0_ , \g23714/_0_ , \g23715/_0_ , \g23716/_0_ , \g23754/_0_ , \g23755/_0_ , \g23756/_0_ , \g23757/_0_ , \g23758/_0_ , \g23759/_0_ , \g23760/_0_ , \g23761/_0_ , \g23763/_3_ , \g23767/_0_ , \g23768/_0_ , \g23833/_0_ , \g23837/_0_ , \g23838/_0_ , \g23839/_0_ , \g23840/_0_ , \g23841/_0_ , \g23842/_0_ , \g23843/_0_ , \g23844/_0_ , \g23845/_0_ , \g23849/_3_ , \g23851/_3_ , \g23858/_0_ , \g23870/_0_ , \g23871/_0_ , \g23872/_3_ , \g23873/_3_ , \g23874/_3_ , \g23875/_3_ , \g23876/_3_ , \g23877/_3_ , \g23878/_3_ , \g23879/_3_ , \g23880/_3_ , \g23881/_3_ , \g23882/_3_ , \g23883/_3_ , \g23884/_3_ , \g23885/_3_ , \g23886/_3_ , \g23887/_3_ , \g23888/_3_ , \g23889/_3_ , \g23890/_3_ , \g23891/_3_ , \g23892/_3_ , \g23893/_3_ , \g23894/_3_ , \g23895/_3_ , \g23896/_3_ , \g23897/_3_ , \g23898/_3_ , \g23899/_3_ , \g23900/_3_ , \g23901/_3_ , \g23902/_3_ , \g23903/_3_ , \g23904/_3_ , \g23905/_3_ , \g23906/_3_ , \g23907/_3_ , \g23908/_3_ , \g23909/_3_ , \g23910/_3_ , \g23911/_3_ , \g23912/_3_ , \g23913/_3_ , \g23914/_3_ , \g23915/_3_ , \g23959/_0_ , \g23961/_0_ , \g23962/_0_ , \g23966/_0_ , \g23967/_0_ , \g23969/_0_ , \g23970/_0_ , \g23971/_0_ , \g23972/_0_ , \g23979/_0_ , \g23987/_0_ , \g23988/_0_ , \g23989/_0_ , \g23990/_0_ , \g24005/_0_ , \g24010/_0_ , \g24012/_0_ , \g24013/_0_ , \g24014/_0_ , \g24015/_0_ , \g24016/_0_ , \g24017/_0_ , \g24018/_0_ , \g24019/_0_ , \g24020/_0_ , \g24026/_0_ , \g24027/_0_ , \g24028/_0_ , \g24029/_0_ , \g24030/_0_ , \g24031/_0_ , \g24032/_0_ , \g24033/_0_ , \g24034/_0_ , \g24035/_0_ , \g24036/_0_ , \g24037/_0_ , \g24038/_0_ , \g24039/_0_ , \g24042/_0_ , \g24049/_0_ , \g24063/_0_ , \g24119/_0_ , \g24120/_0_ , \g24357/_0_ , \g24432/_0_ , \g24433/_0_ , \g24437/_0_ , \g24438/_0_ , \g24477/_0_ , \g24491/_0_ , \g24530/_2_ , \g24532/_0_ , \g24534/_0_ , \g24537/_0_ , \g24538/_0_ , \g24539/_0_ , \g24540/_0_ , \g24606/_2_ , \g24612/_0_ , \g24677/_0_ , \g24678/_0_ , \g24679/_0_ , \g24688/_0_ , \g24743/_0_ , \g24847/_0_ , \g24849/_0_ , \g24850/_0_ , \g24854/_0_ , \g24862/_0_ , \g24872/_0_ , \g24873/_0_ , \g24874/_0_ , \g24876/_0_ , \g24879/_0_ , \g24880/_0_ , \g24881/_0_ , \g24882/_0_ , \g24952/_2_ , \g24976/_1_ , \g25003/_0_ , \g25004/_0_ , \g25005/_0_ , \g25006/_0_ , \g25011/_0_ , \g25012/_0_ , \g25013/_0_ , \g25031/_0_ , \g25032/_0_ , \g25033/_0_ , \g25034/_0_ , \g25035/_0_ , \g25153/_2_ , \g25183/_0_ , \g25184/_0_ , \g25224/_0_ , \g25232/_0_ , \g25237/_0_ , \g25241/_2_ , \g25243/_2_ , \g25248/_3_ , \g25261/_0_ , \g25262/_0_ , \g25266/_3_ , \g25267/_0_ , \g25269/_0_ , \g25543/_1_ , \g25602/_3_ , \g25610/_0_ , \g25611/_0_ , \g25841/_0_ , \g25843/_0_ , \g25893/_0_ , \g27013/_0_ , \g27060/_0_ , \g27073/_0_ , \g27184/_0_ , \g27186/_0_ , \g27189/_2_ , \g47/_0_ , \u0_u0_ch_done_reg/_05_ , \u2_adr0_cnt_reg[0]/P0000 , \u2_adr1_cnt_reg[0]/P0000 , \u3_u0_mast_we_r_reg/_05_ , \wb0_ack_o_pad , \wb0_addr_o[0]_pad , \wb0_addr_o[10]_pad , \wb0_addr_o[11]_pad , \wb0_addr_o[12]_pad , \wb0_addr_o[13]_pad , \wb0_addr_o[14]_pad , \wb0_addr_o[15]_pad , \wb0_addr_o[16]_pad , \wb0_addr_o[17]_pad , \wb0_addr_o[18]_pad , \wb0_addr_o[19]_pad , \wb0_addr_o[1]_pad , \wb0_addr_o[20]_pad , \wb0_addr_o[21]_pad , \wb0_addr_o[22]_pad , \wb0_addr_o[23]_pad , \wb0_addr_o[24]_pad , \wb0_addr_o[25]_pad , \wb0_addr_o[26]_pad , \wb0_addr_o[27]_pad , \wb0_addr_o[28]_pad , \wb0_addr_o[29]_pad , \wb0_addr_o[2]_pad , \wb0_addr_o[30]_pad , \wb0_addr_o[31]_pad , \wb0_addr_o[3]_pad , \wb0_addr_o[4]_pad , \wb0_addr_o[5]_pad , \wb0_addr_o[6]_pad , \wb0_addr_o[7]_pad , \wb0_addr_o[8]_pad , \wb0_addr_o[9]_pad , \wb0_cyc_o_pad , \wb0_err_o_pad , \wb0_rty_o_pad , \wb0_sel_o[0]_pad , \wb0_sel_o[1]_pad , \wb0_sel_o[2]_pad , \wb0_sel_o[3]_pad , \wb0_stb_o_pad , \wb0_we_o_pad , \wb0m_data_o[0]_pad , \wb0m_data_o[10]_pad , \wb0m_data_o[11]_pad , \wb0m_data_o[12]_pad , \wb0m_data_o[13]_pad , \wb0m_data_o[14]_pad , \wb0m_data_o[15]_pad , \wb0m_data_o[16]_pad , \wb0m_data_o[17]_pad , \wb0m_data_o[18]_pad , \wb0m_data_o[19]_pad , \wb0m_data_o[1]_pad , \wb0m_data_o[20]_pad , \wb0m_data_o[21]_pad , \wb0m_data_o[22]_pad , \wb0m_data_o[23]_pad , \wb0m_data_o[24]_pad , \wb0m_data_o[25]_pad , \wb0m_data_o[26]_pad , \wb0m_data_o[27]_pad , \wb0m_data_o[28]_pad , \wb0m_data_o[29]_pad , \wb0m_data_o[2]_pad , \wb0m_data_o[30]_pad , \wb0m_data_o[31]_pad , \wb0m_data_o[3]_pad , \wb0m_data_o[4]_pad , \wb0m_data_o[5]_pad , \wb0m_data_o[6]_pad , \wb0m_data_o[7]_pad , \wb0m_data_o[8]_pad , \wb0m_data_o[9]_pad , \wb0s_data_o[0]_pad , \wb0s_data_o[10]_pad , \wb0s_data_o[11]_pad , \wb0s_data_o[12]_pad , \wb0s_data_o[13]_pad , \wb0s_data_o[14]_pad , \wb0s_data_o[15]_pad , \wb0s_data_o[16]_pad , \wb0s_data_o[17]_pad , \wb0s_data_o[18]_pad , \wb0s_data_o[19]_pad , \wb0s_data_o[1]_pad , \wb0s_data_o[20]_pad , \wb0s_data_o[21]_pad , \wb0s_data_o[22]_pad , \wb0s_data_o[23]_pad , \wb0s_data_o[24]_pad , \wb0s_data_o[25]_pad , \wb0s_data_o[26]_pad , \wb0s_data_o[27]_pad , \wb0s_data_o[28]_pad , \wb0s_data_o[29]_pad , \wb0s_data_o[2]_pad , \wb0s_data_o[30]_pad , \wb0s_data_o[31]_pad , \wb0s_data_o[3]_pad , \wb0s_data_o[4]_pad , \wb0s_data_o[5]_pad , \wb0s_data_o[6]_pad , \wb0s_data_o[7]_pad , \wb0s_data_o[8]_pad , \wb0s_data_o[9]_pad , \wb1_ack_o_pad , \wb1_addr_o[0]_pad , \wb1_addr_o[10]_pad , \wb1_addr_o[11]_pad , \wb1_addr_o[12]_pad , \wb1_addr_o[13]_pad , \wb1_addr_o[14]_pad , \wb1_addr_o[15]_pad , \wb1_addr_o[16]_pad , \wb1_addr_o[17]_pad , \wb1_addr_o[18]_pad , \wb1_addr_o[19]_pad , \wb1_addr_o[1]_pad , \wb1_addr_o[20]_pad , \wb1_addr_o[21]_pad , \wb1_addr_o[22]_pad , \wb1_addr_o[23]_pad , \wb1_addr_o[24]_pad , \wb1_addr_o[25]_pad , \wb1_addr_o[26]_pad , \wb1_addr_o[27]_pad , \wb1_addr_o[28]_pad , \wb1_addr_o[29]_pad , \wb1_addr_o[2]_pad , \wb1_addr_o[30]_pad , \wb1_addr_o[31]_pad , \wb1_addr_o[3]_pad , \wb1_addr_o[4]_pad , \wb1_addr_o[5]_pad , \wb1_addr_o[6]_pad , \wb1_addr_o[7]_pad , \wb1_addr_o[8]_pad , \wb1_addr_o[9]_pad , \wb1_cyc_o_pad , \wb1_err_o_pad , \wb1_rty_o_pad , \wb1_sel_o[0]_pad , \wb1_sel_o[1]_pad , \wb1_sel_o[2]_pad , \wb1_sel_o[3]_pad , \wb1_stb_o_pad , \wb1_we_o_pad , \wb1m_data_o[0]_pad , \wb1m_data_o[10]_pad , \wb1m_data_o[11]_pad , \wb1m_data_o[12]_pad , \wb1m_data_o[13]_pad , \wb1m_data_o[14]_pad , \wb1m_data_o[15]_pad , \wb1m_data_o[16]_pad , \wb1m_data_o[17]_pad , \wb1m_data_o[18]_pad , \wb1m_data_o[19]_pad , \wb1m_data_o[1]_pad , \wb1m_data_o[20]_pad , \wb1m_data_o[21]_pad , \wb1m_data_o[22]_pad , \wb1m_data_o[23]_pad , \wb1m_data_o[24]_pad , \wb1m_data_o[25]_pad , \wb1m_data_o[26]_pad , \wb1m_data_o[27]_pad , \wb1m_data_o[28]_pad , \wb1m_data_o[29]_pad , \wb1m_data_o[2]_pad , \wb1m_data_o[30]_pad , \wb1m_data_o[31]_pad , \wb1m_data_o[3]_pad , \wb1m_data_o[4]_pad , \wb1m_data_o[5]_pad , \wb1m_data_o[6]_pad , \wb1m_data_o[7]_pad , \wb1m_data_o[8]_pad , \wb1m_data_o[9]_pad , \wb1s_data_o[0]_pad , \wb1s_data_o[10]_pad , \wb1s_data_o[11]_pad , \wb1s_data_o[12]_pad , \wb1s_data_o[13]_pad , \wb1s_data_o[14]_pad , \wb1s_data_o[15]_pad , \wb1s_data_o[16]_pad , \wb1s_data_o[17]_pad , \wb1s_data_o[18]_pad , \wb1s_data_o[19]_pad , \wb1s_data_o[1]_pad , \wb1s_data_o[20]_pad , \wb1s_data_o[21]_pad , \wb1s_data_o[22]_pad , \wb1s_data_o[23]_pad , \wb1s_data_o[24]_pad , \wb1s_data_o[25]_pad , \wb1s_data_o[26]_pad , \wb1s_data_o[27]_pad , \wb1s_data_o[28]_pad , \wb1s_data_o[29]_pad , \wb1s_data_o[2]_pad , \wb1s_data_o[30]_pad , \wb1s_data_o[31]_pad , \wb1s_data_o[3]_pad , \wb1s_data_o[4]_pad , \wb1s_data_o[5]_pad , \wb1s_data_o[6]_pad , \wb1s_data_o[7]_pad , \wb1s_data_o[8]_pad , \wb1s_data_o[9]_pad );
	input dma_ack_o_pad ;
	input dma_nd_i_pad ;
	input dma_req_i_pad ;
	input \u0_csr_r_reg[0]/NET0131  ;
	input \u0_int_maska_r_reg[0]/NET0131  ;
	input \u0_int_maska_r_reg[10]/NET0131  ;
	input \u0_int_maska_r_reg[11]/NET0131  ;
	input \u0_int_maska_r_reg[12]/NET0131  ;
	input \u0_int_maska_r_reg[13]/NET0131  ;
	input \u0_int_maska_r_reg[14]/NET0131  ;
	input \u0_int_maska_r_reg[15]/NET0131  ;
	input \u0_int_maska_r_reg[16]/NET0131  ;
	input \u0_int_maska_r_reg[17]/NET0131  ;
	input \u0_int_maska_r_reg[18]/NET0131  ;
	input \u0_int_maska_r_reg[19]/NET0131  ;
	input \u0_int_maska_r_reg[1]/NET0131  ;
	input \u0_int_maska_r_reg[20]/NET0131  ;
	input \u0_int_maska_r_reg[21]/NET0131  ;
	input \u0_int_maska_r_reg[22]/NET0131  ;
	input \u0_int_maska_r_reg[23]/NET0131  ;
	input \u0_int_maska_r_reg[24]/NET0131  ;
	input \u0_int_maska_r_reg[25]/NET0131  ;
	input \u0_int_maska_r_reg[26]/NET0131  ;
	input \u0_int_maska_r_reg[27]/NET0131  ;
	input \u0_int_maska_r_reg[28]/NET0131  ;
	input \u0_int_maska_r_reg[29]/NET0131  ;
	input \u0_int_maska_r_reg[2]/NET0131  ;
	input \u0_int_maska_r_reg[30]/NET0131  ;
	input \u0_int_maska_r_reg[3]/NET0131  ;
	input \u0_int_maska_r_reg[4]/NET0131  ;
	input \u0_int_maska_r_reg[5]/NET0131  ;
	input \u0_int_maska_r_reg[6]/NET0131  ;
	input \u0_int_maska_r_reg[7]/NET0131  ;
	input \u0_int_maska_r_reg[8]/NET0131  ;
	input \u0_int_maska_r_reg[9]/NET0131  ;
	input \u0_int_maskb_r_reg[0]/NET0131  ;
	input \u0_int_maskb_r_reg[10]/NET0131  ;
	input \u0_int_maskb_r_reg[11]/NET0131  ;
	input \u0_int_maskb_r_reg[12]/NET0131  ;
	input \u0_int_maskb_r_reg[13]/NET0131  ;
	input \u0_int_maskb_r_reg[14]/NET0131  ;
	input \u0_int_maskb_r_reg[15]/NET0131  ;
	input \u0_int_maskb_r_reg[16]/NET0131  ;
	input \u0_int_maskb_r_reg[17]/NET0131  ;
	input \u0_int_maskb_r_reg[18]/NET0131  ;
	input \u0_int_maskb_r_reg[19]/NET0131  ;
	input \u0_int_maskb_r_reg[1]/NET0131  ;
	input \u0_int_maskb_r_reg[20]/NET0131  ;
	input \u0_int_maskb_r_reg[21]/NET0131  ;
	input \u0_int_maskb_r_reg[22]/NET0131  ;
	input \u0_int_maskb_r_reg[23]/NET0131  ;
	input \u0_int_maskb_r_reg[24]/NET0131  ;
	input \u0_int_maskb_r_reg[25]/NET0131  ;
	input \u0_int_maskb_r_reg[26]/NET0131  ;
	input \u0_int_maskb_r_reg[27]/NET0131  ;
	input \u0_int_maskb_r_reg[28]/NET0131  ;
	input \u0_int_maskb_r_reg[29]/NET0131  ;
	input \u0_int_maskb_r_reg[2]/NET0131  ;
	input \u0_int_maskb_r_reg[30]/NET0131  ;
	input \u0_int_maskb_r_reg[3]/NET0131  ;
	input \u0_int_maskb_r_reg[4]/NET0131  ;
	input \u0_int_maskb_r_reg[5]/NET0131  ;
	input \u0_int_maskb_r_reg[6]/NET0131  ;
	input \u0_int_maskb_r_reg[7]/NET0131  ;
	input \u0_int_maskb_r_reg[8]/NET0131  ;
	input \u0_int_maskb_r_reg[9]/NET0131  ;
	input \u0_u0_ch_adr0_r_reg[0]/P0001  ;
	input \u0_u0_ch_adr0_r_reg[10]/P0001  ;
	input \u0_u0_ch_adr0_r_reg[11]/P0001  ;
	input \u0_u0_ch_adr0_r_reg[12]/P0001  ;
	input \u0_u0_ch_adr0_r_reg[13]/P0001  ;
	input \u0_u0_ch_adr0_r_reg[14]/P0001  ;
	input \u0_u0_ch_adr0_r_reg[15]/P0001  ;
	input \u0_u0_ch_adr0_r_reg[16]/P0001  ;
	input \u0_u0_ch_adr0_r_reg[17]/P0001  ;
	input \u0_u0_ch_adr0_r_reg[18]/P0001  ;
	input \u0_u0_ch_adr0_r_reg[19]/P0001  ;
	input \u0_u0_ch_adr0_r_reg[1]/P0001  ;
	input \u0_u0_ch_adr0_r_reg[20]/P0001  ;
	input \u0_u0_ch_adr0_r_reg[21]/P0001  ;
	input \u0_u0_ch_adr0_r_reg[22]/P0001  ;
	input \u0_u0_ch_adr0_r_reg[23]/P0001  ;
	input \u0_u0_ch_adr0_r_reg[24]/P0001  ;
	input \u0_u0_ch_adr0_r_reg[25]/P0001  ;
	input \u0_u0_ch_adr0_r_reg[26]/P0001  ;
	input \u0_u0_ch_adr0_r_reg[27]/P0001  ;
	input \u0_u0_ch_adr0_r_reg[28]/P0001  ;
	input \u0_u0_ch_adr0_r_reg[29]/P0001  ;
	input \u0_u0_ch_adr0_r_reg[2]/P0001  ;
	input \u0_u0_ch_adr0_r_reg[3]/P0001  ;
	input \u0_u0_ch_adr0_r_reg[4]/P0001  ;
	input \u0_u0_ch_adr0_r_reg[5]/P0001  ;
	input \u0_u0_ch_adr0_r_reg[6]/P0001  ;
	input \u0_u0_ch_adr0_r_reg[7]/P0001  ;
	input \u0_u0_ch_adr0_r_reg[8]/P0001  ;
	input \u0_u0_ch_adr0_r_reg[9]/P0001  ;
	input \u0_u0_ch_adr1_r_reg[0]/P0001  ;
	input \u0_u0_ch_adr1_r_reg[10]/P0001  ;
	input \u0_u0_ch_adr1_r_reg[11]/P0001  ;
	input \u0_u0_ch_adr1_r_reg[12]/P0001  ;
	input \u0_u0_ch_adr1_r_reg[13]/P0001  ;
	input \u0_u0_ch_adr1_r_reg[14]/P0001  ;
	input \u0_u0_ch_adr1_r_reg[15]/P0001  ;
	input \u0_u0_ch_adr1_r_reg[16]/P0001  ;
	input \u0_u0_ch_adr1_r_reg[17]/P0001  ;
	input \u0_u0_ch_adr1_r_reg[18]/P0001  ;
	input \u0_u0_ch_adr1_r_reg[19]/P0001  ;
	input \u0_u0_ch_adr1_r_reg[1]/P0001  ;
	input \u0_u0_ch_adr1_r_reg[20]/P0001  ;
	input \u0_u0_ch_adr1_r_reg[21]/P0001  ;
	input \u0_u0_ch_adr1_r_reg[22]/P0001  ;
	input \u0_u0_ch_adr1_r_reg[23]/P0001  ;
	input \u0_u0_ch_adr1_r_reg[24]/P0001  ;
	input \u0_u0_ch_adr1_r_reg[25]/P0001  ;
	input \u0_u0_ch_adr1_r_reg[26]/P0001  ;
	input \u0_u0_ch_adr1_r_reg[27]/P0001  ;
	input \u0_u0_ch_adr1_r_reg[28]/P0001  ;
	input \u0_u0_ch_adr1_r_reg[29]/P0001  ;
	input \u0_u0_ch_adr1_r_reg[2]/P0001  ;
	input \u0_u0_ch_adr1_r_reg[3]/P0001  ;
	input \u0_u0_ch_adr1_r_reg[4]/P0001  ;
	input \u0_u0_ch_adr1_r_reg[5]/P0001  ;
	input \u0_u0_ch_adr1_r_reg[6]/P0001  ;
	input \u0_u0_ch_adr1_r_reg[7]/P0001  ;
	input \u0_u0_ch_adr1_r_reg[8]/P0001  ;
	input \u0_u0_ch_adr1_r_reg[9]/P0001  ;
	input \u0_u0_ch_busy_reg/P0001  ;
	input \u0_u0_ch_chk_sz_r_reg[0]/P0001  ;
	input \u0_u0_ch_chk_sz_r_reg[10]/P0001  ;
	input \u0_u0_ch_chk_sz_r_reg[1]/P0001  ;
	input \u0_u0_ch_chk_sz_r_reg[2]/P0001  ;
	input \u0_u0_ch_chk_sz_r_reg[3]/P0001  ;
	input \u0_u0_ch_chk_sz_r_reg[4]/P0001  ;
	input \u0_u0_ch_chk_sz_r_reg[5]/P0001  ;
	input \u0_u0_ch_chk_sz_r_reg[6]/P0001  ;
	input \u0_u0_ch_chk_sz_r_reg[7]/P0001  ;
	input \u0_u0_ch_chk_sz_r_reg[8]/P0001  ;
	input \u0_u0_ch_chk_sz_r_reg[9]/P0001  ;
	input \u0_u0_ch_csr_r2_reg[0]/NET0131  ;
	input \u0_u0_ch_csr_r2_reg[1]/NET0131  ;
	input \u0_u0_ch_csr_r2_reg[2]/NET0131  ;
	input \u0_u0_ch_csr_r3_reg[0]/NET0131  ;
	input \u0_u0_ch_csr_r3_reg[1]/NET0131  ;
	input \u0_u0_ch_csr_r3_reg[2]/NET0131  ;
	input \u0_u0_ch_csr_r_reg[0]/NET0131  ;
	input \u0_u0_ch_csr_r_reg[1]/NET0131  ;
	input \u0_u0_ch_csr_r_reg[2]/NET0131  ;
	input \u0_u0_ch_csr_r_reg[3]/NET0131  ;
	input \u0_u0_ch_csr_r_reg[4]/NET0131  ;
	input \u0_u0_ch_csr_r_reg[5]/NET0131  ;
	input \u0_u0_ch_csr_r_reg[6]/NET0131  ;
	input \u0_u0_ch_csr_r_reg[7]/NET0131  ;
	input \u0_u0_ch_csr_r_reg[8]/NET0131  ;
	input \u0_u0_ch_done_reg/P0002  ;
	input \u0_u0_ch_err_reg/NET0131  ;
	input \u0_u0_ch_stop_reg/P0001  ;
	input \u0_u0_ch_sz_inf_reg/NET0131  ;
	input \u0_u0_ch_tot_sz_r_reg[0]/P0001  ;
	input \u0_u0_ch_tot_sz_r_reg[10]/P0001  ;
	input \u0_u0_ch_tot_sz_r_reg[11]/P0001  ;
	input \u0_u0_ch_tot_sz_r_reg[1]/P0001  ;
	input \u0_u0_ch_tot_sz_r_reg[2]/P0001  ;
	input \u0_u0_ch_tot_sz_r_reg[3]/P0001  ;
	input \u0_u0_ch_tot_sz_r_reg[4]/P0001  ;
	input \u0_u0_ch_tot_sz_r_reg[5]/P0001  ;
	input \u0_u0_ch_tot_sz_r_reg[6]/P0001  ;
	input \u0_u0_ch_tot_sz_r_reg[7]/P0001  ;
	input \u0_u0_ch_tot_sz_r_reg[8]/P0001  ;
	input \u0_u0_ch_tot_sz_r_reg[9]/P0001  ;
	input \u0_u0_int_src_r_reg[1]/NET0131  ;
	input \u0_u0_int_src_r_reg[2]/NET0131  ;
	input \u0_u0_rest_en_reg/NET0131  ;
	input \u0_wb_rf_dout_reg[0]/P0001  ;
	input \u0_wb_rf_dout_reg[10]/P0001  ;
	input \u0_wb_rf_dout_reg[11]/P0001  ;
	input \u0_wb_rf_dout_reg[12]/P0001  ;
	input \u0_wb_rf_dout_reg[13]/P0001  ;
	input \u0_wb_rf_dout_reg[14]/P0001  ;
	input \u0_wb_rf_dout_reg[15]/P0001  ;
	input \u0_wb_rf_dout_reg[16]/P0001  ;
	input \u0_wb_rf_dout_reg[17]/P0001  ;
	input \u0_wb_rf_dout_reg[18]/P0001  ;
	input \u0_wb_rf_dout_reg[19]/P0001  ;
	input \u0_wb_rf_dout_reg[1]/P0001  ;
	input \u0_wb_rf_dout_reg[20]/P0001  ;
	input \u0_wb_rf_dout_reg[21]/P0001  ;
	input \u0_wb_rf_dout_reg[22]/P0001  ;
	input \u0_wb_rf_dout_reg[23]/P0001  ;
	input \u0_wb_rf_dout_reg[24]/P0001  ;
	input \u0_wb_rf_dout_reg[25]/P0001  ;
	input \u0_wb_rf_dout_reg[26]/P0001  ;
	input \u0_wb_rf_dout_reg[27]/P0001  ;
	input \u0_wb_rf_dout_reg[28]/P0001  ;
	input \u0_wb_rf_dout_reg[29]/P0001  ;
	input \u0_wb_rf_dout_reg[2]/P0001  ;
	input \u0_wb_rf_dout_reg[30]/P0001  ;
	input \u0_wb_rf_dout_reg[31]/P0001  ;
	input \u0_wb_rf_dout_reg[3]/P0001  ;
	input \u0_wb_rf_dout_reg[4]/P0001  ;
	input \u0_wb_rf_dout_reg[5]/P0001  ;
	input \u0_wb_rf_dout_reg[6]/P0001  ;
	input \u0_wb_rf_dout_reg[7]/P0001  ;
	input \u0_wb_rf_dout_reg[8]/P0001  ;
	input \u0_wb_rf_dout_reg[9]/P0001  ;
	input \u1_de_start_r_reg/P0001  ;
	input \u1_ndnr_reg[0]/P0001  ;
	input \u1_ndr_r_reg[0]/NET0131  ;
	input \u1_next_start_reg/P0001  ;
	input \u1_req_r_reg[0]/P0001  ;
	input \u2_adr0_cnt_reg[0]/P0001  ;
	input \u2_adr0_cnt_reg[10]/P0001  ;
	input \u2_adr0_cnt_reg[11]/P0001  ;
	input \u2_adr0_cnt_reg[12]/P0001  ;
	input \u2_adr0_cnt_reg[13]/P0001  ;
	input \u2_adr0_cnt_reg[14]/P0001  ;
	input \u2_adr0_cnt_reg[15]/P0001  ;
	input \u2_adr0_cnt_reg[16]/NET0131  ;
	input \u2_adr0_cnt_reg[17]/P0001  ;
	input \u2_adr0_cnt_reg[18]/P0001  ;
	input \u2_adr0_cnt_reg[19]/P0001  ;
	input \u2_adr0_cnt_reg[1]/P0001  ;
	input \u2_adr0_cnt_reg[20]/P0001  ;
	input \u2_adr0_cnt_reg[21]/P0001  ;
	input \u2_adr0_cnt_reg[22]/P0001  ;
	input \u2_adr0_cnt_reg[23]/P0001  ;
	input \u2_adr0_cnt_reg[24]/P0001  ;
	input \u2_adr0_cnt_reg[25]/P0001  ;
	input \u2_adr0_cnt_reg[26]/P0001  ;
	input \u2_adr0_cnt_reg[27]/P0001  ;
	input \u2_adr0_cnt_reg[28]/P0001  ;
	input \u2_adr0_cnt_reg[29]/P0001  ;
	input \u2_adr0_cnt_reg[2]/P0001  ;
	input \u2_adr0_cnt_reg[3]/P0001  ;
	input \u2_adr0_cnt_reg[4]/P0001  ;
	input \u2_adr0_cnt_reg[5]/P0001  ;
	input \u2_adr0_cnt_reg[6]/P0001  ;
	input \u2_adr0_cnt_reg[7]/P0001  ;
	input \u2_adr0_cnt_reg[8]/P0001  ;
	input \u2_adr0_cnt_reg[9]/P0001  ;
	input \u2_adr1_cnt_reg[0]/P0001  ;
	input \u2_adr1_cnt_reg[10]/P0001  ;
	input \u2_adr1_cnt_reg[11]/P0001  ;
	input \u2_adr1_cnt_reg[12]/P0001  ;
	input \u2_adr1_cnt_reg[13]/P0001  ;
	input \u2_adr1_cnt_reg[14]/P0001  ;
	input \u2_adr1_cnt_reg[15]/P0001  ;
	input \u2_adr1_cnt_reg[16]/NET0131  ;
	input \u2_adr1_cnt_reg[17]/P0001  ;
	input \u2_adr1_cnt_reg[18]/P0001  ;
	input \u2_adr1_cnt_reg[19]/P0001  ;
	input \u2_adr1_cnt_reg[1]/P0001  ;
	input \u2_adr1_cnt_reg[20]/P0001  ;
	input \u2_adr1_cnt_reg[21]/P0001  ;
	input \u2_adr1_cnt_reg[22]/P0001  ;
	input \u2_adr1_cnt_reg[23]/P0001  ;
	input \u2_adr1_cnt_reg[24]/P0001  ;
	input \u2_adr1_cnt_reg[25]/P0001  ;
	input \u2_adr1_cnt_reg[26]/P0001  ;
	input \u2_adr1_cnt_reg[27]/P0001  ;
	input \u2_adr1_cnt_reg[28]/P0001  ;
	input \u2_adr1_cnt_reg[29]/P0001  ;
	input \u2_adr1_cnt_reg[2]/P0001  ;
	input \u2_adr1_cnt_reg[3]/P0001  ;
	input \u2_adr1_cnt_reg[4]/P0001  ;
	input \u2_adr1_cnt_reg[5]/P0001  ;
	input \u2_adr1_cnt_reg[6]/P0001  ;
	input \u2_adr1_cnt_reg[7]/P0001  ;
	input \u2_adr1_cnt_reg[8]/P0001  ;
	input \u2_adr1_cnt_reg[9]/P0001  ;
	input \u2_chunk_0_reg/P0001  ;
	input \u2_chunk_cnt_is_0_r_reg/P0001  ;
	input \u2_chunk_cnt_reg[0]/NET0131  ;
	input \u2_chunk_cnt_reg[1]/NET0131  ;
	input \u2_chunk_cnt_reg[2]/NET0131  ;
	input \u2_chunk_cnt_reg[3]/NET0131  ;
	input \u2_chunk_cnt_reg[4]/NET0131  ;
	input \u2_chunk_cnt_reg[5]/NET0131  ;
	input \u2_chunk_cnt_reg[6]/NET0131  ;
	input \u2_chunk_cnt_reg[7]/NET0131  ;
	input \u2_chunk_cnt_reg[8]/NET0131  ;
	input \u2_chunk_dec_reg/P0001  ;
	input \u2_dma_abort_r_reg/NET0131  ;
	input \u2_mast0_adr_reg[10]/P0001  ;
	input \u2_mast0_adr_reg[11]/P0001  ;
	input \u2_mast0_adr_reg[12]/P0001  ;
	input \u2_mast0_adr_reg[13]/P0001  ;
	input \u2_mast0_adr_reg[14]/P0001  ;
	input \u2_mast0_adr_reg[15]/P0001  ;
	input \u2_mast0_adr_reg[16]/P0001  ;
	input \u2_mast0_adr_reg[17]/P0001  ;
	input \u2_mast0_adr_reg[18]/P0001  ;
	input \u2_mast0_adr_reg[19]/P0001  ;
	input \u2_mast0_adr_reg[20]/P0001  ;
	input \u2_mast0_adr_reg[21]/P0001  ;
	input \u2_mast0_adr_reg[22]/P0001  ;
	input \u2_mast0_adr_reg[23]/P0001  ;
	input \u2_mast0_adr_reg[24]/P0001  ;
	input \u2_mast0_adr_reg[25]/P0001  ;
	input \u2_mast0_adr_reg[26]/P0001  ;
	input \u2_mast0_adr_reg[27]/P0001  ;
	input \u2_mast0_adr_reg[28]/P0001  ;
	input \u2_mast0_adr_reg[29]/P0001  ;
	input \u2_mast0_adr_reg[2]/P0001  ;
	input \u2_mast0_adr_reg[30]/P0001  ;
	input \u2_mast0_adr_reg[31]/P0001  ;
	input \u2_mast0_adr_reg[3]/NET0131  ;
	input \u2_mast0_adr_reg[4]/P0001  ;
	input \u2_mast0_adr_reg[5]/P0001  ;
	input \u2_mast0_adr_reg[6]/P0001  ;
	input \u2_mast0_adr_reg[7]/P0001  ;
	input \u2_mast0_adr_reg[8]/P0001  ;
	input \u2_mast0_adr_reg[9]/P0001  ;
	input \u2_mast0_drdy_r_reg/P0001  ;
	input \u2_mast1_adr_reg[10]/P0001  ;
	input \u2_mast1_adr_reg[11]/P0001  ;
	input \u2_mast1_adr_reg[12]/P0001  ;
	input \u2_mast1_adr_reg[13]/P0001  ;
	input \u2_mast1_adr_reg[14]/P0001  ;
	input \u2_mast1_adr_reg[15]/P0001  ;
	input \u2_mast1_adr_reg[16]/P0001  ;
	input \u2_mast1_adr_reg[17]/P0001  ;
	input \u2_mast1_adr_reg[18]/P0001  ;
	input \u2_mast1_adr_reg[19]/P0001  ;
	input \u2_mast1_adr_reg[20]/P0001  ;
	input \u2_mast1_adr_reg[21]/P0001  ;
	input \u2_mast1_adr_reg[22]/P0001  ;
	input \u2_mast1_adr_reg[23]/P0001  ;
	input \u2_mast1_adr_reg[24]/P0001  ;
	input \u2_mast1_adr_reg[25]/P0001  ;
	input \u2_mast1_adr_reg[26]/P0001  ;
	input \u2_mast1_adr_reg[27]/P0001  ;
	input \u2_mast1_adr_reg[28]/P0001  ;
	input \u2_mast1_adr_reg[29]/P0001  ;
	input \u2_mast1_adr_reg[2]/P0001  ;
	input \u2_mast1_adr_reg[30]/P0001  ;
	input \u2_mast1_adr_reg[31]/P0001  ;
	input \u2_mast1_adr_reg[3]/P0001  ;
	input \u2_mast1_adr_reg[4]/P0001  ;
	input \u2_mast1_adr_reg[5]/P0001  ;
	input \u2_mast1_adr_reg[6]/P0001  ;
	input \u2_mast1_adr_reg[7]/P0001  ;
	input \u2_mast1_adr_reg[8]/P0001  ;
	input \u2_mast1_adr_reg[9]/P0001  ;
	input \u2_next_ch_reg/P0001  ;
	input \u2_read_r_reg/P0001  ;
	input \u2_state_reg[0]/NET0131  ;
	input \u2_state_reg[10]/NET0131  ;
	input \u2_state_reg[1]/NET0131  ;
	input \u2_state_reg[2]/NET0131  ;
	input \u2_state_reg[3]/NET0131  ;
	input \u2_state_reg[4]/NET0131  ;
	input \u2_state_reg[5]/NET0131  ;
	input \u2_state_reg[6]/NET0131  ;
	input \u2_state_reg[7]/NET0131  ;
	input \u2_state_reg[8]/NET0131  ;
	input \u2_state_reg[9]/NET0131  ;
	input \u2_tsz_cnt_is_0_r_reg/P0001  ;
	input \u2_tsz_cnt_reg[0]/NET0131  ;
	input \u2_tsz_cnt_reg[10]/NET0131  ;
	input \u2_tsz_cnt_reg[11]/NET0131  ;
	input \u2_tsz_cnt_reg[1]/NET0131  ;
	input \u2_tsz_cnt_reg[2]/NET0131  ;
	input \u2_tsz_cnt_reg[3]/NET0131  ;
	input \u2_tsz_cnt_reg[4]/NET0131  ;
	input \u2_tsz_cnt_reg[5]/NET0131  ;
	input \u2_tsz_cnt_reg[6]/NET0131  ;
	input \u2_tsz_cnt_reg[7]/NET0131  ;
	input \u2_tsz_cnt_reg[8]/NET0131  ;
	input \u2_tsz_cnt_reg[9]/NET0131  ;
	input \u2_u0_out_r_reg[0]/P0001  ;
	input \u2_u0_out_r_reg[10]/P0001  ;
	input \u2_u0_out_r_reg[11]/P0001  ;
	input \u2_u0_out_r_reg[12]/P0001  ;
	input \u2_u0_out_r_reg[13]/P0001  ;
	input \u2_u0_out_r_reg[14]/P0001  ;
	input \u2_u0_out_r_reg[15]/P0001  ;
	input \u2_u0_out_r_reg[16]/P0001  ;
	input \u2_u0_out_r_reg[1]/P0001  ;
	input \u2_u0_out_r_reg[2]/P0001  ;
	input \u2_u0_out_r_reg[3]/P0001  ;
	input \u2_u0_out_r_reg[4]/P0001  ;
	input \u2_u0_out_r_reg[5]/P0001  ;
	input \u2_u0_out_r_reg[6]/P0001  ;
	input \u2_u0_out_r_reg[7]/P0001  ;
	input \u2_u0_out_r_reg[8]/P0001  ;
	input \u2_u0_out_r_reg[9]/P0001  ;
	input \u2_u1_out_r_reg[0]/P0001  ;
	input \u2_u1_out_r_reg[10]/P0001  ;
	input \u2_u1_out_r_reg[11]/P0001  ;
	input \u2_u1_out_r_reg[12]/P0001  ;
	input \u2_u1_out_r_reg[13]/P0001  ;
	input \u2_u1_out_r_reg[14]/P0001  ;
	input \u2_u1_out_r_reg[15]/P0001  ;
	input \u2_u1_out_r_reg[16]/P0001  ;
	input \u2_u1_out_r_reg[1]/P0001  ;
	input \u2_u1_out_r_reg[2]/P0001  ;
	input \u2_u1_out_r_reg[3]/P0001  ;
	input \u2_u1_out_r_reg[4]/P0001  ;
	input \u2_u1_out_r_reg[5]/P0001  ;
	input \u2_u1_out_r_reg[6]/P0001  ;
	input \u2_u1_out_r_reg[7]/P0001  ;
	input \u2_u1_out_r_reg[8]/P0001  ;
	input \u2_u1_out_r_reg[9]/P0001  ;
	input \u2_write_hold_r_reg/P0001  ;
	input \u2_write_r_reg/P0001  ;
	input \u3_u0_mast_cyc_reg/P0001  ;
	input \u3_u0_mast_dout_reg[0]/P0001  ;
	input \u3_u0_mast_dout_reg[10]/P0001  ;
	input \u3_u0_mast_dout_reg[11]/P0001  ;
	input \u3_u0_mast_dout_reg[12]/P0001  ;
	input \u3_u0_mast_dout_reg[13]/P0001  ;
	input \u3_u0_mast_dout_reg[14]/P0001  ;
	input \u3_u0_mast_dout_reg[15]/P0001  ;
	input \u3_u0_mast_dout_reg[16]/P0001  ;
	input \u3_u0_mast_dout_reg[17]/P0001  ;
	input \u3_u0_mast_dout_reg[18]/P0001  ;
	input \u3_u0_mast_dout_reg[19]/P0001  ;
	input \u3_u0_mast_dout_reg[1]/P0001  ;
	input \u3_u0_mast_dout_reg[20]/P0001  ;
	input \u3_u0_mast_dout_reg[21]/P0001  ;
	input \u3_u0_mast_dout_reg[22]/P0001  ;
	input \u3_u0_mast_dout_reg[23]/P0001  ;
	input \u3_u0_mast_dout_reg[24]/P0001  ;
	input \u3_u0_mast_dout_reg[25]/P0001  ;
	input \u3_u0_mast_dout_reg[26]/P0001  ;
	input \u3_u0_mast_dout_reg[27]/P0001  ;
	input \u3_u0_mast_dout_reg[28]/P0001  ;
	input \u3_u0_mast_dout_reg[29]/P0001  ;
	input \u3_u0_mast_dout_reg[2]/P0001  ;
	input \u3_u0_mast_dout_reg[30]/P0001  ;
	input \u3_u0_mast_dout_reg[31]/P0001  ;
	input \u3_u0_mast_dout_reg[3]/P0001  ;
	input \u3_u0_mast_dout_reg[4]/P0001  ;
	input \u3_u0_mast_dout_reg[5]/P0001  ;
	input \u3_u0_mast_dout_reg[6]/P0001  ;
	input \u3_u0_mast_dout_reg[7]/P0001  ;
	input \u3_u0_mast_dout_reg[8]/P0001  ;
	input \u3_u0_mast_dout_reg[9]/P0001  ;
	input \u3_u0_mast_stb_reg/P0001  ;
	input \u3_u0_mast_we_r_reg/P0002  ;
	input \u3_u1_rf_ack_reg/P0001  ;
	input \u3_u1_slv_adr_reg[2]/NET0131  ;
	input \u3_u1_slv_adr_reg[3]/P0001  ;
	input \u3_u1_slv_adr_reg[4]/NET0131  ;
	input \u3_u1_slv_adr_reg[5]/P0001  ;
	input \u3_u1_slv_adr_reg[6]/NET0131  ;
	input \u3_u1_slv_adr_reg[7]/NET0131  ;
	input \u3_u1_slv_adr_reg[8]/NET0131  ;
	input \u3_u1_slv_adr_reg[9]/NET0131  ;
	input \u3_u1_slv_dout_reg[0]/P0001  ;
	input \u3_u1_slv_dout_reg[10]/P0001  ;
	input \u3_u1_slv_dout_reg[11]/P0001  ;
	input \u3_u1_slv_dout_reg[12]/P0001  ;
	input \u3_u1_slv_dout_reg[13]/P0001  ;
	input \u3_u1_slv_dout_reg[14]/P0001  ;
	input \u3_u1_slv_dout_reg[15]/P0001  ;
	input \u3_u1_slv_dout_reg[16]/P0001  ;
	input \u3_u1_slv_dout_reg[17]/P0001  ;
	input \u3_u1_slv_dout_reg[18]/P0001  ;
	input \u3_u1_slv_dout_reg[19]/P0001  ;
	input \u3_u1_slv_dout_reg[1]/P0001  ;
	input \u3_u1_slv_dout_reg[20]/P0001  ;
	input \u3_u1_slv_dout_reg[21]/P0001  ;
	input \u3_u1_slv_dout_reg[22]/P0001  ;
	input \u3_u1_slv_dout_reg[23]/P0001  ;
	input \u3_u1_slv_dout_reg[24]/P0001  ;
	input \u3_u1_slv_dout_reg[25]/P0001  ;
	input \u3_u1_slv_dout_reg[26]/P0001  ;
	input \u3_u1_slv_dout_reg[27]/P0001  ;
	input \u3_u1_slv_dout_reg[28]/P0001  ;
	input \u3_u1_slv_dout_reg[29]/P0001  ;
	input \u3_u1_slv_dout_reg[2]/P0001  ;
	input \u3_u1_slv_dout_reg[30]/P0001  ;
	input \u3_u1_slv_dout_reg[31]/P0001  ;
	input \u3_u1_slv_dout_reg[3]/P0001  ;
	input \u3_u1_slv_dout_reg[4]/P0001  ;
	input \u3_u1_slv_dout_reg[5]/P0001  ;
	input \u3_u1_slv_dout_reg[6]/P0001  ;
	input \u3_u1_slv_dout_reg[7]/P0001  ;
	input \u3_u1_slv_dout_reg[8]/P0001  ;
	input \u3_u1_slv_dout_reg[9]/P0001  ;
	input \u3_u1_slv_re_reg/P0001  ;
	input \u3_u1_slv_we_reg/P0001  ;
	input \u4_u0_mast_cyc_reg/P0001  ;
	input \u4_u0_mast_dout_reg[0]/P0001  ;
	input \u4_u0_mast_dout_reg[10]/P0001  ;
	input \u4_u0_mast_dout_reg[11]/P0001  ;
	input \u4_u0_mast_dout_reg[12]/P0001  ;
	input \u4_u0_mast_dout_reg[13]/P0001  ;
	input \u4_u0_mast_dout_reg[14]/P0001  ;
	input \u4_u0_mast_dout_reg[15]/P0001  ;
	input \u4_u0_mast_dout_reg[16]/P0001  ;
	input \u4_u0_mast_dout_reg[17]/P0001  ;
	input \u4_u0_mast_dout_reg[18]/P0001  ;
	input \u4_u0_mast_dout_reg[19]/P0001  ;
	input \u4_u0_mast_dout_reg[1]/P0001  ;
	input \u4_u0_mast_dout_reg[20]/P0001  ;
	input \u4_u0_mast_dout_reg[21]/P0001  ;
	input \u4_u0_mast_dout_reg[22]/P0001  ;
	input \u4_u0_mast_dout_reg[23]/P0001  ;
	input \u4_u0_mast_dout_reg[24]/P0001  ;
	input \u4_u0_mast_dout_reg[25]/P0001  ;
	input \u4_u0_mast_dout_reg[26]/P0001  ;
	input \u4_u0_mast_dout_reg[27]/P0001  ;
	input \u4_u0_mast_dout_reg[28]/P0001  ;
	input \u4_u0_mast_dout_reg[29]/P0001  ;
	input \u4_u0_mast_dout_reg[2]/P0001  ;
	input \u4_u0_mast_dout_reg[30]/P0001  ;
	input \u4_u0_mast_dout_reg[31]/P0001  ;
	input \u4_u0_mast_dout_reg[3]/P0001  ;
	input \u4_u0_mast_dout_reg[4]/P0001  ;
	input \u4_u0_mast_dout_reg[5]/P0001  ;
	input \u4_u0_mast_dout_reg[6]/P0001  ;
	input \u4_u0_mast_dout_reg[7]/P0001  ;
	input \u4_u0_mast_dout_reg[8]/P0001  ;
	input \u4_u0_mast_dout_reg[9]/P0001  ;
	input \u4_u0_mast_stb_reg/P0001  ;
	input \u4_u0_mast_we_r_reg/P0001  ;
	input \u4_u1_rf_ack_reg/P0001  ;
	input \u4_u1_slv_re_reg/P0001  ;
	input \u4_u1_slv_we_reg/P0001  ;
	input \wb0_ack_i_pad  ;
	input \wb0_addr_i[0]_pad  ;
	input \wb0_addr_i[10]_pad  ;
	input \wb0_addr_i[11]_pad  ;
	input \wb0_addr_i[12]_pad  ;
	input \wb0_addr_i[13]_pad  ;
	input \wb0_addr_i[14]_pad  ;
	input \wb0_addr_i[15]_pad  ;
	input \wb0_addr_i[16]_pad  ;
	input \wb0_addr_i[17]_pad  ;
	input \wb0_addr_i[18]_pad  ;
	input \wb0_addr_i[19]_pad  ;
	input \wb0_addr_i[1]_pad  ;
	input \wb0_addr_i[20]_pad  ;
	input \wb0_addr_i[21]_pad  ;
	input \wb0_addr_i[22]_pad  ;
	input \wb0_addr_i[23]_pad  ;
	input \wb0_addr_i[24]_pad  ;
	input \wb0_addr_i[25]_pad  ;
	input \wb0_addr_i[26]_pad  ;
	input \wb0_addr_i[27]_pad  ;
	input \wb0_addr_i[28]_pad  ;
	input \wb0_addr_i[29]_pad  ;
	input \wb0_addr_i[2]_pad  ;
	input \wb0_addr_i[30]_pad  ;
	input \wb0_addr_i[31]_pad  ;
	input \wb0_addr_i[3]_pad  ;
	input \wb0_addr_i[4]_pad  ;
	input \wb0_addr_i[5]_pad  ;
	input \wb0_addr_i[6]_pad  ;
	input \wb0_addr_i[7]_pad  ;
	input \wb0_addr_i[8]_pad  ;
	input \wb0_addr_i[9]_pad  ;
	input \wb0_cyc_i_pad  ;
	input \wb0_err_i_pad  ;
	input \wb0_rty_i_pad  ;
	input \wb0_sel_i[0]_pad  ;
	input \wb0_sel_i[1]_pad  ;
	input \wb0_sel_i[2]_pad  ;
	input \wb0_sel_i[3]_pad  ;
	input \wb0_stb_i_pad  ;
	input \wb0_we_i_pad  ;
	input \wb0m_data_i[0]_pad  ;
	input \wb0m_data_i[10]_pad  ;
	input \wb0m_data_i[11]_pad  ;
	input \wb0m_data_i[12]_pad  ;
	input \wb0m_data_i[13]_pad  ;
	input \wb0m_data_i[14]_pad  ;
	input \wb0m_data_i[15]_pad  ;
	input \wb0m_data_i[16]_pad  ;
	input \wb0m_data_i[17]_pad  ;
	input \wb0m_data_i[18]_pad  ;
	input \wb0m_data_i[19]_pad  ;
	input \wb0m_data_i[1]_pad  ;
	input \wb0m_data_i[20]_pad  ;
	input \wb0m_data_i[21]_pad  ;
	input \wb0m_data_i[22]_pad  ;
	input \wb0m_data_i[23]_pad  ;
	input \wb0m_data_i[24]_pad  ;
	input \wb0m_data_i[25]_pad  ;
	input \wb0m_data_i[26]_pad  ;
	input \wb0m_data_i[27]_pad  ;
	input \wb0m_data_i[28]_pad  ;
	input \wb0m_data_i[29]_pad  ;
	input \wb0m_data_i[2]_pad  ;
	input \wb0m_data_i[30]_pad  ;
	input \wb0m_data_i[31]_pad  ;
	input \wb0m_data_i[3]_pad  ;
	input \wb0m_data_i[4]_pad  ;
	input \wb0m_data_i[5]_pad  ;
	input \wb0m_data_i[6]_pad  ;
	input \wb0m_data_i[7]_pad  ;
	input \wb0m_data_i[8]_pad  ;
	input \wb0m_data_i[9]_pad  ;
	input \wb0s_data_i[0]_pad  ;
	input \wb0s_data_i[10]_pad  ;
	input \wb0s_data_i[11]_pad  ;
	input \wb0s_data_i[12]_pad  ;
	input \wb0s_data_i[13]_pad  ;
	input \wb0s_data_i[14]_pad  ;
	input \wb0s_data_i[15]_pad  ;
	input \wb0s_data_i[16]_pad  ;
	input \wb0s_data_i[17]_pad  ;
	input \wb0s_data_i[18]_pad  ;
	input \wb0s_data_i[19]_pad  ;
	input \wb0s_data_i[1]_pad  ;
	input \wb0s_data_i[20]_pad  ;
	input \wb0s_data_i[21]_pad  ;
	input \wb0s_data_i[22]_pad  ;
	input \wb0s_data_i[23]_pad  ;
	input \wb0s_data_i[24]_pad  ;
	input \wb0s_data_i[25]_pad  ;
	input \wb0s_data_i[26]_pad  ;
	input \wb0s_data_i[27]_pad  ;
	input \wb0s_data_i[28]_pad  ;
	input \wb0s_data_i[29]_pad  ;
	input \wb0s_data_i[2]_pad  ;
	input \wb0s_data_i[30]_pad  ;
	input \wb0s_data_i[31]_pad  ;
	input \wb0s_data_i[3]_pad  ;
	input \wb0s_data_i[4]_pad  ;
	input \wb0s_data_i[5]_pad  ;
	input \wb0s_data_i[6]_pad  ;
	input \wb0s_data_i[7]_pad  ;
	input \wb0s_data_i[8]_pad  ;
	input \wb0s_data_i[9]_pad  ;
	input \wb1_ack_i_pad  ;
	input \wb1_addr_i[0]_pad  ;
	input \wb1_addr_i[10]_pad  ;
	input \wb1_addr_i[11]_pad  ;
	input \wb1_addr_i[12]_pad  ;
	input \wb1_addr_i[13]_pad  ;
	input \wb1_addr_i[14]_pad  ;
	input \wb1_addr_i[15]_pad  ;
	input \wb1_addr_i[16]_pad  ;
	input \wb1_addr_i[17]_pad  ;
	input \wb1_addr_i[18]_pad  ;
	input \wb1_addr_i[19]_pad  ;
	input \wb1_addr_i[1]_pad  ;
	input \wb1_addr_i[20]_pad  ;
	input \wb1_addr_i[21]_pad  ;
	input \wb1_addr_i[22]_pad  ;
	input \wb1_addr_i[23]_pad  ;
	input \wb1_addr_i[24]_pad  ;
	input \wb1_addr_i[25]_pad  ;
	input \wb1_addr_i[26]_pad  ;
	input \wb1_addr_i[27]_pad  ;
	input \wb1_addr_i[28]_pad  ;
	input \wb1_addr_i[29]_pad  ;
	input \wb1_addr_i[2]_pad  ;
	input \wb1_addr_i[30]_pad  ;
	input \wb1_addr_i[31]_pad  ;
	input \wb1_addr_i[3]_pad  ;
	input \wb1_addr_i[4]_pad  ;
	input \wb1_addr_i[5]_pad  ;
	input \wb1_addr_i[6]_pad  ;
	input \wb1_addr_i[7]_pad  ;
	input \wb1_addr_i[8]_pad  ;
	input \wb1_addr_i[9]_pad  ;
	input \wb1_cyc_i_pad  ;
	input \wb1_err_i_pad  ;
	input \wb1_rty_i_pad  ;
	input \wb1_sel_i[0]_pad  ;
	input \wb1_sel_i[1]_pad  ;
	input \wb1_sel_i[2]_pad  ;
	input \wb1_sel_i[3]_pad  ;
	input \wb1_stb_i_pad  ;
	input \wb1_we_i_pad  ;
	input \wb1m_data_i[0]_pad  ;
	input \wb1m_data_i[10]_pad  ;
	input \wb1m_data_i[11]_pad  ;
	input \wb1m_data_i[12]_pad  ;
	input \wb1m_data_i[13]_pad  ;
	input \wb1m_data_i[14]_pad  ;
	input \wb1m_data_i[15]_pad  ;
	input \wb1m_data_i[16]_pad  ;
	input \wb1m_data_i[17]_pad  ;
	input \wb1m_data_i[18]_pad  ;
	input \wb1m_data_i[19]_pad  ;
	input \wb1m_data_i[1]_pad  ;
	input \wb1m_data_i[20]_pad  ;
	input \wb1m_data_i[21]_pad  ;
	input \wb1m_data_i[22]_pad  ;
	input \wb1m_data_i[23]_pad  ;
	input \wb1m_data_i[24]_pad  ;
	input \wb1m_data_i[25]_pad  ;
	input \wb1m_data_i[26]_pad  ;
	input \wb1m_data_i[27]_pad  ;
	input \wb1m_data_i[28]_pad  ;
	input \wb1m_data_i[29]_pad  ;
	input \wb1m_data_i[2]_pad  ;
	input \wb1m_data_i[30]_pad  ;
	input \wb1m_data_i[31]_pad  ;
	input \wb1m_data_i[3]_pad  ;
	input \wb1m_data_i[4]_pad  ;
	input \wb1m_data_i[5]_pad  ;
	input \wb1m_data_i[6]_pad  ;
	input \wb1m_data_i[7]_pad  ;
	input \wb1m_data_i[8]_pad  ;
	input \wb1m_data_i[9]_pad  ;
	input \wb1s_data_i[0]_pad  ;
	input \wb1s_data_i[10]_pad  ;
	input \wb1s_data_i[11]_pad  ;
	input \wb1s_data_i[12]_pad  ;
	input \wb1s_data_i[13]_pad  ;
	input \wb1s_data_i[14]_pad  ;
	input \wb1s_data_i[15]_pad  ;
	input \wb1s_data_i[16]_pad  ;
	input \wb1s_data_i[17]_pad  ;
	input \wb1s_data_i[18]_pad  ;
	input \wb1s_data_i[19]_pad  ;
	input \wb1s_data_i[1]_pad  ;
	input \wb1s_data_i[20]_pad  ;
	input \wb1s_data_i[21]_pad  ;
	input \wb1s_data_i[22]_pad  ;
	input \wb1s_data_i[23]_pad  ;
	input \wb1s_data_i[24]_pad  ;
	input \wb1s_data_i[25]_pad  ;
	input \wb1s_data_i[26]_pad  ;
	input \wb1s_data_i[27]_pad  ;
	input \wb1s_data_i[28]_pad  ;
	input \wb1s_data_i[29]_pad  ;
	input \wb1s_data_i[2]_pad  ;
	input \wb1s_data_i[30]_pad  ;
	input \wb1s_data_i[31]_pad  ;
	input \wb1s_data_i[3]_pad  ;
	input \wb1s_data_i[4]_pad  ;
	input \wb1s_data_i[5]_pad  ;
	input \wb1s_data_i[6]_pad  ;
	input \wb1s_data_i[7]_pad  ;
	input \wb1s_data_i[8]_pad  ;
	input \wb1s_data_i[9]_pad  ;
	output \_al_n0  ;
	output \_al_n1  ;
	output \g22594/_0_  ;
	output \g22595/_0_  ;
	output \g22599/_0_  ;
	output \g22600/_0_  ;
	output \g22606/_0_  ;
	output \g22607/_0_  ;
	output \g22610/_0_  ;
	output \g22614/_0_  ;
	output \g22615/_0_  ;
	output \g22616/_0_  ;
	output \g22619/_0_  ;
	output \g22620/_0_  ;
	output \g22626/_0_  ;
	output \g22635/_0_  ;
	output \g22650/_0_  ;
	output \g22651/_0_  ;
	output \g22692/_0_  ;
	output \g22727/_0_  ;
	output \g22729/_3_  ;
	output \g22774/_0_  ;
	output \g22775/_0_  ;
	output \g22776/_0_  ;
	output \g22777/_0_  ;
	output \g22779/_3_  ;
	output \g22780/_0_  ;
	output \g22781/_0_  ;
	output \g22782/_0_  ;
	output \g22784/_0_  ;
	output \g22785/_0_  ;
	output \g22786/_0_  ;
	output \g22787/_0_  ;
	output \g22789/_3_  ;
	output \g22790/_0_  ;
	output \g22791/_0_  ;
	output \g22792/_0_  ;
	output \g22793/_0_  ;
	output \g22794/_0_  ;
	output \g22795/_0_  ;
	output \g22796/_0_  ;
	output \g22797/_0_  ;
	output \g22798/_0_  ;
	output \g22799/_0_  ;
	output \g22838/_0_  ;
	output \g22839/_0_  ;
	output \g22841/_0_  ;
	output \g22842/_0_  ;
	output \g22847/_0_  ;
	output \g22848/_0_  ;
	output \g22849/_0_  ;
	output \g22850/_0_  ;
	output \g22851/_0_  ;
	output \g22852/_0_  ;
	output \g22853/_0_  ;
	output \g22854/_0_  ;
	output \g22855/_0_  ;
	output \g22856/_0_  ;
	output \g22857/_0_  ;
	output \g22858/_0_  ;
	output \g22859/_0_  ;
	output \g22860/_0_  ;
	output \g22861/_0_  ;
	output \g22862/_0_  ;
	output \g22863/_0_  ;
	output \g22864/_0_  ;
	output \g22865/_0_  ;
	output \g22867/_0_  ;
	output \g22868/_0_  ;
	output \g22869/_0_  ;
	output \g22871/_0_  ;
	output \g22872/_0_  ;
	output \g22873/_0_  ;
	output \g22874/_0_  ;
	output \g22875/_0_  ;
	output \g22876/_0_  ;
	output \g22878/_0_  ;
	output \g22882/_2_  ;
	output \g22995/_0_  ;
	output \g23030/_0_  ;
	output \g23046/_0_  ;
	output \g23077/_0_  ;
	output \g23111/_0_  ;
	output \g23115/_1_  ;
	output \g23124/_2_  ;
	output \g23126/_2_  ;
	output \g23128/_2_  ;
	output \g23130/_2_  ;
	output \g23132/_2_  ;
	output \g23134/_2_  ;
	output \g23136/_2_  ;
	output \g23137/_0_  ;
	output \g23140/_2_  ;
	output \g23142/_2_  ;
	output \g23144/_2_  ;
	output \g23146/_2_  ;
	output \g23148/_2_  ;
	output \g23150/_2_  ;
	output \g23152/_2_  ;
	output \g23154/_2_  ;
	output \g23156/_2_  ;
	output \g23158/_2_  ;
	output \g23160/_2_  ;
	output \g23162/_2_  ;
	output \g23163/_3_  ;
	output \g23164/_0_  ;
	output \g23166/_0_  ;
	output \g23168/_0_  ;
	output \g23170/_2_  ;
	output \g23172/_2_  ;
	output \g23174/_2_  ;
	output \g23175/_0_  ;
	output \g23177/_0_  ;
	output \g23180/_2_  ;
	output \g23220/_0_  ;
	output \g23238/_0_  ;
	output \g23239/_0_  ;
	output \g23240/_0_  ;
	output \g23241/_0_  ;
	output \g23242/_0_  ;
	output \g23243/_0_  ;
	output \g23244/_0_  ;
	output \g23245/_0_  ;
	output \g23247/_3_  ;
	output \g23248/_0_  ;
	output \g23249/_0_  ;
	output \g23250/_0_  ;
	output \g23251/_0_  ;
	output \g23252/_0_  ;
	output \g23253/_0_  ;
	output \g23255/_3_  ;
	output \g23260/_0_  ;
	output \g23284/_3_  ;
	output \g23285/_0_  ;
	output \g23334/_0_  ;
	output \g23343/_0_  ;
	output \g23366/_0_  ;
	output \g23402/_0_  ;
	output \g23403/_0_  ;
	output \g23404/_0_  ;
	output \g23405/_0_  ;
	output \g23407/_0_  ;
	output \g23408/_0_  ;
	output \g23409/_0_  ;
	output \g23410/_0_  ;
	output \g23411/_0_  ;
	output \g23413/_2_  ;
	output \g23415/_2_  ;
	output \g23417/_2_  ;
	output \g23542/_0_  ;
	output \g23607/_0_  ;
	output \g23608/_0_  ;
	output \g23609/_3_  ;
	output \g23707/_0_  ;
	output \g23708/_0_  ;
	output \g23709/_0_  ;
	output \g23710/_0_  ;
	output \g23711/_0_  ;
	output \g23712/_0_  ;
	output \g23713/_0_  ;
	output \g23714/_0_  ;
	output \g23715/_0_  ;
	output \g23716/_0_  ;
	output \g23754/_0_  ;
	output \g23755/_0_  ;
	output \g23756/_0_  ;
	output \g23757/_0_  ;
	output \g23758/_0_  ;
	output \g23759/_0_  ;
	output \g23760/_0_  ;
	output \g23761/_0_  ;
	output \g23763/_3_  ;
	output \g23767/_0_  ;
	output \g23768/_0_  ;
	output \g23833/_0_  ;
	output \g23837/_0_  ;
	output \g23838/_0_  ;
	output \g23839/_0_  ;
	output \g23840/_0_  ;
	output \g23841/_0_  ;
	output \g23842/_0_  ;
	output \g23843/_0_  ;
	output \g23844/_0_  ;
	output \g23845/_0_  ;
	output \g23849/_3_  ;
	output \g23851/_3_  ;
	output \g23858/_0_  ;
	output \g23870/_0_  ;
	output \g23871/_0_  ;
	output \g23872/_3_  ;
	output \g23873/_3_  ;
	output \g23874/_3_  ;
	output \g23875/_3_  ;
	output \g23876/_3_  ;
	output \g23877/_3_  ;
	output \g23878/_3_  ;
	output \g23879/_3_  ;
	output \g23880/_3_  ;
	output \g23881/_3_  ;
	output \g23882/_3_  ;
	output \g23883/_3_  ;
	output \g23884/_3_  ;
	output \g23885/_3_  ;
	output \g23886/_3_  ;
	output \g23887/_3_  ;
	output \g23888/_3_  ;
	output \g23889/_3_  ;
	output \g23890/_3_  ;
	output \g23891/_3_  ;
	output \g23892/_3_  ;
	output \g23893/_3_  ;
	output \g23894/_3_  ;
	output \g23895/_3_  ;
	output \g23896/_3_  ;
	output \g23897/_3_  ;
	output \g23898/_3_  ;
	output \g23899/_3_  ;
	output \g23900/_3_  ;
	output \g23901/_3_  ;
	output \g23902/_3_  ;
	output \g23903/_3_  ;
	output \g23904/_3_  ;
	output \g23905/_3_  ;
	output \g23906/_3_  ;
	output \g23907/_3_  ;
	output \g23908/_3_  ;
	output \g23909/_3_  ;
	output \g23910/_3_  ;
	output \g23911/_3_  ;
	output \g23912/_3_  ;
	output \g23913/_3_  ;
	output \g23914/_3_  ;
	output \g23915/_3_  ;
	output \g23959/_0_  ;
	output \g23961/_0_  ;
	output \g23962/_0_  ;
	output \g23966/_0_  ;
	output \g23967/_0_  ;
	output \g23969/_0_  ;
	output \g23970/_0_  ;
	output \g23971/_0_  ;
	output \g23972/_0_  ;
	output \g23979/_0_  ;
	output \g23987/_0_  ;
	output \g23988/_0_  ;
	output \g23989/_0_  ;
	output \g23990/_0_  ;
	output \g24005/_0_  ;
	output \g24010/_0_  ;
	output \g24012/_0_  ;
	output \g24013/_0_  ;
	output \g24014/_0_  ;
	output \g24015/_0_  ;
	output \g24016/_0_  ;
	output \g24017/_0_  ;
	output \g24018/_0_  ;
	output \g24019/_0_  ;
	output \g24020/_0_  ;
	output \g24026/_0_  ;
	output \g24027/_0_  ;
	output \g24028/_0_  ;
	output \g24029/_0_  ;
	output \g24030/_0_  ;
	output \g24031/_0_  ;
	output \g24032/_0_  ;
	output \g24033/_0_  ;
	output \g24034/_0_  ;
	output \g24035/_0_  ;
	output \g24036/_0_  ;
	output \g24037/_0_  ;
	output \g24038/_0_  ;
	output \g24039/_0_  ;
	output \g24042/_0_  ;
	output \g24049/_0_  ;
	output \g24063/_0_  ;
	output \g24119/_0_  ;
	output \g24120/_0_  ;
	output \g24357/_0_  ;
	output \g24432/_0_  ;
	output \g24433/_0_  ;
	output \g24437/_0_  ;
	output \g24438/_0_  ;
	output \g24477/_0_  ;
	output \g24491/_0_  ;
	output \g24530/_2_  ;
	output \g24532/_0_  ;
	output \g24534/_0_  ;
	output \g24537/_0_  ;
	output \g24538/_0_  ;
	output \g24539/_0_  ;
	output \g24540/_0_  ;
	output \g24606/_2_  ;
	output \g24612/_0_  ;
	output \g24677/_0_  ;
	output \g24678/_0_  ;
	output \g24679/_0_  ;
	output \g24688/_0_  ;
	output \g24743/_0_  ;
	output \g24847/_0_  ;
	output \g24849/_0_  ;
	output \g24850/_0_  ;
	output \g24854/_0_  ;
	output \g24862/_0_  ;
	output \g24872/_0_  ;
	output \g24873/_0_  ;
	output \g24874/_0_  ;
	output \g24876/_0_  ;
	output \g24879/_0_  ;
	output \g24880/_0_  ;
	output \g24881/_0_  ;
	output \g24882/_0_  ;
	output \g24952/_2_  ;
	output \g24976/_1_  ;
	output \g25003/_0_  ;
	output \g25004/_0_  ;
	output \g25005/_0_  ;
	output \g25006/_0_  ;
	output \g25011/_0_  ;
	output \g25012/_0_  ;
	output \g25013/_0_  ;
	output \g25031/_0_  ;
	output \g25032/_0_  ;
	output \g25033/_0_  ;
	output \g25034/_0_  ;
	output \g25035/_0_  ;
	output \g25153/_2_  ;
	output \g25183/_0_  ;
	output \g25184/_0_  ;
	output \g25224/_0_  ;
	output \g25232/_0_  ;
	output \g25237/_0_  ;
	output \g25241/_2_  ;
	output \g25243/_2_  ;
	output \g25248/_3_  ;
	output \g25261/_0_  ;
	output \g25262/_0_  ;
	output \g25266/_3_  ;
	output \g25267/_0_  ;
	output \g25269/_0_  ;
	output \g25543/_1_  ;
	output \g25602/_3_  ;
	output \g25610/_0_  ;
	output \g25611/_0_  ;
	output \g25841/_0_  ;
	output \g25843/_0_  ;
	output \g25893/_0_  ;
	output \g27013/_0_  ;
	output \g27060/_0_  ;
	output \g27073/_0_  ;
	output \g27184/_0_  ;
	output \g27186/_0_  ;
	output \g27189/_2_  ;
	output \g47/_0_  ;
	output \u0_u0_ch_done_reg/_05_  ;
	output \u2_adr0_cnt_reg[0]/P0000  ;
	output \u2_adr1_cnt_reg[0]/P0000  ;
	output \u3_u0_mast_we_r_reg/_05_  ;
	output \wb0_ack_o_pad  ;
	output \wb0_addr_o[0]_pad  ;
	output \wb0_addr_o[10]_pad  ;
	output \wb0_addr_o[11]_pad  ;
	output \wb0_addr_o[12]_pad  ;
	output \wb0_addr_o[13]_pad  ;
	output \wb0_addr_o[14]_pad  ;
	output \wb0_addr_o[15]_pad  ;
	output \wb0_addr_o[16]_pad  ;
	output \wb0_addr_o[17]_pad  ;
	output \wb0_addr_o[18]_pad  ;
	output \wb0_addr_o[19]_pad  ;
	output \wb0_addr_o[1]_pad  ;
	output \wb0_addr_o[20]_pad  ;
	output \wb0_addr_o[21]_pad  ;
	output \wb0_addr_o[22]_pad  ;
	output \wb0_addr_o[23]_pad  ;
	output \wb0_addr_o[24]_pad  ;
	output \wb0_addr_o[25]_pad  ;
	output \wb0_addr_o[26]_pad  ;
	output \wb0_addr_o[27]_pad  ;
	output \wb0_addr_o[28]_pad  ;
	output \wb0_addr_o[29]_pad  ;
	output \wb0_addr_o[2]_pad  ;
	output \wb0_addr_o[30]_pad  ;
	output \wb0_addr_o[31]_pad  ;
	output \wb0_addr_o[3]_pad  ;
	output \wb0_addr_o[4]_pad  ;
	output \wb0_addr_o[5]_pad  ;
	output \wb0_addr_o[6]_pad  ;
	output \wb0_addr_o[7]_pad  ;
	output \wb0_addr_o[8]_pad  ;
	output \wb0_addr_o[9]_pad  ;
	output \wb0_cyc_o_pad  ;
	output \wb0_err_o_pad  ;
	output \wb0_rty_o_pad  ;
	output \wb0_sel_o[0]_pad  ;
	output \wb0_sel_o[1]_pad  ;
	output \wb0_sel_o[2]_pad  ;
	output \wb0_sel_o[3]_pad  ;
	output \wb0_stb_o_pad  ;
	output \wb0_we_o_pad  ;
	output \wb0m_data_o[0]_pad  ;
	output \wb0m_data_o[10]_pad  ;
	output \wb0m_data_o[11]_pad  ;
	output \wb0m_data_o[12]_pad  ;
	output \wb0m_data_o[13]_pad  ;
	output \wb0m_data_o[14]_pad  ;
	output \wb0m_data_o[15]_pad  ;
	output \wb0m_data_o[16]_pad  ;
	output \wb0m_data_o[17]_pad  ;
	output \wb0m_data_o[18]_pad  ;
	output \wb0m_data_o[19]_pad  ;
	output \wb0m_data_o[1]_pad  ;
	output \wb0m_data_o[20]_pad  ;
	output \wb0m_data_o[21]_pad  ;
	output \wb0m_data_o[22]_pad  ;
	output \wb0m_data_o[23]_pad  ;
	output \wb0m_data_o[24]_pad  ;
	output \wb0m_data_o[25]_pad  ;
	output \wb0m_data_o[26]_pad  ;
	output \wb0m_data_o[27]_pad  ;
	output \wb0m_data_o[28]_pad  ;
	output \wb0m_data_o[29]_pad  ;
	output \wb0m_data_o[2]_pad  ;
	output \wb0m_data_o[30]_pad  ;
	output \wb0m_data_o[31]_pad  ;
	output \wb0m_data_o[3]_pad  ;
	output \wb0m_data_o[4]_pad  ;
	output \wb0m_data_o[5]_pad  ;
	output \wb0m_data_o[6]_pad  ;
	output \wb0m_data_o[7]_pad  ;
	output \wb0m_data_o[8]_pad  ;
	output \wb0m_data_o[9]_pad  ;
	output \wb0s_data_o[0]_pad  ;
	output \wb0s_data_o[10]_pad  ;
	output \wb0s_data_o[11]_pad  ;
	output \wb0s_data_o[12]_pad  ;
	output \wb0s_data_o[13]_pad  ;
	output \wb0s_data_o[14]_pad  ;
	output \wb0s_data_o[15]_pad  ;
	output \wb0s_data_o[16]_pad  ;
	output \wb0s_data_o[17]_pad  ;
	output \wb0s_data_o[18]_pad  ;
	output \wb0s_data_o[19]_pad  ;
	output \wb0s_data_o[1]_pad  ;
	output \wb0s_data_o[20]_pad  ;
	output \wb0s_data_o[21]_pad  ;
	output \wb0s_data_o[22]_pad  ;
	output \wb0s_data_o[23]_pad  ;
	output \wb0s_data_o[24]_pad  ;
	output \wb0s_data_o[25]_pad  ;
	output \wb0s_data_o[26]_pad  ;
	output \wb0s_data_o[27]_pad  ;
	output \wb0s_data_o[28]_pad  ;
	output \wb0s_data_o[29]_pad  ;
	output \wb0s_data_o[2]_pad  ;
	output \wb0s_data_o[30]_pad  ;
	output \wb0s_data_o[31]_pad  ;
	output \wb0s_data_o[3]_pad  ;
	output \wb0s_data_o[4]_pad  ;
	output \wb0s_data_o[5]_pad  ;
	output \wb0s_data_o[6]_pad  ;
	output \wb0s_data_o[7]_pad  ;
	output \wb0s_data_o[8]_pad  ;
	output \wb0s_data_o[9]_pad  ;
	output \wb1_ack_o_pad  ;
	output \wb1_addr_o[0]_pad  ;
	output \wb1_addr_o[10]_pad  ;
	output \wb1_addr_o[11]_pad  ;
	output \wb1_addr_o[12]_pad  ;
	output \wb1_addr_o[13]_pad  ;
	output \wb1_addr_o[14]_pad  ;
	output \wb1_addr_o[15]_pad  ;
	output \wb1_addr_o[16]_pad  ;
	output \wb1_addr_o[17]_pad  ;
	output \wb1_addr_o[18]_pad  ;
	output \wb1_addr_o[19]_pad  ;
	output \wb1_addr_o[1]_pad  ;
	output \wb1_addr_o[20]_pad  ;
	output \wb1_addr_o[21]_pad  ;
	output \wb1_addr_o[22]_pad  ;
	output \wb1_addr_o[23]_pad  ;
	output \wb1_addr_o[24]_pad  ;
	output \wb1_addr_o[25]_pad  ;
	output \wb1_addr_o[26]_pad  ;
	output \wb1_addr_o[27]_pad  ;
	output \wb1_addr_o[28]_pad  ;
	output \wb1_addr_o[29]_pad  ;
	output \wb1_addr_o[2]_pad  ;
	output \wb1_addr_o[30]_pad  ;
	output \wb1_addr_o[31]_pad  ;
	output \wb1_addr_o[3]_pad  ;
	output \wb1_addr_o[4]_pad  ;
	output \wb1_addr_o[5]_pad  ;
	output \wb1_addr_o[6]_pad  ;
	output \wb1_addr_o[7]_pad  ;
	output \wb1_addr_o[8]_pad  ;
	output \wb1_addr_o[9]_pad  ;
	output \wb1_cyc_o_pad  ;
	output \wb1_err_o_pad  ;
	output \wb1_rty_o_pad  ;
	output \wb1_sel_o[0]_pad  ;
	output \wb1_sel_o[1]_pad  ;
	output \wb1_sel_o[2]_pad  ;
	output \wb1_sel_o[3]_pad  ;
	output \wb1_stb_o_pad  ;
	output \wb1_we_o_pad  ;
	output \wb1m_data_o[0]_pad  ;
	output \wb1m_data_o[10]_pad  ;
	output \wb1m_data_o[11]_pad  ;
	output \wb1m_data_o[12]_pad  ;
	output \wb1m_data_o[13]_pad  ;
	output \wb1m_data_o[14]_pad  ;
	output \wb1m_data_o[15]_pad  ;
	output \wb1m_data_o[16]_pad  ;
	output \wb1m_data_o[17]_pad  ;
	output \wb1m_data_o[18]_pad  ;
	output \wb1m_data_o[19]_pad  ;
	output \wb1m_data_o[1]_pad  ;
	output \wb1m_data_o[20]_pad  ;
	output \wb1m_data_o[21]_pad  ;
	output \wb1m_data_o[22]_pad  ;
	output \wb1m_data_o[23]_pad  ;
	output \wb1m_data_o[24]_pad  ;
	output \wb1m_data_o[25]_pad  ;
	output \wb1m_data_o[26]_pad  ;
	output \wb1m_data_o[27]_pad  ;
	output \wb1m_data_o[28]_pad  ;
	output \wb1m_data_o[29]_pad  ;
	output \wb1m_data_o[2]_pad  ;
	output \wb1m_data_o[30]_pad  ;
	output \wb1m_data_o[31]_pad  ;
	output \wb1m_data_o[3]_pad  ;
	output \wb1m_data_o[4]_pad  ;
	output \wb1m_data_o[5]_pad  ;
	output \wb1m_data_o[6]_pad  ;
	output \wb1m_data_o[7]_pad  ;
	output \wb1m_data_o[8]_pad  ;
	output \wb1m_data_o[9]_pad  ;
	output \wb1s_data_o[0]_pad  ;
	output \wb1s_data_o[10]_pad  ;
	output \wb1s_data_o[11]_pad  ;
	output \wb1s_data_o[12]_pad  ;
	output \wb1s_data_o[13]_pad  ;
	output \wb1s_data_o[14]_pad  ;
	output \wb1s_data_o[15]_pad  ;
	output \wb1s_data_o[16]_pad  ;
	output \wb1s_data_o[17]_pad  ;
	output \wb1s_data_o[18]_pad  ;
	output \wb1s_data_o[19]_pad  ;
	output \wb1s_data_o[1]_pad  ;
	output \wb1s_data_o[20]_pad  ;
	output \wb1s_data_o[21]_pad  ;
	output \wb1s_data_o[22]_pad  ;
	output \wb1s_data_o[23]_pad  ;
	output \wb1s_data_o[24]_pad  ;
	output \wb1s_data_o[25]_pad  ;
	output \wb1s_data_o[26]_pad  ;
	output \wb1s_data_o[27]_pad  ;
	output \wb1s_data_o[28]_pad  ;
	output \wb1s_data_o[29]_pad  ;
	output \wb1s_data_o[2]_pad  ;
	output \wb1s_data_o[30]_pad  ;
	output \wb1s_data_o[31]_pad  ;
	output \wb1s_data_o[3]_pad  ;
	output \wb1s_data_o[4]_pad  ;
	output \wb1s_data_o[5]_pad  ;
	output \wb1s_data_o[6]_pad  ;
	output \wb1s_data_o[7]_pad  ;
	output \wb1s_data_o[8]_pad  ;
	output \wb1s_data_o[9]_pad  ;
	wire _w2765_ ;
	wire _w2764_ ;
	wire _w2763_ ;
	wire _w2762_ ;
	wire _w2761_ ;
	wire _w2760_ ;
	wire _w2759_ ;
	wire _w2758_ ;
	wire _w2757_ ;
	wire _w2756_ ;
	wire _w2755_ ;
	wire _w2754_ ;
	wire _w2753_ ;
	wire _w2752_ ;
	wire _w2751_ ;
	wire _w2750_ ;
	wire _w2749_ ;
	wire _w2748_ ;
	wire _w2747_ ;
	wire _w2746_ ;
	wire _w2745_ ;
	wire _w2744_ ;
	wire _w2743_ ;
	wire _w2742_ ;
	wire _w2741_ ;
	wire _w2740_ ;
	wire _w2739_ ;
	wire _w2738_ ;
	wire _w2737_ ;
	wire _w2736_ ;
	wire _w2735_ ;
	wire _w2734_ ;
	wire _w2733_ ;
	wire _w2732_ ;
	wire _w2731_ ;
	wire _w2730_ ;
	wire _w2729_ ;
	wire _w2728_ ;
	wire _w2727_ ;
	wire _w2726_ ;
	wire _w2725_ ;
	wire _w2724_ ;
	wire _w2723_ ;
	wire _w2722_ ;
	wire _w2721_ ;
	wire _w2720_ ;
	wire _w2719_ ;
	wire _w2718_ ;
	wire _w2717_ ;
	wire _w2716_ ;
	wire _w2715_ ;
	wire _w2714_ ;
	wire _w2713_ ;
	wire _w2712_ ;
	wire _w2711_ ;
	wire _w2710_ ;
	wire _w2709_ ;
	wire _w2708_ ;
	wire _w2707_ ;
	wire _w2706_ ;
	wire _w2705_ ;
	wire _w2704_ ;
	wire _w2703_ ;
	wire _w2702_ ;
	wire _w2701_ ;
	wire _w2700_ ;
	wire _w2699_ ;
	wire _w2698_ ;
	wire _w2697_ ;
	wire _w2696_ ;
	wire _w2695_ ;
	wire _w2694_ ;
	wire _w2693_ ;
	wire _w2692_ ;
	wire _w2691_ ;
	wire _w2690_ ;
	wire _w2689_ ;
	wire _w2688_ ;
	wire _w2687_ ;
	wire _w2686_ ;
	wire _w2685_ ;
	wire _w2684_ ;
	wire _w2683_ ;
	wire _w2682_ ;
	wire _w2681_ ;
	wire _w2680_ ;
	wire _w2679_ ;
	wire _w2678_ ;
	wire _w2677_ ;
	wire _w2676_ ;
	wire _w2675_ ;
	wire _w2674_ ;
	wire _w2673_ ;
	wire _w2672_ ;
	wire _w2671_ ;
	wire _w2670_ ;
	wire _w2669_ ;
	wire _w2668_ ;
	wire _w2667_ ;
	wire _w2666_ ;
	wire _w2665_ ;
	wire _w2664_ ;
	wire _w2663_ ;
	wire _w2662_ ;
	wire _w2661_ ;
	wire _w2660_ ;
	wire _w2659_ ;
	wire _w2658_ ;
	wire _w2657_ ;
	wire _w2656_ ;
	wire _w2655_ ;
	wire _w2654_ ;
	wire _w2653_ ;
	wire _w2652_ ;
	wire _w2651_ ;
	wire _w2650_ ;
	wire _w2649_ ;
	wire _w2648_ ;
	wire _w2647_ ;
	wire _w2646_ ;
	wire _w2645_ ;
	wire _w2644_ ;
	wire _w2643_ ;
	wire _w2642_ ;
	wire _w2641_ ;
	wire _w2640_ ;
	wire _w2639_ ;
	wire _w2638_ ;
	wire _w2637_ ;
	wire _w2636_ ;
	wire _w2635_ ;
	wire _w2634_ ;
	wire _w2633_ ;
	wire _w2632_ ;
	wire _w2631_ ;
	wire _w2630_ ;
	wire _w2629_ ;
	wire _w2628_ ;
	wire _w2627_ ;
	wire _w2626_ ;
	wire _w2625_ ;
	wire _w2624_ ;
	wire _w2623_ ;
	wire _w2622_ ;
	wire _w2621_ ;
	wire _w2620_ ;
	wire _w2619_ ;
	wire _w2618_ ;
	wire _w2617_ ;
	wire _w2616_ ;
	wire _w2615_ ;
	wire _w2614_ ;
	wire _w2613_ ;
	wire _w2612_ ;
	wire _w2611_ ;
	wire _w2610_ ;
	wire _w2609_ ;
	wire _w2608_ ;
	wire _w2607_ ;
	wire _w2606_ ;
	wire _w2605_ ;
	wire _w2604_ ;
	wire _w2603_ ;
	wire _w2602_ ;
	wire _w2601_ ;
	wire _w2599_ ;
	wire _w2598_ ;
	wire _w2597_ ;
	wire _w2596_ ;
	wire _w2595_ ;
	wire _w2594_ ;
	wire _w2593_ ;
	wire _w2592_ ;
	wire _w2591_ ;
	wire _w2590_ ;
	wire _w2589_ ;
	wire _w2588_ ;
	wire _w2587_ ;
	wire _w2586_ ;
	wire _w2585_ ;
	wire _w2584_ ;
	wire _w2583_ ;
	wire _w2582_ ;
	wire _w2581_ ;
	wire _w2580_ ;
	wire _w2579_ ;
	wire _w2578_ ;
	wire _w2577_ ;
	wire _w2576_ ;
	wire _w2575_ ;
	wire _w2574_ ;
	wire _w2573_ ;
	wire _w2572_ ;
	wire _w2571_ ;
	wire _w2570_ ;
	wire _w2568_ ;
	wire _w2567_ ;
	wire _w2566_ ;
	wire _w2565_ ;
	wire _w2564_ ;
	wire _w2563_ ;
	wire _w2562_ ;
	wire _w2561_ ;
	wire _w2560_ ;
	wire _w2559_ ;
	wire _w2558_ ;
	wire _w2557_ ;
	wire _w2556_ ;
	wire _w2555_ ;
	wire _w2554_ ;
	wire _w2553_ ;
	wire _w2552_ ;
	wire _w2551_ ;
	wire _w2550_ ;
	wire _w2549_ ;
	wire _w2548_ ;
	wire _w2547_ ;
	wire _w2546_ ;
	wire _w2545_ ;
	wire _w2544_ ;
	wire _w2543_ ;
	wire _w2542_ ;
	wire _w2541_ ;
	wire _w2540_ ;
	wire _w2539_ ;
	wire _w2538_ ;
	wire _w2537_ ;
	wire _w2536_ ;
	wire _w2535_ ;
	wire _w2534_ ;
	wire _w2533_ ;
	wire _w2532_ ;
	wire _w2531_ ;
	wire _w2530_ ;
	wire _w2529_ ;
	wire _w2528_ ;
	wire _w2527_ ;
	wire _w2526_ ;
	wire _w2525_ ;
	wire _w2524_ ;
	wire _w2523_ ;
	wire _w2522_ ;
	wire _w2521_ ;
	wire _w2520_ ;
	wire _w2519_ ;
	wire _w2518_ ;
	wire _w2517_ ;
	wire _w2516_ ;
	wire _w2515_ ;
	wire _w2514_ ;
	wire _w2513_ ;
	wire _w2512_ ;
	wire _w2511_ ;
	wire _w2510_ ;
	wire _w2509_ ;
	wire _w2508_ ;
	wire _w2507_ ;
	wire _w2506_ ;
	wire _w2505_ ;
	wire _w2504_ ;
	wire _w2503_ ;
	wire _w2502_ ;
	wire _w2501_ ;
	wire _w2500_ ;
	wire _w2499_ ;
	wire _w2498_ ;
	wire _w2497_ ;
	wire _w2496_ ;
	wire _w2495_ ;
	wire _w2494_ ;
	wire _w2493_ ;
	wire _w2492_ ;
	wire _w2491_ ;
	wire _w2490_ ;
	wire _w2489_ ;
	wire _w2488_ ;
	wire _w2487_ ;
	wire _w2486_ ;
	wire _w2485_ ;
	wire _w2484_ ;
	wire _w2483_ ;
	wire _w2482_ ;
	wire _w2481_ ;
	wire _w2480_ ;
	wire _w2479_ ;
	wire _w2478_ ;
	wire _w2477_ ;
	wire _w2476_ ;
	wire _w2475_ ;
	wire _w2474_ ;
	wire _w2473_ ;
	wire _w2472_ ;
	wire _w2471_ ;
	wire _w2470_ ;
	wire _w2469_ ;
	wire _w2468_ ;
	wire _w2467_ ;
	wire _w2466_ ;
	wire _w2465_ ;
	wire _w2464_ ;
	wire _w2463_ ;
	wire _w2462_ ;
	wire _w2461_ ;
	wire _w2460_ ;
	wire _w2459_ ;
	wire _w2458_ ;
	wire _w2457_ ;
	wire _w2456_ ;
	wire _w2455_ ;
	wire _w2454_ ;
	wire _w2453_ ;
	wire _w2452_ ;
	wire _w2451_ ;
	wire _w2450_ ;
	wire _w2449_ ;
	wire _w2448_ ;
	wire _w2447_ ;
	wire _w2446_ ;
	wire _w2445_ ;
	wire _w2444_ ;
	wire _w2443_ ;
	wire _w2442_ ;
	wire _w2441_ ;
	wire _w2440_ ;
	wire _w2439_ ;
	wire _w2438_ ;
	wire _w2437_ ;
	wire _w2436_ ;
	wire _w2435_ ;
	wire _w2434_ ;
	wire _w2433_ ;
	wire _w2432_ ;
	wire _w2431_ ;
	wire _w2430_ ;
	wire _w2429_ ;
	wire _w2428_ ;
	wire _w2427_ ;
	wire _w2426_ ;
	wire _w2425_ ;
	wire _w2424_ ;
	wire _w2423_ ;
	wire _w2422_ ;
	wire _w2421_ ;
	wire _w2420_ ;
	wire _w2419_ ;
	wire _w2418_ ;
	wire _w2417_ ;
	wire _w2416_ ;
	wire _w2415_ ;
	wire _w2414_ ;
	wire _w2413_ ;
	wire _w2412_ ;
	wire _w2411_ ;
	wire _w2410_ ;
	wire _w2409_ ;
	wire _w2408_ ;
	wire _w2407_ ;
	wire _w2406_ ;
	wire _w2405_ ;
	wire _w2404_ ;
	wire _w2403_ ;
	wire _w2402_ ;
	wire _w2401_ ;
	wire _w2400_ ;
	wire _w2399_ ;
	wire _w2398_ ;
	wire _w2397_ ;
	wire _w2396_ ;
	wire _w2395_ ;
	wire _w2394_ ;
	wire _w2393_ ;
	wire _w2392_ ;
	wire _w2391_ ;
	wire _w2390_ ;
	wire _w2389_ ;
	wire _w2388_ ;
	wire _w2387_ ;
	wire _w2386_ ;
	wire _w2385_ ;
	wire _w2384_ ;
	wire _w2383_ ;
	wire _w2382_ ;
	wire _w2381_ ;
	wire _w2380_ ;
	wire _w2379_ ;
	wire _w2378_ ;
	wire _w2377_ ;
	wire _w2376_ ;
	wire _w2375_ ;
	wire _w2374_ ;
	wire _w2373_ ;
	wire _w2372_ ;
	wire _w2371_ ;
	wire _w2370_ ;
	wire _w2369_ ;
	wire _w2368_ ;
	wire _w2367_ ;
	wire _w2366_ ;
	wire _w2365_ ;
	wire _w2364_ ;
	wire _w2363_ ;
	wire _w2362_ ;
	wire _w2361_ ;
	wire _w2360_ ;
	wire _w2359_ ;
	wire _w2358_ ;
	wire _w2357_ ;
	wire _w2356_ ;
	wire _w2355_ ;
	wire _w2354_ ;
	wire _w2353_ ;
	wire _w2352_ ;
	wire _w2351_ ;
	wire _w2350_ ;
	wire _w2349_ ;
	wire _w2348_ ;
	wire _w2347_ ;
	wire _w2346_ ;
	wire _w2345_ ;
	wire _w2344_ ;
	wire _w2343_ ;
	wire _w2342_ ;
	wire _w2341_ ;
	wire _w2340_ ;
	wire _w2339_ ;
	wire _w2338_ ;
	wire _w2337_ ;
	wire _w2336_ ;
	wire _w2335_ ;
	wire _w2334_ ;
	wire _w2333_ ;
	wire _w2332_ ;
	wire _w2331_ ;
	wire _w2330_ ;
	wire _w2329_ ;
	wire _w2328_ ;
	wire _w2327_ ;
	wire _w2326_ ;
	wire _w2325_ ;
	wire _w2324_ ;
	wire _w2323_ ;
	wire _w2322_ ;
	wire _w2321_ ;
	wire _w2320_ ;
	wire _w2319_ ;
	wire _w2318_ ;
	wire _w2317_ ;
	wire _w2316_ ;
	wire _w2315_ ;
	wire _w2314_ ;
	wire _w2313_ ;
	wire _w2312_ ;
	wire _w2311_ ;
	wire _w2310_ ;
	wire _w2309_ ;
	wire _w2308_ ;
	wire _w2307_ ;
	wire _w2306_ ;
	wire _w2305_ ;
	wire _w2304_ ;
	wire _w2303_ ;
	wire _w2302_ ;
	wire _w2301_ ;
	wire _w2300_ ;
	wire _w2299_ ;
	wire _w2298_ ;
	wire _w2297_ ;
	wire _w2296_ ;
	wire _w2295_ ;
	wire _w2294_ ;
	wire _w2293_ ;
	wire _w2292_ ;
	wire _w2291_ ;
	wire _w2290_ ;
	wire _w2289_ ;
	wire _w2288_ ;
	wire _w2287_ ;
	wire _w2286_ ;
	wire _w2285_ ;
	wire _w2284_ ;
	wire _w2283_ ;
	wire _w2282_ ;
	wire _w2281_ ;
	wire _w2280_ ;
	wire _w2279_ ;
	wire _w2278_ ;
	wire _w2277_ ;
	wire _w2276_ ;
	wire _w2275_ ;
	wire _w2274_ ;
	wire _w2273_ ;
	wire _w2272_ ;
	wire _w2271_ ;
	wire _w2270_ ;
	wire _w2269_ ;
	wire _w2268_ ;
	wire _w2267_ ;
	wire _w2266_ ;
	wire _w2265_ ;
	wire _w2264_ ;
	wire _w2263_ ;
	wire _w2262_ ;
	wire _w2261_ ;
	wire _w2260_ ;
	wire _w2259_ ;
	wire _w2258_ ;
	wire _w2257_ ;
	wire _w2256_ ;
	wire _w2255_ ;
	wire _w2254_ ;
	wire _w2253_ ;
	wire _w2252_ ;
	wire _w2251_ ;
	wire _w2250_ ;
	wire _w2249_ ;
	wire _w2248_ ;
	wire _w2247_ ;
	wire _w2246_ ;
	wire _w2245_ ;
	wire _w2244_ ;
	wire _w2243_ ;
	wire _w2242_ ;
	wire _w2241_ ;
	wire _w2240_ ;
	wire _w2239_ ;
	wire _w2238_ ;
	wire _w2237_ ;
	wire _w2236_ ;
	wire _w2235_ ;
	wire _w2234_ ;
	wire _w2233_ ;
	wire _w2232_ ;
	wire _w2231_ ;
	wire _w2230_ ;
	wire _w2229_ ;
	wire _w2228_ ;
	wire _w2227_ ;
	wire _w2226_ ;
	wire _w2225_ ;
	wire _w2224_ ;
	wire _w2223_ ;
	wire _w2222_ ;
	wire _w2221_ ;
	wire _w2220_ ;
	wire _w2219_ ;
	wire _w2218_ ;
	wire _w2217_ ;
	wire _w2216_ ;
	wire _w2215_ ;
	wire _w2214_ ;
	wire _w2213_ ;
	wire _w2212_ ;
	wire _w2211_ ;
	wire _w2210_ ;
	wire _w2209_ ;
	wire _w2208_ ;
	wire _w2207_ ;
	wire _w2206_ ;
	wire _w2205_ ;
	wire _w2204_ ;
	wire _w2203_ ;
	wire _w2202_ ;
	wire _w2201_ ;
	wire _w2200_ ;
	wire _w2199_ ;
	wire _w2198_ ;
	wire _w2197_ ;
	wire _w2196_ ;
	wire _w2195_ ;
	wire _w2194_ ;
	wire _w2193_ ;
	wire _w2192_ ;
	wire _w2191_ ;
	wire _w2190_ ;
	wire _w2189_ ;
	wire _w2188_ ;
	wire _w2187_ ;
	wire _w2186_ ;
	wire _w2185_ ;
	wire _w2184_ ;
	wire _w2183_ ;
	wire _w2182_ ;
	wire _w2181_ ;
	wire _w2180_ ;
	wire _w2179_ ;
	wire _w2178_ ;
	wire _w2177_ ;
	wire _w2176_ ;
	wire _w2175_ ;
	wire _w2174_ ;
	wire _w2173_ ;
	wire _w2172_ ;
	wire _w2171_ ;
	wire _w2170_ ;
	wire _w2169_ ;
	wire _w2168_ ;
	wire _w2167_ ;
	wire _w2166_ ;
	wire _w2165_ ;
	wire _w2164_ ;
	wire _w2163_ ;
	wire _w2162_ ;
	wire _w2161_ ;
	wire _w2160_ ;
	wire _w2159_ ;
	wire _w2158_ ;
	wire _w2157_ ;
	wire _w2156_ ;
	wire _w2155_ ;
	wire _w2154_ ;
	wire _w2153_ ;
	wire _w2152_ ;
	wire _w2151_ ;
	wire _w2150_ ;
	wire _w2149_ ;
	wire _w2148_ ;
	wire _w2147_ ;
	wire _w2146_ ;
	wire _w2145_ ;
	wire _w2144_ ;
	wire _w2143_ ;
	wire _w2142_ ;
	wire _w2141_ ;
	wire _w2140_ ;
	wire _w2139_ ;
	wire _w2138_ ;
	wire _w2137_ ;
	wire _w2136_ ;
	wire _w2135_ ;
	wire _w2134_ ;
	wire _w2133_ ;
	wire _w2132_ ;
	wire _w2131_ ;
	wire _w2130_ ;
	wire _w2129_ ;
	wire _w2128_ ;
	wire _w2127_ ;
	wire _w2126_ ;
	wire _w2125_ ;
	wire _w2124_ ;
	wire _w2123_ ;
	wire _w2122_ ;
	wire _w2121_ ;
	wire _w2120_ ;
	wire _w2119_ ;
	wire _w2118_ ;
	wire _w2117_ ;
	wire _w2116_ ;
	wire _w2115_ ;
	wire _w2114_ ;
	wire _w2113_ ;
	wire _w2112_ ;
	wire _w2111_ ;
	wire _w2110_ ;
	wire _w2109_ ;
	wire _w2108_ ;
	wire _w2107_ ;
	wire _w2106_ ;
	wire _w2105_ ;
	wire _w2104_ ;
	wire _w2103_ ;
	wire _w2102_ ;
	wire _w2101_ ;
	wire _w2100_ ;
	wire _w2099_ ;
	wire _w2098_ ;
	wire _w2097_ ;
	wire _w2096_ ;
	wire _w2095_ ;
	wire _w2094_ ;
	wire _w2093_ ;
	wire _w2092_ ;
	wire _w2091_ ;
	wire _w2090_ ;
	wire _w2089_ ;
	wire _w2088_ ;
	wire _w2087_ ;
	wire _w2086_ ;
	wire _w2085_ ;
	wire _w2084_ ;
	wire _w2083_ ;
	wire _w2082_ ;
	wire _w2081_ ;
	wire _w2080_ ;
	wire _w2079_ ;
	wire _w2078_ ;
	wire _w2077_ ;
	wire _w2076_ ;
	wire _w2075_ ;
	wire _w2074_ ;
	wire _w2073_ ;
	wire _w2072_ ;
	wire _w2071_ ;
	wire _w2070_ ;
	wire _w2069_ ;
	wire _w2068_ ;
	wire _w2067_ ;
	wire _w2066_ ;
	wire _w2065_ ;
	wire _w2064_ ;
	wire _w2063_ ;
	wire _w2062_ ;
	wire _w2061_ ;
	wire _w2060_ ;
	wire _w2059_ ;
	wire _w2058_ ;
	wire _w2057_ ;
	wire _w2056_ ;
	wire _w2055_ ;
	wire _w2054_ ;
	wire _w2053_ ;
	wire _w2052_ ;
	wire _w2051_ ;
	wire _w2050_ ;
	wire _w2049_ ;
	wire _w2048_ ;
	wire _w2047_ ;
	wire _w2046_ ;
	wire _w2045_ ;
	wire _w2044_ ;
	wire _w2043_ ;
	wire _w2042_ ;
	wire _w2041_ ;
	wire _w2040_ ;
	wire _w2039_ ;
	wire _w2038_ ;
	wire _w2037_ ;
	wire _w2036_ ;
	wire _w2035_ ;
	wire _w2034_ ;
	wire _w2033_ ;
	wire _w2032_ ;
	wire _w2031_ ;
	wire _w2030_ ;
	wire _w2029_ ;
	wire _w2028_ ;
	wire _w2027_ ;
	wire _w2026_ ;
	wire _w2025_ ;
	wire _w2024_ ;
	wire _w2023_ ;
	wire _w2022_ ;
	wire _w2021_ ;
	wire _w2020_ ;
	wire _w2019_ ;
	wire _w2018_ ;
	wire _w2017_ ;
	wire _w2016_ ;
	wire _w2015_ ;
	wire _w2014_ ;
	wire _w2013_ ;
	wire _w2012_ ;
	wire _w2011_ ;
	wire _w2010_ ;
	wire _w2009_ ;
	wire _w2008_ ;
	wire _w2007_ ;
	wire _w2006_ ;
	wire _w2005_ ;
	wire _w2004_ ;
	wire _w2003_ ;
	wire _w2002_ ;
	wire _w2001_ ;
	wire _w2000_ ;
	wire _w1999_ ;
	wire _w1998_ ;
	wire _w1997_ ;
	wire _w1996_ ;
	wire _w1995_ ;
	wire _w1994_ ;
	wire _w1993_ ;
	wire _w1992_ ;
	wire _w1991_ ;
	wire _w1990_ ;
	wire _w1989_ ;
	wire _w1988_ ;
	wire _w1987_ ;
	wire _w1986_ ;
	wire _w1985_ ;
	wire _w1984_ ;
	wire _w1983_ ;
	wire _w1982_ ;
	wire _w1981_ ;
	wire _w1980_ ;
	wire _w1979_ ;
	wire _w1978_ ;
	wire _w1977_ ;
	wire _w1976_ ;
	wire _w1975_ ;
	wire _w1974_ ;
	wire _w1973_ ;
	wire _w1972_ ;
	wire _w1971_ ;
	wire _w1970_ ;
	wire _w1969_ ;
	wire _w1968_ ;
	wire _w1967_ ;
	wire _w1966_ ;
	wire _w1965_ ;
	wire _w1964_ ;
	wire _w1963_ ;
	wire _w1962_ ;
	wire _w1961_ ;
	wire _w1960_ ;
	wire _w1959_ ;
	wire _w1958_ ;
	wire _w1957_ ;
	wire _w1956_ ;
	wire _w1955_ ;
	wire _w1954_ ;
	wire _w1953_ ;
	wire _w1952_ ;
	wire _w1951_ ;
	wire _w1950_ ;
	wire _w1949_ ;
	wire _w1948_ ;
	wire _w1947_ ;
	wire _w1946_ ;
	wire _w1945_ ;
	wire _w1944_ ;
	wire _w1943_ ;
	wire _w1942_ ;
	wire _w1941_ ;
	wire _w1940_ ;
	wire _w1939_ ;
	wire _w1938_ ;
	wire _w1937_ ;
	wire _w1936_ ;
	wire _w1935_ ;
	wire _w1934_ ;
	wire _w1933_ ;
	wire _w1932_ ;
	wire _w1931_ ;
	wire _w1930_ ;
	wire _w1929_ ;
	wire _w1928_ ;
	wire _w1927_ ;
	wire _w1926_ ;
	wire _w1925_ ;
	wire _w1924_ ;
	wire _w1923_ ;
	wire _w1922_ ;
	wire _w1921_ ;
	wire _w1920_ ;
	wire _w1919_ ;
	wire _w1918_ ;
	wire _w1917_ ;
	wire _w1916_ ;
	wire _w1915_ ;
	wire _w1914_ ;
	wire _w1913_ ;
	wire _w1912_ ;
	wire _w1911_ ;
	wire _w1910_ ;
	wire _w1909_ ;
	wire _w1908_ ;
	wire _w1907_ ;
	wire _w1906_ ;
	wire _w1905_ ;
	wire _w1904_ ;
	wire _w1903_ ;
	wire _w1902_ ;
	wire _w1901_ ;
	wire _w1900_ ;
	wire _w1899_ ;
	wire _w1898_ ;
	wire _w1897_ ;
	wire _w1896_ ;
	wire _w1895_ ;
	wire _w1894_ ;
	wire _w1893_ ;
	wire _w1892_ ;
	wire _w1891_ ;
	wire _w1890_ ;
	wire _w1889_ ;
	wire _w1888_ ;
	wire _w1887_ ;
	wire _w1886_ ;
	wire _w1885_ ;
	wire _w1884_ ;
	wire _w1883_ ;
	wire _w1882_ ;
	wire _w1881_ ;
	wire _w1880_ ;
	wire _w1879_ ;
	wire _w1878_ ;
	wire _w1877_ ;
	wire _w1876_ ;
	wire _w1875_ ;
	wire _w1874_ ;
	wire _w1873_ ;
	wire _w1872_ ;
	wire _w1871_ ;
	wire _w1870_ ;
	wire _w1869_ ;
	wire _w1868_ ;
	wire _w1867_ ;
	wire _w1866_ ;
	wire _w1865_ ;
	wire _w1864_ ;
	wire _w1863_ ;
	wire _w1862_ ;
	wire _w1861_ ;
	wire _w1860_ ;
	wire _w1859_ ;
	wire _w1858_ ;
	wire _w1857_ ;
	wire _w1856_ ;
	wire _w1855_ ;
	wire _w1854_ ;
	wire _w1853_ ;
	wire _w1852_ ;
	wire _w1851_ ;
	wire _w1850_ ;
	wire _w1849_ ;
	wire _w1848_ ;
	wire _w1847_ ;
	wire _w1846_ ;
	wire _w1845_ ;
	wire _w1844_ ;
	wire _w1275_ ;
	wire _w1274_ ;
	wire _w1273_ ;
	wire _w1272_ ;
	wire _w1271_ ;
	wire _w1270_ ;
	wire _w1269_ ;
	wire _w1268_ ;
	wire _w1267_ ;
	wire _w1266_ ;
	wire _w1265_ ;
	wire _w1264_ ;
	wire _w1263_ ;
	wire _w1262_ ;
	wire _w1261_ ;
	wire _w1260_ ;
	wire _w1259_ ;
	wire _w1258_ ;
	wire _w1257_ ;
	wire _w1256_ ;
	wire _w1255_ ;
	wire _w1254_ ;
	wire _w1253_ ;
	wire _w1252_ ;
	wire _w1251_ ;
	wire _w1250_ ;
	wire _w1249_ ;
	wire _w1248_ ;
	wire _w1247_ ;
	wire _w1246_ ;
	wire _w1245_ ;
	wire _w1244_ ;
	wire _w1243_ ;
	wire _w1242_ ;
	wire _w1241_ ;
	wire _w1240_ ;
	wire _w1239_ ;
	wire _w1238_ ;
	wire _w1237_ ;
	wire _w1236_ ;
	wire _w1235_ ;
	wire _w1234_ ;
	wire _w1233_ ;
	wire _w1232_ ;
	wire _w1231_ ;
	wire _w1230_ ;
	wire _w1229_ ;
	wire _w1228_ ;
	wire _w1227_ ;
	wire _w1226_ ;
	wire _w1225_ ;
	wire _w1224_ ;
	wire _w1223_ ;
	wire _w1222_ ;
	wire _w1221_ ;
	wire _w1220_ ;
	wire _w1219_ ;
	wire _w1218_ ;
	wire _w1217_ ;
	wire _w1216_ ;
	wire _w1215_ ;
	wire _w1214_ ;
	wire _w1213_ ;
	wire _w1212_ ;
	wire _w1211_ ;
	wire _w1210_ ;
	wire _w1209_ ;
	wire _w1208_ ;
	wire _w1207_ ;
	wire _w1206_ ;
	wire _w1205_ ;
	wire _w1204_ ;
	wire _w1203_ ;
	wire _w1202_ ;
	wire _w1201_ ;
	wire _w1200_ ;
	wire _w1199_ ;
	wire _w1198_ ;
	wire _w1197_ ;
	wire _w1196_ ;
	wire _w1195_ ;
	wire _w1194_ ;
	wire _w1193_ ;
	wire _w1192_ ;
	wire _w1191_ ;
	wire _w1190_ ;
	wire _w1189_ ;
	wire _w1188_ ;
	wire _w1187_ ;
	wire _w1186_ ;
	wire _w1185_ ;
	wire _w1184_ ;
	wire _w1183_ ;
	wire _w1182_ ;
	wire _w1181_ ;
	wire _w1180_ ;
	wire _w1179_ ;
	wire _w1178_ ;
	wire _w1177_ ;
	wire _w1176_ ;
	wire _w1175_ ;
	wire _w1174_ ;
	wire _w1173_ ;
	wire _w1172_ ;
	wire _w1171_ ;
	wire _w1170_ ;
	wire _w1169_ ;
	wire _w1168_ ;
	wire _w1167_ ;
	wire _w1166_ ;
	wire _w1165_ ;
	wire _w1164_ ;
	wire _w1163_ ;
	wire _w1162_ ;
	wire _w1161_ ;
	wire _w1160_ ;
	wire _w1159_ ;
	wire _w1158_ ;
	wire _w1157_ ;
	wire _w1156_ ;
	wire _w1155_ ;
	wire _w1154_ ;
	wire _w1153_ ;
	wire _w1152_ ;
	wire _w1151_ ;
	wire _w1150_ ;
	wire _w1149_ ;
	wire _w1148_ ;
	wire _w1147_ ;
	wire _w1146_ ;
	wire _w1145_ ;
	wire _w1144_ ;
	wire _w1143_ ;
	wire _w1142_ ;
	wire _w1141_ ;
	wire _w1140_ ;
	wire _w1139_ ;
	wire _w1138_ ;
	wire _w1137_ ;
	wire _w1136_ ;
	wire _w1135_ ;
	wire _w1134_ ;
	wire _w1133_ ;
	wire _w1132_ ;
	wire _w1131_ ;
	wire _w1130_ ;
	wire _w1129_ ;
	wire _w1128_ ;
	wire _w1127_ ;
	wire _w1126_ ;
	wire _w1125_ ;
	wire _w1124_ ;
	wire _w1123_ ;
	wire _w1122_ ;
	wire _w1121_ ;
	wire _w1120_ ;
	wire _w1119_ ;
	wire _w1118_ ;
	wire _w1117_ ;
	wire _w1116_ ;
	wire _w1115_ ;
	wire _w1114_ ;
	wire _w1113_ ;
	wire _w1112_ ;
	wire _w1111_ ;
	wire _w1110_ ;
	wire _w1109_ ;
	wire _w1108_ ;
	wire _w1107_ ;
	wire _w1106_ ;
	wire _w1105_ ;
	wire _w1104_ ;
	wire _w1103_ ;
	wire _w1102_ ;
	wire _w1101_ ;
	wire _w1100_ ;
	wire _w1099_ ;
	wire _w1098_ ;
	wire _w1097_ ;
	wire _w1096_ ;
	wire _w1095_ ;
	wire _w1094_ ;
	wire _w1093_ ;
	wire _w1092_ ;
	wire _w1091_ ;
	wire _w1090_ ;
	wire _w1089_ ;
	wire _w1088_ ;
	wire _w1087_ ;
	wire _w1086_ ;
	wire _w1085_ ;
	wire _w1084_ ;
	wire _w1083_ ;
	wire _w1082_ ;
	wire _w1081_ ;
	wire _w1080_ ;
	wire _w1079_ ;
	wire _w1078_ ;
	wire _w1077_ ;
	wire _w1076_ ;
	wire _w1075_ ;
	wire _w1074_ ;
	wire _w1073_ ;
	wire _w1072_ ;
	wire _w1071_ ;
	wire _w1070_ ;
	wire _w1069_ ;
	wire _w1068_ ;
	wire _w1067_ ;
	wire _w1066_ ;
	wire _w1065_ ;
	wire _w1064_ ;
	wire _w1063_ ;
	wire _w1062_ ;
	wire _w1061_ ;
	wire _w1060_ ;
	wire _w1059_ ;
	wire _w1058_ ;
	wire _w1057_ ;
	wire _w1056_ ;
	wire _w1055_ ;
	wire _w1054_ ;
	wire _w1053_ ;
	wire _w1052_ ;
	wire _w1051_ ;
	wire _w1050_ ;
	wire _w1049_ ;
	wire _w1048_ ;
	wire _w1047_ ;
	wire _w1046_ ;
	wire _w1045_ ;
	wire _w1044_ ;
	wire _w1043_ ;
	wire _w1042_ ;
	wire _w1041_ ;
	wire _w1040_ ;
	wire _w1039_ ;
	wire _w1038_ ;
	wire _w1037_ ;
	wire _w1036_ ;
	wire _w1035_ ;
	wire _w1034_ ;
	wire _w1033_ ;
	wire _w1032_ ;
	wire _w1031_ ;
	wire _w1030_ ;
	wire _w1029_ ;
	wire _w1028_ ;
	wire _w1027_ ;
	wire _w1026_ ;
	wire _w1025_ ;
	wire _w1024_ ;
	wire _w1023_ ;
	wire _w1022_ ;
	wire _w1021_ ;
	wire _w1020_ ;
	wire _w1019_ ;
	wire _w1018_ ;
	wire _w1017_ ;
	wire _w1016_ ;
	wire _w1015_ ;
	wire _w1014_ ;
	wire _w1013_ ;
	wire _w1012_ ;
	wire _w1011_ ;
	wire _w1010_ ;
	wire _w1009_ ;
	wire _w1008_ ;
	wire _w1007_ ;
	wire _w1006_ ;
	wire _w1005_ ;
	wire _w1004_ ;
	wire _w1003_ ;
	wire _w1002_ ;
	wire _w1001_ ;
	wire _w1000_ ;
	wire _w999_ ;
	wire _w998_ ;
	wire _w997_ ;
	wire _w996_ ;
	wire _w995_ ;
	wire _w994_ ;
	wire _w993_ ;
	wire _w992_ ;
	wire _w861_ ;
	wire _w860_ ;
	wire _w859_ ;
	wire _w858_ ;
	wire _w857_ ;
	wire _w856_ ;
	wire _w855_ ;
	wire _w854_ ;
	wire _w853_ ;
	wire _w852_ ;
	wire _w851_ ;
	wire _w850_ ;
	wire _w849_ ;
	wire _w848_ ;
	wire _w846_ ;
	wire _w845_ ;
	wire _w844_ ;
	wire _w843_ ;
	wire _w842_ ;
	wire _w841_ ;
	wire _w840_ ;
	wire _w839_ ;
	wire _w838_ ;
	wire _w837_ ;
	wire _w836_ ;
	wire _w835_ ;
	wire _w834_ ;
	wire _w833_ ;
	wire _w832_ ;
	wire _w831_ ;
	wire _w830_ ;
	wire _w829_ ;
	wire _w828_ ;
	wire _w827_ ;
	wire _w826_ ;
	wire _w825_ ;
	wire _w824_ ;
	wire _w823_ ;
	wire _w822_ ;
	wire _w821_ ;
	wire _w820_ ;
	wire _w819_ ;
	wire _w818_ ;
	wire _w817_ ;
	wire _w816_ ;
	wire _w815_ ;
	wire _w814_ ;
	wire _w813_ ;
	wire _w812_ ;
	wire _w811_ ;
	wire _w810_ ;
	wire _w809_ ;
	wire _w808_ ;
	wire _w807_ ;
	wire _w806_ ;
	wire _w805_ ;
	wire _w804_ ;
	wire _w803_ ;
	wire _w802_ ;
	wire _w801_ ;
	wire _w800_ ;
	wire _w799_ ;
	wire _w798_ ;
	wire _w797_ ;
	wire _w796_ ;
	wire _w795_ ;
	wire _w794_ ;
	wire _w762_ ;
	wire _w761_ ;
	wire _w760_ ;
	wire _w759_ ;
	wire _w758_ ;
	wire _w757_ ;
	wire _w756_ ;
	wire _w755_ ;
	wire _w754_ ;
	wire _w752_ ;
	wire _w750_ ;
	wire _w749_ ;
	wire _w748_ ;
	wire _w763_ ;
	wire _w847_ ;
	wire _w753_ ;
	wire _w2569_ ;
	wire _w212_ ;
	wire _w1321_ ;
	wire _w983_ ;
	wire _w743_ ;
	wire _w745_ ;
	wire _w751_ ;
	wire _w774_ ;
	wire _w737_ ;
	wire _w738_ ;
	wire _w739_ ;
	wire _w740_ ;
	wire _w741_ ;
	wire _w742_ ;
	wire _w744_ ;
	wire _w746_ ;
	wire _w747_ ;
	wire _w764_ ;
	wire _w765_ ;
	wire _w766_ ;
	wire _w767_ ;
	wire _w768_ ;
	wire _w769_ ;
	wire _w770_ ;
	wire _w771_ ;
	wire _w772_ ;
	wire _w773_ ;
	wire _w775_ ;
	wire _w776_ ;
	wire _w777_ ;
	wire _w778_ ;
	wire _w779_ ;
	wire _w780_ ;
	wire _w781_ ;
	wire _w782_ ;
	wire _w783_ ;
	wire _w2600_ ;
	wire _w243_ ;
	wire _w1352_ ;
	wire _w784_ ;
	wire _w785_ ;
	wire _w786_ ;
	wire _w787_ ;
	wire _w788_ ;
	wire _w789_ ;
	wire _w790_ ;
	wire _w791_ ;
	wire _w792_ ;
	wire _w793_ ;
	wire _w862_ ;
	wire _w863_ ;
	wire _w864_ ;
	wire _w865_ ;
	wire _w866_ ;
	wire _w867_ ;
	wire _w868_ ;
	wire _w869_ ;
	wire _w870_ ;
	wire _w871_ ;
	wire _w872_ ;
	wire _w873_ ;
	wire _w874_ ;
	wire _w875_ ;
	wire _w876_ ;
	wire _w877_ ;
	wire _w878_ ;
	wire _w879_ ;
	wire _w880_ ;
	wire _w881_ ;
	wire _w882_ ;
	wire _w883_ ;
	wire _w884_ ;
	wire _w885_ ;
	wire _w886_ ;
	wire _w887_ ;
	wire _w888_ ;
	wire _w889_ ;
	wire _w890_ ;
	wire _w891_ ;
	wire _w892_ ;
	wire _w893_ ;
	wire _w894_ ;
	wire _w895_ ;
	wire _w896_ ;
	wire _w897_ ;
	wire _w898_ ;
	wire _w899_ ;
	wire _w900_ ;
	wire _w901_ ;
	wire _w902_ ;
	wire _w903_ ;
	wire _w904_ ;
	wire _w905_ ;
	wire _w906_ ;
	wire _w907_ ;
	wire _w908_ ;
	wire _w909_ ;
	wire _w910_ ;
	wire _w911_ ;
	wire _w912_ ;
	wire _w913_ ;
	wire _w914_ ;
	wire _w915_ ;
	wire _w916_ ;
	wire _w917_ ;
	wire _w918_ ;
	wire _w919_ ;
	wire _w920_ ;
	wire _w921_ ;
	wire _w922_ ;
	wire _w923_ ;
	wire _w924_ ;
	wire _w925_ ;
	wire _w926_ ;
	wire _w927_ ;
	wire _w928_ ;
	wire _w929_ ;
	wire _w930_ ;
	wire _w931_ ;
	wire _w932_ ;
	wire _w933_ ;
	wire _w934_ ;
	wire _w935_ ;
	wire _w936_ ;
	wire _w937_ ;
	wire _w938_ ;
	wire _w939_ ;
	wire _w940_ ;
	wire _w941_ ;
	wire _w942_ ;
	wire _w943_ ;
	wire _w944_ ;
	wire _w945_ ;
	wire _w946_ ;
	wire _w947_ ;
	wire _w948_ ;
	wire _w949_ ;
	wire _w950_ ;
	wire _w951_ ;
	wire _w952_ ;
	wire _w953_ ;
	wire _w954_ ;
	wire _w955_ ;
	wire _w956_ ;
	wire _w957_ ;
	wire _w958_ ;
	wire _w959_ ;
	wire _w960_ ;
	wire _w961_ ;
	wire _w962_ ;
	wire _w963_ ;
	wire _w964_ ;
	wire _w965_ ;
	wire _w966_ ;
	wire _w967_ ;
	wire _w968_ ;
	wire _w969_ ;
	wire _w970_ ;
	wire _w971_ ;
	wire _w972_ ;
	wire _w973_ ;
	wire _w974_ ;
	wire _w975_ ;
	wire _w976_ ;
	wire _w977_ ;
	wire _w978_ ;
	wire _w979_ ;
	wire _w980_ ;
	wire _w981_ ;
	wire _w982_ ;
	wire _w984_ ;
	wire _w985_ ;
	wire _w986_ ;
	wire _w987_ ;
	wire _w988_ ;
	wire _w989_ ;
	wire _w990_ ;
	wire _w991_ ;
	wire _w1276_ ;
	wire _w1277_ ;
	wire _w1278_ ;
	wire _w1279_ ;
	wire _w1280_ ;
	wire _w1281_ ;
	wire _w1282_ ;
	wire _w1283_ ;
	wire _w1284_ ;
	wire _w1285_ ;
	wire _w1286_ ;
	wire _w1287_ ;
	wire _w1288_ ;
	wire _w1289_ ;
	wire _w1290_ ;
	wire _w1291_ ;
	wire _w1292_ ;
	wire _w1293_ ;
	wire _w1294_ ;
	wire _w1295_ ;
	wire _w1296_ ;
	wire _w1297_ ;
	wire _w1298_ ;
	wire _w1299_ ;
	wire _w1300_ ;
	wire _w1301_ ;
	wire _w1302_ ;
	wire _w1303_ ;
	wire _w1304_ ;
	wire _w1305_ ;
	wire _w1306_ ;
	wire _w1307_ ;
	wire _w1308_ ;
	wire _w1309_ ;
	wire _w1310_ ;
	wire _w1311_ ;
	wire _w1312_ ;
	wire _w1313_ ;
	wire _w1314_ ;
	wire _w1315_ ;
	wire _w1316_ ;
	wire _w1317_ ;
	wire _w1318_ ;
	wire _w1319_ ;
	wire _w1320_ ;
	wire _w1322_ ;
	wire _w1323_ ;
	wire _w1324_ ;
	wire _w1325_ ;
	wire _w1326_ ;
	wire _w1327_ ;
	wire _w1328_ ;
	wire _w1329_ ;
	wire _w1330_ ;
	wire _w1331_ ;
	wire _w1332_ ;
	wire _w1333_ ;
	wire _w1334_ ;
	wire _w1335_ ;
	wire _w1336_ ;
	wire _w1337_ ;
	wire _w1338_ ;
	wire _w1339_ ;
	wire _w1340_ ;
	wire _w1341_ ;
	wire _w1342_ ;
	wire _w1343_ ;
	wire _w1344_ ;
	wire _w1345_ ;
	wire _w1346_ ;
	wire _w1347_ ;
	wire _w1348_ ;
	wire _w1349_ ;
	wire _w1350_ ;
	wire _w1351_ ;
	wire _w1353_ ;
	wire _w1354_ ;
	wire _w1355_ ;
	wire _w1356_ ;
	wire _w1357_ ;
	wire _w1358_ ;
	wire _w1359_ ;
	wire _w1360_ ;
	wire _w1361_ ;
	wire _w1362_ ;
	wire _w1363_ ;
	wire _w1364_ ;
	wire _w1365_ ;
	wire _w1366_ ;
	wire _w1367_ ;
	wire _w1368_ ;
	wire _w1369_ ;
	wire _w1370_ ;
	wire _w1371_ ;
	wire _w1372_ ;
	wire _w1373_ ;
	wire _w1374_ ;
	wire _w1375_ ;
	wire _w1376_ ;
	wire _w1377_ ;
	wire _w1378_ ;
	wire _w1379_ ;
	wire _w1380_ ;
	wire _w1381_ ;
	wire _w1382_ ;
	wire _w1383_ ;
	wire _w1384_ ;
	wire _w1385_ ;
	wire _w1386_ ;
	wire _w1387_ ;
	wire _w1388_ ;
	wire _w1389_ ;
	wire _w1390_ ;
	wire _w1391_ ;
	wire _w1392_ ;
	wire _w1393_ ;
	wire _w1394_ ;
	wire _w1395_ ;
	wire _w1396_ ;
	wire _w1397_ ;
	wire _w1398_ ;
	wire _w1399_ ;
	wire _w1400_ ;
	wire _w1401_ ;
	wire _w1402_ ;
	wire _w1403_ ;
	wire _w1404_ ;
	wire _w1405_ ;
	wire _w1406_ ;
	wire _w1407_ ;
	wire _w1408_ ;
	wire _w1409_ ;
	wire _w1410_ ;
	wire _w1411_ ;
	wire _w1412_ ;
	wire _w1413_ ;
	wire _w1414_ ;
	wire _w1415_ ;
	wire _w1416_ ;
	wire _w1417_ ;
	wire _w1418_ ;
	wire _w1419_ ;
	wire _w1420_ ;
	wire _w1421_ ;
	wire _w1422_ ;
	wire _w1423_ ;
	wire _w1424_ ;
	wire _w1425_ ;
	wire _w1426_ ;
	wire _w1427_ ;
	wire _w1428_ ;
	wire _w1429_ ;
	wire _w1430_ ;
	wire _w1431_ ;
	wire _w1432_ ;
	wire _w1433_ ;
	wire _w1434_ ;
	wire _w1435_ ;
	wire _w1436_ ;
	wire _w1437_ ;
	wire _w1438_ ;
	wire _w1439_ ;
	wire _w1440_ ;
	wire _w1441_ ;
	wire _w1442_ ;
	wire _w1443_ ;
	wire _w1444_ ;
	wire _w1445_ ;
	wire _w1446_ ;
	wire _w1447_ ;
	wire _w1448_ ;
	wire _w1449_ ;
	wire _w1450_ ;
	wire _w1451_ ;
	wire _w1452_ ;
	wire _w1453_ ;
	wire _w1454_ ;
	wire _w1455_ ;
	wire _w1456_ ;
	wire _w1457_ ;
	wire _w1458_ ;
	wire _w1459_ ;
	wire _w1460_ ;
	wire _w1461_ ;
	wire _w1462_ ;
	wire _w1463_ ;
	wire _w1464_ ;
	wire _w1465_ ;
	wire _w1466_ ;
	wire _w1467_ ;
	wire _w1468_ ;
	wire _w1469_ ;
	wire _w1470_ ;
	wire _w1471_ ;
	wire _w1472_ ;
	wire _w1473_ ;
	wire _w1474_ ;
	wire _w1475_ ;
	wire _w1476_ ;
	wire _w1477_ ;
	wire _w1478_ ;
	wire _w1479_ ;
	wire _w1480_ ;
	wire _w1481_ ;
	wire _w1482_ ;
	wire _w1483_ ;
	wire _w1484_ ;
	wire _w1485_ ;
	wire _w1486_ ;
	wire _w1487_ ;
	wire _w1488_ ;
	wire _w1489_ ;
	wire _w1490_ ;
	wire _w1491_ ;
	wire _w1492_ ;
	wire _w1493_ ;
	wire _w1494_ ;
	wire _w1495_ ;
	wire _w1496_ ;
	wire _w1497_ ;
	wire _w1498_ ;
	wire _w1499_ ;
	wire _w1500_ ;
	wire _w1501_ ;
	wire _w1502_ ;
	wire _w1503_ ;
	wire _w1504_ ;
	wire _w1505_ ;
	wire _w1506_ ;
	wire _w1507_ ;
	wire _w1508_ ;
	wire _w1509_ ;
	wire _w1510_ ;
	wire _w1511_ ;
	wire _w1512_ ;
	wire _w1513_ ;
	wire _w1514_ ;
	wire _w1515_ ;
	wire _w1516_ ;
	wire _w1517_ ;
	wire _w1518_ ;
	wire _w1519_ ;
	wire _w1520_ ;
	wire _w1521_ ;
	wire _w1522_ ;
	wire _w1523_ ;
	wire _w1524_ ;
	wire _w1525_ ;
	wire _w1526_ ;
	wire _w1527_ ;
	wire _w1528_ ;
	wire _w1529_ ;
	wire _w1530_ ;
	wire _w1531_ ;
	wire _w1532_ ;
	wire _w1533_ ;
	wire _w1534_ ;
	wire _w1535_ ;
	wire _w1536_ ;
	wire _w1537_ ;
	wire _w1538_ ;
	wire _w1539_ ;
	wire _w1540_ ;
	wire _w1541_ ;
	wire _w1542_ ;
	wire _w1543_ ;
	wire _w1544_ ;
	wire _w1545_ ;
	wire _w1546_ ;
	wire _w1547_ ;
	wire _w1548_ ;
	wire _w1549_ ;
	wire _w1550_ ;
	wire _w1551_ ;
	wire _w1552_ ;
	wire _w1553_ ;
	wire _w1554_ ;
	wire _w1555_ ;
	wire _w1556_ ;
	wire _w1557_ ;
	wire _w1558_ ;
	wire _w1559_ ;
	wire _w1560_ ;
	wire _w1561_ ;
	wire _w1562_ ;
	wire _w1563_ ;
	wire _w1564_ ;
	wire _w1565_ ;
	wire _w1566_ ;
	wire _w1567_ ;
	wire _w1568_ ;
	wire _w1569_ ;
	wire _w1570_ ;
	wire _w1571_ ;
	wire _w1572_ ;
	wire _w1573_ ;
	wire _w1574_ ;
	wire _w1575_ ;
	wire _w1576_ ;
	wire _w1577_ ;
	wire _w1578_ ;
	wire _w1579_ ;
	wire _w1580_ ;
	wire _w1581_ ;
	wire _w1582_ ;
	wire _w1583_ ;
	wire _w1584_ ;
	wire _w1585_ ;
	wire _w1586_ ;
	wire _w1587_ ;
	wire _w1588_ ;
	wire _w1589_ ;
	wire _w1590_ ;
	wire _w1591_ ;
	wire _w1592_ ;
	wire _w1593_ ;
	wire _w1594_ ;
	wire _w1595_ ;
	wire _w1596_ ;
	wire _w1597_ ;
	wire _w1598_ ;
	wire _w1599_ ;
	wire _w1600_ ;
	wire _w1601_ ;
	wire _w1602_ ;
	wire _w1603_ ;
	wire _w1604_ ;
	wire _w1605_ ;
	wire _w1606_ ;
	wire _w1607_ ;
	wire _w1608_ ;
	wire _w1609_ ;
	wire _w1610_ ;
	wire _w1611_ ;
	wire _w1612_ ;
	wire _w1613_ ;
	wire _w1614_ ;
	wire _w1615_ ;
	wire _w1616_ ;
	wire _w1617_ ;
	wire _w1618_ ;
	wire _w1619_ ;
	wire _w1620_ ;
	wire _w1621_ ;
	wire _w1622_ ;
	wire _w1623_ ;
	wire _w1624_ ;
	wire _w1625_ ;
	wire _w1626_ ;
	wire _w1627_ ;
	wire _w1628_ ;
	wire _w1629_ ;
	wire _w1630_ ;
	wire _w1631_ ;
	wire _w1632_ ;
	wire _w1633_ ;
	wire _w1634_ ;
	wire _w1635_ ;
	wire _w1636_ ;
	wire _w1637_ ;
	wire _w1638_ ;
	wire _w1639_ ;
	wire _w1640_ ;
	wire _w1641_ ;
	wire _w1642_ ;
	wire _w1643_ ;
	wire _w1644_ ;
	wire _w1645_ ;
	wire _w1646_ ;
	wire _w1647_ ;
	wire _w1648_ ;
	wire _w1649_ ;
	wire _w1650_ ;
	wire _w1651_ ;
	wire _w1652_ ;
	wire _w1653_ ;
	wire _w1654_ ;
	wire _w1655_ ;
	wire _w1656_ ;
	wire _w1657_ ;
	wire _w1658_ ;
	wire _w1659_ ;
	wire _w1660_ ;
	wire _w1661_ ;
	wire _w1662_ ;
	wire _w1663_ ;
	wire _w1664_ ;
	wire _w1665_ ;
	wire _w1666_ ;
	wire _w1667_ ;
	wire _w1668_ ;
	wire _w1669_ ;
	wire _w1670_ ;
	wire _w1671_ ;
	wire _w1672_ ;
	wire _w1673_ ;
	wire _w1674_ ;
	wire _w1675_ ;
	wire _w1676_ ;
	wire _w1677_ ;
	wire _w1678_ ;
	wire _w1679_ ;
	wire _w1680_ ;
	wire _w1681_ ;
	wire _w1682_ ;
	wire _w1683_ ;
	wire _w1684_ ;
	wire _w1685_ ;
	wire _w1686_ ;
	wire _w1687_ ;
	wire _w1688_ ;
	wire _w1689_ ;
	wire _w1690_ ;
	wire _w1691_ ;
	wire _w1692_ ;
	wire _w1693_ ;
	wire _w1694_ ;
	wire _w1695_ ;
	wire _w1696_ ;
	wire _w1697_ ;
	wire _w1698_ ;
	wire _w1699_ ;
	wire _w1700_ ;
	wire _w1701_ ;
	wire _w1702_ ;
	wire _w1703_ ;
	wire _w1704_ ;
	wire _w1705_ ;
	wire _w1706_ ;
	wire _w1707_ ;
	wire _w1708_ ;
	wire _w1709_ ;
	wire _w1710_ ;
	wire _w1711_ ;
	wire _w1712_ ;
	wire _w1713_ ;
	wire _w1714_ ;
	wire _w1715_ ;
	wire _w1716_ ;
	wire _w1717_ ;
	wire _w1718_ ;
	wire _w1719_ ;
	wire _w1720_ ;
	wire _w1721_ ;
	wire _w1722_ ;
	wire _w1723_ ;
	wire _w1724_ ;
	wire _w1725_ ;
	wire _w1726_ ;
	wire _w1727_ ;
	wire _w1728_ ;
	wire _w1729_ ;
	wire _w1730_ ;
	wire _w1731_ ;
	wire _w1732_ ;
	wire _w1733_ ;
	wire _w1734_ ;
	wire _w1735_ ;
	wire _w1736_ ;
	wire _w1737_ ;
	wire _w1738_ ;
	wire _w1739_ ;
	wire _w1740_ ;
	wire _w1741_ ;
	wire _w1742_ ;
	wire _w1743_ ;
	wire _w1744_ ;
	wire _w1745_ ;
	wire _w1746_ ;
	wire _w1747_ ;
	wire _w1748_ ;
	wire _w1749_ ;
	wire _w1750_ ;
	wire _w1751_ ;
	wire _w1752_ ;
	wire _w1753_ ;
	wire _w1754_ ;
	wire _w1755_ ;
	wire _w1756_ ;
	wire _w1757_ ;
	wire _w1758_ ;
	wire _w1759_ ;
	wire _w1760_ ;
	wire _w1761_ ;
	wire _w1762_ ;
	wire _w1763_ ;
	wire _w1764_ ;
	wire _w1765_ ;
	wire _w1766_ ;
	wire _w1767_ ;
	wire _w1768_ ;
	wire _w1769_ ;
	wire _w1770_ ;
	wire _w1771_ ;
	wire _w1772_ ;
	wire _w1773_ ;
	wire _w1774_ ;
	wire _w1775_ ;
	wire _w1776_ ;
	wire _w1777_ ;
	wire _w1778_ ;
	wire _w1779_ ;
	wire _w1780_ ;
	wire _w1781_ ;
	wire _w1782_ ;
	wire _w1783_ ;
	wire _w1784_ ;
	wire _w1785_ ;
	wire _w1786_ ;
	wire _w1787_ ;
	wire _w1788_ ;
	wire _w1789_ ;
	wire _w1790_ ;
	wire _w1791_ ;
	wire _w1792_ ;
	wire _w1793_ ;
	wire _w1794_ ;
	wire _w1795_ ;
	wire _w1796_ ;
	wire _w1797_ ;
	wire _w1798_ ;
	wire _w1799_ ;
	wire _w1800_ ;
	wire _w1801_ ;
	wire _w1802_ ;
	wire _w1803_ ;
	wire _w1804_ ;
	wire _w1805_ ;
	wire _w1806_ ;
	wire _w1807_ ;
	wire _w1808_ ;
	wire _w1809_ ;
	wire _w1810_ ;
	wire _w1811_ ;
	wire _w1812_ ;
	wire _w1813_ ;
	wire _w1814_ ;
	wire _w1815_ ;
	wire _w1816_ ;
	wire _w1817_ ;
	wire _w1818_ ;
	wire _w1819_ ;
	wire _w1820_ ;
	wire _w1821_ ;
	wire _w1822_ ;
	wire _w1823_ ;
	wire _w1824_ ;
	wire _w1825_ ;
	wire _w1826_ ;
	wire _w1827_ ;
	wire _w1828_ ;
	wire _w1829_ ;
	wire _w1830_ ;
	wire _w1831_ ;
	wire _w1832_ ;
	wire _w1833_ ;
	wire _w1834_ ;
	wire _w1835_ ;
	wire _w1836_ ;
	wire _w1837_ ;
	wire _w1838_ ;
	wire _w1839_ ;
	wire _w1840_ ;
	wire _w1841_ ;
	wire _w1842_ ;
	wire _w1843_ ;
	LUT1 #(
		.INIT('h1)
	) name0 (
		\u2_adr0_cnt_reg[0]/P0001 ,
		_w212_
	);
	LUT1 #(
		.INIT('h1)
	) name1 (
		\u2_adr1_cnt_reg[0]/P0001 ,
		_w243_
	);
	LUT3 #(
		.INIT('h1b)
	) name2 (
		\u0_u0_ch_csr_r_reg[1]/NET0131 ,
		\wb0_ack_i_pad ,
		\wb1_ack_i_pad ,
		_w737_
	);
	LUT2 #(
		.INIT('h8)
	) name3 (
		\u0_u0_ch_csr_r_reg[3]/NET0131 ,
		\u2_write_r_reg/P0001 ,
		_w738_
	);
	LUT2 #(
		.INIT('h8)
	) name4 (
		\u2_adr1_cnt_reg[16]/NET0131 ,
		\u2_u1_out_r_reg[16]/P0001 ,
		_w739_
	);
	LUT3 #(
		.INIT('h80)
	) name5 (
		\u2_adr1_cnt_reg[16]/NET0131 ,
		\u2_adr1_cnt_reg[17]/P0001 ,
		\u2_u1_out_r_reg[16]/P0001 ,
		_w740_
	);
	LUT3 #(
		.INIT('h80)
	) name6 (
		\u2_adr1_cnt_reg[18]/P0001 ,
		\u2_adr1_cnt_reg[19]/P0001 ,
		\u2_adr1_cnt_reg[20]/P0001 ,
		_w741_
	);
	LUT4 #(
		.INIT('h4000)
	) name7 (
		_w737_,
		_w738_,
		_w740_,
		_w741_,
		_w742_
	);
	LUT3 #(
		.INIT('h80)
	) name8 (
		\u2_adr1_cnt_reg[23]/P0001 ,
		\u2_adr1_cnt_reg[24]/P0001 ,
		\u2_adr1_cnt_reg[25]/P0001 ,
		_w743_
	);
	LUT2 #(
		.INIT('h8)
	) name9 (
		\u2_adr1_cnt_reg[21]/P0001 ,
		\u2_adr1_cnt_reg[22]/P0001 ,
		_w744_
	);
	LUT3 #(
		.INIT('h80)
	) name10 (
		\u2_adr1_cnt_reg[21]/P0001 ,
		\u2_adr1_cnt_reg[22]/P0001 ,
		\u2_adr1_cnt_reg[26]/P0001 ,
		_w745_
	);
	LUT2 #(
		.INIT('h8)
	) name11 (
		_w743_,
		_w745_,
		_w746_
	);
	LUT3 #(
		.INIT('h8c)
	) name12 (
		dma_ack_o_pad,
		\u0_u0_ch_csr_r_reg[5]/NET0131 ,
		\u1_req_r_reg[0]/P0001 ,
		_w747_
	);
	LUT2 #(
		.INIT('h2)
	) name13 (
		\u0_u0_ch_csr_r_reg[0]/NET0131 ,
		\u1_de_start_r_reg/P0001 ,
		_w748_
	);
	LUT2 #(
		.INIT('h1)
	) name14 (
		\u1_next_start_reg/P0001 ,
		\u2_state_reg[8]/NET0131 ,
		_w749_
	);
	LUT3 #(
		.INIT('hb0)
	) name15 (
		_w747_,
		_w748_,
		_w749_,
		_w750_
	);
	LUT4 #(
		.INIT('h8a00)
	) name16 (
		\u2_adr1_cnt_reg[28]/P0001 ,
		_w747_,
		_w748_,
		_w749_,
		_w751_
	);
	LUT4 #(
		.INIT('h7f00)
	) name17 (
		\u2_adr1_cnt_reg[27]/P0001 ,
		_w742_,
		_w746_,
		_w751_,
		_w752_
	);
	LUT4 #(
		.INIT('h4500)
	) name18 (
		\u2_adr1_cnt_reg[28]/P0001 ,
		_w747_,
		_w748_,
		_w749_,
		_w753_
	);
	LUT4 #(
		.INIT('h8000)
	) name19 (
		\u2_adr1_cnt_reg[27]/P0001 ,
		_w742_,
		_w746_,
		_w753_,
		_w754_
	);
	LUT4 #(
		.INIT('h20aa)
	) name20 (
		\u0_u0_ch_adr1_r_reg[28]/P0001 ,
		_w747_,
		_w748_,
		_w749_,
		_w755_
	);
	LUT3 #(
		.INIT('hfe)
	) name21 (
		_w752_,
		_w754_,
		_w755_,
		_w756_
	);
	LUT3 #(
		.INIT('h1b)
	) name22 (
		\u0_u0_ch_csr_r_reg[2]/NET0131 ,
		\wb0_ack_i_pad ,
		\wb1_ack_i_pad ,
		_w757_
	);
	LUT2 #(
		.INIT('h8)
	) name23 (
		\u0_u0_ch_csr_r_reg[4]/NET0131 ,
		\u2_read_r_reg/P0001 ,
		_w758_
	);
	LUT3 #(
		.INIT('h80)
	) name24 (
		\u0_u0_ch_csr_r_reg[4]/NET0131 ,
		\u2_read_r_reg/P0001 ,
		\u2_u0_out_r_reg[16]/P0001 ,
		_w759_
	);
	LUT4 #(
		.INIT('h8000)
	) name25 (
		\u2_adr0_cnt_reg[16]/NET0131 ,
		\u2_adr0_cnt_reg[17]/P0001 ,
		\u2_adr0_cnt_reg[18]/P0001 ,
		\u2_adr0_cnt_reg[19]/P0001 ,
		_w760_
	);
	LUT4 #(
		.INIT('h2000)
	) name26 (
		\u2_adr0_cnt_reg[20]/P0001 ,
		_w757_,
		_w759_,
		_w760_,
		_w761_
	);
	LUT3 #(
		.INIT('h80)
	) name27 (
		\u2_adr0_cnt_reg[21]/P0001 ,
		\u2_adr0_cnt_reg[22]/P0001 ,
		\u2_adr0_cnt_reg[23]/P0001 ,
		_w762_
	);
	LUT2 #(
		.INIT('h8)
	) name28 (
		\u2_adr0_cnt_reg[24]/P0001 ,
		\u2_adr0_cnt_reg[25]/P0001 ,
		_w763_
	);
	LUT4 #(
		.INIT('h8000)
	) name29 (
		\u2_adr0_cnt_reg[24]/P0001 ,
		\u2_adr0_cnt_reg[25]/P0001 ,
		\u2_adr0_cnt_reg[26]/P0001 ,
		\u2_adr0_cnt_reg[27]/P0001 ,
		_w764_
	);
	LUT2 #(
		.INIT('h8)
	) name30 (
		_w762_,
		_w764_,
		_w765_
	);
	LUT4 #(
		.INIT('hb777)
	) name31 (
		\u2_adr0_cnt_reg[28]/P0001 ,
		_w750_,
		_w761_,
		_w765_,
		_w766_
	);
	LUT4 #(
		.INIT('h20aa)
	) name32 (
		\u0_u0_ch_adr0_r_reg[28]/P0001 ,
		_w747_,
		_w748_,
		_w749_,
		_w767_
	);
	LUT2 #(
		.INIT('hd)
	) name33 (
		_w766_,
		_w767_,
		_w768_
	);
	LUT4 #(
		.INIT('h95ff)
	) name34 (
		\u2_adr1_cnt_reg[27]/P0001 ,
		_w742_,
		_w746_,
		_w750_,
		_w769_
	);
	LUT4 #(
		.INIT('h20aa)
	) name35 (
		\u0_u0_ch_adr1_r_reg[27]/P0001 ,
		_w747_,
		_w748_,
		_w749_,
		_w770_
	);
	LUT2 #(
		.INIT('hd)
	) name36 (
		_w769_,
		_w770_,
		_w771_
	);
	LUT4 #(
		.INIT('h20aa)
	) name37 (
		\u0_u0_ch_adr0_r_reg[27]/P0001 ,
		_w747_,
		_w748_,
		_w749_,
		_w772_
	);
	LUT3 #(
		.INIT('h80)
	) name38 (
		\u2_adr0_cnt_reg[24]/P0001 ,
		\u2_adr0_cnt_reg[25]/P0001 ,
		\u2_adr0_cnt_reg[26]/P0001 ,
		_w773_
	);
	LUT2 #(
		.INIT('h8)
	) name39 (
		_w762_,
		_w773_,
		_w774_
	);
	LUT3 #(
		.INIT('h15)
	) name40 (
		\u2_adr0_cnt_reg[27]/P0001 ,
		_w761_,
		_w774_,
		_w775_
	);
	LUT3 #(
		.INIT('h2a)
	) name41 (
		_w750_,
		_w761_,
		_w765_,
		_w776_
	);
	LUT3 #(
		.INIT('hba)
	) name42 (
		_w772_,
		_w775_,
		_w776_,
		_w777_
	);
	LUT2 #(
		.INIT('h8)
	) name43 (
		_w743_,
		_w744_,
		_w778_
	);
	LUT3 #(
		.INIT('h15)
	) name44 (
		\u2_adr1_cnt_reg[26]/P0001 ,
		_w742_,
		_w778_,
		_w779_
	);
	LUT3 #(
		.INIT('h70)
	) name45 (
		_w742_,
		_w746_,
		_w750_,
		_w780_
	);
	LUT4 #(
		.INIT('h20aa)
	) name46 (
		\u0_u0_ch_adr1_r_reg[26]/P0001 ,
		_w747_,
		_w748_,
		_w749_,
		_w781_
	);
	LUT3 #(
		.INIT('hf4)
	) name47 (
		_w779_,
		_w780_,
		_w781_,
		_w782_
	);
	LUT2 #(
		.INIT('h8)
	) name48 (
		_w762_,
		_w763_,
		_w783_
	);
	LUT3 #(
		.INIT('h15)
	) name49 (
		\u2_adr0_cnt_reg[26]/P0001 ,
		_w761_,
		_w783_,
		_w784_
	);
	LUT3 #(
		.INIT('h2a)
	) name50 (
		_w750_,
		_w761_,
		_w774_,
		_w785_
	);
	LUT4 #(
		.INIT('h20aa)
	) name51 (
		\u0_u0_ch_adr0_r_reg[26]/P0001 ,
		_w747_,
		_w748_,
		_w749_,
		_w786_
	);
	LUT3 #(
		.INIT('hf4)
	) name52 (
		_w784_,
		_w785_,
		_w786_,
		_w787_
	);
	LUT4 #(
		.INIT('h8000)
	) name53 (
		\u2_adr0_cnt_reg[21]/P0001 ,
		\u2_adr0_cnt_reg[22]/P0001 ,
		\u2_adr0_cnt_reg[23]/P0001 ,
		\u2_adr0_cnt_reg[24]/P0001 ,
		_w788_
	);
	LUT4 #(
		.INIT('h4888)
	) name54 (
		\u2_adr0_cnt_reg[24]/P0001 ,
		_w750_,
		_w761_,
		_w762_,
		_w789_
	);
	LUT4 #(
		.INIT('h20aa)
	) name55 (
		\u0_u0_ch_adr0_r_reg[24]/P0001 ,
		_w747_,
		_w748_,
		_w749_,
		_w790_
	);
	LUT2 #(
		.INIT('he)
	) name56 (
		_w789_,
		_w790_,
		_w791_
	);
	LUT3 #(
		.INIT('h80)
	) name57 (
		\u2_adr1_cnt_reg[21]/P0001 ,
		\u2_adr1_cnt_reg[22]/P0001 ,
		\u2_adr1_cnt_reg[23]/P0001 ,
		_w792_
	);
	LUT3 #(
		.INIT('h15)
	) name58 (
		\u2_adr1_cnt_reg[24]/P0001 ,
		_w742_,
		_w792_,
		_w793_
	);
	LUT4 #(
		.INIT('h8000)
	) name59 (
		\u2_adr1_cnt_reg[21]/P0001 ,
		\u2_adr1_cnt_reg[22]/P0001 ,
		\u2_adr1_cnt_reg[23]/P0001 ,
		\u2_adr1_cnt_reg[24]/P0001 ,
		_w794_
	);
	LUT3 #(
		.INIT('h4c)
	) name60 (
		_w742_,
		_w750_,
		_w794_,
		_w795_
	);
	LUT4 #(
		.INIT('h20aa)
	) name61 (
		\u0_u0_ch_adr1_r_reg[24]/P0001 ,
		_w747_,
		_w748_,
		_w749_,
		_w796_
	);
	LUT3 #(
		.INIT('hf4)
	) name62 (
		_w793_,
		_w795_,
		_w796_,
		_w797_
	);
	LUT4 #(
		.INIT('h20aa)
	) name63 (
		\u0_u0_ch_adr0_r_reg[23]/P0001 ,
		_w747_,
		_w748_,
		_w749_,
		_w798_
	);
	LUT2 #(
		.INIT('h8)
	) name64 (
		\u2_adr0_cnt_reg[20]/P0001 ,
		\u2_adr0_cnt_reg[21]/P0001 ,
		_w799_
	);
	LUT4 #(
		.INIT('h4000)
	) name65 (
		_w757_,
		_w759_,
		_w760_,
		_w799_,
		_w800_
	);
	LUT3 #(
		.INIT('h13)
	) name66 (
		\u2_adr0_cnt_reg[22]/P0001 ,
		\u2_adr0_cnt_reg[23]/P0001 ,
		_w800_,
		_w801_
	);
	LUT3 #(
		.INIT('h2a)
	) name67 (
		_w750_,
		_w761_,
		_w762_,
		_w802_
	);
	LUT3 #(
		.INIT('hba)
	) name68 (
		_w798_,
		_w801_,
		_w802_,
		_w803_
	);
	LUT4 #(
		.INIT('h6a00)
	) name69 (
		\u2_adr1_cnt_reg[23]/P0001 ,
		_w742_,
		_w744_,
		_w750_,
		_w804_
	);
	LUT4 #(
		.INIT('h20aa)
	) name70 (
		\u0_u0_ch_adr1_r_reg[23]/P0001 ,
		_w747_,
		_w748_,
		_w749_,
		_w805_
	);
	LUT2 #(
		.INIT('he)
	) name71 (
		_w804_,
		_w805_,
		_w806_
	);
	LUT4 #(
		.INIT('h3aca)
	) name72 (
		\u0_u0_ch_adr0_r_reg[22]/P0001 ,
		\u2_adr0_cnt_reg[22]/P0001 ,
		_w750_,
		_w800_,
		_w807_
	);
	LUT4 #(
		.INIT('h20aa)
	) name73 (
		\u0_u0_ch_adr1_r_reg[22]/P0001 ,
		_w747_,
		_w748_,
		_w749_,
		_w808_
	);
	LUT4 #(
		.INIT('h6c00)
	) name74 (
		\u2_adr1_cnt_reg[21]/P0001 ,
		\u2_adr1_cnt_reg[22]/P0001 ,
		_w742_,
		_w750_,
		_w809_
	);
	LUT2 #(
		.INIT('he)
	) name75 (
		_w808_,
		_w809_,
		_w810_
	);
	LUT3 #(
		.INIT('h40)
	) name76 (
		_w757_,
		_w759_,
		_w760_,
		_w811_
	);
	LUT4 #(
		.INIT('h4555)
	) name77 (
		\u2_adr0_cnt_reg[20]/P0001 ,
		_w757_,
		_w759_,
		_w760_,
		_w812_
	);
	LUT4 #(
		.INIT('h222e)
	) name78 (
		\u0_u0_ch_adr0_r_reg[20]/P0001 ,
		_w750_,
		_w761_,
		_w812_,
		_w813_
	);
	LUT4 #(
		.INIT('h20aa)
	) name79 (
		\u0_u0_ch_adr1_r_reg[20]/P0001 ,
		_w747_,
		_w748_,
		_w749_,
		_w814_
	);
	LUT2 #(
		.INIT('h8)
	) name80 (
		\u2_adr1_cnt_reg[18]/P0001 ,
		\u2_adr1_cnt_reg[19]/P0001 ,
		_w815_
	);
	LUT4 #(
		.INIT('h4000)
	) name81 (
		_w737_,
		_w738_,
		_w740_,
		_w815_,
		_w816_
	);
	LUT4 #(
		.INIT('h3020)
	) name82 (
		\u2_adr1_cnt_reg[20]/P0001 ,
		_w742_,
		_w750_,
		_w816_,
		_w817_
	);
	LUT2 #(
		.INIT('he)
	) name83 (
		_w814_,
		_w817_,
		_w818_
	);
	LUT4 #(
		.INIT('h8000)
	) name84 (
		\u0_u0_ch_csr_r_reg[4]/NET0131 ,
		\u2_adr0_cnt_reg[16]/NET0131 ,
		\u2_read_r_reg/P0001 ,
		\u2_u0_out_r_reg[16]/P0001 ,
		_w819_
	);
	LUT2 #(
		.INIT('h4)
	) name85 (
		_w757_,
		_w819_,
		_w820_
	);
	LUT2 #(
		.INIT('h8)
	) name86 (
		\u2_adr0_cnt_reg[17]/P0001 ,
		\u2_adr0_cnt_reg[18]/P0001 ,
		_w821_
	);
	LUT3 #(
		.INIT('h40)
	) name87 (
		_w757_,
		_w819_,
		_w821_,
		_w822_
	);
	LUT4 #(
		.INIT('h4555)
	) name88 (
		\u2_adr0_cnt_reg[19]/P0001 ,
		_w757_,
		_w819_,
		_w821_,
		_w823_
	);
	LUT4 #(
		.INIT('h222e)
	) name89 (
		\u0_u0_ch_adr0_r_reg[19]/P0001 ,
		_w750_,
		_w811_,
		_w823_,
		_w824_
	);
	LUT4 #(
		.INIT('h8000)
	) name90 (
		\u2_adr1_cnt_reg[16]/NET0131 ,
		\u2_adr1_cnt_reg[17]/P0001 ,
		\u2_adr1_cnt_reg[18]/P0001 ,
		\u2_u1_out_r_reg[16]/P0001 ,
		_w825_
	);
	LUT3 #(
		.INIT('h40)
	) name91 (
		_w737_,
		_w738_,
		_w825_,
		_w826_
	);
	LUT4 #(
		.INIT('h4555)
	) name92 (
		\u2_adr1_cnt_reg[19]/P0001 ,
		_w737_,
		_w738_,
		_w825_,
		_w827_
	);
	LUT4 #(
		.INIT('h222e)
	) name93 (
		\u0_u0_ch_adr1_r_reg[19]/P0001 ,
		_w750_,
		_w816_,
		_w827_,
		_w828_
	);
	LUT4 #(
		.INIT('h3133)
	) name94 (
		\u2_adr0_cnt_reg[17]/P0001 ,
		\u2_adr0_cnt_reg[18]/P0001 ,
		_w757_,
		_w819_,
		_w829_
	);
	LUT4 #(
		.INIT('h222e)
	) name95 (
		\u0_u0_ch_adr0_r_reg[18]/P0001 ,
		_w750_,
		_w822_,
		_w829_,
		_w830_
	);
	LUT4 #(
		.INIT('h4555)
	) name96 (
		\u2_adr1_cnt_reg[18]/P0001 ,
		_w737_,
		_w738_,
		_w740_,
		_w831_
	);
	LUT4 #(
		.INIT('h222e)
	) name97 (
		\u0_u0_ch_adr1_r_reg[18]/P0001 ,
		_w750_,
		_w826_,
		_w831_,
		_w832_
	);
	LUT4 #(
		.INIT('h4500)
	) name98 (
		\u2_adr0_cnt_reg[29]/P0001 ,
		_w747_,
		_w748_,
		_w749_,
		_w833_
	);
	LUT4 #(
		.INIT('h7f00)
	) name99 (
		\u2_adr0_cnt_reg[28]/P0001 ,
		_w761_,
		_w765_,
		_w833_,
		_w834_
	);
	LUT4 #(
		.INIT('h8a00)
	) name100 (
		\u2_adr0_cnt_reg[29]/P0001 ,
		_w747_,
		_w748_,
		_w749_,
		_w835_
	);
	LUT4 #(
		.INIT('h8000)
	) name101 (
		\u2_adr0_cnt_reg[28]/P0001 ,
		_w761_,
		_w765_,
		_w835_,
		_w836_
	);
	LUT4 #(
		.INIT('h1055)
	) name102 (
		\u0_u0_ch_adr0_r_reg[29]/P0001 ,
		_w747_,
		_w748_,
		_w749_,
		_w837_
	);
	LUT3 #(
		.INIT('h01)
	) name103 (
		_w834_,
		_w836_,
		_w837_,
		_w838_
	);
	LUT2 #(
		.INIT('h1)
	) name104 (
		\u2_chunk_cnt_reg[6]/NET0131 ,
		\u2_chunk_cnt_reg[7]/NET0131 ,
		_w839_
	);
	LUT4 #(
		.INIT('h0001)
	) name105 (
		\u2_chunk_cnt_reg[0]/NET0131 ,
		\u2_chunk_cnt_reg[1]/NET0131 ,
		\u2_chunk_cnt_reg[2]/NET0131 ,
		\u2_chunk_cnt_reg[3]/NET0131 ,
		_w840_
	);
	LUT3 #(
		.INIT('h01)
	) name106 (
		\u2_chunk_cnt_reg[4]/NET0131 ,
		\u2_chunk_cnt_reg[5]/NET0131 ,
		\u2_chunk_cnt_reg[8]/NET0131 ,
		_w841_
	);
	LUT4 #(
		.INIT('h0001)
	) name107 (
		\u2_chunk_0_reg/P0001 ,
		\u2_chunk_cnt_reg[4]/NET0131 ,
		\u2_chunk_cnt_reg[5]/NET0131 ,
		\u2_chunk_cnt_reg[8]/NET0131 ,
		_w842_
	);
	LUT3 #(
		.INIT('h80)
	) name108 (
		_w839_,
		_w840_,
		_w842_,
		_w843_
	);
	LUT2 #(
		.INIT('h1)
	) name109 (
		\u0_u0_ch_sz_inf_reg/NET0131 ,
		\u2_tsz_cnt_reg[0]/NET0131 ,
		_w844_
	);
	LUT4 #(
		.INIT('h0001)
	) name110 (
		\u2_tsz_cnt_reg[10]/NET0131 ,
		\u2_tsz_cnt_reg[11]/NET0131 ,
		\u2_tsz_cnt_reg[1]/NET0131 ,
		\u2_tsz_cnt_reg[2]/NET0131 ,
		_w845_
	);
	LUT3 #(
		.INIT('h01)
	) name111 (
		\u2_tsz_cnt_reg[7]/NET0131 ,
		\u2_tsz_cnt_reg[8]/NET0131 ,
		\u2_tsz_cnt_reg[9]/NET0131 ,
		_w846_
	);
	LUT2 #(
		.INIT('h1)
	) name112 (
		\u2_tsz_cnt_reg[5]/NET0131 ,
		\u2_tsz_cnt_reg[6]/NET0131 ,
		_w847_
	);
	LUT4 #(
		.INIT('h0001)
	) name113 (
		\u2_tsz_cnt_reg[3]/NET0131 ,
		\u2_tsz_cnt_reg[4]/NET0131 ,
		\u2_tsz_cnt_reg[5]/NET0131 ,
		\u2_tsz_cnt_reg[6]/NET0131 ,
		_w848_
	);
	LUT4 #(
		.INIT('h8000)
	) name114 (
		_w844_,
		_w845_,
		_w846_,
		_w848_,
		_w849_
	);
	LUT2 #(
		.INIT('h4)
	) name115 (
		\u2_state_reg[1]/NET0131 ,
		\u2_state_reg[2]/NET0131 ,
		_w850_
	);
	LUT3 #(
		.INIT('h10)
	) name116 (
		\u2_dma_abort_r_reg/NET0131 ,
		\u2_state_reg[1]/NET0131 ,
		\u2_state_reg[2]/NET0131 ,
		_w851_
	);
	LUT2 #(
		.INIT('h4)
	) name117 (
		_w737_,
		_w851_,
		_w852_
	);
	LUT3 #(
		.INIT('h10)
	) name118 (
		_w843_,
		_w849_,
		_w852_,
		_w853_
	);
	LUT3 #(
		.INIT('h04)
	) name119 (
		\u2_dma_abort_r_reg/NET0131 ,
		\u2_state_reg[1]/NET0131 ,
		\u2_state_reg[2]/NET0131 ,
		_w854_
	);
	LUT2 #(
		.INIT('h8)
	) name120 (
		_w757_,
		_w854_,
		_w855_
	);
	LUT4 #(
		.INIT('h00ef)
	) name121 (
		_w843_,
		_w849_,
		_w852_,
		_w855_,
		_w856_
	);
	LUT4 #(
		.INIT('hff10)
	) name122 (
		_w843_,
		_w849_,
		_w852_,
		_w855_,
		_w857_
	);
	LUT4 #(
		.INIT('h4c5f)
	) name123 (
		_w737_,
		_w757_,
		_w851_,
		_w854_,
		_w858_
	);
	LUT4 #(
		.INIT('hb3a0)
	) name124 (
		_w737_,
		_w757_,
		_w851_,
		_w854_,
		_w859_
	);
	LUT2 #(
		.INIT('h1)
	) name125 (
		\u0_u0_ch_csr_r_reg[1]/NET0131 ,
		_w858_,
		_w860_
	);
	LUT4 #(
		.INIT('h0001)
	) name126 (
		\u2_state_reg[10]/NET0131 ,
		\u2_state_reg[3]/NET0131 ,
		\u2_state_reg[8]/NET0131 ,
		\u2_state_reg[9]/NET0131 ,
		_w861_
	);
	LUT2 #(
		.INIT('h4)
	) name127 (
		\u2_state_reg[7]/NET0131 ,
		_w861_,
		_w862_
	);
	LUT3 #(
		.INIT('h01)
	) name128 (
		\u2_state_reg[0]/NET0131 ,
		\u2_state_reg[1]/NET0131 ,
		\u2_state_reg[2]/NET0131 ,
		_w863_
	);
	LUT2 #(
		.INIT('h8)
	) name129 (
		\u2_state_reg[4]/NET0131 ,
		\u2_state_reg[6]/NET0131 ,
		_w864_
	);
	LUT3 #(
		.INIT('h01)
	) name130 (
		\u2_state_reg[4]/NET0131 ,
		\u2_state_reg[5]/NET0131 ,
		\u2_state_reg[6]/NET0131 ,
		_w865_
	);
	LUT3 #(
		.INIT('h36)
	) name131 (
		\u2_state_reg[4]/NET0131 ,
		\u2_state_reg[5]/NET0131 ,
		\u2_state_reg[6]/NET0131 ,
		_w866_
	);
	LUT3 #(
		.INIT('h20)
	) name132 (
		_w863_,
		_w864_,
		_w866_,
		_w867_
	);
	LUT2 #(
		.INIT('h1)
	) name133 (
		\u2_state_reg[7]/NET0131 ,
		\u2_state_reg[9]/NET0131 ,
		_w868_
	);
	LUT4 #(
		.INIT('h8000)
	) name134 (
		\u0_u0_ch_csr_r_reg[7]/NET0131 ,
		\u0_u0_ch_csr_r_reg[8]/NET0131 ,
		\u1_ndr_r_reg[0]/NET0131 ,
		\u2_state_reg[3]/NET0131 ,
		_w869_
	);
	LUT3 #(
		.INIT('h0e)
	) name135 (
		\u2_state_reg[7]/NET0131 ,
		\u2_state_reg[9]/NET0131 ,
		\wb0_ack_i_pad ,
		_w870_
	);
	LUT3 #(
		.INIT('h2e)
	) name136 (
		\wb0_ack_i_pad ,
		_w868_,
		_w869_,
		_w871_
	);
	LUT3 #(
		.INIT('h70)
	) name137 (
		_w862_,
		_w867_,
		_w871_,
		_w872_
	);
	LUT4 #(
		.INIT('h0e00)
	) name138 (
		\u0_u0_ch_csr_r_reg[2]/NET0131 ,
		_w856_,
		_w860_,
		_w872_,
		_w873_
	);
	LUT4 #(
		.INIT('h005f)
	) name139 (
		_w737_,
		_w757_,
		_w851_,
		_w854_,
		_w874_
	);
	LUT4 #(
		.INIT('hef00)
	) name140 (
		_w843_,
		_w849_,
		_w852_,
		_w874_,
		_w875_
	);
	LUT4 #(
		.INIT('h10ff)
	) name141 (
		_w843_,
		_w849_,
		_w852_,
		_w874_,
		_w876_
	);
	LUT2 #(
		.INIT('h4)
	) name142 (
		\u0_u0_ch_csr_r_reg[1]/NET0131 ,
		\u2_write_hold_r_reg/P0001 ,
		_w877_
	);
	LUT2 #(
		.INIT('h4)
	) name143 (
		_w875_,
		_w877_,
		_w878_
	);
	LUT3 #(
		.INIT('h01)
	) name144 (
		_w843_,
		_w849_,
		_w858_,
		_w879_
	);
	LUT4 #(
		.INIT('h5f1f)
	) name145 (
		\u0_u0_ch_csr_r_reg[2]/NET0131 ,
		_w856_,
		_w872_,
		_w879_,
		_w880_
	);
	LUT2 #(
		.INIT('he)
	) name146 (
		_w878_,
		_w880_,
		_w881_
	);
	LUT3 #(
		.INIT('h54)
	) name147 (
		_w873_,
		_w878_,
		_w880_,
		_w882_
	);
	LUT4 #(
		.INIT('h8000)
	) name148 (
		\u2_adr1_cnt_reg[25]/P0001 ,
		\u2_adr1_cnt_reg[26]/P0001 ,
		\u2_adr1_cnt_reg[27]/P0001 ,
		\u2_adr1_cnt_reg[28]/P0001 ,
		_w883_
	);
	LUT4 #(
		.INIT('h4500)
	) name149 (
		\u2_adr1_cnt_reg[29]/P0001 ,
		_w747_,
		_w748_,
		_w749_,
		_w884_
	);
	LUT4 #(
		.INIT('h7f00)
	) name150 (
		_w742_,
		_w794_,
		_w883_,
		_w884_,
		_w885_
	);
	LUT4 #(
		.INIT('h8a00)
	) name151 (
		\u2_adr1_cnt_reg[29]/P0001 ,
		_w747_,
		_w748_,
		_w749_,
		_w886_
	);
	LUT4 #(
		.INIT('h8000)
	) name152 (
		_w742_,
		_w794_,
		_w883_,
		_w886_,
		_w887_
	);
	LUT4 #(
		.INIT('h1055)
	) name153 (
		\u0_u0_ch_adr1_r_reg[29]/P0001 ,
		_w747_,
		_w748_,
		_w749_,
		_w888_
	);
	LUT3 #(
		.INIT('h01)
	) name154 (
		_w885_,
		_w887_,
		_w888_,
		_w889_
	);
	LUT3 #(
		.INIT('h2a)
	) name155 (
		\u2_adr1_cnt_reg[0]/P0001 ,
		_w757_,
		_w854_,
		_w890_
	);
	LUT4 #(
		.INIT('hef00)
	) name156 (
		_w843_,
		_w849_,
		_w852_,
		_w890_,
		_w891_
	);
	LUT4 #(
		.INIT('h0fdf)
	) name157 (
		\u2_adr0_cnt_reg[0]/P0001 ,
		_w856_,
		_w872_,
		_w891_,
		_w892_
	);
	LUT3 #(
		.INIT('h07)
	) name158 (
		_w862_,
		_w867_,
		_w870_,
		_w893_
	);
	LUT4 #(
		.INIT('h0001)
	) name159 (
		\u2_state_reg[0]/NET0131 ,
		\u2_state_reg[1]/NET0131 ,
		\u2_state_reg[2]/NET0131 ,
		\u2_state_reg[3]/NET0131 ,
		_w894_
	);
	LUT4 #(
		.INIT('h0001)
	) name160 (
		\u2_state_reg[4]/NET0131 ,
		\u2_state_reg[5]/NET0131 ,
		\u2_state_reg[6]/NET0131 ,
		\u2_state_reg[7]/NET0131 ,
		_w895_
	);
	LUT3 #(
		.INIT('h10)
	) name161 (
		\u2_state_reg[10]/NET0131 ,
		\u2_state_reg[8]/NET0131 ,
		\u2_state_reg[9]/NET0131 ,
		_w896_
	);
	LUT3 #(
		.INIT('h80)
	) name162 (
		_w894_,
		_w895_,
		_w896_,
		_w897_
	);
	LUT4 #(
		.INIT('h1555)
	) name163 (
		_w869_,
		_w894_,
		_w895_,
		_w896_,
		_w898_
	);
	LUT2 #(
		.INIT('h1)
	) name164 (
		\u2_state_reg[1]/NET0131 ,
		\u2_state_reg[2]/NET0131 ,
		_w899_
	);
	LUT2 #(
		.INIT('h1)
	) name165 (
		\u2_state_reg[0]/NET0131 ,
		\u2_state_reg[5]/NET0131 ,
		_w900_
	);
	LUT3 #(
		.INIT('h10)
	) name166 (
		\u2_state_reg[4]/NET0131 ,
		\u2_state_reg[6]/NET0131 ,
		\u2_state_reg[7]/NET0131 ,
		_w901_
	);
	LUT4 #(
		.INIT('h8000)
	) name167 (
		_w861_,
		_w899_,
		_w900_,
		_w901_,
		_w902_
	);
	LUT4 #(
		.INIT('h05fb)
	) name168 (
		\u2_state_reg[4]/NET0131 ,
		\u2_state_reg[5]/NET0131 ,
		\u2_state_reg[6]/NET0131 ,
		\wb0_ack_i_pad ,
		_w903_
	);
	LUT3 #(
		.INIT('h8a)
	) name169 (
		_w898_,
		_w902_,
		_w903_,
		_w904_
	);
	LUT2 #(
		.INIT('h4)
	) name170 (
		_w893_,
		_w904_,
		_w905_
	);
	LUT2 #(
		.INIT('hd)
	) name171 (
		_w892_,
		_w905_,
		_w906_
	);
	LUT3 #(
		.INIT('h2a)
	) name172 (
		\u2_adr1_cnt_reg[1]/P0001 ,
		_w757_,
		_w854_,
		_w907_
	);
	LUT4 #(
		.INIT('hef00)
	) name173 (
		_w843_,
		_w849_,
		_w852_,
		_w907_,
		_w908_
	);
	LUT4 #(
		.INIT('h0fdf)
	) name174 (
		\u2_adr0_cnt_reg[1]/P0001 ,
		_w856_,
		_w872_,
		_w908_,
		_w909_
	);
	LUT2 #(
		.INIT('h1)
	) name175 (
		\u2_state_reg[5]/NET0131 ,
		\u2_state_reg[6]/NET0131 ,
		_w910_
	);
	LUT4 #(
		.INIT('hfcf8)
	) name176 (
		\u2_state_reg[4]/NET0131 ,
		\u2_state_reg[5]/NET0131 ,
		\u2_state_reg[6]/NET0131 ,
		\wb0_ack_i_pad ,
		_w911_
	);
	LUT3 #(
		.INIT('ha8)
	) name177 (
		_w898_,
		_w902_,
		_w911_,
		_w912_
	);
	LUT2 #(
		.INIT('h4)
	) name178 (
		_w893_,
		_w912_,
		_w913_
	);
	LUT2 #(
		.INIT('hd)
	) name179 (
		_w909_,
		_w913_,
		_w914_
	);
	LUT4 #(
		.INIT('h5355)
	) name180 (
		\u2_adr0_cnt_reg[0]/P0001 ,
		\u2_u0_out_r_reg[0]/P0001 ,
		_w757_,
		_w758_,
		_w915_
	);
	LUT3 #(
		.INIT('h2e)
	) name181 (
		\u0_u0_ch_adr0_r_reg[0]/P0001 ,
		_w750_,
		_w915_,
		_w916_
	);
	LUT4 #(
		.INIT('h5355)
	) name182 (
		\u2_adr0_cnt_reg[10]/P0001 ,
		\u2_u0_out_r_reg[10]/P0001 ,
		_w757_,
		_w758_,
		_w917_
	);
	LUT3 #(
		.INIT('h2e)
	) name183 (
		\u0_u0_ch_adr0_r_reg[10]/P0001 ,
		_w750_,
		_w917_,
		_w918_
	);
	LUT4 #(
		.INIT('h5355)
	) name184 (
		\u2_adr0_cnt_reg[11]/P0001 ,
		\u2_u0_out_r_reg[11]/P0001 ,
		_w757_,
		_w758_,
		_w919_
	);
	LUT3 #(
		.INIT('h2e)
	) name185 (
		\u0_u0_ch_adr0_r_reg[11]/P0001 ,
		_w750_,
		_w919_,
		_w920_
	);
	LUT4 #(
		.INIT('h5355)
	) name186 (
		\u2_adr0_cnt_reg[12]/P0001 ,
		\u2_u0_out_r_reg[12]/P0001 ,
		_w757_,
		_w758_,
		_w921_
	);
	LUT3 #(
		.INIT('h2e)
	) name187 (
		\u0_u0_ch_adr0_r_reg[12]/P0001 ,
		_w750_,
		_w921_,
		_w922_
	);
	LUT4 #(
		.INIT('h5355)
	) name188 (
		\u2_adr0_cnt_reg[14]/P0001 ,
		\u2_u0_out_r_reg[14]/P0001 ,
		_w757_,
		_w758_,
		_w923_
	);
	LUT3 #(
		.INIT('h2e)
	) name189 (
		\u0_u0_ch_adr0_r_reg[14]/P0001 ,
		_w750_,
		_w923_,
		_w924_
	);
	LUT4 #(
		.INIT('h5355)
	) name190 (
		\u2_adr0_cnt_reg[15]/P0001 ,
		\u2_u0_out_r_reg[15]/P0001 ,
		_w757_,
		_w758_,
		_w925_
	);
	LUT3 #(
		.INIT('h2e)
	) name191 (
		\u0_u0_ch_adr0_r_reg[15]/P0001 ,
		_w750_,
		_w925_,
		_w926_
	);
	LUT4 #(
		.INIT('ha6aa)
	) name192 (
		\u2_adr0_cnt_reg[16]/NET0131 ,
		\u2_u0_out_r_reg[16]/P0001 ,
		_w757_,
		_w758_,
		_w927_
	);
	LUT3 #(
		.INIT('he2)
	) name193 (
		\u0_u0_ch_adr0_r_reg[16]/P0001 ,
		_w750_,
		_w927_,
		_w928_
	);
	LUT4 #(
		.INIT('h3aca)
	) name194 (
		\u0_u0_ch_adr0_r_reg[17]/P0001 ,
		\u2_adr0_cnt_reg[17]/P0001 ,
		_w750_,
		_w820_,
		_w929_
	);
	LUT4 #(
		.INIT('h5355)
	) name195 (
		\u2_adr0_cnt_reg[1]/P0001 ,
		\u2_u0_out_r_reg[1]/P0001 ,
		_w757_,
		_w758_,
		_w930_
	);
	LUT3 #(
		.INIT('h2e)
	) name196 (
		\u0_u0_ch_adr0_r_reg[1]/P0001 ,
		_w750_,
		_w930_,
		_w931_
	);
	LUT4 #(
		.INIT('h00c8)
	) name197 (
		\u2_adr0_cnt_reg[21]/P0001 ,
		_w750_,
		_w761_,
		_w800_,
		_w932_
	);
	LUT4 #(
		.INIT('h20aa)
	) name198 (
		\u0_u0_ch_adr0_r_reg[21]/P0001 ,
		_w747_,
		_w748_,
		_w749_,
		_w933_
	);
	LUT2 #(
		.INIT('he)
	) name199 (
		_w932_,
		_w933_,
		_w934_
	);
	LUT4 #(
		.INIT('h20aa)
	) name200 (
		\u0_u0_ch_adr0_r_reg[25]/P0001 ,
		_w747_,
		_w748_,
		_w749_,
		_w935_
	);
	LUT3 #(
		.INIT('h15)
	) name201 (
		\u2_adr0_cnt_reg[25]/P0001 ,
		_w761_,
		_w788_,
		_w936_
	);
	LUT3 #(
		.INIT('h2a)
	) name202 (
		_w750_,
		_w761_,
		_w783_,
		_w937_
	);
	LUT3 #(
		.INIT('hba)
	) name203 (
		_w935_,
		_w936_,
		_w937_,
		_w938_
	);
	LUT4 #(
		.INIT('h5355)
	) name204 (
		\u2_adr0_cnt_reg[2]/P0001 ,
		\u2_u0_out_r_reg[2]/P0001 ,
		_w757_,
		_w758_,
		_w939_
	);
	LUT3 #(
		.INIT('h2e)
	) name205 (
		\u0_u0_ch_adr0_r_reg[2]/P0001 ,
		_w750_,
		_w939_,
		_w940_
	);
	LUT4 #(
		.INIT('h5355)
	) name206 (
		\u2_adr0_cnt_reg[3]/P0001 ,
		\u2_u0_out_r_reg[3]/P0001 ,
		_w757_,
		_w758_,
		_w941_
	);
	LUT3 #(
		.INIT('h2e)
	) name207 (
		\u0_u0_ch_adr0_r_reg[3]/P0001 ,
		_w750_,
		_w941_,
		_w942_
	);
	LUT4 #(
		.INIT('h5355)
	) name208 (
		\u2_adr0_cnt_reg[4]/P0001 ,
		\u2_u0_out_r_reg[4]/P0001 ,
		_w757_,
		_w758_,
		_w943_
	);
	LUT3 #(
		.INIT('h2e)
	) name209 (
		\u0_u0_ch_adr0_r_reg[4]/P0001 ,
		_w750_,
		_w943_,
		_w944_
	);
	LUT4 #(
		.INIT('h5355)
	) name210 (
		\u2_adr0_cnt_reg[5]/P0001 ,
		\u2_u0_out_r_reg[5]/P0001 ,
		_w757_,
		_w758_,
		_w945_
	);
	LUT3 #(
		.INIT('h2e)
	) name211 (
		\u0_u0_ch_adr0_r_reg[5]/P0001 ,
		_w750_,
		_w945_,
		_w946_
	);
	LUT4 #(
		.INIT('h5355)
	) name212 (
		\u2_adr0_cnt_reg[6]/P0001 ,
		\u2_u0_out_r_reg[6]/P0001 ,
		_w757_,
		_w758_,
		_w947_
	);
	LUT3 #(
		.INIT('h2e)
	) name213 (
		\u0_u0_ch_adr0_r_reg[6]/P0001 ,
		_w750_,
		_w947_,
		_w948_
	);
	LUT4 #(
		.INIT('h5355)
	) name214 (
		\u2_adr0_cnt_reg[7]/P0001 ,
		\u2_u0_out_r_reg[7]/P0001 ,
		_w757_,
		_w758_,
		_w949_
	);
	LUT3 #(
		.INIT('h2e)
	) name215 (
		\u0_u0_ch_adr0_r_reg[7]/P0001 ,
		_w750_,
		_w949_,
		_w950_
	);
	LUT4 #(
		.INIT('h5355)
	) name216 (
		\u2_adr0_cnt_reg[8]/P0001 ,
		\u2_u0_out_r_reg[8]/P0001 ,
		_w757_,
		_w758_,
		_w951_
	);
	LUT3 #(
		.INIT('h2e)
	) name217 (
		\u0_u0_ch_adr0_r_reg[8]/P0001 ,
		_w750_,
		_w951_,
		_w952_
	);
	LUT4 #(
		.INIT('h5355)
	) name218 (
		\u2_adr0_cnt_reg[9]/P0001 ,
		\u2_u0_out_r_reg[9]/P0001 ,
		_w757_,
		_w758_,
		_w953_
	);
	LUT3 #(
		.INIT('h2e)
	) name219 (
		\u0_u0_ch_adr0_r_reg[9]/P0001 ,
		_w750_,
		_w953_,
		_w954_
	);
	LUT2 #(
		.INIT('h2)
	) name220 (
		\u0_u0_ch_csr_r_reg[1]/NET0131 ,
		_w858_,
		_w955_
	);
	LUT3 #(
		.INIT('h31)
	) name221 (
		\u0_u0_ch_csr_r_reg[1]/NET0131 ,
		\u0_u0_ch_csr_r_reg[2]/NET0131 ,
		_w858_,
		_w956_
	);
	LUT3 #(
		.INIT('h31)
	) name222 (
		\u0_u0_ch_csr_r_reg[1]/NET0131 ,
		_w855_,
		_w858_,
		_w957_
	);
	LUT3 #(
		.INIT('h23)
	) name223 (
		_w853_,
		_w956_,
		_w957_,
		_w958_
	);
	LUT3 #(
		.INIT('ha2)
	) name224 (
		\u0_u0_ch_csr_r_reg[2]/NET0131 ,
		_w856_,
		_w879_,
		_w959_
	);
	LUT2 #(
		.INIT('h8)
	) name225 (
		\u0_u0_ch_csr_r_reg[1]/NET0131 ,
		\u2_write_hold_r_reg/P0001 ,
		_w960_
	);
	LUT2 #(
		.INIT('h4)
	) name226 (
		_w875_,
		_w960_,
		_w961_
	);
	LUT2 #(
		.INIT('he)
	) name227 (
		_w959_,
		_w961_,
		_w962_
	);
	LUT3 #(
		.INIT('ha8)
	) name228 (
		_w958_,
		_w959_,
		_w961_,
		_w963_
	);
	LUT4 #(
		.INIT('h9aaa)
	) name229 (
		\u2_adr1_cnt_reg[17]/P0001 ,
		_w737_,
		_w738_,
		_w739_,
		_w964_
	);
	LUT3 #(
		.INIT('he2)
	) name230 (
		\u0_u0_ch_adr1_r_reg[17]/P0001 ,
		_w750_,
		_w964_,
		_w965_
	);
	LUT4 #(
		.INIT('h3caa)
	) name231 (
		\u0_u0_ch_adr1_r_reg[21]/P0001 ,
		\u2_adr1_cnt_reg[21]/P0001 ,
		_w742_,
		_w750_,
		_w966_
	);
	LUT3 #(
		.INIT('h2a)
	) name232 (
		\u2_adr1_cnt_reg[9]/P0001 ,
		_w757_,
		_w854_,
		_w967_
	);
	LUT4 #(
		.INIT('hef00)
	) name233 (
		_w843_,
		_w849_,
		_w852_,
		_w967_,
		_w968_
	);
	LUT4 #(
		.INIT('hf020)
	) name234 (
		\u2_adr0_cnt_reg[9]/P0001 ,
		_w856_,
		_w872_,
		_w968_,
		_w969_
	);
	LUT3 #(
		.INIT('h2a)
	) name235 (
		\u2_adr1_cnt_reg[10]/P0001 ,
		_w757_,
		_w854_,
		_w970_
	);
	LUT4 #(
		.INIT('hef00)
	) name236 (
		_w843_,
		_w849_,
		_w852_,
		_w970_,
		_w971_
	);
	LUT4 #(
		.INIT('hf020)
	) name237 (
		\u2_adr0_cnt_reg[10]/P0001 ,
		_w856_,
		_w872_,
		_w971_,
		_w972_
	);
	LUT3 #(
		.INIT('h2a)
	) name238 (
		\u2_adr1_cnt_reg[11]/P0001 ,
		_w757_,
		_w854_,
		_w973_
	);
	LUT4 #(
		.INIT('hef00)
	) name239 (
		_w843_,
		_w849_,
		_w852_,
		_w973_,
		_w974_
	);
	LUT4 #(
		.INIT('hf020)
	) name240 (
		\u2_adr0_cnt_reg[11]/P0001 ,
		_w856_,
		_w872_,
		_w974_,
		_w975_
	);
	LUT3 #(
		.INIT('h2a)
	) name241 (
		\u2_adr1_cnt_reg[12]/P0001 ,
		_w757_,
		_w854_,
		_w976_
	);
	LUT4 #(
		.INIT('hef00)
	) name242 (
		_w843_,
		_w849_,
		_w852_,
		_w976_,
		_w977_
	);
	LUT4 #(
		.INIT('hf020)
	) name243 (
		\u2_adr0_cnt_reg[12]/P0001 ,
		_w856_,
		_w872_,
		_w977_,
		_w978_
	);
	LUT3 #(
		.INIT('h2a)
	) name244 (
		\u2_adr1_cnt_reg[13]/P0001 ,
		_w757_,
		_w854_,
		_w979_
	);
	LUT4 #(
		.INIT('hef00)
	) name245 (
		_w843_,
		_w849_,
		_w852_,
		_w979_,
		_w980_
	);
	LUT4 #(
		.INIT('hf020)
	) name246 (
		\u2_adr0_cnt_reg[13]/P0001 ,
		_w856_,
		_w872_,
		_w980_,
		_w981_
	);
	LUT3 #(
		.INIT('h2a)
	) name247 (
		\u2_adr1_cnt_reg[14]/P0001 ,
		_w757_,
		_w854_,
		_w982_
	);
	LUT4 #(
		.INIT('hef00)
	) name248 (
		_w843_,
		_w849_,
		_w852_,
		_w982_,
		_w983_
	);
	LUT4 #(
		.INIT('hf020)
	) name249 (
		\u2_adr0_cnt_reg[14]/P0001 ,
		_w856_,
		_w872_,
		_w983_,
		_w984_
	);
	LUT3 #(
		.INIT('h2a)
	) name250 (
		\u2_adr1_cnt_reg[15]/P0001 ,
		_w757_,
		_w854_,
		_w985_
	);
	LUT4 #(
		.INIT('hef00)
	) name251 (
		_w843_,
		_w849_,
		_w852_,
		_w985_,
		_w986_
	);
	LUT4 #(
		.INIT('hf020)
	) name252 (
		\u2_adr0_cnt_reg[15]/P0001 ,
		_w856_,
		_w872_,
		_w986_,
		_w987_
	);
	LUT3 #(
		.INIT('h2a)
	) name253 (
		\u2_adr1_cnt_reg[16]/NET0131 ,
		_w757_,
		_w854_,
		_w988_
	);
	LUT4 #(
		.INIT('hef00)
	) name254 (
		_w843_,
		_w849_,
		_w852_,
		_w988_,
		_w989_
	);
	LUT4 #(
		.INIT('hf020)
	) name255 (
		\u2_adr0_cnt_reg[16]/NET0131 ,
		_w856_,
		_w872_,
		_w989_,
		_w990_
	);
	LUT3 #(
		.INIT('h2a)
	) name256 (
		\u2_adr1_cnt_reg[17]/P0001 ,
		_w757_,
		_w854_,
		_w991_
	);
	LUT4 #(
		.INIT('hef00)
	) name257 (
		_w843_,
		_w849_,
		_w852_,
		_w991_,
		_w992_
	);
	LUT4 #(
		.INIT('hf020)
	) name258 (
		\u2_adr0_cnt_reg[17]/P0001 ,
		_w856_,
		_w872_,
		_w992_,
		_w993_
	);
	LUT3 #(
		.INIT('h2a)
	) name259 (
		\u2_adr1_cnt_reg[18]/P0001 ,
		_w757_,
		_w854_,
		_w994_
	);
	LUT4 #(
		.INIT('hef00)
	) name260 (
		_w843_,
		_w849_,
		_w852_,
		_w994_,
		_w995_
	);
	LUT4 #(
		.INIT('hf020)
	) name261 (
		\u2_adr0_cnt_reg[18]/P0001 ,
		_w856_,
		_w872_,
		_w995_,
		_w996_
	);
	LUT3 #(
		.INIT('h2a)
	) name262 (
		\u2_adr1_cnt_reg[19]/P0001 ,
		_w757_,
		_w854_,
		_w997_
	);
	LUT4 #(
		.INIT('hef00)
	) name263 (
		_w843_,
		_w849_,
		_w852_,
		_w997_,
		_w998_
	);
	LUT4 #(
		.INIT('hf020)
	) name264 (
		\u2_adr0_cnt_reg[19]/P0001 ,
		_w856_,
		_w872_,
		_w998_,
		_w999_
	);
	LUT3 #(
		.INIT('h2a)
	) name265 (
		\u2_adr1_cnt_reg[20]/P0001 ,
		_w757_,
		_w854_,
		_w1000_
	);
	LUT4 #(
		.INIT('hef00)
	) name266 (
		_w843_,
		_w849_,
		_w852_,
		_w1000_,
		_w1001_
	);
	LUT4 #(
		.INIT('hf020)
	) name267 (
		\u2_adr0_cnt_reg[20]/P0001 ,
		_w856_,
		_w872_,
		_w1001_,
		_w1002_
	);
	LUT3 #(
		.INIT('h2a)
	) name268 (
		\u2_adr1_cnt_reg[21]/P0001 ,
		_w757_,
		_w854_,
		_w1003_
	);
	LUT4 #(
		.INIT('hef00)
	) name269 (
		_w843_,
		_w849_,
		_w852_,
		_w1003_,
		_w1004_
	);
	LUT4 #(
		.INIT('hf020)
	) name270 (
		\u2_adr0_cnt_reg[21]/P0001 ,
		_w856_,
		_w872_,
		_w1004_,
		_w1005_
	);
	LUT3 #(
		.INIT('h2a)
	) name271 (
		\u2_adr1_cnt_reg[22]/P0001 ,
		_w757_,
		_w854_,
		_w1006_
	);
	LUT4 #(
		.INIT('hef00)
	) name272 (
		_w843_,
		_w849_,
		_w852_,
		_w1006_,
		_w1007_
	);
	LUT4 #(
		.INIT('hf020)
	) name273 (
		\u2_adr0_cnt_reg[22]/P0001 ,
		_w856_,
		_w872_,
		_w1007_,
		_w1008_
	);
	LUT3 #(
		.INIT('h2a)
	) name274 (
		\u2_adr1_cnt_reg[23]/P0001 ,
		_w757_,
		_w854_,
		_w1009_
	);
	LUT4 #(
		.INIT('hef00)
	) name275 (
		_w843_,
		_w849_,
		_w852_,
		_w1009_,
		_w1010_
	);
	LUT4 #(
		.INIT('hf020)
	) name276 (
		\u2_adr0_cnt_reg[23]/P0001 ,
		_w856_,
		_w872_,
		_w1010_,
		_w1011_
	);
	LUT3 #(
		.INIT('h2a)
	) name277 (
		\u2_adr1_cnt_reg[24]/P0001 ,
		_w757_,
		_w854_,
		_w1012_
	);
	LUT4 #(
		.INIT('hef00)
	) name278 (
		_w843_,
		_w849_,
		_w852_,
		_w1012_,
		_w1013_
	);
	LUT4 #(
		.INIT('hf020)
	) name279 (
		\u2_adr0_cnt_reg[24]/P0001 ,
		_w856_,
		_w872_,
		_w1013_,
		_w1014_
	);
	LUT3 #(
		.INIT('h2a)
	) name280 (
		\u2_adr1_cnt_reg[25]/P0001 ,
		_w757_,
		_w854_,
		_w1015_
	);
	LUT4 #(
		.INIT('hef00)
	) name281 (
		_w843_,
		_w849_,
		_w852_,
		_w1015_,
		_w1016_
	);
	LUT4 #(
		.INIT('hf020)
	) name282 (
		\u2_adr0_cnt_reg[25]/P0001 ,
		_w856_,
		_w872_,
		_w1016_,
		_w1017_
	);
	LUT3 #(
		.INIT('h2a)
	) name283 (
		\u2_adr1_cnt_reg[26]/P0001 ,
		_w757_,
		_w854_,
		_w1018_
	);
	LUT4 #(
		.INIT('hef00)
	) name284 (
		_w843_,
		_w849_,
		_w852_,
		_w1018_,
		_w1019_
	);
	LUT4 #(
		.INIT('hf020)
	) name285 (
		\u2_adr0_cnt_reg[26]/P0001 ,
		_w856_,
		_w872_,
		_w1019_,
		_w1020_
	);
	LUT3 #(
		.INIT('h2a)
	) name286 (
		\u2_adr1_cnt_reg[27]/P0001 ,
		_w757_,
		_w854_,
		_w1021_
	);
	LUT4 #(
		.INIT('hef00)
	) name287 (
		_w843_,
		_w849_,
		_w852_,
		_w1021_,
		_w1022_
	);
	LUT4 #(
		.INIT('hf020)
	) name288 (
		\u2_adr0_cnt_reg[27]/P0001 ,
		_w856_,
		_w872_,
		_w1022_,
		_w1023_
	);
	LUT3 #(
		.INIT('h2a)
	) name289 (
		\u2_adr1_cnt_reg[28]/P0001 ,
		_w757_,
		_w854_,
		_w1024_
	);
	LUT4 #(
		.INIT('hef00)
	) name290 (
		_w843_,
		_w849_,
		_w852_,
		_w1024_,
		_w1025_
	);
	LUT4 #(
		.INIT('hf020)
	) name291 (
		\u2_adr0_cnt_reg[28]/P0001 ,
		_w856_,
		_w872_,
		_w1025_,
		_w1026_
	);
	LUT3 #(
		.INIT('h2a)
	) name292 (
		\u2_adr1_cnt_reg[29]/P0001 ,
		_w757_,
		_w854_,
		_w1027_
	);
	LUT4 #(
		.INIT('hef00)
	) name293 (
		_w843_,
		_w849_,
		_w852_,
		_w1027_,
		_w1028_
	);
	LUT4 #(
		.INIT('hf020)
	) name294 (
		\u2_adr0_cnt_reg[29]/P0001 ,
		_w856_,
		_w872_,
		_w1028_,
		_w1029_
	);
	LUT3 #(
		.INIT('h2a)
	) name295 (
		\u2_adr1_cnt_reg[8]/P0001 ,
		_w757_,
		_w854_,
		_w1030_
	);
	LUT4 #(
		.INIT('hef00)
	) name296 (
		_w843_,
		_w849_,
		_w852_,
		_w1030_,
		_w1031_
	);
	LUT4 #(
		.INIT('hf020)
	) name297 (
		\u2_adr0_cnt_reg[8]/P0001 ,
		_w856_,
		_w872_,
		_w1031_,
		_w1032_
	);
	LUT3 #(
		.INIT('h2a)
	) name298 (
		\u2_adr1_cnt_reg[2]/P0001 ,
		_w757_,
		_w854_,
		_w1033_
	);
	LUT4 #(
		.INIT('hef00)
	) name299 (
		_w843_,
		_w849_,
		_w852_,
		_w1033_,
		_w1034_
	);
	LUT4 #(
		.INIT('hf020)
	) name300 (
		\u2_adr0_cnt_reg[2]/P0001 ,
		_w856_,
		_w872_,
		_w1034_,
		_w1035_
	);
	LUT3 #(
		.INIT('h2a)
	) name301 (
		\u2_adr1_cnt_reg[3]/P0001 ,
		_w757_,
		_w854_,
		_w1036_
	);
	LUT4 #(
		.INIT('hef00)
	) name302 (
		_w843_,
		_w849_,
		_w852_,
		_w1036_,
		_w1037_
	);
	LUT4 #(
		.INIT('hf020)
	) name303 (
		\u2_adr0_cnt_reg[3]/P0001 ,
		_w856_,
		_w872_,
		_w1037_,
		_w1038_
	);
	LUT3 #(
		.INIT('h2a)
	) name304 (
		\u2_adr1_cnt_reg[4]/P0001 ,
		_w757_,
		_w854_,
		_w1039_
	);
	LUT4 #(
		.INIT('hef00)
	) name305 (
		_w843_,
		_w849_,
		_w852_,
		_w1039_,
		_w1040_
	);
	LUT4 #(
		.INIT('hf020)
	) name306 (
		\u2_adr0_cnt_reg[4]/P0001 ,
		_w856_,
		_w872_,
		_w1040_,
		_w1041_
	);
	LUT3 #(
		.INIT('h2a)
	) name307 (
		\u2_adr1_cnt_reg[5]/P0001 ,
		_w757_,
		_w854_,
		_w1042_
	);
	LUT4 #(
		.INIT('hef00)
	) name308 (
		_w843_,
		_w849_,
		_w852_,
		_w1042_,
		_w1043_
	);
	LUT4 #(
		.INIT('hf020)
	) name309 (
		\u2_adr0_cnt_reg[5]/P0001 ,
		_w856_,
		_w872_,
		_w1043_,
		_w1044_
	);
	LUT3 #(
		.INIT('h2a)
	) name310 (
		\u2_adr1_cnt_reg[6]/P0001 ,
		_w757_,
		_w854_,
		_w1045_
	);
	LUT4 #(
		.INIT('hef00)
	) name311 (
		_w843_,
		_w849_,
		_w852_,
		_w1045_,
		_w1046_
	);
	LUT4 #(
		.INIT('hf020)
	) name312 (
		\u2_adr0_cnt_reg[6]/P0001 ,
		_w856_,
		_w872_,
		_w1046_,
		_w1047_
	);
	LUT3 #(
		.INIT('h2a)
	) name313 (
		\u2_adr1_cnt_reg[7]/P0001 ,
		_w757_,
		_w854_,
		_w1048_
	);
	LUT4 #(
		.INIT('hef00)
	) name314 (
		_w843_,
		_w849_,
		_w852_,
		_w1048_,
		_w1049_
	);
	LUT4 #(
		.INIT('hf020)
	) name315 (
		\u2_adr0_cnt_reg[7]/P0001 ,
		_w856_,
		_w872_,
		_w1049_,
		_w1050_
	);
	LUT4 #(
		.INIT('h0001)
	) name316 (
		\u3_u1_slv_adr_reg[6]/NET0131 ,
		\u3_u1_slv_adr_reg[7]/NET0131 ,
		\u3_u1_slv_adr_reg[8]/NET0131 ,
		\u3_u1_slv_adr_reg[9]/NET0131 ,
		_w1051_
	);
	LUT2 #(
		.INIT('h1)
	) name317 (
		\u3_u1_slv_adr_reg[2]/NET0131 ,
		\u3_u1_slv_adr_reg[3]/P0001 ,
		_w1052_
	);
	LUT3 #(
		.INIT('h10)
	) name318 (
		\u3_u1_slv_adr_reg[2]/NET0131 ,
		\u3_u1_slv_adr_reg[3]/P0001 ,
		\u3_u1_slv_adr_reg[5]/P0001 ,
		_w1053_
	);
	LUT2 #(
		.INIT('h4)
	) name319 (
		\u3_u1_slv_adr_reg[4]/NET0131 ,
		\u3_u1_slv_we_reg/P0001 ,
		_w1054_
	);
	LUT3 #(
		.INIT('h10)
	) name320 (
		\u3_u1_slv_adr_reg[4]/NET0131 ,
		\u3_u1_slv_dout_reg[0]/P0001 ,
		\u3_u1_slv_we_reg/P0001 ,
		_w1055_
	);
	LUT3 #(
		.INIT('h80)
	) name321 (
		_w1051_,
		_w1053_,
		_w1055_,
		_w1056_
	);
	LUT3 #(
		.INIT('h80)
	) name322 (
		_w1051_,
		_w1053_,
		_w1054_,
		_w1057_
	);
	LUT4 #(
		.INIT('h1555)
	) name323 (
		\u0_u0_ch_csr_r_reg[0]/NET0131 ,
		_w1051_,
		_w1053_,
		_w1054_,
		_w1058_
	);
	LUT2 #(
		.INIT('h1)
	) name324 (
		\u1_ndnr_reg[0]/P0001 ,
		\u2_state_reg[3]/NET0131 ,
		_w1059_
	);
	LUT4 #(
		.INIT('h0002)
	) name325 (
		\u1_ndr_r_reg[0]/NET0131 ,
		\u2_chunk_cnt_reg[4]/NET0131 ,
		\u2_chunk_cnt_reg[5]/NET0131 ,
		\u2_chunk_cnt_reg[8]/NET0131 ,
		_w1060_
	);
	LUT2 #(
		.INIT('h1)
	) name326 (
		\u1_ndnr_reg[0]/P0001 ,
		\u2_tsz_cnt_is_0_r_reg/P0001 ,
		_w1061_
	);
	LUT4 #(
		.INIT('h7f00)
	) name327 (
		_w839_,
		_w840_,
		_w1060_,
		_w1061_,
		_w1062_
	);
	LUT2 #(
		.INIT('h1)
	) name328 (
		\u0_u0_ch_csr_r_reg[6]/NET0131 ,
		\u0_u0_ch_csr_r_reg[7]/NET0131 ,
		_w1063_
	);
	LUT4 #(
		.INIT('h7f00)
	) name329 (
		_w1051_,
		_w1053_,
		_w1054_,
		_w1063_,
		_w1064_
	);
	LUT4 #(
		.INIT('h5455)
	) name330 (
		_w1058_,
		_w1059_,
		_w1062_,
		_w1064_,
		_w1065_
	);
	LUT2 #(
		.INIT('h4)
	) name331 (
		_w1056_,
		_w1065_,
		_w1066_
	);
	LUT4 #(
		.INIT('h0001)
	) name332 (
		\u2_state_reg[10]/NET0131 ,
		\u2_state_reg[7]/NET0131 ,
		\u2_state_reg[8]/NET0131 ,
		\u2_state_reg[9]/NET0131 ,
		_w1067_
	);
	LUT4 #(
		.INIT('h0001)
	) name333 (
		\u2_state_reg[3]/NET0131 ,
		\u2_state_reg[4]/NET0131 ,
		\u2_state_reg[5]/NET0131 ,
		\u2_state_reg[6]/NET0131 ,
		_w1068_
	);
	LUT3 #(
		.INIT('h40)
	) name334 (
		\u2_state_reg[0]/NET0131 ,
		_w1067_,
		_w1068_,
		_w1069_
	);
	LUT4 #(
		.INIT('h048c)
	) name335 (
		\u0_u0_ch_csr_r_reg[1]/NET0131 ,
		\u2_state_reg[1]/NET0131 ,
		\wb0_ack_i_pad ,
		\wb1_ack_i_pad ,
		_w1070_
	);
	LUT2 #(
		.INIT('h8)
	) name336 (
		_w851_,
		_w1070_,
		_w1071_
	);
	LUT4 #(
		.INIT('h00ef)
	) name337 (
		_w843_,
		_w849_,
		_w852_,
		_w1071_,
		_w1072_
	);
	LUT4 #(
		.INIT('h0010)
	) name338 (
		\u2_state_reg[10]/NET0131 ,
		\u2_state_reg[7]/NET0131 ,
		\u2_state_reg[8]/NET0131 ,
		\u2_state_reg[9]/NET0131 ,
		_w1073_
	);
	LUT3 #(
		.INIT('h80)
	) name339 (
		_w865_,
		_w894_,
		_w1073_,
		_w1074_
	);
	LUT3 #(
		.INIT('h45)
	) name340 (
		\u1_next_start_reg/P0001 ,
		_w747_,
		_w748_,
		_w1075_
	);
	LUT2 #(
		.INIT('h2)
	) name341 (
		\u0_u0_ch_csr_r_reg[7]/NET0131 ,
		\u0_u0_ch_err_reg/NET0131 ,
		_w1076_
	);
	LUT4 #(
		.INIT('hba00)
	) name342 (
		\u1_next_start_reg/P0001 ,
		_w747_,
		_w748_,
		_w1076_,
		_w1077_
	);
	LUT3 #(
		.INIT('h02)
	) name343 (
		\u2_state_reg[0]/NET0131 ,
		\u2_state_reg[1]/NET0131 ,
		\u2_state_reg[2]/NET0131 ,
		_w1078_
	);
	LUT4 #(
		.INIT('h0004)
	) name344 (
		\u0_csr_r_reg[0]/NET0131 ,
		\u2_state_reg[0]/NET0131 ,
		\u2_state_reg[1]/NET0131 ,
		\u2_state_reg[2]/NET0131 ,
		_w1079_
	);
	LUT3 #(
		.INIT('h80)
	) name345 (
		_w1067_,
		_w1068_,
		_w1079_,
		_w1080_
	);
	LUT2 #(
		.INIT('h2)
	) name346 (
		\u0_u0_ch_err_reg/NET0131 ,
		\u2_state_reg[1]/NET0131 ,
		_w1081_
	);
	LUT2 #(
		.INIT('h1)
	) name347 (
		\u1_next_start_reg/P0001 ,
		\u2_state_reg[1]/NET0131 ,
		_w1082_
	);
	LUT4 #(
		.INIT('h040f)
	) name348 (
		_w747_,
		_w748_,
		_w1081_,
		_w1082_,
		_w1083_
	);
	LUT4 #(
		.INIT('h4555)
	) name349 (
		_w1074_,
		_w1077_,
		_w1080_,
		_w1083_,
		_w1084_
	);
	LUT4 #(
		.INIT('h8cff)
	) name350 (
		_w855_,
		_w1069_,
		_w1072_,
		_w1084_,
		_w1085_
	);
	LUT4 #(
		.INIT('h4544)
	) name351 (
		\u0_u0_ch_err_reg/NET0131 ,
		\u1_next_start_reg/P0001 ,
		_w747_,
		_w748_,
		_w1086_
	);
	LUT2 #(
		.INIT('h2)
	) name352 (
		_w1080_,
		_w1086_,
		_w1087_
	);
	LUT3 #(
		.INIT('h80)
	) name353 (
		\u0_u0_ch_csr_r_reg[7]/NET0131 ,
		\u0_u0_ch_csr_r_reg[8]/NET0131 ,
		\u1_ndr_r_reg[0]/NET0131 ,
		_w1088_
	);
	LUT2 #(
		.INIT('h2)
	) name354 (
		\u2_state_reg[3]/NET0131 ,
		\u2_state_reg[4]/NET0131 ,
		_w1089_
	);
	LUT4 #(
		.INIT('h8000)
	) name355 (
		_w863_,
		_w910_,
		_w1067_,
		_w1089_,
		_w1090_
	);
	LUT4 #(
		.INIT('h8000)
	) name356 (
		\wb0_ack_i_pad ,
		_w894_,
		_w895_,
		_w896_,
		_w1091_
	);
	LUT2 #(
		.INIT('h2)
	) name357 (
		\u2_state_reg[10]/NET0131 ,
		\u2_state_reg[8]/NET0131 ,
		_w1092_
	);
	LUT4 #(
		.INIT('h000d)
	) name358 (
		\u0_csr_r_reg[0]/NET0131 ,
		\u2_state_reg[0]/NET0131 ,
		\u2_state_reg[7]/NET0131 ,
		\u2_state_reg[9]/NET0131 ,
		_w1093_
	);
	LUT4 #(
		.INIT('h8000)
	) name359 (
		_w865_,
		_w894_,
		_w1092_,
		_w1093_,
		_w1094_
	);
	LUT4 #(
		.INIT('h000b)
	) name360 (
		_w1088_,
		_w1090_,
		_w1091_,
		_w1094_,
		_w1095_
	);
	LUT2 #(
		.INIT('hb)
	) name361 (
		_w1087_,
		_w1095_,
		_w1096_
	);
	LUT3 #(
		.INIT('h10)
	) name362 (
		\u3_u1_slv_adr_reg[3]/P0001 ,
		\u3_u1_slv_adr_reg[4]/NET0131 ,
		\u3_u1_slv_adr_reg[5]/P0001 ,
		_w1097_
	);
	LUT2 #(
		.INIT('h4)
	) name363 (
		\u3_u1_slv_adr_reg[2]/NET0131 ,
		\u3_u1_slv_re_reg/P0001 ,
		_w1098_
	);
	LUT4 #(
		.INIT('h2aaa)
	) name364 (
		\u0_u0_int_src_r_reg[1]/NET0131 ,
		_w1051_,
		_w1097_,
		_w1098_,
		_w1099_
	);
	LUT4 #(
		.INIT('hff10)
	) name365 (
		_w1059_,
		_w1062_,
		_w1063_,
		_w1099_,
		_w1100_
	);
	LUT4 #(
		.INIT('ha6aa)
	) name366 (
		\u2_adr1_cnt_reg[16]/NET0131 ,
		\u2_u1_out_r_reg[16]/P0001 ,
		_w737_,
		_w738_,
		_w1101_
	);
	LUT3 #(
		.INIT('he2)
	) name367 (
		\u0_u0_ch_adr1_r_reg[16]/P0001 ,
		_w750_,
		_w1101_,
		_w1102_
	);
	LUT2 #(
		.INIT('h1)
	) name368 (
		\u2_read_r_reg/P0001 ,
		_w856_,
		_w1103_
	);
	LUT3 #(
		.INIT('h08)
	) name369 (
		\u2_dma_abort_r_reg/NET0131 ,
		\u2_state_reg[1]/NET0131 ,
		\u2_state_reg[2]/NET0131 ,
		_w1104_
	);
	LUT3 #(
		.INIT('h20)
	) name370 (
		\u2_state_reg[1]/NET0131 ,
		\u2_state_reg[2]/NET0131 ,
		\u2_state_reg[3]/NET0131 ,
		_w1105_
	);
	LUT3 #(
		.INIT('h13)
	) name371 (
		_w757_,
		_w1104_,
		_w1105_,
		_w1106_
	);
	LUT2 #(
		.INIT('h2)
	) name372 (
		_w1069_,
		_w1106_,
		_w1107_
	);
	LUT4 #(
		.INIT('h0123)
	) name373 (
		\u0_u0_ch_csr_r_reg[1]/NET0131 ,
		\u2_state_reg[3]/NET0131 ,
		\wb0_ack_i_pad ,
		\wb1_ack_i_pad ,
		_w1108_
	);
	LUT2 #(
		.INIT('h4)
	) name374 (
		\u2_dma_abort_r_reg/NET0131 ,
		_w1108_,
		_w1109_
	);
	LUT4 #(
		.INIT('h3210)
	) name375 (
		\u0_u0_ch_csr_r_reg[1]/NET0131 ,
		\u2_dma_abort_r_reg/NET0131 ,
		\wb0_ack_i_pad ,
		\wb1_ack_i_pad ,
		_w1110_
	);
	LUT4 #(
		.INIT('h0e0f)
	) name376 (
		_w843_,
		_w849_,
		_w1109_,
		_w1110_,
		_w1111_
	);
	LUT4 #(
		.INIT('h4000)
	) name377 (
		\u2_state_reg[0]/NET0131 ,
		_w850_,
		_w1067_,
		_w1068_,
		_w1112_
	);
	LUT3 #(
		.INIT('hea)
	) name378 (
		_w1107_,
		_w1111_,
		_w1112_,
		_w1113_
	);
	LUT3 #(
		.INIT('hf2)
	) name379 (
		\u2_adr0_cnt_reg[9]/P0001 ,
		_w856_,
		_w968_,
		_w1114_
	);
	LUT3 #(
		.INIT('hf2)
	) name380 (
		\u2_adr0_cnt_reg[8]/P0001 ,
		_w856_,
		_w1031_,
		_w1115_
	);
	LUT3 #(
		.INIT('hf2)
	) name381 (
		\u2_adr0_cnt_reg[10]/P0001 ,
		_w856_,
		_w971_,
		_w1116_
	);
	LUT3 #(
		.INIT('hf2)
	) name382 (
		\u2_adr0_cnt_reg[11]/P0001 ,
		_w856_,
		_w974_,
		_w1117_
	);
	LUT3 #(
		.INIT('hf2)
	) name383 (
		\u2_adr0_cnt_reg[12]/P0001 ,
		_w856_,
		_w977_,
		_w1118_
	);
	LUT3 #(
		.INIT('hf2)
	) name384 (
		\u2_adr0_cnt_reg[13]/P0001 ,
		_w856_,
		_w980_,
		_w1119_
	);
	LUT3 #(
		.INIT('hf2)
	) name385 (
		\u2_adr0_cnt_reg[14]/P0001 ,
		_w856_,
		_w983_,
		_w1120_
	);
	LUT3 #(
		.INIT('hf2)
	) name386 (
		\u2_adr0_cnt_reg[15]/P0001 ,
		_w856_,
		_w986_,
		_w1121_
	);
	LUT3 #(
		.INIT('hf2)
	) name387 (
		\u2_adr0_cnt_reg[16]/NET0131 ,
		_w856_,
		_w989_,
		_w1122_
	);
	LUT3 #(
		.INIT('hf2)
	) name388 (
		\u2_adr0_cnt_reg[17]/P0001 ,
		_w856_,
		_w992_,
		_w1123_
	);
	LUT3 #(
		.INIT('hf2)
	) name389 (
		\u2_adr0_cnt_reg[18]/P0001 ,
		_w856_,
		_w995_,
		_w1124_
	);
	LUT3 #(
		.INIT('hf2)
	) name390 (
		\u2_adr0_cnt_reg[19]/P0001 ,
		_w856_,
		_w998_,
		_w1125_
	);
	LUT3 #(
		.INIT('hf2)
	) name391 (
		\u2_adr0_cnt_reg[20]/P0001 ,
		_w856_,
		_w1001_,
		_w1126_
	);
	LUT3 #(
		.INIT('hf2)
	) name392 (
		\u2_adr0_cnt_reg[21]/P0001 ,
		_w856_,
		_w1004_,
		_w1127_
	);
	LUT3 #(
		.INIT('hf2)
	) name393 (
		\u2_adr0_cnt_reg[22]/P0001 ,
		_w856_,
		_w1007_,
		_w1128_
	);
	LUT3 #(
		.INIT('hf2)
	) name394 (
		\u2_adr0_cnt_reg[23]/P0001 ,
		_w856_,
		_w1010_,
		_w1129_
	);
	LUT3 #(
		.INIT('hf2)
	) name395 (
		\u2_adr0_cnt_reg[24]/P0001 ,
		_w856_,
		_w1013_,
		_w1130_
	);
	LUT3 #(
		.INIT('hf2)
	) name396 (
		\u2_adr0_cnt_reg[25]/P0001 ,
		_w856_,
		_w1016_,
		_w1131_
	);
	LUT3 #(
		.INIT('hf2)
	) name397 (
		\u2_adr0_cnt_reg[26]/P0001 ,
		_w856_,
		_w1019_,
		_w1132_
	);
	LUT3 #(
		.INIT('hf2)
	) name398 (
		\u2_adr0_cnt_reg[27]/P0001 ,
		_w856_,
		_w1022_,
		_w1133_
	);
	LUT3 #(
		.INIT('hf2)
	) name399 (
		\u2_adr0_cnt_reg[0]/P0001 ,
		_w856_,
		_w891_,
		_w1134_
	);
	LUT3 #(
		.INIT('hf2)
	) name400 (
		\u2_adr0_cnt_reg[28]/P0001 ,
		_w856_,
		_w1025_,
		_w1135_
	);
	LUT3 #(
		.INIT('hf2)
	) name401 (
		\u2_adr0_cnt_reg[29]/P0001 ,
		_w856_,
		_w1028_,
		_w1136_
	);
	LUT3 #(
		.INIT('hf2)
	) name402 (
		\u2_adr0_cnt_reg[1]/P0001 ,
		_w856_,
		_w908_,
		_w1137_
	);
	LUT3 #(
		.INIT('hf2)
	) name403 (
		\u2_adr0_cnt_reg[2]/P0001 ,
		_w856_,
		_w1034_,
		_w1138_
	);
	LUT3 #(
		.INIT('hf2)
	) name404 (
		\u2_adr0_cnt_reg[3]/P0001 ,
		_w856_,
		_w1037_,
		_w1139_
	);
	LUT3 #(
		.INIT('hf2)
	) name405 (
		\u2_adr0_cnt_reg[4]/P0001 ,
		_w856_,
		_w1040_,
		_w1140_
	);
	LUT3 #(
		.INIT('hf2)
	) name406 (
		\u2_adr0_cnt_reg[5]/P0001 ,
		_w856_,
		_w1043_,
		_w1141_
	);
	LUT3 #(
		.INIT('hf2)
	) name407 (
		\u2_adr0_cnt_reg[6]/P0001 ,
		_w856_,
		_w1046_,
		_w1142_
	);
	LUT3 #(
		.INIT('hf2)
	) name408 (
		\u2_adr0_cnt_reg[7]/P0001 ,
		_w856_,
		_w1049_,
		_w1143_
	);
	LUT2 #(
		.INIT('h8)
	) name409 (
		_w1088_,
		_w1090_,
		_w1144_
	);
	LUT4 #(
		.INIT('h0001)
	) name410 (
		\u2_state_reg[0]/NET0131 ,
		\u2_state_reg[1]/NET0131 ,
		\u2_state_reg[2]/NET0131 ,
		\u2_state_reg[5]/NET0131 ,
		_w1145_
	);
	LUT3 #(
		.INIT('h10)
	) name411 (
		\u2_state_reg[3]/NET0131 ,
		\u2_state_reg[4]/NET0131 ,
		\u2_state_reg[6]/NET0131 ,
		_w1146_
	);
	LUT3 #(
		.INIT('h80)
	) name412 (
		_w1067_,
		_w1145_,
		_w1146_,
		_w1147_
	);
	LUT2 #(
		.INIT('h2)
	) name413 (
		\u2_state_reg[9]/NET0131 ,
		\wb0_ack_i_pad ,
		_w1148_
	);
	LUT3 #(
		.INIT('he0)
	) name414 (
		_w897_,
		_w1147_,
		_w1148_,
		_w1149_
	);
	LUT2 #(
		.INIT('he)
	) name415 (
		_w1144_,
		_w1149_,
		_w1150_
	);
	LUT4 #(
		.INIT('h5355)
	) name416 (
		\u2_adr1_cnt_reg[2]/P0001 ,
		\u2_u1_out_r_reg[2]/P0001 ,
		_w737_,
		_w738_,
		_w1151_
	);
	LUT3 #(
		.INIT('h2e)
	) name417 (
		\u0_u0_ch_adr1_r_reg[2]/P0001 ,
		_w750_,
		_w1151_,
		_w1152_
	);
	LUT4 #(
		.INIT('h5355)
	) name418 (
		\u2_adr1_cnt_reg[3]/P0001 ,
		\u2_u1_out_r_reg[3]/P0001 ,
		_w737_,
		_w738_,
		_w1153_
	);
	LUT3 #(
		.INIT('h2e)
	) name419 (
		\u0_u0_ch_adr1_r_reg[3]/P0001 ,
		_w750_,
		_w1153_,
		_w1154_
	);
	LUT4 #(
		.INIT('h5355)
	) name420 (
		\u2_adr1_cnt_reg[4]/P0001 ,
		\u2_u1_out_r_reg[4]/P0001 ,
		_w737_,
		_w738_,
		_w1155_
	);
	LUT3 #(
		.INIT('h2e)
	) name421 (
		\u0_u0_ch_adr1_r_reg[4]/P0001 ,
		_w750_,
		_w1155_,
		_w1156_
	);
	LUT4 #(
		.INIT('h5355)
	) name422 (
		\u2_adr1_cnt_reg[5]/P0001 ,
		\u2_u1_out_r_reg[5]/P0001 ,
		_w737_,
		_w738_,
		_w1157_
	);
	LUT3 #(
		.INIT('h2e)
	) name423 (
		\u0_u0_ch_adr1_r_reg[5]/P0001 ,
		_w750_,
		_w1157_,
		_w1158_
	);
	LUT4 #(
		.INIT('h5355)
	) name424 (
		\u2_adr1_cnt_reg[6]/P0001 ,
		\u2_u1_out_r_reg[6]/P0001 ,
		_w737_,
		_w738_,
		_w1159_
	);
	LUT3 #(
		.INIT('h2e)
	) name425 (
		\u0_u0_ch_adr1_r_reg[6]/P0001 ,
		_w750_,
		_w1159_,
		_w1160_
	);
	LUT4 #(
		.INIT('h5355)
	) name426 (
		\u2_adr1_cnt_reg[7]/P0001 ,
		\u2_u1_out_r_reg[7]/P0001 ,
		_w737_,
		_w738_,
		_w1161_
	);
	LUT3 #(
		.INIT('h2e)
	) name427 (
		\u0_u0_ch_adr1_r_reg[7]/P0001 ,
		_w750_,
		_w1161_,
		_w1162_
	);
	LUT4 #(
		.INIT('h5355)
	) name428 (
		\u2_adr1_cnt_reg[8]/P0001 ,
		\u2_u1_out_r_reg[8]/P0001 ,
		_w737_,
		_w738_,
		_w1163_
	);
	LUT3 #(
		.INIT('h2e)
	) name429 (
		\u0_u0_ch_adr1_r_reg[8]/P0001 ,
		_w750_,
		_w1163_,
		_w1164_
	);
	LUT4 #(
		.INIT('h5355)
	) name430 (
		\u2_adr1_cnt_reg[9]/P0001 ,
		\u2_u1_out_r_reg[9]/P0001 ,
		_w737_,
		_w738_,
		_w1165_
	);
	LUT3 #(
		.INIT('h2e)
	) name431 (
		\u0_u0_ch_adr1_r_reg[9]/P0001 ,
		_w750_,
		_w1165_,
		_w1166_
	);
	LUT4 #(
		.INIT('h5355)
	) name432 (
		\u2_adr1_cnt_reg[0]/P0001 ,
		\u2_u1_out_r_reg[0]/P0001 ,
		_w737_,
		_w738_,
		_w1167_
	);
	LUT3 #(
		.INIT('h2e)
	) name433 (
		\u0_u0_ch_adr1_r_reg[0]/P0001 ,
		_w750_,
		_w1167_,
		_w1168_
	);
	LUT4 #(
		.INIT('h5355)
	) name434 (
		\u2_adr1_cnt_reg[10]/P0001 ,
		\u2_u1_out_r_reg[10]/P0001 ,
		_w737_,
		_w738_,
		_w1169_
	);
	LUT3 #(
		.INIT('h2e)
	) name435 (
		\u0_u0_ch_adr1_r_reg[10]/P0001 ,
		_w750_,
		_w1169_,
		_w1170_
	);
	LUT4 #(
		.INIT('h5355)
	) name436 (
		\u2_adr1_cnt_reg[11]/P0001 ,
		\u2_u1_out_r_reg[11]/P0001 ,
		_w737_,
		_w738_,
		_w1171_
	);
	LUT3 #(
		.INIT('h2e)
	) name437 (
		\u0_u0_ch_adr1_r_reg[11]/P0001 ,
		_w750_,
		_w1171_,
		_w1172_
	);
	LUT4 #(
		.INIT('h5355)
	) name438 (
		\u2_adr1_cnt_reg[12]/P0001 ,
		\u2_u1_out_r_reg[12]/P0001 ,
		_w737_,
		_w738_,
		_w1173_
	);
	LUT3 #(
		.INIT('h2e)
	) name439 (
		\u0_u0_ch_adr1_r_reg[12]/P0001 ,
		_w750_,
		_w1173_,
		_w1174_
	);
	LUT4 #(
		.INIT('h5355)
	) name440 (
		\u2_adr1_cnt_reg[13]/P0001 ,
		\u2_u1_out_r_reg[13]/P0001 ,
		_w737_,
		_w738_,
		_w1175_
	);
	LUT3 #(
		.INIT('h2e)
	) name441 (
		\u0_u0_ch_adr1_r_reg[13]/P0001 ,
		_w750_,
		_w1175_,
		_w1176_
	);
	LUT4 #(
		.INIT('h5355)
	) name442 (
		\u2_adr1_cnt_reg[14]/P0001 ,
		\u2_u1_out_r_reg[14]/P0001 ,
		_w737_,
		_w738_,
		_w1177_
	);
	LUT3 #(
		.INIT('h2e)
	) name443 (
		\u0_u0_ch_adr1_r_reg[14]/P0001 ,
		_w750_,
		_w1177_,
		_w1178_
	);
	LUT4 #(
		.INIT('h5355)
	) name444 (
		\u2_adr1_cnt_reg[15]/P0001 ,
		\u2_u1_out_r_reg[15]/P0001 ,
		_w737_,
		_w738_,
		_w1179_
	);
	LUT3 #(
		.INIT('h2e)
	) name445 (
		\u0_u0_ch_adr1_r_reg[15]/P0001 ,
		_w750_,
		_w1179_,
		_w1180_
	);
	LUT4 #(
		.INIT('h5355)
	) name446 (
		\u2_adr1_cnt_reg[1]/P0001 ,
		\u2_u1_out_r_reg[1]/P0001 ,
		_w737_,
		_w738_,
		_w1181_
	);
	LUT3 #(
		.INIT('h2e)
	) name447 (
		\u0_u0_ch_adr1_r_reg[1]/P0001 ,
		_w750_,
		_w1181_,
		_w1182_
	);
	LUT2 #(
		.INIT('h8)
	) name448 (
		\u0_u0_ch_csr_r_reg[0]/NET0131 ,
		\u2_next_ch_reg/P0001 ,
		_w1183_
	);
	LUT2 #(
		.INIT('h4)
	) name449 (
		_w747_,
		_w1183_,
		_w1184_
	);
	LUT2 #(
		.INIT('h8)
	) name450 (
		\u0_u0_ch_csr_r_reg[5]/NET0131 ,
		\u2_state_reg[3]/NET0131 ,
		_w1185_
	);
	LUT3 #(
		.INIT('he0)
	) name451 (
		_w843_,
		_w849_,
		_w1185_,
		_w1186_
	);
	LUT3 #(
		.INIT('ha8)
	) name452 (
		\u2_state_reg[3]/NET0131 ,
		_w843_,
		_w849_,
		_w1187_
	);
	LUT4 #(
		.INIT('h2aaa)
	) name453 (
		\u0_u0_int_src_r_reg[2]/NET0131 ,
		_w1051_,
		_w1097_,
		_w1098_,
		_w1188_
	);
	LUT4 #(
		.INIT('hffa8)
	) name454 (
		\u2_state_reg[3]/NET0131 ,
		_w843_,
		_w849_,
		_w1188_,
		_w1189_
	);
	LUT3 #(
		.INIT('h80)
	) name455 (
		_w1067_,
		_w1068_,
		_w1078_,
		_w1190_
	);
	LUT3 #(
		.INIT('h7f)
	) name456 (
		_w1067_,
		_w1068_,
		_w1078_,
		_w1191_
	);
	LUT4 #(
		.INIT('h0002)
	) name457 (
		\u2_state_reg[10]/NET0131 ,
		\u2_state_reg[7]/NET0131 ,
		\u2_state_reg[8]/NET0131 ,
		\u2_state_reg[9]/NET0131 ,
		_w1192_
	);
	LUT3 #(
		.INIT('h80)
	) name458 (
		_w865_,
		_w894_,
		_w1192_,
		_w1193_
	);
	LUT3 #(
		.INIT('ha8)
	) name459 (
		\u0_csr_r_reg[0]/NET0131 ,
		_w1190_,
		_w1193_,
		_w1194_
	);
	LUT4 #(
		.INIT('h0008)
	) name460 (
		\u2_state_reg[0]/NET0131 ,
		\u2_state_reg[10]/NET0131 ,
		\u2_state_reg[1]/NET0131 ,
		\u2_state_reg[2]/NET0131 ,
		_w1195_
	);
	LUT3 #(
		.INIT('h80)
	) name461 (
		_w1067_,
		_w1068_,
		_w1195_,
		_w1196_
	);
	LUT2 #(
		.INIT('h4)
	) name462 (
		_w1086_,
		_w1196_,
		_w1197_
	);
	LUT2 #(
		.INIT('he)
	) name463 (
		_w1194_,
		_w1197_,
		_w1198_
	);
	LUT2 #(
		.INIT('h8)
	) name464 (
		\u0_u0_ch_err_reg/NET0131 ,
		\u2_state_reg[4]/NET0131 ,
		_w1199_
	);
	LUT2 #(
		.INIT('h4)
	) name465 (
		\u1_next_start_reg/P0001 ,
		\u2_state_reg[4]/NET0131 ,
		_w1200_
	);
	LUT4 #(
		.INIT('h040f)
	) name466 (
		_w747_,
		_w748_,
		_w1199_,
		_w1200_,
		_w1201_
	);
	LUT3 #(
		.INIT('h8c)
	) name467 (
		_w1077_,
		_w1080_,
		_w1201_,
		_w1202_
	);
	LUT2 #(
		.INIT('h4)
	) name468 (
		\u2_state_reg[3]/NET0131 ,
		\u2_state_reg[4]/NET0131 ,
		_w1203_
	);
	LUT4 #(
		.INIT('h8000)
	) name469 (
		_w863_,
		_w910_,
		_w1067_,
		_w1203_,
		_w1204_
	);
	LUT2 #(
		.INIT('h2)
	) name470 (
		\u2_state_reg[4]/NET0131 ,
		\wb0_ack_i_pad ,
		_w1205_
	);
	LUT4 #(
		.INIT('hfe00)
	) name471 (
		_w897_,
		_w1147_,
		_w1204_,
		_w1205_,
		_w1206_
	);
	LUT2 #(
		.INIT('he)
	) name472 (
		_w1202_,
		_w1206_,
		_w1207_
	);
	LUT2 #(
		.INIT('h4)
	) name473 (
		_w858_,
		_w1069_,
		_w1208_
	);
	LUT4 #(
		.INIT('h0002)
	) name474 (
		\u2_chunk_dec_reg/P0001 ,
		\u2_tsz_cnt_is_0_r_reg/P0001 ,
		\u2_tsz_cnt_reg[0]/NET0131 ,
		\u2_tsz_cnt_reg[1]/NET0131 ,
		_w1209_
	);
	LUT3 #(
		.INIT('h01)
	) name475 (
		\u2_tsz_cnt_reg[2]/NET0131 ,
		\u2_tsz_cnt_reg[3]/NET0131 ,
		\u2_tsz_cnt_reg[4]/NET0131 ,
		_w1210_
	);
	LUT4 #(
		.INIT('h8000)
	) name476 (
		_w846_,
		_w847_,
		_w1209_,
		_w1210_,
		_w1211_
	);
	LUT4 #(
		.INIT('h3aca)
	) name477 (
		\u0_u0_ch_tot_sz_r_reg[10]/P0001 ,
		\u2_tsz_cnt_reg[10]/NET0131 ,
		_w750_,
		_w1211_,
		_w1212_
	);
	LUT4 #(
		.INIT('h9fcf)
	) name478 (
		\u2_tsz_cnt_reg[10]/NET0131 ,
		\u2_tsz_cnt_reg[11]/NET0131 ,
		_w750_,
		_w1211_,
		_w1213_
	);
	LUT4 #(
		.INIT('h1055)
	) name479 (
		\u0_u0_ch_tot_sz_r_reg[11]/P0001 ,
		_w747_,
		_w748_,
		_w749_,
		_w1214_
	);
	LUT2 #(
		.INIT('h2)
	) name480 (
		_w1213_,
		_w1214_,
		_w1215_
	);
	LUT4 #(
		.INIT('h02fd)
	) name481 (
		\u2_chunk_dec_reg/P0001 ,
		\u2_tsz_cnt_is_0_r_reg/P0001 ,
		\u2_tsz_cnt_reg[0]/NET0131 ,
		\u2_tsz_cnt_reg[1]/NET0131 ,
		_w1216_
	);
	LUT4 #(
		.INIT('h00b0)
	) name482 (
		_w747_,
		_w748_,
		_w749_,
		_w1216_,
		_w1217_
	);
	LUT4 #(
		.INIT('h20aa)
	) name483 (
		\u0_u0_ch_tot_sz_r_reg[1]/P0001 ,
		_w747_,
		_w748_,
		_w749_,
		_w1218_
	);
	LUT2 #(
		.INIT('he)
	) name484 (
		_w1217_,
		_w1218_,
		_w1219_
	);
	LUT3 #(
		.INIT('h63)
	) name485 (
		\u2_tsz_cnt_reg[2]/NET0131 ,
		\u2_tsz_cnt_reg[3]/NET0131 ,
		_w1209_,
		_w1220_
	);
	LUT3 #(
		.INIT('h2e)
	) name486 (
		\u0_u0_ch_tot_sz_r_reg[3]/P0001 ,
		_w750_,
		_w1220_,
		_w1221_
	);
	LUT4 #(
		.INIT('h0001)
	) name487 (
		\u2_tsz_cnt_reg[5]/NET0131 ,
		\u2_tsz_cnt_reg[6]/NET0131 ,
		\u2_tsz_cnt_reg[7]/NET0131 ,
		\u2_tsz_cnt_reg[8]/NET0131 ,
		_w1222_
	);
	LUT3 #(
		.INIT('h80)
	) name488 (
		_w1209_,
		_w1210_,
		_w1222_,
		_w1223_
	);
	LUT4 #(
		.INIT('h2aaa)
	) name489 (
		\u2_tsz_cnt_reg[9]/NET0131 ,
		_w1209_,
		_w1210_,
		_w1222_,
		_w1224_
	);
	LUT4 #(
		.INIT('heee2)
	) name490 (
		\u0_u0_ch_tot_sz_r_reg[9]/P0001 ,
		_w750_,
		_w1211_,
		_w1224_,
		_w1225_
	);
	LUT3 #(
		.INIT('h95)
	) name491 (
		\u2_tsz_cnt_reg[5]/NET0131 ,
		_w1209_,
		_w1210_,
		_w1226_
	);
	LUT3 #(
		.INIT('h2e)
	) name492 (
		\u0_u0_ch_tot_sz_r_reg[5]/P0001 ,
		_w750_,
		_w1226_,
		_w1227_
	);
	LUT4 #(
		.INIT('h6333)
	) name493 (
		\u2_tsz_cnt_reg[5]/NET0131 ,
		\u2_tsz_cnt_reg[6]/NET0131 ,
		_w1209_,
		_w1210_,
		_w1228_
	);
	LUT3 #(
		.INIT('h2e)
	) name494 (
		\u0_u0_ch_tot_sz_r_reg[6]/P0001 ,
		_w750_,
		_w1228_,
		_w1229_
	);
	LUT3 #(
		.INIT('h01)
	) name495 (
		\u2_tsz_cnt_reg[5]/NET0131 ,
		\u2_tsz_cnt_reg[6]/NET0131 ,
		\u2_tsz_cnt_reg[7]/NET0131 ,
		_w1230_
	);
	LUT3 #(
		.INIT('h80)
	) name496 (
		_w1209_,
		_w1210_,
		_w1230_,
		_w1231_
	);
	LUT4 #(
		.INIT('h2aaa)
	) name497 (
		\u2_tsz_cnt_reg[7]/NET0131 ,
		_w847_,
		_w1209_,
		_w1210_,
		_w1232_
	);
	LUT4 #(
		.INIT('heee2)
	) name498 (
		\u0_u0_ch_tot_sz_r_reg[7]/P0001 ,
		_w750_,
		_w1231_,
		_w1232_,
		_w1233_
	);
	LUT4 #(
		.INIT('h20aa)
	) name499 (
		\u0_u0_ch_tot_sz_r_reg[0]/P0001 ,
		_w747_,
		_w748_,
		_w749_,
		_w1234_
	);
	LUT3 #(
		.INIT('h2d)
	) name500 (
		\u2_chunk_dec_reg/P0001 ,
		\u2_tsz_cnt_is_0_r_reg/P0001 ,
		\u2_tsz_cnt_reg[0]/NET0131 ,
		_w1235_
	);
	LUT4 #(
		.INIT('h00b0)
	) name501 (
		_w747_,
		_w748_,
		_w749_,
		_w1235_,
		_w1236_
	);
	LUT2 #(
		.INIT('he)
	) name502 (
		_w1234_,
		_w1236_,
		_w1237_
	);
	LUT4 #(
		.INIT('h1e0f)
	) name503 (
		\u2_tsz_cnt_reg[2]/NET0131 ,
		\u2_tsz_cnt_reg[3]/NET0131 ,
		\u2_tsz_cnt_reg[4]/NET0131 ,
		_w1209_,
		_w1238_
	);
	LUT3 #(
		.INIT('h2e)
	) name504 (
		\u0_u0_ch_tot_sz_r_reg[4]/P0001 ,
		_w750_,
		_w1238_,
		_w1239_
	);
	LUT4 #(
		.INIT('h2aaa)
	) name505 (
		\u2_tsz_cnt_reg[8]/NET0131 ,
		_w1209_,
		_w1210_,
		_w1230_,
		_w1240_
	);
	LUT4 #(
		.INIT('heee2)
	) name506 (
		\u0_u0_ch_tot_sz_r_reg[8]/P0001 ,
		_w750_,
		_w1223_,
		_w1240_,
		_w1241_
	);
	LUT4 #(
		.INIT('h0100)
	) name507 (
		\u2_chunk_cnt_is_0_r_reg/P0001 ,
		\u2_chunk_cnt_reg[0]/NET0131 ,
		\u2_chunk_cnt_reg[1]/NET0131 ,
		\u2_chunk_dec_reg/P0001 ,
		_w1242_
	);
	LUT3 #(
		.INIT('h01)
	) name508 (
		\u2_chunk_cnt_reg[2]/NET0131 ,
		\u2_chunk_cnt_reg[3]/NET0131 ,
		\u2_chunk_cnt_reg[4]/NET0131 ,
		_w1243_
	);
	LUT3 #(
		.INIT('h01)
	) name509 (
		\u2_chunk_cnt_reg[5]/NET0131 ,
		\u2_chunk_cnt_reg[6]/NET0131 ,
		\u2_chunk_cnt_reg[7]/NET0131 ,
		_w1244_
	);
	LUT3 #(
		.INIT('h80)
	) name510 (
		_w1242_,
		_w1243_,
		_w1244_,
		_w1245_
	);
	LUT2 #(
		.INIT('h4)
	) name511 (
		\u1_next_start_reg/P0001 ,
		\u2_chunk_cnt_reg[8]/NET0131 ,
		_w1246_
	);
	LUT3 #(
		.INIT('hb0)
	) name512 (
		_w747_,
		_w748_,
		_w1246_,
		_w1247_
	);
	LUT2 #(
		.INIT('h1)
	) name513 (
		\u1_next_start_reg/P0001 ,
		\u2_chunk_cnt_reg[8]/NET0131 ,
		_w1248_
	);
	LUT3 #(
		.INIT('hb0)
	) name514 (
		_w747_,
		_w748_,
		_w1248_,
		_w1249_
	);
	LUT4 #(
		.INIT('h8a88)
	) name515 (
		\u0_u0_ch_chk_sz_r_reg[8]/P0001 ,
		\u1_next_start_reg/P0001 ,
		_w747_,
		_w748_,
		_w1250_
	);
	LUT4 #(
		.INIT('hffe4)
	) name516 (
		_w1245_,
		_w1247_,
		_w1249_,
		_w1250_,
		_w1251_
	);
	LUT3 #(
		.INIT('h40)
	) name517 (
		\u3_u1_slv_adr_reg[4]/NET0131 ,
		\u3_u1_slv_adr_reg[5]/P0001 ,
		\u3_u1_slv_we_reg/P0001 ,
		_w1252_
	);
	LUT2 #(
		.INIT('h2)
	) name518 (
		\u3_u1_slv_adr_reg[2]/NET0131 ,
		\u3_u1_slv_adr_reg[3]/P0001 ,
		_w1253_
	);
	LUT3 #(
		.INIT('h80)
	) name519 (
		_w1051_,
		_w1252_,
		_w1253_,
		_w1254_
	);
	LUT2 #(
		.INIT('h9)
	) name520 (
		\u2_state_reg[3]/NET0131 ,
		\u2_state_reg[4]/NET0131 ,
		_w1255_
	);
	LUT4 #(
		.INIT('h0080)
	) name521 (
		_w910_,
		_w1067_,
		_w1145_,
		_w1255_,
		_w1256_
	);
	LUT2 #(
		.INIT('h8)
	) name522 (
		\u2_mast0_drdy_r_reg/P0001 ,
		\u2_state_reg[5]/NET0131 ,
		_w1257_
	);
	LUT3 #(
		.INIT('h2a)
	) name523 (
		\u0_u0_ch_tot_sz_r_reg[0]/P0001 ,
		\u2_mast0_drdy_r_reg/P0001 ,
		\u2_state_reg[5]/NET0131 ,
		_w1258_
	);
	LUT3 #(
		.INIT('h10)
	) name524 (
		_w1254_,
		_w1256_,
		_w1258_,
		_w1259_
	);
	LUT3 #(
		.INIT('h53)
	) name525 (
		\u2_tsz_cnt_reg[0]/NET0131 ,
		\u3_u0_mast_dout_reg[0]/P0001 ,
		_w895_,
		_w1260_
	);
	LUT4 #(
		.INIT('h0054)
	) name526 (
		_w1254_,
		_w1256_,
		_w1257_,
		_w1260_,
		_w1261_
	);
	LUT3 #(
		.INIT('h20)
	) name527 (
		\u3_u1_slv_adr_reg[2]/NET0131 ,
		\u3_u1_slv_adr_reg[3]/P0001 ,
		\u3_u1_slv_dout_reg[0]/P0001 ,
		_w1262_
	);
	LUT3 #(
		.INIT('h80)
	) name528 (
		_w1051_,
		_w1252_,
		_w1262_,
		_w1263_
	);
	LUT3 #(
		.INIT('hfe)
	) name529 (
		_w1259_,
		_w1261_,
		_w1263_,
		_w1264_
	);
	LUT3 #(
		.INIT('h2a)
	) name530 (
		\u0_u0_ch_tot_sz_r_reg[1]/P0001 ,
		\u2_mast0_drdy_r_reg/P0001 ,
		\u2_state_reg[5]/NET0131 ,
		_w1265_
	);
	LUT3 #(
		.INIT('h10)
	) name531 (
		_w1254_,
		_w1256_,
		_w1265_,
		_w1266_
	);
	LUT3 #(
		.INIT('h53)
	) name532 (
		\u2_tsz_cnt_reg[1]/NET0131 ,
		\u3_u0_mast_dout_reg[1]/P0001 ,
		_w895_,
		_w1267_
	);
	LUT4 #(
		.INIT('h0054)
	) name533 (
		_w1254_,
		_w1256_,
		_w1257_,
		_w1267_,
		_w1268_
	);
	LUT3 #(
		.INIT('h20)
	) name534 (
		\u3_u1_slv_adr_reg[2]/NET0131 ,
		\u3_u1_slv_adr_reg[3]/P0001 ,
		\u3_u1_slv_dout_reg[1]/P0001 ,
		_w1269_
	);
	LUT3 #(
		.INIT('h80)
	) name535 (
		_w1051_,
		_w1252_,
		_w1269_,
		_w1270_
	);
	LUT3 #(
		.INIT('hfe)
	) name536 (
		_w1266_,
		_w1268_,
		_w1270_,
		_w1271_
	);
	LUT3 #(
		.INIT('h53)
	) name537 (
		\u2_tsz_cnt_reg[10]/NET0131 ,
		\u3_u0_mast_dout_reg[10]/P0001 ,
		_w895_,
		_w1272_
	);
	LUT4 #(
		.INIT('h0054)
	) name538 (
		_w1254_,
		_w1256_,
		_w1257_,
		_w1272_,
		_w1273_
	);
	LUT3 #(
		.INIT('h20)
	) name539 (
		\u3_u1_slv_adr_reg[2]/NET0131 ,
		\u3_u1_slv_adr_reg[3]/P0001 ,
		\u3_u1_slv_dout_reg[10]/P0001 ,
		_w1274_
	);
	LUT3 #(
		.INIT('h80)
	) name540 (
		_w1051_,
		_w1252_,
		_w1274_,
		_w1275_
	);
	LUT4 #(
		.INIT('h2aaa)
	) name541 (
		\u0_u0_ch_tot_sz_r_reg[10]/P0001 ,
		_w1051_,
		_w1252_,
		_w1253_,
		_w1276_
	);
	LUT4 #(
		.INIT('h0e0f)
	) name542 (
		_w1256_,
		_w1257_,
		_w1275_,
		_w1276_,
		_w1277_
	);
	LUT2 #(
		.INIT('hb)
	) name543 (
		_w1273_,
		_w1277_,
		_w1278_
	);
	LUT3 #(
		.INIT('h53)
	) name544 (
		\u2_tsz_cnt_reg[11]/NET0131 ,
		\u3_u0_mast_dout_reg[11]/P0001 ,
		_w895_,
		_w1279_
	);
	LUT4 #(
		.INIT('h0054)
	) name545 (
		_w1254_,
		_w1256_,
		_w1257_,
		_w1279_,
		_w1280_
	);
	LUT3 #(
		.INIT('h20)
	) name546 (
		\u3_u1_slv_adr_reg[2]/NET0131 ,
		\u3_u1_slv_adr_reg[3]/P0001 ,
		\u3_u1_slv_dout_reg[11]/P0001 ,
		_w1281_
	);
	LUT3 #(
		.INIT('h80)
	) name547 (
		_w1051_,
		_w1252_,
		_w1281_,
		_w1282_
	);
	LUT4 #(
		.INIT('h2aaa)
	) name548 (
		\u0_u0_ch_tot_sz_r_reg[11]/P0001 ,
		_w1051_,
		_w1252_,
		_w1253_,
		_w1283_
	);
	LUT4 #(
		.INIT('h0e0f)
	) name549 (
		_w1256_,
		_w1257_,
		_w1282_,
		_w1283_,
		_w1284_
	);
	LUT2 #(
		.INIT('hb)
	) name550 (
		_w1280_,
		_w1284_,
		_w1285_
	);
	LUT3 #(
		.INIT('h53)
	) name551 (
		\u2_tsz_cnt_reg[2]/NET0131 ,
		\u3_u0_mast_dout_reg[2]/P0001 ,
		_w895_,
		_w1286_
	);
	LUT4 #(
		.INIT('h0054)
	) name552 (
		_w1254_,
		_w1256_,
		_w1257_,
		_w1286_,
		_w1287_
	);
	LUT3 #(
		.INIT('h20)
	) name553 (
		\u3_u1_slv_adr_reg[2]/NET0131 ,
		\u3_u1_slv_adr_reg[3]/P0001 ,
		\u3_u1_slv_dout_reg[2]/P0001 ,
		_w1288_
	);
	LUT3 #(
		.INIT('h80)
	) name554 (
		_w1051_,
		_w1252_,
		_w1288_,
		_w1289_
	);
	LUT4 #(
		.INIT('h2aaa)
	) name555 (
		\u0_u0_ch_tot_sz_r_reg[2]/P0001 ,
		_w1051_,
		_w1252_,
		_w1253_,
		_w1290_
	);
	LUT4 #(
		.INIT('h0e0f)
	) name556 (
		_w1256_,
		_w1257_,
		_w1289_,
		_w1290_,
		_w1291_
	);
	LUT2 #(
		.INIT('hb)
	) name557 (
		_w1287_,
		_w1291_,
		_w1292_
	);
	LUT3 #(
		.INIT('h53)
	) name558 (
		\u2_tsz_cnt_reg[3]/NET0131 ,
		\u3_u0_mast_dout_reg[3]/P0001 ,
		_w895_,
		_w1293_
	);
	LUT4 #(
		.INIT('h0054)
	) name559 (
		_w1254_,
		_w1256_,
		_w1257_,
		_w1293_,
		_w1294_
	);
	LUT3 #(
		.INIT('h20)
	) name560 (
		\u3_u1_slv_adr_reg[2]/NET0131 ,
		\u3_u1_slv_adr_reg[3]/P0001 ,
		\u3_u1_slv_dout_reg[3]/P0001 ,
		_w1295_
	);
	LUT3 #(
		.INIT('h80)
	) name561 (
		_w1051_,
		_w1252_,
		_w1295_,
		_w1296_
	);
	LUT4 #(
		.INIT('h2aaa)
	) name562 (
		\u0_u0_ch_tot_sz_r_reg[3]/P0001 ,
		_w1051_,
		_w1252_,
		_w1253_,
		_w1297_
	);
	LUT4 #(
		.INIT('h0e0f)
	) name563 (
		_w1256_,
		_w1257_,
		_w1296_,
		_w1297_,
		_w1298_
	);
	LUT2 #(
		.INIT('hb)
	) name564 (
		_w1294_,
		_w1298_,
		_w1299_
	);
	LUT3 #(
		.INIT('h53)
	) name565 (
		\u2_tsz_cnt_reg[4]/NET0131 ,
		\u3_u0_mast_dout_reg[4]/P0001 ,
		_w895_,
		_w1300_
	);
	LUT4 #(
		.INIT('h0054)
	) name566 (
		_w1254_,
		_w1256_,
		_w1257_,
		_w1300_,
		_w1301_
	);
	LUT3 #(
		.INIT('h20)
	) name567 (
		\u3_u1_slv_adr_reg[2]/NET0131 ,
		\u3_u1_slv_adr_reg[3]/P0001 ,
		\u3_u1_slv_dout_reg[4]/P0001 ,
		_w1302_
	);
	LUT3 #(
		.INIT('h80)
	) name568 (
		_w1051_,
		_w1252_,
		_w1302_,
		_w1303_
	);
	LUT4 #(
		.INIT('h2aaa)
	) name569 (
		\u0_u0_ch_tot_sz_r_reg[4]/P0001 ,
		_w1051_,
		_w1252_,
		_w1253_,
		_w1304_
	);
	LUT4 #(
		.INIT('h0e0f)
	) name570 (
		_w1256_,
		_w1257_,
		_w1303_,
		_w1304_,
		_w1305_
	);
	LUT2 #(
		.INIT('hb)
	) name571 (
		_w1301_,
		_w1305_,
		_w1306_
	);
	LUT3 #(
		.INIT('h53)
	) name572 (
		\u2_tsz_cnt_reg[5]/NET0131 ,
		\u3_u0_mast_dout_reg[5]/P0001 ,
		_w895_,
		_w1307_
	);
	LUT4 #(
		.INIT('h0054)
	) name573 (
		_w1254_,
		_w1256_,
		_w1257_,
		_w1307_,
		_w1308_
	);
	LUT3 #(
		.INIT('h20)
	) name574 (
		\u3_u1_slv_adr_reg[2]/NET0131 ,
		\u3_u1_slv_adr_reg[3]/P0001 ,
		\u3_u1_slv_dout_reg[5]/P0001 ,
		_w1309_
	);
	LUT3 #(
		.INIT('h80)
	) name575 (
		_w1051_,
		_w1252_,
		_w1309_,
		_w1310_
	);
	LUT4 #(
		.INIT('h2aaa)
	) name576 (
		\u0_u0_ch_tot_sz_r_reg[5]/P0001 ,
		_w1051_,
		_w1252_,
		_w1253_,
		_w1311_
	);
	LUT4 #(
		.INIT('h0e0f)
	) name577 (
		_w1256_,
		_w1257_,
		_w1310_,
		_w1311_,
		_w1312_
	);
	LUT2 #(
		.INIT('hb)
	) name578 (
		_w1308_,
		_w1312_,
		_w1313_
	);
	LUT3 #(
		.INIT('h53)
	) name579 (
		\u2_tsz_cnt_reg[6]/NET0131 ,
		\u3_u0_mast_dout_reg[6]/P0001 ,
		_w895_,
		_w1314_
	);
	LUT4 #(
		.INIT('h0054)
	) name580 (
		_w1254_,
		_w1256_,
		_w1257_,
		_w1314_,
		_w1315_
	);
	LUT3 #(
		.INIT('h20)
	) name581 (
		\u3_u1_slv_adr_reg[2]/NET0131 ,
		\u3_u1_slv_adr_reg[3]/P0001 ,
		\u3_u1_slv_dout_reg[6]/P0001 ,
		_w1316_
	);
	LUT3 #(
		.INIT('h80)
	) name582 (
		_w1051_,
		_w1252_,
		_w1316_,
		_w1317_
	);
	LUT4 #(
		.INIT('h2aaa)
	) name583 (
		\u0_u0_ch_tot_sz_r_reg[6]/P0001 ,
		_w1051_,
		_w1252_,
		_w1253_,
		_w1318_
	);
	LUT4 #(
		.INIT('h0e0f)
	) name584 (
		_w1256_,
		_w1257_,
		_w1317_,
		_w1318_,
		_w1319_
	);
	LUT2 #(
		.INIT('hb)
	) name585 (
		_w1315_,
		_w1319_,
		_w1320_
	);
	LUT3 #(
		.INIT('h53)
	) name586 (
		\u2_tsz_cnt_reg[7]/NET0131 ,
		\u3_u0_mast_dout_reg[7]/P0001 ,
		_w895_,
		_w1321_
	);
	LUT4 #(
		.INIT('h0054)
	) name587 (
		_w1254_,
		_w1256_,
		_w1257_,
		_w1321_,
		_w1322_
	);
	LUT3 #(
		.INIT('h20)
	) name588 (
		\u3_u1_slv_adr_reg[2]/NET0131 ,
		\u3_u1_slv_adr_reg[3]/P0001 ,
		\u3_u1_slv_dout_reg[7]/P0001 ,
		_w1323_
	);
	LUT3 #(
		.INIT('h80)
	) name589 (
		_w1051_,
		_w1252_,
		_w1323_,
		_w1324_
	);
	LUT4 #(
		.INIT('h2aaa)
	) name590 (
		\u0_u0_ch_tot_sz_r_reg[7]/P0001 ,
		_w1051_,
		_w1252_,
		_w1253_,
		_w1325_
	);
	LUT4 #(
		.INIT('h0e0f)
	) name591 (
		_w1256_,
		_w1257_,
		_w1324_,
		_w1325_,
		_w1326_
	);
	LUT2 #(
		.INIT('hb)
	) name592 (
		_w1322_,
		_w1326_,
		_w1327_
	);
	LUT3 #(
		.INIT('h53)
	) name593 (
		\u2_tsz_cnt_reg[8]/NET0131 ,
		\u3_u0_mast_dout_reg[8]/P0001 ,
		_w895_,
		_w1328_
	);
	LUT4 #(
		.INIT('h0054)
	) name594 (
		_w1254_,
		_w1256_,
		_w1257_,
		_w1328_,
		_w1329_
	);
	LUT3 #(
		.INIT('h20)
	) name595 (
		\u3_u1_slv_adr_reg[2]/NET0131 ,
		\u3_u1_slv_adr_reg[3]/P0001 ,
		\u3_u1_slv_dout_reg[8]/P0001 ,
		_w1330_
	);
	LUT3 #(
		.INIT('h80)
	) name596 (
		_w1051_,
		_w1252_,
		_w1330_,
		_w1331_
	);
	LUT4 #(
		.INIT('h2aaa)
	) name597 (
		\u0_u0_ch_tot_sz_r_reg[8]/P0001 ,
		_w1051_,
		_w1252_,
		_w1253_,
		_w1332_
	);
	LUT4 #(
		.INIT('h0e0f)
	) name598 (
		_w1256_,
		_w1257_,
		_w1331_,
		_w1332_,
		_w1333_
	);
	LUT2 #(
		.INIT('hb)
	) name599 (
		_w1329_,
		_w1333_,
		_w1334_
	);
	LUT3 #(
		.INIT('h53)
	) name600 (
		\u2_tsz_cnt_reg[9]/NET0131 ,
		\u3_u0_mast_dout_reg[9]/P0001 ,
		_w895_,
		_w1335_
	);
	LUT4 #(
		.INIT('h0054)
	) name601 (
		_w1254_,
		_w1256_,
		_w1257_,
		_w1335_,
		_w1336_
	);
	LUT3 #(
		.INIT('h20)
	) name602 (
		\u3_u1_slv_adr_reg[2]/NET0131 ,
		\u3_u1_slv_adr_reg[3]/P0001 ,
		\u3_u1_slv_dout_reg[9]/P0001 ,
		_w1337_
	);
	LUT3 #(
		.INIT('h80)
	) name603 (
		_w1051_,
		_w1252_,
		_w1337_,
		_w1338_
	);
	LUT4 #(
		.INIT('h2aaa)
	) name604 (
		\u0_u0_ch_tot_sz_r_reg[9]/P0001 ,
		_w1051_,
		_w1252_,
		_w1253_,
		_w1339_
	);
	LUT4 #(
		.INIT('h0e0f)
	) name605 (
		_w1256_,
		_w1257_,
		_w1338_,
		_w1339_,
		_w1340_
	);
	LUT2 #(
		.INIT('hb)
	) name606 (
		_w1336_,
		_w1340_,
		_w1341_
	);
	LUT4 #(
		.INIT('h8a88)
	) name607 (
		\u0_u0_ch_chk_sz_r_reg[0]/P0001 ,
		\u1_next_start_reg/P0001 ,
		_w747_,
		_w748_,
		_w1342_
	);
	LUT3 #(
		.INIT('h63)
	) name608 (
		\u2_chunk_cnt_is_0_r_reg/P0001 ,
		\u2_chunk_cnt_reg[0]/NET0131 ,
		\u2_chunk_dec_reg/P0001 ,
		_w1343_
	);
	LUT4 #(
		.INIT('h0045)
	) name609 (
		\u1_next_start_reg/P0001 ,
		_w747_,
		_w748_,
		_w1343_,
		_w1344_
	);
	LUT2 #(
		.INIT('he)
	) name610 (
		_w1342_,
		_w1344_,
		_w1345_
	);
	LUT4 #(
		.INIT('h8a88)
	) name611 (
		\u0_u0_ch_chk_sz_r_reg[1]/P0001 ,
		\u1_next_start_reg/P0001 ,
		_w747_,
		_w748_,
		_w1346_
	);
	LUT4 #(
		.INIT('h1e0f)
	) name612 (
		\u2_chunk_cnt_is_0_r_reg/P0001 ,
		\u2_chunk_cnt_reg[0]/NET0131 ,
		\u2_chunk_cnt_reg[1]/NET0131 ,
		\u2_chunk_dec_reg/P0001 ,
		_w1347_
	);
	LUT4 #(
		.INIT('h0045)
	) name613 (
		\u1_next_start_reg/P0001 ,
		_w747_,
		_w748_,
		_w1347_,
		_w1348_
	);
	LUT2 #(
		.INIT('he)
	) name614 (
		_w1346_,
		_w1348_,
		_w1349_
	);
	LUT2 #(
		.INIT('h9)
	) name615 (
		\u2_chunk_cnt_reg[2]/NET0131 ,
		_w1242_,
		_w1350_
	);
	LUT3 #(
		.INIT('h2e)
	) name616 (
		\u0_u0_ch_chk_sz_r_reg[2]/P0001 ,
		_w1075_,
		_w1350_,
		_w1351_
	);
	LUT3 #(
		.INIT('h63)
	) name617 (
		\u2_chunk_cnt_reg[2]/NET0131 ,
		\u2_chunk_cnt_reg[3]/NET0131 ,
		_w1242_,
		_w1352_
	);
	LUT3 #(
		.INIT('h2e)
	) name618 (
		\u0_u0_ch_chk_sz_r_reg[3]/P0001 ,
		_w1075_,
		_w1352_,
		_w1353_
	);
	LUT4 #(
		.INIT('h1e0f)
	) name619 (
		\u2_chunk_cnt_reg[2]/NET0131 ,
		\u2_chunk_cnt_reg[3]/NET0131 ,
		\u2_chunk_cnt_reg[4]/NET0131 ,
		_w1242_,
		_w1354_
	);
	LUT3 #(
		.INIT('h2e)
	) name620 (
		\u0_u0_ch_chk_sz_r_reg[4]/P0001 ,
		_w1075_,
		_w1354_,
		_w1355_
	);
	LUT3 #(
		.INIT('h40)
	) name621 (
		\u2_chunk_cnt_reg[5]/NET0131 ,
		_w1242_,
		_w1243_,
		_w1356_
	);
	LUT3 #(
		.INIT('h95)
	) name622 (
		\u2_chunk_cnt_reg[5]/NET0131 ,
		_w1242_,
		_w1243_,
		_w1357_
	);
	LUT3 #(
		.INIT('h2e)
	) name623 (
		\u0_u0_ch_chk_sz_r_reg[5]/P0001 ,
		_w1075_,
		_w1357_,
		_w1358_
	);
	LUT4 #(
		.INIT('h8a88)
	) name624 (
		\u0_u0_ch_chk_sz_r_reg[6]/P0001 ,
		\u1_next_start_reg/P0001 ,
		_w747_,
		_w748_,
		_w1359_
	);
	LUT2 #(
		.INIT('h4)
	) name625 (
		\u1_next_start_reg/P0001 ,
		\u2_chunk_cnt_reg[6]/NET0131 ,
		_w1360_
	);
	LUT3 #(
		.INIT('hb0)
	) name626 (
		_w747_,
		_w748_,
		_w1360_,
		_w1361_
	);
	LUT2 #(
		.INIT('h1)
	) name627 (
		\u1_next_start_reg/P0001 ,
		\u2_chunk_cnt_reg[6]/NET0131 ,
		_w1362_
	);
	LUT3 #(
		.INIT('hb0)
	) name628 (
		_w747_,
		_w748_,
		_w1362_,
		_w1363_
	);
	LUT4 #(
		.INIT('hfedc)
	) name629 (
		_w1356_,
		_w1359_,
		_w1361_,
		_w1363_,
		_w1364_
	);
	LUT2 #(
		.INIT('h1)
	) name630 (
		\u2_chunk_cnt_reg[5]/NET0131 ,
		\u2_chunk_cnt_reg[6]/NET0131 ,
		_w1365_
	);
	LUT4 #(
		.INIT('h2aaa)
	) name631 (
		\u2_chunk_cnt_reg[7]/NET0131 ,
		_w1242_,
		_w1243_,
		_w1365_,
		_w1366_
	);
	LUT4 #(
		.INIT('heee2)
	) name632 (
		\u0_u0_ch_chk_sz_r_reg[7]/P0001 ,
		_w1075_,
		_w1245_,
		_w1366_,
		_w1367_
	);
	LUT3 #(
		.INIT('h01)
	) name633 (
		\u0_u0_ch_chk_sz_r_reg[6]/P0001 ,
		\u0_u0_ch_chk_sz_r_reg[7]/P0001 ,
		\u0_u0_ch_chk_sz_r_reg[8]/P0001 ,
		_w1368_
	);
	LUT2 #(
		.INIT('h1)
	) name634 (
		\u0_u0_ch_chk_sz_r_reg[0]/P0001 ,
		\u0_u0_ch_chk_sz_r_reg[1]/P0001 ,
		_w1369_
	);
	LUT4 #(
		.INIT('h0001)
	) name635 (
		\u0_u0_ch_chk_sz_r_reg[2]/P0001 ,
		\u0_u0_ch_chk_sz_r_reg[3]/P0001 ,
		\u0_u0_ch_chk_sz_r_reg[4]/P0001 ,
		\u0_u0_ch_chk_sz_r_reg[5]/P0001 ,
		_w1370_
	);
	LUT3 #(
		.INIT('h80)
	) name636 (
		_w1368_,
		_w1369_,
		_w1370_,
		_w1371_
	);
	LUT4 #(
		.INIT('h8000)
	) name637 (
		\u2_adr0_cnt_reg[0]/P0001 ,
		\u2_adr0_cnt_reg[1]/P0001 ,
		\u2_adr0_cnt_reg[2]/P0001 ,
		\u2_adr0_cnt_reg[3]/P0001 ,
		_w1372_
	);
	LUT3 #(
		.INIT('h80)
	) name638 (
		\u2_adr0_cnt_reg[4]/P0001 ,
		\u2_adr0_cnt_reg[5]/P0001 ,
		\u2_adr0_cnt_reg[6]/P0001 ,
		_w1373_
	);
	LUT3 #(
		.INIT('h80)
	) name639 (
		\u2_adr0_cnt_reg[7]/P0001 ,
		\u2_adr0_cnt_reg[8]/P0001 ,
		\u2_adr0_cnt_reg[9]/P0001 ,
		_w1374_
	);
	LUT3 #(
		.INIT('h80)
	) name640 (
		_w1372_,
		_w1373_,
		_w1374_,
		_w1375_
	);
	LUT2 #(
		.INIT('h8)
	) name641 (
		\u2_adr0_cnt_reg[10]/P0001 ,
		\u2_adr0_cnt_reg[11]/P0001 ,
		_w1376_
	);
	LUT4 #(
		.INIT('h8000)
	) name642 (
		_w1372_,
		_w1373_,
		_w1374_,
		_w1376_,
		_w1377_
	);
	LUT3 #(
		.INIT('h80)
	) name643 (
		\u2_adr0_cnt_reg[10]/P0001 ,
		\u2_adr0_cnt_reg[11]/P0001 ,
		\u2_adr0_cnt_reg[12]/P0001 ,
		_w1378_
	);
	LUT4 #(
		.INIT('h8000)
	) name644 (
		_w1372_,
		_w1373_,
		_w1374_,
		_w1378_,
		_w1379_
	);
	LUT3 #(
		.INIT('h0e)
	) name645 (
		\u2_adr0_cnt_reg[12]/P0001 ,
		_w1377_,
		_w1379_,
		_w1380_
	);
	LUT4 #(
		.INIT('h8000)
	) name646 (
		\u2_adr1_cnt_reg[0]/P0001 ,
		\u2_adr1_cnt_reg[1]/P0001 ,
		\u2_adr1_cnt_reg[2]/P0001 ,
		\u2_adr1_cnt_reg[3]/P0001 ,
		_w1381_
	);
	LUT3 #(
		.INIT('h80)
	) name647 (
		\u2_adr1_cnt_reg[4]/P0001 ,
		\u2_adr1_cnt_reg[5]/P0001 ,
		\u2_adr1_cnt_reg[6]/P0001 ,
		_w1382_
	);
	LUT3 #(
		.INIT('h80)
	) name648 (
		\u2_adr1_cnt_reg[7]/P0001 ,
		\u2_adr1_cnt_reg[8]/P0001 ,
		\u2_adr1_cnt_reg[9]/P0001 ,
		_w1383_
	);
	LUT3 #(
		.INIT('h80)
	) name649 (
		_w1381_,
		_w1382_,
		_w1383_,
		_w1384_
	);
	LUT2 #(
		.INIT('h8)
	) name650 (
		\u2_adr1_cnt_reg[10]/P0001 ,
		\u2_adr1_cnt_reg[11]/P0001 ,
		_w1385_
	);
	LUT4 #(
		.INIT('h8000)
	) name651 (
		_w1381_,
		_w1382_,
		_w1383_,
		_w1385_,
		_w1386_
	);
	LUT3 #(
		.INIT('h80)
	) name652 (
		\u2_adr1_cnt_reg[10]/P0001 ,
		\u2_adr1_cnt_reg[11]/P0001 ,
		\u2_adr1_cnt_reg[12]/P0001 ,
		_w1387_
	);
	LUT4 #(
		.INIT('h8000)
	) name653 (
		_w1381_,
		_w1382_,
		_w1383_,
		_w1387_,
		_w1388_
	);
	LUT3 #(
		.INIT('h0e)
	) name654 (
		\u2_adr1_cnt_reg[12]/P0001 ,
		_w1386_,
		_w1388_,
		_w1389_
	);
	LUT3 #(
		.INIT('h07)
	) name655 (
		\u3_u1_slv_adr_reg[2]/NET0131 ,
		\u3_u1_slv_adr_reg[3]/P0001 ,
		\u3_u1_slv_adr_reg[4]/NET0131 ,
		_w1390_
	);
	LUT3 #(
		.INIT('h04)
	) name656 (
		\u3_u1_slv_adr_reg[5]/P0001 ,
		_w1051_,
		_w1390_,
		_w1391_
	);
	LUT2 #(
		.INIT('h8)
	) name657 (
		\u3_u1_slv_adr_reg[3]/P0001 ,
		\u3_u1_slv_adr_reg[4]/NET0131 ,
		_w1392_
	);
	LUT3 #(
		.INIT('h57)
	) name658 (
		_w1051_,
		_w1097_,
		_w1392_,
		_w1393_
	);
	LUT2 #(
		.INIT('h4)
	) name659 (
		_w1391_,
		_w1393_,
		_w1394_
	);
	LUT2 #(
		.INIT('h1)
	) name660 (
		\u3_u1_slv_adr_reg[2]/NET0131 ,
		\u3_u1_slv_adr_reg[5]/P0001 ,
		_w1395_
	);
	LUT3 #(
		.INIT('h84)
	) name661 (
		\u3_u1_slv_adr_reg[3]/P0001 ,
		_w1051_,
		_w1395_,
		_w1396_
	);
	LUT4 #(
		.INIT('h5400)
	) name662 (
		\u3_u1_slv_adr_reg[2]/NET0131 ,
		\u3_u1_slv_adr_reg[3]/P0001 ,
		\u3_u1_slv_adr_reg[4]/NET0131 ,
		\u3_u1_slv_adr_reg[5]/P0001 ,
		_w1397_
	);
	LUT3 #(
		.INIT('h80)
	) name663 (
		\u0_u0_ch_adr1_r_reg[7]/P0001 ,
		_w1051_,
		_w1397_,
		_w1398_
	);
	LUT4 #(
		.INIT('h4000)
	) name664 (
		_w1391_,
		_w1393_,
		_w1396_,
		_w1398_,
		_w1399_
	);
	LUT4 #(
		.INIT('ha800)
	) name665 (
		\u3_u1_slv_adr_reg[2]/NET0131 ,
		\u3_u1_slv_adr_reg[3]/P0001 ,
		\u3_u1_slv_adr_reg[4]/NET0131 ,
		\u3_u1_slv_adr_reg[5]/P0001 ,
		_w1400_
	);
	LUT2 #(
		.INIT('h8)
	) name666 (
		_w1051_,
		_w1400_,
		_w1401_
	);
	LUT3 #(
		.INIT('h40)
	) name667 (
		_w1391_,
		_w1393_,
		_w1401_,
		_w1402_
	);
	LUT2 #(
		.INIT('h1)
	) name668 (
		_w1399_,
		_w1402_,
		_w1403_
	);
	LUT3 #(
		.INIT('he0)
	) name669 (
		\u3_u1_slv_adr_reg[3]/P0001 ,
		\u3_u1_slv_adr_reg[4]/NET0131 ,
		\u3_u1_slv_adr_reg[5]/P0001 ,
		_w1404_
	);
	LUT2 #(
		.INIT('h6)
	) name670 (
		\u3_u1_slv_adr_reg[2]/NET0131 ,
		\u3_u1_slv_adr_reg[5]/P0001 ,
		_w1405_
	);
	LUT3 #(
		.INIT('h02)
	) name671 (
		_w1051_,
		_w1404_,
		_w1405_,
		_w1406_
	);
	LUT2 #(
		.INIT('h8)
	) name672 (
		_w1396_,
		_w1406_,
		_w1407_
	);
	LUT4 #(
		.INIT('hb000)
	) name673 (
		_w1391_,
		_w1393_,
		_w1396_,
		_w1406_,
		_w1408_
	);
	LUT3 #(
		.INIT('h75)
	) name674 (
		_w1051_,
		_w1404_,
		_w1405_,
		_w1409_
	);
	LUT2 #(
		.INIT('h8)
	) name675 (
		_w1396_,
		_w1409_,
		_w1410_
	);
	LUT4 #(
		.INIT('h4000)
	) name676 (
		_w1391_,
		_w1393_,
		_w1396_,
		_w1409_,
		_w1411_
	);
	LUT4 #(
		.INIT('h153f)
	) name677 (
		\u0_int_maska_r_reg[9]/NET0131 ,
		\u0_u0_ch_tot_sz_r_reg[9]/P0001 ,
		_w1408_,
		_w1411_,
		_w1412_
	);
	LUT4 #(
		.INIT('h4000)
	) name678 (
		_w1391_,
		_w1393_,
		_w1396_,
		_w1406_,
		_w1413_
	);
	LUT3 #(
		.INIT('h80)
	) name679 (
		\u0_u0_ch_adr0_r_reg[7]/P0001 ,
		_w1051_,
		_w1397_,
		_w1414_
	);
	LUT4 #(
		.INIT('h0400)
	) name680 (
		_w1391_,
		_w1393_,
		_w1396_,
		_w1414_,
		_w1415_
	);
	LUT3 #(
		.INIT('h07)
	) name681 (
		\u0_int_maskb_r_reg[9]/NET0131 ,
		_w1413_,
		_w1415_,
		_w1416_
	);
	LUT3 #(
		.INIT('h7f)
	) name682 (
		_w1403_,
		_w1412_,
		_w1416_,
		_w1417_
	);
	LUT4 #(
		.INIT('hb000)
	) name683 (
		_w1391_,
		_w1393_,
		_w1396_,
		_w1409_,
		_w1418_
	);
	LUT3 #(
		.INIT('h13)
	) name684 (
		\u0_u0_ch_err_reg/NET0131 ,
		_w1402_,
		_w1418_,
		_w1419_
	);
	LUT3 #(
		.INIT('h80)
	) name685 (
		\u0_u0_ch_adr1_r_reg[10]/P0001 ,
		_w1051_,
		_w1397_,
		_w1420_
	);
	LUT4 #(
		.INIT('h4000)
	) name686 (
		_w1391_,
		_w1393_,
		_w1396_,
		_w1420_,
		_w1421_
	);
	LUT3 #(
		.INIT('h80)
	) name687 (
		\u0_u0_ch_adr0_r_reg[10]/P0001 ,
		_w1051_,
		_w1397_,
		_w1422_
	);
	LUT4 #(
		.INIT('h0400)
	) name688 (
		_w1391_,
		_w1393_,
		_w1396_,
		_w1422_,
		_w1423_
	);
	LUT2 #(
		.INIT('h1)
	) name689 (
		_w1421_,
		_w1423_,
		_w1424_
	);
	LUT4 #(
		.INIT('h135f)
	) name690 (
		\u0_int_maska_r_reg[12]/NET0131 ,
		\u0_int_maskb_r_reg[12]/NET0131 ,
		_w1411_,
		_w1413_,
		_w1425_
	);
	LUT3 #(
		.INIT('h7f)
	) name691 (
		_w1419_,
		_w1424_,
		_w1425_,
		_w1426_
	);
	LUT3 #(
		.INIT('h80)
	) name692 (
		\u0_u0_ch_adr0_r_reg[11]/P0001 ,
		_w1051_,
		_w1397_,
		_w1427_
	);
	LUT4 #(
		.INIT('h0400)
	) name693 (
		_w1391_,
		_w1393_,
		_w1396_,
		_w1427_,
		_w1428_
	);
	LUT2 #(
		.INIT('h1)
	) name694 (
		_w1402_,
		_w1428_,
		_w1429_
	);
	LUT4 #(
		.INIT('h53ff)
	) name695 (
		\u0_int_maska_r_reg[13]/NET0131 ,
		\u0_u0_ch_csr_r2_reg[0]/NET0131 ,
		_w1394_,
		_w1410_,
		_w1430_
	);
	LUT3 #(
		.INIT('h80)
	) name696 (
		\u0_u0_ch_adr1_r_reg[11]/P0001 ,
		_w1051_,
		_w1397_,
		_w1431_
	);
	LUT4 #(
		.INIT('h4000)
	) name697 (
		_w1391_,
		_w1393_,
		_w1396_,
		_w1431_,
		_w1432_
	);
	LUT3 #(
		.INIT('h07)
	) name698 (
		\u0_int_maskb_r_reg[13]/NET0131 ,
		_w1413_,
		_w1432_,
		_w1433_
	);
	LUT3 #(
		.INIT('h7f)
	) name699 (
		_w1429_,
		_w1430_,
		_w1433_,
		_w1434_
	);
	LUT3 #(
		.INIT('h80)
	) name700 (
		\u0_u0_ch_adr0_r_reg[12]/P0001 ,
		_w1051_,
		_w1397_,
		_w1435_
	);
	LUT4 #(
		.INIT('h0400)
	) name701 (
		_w1391_,
		_w1393_,
		_w1396_,
		_w1435_,
		_w1436_
	);
	LUT2 #(
		.INIT('h1)
	) name702 (
		_w1402_,
		_w1436_,
		_w1437_
	);
	LUT4 #(
		.INIT('h53ff)
	) name703 (
		\u0_int_maska_r_reg[14]/NET0131 ,
		\u0_u0_ch_csr_r2_reg[1]/NET0131 ,
		_w1394_,
		_w1410_,
		_w1438_
	);
	LUT3 #(
		.INIT('h80)
	) name704 (
		\u0_u0_ch_adr1_r_reg[12]/P0001 ,
		_w1051_,
		_w1397_,
		_w1439_
	);
	LUT4 #(
		.INIT('h4000)
	) name705 (
		_w1391_,
		_w1393_,
		_w1396_,
		_w1439_,
		_w1440_
	);
	LUT3 #(
		.INIT('h07)
	) name706 (
		\u0_int_maskb_r_reg[14]/NET0131 ,
		_w1413_,
		_w1440_,
		_w1441_
	);
	LUT3 #(
		.INIT('h7f)
	) name707 (
		_w1437_,
		_w1438_,
		_w1441_,
		_w1442_
	);
	LUT3 #(
		.INIT('h80)
	) name708 (
		\u0_u0_ch_adr0_r_reg[21]/P0001 ,
		_w1051_,
		_w1397_,
		_w1443_
	);
	LUT4 #(
		.INIT('h0400)
	) name709 (
		_w1391_,
		_w1393_,
		_w1396_,
		_w1443_,
		_w1444_
	);
	LUT2 #(
		.INIT('h1)
	) name710 (
		_w1402_,
		_w1444_,
		_w1445_
	);
	LUT3 #(
		.INIT('h80)
	) name711 (
		\u0_u0_ch_adr1_r_reg[21]/P0001 ,
		_w1051_,
		_w1397_,
		_w1446_
	);
	LUT4 #(
		.INIT('h4000)
	) name712 (
		_w1391_,
		_w1393_,
		_w1396_,
		_w1446_,
		_w1447_
	);
	LUT3 #(
		.INIT('h07)
	) name713 (
		\u0_int_maskb_r_reg[23]/NET0131 ,
		_w1413_,
		_w1447_,
		_w1448_
	);
	LUT4 #(
		.INIT('h153f)
	) name714 (
		\u0_int_maska_r_reg[23]/NET0131 ,
		\u0_u0_ch_chk_sz_r_reg[7]/P0001 ,
		_w1408_,
		_w1411_,
		_w1449_
	);
	LUT3 #(
		.INIT('h7f)
	) name715 (
		_w1445_,
		_w1448_,
		_w1449_,
		_w1450_
	);
	LUT3 #(
		.INIT('h80)
	) name716 (
		\u0_u0_ch_adr0_r_reg[22]/P0001 ,
		_w1051_,
		_w1397_,
		_w1451_
	);
	LUT4 #(
		.INIT('h0400)
	) name717 (
		_w1391_,
		_w1393_,
		_w1396_,
		_w1451_,
		_w1452_
	);
	LUT2 #(
		.INIT('h1)
	) name718 (
		_w1402_,
		_w1452_,
		_w1453_
	);
	LUT3 #(
		.INIT('h80)
	) name719 (
		\u0_u0_ch_adr1_r_reg[22]/P0001 ,
		_w1051_,
		_w1397_,
		_w1454_
	);
	LUT4 #(
		.INIT('h4000)
	) name720 (
		_w1391_,
		_w1393_,
		_w1396_,
		_w1454_,
		_w1455_
	);
	LUT3 #(
		.INIT('h07)
	) name721 (
		\u0_int_maskb_r_reg[24]/NET0131 ,
		_w1413_,
		_w1455_,
		_w1456_
	);
	LUT4 #(
		.INIT('h153f)
	) name722 (
		\u0_int_maska_r_reg[24]/NET0131 ,
		\u0_u0_ch_chk_sz_r_reg[8]/P0001 ,
		_w1408_,
		_w1411_,
		_w1457_
	);
	LUT3 #(
		.INIT('h7f)
	) name723 (
		_w1453_,
		_w1456_,
		_w1457_,
		_w1458_
	);
	LUT3 #(
		.INIT('h80)
	) name724 (
		\u0_u0_ch_adr0_r_reg[23]/P0001 ,
		_w1051_,
		_w1397_,
		_w1459_
	);
	LUT4 #(
		.INIT('h0400)
	) name725 (
		_w1391_,
		_w1393_,
		_w1396_,
		_w1459_,
		_w1460_
	);
	LUT2 #(
		.INIT('h1)
	) name726 (
		_w1402_,
		_w1460_,
		_w1461_
	);
	LUT4 #(
		.INIT('h153f)
	) name727 (
		\u0_int_maska_r_reg[25]/NET0131 ,
		\u0_u0_ch_chk_sz_r_reg[9]/P0001 ,
		_w1408_,
		_w1411_,
		_w1462_
	);
	LUT3 #(
		.INIT('h80)
	) name728 (
		\u0_u0_ch_adr1_r_reg[23]/P0001 ,
		_w1051_,
		_w1397_,
		_w1463_
	);
	LUT4 #(
		.INIT('h4000)
	) name729 (
		_w1391_,
		_w1393_,
		_w1396_,
		_w1463_,
		_w1464_
	);
	LUT3 #(
		.INIT('h07)
	) name730 (
		\u0_int_maskb_r_reg[25]/NET0131 ,
		_w1413_,
		_w1464_,
		_w1465_
	);
	LUT3 #(
		.INIT('h7f)
	) name731 (
		_w1461_,
		_w1462_,
		_w1465_,
		_w1466_
	);
	LUT3 #(
		.INIT('h80)
	) name732 (
		\u0_u0_ch_adr0_r_reg[24]/P0001 ,
		_w1051_,
		_w1397_,
		_w1467_
	);
	LUT4 #(
		.INIT('h0400)
	) name733 (
		_w1391_,
		_w1393_,
		_w1396_,
		_w1467_,
		_w1468_
	);
	LUT2 #(
		.INIT('h1)
	) name734 (
		_w1402_,
		_w1468_,
		_w1469_
	);
	LUT4 #(
		.INIT('h153f)
	) name735 (
		\u0_int_maska_r_reg[26]/NET0131 ,
		\u0_u0_ch_chk_sz_r_reg[10]/P0001 ,
		_w1408_,
		_w1411_,
		_w1470_
	);
	LUT3 #(
		.INIT('h80)
	) name736 (
		\u0_u0_ch_adr1_r_reg[24]/P0001 ,
		_w1051_,
		_w1397_,
		_w1471_
	);
	LUT4 #(
		.INIT('h4000)
	) name737 (
		_w1391_,
		_w1393_,
		_w1396_,
		_w1471_,
		_w1472_
	);
	LUT3 #(
		.INIT('h07)
	) name738 (
		\u0_int_maskb_r_reg[26]/NET0131 ,
		_w1413_,
		_w1472_,
		_w1473_
	);
	LUT3 #(
		.INIT('h7f)
	) name739 (
		_w1469_,
		_w1470_,
		_w1473_,
		_w1474_
	);
	LUT3 #(
		.INIT('h80)
	) name740 (
		\u0_u0_ch_adr0_r_reg[0]/P0001 ,
		_w1051_,
		_w1397_,
		_w1475_
	);
	LUT4 #(
		.INIT('h0400)
	) name741 (
		_w1391_,
		_w1393_,
		_w1396_,
		_w1475_,
		_w1476_
	);
	LUT3 #(
		.INIT('h80)
	) name742 (
		\u0_u0_ch_adr1_r_reg[0]/P0001 ,
		_w1051_,
		_w1397_,
		_w1477_
	);
	LUT4 #(
		.INIT('h4000)
	) name743 (
		_w1391_,
		_w1393_,
		_w1396_,
		_w1477_,
		_w1478_
	);
	LUT2 #(
		.INIT('h1)
	) name744 (
		_w1476_,
		_w1478_,
		_w1479_
	);
	LUT4 #(
		.INIT('h53ff)
	) name745 (
		\u0_int_maska_r_reg[2]/NET0131 ,
		\u0_u0_ch_csr_r_reg[2]/NET0131 ,
		_w1394_,
		_w1410_,
		_w1480_
	);
	LUT4 #(
		.INIT('h53ff)
	) name746 (
		\u0_int_maskb_r_reg[2]/NET0131 ,
		\u0_u0_ch_tot_sz_r_reg[2]/P0001 ,
		_w1394_,
		_w1407_,
		_w1481_
	);
	LUT3 #(
		.INIT('h7f)
	) name747 (
		_w1479_,
		_w1480_,
		_w1481_,
		_w1482_
	);
	LUT3 #(
		.INIT('h80)
	) name748 (
		\u0_u0_ch_adr0_r_reg[1]/P0001 ,
		_w1051_,
		_w1397_,
		_w1483_
	);
	LUT4 #(
		.INIT('h0400)
	) name749 (
		_w1391_,
		_w1393_,
		_w1396_,
		_w1483_,
		_w1484_
	);
	LUT3 #(
		.INIT('h80)
	) name750 (
		\u0_u0_ch_adr1_r_reg[1]/P0001 ,
		_w1051_,
		_w1397_,
		_w1485_
	);
	LUT4 #(
		.INIT('h4000)
	) name751 (
		_w1391_,
		_w1393_,
		_w1396_,
		_w1485_,
		_w1486_
	);
	LUT2 #(
		.INIT('h1)
	) name752 (
		_w1484_,
		_w1486_,
		_w1487_
	);
	LUT4 #(
		.INIT('h53ff)
	) name753 (
		\u0_int_maska_r_reg[3]/NET0131 ,
		\u0_u0_ch_csr_r_reg[3]/NET0131 ,
		_w1394_,
		_w1410_,
		_w1488_
	);
	LUT4 #(
		.INIT('h53ff)
	) name754 (
		\u0_int_maskb_r_reg[3]/NET0131 ,
		\u0_u0_ch_tot_sz_r_reg[3]/P0001 ,
		_w1394_,
		_w1407_,
		_w1489_
	);
	LUT3 #(
		.INIT('h7f)
	) name755 (
		_w1487_,
		_w1488_,
		_w1489_,
		_w1490_
	);
	LUT2 #(
		.INIT('h8)
	) name756 (
		\u2_adr0_cnt_reg[13]/P0001 ,
		\u2_adr0_cnt_reg[14]/P0001 ,
		_w1491_
	);
	LUT2 #(
		.INIT('h8)
	) name757 (
		_w1378_,
		_w1491_,
		_w1492_
	);
	LUT3 #(
		.INIT('h80)
	) name758 (
		\u2_adr0_cnt_reg[15]/P0001 ,
		_w1375_,
		_w1492_,
		_w1493_
	);
	LUT2 #(
		.INIT('h8)
	) name759 (
		\u2_adr1_cnt_reg[13]/P0001 ,
		\u2_adr1_cnt_reg[14]/P0001 ,
		_w1494_
	);
	LUT2 #(
		.INIT('h8)
	) name760 (
		_w1387_,
		_w1494_,
		_w1495_
	);
	LUT3 #(
		.INIT('h80)
	) name761 (
		\u2_adr1_cnt_reg[15]/P0001 ,
		_w1384_,
		_w1495_,
		_w1496_
	);
	LUT2 #(
		.INIT('h8)
	) name762 (
		\u0_int_maskb_r_reg[0]/NET0131 ,
		_w1413_,
		_w1497_
	);
	LUT4 #(
		.INIT('h0008)
	) name763 (
		\u2_state_reg[10]/NET0131 ,
		_w1051_,
		_w1404_,
		_w1405_,
		_w1498_
	);
	LUT4 #(
		.INIT('h0400)
	) name764 (
		_w1391_,
		_w1393_,
		_w1396_,
		_w1498_,
		_w1499_
	);
	LUT2 #(
		.INIT('h8)
	) name765 (
		\u0_u0_ch_csr_r3_reg[2]/NET0131 ,
		\u0_u0_int_src_r_reg[2]/NET0131 ,
		_w1500_
	);
	LUT4 #(
		.INIT('h135f)
	) name766 (
		\u0_u0_ch_csr_r3_reg[0]/NET0131 ,
		\u0_u0_ch_csr_r3_reg[1]/NET0131 ,
		\u0_u0_ch_err_reg/NET0131 ,
		\u0_u0_int_src_r_reg[1]/NET0131 ,
		_w1501_
	);
	LUT3 #(
		.INIT('h8a)
	) name767 (
		\u0_int_maska_r_reg[0]/NET0131 ,
		_w1500_,
		_w1501_,
		_w1502_
	);
	LUT3 #(
		.INIT('h8a)
	) name768 (
		\u0_int_maskb_r_reg[0]/NET0131 ,
		_w1500_,
		_w1501_,
		_w1503_
	);
	LUT4 #(
		.INIT('h153f)
	) name769 (
		_w1406_,
		_w1409_,
		_w1502_,
		_w1503_,
		_w1504_
	);
	LUT3 #(
		.INIT('h0b)
	) name770 (
		_w1391_,
		_w1393_,
		_w1396_,
		_w1505_
	);
	LUT3 #(
		.INIT('h45)
	) name771 (
		_w1499_,
		_w1504_,
		_w1505_,
		_w1506_
	);
	LUT2 #(
		.INIT('h8)
	) name772 (
		\u0_int_maska_r_reg[0]/NET0131 ,
		_w1411_,
		_w1507_
	);
	LUT4 #(
		.INIT('h153f)
	) name773 (
		\u0_u0_ch_csr_r_reg[0]/NET0131 ,
		\u0_u0_ch_tot_sz_r_reg[0]/P0001 ,
		_w1408_,
		_w1418_,
		_w1508_
	);
	LUT4 #(
		.INIT('hfbff)
	) name774 (
		_w1497_,
		_w1506_,
		_w1507_,
		_w1508_,
		_w1509_
	);
	LUT2 #(
		.INIT('h8)
	) name775 (
		\u2_adr0_cnt_reg[7]/P0001 ,
		\u2_adr0_cnt_reg[8]/P0001 ,
		_w1510_
	);
	LUT4 #(
		.INIT('h6ccc)
	) name776 (
		\u2_adr0_cnt_reg[7]/P0001 ,
		\u2_adr0_cnt_reg[8]/P0001 ,
		_w1372_,
		_w1373_,
		_w1511_
	);
	LUT2 #(
		.INIT('h8)
	) name777 (
		\u2_adr1_cnt_reg[7]/P0001 ,
		\u2_adr1_cnt_reg[8]/P0001 ,
		_w1512_
	);
	LUT4 #(
		.INIT('h6ccc)
	) name778 (
		\u2_adr1_cnt_reg[7]/P0001 ,
		\u2_adr1_cnt_reg[8]/P0001 ,
		_w1381_,
		_w1382_,
		_w1513_
	);
	LUT2 #(
		.INIT('h4)
	) name779 (
		\u3_u1_slv_adr_reg[2]/NET0131 ,
		\u3_u1_slv_adr_reg[3]/P0001 ,
		_w1514_
	);
	LUT3 #(
		.INIT('h80)
	) name780 (
		_w1051_,
		_w1252_,
		_w1514_,
		_w1515_
	);
	LUT2 #(
		.INIT('h8)
	) name781 (
		\u2_mast0_drdy_r_reg/P0001 ,
		\u2_state_reg[6]/NET0131 ,
		_w1516_
	);
	LUT3 #(
		.INIT('h15)
	) name782 (
		\u0_u0_ch_adr0_r_reg[10]/P0001 ,
		\u2_mast0_drdy_r_reg/P0001 ,
		\u2_state_reg[6]/NET0131 ,
		_w1517_
	);
	LUT3 #(
		.INIT('h10)
	) name783 (
		_w1090_,
		_w1515_,
		_w1517_,
		_w1518_
	);
	LUT3 #(
		.INIT('h53)
	) name784 (
		\u2_adr0_cnt_reg[10]/P0001 ,
		\u3_u0_mast_dout_reg[12]/P0001 ,
		_w895_,
		_w1519_
	);
	LUT4 #(
		.INIT('h3200)
	) name785 (
		_w1090_,
		_w1515_,
		_w1516_,
		_w1519_,
		_w1520_
	);
	LUT3 #(
		.INIT('h04)
	) name786 (
		\u3_u1_slv_adr_reg[2]/NET0131 ,
		\u3_u1_slv_adr_reg[3]/P0001 ,
		\u3_u1_slv_dout_reg[12]/P0001 ,
		_w1521_
	);
	LUT3 #(
		.INIT('h80)
	) name787 (
		_w1051_,
		_w1252_,
		_w1521_,
		_w1522_
	);
	LUT3 #(
		.INIT('h01)
	) name788 (
		_w1518_,
		_w1520_,
		_w1522_,
		_w1523_
	);
	LUT3 #(
		.INIT('h15)
	) name789 (
		\u0_u0_ch_adr0_r_reg[11]/P0001 ,
		\u2_mast0_drdy_r_reg/P0001 ,
		\u2_state_reg[6]/NET0131 ,
		_w1524_
	);
	LUT3 #(
		.INIT('h10)
	) name790 (
		_w1090_,
		_w1515_,
		_w1524_,
		_w1525_
	);
	LUT3 #(
		.INIT('h53)
	) name791 (
		\u2_adr0_cnt_reg[11]/P0001 ,
		\u3_u0_mast_dout_reg[13]/P0001 ,
		_w895_,
		_w1526_
	);
	LUT4 #(
		.INIT('h3200)
	) name792 (
		_w1090_,
		_w1515_,
		_w1516_,
		_w1526_,
		_w1527_
	);
	LUT3 #(
		.INIT('h04)
	) name793 (
		\u3_u1_slv_adr_reg[2]/NET0131 ,
		\u3_u1_slv_adr_reg[3]/P0001 ,
		\u3_u1_slv_dout_reg[13]/P0001 ,
		_w1528_
	);
	LUT3 #(
		.INIT('h80)
	) name794 (
		_w1051_,
		_w1252_,
		_w1528_,
		_w1529_
	);
	LUT3 #(
		.INIT('h01)
	) name795 (
		_w1525_,
		_w1527_,
		_w1529_,
		_w1530_
	);
	LUT3 #(
		.INIT('h15)
	) name796 (
		\u0_u0_ch_adr0_r_reg[12]/P0001 ,
		\u2_mast0_drdy_r_reg/P0001 ,
		\u2_state_reg[6]/NET0131 ,
		_w1531_
	);
	LUT3 #(
		.INIT('h10)
	) name797 (
		_w1090_,
		_w1515_,
		_w1531_,
		_w1532_
	);
	LUT3 #(
		.INIT('h53)
	) name798 (
		\u2_adr0_cnt_reg[12]/P0001 ,
		\u3_u0_mast_dout_reg[14]/P0001 ,
		_w895_,
		_w1533_
	);
	LUT4 #(
		.INIT('h3200)
	) name799 (
		_w1090_,
		_w1515_,
		_w1516_,
		_w1533_,
		_w1534_
	);
	LUT3 #(
		.INIT('h04)
	) name800 (
		\u3_u1_slv_adr_reg[2]/NET0131 ,
		\u3_u1_slv_adr_reg[3]/P0001 ,
		\u3_u1_slv_dout_reg[14]/P0001 ,
		_w1535_
	);
	LUT3 #(
		.INIT('h80)
	) name801 (
		_w1051_,
		_w1252_,
		_w1535_,
		_w1536_
	);
	LUT3 #(
		.INIT('h01)
	) name802 (
		_w1532_,
		_w1534_,
		_w1536_,
		_w1537_
	);
	LUT3 #(
		.INIT('h15)
	) name803 (
		\u0_u0_ch_adr0_r_reg[13]/P0001 ,
		\u2_mast0_drdy_r_reg/P0001 ,
		\u2_state_reg[6]/NET0131 ,
		_w1538_
	);
	LUT3 #(
		.INIT('h10)
	) name804 (
		_w1090_,
		_w1515_,
		_w1538_,
		_w1539_
	);
	LUT3 #(
		.INIT('h53)
	) name805 (
		\u2_adr0_cnt_reg[13]/P0001 ,
		\u3_u0_mast_dout_reg[15]/P0001 ,
		_w895_,
		_w1540_
	);
	LUT4 #(
		.INIT('h3200)
	) name806 (
		_w1090_,
		_w1515_,
		_w1516_,
		_w1540_,
		_w1541_
	);
	LUT3 #(
		.INIT('h04)
	) name807 (
		\u3_u1_slv_adr_reg[2]/NET0131 ,
		\u3_u1_slv_adr_reg[3]/P0001 ,
		\u3_u1_slv_dout_reg[15]/P0001 ,
		_w1542_
	);
	LUT3 #(
		.INIT('h80)
	) name808 (
		_w1051_,
		_w1252_,
		_w1542_,
		_w1543_
	);
	LUT3 #(
		.INIT('h01)
	) name809 (
		_w1539_,
		_w1541_,
		_w1543_,
		_w1544_
	);
	LUT3 #(
		.INIT('h15)
	) name810 (
		\u0_u0_ch_adr0_r_reg[14]/P0001 ,
		\u2_mast0_drdy_r_reg/P0001 ,
		\u2_state_reg[6]/NET0131 ,
		_w1545_
	);
	LUT3 #(
		.INIT('h10)
	) name811 (
		_w1090_,
		_w1515_,
		_w1545_,
		_w1546_
	);
	LUT3 #(
		.INIT('h53)
	) name812 (
		\u2_adr0_cnt_reg[14]/P0001 ,
		\u3_u0_mast_dout_reg[16]/P0001 ,
		_w895_,
		_w1547_
	);
	LUT4 #(
		.INIT('h3200)
	) name813 (
		_w1090_,
		_w1515_,
		_w1516_,
		_w1547_,
		_w1548_
	);
	LUT3 #(
		.INIT('h04)
	) name814 (
		\u3_u1_slv_adr_reg[2]/NET0131 ,
		\u3_u1_slv_adr_reg[3]/P0001 ,
		\u3_u1_slv_dout_reg[16]/P0001 ,
		_w1549_
	);
	LUT3 #(
		.INIT('h80)
	) name815 (
		_w1051_,
		_w1252_,
		_w1549_,
		_w1550_
	);
	LUT3 #(
		.INIT('h01)
	) name816 (
		_w1546_,
		_w1548_,
		_w1550_,
		_w1551_
	);
	LUT3 #(
		.INIT('h15)
	) name817 (
		\u0_u0_ch_adr0_r_reg[15]/P0001 ,
		\u2_mast0_drdy_r_reg/P0001 ,
		\u2_state_reg[6]/NET0131 ,
		_w1552_
	);
	LUT3 #(
		.INIT('h10)
	) name818 (
		_w1090_,
		_w1515_,
		_w1552_,
		_w1553_
	);
	LUT3 #(
		.INIT('h53)
	) name819 (
		\u2_adr0_cnt_reg[15]/P0001 ,
		\u3_u0_mast_dout_reg[17]/P0001 ,
		_w895_,
		_w1554_
	);
	LUT4 #(
		.INIT('h3200)
	) name820 (
		_w1090_,
		_w1515_,
		_w1516_,
		_w1554_,
		_w1555_
	);
	LUT3 #(
		.INIT('h04)
	) name821 (
		\u3_u1_slv_adr_reg[2]/NET0131 ,
		\u3_u1_slv_adr_reg[3]/P0001 ,
		\u3_u1_slv_dout_reg[17]/P0001 ,
		_w1556_
	);
	LUT3 #(
		.INIT('h80)
	) name822 (
		_w1051_,
		_w1252_,
		_w1556_,
		_w1557_
	);
	LUT3 #(
		.INIT('h01)
	) name823 (
		_w1553_,
		_w1555_,
		_w1557_,
		_w1558_
	);
	LUT3 #(
		.INIT('h15)
	) name824 (
		\u0_u0_ch_adr0_r_reg[16]/P0001 ,
		\u2_mast0_drdy_r_reg/P0001 ,
		\u2_state_reg[6]/NET0131 ,
		_w1559_
	);
	LUT3 #(
		.INIT('h10)
	) name825 (
		_w1090_,
		_w1515_,
		_w1559_,
		_w1560_
	);
	LUT3 #(
		.INIT('h53)
	) name826 (
		\u2_adr0_cnt_reg[16]/NET0131 ,
		\u3_u0_mast_dout_reg[18]/P0001 ,
		_w895_,
		_w1561_
	);
	LUT4 #(
		.INIT('h3200)
	) name827 (
		_w1090_,
		_w1515_,
		_w1516_,
		_w1561_,
		_w1562_
	);
	LUT3 #(
		.INIT('h04)
	) name828 (
		\u3_u1_slv_adr_reg[2]/NET0131 ,
		\u3_u1_slv_adr_reg[3]/P0001 ,
		\u3_u1_slv_dout_reg[18]/P0001 ,
		_w1563_
	);
	LUT3 #(
		.INIT('h80)
	) name829 (
		_w1051_,
		_w1252_,
		_w1563_,
		_w1564_
	);
	LUT3 #(
		.INIT('h01)
	) name830 (
		_w1560_,
		_w1562_,
		_w1564_,
		_w1565_
	);
	LUT3 #(
		.INIT('h15)
	) name831 (
		\u0_u0_ch_adr0_r_reg[17]/P0001 ,
		\u2_mast0_drdy_r_reg/P0001 ,
		\u2_state_reg[6]/NET0131 ,
		_w1566_
	);
	LUT3 #(
		.INIT('h10)
	) name832 (
		_w1090_,
		_w1515_,
		_w1566_,
		_w1567_
	);
	LUT3 #(
		.INIT('h53)
	) name833 (
		\u2_adr0_cnt_reg[17]/P0001 ,
		\u3_u0_mast_dout_reg[19]/P0001 ,
		_w895_,
		_w1568_
	);
	LUT4 #(
		.INIT('h3200)
	) name834 (
		_w1090_,
		_w1515_,
		_w1516_,
		_w1568_,
		_w1569_
	);
	LUT3 #(
		.INIT('h04)
	) name835 (
		\u3_u1_slv_adr_reg[2]/NET0131 ,
		\u3_u1_slv_adr_reg[3]/P0001 ,
		\u3_u1_slv_dout_reg[19]/P0001 ,
		_w1570_
	);
	LUT3 #(
		.INIT('h80)
	) name836 (
		_w1051_,
		_w1252_,
		_w1570_,
		_w1571_
	);
	LUT3 #(
		.INIT('h01)
	) name837 (
		_w1567_,
		_w1569_,
		_w1571_,
		_w1572_
	);
	LUT3 #(
		.INIT('h15)
	) name838 (
		\u0_u0_ch_adr0_r_reg[18]/P0001 ,
		\u2_mast0_drdy_r_reg/P0001 ,
		\u2_state_reg[6]/NET0131 ,
		_w1573_
	);
	LUT3 #(
		.INIT('h10)
	) name839 (
		_w1090_,
		_w1515_,
		_w1573_,
		_w1574_
	);
	LUT3 #(
		.INIT('h53)
	) name840 (
		\u2_adr0_cnt_reg[18]/P0001 ,
		\u3_u0_mast_dout_reg[20]/P0001 ,
		_w895_,
		_w1575_
	);
	LUT4 #(
		.INIT('h3200)
	) name841 (
		_w1090_,
		_w1515_,
		_w1516_,
		_w1575_,
		_w1576_
	);
	LUT3 #(
		.INIT('h04)
	) name842 (
		\u3_u1_slv_adr_reg[2]/NET0131 ,
		\u3_u1_slv_adr_reg[3]/P0001 ,
		\u3_u1_slv_dout_reg[20]/P0001 ,
		_w1577_
	);
	LUT3 #(
		.INIT('h80)
	) name843 (
		_w1051_,
		_w1252_,
		_w1577_,
		_w1578_
	);
	LUT3 #(
		.INIT('h01)
	) name844 (
		_w1574_,
		_w1576_,
		_w1578_,
		_w1579_
	);
	LUT3 #(
		.INIT('h15)
	) name845 (
		\u0_u0_ch_adr0_r_reg[19]/P0001 ,
		\u2_mast0_drdy_r_reg/P0001 ,
		\u2_state_reg[6]/NET0131 ,
		_w1580_
	);
	LUT3 #(
		.INIT('h10)
	) name846 (
		_w1090_,
		_w1515_,
		_w1580_,
		_w1581_
	);
	LUT3 #(
		.INIT('h53)
	) name847 (
		\u2_adr0_cnt_reg[19]/P0001 ,
		\u3_u0_mast_dout_reg[21]/P0001 ,
		_w895_,
		_w1582_
	);
	LUT4 #(
		.INIT('h3200)
	) name848 (
		_w1090_,
		_w1515_,
		_w1516_,
		_w1582_,
		_w1583_
	);
	LUT3 #(
		.INIT('h04)
	) name849 (
		\u3_u1_slv_adr_reg[2]/NET0131 ,
		\u3_u1_slv_adr_reg[3]/P0001 ,
		\u3_u1_slv_dout_reg[21]/P0001 ,
		_w1584_
	);
	LUT3 #(
		.INIT('h80)
	) name850 (
		_w1051_,
		_w1252_,
		_w1584_,
		_w1585_
	);
	LUT3 #(
		.INIT('h01)
	) name851 (
		_w1581_,
		_w1583_,
		_w1585_,
		_w1586_
	);
	LUT3 #(
		.INIT('h15)
	) name852 (
		\u0_u0_ch_adr0_r_reg[20]/P0001 ,
		\u2_mast0_drdy_r_reg/P0001 ,
		\u2_state_reg[6]/NET0131 ,
		_w1587_
	);
	LUT3 #(
		.INIT('h10)
	) name853 (
		_w1090_,
		_w1515_,
		_w1587_,
		_w1588_
	);
	LUT3 #(
		.INIT('h53)
	) name854 (
		\u2_adr0_cnt_reg[20]/P0001 ,
		\u3_u0_mast_dout_reg[22]/P0001 ,
		_w895_,
		_w1589_
	);
	LUT4 #(
		.INIT('h3200)
	) name855 (
		_w1090_,
		_w1515_,
		_w1516_,
		_w1589_,
		_w1590_
	);
	LUT3 #(
		.INIT('h04)
	) name856 (
		\u3_u1_slv_adr_reg[2]/NET0131 ,
		\u3_u1_slv_adr_reg[3]/P0001 ,
		\u3_u1_slv_dout_reg[22]/P0001 ,
		_w1591_
	);
	LUT3 #(
		.INIT('h80)
	) name857 (
		_w1051_,
		_w1252_,
		_w1591_,
		_w1592_
	);
	LUT3 #(
		.INIT('h01)
	) name858 (
		_w1588_,
		_w1590_,
		_w1592_,
		_w1593_
	);
	LUT3 #(
		.INIT('h15)
	) name859 (
		\u0_u0_ch_adr0_r_reg[21]/P0001 ,
		\u2_mast0_drdy_r_reg/P0001 ,
		\u2_state_reg[6]/NET0131 ,
		_w1594_
	);
	LUT3 #(
		.INIT('h10)
	) name860 (
		_w1090_,
		_w1515_,
		_w1594_,
		_w1595_
	);
	LUT3 #(
		.INIT('h53)
	) name861 (
		\u2_adr0_cnt_reg[21]/P0001 ,
		\u3_u0_mast_dout_reg[23]/P0001 ,
		_w895_,
		_w1596_
	);
	LUT4 #(
		.INIT('h3200)
	) name862 (
		_w1090_,
		_w1515_,
		_w1516_,
		_w1596_,
		_w1597_
	);
	LUT3 #(
		.INIT('h04)
	) name863 (
		\u3_u1_slv_adr_reg[2]/NET0131 ,
		\u3_u1_slv_adr_reg[3]/P0001 ,
		\u3_u1_slv_dout_reg[23]/P0001 ,
		_w1598_
	);
	LUT3 #(
		.INIT('h80)
	) name864 (
		_w1051_,
		_w1252_,
		_w1598_,
		_w1599_
	);
	LUT3 #(
		.INIT('h01)
	) name865 (
		_w1595_,
		_w1597_,
		_w1599_,
		_w1600_
	);
	LUT3 #(
		.INIT('h15)
	) name866 (
		\u0_u0_ch_adr0_r_reg[22]/P0001 ,
		\u2_mast0_drdy_r_reg/P0001 ,
		\u2_state_reg[6]/NET0131 ,
		_w1601_
	);
	LUT3 #(
		.INIT('h10)
	) name867 (
		_w1090_,
		_w1515_,
		_w1601_,
		_w1602_
	);
	LUT3 #(
		.INIT('h53)
	) name868 (
		\u2_adr0_cnt_reg[22]/P0001 ,
		\u3_u0_mast_dout_reg[24]/P0001 ,
		_w895_,
		_w1603_
	);
	LUT4 #(
		.INIT('h3200)
	) name869 (
		_w1090_,
		_w1515_,
		_w1516_,
		_w1603_,
		_w1604_
	);
	LUT3 #(
		.INIT('h04)
	) name870 (
		\u3_u1_slv_adr_reg[2]/NET0131 ,
		\u3_u1_slv_adr_reg[3]/P0001 ,
		\u3_u1_slv_dout_reg[24]/P0001 ,
		_w1605_
	);
	LUT3 #(
		.INIT('h80)
	) name871 (
		_w1051_,
		_w1252_,
		_w1605_,
		_w1606_
	);
	LUT3 #(
		.INIT('h01)
	) name872 (
		_w1602_,
		_w1604_,
		_w1606_,
		_w1607_
	);
	LUT3 #(
		.INIT('h15)
	) name873 (
		\u0_u0_ch_adr0_r_reg[23]/P0001 ,
		\u2_mast0_drdy_r_reg/P0001 ,
		\u2_state_reg[6]/NET0131 ,
		_w1608_
	);
	LUT3 #(
		.INIT('h10)
	) name874 (
		_w1090_,
		_w1515_,
		_w1608_,
		_w1609_
	);
	LUT3 #(
		.INIT('h53)
	) name875 (
		\u2_adr0_cnt_reg[23]/P0001 ,
		\u3_u0_mast_dout_reg[25]/P0001 ,
		_w895_,
		_w1610_
	);
	LUT4 #(
		.INIT('h3200)
	) name876 (
		_w1090_,
		_w1515_,
		_w1516_,
		_w1610_,
		_w1611_
	);
	LUT3 #(
		.INIT('h04)
	) name877 (
		\u3_u1_slv_adr_reg[2]/NET0131 ,
		\u3_u1_slv_adr_reg[3]/P0001 ,
		\u3_u1_slv_dout_reg[25]/P0001 ,
		_w1612_
	);
	LUT3 #(
		.INIT('h80)
	) name878 (
		_w1051_,
		_w1252_,
		_w1612_,
		_w1613_
	);
	LUT3 #(
		.INIT('h01)
	) name879 (
		_w1609_,
		_w1611_,
		_w1613_,
		_w1614_
	);
	LUT3 #(
		.INIT('h15)
	) name880 (
		\u0_u0_ch_adr0_r_reg[24]/P0001 ,
		\u2_mast0_drdy_r_reg/P0001 ,
		\u2_state_reg[6]/NET0131 ,
		_w1615_
	);
	LUT3 #(
		.INIT('h10)
	) name881 (
		_w1090_,
		_w1515_,
		_w1615_,
		_w1616_
	);
	LUT3 #(
		.INIT('h53)
	) name882 (
		\u2_adr0_cnt_reg[24]/P0001 ,
		\u3_u0_mast_dout_reg[26]/P0001 ,
		_w895_,
		_w1617_
	);
	LUT4 #(
		.INIT('h3200)
	) name883 (
		_w1090_,
		_w1515_,
		_w1516_,
		_w1617_,
		_w1618_
	);
	LUT3 #(
		.INIT('h04)
	) name884 (
		\u3_u1_slv_adr_reg[2]/NET0131 ,
		\u3_u1_slv_adr_reg[3]/P0001 ,
		\u3_u1_slv_dout_reg[26]/P0001 ,
		_w1619_
	);
	LUT3 #(
		.INIT('h80)
	) name885 (
		_w1051_,
		_w1252_,
		_w1619_,
		_w1620_
	);
	LUT3 #(
		.INIT('h01)
	) name886 (
		_w1616_,
		_w1618_,
		_w1620_,
		_w1621_
	);
	LUT3 #(
		.INIT('h15)
	) name887 (
		\u0_u0_ch_adr0_r_reg[25]/P0001 ,
		\u2_mast0_drdy_r_reg/P0001 ,
		\u2_state_reg[6]/NET0131 ,
		_w1622_
	);
	LUT3 #(
		.INIT('h10)
	) name888 (
		_w1090_,
		_w1515_,
		_w1622_,
		_w1623_
	);
	LUT3 #(
		.INIT('h53)
	) name889 (
		\u2_adr0_cnt_reg[25]/P0001 ,
		\u3_u0_mast_dout_reg[27]/P0001 ,
		_w895_,
		_w1624_
	);
	LUT4 #(
		.INIT('h3200)
	) name890 (
		_w1090_,
		_w1515_,
		_w1516_,
		_w1624_,
		_w1625_
	);
	LUT3 #(
		.INIT('h04)
	) name891 (
		\u3_u1_slv_adr_reg[2]/NET0131 ,
		\u3_u1_slv_adr_reg[3]/P0001 ,
		\u3_u1_slv_dout_reg[27]/P0001 ,
		_w1626_
	);
	LUT3 #(
		.INIT('h80)
	) name892 (
		_w1051_,
		_w1252_,
		_w1626_,
		_w1627_
	);
	LUT3 #(
		.INIT('h01)
	) name893 (
		_w1623_,
		_w1625_,
		_w1627_,
		_w1628_
	);
	LUT3 #(
		.INIT('h15)
	) name894 (
		\u0_u0_ch_adr0_r_reg[26]/P0001 ,
		\u2_mast0_drdy_r_reg/P0001 ,
		\u2_state_reg[6]/NET0131 ,
		_w1629_
	);
	LUT3 #(
		.INIT('h10)
	) name895 (
		_w1090_,
		_w1515_,
		_w1629_,
		_w1630_
	);
	LUT3 #(
		.INIT('h53)
	) name896 (
		\u2_adr0_cnt_reg[26]/P0001 ,
		\u3_u0_mast_dout_reg[28]/P0001 ,
		_w895_,
		_w1631_
	);
	LUT4 #(
		.INIT('h3200)
	) name897 (
		_w1090_,
		_w1515_,
		_w1516_,
		_w1631_,
		_w1632_
	);
	LUT3 #(
		.INIT('h04)
	) name898 (
		\u3_u1_slv_adr_reg[2]/NET0131 ,
		\u3_u1_slv_adr_reg[3]/P0001 ,
		\u3_u1_slv_dout_reg[28]/P0001 ,
		_w1633_
	);
	LUT3 #(
		.INIT('h80)
	) name899 (
		_w1051_,
		_w1252_,
		_w1633_,
		_w1634_
	);
	LUT3 #(
		.INIT('h01)
	) name900 (
		_w1630_,
		_w1632_,
		_w1634_,
		_w1635_
	);
	LUT3 #(
		.INIT('h15)
	) name901 (
		\u0_u0_ch_adr0_r_reg[27]/P0001 ,
		\u2_mast0_drdy_r_reg/P0001 ,
		\u2_state_reg[6]/NET0131 ,
		_w1636_
	);
	LUT3 #(
		.INIT('h10)
	) name902 (
		_w1090_,
		_w1515_,
		_w1636_,
		_w1637_
	);
	LUT3 #(
		.INIT('h53)
	) name903 (
		\u2_adr0_cnt_reg[27]/P0001 ,
		\u3_u0_mast_dout_reg[29]/P0001 ,
		_w895_,
		_w1638_
	);
	LUT4 #(
		.INIT('h3200)
	) name904 (
		_w1090_,
		_w1515_,
		_w1516_,
		_w1638_,
		_w1639_
	);
	LUT3 #(
		.INIT('h04)
	) name905 (
		\u3_u1_slv_adr_reg[2]/NET0131 ,
		\u3_u1_slv_adr_reg[3]/P0001 ,
		\u3_u1_slv_dout_reg[29]/P0001 ,
		_w1640_
	);
	LUT3 #(
		.INIT('h80)
	) name906 (
		_w1051_,
		_w1252_,
		_w1640_,
		_w1641_
	);
	LUT3 #(
		.INIT('h01)
	) name907 (
		_w1637_,
		_w1639_,
		_w1641_,
		_w1642_
	);
	LUT3 #(
		.INIT('h15)
	) name908 (
		\u0_u0_ch_adr0_r_reg[28]/P0001 ,
		\u2_mast0_drdy_r_reg/P0001 ,
		\u2_state_reg[6]/NET0131 ,
		_w1643_
	);
	LUT3 #(
		.INIT('h10)
	) name909 (
		_w1090_,
		_w1515_,
		_w1643_,
		_w1644_
	);
	LUT3 #(
		.INIT('h53)
	) name910 (
		\u2_adr0_cnt_reg[28]/P0001 ,
		\u3_u0_mast_dout_reg[30]/P0001 ,
		_w895_,
		_w1645_
	);
	LUT4 #(
		.INIT('h3200)
	) name911 (
		_w1090_,
		_w1515_,
		_w1516_,
		_w1645_,
		_w1646_
	);
	LUT3 #(
		.INIT('h04)
	) name912 (
		\u3_u1_slv_adr_reg[2]/NET0131 ,
		\u3_u1_slv_adr_reg[3]/P0001 ,
		\u3_u1_slv_dout_reg[30]/P0001 ,
		_w1647_
	);
	LUT3 #(
		.INIT('h80)
	) name913 (
		_w1051_,
		_w1252_,
		_w1647_,
		_w1648_
	);
	LUT3 #(
		.INIT('h01)
	) name914 (
		_w1644_,
		_w1646_,
		_w1648_,
		_w1649_
	);
	LUT3 #(
		.INIT('h15)
	) name915 (
		\u0_u0_ch_adr0_r_reg[29]/P0001 ,
		\u2_mast0_drdy_r_reg/P0001 ,
		\u2_state_reg[6]/NET0131 ,
		_w1650_
	);
	LUT3 #(
		.INIT('h10)
	) name916 (
		_w1090_,
		_w1515_,
		_w1650_,
		_w1651_
	);
	LUT3 #(
		.INIT('h53)
	) name917 (
		\u2_adr0_cnt_reg[29]/P0001 ,
		\u3_u0_mast_dout_reg[31]/P0001 ,
		_w895_,
		_w1652_
	);
	LUT4 #(
		.INIT('h3200)
	) name918 (
		_w1090_,
		_w1515_,
		_w1516_,
		_w1652_,
		_w1653_
	);
	LUT3 #(
		.INIT('h04)
	) name919 (
		\u3_u1_slv_adr_reg[2]/NET0131 ,
		\u3_u1_slv_adr_reg[3]/P0001 ,
		\u3_u1_slv_dout_reg[31]/P0001 ,
		_w1654_
	);
	LUT3 #(
		.INIT('h80)
	) name920 (
		_w1051_,
		_w1252_,
		_w1654_,
		_w1655_
	);
	LUT3 #(
		.INIT('h01)
	) name921 (
		_w1651_,
		_w1653_,
		_w1655_,
		_w1656_
	);
	LUT2 #(
		.INIT('h8)
	) name922 (
		\u3_u1_slv_adr_reg[4]/NET0131 ,
		\u3_u1_slv_we_reg/P0001 ,
		_w1657_
	);
	LUT3 #(
		.INIT('h80)
	) name923 (
		_w1051_,
		_w1053_,
		_w1657_,
		_w1658_
	);
	LUT2 #(
		.INIT('h4)
	) name924 (
		\u2_mast0_drdy_r_reg/P0001 ,
		\u2_state_reg[7]/NET0131 ,
		_w1659_
	);
	LUT3 #(
		.INIT('h10)
	) name925 (
		\u0_u0_ch_adr1_r_reg[10]/P0001 ,
		\u2_mast0_drdy_r_reg/P0001 ,
		\u2_state_reg[7]/NET0131 ,
		_w1660_
	);
	LUT2 #(
		.INIT('h1)
	) name926 (
		\u0_u0_ch_adr1_r_reg[10]/P0001 ,
		\u2_state_reg[7]/NET0131 ,
		_w1661_
	);
	LUT3 #(
		.INIT('h23)
	) name927 (
		_w1090_,
		_w1660_,
		_w1661_,
		_w1662_
	);
	LUT4 #(
		.INIT('h0053)
	) name928 (
		\u2_adr1_cnt_reg[10]/P0001 ,
		\u3_u0_mast_dout_reg[12]/P0001 ,
		_w895_,
		_w1659_,
		_w1663_
	);
	LUT3 #(
		.INIT('he0)
	) name929 (
		\u2_state_reg[7]/NET0131 ,
		_w1090_,
		_w1663_,
		_w1664_
	);
	LUT3 #(
		.INIT('h20)
	) name930 (
		\u3_u1_slv_adr_reg[4]/NET0131 ,
		\u3_u1_slv_dout_reg[12]/P0001 ,
		\u3_u1_slv_we_reg/P0001 ,
		_w1665_
	);
	LUT3 #(
		.INIT('h80)
	) name931 (
		_w1051_,
		_w1053_,
		_w1665_,
		_w1666_
	);
	LUT4 #(
		.INIT('h00ae)
	) name932 (
		_w1658_,
		_w1662_,
		_w1664_,
		_w1666_,
		_w1667_
	);
	LUT3 #(
		.INIT('h10)
	) name933 (
		\u0_u0_ch_adr1_r_reg[11]/P0001 ,
		\u2_mast0_drdy_r_reg/P0001 ,
		\u2_state_reg[7]/NET0131 ,
		_w1668_
	);
	LUT2 #(
		.INIT('h1)
	) name934 (
		\u0_u0_ch_adr1_r_reg[11]/P0001 ,
		\u2_state_reg[7]/NET0131 ,
		_w1669_
	);
	LUT3 #(
		.INIT('h23)
	) name935 (
		_w1090_,
		_w1668_,
		_w1669_,
		_w1670_
	);
	LUT4 #(
		.INIT('h0053)
	) name936 (
		\u2_adr1_cnt_reg[11]/P0001 ,
		\u3_u0_mast_dout_reg[13]/P0001 ,
		_w895_,
		_w1659_,
		_w1671_
	);
	LUT3 #(
		.INIT('he0)
	) name937 (
		\u2_state_reg[7]/NET0131 ,
		_w1090_,
		_w1671_,
		_w1672_
	);
	LUT3 #(
		.INIT('h20)
	) name938 (
		\u3_u1_slv_adr_reg[4]/NET0131 ,
		\u3_u1_slv_dout_reg[13]/P0001 ,
		\u3_u1_slv_we_reg/P0001 ,
		_w1673_
	);
	LUT3 #(
		.INIT('h80)
	) name939 (
		_w1051_,
		_w1053_,
		_w1673_,
		_w1674_
	);
	LUT4 #(
		.INIT('h00ae)
	) name940 (
		_w1658_,
		_w1670_,
		_w1672_,
		_w1674_,
		_w1675_
	);
	LUT3 #(
		.INIT('h10)
	) name941 (
		\u0_u0_ch_adr1_r_reg[12]/P0001 ,
		\u2_mast0_drdy_r_reg/P0001 ,
		\u2_state_reg[7]/NET0131 ,
		_w1676_
	);
	LUT2 #(
		.INIT('h1)
	) name942 (
		\u0_u0_ch_adr1_r_reg[12]/P0001 ,
		\u2_state_reg[7]/NET0131 ,
		_w1677_
	);
	LUT3 #(
		.INIT('h23)
	) name943 (
		_w1090_,
		_w1676_,
		_w1677_,
		_w1678_
	);
	LUT4 #(
		.INIT('h0053)
	) name944 (
		\u2_adr1_cnt_reg[12]/P0001 ,
		\u3_u0_mast_dout_reg[14]/P0001 ,
		_w895_,
		_w1659_,
		_w1679_
	);
	LUT3 #(
		.INIT('he0)
	) name945 (
		\u2_state_reg[7]/NET0131 ,
		_w1090_,
		_w1679_,
		_w1680_
	);
	LUT3 #(
		.INIT('h20)
	) name946 (
		\u3_u1_slv_adr_reg[4]/NET0131 ,
		\u3_u1_slv_dout_reg[14]/P0001 ,
		\u3_u1_slv_we_reg/P0001 ,
		_w1681_
	);
	LUT3 #(
		.INIT('h80)
	) name947 (
		_w1051_,
		_w1053_,
		_w1681_,
		_w1682_
	);
	LUT4 #(
		.INIT('h00ae)
	) name948 (
		_w1658_,
		_w1678_,
		_w1680_,
		_w1682_,
		_w1683_
	);
	LUT3 #(
		.INIT('h10)
	) name949 (
		\u0_u0_ch_adr1_r_reg[13]/P0001 ,
		\u2_mast0_drdy_r_reg/P0001 ,
		\u2_state_reg[7]/NET0131 ,
		_w1684_
	);
	LUT2 #(
		.INIT('h1)
	) name950 (
		\u0_u0_ch_adr1_r_reg[13]/P0001 ,
		\u2_state_reg[7]/NET0131 ,
		_w1685_
	);
	LUT3 #(
		.INIT('h23)
	) name951 (
		_w1090_,
		_w1684_,
		_w1685_,
		_w1686_
	);
	LUT4 #(
		.INIT('h0053)
	) name952 (
		\u2_adr1_cnt_reg[13]/P0001 ,
		\u3_u0_mast_dout_reg[15]/P0001 ,
		_w895_,
		_w1659_,
		_w1687_
	);
	LUT3 #(
		.INIT('he0)
	) name953 (
		\u2_state_reg[7]/NET0131 ,
		_w1090_,
		_w1687_,
		_w1688_
	);
	LUT3 #(
		.INIT('h20)
	) name954 (
		\u3_u1_slv_adr_reg[4]/NET0131 ,
		\u3_u1_slv_dout_reg[15]/P0001 ,
		\u3_u1_slv_we_reg/P0001 ,
		_w1689_
	);
	LUT3 #(
		.INIT('h80)
	) name955 (
		_w1051_,
		_w1053_,
		_w1689_,
		_w1690_
	);
	LUT4 #(
		.INIT('h00ae)
	) name956 (
		_w1658_,
		_w1686_,
		_w1688_,
		_w1690_,
		_w1691_
	);
	LUT3 #(
		.INIT('h10)
	) name957 (
		\u0_u0_ch_adr1_r_reg[14]/P0001 ,
		\u2_mast0_drdy_r_reg/P0001 ,
		\u2_state_reg[7]/NET0131 ,
		_w1692_
	);
	LUT2 #(
		.INIT('h1)
	) name958 (
		\u0_u0_ch_adr1_r_reg[14]/P0001 ,
		\u2_state_reg[7]/NET0131 ,
		_w1693_
	);
	LUT3 #(
		.INIT('h23)
	) name959 (
		_w1090_,
		_w1692_,
		_w1693_,
		_w1694_
	);
	LUT4 #(
		.INIT('h0053)
	) name960 (
		\u2_adr1_cnt_reg[14]/P0001 ,
		\u3_u0_mast_dout_reg[16]/P0001 ,
		_w895_,
		_w1659_,
		_w1695_
	);
	LUT3 #(
		.INIT('he0)
	) name961 (
		\u2_state_reg[7]/NET0131 ,
		_w1090_,
		_w1695_,
		_w1696_
	);
	LUT3 #(
		.INIT('h20)
	) name962 (
		\u3_u1_slv_adr_reg[4]/NET0131 ,
		\u3_u1_slv_dout_reg[16]/P0001 ,
		\u3_u1_slv_we_reg/P0001 ,
		_w1697_
	);
	LUT3 #(
		.INIT('h80)
	) name963 (
		_w1051_,
		_w1053_,
		_w1697_,
		_w1698_
	);
	LUT4 #(
		.INIT('h00ae)
	) name964 (
		_w1658_,
		_w1694_,
		_w1696_,
		_w1698_,
		_w1699_
	);
	LUT3 #(
		.INIT('h10)
	) name965 (
		\u0_u0_ch_adr1_r_reg[15]/P0001 ,
		\u2_mast0_drdy_r_reg/P0001 ,
		\u2_state_reg[7]/NET0131 ,
		_w1700_
	);
	LUT2 #(
		.INIT('h1)
	) name966 (
		\u0_u0_ch_adr1_r_reg[15]/P0001 ,
		\u2_state_reg[7]/NET0131 ,
		_w1701_
	);
	LUT3 #(
		.INIT('h23)
	) name967 (
		_w1090_,
		_w1700_,
		_w1701_,
		_w1702_
	);
	LUT4 #(
		.INIT('h0053)
	) name968 (
		\u2_adr1_cnt_reg[15]/P0001 ,
		\u3_u0_mast_dout_reg[17]/P0001 ,
		_w895_,
		_w1659_,
		_w1703_
	);
	LUT3 #(
		.INIT('he0)
	) name969 (
		\u2_state_reg[7]/NET0131 ,
		_w1090_,
		_w1703_,
		_w1704_
	);
	LUT3 #(
		.INIT('h20)
	) name970 (
		\u3_u1_slv_adr_reg[4]/NET0131 ,
		\u3_u1_slv_dout_reg[17]/P0001 ,
		\u3_u1_slv_we_reg/P0001 ,
		_w1705_
	);
	LUT3 #(
		.INIT('h80)
	) name971 (
		_w1051_,
		_w1053_,
		_w1705_,
		_w1706_
	);
	LUT4 #(
		.INIT('h00ae)
	) name972 (
		_w1658_,
		_w1702_,
		_w1704_,
		_w1706_,
		_w1707_
	);
	LUT3 #(
		.INIT('h10)
	) name973 (
		\u0_u0_ch_adr1_r_reg[16]/P0001 ,
		\u2_mast0_drdy_r_reg/P0001 ,
		\u2_state_reg[7]/NET0131 ,
		_w1708_
	);
	LUT2 #(
		.INIT('h1)
	) name974 (
		\u0_u0_ch_adr1_r_reg[16]/P0001 ,
		\u2_state_reg[7]/NET0131 ,
		_w1709_
	);
	LUT3 #(
		.INIT('h23)
	) name975 (
		_w1090_,
		_w1708_,
		_w1709_,
		_w1710_
	);
	LUT4 #(
		.INIT('h0053)
	) name976 (
		\u2_adr1_cnt_reg[16]/NET0131 ,
		\u3_u0_mast_dout_reg[18]/P0001 ,
		_w895_,
		_w1659_,
		_w1711_
	);
	LUT3 #(
		.INIT('he0)
	) name977 (
		\u2_state_reg[7]/NET0131 ,
		_w1090_,
		_w1711_,
		_w1712_
	);
	LUT3 #(
		.INIT('h20)
	) name978 (
		\u3_u1_slv_adr_reg[4]/NET0131 ,
		\u3_u1_slv_dout_reg[18]/P0001 ,
		\u3_u1_slv_we_reg/P0001 ,
		_w1713_
	);
	LUT3 #(
		.INIT('h80)
	) name979 (
		_w1051_,
		_w1053_,
		_w1713_,
		_w1714_
	);
	LUT4 #(
		.INIT('h00ae)
	) name980 (
		_w1658_,
		_w1710_,
		_w1712_,
		_w1714_,
		_w1715_
	);
	LUT3 #(
		.INIT('h10)
	) name981 (
		\u0_u0_ch_adr1_r_reg[17]/P0001 ,
		\u2_mast0_drdy_r_reg/P0001 ,
		\u2_state_reg[7]/NET0131 ,
		_w1716_
	);
	LUT2 #(
		.INIT('h1)
	) name982 (
		\u0_u0_ch_adr1_r_reg[17]/P0001 ,
		\u2_state_reg[7]/NET0131 ,
		_w1717_
	);
	LUT3 #(
		.INIT('h23)
	) name983 (
		_w1090_,
		_w1716_,
		_w1717_,
		_w1718_
	);
	LUT4 #(
		.INIT('h0053)
	) name984 (
		\u2_adr1_cnt_reg[17]/P0001 ,
		\u3_u0_mast_dout_reg[19]/P0001 ,
		_w895_,
		_w1659_,
		_w1719_
	);
	LUT3 #(
		.INIT('he0)
	) name985 (
		\u2_state_reg[7]/NET0131 ,
		_w1090_,
		_w1719_,
		_w1720_
	);
	LUT3 #(
		.INIT('h20)
	) name986 (
		\u3_u1_slv_adr_reg[4]/NET0131 ,
		\u3_u1_slv_dout_reg[19]/P0001 ,
		\u3_u1_slv_we_reg/P0001 ,
		_w1721_
	);
	LUT3 #(
		.INIT('h80)
	) name987 (
		_w1051_,
		_w1053_,
		_w1721_,
		_w1722_
	);
	LUT4 #(
		.INIT('h00ae)
	) name988 (
		_w1658_,
		_w1718_,
		_w1720_,
		_w1722_,
		_w1723_
	);
	LUT3 #(
		.INIT('h10)
	) name989 (
		\u0_u0_ch_adr1_r_reg[18]/P0001 ,
		\u2_mast0_drdy_r_reg/P0001 ,
		\u2_state_reg[7]/NET0131 ,
		_w1724_
	);
	LUT2 #(
		.INIT('h1)
	) name990 (
		\u0_u0_ch_adr1_r_reg[18]/P0001 ,
		\u2_state_reg[7]/NET0131 ,
		_w1725_
	);
	LUT3 #(
		.INIT('h23)
	) name991 (
		_w1090_,
		_w1724_,
		_w1725_,
		_w1726_
	);
	LUT4 #(
		.INIT('h0053)
	) name992 (
		\u2_adr1_cnt_reg[18]/P0001 ,
		\u3_u0_mast_dout_reg[20]/P0001 ,
		_w895_,
		_w1659_,
		_w1727_
	);
	LUT3 #(
		.INIT('he0)
	) name993 (
		\u2_state_reg[7]/NET0131 ,
		_w1090_,
		_w1727_,
		_w1728_
	);
	LUT3 #(
		.INIT('h20)
	) name994 (
		\u3_u1_slv_adr_reg[4]/NET0131 ,
		\u3_u1_slv_dout_reg[20]/P0001 ,
		\u3_u1_slv_we_reg/P0001 ,
		_w1729_
	);
	LUT3 #(
		.INIT('h80)
	) name995 (
		_w1051_,
		_w1053_,
		_w1729_,
		_w1730_
	);
	LUT4 #(
		.INIT('h00ae)
	) name996 (
		_w1658_,
		_w1726_,
		_w1728_,
		_w1730_,
		_w1731_
	);
	LUT3 #(
		.INIT('h10)
	) name997 (
		\u0_u0_ch_adr1_r_reg[19]/P0001 ,
		\u2_mast0_drdy_r_reg/P0001 ,
		\u2_state_reg[7]/NET0131 ,
		_w1732_
	);
	LUT2 #(
		.INIT('h1)
	) name998 (
		\u0_u0_ch_adr1_r_reg[19]/P0001 ,
		\u2_state_reg[7]/NET0131 ,
		_w1733_
	);
	LUT3 #(
		.INIT('h23)
	) name999 (
		_w1090_,
		_w1732_,
		_w1733_,
		_w1734_
	);
	LUT4 #(
		.INIT('h0053)
	) name1000 (
		\u2_adr1_cnt_reg[19]/P0001 ,
		\u3_u0_mast_dout_reg[21]/P0001 ,
		_w895_,
		_w1659_,
		_w1735_
	);
	LUT3 #(
		.INIT('he0)
	) name1001 (
		\u2_state_reg[7]/NET0131 ,
		_w1090_,
		_w1735_,
		_w1736_
	);
	LUT3 #(
		.INIT('h20)
	) name1002 (
		\u3_u1_slv_adr_reg[4]/NET0131 ,
		\u3_u1_slv_dout_reg[21]/P0001 ,
		\u3_u1_slv_we_reg/P0001 ,
		_w1737_
	);
	LUT3 #(
		.INIT('h80)
	) name1003 (
		_w1051_,
		_w1053_,
		_w1737_,
		_w1738_
	);
	LUT4 #(
		.INIT('h00ae)
	) name1004 (
		_w1658_,
		_w1734_,
		_w1736_,
		_w1738_,
		_w1739_
	);
	LUT3 #(
		.INIT('h10)
	) name1005 (
		\u0_u0_ch_adr1_r_reg[20]/P0001 ,
		\u2_mast0_drdy_r_reg/P0001 ,
		\u2_state_reg[7]/NET0131 ,
		_w1740_
	);
	LUT2 #(
		.INIT('h1)
	) name1006 (
		\u0_u0_ch_adr1_r_reg[20]/P0001 ,
		\u2_state_reg[7]/NET0131 ,
		_w1741_
	);
	LUT3 #(
		.INIT('h23)
	) name1007 (
		_w1090_,
		_w1740_,
		_w1741_,
		_w1742_
	);
	LUT4 #(
		.INIT('h0053)
	) name1008 (
		\u2_adr1_cnt_reg[20]/P0001 ,
		\u3_u0_mast_dout_reg[22]/P0001 ,
		_w895_,
		_w1659_,
		_w1743_
	);
	LUT3 #(
		.INIT('he0)
	) name1009 (
		\u2_state_reg[7]/NET0131 ,
		_w1090_,
		_w1743_,
		_w1744_
	);
	LUT3 #(
		.INIT('h20)
	) name1010 (
		\u3_u1_slv_adr_reg[4]/NET0131 ,
		\u3_u1_slv_dout_reg[22]/P0001 ,
		\u3_u1_slv_we_reg/P0001 ,
		_w1745_
	);
	LUT3 #(
		.INIT('h80)
	) name1011 (
		_w1051_,
		_w1053_,
		_w1745_,
		_w1746_
	);
	LUT4 #(
		.INIT('h00ae)
	) name1012 (
		_w1658_,
		_w1742_,
		_w1744_,
		_w1746_,
		_w1747_
	);
	LUT3 #(
		.INIT('h10)
	) name1013 (
		\u0_u0_ch_adr1_r_reg[21]/P0001 ,
		\u2_mast0_drdy_r_reg/P0001 ,
		\u2_state_reg[7]/NET0131 ,
		_w1748_
	);
	LUT2 #(
		.INIT('h1)
	) name1014 (
		\u0_u0_ch_adr1_r_reg[21]/P0001 ,
		\u2_state_reg[7]/NET0131 ,
		_w1749_
	);
	LUT3 #(
		.INIT('h23)
	) name1015 (
		_w1090_,
		_w1748_,
		_w1749_,
		_w1750_
	);
	LUT4 #(
		.INIT('h0053)
	) name1016 (
		\u2_adr1_cnt_reg[21]/P0001 ,
		\u3_u0_mast_dout_reg[23]/P0001 ,
		_w895_,
		_w1659_,
		_w1751_
	);
	LUT3 #(
		.INIT('he0)
	) name1017 (
		\u2_state_reg[7]/NET0131 ,
		_w1090_,
		_w1751_,
		_w1752_
	);
	LUT3 #(
		.INIT('h20)
	) name1018 (
		\u3_u1_slv_adr_reg[4]/NET0131 ,
		\u3_u1_slv_dout_reg[23]/P0001 ,
		\u3_u1_slv_we_reg/P0001 ,
		_w1753_
	);
	LUT3 #(
		.INIT('h80)
	) name1019 (
		_w1051_,
		_w1053_,
		_w1753_,
		_w1754_
	);
	LUT4 #(
		.INIT('h00ae)
	) name1020 (
		_w1658_,
		_w1750_,
		_w1752_,
		_w1754_,
		_w1755_
	);
	LUT3 #(
		.INIT('h10)
	) name1021 (
		\u0_u0_ch_adr1_r_reg[22]/P0001 ,
		\u2_mast0_drdy_r_reg/P0001 ,
		\u2_state_reg[7]/NET0131 ,
		_w1756_
	);
	LUT2 #(
		.INIT('h1)
	) name1022 (
		\u0_u0_ch_adr1_r_reg[22]/P0001 ,
		\u2_state_reg[7]/NET0131 ,
		_w1757_
	);
	LUT3 #(
		.INIT('h23)
	) name1023 (
		_w1090_,
		_w1756_,
		_w1757_,
		_w1758_
	);
	LUT4 #(
		.INIT('h0053)
	) name1024 (
		\u2_adr1_cnt_reg[22]/P0001 ,
		\u3_u0_mast_dout_reg[24]/P0001 ,
		_w895_,
		_w1659_,
		_w1759_
	);
	LUT3 #(
		.INIT('he0)
	) name1025 (
		\u2_state_reg[7]/NET0131 ,
		_w1090_,
		_w1759_,
		_w1760_
	);
	LUT3 #(
		.INIT('h20)
	) name1026 (
		\u3_u1_slv_adr_reg[4]/NET0131 ,
		\u3_u1_slv_dout_reg[24]/P0001 ,
		\u3_u1_slv_we_reg/P0001 ,
		_w1761_
	);
	LUT3 #(
		.INIT('h80)
	) name1027 (
		_w1051_,
		_w1053_,
		_w1761_,
		_w1762_
	);
	LUT4 #(
		.INIT('h00ae)
	) name1028 (
		_w1658_,
		_w1758_,
		_w1760_,
		_w1762_,
		_w1763_
	);
	LUT3 #(
		.INIT('h10)
	) name1029 (
		\u0_u0_ch_adr1_r_reg[23]/P0001 ,
		\u2_mast0_drdy_r_reg/P0001 ,
		\u2_state_reg[7]/NET0131 ,
		_w1764_
	);
	LUT2 #(
		.INIT('h1)
	) name1030 (
		\u0_u0_ch_adr1_r_reg[23]/P0001 ,
		\u2_state_reg[7]/NET0131 ,
		_w1765_
	);
	LUT3 #(
		.INIT('h23)
	) name1031 (
		_w1090_,
		_w1764_,
		_w1765_,
		_w1766_
	);
	LUT4 #(
		.INIT('h0053)
	) name1032 (
		\u2_adr1_cnt_reg[23]/P0001 ,
		\u3_u0_mast_dout_reg[25]/P0001 ,
		_w895_,
		_w1659_,
		_w1767_
	);
	LUT3 #(
		.INIT('he0)
	) name1033 (
		\u2_state_reg[7]/NET0131 ,
		_w1090_,
		_w1767_,
		_w1768_
	);
	LUT3 #(
		.INIT('h20)
	) name1034 (
		\u3_u1_slv_adr_reg[4]/NET0131 ,
		\u3_u1_slv_dout_reg[25]/P0001 ,
		\u3_u1_slv_we_reg/P0001 ,
		_w1769_
	);
	LUT3 #(
		.INIT('h80)
	) name1035 (
		_w1051_,
		_w1053_,
		_w1769_,
		_w1770_
	);
	LUT4 #(
		.INIT('h00ae)
	) name1036 (
		_w1658_,
		_w1766_,
		_w1768_,
		_w1770_,
		_w1771_
	);
	LUT3 #(
		.INIT('h10)
	) name1037 (
		\u0_u0_ch_adr1_r_reg[24]/P0001 ,
		\u2_mast0_drdy_r_reg/P0001 ,
		\u2_state_reg[7]/NET0131 ,
		_w1772_
	);
	LUT2 #(
		.INIT('h1)
	) name1038 (
		\u0_u0_ch_adr1_r_reg[24]/P0001 ,
		\u2_state_reg[7]/NET0131 ,
		_w1773_
	);
	LUT3 #(
		.INIT('h23)
	) name1039 (
		_w1090_,
		_w1772_,
		_w1773_,
		_w1774_
	);
	LUT4 #(
		.INIT('h0053)
	) name1040 (
		\u2_adr1_cnt_reg[24]/P0001 ,
		\u3_u0_mast_dout_reg[26]/P0001 ,
		_w895_,
		_w1659_,
		_w1775_
	);
	LUT3 #(
		.INIT('he0)
	) name1041 (
		\u2_state_reg[7]/NET0131 ,
		_w1090_,
		_w1775_,
		_w1776_
	);
	LUT3 #(
		.INIT('h20)
	) name1042 (
		\u3_u1_slv_adr_reg[4]/NET0131 ,
		\u3_u1_slv_dout_reg[26]/P0001 ,
		\u3_u1_slv_we_reg/P0001 ,
		_w1777_
	);
	LUT3 #(
		.INIT('h80)
	) name1043 (
		_w1051_,
		_w1053_,
		_w1777_,
		_w1778_
	);
	LUT4 #(
		.INIT('h00ae)
	) name1044 (
		_w1658_,
		_w1774_,
		_w1776_,
		_w1778_,
		_w1779_
	);
	LUT3 #(
		.INIT('h10)
	) name1045 (
		\u0_u0_ch_adr1_r_reg[25]/P0001 ,
		\u2_mast0_drdy_r_reg/P0001 ,
		\u2_state_reg[7]/NET0131 ,
		_w1780_
	);
	LUT2 #(
		.INIT('h1)
	) name1046 (
		\u0_u0_ch_adr1_r_reg[25]/P0001 ,
		\u2_state_reg[7]/NET0131 ,
		_w1781_
	);
	LUT3 #(
		.INIT('h23)
	) name1047 (
		_w1090_,
		_w1780_,
		_w1781_,
		_w1782_
	);
	LUT4 #(
		.INIT('h0053)
	) name1048 (
		\u2_adr1_cnt_reg[25]/P0001 ,
		\u3_u0_mast_dout_reg[27]/P0001 ,
		_w895_,
		_w1659_,
		_w1783_
	);
	LUT3 #(
		.INIT('he0)
	) name1049 (
		\u2_state_reg[7]/NET0131 ,
		_w1090_,
		_w1783_,
		_w1784_
	);
	LUT3 #(
		.INIT('h20)
	) name1050 (
		\u3_u1_slv_adr_reg[4]/NET0131 ,
		\u3_u1_slv_dout_reg[27]/P0001 ,
		\u3_u1_slv_we_reg/P0001 ,
		_w1785_
	);
	LUT3 #(
		.INIT('h80)
	) name1051 (
		_w1051_,
		_w1053_,
		_w1785_,
		_w1786_
	);
	LUT4 #(
		.INIT('h00ae)
	) name1052 (
		_w1658_,
		_w1782_,
		_w1784_,
		_w1786_,
		_w1787_
	);
	LUT3 #(
		.INIT('h10)
	) name1053 (
		\u0_u0_ch_adr1_r_reg[26]/P0001 ,
		\u2_mast0_drdy_r_reg/P0001 ,
		\u2_state_reg[7]/NET0131 ,
		_w1788_
	);
	LUT2 #(
		.INIT('h1)
	) name1054 (
		\u0_u0_ch_adr1_r_reg[26]/P0001 ,
		\u2_state_reg[7]/NET0131 ,
		_w1789_
	);
	LUT3 #(
		.INIT('h23)
	) name1055 (
		_w1090_,
		_w1788_,
		_w1789_,
		_w1790_
	);
	LUT4 #(
		.INIT('h0053)
	) name1056 (
		\u2_adr1_cnt_reg[26]/P0001 ,
		\u3_u0_mast_dout_reg[28]/P0001 ,
		_w895_,
		_w1659_,
		_w1791_
	);
	LUT3 #(
		.INIT('he0)
	) name1057 (
		\u2_state_reg[7]/NET0131 ,
		_w1090_,
		_w1791_,
		_w1792_
	);
	LUT3 #(
		.INIT('h20)
	) name1058 (
		\u3_u1_slv_adr_reg[4]/NET0131 ,
		\u3_u1_slv_dout_reg[28]/P0001 ,
		\u3_u1_slv_we_reg/P0001 ,
		_w1793_
	);
	LUT3 #(
		.INIT('h80)
	) name1059 (
		_w1051_,
		_w1053_,
		_w1793_,
		_w1794_
	);
	LUT4 #(
		.INIT('h00ae)
	) name1060 (
		_w1658_,
		_w1790_,
		_w1792_,
		_w1794_,
		_w1795_
	);
	LUT3 #(
		.INIT('h10)
	) name1061 (
		\u0_u0_ch_adr1_r_reg[27]/P0001 ,
		\u2_mast0_drdy_r_reg/P0001 ,
		\u2_state_reg[7]/NET0131 ,
		_w1796_
	);
	LUT2 #(
		.INIT('h1)
	) name1062 (
		\u0_u0_ch_adr1_r_reg[27]/P0001 ,
		\u2_state_reg[7]/NET0131 ,
		_w1797_
	);
	LUT3 #(
		.INIT('h23)
	) name1063 (
		_w1090_,
		_w1796_,
		_w1797_,
		_w1798_
	);
	LUT4 #(
		.INIT('h0053)
	) name1064 (
		\u2_adr1_cnt_reg[27]/P0001 ,
		\u3_u0_mast_dout_reg[29]/P0001 ,
		_w895_,
		_w1659_,
		_w1799_
	);
	LUT3 #(
		.INIT('he0)
	) name1065 (
		\u2_state_reg[7]/NET0131 ,
		_w1090_,
		_w1799_,
		_w1800_
	);
	LUT3 #(
		.INIT('h20)
	) name1066 (
		\u3_u1_slv_adr_reg[4]/NET0131 ,
		\u3_u1_slv_dout_reg[29]/P0001 ,
		\u3_u1_slv_we_reg/P0001 ,
		_w1801_
	);
	LUT3 #(
		.INIT('h80)
	) name1067 (
		_w1051_,
		_w1053_,
		_w1801_,
		_w1802_
	);
	LUT4 #(
		.INIT('h00ae)
	) name1068 (
		_w1658_,
		_w1798_,
		_w1800_,
		_w1802_,
		_w1803_
	);
	LUT3 #(
		.INIT('h10)
	) name1069 (
		\u0_u0_ch_adr1_r_reg[28]/P0001 ,
		\u2_mast0_drdy_r_reg/P0001 ,
		\u2_state_reg[7]/NET0131 ,
		_w1804_
	);
	LUT2 #(
		.INIT('h1)
	) name1070 (
		\u0_u0_ch_adr1_r_reg[28]/P0001 ,
		\u2_state_reg[7]/NET0131 ,
		_w1805_
	);
	LUT3 #(
		.INIT('h23)
	) name1071 (
		_w1090_,
		_w1804_,
		_w1805_,
		_w1806_
	);
	LUT4 #(
		.INIT('h0053)
	) name1072 (
		\u2_adr1_cnt_reg[28]/P0001 ,
		\u3_u0_mast_dout_reg[30]/P0001 ,
		_w895_,
		_w1659_,
		_w1807_
	);
	LUT3 #(
		.INIT('he0)
	) name1073 (
		\u2_state_reg[7]/NET0131 ,
		_w1090_,
		_w1807_,
		_w1808_
	);
	LUT3 #(
		.INIT('h20)
	) name1074 (
		\u3_u1_slv_adr_reg[4]/NET0131 ,
		\u3_u1_slv_dout_reg[30]/P0001 ,
		\u3_u1_slv_we_reg/P0001 ,
		_w1809_
	);
	LUT3 #(
		.INIT('h80)
	) name1075 (
		_w1051_,
		_w1053_,
		_w1809_,
		_w1810_
	);
	LUT4 #(
		.INIT('h00ae)
	) name1076 (
		_w1658_,
		_w1806_,
		_w1808_,
		_w1810_,
		_w1811_
	);
	LUT3 #(
		.INIT('h10)
	) name1077 (
		\u0_u0_ch_adr1_r_reg[29]/P0001 ,
		\u2_mast0_drdy_r_reg/P0001 ,
		\u2_state_reg[7]/NET0131 ,
		_w1812_
	);
	LUT2 #(
		.INIT('h1)
	) name1078 (
		\u0_u0_ch_adr1_r_reg[29]/P0001 ,
		\u2_state_reg[7]/NET0131 ,
		_w1813_
	);
	LUT3 #(
		.INIT('h23)
	) name1079 (
		_w1090_,
		_w1812_,
		_w1813_,
		_w1814_
	);
	LUT4 #(
		.INIT('h0053)
	) name1080 (
		\u2_adr1_cnt_reg[29]/P0001 ,
		\u3_u0_mast_dout_reg[31]/P0001 ,
		_w895_,
		_w1659_,
		_w1815_
	);
	LUT3 #(
		.INIT('he0)
	) name1081 (
		\u2_state_reg[7]/NET0131 ,
		_w1090_,
		_w1815_,
		_w1816_
	);
	LUT3 #(
		.INIT('h20)
	) name1082 (
		\u3_u1_slv_adr_reg[4]/NET0131 ,
		\u3_u1_slv_dout_reg[31]/P0001 ,
		\u3_u1_slv_we_reg/P0001 ,
		_w1817_
	);
	LUT3 #(
		.INIT('h80)
	) name1083 (
		_w1051_,
		_w1053_,
		_w1817_,
		_w1818_
	);
	LUT4 #(
		.INIT('h00ae)
	) name1084 (
		_w1658_,
		_w1814_,
		_w1816_,
		_w1818_,
		_w1819_
	);
	LUT3 #(
		.INIT('h02)
	) name1085 (
		\u2_state_reg[4]/NET0131 ,
		\u2_state_reg[6]/NET0131 ,
		\u2_state_reg[7]/NET0131 ,
		_w1820_
	);
	LUT4 #(
		.INIT('h8000)
	) name1086 (
		_w861_,
		_w899_,
		_w900_,
		_w1820_,
		_w1821_
	);
	LUT3 #(
		.INIT('h2a)
	) name1087 (
		\u0_u0_ch_csr_r_reg[1]/NET0131 ,
		\u2_mast0_drdy_r_reg/P0001 ,
		\u2_state_reg[5]/NET0131 ,
		_w1822_
	);
	LUT3 #(
		.INIT('h10)
	) name1088 (
		_w1057_,
		_w1821_,
		_w1822_,
		_w1823_
	);
	LUT4 #(
		.INIT('h2aaa)
	) name1089 (
		\u3_u0_mast_dout_reg[16]/P0001 ,
		_w1051_,
		_w1053_,
		_w1054_,
		_w1824_
	);
	LUT3 #(
		.INIT('he0)
	) name1090 (
		_w1257_,
		_w1821_,
		_w1824_,
		_w1825_
	);
	LUT3 #(
		.INIT('h40)
	) name1091 (
		\u3_u1_slv_adr_reg[4]/NET0131 ,
		\u3_u1_slv_dout_reg[1]/P0001 ,
		\u3_u1_slv_we_reg/P0001 ,
		_w1826_
	);
	LUT3 #(
		.INIT('h80)
	) name1092 (
		_w1051_,
		_w1053_,
		_w1826_,
		_w1827_
	);
	LUT3 #(
		.INIT('hfe)
	) name1093 (
		_w1823_,
		_w1825_,
		_w1827_,
		_w1828_
	);
	LUT3 #(
		.INIT('h2a)
	) name1094 (
		\u0_u0_ch_csr_r_reg[2]/NET0131 ,
		\u2_mast0_drdy_r_reg/P0001 ,
		\u2_state_reg[5]/NET0131 ,
		_w1829_
	);
	LUT3 #(
		.INIT('h10)
	) name1095 (
		_w1057_,
		_w1821_,
		_w1829_,
		_w1830_
	);
	LUT4 #(
		.INIT('h2aaa)
	) name1096 (
		\u3_u0_mast_dout_reg[17]/P0001 ,
		_w1051_,
		_w1053_,
		_w1054_,
		_w1831_
	);
	LUT3 #(
		.INIT('he0)
	) name1097 (
		_w1257_,
		_w1821_,
		_w1831_,
		_w1832_
	);
	LUT3 #(
		.INIT('h40)
	) name1098 (
		\u3_u1_slv_adr_reg[4]/NET0131 ,
		\u3_u1_slv_dout_reg[2]/P0001 ,
		\u3_u1_slv_we_reg/P0001 ,
		_w1833_
	);
	LUT3 #(
		.INIT('h80)
	) name1099 (
		_w1051_,
		_w1053_,
		_w1833_,
		_w1834_
	);
	LUT3 #(
		.INIT('hfe)
	) name1100 (
		_w1830_,
		_w1832_,
		_w1834_,
		_w1835_
	);
	LUT3 #(
		.INIT('h2a)
	) name1101 (
		\u0_u0_ch_csr_r_reg[3]/NET0131 ,
		\u2_mast0_drdy_r_reg/P0001 ,
		\u2_state_reg[5]/NET0131 ,
		_w1836_
	);
	LUT3 #(
		.INIT('h10)
	) name1102 (
		_w1057_,
		_w1821_,
		_w1836_,
		_w1837_
	);
	LUT4 #(
		.INIT('h2aaa)
	) name1103 (
		\u3_u0_mast_dout_reg[18]/P0001 ,
		_w1051_,
		_w1053_,
		_w1054_,
		_w1838_
	);
	LUT3 #(
		.INIT('he0)
	) name1104 (
		_w1257_,
		_w1821_,
		_w1838_,
		_w1839_
	);
	LUT3 #(
		.INIT('h40)
	) name1105 (
		\u3_u1_slv_adr_reg[4]/NET0131 ,
		\u3_u1_slv_dout_reg[3]/P0001 ,
		\u3_u1_slv_we_reg/P0001 ,
		_w1840_
	);
	LUT3 #(
		.INIT('h80)
	) name1106 (
		_w1051_,
		_w1053_,
		_w1840_,
		_w1841_
	);
	LUT3 #(
		.INIT('hfe)
	) name1107 (
		_w1837_,
		_w1839_,
		_w1841_,
		_w1842_
	);
	LUT3 #(
		.INIT('h2a)
	) name1108 (
		\u0_u0_ch_csr_r_reg[4]/NET0131 ,
		\u2_mast0_drdy_r_reg/P0001 ,
		\u2_state_reg[5]/NET0131 ,
		_w1843_
	);
	LUT3 #(
		.INIT('h10)
	) name1109 (
		_w1057_,
		_w1821_,
		_w1843_,
		_w1844_
	);
	LUT4 #(
		.INIT('h2aaa)
	) name1110 (
		\u3_u0_mast_dout_reg[19]/P0001 ,
		_w1051_,
		_w1053_,
		_w1054_,
		_w1845_
	);
	LUT3 #(
		.INIT('he0)
	) name1111 (
		_w1257_,
		_w1821_,
		_w1845_,
		_w1846_
	);
	LUT3 #(
		.INIT('h40)
	) name1112 (
		\u3_u1_slv_adr_reg[4]/NET0131 ,
		\u3_u1_slv_dout_reg[4]/P0001 ,
		\u3_u1_slv_we_reg/P0001 ,
		_w1847_
	);
	LUT3 #(
		.INIT('h80)
	) name1113 (
		_w1051_,
		_w1053_,
		_w1847_,
		_w1848_
	);
	LUT3 #(
		.INIT('hfe)
	) name1114 (
		_w1844_,
		_w1846_,
		_w1848_,
		_w1849_
	);
	LUT3 #(
		.INIT('h53)
	) name1115 (
		\u2_adr1_cnt_reg[0]/P0001 ,
		\u3_u0_mast_dout_reg[2]/P0001 ,
		_w895_,
		_w1850_
	);
	LUT4 #(
		.INIT('h007f)
	) name1116 (
		_w1051_,
		_w1053_,
		_w1657_,
		_w1659_,
		_w1851_
	);
	LUT4 #(
		.INIT('h0e00)
	) name1117 (
		\u2_state_reg[7]/NET0131 ,
		_w1090_,
		_w1850_,
		_w1851_,
		_w1852_
	);
	LUT3 #(
		.INIT('h80)
	) name1118 (
		\u3_u1_slv_adr_reg[4]/NET0131 ,
		\u3_u1_slv_dout_reg[2]/P0001 ,
		\u3_u1_slv_we_reg/P0001 ,
		_w1853_
	);
	LUT3 #(
		.INIT('h80)
	) name1119 (
		_w1051_,
		_w1053_,
		_w1853_,
		_w1854_
	);
	LUT4 #(
		.INIT('h2aaa)
	) name1120 (
		\u0_u0_ch_adr1_r_reg[0]/P0001 ,
		_w1051_,
		_w1053_,
		_w1657_,
		_w1855_
	);
	LUT4 #(
		.INIT('h4700)
	) name1121 (
		\u2_mast0_drdy_r_reg/P0001 ,
		\u2_state_reg[7]/NET0131 ,
		_w1090_,
		_w1855_,
		_w1856_
	);
	LUT3 #(
		.INIT('hfe)
	) name1122 (
		_w1852_,
		_w1854_,
		_w1856_,
		_w1857_
	);
	LUT3 #(
		.INIT('h53)
	) name1123 (
		\u2_adr1_cnt_reg[2]/P0001 ,
		\u3_u0_mast_dout_reg[4]/P0001 ,
		_w895_,
		_w1858_
	);
	LUT4 #(
		.INIT('h00e0)
	) name1124 (
		\u2_state_reg[7]/NET0131 ,
		_w1090_,
		_w1851_,
		_w1858_,
		_w1859_
	);
	LUT3 #(
		.INIT('h80)
	) name1125 (
		\u3_u1_slv_adr_reg[4]/NET0131 ,
		\u3_u1_slv_dout_reg[4]/P0001 ,
		\u3_u1_slv_we_reg/P0001 ,
		_w1860_
	);
	LUT3 #(
		.INIT('h80)
	) name1126 (
		_w1051_,
		_w1053_,
		_w1860_,
		_w1861_
	);
	LUT4 #(
		.INIT('h2aaa)
	) name1127 (
		\u0_u0_ch_adr1_r_reg[2]/P0001 ,
		_w1051_,
		_w1053_,
		_w1657_,
		_w1862_
	);
	LUT4 #(
		.INIT('h4700)
	) name1128 (
		\u2_mast0_drdy_r_reg/P0001 ,
		\u2_state_reg[7]/NET0131 ,
		_w1090_,
		_w1862_,
		_w1863_
	);
	LUT3 #(
		.INIT('hfe)
	) name1129 (
		_w1859_,
		_w1861_,
		_w1863_,
		_w1864_
	);
	LUT3 #(
		.INIT('h53)
	) name1130 (
		\u2_adr1_cnt_reg[1]/P0001 ,
		\u3_u0_mast_dout_reg[3]/P0001 ,
		_w895_,
		_w1865_
	);
	LUT4 #(
		.INIT('h00e0)
	) name1131 (
		\u2_state_reg[7]/NET0131 ,
		_w1090_,
		_w1851_,
		_w1865_,
		_w1866_
	);
	LUT3 #(
		.INIT('h80)
	) name1132 (
		\u3_u1_slv_adr_reg[4]/NET0131 ,
		\u3_u1_slv_dout_reg[3]/P0001 ,
		\u3_u1_slv_we_reg/P0001 ,
		_w1867_
	);
	LUT3 #(
		.INIT('h80)
	) name1133 (
		_w1051_,
		_w1053_,
		_w1867_,
		_w1868_
	);
	LUT4 #(
		.INIT('h2aaa)
	) name1134 (
		\u0_u0_ch_adr1_r_reg[1]/P0001 ,
		_w1051_,
		_w1053_,
		_w1657_,
		_w1869_
	);
	LUT4 #(
		.INIT('h4700)
	) name1135 (
		\u2_mast0_drdy_r_reg/P0001 ,
		\u2_state_reg[7]/NET0131 ,
		_w1090_,
		_w1869_,
		_w1870_
	);
	LUT3 #(
		.INIT('hfe)
	) name1136 (
		_w1866_,
		_w1868_,
		_w1870_,
		_w1871_
	);
	LUT3 #(
		.INIT('h53)
	) name1137 (
		\u2_adr1_cnt_reg[3]/P0001 ,
		\u3_u0_mast_dout_reg[5]/P0001 ,
		_w895_,
		_w1872_
	);
	LUT4 #(
		.INIT('h00e0)
	) name1138 (
		\u2_state_reg[7]/NET0131 ,
		_w1090_,
		_w1851_,
		_w1872_,
		_w1873_
	);
	LUT3 #(
		.INIT('h80)
	) name1139 (
		\u3_u1_slv_adr_reg[4]/NET0131 ,
		\u3_u1_slv_dout_reg[5]/P0001 ,
		\u3_u1_slv_we_reg/P0001 ,
		_w1874_
	);
	LUT3 #(
		.INIT('h80)
	) name1140 (
		_w1051_,
		_w1053_,
		_w1874_,
		_w1875_
	);
	LUT4 #(
		.INIT('h2aaa)
	) name1141 (
		\u0_u0_ch_adr1_r_reg[3]/P0001 ,
		_w1051_,
		_w1053_,
		_w1657_,
		_w1876_
	);
	LUT4 #(
		.INIT('h4700)
	) name1142 (
		\u2_mast0_drdy_r_reg/P0001 ,
		\u2_state_reg[7]/NET0131 ,
		_w1090_,
		_w1876_,
		_w1877_
	);
	LUT3 #(
		.INIT('hfe)
	) name1143 (
		_w1873_,
		_w1875_,
		_w1877_,
		_w1878_
	);
	LUT3 #(
		.INIT('h53)
	) name1144 (
		\u2_adr1_cnt_reg[4]/P0001 ,
		\u3_u0_mast_dout_reg[6]/P0001 ,
		_w895_,
		_w1879_
	);
	LUT4 #(
		.INIT('h00e0)
	) name1145 (
		\u2_state_reg[7]/NET0131 ,
		_w1090_,
		_w1851_,
		_w1879_,
		_w1880_
	);
	LUT3 #(
		.INIT('h80)
	) name1146 (
		\u3_u1_slv_adr_reg[4]/NET0131 ,
		\u3_u1_slv_dout_reg[6]/P0001 ,
		\u3_u1_slv_we_reg/P0001 ,
		_w1881_
	);
	LUT3 #(
		.INIT('h80)
	) name1147 (
		_w1051_,
		_w1053_,
		_w1881_,
		_w1882_
	);
	LUT4 #(
		.INIT('h2aaa)
	) name1148 (
		\u0_u0_ch_adr1_r_reg[4]/P0001 ,
		_w1051_,
		_w1053_,
		_w1657_,
		_w1883_
	);
	LUT4 #(
		.INIT('h4700)
	) name1149 (
		\u2_mast0_drdy_r_reg/P0001 ,
		\u2_state_reg[7]/NET0131 ,
		_w1090_,
		_w1883_,
		_w1884_
	);
	LUT3 #(
		.INIT('hfe)
	) name1150 (
		_w1880_,
		_w1882_,
		_w1884_,
		_w1885_
	);
	LUT3 #(
		.INIT('h53)
	) name1151 (
		\u2_adr1_cnt_reg[5]/P0001 ,
		\u3_u0_mast_dout_reg[7]/P0001 ,
		_w895_,
		_w1886_
	);
	LUT4 #(
		.INIT('h00e0)
	) name1152 (
		\u2_state_reg[7]/NET0131 ,
		_w1090_,
		_w1851_,
		_w1886_,
		_w1887_
	);
	LUT3 #(
		.INIT('h80)
	) name1153 (
		\u3_u1_slv_adr_reg[4]/NET0131 ,
		\u3_u1_slv_dout_reg[7]/P0001 ,
		\u3_u1_slv_we_reg/P0001 ,
		_w1888_
	);
	LUT3 #(
		.INIT('h80)
	) name1154 (
		_w1051_,
		_w1053_,
		_w1888_,
		_w1889_
	);
	LUT4 #(
		.INIT('h2aaa)
	) name1155 (
		\u0_u0_ch_adr1_r_reg[5]/P0001 ,
		_w1051_,
		_w1053_,
		_w1657_,
		_w1890_
	);
	LUT4 #(
		.INIT('h4700)
	) name1156 (
		\u2_mast0_drdy_r_reg/P0001 ,
		\u2_state_reg[7]/NET0131 ,
		_w1090_,
		_w1890_,
		_w1891_
	);
	LUT3 #(
		.INIT('hfe)
	) name1157 (
		_w1887_,
		_w1889_,
		_w1891_,
		_w1892_
	);
	LUT3 #(
		.INIT('h53)
	) name1158 (
		\u2_adr1_cnt_reg[6]/P0001 ,
		\u3_u0_mast_dout_reg[8]/P0001 ,
		_w895_,
		_w1893_
	);
	LUT4 #(
		.INIT('h00e0)
	) name1159 (
		\u2_state_reg[7]/NET0131 ,
		_w1090_,
		_w1851_,
		_w1893_,
		_w1894_
	);
	LUT3 #(
		.INIT('h80)
	) name1160 (
		\u3_u1_slv_adr_reg[4]/NET0131 ,
		\u3_u1_slv_dout_reg[8]/P0001 ,
		\u3_u1_slv_we_reg/P0001 ,
		_w1895_
	);
	LUT3 #(
		.INIT('h80)
	) name1161 (
		_w1051_,
		_w1053_,
		_w1895_,
		_w1896_
	);
	LUT4 #(
		.INIT('h2aaa)
	) name1162 (
		\u0_u0_ch_adr1_r_reg[6]/P0001 ,
		_w1051_,
		_w1053_,
		_w1657_,
		_w1897_
	);
	LUT4 #(
		.INIT('h4700)
	) name1163 (
		\u2_mast0_drdy_r_reg/P0001 ,
		\u2_state_reg[7]/NET0131 ,
		_w1090_,
		_w1897_,
		_w1898_
	);
	LUT3 #(
		.INIT('hfe)
	) name1164 (
		_w1894_,
		_w1896_,
		_w1898_,
		_w1899_
	);
	LUT3 #(
		.INIT('h53)
	) name1165 (
		\u2_adr1_cnt_reg[7]/P0001 ,
		\u3_u0_mast_dout_reg[9]/P0001 ,
		_w895_,
		_w1900_
	);
	LUT4 #(
		.INIT('h00e0)
	) name1166 (
		\u2_state_reg[7]/NET0131 ,
		_w1090_,
		_w1851_,
		_w1900_,
		_w1901_
	);
	LUT3 #(
		.INIT('h80)
	) name1167 (
		\u3_u1_slv_adr_reg[4]/NET0131 ,
		\u3_u1_slv_dout_reg[9]/P0001 ,
		\u3_u1_slv_we_reg/P0001 ,
		_w1902_
	);
	LUT3 #(
		.INIT('h80)
	) name1168 (
		_w1051_,
		_w1053_,
		_w1902_,
		_w1903_
	);
	LUT4 #(
		.INIT('h2aaa)
	) name1169 (
		\u0_u0_ch_adr1_r_reg[7]/P0001 ,
		_w1051_,
		_w1053_,
		_w1657_,
		_w1904_
	);
	LUT4 #(
		.INIT('h4700)
	) name1170 (
		\u2_mast0_drdy_r_reg/P0001 ,
		\u2_state_reg[7]/NET0131 ,
		_w1090_,
		_w1904_,
		_w1905_
	);
	LUT3 #(
		.INIT('hfe)
	) name1171 (
		_w1901_,
		_w1903_,
		_w1905_,
		_w1906_
	);
	LUT3 #(
		.INIT('h53)
	) name1172 (
		\u2_adr1_cnt_reg[8]/P0001 ,
		\u3_u0_mast_dout_reg[10]/P0001 ,
		_w895_,
		_w1907_
	);
	LUT4 #(
		.INIT('h00e0)
	) name1173 (
		\u2_state_reg[7]/NET0131 ,
		_w1090_,
		_w1851_,
		_w1907_,
		_w1908_
	);
	LUT3 #(
		.INIT('h80)
	) name1174 (
		\u3_u1_slv_adr_reg[4]/NET0131 ,
		\u3_u1_slv_dout_reg[10]/P0001 ,
		\u3_u1_slv_we_reg/P0001 ,
		_w1909_
	);
	LUT3 #(
		.INIT('h80)
	) name1175 (
		_w1051_,
		_w1053_,
		_w1909_,
		_w1910_
	);
	LUT4 #(
		.INIT('h2aaa)
	) name1176 (
		\u0_u0_ch_adr1_r_reg[8]/P0001 ,
		_w1051_,
		_w1053_,
		_w1657_,
		_w1911_
	);
	LUT4 #(
		.INIT('h4700)
	) name1177 (
		\u2_mast0_drdy_r_reg/P0001 ,
		\u2_state_reg[7]/NET0131 ,
		_w1090_,
		_w1911_,
		_w1912_
	);
	LUT3 #(
		.INIT('hfe)
	) name1178 (
		_w1908_,
		_w1910_,
		_w1912_,
		_w1913_
	);
	LUT3 #(
		.INIT('h53)
	) name1179 (
		\u2_adr1_cnt_reg[9]/P0001 ,
		\u3_u0_mast_dout_reg[11]/P0001 ,
		_w895_,
		_w1914_
	);
	LUT4 #(
		.INIT('h00e0)
	) name1180 (
		\u2_state_reg[7]/NET0131 ,
		_w1090_,
		_w1851_,
		_w1914_,
		_w1915_
	);
	LUT3 #(
		.INIT('h80)
	) name1181 (
		\u3_u1_slv_adr_reg[4]/NET0131 ,
		\u3_u1_slv_dout_reg[11]/P0001 ,
		\u3_u1_slv_we_reg/P0001 ,
		_w1916_
	);
	LUT3 #(
		.INIT('h80)
	) name1182 (
		_w1051_,
		_w1053_,
		_w1916_,
		_w1917_
	);
	LUT4 #(
		.INIT('h2aaa)
	) name1183 (
		\u0_u0_ch_adr1_r_reg[9]/P0001 ,
		_w1051_,
		_w1053_,
		_w1657_,
		_w1918_
	);
	LUT4 #(
		.INIT('h4700)
	) name1184 (
		\u2_mast0_drdy_r_reg/P0001 ,
		\u2_state_reg[7]/NET0131 ,
		_w1090_,
		_w1918_,
		_w1919_
	);
	LUT3 #(
		.INIT('hfe)
	) name1185 (
		_w1915_,
		_w1917_,
		_w1919_,
		_w1920_
	);
	LUT4 #(
		.INIT('h135f)
	) name1186 (
		\u0_int_maska_r_reg[27]/NET0131 ,
		\u0_int_maskb_r_reg[27]/NET0131 ,
		_w1411_,
		_w1413_,
		_w1921_
	);
	LUT3 #(
		.INIT('h80)
	) name1187 (
		\u0_u0_ch_adr1_r_reg[25]/P0001 ,
		_w1051_,
		_w1397_,
		_w1922_
	);
	LUT4 #(
		.INIT('h4000)
	) name1188 (
		_w1391_,
		_w1393_,
		_w1396_,
		_w1922_,
		_w1923_
	);
	LUT3 #(
		.INIT('h80)
	) name1189 (
		\u0_u0_ch_adr0_r_reg[25]/P0001 ,
		_w1051_,
		_w1397_,
		_w1924_
	);
	LUT4 #(
		.INIT('h0400)
	) name1190 (
		_w1391_,
		_w1393_,
		_w1396_,
		_w1924_,
		_w1925_
	);
	LUT3 #(
		.INIT('h01)
	) name1191 (
		_w1402_,
		_w1923_,
		_w1925_,
		_w1926_
	);
	LUT2 #(
		.INIT('h7)
	) name1192 (
		_w1921_,
		_w1926_,
		_w1927_
	);
	LUT4 #(
		.INIT('h135f)
	) name1193 (
		\u0_int_maska_r_reg[28]/NET0131 ,
		\u0_int_maskb_r_reg[28]/NET0131 ,
		_w1411_,
		_w1413_,
		_w1928_
	);
	LUT3 #(
		.INIT('h80)
	) name1194 (
		\u0_u0_ch_adr1_r_reg[26]/P0001 ,
		_w1051_,
		_w1397_,
		_w1929_
	);
	LUT4 #(
		.INIT('h4000)
	) name1195 (
		_w1391_,
		_w1393_,
		_w1396_,
		_w1929_,
		_w1930_
	);
	LUT3 #(
		.INIT('h80)
	) name1196 (
		\u0_u0_ch_adr0_r_reg[26]/P0001 ,
		_w1051_,
		_w1397_,
		_w1931_
	);
	LUT4 #(
		.INIT('h0400)
	) name1197 (
		_w1391_,
		_w1393_,
		_w1396_,
		_w1931_,
		_w1932_
	);
	LUT3 #(
		.INIT('h01)
	) name1198 (
		_w1402_,
		_w1930_,
		_w1932_,
		_w1933_
	);
	LUT2 #(
		.INIT('h7)
	) name1199 (
		_w1928_,
		_w1933_,
		_w1934_
	);
	LUT4 #(
		.INIT('h135f)
	) name1200 (
		\u0_int_maska_r_reg[29]/NET0131 ,
		\u0_int_maskb_r_reg[29]/NET0131 ,
		_w1411_,
		_w1413_,
		_w1935_
	);
	LUT3 #(
		.INIT('h80)
	) name1201 (
		\u0_u0_ch_adr1_r_reg[27]/P0001 ,
		_w1051_,
		_w1397_,
		_w1936_
	);
	LUT4 #(
		.INIT('h4000)
	) name1202 (
		_w1391_,
		_w1393_,
		_w1396_,
		_w1936_,
		_w1937_
	);
	LUT3 #(
		.INIT('h80)
	) name1203 (
		\u0_u0_ch_adr0_r_reg[27]/P0001 ,
		_w1051_,
		_w1397_,
		_w1938_
	);
	LUT4 #(
		.INIT('h0400)
	) name1204 (
		_w1391_,
		_w1393_,
		_w1396_,
		_w1938_,
		_w1939_
	);
	LUT3 #(
		.INIT('h01)
	) name1205 (
		_w1402_,
		_w1937_,
		_w1939_,
		_w1940_
	);
	LUT2 #(
		.INIT('h7)
	) name1206 (
		_w1935_,
		_w1940_,
		_w1941_
	);
	LUT4 #(
		.INIT('h135f)
	) name1207 (
		\u0_int_maska_r_reg[30]/NET0131 ,
		\u0_int_maskb_r_reg[30]/NET0131 ,
		_w1411_,
		_w1413_,
		_w1942_
	);
	LUT3 #(
		.INIT('h80)
	) name1208 (
		\u0_u0_ch_adr1_r_reg[28]/P0001 ,
		_w1051_,
		_w1397_,
		_w1943_
	);
	LUT4 #(
		.INIT('h4000)
	) name1209 (
		_w1391_,
		_w1393_,
		_w1396_,
		_w1943_,
		_w1944_
	);
	LUT3 #(
		.INIT('h80)
	) name1210 (
		\u0_u0_ch_adr0_r_reg[28]/P0001 ,
		_w1051_,
		_w1397_,
		_w1945_
	);
	LUT4 #(
		.INIT('h0400)
	) name1211 (
		_w1391_,
		_w1393_,
		_w1396_,
		_w1945_,
		_w1946_
	);
	LUT3 #(
		.INIT('h01)
	) name1212 (
		_w1402_,
		_w1944_,
		_w1946_,
		_w1947_
	);
	LUT2 #(
		.INIT('h7)
	) name1213 (
		_w1942_,
		_w1947_,
		_w1948_
	);
	LUT3 #(
		.INIT('h53)
	) name1214 (
		\u2_adr0_cnt_reg[9]/P0001 ,
		\u3_u0_mast_dout_reg[11]/P0001 ,
		_w895_,
		_w1949_
	);
	LUT4 #(
		.INIT('h0032)
	) name1215 (
		_w1090_,
		_w1515_,
		_w1516_,
		_w1949_,
		_w1950_
	);
	LUT3 #(
		.INIT('h40)
	) name1216 (
		\u3_u1_slv_adr_reg[2]/NET0131 ,
		\u3_u1_slv_adr_reg[3]/P0001 ,
		\u3_u1_slv_dout_reg[11]/P0001 ,
		_w1951_
	);
	LUT3 #(
		.INIT('h80)
	) name1217 (
		_w1051_,
		_w1252_,
		_w1951_,
		_w1952_
	);
	LUT4 #(
		.INIT('h2aaa)
	) name1218 (
		\u0_u0_ch_adr0_r_reg[9]/P0001 ,
		_w1051_,
		_w1252_,
		_w1514_,
		_w1953_
	);
	LUT4 #(
		.INIT('h0e0f)
	) name1219 (
		_w1090_,
		_w1516_,
		_w1952_,
		_w1953_,
		_w1954_
	);
	LUT2 #(
		.INIT('hb)
	) name1220 (
		_w1950_,
		_w1954_,
		_w1955_
	);
	LUT3 #(
		.INIT('h53)
	) name1221 (
		\u2_adr0_cnt_reg[0]/P0001 ,
		\u3_u0_mast_dout_reg[2]/P0001 ,
		_w895_,
		_w1956_
	);
	LUT4 #(
		.INIT('h0032)
	) name1222 (
		_w1090_,
		_w1515_,
		_w1516_,
		_w1956_,
		_w1957_
	);
	LUT3 #(
		.INIT('h40)
	) name1223 (
		\u3_u1_slv_adr_reg[2]/NET0131 ,
		\u3_u1_slv_adr_reg[3]/P0001 ,
		\u3_u1_slv_dout_reg[2]/P0001 ,
		_w1958_
	);
	LUT3 #(
		.INIT('h80)
	) name1224 (
		_w1051_,
		_w1252_,
		_w1958_,
		_w1959_
	);
	LUT4 #(
		.INIT('h2aaa)
	) name1225 (
		\u0_u0_ch_adr0_r_reg[0]/P0001 ,
		_w1051_,
		_w1252_,
		_w1514_,
		_w1960_
	);
	LUT4 #(
		.INIT('h0e0f)
	) name1226 (
		_w1090_,
		_w1516_,
		_w1959_,
		_w1960_,
		_w1961_
	);
	LUT2 #(
		.INIT('hb)
	) name1227 (
		_w1957_,
		_w1961_,
		_w1962_
	);
	LUT3 #(
		.INIT('h53)
	) name1228 (
		\u2_adr0_cnt_reg[1]/P0001 ,
		\u3_u0_mast_dout_reg[3]/P0001 ,
		_w895_,
		_w1963_
	);
	LUT4 #(
		.INIT('h0032)
	) name1229 (
		_w1090_,
		_w1515_,
		_w1516_,
		_w1963_,
		_w1964_
	);
	LUT3 #(
		.INIT('h40)
	) name1230 (
		\u3_u1_slv_adr_reg[2]/NET0131 ,
		\u3_u1_slv_adr_reg[3]/P0001 ,
		\u3_u1_slv_dout_reg[3]/P0001 ,
		_w1965_
	);
	LUT3 #(
		.INIT('h80)
	) name1231 (
		_w1051_,
		_w1252_,
		_w1965_,
		_w1966_
	);
	LUT4 #(
		.INIT('h2aaa)
	) name1232 (
		\u0_u0_ch_adr0_r_reg[1]/P0001 ,
		_w1051_,
		_w1252_,
		_w1514_,
		_w1967_
	);
	LUT4 #(
		.INIT('h0e0f)
	) name1233 (
		_w1090_,
		_w1516_,
		_w1966_,
		_w1967_,
		_w1968_
	);
	LUT2 #(
		.INIT('hb)
	) name1234 (
		_w1964_,
		_w1968_,
		_w1969_
	);
	LUT3 #(
		.INIT('h53)
	) name1235 (
		\u2_adr0_cnt_reg[2]/P0001 ,
		\u3_u0_mast_dout_reg[4]/P0001 ,
		_w895_,
		_w1970_
	);
	LUT4 #(
		.INIT('h0032)
	) name1236 (
		_w1090_,
		_w1515_,
		_w1516_,
		_w1970_,
		_w1971_
	);
	LUT3 #(
		.INIT('h40)
	) name1237 (
		\u3_u1_slv_adr_reg[2]/NET0131 ,
		\u3_u1_slv_adr_reg[3]/P0001 ,
		\u3_u1_slv_dout_reg[4]/P0001 ,
		_w1972_
	);
	LUT3 #(
		.INIT('h80)
	) name1238 (
		_w1051_,
		_w1252_,
		_w1972_,
		_w1973_
	);
	LUT4 #(
		.INIT('h2aaa)
	) name1239 (
		\u0_u0_ch_adr0_r_reg[2]/P0001 ,
		_w1051_,
		_w1252_,
		_w1514_,
		_w1974_
	);
	LUT4 #(
		.INIT('h0e0f)
	) name1240 (
		_w1090_,
		_w1516_,
		_w1973_,
		_w1974_,
		_w1975_
	);
	LUT2 #(
		.INIT('hb)
	) name1241 (
		_w1971_,
		_w1975_,
		_w1976_
	);
	LUT3 #(
		.INIT('h53)
	) name1242 (
		\u2_adr0_cnt_reg[3]/P0001 ,
		\u3_u0_mast_dout_reg[5]/P0001 ,
		_w895_,
		_w1977_
	);
	LUT4 #(
		.INIT('h0032)
	) name1243 (
		_w1090_,
		_w1515_,
		_w1516_,
		_w1977_,
		_w1978_
	);
	LUT3 #(
		.INIT('h40)
	) name1244 (
		\u3_u1_slv_adr_reg[2]/NET0131 ,
		\u3_u1_slv_adr_reg[3]/P0001 ,
		\u3_u1_slv_dout_reg[5]/P0001 ,
		_w1979_
	);
	LUT3 #(
		.INIT('h80)
	) name1245 (
		_w1051_,
		_w1252_,
		_w1979_,
		_w1980_
	);
	LUT4 #(
		.INIT('h2aaa)
	) name1246 (
		\u0_u0_ch_adr0_r_reg[3]/P0001 ,
		_w1051_,
		_w1252_,
		_w1514_,
		_w1981_
	);
	LUT4 #(
		.INIT('h0e0f)
	) name1247 (
		_w1090_,
		_w1516_,
		_w1980_,
		_w1981_,
		_w1982_
	);
	LUT2 #(
		.INIT('hb)
	) name1248 (
		_w1978_,
		_w1982_,
		_w1983_
	);
	LUT3 #(
		.INIT('h53)
	) name1249 (
		\u2_adr0_cnt_reg[4]/P0001 ,
		\u3_u0_mast_dout_reg[6]/P0001 ,
		_w895_,
		_w1984_
	);
	LUT4 #(
		.INIT('h0032)
	) name1250 (
		_w1090_,
		_w1515_,
		_w1516_,
		_w1984_,
		_w1985_
	);
	LUT3 #(
		.INIT('h40)
	) name1251 (
		\u3_u1_slv_adr_reg[2]/NET0131 ,
		\u3_u1_slv_adr_reg[3]/P0001 ,
		\u3_u1_slv_dout_reg[6]/P0001 ,
		_w1986_
	);
	LUT3 #(
		.INIT('h80)
	) name1252 (
		_w1051_,
		_w1252_,
		_w1986_,
		_w1987_
	);
	LUT4 #(
		.INIT('h2aaa)
	) name1253 (
		\u0_u0_ch_adr0_r_reg[4]/P0001 ,
		_w1051_,
		_w1252_,
		_w1514_,
		_w1988_
	);
	LUT4 #(
		.INIT('h0e0f)
	) name1254 (
		_w1090_,
		_w1516_,
		_w1987_,
		_w1988_,
		_w1989_
	);
	LUT2 #(
		.INIT('hb)
	) name1255 (
		_w1985_,
		_w1989_,
		_w1990_
	);
	LUT3 #(
		.INIT('h53)
	) name1256 (
		\u2_adr0_cnt_reg[5]/P0001 ,
		\u3_u0_mast_dout_reg[7]/P0001 ,
		_w895_,
		_w1991_
	);
	LUT4 #(
		.INIT('h0032)
	) name1257 (
		_w1090_,
		_w1515_,
		_w1516_,
		_w1991_,
		_w1992_
	);
	LUT3 #(
		.INIT('h40)
	) name1258 (
		\u3_u1_slv_adr_reg[2]/NET0131 ,
		\u3_u1_slv_adr_reg[3]/P0001 ,
		\u3_u1_slv_dout_reg[7]/P0001 ,
		_w1993_
	);
	LUT3 #(
		.INIT('h80)
	) name1259 (
		_w1051_,
		_w1252_,
		_w1993_,
		_w1994_
	);
	LUT4 #(
		.INIT('h2aaa)
	) name1260 (
		\u0_u0_ch_adr0_r_reg[5]/P0001 ,
		_w1051_,
		_w1252_,
		_w1514_,
		_w1995_
	);
	LUT4 #(
		.INIT('h0e0f)
	) name1261 (
		_w1090_,
		_w1516_,
		_w1994_,
		_w1995_,
		_w1996_
	);
	LUT2 #(
		.INIT('hb)
	) name1262 (
		_w1992_,
		_w1996_,
		_w1997_
	);
	LUT3 #(
		.INIT('h53)
	) name1263 (
		\u2_adr0_cnt_reg[6]/P0001 ,
		\u3_u0_mast_dout_reg[8]/P0001 ,
		_w895_,
		_w1998_
	);
	LUT4 #(
		.INIT('h0032)
	) name1264 (
		_w1090_,
		_w1515_,
		_w1516_,
		_w1998_,
		_w1999_
	);
	LUT3 #(
		.INIT('h40)
	) name1265 (
		\u3_u1_slv_adr_reg[2]/NET0131 ,
		\u3_u1_slv_adr_reg[3]/P0001 ,
		\u3_u1_slv_dout_reg[8]/P0001 ,
		_w2000_
	);
	LUT3 #(
		.INIT('h80)
	) name1266 (
		_w1051_,
		_w1252_,
		_w2000_,
		_w2001_
	);
	LUT4 #(
		.INIT('h2aaa)
	) name1267 (
		\u0_u0_ch_adr0_r_reg[6]/P0001 ,
		_w1051_,
		_w1252_,
		_w1514_,
		_w2002_
	);
	LUT4 #(
		.INIT('h0e0f)
	) name1268 (
		_w1090_,
		_w1516_,
		_w2001_,
		_w2002_,
		_w2003_
	);
	LUT2 #(
		.INIT('hb)
	) name1269 (
		_w1999_,
		_w2003_,
		_w2004_
	);
	LUT3 #(
		.INIT('h53)
	) name1270 (
		\u2_adr0_cnt_reg[7]/P0001 ,
		\u3_u0_mast_dout_reg[9]/P0001 ,
		_w895_,
		_w2005_
	);
	LUT4 #(
		.INIT('h0032)
	) name1271 (
		_w1090_,
		_w1515_,
		_w1516_,
		_w2005_,
		_w2006_
	);
	LUT3 #(
		.INIT('h40)
	) name1272 (
		\u3_u1_slv_adr_reg[2]/NET0131 ,
		\u3_u1_slv_adr_reg[3]/P0001 ,
		\u3_u1_slv_dout_reg[9]/P0001 ,
		_w2007_
	);
	LUT3 #(
		.INIT('h80)
	) name1273 (
		_w1051_,
		_w1252_,
		_w2007_,
		_w2008_
	);
	LUT4 #(
		.INIT('h2aaa)
	) name1274 (
		\u0_u0_ch_adr0_r_reg[7]/P0001 ,
		_w1051_,
		_w1252_,
		_w1514_,
		_w2009_
	);
	LUT4 #(
		.INIT('h0e0f)
	) name1275 (
		_w1090_,
		_w1516_,
		_w2008_,
		_w2009_,
		_w2010_
	);
	LUT2 #(
		.INIT('hb)
	) name1276 (
		_w2006_,
		_w2010_,
		_w2011_
	);
	LUT3 #(
		.INIT('h53)
	) name1277 (
		\u2_adr0_cnt_reg[8]/P0001 ,
		\u3_u0_mast_dout_reg[10]/P0001 ,
		_w895_,
		_w2012_
	);
	LUT4 #(
		.INIT('h0032)
	) name1278 (
		_w1090_,
		_w1515_,
		_w1516_,
		_w2012_,
		_w2013_
	);
	LUT3 #(
		.INIT('h40)
	) name1279 (
		\u3_u1_slv_adr_reg[2]/NET0131 ,
		\u3_u1_slv_adr_reg[3]/P0001 ,
		\u3_u1_slv_dout_reg[10]/P0001 ,
		_w2014_
	);
	LUT3 #(
		.INIT('h80)
	) name1280 (
		_w1051_,
		_w1252_,
		_w2014_,
		_w2015_
	);
	LUT4 #(
		.INIT('h2aaa)
	) name1281 (
		\u0_u0_ch_adr0_r_reg[8]/P0001 ,
		_w1051_,
		_w1252_,
		_w1514_,
		_w2016_
	);
	LUT4 #(
		.INIT('h0e0f)
	) name1282 (
		_w1090_,
		_w1516_,
		_w2015_,
		_w2016_,
		_w2017_
	);
	LUT2 #(
		.INIT('hb)
	) name1283 (
		_w2013_,
		_w2017_,
		_w2018_
	);
	LUT2 #(
		.INIT('h8)
	) name1284 (
		\u0_u0_ch_tot_sz_r_reg[11]/P0001 ,
		_w1408_,
		_w2019_
	);
	LUT3 #(
		.INIT('h80)
	) name1285 (
		\u0_u0_ch_adr0_r_reg[9]/P0001 ,
		_w1051_,
		_w1397_,
		_w2020_
	);
	LUT4 #(
		.INIT('h0400)
	) name1286 (
		_w1391_,
		_w1393_,
		_w1396_,
		_w2020_,
		_w2021_
	);
	LUT3 #(
		.INIT('h07)
	) name1287 (
		\u0_int_maskb_r_reg[11]/NET0131 ,
		_w1413_,
		_w2021_,
		_w2022_
	);
	LUT3 #(
		.INIT('h13)
	) name1288 (
		\u0_int_maska_r_reg[11]/NET0131 ,
		_w1402_,
		_w1411_,
		_w2023_
	);
	LUT3 #(
		.INIT('h80)
	) name1289 (
		\u0_u0_ch_adr1_r_reg[9]/P0001 ,
		_w1051_,
		_w1397_,
		_w2024_
	);
	LUT4 #(
		.INIT('h4000)
	) name1290 (
		_w1391_,
		_w1393_,
		_w1396_,
		_w2024_,
		_w2025_
	);
	LUT3 #(
		.INIT('h07)
	) name1291 (
		\u0_u0_ch_done_reg/P0002 ,
		_w1418_,
		_w2025_,
		_w2026_
	);
	LUT4 #(
		.INIT('hbfff)
	) name1292 (
		_w2019_,
		_w2022_,
		_w2023_,
		_w2026_,
		_w2027_
	);
	LUT2 #(
		.INIT('h8)
	) name1293 (
		\u0_u0_ch_csr_r2_reg[2]/NET0131 ,
		_w1418_,
		_w2028_
	);
	LUT4 #(
		.INIT('h135f)
	) name1294 (
		\u0_int_maska_r_reg[15]/NET0131 ,
		\u0_int_maskb_r_reg[15]/NET0131 ,
		_w1411_,
		_w1413_,
		_w2029_
	);
	LUT3 #(
		.INIT('h80)
	) name1295 (
		\u0_u0_ch_adr1_r_reg[13]/P0001 ,
		_w1051_,
		_w1397_,
		_w2030_
	);
	LUT4 #(
		.INIT('h4000)
	) name1296 (
		_w1391_,
		_w1393_,
		_w1396_,
		_w2030_,
		_w2031_
	);
	LUT2 #(
		.INIT('h1)
	) name1297 (
		_w1402_,
		_w2031_,
		_w2032_
	);
	LUT3 #(
		.INIT('h80)
	) name1298 (
		\u0_u0_ch_adr0_r_reg[13]/P0001 ,
		_w1051_,
		_w1397_,
		_w2033_
	);
	LUT4 #(
		.INIT('h0400)
	) name1299 (
		_w1391_,
		_w1393_,
		_w1396_,
		_w2033_,
		_w2034_
	);
	LUT3 #(
		.INIT('h07)
	) name1300 (
		\u0_u0_ch_sz_inf_reg/NET0131 ,
		_w1408_,
		_w2034_,
		_w2035_
	);
	LUT4 #(
		.INIT('hbfff)
	) name1301 (
		_w2028_,
		_w2029_,
		_w2032_,
		_w2035_,
		_w2036_
	);
	LUT2 #(
		.INIT('h8)
	) name1302 (
		\u0_int_maskb_r_reg[16]/NET0131 ,
		_w1413_,
		_w2037_
	);
	LUT4 #(
		.INIT('h53ff)
	) name1303 (
		\u0_int_maska_r_reg[16]/NET0131 ,
		\u0_u0_rest_en_reg/NET0131 ,
		_w1394_,
		_w1410_,
		_w2038_
	);
	LUT3 #(
		.INIT('h80)
	) name1304 (
		\u0_u0_ch_adr1_r_reg[14]/P0001 ,
		_w1051_,
		_w1397_,
		_w2039_
	);
	LUT4 #(
		.INIT('h4000)
	) name1305 (
		_w1391_,
		_w1393_,
		_w1396_,
		_w2039_,
		_w2040_
	);
	LUT2 #(
		.INIT('h1)
	) name1306 (
		_w1402_,
		_w2040_,
		_w2041_
	);
	LUT3 #(
		.INIT('h80)
	) name1307 (
		\u0_u0_ch_adr0_r_reg[14]/P0001 ,
		_w1051_,
		_w1397_,
		_w2042_
	);
	LUT4 #(
		.INIT('h0400)
	) name1308 (
		_w1391_,
		_w1393_,
		_w1396_,
		_w2042_,
		_w2043_
	);
	LUT3 #(
		.INIT('h07)
	) name1309 (
		\u0_u0_ch_chk_sz_r_reg[0]/P0001 ,
		_w1408_,
		_w2043_,
		_w2044_
	);
	LUT4 #(
		.INIT('hbfff)
	) name1310 (
		_w2037_,
		_w2038_,
		_w2041_,
		_w2044_,
		_w2045_
	);
	LUT3 #(
		.INIT('h80)
	) name1311 (
		\u0_u0_ch_adr1_r_reg[15]/P0001 ,
		_w1051_,
		_w1397_,
		_w2046_
	);
	LUT4 #(
		.INIT('h4000)
	) name1312 (
		_w1391_,
		_w1393_,
		_w1396_,
		_w2046_,
		_w2047_
	);
	LUT4 #(
		.INIT('h135f)
	) name1313 (
		\u0_int_maska_r_reg[17]/NET0131 ,
		\u0_int_maskb_r_reg[17]/NET0131 ,
		_w1411_,
		_w1413_,
		_w2048_
	);
	LUT3 #(
		.INIT('h13)
	) name1314 (
		\u0_u0_ch_chk_sz_r_reg[1]/P0001 ,
		_w1402_,
		_w1408_,
		_w2049_
	);
	LUT3 #(
		.INIT('h80)
	) name1315 (
		\u0_u0_ch_adr0_r_reg[15]/P0001 ,
		_w1051_,
		_w1397_,
		_w2050_
	);
	LUT4 #(
		.INIT('h0400)
	) name1316 (
		_w1391_,
		_w1393_,
		_w1396_,
		_w2050_,
		_w2051_
	);
	LUT3 #(
		.INIT('h07)
	) name1317 (
		\u0_u0_ch_csr_r3_reg[0]/NET0131 ,
		_w1418_,
		_w2051_,
		_w2052_
	);
	LUT4 #(
		.INIT('hbfff)
	) name1318 (
		_w2047_,
		_w2048_,
		_w2049_,
		_w2052_,
		_w2053_
	);
	LUT3 #(
		.INIT('h80)
	) name1319 (
		\u0_u0_ch_adr1_r_reg[16]/P0001 ,
		_w1051_,
		_w1397_,
		_w2054_
	);
	LUT4 #(
		.INIT('h4000)
	) name1320 (
		_w1391_,
		_w1393_,
		_w1396_,
		_w2054_,
		_w2055_
	);
	LUT4 #(
		.INIT('h135f)
	) name1321 (
		\u0_int_maska_r_reg[18]/NET0131 ,
		\u0_int_maskb_r_reg[18]/NET0131 ,
		_w1411_,
		_w1413_,
		_w2056_
	);
	LUT3 #(
		.INIT('h13)
	) name1322 (
		\u0_u0_ch_chk_sz_r_reg[2]/P0001 ,
		_w1402_,
		_w1408_,
		_w2057_
	);
	LUT3 #(
		.INIT('h80)
	) name1323 (
		\u0_u0_ch_adr0_r_reg[16]/P0001 ,
		_w1051_,
		_w1397_,
		_w2058_
	);
	LUT4 #(
		.INIT('h0400)
	) name1324 (
		_w1391_,
		_w1393_,
		_w1396_,
		_w2058_,
		_w2059_
	);
	LUT3 #(
		.INIT('h07)
	) name1325 (
		\u0_u0_ch_csr_r3_reg[1]/NET0131 ,
		_w1418_,
		_w2059_,
		_w2060_
	);
	LUT4 #(
		.INIT('hbfff)
	) name1326 (
		_w2055_,
		_w2056_,
		_w2057_,
		_w2060_,
		_w2061_
	);
	LUT3 #(
		.INIT('h80)
	) name1327 (
		\u0_u0_ch_adr1_r_reg[17]/P0001 ,
		_w1051_,
		_w1397_,
		_w2062_
	);
	LUT4 #(
		.INIT('h4000)
	) name1328 (
		_w1391_,
		_w1393_,
		_w1396_,
		_w2062_,
		_w2063_
	);
	LUT4 #(
		.INIT('h135f)
	) name1329 (
		\u0_int_maska_r_reg[19]/NET0131 ,
		\u0_int_maskb_r_reg[19]/NET0131 ,
		_w1411_,
		_w1413_,
		_w2064_
	);
	LUT3 #(
		.INIT('h13)
	) name1330 (
		\u0_u0_ch_chk_sz_r_reg[3]/P0001 ,
		_w1402_,
		_w1408_,
		_w2065_
	);
	LUT3 #(
		.INIT('h80)
	) name1331 (
		\u0_u0_ch_adr0_r_reg[17]/P0001 ,
		_w1051_,
		_w1397_,
		_w2066_
	);
	LUT4 #(
		.INIT('h0400)
	) name1332 (
		_w1391_,
		_w1393_,
		_w1396_,
		_w2066_,
		_w2067_
	);
	LUT3 #(
		.INIT('h07)
	) name1333 (
		\u0_u0_ch_csr_r3_reg[2]/NET0131 ,
		_w1418_,
		_w2067_,
		_w2068_
	);
	LUT4 #(
		.INIT('hbfff)
	) name1334 (
		_w2063_,
		_w2064_,
		_w2065_,
		_w2068_,
		_w2069_
	);
	LUT2 #(
		.INIT('h8)
	) name1335 (
		\u0_int_maskb_r_reg[20]/NET0131 ,
		_w1413_,
		_w2070_
	);
	LUT3 #(
		.INIT('h80)
	) name1336 (
		\u0_u0_ch_adr1_r_reg[18]/P0001 ,
		_w1051_,
		_w1397_,
		_w2071_
	);
	LUT4 #(
		.INIT('h4000)
	) name1337 (
		_w1391_,
		_w1393_,
		_w1396_,
		_w2071_,
		_w2072_
	);
	LUT3 #(
		.INIT('h07)
	) name1338 (
		\u0_int_maska_r_reg[20]/NET0131 ,
		_w1411_,
		_w2072_,
		_w2073_
	);
	LUT3 #(
		.INIT('h80)
	) name1339 (
		\u0_u0_ch_adr0_r_reg[18]/P0001 ,
		_w1051_,
		_w1397_,
		_w2074_
	);
	LUT4 #(
		.INIT('h0400)
	) name1340 (
		_w1391_,
		_w1393_,
		_w1396_,
		_w2074_,
		_w2075_
	);
	LUT3 #(
		.INIT('h07)
	) name1341 (
		\u0_u0_ch_chk_sz_r_reg[4]/P0001 ,
		_w1408_,
		_w2075_,
		_w2076_
	);
	LUT4 #(
		.INIT('hdfff)
	) name1342 (
		_w1419_,
		_w2070_,
		_w2073_,
		_w2076_,
		_w2077_
	);
	LUT3 #(
		.INIT('h80)
	) name1343 (
		\u0_u0_ch_adr1_r_reg[19]/P0001 ,
		_w1051_,
		_w1397_,
		_w2078_
	);
	LUT4 #(
		.INIT('h4000)
	) name1344 (
		_w1391_,
		_w1393_,
		_w1396_,
		_w2078_,
		_w2079_
	);
	LUT4 #(
		.INIT('h135f)
	) name1345 (
		\u0_int_maska_r_reg[21]/NET0131 ,
		\u0_int_maskb_r_reg[21]/NET0131 ,
		_w1411_,
		_w1413_,
		_w2080_
	);
	LUT3 #(
		.INIT('h13)
	) name1346 (
		\u0_u0_ch_chk_sz_r_reg[5]/P0001 ,
		_w1402_,
		_w1408_,
		_w2081_
	);
	LUT3 #(
		.INIT('h80)
	) name1347 (
		\u0_u0_ch_adr0_r_reg[19]/P0001 ,
		_w1051_,
		_w1397_,
		_w2082_
	);
	LUT4 #(
		.INIT('h0400)
	) name1348 (
		_w1391_,
		_w1393_,
		_w1396_,
		_w2082_,
		_w2083_
	);
	LUT3 #(
		.INIT('h07)
	) name1349 (
		\u0_u0_int_src_r_reg[1]/NET0131 ,
		_w1418_,
		_w2083_,
		_w2084_
	);
	LUT4 #(
		.INIT('hbfff)
	) name1350 (
		_w2079_,
		_w2080_,
		_w2081_,
		_w2084_,
		_w2085_
	);
	LUT3 #(
		.INIT('h80)
	) name1351 (
		\u0_u0_ch_adr1_r_reg[20]/P0001 ,
		_w1051_,
		_w1397_,
		_w2086_
	);
	LUT4 #(
		.INIT('h4000)
	) name1352 (
		_w1391_,
		_w1393_,
		_w1396_,
		_w2086_,
		_w2087_
	);
	LUT4 #(
		.INIT('h135f)
	) name1353 (
		\u0_int_maska_r_reg[22]/NET0131 ,
		\u0_int_maskb_r_reg[22]/NET0131 ,
		_w1411_,
		_w1413_,
		_w2088_
	);
	LUT3 #(
		.INIT('h13)
	) name1354 (
		\u0_u0_ch_chk_sz_r_reg[6]/P0001 ,
		_w1402_,
		_w1408_,
		_w2089_
	);
	LUT3 #(
		.INIT('h80)
	) name1355 (
		\u0_u0_ch_adr0_r_reg[20]/P0001 ,
		_w1051_,
		_w1397_,
		_w2090_
	);
	LUT4 #(
		.INIT('h0400)
	) name1356 (
		_w1391_,
		_w1393_,
		_w1396_,
		_w2090_,
		_w2091_
	);
	LUT3 #(
		.INIT('h07)
	) name1357 (
		\u0_u0_int_src_r_reg[2]/NET0131 ,
		_w1418_,
		_w2091_,
		_w2092_
	);
	LUT4 #(
		.INIT('hbfff)
	) name1358 (
		_w2087_,
		_w2088_,
		_w2089_,
		_w2092_,
		_w2093_
	);
	LUT3 #(
		.INIT('h80)
	) name1359 (
		\u0_u0_ch_adr0_r_reg[2]/P0001 ,
		_w1051_,
		_w1397_,
		_w2094_
	);
	LUT4 #(
		.INIT('h0400)
	) name1360 (
		_w1391_,
		_w1393_,
		_w1396_,
		_w2094_,
		_w2095_
	);
	LUT4 #(
		.INIT('h135f)
	) name1361 (
		\u0_int_maska_r_reg[4]/NET0131 ,
		\u0_int_maskb_r_reg[4]/NET0131 ,
		_w1411_,
		_w1413_,
		_w2096_
	);
	LUT3 #(
		.INIT('h13)
	) name1362 (
		\u0_u0_ch_csr_r_reg[4]/NET0131 ,
		_w1402_,
		_w1418_,
		_w2097_
	);
	LUT3 #(
		.INIT('h80)
	) name1363 (
		\u0_u0_ch_adr1_r_reg[2]/P0001 ,
		_w1051_,
		_w1397_,
		_w2098_
	);
	LUT4 #(
		.INIT('h4000)
	) name1364 (
		_w1391_,
		_w1393_,
		_w1396_,
		_w2098_,
		_w2099_
	);
	LUT3 #(
		.INIT('h07)
	) name1365 (
		\u0_u0_ch_tot_sz_r_reg[4]/P0001 ,
		_w1408_,
		_w2099_,
		_w2100_
	);
	LUT4 #(
		.INIT('hbfff)
	) name1366 (
		_w2095_,
		_w2096_,
		_w2097_,
		_w2100_,
		_w2101_
	);
	LUT2 #(
		.INIT('h8)
	) name1367 (
		\u0_u0_ch_tot_sz_r_reg[5]/P0001 ,
		_w1408_,
		_w2102_
	);
	LUT3 #(
		.INIT('h80)
	) name1368 (
		\u0_u0_ch_adr0_r_reg[3]/P0001 ,
		_w1051_,
		_w1397_,
		_w2103_
	);
	LUT4 #(
		.INIT('h0400)
	) name1369 (
		_w1391_,
		_w1393_,
		_w1396_,
		_w2103_,
		_w2104_
	);
	LUT3 #(
		.INIT('h07)
	) name1370 (
		\u0_int_maskb_r_reg[5]/NET0131 ,
		_w1413_,
		_w2104_,
		_w2105_
	);
	LUT3 #(
		.INIT('h13)
	) name1371 (
		\u0_u0_ch_csr_r_reg[5]/NET0131 ,
		_w1402_,
		_w1418_,
		_w2106_
	);
	LUT3 #(
		.INIT('h80)
	) name1372 (
		\u0_u0_ch_adr1_r_reg[3]/P0001 ,
		_w1051_,
		_w1397_,
		_w2107_
	);
	LUT4 #(
		.INIT('h4000)
	) name1373 (
		_w1391_,
		_w1393_,
		_w1396_,
		_w2107_,
		_w2108_
	);
	LUT3 #(
		.INIT('h07)
	) name1374 (
		\u0_int_maska_r_reg[5]/NET0131 ,
		_w1411_,
		_w2108_,
		_w2109_
	);
	LUT4 #(
		.INIT('hbfff)
	) name1375 (
		_w2102_,
		_w2105_,
		_w2106_,
		_w2109_,
		_w2110_
	);
	LUT2 #(
		.INIT('h8)
	) name1376 (
		\u0_u0_ch_tot_sz_r_reg[6]/P0001 ,
		_w1408_,
		_w2111_
	);
	LUT3 #(
		.INIT('h80)
	) name1377 (
		\u0_u0_ch_adr0_r_reg[4]/P0001 ,
		_w1051_,
		_w1397_,
		_w2112_
	);
	LUT4 #(
		.INIT('h0400)
	) name1378 (
		_w1391_,
		_w1393_,
		_w1396_,
		_w2112_,
		_w2113_
	);
	LUT3 #(
		.INIT('h07)
	) name1379 (
		\u0_int_maskb_r_reg[6]/NET0131 ,
		_w1413_,
		_w2113_,
		_w2114_
	);
	LUT3 #(
		.INIT('h13)
	) name1380 (
		\u0_u0_ch_csr_r_reg[6]/NET0131 ,
		_w1402_,
		_w1418_,
		_w2115_
	);
	LUT3 #(
		.INIT('h80)
	) name1381 (
		\u0_u0_ch_adr1_r_reg[4]/P0001 ,
		_w1051_,
		_w1397_,
		_w2116_
	);
	LUT4 #(
		.INIT('h4000)
	) name1382 (
		_w1391_,
		_w1393_,
		_w1396_,
		_w2116_,
		_w2117_
	);
	LUT3 #(
		.INIT('h07)
	) name1383 (
		\u0_int_maska_r_reg[6]/NET0131 ,
		_w1411_,
		_w2117_,
		_w2118_
	);
	LUT4 #(
		.INIT('hbfff)
	) name1384 (
		_w2111_,
		_w2114_,
		_w2115_,
		_w2118_,
		_w2119_
	);
	LUT2 #(
		.INIT('h8)
	) name1385 (
		\u0_u0_ch_tot_sz_r_reg[7]/P0001 ,
		_w1408_,
		_w2120_
	);
	LUT3 #(
		.INIT('h80)
	) name1386 (
		\u0_u0_ch_adr0_r_reg[5]/P0001 ,
		_w1051_,
		_w1397_,
		_w2121_
	);
	LUT4 #(
		.INIT('h0400)
	) name1387 (
		_w1391_,
		_w1393_,
		_w1396_,
		_w2121_,
		_w2122_
	);
	LUT3 #(
		.INIT('h07)
	) name1388 (
		\u0_int_maskb_r_reg[7]/NET0131 ,
		_w1413_,
		_w2122_,
		_w2123_
	);
	LUT3 #(
		.INIT('h13)
	) name1389 (
		\u0_u0_ch_csr_r_reg[7]/NET0131 ,
		_w1402_,
		_w1418_,
		_w2124_
	);
	LUT3 #(
		.INIT('h80)
	) name1390 (
		\u0_u0_ch_adr1_r_reg[5]/P0001 ,
		_w1051_,
		_w1397_,
		_w2125_
	);
	LUT4 #(
		.INIT('h4000)
	) name1391 (
		_w1391_,
		_w1393_,
		_w1396_,
		_w2125_,
		_w2126_
	);
	LUT3 #(
		.INIT('h07)
	) name1392 (
		\u0_int_maska_r_reg[7]/NET0131 ,
		_w1411_,
		_w2126_,
		_w2127_
	);
	LUT4 #(
		.INIT('hbfff)
	) name1393 (
		_w2120_,
		_w2123_,
		_w2124_,
		_w2127_,
		_w2128_
	);
	LUT2 #(
		.INIT('h8)
	) name1394 (
		\u0_u0_ch_tot_sz_r_reg[8]/P0001 ,
		_w1408_,
		_w2129_
	);
	LUT3 #(
		.INIT('h80)
	) name1395 (
		\u0_u0_ch_adr0_r_reg[6]/P0001 ,
		_w1051_,
		_w1397_,
		_w2130_
	);
	LUT4 #(
		.INIT('h0400)
	) name1396 (
		_w1391_,
		_w1393_,
		_w1396_,
		_w2130_,
		_w2131_
	);
	LUT3 #(
		.INIT('h07)
	) name1397 (
		\u0_int_maskb_r_reg[8]/NET0131 ,
		_w1413_,
		_w2131_,
		_w2132_
	);
	LUT3 #(
		.INIT('h13)
	) name1398 (
		\u0_int_maska_r_reg[8]/NET0131 ,
		_w1402_,
		_w1411_,
		_w2133_
	);
	LUT3 #(
		.INIT('h80)
	) name1399 (
		\u0_u0_ch_adr1_r_reg[6]/P0001 ,
		_w1051_,
		_w1397_,
		_w2134_
	);
	LUT4 #(
		.INIT('h4000)
	) name1400 (
		_w1391_,
		_w1393_,
		_w1396_,
		_w2134_,
		_w2135_
	);
	LUT3 #(
		.INIT('h07)
	) name1401 (
		\u0_u0_ch_csr_r_reg[8]/NET0131 ,
		_w1418_,
		_w2135_,
		_w2136_
	);
	LUT4 #(
		.INIT('hbfff)
	) name1402 (
		_w2129_,
		_w2132_,
		_w2133_,
		_w2136_,
		_w2137_
	);
	LUT3 #(
		.INIT('h80)
	) name1403 (
		\u0_u0_ch_adr0_r_reg[29]/P0001 ,
		_w1051_,
		_w1397_,
		_w2138_
	);
	LUT4 #(
		.INIT('h0400)
	) name1404 (
		_w1391_,
		_w1393_,
		_w1396_,
		_w2138_,
		_w2139_
	);
	LUT3 #(
		.INIT('h80)
	) name1405 (
		\u0_u0_ch_adr1_r_reg[29]/P0001 ,
		_w1051_,
		_w1397_,
		_w2140_
	);
	LUT4 #(
		.INIT('h4000)
	) name1406 (
		_w1391_,
		_w1393_,
		_w1396_,
		_w2140_,
		_w2141_
	);
	LUT3 #(
		.INIT('hfe)
	) name1407 (
		_w1402_,
		_w2139_,
		_w2141_,
		_w2142_
	);
	LUT4 #(
		.INIT('h153f)
	) name1408 (
		\u0_u0_ch_csr_r_reg[1]/NET0131 ,
		\u0_u0_ch_tot_sz_r_reg[1]/P0001 ,
		_w1408_,
		_w1418_,
		_w2143_
	);
	LUT4 #(
		.INIT('h135f)
	) name1409 (
		\u0_int_maska_r_reg[1]/NET0131 ,
		\u0_int_maskb_r_reg[1]/NET0131 ,
		_w1411_,
		_w1413_,
		_w2144_
	);
	LUT2 #(
		.INIT('h7)
	) name1410 (
		_w2143_,
		_w2144_,
		_w2145_
	);
	LUT2 #(
		.INIT('h1)
	) name1411 (
		\u0_u0_ch_err_reg/NET0131 ,
		\u2_dma_abort_r_reg/NET0131 ,
		_w2146_
	);
	LUT3 #(
		.INIT('h10)
	) name1412 (
		\u2_dma_abort_r_reg/NET0131 ,
		\u3_u1_slv_adr_reg[2]/NET0131 ,
		\u3_u1_slv_re_reg/P0001 ,
		_w2147_
	);
	LUT4 #(
		.INIT('h070f)
	) name1413 (
		_w1051_,
		_w1097_,
		_w2146_,
		_w2147_,
		_w2148_
	);
	LUT3 #(
		.INIT('h6a)
	) name1414 (
		\u2_adr0_cnt_reg[15]/P0001 ,
		_w1375_,
		_w1492_,
		_w2149_
	);
	LUT3 #(
		.INIT('h6a)
	) name1415 (
		\u2_adr1_cnt_reg[15]/P0001 ,
		_w1384_,
		_w1495_,
		_w2150_
	);
	LUT3 #(
		.INIT('h6c)
	) name1416 (
		\u2_adr0_cnt_reg[10]/P0001 ,
		\u2_adr0_cnt_reg[11]/P0001 ,
		_w1375_,
		_w2151_
	);
	LUT3 #(
		.INIT('h6c)
	) name1417 (
		\u2_adr1_cnt_reg[10]/P0001 ,
		\u2_adr1_cnt_reg[11]/P0001 ,
		_w1384_,
		_w2152_
	);
	LUT2 #(
		.INIT('h6)
	) name1418 (
		\u2_adr0_cnt_reg[4]/P0001 ,
		_w1372_,
		_w2153_
	);
	LUT2 #(
		.INIT('h6)
	) name1419 (
		\u2_adr1_cnt_reg[4]/P0001 ,
		_w1381_,
		_w2154_
	);
	LUT3 #(
		.INIT('hfe)
	) name1420 (
		\u0_u0_ch_stop_reg/P0001 ,
		\wb0_err_i_pad ,
		\wb1_err_i_pad ,
		_w2155_
	);
	LUT2 #(
		.INIT('h1)
	) name1421 (
		\u2_state_reg[7]/NET0131 ,
		\wb0_ack_i_pad ,
		_w2156_
	);
	LUT4 #(
		.INIT('h0080)
	) name1422 (
		_w1067_,
		_w1145_,
		_w1146_,
		_w2156_,
		_w2157_
	);
	LUT4 #(
		.INIT('h0004)
	) name1423 (
		\u2_state_reg[10]/NET0131 ,
		\u2_state_reg[7]/NET0131 ,
		\u2_state_reg[8]/NET0131 ,
		\u2_state_reg[9]/NET0131 ,
		_w2158_
	);
	LUT4 #(
		.INIT('h4000)
	) name1424 (
		\wb0_ack_i_pad ,
		_w865_,
		_w894_,
		_w2158_,
		_w2159_
	);
	LUT2 #(
		.INIT('he)
	) name1425 (
		_w2157_,
		_w2159_,
		_w2160_
	);
	LUT2 #(
		.INIT('h1)
	) name1426 (
		\u2_state_reg[5]/NET0131 ,
		\wb0_ack_i_pad ,
		_w2161_
	);
	LUT3 #(
		.INIT('h04)
	) name1427 (
		\u2_state_reg[4]/NET0131 ,
		\u2_state_reg[5]/NET0131 ,
		\u2_state_reg[6]/NET0131 ,
		_w2162_
	);
	LUT4 #(
		.INIT('h8000)
	) name1428 (
		_w861_,
		_w863_,
		_w2156_,
		_w2162_,
		_w2163_
	);
	LUT3 #(
		.INIT('h32)
	) name1429 (
		_w1204_,
		_w2161_,
		_w2163_,
		_w2164_
	);
	LUT4 #(
		.INIT('h8000)
	) name1430 (
		\wb0_ack_i_pad ,
		_w865_,
		_w894_,
		_w2158_,
		_w2165_
	);
	LUT3 #(
		.INIT('h32)
	) name1431 (
		\u2_state_reg[6]/NET0131 ,
		\u2_state_reg[7]/NET0131 ,
		\wb0_ack_i_pad ,
		_w2166_
	);
	LUT4 #(
		.INIT('h8000)
	) name1432 (
		_w861_,
		_w863_,
		_w2162_,
		_w2166_,
		_w2167_
	);
	LUT4 #(
		.INIT('h4000)
	) name1433 (
		\wb0_ack_i_pad ,
		_w1067_,
		_w1145_,
		_w1146_,
		_w2168_
	);
	LUT2 #(
		.INIT('he)
	) name1434 (
		_w2167_,
		_w2168_,
		_w2169_
	);
	LUT4 #(
		.INIT('h8000)
	) name1435 (
		\u2_adr0_cnt_reg[10]/P0001 ,
		\u2_adr0_cnt_reg[11]/P0001 ,
		\u2_adr0_cnt_reg[12]/P0001 ,
		\u2_adr0_cnt_reg[13]/P0001 ,
		_w2170_
	);
	LUT4 #(
		.INIT('h8000)
	) name1436 (
		_w1372_,
		_w1373_,
		_w1374_,
		_w2170_,
		_w2171_
	);
	LUT4 #(
		.INIT('h2e2a)
	) name1437 (
		\u2_adr0_cnt_reg[14]/P0001 ,
		_w1375_,
		_w1492_,
		_w2170_,
		_w2172_
	);
	LUT4 #(
		.INIT('h8000)
	) name1438 (
		\u2_adr1_cnt_reg[10]/P0001 ,
		\u2_adr1_cnt_reg[11]/P0001 ,
		\u2_adr1_cnt_reg[12]/P0001 ,
		\u2_adr1_cnt_reg[13]/P0001 ,
		_w2173_
	);
	LUT4 #(
		.INIT('h8000)
	) name1439 (
		_w1381_,
		_w1382_,
		_w1383_,
		_w2173_,
		_w2174_
	);
	LUT4 #(
		.INIT('h2e2a)
	) name1440 (
		\u2_adr1_cnt_reg[14]/P0001 ,
		_w1384_,
		_w1495_,
		_w2173_,
		_w2175_
	);
	LUT3 #(
		.INIT('h6a)
	) name1441 (
		\u2_adr0_cnt_reg[7]/P0001 ,
		_w1372_,
		_w1373_,
		_w2176_
	);
	LUT3 #(
		.INIT('h6a)
	) name1442 (
		\u2_adr1_cnt_reg[7]/P0001 ,
		_w1381_,
		_w1382_,
		_w2177_
	);
	LUT2 #(
		.INIT('h4)
	) name1443 (
		\u4_u1_rf_ack_reg/P0001 ,
		\wb1_stb_i_pad ,
		_w2178_
	);
	LUT3 #(
		.INIT('he0)
	) name1444 (
		\u4_u1_slv_re_reg/P0001 ,
		\u4_u1_slv_we_reg/P0001 ,
		\wb1_cyc_i_pad ,
		_w2179_
	);
	LUT2 #(
		.INIT('h8)
	) name1445 (
		_w2178_,
		_w2179_,
		_w2180_
	);
	LUT3 #(
		.INIT('h80)
	) name1446 (
		_w839_,
		_w840_,
		_w841_,
		_w2181_
	);
	LUT4 #(
		.INIT('h2aaa)
	) name1447 (
		\u0_u0_ch_csr_r_reg[5]/NET0131 ,
		_w1051_,
		_w1053_,
		_w1054_,
		_w2182_
	);
	LUT3 #(
		.INIT('h40)
	) name1448 (
		\u3_u1_slv_adr_reg[4]/NET0131 ,
		\u3_u1_slv_dout_reg[5]/P0001 ,
		\u3_u1_slv_we_reg/P0001 ,
		_w2183_
	);
	LUT3 #(
		.INIT('h80)
	) name1449 (
		_w1051_,
		_w1053_,
		_w2183_,
		_w2184_
	);
	LUT2 #(
		.INIT('he)
	) name1450 (
		_w2182_,
		_w2184_,
		_w2185_
	);
	LUT4 #(
		.INIT('h2aaa)
	) name1451 (
		\u0_u0_ch_csr_r_reg[6]/NET0131 ,
		_w1051_,
		_w1053_,
		_w1054_,
		_w2186_
	);
	LUT3 #(
		.INIT('h40)
	) name1452 (
		\u3_u1_slv_adr_reg[4]/NET0131 ,
		\u3_u1_slv_dout_reg[6]/P0001 ,
		\u3_u1_slv_we_reg/P0001 ,
		_w2187_
	);
	LUT3 #(
		.INIT('h80)
	) name1453 (
		_w1051_,
		_w1053_,
		_w2187_,
		_w2188_
	);
	LUT2 #(
		.INIT('he)
	) name1454 (
		_w2186_,
		_w2188_,
		_w2189_
	);
	LUT4 #(
		.INIT('h2aaa)
	) name1455 (
		\u0_u0_ch_csr_r_reg[7]/NET0131 ,
		_w1051_,
		_w1053_,
		_w1054_,
		_w2190_
	);
	LUT3 #(
		.INIT('h40)
	) name1456 (
		\u3_u1_slv_adr_reg[4]/NET0131 ,
		\u3_u1_slv_dout_reg[7]/P0001 ,
		\u3_u1_slv_we_reg/P0001 ,
		_w2191_
	);
	LUT3 #(
		.INIT('h80)
	) name1457 (
		_w1051_,
		_w1053_,
		_w2191_,
		_w2192_
	);
	LUT2 #(
		.INIT('he)
	) name1458 (
		_w2190_,
		_w2192_,
		_w2193_
	);
	LUT4 #(
		.INIT('h2aaa)
	) name1459 (
		\u0_u0_ch_csr_r_reg[8]/NET0131 ,
		_w1051_,
		_w1053_,
		_w1054_,
		_w2194_
	);
	LUT3 #(
		.INIT('h40)
	) name1460 (
		\u3_u1_slv_adr_reg[4]/NET0131 ,
		\u3_u1_slv_dout_reg[8]/P0001 ,
		\u3_u1_slv_we_reg/P0001 ,
		_w2195_
	);
	LUT3 #(
		.INIT('h80)
	) name1461 (
		_w1051_,
		_w1053_,
		_w2195_,
		_w2196_
	);
	LUT2 #(
		.INIT('he)
	) name1462 (
		_w2194_,
		_w2196_,
		_w2197_
	);
	LUT3 #(
		.INIT('h40)
	) name1463 (
		\u3_u1_slv_adr_reg[4]/NET0131 ,
		\u3_u1_slv_dout_reg[9]/P0001 ,
		\u3_u1_slv_we_reg/P0001 ,
		_w2198_
	);
	LUT3 #(
		.INIT('h80)
	) name1464 (
		_w1051_,
		_w1053_,
		_w2198_,
		_w2199_
	);
	LUT4 #(
		.INIT('h7f80)
	) name1465 (
		\u2_adr1_cnt_reg[0]/P0001 ,
		\u2_adr1_cnt_reg[1]/P0001 ,
		\u2_adr1_cnt_reg[2]/P0001 ,
		\u2_adr1_cnt_reg[3]/P0001 ,
		_w2200_
	);
	LUT3 #(
		.INIT('h10)
	) name1466 (
		\u3_u1_slv_adr_reg[4]/NET0131 ,
		\u3_u1_slv_adr_reg[5]/P0001 ,
		\u3_u1_slv_we_reg/P0001 ,
		_w2201_
	);
	LUT3 #(
		.INIT('h80)
	) name1467 (
		_w1051_,
		_w1253_,
		_w2201_,
		_w2202_
	);
	LUT4 #(
		.INIT('h2aaa)
	) name1468 (
		\u0_int_maska_r_reg[0]/NET0131 ,
		_w1051_,
		_w1253_,
		_w2201_,
		_w2203_
	);
	LUT3 #(
		.INIT('h80)
	) name1469 (
		_w1051_,
		_w1262_,
		_w2201_,
		_w2204_
	);
	LUT2 #(
		.INIT('he)
	) name1470 (
		_w2203_,
		_w2204_,
		_w2205_
	);
	LUT4 #(
		.INIT('h2aaa)
	) name1471 (
		\u0_int_maska_r_reg[10]/NET0131 ,
		_w1051_,
		_w1253_,
		_w2201_,
		_w2206_
	);
	LUT3 #(
		.INIT('h80)
	) name1472 (
		_w1051_,
		_w1274_,
		_w2201_,
		_w2207_
	);
	LUT2 #(
		.INIT('he)
	) name1473 (
		_w2206_,
		_w2207_,
		_w2208_
	);
	LUT4 #(
		.INIT('h2aaa)
	) name1474 (
		\u0_int_maska_r_reg[11]/NET0131 ,
		_w1051_,
		_w1253_,
		_w2201_,
		_w2209_
	);
	LUT3 #(
		.INIT('h80)
	) name1475 (
		_w1051_,
		_w1281_,
		_w2201_,
		_w2210_
	);
	LUT2 #(
		.INIT('he)
	) name1476 (
		_w2209_,
		_w2210_,
		_w2211_
	);
	LUT4 #(
		.INIT('h2aaa)
	) name1477 (
		\u0_int_maska_r_reg[8]/NET0131 ,
		_w1051_,
		_w1253_,
		_w2201_,
		_w2212_
	);
	LUT3 #(
		.INIT('h80)
	) name1478 (
		_w1051_,
		_w1330_,
		_w2201_,
		_w2213_
	);
	LUT2 #(
		.INIT('he)
	) name1479 (
		_w2212_,
		_w2213_,
		_w2214_
	);
	LUT4 #(
		.INIT('h2aaa)
	) name1480 (
		\u0_int_maska_r_reg[5]/NET0131 ,
		_w1051_,
		_w1253_,
		_w2201_,
		_w2215_
	);
	LUT3 #(
		.INIT('h80)
	) name1481 (
		_w1051_,
		_w1309_,
		_w2201_,
		_w2216_
	);
	LUT2 #(
		.INIT('he)
	) name1482 (
		_w2215_,
		_w2216_,
		_w2217_
	);
	LUT4 #(
		.INIT('h2aaa)
	) name1483 (
		\u0_int_maska_r_reg[6]/NET0131 ,
		_w1051_,
		_w1253_,
		_w2201_,
		_w2218_
	);
	LUT3 #(
		.INIT('h80)
	) name1484 (
		_w1051_,
		_w1316_,
		_w2201_,
		_w2219_
	);
	LUT2 #(
		.INIT('he)
	) name1485 (
		_w2218_,
		_w2219_,
		_w2220_
	);
	LUT4 #(
		.INIT('h2aaa)
	) name1486 (
		\u0_int_maska_r_reg[7]/NET0131 ,
		_w1051_,
		_w1253_,
		_w2201_,
		_w2221_
	);
	LUT3 #(
		.INIT('h80)
	) name1487 (
		_w1051_,
		_w1323_,
		_w2201_,
		_w2222_
	);
	LUT2 #(
		.INIT('he)
	) name1488 (
		_w2221_,
		_w2222_,
		_w2223_
	);
	LUT4 #(
		.INIT('h2aaa)
	) name1489 (
		\u0_int_maska_r_reg[9]/NET0131 ,
		_w1051_,
		_w1253_,
		_w2201_,
		_w2224_
	);
	LUT3 #(
		.INIT('h80)
	) name1490 (
		_w1051_,
		_w1337_,
		_w2201_,
		_w2225_
	);
	LUT2 #(
		.INIT('he)
	) name1491 (
		_w2224_,
		_w2225_,
		_w2226_
	);
	LUT3 #(
		.INIT('h10)
	) name1492 (
		\u3_u1_slv_adr_reg[2]/NET0131 ,
		\u3_u1_slv_adr_reg[3]/P0001 ,
		\u3_u1_slv_dout_reg[0]/P0001 ,
		_w2227_
	);
	LUT3 #(
		.INIT('h80)
	) name1493 (
		_w1051_,
		_w2201_,
		_w2227_,
		_w2228_
	);
	LUT4 #(
		.INIT('h2aaa)
	) name1494 (
		\u0_csr_r_reg[0]/NET0131 ,
		_w1051_,
		_w1052_,
		_w2201_,
		_w2229_
	);
	LUT2 #(
		.INIT('he)
	) name1495 (
		_w2228_,
		_w2229_,
		_w2230_
	);
	LUT4 #(
		.INIT('h7f80)
	) name1496 (
		\u2_adr0_cnt_reg[0]/P0001 ,
		\u2_adr0_cnt_reg[1]/P0001 ,
		\u2_adr0_cnt_reg[2]/P0001 ,
		\u2_adr0_cnt_reg[3]/P0001 ,
		_w2231_
	);
	LUT4 #(
		.INIT('h6aaa)
	) name1497 (
		\u2_adr1_cnt_reg[10]/P0001 ,
		_w1381_,
		_w1382_,
		_w1383_,
		_w2232_
	);
	LUT4 #(
		.INIT('h6aaa)
	) name1498 (
		\u2_adr0_cnt_reg[10]/P0001 ,
		_w1372_,
		_w1373_,
		_w1374_,
		_w2233_
	);
	LUT4 #(
		.INIT('h78f0)
	) name1499 (
		\u2_adr0_cnt_reg[4]/P0001 ,
		\u2_adr0_cnt_reg[5]/P0001 ,
		\u2_adr0_cnt_reg[6]/P0001 ,
		_w1372_,
		_w2234_
	);
	LUT3 #(
		.INIT('h0e)
	) name1500 (
		\u2_adr0_cnt_reg[13]/P0001 ,
		_w1379_,
		_w2171_,
		_w2235_
	);
	LUT3 #(
		.INIT('h0e)
	) name1501 (
		\u2_adr1_cnt_reg[13]/P0001 ,
		_w1388_,
		_w2174_,
		_w2236_
	);
	LUT4 #(
		.INIT('h78f0)
	) name1502 (
		\u2_adr1_cnt_reg[4]/P0001 ,
		\u2_adr1_cnt_reg[5]/P0001 ,
		\u2_adr1_cnt_reg[6]/P0001 ,
		_w1381_,
		_w2237_
	);
	LUT3 #(
		.INIT('h80)
	) name1503 (
		_w1051_,
		_w1514_,
		_w2201_,
		_w2238_
	);
	LUT4 #(
		.INIT('h2aaa)
	) name1504 (
		\u0_int_maskb_r_reg[11]/NET0131 ,
		_w1051_,
		_w1514_,
		_w2201_,
		_w2239_
	);
	LUT3 #(
		.INIT('h80)
	) name1505 (
		_w1051_,
		_w1951_,
		_w2201_,
		_w2240_
	);
	LUT2 #(
		.INIT('he)
	) name1506 (
		_w2239_,
		_w2240_,
		_w2241_
	);
	LUT4 #(
		.INIT('h2aaa)
	) name1507 (
		\u0_int_maskb_r_reg[10]/NET0131 ,
		_w1051_,
		_w1514_,
		_w2201_,
		_w2242_
	);
	LUT3 #(
		.INIT('h80)
	) name1508 (
		_w1051_,
		_w2014_,
		_w2201_,
		_w2243_
	);
	LUT2 #(
		.INIT('he)
	) name1509 (
		_w2242_,
		_w2243_,
		_w2244_
	);
	LUT4 #(
		.INIT('h2aaa)
	) name1510 (
		\u0_int_maskb_r_reg[0]/NET0131 ,
		_w1051_,
		_w1514_,
		_w2201_,
		_w2245_
	);
	LUT3 #(
		.INIT('h40)
	) name1511 (
		\u3_u1_slv_adr_reg[2]/NET0131 ,
		\u3_u1_slv_adr_reg[3]/P0001 ,
		\u3_u1_slv_dout_reg[0]/P0001 ,
		_w2246_
	);
	LUT3 #(
		.INIT('h80)
	) name1512 (
		_w1051_,
		_w2201_,
		_w2246_,
		_w2247_
	);
	LUT2 #(
		.INIT('he)
	) name1513 (
		_w2245_,
		_w2247_,
		_w2248_
	);
	LUT4 #(
		.INIT('h2aaa)
	) name1514 (
		\u0_int_maskb_r_reg[5]/NET0131 ,
		_w1051_,
		_w1514_,
		_w2201_,
		_w2249_
	);
	LUT3 #(
		.INIT('h80)
	) name1515 (
		_w1051_,
		_w1979_,
		_w2201_,
		_w2250_
	);
	LUT2 #(
		.INIT('he)
	) name1516 (
		_w2249_,
		_w2250_,
		_w2251_
	);
	LUT4 #(
		.INIT('h2aaa)
	) name1517 (
		\u0_int_maskb_r_reg[6]/NET0131 ,
		_w1051_,
		_w1514_,
		_w2201_,
		_w2252_
	);
	LUT3 #(
		.INIT('h80)
	) name1518 (
		_w1051_,
		_w1986_,
		_w2201_,
		_w2253_
	);
	LUT2 #(
		.INIT('he)
	) name1519 (
		_w2252_,
		_w2253_,
		_w2254_
	);
	LUT4 #(
		.INIT('h2aaa)
	) name1520 (
		\u0_int_maskb_r_reg[7]/NET0131 ,
		_w1051_,
		_w1514_,
		_w2201_,
		_w2255_
	);
	LUT3 #(
		.INIT('h80)
	) name1521 (
		_w1051_,
		_w1993_,
		_w2201_,
		_w2256_
	);
	LUT2 #(
		.INIT('he)
	) name1522 (
		_w2255_,
		_w2256_,
		_w2257_
	);
	LUT4 #(
		.INIT('h2aaa)
	) name1523 (
		\u0_int_maskb_r_reg[8]/NET0131 ,
		_w1051_,
		_w1514_,
		_w2201_,
		_w2258_
	);
	LUT3 #(
		.INIT('h80)
	) name1524 (
		_w1051_,
		_w2000_,
		_w2201_,
		_w2259_
	);
	LUT2 #(
		.INIT('he)
	) name1525 (
		_w2258_,
		_w2259_,
		_w2260_
	);
	LUT4 #(
		.INIT('h2aaa)
	) name1526 (
		\u0_int_maskb_r_reg[9]/NET0131 ,
		_w1051_,
		_w1514_,
		_w2201_,
		_w2261_
	);
	LUT3 #(
		.INIT('h80)
	) name1527 (
		_w1051_,
		_w2007_,
		_w2201_,
		_w2262_
	);
	LUT2 #(
		.INIT('he)
	) name1528 (
		_w2261_,
		_w2262_,
		_w2263_
	);
	LUT4 #(
		.INIT('h1555)
	) name1529 (
		\u2_adr0_cnt_reg[9]/P0001 ,
		_w1372_,
		_w1373_,
		_w1510_,
		_w2264_
	);
	LUT2 #(
		.INIT('h1)
	) name1530 (
		_w1375_,
		_w2264_,
		_w2265_
	);
	LUT4 #(
		.INIT('h1555)
	) name1531 (
		\u2_adr1_cnt_reg[9]/P0001 ,
		_w1381_,
		_w1382_,
		_w1512_,
		_w2266_
	);
	LUT2 #(
		.INIT('h1)
	) name1532 (
		_w1384_,
		_w2266_,
		_w2267_
	);
	LUT4 #(
		.INIT('h0001)
	) name1533 (
		\wb1_addr_i[28]_pad ,
		\wb1_addr_i[29]_pad ,
		\wb1_addr_i[30]_pad ,
		\wb1_addr_i[31]_pad ,
		_w2268_
	);
	LUT4 #(
		.INIT('h0010)
	) name1534 (
		\u4_u1_rf_ack_reg/P0001 ,
		\u4_u1_slv_re_reg/P0001 ,
		\wb1_stb_i_pad ,
		\wb1_we_i_pad ,
		_w2269_
	);
	LUT3 #(
		.INIT('h80)
	) name1535 (
		\wb1_cyc_i_pad ,
		_w2268_,
		_w2269_,
		_w2270_
	);
	LUT4 #(
		.INIT('h0001)
	) name1536 (
		\wb0_addr_i[28]_pad ,
		\wb0_addr_i[29]_pad ,
		\wb0_addr_i[30]_pad ,
		\wb0_addr_i[31]_pad ,
		_w2271_
	);
	LUT3 #(
		.INIT('h40)
	) name1537 (
		\u3_u1_rf_ack_reg/P0001 ,
		\wb0_cyc_i_pad ,
		\wb0_stb_i_pad ,
		_w2272_
	);
	LUT2 #(
		.INIT('h1)
	) name1538 (
		\u3_u1_slv_re_reg/P0001 ,
		\wb0_we_i_pad ,
		_w2273_
	);
	LUT3 #(
		.INIT('h80)
	) name1539 (
		_w2271_,
		_w2272_,
		_w2273_,
		_w2274_
	);
	LUT4 #(
		.INIT('h4000)
	) name1540 (
		\u4_u1_rf_ack_reg/P0001 ,
		\wb1_cyc_i_pad ,
		\wb1_stb_i_pad ,
		\wb1_we_i_pad ,
		_w2275_
	);
	LUT2 #(
		.INIT('h8)
	) name1541 (
		_w2268_,
		_w2275_,
		_w2276_
	);
	LUT3 #(
		.INIT('h6c)
	) name1542 (
		\u2_adr0_cnt_reg[4]/P0001 ,
		\u2_adr0_cnt_reg[5]/P0001 ,
		_w1372_,
		_w2277_
	);
	LUT3 #(
		.INIT('h6c)
	) name1543 (
		\u2_adr1_cnt_reg[4]/P0001 ,
		\u2_adr1_cnt_reg[5]/P0001 ,
		_w1381_,
		_w2278_
	);
	LUT4 #(
		.INIT('h4000)
	) name1544 (
		\u3_u1_rf_ack_reg/P0001 ,
		\wb0_cyc_i_pad ,
		\wb0_stb_i_pad ,
		\wb0_we_i_pad ,
		_w2279_
	);
	LUT2 #(
		.INIT('h8)
	) name1545 (
		_w2271_,
		_w2279_,
		_w2280_
	);
	LUT3 #(
		.INIT('h78)
	) name1546 (
		\u2_adr0_cnt_reg[0]/P0001 ,
		\u2_adr0_cnt_reg[1]/P0001 ,
		\u2_adr0_cnt_reg[2]/P0001 ,
		_w2281_
	);
	LUT3 #(
		.INIT('h78)
	) name1547 (
		\u2_adr1_cnt_reg[0]/P0001 ,
		\u2_adr1_cnt_reg[1]/P0001 ,
		\u2_adr1_cnt_reg[2]/P0001 ,
		_w2282_
	);
	LUT4 #(
		.INIT('h4c0c)
	) name1548 (
		dma_ack_o_pad,
		\u0_u0_ch_csr_r_reg[0]/NET0131 ,
		\u0_u0_ch_csr_r_reg[5]/NET0131 ,
		\u1_req_r_reg[0]/P0001 ,
		_w2283_
	);
	LUT2 #(
		.INIT('h1)
	) name1549 (
		\u3_u1_slv_re_reg/P0001 ,
		\u3_u1_slv_we_reg/P0001 ,
		_w2284_
	);
	LUT2 #(
		.INIT('h2)
	) name1550 (
		_w2272_,
		_w2284_,
		_w2285_
	);
	LUT2 #(
		.INIT('h6)
	) name1551 (
		\u2_adr0_cnt_reg[0]/P0001 ,
		\u2_adr0_cnt_reg[1]/P0001 ,
		_w2286_
	);
	LUT2 #(
		.INIT('h6)
	) name1552 (
		\u2_adr1_cnt_reg[0]/P0001 ,
		\u2_adr1_cnt_reg[1]/P0001 ,
		_w2287_
	);
	LUT2 #(
		.INIT('h2)
	) name1553 (
		dma_nd_i_pad,
		dma_req_i_pad,
		_w2288_
	);
	LUT2 #(
		.INIT('h4)
	) name1554 (
		dma_ack_o_pad,
		dma_req_i_pad,
		_w2289_
	);
	LUT2 #(
		.INIT('h8)
	) name1555 (
		dma_nd_i_pad,
		dma_req_i_pad,
		_w2290_
	);
	LUT2 #(
		.INIT('h9)
	) name1556 (
		\u2_tsz_cnt_reg[2]/NET0131 ,
		_w1209_,
		_w2291_
	);
	LUT3 #(
		.INIT('h2e)
	) name1557 (
		\u0_u0_ch_tot_sz_r_reg[2]/P0001 ,
		_w750_,
		_w2291_,
		_w2292_
	);
	LUT4 #(
		.INIT('h20aa)
	) name1558 (
		\u0_u0_ch_adr1_r_reg[25]/P0001 ,
		_w747_,
		_w748_,
		_w749_,
		_w2293_
	);
	LUT3 #(
		.INIT('h15)
	) name1559 (
		\u2_adr1_cnt_reg[25]/P0001 ,
		_w742_,
		_w794_,
		_w2294_
	);
	LUT3 #(
		.INIT('h4c)
	) name1560 (
		_w742_,
		_w750_,
		_w778_,
		_w2295_
	);
	LUT3 #(
		.INIT('hba)
	) name1561 (
		_w2293_,
		_w2294_,
		_w2295_,
		_w2296_
	);
	LUT4 #(
		.INIT('h5355)
	) name1562 (
		\u2_adr0_cnt_reg[13]/P0001 ,
		\u2_u0_out_r_reg[13]/P0001 ,
		_w757_,
		_w758_,
		_w2297_
	);
	LUT3 #(
		.INIT('h2e)
	) name1563 (
		\u0_u0_ch_adr0_r_reg[13]/P0001 ,
		_w750_,
		_w2297_,
		_w2298_
	);
	LUT2 #(
		.INIT('h8)
	) name1564 (
		\u0_u0_ch_tot_sz_r_reg[10]/P0001 ,
		_w1408_,
		_w2299_
	);
	LUT4 #(
		.INIT('h135f)
	) name1565 (
		\u0_int_maskb_r_reg[10]/NET0131 ,
		\u0_u0_ch_busy_reg/P0001 ,
		_w1413_,
		_w1418_,
		_w2300_
	);
	LUT3 #(
		.INIT('h13)
	) name1566 (
		\u0_int_maska_r_reg[10]/NET0131 ,
		_w1402_,
		_w1411_,
		_w2301_
	);
	LUT3 #(
		.INIT('h80)
	) name1567 (
		\u0_u0_ch_adr0_r_reg[8]/P0001 ,
		_w1051_,
		_w1397_,
		_w2302_
	);
	LUT4 #(
		.INIT('h0400)
	) name1568 (
		_w1391_,
		_w1393_,
		_w1396_,
		_w2302_,
		_w2303_
	);
	LUT3 #(
		.INIT('h80)
	) name1569 (
		\u0_u0_ch_adr1_r_reg[8]/P0001 ,
		_w1051_,
		_w1397_,
		_w2304_
	);
	LUT4 #(
		.INIT('h4000)
	) name1570 (
		_w1391_,
		_w1393_,
		_w1396_,
		_w2304_,
		_w2305_
	);
	LUT2 #(
		.INIT('h1)
	) name1571 (
		_w2303_,
		_w2305_,
		_w2306_
	);
	LUT4 #(
		.INIT('hbfff)
	) name1572 (
		_w2299_,
		_w2300_,
		_w2301_,
		_w2306_,
		_w2307_
	);
	LUT4 #(
		.INIT('h2aaa)
	) name1573 (
		\u0_u0_ch_done_reg/P0002 ,
		_w1051_,
		_w1053_,
		_w1054_,
		_w2308_
	);
	LUT4 #(
		.INIT('h00ef)
	) name1574 (
		_w1059_,
		_w1062_,
		_w1064_,
		_w2308_,
		_w2309_
	);
	LUT2 #(
		.INIT('hb)
	) name1575 (
		_w1056_,
		_w2309_,
		_w2310_
	);
	LUT4 #(
		.INIT('hf800)
	) name1576 (
		_w862_,
		_w867_,
		_w870_,
		_w898_,
		_w2311_
	);
	LUT3 #(
		.INIT('h0b)
	) name1577 (
		_w860_,
		_w872_,
		_w2311_,
		_w2312_
	);
	LUT4 #(
		.INIT('haae2)
	) name1578 (
		\u3_u1_rf_ack_reg/P0001 ,
		\wb0_cyc_i_pad ,
		\wb1_ack_i_pad ,
		_w2271_,
		_w2313_
	);
	LUT2 #(
		.INIT('h8)
	) name1579 (
		\wb1_addr_i[0]_pad ,
		\wb1_cyc_i_pad ,
		_w2314_
	);
	LUT2 #(
		.INIT('h4)
	) name1580 (
		_w2268_,
		_w2314_,
		_w2315_
	);
	LUT2 #(
		.INIT('h2)
	) name1581 (
		\wb1_cyc_i_pad ,
		_w2268_,
		_w2316_
	);
	LUT4 #(
		.INIT('haaca)
	) name1582 (
		\u2_mast0_adr_reg[10]/P0001 ,
		\wb1_addr_i[10]_pad ,
		\wb1_cyc_i_pad ,
		_w2268_,
		_w2317_
	);
	LUT4 #(
		.INIT('haaca)
	) name1583 (
		\u2_mast0_adr_reg[11]/P0001 ,
		\wb1_addr_i[11]_pad ,
		\wb1_cyc_i_pad ,
		_w2268_,
		_w2318_
	);
	LUT4 #(
		.INIT('haaca)
	) name1584 (
		\u2_mast0_adr_reg[12]/P0001 ,
		\wb1_addr_i[12]_pad ,
		\wb1_cyc_i_pad ,
		_w2268_,
		_w2319_
	);
	LUT4 #(
		.INIT('haaca)
	) name1585 (
		\u2_mast0_adr_reg[13]/P0001 ,
		\wb1_addr_i[13]_pad ,
		\wb1_cyc_i_pad ,
		_w2268_,
		_w2320_
	);
	LUT4 #(
		.INIT('haaca)
	) name1586 (
		\u2_mast0_adr_reg[14]/P0001 ,
		\wb1_addr_i[14]_pad ,
		\wb1_cyc_i_pad ,
		_w2268_,
		_w2321_
	);
	LUT4 #(
		.INIT('haaca)
	) name1587 (
		\u2_mast0_adr_reg[15]/P0001 ,
		\wb1_addr_i[15]_pad ,
		\wb1_cyc_i_pad ,
		_w2268_,
		_w2322_
	);
	LUT4 #(
		.INIT('haaca)
	) name1588 (
		\u2_mast0_adr_reg[16]/P0001 ,
		\wb1_addr_i[16]_pad ,
		\wb1_cyc_i_pad ,
		_w2268_,
		_w2323_
	);
	LUT4 #(
		.INIT('haaca)
	) name1589 (
		\u2_mast0_adr_reg[17]/P0001 ,
		\wb1_addr_i[17]_pad ,
		\wb1_cyc_i_pad ,
		_w2268_,
		_w2324_
	);
	LUT4 #(
		.INIT('haaca)
	) name1590 (
		\u2_mast0_adr_reg[18]/P0001 ,
		\wb1_addr_i[18]_pad ,
		\wb1_cyc_i_pad ,
		_w2268_,
		_w2325_
	);
	LUT4 #(
		.INIT('haaca)
	) name1591 (
		\u2_mast0_adr_reg[19]/P0001 ,
		\wb1_addr_i[19]_pad ,
		\wb1_cyc_i_pad ,
		_w2268_,
		_w2326_
	);
	LUT2 #(
		.INIT('h8)
	) name1592 (
		\wb1_addr_i[1]_pad ,
		\wb1_cyc_i_pad ,
		_w2327_
	);
	LUT2 #(
		.INIT('h4)
	) name1593 (
		_w2268_,
		_w2327_,
		_w2328_
	);
	LUT4 #(
		.INIT('haaca)
	) name1594 (
		\u2_mast0_adr_reg[20]/P0001 ,
		\wb1_addr_i[20]_pad ,
		\wb1_cyc_i_pad ,
		_w2268_,
		_w2329_
	);
	LUT4 #(
		.INIT('haaca)
	) name1595 (
		\u2_mast0_adr_reg[21]/P0001 ,
		\wb1_addr_i[21]_pad ,
		\wb1_cyc_i_pad ,
		_w2268_,
		_w2330_
	);
	LUT4 #(
		.INIT('haaca)
	) name1596 (
		\u2_mast0_adr_reg[22]/P0001 ,
		\wb1_addr_i[22]_pad ,
		\wb1_cyc_i_pad ,
		_w2268_,
		_w2331_
	);
	LUT4 #(
		.INIT('haaca)
	) name1597 (
		\u2_mast0_adr_reg[23]/P0001 ,
		\wb1_addr_i[23]_pad ,
		\wb1_cyc_i_pad ,
		_w2268_,
		_w2332_
	);
	LUT4 #(
		.INIT('haaca)
	) name1598 (
		\u2_mast0_adr_reg[24]/P0001 ,
		\wb1_addr_i[24]_pad ,
		\wb1_cyc_i_pad ,
		_w2268_,
		_w2333_
	);
	LUT4 #(
		.INIT('haaca)
	) name1599 (
		\u2_mast0_adr_reg[25]/P0001 ,
		\wb1_addr_i[25]_pad ,
		\wb1_cyc_i_pad ,
		_w2268_,
		_w2334_
	);
	LUT4 #(
		.INIT('haaca)
	) name1600 (
		\u2_mast0_adr_reg[26]/P0001 ,
		\wb1_addr_i[26]_pad ,
		\wb1_cyc_i_pad ,
		_w2268_,
		_w2335_
	);
	LUT4 #(
		.INIT('haaca)
	) name1601 (
		\u2_mast0_adr_reg[27]/P0001 ,
		\wb1_addr_i[27]_pad ,
		\wb1_cyc_i_pad ,
		_w2268_,
		_w2336_
	);
	LUT3 #(
		.INIT('h15)
	) name1602 (
		\u2_mast0_adr_reg[28]/P0001 ,
		\wb1_addr_i[28]_pad ,
		\wb1_cyc_i_pad ,
		_w2337_
	);
	LUT2 #(
		.INIT('h4)
	) name1603 (
		\wb1_addr_i[28]_pad ,
		\wb1_cyc_i_pad ,
		_w2338_
	);
	LUT3 #(
		.INIT('h23)
	) name1604 (
		_w2268_,
		_w2337_,
		_w2338_,
		_w2339_
	);
	LUT3 #(
		.INIT('h15)
	) name1605 (
		\u2_mast0_adr_reg[29]/P0001 ,
		\wb1_addr_i[29]_pad ,
		\wb1_cyc_i_pad ,
		_w2340_
	);
	LUT2 #(
		.INIT('h4)
	) name1606 (
		\wb1_addr_i[29]_pad ,
		\wb1_cyc_i_pad ,
		_w2341_
	);
	LUT3 #(
		.INIT('h23)
	) name1607 (
		_w2268_,
		_w2340_,
		_w2341_,
		_w2342_
	);
	LUT4 #(
		.INIT('haaca)
	) name1608 (
		\u2_mast0_adr_reg[2]/P0001 ,
		\wb1_addr_i[2]_pad ,
		\wb1_cyc_i_pad ,
		_w2268_,
		_w2343_
	);
	LUT3 #(
		.INIT('h15)
	) name1609 (
		\u2_mast0_adr_reg[30]/P0001 ,
		\wb1_addr_i[30]_pad ,
		\wb1_cyc_i_pad ,
		_w2344_
	);
	LUT2 #(
		.INIT('h4)
	) name1610 (
		\wb1_addr_i[30]_pad ,
		\wb1_cyc_i_pad ,
		_w2345_
	);
	LUT3 #(
		.INIT('h23)
	) name1611 (
		_w2268_,
		_w2344_,
		_w2345_,
		_w2346_
	);
	LUT3 #(
		.INIT('h15)
	) name1612 (
		\u2_mast0_adr_reg[31]/P0001 ,
		\wb1_addr_i[31]_pad ,
		\wb1_cyc_i_pad ,
		_w2347_
	);
	LUT2 #(
		.INIT('h4)
	) name1613 (
		\wb1_addr_i[31]_pad ,
		\wb1_cyc_i_pad ,
		_w2348_
	);
	LUT3 #(
		.INIT('h23)
	) name1614 (
		_w2268_,
		_w2347_,
		_w2348_,
		_w2349_
	);
	LUT4 #(
		.INIT('haaca)
	) name1615 (
		\u2_mast0_adr_reg[3]/NET0131 ,
		\wb1_addr_i[3]_pad ,
		\wb1_cyc_i_pad ,
		_w2268_,
		_w2350_
	);
	LUT4 #(
		.INIT('haaca)
	) name1616 (
		\u2_mast0_adr_reg[4]/P0001 ,
		\wb1_addr_i[4]_pad ,
		\wb1_cyc_i_pad ,
		_w2268_,
		_w2351_
	);
	LUT4 #(
		.INIT('haaca)
	) name1617 (
		\u2_mast0_adr_reg[5]/P0001 ,
		\wb1_addr_i[5]_pad ,
		\wb1_cyc_i_pad ,
		_w2268_,
		_w2352_
	);
	LUT4 #(
		.INIT('haaca)
	) name1618 (
		\u2_mast0_adr_reg[6]/P0001 ,
		\wb1_addr_i[6]_pad ,
		\wb1_cyc_i_pad ,
		_w2268_,
		_w2353_
	);
	LUT4 #(
		.INIT('haaca)
	) name1619 (
		\u2_mast0_adr_reg[7]/P0001 ,
		\wb1_addr_i[7]_pad ,
		\wb1_cyc_i_pad ,
		_w2268_,
		_w2354_
	);
	LUT4 #(
		.INIT('haaca)
	) name1620 (
		\u2_mast0_adr_reg[8]/P0001 ,
		\wb1_addr_i[8]_pad ,
		\wb1_cyc_i_pad ,
		_w2268_,
		_w2355_
	);
	LUT4 #(
		.INIT('haaca)
	) name1621 (
		\u2_mast0_adr_reg[9]/P0001 ,
		\wb1_addr_i[9]_pad ,
		\wb1_cyc_i_pad ,
		_w2268_,
		_w2356_
	);
	LUT3 #(
		.INIT('hae)
	) name1622 (
		\u3_u0_mast_cyc_reg/P0001 ,
		\wb1_cyc_i_pad ,
		_w2268_,
		_w2357_
	);
	LUT2 #(
		.INIT('h8)
	) name1623 (
		\wb0_cyc_i_pad ,
		\wb1_err_i_pad ,
		_w2358_
	);
	LUT2 #(
		.INIT('h4)
	) name1624 (
		_w2271_,
		_w2358_,
		_w2359_
	);
	LUT2 #(
		.INIT('h8)
	) name1625 (
		\wb0_cyc_i_pad ,
		\wb1_rty_i_pad ,
		_w2360_
	);
	LUT2 #(
		.INIT('h4)
	) name1626 (
		_w2271_,
		_w2360_,
		_w2361_
	);
	LUT2 #(
		.INIT('h2)
	) name1627 (
		\wb1_cyc_i_pad ,
		\wb1_sel_i[0]_pad ,
		_w2362_
	);
	LUT2 #(
		.INIT('hb)
	) name1628 (
		_w2268_,
		_w2362_,
		_w2363_
	);
	LUT2 #(
		.INIT('h2)
	) name1629 (
		\wb1_cyc_i_pad ,
		\wb1_sel_i[1]_pad ,
		_w2364_
	);
	LUT2 #(
		.INIT('hb)
	) name1630 (
		_w2268_,
		_w2364_,
		_w2365_
	);
	LUT2 #(
		.INIT('h2)
	) name1631 (
		\wb1_cyc_i_pad ,
		\wb1_sel_i[2]_pad ,
		_w2366_
	);
	LUT2 #(
		.INIT('hb)
	) name1632 (
		_w2268_,
		_w2366_,
		_w2367_
	);
	LUT2 #(
		.INIT('h2)
	) name1633 (
		\wb1_cyc_i_pad ,
		\wb1_sel_i[3]_pad ,
		_w2368_
	);
	LUT2 #(
		.INIT('hb)
	) name1634 (
		_w2268_,
		_w2368_,
		_w2369_
	);
	LUT4 #(
		.INIT('haae2)
	) name1635 (
		\u3_u0_mast_stb_reg/P0001 ,
		\wb1_cyc_i_pad ,
		\wb1_stb_i_pad ,
		_w2268_,
		_w2370_
	);
	LUT4 #(
		.INIT('haae2)
	) name1636 (
		\u3_u0_mast_we_r_reg/P0002 ,
		\wb1_cyc_i_pad ,
		\wb1_we_i_pad ,
		_w2268_,
		_w2371_
	);
	LUT4 #(
		.INIT('haae2)
	) name1637 (
		\u0_wb_rf_dout_reg[0]/P0001 ,
		\wb0_cyc_i_pad ,
		\wb1s_data_i[0]_pad ,
		_w2271_,
		_w2372_
	);
	LUT4 #(
		.INIT('haae2)
	) name1638 (
		\u0_wb_rf_dout_reg[10]/P0001 ,
		\wb0_cyc_i_pad ,
		\wb1s_data_i[10]_pad ,
		_w2271_,
		_w2373_
	);
	LUT4 #(
		.INIT('haae2)
	) name1639 (
		\u0_wb_rf_dout_reg[11]/P0001 ,
		\wb0_cyc_i_pad ,
		\wb1s_data_i[11]_pad ,
		_w2271_,
		_w2374_
	);
	LUT4 #(
		.INIT('haae2)
	) name1640 (
		\u0_wb_rf_dout_reg[12]/P0001 ,
		\wb0_cyc_i_pad ,
		\wb1s_data_i[12]_pad ,
		_w2271_,
		_w2375_
	);
	LUT4 #(
		.INIT('haae2)
	) name1641 (
		\u0_wb_rf_dout_reg[13]/P0001 ,
		\wb0_cyc_i_pad ,
		\wb1s_data_i[13]_pad ,
		_w2271_,
		_w2376_
	);
	LUT4 #(
		.INIT('haae2)
	) name1642 (
		\u0_wb_rf_dout_reg[14]/P0001 ,
		\wb0_cyc_i_pad ,
		\wb1s_data_i[14]_pad ,
		_w2271_,
		_w2377_
	);
	LUT4 #(
		.INIT('haae2)
	) name1643 (
		\u0_wb_rf_dout_reg[15]/P0001 ,
		\wb0_cyc_i_pad ,
		\wb1s_data_i[15]_pad ,
		_w2271_,
		_w2378_
	);
	LUT4 #(
		.INIT('haae2)
	) name1644 (
		\u0_wb_rf_dout_reg[16]/P0001 ,
		\wb0_cyc_i_pad ,
		\wb1s_data_i[16]_pad ,
		_w2271_,
		_w2379_
	);
	LUT4 #(
		.INIT('haae2)
	) name1645 (
		\u0_wb_rf_dout_reg[17]/P0001 ,
		\wb0_cyc_i_pad ,
		\wb1s_data_i[17]_pad ,
		_w2271_,
		_w2380_
	);
	LUT4 #(
		.INIT('haae2)
	) name1646 (
		\u0_wb_rf_dout_reg[18]/P0001 ,
		\wb0_cyc_i_pad ,
		\wb1s_data_i[18]_pad ,
		_w2271_,
		_w2381_
	);
	LUT4 #(
		.INIT('haae2)
	) name1647 (
		\u0_wb_rf_dout_reg[19]/P0001 ,
		\wb0_cyc_i_pad ,
		\wb1s_data_i[19]_pad ,
		_w2271_,
		_w2382_
	);
	LUT4 #(
		.INIT('haae2)
	) name1648 (
		\u0_wb_rf_dout_reg[1]/P0001 ,
		\wb0_cyc_i_pad ,
		\wb1s_data_i[1]_pad ,
		_w2271_,
		_w2383_
	);
	LUT4 #(
		.INIT('haae2)
	) name1649 (
		\u0_wb_rf_dout_reg[20]/P0001 ,
		\wb0_cyc_i_pad ,
		\wb1s_data_i[20]_pad ,
		_w2271_,
		_w2384_
	);
	LUT4 #(
		.INIT('haae2)
	) name1650 (
		\u0_wb_rf_dout_reg[21]/P0001 ,
		\wb0_cyc_i_pad ,
		\wb1s_data_i[21]_pad ,
		_w2271_,
		_w2385_
	);
	LUT4 #(
		.INIT('haae2)
	) name1651 (
		\u0_wb_rf_dout_reg[22]/P0001 ,
		\wb0_cyc_i_pad ,
		\wb1s_data_i[22]_pad ,
		_w2271_,
		_w2386_
	);
	LUT4 #(
		.INIT('haae2)
	) name1652 (
		\u0_wb_rf_dout_reg[23]/P0001 ,
		\wb0_cyc_i_pad ,
		\wb1s_data_i[23]_pad ,
		_w2271_,
		_w2387_
	);
	LUT4 #(
		.INIT('haae2)
	) name1653 (
		\u0_wb_rf_dout_reg[24]/P0001 ,
		\wb0_cyc_i_pad ,
		\wb1s_data_i[24]_pad ,
		_w2271_,
		_w2388_
	);
	LUT4 #(
		.INIT('haae2)
	) name1654 (
		\u0_wb_rf_dout_reg[25]/P0001 ,
		\wb0_cyc_i_pad ,
		\wb1s_data_i[25]_pad ,
		_w2271_,
		_w2389_
	);
	LUT4 #(
		.INIT('haae2)
	) name1655 (
		\u0_wb_rf_dout_reg[26]/P0001 ,
		\wb0_cyc_i_pad ,
		\wb1s_data_i[26]_pad ,
		_w2271_,
		_w2390_
	);
	LUT4 #(
		.INIT('haae2)
	) name1656 (
		\u0_wb_rf_dout_reg[27]/P0001 ,
		\wb0_cyc_i_pad ,
		\wb1s_data_i[27]_pad ,
		_w2271_,
		_w2391_
	);
	LUT4 #(
		.INIT('haae2)
	) name1657 (
		\u0_wb_rf_dout_reg[28]/P0001 ,
		\wb0_cyc_i_pad ,
		\wb1s_data_i[28]_pad ,
		_w2271_,
		_w2392_
	);
	LUT4 #(
		.INIT('haae2)
	) name1658 (
		\u0_wb_rf_dout_reg[29]/P0001 ,
		\wb0_cyc_i_pad ,
		\wb1s_data_i[29]_pad ,
		_w2271_,
		_w2393_
	);
	LUT4 #(
		.INIT('haae2)
	) name1659 (
		\u0_wb_rf_dout_reg[2]/P0001 ,
		\wb0_cyc_i_pad ,
		\wb1s_data_i[2]_pad ,
		_w2271_,
		_w2394_
	);
	LUT4 #(
		.INIT('haae2)
	) name1660 (
		\u0_wb_rf_dout_reg[30]/P0001 ,
		\wb0_cyc_i_pad ,
		\wb1s_data_i[30]_pad ,
		_w2271_,
		_w2395_
	);
	LUT4 #(
		.INIT('haae2)
	) name1661 (
		\u0_wb_rf_dout_reg[31]/P0001 ,
		\wb0_cyc_i_pad ,
		\wb1s_data_i[31]_pad ,
		_w2271_,
		_w2396_
	);
	LUT4 #(
		.INIT('haae2)
	) name1662 (
		\u0_wb_rf_dout_reg[3]/P0001 ,
		\wb0_cyc_i_pad ,
		\wb1s_data_i[3]_pad ,
		_w2271_,
		_w2397_
	);
	LUT4 #(
		.INIT('haae2)
	) name1663 (
		\u0_wb_rf_dout_reg[4]/P0001 ,
		\wb0_cyc_i_pad ,
		\wb1s_data_i[4]_pad ,
		_w2271_,
		_w2398_
	);
	LUT4 #(
		.INIT('haae2)
	) name1664 (
		\u0_wb_rf_dout_reg[5]/P0001 ,
		\wb0_cyc_i_pad ,
		\wb1s_data_i[5]_pad ,
		_w2271_,
		_w2399_
	);
	LUT4 #(
		.INIT('haae2)
	) name1665 (
		\u0_wb_rf_dout_reg[6]/P0001 ,
		\wb0_cyc_i_pad ,
		\wb1s_data_i[6]_pad ,
		_w2271_,
		_w2400_
	);
	LUT4 #(
		.INIT('haae2)
	) name1666 (
		\u0_wb_rf_dout_reg[7]/P0001 ,
		\wb0_cyc_i_pad ,
		\wb1s_data_i[7]_pad ,
		_w2271_,
		_w2401_
	);
	LUT4 #(
		.INIT('haae2)
	) name1667 (
		\u0_wb_rf_dout_reg[8]/P0001 ,
		\wb0_cyc_i_pad ,
		\wb1s_data_i[8]_pad ,
		_w2271_,
		_w2402_
	);
	LUT4 #(
		.INIT('haae2)
	) name1668 (
		\u0_wb_rf_dout_reg[9]/P0001 ,
		\wb0_cyc_i_pad ,
		\wb1s_data_i[9]_pad ,
		_w2271_,
		_w2403_
	);
	LUT2 #(
		.INIT('h8)
	) name1669 (
		\wb1_cyc_i_pad ,
		\wb1m_data_i[0]_pad ,
		_w2404_
	);
	LUT2 #(
		.INIT('h4)
	) name1670 (
		_w2268_,
		_w2404_,
		_w2405_
	);
	LUT3 #(
		.INIT('h1b)
	) name1671 (
		\u0_u0_ch_csr_r_reg[2]/NET0131 ,
		\u3_u0_mast_dout_reg[0]/P0001 ,
		\u4_u0_mast_dout_reg[0]/P0001 ,
		_w2406_
	);
	LUT2 #(
		.INIT('h4)
	) name1672 (
		_w869_,
		_w2406_,
		_w2407_
	);
	LUT2 #(
		.INIT('h4)
	) name1673 (
		_w897_,
		_w2407_,
		_w2408_
	);
	LUT2 #(
		.INIT('h4)
	) name1674 (
		\u2_tsz_cnt_reg[0]/NET0131 ,
		_w869_,
		_w2409_
	);
	LUT4 #(
		.INIT('h4000)
	) name1675 (
		\u2_tsz_cnt_reg[0]/NET0131 ,
		_w894_,
		_w895_,
		_w896_,
		_w2410_
	);
	LUT3 #(
		.INIT('h01)
	) name1676 (
		_w2316_,
		_w2409_,
		_w2410_,
		_w2411_
	);
	LUT3 #(
		.INIT('hba)
	) name1677 (
		_w2405_,
		_w2408_,
		_w2411_,
		_w2412_
	);
	LUT2 #(
		.INIT('h8)
	) name1678 (
		\wb1_cyc_i_pad ,
		\wb1m_data_i[10]_pad ,
		_w2413_
	);
	LUT2 #(
		.INIT('h4)
	) name1679 (
		_w2268_,
		_w2413_,
		_w2414_
	);
	LUT3 #(
		.INIT('h1b)
	) name1680 (
		\u0_u0_ch_csr_r_reg[2]/NET0131 ,
		\u3_u0_mast_dout_reg[10]/P0001 ,
		\u4_u0_mast_dout_reg[10]/P0001 ,
		_w2415_
	);
	LUT2 #(
		.INIT('h4)
	) name1681 (
		_w869_,
		_w2415_,
		_w2416_
	);
	LUT2 #(
		.INIT('h4)
	) name1682 (
		_w897_,
		_w2416_,
		_w2417_
	);
	LUT2 #(
		.INIT('h4)
	) name1683 (
		\u2_tsz_cnt_reg[10]/NET0131 ,
		_w869_,
		_w2418_
	);
	LUT4 #(
		.INIT('h4000)
	) name1684 (
		\u2_tsz_cnt_reg[10]/NET0131 ,
		_w894_,
		_w895_,
		_w896_,
		_w2419_
	);
	LUT3 #(
		.INIT('h01)
	) name1685 (
		_w2316_,
		_w2418_,
		_w2419_,
		_w2420_
	);
	LUT3 #(
		.INIT('hba)
	) name1686 (
		_w2414_,
		_w2417_,
		_w2420_,
		_w2421_
	);
	LUT2 #(
		.INIT('h8)
	) name1687 (
		\wb1_cyc_i_pad ,
		\wb1m_data_i[11]_pad ,
		_w2422_
	);
	LUT2 #(
		.INIT('h4)
	) name1688 (
		_w2268_,
		_w2422_,
		_w2423_
	);
	LUT3 #(
		.INIT('h1b)
	) name1689 (
		\u0_u0_ch_csr_r_reg[2]/NET0131 ,
		\u3_u0_mast_dout_reg[11]/P0001 ,
		\u4_u0_mast_dout_reg[11]/P0001 ,
		_w2424_
	);
	LUT2 #(
		.INIT('h4)
	) name1690 (
		_w869_,
		_w2424_,
		_w2425_
	);
	LUT2 #(
		.INIT('h4)
	) name1691 (
		_w897_,
		_w2425_,
		_w2426_
	);
	LUT2 #(
		.INIT('h4)
	) name1692 (
		\u2_tsz_cnt_reg[11]/NET0131 ,
		_w869_,
		_w2427_
	);
	LUT4 #(
		.INIT('h4000)
	) name1693 (
		\u2_tsz_cnt_reg[11]/NET0131 ,
		_w894_,
		_w895_,
		_w896_,
		_w2428_
	);
	LUT3 #(
		.INIT('h01)
	) name1694 (
		_w2316_,
		_w2427_,
		_w2428_,
		_w2429_
	);
	LUT3 #(
		.INIT('hba)
	) name1695 (
		_w2423_,
		_w2426_,
		_w2429_,
		_w2430_
	);
	LUT2 #(
		.INIT('h8)
	) name1696 (
		\wb1_cyc_i_pad ,
		\wb1m_data_i[12]_pad ,
		_w2431_
	);
	LUT2 #(
		.INIT('h4)
	) name1697 (
		_w2268_,
		_w2431_,
		_w2432_
	);
	LUT3 #(
		.INIT('h1b)
	) name1698 (
		\u0_u0_ch_csr_r_reg[2]/NET0131 ,
		\u3_u0_mast_dout_reg[12]/P0001 ,
		\u4_u0_mast_dout_reg[12]/P0001 ,
		_w2433_
	);
	LUT4 #(
		.INIT('h0031)
	) name1699 (
		\wb1_cyc_i_pad ,
		_w869_,
		_w2268_,
		_w2433_,
		_w2434_
	);
	LUT3 #(
		.INIT('hdc)
	) name1700 (
		_w897_,
		_w2432_,
		_w2434_,
		_w2435_
	);
	LUT2 #(
		.INIT('h8)
	) name1701 (
		\wb1_cyc_i_pad ,
		\wb1m_data_i[13]_pad ,
		_w2436_
	);
	LUT2 #(
		.INIT('h4)
	) name1702 (
		_w2268_,
		_w2436_,
		_w2437_
	);
	LUT3 #(
		.INIT('h1b)
	) name1703 (
		\u0_u0_ch_csr_r_reg[2]/NET0131 ,
		\u3_u0_mast_dout_reg[13]/P0001 ,
		\u4_u0_mast_dout_reg[13]/P0001 ,
		_w2438_
	);
	LUT4 #(
		.INIT('h0031)
	) name1704 (
		\wb1_cyc_i_pad ,
		_w869_,
		_w2268_,
		_w2438_,
		_w2439_
	);
	LUT3 #(
		.INIT('hdc)
	) name1705 (
		_w897_,
		_w2437_,
		_w2439_,
		_w2440_
	);
	LUT2 #(
		.INIT('h8)
	) name1706 (
		\wb1_cyc_i_pad ,
		\wb1m_data_i[14]_pad ,
		_w2441_
	);
	LUT2 #(
		.INIT('h4)
	) name1707 (
		_w2268_,
		_w2441_,
		_w2442_
	);
	LUT3 #(
		.INIT('h1b)
	) name1708 (
		\u0_u0_ch_csr_r_reg[2]/NET0131 ,
		\u3_u0_mast_dout_reg[14]/P0001 ,
		\u4_u0_mast_dout_reg[14]/P0001 ,
		_w2443_
	);
	LUT4 #(
		.INIT('h0031)
	) name1709 (
		\wb1_cyc_i_pad ,
		_w869_,
		_w2268_,
		_w2443_,
		_w2444_
	);
	LUT3 #(
		.INIT('hdc)
	) name1710 (
		_w897_,
		_w2442_,
		_w2444_,
		_w2445_
	);
	LUT2 #(
		.INIT('h8)
	) name1711 (
		\wb1_cyc_i_pad ,
		\wb1m_data_i[15]_pad ,
		_w2446_
	);
	LUT2 #(
		.INIT('h4)
	) name1712 (
		_w2268_,
		_w2446_,
		_w2447_
	);
	LUT3 #(
		.INIT('h1b)
	) name1713 (
		\u0_u0_ch_csr_r_reg[2]/NET0131 ,
		\u3_u0_mast_dout_reg[15]/P0001 ,
		\u4_u0_mast_dout_reg[15]/P0001 ,
		_w2448_
	);
	LUT4 #(
		.INIT('h0031)
	) name1714 (
		\wb1_cyc_i_pad ,
		_w869_,
		_w2268_,
		_w2448_,
		_w2449_
	);
	LUT3 #(
		.INIT('hdc)
	) name1715 (
		_w897_,
		_w2447_,
		_w2449_,
		_w2450_
	);
	LUT2 #(
		.INIT('h8)
	) name1716 (
		\wb1_cyc_i_pad ,
		\wb1m_data_i[16]_pad ,
		_w2451_
	);
	LUT2 #(
		.INIT('h4)
	) name1717 (
		_w2268_,
		_w2451_,
		_w2452_
	);
	LUT3 #(
		.INIT('h1b)
	) name1718 (
		\u0_u0_ch_csr_r_reg[2]/NET0131 ,
		\u3_u0_mast_dout_reg[16]/P0001 ,
		\u4_u0_mast_dout_reg[16]/P0001 ,
		_w2453_
	);
	LUT4 #(
		.INIT('h0031)
	) name1719 (
		\wb1_cyc_i_pad ,
		_w869_,
		_w2268_,
		_w2453_,
		_w2454_
	);
	LUT3 #(
		.INIT('hdc)
	) name1720 (
		_w897_,
		_w2452_,
		_w2454_,
		_w2455_
	);
	LUT2 #(
		.INIT('h8)
	) name1721 (
		\wb1_cyc_i_pad ,
		\wb1m_data_i[17]_pad ,
		_w2456_
	);
	LUT2 #(
		.INIT('h4)
	) name1722 (
		_w2268_,
		_w2456_,
		_w2457_
	);
	LUT3 #(
		.INIT('h1b)
	) name1723 (
		\u0_u0_ch_csr_r_reg[2]/NET0131 ,
		\u3_u0_mast_dout_reg[17]/P0001 ,
		\u4_u0_mast_dout_reg[17]/P0001 ,
		_w2458_
	);
	LUT4 #(
		.INIT('h0031)
	) name1724 (
		\wb1_cyc_i_pad ,
		_w869_,
		_w2268_,
		_w2458_,
		_w2459_
	);
	LUT3 #(
		.INIT('hdc)
	) name1725 (
		_w897_,
		_w2457_,
		_w2459_,
		_w2460_
	);
	LUT2 #(
		.INIT('h8)
	) name1726 (
		\wb1_cyc_i_pad ,
		\wb1m_data_i[18]_pad ,
		_w2461_
	);
	LUT2 #(
		.INIT('h4)
	) name1727 (
		_w2268_,
		_w2461_,
		_w2462_
	);
	LUT3 #(
		.INIT('h1b)
	) name1728 (
		\u0_u0_ch_csr_r_reg[2]/NET0131 ,
		\u3_u0_mast_dout_reg[18]/P0001 ,
		\u4_u0_mast_dout_reg[18]/P0001 ,
		_w2463_
	);
	LUT4 #(
		.INIT('h0031)
	) name1729 (
		\wb1_cyc_i_pad ,
		_w869_,
		_w2268_,
		_w2463_,
		_w2464_
	);
	LUT3 #(
		.INIT('hdc)
	) name1730 (
		_w897_,
		_w2462_,
		_w2464_,
		_w2465_
	);
	LUT2 #(
		.INIT('h8)
	) name1731 (
		\wb1_cyc_i_pad ,
		\wb1m_data_i[19]_pad ,
		_w2466_
	);
	LUT2 #(
		.INIT('h4)
	) name1732 (
		_w2268_,
		_w2466_,
		_w2467_
	);
	LUT3 #(
		.INIT('h1b)
	) name1733 (
		\u0_u0_ch_csr_r_reg[2]/NET0131 ,
		\u3_u0_mast_dout_reg[19]/P0001 ,
		\u4_u0_mast_dout_reg[19]/P0001 ,
		_w2468_
	);
	LUT4 #(
		.INIT('h0031)
	) name1734 (
		\wb1_cyc_i_pad ,
		_w869_,
		_w2268_,
		_w2468_,
		_w2469_
	);
	LUT3 #(
		.INIT('hdc)
	) name1735 (
		_w897_,
		_w2467_,
		_w2469_,
		_w2470_
	);
	LUT2 #(
		.INIT('h8)
	) name1736 (
		\wb1_cyc_i_pad ,
		\wb1m_data_i[1]_pad ,
		_w2471_
	);
	LUT2 #(
		.INIT('h4)
	) name1737 (
		_w2268_,
		_w2471_,
		_w2472_
	);
	LUT3 #(
		.INIT('h1b)
	) name1738 (
		\u0_u0_ch_csr_r_reg[2]/NET0131 ,
		\u3_u0_mast_dout_reg[1]/P0001 ,
		\u4_u0_mast_dout_reg[1]/P0001 ,
		_w2473_
	);
	LUT2 #(
		.INIT('h4)
	) name1739 (
		_w869_,
		_w2473_,
		_w2474_
	);
	LUT2 #(
		.INIT('h4)
	) name1740 (
		_w897_,
		_w2474_,
		_w2475_
	);
	LUT2 #(
		.INIT('h4)
	) name1741 (
		\u2_tsz_cnt_reg[1]/NET0131 ,
		_w869_,
		_w2476_
	);
	LUT4 #(
		.INIT('h4000)
	) name1742 (
		\u2_tsz_cnt_reg[1]/NET0131 ,
		_w894_,
		_w895_,
		_w896_,
		_w2477_
	);
	LUT3 #(
		.INIT('h01)
	) name1743 (
		_w2316_,
		_w2476_,
		_w2477_,
		_w2478_
	);
	LUT3 #(
		.INIT('hba)
	) name1744 (
		_w2472_,
		_w2475_,
		_w2478_,
		_w2479_
	);
	LUT2 #(
		.INIT('h8)
	) name1745 (
		\wb1_cyc_i_pad ,
		\wb1m_data_i[20]_pad ,
		_w2480_
	);
	LUT2 #(
		.INIT('h4)
	) name1746 (
		_w2268_,
		_w2480_,
		_w2481_
	);
	LUT3 #(
		.INIT('h1b)
	) name1747 (
		\u0_u0_ch_csr_r_reg[2]/NET0131 ,
		\u3_u0_mast_dout_reg[20]/P0001 ,
		\u4_u0_mast_dout_reg[20]/P0001 ,
		_w2482_
	);
	LUT4 #(
		.INIT('h0031)
	) name1748 (
		\wb1_cyc_i_pad ,
		_w869_,
		_w2268_,
		_w2482_,
		_w2483_
	);
	LUT3 #(
		.INIT('hdc)
	) name1749 (
		_w897_,
		_w2481_,
		_w2483_,
		_w2484_
	);
	LUT2 #(
		.INIT('h8)
	) name1750 (
		\wb1_cyc_i_pad ,
		\wb1m_data_i[21]_pad ,
		_w2485_
	);
	LUT2 #(
		.INIT('h4)
	) name1751 (
		_w2268_,
		_w2485_,
		_w2486_
	);
	LUT3 #(
		.INIT('h1b)
	) name1752 (
		\u0_u0_ch_csr_r_reg[2]/NET0131 ,
		\u3_u0_mast_dout_reg[21]/P0001 ,
		\u4_u0_mast_dout_reg[21]/P0001 ,
		_w2487_
	);
	LUT4 #(
		.INIT('h0031)
	) name1753 (
		\wb1_cyc_i_pad ,
		_w869_,
		_w2268_,
		_w2487_,
		_w2488_
	);
	LUT3 #(
		.INIT('hdc)
	) name1754 (
		_w897_,
		_w2486_,
		_w2488_,
		_w2489_
	);
	LUT2 #(
		.INIT('h8)
	) name1755 (
		\wb1_cyc_i_pad ,
		\wb1m_data_i[22]_pad ,
		_w2490_
	);
	LUT2 #(
		.INIT('h4)
	) name1756 (
		_w2268_,
		_w2490_,
		_w2491_
	);
	LUT3 #(
		.INIT('h1b)
	) name1757 (
		\u0_u0_ch_csr_r_reg[2]/NET0131 ,
		\u3_u0_mast_dout_reg[22]/P0001 ,
		\u4_u0_mast_dout_reg[22]/P0001 ,
		_w2492_
	);
	LUT4 #(
		.INIT('h0031)
	) name1758 (
		\wb1_cyc_i_pad ,
		_w869_,
		_w2268_,
		_w2492_,
		_w2493_
	);
	LUT3 #(
		.INIT('hdc)
	) name1759 (
		_w897_,
		_w2491_,
		_w2493_,
		_w2494_
	);
	LUT2 #(
		.INIT('h8)
	) name1760 (
		\wb1_cyc_i_pad ,
		\wb1m_data_i[23]_pad ,
		_w2495_
	);
	LUT2 #(
		.INIT('h4)
	) name1761 (
		_w2268_,
		_w2495_,
		_w2496_
	);
	LUT3 #(
		.INIT('h1b)
	) name1762 (
		\u0_u0_ch_csr_r_reg[2]/NET0131 ,
		\u3_u0_mast_dout_reg[23]/P0001 ,
		\u4_u0_mast_dout_reg[23]/P0001 ,
		_w2497_
	);
	LUT4 #(
		.INIT('h0031)
	) name1763 (
		\wb1_cyc_i_pad ,
		_w869_,
		_w2268_,
		_w2497_,
		_w2498_
	);
	LUT3 #(
		.INIT('hdc)
	) name1764 (
		_w897_,
		_w2496_,
		_w2498_,
		_w2499_
	);
	LUT2 #(
		.INIT('h8)
	) name1765 (
		\wb1_cyc_i_pad ,
		\wb1m_data_i[24]_pad ,
		_w2500_
	);
	LUT2 #(
		.INIT('h4)
	) name1766 (
		_w2268_,
		_w2500_,
		_w2501_
	);
	LUT3 #(
		.INIT('h1b)
	) name1767 (
		\u0_u0_ch_csr_r_reg[2]/NET0131 ,
		\u3_u0_mast_dout_reg[24]/P0001 ,
		\u4_u0_mast_dout_reg[24]/P0001 ,
		_w2502_
	);
	LUT4 #(
		.INIT('h0031)
	) name1768 (
		\wb1_cyc_i_pad ,
		_w869_,
		_w2268_,
		_w2502_,
		_w2503_
	);
	LUT3 #(
		.INIT('hdc)
	) name1769 (
		_w897_,
		_w2501_,
		_w2503_,
		_w2504_
	);
	LUT2 #(
		.INIT('h8)
	) name1770 (
		\wb1_cyc_i_pad ,
		\wb1m_data_i[25]_pad ,
		_w2505_
	);
	LUT2 #(
		.INIT('h4)
	) name1771 (
		_w2268_,
		_w2505_,
		_w2506_
	);
	LUT3 #(
		.INIT('h1b)
	) name1772 (
		\u0_u0_ch_csr_r_reg[2]/NET0131 ,
		\u3_u0_mast_dout_reg[25]/P0001 ,
		\u4_u0_mast_dout_reg[25]/P0001 ,
		_w2507_
	);
	LUT4 #(
		.INIT('h0031)
	) name1773 (
		\wb1_cyc_i_pad ,
		_w869_,
		_w2268_,
		_w2507_,
		_w2508_
	);
	LUT3 #(
		.INIT('hdc)
	) name1774 (
		_w897_,
		_w2506_,
		_w2508_,
		_w2509_
	);
	LUT2 #(
		.INIT('h8)
	) name1775 (
		\wb1_cyc_i_pad ,
		\wb1m_data_i[26]_pad ,
		_w2510_
	);
	LUT2 #(
		.INIT('h4)
	) name1776 (
		_w2268_,
		_w2510_,
		_w2511_
	);
	LUT3 #(
		.INIT('h1b)
	) name1777 (
		\u0_u0_ch_csr_r_reg[2]/NET0131 ,
		\u3_u0_mast_dout_reg[26]/P0001 ,
		\u4_u0_mast_dout_reg[26]/P0001 ,
		_w2512_
	);
	LUT4 #(
		.INIT('h0031)
	) name1778 (
		\wb1_cyc_i_pad ,
		_w869_,
		_w2268_,
		_w2512_,
		_w2513_
	);
	LUT3 #(
		.INIT('hdc)
	) name1779 (
		_w897_,
		_w2511_,
		_w2513_,
		_w2514_
	);
	LUT2 #(
		.INIT('h8)
	) name1780 (
		\wb1_cyc_i_pad ,
		\wb1m_data_i[27]_pad ,
		_w2515_
	);
	LUT2 #(
		.INIT('h4)
	) name1781 (
		_w2268_,
		_w2515_,
		_w2516_
	);
	LUT3 #(
		.INIT('h1b)
	) name1782 (
		\u0_u0_ch_csr_r_reg[2]/NET0131 ,
		\u3_u0_mast_dout_reg[27]/P0001 ,
		\u4_u0_mast_dout_reg[27]/P0001 ,
		_w2517_
	);
	LUT4 #(
		.INIT('h0031)
	) name1783 (
		\wb1_cyc_i_pad ,
		_w869_,
		_w2268_,
		_w2517_,
		_w2518_
	);
	LUT3 #(
		.INIT('hdc)
	) name1784 (
		_w897_,
		_w2516_,
		_w2518_,
		_w2519_
	);
	LUT2 #(
		.INIT('h8)
	) name1785 (
		\wb1_cyc_i_pad ,
		\wb1m_data_i[28]_pad ,
		_w2520_
	);
	LUT2 #(
		.INIT('h4)
	) name1786 (
		_w2268_,
		_w2520_,
		_w2521_
	);
	LUT3 #(
		.INIT('h1b)
	) name1787 (
		\u0_u0_ch_csr_r_reg[2]/NET0131 ,
		\u3_u0_mast_dout_reg[28]/P0001 ,
		\u4_u0_mast_dout_reg[28]/P0001 ,
		_w2522_
	);
	LUT4 #(
		.INIT('h0031)
	) name1788 (
		\wb1_cyc_i_pad ,
		_w869_,
		_w2268_,
		_w2522_,
		_w2523_
	);
	LUT3 #(
		.INIT('hdc)
	) name1789 (
		_w897_,
		_w2521_,
		_w2523_,
		_w2524_
	);
	LUT2 #(
		.INIT('h8)
	) name1790 (
		\wb1_cyc_i_pad ,
		\wb1m_data_i[29]_pad ,
		_w2525_
	);
	LUT2 #(
		.INIT('h4)
	) name1791 (
		_w2268_,
		_w2525_,
		_w2526_
	);
	LUT3 #(
		.INIT('h1b)
	) name1792 (
		\u0_u0_ch_csr_r_reg[2]/NET0131 ,
		\u3_u0_mast_dout_reg[29]/P0001 ,
		\u4_u0_mast_dout_reg[29]/P0001 ,
		_w2527_
	);
	LUT4 #(
		.INIT('h0031)
	) name1793 (
		\wb1_cyc_i_pad ,
		_w869_,
		_w2268_,
		_w2527_,
		_w2528_
	);
	LUT3 #(
		.INIT('hdc)
	) name1794 (
		_w897_,
		_w2526_,
		_w2528_,
		_w2529_
	);
	LUT2 #(
		.INIT('h8)
	) name1795 (
		\wb1_cyc_i_pad ,
		\wb1m_data_i[2]_pad ,
		_w2530_
	);
	LUT2 #(
		.INIT('h4)
	) name1796 (
		_w2268_,
		_w2530_,
		_w2531_
	);
	LUT3 #(
		.INIT('h1b)
	) name1797 (
		\u0_u0_ch_csr_r_reg[2]/NET0131 ,
		\u3_u0_mast_dout_reg[2]/P0001 ,
		\u4_u0_mast_dout_reg[2]/P0001 ,
		_w2532_
	);
	LUT2 #(
		.INIT('h4)
	) name1798 (
		_w869_,
		_w2532_,
		_w2533_
	);
	LUT2 #(
		.INIT('h4)
	) name1799 (
		_w897_,
		_w2533_,
		_w2534_
	);
	LUT2 #(
		.INIT('h4)
	) name1800 (
		\u2_tsz_cnt_reg[2]/NET0131 ,
		_w869_,
		_w2535_
	);
	LUT4 #(
		.INIT('h4000)
	) name1801 (
		\u2_tsz_cnt_reg[2]/NET0131 ,
		_w894_,
		_w895_,
		_w896_,
		_w2536_
	);
	LUT3 #(
		.INIT('h01)
	) name1802 (
		_w2316_,
		_w2535_,
		_w2536_,
		_w2537_
	);
	LUT3 #(
		.INIT('hba)
	) name1803 (
		_w2531_,
		_w2534_,
		_w2537_,
		_w2538_
	);
	LUT2 #(
		.INIT('h8)
	) name1804 (
		\wb1_cyc_i_pad ,
		\wb1m_data_i[30]_pad ,
		_w2539_
	);
	LUT2 #(
		.INIT('h4)
	) name1805 (
		_w2268_,
		_w2539_,
		_w2540_
	);
	LUT3 #(
		.INIT('h1b)
	) name1806 (
		\u0_u0_ch_csr_r_reg[2]/NET0131 ,
		\u3_u0_mast_dout_reg[30]/P0001 ,
		\u4_u0_mast_dout_reg[30]/P0001 ,
		_w2541_
	);
	LUT4 #(
		.INIT('h0031)
	) name1807 (
		\wb1_cyc_i_pad ,
		_w869_,
		_w2268_,
		_w2541_,
		_w2542_
	);
	LUT3 #(
		.INIT('hdc)
	) name1808 (
		_w897_,
		_w2540_,
		_w2542_,
		_w2543_
	);
	LUT2 #(
		.INIT('h8)
	) name1809 (
		\wb1_cyc_i_pad ,
		\wb1m_data_i[31]_pad ,
		_w2544_
	);
	LUT2 #(
		.INIT('h4)
	) name1810 (
		_w2268_,
		_w2544_,
		_w2545_
	);
	LUT3 #(
		.INIT('h1b)
	) name1811 (
		\u0_u0_ch_csr_r_reg[2]/NET0131 ,
		\u3_u0_mast_dout_reg[31]/P0001 ,
		\u4_u0_mast_dout_reg[31]/P0001 ,
		_w2546_
	);
	LUT4 #(
		.INIT('h0031)
	) name1812 (
		\wb1_cyc_i_pad ,
		_w869_,
		_w2268_,
		_w2546_,
		_w2547_
	);
	LUT3 #(
		.INIT('hdc)
	) name1813 (
		_w897_,
		_w2545_,
		_w2547_,
		_w2548_
	);
	LUT2 #(
		.INIT('h8)
	) name1814 (
		\wb1_cyc_i_pad ,
		\wb1m_data_i[3]_pad ,
		_w2549_
	);
	LUT2 #(
		.INIT('h4)
	) name1815 (
		_w2268_,
		_w2549_,
		_w2550_
	);
	LUT3 #(
		.INIT('h1b)
	) name1816 (
		\u0_u0_ch_csr_r_reg[2]/NET0131 ,
		\u3_u0_mast_dout_reg[3]/P0001 ,
		\u4_u0_mast_dout_reg[3]/P0001 ,
		_w2551_
	);
	LUT2 #(
		.INIT('h4)
	) name1817 (
		_w869_,
		_w2551_,
		_w2552_
	);
	LUT2 #(
		.INIT('h4)
	) name1818 (
		_w897_,
		_w2552_,
		_w2553_
	);
	LUT2 #(
		.INIT('h4)
	) name1819 (
		\u2_tsz_cnt_reg[3]/NET0131 ,
		_w869_,
		_w2554_
	);
	LUT4 #(
		.INIT('h4000)
	) name1820 (
		\u2_tsz_cnt_reg[3]/NET0131 ,
		_w894_,
		_w895_,
		_w896_,
		_w2555_
	);
	LUT3 #(
		.INIT('h01)
	) name1821 (
		_w2316_,
		_w2554_,
		_w2555_,
		_w2556_
	);
	LUT3 #(
		.INIT('hba)
	) name1822 (
		_w2550_,
		_w2553_,
		_w2556_,
		_w2557_
	);
	LUT2 #(
		.INIT('h8)
	) name1823 (
		\wb1_cyc_i_pad ,
		\wb1m_data_i[4]_pad ,
		_w2558_
	);
	LUT2 #(
		.INIT('h4)
	) name1824 (
		_w2268_,
		_w2558_,
		_w2559_
	);
	LUT3 #(
		.INIT('h1b)
	) name1825 (
		\u0_u0_ch_csr_r_reg[2]/NET0131 ,
		\u3_u0_mast_dout_reg[4]/P0001 ,
		\u4_u0_mast_dout_reg[4]/P0001 ,
		_w2560_
	);
	LUT2 #(
		.INIT('h4)
	) name1826 (
		_w869_,
		_w2560_,
		_w2561_
	);
	LUT2 #(
		.INIT('h4)
	) name1827 (
		_w897_,
		_w2561_,
		_w2562_
	);
	LUT2 #(
		.INIT('h4)
	) name1828 (
		\u2_tsz_cnt_reg[4]/NET0131 ,
		_w869_,
		_w2563_
	);
	LUT4 #(
		.INIT('h4000)
	) name1829 (
		\u2_tsz_cnt_reg[4]/NET0131 ,
		_w894_,
		_w895_,
		_w896_,
		_w2564_
	);
	LUT3 #(
		.INIT('h01)
	) name1830 (
		_w2316_,
		_w2563_,
		_w2564_,
		_w2565_
	);
	LUT3 #(
		.INIT('hba)
	) name1831 (
		_w2559_,
		_w2562_,
		_w2565_,
		_w2566_
	);
	LUT2 #(
		.INIT('h8)
	) name1832 (
		\wb1_cyc_i_pad ,
		\wb1m_data_i[5]_pad ,
		_w2567_
	);
	LUT2 #(
		.INIT('h4)
	) name1833 (
		_w2268_,
		_w2567_,
		_w2568_
	);
	LUT3 #(
		.INIT('h1b)
	) name1834 (
		\u0_u0_ch_csr_r_reg[2]/NET0131 ,
		\u3_u0_mast_dout_reg[5]/P0001 ,
		\u4_u0_mast_dout_reg[5]/P0001 ,
		_w2569_
	);
	LUT2 #(
		.INIT('h4)
	) name1835 (
		_w869_,
		_w2569_,
		_w2570_
	);
	LUT2 #(
		.INIT('h4)
	) name1836 (
		_w897_,
		_w2570_,
		_w2571_
	);
	LUT2 #(
		.INIT('h4)
	) name1837 (
		\u2_tsz_cnt_reg[5]/NET0131 ,
		_w869_,
		_w2572_
	);
	LUT4 #(
		.INIT('h4000)
	) name1838 (
		\u2_tsz_cnt_reg[5]/NET0131 ,
		_w894_,
		_w895_,
		_w896_,
		_w2573_
	);
	LUT3 #(
		.INIT('h01)
	) name1839 (
		_w2316_,
		_w2572_,
		_w2573_,
		_w2574_
	);
	LUT3 #(
		.INIT('hba)
	) name1840 (
		_w2568_,
		_w2571_,
		_w2574_,
		_w2575_
	);
	LUT2 #(
		.INIT('h8)
	) name1841 (
		\wb1_cyc_i_pad ,
		\wb1m_data_i[6]_pad ,
		_w2576_
	);
	LUT2 #(
		.INIT('h4)
	) name1842 (
		_w2268_,
		_w2576_,
		_w2577_
	);
	LUT3 #(
		.INIT('h1b)
	) name1843 (
		\u0_u0_ch_csr_r_reg[2]/NET0131 ,
		\u3_u0_mast_dout_reg[6]/P0001 ,
		\u4_u0_mast_dout_reg[6]/P0001 ,
		_w2578_
	);
	LUT2 #(
		.INIT('h4)
	) name1844 (
		_w869_,
		_w2578_,
		_w2579_
	);
	LUT2 #(
		.INIT('h4)
	) name1845 (
		_w897_,
		_w2579_,
		_w2580_
	);
	LUT2 #(
		.INIT('h4)
	) name1846 (
		\u2_tsz_cnt_reg[6]/NET0131 ,
		_w869_,
		_w2581_
	);
	LUT4 #(
		.INIT('h4000)
	) name1847 (
		\u2_tsz_cnt_reg[6]/NET0131 ,
		_w894_,
		_w895_,
		_w896_,
		_w2582_
	);
	LUT3 #(
		.INIT('h01)
	) name1848 (
		_w2316_,
		_w2581_,
		_w2582_,
		_w2583_
	);
	LUT3 #(
		.INIT('hba)
	) name1849 (
		_w2577_,
		_w2580_,
		_w2583_,
		_w2584_
	);
	LUT2 #(
		.INIT('h8)
	) name1850 (
		\wb1_cyc_i_pad ,
		\wb1m_data_i[7]_pad ,
		_w2585_
	);
	LUT2 #(
		.INIT('h4)
	) name1851 (
		_w2268_,
		_w2585_,
		_w2586_
	);
	LUT3 #(
		.INIT('h1b)
	) name1852 (
		\u0_u0_ch_csr_r_reg[2]/NET0131 ,
		\u3_u0_mast_dout_reg[7]/P0001 ,
		\u4_u0_mast_dout_reg[7]/P0001 ,
		_w2587_
	);
	LUT2 #(
		.INIT('h4)
	) name1853 (
		_w869_,
		_w2587_,
		_w2588_
	);
	LUT2 #(
		.INIT('h4)
	) name1854 (
		_w897_,
		_w2588_,
		_w2589_
	);
	LUT2 #(
		.INIT('h4)
	) name1855 (
		\u2_tsz_cnt_reg[7]/NET0131 ,
		_w869_,
		_w2590_
	);
	LUT4 #(
		.INIT('h4000)
	) name1856 (
		\u2_tsz_cnt_reg[7]/NET0131 ,
		_w894_,
		_w895_,
		_w896_,
		_w2591_
	);
	LUT3 #(
		.INIT('h01)
	) name1857 (
		_w2316_,
		_w2590_,
		_w2591_,
		_w2592_
	);
	LUT3 #(
		.INIT('hba)
	) name1858 (
		_w2586_,
		_w2589_,
		_w2592_,
		_w2593_
	);
	LUT2 #(
		.INIT('h8)
	) name1859 (
		\wb1_cyc_i_pad ,
		\wb1m_data_i[8]_pad ,
		_w2594_
	);
	LUT2 #(
		.INIT('h4)
	) name1860 (
		_w2268_,
		_w2594_,
		_w2595_
	);
	LUT3 #(
		.INIT('h1b)
	) name1861 (
		\u0_u0_ch_csr_r_reg[2]/NET0131 ,
		\u3_u0_mast_dout_reg[8]/P0001 ,
		\u4_u0_mast_dout_reg[8]/P0001 ,
		_w2596_
	);
	LUT2 #(
		.INIT('h4)
	) name1862 (
		_w869_,
		_w2596_,
		_w2597_
	);
	LUT2 #(
		.INIT('h4)
	) name1863 (
		_w897_,
		_w2597_,
		_w2598_
	);
	LUT2 #(
		.INIT('h4)
	) name1864 (
		\u2_tsz_cnt_reg[8]/NET0131 ,
		_w869_,
		_w2599_
	);
	LUT4 #(
		.INIT('h4000)
	) name1865 (
		\u2_tsz_cnt_reg[8]/NET0131 ,
		_w894_,
		_w895_,
		_w896_,
		_w2600_
	);
	LUT3 #(
		.INIT('h01)
	) name1866 (
		_w2316_,
		_w2599_,
		_w2600_,
		_w2601_
	);
	LUT3 #(
		.INIT('hba)
	) name1867 (
		_w2595_,
		_w2598_,
		_w2601_,
		_w2602_
	);
	LUT2 #(
		.INIT('h8)
	) name1868 (
		\wb1_cyc_i_pad ,
		\wb1m_data_i[9]_pad ,
		_w2603_
	);
	LUT2 #(
		.INIT('h4)
	) name1869 (
		_w2268_,
		_w2603_,
		_w2604_
	);
	LUT3 #(
		.INIT('h1b)
	) name1870 (
		\u0_u0_ch_csr_r_reg[2]/NET0131 ,
		\u3_u0_mast_dout_reg[9]/P0001 ,
		\u4_u0_mast_dout_reg[9]/P0001 ,
		_w2605_
	);
	LUT2 #(
		.INIT('h4)
	) name1871 (
		_w869_,
		_w2605_,
		_w2606_
	);
	LUT2 #(
		.INIT('h4)
	) name1872 (
		_w897_,
		_w2606_,
		_w2607_
	);
	LUT2 #(
		.INIT('h4)
	) name1873 (
		\u2_tsz_cnt_reg[9]/NET0131 ,
		_w869_,
		_w2608_
	);
	LUT4 #(
		.INIT('h4000)
	) name1874 (
		\u2_tsz_cnt_reg[9]/NET0131 ,
		_w894_,
		_w895_,
		_w896_,
		_w2609_
	);
	LUT3 #(
		.INIT('h01)
	) name1875 (
		_w2316_,
		_w2608_,
		_w2609_,
		_w2610_
	);
	LUT3 #(
		.INIT('hba)
	) name1876 (
		_w2604_,
		_w2607_,
		_w2610_,
		_w2611_
	);
	LUT4 #(
		.INIT('haaca)
	) name1877 (
		\u4_u1_rf_ack_reg/P0001 ,
		\wb0_ack_i_pad ,
		\wb1_cyc_i_pad ,
		_w2268_,
		_w2612_
	);
	LUT2 #(
		.INIT('h8)
	) name1878 (
		\wb0_addr_i[0]_pad ,
		\wb0_cyc_i_pad ,
		_w2613_
	);
	LUT2 #(
		.INIT('h4)
	) name1879 (
		_w2271_,
		_w2613_,
		_w2614_
	);
	LUT4 #(
		.INIT('haaca)
	) name1880 (
		\u2_mast1_adr_reg[10]/P0001 ,
		\wb0_addr_i[10]_pad ,
		\wb0_cyc_i_pad ,
		_w2271_,
		_w2615_
	);
	LUT4 #(
		.INIT('haaca)
	) name1881 (
		\u2_mast1_adr_reg[11]/P0001 ,
		\wb0_addr_i[11]_pad ,
		\wb0_cyc_i_pad ,
		_w2271_,
		_w2616_
	);
	LUT4 #(
		.INIT('haaca)
	) name1882 (
		\u2_mast1_adr_reg[12]/P0001 ,
		\wb0_addr_i[12]_pad ,
		\wb0_cyc_i_pad ,
		_w2271_,
		_w2617_
	);
	LUT4 #(
		.INIT('haaca)
	) name1883 (
		\u2_mast1_adr_reg[13]/P0001 ,
		\wb0_addr_i[13]_pad ,
		\wb0_cyc_i_pad ,
		_w2271_,
		_w2618_
	);
	LUT4 #(
		.INIT('haaca)
	) name1884 (
		\u2_mast1_adr_reg[14]/P0001 ,
		\wb0_addr_i[14]_pad ,
		\wb0_cyc_i_pad ,
		_w2271_,
		_w2619_
	);
	LUT4 #(
		.INIT('haaca)
	) name1885 (
		\u2_mast1_adr_reg[15]/P0001 ,
		\wb0_addr_i[15]_pad ,
		\wb0_cyc_i_pad ,
		_w2271_,
		_w2620_
	);
	LUT4 #(
		.INIT('haaca)
	) name1886 (
		\u2_mast1_adr_reg[16]/P0001 ,
		\wb0_addr_i[16]_pad ,
		\wb0_cyc_i_pad ,
		_w2271_,
		_w2621_
	);
	LUT4 #(
		.INIT('haaca)
	) name1887 (
		\u2_mast1_adr_reg[17]/P0001 ,
		\wb0_addr_i[17]_pad ,
		\wb0_cyc_i_pad ,
		_w2271_,
		_w2622_
	);
	LUT4 #(
		.INIT('haaca)
	) name1888 (
		\u2_mast1_adr_reg[18]/P0001 ,
		\wb0_addr_i[18]_pad ,
		\wb0_cyc_i_pad ,
		_w2271_,
		_w2623_
	);
	LUT4 #(
		.INIT('haaca)
	) name1889 (
		\u2_mast1_adr_reg[19]/P0001 ,
		\wb0_addr_i[19]_pad ,
		\wb0_cyc_i_pad ,
		_w2271_,
		_w2624_
	);
	LUT2 #(
		.INIT('h8)
	) name1890 (
		\wb0_addr_i[1]_pad ,
		\wb0_cyc_i_pad ,
		_w2625_
	);
	LUT2 #(
		.INIT('h4)
	) name1891 (
		_w2271_,
		_w2625_,
		_w2626_
	);
	LUT4 #(
		.INIT('haaca)
	) name1892 (
		\u2_mast1_adr_reg[20]/P0001 ,
		\wb0_addr_i[20]_pad ,
		\wb0_cyc_i_pad ,
		_w2271_,
		_w2627_
	);
	LUT4 #(
		.INIT('haaca)
	) name1893 (
		\u2_mast1_adr_reg[21]/P0001 ,
		\wb0_addr_i[21]_pad ,
		\wb0_cyc_i_pad ,
		_w2271_,
		_w2628_
	);
	LUT4 #(
		.INIT('haaca)
	) name1894 (
		\u2_mast1_adr_reg[22]/P0001 ,
		\wb0_addr_i[22]_pad ,
		\wb0_cyc_i_pad ,
		_w2271_,
		_w2629_
	);
	LUT4 #(
		.INIT('haaca)
	) name1895 (
		\u2_mast1_adr_reg[23]/P0001 ,
		\wb0_addr_i[23]_pad ,
		\wb0_cyc_i_pad ,
		_w2271_,
		_w2630_
	);
	LUT4 #(
		.INIT('haaca)
	) name1896 (
		\u2_mast1_adr_reg[24]/P0001 ,
		\wb0_addr_i[24]_pad ,
		\wb0_cyc_i_pad ,
		_w2271_,
		_w2631_
	);
	LUT4 #(
		.INIT('haaca)
	) name1897 (
		\u2_mast1_adr_reg[25]/P0001 ,
		\wb0_addr_i[25]_pad ,
		\wb0_cyc_i_pad ,
		_w2271_,
		_w2632_
	);
	LUT4 #(
		.INIT('haaca)
	) name1898 (
		\u2_mast1_adr_reg[26]/P0001 ,
		\wb0_addr_i[26]_pad ,
		\wb0_cyc_i_pad ,
		_w2271_,
		_w2633_
	);
	LUT4 #(
		.INIT('haaca)
	) name1899 (
		\u2_mast1_adr_reg[27]/P0001 ,
		\wb0_addr_i[27]_pad ,
		\wb0_cyc_i_pad ,
		_w2271_,
		_w2634_
	);
	LUT3 #(
		.INIT('h15)
	) name1900 (
		\u2_mast1_adr_reg[28]/P0001 ,
		\wb0_addr_i[28]_pad ,
		\wb0_cyc_i_pad ,
		_w2635_
	);
	LUT2 #(
		.INIT('h4)
	) name1901 (
		\wb0_addr_i[28]_pad ,
		\wb0_cyc_i_pad ,
		_w2636_
	);
	LUT3 #(
		.INIT('h23)
	) name1902 (
		_w2271_,
		_w2635_,
		_w2636_,
		_w2637_
	);
	LUT3 #(
		.INIT('h15)
	) name1903 (
		\u2_mast1_adr_reg[29]/P0001 ,
		\wb0_addr_i[29]_pad ,
		\wb0_cyc_i_pad ,
		_w2638_
	);
	LUT2 #(
		.INIT('h4)
	) name1904 (
		\wb0_addr_i[29]_pad ,
		\wb0_cyc_i_pad ,
		_w2639_
	);
	LUT3 #(
		.INIT('h23)
	) name1905 (
		_w2271_,
		_w2638_,
		_w2639_,
		_w2640_
	);
	LUT4 #(
		.INIT('haaca)
	) name1906 (
		\u2_mast1_adr_reg[2]/P0001 ,
		\wb0_addr_i[2]_pad ,
		\wb0_cyc_i_pad ,
		_w2271_,
		_w2641_
	);
	LUT3 #(
		.INIT('h15)
	) name1907 (
		\u2_mast1_adr_reg[30]/P0001 ,
		\wb0_addr_i[30]_pad ,
		\wb0_cyc_i_pad ,
		_w2642_
	);
	LUT2 #(
		.INIT('h4)
	) name1908 (
		\wb0_addr_i[30]_pad ,
		\wb0_cyc_i_pad ,
		_w2643_
	);
	LUT3 #(
		.INIT('h23)
	) name1909 (
		_w2271_,
		_w2642_,
		_w2643_,
		_w2644_
	);
	LUT3 #(
		.INIT('h15)
	) name1910 (
		\u2_mast1_adr_reg[31]/P0001 ,
		\wb0_addr_i[31]_pad ,
		\wb0_cyc_i_pad ,
		_w2645_
	);
	LUT2 #(
		.INIT('h4)
	) name1911 (
		\wb0_addr_i[31]_pad ,
		\wb0_cyc_i_pad ,
		_w2646_
	);
	LUT3 #(
		.INIT('h23)
	) name1912 (
		_w2271_,
		_w2645_,
		_w2646_,
		_w2647_
	);
	LUT4 #(
		.INIT('haaca)
	) name1913 (
		\u2_mast1_adr_reg[3]/P0001 ,
		\wb0_addr_i[3]_pad ,
		\wb0_cyc_i_pad ,
		_w2271_,
		_w2648_
	);
	LUT4 #(
		.INIT('haaca)
	) name1914 (
		\u2_mast1_adr_reg[4]/P0001 ,
		\wb0_addr_i[4]_pad ,
		\wb0_cyc_i_pad ,
		_w2271_,
		_w2649_
	);
	LUT4 #(
		.INIT('haaca)
	) name1915 (
		\u2_mast1_adr_reg[5]/P0001 ,
		\wb0_addr_i[5]_pad ,
		\wb0_cyc_i_pad ,
		_w2271_,
		_w2650_
	);
	LUT4 #(
		.INIT('haaca)
	) name1916 (
		\u2_mast1_adr_reg[6]/P0001 ,
		\wb0_addr_i[6]_pad ,
		\wb0_cyc_i_pad ,
		_w2271_,
		_w2651_
	);
	LUT4 #(
		.INIT('haaca)
	) name1917 (
		\u2_mast1_adr_reg[7]/P0001 ,
		\wb0_addr_i[7]_pad ,
		\wb0_cyc_i_pad ,
		_w2271_,
		_w2652_
	);
	LUT4 #(
		.INIT('haaca)
	) name1918 (
		\u2_mast1_adr_reg[8]/P0001 ,
		\wb0_addr_i[8]_pad ,
		\wb0_cyc_i_pad ,
		_w2271_,
		_w2653_
	);
	LUT4 #(
		.INIT('haaca)
	) name1919 (
		\u2_mast1_adr_reg[9]/P0001 ,
		\wb0_addr_i[9]_pad ,
		\wb0_cyc_i_pad ,
		_w2271_,
		_w2654_
	);
	LUT3 #(
		.INIT('hae)
	) name1920 (
		\u4_u0_mast_cyc_reg/P0001 ,
		\wb0_cyc_i_pad ,
		_w2271_,
		_w2655_
	);
	LUT2 #(
		.INIT('h8)
	) name1921 (
		\wb0_err_i_pad ,
		\wb1_cyc_i_pad ,
		_w2656_
	);
	LUT2 #(
		.INIT('h4)
	) name1922 (
		_w2268_,
		_w2656_,
		_w2657_
	);
	LUT2 #(
		.INIT('h8)
	) name1923 (
		\wb0_rty_i_pad ,
		\wb1_cyc_i_pad ,
		_w2658_
	);
	LUT2 #(
		.INIT('h4)
	) name1924 (
		_w2268_,
		_w2658_,
		_w2659_
	);
	LUT2 #(
		.INIT('h2)
	) name1925 (
		\wb0_cyc_i_pad ,
		\wb0_sel_i[0]_pad ,
		_w2660_
	);
	LUT2 #(
		.INIT('hb)
	) name1926 (
		_w2271_,
		_w2660_,
		_w2661_
	);
	LUT2 #(
		.INIT('h2)
	) name1927 (
		\wb0_cyc_i_pad ,
		\wb0_sel_i[1]_pad ,
		_w2662_
	);
	LUT2 #(
		.INIT('hb)
	) name1928 (
		_w2271_,
		_w2662_,
		_w2663_
	);
	LUT2 #(
		.INIT('h2)
	) name1929 (
		\wb0_cyc_i_pad ,
		\wb0_sel_i[2]_pad ,
		_w2664_
	);
	LUT2 #(
		.INIT('hb)
	) name1930 (
		_w2271_,
		_w2664_,
		_w2665_
	);
	LUT2 #(
		.INIT('h2)
	) name1931 (
		\wb0_cyc_i_pad ,
		\wb0_sel_i[3]_pad ,
		_w2666_
	);
	LUT2 #(
		.INIT('hb)
	) name1932 (
		_w2271_,
		_w2666_,
		_w2667_
	);
	LUT4 #(
		.INIT('haae2)
	) name1933 (
		\u4_u0_mast_stb_reg/P0001 ,
		\wb0_cyc_i_pad ,
		\wb0_stb_i_pad ,
		_w2271_,
		_w2668_
	);
	LUT4 #(
		.INIT('haae2)
	) name1934 (
		\u4_u0_mast_we_r_reg/P0001 ,
		\wb0_cyc_i_pad ,
		\wb0_we_i_pad ,
		_w2271_,
		_w2669_
	);
	LUT2 #(
		.INIT('h8)
	) name1935 (
		\wb0s_data_i[0]_pad ,
		\wb1_cyc_i_pad ,
		_w2670_
	);
	LUT2 #(
		.INIT('h4)
	) name1936 (
		_w2268_,
		_w2670_,
		_w2671_
	);
	LUT2 #(
		.INIT('h8)
	) name1937 (
		\wb0s_data_i[10]_pad ,
		\wb1_cyc_i_pad ,
		_w2672_
	);
	LUT2 #(
		.INIT('h4)
	) name1938 (
		_w2268_,
		_w2672_,
		_w2673_
	);
	LUT2 #(
		.INIT('h8)
	) name1939 (
		\wb0s_data_i[11]_pad ,
		\wb1_cyc_i_pad ,
		_w2674_
	);
	LUT2 #(
		.INIT('h4)
	) name1940 (
		_w2268_,
		_w2674_,
		_w2675_
	);
	LUT2 #(
		.INIT('h8)
	) name1941 (
		\wb0s_data_i[12]_pad ,
		\wb1_cyc_i_pad ,
		_w2676_
	);
	LUT2 #(
		.INIT('h4)
	) name1942 (
		_w2268_,
		_w2676_,
		_w2677_
	);
	LUT2 #(
		.INIT('h8)
	) name1943 (
		\wb0s_data_i[13]_pad ,
		\wb1_cyc_i_pad ,
		_w2678_
	);
	LUT2 #(
		.INIT('h4)
	) name1944 (
		_w2268_,
		_w2678_,
		_w2679_
	);
	LUT2 #(
		.INIT('h8)
	) name1945 (
		\wb0s_data_i[14]_pad ,
		\wb1_cyc_i_pad ,
		_w2680_
	);
	LUT2 #(
		.INIT('h4)
	) name1946 (
		_w2268_,
		_w2680_,
		_w2681_
	);
	LUT2 #(
		.INIT('h8)
	) name1947 (
		\wb0s_data_i[15]_pad ,
		\wb1_cyc_i_pad ,
		_w2682_
	);
	LUT2 #(
		.INIT('h4)
	) name1948 (
		_w2268_,
		_w2682_,
		_w2683_
	);
	LUT2 #(
		.INIT('h8)
	) name1949 (
		\wb0s_data_i[16]_pad ,
		\wb1_cyc_i_pad ,
		_w2684_
	);
	LUT2 #(
		.INIT('h4)
	) name1950 (
		_w2268_,
		_w2684_,
		_w2685_
	);
	LUT2 #(
		.INIT('h8)
	) name1951 (
		\wb0s_data_i[17]_pad ,
		\wb1_cyc_i_pad ,
		_w2686_
	);
	LUT2 #(
		.INIT('h4)
	) name1952 (
		_w2268_,
		_w2686_,
		_w2687_
	);
	LUT2 #(
		.INIT('h8)
	) name1953 (
		\wb0s_data_i[18]_pad ,
		\wb1_cyc_i_pad ,
		_w2688_
	);
	LUT2 #(
		.INIT('h4)
	) name1954 (
		_w2268_,
		_w2688_,
		_w2689_
	);
	LUT2 #(
		.INIT('h8)
	) name1955 (
		\wb0s_data_i[19]_pad ,
		\wb1_cyc_i_pad ,
		_w2690_
	);
	LUT2 #(
		.INIT('h4)
	) name1956 (
		_w2268_,
		_w2690_,
		_w2691_
	);
	LUT2 #(
		.INIT('h8)
	) name1957 (
		\wb0s_data_i[1]_pad ,
		\wb1_cyc_i_pad ,
		_w2692_
	);
	LUT2 #(
		.INIT('h4)
	) name1958 (
		_w2268_,
		_w2692_,
		_w2693_
	);
	LUT2 #(
		.INIT('h8)
	) name1959 (
		\wb0s_data_i[20]_pad ,
		\wb1_cyc_i_pad ,
		_w2694_
	);
	LUT2 #(
		.INIT('h4)
	) name1960 (
		_w2268_,
		_w2694_,
		_w2695_
	);
	LUT2 #(
		.INIT('h8)
	) name1961 (
		\wb0s_data_i[21]_pad ,
		\wb1_cyc_i_pad ,
		_w2696_
	);
	LUT2 #(
		.INIT('h4)
	) name1962 (
		_w2268_,
		_w2696_,
		_w2697_
	);
	LUT2 #(
		.INIT('h8)
	) name1963 (
		\wb0s_data_i[22]_pad ,
		\wb1_cyc_i_pad ,
		_w2698_
	);
	LUT2 #(
		.INIT('h4)
	) name1964 (
		_w2268_,
		_w2698_,
		_w2699_
	);
	LUT2 #(
		.INIT('h8)
	) name1965 (
		\wb0s_data_i[23]_pad ,
		\wb1_cyc_i_pad ,
		_w2700_
	);
	LUT2 #(
		.INIT('h4)
	) name1966 (
		_w2268_,
		_w2700_,
		_w2701_
	);
	LUT2 #(
		.INIT('h8)
	) name1967 (
		\wb0s_data_i[24]_pad ,
		\wb1_cyc_i_pad ,
		_w2702_
	);
	LUT2 #(
		.INIT('h4)
	) name1968 (
		_w2268_,
		_w2702_,
		_w2703_
	);
	LUT2 #(
		.INIT('h8)
	) name1969 (
		\wb0s_data_i[25]_pad ,
		\wb1_cyc_i_pad ,
		_w2704_
	);
	LUT2 #(
		.INIT('h4)
	) name1970 (
		_w2268_,
		_w2704_,
		_w2705_
	);
	LUT2 #(
		.INIT('h8)
	) name1971 (
		\wb0s_data_i[26]_pad ,
		\wb1_cyc_i_pad ,
		_w2706_
	);
	LUT2 #(
		.INIT('h4)
	) name1972 (
		_w2268_,
		_w2706_,
		_w2707_
	);
	LUT2 #(
		.INIT('h8)
	) name1973 (
		\wb0s_data_i[27]_pad ,
		\wb1_cyc_i_pad ,
		_w2708_
	);
	LUT2 #(
		.INIT('h4)
	) name1974 (
		_w2268_,
		_w2708_,
		_w2709_
	);
	LUT2 #(
		.INIT('h8)
	) name1975 (
		\wb0s_data_i[28]_pad ,
		\wb1_cyc_i_pad ,
		_w2710_
	);
	LUT2 #(
		.INIT('h4)
	) name1976 (
		_w2268_,
		_w2710_,
		_w2711_
	);
	LUT2 #(
		.INIT('h8)
	) name1977 (
		\wb0s_data_i[29]_pad ,
		\wb1_cyc_i_pad ,
		_w2712_
	);
	LUT2 #(
		.INIT('h4)
	) name1978 (
		_w2268_,
		_w2712_,
		_w2713_
	);
	LUT2 #(
		.INIT('h8)
	) name1979 (
		\wb0s_data_i[2]_pad ,
		\wb1_cyc_i_pad ,
		_w2714_
	);
	LUT2 #(
		.INIT('h4)
	) name1980 (
		_w2268_,
		_w2714_,
		_w2715_
	);
	LUT2 #(
		.INIT('h8)
	) name1981 (
		\wb0s_data_i[30]_pad ,
		\wb1_cyc_i_pad ,
		_w2716_
	);
	LUT2 #(
		.INIT('h4)
	) name1982 (
		_w2268_,
		_w2716_,
		_w2717_
	);
	LUT2 #(
		.INIT('h8)
	) name1983 (
		\wb0s_data_i[31]_pad ,
		\wb1_cyc_i_pad ,
		_w2718_
	);
	LUT2 #(
		.INIT('h4)
	) name1984 (
		_w2268_,
		_w2718_,
		_w2719_
	);
	LUT2 #(
		.INIT('h8)
	) name1985 (
		\wb0s_data_i[3]_pad ,
		\wb1_cyc_i_pad ,
		_w2720_
	);
	LUT2 #(
		.INIT('h4)
	) name1986 (
		_w2268_,
		_w2720_,
		_w2721_
	);
	LUT2 #(
		.INIT('h8)
	) name1987 (
		\wb0s_data_i[4]_pad ,
		\wb1_cyc_i_pad ,
		_w2722_
	);
	LUT2 #(
		.INIT('h4)
	) name1988 (
		_w2268_,
		_w2722_,
		_w2723_
	);
	LUT2 #(
		.INIT('h8)
	) name1989 (
		\wb0s_data_i[5]_pad ,
		\wb1_cyc_i_pad ,
		_w2724_
	);
	LUT2 #(
		.INIT('h4)
	) name1990 (
		_w2268_,
		_w2724_,
		_w2725_
	);
	LUT2 #(
		.INIT('h8)
	) name1991 (
		\wb0s_data_i[6]_pad ,
		\wb1_cyc_i_pad ,
		_w2726_
	);
	LUT2 #(
		.INIT('h4)
	) name1992 (
		_w2268_,
		_w2726_,
		_w2727_
	);
	LUT2 #(
		.INIT('h8)
	) name1993 (
		\wb0s_data_i[7]_pad ,
		\wb1_cyc_i_pad ,
		_w2728_
	);
	LUT2 #(
		.INIT('h4)
	) name1994 (
		_w2268_,
		_w2728_,
		_w2729_
	);
	LUT2 #(
		.INIT('h8)
	) name1995 (
		\wb0s_data_i[8]_pad ,
		\wb1_cyc_i_pad ,
		_w2730_
	);
	LUT2 #(
		.INIT('h4)
	) name1996 (
		_w2268_,
		_w2730_,
		_w2731_
	);
	LUT2 #(
		.INIT('h8)
	) name1997 (
		\wb0s_data_i[9]_pad ,
		\wb1_cyc_i_pad ,
		_w2732_
	);
	LUT2 #(
		.INIT('h4)
	) name1998 (
		_w2268_,
		_w2732_,
		_w2733_
	);
	LUT4 #(
		.INIT('h08fd)
	) name1999 (
		\wb0_cyc_i_pad ,
		\wb0m_data_i[0]_pad ,
		_w2271_,
		_w2406_,
		_w2734_
	);
	LUT4 #(
		.INIT('h08fd)
	) name2000 (
		\wb0_cyc_i_pad ,
		\wb0m_data_i[10]_pad ,
		_w2271_,
		_w2415_,
		_w2735_
	);
	LUT4 #(
		.INIT('h08fd)
	) name2001 (
		\wb0_cyc_i_pad ,
		\wb0m_data_i[11]_pad ,
		_w2271_,
		_w2424_,
		_w2736_
	);
	LUT4 #(
		.INIT('h08fd)
	) name2002 (
		\wb0_cyc_i_pad ,
		\wb0m_data_i[12]_pad ,
		_w2271_,
		_w2433_,
		_w2737_
	);
	LUT4 #(
		.INIT('h08fd)
	) name2003 (
		\wb0_cyc_i_pad ,
		\wb0m_data_i[13]_pad ,
		_w2271_,
		_w2438_,
		_w2738_
	);
	LUT4 #(
		.INIT('h08fd)
	) name2004 (
		\wb0_cyc_i_pad ,
		\wb0m_data_i[14]_pad ,
		_w2271_,
		_w2443_,
		_w2739_
	);
	LUT4 #(
		.INIT('h08fd)
	) name2005 (
		\wb0_cyc_i_pad ,
		\wb0m_data_i[15]_pad ,
		_w2271_,
		_w2448_,
		_w2740_
	);
	LUT4 #(
		.INIT('h08fd)
	) name2006 (
		\wb0_cyc_i_pad ,
		\wb0m_data_i[16]_pad ,
		_w2271_,
		_w2453_,
		_w2741_
	);
	LUT4 #(
		.INIT('h08fd)
	) name2007 (
		\wb0_cyc_i_pad ,
		\wb0m_data_i[17]_pad ,
		_w2271_,
		_w2458_,
		_w2742_
	);
	LUT4 #(
		.INIT('h08fd)
	) name2008 (
		\wb0_cyc_i_pad ,
		\wb0m_data_i[18]_pad ,
		_w2271_,
		_w2463_,
		_w2743_
	);
	LUT4 #(
		.INIT('h08fd)
	) name2009 (
		\wb0_cyc_i_pad ,
		\wb0m_data_i[19]_pad ,
		_w2271_,
		_w2468_,
		_w2744_
	);
	LUT4 #(
		.INIT('h08fd)
	) name2010 (
		\wb0_cyc_i_pad ,
		\wb0m_data_i[1]_pad ,
		_w2271_,
		_w2473_,
		_w2745_
	);
	LUT4 #(
		.INIT('h08fd)
	) name2011 (
		\wb0_cyc_i_pad ,
		\wb0m_data_i[20]_pad ,
		_w2271_,
		_w2482_,
		_w2746_
	);
	LUT4 #(
		.INIT('h08fd)
	) name2012 (
		\wb0_cyc_i_pad ,
		\wb0m_data_i[21]_pad ,
		_w2271_,
		_w2487_,
		_w2747_
	);
	LUT4 #(
		.INIT('h08fd)
	) name2013 (
		\wb0_cyc_i_pad ,
		\wb0m_data_i[22]_pad ,
		_w2271_,
		_w2492_,
		_w2748_
	);
	LUT4 #(
		.INIT('h08fd)
	) name2014 (
		\wb0_cyc_i_pad ,
		\wb0m_data_i[23]_pad ,
		_w2271_,
		_w2497_,
		_w2749_
	);
	LUT4 #(
		.INIT('h08fd)
	) name2015 (
		\wb0_cyc_i_pad ,
		\wb0m_data_i[24]_pad ,
		_w2271_,
		_w2502_,
		_w2750_
	);
	LUT4 #(
		.INIT('h08fd)
	) name2016 (
		\wb0_cyc_i_pad ,
		\wb0m_data_i[25]_pad ,
		_w2271_,
		_w2507_,
		_w2751_
	);
	LUT4 #(
		.INIT('h08fd)
	) name2017 (
		\wb0_cyc_i_pad ,
		\wb0m_data_i[26]_pad ,
		_w2271_,
		_w2512_,
		_w2752_
	);
	LUT4 #(
		.INIT('h08fd)
	) name2018 (
		\wb0_cyc_i_pad ,
		\wb0m_data_i[27]_pad ,
		_w2271_,
		_w2517_,
		_w2753_
	);
	LUT4 #(
		.INIT('h08fd)
	) name2019 (
		\wb0_cyc_i_pad ,
		\wb0m_data_i[28]_pad ,
		_w2271_,
		_w2522_,
		_w2754_
	);
	LUT4 #(
		.INIT('h08fd)
	) name2020 (
		\wb0_cyc_i_pad ,
		\wb0m_data_i[29]_pad ,
		_w2271_,
		_w2527_,
		_w2755_
	);
	LUT4 #(
		.INIT('h08fd)
	) name2021 (
		\wb0_cyc_i_pad ,
		\wb0m_data_i[2]_pad ,
		_w2271_,
		_w2532_,
		_w2756_
	);
	LUT4 #(
		.INIT('h08fd)
	) name2022 (
		\wb0_cyc_i_pad ,
		\wb0m_data_i[30]_pad ,
		_w2271_,
		_w2541_,
		_w2757_
	);
	LUT4 #(
		.INIT('h08fd)
	) name2023 (
		\wb0_cyc_i_pad ,
		\wb0m_data_i[31]_pad ,
		_w2271_,
		_w2546_,
		_w2758_
	);
	LUT4 #(
		.INIT('h08fd)
	) name2024 (
		\wb0_cyc_i_pad ,
		\wb0m_data_i[3]_pad ,
		_w2271_,
		_w2551_,
		_w2759_
	);
	LUT4 #(
		.INIT('h08fd)
	) name2025 (
		\wb0_cyc_i_pad ,
		\wb0m_data_i[4]_pad ,
		_w2271_,
		_w2560_,
		_w2760_
	);
	LUT4 #(
		.INIT('h08fd)
	) name2026 (
		\wb0_cyc_i_pad ,
		\wb0m_data_i[5]_pad ,
		_w2271_,
		_w2569_,
		_w2761_
	);
	LUT4 #(
		.INIT('h08fd)
	) name2027 (
		\wb0_cyc_i_pad ,
		\wb0m_data_i[6]_pad ,
		_w2271_,
		_w2578_,
		_w2762_
	);
	LUT4 #(
		.INIT('h08fd)
	) name2028 (
		\wb0_cyc_i_pad ,
		\wb0m_data_i[7]_pad ,
		_w2271_,
		_w2587_,
		_w2763_
	);
	LUT4 #(
		.INIT('h08fd)
	) name2029 (
		\wb0_cyc_i_pad ,
		\wb0m_data_i[8]_pad ,
		_w2271_,
		_w2596_,
		_w2764_
	);
	LUT4 #(
		.INIT('h08fd)
	) name2030 (
		\wb0_cyc_i_pad ,
		\wb0m_data_i[9]_pad ,
		_w2271_,
		_w2605_,
		_w2765_
	);
	assign \_al_n0  = 1'b0;
	assign \_al_n1  = 1'b1;
	assign \g22594/_0_  = _w756_ ;
	assign \g22595/_0_  = _w768_ ;
	assign \g22599/_0_  = _w771_ ;
	assign \g22600/_0_  = _w777_ ;
	assign \g22606/_0_  = _w782_ ;
	assign \g22607/_0_  = _w787_ ;
	assign \g22610/_0_  = _w791_ ;
	assign \g22614/_0_  = _w797_ ;
	assign \g22615/_0_  = _w803_ ;
	assign \g22616/_0_  = _w806_ ;
	assign \g22619/_0_  = _w807_ ;
	assign \g22620/_0_  = _w810_ ;
	assign \g22626/_0_  = _w813_ ;
	assign \g22635/_0_  = _w818_ ;
	assign \g22650/_0_  = _w824_ ;
	assign \g22651/_0_  = _w828_ ;
	assign \g22692/_0_  = _w830_ ;
	assign \g22727/_0_  = _w832_ ;
	assign \g22729/_3_  = _w838_ ;
	assign \g22774/_0_  = _w882_ ;
	assign \g22775/_0_  = _w889_ ;
	assign \g22776/_0_  = _w906_ ;
	assign \g22777/_0_  = _w914_ ;
	assign \g22779/_3_  = _w916_ ;
	assign \g22780/_0_  = _w918_ ;
	assign \g22781/_0_  = _w920_ ;
	assign \g22782/_0_  = _w922_ ;
	assign \g22784/_0_  = _w924_ ;
	assign \g22785/_0_  = _w926_ ;
	assign \g22786/_0_  = _w928_ ;
	assign \g22787/_0_  = _w929_ ;
	assign \g22789/_3_  = _w931_ ;
	assign \g22790/_0_  = _w934_ ;
	assign \g22791/_0_  = _w938_ ;
	assign \g22792/_0_  = _w940_ ;
	assign \g22793/_0_  = _w942_ ;
	assign \g22794/_0_  = _w944_ ;
	assign \g22795/_0_  = _w946_ ;
	assign \g22796/_0_  = _w948_ ;
	assign \g22797/_0_  = _w950_ ;
	assign \g22798/_0_  = _w952_ ;
	assign \g22799/_0_  = _w954_ ;
	assign \g22838/_0_  = _w881_ ;
	assign \g22839/_0_  = _w963_ ;
	assign \g22841/_0_  = _w965_ ;
	assign \g22842/_0_  = _w966_ ;
	assign \g22847/_0_  = _w969_ ;
	assign \g22848/_0_  = _w972_ ;
	assign \g22849/_0_  = _w975_ ;
	assign \g22850/_0_  = _w978_ ;
	assign \g22851/_0_  = _w981_ ;
	assign \g22852/_0_  = _w984_ ;
	assign \g22853/_0_  = _w987_ ;
	assign \g22854/_0_  = _w990_ ;
	assign \g22855/_0_  = _w993_ ;
	assign \g22856/_0_  = _w996_ ;
	assign \g22857/_0_  = _w999_ ;
	assign \g22858/_0_  = _w1002_ ;
	assign \g22859/_0_  = _w1005_ ;
	assign \g22860/_0_  = _w1008_ ;
	assign \g22861/_0_  = _w1011_ ;
	assign \g22862/_0_  = _w1014_ ;
	assign \g22863/_0_  = _w1017_ ;
	assign \g22864/_0_  = _w1020_ ;
	assign \g22865/_0_  = _w1023_ ;
	assign \g22867/_0_  = _w1026_ ;
	assign \g22868/_0_  = _w1029_ ;
	assign \g22869/_0_  = _w1032_ ;
	assign \g22871/_0_  = _w1035_ ;
	assign \g22872/_0_  = _w1038_ ;
	assign \g22873/_0_  = _w1041_ ;
	assign \g22874/_0_  = _w1044_ ;
	assign \g22875/_0_  = _w1047_ ;
	assign \g22876/_0_  = _w1050_ ;
	assign \g22878/_0_  = _w1066_ ;
	assign \g22882/_2_  = _w962_ ;
	assign \g22995/_0_  = _w1085_ ;
	assign \g23030/_0_  = _w1096_ ;
	assign \g23046/_0_  = _w1100_ ;
	assign \g23077/_0_  = _w1102_ ;
	assign \g23111/_0_  = _w1103_ ;
	assign \g23115/_1_  = _w1113_ ;
	assign \g23124/_2_  = _w1114_ ;
	assign \g23126/_2_  = _w1115_ ;
	assign \g23128/_2_  = _w1116_ ;
	assign \g23130/_2_  = _w1117_ ;
	assign \g23132/_2_  = _w1118_ ;
	assign \g23134/_2_  = _w1119_ ;
	assign \g23136/_2_  = _w1120_ ;
	assign \g23137/_0_  = _w1121_ ;
	assign \g23140/_2_  = _w1122_ ;
	assign \g23142/_2_  = _w1123_ ;
	assign \g23144/_2_  = _w1124_ ;
	assign \g23146/_2_  = _w1125_ ;
	assign \g23148/_2_  = _w1126_ ;
	assign \g23150/_2_  = _w1127_ ;
	assign \g23152/_2_  = _w1128_ ;
	assign \g23154/_2_  = _w1129_ ;
	assign \g23156/_2_  = _w1130_ ;
	assign \g23158/_2_  = _w1131_ ;
	assign \g23160/_2_  = _w1132_ ;
	assign \g23162/_2_  = _w1133_ ;
	assign \g23163/_3_  = _w1134_ ;
	assign \g23164/_0_  = _w1135_ ;
	assign \g23166/_0_  = _w1136_ ;
	assign \g23168/_0_  = _w1137_ ;
	assign \g23170/_2_  = _w1138_ ;
	assign \g23172/_2_  = _w1139_ ;
	assign \g23174/_2_  = _w1140_ ;
	assign \g23175/_0_  = _w1141_ ;
	assign \g23177/_0_  = _w1142_ ;
	assign \g23180/_2_  = _w1143_ ;
	assign \g23220/_0_  = _w1150_ ;
	assign \g23238/_0_  = _w1152_ ;
	assign \g23239/_0_  = _w1154_ ;
	assign \g23240/_0_  = _w1156_ ;
	assign \g23241/_0_  = _w1158_ ;
	assign \g23242/_0_  = _w1160_ ;
	assign \g23243/_0_  = _w1162_ ;
	assign \g23244/_0_  = _w1164_ ;
	assign \g23245/_0_  = _w1166_ ;
	assign \g23247/_3_  = _w1168_ ;
	assign \g23248/_0_  = _w1170_ ;
	assign \g23249/_0_  = _w1172_ ;
	assign \g23250/_0_  = _w1174_ ;
	assign \g23251/_0_  = _w1176_ ;
	assign \g23252/_0_  = _w1178_ ;
	assign \g23253/_0_  = _w1180_ ;
	assign \g23255/_3_  = _w1182_ ;
	assign \g23260/_0_  = _w1184_ ;
	assign \g23284/_3_  = _w1186_ ;
	assign \g23285/_0_  = _w1189_ ;
	assign \g23334/_0_  = _w1198_ ;
	assign \g23343/_0_  = _w1187_ ;
	assign \g23366/_0_  = _w1207_ ;
	assign \g23402/_0_  = _w1208_ ;
	assign \g23403/_0_  = _w1212_ ;
	assign \g23404/_0_  = _w1215_ ;
	assign \g23405/_0_  = _w1219_ ;
	assign \g23407/_0_  = _w1221_ ;
	assign \g23408/_0_  = _w1225_ ;
	assign \g23409/_0_  = _w1227_ ;
	assign \g23410/_0_  = _w1229_ ;
	assign \g23411/_0_  = _w1233_ ;
	assign \g23413/_2_  = _w1237_ ;
	assign \g23415/_2_  = _w1239_ ;
	assign \g23417/_2_  = _w1241_ ;
	assign \g23542/_0_  = _w955_ ;
	assign \g23607/_0_  = _w1251_ ;
	assign \g23608/_0_  = _w1264_ ;
	assign \g23609/_3_  = _w1271_ ;
	assign \g23707/_0_  = _w1278_ ;
	assign \g23708/_0_  = _w1285_ ;
	assign \g23709/_0_  = _w1292_ ;
	assign \g23710/_0_  = _w1299_ ;
	assign \g23711/_0_  = _w1306_ ;
	assign \g23712/_0_  = _w1313_ ;
	assign \g23713/_0_  = _w1320_ ;
	assign \g23714/_0_  = _w1327_ ;
	assign \g23715/_0_  = _w1334_ ;
	assign \g23716/_0_  = _w1341_ ;
	assign \g23754/_0_  = _w1345_ ;
	assign \g23755/_0_  = _w1349_ ;
	assign \g23756/_0_  = _w1351_ ;
	assign \g23757/_0_  = _w1353_ ;
	assign \g23758/_0_  = _w1355_ ;
	assign \g23759/_0_  = _w1358_ ;
	assign \g23760/_0_  = _w1364_ ;
	assign \g23761/_0_  = _w1367_ ;
	assign \g23763/_3_  = _w1371_ ;
	assign \g23767/_0_  = _w1380_ ;
	assign \g23768/_0_  = _w1389_ ;
	assign \g23833/_0_  = _w1417_ ;
	assign \g23837/_0_  = _w1426_ ;
	assign \g23838/_0_  = _w1434_ ;
	assign \g23839/_0_  = _w1442_ ;
	assign \g23840/_0_  = _w1450_ ;
	assign \g23841/_0_  = _w1458_ ;
	assign \g23842/_0_  = _w1466_ ;
	assign \g23843/_0_  = _w1474_ ;
	assign \g23844/_0_  = _w1482_ ;
	assign \g23845/_0_  = _w1490_ ;
	assign \g23849/_3_  = _w1493_ ;
	assign \g23851/_3_  = _w1496_ ;
	assign \g23858/_0_  = _w1509_ ;
	assign \g23870/_0_  = _w1511_ ;
	assign \g23871/_0_  = _w1513_ ;
	assign \g23872/_3_  = _w1523_ ;
	assign \g23873/_3_  = _w1530_ ;
	assign \g23874/_3_  = _w1537_ ;
	assign \g23875/_3_  = _w1544_ ;
	assign \g23876/_3_  = _w1551_ ;
	assign \g23877/_3_  = _w1558_ ;
	assign \g23878/_3_  = _w1565_ ;
	assign \g23879/_3_  = _w1572_ ;
	assign \g23880/_3_  = _w1579_ ;
	assign \g23881/_3_  = _w1586_ ;
	assign \g23882/_3_  = _w1593_ ;
	assign \g23883/_3_  = _w1600_ ;
	assign \g23884/_3_  = _w1607_ ;
	assign \g23885/_3_  = _w1614_ ;
	assign \g23886/_3_  = _w1621_ ;
	assign \g23887/_3_  = _w1628_ ;
	assign \g23888/_3_  = _w1635_ ;
	assign \g23889/_3_  = _w1642_ ;
	assign \g23890/_3_  = _w1649_ ;
	assign \g23891/_3_  = _w1656_ ;
	assign \g23892/_3_  = _w1667_ ;
	assign \g23893/_3_  = _w1675_ ;
	assign \g23894/_3_  = _w1683_ ;
	assign \g23895/_3_  = _w1691_ ;
	assign \g23896/_3_  = _w1699_ ;
	assign \g23897/_3_  = _w1707_ ;
	assign \g23898/_3_  = _w1715_ ;
	assign \g23899/_3_  = _w1723_ ;
	assign \g23900/_3_  = _w1731_ ;
	assign \g23901/_3_  = _w1739_ ;
	assign \g23902/_3_  = _w1747_ ;
	assign \g23903/_3_  = _w1755_ ;
	assign \g23904/_3_  = _w1763_ ;
	assign \g23905/_3_  = _w1771_ ;
	assign \g23906/_3_  = _w1779_ ;
	assign \g23907/_3_  = _w1787_ ;
	assign \g23908/_3_  = _w1795_ ;
	assign \g23909/_3_  = _w1803_ ;
	assign \g23910/_3_  = _w1811_ ;
	assign \g23911/_3_  = _w1819_ ;
	assign \g23912/_3_  = _w1828_ ;
	assign \g23913/_3_  = _w1835_ ;
	assign \g23914/_3_  = _w1842_ ;
	assign \g23915/_3_  = _w1849_ ;
	assign \g23959/_0_  = _w1857_ ;
	assign \g23961/_0_  = _w1864_ ;
	assign \g23962/_0_  = _w1871_ ;
	assign \g23966/_0_  = _w1878_ ;
	assign \g23967/_0_  = _w1885_ ;
	assign \g23969/_0_  = _w1892_ ;
	assign \g23970/_0_  = _w1899_ ;
	assign \g23971/_0_  = _w1906_ ;
	assign \g23972/_0_  = _w1913_ ;
	assign \g23979/_0_  = _w1920_ ;
	assign \g23987/_0_  = _w1927_ ;
	assign \g23988/_0_  = _w1934_ ;
	assign \g23989/_0_  = _w1941_ ;
	assign \g23990/_0_  = _w1948_ ;
	assign \g24005/_0_  = _w1955_ ;
	assign \g24010/_0_  = _w849_ ;
	assign \g24012/_0_  = _w1962_ ;
	assign \g24013/_0_  = _w1969_ ;
	assign \g24014/_0_  = _w1976_ ;
	assign \g24015/_0_  = _w1983_ ;
	assign \g24016/_0_  = _w1990_ ;
	assign \g24017/_0_  = _w1997_ ;
	assign \g24018/_0_  = _w2004_ ;
	assign \g24019/_0_  = _w2011_ ;
	assign \g24020/_0_  = _w2018_ ;
	assign \g24026/_0_  = _w2027_ ;
	assign \g24027/_0_  = _w2036_ ;
	assign \g24028/_0_  = _w2045_ ;
	assign \g24029/_0_  = _w2053_ ;
	assign \g24030/_0_  = _w2061_ ;
	assign \g24031/_0_  = _w2069_ ;
	assign \g24032/_0_  = _w2077_ ;
	assign \g24033/_0_  = _w2085_ ;
	assign \g24034/_0_  = _w2093_ ;
	assign \g24035/_0_  = _w2101_ ;
	assign \g24036/_0_  = _w2110_ ;
	assign \g24037/_0_  = _w2119_ ;
	assign \g24038/_0_  = _w2128_ ;
	assign \g24039/_0_  = _w2137_ ;
	assign \g24042/_0_  = _w2142_ ;
	assign \g24049/_0_  = _w2145_ ;
	assign \g24063/_0_  = _w2148_ ;
	assign \g24119/_0_  = _w2149_ ;
	assign \g24120/_0_  = _w2150_ ;
	assign \g24357/_0_  = _w1191_ ;
	assign \g24432/_0_  = _w2151_ ;
	assign \g24433/_0_  = _w2152_ ;
	assign \g24437/_0_  = _w2153_ ;
	assign \g24438/_0_  = _w2154_ ;
	assign \g24477/_0_  = _w2155_ ;
	assign \g24491/_0_  = _w2160_ ;
	assign \g24530/_2_  = _w2164_ ;
	assign \g24532/_0_  = _w2165_ ;
	assign \g24534/_0_  = _w2169_ ;
	assign \g24537/_0_  = _w2172_ ;
	assign \g24538/_0_  = _w2175_ ;
	assign \g24539/_0_  = _w2176_ ;
	assign \g24540/_0_  = _w2177_ ;
	assign \g24606/_2_  = _w2180_ ;
	assign \g24612/_0_  = _w2181_ ;
	assign \g24677/_0_  = _w2185_ ;
	assign \g24678/_0_  = _w2189_ ;
	assign \g24679/_0_  = _w2193_ ;
	assign \g24688/_0_  = _w2197_ ;
	assign \g24743/_0_  = _w2199_ ;
	assign \g24847/_0_  = _w2200_ ;
	assign \g24849/_0_  = _w2205_ ;
	assign \g24850/_0_  = _w2208_ ;
	assign \g24854/_0_  = _w2211_ ;
	assign \g24862/_0_  = _w2214_ ;
	assign \g24872/_0_  = _w2217_ ;
	assign \g24873/_0_  = _w2220_ ;
	assign \g24874/_0_  = _w2223_ ;
	assign \g24876/_0_  = _w2226_ ;
	assign \g24879/_0_  = _w2230_ ;
	assign \g24880/_0_  = _w2231_ ;
	assign \g24881/_0_  = _w2232_ ;
	assign \g24882/_0_  = _w2233_ ;
	assign \g24952/_2_  = _w1057_ ;
	assign \g24976/_1_  = _w1254_ ;
	assign \g25003/_0_  = _w2234_ ;
	assign \g25004/_0_  = _w2235_ ;
	assign \g25005/_0_  = _w2236_ ;
	assign \g25006/_0_  = _w2237_ ;
	assign \g25011/_0_  = _w2241_ ;
	assign \g25012/_0_  = _w2244_ ;
	assign \g25013/_0_  = _w2248_ ;
	assign \g25031/_0_  = _w2251_ ;
	assign \g25032/_0_  = _w2254_ ;
	assign \g25033/_0_  = _w2257_ ;
	assign \g25034/_0_  = _w2260_ ;
	assign \g25035/_0_  = _w2263_ ;
	assign \g25153/_2_  = _w2202_ ;
	assign \g25183/_0_  = _w2265_ ;
	assign \g25184/_0_  = _w2267_ ;
	assign \g25224/_0_  = _w2270_ ;
	assign \g25232/_0_  = _w2274_ ;
	assign \g25237/_0_  = _w2276_ ;
	assign \g25241/_2_  = _w1502_ ;
	assign \g25243/_2_  = _w1503_ ;
	assign \g25248/_3_  = _w2238_ ;
	assign \g25261/_0_  = _w2277_ ;
	assign \g25262/_0_  = _w2278_ ;
	assign \g25266/_3_  = _w2280_ ;
	assign \g25267/_0_  = _w2281_ ;
	assign \g25269/_0_  = _w2282_ ;
	assign \g25543/_1_  = _w2283_ ;
	assign \g25602/_3_  = _w2285_ ;
	assign \g25610/_0_  = _w2286_ ;
	assign \g25611/_0_  = _w2287_ ;
	assign \g25841/_0_  = _w2288_ ;
	assign \g25843/_0_  = _w2289_ ;
	assign \g25893/_0_  = _w2290_ ;
	assign \g27013/_0_  = _w2292_ ;
	assign \g27060/_0_  = _w2296_ ;
	assign \g27073/_0_  = _w2298_ ;
	assign \g27184/_0_  = _w876_ ;
	assign \g27186/_0_  = _w857_ ;
	assign \g27189/_2_  = _w859_ ;
	assign \g47/_0_  = _w2307_ ;
	assign \u0_u0_ch_done_reg/_05_  = _w2310_ ;
	assign \u2_adr0_cnt_reg[0]/P0000  = _w212_ ;
	assign \u2_adr1_cnt_reg[0]/P0000  = _w243_ ;
	assign \u3_u0_mast_we_r_reg/_05_  = _w2312_ ;
	assign \wb0_ack_o_pad  = _w2313_ ;
	assign \wb0_addr_o[0]_pad  = _w2315_ ;
	assign \wb0_addr_o[10]_pad  = _w2317_ ;
	assign \wb0_addr_o[11]_pad  = _w2318_ ;
	assign \wb0_addr_o[12]_pad  = _w2319_ ;
	assign \wb0_addr_o[13]_pad  = _w2320_ ;
	assign \wb0_addr_o[14]_pad  = _w2321_ ;
	assign \wb0_addr_o[15]_pad  = _w2322_ ;
	assign \wb0_addr_o[16]_pad  = _w2323_ ;
	assign \wb0_addr_o[17]_pad  = _w2324_ ;
	assign \wb0_addr_o[18]_pad  = _w2325_ ;
	assign \wb0_addr_o[19]_pad  = _w2326_ ;
	assign \wb0_addr_o[1]_pad  = _w2328_ ;
	assign \wb0_addr_o[20]_pad  = _w2329_ ;
	assign \wb0_addr_o[21]_pad  = _w2330_ ;
	assign \wb0_addr_o[22]_pad  = _w2331_ ;
	assign \wb0_addr_o[23]_pad  = _w2332_ ;
	assign \wb0_addr_o[24]_pad  = _w2333_ ;
	assign \wb0_addr_o[25]_pad  = _w2334_ ;
	assign \wb0_addr_o[26]_pad  = _w2335_ ;
	assign \wb0_addr_o[27]_pad  = _w2336_ ;
	assign \wb0_addr_o[28]_pad  = _w2339_ ;
	assign \wb0_addr_o[29]_pad  = _w2342_ ;
	assign \wb0_addr_o[2]_pad  = _w2343_ ;
	assign \wb0_addr_o[30]_pad  = _w2346_ ;
	assign \wb0_addr_o[31]_pad  = _w2349_ ;
	assign \wb0_addr_o[3]_pad  = _w2350_ ;
	assign \wb0_addr_o[4]_pad  = _w2351_ ;
	assign \wb0_addr_o[5]_pad  = _w2352_ ;
	assign \wb0_addr_o[6]_pad  = _w2353_ ;
	assign \wb0_addr_o[7]_pad  = _w2354_ ;
	assign \wb0_addr_o[8]_pad  = _w2355_ ;
	assign \wb0_addr_o[9]_pad  = _w2356_ ;
	assign \wb0_cyc_o_pad  = _w2357_ ;
	assign \wb0_err_o_pad  = _w2359_ ;
	assign \wb0_rty_o_pad  = _w2361_ ;
	assign \wb0_sel_o[0]_pad  = _w2363_ ;
	assign \wb0_sel_o[1]_pad  = _w2365_ ;
	assign \wb0_sel_o[2]_pad  = _w2367_ ;
	assign \wb0_sel_o[3]_pad  = _w2369_ ;
	assign \wb0_stb_o_pad  = _w2370_ ;
	assign \wb0_we_o_pad  = _w2371_ ;
	assign \wb0m_data_o[0]_pad  = _w2372_ ;
	assign \wb0m_data_o[10]_pad  = _w2373_ ;
	assign \wb0m_data_o[11]_pad  = _w2374_ ;
	assign \wb0m_data_o[12]_pad  = _w2375_ ;
	assign \wb0m_data_o[13]_pad  = _w2376_ ;
	assign \wb0m_data_o[14]_pad  = _w2377_ ;
	assign \wb0m_data_o[15]_pad  = _w2378_ ;
	assign \wb0m_data_o[16]_pad  = _w2379_ ;
	assign \wb0m_data_o[17]_pad  = _w2380_ ;
	assign \wb0m_data_o[18]_pad  = _w2381_ ;
	assign \wb0m_data_o[19]_pad  = _w2382_ ;
	assign \wb0m_data_o[1]_pad  = _w2383_ ;
	assign \wb0m_data_o[20]_pad  = _w2384_ ;
	assign \wb0m_data_o[21]_pad  = _w2385_ ;
	assign \wb0m_data_o[22]_pad  = _w2386_ ;
	assign \wb0m_data_o[23]_pad  = _w2387_ ;
	assign \wb0m_data_o[24]_pad  = _w2388_ ;
	assign \wb0m_data_o[25]_pad  = _w2389_ ;
	assign \wb0m_data_o[26]_pad  = _w2390_ ;
	assign \wb0m_data_o[27]_pad  = _w2391_ ;
	assign \wb0m_data_o[28]_pad  = _w2392_ ;
	assign \wb0m_data_o[29]_pad  = _w2393_ ;
	assign \wb0m_data_o[2]_pad  = _w2394_ ;
	assign \wb0m_data_o[30]_pad  = _w2395_ ;
	assign \wb0m_data_o[31]_pad  = _w2396_ ;
	assign \wb0m_data_o[3]_pad  = _w2397_ ;
	assign \wb0m_data_o[4]_pad  = _w2398_ ;
	assign \wb0m_data_o[5]_pad  = _w2399_ ;
	assign \wb0m_data_o[6]_pad  = _w2400_ ;
	assign \wb0m_data_o[7]_pad  = _w2401_ ;
	assign \wb0m_data_o[8]_pad  = _w2402_ ;
	assign \wb0m_data_o[9]_pad  = _w2403_ ;
	assign \wb0s_data_o[0]_pad  = _w2412_ ;
	assign \wb0s_data_o[10]_pad  = _w2421_ ;
	assign \wb0s_data_o[11]_pad  = _w2430_ ;
	assign \wb0s_data_o[12]_pad  = _w2435_ ;
	assign \wb0s_data_o[13]_pad  = _w2440_ ;
	assign \wb0s_data_o[14]_pad  = _w2445_ ;
	assign \wb0s_data_o[15]_pad  = _w2450_ ;
	assign \wb0s_data_o[16]_pad  = _w2455_ ;
	assign \wb0s_data_o[17]_pad  = _w2460_ ;
	assign \wb0s_data_o[18]_pad  = _w2465_ ;
	assign \wb0s_data_o[19]_pad  = _w2470_ ;
	assign \wb0s_data_o[1]_pad  = _w2479_ ;
	assign \wb0s_data_o[20]_pad  = _w2484_ ;
	assign \wb0s_data_o[21]_pad  = _w2489_ ;
	assign \wb0s_data_o[22]_pad  = _w2494_ ;
	assign \wb0s_data_o[23]_pad  = _w2499_ ;
	assign \wb0s_data_o[24]_pad  = _w2504_ ;
	assign \wb0s_data_o[25]_pad  = _w2509_ ;
	assign \wb0s_data_o[26]_pad  = _w2514_ ;
	assign \wb0s_data_o[27]_pad  = _w2519_ ;
	assign \wb0s_data_o[28]_pad  = _w2524_ ;
	assign \wb0s_data_o[29]_pad  = _w2529_ ;
	assign \wb0s_data_o[2]_pad  = _w2538_ ;
	assign \wb0s_data_o[30]_pad  = _w2543_ ;
	assign \wb0s_data_o[31]_pad  = _w2548_ ;
	assign \wb0s_data_o[3]_pad  = _w2557_ ;
	assign \wb0s_data_o[4]_pad  = _w2566_ ;
	assign \wb0s_data_o[5]_pad  = _w2575_ ;
	assign \wb0s_data_o[6]_pad  = _w2584_ ;
	assign \wb0s_data_o[7]_pad  = _w2593_ ;
	assign \wb0s_data_o[8]_pad  = _w2602_ ;
	assign \wb0s_data_o[9]_pad  = _w2611_ ;
	assign \wb1_ack_o_pad  = _w2612_ ;
	assign \wb1_addr_o[0]_pad  = _w2614_ ;
	assign \wb1_addr_o[10]_pad  = _w2615_ ;
	assign \wb1_addr_o[11]_pad  = _w2616_ ;
	assign \wb1_addr_o[12]_pad  = _w2617_ ;
	assign \wb1_addr_o[13]_pad  = _w2618_ ;
	assign \wb1_addr_o[14]_pad  = _w2619_ ;
	assign \wb1_addr_o[15]_pad  = _w2620_ ;
	assign \wb1_addr_o[16]_pad  = _w2621_ ;
	assign \wb1_addr_o[17]_pad  = _w2622_ ;
	assign \wb1_addr_o[18]_pad  = _w2623_ ;
	assign \wb1_addr_o[19]_pad  = _w2624_ ;
	assign \wb1_addr_o[1]_pad  = _w2626_ ;
	assign \wb1_addr_o[20]_pad  = _w2627_ ;
	assign \wb1_addr_o[21]_pad  = _w2628_ ;
	assign \wb1_addr_o[22]_pad  = _w2629_ ;
	assign \wb1_addr_o[23]_pad  = _w2630_ ;
	assign \wb1_addr_o[24]_pad  = _w2631_ ;
	assign \wb1_addr_o[25]_pad  = _w2632_ ;
	assign \wb1_addr_o[26]_pad  = _w2633_ ;
	assign \wb1_addr_o[27]_pad  = _w2634_ ;
	assign \wb1_addr_o[28]_pad  = _w2637_ ;
	assign \wb1_addr_o[29]_pad  = _w2640_ ;
	assign \wb1_addr_o[2]_pad  = _w2641_ ;
	assign \wb1_addr_o[30]_pad  = _w2644_ ;
	assign \wb1_addr_o[31]_pad  = _w2647_ ;
	assign \wb1_addr_o[3]_pad  = _w2648_ ;
	assign \wb1_addr_o[4]_pad  = _w2649_ ;
	assign \wb1_addr_o[5]_pad  = _w2650_ ;
	assign \wb1_addr_o[6]_pad  = _w2651_ ;
	assign \wb1_addr_o[7]_pad  = _w2652_ ;
	assign \wb1_addr_o[8]_pad  = _w2653_ ;
	assign \wb1_addr_o[9]_pad  = _w2654_ ;
	assign \wb1_cyc_o_pad  = _w2655_ ;
	assign \wb1_err_o_pad  = _w2657_ ;
	assign \wb1_rty_o_pad  = _w2659_ ;
	assign \wb1_sel_o[0]_pad  = _w2661_ ;
	assign \wb1_sel_o[1]_pad  = _w2663_ ;
	assign \wb1_sel_o[2]_pad  = _w2665_ ;
	assign \wb1_sel_o[3]_pad  = _w2667_ ;
	assign \wb1_stb_o_pad  = _w2668_ ;
	assign \wb1_we_o_pad  = _w2669_ ;
	assign \wb1m_data_o[0]_pad  = _w2671_ ;
	assign \wb1m_data_o[10]_pad  = _w2673_ ;
	assign \wb1m_data_o[11]_pad  = _w2675_ ;
	assign \wb1m_data_o[12]_pad  = _w2677_ ;
	assign \wb1m_data_o[13]_pad  = _w2679_ ;
	assign \wb1m_data_o[14]_pad  = _w2681_ ;
	assign \wb1m_data_o[15]_pad  = _w2683_ ;
	assign \wb1m_data_o[16]_pad  = _w2685_ ;
	assign \wb1m_data_o[17]_pad  = _w2687_ ;
	assign \wb1m_data_o[18]_pad  = _w2689_ ;
	assign \wb1m_data_o[19]_pad  = _w2691_ ;
	assign \wb1m_data_o[1]_pad  = _w2693_ ;
	assign \wb1m_data_o[20]_pad  = _w2695_ ;
	assign \wb1m_data_o[21]_pad  = _w2697_ ;
	assign \wb1m_data_o[22]_pad  = _w2699_ ;
	assign \wb1m_data_o[23]_pad  = _w2701_ ;
	assign \wb1m_data_o[24]_pad  = _w2703_ ;
	assign \wb1m_data_o[25]_pad  = _w2705_ ;
	assign \wb1m_data_o[26]_pad  = _w2707_ ;
	assign \wb1m_data_o[27]_pad  = _w2709_ ;
	assign \wb1m_data_o[28]_pad  = _w2711_ ;
	assign \wb1m_data_o[29]_pad  = _w2713_ ;
	assign \wb1m_data_o[2]_pad  = _w2715_ ;
	assign \wb1m_data_o[30]_pad  = _w2717_ ;
	assign \wb1m_data_o[31]_pad  = _w2719_ ;
	assign \wb1m_data_o[3]_pad  = _w2721_ ;
	assign \wb1m_data_o[4]_pad  = _w2723_ ;
	assign \wb1m_data_o[5]_pad  = _w2725_ ;
	assign \wb1m_data_o[6]_pad  = _w2727_ ;
	assign \wb1m_data_o[7]_pad  = _w2729_ ;
	assign \wb1m_data_o[8]_pad  = _w2731_ ;
	assign \wb1m_data_o[9]_pad  = _w2733_ ;
	assign \wb1s_data_o[0]_pad  = _w2734_ ;
	assign \wb1s_data_o[10]_pad  = _w2735_ ;
	assign \wb1s_data_o[11]_pad  = _w2736_ ;
	assign \wb1s_data_o[12]_pad  = _w2737_ ;
	assign \wb1s_data_o[13]_pad  = _w2738_ ;
	assign \wb1s_data_o[14]_pad  = _w2739_ ;
	assign \wb1s_data_o[15]_pad  = _w2740_ ;
	assign \wb1s_data_o[16]_pad  = _w2741_ ;
	assign \wb1s_data_o[17]_pad  = _w2742_ ;
	assign \wb1s_data_o[18]_pad  = _w2743_ ;
	assign \wb1s_data_o[19]_pad  = _w2744_ ;
	assign \wb1s_data_o[1]_pad  = _w2745_ ;
	assign \wb1s_data_o[20]_pad  = _w2746_ ;
	assign \wb1s_data_o[21]_pad  = _w2747_ ;
	assign \wb1s_data_o[22]_pad  = _w2748_ ;
	assign \wb1s_data_o[23]_pad  = _w2749_ ;
	assign \wb1s_data_o[24]_pad  = _w2750_ ;
	assign \wb1s_data_o[25]_pad  = _w2751_ ;
	assign \wb1s_data_o[26]_pad  = _w2752_ ;
	assign \wb1s_data_o[27]_pad  = _w2753_ ;
	assign \wb1s_data_o[28]_pad  = _w2754_ ;
	assign \wb1s_data_o[29]_pad  = _w2755_ ;
	assign \wb1s_data_o[2]_pad  = _w2756_ ;
	assign \wb1s_data_o[30]_pad  = _w2757_ ;
	assign \wb1s_data_o[31]_pad  = _w2758_ ;
	assign \wb1s_data_o[3]_pad  = _w2759_ ;
	assign \wb1s_data_o[4]_pad  = _w2760_ ;
	assign \wb1s_data_o[5]_pad  = _w2761_ ;
	assign \wb1s_data_o[6]_pad  = _w2762_ ;
	assign \wb1s_data_o[7]_pad  = _w2763_ ;
	assign \wb1s_data_o[8]_pad  = _w2764_ ;
	assign \wb1s_data_o[9]_pad  = _w2765_ ;
endmodule;