module top( \a0_pad  , a_pad , \b0_pad  , b_pad , \c0_pad  , c_pad , \d0_pad  , d_pad , \e0_pad  , e_pad , \f0_pad  , f_pad , g_pad , h_pad , i_pad , j_pad , k_pad , l_pad , m_pad , n_pad , o_pad , p_pad , q_pad , r_pad , s_pad , t_pad , u_pad , v_pad , w_pad , x_pad , y_pad , z_pad , \g0_pad  , \h0_pad  , \i0_pad  );
  input \a0_pad  ;
  input a_pad ;
  input \b0_pad  ;
  input b_pad ;
  input \c0_pad  ;
  input c_pad ;
  input \d0_pad  ;
  input d_pad ;
  input \e0_pad  ;
  input e_pad ;
  input \f0_pad  ;
  input f_pad ;
  input g_pad ;
  input h_pad ;
  input i_pad ;
  input j_pad ;
  input k_pad ;
  input l_pad ;
  input m_pad ;
  input n_pad ;
  input o_pad ;
  input p_pad ;
  input q_pad ;
  input r_pad ;
  input s_pad ;
  input t_pad ;
  input u_pad ;
  input v_pad ;
  input w_pad ;
  input x_pad ;
  input y_pad ;
  input z_pad ;
  output \g0_pad  ;
  output \h0_pad  ;
  output \i0_pad  ;
  wire n33 , n34 , n35 , n36 , n37 , n38 , n39 , n40 , n41 , n42 , n43 , n44 , n45 , n46 , n47 , n48 , n49 , n50 , n51 , n52 , n53 , n54 , n55 , n56 , n57 , n58 , n59 , n60 , n61 , n62 , n63 , n64 , n65 , n66 , n67 , n68 , n69 , n70 , n71 , n72 , n73 , n74 , n75 , n76 , n77 , n78 , n79 , n80 , n81 , n82 , n83 , n84 , n85 , n86 , n87 , n88 , n89 , n90 , n91 , n92 , n93 , n94 , n95 , n96 , n97 , n98 , n99 , n100 , n101 , n102 , n103 , n104 , n105 , n106 , n107 , n108 , n109 , n110 , n111 , n112 , n113 , n114 , n115 , n116 ;
  assign n38 = ~i_pad & y_pad ;
  assign n36 = \b0_pad  & ~l_pad ;
  assign n37 = \c0_pad  & ~m_pad ;
  assign n45 = ~n36 & ~n37 ;
  assign n46 = ~n38 & n45 ;
  assign n42 = ~\a0_pad  & k_pad ;
  assign n43 = ~\b0_pad  & l_pad ;
  assign n44 = ~n42 & ~n43 ;
  assign n33 = j_pad & ~z_pad ;
  assign n34 = i_pad & ~y_pad ;
  assign n35 = ~n33 & ~n34 ;
  assign n39 = \a0_pad  & ~k_pad ;
  assign n40 = ~j_pad & z_pad ;
  assign n41 = ~n39 & ~n40 ;
  assign n47 = n35 & n41 ;
  assign n48 = n44 & n47 ;
  assign n49 = n46 & n48 ;
  assign n51 = ~\e0_pad  & o_pad ;
  assign n52 = ~\f0_pad  & p_pad ;
  assign n53 = ~n51 & ~n52 ;
  assign n54 = \e0_pad  & ~o_pad ;
  assign n55 = \d0_pad  & ~n_pad ;
  assign n56 = ~n54 & ~n55 ;
  assign n57 = ~n53 & n56 ;
  assign n50 = ~\c0_pad  & m_pad ;
  assign n58 = ~\d0_pad  & n_pad ;
  assign n59 = ~n50 & ~n58 ;
  assign n60 = ~n57 & n59 ;
  assign n61 = n49 & ~n60 ;
  assign n62 = n41 & ~n44 ;
  assign n63 = n35 & ~n62 ;
  assign n64 = ~n38 & ~n63 ;
  assign n65 = ~n61 & ~n64 ;
  assign n82 = ~a_pad & q_pad ;
  assign n79 = b_pad & ~r_pad ;
  assign n80 = a_pad & ~q_pad ;
  assign n81 = ~n79 & ~n80 ;
  assign n84 = c_pad & ~s_pad ;
  assign n85 = d_pad & ~t_pad ;
  assign n86 = ~n84 & ~n85 ;
  assign n87 = ~c_pad & s_pad ;
  assign n88 = ~b_pad & r_pad ;
  assign n89 = ~n87 & ~n88 ;
  assign n94 = ~n86 & n89 ;
  assign n95 = n81 & ~n94 ;
  assign n96 = ~n82 & ~n95 ;
  assign n66 = ~e_pad & u_pad ;
  assign n67 = e_pad & ~u_pad ;
  assign n68 = f_pad & ~v_pad ;
  assign n69 = ~n67 & ~n68 ;
  assign n70 = g_pad & ~w_pad ;
  assign n71 = h_pad & ~x_pad ;
  assign n72 = ~n70 & ~n71 ;
  assign n73 = ~f_pad & v_pad ;
  assign n74 = ~g_pad & w_pad ;
  assign n75 = ~n73 & ~n74 ;
  assign n76 = ~n72 & n75 ;
  assign n77 = n69 & ~n76 ;
  assign n78 = ~n66 & ~n77 ;
  assign n83 = ~d_pad & t_pad ;
  assign n90 = ~n82 & ~n83 ;
  assign n91 = n81 & n90 ;
  assign n92 = n86 & n89 ;
  assign n93 = n91 & n92 ;
  assign n97 = ~h_pad & x_pad ;
  assign n98 = ~n66 & ~n97 ;
  assign n99 = n69 & n98 ;
  assign n100 = n72 & n75 ;
  assign n101 = n99 & n100 ;
  assign n102 = n93 & n101 ;
  assign n103 = ~n78 & n102 ;
  assign n104 = ~n96 & n103 ;
  assign n105 = ~n65 & n104 ;
  assign n106 = n78 & n93 ;
  assign n107 = ~n96 & ~n106 ;
  assign n108 = ~n105 & n107 ;
  assign n109 = \f0_pad  & ~p_pad ;
  assign n110 = n53 & ~n109 ;
  assign n111 = n56 & n110 ;
  assign n112 = n60 & n111 ;
  assign n113 = n49 & n112 ;
  assign n114 = ~n64 & n113 ;
  assign n115 = n104 & n114 ;
  assign n116 = n108 & ~n115 ;
  assign \g0_pad  = n116 ;
  assign \h0_pad  = n115 ;
  assign \i0_pad  = ~n108 ;
endmodule
