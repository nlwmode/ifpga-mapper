module top( \g102_pad  , \g10_reg/NET0131  , \g11_reg/NET0131  , \g1293_pad  , \g14_reg/NET0131  , \g15_reg/NET0131  , \g18_reg/NET0131  , \g197_reg/NET0131  , \g19_reg/NET0131  , \g1_reg/NET0131  , \g204_reg/NET0131  , \g205_reg/NET0131  , \g206_reg/NET0131  , \g207_reg/NET0131  , \g208_reg/NET0131  , \g209_reg/NET0131  , \g210_reg/NET0131  , \g211_reg/NET0131  , \g212_reg/NET0131  , \g218_reg/NET0131  , \g224_reg/NET0131  , \g230_reg/NET0131  , \g236_reg/NET0131  , \g242_reg/NET0131  , \g248_reg/NET0131  , \g24_reg/NET0131  , \g254_reg/NET0131  , \g25_reg/NET0131  , \g260_reg/NET0131  , \g266_reg/NET0131  , \g269_reg/NET0131  , \g276_reg/NET0131  , \g277_reg/NET0131  , \g278_reg/NET0131  , \g279_reg/NET0131  , \g280_reg/NET0131  , \g281_reg/NET0131  , \g282_reg/NET0131  , \g283_reg/NET0131  , \g28_reg/NET0131  , \g293_reg/NET0131  , \g297_reg/NET0131  , \g29_reg/NET0131  , \g2_reg/NET0131  , \g33_reg/NET0131  , \g3_reg/NET0131  , \g402_reg/NET0131  , \g406_reg/NET0131  , \g4099_pad  , \g4100_pad  , \g4101_pad  , \g4102_pad  , \g4103_pad  , \g4104_pad  , \g4105_pad  , \g4108_pad  , \g410_reg/NET0131  , \g4110_pad  , \g4112_pad  , \g414_reg/NET0131  , \g418_reg/NET0131  , \g422_reg/NET0131  , \g426_reg/NET0131  , \g430_reg/NET0131  , \g434_reg/NET0131  , \g437_reg/NET0131  , \g441_reg/NET0131  , \g4422_pad  , \g445_reg/NET0131  , \g449_reg/NET0131  , \g453_reg/NET0131  , \g457_reg/NET0131  , \g461_reg/NET0131  , \g465_reg/NET0131  , \g471_reg/NET0131  , \g478_reg/NET0131  , \g486_reg/NET0131  , \g489_reg/NET0131  , \g48_reg/NET0131  , \g492_reg/NET0131  , \g496_reg/NET0131  , \g500_reg/NET0131  , \g504_reg/NET0131  , \g508_reg/NET0131  , \g512_reg/NET0131  , \g536_reg/NET0131  , \g541_reg/NET0131  , \g545_reg/NET0131  , \g548_reg/NET0131  , \g551_reg/NET0131  , \g554_reg/NET0131  , \g557_pad  , \g558_pad  , \g559_pad  , \g560_pad  , \g561_pad  , \g562_pad  , \g563_pad  , \g567_pad  , \g571_reg/NET0131  , \g574_reg/NET0131  , \g578_reg/NET0131  , \g582_reg/NET0131  , \g586_reg/NET0131  , \g590_reg/NET0131  , \g594_reg/NET0131  , \g598_reg/NET0131  , \g602_reg/NET0131  , \g606_reg/NET0131  , \g610_reg/NET0131  , \g613_reg/NET0131  , \g616_reg/NET0131  , \g619_reg/NET0131  , \g622_reg/NET0131  , \g625_reg/NET0131  , \g628_reg/NET0131  , \g631_reg/NET0131  , \g634_reg/NET0131  , \g638_reg/NET0131  , \g639_pad  , \g642_reg/NET0131  , \g646_reg/NET0131  , \g650_reg/NET0131  , \g654_reg/NET0131  , \g662_reg/NET0131  , \g669_reg/NET0131  , \g672_reg/NET0131  , \g675_reg/NET0131  , \g676_reg/NET0131  , \g677_reg/NET0131  , \g678_reg/NET0131  , \g679_reg/NET0131  , \g680_reg/NET0131  , \g681_reg/NET0131  , \g682_reg/NET0131  , \g683_reg/NET0131  , \g684_reg/NET0131  , \g685_reg/NET0131  , \g687_reg/NET0131  , \g688_reg/NET0131  , \g689_reg/NET0131  , \g698_reg/NET0131  , \g6_reg/NET0131  , \g702_pad  , \g7_reg/NET0131  , \g89_pad  , \_al_n1  , \g10560/_0_  , \g10562/_1_  , \g10564/_1_  , \g10566/_1_  , \g10567/_0_  , \g10569/_1_  , \g10580/_0_  , \g10616/_2_  , \g10627/_2_  , \g10628/_0_  , \g10629/_2_  , \g10630/_2_  , \g10633/_2_  , \g10635/_2_  , \g10636/_2_  , \g10637/_2_  , \g10641/_0_  , \g10649/_0_  , \g10672/_0_  , \g10673/_0_  , \g10680/_0_  , \g10683/_0_  , \g10686/_0_  , \g10695/_0_  , \g10700/_0_  , \g10703/_0_  , \g10704/_0_  , \g10748/_0_  , \g10750/_2_  , \g10757/_0_  , \g10758/_0_  , \g10782/_0_  , \g10826/_0_  , \g10827/_0_  , \g10828/_1_  , \g10832/_2_  , \g10834/_2_  , \g10836/_0_  , \g10837/_1__syn_2  , \g10868/_0_  , \g10904/_0_  , \g10913/_0_  , \g10915/_0_  , \g10922/_0_  , \g10938/_0_  , \g10939/_0_  , \g10940/_0_  , \g10941/_0_  , \g10942/_0_  , \g10944/_2_  , \g10977/_0_  , \g10980/_0_  , \g11020/_0_  , \g11028/_0_  , \g11051/_0_  , \g11057/_0_  , \g11109/_0_  , \g11113/_2_  , \g11156/_0_  , \g11172/_3_  , \g11193/_0_  , \g11219/_0_  , \g11355/_0_  , \g11384/_0_  , \g11442/_0_  , \g11448/_0_  , \g11558/_0_  , \g11559/_0_  , \g11824/_1_  , \g11853/_0_  , \g11854/_0_  , \g11977/_0_  , \g11981/_0_  , \g2584_pad  , \g4121_pad  , \g4809_pad  , \g5692_pad  , \g6282_pad  , \g6284_pad  , \g6360_pad  , \g6362_pad  , \g6364_pad  , \g6366_pad  , \g6368_pad  , \g6370_pad  , \g6372_pad  , \g6374_pad  );
  input \g102_pad  ;
  input \g10_reg/NET0131  ;
  input \g11_reg/NET0131  ;
  input \g1293_pad  ;
  input \g14_reg/NET0131  ;
  input \g15_reg/NET0131  ;
  input \g18_reg/NET0131  ;
  input \g197_reg/NET0131  ;
  input \g19_reg/NET0131  ;
  input \g1_reg/NET0131  ;
  input \g204_reg/NET0131  ;
  input \g205_reg/NET0131  ;
  input \g206_reg/NET0131  ;
  input \g207_reg/NET0131  ;
  input \g208_reg/NET0131  ;
  input \g209_reg/NET0131  ;
  input \g210_reg/NET0131  ;
  input \g211_reg/NET0131  ;
  input \g212_reg/NET0131  ;
  input \g218_reg/NET0131  ;
  input \g224_reg/NET0131  ;
  input \g230_reg/NET0131  ;
  input \g236_reg/NET0131  ;
  input \g242_reg/NET0131  ;
  input \g248_reg/NET0131  ;
  input \g24_reg/NET0131  ;
  input \g254_reg/NET0131  ;
  input \g25_reg/NET0131  ;
  input \g260_reg/NET0131  ;
  input \g266_reg/NET0131  ;
  input \g269_reg/NET0131  ;
  input \g276_reg/NET0131  ;
  input \g277_reg/NET0131  ;
  input \g278_reg/NET0131  ;
  input \g279_reg/NET0131  ;
  input \g280_reg/NET0131  ;
  input \g281_reg/NET0131  ;
  input \g282_reg/NET0131  ;
  input \g283_reg/NET0131  ;
  input \g28_reg/NET0131  ;
  input \g293_reg/NET0131  ;
  input \g297_reg/NET0131  ;
  input \g29_reg/NET0131  ;
  input \g2_reg/NET0131  ;
  input \g33_reg/NET0131  ;
  input \g3_reg/NET0131  ;
  input \g402_reg/NET0131  ;
  input \g406_reg/NET0131  ;
  input \g4099_pad  ;
  input \g4100_pad  ;
  input \g4101_pad  ;
  input \g4102_pad  ;
  input \g4103_pad  ;
  input \g4104_pad  ;
  input \g4105_pad  ;
  input \g4108_pad  ;
  input \g410_reg/NET0131  ;
  input \g4110_pad  ;
  input \g4112_pad  ;
  input \g414_reg/NET0131  ;
  input \g418_reg/NET0131  ;
  input \g422_reg/NET0131  ;
  input \g426_reg/NET0131  ;
  input \g430_reg/NET0131  ;
  input \g434_reg/NET0131  ;
  input \g437_reg/NET0131  ;
  input \g441_reg/NET0131  ;
  input \g4422_pad  ;
  input \g445_reg/NET0131  ;
  input \g449_reg/NET0131  ;
  input \g453_reg/NET0131  ;
  input \g457_reg/NET0131  ;
  input \g461_reg/NET0131  ;
  input \g465_reg/NET0131  ;
  input \g471_reg/NET0131  ;
  input \g478_reg/NET0131  ;
  input \g486_reg/NET0131  ;
  input \g489_reg/NET0131  ;
  input \g48_reg/NET0131  ;
  input \g492_reg/NET0131  ;
  input \g496_reg/NET0131  ;
  input \g500_reg/NET0131  ;
  input \g504_reg/NET0131  ;
  input \g508_reg/NET0131  ;
  input \g512_reg/NET0131  ;
  input \g536_reg/NET0131  ;
  input \g541_reg/NET0131  ;
  input \g545_reg/NET0131  ;
  input \g548_reg/NET0131  ;
  input \g551_reg/NET0131  ;
  input \g554_reg/NET0131  ;
  input \g557_pad  ;
  input \g558_pad  ;
  input \g559_pad  ;
  input \g560_pad  ;
  input \g561_pad  ;
  input \g562_pad  ;
  input \g563_pad  ;
  input \g567_pad  ;
  input \g571_reg/NET0131  ;
  input \g574_reg/NET0131  ;
  input \g578_reg/NET0131  ;
  input \g582_reg/NET0131  ;
  input \g586_reg/NET0131  ;
  input \g590_reg/NET0131  ;
  input \g594_reg/NET0131  ;
  input \g598_reg/NET0131  ;
  input \g602_reg/NET0131  ;
  input \g606_reg/NET0131  ;
  input \g610_reg/NET0131  ;
  input \g613_reg/NET0131  ;
  input \g616_reg/NET0131  ;
  input \g619_reg/NET0131  ;
  input \g622_reg/NET0131  ;
  input \g625_reg/NET0131  ;
  input \g628_reg/NET0131  ;
  input \g631_reg/NET0131  ;
  input \g634_reg/NET0131  ;
  input \g638_reg/NET0131  ;
  input \g639_pad  ;
  input \g642_reg/NET0131  ;
  input \g646_reg/NET0131  ;
  input \g650_reg/NET0131  ;
  input \g654_reg/NET0131  ;
  input \g662_reg/NET0131  ;
  input \g669_reg/NET0131  ;
  input \g672_reg/NET0131  ;
  input \g675_reg/NET0131  ;
  input \g676_reg/NET0131  ;
  input \g677_reg/NET0131  ;
  input \g678_reg/NET0131  ;
  input \g679_reg/NET0131  ;
  input \g680_reg/NET0131  ;
  input \g681_reg/NET0131  ;
  input \g682_reg/NET0131  ;
  input \g683_reg/NET0131  ;
  input \g684_reg/NET0131  ;
  input \g685_reg/NET0131  ;
  input \g687_reg/NET0131  ;
  input \g688_reg/NET0131  ;
  input \g689_reg/NET0131  ;
  input \g698_reg/NET0131  ;
  input \g6_reg/NET0131  ;
  input \g702_pad  ;
  input \g7_reg/NET0131  ;
  input \g89_pad  ;
  output \_al_n1  ;
  output \g10560/_0_  ;
  output \g10562/_1_  ;
  output \g10564/_1_  ;
  output \g10566/_1_  ;
  output \g10567/_0_  ;
  output \g10569/_1_  ;
  output \g10580/_0_  ;
  output \g10616/_2_  ;
  output \g10627/_2_  ;
  output \g10628/_0_  ;
  output \g10629/_2_  ;
  output \g10630/_2_  ;
  output \g10633/_2_  ;
  output \g10635/_2_  ;
  output \g10636/_2_  ;
  output \g10637/_2_  ;
  output \g10641/_0_  ;
  output \g10649/_0_  ;
  output \g10672/_0_  ;
  output \g10673/_0_  ;
  output \g10680/_0_  ;
  output \g10683/_0_  ;
  output \g10686/_0_  ;
  output \g10695/_0_  ;
  output \g10700/_0_  ;
  output \g10703/_0_  ;
  output \g10704/_0_  ;
  output \g10748/_0_  ;
  output \g10750/_2_  ;
  output \g10757/_0_  ;
  output \g10758/_0_  ;
  output \g10782/_0_  ;
  output \g10826/_0_  ;
  output \g10827/_0_  ;
  output \g10828/_1_  ;
  output \g10832/_2_  ;
  output \g10834/_2_  ;
  output \g10836/_0_  ;
  output \g10837/_1__syn_2  ;
  output \g10868/_0_  ;
  output \g10904/_0_  ;
  output \g10913/_0_  ;
  output \g10915/_0_  ;
  output \g10922/_0_  ;
  output \g10938/_0_  ;
  output \g10939/_0_  ;
  output \g10940/_0_  ;
  output \g10941/_0_  ;
  output \g10942/_0_  ;
  output \g10944/_2_  ;
  output \g10977/_0_  ;
  output \g10980/_0_  ;
  output \g11020/_0_  ;
  output \g11028/_0_  ;
  output \g11051/_0_  ;
  output \g11057/_0_  ;
  output \g11109/_0_  ;
  output \g11113/_2_  ;
  output \g11156/_0_  ;
  output \g11172/_3_  ;
  output \g11193/_0_  ;
  output \g11219/_0_  ;
  output \g11355/_0_  ;
  output \g11384/_0_  ;
  output \g11442/_0_  ;
  output \g11448/_0_  ;
  output \g11558/_0_  ;
  output \g11559/_0_  ;
  output \g11824/_1_  ;
  output \g11853/_0_  ;
  output \g11854/_0_  ;
  output \g11977/_0_  ;
  output \g11981/_0_  ;
  output \g2584_pad  ;
  output \g4121_pad  ;
  output \g4809_pad  ;
  output \g5692_pad  ;
  output \g6282_pad  ;
  output \g6284_pad  ;
  output \g6360_pad  ;
  output \g6362_pad  ;
  output \g6364_pad  ;
  output \g6366_pad  ;
  output \g6368_pad  ;
  output \g6370_pad  ;
  output \g6372_pad  ;
  output \g6374_pad  ;
  wire n147 , n148 , n149 , n150 , n151 , n152 , n153 , n154 , n155 , n156 , n157 , n158 , n159 , n160 , n161 , n162 , n163 , n164 , n165 , n166 , n167 , n168 , n169 , n170 , n171 , n172 , n173 , n174 , n175 , n176 , n177 , n178 , n179 , n180 , n181 , n182 , n183 , n184 , n185 , n186 , n187 , n188 , n189 , n190 , n191 , n192 , n193 , n194 , n195 , n196 , n197 , n198 , n199 , n200 , n201 , n202 , n203 , n204 , n205 , n206 , n207 , n208 , n209 , n210 , n211 , n212 , n213 , n214 , n215 , n216 , n217 , n218 , n219 , n220 , n221 , n222 , n223 , n224 , n225 , n226 , n227 , n228 , n229 , n230 , n231 , n232 , n233 , n234 , n235 , n236 , n237 , n238 , n239 , n240 , n241 , n242 , n243 , n244 , n245 , n246 , n247 , n248 , n249 , n250 , n251 , n252 , n253 , n254 , n255 , n256 , n257 , n258 , n259 , n260 , n261 , n262 , n263 , n264 , n265 , n266 , n267 , n268 , n269 , n270 , n271 , n272 , n273 , n274 , n275 , n276 , n277 , n278 , n279 , n280 , n281 , n282 , n283 , n284 , n285 , n286 , n287 , n288 , n289 , n290 , n291 , n292 , n293 , n294 , n295 , n296 , n297 , n298 , n299 , n300 , n301 , n302 , n303 , n304 , n305 , n306 , n307 , n308 , n309 , n310 , n311 , n312 , n313 , n314 , n315 , n316 , n317 , n318 , n319 , n320 , n321 , n322 , n323 , n324 , n325 , n326 , n327 , n328 , n329 , n330 , n331 , n332 , n333 , n334 , n335 , n336 , n337 , n338 , n339 , n340 , n341 , n342 , n343 , n344 , n345 , n346 , n347 , n348 , n349 , n350 , n351 , n352 , n353 , n354 , n355 , n356 , n357 , n358 , n359 , n360 , n361 , n362 , n363 , n364 , n365 , n366 , n367 , n368 , n369 , n370 , n371 , n372 , n373 , n374 , n375 , n376 , n377 , n378 , n379 , n380 , n381 , n382 , n383 , n384 , n385 , n386 , n387 , n388 , n389 , n390 , n391 , n392 , n393 , n394 , n395 , n396 , n397 , n398 , n399 , n400 , n401 , n402 , n403 , n404 , n405 , n406 , n407 , n408 , n409 , n410 , n411 , n412 , n413 , n414 , n415 , n416 , n417 , n418 , n419 , n420 , n421 , n422 , n423 , n424 , n425 , n426 , n427 , n428 , n429 , n430 , n431 , n432 , n433 , n434 , n435 , n436 , n437 , n438 , n439 , n440 , n441 , n442 , n443 , n444 , n445 , n446 , n447 , n448 , n449 , n450 , n451 , n452 , n453 , n454 , n455 , n456 , n457 , n458 , n459 , n460 , n461 , n462 , n463 , n464 , n465 , n466 , n467 , n468 , n469 , n470 , n471 , n472 , n473 , n474 , n475 , n476 , n477 , n478 , n479 , n480 , n481 , n482 , n483 , n484 , n485 , n486 , n487 , n488 , n489 , n490 , n491 , n492 , n493 , n494 , n495 , n496 , n497 , n498 , n499 , n500 , n501 , n502 , n503 , n504 , n505 , n506 , n507 , n508 , n509 , n510 , n511 , n512 , n513 , n514 , n515 , n516 , n517 , n518 , n519 , n520 , n521 , n522 , n523 , n524 , n525 , n526 , n527 , n528 , n529 , n530 , n531 , n532 , n533 , n534 , n535 , n536 , n537 , n538 , n539 , n540 , n541 , n542 , n543 , n544 , n545 , n546 , n547 , n548 , n549 , n550 , n551 , n552 , n553 , n554 , n555 , n556 , n557 , n558 , n559 , n560 , n561 , n562 , n563 , n564 , n565 , n566 , n567 , n568 , n569 , n570 , n571 , n572 , n573 , n574 , n575 , n576 , n577 , n578 , n579 , n580 , n581 , n582 , n583 , n584 , n585 , n586 , n587 , n588 , n589 , n590 , n591 , n592 , n593 , n594 , n595 , n596 , n597 , n598 , n599 , n600 , n601 , n602 , n603 , n604 , n605 , n606 , n607 , n608 , n609 , n610 , n611 , n612 , n613 , n614 , n615 , n616 , n617 , n618 , n619 , n620 , n621 , n622 , n623 , n624 , n625 , n626 , n627 , n628 , n629 , n630 , n631 , n632 , n633 , n634 , n635 , n636 , n637 , n638 , n639 , n640 , n641 , n642 , n643 , n644 , n645 , n646 , n647 , n648 , n649 , n650 , n651 , n652 , n653 , n654 , n655 , n656 , n657 , n658 , n659 , n660 , n661 , n662 , n663 , n664 , n665 , n666 , n667 , n668 , n669 , n670 , n671 , n672 , n673 , n674 , n675 , n676 , n677 , n678 , n679 , n680 , n681 , n682 , n683 , n684 , n685 , n686 , n687 , n688 , n689 , n690 , n691 , n692 , n693 , n694 , n695 , n696 , n697 , n698 , n699 , n700 , n701 , n702 , n703 , n704 , n705 , n706 , n707 , n708 , n709 , n710 , n711 , n712 , n713 , n714 , n715 , n716 , n717 , n718 , n719 , n720 , n721 , n722 , n723 , n724 , n725 , n726 , n727 , n728 , n729 , n730 , n731 , n732 , n733 , n734 , n735 , n736 , n737 , n738 , n739 , n740 , n741 , n742 , n743 , n744 , n745 , n746 , n747 , n748 , n749 , n750 , n751 , n752 , n753 , n754 , n755 , n756 , n757 , n758 , n759 , n760 , n761 , n762 , n763 , n764 , n765 , n766 , n767 , n768 , n769 , n770 , n771 , n772 , n773 , n774 , n775 , n776 , n777 , n778 , n779 , n780 , n781 , n782 , n783 , n784 , n785 , n786 , n787 , n788 , n789 , n790 , n791 , n792 , n793 , n794 , n795 , n796 , n797 , n798 , n799 , n800 , n801 , n802 , n803 , n804 , n805 , n806 , n807 , n808 , n809 , n810 , n811 , n812 , n813 ;
  assign n147 = \g602_reg/NET0131  & \g610_reg/NET0131  ;
  assign n148 = \g613_reg/NET0131  & n147 ;
  assign n149 = \g616_reg/NET0131  & n148 ;
  assign n150 = \g619_reg/NET0131  & n149 ;
  assign n151 = \g622_reg/NET0131  & n150 ;
  assign n152 = \g625_reg/NET0131  & n151 ;
  assign n153 = \g628_reg/NET0131  & n152 ;
  assign n154 = \g631_reg/NET0131  & n153 ;
  assign n155 = \g578_reg/NET0131  & n154 ;
  assign n156 = \g582_reg/NET0131  & n155 ;
  assign n157 = \g586_reg/NET0131  & n156 ;
  assign n158 = \g574_reg/NET0131  & n157 ;
  assign n159 = ~\g590_reg/NET0131  & ~n158 ;
  assign n160 = \g590_reg/NET0131  & n158 ;
  assign n161 = ~n159 & ~n160 ;
  assign n162 = \g594_reg/NET0131  & n160 ;
  assign n163 = \g639_pad  & ~n162 ;
  assign n164 = ~n161 & n163 ;
  assign n165 = ~\g582_reg/NET0131  & ~n155 ;
  assign n166 = ~n156 & ~n165 ;
  assign n167 = n163 & n166 ;
  assign n168 = ~\g586_reg/NET0131  & ~n156 ;
  assign n169 = ~n157 & ~n168 ;
  assign n170 = n163 & n169 ;
  assign n171 = ~\g594_reg/NET0131  & ~n160 ;
  assign n172 = n163 & ~n171 ;
  assign n173 = ~\g574_reg/NET0131  & ~n157 ;
  assign n174 = ~n158 & ~n173 ;
  assign n175 = n163 & ~n174 ;
  assign n176 = ~\g578_reg/NET0131  & ~n154 ;
  assign n177 = ~n155 & ~n176 ;
  assign n178 = n163 & n177 ;
  assign n179 = \g19_reg/NET0131  & ~\g25_reg/NET0131  ;
  assign n180 = ~\g19_reg/NET0131  & \g25_reg/NET0131  ;
  assign n181 = ~n179 & ~n180 ;
  assign n182 = ~\g3_reg/NET0131  & ~\g7_reg/NET0131  ;
  assign n183 = \g3_reg/NET0131  & \g7_reg/NET0131  ;
  assign n184 = ~n182 & ~n183 ;
  assign n185 = \g33_reg/NET0131  & n184 ;
  assign n186 = ~\g33_reg/NET0131  & ~n184 ;
  assign n187 = ~n185 & ~n186 ;
  assign n188 = \g11_reg/NET0131  & ~\g15_reg/NET0131  ;
  assign n189 = ~\g11_reg/NET0131  & \g15_reg/NET0131  ;
  assign n190 = ~n188 & ~n189 ;
  assign n191 = \g29_reg/NET0131  & n190 ;
  assign n192 = ~\g29_reg/NET0131  & ~n190 ;
  assign n193 = ~n191 & ~n192 ;
  assign n194 = n187 & ~n193 ;
  assign n195 = ~n187 & n193 ;
  assign n196 = ~n194 & ~n195 ;
  assign n197 = n181 & n196 ;
  assign n198 = ~n181 & ~n196 ;
  assign n199 = ~n197 & ~n198 ;
  assign n200 = \g1293_pad  & \g702_pad  ;
  assign n201 = ~\g266_reg/NET0131  & \g4110_pad  ;
  assign n202 = \g662_reg/NET0131  & n201 ;
  assign n203 = n200 & n202 ;
  assign n204 = \g676_reg/NET0131  & n203 ;
  assign n205 = ~\g698_reg/NET0131  & n204 ;
  assign n206 = ~\g688_reg/NET0131  & ~\g689_reg/NET0131  ;
  assign n207 = n205 & n206 ;
  assign n208 = ~\g687_reg/NET0131  & n207 ;
  assign n209 = \g204_reg/NET0131  & \g205_reg/NET0131  ;
  assign n210 = \g206_reg/NET0131  & n209 ;
  assign n211 = \g207_reg/NET0131  & n210 ;
  assign n212 = \g208_reg/NET0131  & n211 ;
  assign n213 = \g209_reg/NET0131  & n212 ;
  assign n214 = \g208_reg/NET0131  & ~\g209_reg/NET0131  ;
  assign n215 = ~\g208_reg/NET0131  & \g209_reg/NET0131  ;
  assign n216 = ~n214 & ~n215 ;
  assign n217 = n211 & n215 ;
  assign n218 = ~n216 & ~n217 ;
  assign n219 = ~\g471_reg/NET0131  & ~n218 ;
  assign n220 = \g471_reg/NET0131  & ~n217 ;
  assign n221 = ~n219 & ~n220 ;
  assign n223 = \g204_reg/NET0131  & \g679_reg/NET0131  ;
  assign n222 = ~\g204_reg/NET0131  & \g680_reg/NET0131  ;
  assign n224 = ~\g205_reg/NET0131  & ~n222 ;
  assign n225 = ~n223 & n224 ;
  assign n227 = ~\g204_reg/NET0131  & \g678_reg/NET0131  ;
  assign n226 = \g204_reg/NET0131  & \g677_reg/NET0131  ;
  assign n228 = \g205_reg/NET0131  & ~n226 ;
  assign n229 = ~n227 & n228 ;
  assign n230 = ~n225 & ~n229 ;
  assign n231 = \g206_reg/NET0131  & ~n230 ;
  assign n233 = \g204_reg/NET0131  & \g683_reg/NET0131  ;
  assign n232 = ~\g204_reg/NET0131  & \g684_reg/NET0131  ;
  assign n234 = ~\g205_reg/NET0131  & ~n232 ;
  assign n235 = ~n233 & n234 ;
  assign n237 = ~\g204_reg/NET0131  & \g682_reg/NET0131  ;
  assign n236 = \g204_reg/NET0131  & \g681_reg/NET0131  ;
  assign n238 = \g205_reg/NET0131  & ~n236 ;
  assign n239 = ~n237 & n238 ;
  assign n240 = ~n235 & ~n239 ;
  assign n241 = ~\g206_reg/NET0131  & ~n240 ;
  assign n242 = ~n231 & ~n241 ;
  assign n244 = \g471_reg/NET0131  & n242 ;
  assign n243 = ~\g471_reg/NET0131  & ~n242 ;
  assign n245 = n216 & ~n243 ;
  assign n246 = ~n244 & n245 ;
  assign n247 = ~n221 & ~n246 ;
  assign n248 = \g210_reg/NET0131  & \g211_reg/NET0131  ;
  assign n249 = ~n247 & n248 ;
  assign n250 = n213 & n249 ;
  assign n253 = \g210_reg/NET0131  & ~\g211_reg/NET0131  ;
  assign n254 = n213 & n253 ;
  assign n255 = n246 & n254 ;
  assign n251 = ~\g210_reg/NET0131  & \g211_reg/NET0131  ;
  assign n252 = n213 & n251 ;
  assign n256 = ~\g210_reg/NET0131  & ~\g211_reg/NET0131  ;
  assign n257 = ~\g471_reg/NET0131  & n256 ;
  assign n258 = ~n218 & n257 ;
  assign n259 = ~n252 & ~n258 ;
  assign n260 = ~n255 & n259 ;
  assign n261 = ~n250 & n260 ;
  assign n262 = \g211_reg/NET0131  & n261 ;
  assign n263 = ~n246 & n254 ;
  assign n264 = ~n213 & n248 ;
  assign n265 = ~n247 & n264 ;
  assign n266 = ~n212 & n253 ;
  assign n267 = n246 & n266 ;
  assign n268 = ~n265 & ~n267 ;
  assign n269 = ~n263 & n268 ;
  assign n270 = ~n262 & n269 ;
  assign n271 = \g197_reg/NET0131  & ~n270 ;
  assign n272 = ~\g197_reg/NET0131  & \g684_reg/NET0131  ;
  assign n273 = ~n271 & ~n272 ;
  assign n274 = n208 & ~n273 ;
  assign n275 = \g687_reg/NET0131  & n207 ;
  assign n276 = \g276_reg/NET0131  & \g277_reg/NET0131  ;
  assign n277 = \g278_reg/NET0131  & n276 ;
  assign n278 = \g279_reg/NET0131  & n277 ;
  assign n279 = \g280_reg/NET0131  & n278 ;
  assign n280 = \g281_reg/NET0131  & n279 ;
  assign n281 = ~\g280_reg/NET0131  & \g281_reg/NET0131  ;
  assign n282 = \g280_reg/NET0131  & ~\g281_reg/NET0131  ;
  assign n283 = ~n281 & ~n282 ;
  assign n285 = \g276_reg/NET0131  & \g679_reg/NET0131  ;
  assign n284 = ~\g276_reg/NET0131  & \g680_reg/NET0131  ;
  assign n286 = ~\g277_reg/NET0131  & ~n284 ;
  assign n287 = ~n285 & n286 ;
  assign n289 = ~\g276_reg/NET0131  & \g678_reg/NET0131  ;
  assign n288 = \g276_reg/NET0131  & \g677_reg/NET0131  ;
  assign n290 = \g277_reg/NET0131  & ~n288 ;
  assign n291 = ~n289 & n290 ;
  assign n292 = ~n287 & ~n291 ;
  assign n293 = \g278_reg/NET0131  & ~n292 ;
  assign n295 = \g276_reg/NET0131  & \g683_reg/NET0131  ;
  assign n294 = ~\g276_reg/NET0131  & \g684_reg/NET0131  ;
  assign n296 = ~\g277_reg/NET0131  & ~n294 ;
  assign n297 = ~n295 & n296 ;
  assign n299 = \g276_reg/NET0131  & \g681_reg/NET0131  ;
  assign n298 = ~\g276_reg/NET0131  & \g682_reg/NET0131  ;
  assign n300 = \g277_reg/NET0131  & ~n298 ;
  assign n301 = ~n299 & n300 ;
  assign n302 = ~n297 & ~n301 ;
  assign n303 = ~\g278_reg/NET0131  & ~n302 ;
  assign n304 = ~n293 & ~n303 ;
  assign n305 = \g478_reg/NET0131  & ~n304 ;
  assign n306 = ~\g478_reg/NET0131  & n304 ;
  assign n307 = ~n305 & ~n306 ;
  assign n308 = n283 & n307 ;
  assign n309 = n278 & n281 ;
  assign n310 = ~n283 & ~n309 ;
  assign n311 = \g478_reg/NET0131  & ~n310 ;
  assign n312 = ~\g478_reg/NET0131  & n310 ;
  assign n313 = ~n311 & ~n312 ;
  assign n314 = ~n283 & n313 ;
  assign n315 = \g282_reg/NET0131  & \g283_reg/NET0131  ;
  assign n316 = ~n314 & n315 ;
  assign n317 = ~n308 & n316 ;
  assign n318 = \g282_reg/NET0131  & ~n317 ;
  assign n319 = n280 & ~n318 ;
  assign n320 = \g283_reg/NET0131  & ~n319 ;
  assign n321 = n283 & ~n307 ;
  assign n322 = \g282_reg/NET0131  & ~\g283_reg/NET0131  ;
  assign n323 = n321 & n322 ;
  assign n324 = ~n317 & ~n323 ;
  assign n325 = ~n280 & ~n324 ;
  assign n326 = n280 & n322 ;
  assign n327 = ~n321 & n326 ;
  assign n328 = ~n325 & ~n327 ;
  assign n329 = ~n320 & n328 ;
  assign n330 = \g269_reg/NET0131  & ~n329 ;
  assign n331 = ~\g269_reg/NET0131  & \g684_reg/NET0131  ;
  assign n332 = ~n330 & ~n331 ;
  assign n333 = n275 & ~n332 ;
  assign n335 = \g689_reg/NET0131  & \g698_reg/NET0131  ;
  assign n336 = ~\g688_reg/NET0131  & n335 ;
  assign n341 = \g685_reg/NET0131  & n336 ;
  assign n342 = ~\g682_reg/NET0131  & n341 ;
  assign n343 = \g683_reg/NET0131  & \g684_reg/NET0131  ;
  assign n344 = ~\g681_reg/NET0131  & n343 ;
  assign n345 = n342 & n344 ;
  assign n346 = n203 & n345 ;
  assign n347 = \g677_reg/NET0131  & n346 ;
  assign n348 = \g500_reg/NET0131  & n347 ;
  assign n350 = \g688_reg/NET0131  & n335 ;
  assign n351 = n203 & n350 ;
  assign n356 = ~\g680_reg/NET0131  & n351 ;
  assign n357 = ~\g679_reg/NET0131  & n356 ;
  assign n349 = ~\g678_reg/NET0131  & ~\g679_reg/NET0131  ;
  assign n352 = \g680_reg/NET0131  & n349 ;
  assign n353 = n351 & n352 ;
  assign n354 = \g684_reg/NET0131  & n341 ;
  assign n355 = n203 & n354 ;
  assign n360 = ~n353 & ~n355 ;
  assign n361 = ~n207 & n360 ;
  assign n362 = ~n357 & n361 ;
  assign n334 = \g689_reg/NET0131  & n205 ;
  assign n337 = ~\g685_reg/NET0131  & n336 ;
  assign n338 = n204 & n337 ;
  assign n339 = ~n334 & ~n338 ;
  assign n358 = \g678_reg/NET0131  & n356 ;
  assign n359 = \g679_reg/NET0131  & n358 ;
  assign n363 = n339 & ~n359 ;
  assign n364 = n362 & n363 ;
  assign n365 = ~n348 & ~n364 ;
  assign n373 = \g557_pad  & n359 ;
  assign n340 = \g684_reg/NET0131  & ~n339 ;
  assign n366 = n203 & n343 ;
  assign n367 = \g682_reg/NET0131  & n341 ;
  assign n368 = n366 & n367 ;
  assign n369 = ~\g677_reg/NET0131  & n368 ;
  assign n370 = \g434_reg/NET0131  & n369 ;
  assign n371 = \g677_reg/NET0131  & n368 ;
  assign n372 = \g430_reg/NET0131  & n371 ;
  assign n374 = ~n370 & ~n372 ;
  assign n375 = ~n340 & n374 ;
  assign n376 = ~n373 & n375 ;
  assign n377 = n365 & n376 ;
  assign n378 = ~n333 & n377 ;
  assign n379 = ~n274 & n378 ;
  assign n380 = ~\g197_reg/NET0131  & \g683_reg/NET0131  ;
  assign n381 = ~\g211_reg/NET0131  & n221 ;
  assign n382 = \g210_reg/NET0131  & ~n381 ;
  assign n383 = n268 & n382 ;
  assign n384 = n261 & ~n383 ;
  assign n385 = ~n263 & n384 ;
  assign n386 = \g197_reg/NET0131  & ~n385 ;
  assign n387 = ~n380 & ~n386 ;
  assign n388 = n208 & ~n387 ;
  assign n389 = ~\g283_reg/NET0131  & ~n283 ;
  assign n390 = ~n313 & n389 ;
  assign n391 = \g282_reg/NET0131  & ~n390 ;
  assign n392 = n324 & ~n391 ;
  assign n393 = ~n325 & ~n392 ;
  assign n394 = ~\g282_reg/NET0131  & ~\g283_reg/NET0131  ;
  assign n395 = ~\g478_reg/NET0131  & n394 ;
  assign n396 = ~n310 & n395 ;
  assign n397 = ~\g282_reg/NET0131  & \g283_reg/NET0131  ;
  assign n398 = n280 & n397 ;
  assign n399 = ~n396 & ~n398 ;
  assign n400 = ~n393 & n399 ;
  assign n401 = \g269_reg/NET0131  & ~n400 ;
  assign n402 = ~\g269_reg/NET0131  & \g683_reg/NET0131  ;
  assign n403 = ~n401 & ~n402 ;
  assign n404 = n275 & ~n403 ;
  assign n408 = \g558_pad  & n359 ;
  assign n405 = \g683_reg/NET0131  & ~n339 ;
  assign n406 = \g426_reg/NET0131  & n371 ;
  assign n407 = \g437_reg/NET0131  & n369 ;
  assign n409 = ~n406 & ~n407 ;
  assign n410 = ~n405 & n409 ;
  assign n411 = ~n408 & n410 ;
  assign n412 = n365 & n411 ;
  assign n413 = ~n404 & n412 ;
  assign n414 = ~n388 & n413 ;
  assign n415 = \g567_pad  & \g598_reg/NET0131  ;
  assign n416 = \g634_reg/NET0131  & n415 ;
  assign n417 = \g642_reg/NET0131  & n416 ;
  assign n418 = \g606_reg/NET0131  & n417 ;
  assign n419 = \g646_reg/NET0131  & n418 ;
  assign n420 = \g650_reg/NET0131  & n419 ;
  assign n421 = \g654_reg/NET0131  & n420 ;
  assign n423 = \g571_reg/NET0131  & n421 ;
  assign n422 = ~\g571_reg/NET0131  & ~n421 ;
  assign n424 = \g638_reg/NET0131  & ~n422 ;
  assign n425 = ~n423 & n424 ;
  assign n445 = ~\g197_reg/NET0131  & \g679_reg/NET0131  ;
  assign n446 = \g197_reg/NET0131  & ~n258 ;
  assign n447 = ~n213 & ~n257 ;
  assign n448 = ~n213 & ~n218 ;
  assign n449 = ~n447 & ~n448 ;
  assign n450 = n446 & ~n449 ;
  assign n451 = ~\g206_reg/NET0131  & ~n209 ;
  assign n452 = ~n210 & ~n451 ;
  assign n453 = n450 & n452 ;
  assign n454 = ~n445 & ~n453 ;
  assign n455 = n208 & ~n454 ;
  assign n426 = ~\g269_reg/NET0131  & \g679_reg/NET0131  ;
  assign n427 = ~n280 & ~n395 ;
  assign n428 = \g269_reg/NET0131  & n427 ;
  assign n429 = ~\g278_reg/NET0131  & ~n276 ;
  assign n430 = ~n277 & ~n429 ;
  assign n431 = n428 & n430 ;
  assign n432 = ~n426 & ~n431 ;
  assign n433 = n275 & ~n432 ;
  assign n434 = \g410_reg/NET0131  & n371 ;
  assign n435 = \g681_reg/NET0131  & n342 ;
  assign n436 = n366 & n435 ;
  assign n437 = \g551_reg/NET0131  & n436 ;
  assign n459 = ~n434 & ~n437 ;
  assign n438 = ~\g683_reg/NET0131  & n354 ;
  assign n439 = n203 & n438 ;
  assign n440 = \g293_reg/NET0131  & n439 ;
  assign n441 = \g453_reg/NET0131  & n369 ;
  assign n460 = ~n440 & ~n441 ;
  assign n461 = n459 & n460 ;
  assign n442 = ~\g677_reg/NET0131  & n346 ;
  assign n443 = \g536_reg/NET0131  & n442 ;
  assign n444 = \g508_reg/NET0131  & n347 ;
  assign n462 = ~n443 & ~n444 ;
  assign n463 = n461 & n462 ;
  assign n456 = \g562_pad  & n358 ;
  assign n457 = n339 & ~n456 ;
  assign n458 = \g679_reg/NET0131  & ~n457 ;
  assign n464 = ~n364 & ~n458 ;
  assign n465 = n463 & n464 ;
  assign n466 = ~n433 & n465 ;
  assign n467 = ~n455 & n466 ;
  assign n475 = ~\g269_reg/NET0131  & \g680_reg/NET0131  ;
  assign n476 = ~\g279_reg/NET0131  & ~n277 ;
  assign n477 = ~n278 & ~n476 ;
  assign n478 = n310 & n395 ;
  assign n479 = ~n280 & ~n478 ;
  assign n480 = ~n477 & n479 ;
  assign n481 = \g269_reg/NET0131  & ~n396 ;
  assign n482 = ~n480 & n481 ;
  assign n483 = ~n475 & ~n482 ;
  assign n484 = n275 & ~n483 ;
  assign n468 = ~\g197_reg/NET0131  & \g680_reg/NET0131  ;
  assign n469 = ~\g207_reg/NET0131  & ~n210 ;
  assign n470 = ~n211 & ~n469 ;
  assign n471 = ~n449 & ~n470 ;
  assign n472 = n446 & ~n471 ;
  assign n473 = ~n468 & ~n472 ;
  assign n474 = n208 & ~n473 ;
  assign n487 = \g512_reg/NET0131  & n347 ;
  assign n488 = \g680_reg/NET0131  & ~n339 ;
  assign n496 = ~n487 & ~n488 ;
  assign n489 = \g541_reg/NET0131  & n442 ;
  assign n492 = \g561_pad  & n359 ;
  assign n497 = ~n489 & ~n492 ;
  assign n498 = n496 & n497 ;
  assign n485 = \g414_reg/NET0131  & n371 ;
  assign n486 = \g449_reg/NET0131  & n369 ;
  assign n493 = ~n485 & ~n486 ;
  assign n490 = \g554_reg/NET0131  & n436 ;
  assign n491 = \g297_reg/NET0131  & n439 ;
  assign n494 = ~n490 & ~n491 ;
  assign n495 = n493 & n494 ;
  assign n499 = ~n364 & n495 ;
  assign n500 = n498 & n499 ;
  assign n501 = ~n474 & n500 ;
  assign n502 = ~n484 & n501 ;
  assign n511 = ~\g281_reg/NET0131  & ~n395 ;
  assign n512 = ~n279 & n511 ;
  assign n513 = n479 & ~n512 ;
  assign n514 = \g269_reg/NET0131  & ~n513 ;
  assign n515 = ~\g269_reg/NET0131  & ~\g682_reg/NET0131  ;
  assign n516 = ~n514 & ~n515 ;
  assign n517 = n275 & n516 ;
  assign n503 = ~\g197_reg/NET0131  & \g682_reg/NET0131  ;
  assign n504 = ~\g209_reg/NET0131  & ~n212 ;
  assign n505 = ~n213 & ~n504 ;
  assign n506 = ~n258 & ~n505 ;
  assign n507 = \g197_reg/NET0131  & ~n449 ;
  assign n508 = ~n506 & n507 ;
  assign n509 = ~n503 & ~n508 ;
  assign n510 = n208 & ~n509 ;
  assign n521 = \g559_pad  & n359 ;
  assign n518 = \g682_reg/NET0131  & ~n339 ;
  assign n519 = \g422_reg/NET0131  & n371 ;
  assign n520 = \g441_reg/NET0131  & n369 ;
  assign n522 = ~n519 & ~n520 ;
  assign n523 = ~n518 & n522 ;
  assign n524 = ~n521 & n523 ;
  assign n525 = ~n364 & n524 ;
  assign n526 = ~n510 & n525 ;
  assign n527 = ~n517 & n526 ;
  assign n544 = ~\g197_reg/NET0131  & \g678_reg/NET0131  ;
  assign n545 = ~\g204_reg/NET0131  & ~\g205_reg/NET0131  ;
  assign n546 = ~n209 & ~n545 ;
  assign n547 = n450 & n546 ;
  assign n548 = ~n544 & ~n547 ;
  assign n549 = n208 & ~n548 ;
  assign n550 = ~\g489_reg/NET0131  & n357 ;
  assign n551 = n339 & ~n550 ;
  assign n552 = \g678_reg/NET0131  & ~n551 ;
  assign n535 = \g457_reg/NET0131  & n369 ;
  assign n536 = \g406_reg/NET0131  & n371 ;
  assign n554 = ~n535 & ~n536 ;
  assign n541 = \g269_reg/NET0131  & n439 ;
  assign n542 = n349 & n356 ;
  assign n543 = \g492_reg/NET0131  & n542 ;
  assign n555 = ~n541 & ~n543 ;
  assign n556 = n554 & n555 ;
  assign n560 = ~n364 & n556 ;
  assign n561 = ~n552 & n560 ;
  assign n528 = ~\g269_reg/NET0131  & \g678_reg/NET0131  ;
  assign n529 = ~\g276_reg/NET0131  & ~\g277_reg/NET0131  ;
  assign n530 = ~n276 & ~n529 ;
  assign n531 = n428 & n530 ;
  assign n532 = ~n528 & ~n531 ;
  assign n533 = n275 & ~n532 ;
  assign n537 = \g465_reg/NET0131  & n442 ;
  assign n534 = \g548_reg/NET0131  & n436 ;
  assign n540 = \g672_reg/NET0131  & n353 ;
  assign n553 = ~n534 & ~n540 ;
  assign n557 = ~n537 & n553 ;
  assign n538 = \g563_pad  & n359 ;
  assign n539 = \g504_reg/NET0131  & n347 ;
  assign n558 = ~n538 & ~n539 ;
  assign n559 = n557 & n558 ;
  assign n562 = ~n533 & n559 ;
  assign n563 = n561 & n562 ;
  assign n564 = ~n549 & n563 ;
  assign n569 = ~\g197_reg/NET0131  & \g677_reg/NET0131  ;
  assign n570 = ~\g204_reg/NET0131  & n450 ;
  assign n571 = ~n569 & ~n570 ;
  assign n572 = n208 & ~n571 ;
  assign n582 = \g461_reg/NET0131  & n369 ;
  assign n579 = \g197_reg/NET0131  & n439 ;
  assign n580 = ~\g486_reg/NET0131  & ~\g679_reg/NET0131  ;
  assign n581 = n358 & n580 ;
  assign n585 = ~n579 & ~n581 ;
  assign n586 = ~n582 & n585 ;
  assign n573 = \g669_reg/NET0131  & n353 ;
  assign n574 = \g545_reg/NET0131  & n436 ;
  assign n583 = ~n573 & ~n574 ;
  assign n575 = \g402_reg/NET0131  & n371 ;
  assign n576 = \g496_reg/NET0131  & n542 ;
  assign n584 = ~n575 & ~n576 ;
  assign n587 = n583 & n584 ;
  assign n590 = n586 & n587 ;
  assign n591 = ~n364 & n590 ;
  assign n565 = ~\g269_reg/NET0131  & \g677_reg/NET0131  ;
  assign n566 = ~\g276_reg/NET0131  & n428 ;
  assign n567 = ~n565 & ~n566 ;
  assign n568 = n275 & ~n567 ;
  assign n578 = \g4422_pad  & n359 ;
  assign n577 = \g677_reg/NET0131  & ~n339 ;
  assign n588 = ~n348 & ~n577 ;
  assign n589 = ~n578 & n588 ;
  assign n592 = ~n568 & n589 ;
  assign n593 = n591 & n592 ;
  assign n594 = ~n572 & n593 ;
  assign n611 = \g681_reg/NET0131  & ~n339 ;
  assign n609 = \g560_pad  & n359 ;
  assign n610 = \g445_reg/NET0131  & n369 ;
  assign n612 = \g418_reg/NET0131  & n371 ;
  assign n613 = ~n610 & ~n612 ;
  assign n614 = ~n609 & n613 ;
  assign n615 = ~n611 & n614 ;
  assign n616 = ~n364 & n615 ;
  assign n595 = ~\g269_reg/NET0131  & \g681_reg/NET0131  ;
  assign n596 = ~\g280_reg/NET0131  & ~n278 ;
  assign n597 = ~n279 & ~n596 ;
  assign n598 = n427 & ~n597 ;
  assign n599 = \g269_reg/NET0131  & ~n598 ;
  assign n600 = ~n595 & ~n599 ;
  assign n601 = n275 & ~n600 ;
  assign n602 = ~\g197_reg/NET0131  & \g681_reg/NET0131  ;
  assign n603 = ~\g208_reg/NET0131  & ~n211 ;
  assign n604 = ~n212 & ~n603 ;
  assign n605 = n447 & ~n604 ;
  assign n606 = \g197_reg/NET0131  & ~n605 ;
  assign n607 = ~n602 & ~n606 ;
  assign n608 = n208 & ~n607 ;
  assign n617 = ~n601 & ~n608 ;
  assign n618 = n616 & n617 ;
  assign n619 = ~\g631_reg/NET0131  & ~n153 ;
  assign n620 = \g639_pad  & ~n154 ;
  assign n621 = ~n619 & n620 ;
  assign n622 = ~\g654_reg/NET0131  & ~n420 ;
  assign n623 = \g638_reg/NET0131  & ~n421 ;
  assign n624 = ~n622 & n623 ;
  assign n625 = ~\g628_reg/NET0131  & ~n152 ;
  assign n626 = \g639_pad  & ~n153 ;
  assign n627 = ~n625 & n626 ;
  assign n628 = ~n270 & ~n384 ;
  assign n629 = ~n329 & ~n400 ;
  assign n630 = ~\g650_reg/NET0131  & ~n419 ;
  assign n631 = \g638_reg/NET0131  & ~n420 ;
  assign n632 = ~n630 & n631 ;
  assign n633 = \g18_reg/NET0131  & ~\g28_reg/NET0131  ;
  assign n634 = ~\g18_reg/NET0131  & \g28_reg/NET0131  ;
  assign n635 = ~n633 & ~n634 ;
  assign n636 = ~\g10_reg/NET0131  & ~\g1_reg/NET0131  ;
  assign n637 = \g10_reg/NET0131  & \g1_reg/NET0131  ;
  assign n638 = ~n636 & ~n637 ;
  assign n639 = n635 & ~n638 ;
  assign n640 = ~n635 & n638 ;
  assign n641 = ~n639 & ~n640 ;
  assign n642 = ~\g14_reg/NET0131  & ~\g48_reg/NET0131  ;
  assign n643 = \g14_reg/NET0131  & \g48_reg/NET0131  ;
  assign n644 = ~n642 & ~n643 ;
  assign n645 = \g2_reg/NET0131  & n644 ;
  assign n646 = ~\g2_reg/NET0131  & ~n644 ;
  assign n647 = ~n645 & ~n646 ;
  assign n648 = \g24_reg/NET0131  & ~\g6_reg/NET0131  ;
  assign n649 = ~\g24_reg/NET0131  & \g6_reg/NET0131  ;
  assign n650 = ~n648 & ~n649 ;
  assign n651 = n647 & ~n650 ;
  assign n652 = ~n647 & n650 ;
  assign n653 = ~n651 & ~n652 ;
  assign n654 = n641 & n653 ;
  assign n655 = ~n641 & ~n653 ;
  assign n656 = ~n654 & ~n655 ;
  assign n657 = ~\g4110_pad  & ~n656 ;
  assign n658 = \g676_reg/NET0131  & ~n657 ;
  assign n659 = ~\g4110_pad  & n200 ;
  assign n660 = n658 & n659 ;
  assign n661 = n345 & n660 ;
  assign n662 = ~\g677_reg/NET0131  & n661 ;
  assign n663 = \g679_reg/NET0131  & n662 ;
  assign n687 = \g465_reg/NET0131  & ~n309 ;
  assign n673 = ~\g212_reg/NET0131  & ~\g248_reg/NET0131  ;
  assign n674 = ~\g254_reg/NET0131  & ~\g500_reg/NET0131  ;
  assign n675 = n673 & n674 ;
  assign n676 = \g212_reg/NET0131  & \g248_reg/NET0131  ;
  assign n677 = \g254_reg/NET0131  & \g500_reg/NET0131  ;
  assign n678 = n676 & n677 ;
  assign n679 = ~n675 & ~n678 ;
  assign n664 = ~\g218_reg/NET0131  & ~\g504_reg/NET0131  ;
  assign n665 = \g218_reg/NET0131  & \g504_reg/NET0131  ;
  assign n666 = ~n664 & ~n665 ;
  assign n680 = ~\g236_reg/NET0131  & ~\g242_reg/NET0131  ;
  assign n681 = ~\g260_reg/NET0131  & n680 ;
  assign n682 = ~n666 & n681 ;
  assign n667 = ~\g230_reg/NET0131  & ~\g512_reg/NET0131  ;
  assign n668 = \g230_reg/NET0131  & \g512_reg/NET0131  ;
  assign n669 = ~n667 & ~n668 ;
  assign n670 = ~\g224_reg/NET0131  & ~\g508_reg/NET0131  ;
  assign n671 = \g224_reg/NET0131  & \g508_reg/NET0131  ;
  assign n672 = ~n670 & ~n671 ;
  assign n683 = ~n669 & ~n672 ;
  assign n684 = n682 & n683 ;
  assign n685 = ~n679 & n684 ;
  assign n686 = ~\g465_reg/NET0131  & ~n217 ;
  assign n688 = n685 & ~n686 ;
  assign n689 = ~n687 & n688 ;
  assign n690 = \g536_reg/NET0131  & ~n689 ;
  assign n691 = ~n662 & n690 ;
  assign n692 = ~n663 & ~n691 ;
  assign n693 = ~\g625_reg/NET0131  & ~n151 ;
  assign n694 = \g639_pad  & ~n152 ;
  assign n695 = ~n693 & n694 ;
  assign n696 = ~\g646_reg/NET0131  & ~n418 ;
  assign n697 = \g638_reg/NET0131  & ~n419 ;
  assign n698 = ~n696 & n697 ;
  assign n699 = ~\g492_reg/NET0131  & ~n317 ;
  assign n700 = ~\g496_reg/NET0131  & ~n249 ;
  assign n701 = \g677_reg/NET0131  & n661 ;
  assign n702 = ~\g622_reg/NET0131  & ~n150 ;
  assign n703 = \g639_pad  & ~n151 ;
  assign n704 = ~n702 & n703 ;
  assign n705 = n438 & n660 ;
  assign n706 = ~\g606_reg/NET0131  & ~n417 ;
  assign n707 = \g638_reg/NET0131  & ~n418 ;
  assign n708 = ~n706 & n707 ;
  assign n709 = \g4101_pad  & ~\g4105_pad  ;
  assign n710 = ~\g4101_pad  & \g4105_pad  ;
  assign n711 = ~n709 & ~n710 ;
  assign n712 = \g4103_pad  & n711 ;
  assign n713 = ~\g4103_pad  & ~n711 ;
  assign n714 = ~n712 & ~n713 ;
  assign n715 = \g4099_pad  & ~n714 ;
  assign n716 = ~\g4099_pad  & n714 ;
  assign n717 = ~n715 & ~n716 ;
  assign n718 = ~\g4100_pad  & ~\g4102_pad  ;
  assign n719 = \g4100_pad  & \g4102_pad  ;
  assign n720 = ~n718 & ~n719 ;
  assign n721 = ~n656 & n720 ;
  assign n722 = n656 & ~n720 ;
  assign n723 = ~n721 & ~n722 ;
  assign n724 = n717 & n723 ;
  assign n725 = ~n717 & ~n723 ;
  assign n726 = ~n724 & ~n725 ;
  assign n727 = ~\g4104_pad  & n726 ;
  assign n728 = ~\g669_reg/NET0131  & ~n727 ;
  assign n729 = ~\g619_reg/NET0131  & ~n149 ;
  assign n730 = \g639_pad  & ~n150 ;
  assign n731 = ~n729 & n730 ;
  assign n732 = ~\g642_reg/NET0131  & ~n416 ;
  assign n733 = \g638_reg/NET0131  & ~n417 ;
  assign n734 = ~n732 & n733 ;
  assign n735 = ~\g4104_pad  & n657 ;
  assign n736 = ~\g672_reg/NET0131  & ~n735 ;
  assign n737 = ~\g536_reg/NET0131  & n685 ;
  assign n738 = ~\g541_reg/NET0131  & n737 ;
  assign n742 = \g578_reg/NET0131  & \g681_reg/NET0131  ;
  assign n741 = ~\g578_reg/NET0131  & \g682_reg/NET0131  ;
  assign n743 = \g582_reg/NET0131  & ~n741 ;
  assign n744 = ~n742 & n743 ;
  assign n746 = \g578_reg/NET0131  & \g683_reg/NET0131  ;
  assign n745 = ~\g578_reg/NET0131  & \g684_reg/NET0131  ;
  assign n747 = ~\g582_reg/NET0131  & ~n745 ;
  assign n748 = ~n746 & n747 ;
  assign n749 = ~n744 & ~n748 ;
  assign n750 = ~\g586_reg/NET0131  & ~n749 ;
  assign n752 = \g578_reg/NET0131  & \g679_reg/NET0131  ;
  assign n751 = ~\g578_reg/NET0131  & \g680_reg/NET0131  ;
  assign n753 = ~\g582_reg/NET0131  & ~n751 ;
  assign n754 = ~n752 & n753 ;
  assign n756 = \g578_reg/NET0131  & \g677_reg/NET0131  ;
  assign n755 = ~\g578_reg/NET0131  & \g678_reg/NET0131  ;
  assign n757 = \g582_reg/NET0131  & ~n755 ;
  assign n758 = ~n756 & n757 ;
  assign n759 = ~n754 & ~n758 ;
  assign n760 = \g586_reg/NET0131  & ~n759 ;
  assign n761 = ~n750 & ~n760 ;
  assign n739 = ~\g590_reg/NET0131  & \g594_reg/NET0131  ;
  assign n740 = \g590_reg/NET0131  & ~\g594_reg/NET0131  ;
  assign n762 = ~n739 & ~n740 ;
  assign n763 = ~n761 & n762 ;
  assign n764 = \g574_reg/NET0131  & \g578_reg/NET0131  ;
  assign n765 = \g582_reg/NET0131  & \g586_reg/NET0131  ;
  assign n766 = n764 & n765 ;
  assign n767 = n739 & n766 ;
  assign n768 = ~n763 & ~n767 ;
  assign n769 = ~\g616_reg/NET0131  & ~n148 ;
  assign n770 = \g639_pad  & ~n149 ;
  assign n771 = ~n769 & n770 ;
  assign n772 = ~\g634_reg/NET0131  & ~n415 ;
  assign n773 = \g638_reg/NET0131  & ~n416 ;
  assign n774 = ~n772 & n773 ;
  assign n775 = ~\g613_reg/NET0131  & ~n147 ;
  assign n776 = ~n148 & ~n775 ;
  assign n777 = \g639_pad  & ~n776 ;
  assign n778 = \g465_reg/NET0131  & \g478_reg/NET0131  ;
  assign n779 = ~\g465_reg/NET0131  & \g471_reg/NET0131  ;
  assign n780 = ~n778 & ~n779 ;
  assign n781 = ~\g567_pad  & ~\g598_reg/NET0131  ;
  assign n782 = \g638_reg/NET0131  & ~n415 ;
  assign n783 = ~n781 & n782 ;
  assign n784 = ~\g602_reg/NET0131  & ~\g610_reg/NET0131  ;
  assign n785 = \g639_pad  & ~n147 ;
  assign n786 = ~n784 & n785 ;
  assign n787 = ~\g266_reg/NET0131  & \g4108_pad  ;
  assign n788 = ~\g602_reg/NET0131  & \g639_pad  ;
  assign n789 = ~\g680_reg/NET0131  & n662 ;
  assign n791 = \g465_reg/NET0131  & ~n280 ;
  assign n790 = ~\g465_reg/NET0131  & ~n213 ;
  assign n792 = n737 & ~n790 ;
  assign n793 = ~n791 & n792 ;
  assign n794 = ~\g541_reg/NET0131  & ~n793 ;
  assign n795 = ~n662 & n794 ;
  assign n796 = ~n789 & ~n795 ;
  assign n797 = ~\g102_pad  & \g89_pad  ;
  assign n798 = \g567_pad  & \g638_reg/NET0131  ;
  assign n799 = ~\g489_reg/NET0131  & \g492_reg/NET0131  ;
  assign n800 = ~\g486_reg/NET0131  & \g496_reg/NET0131  ;
  assign n801 = ~n799 & ~n800 ;
  assign n802 = ~\g4104_pad  & \g675_reg/NET0131  ;
  assign n803 = n658 & n802 ;
  assign n804 = \g4110_pad  & n803 ;
  assign n805 = ~n199 & n804 ;
  assign n806 = ~\g25_reg/NET0131  & n804 ;
  assign n807 = ~\g29_reg/NET0131  & n804 ;
  assign n808 = ~\g3_reg/NET0131  & n804 ;
  assign n809 = ~\g33_reg/NET0131  & n804 ;
  assign n810 = ~\g7_reg/NET0131  & n804 ;
  assign n811 = ~\g11_reg/NET0131  & n804 ;
  assign n812 = ~\g15_reg/NET0131  & n804 ;
  assign n813 = ~\g19_reg/NET0131  & n804 ;
  assign \_al_n1  = ~1'b0 ;
  assign \g10560/_0_  = ~n164 ;
  assign \g10562/_1_  = n167 ;
  assign \g10564/_1_  = n170 ;
  assign \g10566/_1_  = n172 ;
  assign \g10567/_0_  = ~n175 ;
  assign \g10569/_1_  = n178 ;
  assign \g10580/_0_  = n199 ;
  assign \g10616/_2_  = ~n379 ;
  assign \g10627/_2_  = ~n414 ;
  assign \g10628/_0_  = n425 ;
  assign \g10629/_2_  = ~n467 ;
  assign \g10630/_2_  = ~n502 ;
  assign \g10633/_2_  = ~n527 ;
  assign \g10635/_2_  = ~n564 ;
  assign \g10636/_2_  = ~n594 ;
  assign \g10637/_2_  = ~n618 ;
  assign \g10641/_0_  = n621 ;
  assign \g10649/_0_  = n624 ;
  assign \g10672/_0_  = ~n332 ;
  assign \g10673/_0_  = ~n273 ;
  assign \g10680/_0_  = n627 ;
  assign \g10683/_0_  = ~n628 ;
  assign \g10686/_0_  = ~n629 ;
  assign \g10695/_0_  = ~n403 ;
  assign \g10700/_0_  = n632 ;
  assign \g10703/_0_  = ~n270 ;
  assign \g10704/_0_  = ~n692 ;
  assign \g10748/_0_  = n695 ;
  assign \g10750/_2_  = ~n384 ;
  assign \g10757/_0_  = n516 ;
  assign \g10758/_0_  = ~n509 ;
  assign \g10782/_0_  = n698 ;
  assign \g10826/_0_  = ~n699 ;
  assign \g10827/_0_  = ~n700 ;
  assign \g10828/_1_  = n701 ;
  assign \g10832/_2_  = ~n607 ;
  assign \g10834/_2_  = ~n600 ;
  assign \g10836/_0_  = n704 ;
  assign \g10837/_1__syn_2  = n705 ;
  assign \g10868/_0_  = n708 ;
  assign \g10904/_0_  = ~n728 ;
  assign \g10913/_0_  = ~n483 ;
  assign \g10915/_0_  = ~n473 ;
  assign \g10922/_0_  = n731 ;
  assign \g10938/_0_  = ~n567 ;
  assign \g10939/_0_  = ~n532 ;
  assign \g10940/_0_  = ~n571 ;
  assign \g10941/_0_  = ~n548 ;
  assign \g10942/_0_  = ~n432 ;
  assign \g10944/_2_  = ~n454 ;
  assign \g10977/_0_  = n734 ;
  assign \g10980/_0_  = ~n736 ;
  assign \g11020/_0_  = ~n726 ;
  assign \g11028/_0_  = n738 ;
  assign \g11051/_0_  = n768 ;
  assign \g11057/_0_  = n771 ;
  assign \g11109/_0_  = n774 ;
  assign \g11113/_2_  = n685 ;
  assign \g11156/_0_  = ~n777 ;
  assign \g11172/_3_  = ~n780 ;
  assign \g11193/_0_  = n783 ;
  assign \g11219/_0_  = n786 ;
  assign \g11355/_0_  = ~\g678_reg/NET0131  ;
  assign \g11384/_0_  = ~\g677_reg/NET0131  ;
  assign \g11442/_0_  = n787 ;
  assign \g11448/_0_  = n788 ;
  assign \g11558/_0_  = ~\g266_reg/NET0131  ;
  assign \g11559/_0_  = ~\g4112_pad  ;
  assign \g11824/_1_  = ~n387 ;
  assign \g11853/_0_  = n796 ;
  assign \g11854/_0_  = n662 ;
  assign \g11977/_0_  = ~n329 ;
  assign \g11981/_0_  = ~n400 ;
  assign \g2584_pad  = n797 ;
  assign \g4121_pad  = ~n798 ;
  assign \g4809_pad  = n801 ;
  assign \g5692_pad  = 1'b0 ;
  assign \g6282_pad  = ~n803 ;
  assign \g6284_pad  = ~n805 ;
  assign \g6360_pad  = ~n806 ;
  assign \g6362_pad  = ~n807 ;
  assign \g6364_pad  = ~n808 ;
  assign \g6366_pad  = ~n809 ;
  assign \g6368_pad  = ~n810 ;
  assign \g6370_pad  = ~n811 ;
  assign \g6372_pad  = ~n812 ;
  assign \g6374_pad  = ~n813 ;
endmodule
