module top( \P1_P1_ADS_n_reg/NET0131  , \P1_P1_Address_reg[0]/NET0131  , \P1_P1_Address_reg[10]/NET0131  , \P1_P1_Address_reg[11]/NET0131  , \P1_P1_Address_reg[12]/NET0131  , \P1_P1_Address_reg[13]/NET0131  , \P1_P1_Address_reg[14]/NET0131  , \P1_P1_Address_reg[15]/NET0131  , \P1_P1_Address_reg[16]/NET0131  , \P1_P1_Address_reg[17]/NET0131  , \P1_P1_Address_reg[18]/NET0131  , \P1_P1_Address_reg[19]/NET0131  , \P1_P1_Address_reg[1]/NET0131  , \P1_P1_Address_reg[20]/NET0131  , \P1_P1_Address_reg[21]/NET0131  , \P1_P1_Address_reg[22]/NET0131  , \P1_P1_Address_reg[23]/NET0131  , \P1_P1_Address_reg[24]/NET0131  , \P1_P1_Address_reg[25]/NET0131  , \P1_P1_Address_reg[26]/NET0131  , \P1_P1_Address_reg[27]/NET0131  , \P1_P1_Address_reg[28]/NET0131  , \P1_P1_Address_reg[29]/NET0131  , \P1_P1_Address_reg[2]/NET0131  , \P1_P1_Address_reg[3]/NET0131  , \P1_P1_Address_reg[4]/NET0131  , \P1_P1_Address_reg[5]/NET0131  , \P1_P1_Address_reg[6]/NET0131  , \P1_P1_Address_reg[7]/NET0131  , \P1_P1_Address_reg[8]/NET0131  , \P1_P1_Address_reg[9]/NET0131  , \P1_P1_BE_n_reg[0]/NET0131  , \P1_P1_BE_n_reg[1]/NET0131  , \P1_P1_BE_n_reg[2]/NET0131  , \P1_P1_BE_n_reg[3]/NET0131  , \P1_P1_ByteEnable_reg[0]/NET0131  , \P1_P1_ByteEnable_reg[1]/NET0131  , \P1_P1_ByteEnable_reg[2]/NET0131  , \P1_P1_ByteEnable_reg[3]/NET0131  , \P1_P1_CodeFetch_reg/NET0131  , \P1_P1_D_C_n_reg/NET0131  , \P1_P1_DataWidth_reg[0]/NET0131  , \P1_P1_DataWidth_reg[1]/NET0131  , \P1_P1_Datao_reg[0]/NET0131  , \P1_P1_Datao_reg[10]/NET0131  , \P1_P1_Datao_reg[11]/NET0131  , \P1_P1_Datao_reg[12]/NET0131  , \P1_P1_Datao_reg[13]/NET0131  , \P1_P1_Datao_reg[14]/NET0131  , \P1_P1_Datao_reg[15]/NET0131  , \P1_P1_Datao_reg[16]/NET0131  , \P1_P1_Datao_reg[17]/NET0131  , \P1_P1_Datao_reg[18]/NET0131  , \P1_P1_Datao_reg[19]/NET0131  , \P1_P1_Datao_reg[1]/NET0131  , \P1_P1_Datao_reg[20]/NET0131  , \P1_P1_Datao_reg[21]/NET0131  , \P1_P1_Datao_reg[22]/NET0131  , \P1_P1_Datao_reg[23]/NET0131  , \P1_P1_Datao_reg[24]/NET0131  , \P1_P1_Datao_reg[25]/NET0131  , \P1_P1_Datao_reg[26]/NET0131  , \P1_P1_Datao_reg[27]/NET0131  , \P1_P1_Datao_reg[28]/NET0131  , \P1_P1_Datao_reg[29]/NET0131  , \P1_P1_Datao_reg[2]/NET0131  , \P1_P1_Datao_reg[30]/NET0131  , \P1_P1_Datao_reg[3]/NET0131  , \P1_P1_Datao_reg[4]/NET0131  , \P1_P1_Datao_reg[5]/NET0131  , \P1_P1_Datao_reg[6]/NET0131  , \P1_P1_Datao_reg[7]/NET0131  , \P1_P1_Datao_reg[8]/NET0131  , \P1_P1_Datao_reg[9]/NET0131  , \P1_P1_EAX_reg[0]/NET0131  , \P1_P1_EAX_reg[10]/NET0131  , \P1_P1_EAX_reg[11]/NET0131  , \P1_P1_EAX_reg[12]/NET0131  , \P1_P1_EAX_reg[13]/NET0131  , \P1_P1_EAX_reg[14]/NET0131  , \P1_P1_EAX_reg[15]/NET0131  , \P1_P1_EAX_reg[16]/NET0131  , \P1_P1_EAX_reg[17]/NET0131  , \P1_P1_EAX_reg[18]/NET0131  , \P1_P1_EAX_reg[19]/NET0131  , \P1_P1_EAX_reg[1]/NET0131  , \P1_P1_EAX_reg[20]/NET0131  , \P1_P1_EAX_reg[21]/NET0131  , \P1_P1_EAX_reg[22]/NET0131  , \P1_P1_EAX_reg[23]/NET0131  , \P1_P1_EAX_reg[24]/NET0131  , \P1_P1_EAX_reg[25]/NET0131  , \P1_P1_EAX_reg[26]/NET0131  , \P1_P1_EAX_reg[27]/NET0131  , \P1_P1_EAX_reg[28]/NET0131  , \P1_P1_EAX_reg[29]/NET0131  , \P1_P1_EAX_reg[2]/NET0131  , \P1_P1_EAX_reg[30]/NET0131  , \P1_P1_EAX_reg[31]/NET0131  , \P1_P1_EAX_reg[3]/NET0131  , \P1_P1_EAX_reg[4]/NET0131  , \P1_P1_EAX_reg[5]/NET0131  , \P1_P1_EAX_reg[6]/NET0131  , \P1_P1_EAX_reg[7]/NET0131  , \P1_P1_EAX_reg[8]/NET0131  , \P1_P1_EAX_reg[9]/NET0131  , \P1_P1_EBX_reg[0]/NET0131  , \P1_P1_EBX_reg[10]/NET0131  , \P1_P1_EBX_reg[11]/NET0131  , \P1_P1_EBX_reg[12]/NET0131  , \P1_P1_EBX_reg[13]/NET0131  , \P1_P1_EBX_reg[14]/NET0131  , \P1_P1_EBX_reg[15]/NET0131  , \P1_P1_EBX_reg[16]/NET0131  , \P1_P1_EBX_reg[17]/NET0131  , \P1_P1_EBX_reg[18]/NET0131  , \P1_P1_EBX_reg[19]/NET0131  , \P1_P1_EBX_reg[1]/NET0131  , \P1_P1_EBX_reg[20]/NET0131  , \P1_P1_EBX_reg[21]/NET0131  , \P1_P1_EBX_reg[22]/NET0131  , \P1_P1_EBX_reg[23]/NET0131  , \P1_P1_EBX_reg[24]/NET0131  , \P1_P1_EBX_reg[25]/NET0131  , \P1_P1_EBX_reg[26]/NET0131  , \P1_P1_EBX_reg[27]/NET0131  , \P1_P1_EBX_reg[28]/NET0131  , \P1_P1_EBX_reg[29]/NET0131  , \P1_P1_EBX_reg[2]/NET0131  , \P1_P1_EBX_reg[30]/NET0131  , \P1_P1_EBX_reg[31]/NET0131  , \P1_P1_EBX_reg[3]/NET0131  , \P1_P1_EBX_reg[4]/NET0131  , \P1_P1_EBX_reg[5]/NET0131  , \P1_P1_EBX_reg[6]/NET0131  , \P1_P1_EBX_reg[7]/NET0131  , \P1_P1_EBX_reg[8]/NET0131  , \P1_P1_EBX_reg[9]/NET0131  , \P1_P1_Flush_reg/NET0131  , \P1_P1_InstAddrPointer_reg[0]/NET0131  , \P1_P1_InstAddrPointer_reg[10]/NET0131  , \P1_P1_InstAddrPointer_reg[11]/NET0131  , \P1_P1_InstAddrPointer_reg[12]/NET0131  , \P1_P1_InstAddrPointer_reg[13]/NET0131  , \P1_P1_InstAddrPointer_reg[14]/NET0131  , \P1_P1_InstAddrPointer_reg[15]/NET0131  , \P1_P1_InstAddrPointer_reg[16]/NET0131  , \P1_P1_InstAddrPointer_reg[17]/NET0131  , \P1_P1_InstAddrPointer_reg[18]/NET0131  , \P1_P1_InstAddrPointer_reg[19]/NET0131  , \P1_P1_InstAddrPointer_reg[1]/NET0131  , \P1_P1_InstAddrPointer_reg[20]/NET0131  , \P1_P1_InstAddrPointer_reg[21]/NET0131  , \P1_P1_InstAddrPointer_reg[22]/NET0131  , \P1_P1_InstAddrPointer_reg[23]/NET0131  , \P1_P1_InstAddrPointer_reg[24]/NET0131  , \P1_P1_InstAddrPointer_reg[25]/NET0131  , \P1_P1_InstAddrPointer_reg[26]/NET0131  , \P1_P1_InstAddrPointer_reg[27]/NET0131  , \P1_P1_InstAddrPointer_reg[28]/NET0131  , \P1_P1_InstAddrPointer_reg[29]/NET0131  , \P1_P1_InstAddrPointer_reg[2]/NET0131  , \P1_P1_InstAddrPointer_reg[30]/NET0131  , \P1_P1_InstAddrPointer_reg[31]/NET0131  , \P1_P1_InstAddrPointer_reg[3]/NET0131  , \P1_P1_InstAddrPointer_reg[4]/NET0131  , \P1_P1_InstAddrPointer_reg[5]/NET0131  , \P1_P1_InstAddrPointer_reg[6]/NET0131  , \P1_P1_InstAddrPointer_reg[7]/NET0131  , \P1_P1_InstAddrPointer_reg[8]/NET0131  , \P1_P1_InstAddrPointer_reg[9]/NET0131  , \P1_P1_InstQueueRd_Addr_reg[0]/NET0131  , \P1_P1_InstQueueRd_Addr_reg[1]/NET0131  , \P1_P1_InstQueueRd_Addr_reg[2]/NET0131  , \P1_P1_InstQueueRd_Addr_reg[3]/NET0131  , \P1_P1_InstQueueWr_Addr_reg[0]/NET0131  , \P1_P1_InstQueueWr_Addr_reg[1]/NET0131  , \P1_P1_InstQueueWr_Addr_reg[2]/NET0131  , \P1_P1_InstQueueWr_Addr_reg[3]/NET0131  , \P1_P1_InstQueue_reg[0][0]/NET0131  , \P1_P1_InstQueue_reg[0][1]/NET0131  , \P1_P1_InstQueue_reg[0][2]/NET0131  , \P1_P1_InstQueue_reg[0][3]/NET0131  , \P1_P1_InstQueue_reg[0][4]/NET0131  , \P1_P1_InstQueue_reg[0][5]/NET0131  , \P1_P1_InstQueue_reg[0][6]/NET0131  , \P1_P1_InstQueue_reg[0][7]/NET0131  , \P1_P1_InstQueue_reg[10][0]/NET0131  , \P1_P1_InstQueue_reg[10][1]/NET0131  , \P1_P1_InstQueue_reg[10][2]/NET0131  , \P1_P1_InstQueue_reg[10][3]/NET0131  , \P1_P1_InstQueue_reg[10][4]/NET0131  , \P1_P1_InstQueue_reg[10][5]/NET0131  , \P1_P1_InstQueue_reg[10][6]/NET0131  , \P1_P1_InstQueue_reg[10][7]/NET0131  , \P1_P1_InstQueue_reg[11][0]/NET0131  , \P1_P1_InstQueue_reg[11][1]/NET0131  , \P1_P1_InstQueue_reg[11][2]/NET0131  , \P1_P1_InstQueue_reg[11][3]/NET0131  , \P1_P1_InstQueue_reg[11][4]/NET0131  , \P1_P1_InstQueue_reg[11][5]/NET0131  , \P1_P1_InstQueue_reg[11][6]/NET0131  , \P1_P1_InstQueue_reg[11][7]/NET0131  , \P1_P1_InstQueue_reg[12][0]/NET0131  , \P1_P1_InstQueue_reg[12][1]/NET0131  , \P1_P1_InstQueue_reg[12][2]/NET0131  , \P1_P1_InstQueue_reg[12][3]/NET0131  , \P1_P1_InstQueue_reg[12][4]/NET0131  , \P1_P1_InstQueue_reg[12][5]/NET0131  , \P1_P1_InstQueue_reg[12][6]/NET0131  , \P1_P1_InstQueue_reg[12][7]/NET0131  , \P1_P1_InstQueue_reg[13][0]/NET0131  , \P1_P1_InstQueue_reg[13][1]/NET0131  , \P1_P1_InstQueue_reg[13][2]/NET0131  , \P1_P1_InstQueue_reg[13][3]/NET0131  , \P1_P1_InstQueue_reg[13][4]/NET0131  , \P1_P1_InstQueue_reg[13][5]/NET0131  , \P1_P1_InstQueue_reg[13][6]/NET0131  , \P1_P1_InstQueue_reg[13][7]/NET0131  , \P1_P1_InstQueue_reg[14][0]/NET0131  , \P1_P1_InstQueue_reg[14][1]/NET0131  , \P1_P1_InstQueue_reg[14][2]/NET0131  , \P1_P1_InstQueue_reg[14][3]/NET0131  , \P1_P1_InstQueue_reg[14][4]/NET0131  , \P1_P1_InstQueue_reg[14][5]/NET0131  , \P1_P1_InstQueue_reg[14][6]/NET0131  , \P1_P1_InstQueue_reg[14][7]/NET0131  , \P1_P1_InstQueue_reg[15][0]/NET0131  , \P1_P1_InstQueue_reg[15][1]/NET0131  , \P1_P1_InstQueue_reg[15][2]/NET0131  , \P1_P1_InstQueue_reg[15][3]/NET0131  , \P1_P1_InstQueue_reg[15][4]/NET0131  , \P1_P1_InstQueue_reg[15][5]/NET0131  , \P1_P1_InstQueue_reg[15][6]/NET0131  , \P1_P1_InstQueue_reg[15][7]/NET0131  , \P1_P1_InstQueue_reg[1][0]/NET0131  , \P1_P1_InstQueue_reg[1][1]/NET0131  , \P1_P1_InstQueue_reg[1][2]/NET0131  , \P1_P1_InstQueue_reg[1][3]/NET0131  , \P1_P1_InstQueue_reg[1][4]/NET0131  , \P1_P1_InstQueue_reg[1][5]/NET0131  , \P1_P1_InstQueue_reg[1][6]/NET0131  , \P1_P1_InstQueue_reg[1][7]/NET0131  , \P1_P1_InstQueue_reg[2][0]/NET0131  , \P1_P1_InstQueue_reg[2][1]/NET0131  , \P1_P1_InstQueue_reg[2][2]/NET0131  , \P1_P1_InstQueue_reg[2][3]/NET0131  , \P1_P1_InstQueue_reg[2][4]/NET0131  , \P1_P1_InstQueue_reg[2][5]/NET0131  , \P1_P1_InstQueue_reg[2][6]/NET0131  , \P1_P1_InstQueue_reg[2][7]/NET0131  , \P1_P1_InstQueue_reg[3][0]/NET0131  , \P1_P1_InstQueue_reg[3][1]/NET0131  , \P1_P1_InstQueue_reg[3][2]/NET0131  , \P1_P1_InstQueue_reg[3][3]/NET0131  , \P1_P1_InstQueue_reg[3][4]/NET0131  , \P1_P1_InstQueue_reg[3][5]/NET0131  , \P1_P1_InstQueue_reg[3][6]/NET0131  , \P1_P1_InstQueue_reg[3][7]/NET0131  , \P1_P1_InstQueue_reg[4][0]/NET0131  , \P1_P1_InstQueue_reg[4][1]/NET0131  , \P1_P1_InstQueue_reg[4][2]/NET0131  , \P1_P1_InstQueue_reg[4][3]/NET0131  , \P1_P1_InstQueue_reg[4][4]/NET0131  , \P1_P1_InstQueue_reg[4][5]/NET0131  , \P1_P1_InstQueue_reg[4][6]/NET0131  , \P1_P1_InstQueue_reg[4][7]/NET0131  , \P1_P1_InstQueue_reg[5][0]/NET0131  , \P1_P1_InstQueue_reg[5][1]/NET0131  , \P1_P1_InstQueue_reg[5][2]/NET0131  , \P1_P1_InstQueue_reg[5][3]/NET0131  , \P1_P1_InstQueue_reg[5][4]/NET0131  , \P1_P1_InstQueue_reg[5][5]/NET0131  , \P1_P1_InstQueue_reg[5][6]/NET0131  , \P1_P1_InstQueue_reg[5][7]/NET0131  , \P1_P1_InstQueue_reg[6][0]/NET0131  , \P1_P1_InstQueue_reg[6][1]/NET0131  , \P1_P1_InstQueue_reg[6][2]/NET0131  , \P1_P1_InstQueue_reg[6][3]/NET0131  , \P1_P1_InstQueue_reg[6][4]/NET0131  , \P1_P1_InstQueue_reg[6][5]/NET0131  , \P1_P1_InstQueue_reg[6][6]/NET0131  , \P1_P1_InstQueue_reg[6][7]/NET0131  , \P1_P1_InstQueue_reg[7][0]/NET0131  , \P1_P1_InstQueue_reg[7][1]/NET0131  , \P1_P1_InstQueue_reg[7][2]/NET0131  , \P1_P1_InstQueue_reg[7][3]/NET0131  , \P1_P1_InstQueue_reg[7][4]/NET0131  , \P1_P1_InstQueue_reg[7][5]/NET0131  , \P1_P1_InstQueue_reg[7][6]/NET0131  , \P1_P1_InstQueue_reg[7][7]/NET0131  , \P1_P1_InstQueue_reg[8][0]/NET0131  , \P1_P1_InstQueue_reg[8][1]/NET0131  , \P1_P1_InstQueue_reg[8][2]/NET0131  , \P1_P1_InstQueue_reg[8][3]/NET0131  , \P1_P1_InstQueue_reg[8][4]/NET0131  , \P1_P1_InstQueue_reg[8][5]/NET0131  , \P1_P1_InstQueue_reg[8][6]/NET0131  , \P1_P1_InstQueue_reg[8][7]/NET0131  , \P1_P1_InstQueue_reg[9][0]/NET0131  , \P1_P1_InstQueue_reg[9][1]/NET0131  , \P1_P1_InstQueue_reg[9][2]/NET0131  , \P1_P1_InstQueue_reg[9][3]/NET0131  , \P1_P1_InstQueue_reg[9][4]/NET0131  , \P1_P1_InstQueue_reg[9][5]/NET0131  , \P1_P1_InstQueue_reg[9][6]/NET0131  , \P1_P1_InstQueue_reg[9][7]/NET0131  , \P1_P1_M_IO_n_reg/NET0131  , \P1_P1_MemoryFetch_reg/NET0131  , \P1_P1_More_reg/NET0131  , \P1_P1_PhyAddrPointer_reg[0]/NET0131  , \P1_P1_PhyAddrPointer_reg[10]/NET0131  , \P1_P1_PhyAddrPointer_reg[11]/NET0131  , \P1_P1_PhyAddrPointer_reg[12]/NET0131  , \P1_P1_PhyAddrPointer_reg[13]/NET0131  , \P1_P1_PhyAddrPointer_reg[14]/NET0131  , \P1_P1_PhyAddrPointer_reg[15]/NET0131  , \P1_P1_PhyAddrPointer_reg[16]/NET0131  , \P1_P1_PhyAddrPointer_reg[17]/NET0131  , \P1_P1_PhyAddrPointer_reg[18]/NET0131  , \P1_P1_PhyAddrPointer_reg[19]/NET0131  , \P1_P1_PhyAddrPointer_reg[1]/NET0131  , \P1_P1_PhyAddrPointer_reg[20]/NET0131  , \P1_P1_PhyAddrPointer_reg[21]/NET0131  , \P1_P1_PhyAddrPointer_reg[22]/NET0131  , \P1_P1_PhyAddrPointer_reg[23]/NET0131  , \P1_P1_PhyAddrPointer_reg[24]/NET0131  , \P1_P1_PhyAddrPointer_reg[25]/NET0131  , \P1_P1_PhyAddrPointer_reg[26]/NET0131  , \P1_P1_PhyAddrPointer_reg[27]/NET0131  , \P1_P1_PhyAddrPointer_reg[28]/NET0131  , \P1_P1_PhyAddrPointer_reg[29]/NET0131  , \P1_P1_PhyAddrPointer_reg[2]/NET0131  , \P1_P1_PhyAddrPointer_reg[30]/NET0131  , \P1_P1_PhyAddrPointer_reg[31]/NET0131  , \P1_P1_PhyAddrPointer_reg[3]/NET0131  , \P1_P1_PhyAddrPointer_reg[4]/NET0131  , \P1_P1_PhyAddrPointer_reg[5]/NET0131  , \P1_P1_PhyAddrPointer_reg[6]/NET0131  , \P1_P1_PhyAddrPointer_reg[7]/NET0131  , \P1_P1_PhyAddrPointer_reg[8]/NET0131  , \P1_P1_PhyAddrPointer_reg[9]/NET0131  , \P1_P1_ReadRequest_reg/NET0131  , \P1_P1_RequestPending_reg/NET0131  , \P1_P1_State2_reg[0]/NET0131  , \P1_P1_State2_reg[1]/NET0131  , \P1_P1_State2_reg[2]/NET0131  , \P1_P1_State2_reg[3]/NET0131  , \P1_P1_State_reg[0]/NET0131  , \P1_P1_State_reg[1]/NET0131  , \P1_P1_State_reg[2]/NET0131  , \P1_P1_W_R_n_reg/NET0131  , \P1_P1_lWord_reg[0]/NET0131  , \P1_P1_lWord_reg[10]/NET0131  , \P1_P1_lWord_reg[11]/NET0131  , \P1_P1_lWord_reg[12]/NET0131  , \P1_P1_lWord_reg[13]/NET0131  , \P1_P1_lWord_reg[14]/NET0131  , \P1_P1_lWord_reg[15]/NET0131  , \P1_P1_lWord_reg[1]/NET0131  , \P1_P1_lWord_reg[2]/NET0131  , \P1_P1_lWord_reg[3]/NET0131  , \P1_P1_lWord_reg[4]/NET0131  , \P1_P1_lWord_reg[5]/NET0131  , \P1_P1_lWord_reg[6]/NET0131  , \P1_P1_lWord_reg[7]/NET0131  , \P1_P1_lWord_reg[8]/NET0131  , \P1_P1_lWord_reg[9]/NET0131  , \P1_P1_rEIP_reg[0]/NET0131  , \P1_P1_rEIP_reg[10]/NET0131  , \P1_P1_rEIP_reg[11]/NET0131  , \P1_P1_rEIP_reg[12]/NET0131  , \P1_P1_rEIP_reg[13]/NET0131  , \P1_P1_rEIP_reg[14]/NET0131  , \P1_P1_rEIP_reg[15]/NET0131  , \P1_P1_rEIP_reg[16]/NET0131  , \P1_P1_rEIP_reg[17]/NET0131  , \P1_P1_rEIP_reg[18]/NET0131  , \P1_P1_rEIP_reg[19]/NET0131  , \P1_P1_rEIP_reg[1]/NET0131  , \P1_P1_rEIP_reg[20]/NET0131  , \P1_P1_rEIP_reg[21]/NET0131  , \P1_P1_rEIP_reg[22]/NET0131  , \P1_P1_rEIP_reg[23]/NET0131  , \P1_P1_rEIP_reg[24]/NET0131  , \P1_P1_rEIP_reg[25]/NET0131  , \P1_P1_rEIP_reg[26]/NET0131  , \P1_P1_rEIP_reg[27]/NET0131  , \P1_P1_rEIP_reg[28]/NET0131  , \P1_P1_rEIP_reg[29]/NET0131  , \P1_P1_rEIP_reg[2]/NET0131  , \P1_P1_rEIP_reg[30]/NET0131  , \P1_P1_rEIP_reg[31]/NET0131  , \P1_P1_rEIP_reg[3]/NET0131  , \P1_P1_rEIP_reg[4]/NET0131  , \P1_P1_rEIP_reg[5]/NET0131  , \P1_P1_rEIP_reg[6]/NET0131  , \P1_P1_rEIP_reg[7]/NET0131  , \P1_P1_rEIP_reg[8]/NET0131  , \P1_P1_rEIP_reg[9]/NET0131  , \P1_P1_uWord_reg[0]/NET0131  , \P1_P1_uWord_reg[10]/NET0131  , \P1_P1_uWord_reg[11]/NET0131  , \P1_P1_uWord_reg[12]/NET0131  , \P1_P1_uWord_reg[13]/NET0131  , \P1_P1_uWord_reg[14]/NET0131  , \P1_P1_uWord_reg[1]/NET0131  , \P1_P1_uWord_reg[2]/NET0131  , \P1_P1_uWord_reg[3]/NET0131  , \P1_P1_uWord_reg[4]/NET0131  , \P1_P1_uWord_reg[5]/NET0131  , \P1_P1_uWord_reg[6]/NET0131  , \P1_P1_uWord_reg[7]/NET0131  , \P1_P1_uWord_reg[8]/NET0131  , \P1_P1_uWord_reg[9]/NET0131  , \P1_P2_ADS_n_reg/NET0131  , \P1_P2_Address_reg[0]/NET0131  , \P1_P2_Address_reg[10]/NET0131  , \P1_P2_Address_reg[11]/NET0131  , \P1_P2_Address_reg[12]/NET0131  , \P1_P2_Address_reg[13]/NET0131  , \P1_P2_Address_reg[14]/NET0131  , \P1_P2_Address_reg[15]/NET0131  , \P1_P2_Address_reg[16]/NET0131  , \P1_P2_Address_reg[17]/NET0131  , \P1_P2_Address_reg[18]/NET0131  , \P1_P2_Address_reg[19]/NET0131  , \P1_P2_Address_reg[1]/NET0131  , \P1_P2_Address_reg[20]/NET0131  , \P1_P2_Address_reg[21]/NET0131  , \P1_P2_Address_reg[22]/NET0131  , \P1_P2_Address_reg[23]/NET0131  , \P1_P2_Address_reg[24]/NET0131  , \P1_P2_Address_reg[25]/NET0131  , \P1_P2_Address_reg[26]/NET0131  , \P1_P2_Address_reg[27]/NET0131  , \P1_P2_Address_reg[28]/NET0131  , \P1_P2_Address_reg[29]/NET0131  , \P1_P2_Address_reg[2]/NET0131  , \P1_P2_Address_reg[3]/NET0131  , \P1_P2_Address_reg[4]/NET0131  , \P1_P2_Address_reg[5]/NET0131  , \P1_P2_Address_reg[6]/NET0131  , \P1_P2_Address_reg[7]/NET0131  , \P1_P2_Address_reg[8]/NET0131  , \P1_P2_Address_reg[9]/NET0131  , \P1_P2_BE_n_reg[0]/NET0131  , \P1_P2_BE_n_reg[1]/NET0131  , \P1_P2_BE_n_reg[2]/NET0131  , \P1_P2_BE_n_reg[3]/NET0131  , \P1_P2_ByteEnable_reg[0]/NET0131  , \P1_P2_ByteEnable_reg[1]/NET0131  , \P1_P2_ByteEnable_reg[2]/NET0131  , \P1_P2_ByteEnable_reg[3]/NET0131  , \P1_P2_CodeFetch_reg/NET0131  , \P1_P2_D_C_n_reg/NET0131  , \P1_P2_DataWidth_reg[0]/NET0131  , \P1_P2_DataWidth_reg[1]/NET0131  , \P1_P2_Datao_reg[0]/NET0131  , \P1_P2_Datao_reg[10]/NET0131  , \P1_P2_Datao_reg[11]/NET0131  , \P1_P2_Datao_reg[12]/NET0131  , \P1_P2_Datao_reg[13]/NET0131  , \P1_P2_Datao_reg[14]/NET0131  , \P1_P2_Datao_reg[15]/NET0131  , \P1_P2_Datao_reg[16]/NET0131  , \P1_P2_Datao_reg[17]/NET0131  , \P1_P2_Datao_reg[18]/NET0131  , \P1_P2_Datao_reg[19]/NET0131  , \P1_P2_Datao_reg[1]/NET0131  , \P1_P2_Datao_reg[20]/NET0131  , \P1_P2_Datao_reg[21]/NET0131  , \P1_P2_Datao_reg[22]/NET0131  , \P1_P2_Datao_reg[23]/NET0131  , \P1_P2_Datao_reg[24]/NET0131  , \P1_P2_Datao_reg[25]/NET0131  , \P1_P2_Datao_reg[26]/NET0131  , \P1_P2_Datao_reg[27]/NET0131  , \P1_P2_Datao_reg[28]/NET0131  , \P1_P2_Datao_reg[29]/NET0131  , \P1_P2_Datao_reg[2]/NET0131  , \P1_P2_Datao_reg[30]/NET0131  , \P1_P2_Datao_reg[3]/NET0131  , \P1_P2_Datao_reg[4]/NET0131  , \P1_P2_Datao_reg[5]/NET0131  , \P1_P2_Datao_reg[6]/NET0131  , \P1_P2_Datao_reg[7]/NET0131  , \P1_P2_Datao_reg[8]/NET0131  , \P1_P2_Datao_reg[9]/NET0131  , \P1_P2_EAX_reg[0]/NET0131  , \P1_P2_EAX_reg[10]/NET0131  , \P1_P2_EAX_reg[11]/NET0131  , \P1_P2_EAX_reg[12]/NET0131  , \P1_P2_EAX_reg[13]/NET0131  , \P1_P2_EAX_reg[14]/NET0131  , \P1_P2_EAX_reg[15]/NET0131  , \P1_P2_EAX_reg[16]/NET0131  , \P1_P2_EAX_reg[17]/NET0131  , \P1_P2_EAX_reg[18]/NET0131  , \P1_P2_EAX_reg[19]/NET0131  , \P1_P2_EAX_reg[1]/NET0131  , \P1_P2_EAX_reg[20]/NET0131  , \P1_P2_EAX_reg[21]/NET0131  , \P1_P2_EAX_reg[22]/NET0131  , \P1_P2_EAX_reg[23]/NET0131  , \P1_P2_EAX_reg[24]/NET0131  , \P1_P2_EAX_reg[25]/NET0131  , \P1_P2_EAX_reg[26]/NET0131  , \P1_P2_EAX_reg[27]/NET0131  , \P1_P2_EAX_reg[28]/NET0131  , \P1_P2_EAX_reg[29]/NET0131  , \P1_P2_EAX_reg[2]/NET0131  , \P1_P2_EAX_reg[30]/NET0131  , \P1_P2_EAX_reg[31]/NET0131  , \P1_P2_EAX_reg[3]/NET0131  , \P1_P2_EAX_reg[4]/NET0131  , \P1_P2_EAX_reg[5]/NET0131  , \P1_P2_EAX_reg[6]/NET0131  , \P1_P2_EAX_reg[7]/NET0131  , \P1_P2_EAX_reg[8]/NET0131  , \P1_P2_EAX_reg[9]/NET0131  , \P1_P2_EBX_reg[0]/NET0131  , \P1_P2_EBX_reg[10]/NET0131  , \P1_P2_EBX_reg[11]/NET0131  , \P1_P2_EBX_reg[12]/NET0131  , \P1_P2_EBX_reg[13]/NET0131  , \P1_P2_EBX_reg[14]/NET0131  , \P1_P2_EBX_reg[15]/NET0131  , \P1_P2_EBX_reg[16]/NET0131  , \P1_P2_EBX_reg[17]/NET0131  , \P1_P2_EBX_reg[18]/NET0131  , \P1_P2_EBX_reg[19]/NET0131  , \P1_P2_EBX_reg[1]/NET0131  , \P1_P2_EBX_reg[20]/NET0131  , \P1_P2_EBX_reg[21]/NET0131  , \P1_P2_EBX_reg[22]/NET0131  , \P1_P2_EBX_reg[23]/NET0131  , \P1_P2_EBX_reg[24]/NET0131  , \P1_P2_EBX_reg[25]/NET0131  , \P1_P2_EBX_reg[26]/NET0131  , \P1_P2_EBX_reg[27]/NET0131  , \P1_P2_EBX_reg[28]/NET0131  , \P1_P2_EBX_reg[29]/NET0131  , \P1_P2_EBX_reg[2]/NET0131  , \P1_P2_EBX_reg[30]/NET0131  , \P1_P2_EBX_reg[31]/NET0131  , \P1_P2_EBX_reg[3]/NET0131  , \P1_P2_EBX_reg[4]/NET0131  , \P1_P2_EBX_reg[5]/NET0131  , \P1_P2_EBX_reg[6]/NET0131  , \P1_P2_EBX_reg[7]/NET0131  , \P1_P2_EBX_reg[8]/NET0131  , \P1_P2_EBX_reg[9]/NET0131  , \P1_P2_Flush_reg/NET0131  , \P1_P2_InstAddrPointer_reg[0]/NET0131  , \P1_P2_InstAddrPointer_reg[10]/NET0131  , \P1_P2_InstAddrPointer_reg[11]/NET0131  , \P1_P2_InstAddrPointer_reg[12]/NET0131  , \P1_P2_InstAddrPointer_reg[13]/NET0131  , \P1_P2_InstAddrPointer_reg[14]/NET0131  , \P1_P2_InstAddrPointer_reg[15]/NET0131  , \P1_P2_InstAddrPointer_reg[16]/NET0131  , \P1_P2_InstAddrPointer_reg[17]/NET0131  , \P1_P2_InstAddrPointer_reg[18]/NET0131  , \P1_P2_InstAddrPointer_reg[19]/NET0131  , \P1_P2_InstAddrPointer_reg[1]/NET0131  , \P1_P2_InstAddrPointer_reg[20]/NET0131  , \P1_P2_InstAddrPointer_reg[21]/NET0131  , \P1_P2_InstAddrPointer_reg[22]/NET0131  , \P1_P2_InstAddrPointer_reg[23]/NET0131  , \P1_P2_InstAddrPointer_reg[24]/NET0131  , \P1_P2_InstAddrPointer_reg[25]/NET0131  , \P1_P2_InstAddrPointer_reg[26]/NET0131  , \P1_P2_InstAddrPointer_reg[27]/NET0131  , \P1_P2_InstAddrPointer_reg[28]/NET0131  , \P1_P2_InstAddrPointer_reg[29]/NET0131  , \P1_P2_InstAddrPointer_reg[2]/NET0131  , \P1_P2_InstAddrPointer_reg[30]/NET0131  , \P1_P2_InstAddrPointer_reg[31]/NET0131  , \P1_P2_InstAddrPointer_reg[3]/NET0131  , \P1_P2_InstAddrPointer_reg[4]/NET0131  , \P1_P2_InstAddrPointer_reg[5]/NET0131  , \P1_P2_InstAddrPointer_reg[6]/NET0131  , \P1_P2_InstAddrPointer_reg[7]/NET0131  , \P1_P2_InstAddrPointer_reg[8]/NET0131  , \P1_P2_InstAddrPointer_reg[9]/NET0131  , \P1_P2_InstQueueRd_Addr_reg[0]/NET0131  , \P1_P2_InstQueueRd_Addr_reg[1]/NET0131  , \P1_P2_InstQueueRd_Addr_reg[2]/NET0131  , \P1_P2_InstQueueRd_Addr_reg[3]/NET0131  , \P1_P2_InstQueueWr_Addr_reg[0]/NET0131  , \P1_P2_InstQueueWr_Addr_reg[1]/NET0131  , \P1_P2_InstQueueWr_Addr_reg[2]/NET0131  , \P1_P2_InstQueueWr_Addr_reg[3]/NET0131  , \P1_P2_InstQueue_reg[0][0]/NET0131  , \P1_P2_InstQueue_reg[0][1]/NET0131  , \P1_P2_InstQueue_reg[0][2]/NET0131  , \P1_P2_InstQueue_reg[0][3]/NET0131  , \P1_P2_InstQueue_reg[0][4]/NET0131  , \P1_P2_InstQueue_reg[0][5]/NET0131  , \P1_P2_InstQueue_reg[0][6]/NET0131  , \P1_P2_InstQueue_reg[0][7]/NET0131  , \P1_P2_InstQueue_reg[10][0]/NET0131  , \P1_P2_InstQueue_reg[10][1]/NET0131  , \P1_P2_InstQueue_reg[10][2]/NET0131  , \P1_P2_InstQueue_reg[10][3]/NET0131  , \P1_P2_InstQueue_reg[10][4]/NET0131  , \P1_P2_InstQueue_reg[10][5]/NET0131  , \P1_P2_InstQueue_reg[10][6]/NET0131  , \P1_P2_InstQueue_reg[10][7]/NET0131  , \P1_P2_InstQueue_reg[11][0]/NET0131  , \P1_P2_InstQueue_reg[11][1]/NET0131  , \P1_P2_InstQueue_reg[11][2]/NET0131  , \P1_P2_InstQueue_reg[11][3]/NET0131  , \P1_P2_InstQueue_reg[11][4]/NET0131  , \P1_P2_InstQueue_reg[11][5]/NET0131  , \P1_P2_InstQueue_reg[11][6]/NET0131  , \P1_P2_InstQueue_reg[11][7]/NET0131  , \P1_P2_InstQueue_reg[12][0]/NET0131  , \P1_P2_InstQueue_reg[12][1]/NET0131  , \P1_P2_InstQueue_reg[12][2]/NET0131  , \P1_P2_InstQueue_reg[12][3]/NET0131  , \P1_P2_InstQueue_reg[12][4]/NET0131  , \P1_P2_InstQueue_reg[12][5]/NET0131  , \P1_P2_InstQueue_reg[12][6]/NET0131  , \P1_P2_InstQueue_reg[12][7]/NET0131  , \P1_P2_InstQueue_reg[13][0]/NET0131  , \P1_P2_InstQueue_reg[13][1]/NET0131  , \P1_P2_InstQueue_reg[13][2]/NET0131  , \P1_P2_InstQueue_reg[13][3]/NET0131  , \P1_P2_InstQueue_reg[13][4]/NET0131  , \P1_P2_InstQueue_reg[13][5]/NET0131  , \P1_P2_InstQueue_reg[13][6]/NET0131  , \P1_P2_InstQueue_reg[13][7]/NET0131  , \P1_P2_InstQueue_reg[14][0]/NET0131  , \P1_P2_InstQueue_reg[14][1]/NET0131  , \P1_P2_InstQueue_reg[14][2]/NET0131  , \P1_P2_InstQueue_reg[14][3]/NET0131  , \P1_P2_InstQueue_reg[14][4]/NET0131  , \P1_P2_InstQueue_reg[14][5]/NET0131  , \P1_P2_InstQueue_reg[14][6]/NET0131  , \P1_P2_InstQueue_reg[14][7]/NET0131  , \P1_P2_InstQueue_reg[15][0]/NET0131  , \P1_P2_InstQueue_reg[15][1]/NET0131  , \P1_P2_InstQueue_reg[15][2]/NET0131  , \P1_P2_InstQueue_reg[15][3]/NET0131  , \P1_P2_InstQueue_reg[15][4]/NET0131  , \P1_P2_InstQueue_reg[15][5]/NET0131  , \P1_P2_InstQueue_reg[15][6]/NET0131  , \P1_P2_InstQueue_reg[15][7]/NET0131  , \P1_P2_InstQueue_reg[1][0]/NET0131  , \P1_P2_InstQueue_reg[1][1]/NET0131  , \P1_P2_InstQueue_reg[1][2]/NET0131  , \P1_P2_InstQueue_reg[1][3]/NET0131  , \P1_P2_InstQueue_reg[1][4]/NET0131  , \P1_P2_InstQueue_reg[1][5]/NET0131  , \P1_P2_InstQueue_reg[1][6]/NET0131  , \P1_P2_InstQueue_reg[1][7]/NET0131  , \P1_P2_InstQueue_reg[2][0]/NET0131  , \P1_P2_InstQueue_reg[2][1]/NET0131  , \P1_P2_InstQueue_reg[2][2]/NET0131  , \P1_P2_InstQueue_reg[2][3]/NET0131  , \P1_P2_InstQueue_reg[2][4]/NET0131  , \P1_P2_InstQueue_reg[2][5]/NET0131  , \P1_P2_InstQueue_reg[2][6]/NET0131  , \P1_P2_InstQueue_reg[2][7]/NET0131  , \P1_P2_InstQueue_reg[3][0]/NET0131  , \P1_P2_InstQueue_reg[3][1]/NET0131  , \P1_P2_InstQueue_reg[3][2]/NET0131  , \P1_P2_InstQueue_reg[3][3]/NET0131  , \P1_P2_InstQueue_reg[3][4]/NET0131  , \P1_P2_InstQueue_reg[3][5]/NET0131  , \P1_P2_InstQueue_reg[3][6]/NET0131  , \P1_P2_InstQueue_reg[3][7]/NET0131  , \P1_P2_InstQueue_reg[4][0]/NET0131  , \P1_P2_InstQueue_reg[4][1]/NET0131  , \P1_P2_InstQueue_reg[4][2]/NET0131  , \P1_P2_InstQueue_reg[4][3]/NET0131  , \P1_P2_InstQueue_reg[4][4]/NET0131  , \P1_P2_InstQueue_reg[4][5]/NET0131  , \P1_P2_InstQueue_reg[4][6]/NET0131  , \P1_P2_InstQueue_reg[4][7]/NET0131  , \P1_P2_InstQueue_reg[5][0]/NET0131  , \P1_P2_InstQueue_reg[5][1]/NET0131  , \P1_P2_InstQueue_reg[5][2]/NET0131  , \P1_P2_InstQueue_reg[5][3]/NET0131  , \P1_P2_InstQueue_reg[5][4]/NET0131  , \P1_P2_InstQueue_reg[5][5]/NET0131  , \P1_P2_InstQueue_reg[5][6]/NET0131  , \P1_P2_InstQueue_reg[5][7]/NET0131  , \P1_P2_InstQueue_reg[6][0]/NET0131  , \P1_P2_InstQueue_reg[6][1]/NET0131  , \P1_P2_InstQueue_reg[6][2]/NET0131  , \P1_P2_InstQueue_reg[6][3]/NET0131  , \P1_P2_InstQueue_reg[6][4]/NET0131  , \P1_P2_InstQueue_reg[6][5]/NET0131  , \P1_P2_InstQueue_reg[6][6]/NET0131  , \P1_P2_InstQueue_reg[6][7]/NET0131  , \P1_P2_InstQueue_reg[7][0]/NET0131  , \P1_P2_InstQueue_reg[7][1]/NET0131  , \P1_P2_InstQueue_reg[7][2]/NET0131  , \P1_P2_InstQueue_reg[7][3]/NET0131  , \P1_P2_InstQueue_reg[7][4]/NET0131  , \P1_P2_InstQueue_reg[7][5]/NET0131  , \P1_P2_InstQueue_reg[7][6]/NET0131  , \P1_P2_InstQueue_reg[7][7]/NET0131  , \P1_P2_InstQueue_reg[8][0]/NET0131  , \P1_P2_InstQueue_reg[8][1]/NET0131  , \P1_P2_InstQueue_reg[8][2]/NET0131  , \P1_P2_InstQueue_reg[8][3]/NET0131  , \P1_P2_InstQueue_reg[8][4]/NET0131  , \P1_P2_InstQueue_reg[8][5]/NET0131  , \P1_P2_InstQueue_reg[8][6]/NET0131  , \P1_P2_InstQueue_reg[8][7]/NET0131  , \P1_P2_InstQueue_reg[9][0]/NET0131  , \P1_P2_InstQueue_reg[9][1]/NET0131  , \P1_P2_InstQueue_reg[9][2]/NET0131  , \P1_P2_InstQueue_reg[9][3]/NET0131  , \P1_P2_InstQueue_reg[9][4]/NET0131  , \P1_P2_InstQueue_reg[9][5]/NET0131  , \P1_P2_InstQueue_reg[9][6]/NET0131  , \P1_P2_InstQueue_reg[9][7]/NET0131  , \P1_P2_M_IO_n_reg/NET0131  , \P1_P2_MemoryFetch_reg/NET0131  , \P1_P2_More_reg/NET0131  , \P1_P2_PhyAddrPointer_reg[0]/NET0131  , \P1_P2_PhyAddrPointer_reg[10]/NET0131  , \P1_P2_PhyAddrPointer_reg[11]/NET0131  , \P1_P2_PhyAddrPointer_reg[12]/NET0131  , \P1_P2_PhyAddrPointer_reg[13]/NET0131  , \P1_P2_PhyAddrPointer_reg[14]/NET0131  , \P1_P2_PhyAddrPointer_reg[15]/NET0131  , \P1_P2_PhyAddrPointer_reg[16]/NET0131  , \P1_P2_PhyAddrPointer_reg[17]/NET0131  , \P1_P2_PhyAddrPointer_reg[18]/NET0131  , \P1_P2_PhyAddrPointer_reg[19]/NET0131  , \P1_P2_PhyAddrPointer_reg[1]/NET0131  , \P1_P2_PhyAddrPointer_reg[20]/NET0131  , \P1_P2_PhyAddrPointer_reg[21]/NET0131  , \P1_P2_PhyAddrPointer_reg[22]/NET0131  , \P1_P2_PhyAddrPointer_reg[23]/NET0131  , \P1_P2_PhyAddrPointer_reg[24]/NET0131  , \P1_P2_PhyAddrPointer_reg[25]/NET0131  , \P1_P2_PhyAddrPointer_reg[26]/NET0131  , \P1_P2_PhyAddrPointer_reg[27]/NET0131  , \P1_P2_PhyAddrPointer_reg[28]/NET0131  , \P1_P2_PhyAddrPointer_reg[29]/NET0131  , \P1_P2_PhyAddrPointer_reg[2]/NET0131  , \P1_P2_PhyAddrPointer_reg[30]/NET0131  , \P1_P2_PhyAddrPointer_reg[31]/NET0131  , \P1_P2_PhyAddrPointer_reg[3]/NET0131  , \P1_P2_PhyAddrPointer_reg[4]/NET0131  , \P1_P2_PhyAddrPointer_reg[5]/NET0131  , \P1_P2_PhyAddrPointer_reg[6]/NET0131  , \P1_P2_PhyAddrPointer_reg[7]/NET0131  , \P1_P2_PhyAddrPointer_reg[8]/NET0131  , \P1_P2_PhyAddrPointer_reg[9]/NET0131  , \P1_P2_ReadRequest_reg/NET0131  , \P1_P2_RequestPending_reg/NET0131  , \P1_P2_State2_reg[0]/NET0131  , \P1_P2_State2_reg[1]/NET0131  , \P1_P2_State2_reg[2]/NET0131  , \P1_P2_State2_reg[3]/NET0131  , \P1_P2_State_reg[0]/NET0131  , \P1_P2_State_reg[1]/NET0131  , \P1_P2_State_reg[2]/NET0131  , \P1_P2_W_R_n_reg/NET0131  , \P1_P2_lWord_reg[0]/NET0131  , \P1_P2_lWord_reg[10]/NET0131  , \P1_P2_lWord_reg[11]/NET0131  , \P1_P2_lWord_reg[12]/NET0131  , \P1_P2_lWord_reg[13]/NET0131  , \P1_P2_lWord_reg[14]/NET0131  , \P1_P2_lWord_reg[15]/NET0131  , \P1_P2_lWord_reg[1]/NET0131  , \P1_P2_lWord_reg[2]/NET0131  , \P1_P2_lWord_reg[3]/NET0131  , \P1_P2_lWord_reg[4]/NET0131  , \P1_P2_lWord_reg[5]/NET0131  , \P1_P2_lWord_reg[6]/NET0131  , \P1_P2_lWord_reg[7]/NET0131  , \P1_P2_lWord_reg[8]/NET0131  , \P1_P2_lWord_reg[9]/NET0131  , \P1_P2_rEIP_reg[0]/NET0131  , \P1_P2_rEIP_reg[10]/NET0131  , \P1_P2_rEIP_reg[11]/NET0131  , \P1_P2_rEIP_reg[12]/NET0131  , \P1_P2_rEIP_reg[13]/NET0131  , \P1_P2_rEIP_reg[14]/NET0131  , \P1_P2_rEIP_reg[15]/NET0131  , \P1_P2_rEIP_reg[16]/NET0131  , \P1_P2_rEIP_reg[17]/NET0131  , \P1_P2_rEIP_reg[18]/NET0131  , \P1_P2_rEIP_reg[19]/NET0131  , \P1_P2_rEIP_reg[1]/NET0131  , \P1_P2_rEIP_reg[20]/NET0131  , \P1_P2_rEIP_reg[21]/NET0131  , \P1_P2_rEIP_reg[22]/NET0131  , \P1_P2_rEIP_reg[23]/NET0131  , \P1_P2_rEIP_reg[24]/NET0131  , \P1_P2_rEIP_reg[25]/NET0131  , \P1_P2_rEIP_reg[26]/NET0131  , \P1_P2_rEIP_reg[27]/NET0131  , \P1_P2_rEIP_reg[28]/NET0131  , \P1_P2_rEIP_reg[29]/NET0131  , \P1_P2_rEIP_reg[2]/NET0131  , \P1_P2_rEIP_reg[30]/NET0131  , \P1_P2_rEIP_reg[31]/NET0131  , \P1_P2_rEIP_reg[3]/NET0131  , \P1_P2_rEIP_reg[4]/NET0131  , \P1_P2_rEIP_reg[5]/NET0131  , \P1_P2_rEIP_reg[6]/NET0131  , \P1_P2_rEIP_reg[7]/NET0131  , \P1_P2_rEIP_reg[8]/NET0131  , \P1_P2_rEIP_reg[9]/NET0131  , \P1_P2_uWord_reg[0]/NET0131  , \P1_P2_uWord_reg[10]/NET0131  , \P1_P2_uWord_reg[11]/NET0131  , \P1_P2_uWord_reg[12]/NET0131  , \P1_P2_uWord_reg[13]/NET0131  , \P1_P2_uWord_reg[14]/NET0131  , \P1_P2_uWord_reg[1]/NET0131  , \P1_P2_uWord_reg[2]/NET0131  , \P1_P2_uWord_reg[3]/NET0131  , \P1_P2_uWord_reg[4]/NET0131  , \P1_P2_uWord_reg[5]/NET0131  , \P1_P2_uWord_reg[6]/NET0131  , \P1_P2_uWord_reg[7]/NET0131  , \P1_P2_uWord_reg[8]/NET0131  , \P1_P2_uWord_reg[9]/NET0131  , \P1_P3_ADS_n_reg/NET0131  , \P1_P3_Address_reg[0]/NET0131  , \P1_P3_Address_reg[10]/NET0131  , \P1_P3_Address_reg[11]/NET0131  , \P1_P3_Address_reg[12]/NET0131  , \P1_P3_Address_reg[13]/NET0131  , \P1_P3_Address_reg[14]/NET0131  , \P1_P3_Address_reg[15]/NET0131  , \P1_P3_Address_reg[16]/NET0131  , \P1_P3_Address_reg[17]/NET0131  , \P1_P3_Address_reg[18]/NET0131  , \P1_P3_Address_reg[1]/NET0131  , \P1_P3_Address_reg[2]/NET0131  , \P1_P3_Address_reg[3]/NET0131  , \P1_P3_Address_reg[4]/NET0131  , \P1_P3_Address_reg[5]/NET0131  , \P1_P3_Address_reg[6]/NET0131  , \P1_P3_Address_reg[7]/NET0131  , \P1_P3_Address_reg[8]/NET0131  , \P1_P3_Address_reg[9]/NET0131  , \P1_P3_BE_n_reg[0]/NET0131  , \P1_P3_BE_n_reg[1]/NET0131  , \P1_P3_BE_n_reg[2]/NET0131  , \P1_P3_BE_n_reg[3]/NET0131  , \P1_P3_ByteEnable_reg[0]/NET0131  , \P1_P3_ByteEnable_reg[1]/NET0131  , \P1_P3_ByteEnable_reg[2]/NET0131  , \P1_P3_ByteEnable_reg[3]/NET0131  , \P1_P3_CodeFetch_reg/NET0131  , \P1_P3_D_C_n_reg/NET0131  , \P1_P3_DataWidth_reg[0]/NET0131  , \P1_P3_DataWidth_reg[1]/NET0131  , \P1_P3_Datao_reg[30]/NET0131  , \P1_P3_EAX_reg[0]/NET0131  , \P1_P3_EAX_reg[10]/NET0131  , \P1_P3_EAX_reg[11]/NET0131  , \P1_P3_EAX_reg[12]/NET0131  , \P1_P3_EAX_reg[13]/NET0131  , \P1_P3_EAX_reg[14]/NET0131  , \P1_P3_EAX_reg[15]/NET0131  , \P1_P3_EAX_reg[16]/NET0131  , \P1_P3_EAX_reg[17]/NET0131  , \P1_P3_EAX_reg[18]/NET0131  , \P1_P3_EAX_reg[19]/NET0131  , \P1_P3_EAX_reg[1]/NET0131  , \P1_P3_EAX_reg[20]/NET0131  , \P1_P3_EAX_reg[21]/NET0131  , \P1_P3_EAX_reg[22]/NET0131  , \P1_P3_EAX_reg[23]/NET0131  , \P1_P3_EAX_reg[24]/NET0131  , \P1_P3_EAX_reg[25]/NET0131  , \P1_P3_EAX_reg[26]/NET0131  , \P1_P3_EAX_reg[27]/NET0131  , \P1_P3_EAX_reg[28]/NET0131  , \P1_P3_EAX_reg[29]/NET0131  , \P1_P3_EAX_reg[2]/NET0131  , \P1_P3_EAX_reg[30]/NET0131  , \P1_P3_EAX_reg[31]/NET0131  , \P1_P3_EAX_reg[3]/NET0131  , \P1_P3_EAX_reg[4]/NET0131  , \P1_P3_EAX_reg[5]/NET0131  , \P1_P3_EAX_reg[6]/NET0131  , \P1_P3_EAX_reg[7]/NET0131  , \P1_P3_EAX_reg[8]/NET0131  , \P1_P3_EAX_reg[9]/NET0131  , \P1_P3_EBX_reg[0]/NET0131  , \P1_P3_EBX_reg[10]/NET0131  , \P1_P3_EBX_reg[11]/NET0131  , \P1_P3_EBX_reg[12]/NET0131  , \P1_P3_EBX_reg[13]/NET0131  , \P1_P3_EBX_reg[14]/NET0131  , \P1_P3_EBX_reg[15]/NET0131  , \P1_P3_EBX_reg[16]/NET0131  , \P1_P3_EBX_reg[17]/NET0131  , \P1_P3_EBX_reg[18]/NET0131  , \P1_P3_EBX_reg[19]/NET0131  , \P1_P3_EBX_reg[1]/NET0131  , \P1_P3_EBX_reg[20]/NET0131  , \P1_P3_EBX_reg[21]/NET0131  , \P1_P3_EBX_reg[22]/NET0131  , \P1_P3_EBX_reg[23]/NET0131  , \P1_P3_EBX_reg[24]/NET0131  , \P1_P3_EBX_reg[25]/NET0131  , \P1_P3_EBX_reg[26]/NET0131  , \P1_P3_EBX_reg[27]/NET0131  , \P1_P3_EBX_reg[28]/NET0131  , \P1_P3_EBX_reg[29]/NET0131  , \P1_P3_EBX_reg[2]/NET0131  , \P1_P3_EBX_reg[30]/NET0131  , \P1_P3_EBX_reg[31]/NET0131  , \P1_P3_EBX_reg[3]/NET0131  , \P1_P3_EBX_reg[4]/NET0131  , \P1_P3_EBX_reg[5]/NET0131  , \P1_P3_EBX_reg[6]/NET0131  , \P1_P3_EBX_reg[7]/NET0131  , \P1_P3_EBX_reg[8]/NET0131  , \P1_P3_EBX_reg[9]/NET0131  , \P1_P3_Flush_reg/NET0131  , \P1_P3_InstAddrPointer_reg[0]/NET0131  , \P1_P3_InstAddrPointer_reg[10]/NET0131  , \P1_P3_InstAddrPointer_reg[11]/NET0131  , \P1_P3_InstAddrPointer_reg[12]/NET0131  , \P1_P3_InstAddrPointer_reg[13]/NET0131  , \P1_P3_InstAddrPointer_reg[14]/NET0131  , \P1_P3_InstAddrPointer_reg[15]/NET0131  , \P1_P3_InstAddrPointer_reg[16]/NET0131  , \P1_P3_InstAddrPointer_reg[17]/NET0131  , \P1_P3_InstAddrPointer_reg[18]/NET0131  , \P1_P3_InstAddrPointer_reg[19]/NET0131  , \P1_P3_InstAddrPointer_reg[1]/NET0131  , \P1_P3_InstAddrPointer_reg[20]/NET0131  , \P1_P3_InstAddrPointer_reg[21]/NET0131  , \P1_P3_InstAddrPointer_reg[22]/NET0131  , \P1_P3_InstAddrPointer_reg[23]/NET0131  , \P1_P3_InstAddrPointer_reg[24]/NET0131  , \P1_P3_InstAddrPointer_reg[25]/NET0131  , \P1_P3_InstAddrPointer_reg[26]/NET0131  , \P1_P3_InstAddrPointer_reg[27]/NET0131  , \P1_P3_InstAddrPointer_reg[28]/NET0131  , \P1_P3_InstAddrPointer_reg[29]/NET0131  , \P1_P3_InstAddrPointer_reg[2]/NET0131  , \P1_P3_InstAddrPointer_reg[30]/NET0131  , \P1_P3_InstAddrPointer_reg[31]/NET0131  , \P1_P3_InstAddrPointer_reg[3]/NET0131  , \P1_P3_InstAddrPointer_reg[4]/NET0131  , \P1_P3_InstAddrPointer_reg[5]/NET0131  , \P1_P3_InstAddrPointer_reg[6]/NET0131  , \P1_P3_InstAddrPointer_reg[7]/NET0131  , \P1_P3_InstAddrPointer_reg[8]/NET0131  , \P1_P3_InstAddrPointer_reg[9]/NET0131  , \P1_P3_InstQueueRd_Addr_reg[0]/NET0131  , \P1_P3_InstQueueRd_Addr_reg[1]/NET0131  , \P1_P3_InstQueueRd_Addr_reg[2]/NET0131  , \P1_P3_InstQueueRd_Addr_reg[3]/NET0131  , \P1_P3_InstQueueWr_Addr_reg[0]/NET0131  , \P1_P3_InstQueueWr_Addr_reg[1]/NET0131  , \P1_P3_InstQueueWr_Addr_reg[2]/NET0131  , \P1_P3_InstQueueWr_Addr_reg[3]/NET0131  , \P1_P3_InstQueue_reg[0][0]/NET0131  , \P1_P3_InstQueue_reg[0][1]/NET0131  , \P1_P3_InstQueue_reg[0][2]/NET0131  , \P1_P3_InstQueue_reg[0][3]/NET0131  , \P1_P3_InstQueue_reg[0][4]/NET0131  , \P1_P3_InstQueue_reg[0][5]/NET0131  , \P1_P3_InstQueue_reg[0][6]/NET0131  , \P1_P3_InstQueue_reg[0][7]/NET0131  , \P1_P3_InstQueue_reg[10][0]/NET0131  , \P1_P3_InstQueue_reg[10][1]/NET0131  , \P1_P3_InstQueue_reg[10][2]/NET0131  , \P1_P3_InstQueue_reg[10][3]/NET0131  , \P1_P3_InstQueue_reg[10][4]/NET0131  , \P1_P3_InstQueue_reg[10][5]/NET0131  , \P1_P3_InstQueue_reg[10][6]/NET0131  , \P1_P3_InstQueue_reg[10][7]/NET0131  , \P1_P3_InstQueue_reg[11][0]/NET0131  , \P1_P3_InstQueue_reg[11][1]/NET0131  , \P1_P3_InstQueue_reg[11][2]/NET0131  , \P1_P3_InstQueue_reg[11][3]/NET0131  , \P1_P3_InstQueue_reg[11][4]/NET0131  , \P1_P3_InstQueue_reg[11][5]/NET0131  , \P1_P3_InstQueue_reg[11][6]/NET0131  , \P1_P3_InstQueue_reg[11][7]/NET0131  , \P1_P3_InstQueue_reg[12][0]/NET0131  , \P1_P3_InstQueue_reg[12][1]/NET0131  , \P1_P3_InstQueue_reg[12][2]/NET0131  , \P1_P3_InstQueue_reg[12][3]/NET0131  , \P1_P3_InstQueue_reg[12][4]/NET0131  , \P1_P3_InstQueue_reg[12][5]/NET0131  , \P1_P3_InstQueue_reg[12][6]/NET0131  , \P1_P3_InstQueue_reg[12][7]/NET0131  , \P1_P3_InstQueue_reg[13][0]/NET0131  , \P1_P3_InstQueue_reg[13][1]/NET0131  , \P1_P3_InstQueue_reg[13][2]/NET0131  , \P1_P3_InstQueue_reg[13][3]/NET0131  , \P1_P3_InstQueue_reg[13][4]/NET0131  , \P1_P3_InstQueue_reg[13][5]/NET0131  , \P1_P3_InstQueue_reg[13][6]/NET0131  , \P1_P3_InstQueue_reg[13][7]/NET0131  , \P1_P3_InstQueue_reg[14][0]/NET0131  , \P1_P3_InstQueue_reg[14][1]/NET0131  , \P1_P3_InstQueue_reg[14][2]/NET0131  , \P1_P3_InstQueue_reg[14][3]/NET0131  , \P1_P3_InstQueue_reg[14][4]/NET0131  , \P1_P3_InstQueue_reg[14][5]/NET0131  , \P1_P3_InstQueue_reg[14][6]/NET0131  , \P1_P3_InstQueue_reg[14][7]/NET0131  , \P1_P3_InstQueue_reg[15][0]/NET0131  , \P1_P3_InstQueue_reg[15][1]/NET0131  , \P1_P3_InstQueue_reg[15][2]/NET0131  , \P1_P3_InstQueue_reg[15][3]/NET0131  , \P1_P3_InstQueue_reg[15][4]/NET0131  , \P1_P3_InstQueue_reg[15][5]/NET0131  , \P1_P3_InstQueue_reg[15][6]/NET0131  , \P1_P3_InstQueue_reg[15][7]/NET0131  , \P1_P3_InstQueue_reg[1][0]/NET0131  , \P1_P3_InstQueue_reg[1][1]/NET0131  , \P1_P3_InstQueue_reg[1][2]/NET0131  , \P1_P3_InstQueue_reg[1][3]/NET0131  , \P1_P3_InstQueue_reg[1][4]/NET0131  , \P1_P3_InstQueue_reg[1][5]/NET0131  , \P1_P3_InstQueue_reg[1][6]/NET0131  , \P1_P3_InstQueue_reg[1][7]/NET0131  , \P1_P3_InstQueue_reg[2][0]/NET0131  , \P1_P3_InstQueue_reg[2][1]/NET0131  , \P1_P3_InstQueue_reg[2][2]/NET0131  , \P1_P3_InstQueue_reg[2][3]/NET0131  , \P1_P3_InstQueue_reg[2][4]/NET0131  , \P1_P3_InstQueue_reg[2][5]/NET0131  , \P1_P3_InstQueue_reg[2][6]/NET0131  , \P1_P3_InstQueue_reg[2][7]/NET0131  , \P1_P3_InstQueue_reg[3][0]/NET0131  , \P1_P3_InstQueue_reg[3][1]/NET0131  , \P1_P3_InstQueue_reg[3][2]/NET0131  , \P1_P3_InstQueue_reg[3][3]/NET0131  , \P1_P3_InstQueue_reg[3][4]/NET0131  , \P1_P3_InstQueue_reg[3][5]/NET0131  , \P1_P3_InstQueue_reg[3][6]/NET0131  , \P1_P3_InstQueue_reg[3][7]/NET0131  , \P1_P3_InstQueue_reg[4][0]/NET0131  , \P1_P3_InstQueue_reg[4][1]/NET0131  , \P1_P3_InstQueue_reg[4][2]/NET0131  , \P1_P3_InstQueue_reg[4][3]/NET0131  , \P1_P3_InstQueue_reg[4][4]/NET0131  , \P1_P3_InstQueue_reg[4][5]/NET0131  , \P1_P3_InstQueue_reg[4][6]/NET0131  , \P1_P3_InstQueue_reg[4][7]/NET0131  , \P1_P3_InstQueue_reg[5][0]/NET0131  , \P1_P3_InstQueue_reg[5][1]/NET0131  , \P1_P3_InstQueue_reg[5][2]/NET0131  , \P1_P3_InstQueue_reg[5][3]/NET0131  , \P1_P3_InstQueue_reg[5][4]/NET0131  , \P1_P3_InstQueue_reg[5][5]/NET0131  , \P1_P3_InstQueue_reg[5][6]/NET0131  , \P1_P3_InstQueue_reg[5][7]/NET0131  , \P1_P3_InstQueue_reg[6][0]/NET0131  , \P1_P3_InstQueue_reg[6][1]/NET0131  , \P1_P3_InstQueue_reg[6][2]/NET0131  , \P1_P3_InstQueue_reg[6][3]/NET0131  , \P1_P3_InstQueue_reg[6][4]/NET0131  , \P1_P3_InstQueue_reg[6][5]/NET0131  , \P1_P3_InstQueue_reg[6][6]/NET0131  , \P1_P3_InstQueue_reg[6][7]/NET0131  , \P1_P3_InstQueue_reg[7][0]/NET0131  , \P1_P3_InstQueue_reg[7][1]/NET0131  , \P1_P3_InstQueue_reg[7][2]/NET0131  , \P1_P3_InstQueue_reg[7][3]/NET0131  , \P1_P3_InstQueue_reg[7][4]/NET0131  , \P1_P3_InstQueue_reg[7][5]/NET0131  , \P1_P3_InstQueue_reg[7][6]/NET0131  , \P1_P3_InstQueue_reg[7][7]/NET0131  , \P1_P3_InstQueue_reg[8][0]/NET0131  , \P1_P3_InstQueue_reg[8][1]/NET0131  , \P1_P3_InstQueue_reg[8][2]/NET0131  , \P1_P3_InstQueue_reg[8][3]/NET0131  , \P1_P3_InstQueue_reg[8][4]/NET0131  , \P1_P3_InstQueue_reg[8][5]/NET0131  , \P1_P3_InstQueue_reg[8][6]/NET0131  , \P1_P3_InstQueue_reg[8][7]/NET0131  , \P1_P3_InstQueue_reg[9][0]/NET0131  , \P1_P3_InstQueue_reg[9][1]/NET0131  , \P1_P3_InstQueue_reg[9][2]/NET0131  , \P1_P3_InstQueue_reg[9][3]/NET0131  , \P1_P3_InstQueue_reg[9][4]/NET0131  , \P1_P3_InstQueue_reg[9][5]/NET0131  , \P1_P3_InstQueue_reg[9][6]/NET0131  , \P1_P3_InstQueue_reg[9][7]/NET0131  , \P1_P3_M_IO_n_reg/NET0131  , \P1_P3_MemoryFetch_reg/NET0131  , \P1_P3_More_reg/NET0131  , \P1_P3_PhyAddrPointer_reg[0]/NET0131  , \P1_P3_PhyAddrPointer_reg[10]/NET0131  , \P1_P3_PhyAddrPointer_reg[11]/NET0131  , \P1_P3_PhyAddrPointer_reg[12]/NET0131  , \P1_P3_PhyAddrPointer_reg[13]/NET0131  , \P1_P3_PhyAddrPointer_reg[14]/NET0131  , \P1_P3_PhyAddrPointer_reg[15]/NET0131  , \P1_P3_PhyAddrPointer_reg[16]/NET0131  , \P1_P3_PhyAddrPointer_reg[17]/NET0131  , \P1_P3_PhyAddrPointer_reg[18]/NET0131  , \P1_P3_PhyAddrPointer_reg[19]/NET0131  , \P1_P3_PhyAddrPointer_reg[1]/NET0131  , \P1_P3_PhyAddrPointer_reg[20]/NET0131  , \P1_P3_PhyAddrPointer_reg[21]/NET0131  , \P1_P3_PhyAddrPointer_reg[22]/NET0131  , \P1_P3_PhyAddrPointer_reg[23]/NET0131  , \P1_P3_PhyAddrPointer_reg[24]/NET0131  , \P1_P3_PhyAddrPointer_reg[25]/NET0131  , \P1_P3_PhyAddrPointer_reg[26]/NET0131  , \P1_P3_PhyAddrPointer_reg[27]/NET0131  , \P1_P3_PhyAddrPointer_reg[28]/NET0131  , \P1_P3_PhyAddrPointer_reg[29]/NET0131  , \P1_P3_PhyAddrPointer_reg[2]/NET0131  , \P1_P3_PhyAddrPointer_reg[30]/NET0131  , \P1_P3_PhyAddrPointer_reg[31]/NET0131  , \P1_P3_PhyAddrPointer_reg[3]/NET0131  , \P1_P3_PhyAddrPointer_reg[4]/NET0131  , \P1_P3_PhyAddrPointer_reg[5]/NET0131  , \P1_P3_PhyAddrPointer_reg[6]/NET0131  , \P1_P3_PhyAddrPointer_reg[7]/NET0131  , \P1_P3_PhyAddrPointer_reg[8]/NET0131  , \P1_P3_PhyAddrPointer_reg[9]/NET0131  , \P1_P3_ReadRequest_reg/NET0131  , \P1_P3_RequestPending_reg/NET0131  , \P1_P3_State2_reg[0]/NET0131  , \P1_P3_State2_reg[1]/NET0131  , \P1_P3_State2_reg[2]/NET0131  , \P1_P3_State2_reg[3]/NET0131  , \P1_P3_State_reg[0]/NET0131  , \P1_P3_State_reg[1]/NET0131  , \P1_P3_State_reg[2]/NET0131  , \P1_P3_W_R_n_reg/NET0131  , \P1_P3_rEIP_reg[0]/NET0131  , \P1_P3_rEIP_reg[10]/NET0131  , \P1_P3_rEIP_reg[11]/NET0131  , \P1_P3_rEIP_reg[12]/NET0131  , \P1_P3_rEIP_reg[13]/NET0131  , \P1_P3_rEIP_reg[14]/NET0131  , \P1_P3_rEIP_reg[15]/NET0131  , \P1_P3_rEIP_reg[16]/NET0131  , \P1_P3_rEIP_reg[17]/NET0131  , \P1_P3_rEIP_reg[18]/NET0131  , \P1_P3_rEIP_reg[19]/NET0131  , \P1_P3_rEIP_reg[1]/NET0131  , \P1_P3_rEIP_reg[20]/NET0131  , \P1_P3_rEIP_reg[21]/NET0131  , \P1_P3_rEIP_reg[22]/NET0131  , \P1_P3_rEIP_reg[23]/NET0131  , \P1_P3_rEIP_reg[24]/NET0131  , \P1_P3_rEIP_reg[25]/NET0131  , \P1_P3_rEIP_reg[26]/NET0131  , \P1_P3_rEIP_reg[27]/NET0131  , \P1_P3_rEIP_reg[28]/NET0131  , \P1_P3_rEIP_reg[29]/NET0131  , \P1_P3_rEIP_reg[2]/NET0131  , \P1_P3_rEIP_reg[30]/NET0131  , \P1_P3_rEIP_reg[31]/NET0131  , \P1_P3_rEIP_reg[3]/NET0131  , \P1_P3_rEIP_reg[4]/NET0131  , \P1_P3_rEIP_reg[5]/NET0131  , \P1_P3_rEIP_reg[6]/NET0131  , \P1_P3_rEIP_reg[7]/NET0131  , \P1_P3_rEIP_reg[8]/NET0131  , \P1_P3_rEIP_reg[9]/NET0131  , \P1_P3_uWord_reg[14]/NET0131  , \P1_buf1_reg[0]/NET0131  , \P1_buf1_reg[10]/NET0131  , \P1_buf1_reg[11]/NET0131  , \P1_buf1_reg[12]/NET0131  , \P1_buf1_reg[13]/NET0131  , \P1_buf1_reg[14]/NET0131  , \P1_buf1_reg[15]/NET0131  , \P1_buf1_reg[16]/NET0131  , \P1_buf1_reg[17]/NET0131  , \P1_buf1_reg[18]/NET0131  , \P1_buf1_reg[19]/NET0131  , \P1_buf1_reg[1]/NET0131  , \P1_buf1_reg[20]/NET0131  , \P1_buf1_reg[21]/NET0131  , \P1_buf1_reg[22]/NET0131  , \P1_buf1_reg[23]/NET0131  , \P1_buf1_reg[24]/NET0131  , \P1_buf1_reg[25]/NET0131  , \P1_buf1_reg[26]/NET0131  , \P1_buf1_reg[27]/NET0131  , \P1_buf1_reg[28]/NET0131  , \P1_buf1_reg[29]/NET0131  , \P1_buf1_reg[2]/NET0131  , \P1_buf1_reg[30]/NET0131  , \P1_buf1_reg[3]/NET0131  , \P1_buf1_reg[4]/NET0131  , \P1_buf1_reg[5]/NET0131  , \P1_buf1_reg[6]/NET0131  , \P1_buf1_reg[7]/NET0131  , \P1_buf1_reg[8]/NET0131  , \P1_buf1_reg[9]/NET0131  , \P1_buf2_reg[0]/NET0131  , \P1_buf2_reg[10]/NET0131  , \P1_buf2_reg[11]/NET0131  , \P1_buf2_reg[12]/NET0131  , \P1_buf2_reg[13]/NET0131  , \P1_buf2_reg[14]/NET0131  , \P1_buf2_reg[15]/NET0131  , \P1_buf2_reg[16]/NET0131  , \P1_buf2_reg[17]/NET0131  , \P1_buf2_reg[18]/NET0131  , \P1_buf2_reg[19]/NET0131  , \P1_buf2_reg[1]/NET0131  , \P1_buf2_reg[20]/NET0131  , \P1_buf2_reg[21]/NET0131  , \P1_buf2_reg[22]/NET0131  , \P1_buf2_reg[23]/NET0131  , \P1_buf2_reg[24]/NET0131  , \P1_buf2_reg[25]/NET0131  , \P1_buf2_reg[26]/NET0131  , \P1_buf2_reg[27]/NET0131  , \P1_buf2_reg[28]/NET0131  , \P1_buf2_reg[29]/NET0131  , \P1_buf2_reg[2]/NET0131  , \P1_buf2_reg[30]/NET0131  , \P1_buf2_reg[3]/NET0131  , \P1_buf2_reg[4]/NET0131  , \P1_buf2_reg[5]/NET0131  , \P1_buf2_reg[6]/NET0131  , \P1_buf2_reg[7]/NET0131  , \P1_buf2_reg[8]/NET0131  , \P1_buf2_reg[9]/NET0131  , \P1_ready11_reg/NET0131  , \P1_ready12_reg/NET0131  , \P1_ready21_reg/NET0131  , \P1_ready22_reg/NET0131  , \P2_P1_ADS_n_reg/NET0131  , \P2_P1_Address_reg[0]/NET0131  , \P2_P1_Address_reg[10]/NET0131  , \P2_P1_Address_reg[11]/NET0131  , \P2_P1_Address_reg[12]/NET0131  , \P2_P1_Address_reg[13]/NET0131  , \P2_P1_Address_reg[14]/NET0131  , \P2_P1_Address_reg[15]/NET0131  , \P2_P1_Address_reg[16]/NET0131  , \P2_P1_Address_reg[17]/NET0131  , \P2_P1_Address_reg[18]/NET0131  , \P2_P1_Address_reg[19]/NET0131  , \P2_P1_Address_reg[1]/NET0131  , \P2_P1_Address_reg[20]/NET0131  , \P2_P1_Address_reg[21]/NET0131  , \P2_P1_Address_reg[22]/NET0131  , \P2_P1_Address_reg[23]/NET0131  , \P2_P1_Address_reg[24]/NET0131  , \P2_P1_Address_reg[25]/NET0131  , \P2_P1_Address_reg[26]/NET0131  , \P2_P1_Address_reg[27]/NET0131  , \P2_P1_Address_reg[28]/NET0131  , \P2_P1_Address_reg[29]/NET0131  , \P2_P1_Address_reg[2]/NET0131  , \P2_P1_Address_reg[3]/NET0131  , \P2_P1_Address_reg[4]/NET0131  , \P2_P1_Address_reg[5]/NET0131  , \P2_P1_Address_reg[6]/NET0131  , \P2_P1_Address_reg[7]/NET0131  , \P2_P1_Address_reg[8]/NET0131  , \P2_P1_Address_reg[9]/NET0131  , \P2_P1_BE_n_reg[0]/NET0131  , \P2_P1_BE_n_reg[1]/NET0131  , \P2_P1_BE_n_reg[2]/NET0131  , \P2_P1_BE_n_reg[3]/NET0131  , \P2_P1_ByteEnable_reg[0]/NET0131  , \P2_P1_ByteEnable_reg[1]/NET0131  , \P2_P1_ByteEnable_reg[2]/NET0131  , \P2_P1_ByteEnable_reg[3]/NET0131  , \P2_P1_CodeFetch_reg/NET0131  , \P2_P1_D_C_n_reg/NET0131  , \P2_P1_DataWidth_reg[0]/NET0131  , \P2_P1_DataWidth_reg[1]/NET0131  , \P2_P1_Datao_reg[0]/NET0131  , \P2_P1_Datao_reg[10]/NET0131  , \P2_P1_Datao_reg[11]/NET0131  , \P2_P1_Datao_reg[12]/NET0131  , \P2_P1_Datao_reg[13]/NET0131  , \P2_P1_Datao_reg[14]/NET0131  , \P2_P1_Datao_reg[15]/NET0131  , \P2_P1_Datao_reg[16]/NET0131  , \P2_P1_Datao_reg[17]/NET0131  , \P2_P1_Datao_reg[18]/NET0131  , \P2_P1_Datao_reg[19]/NET0131  , \P2_P1_Datao_reg[1]/NET0131  , \P2_P1_Datao_reg[20]/NET0131  , \P2_P1_Datao_reg[21]/NET0131  , \P2_P1_Datao_reg[22]/NET0131  , \P2_P1_Datao_reg[23]/NET0131  , \P2_P1_Datao_reg[24]/NET0131  , \P2_P1_Datao_reg[25]/NET0131  , \P2_P1_Datao_reg[26]/NET0131  , \P2_P1_Datao_reg[27]/NET0131  , \P2_P1_Datao_reg[28]/NET0131  , \P2_P1_Datao_reg[29]/NET0131  , \P2_P1_Datao_reg[2]/NET0131  , \P2_P1_Datao_reg[30]/NET0131  , \P2_P1_Datao_reg[3]/NET0131  , \P2_P1_Datao_reg[4]/NET0131  , \P2_P1_Datao_reg[5]/NET0131  , \P2_P1_Datao_reg[6]/NET0131  , \P2_P1_Datao_reg[7]/NET0131  , \P2_P1_Datao_reg[8]/NET0131  , \P2_P1_Datao_reg[9]/NET0131  , \P2_P1_EAX_reg[0]/NET0131  , \P2_P1_EAX_reg[10]/NET0131  , \P2_P1_EAX_reg[11]/NET0131  , \P2_P1_EAX_reg[12]/NET0131  , \P2_P1_EAX_reg[13]/NET0131  , \P2_P1_EAX_reg[14]/NET0131  , \P2_P1_EAX_reg[15]/NET0131  , \P2_P1_EAX_reg[16]/NET0131  , \P2_P1_EAX_reg[17]/NET0131  , \P2_P1_EAX_reg[18]/NET0131  , \P2_P1_EAX_reg[19]/NET0131  , \P2_P1_EAX_reg[1]/NET0131  , \P2_P1_EAX_reg[20]/NET0131  , \P2_P1_EAX_reg[21]/NET0131  , \P2_P1_EAX_reg[22]/NET0131  , \P2_P1_EAX_reg[23]/NET0131  , \P2_P1_EAX_reg[24]/NET0131  , \P2_P1_EAX_reg[25]/NET0131  , \P2_P1_EAX_reg[26]/NET0131  , \P2_P1_EAX_reg[27]/NET0131  , \P2_P1_EAX_reg[28]/NET0131  , \P2_P1_EAX_reg[29]/NET0131  , \P2_P1_EAX_reg[2]/NET0131  , \P2_P1_EAX_reg[30]/NET0131  , \P2_P1_EAX_reg[31]/NET0131  , \P2_P1_EAX_reg[3]/NET0131  , \P2_P1_EAX_reg[4]/NET0131  , \P2_P1_EAX_reg[5]/NET0131  , \P2_P1_EAX_reg[6]/NET0131  , \P2_P1_EAX_reg[7]/NET0131  , \P2_P1_EAX_reg[8]/NET0131  , \P2_P1_EAX_reg[9]/NET0131  , \P2_P1_EBX_reg[0]/NET0131  , \P2_P1_EBX_reg[10]/NET0131  , \P2_P1_EBX_reg[11]/NET0131  , \P2_P1_EBX_reg[12]/NET0131  , \P2_P1_EBX_reg[13]/NET0131  , \P2_P1_EBX_reg[14]/NET0131  , \P2_P1_EBX_reg[15]/NET0131  , \P2_P1_EBX_reg[16]/NET0131  , \P2_P1_EBX_reg[17]/NET0131  , \P2_P1_EBX_reg[18]/NET0131  , \P2_P1_EBX_reg[19]/NET0131  , \P2_P1_EBX_reg[1]/NET0131  , \P2_P1_EBX_reg[20]/NET0131  , \P2_P1_EBX_reg[21]/NET0131  , \P2_P1_EBX_reg[22]/NET0131  , \P2_P1_EBX_reg[23]/NET0131  , \P2_P1_EBX_reg[24]/NET0131  , \P2_P1_EBX_reg[25]/NET0131  , \P2_P1_EBX_reg[26]/NET0131  , \P2_P1_EBX_reg[27]/NET0131  , \P2_P1_EBX_reg[28]/NET0131  , \P2_P1_EBX_reg[29]/NET0131  , \P2_P1_EBX_reg[2]/NET0131  , \P2_P1_EBX_reg[30]/NET0131  , \P2_P1_EBX_reg[31]/NET0131  , \P2_P1_EBX_reg[3]/NET0131  , \P2_P1_EBX_reg[4]/NET0131  , \P2_P1_EBX_reg[5]/NET0131  , \P2_P1_EBX_reg[6]/NET0131  , \P2_P1_EBX_reg[7]/NET0131  , \P2_P1_EBX_reg[8]/NET0131  , \P2_P1_EBX_reg[9]/NET0131  , \P2_P1_Flush_reg/NET0131  , \P2_P1_InstAddrPointer_reg[0]/NET0131  , \P2_P1_InstAddrPointer_reg[10]/NET0131  , \P2_P1_InstAddrPointer_reg[11]/NET0131  , \P2_P1_InstAddrPointer_reg[12]/NET0131  , \P2_P1_InstAddrPointer_reg[13]/NET0131  , \P2_P1_InstAddrPointer_reg[14]/NET0131  , \P2_P1_InstAddrPointer_reg[15]/NET0131  , \P2_P1_InstAddrPointer_reg[16]/NET0131  , \P2_P1_InstAddrPointer_reg[17]/NET0131  , \P2_P1_InstAddrPointer_reg[18]/NET0131  , \P2_P1_InstAddrPointer_reg[19]/NET0131  , \P2_P1_InstAddrPointer_reg[1]/NET0131  , \P2_P1_InstAddrPointer_reg[20]/NET0131  , \P2_P1_InstAddrPointer_reg[21]/NET0131  , \P2_P1_InstAddrPointer_reg[22]/NET0131  , \P2_P1_InstAddrPointer_reg[23]/NET0131  , \P2_P1_InstAddrPointer_reg[24]/NET0131  , \P2_P1_InstAddrPointer_reg[25]/NET0131  , \P2_P1_InstAddrPointer_reg[26]/NET0131  , \P2_P1_InstAddrPointer_reg[27]/NET0131  , \P2_P1_InstAddrPointer_reg[28]/NET0131  , \P2_P1_InstAddrPointer_reg[29]/NET0131  , \P2_P1_InstAddrPointer_reg[2]/NET0131  , \P2_P1_InstAddrPointer_reg[30]/NET0131  , \P2_P1_InstAddrPointer_reg[31]/NET0131  , \P2_P1_InstAddrPointer_reg[3]/NET0131  , \P2_P1_InstAddrPointer_reg[4]/NET0131  , \P2_P1_InstAddrPointer_reg[5]/NET0131  , \P2_P1_InstAddrPointer_reg[6]/NET0131  , \P2_P1_InstAddrPointer_reg[7]/NET0131  , \P2_P1_InstAddrPointer_reg[8]/NET0131  , \P2_P1_InstAddrPointer_reg[9]/NET0131  , \P2_P1_InstQueueRd_Addr_reg[0]/NET0131  , \P2_P1_InstQueueRd_Addr_reg[1]/NET0131  , \P2_P1_InstQueueRd_Addr_reg[2]/NET0131  , \P2_P1_InstQueueRd_Addr_reg[3]/NET0131  , \P2_P1_InstQueueWr_Addr_reg[0]/NET0131  , \P2_P1_InstQueueWr_Addr_reg[1]/NET0131  , \P2_P1_InstQueueWr_Addr_reg[2]/NET0131  , \P2_P1_InstQueueWr_Addr_reg[3]/NET0131  , \P2_P1_InstQueue_reg[0][0]/NET0131  , \P2_P1_InstQueue_reg[0][1]/NET0131  , \P2_P1_InstQueue_reg[0][2]/NET0131  , \P2_P1_InstQueue_reg[0][3]/NET0131  , \P2_P1_InstQueue_reg[0][4]/NET0131  , \P2_P1_InstQueue_reg[0][5]/NET0131  , \P2_P1_InstQueue_reg[0][6]/NET0131  , \P2_P1_InstQueue_reg[0][7]/NET0131  , \P2_P1_InstQueue_reg[10][0]/NET0131  , \P2_P1_InstQueue_reg[10][1]/NET0131  , \P2_P1_InstQueue_reg[10][2]/NET0131  , \P2_P1_InstQueue_reg[10][3]/NET0131  , \P2_P1_InstQueue_reg[10][4]/NET0131  , \P2_P1_InstQueue_reg[10][5]/NET0131  , \P2_P1_InstQueue_reg[10][6]/NET0131  , \P2_P1_InstQueue_reg[10][7]/NET0131  , \P2_P1_InstQueue_reg[11][0]/NET0131  , \P2_P1_InstQueue_reg[11][1]/NET0131  , \P2_P1_InstQueue_reg[11][2]/NET0131  , \P2_P1_InstQueue_reg[11][3]/NET0131  , \P2_P1_InstQueue_reg[11][4]/NET0131  , \P2_P1_InstQueue_reg[11][5]/NET0131  , \P2_P1_InstQueue_reg[11][6]/NET0131  , \P2_P1_InstQueue_reg[11][7]/NET0131  , \P2_P1_InstQueue_reg[12][0]/NET0131  , \P2_P1_InstQueue_reg[12][1]/NET0131  , \P2_P1_InstQueue_reg[12][2]/NET0131  , \P2_P1_InstQueue_reg[12][3]/NET0131  , \P2_P1_InstQueue_reg[12][4]/NET0131  , \P2_P1_InstQueue_reg[12][5]/NET0131  , \P2_P1_InstQueue_reg[12][6]/NET0131  , \P2_P1_InstQueue_reg[12][7]/NET0131  , \P2_P1_InstQueue_reg[13][0]/NET0131  , \P2_P1_InstQueue_reg[13][1]/NET0131  , \P2_P1_InstQueue_reg[13][2]/NET0131  , \P2_P1_InstQueue_reg[13][3]/NET0131  , \P2_P1_InstQueue_reg[13][4]/NET0131  , \P2_P1_InstQueue_reg[13][5]/NET0131  , \P2_P1_InstQueue_reg[13][6]/NET0131  , \P2_P1_InstQueue_reg[13][7]/NET0131  , \P2_P1_InstQueue_reg[14][0]/NET0131  , \P2_P1_InstQueue_reg[14][1]/NET0131  , \P2_P1_InstQueue_reg[14][2]/NET0131  , \P2_P1_InstQueue_reg[14][3]/NET0131  , \P2_P1_InstQueue_reg[14][4]/NET0131  , \P2_P1_InstQueue_reg[14][5]/NET0131  , \P2_P1_InstQueue_reg[14][6]/NET0131  , \P2_P1_InstQueue_reg[14][7]/NET0131  , \P2_P1_InstQueue_reg[15][0]/NET0131  , \P2_P1_InstQueue_reg[15][1]/NET0131  , \P2_P1_InstQueue_reg[15][2]/NET0131  , \P2_P1_InstQueue_reg[15][3]/NET0131  , \P2_P1_InstQueue_reg[15][4]/NET0131  , \P2_P1_InstQueue_reg[15][5]/NET0131  , \P2_P1_InstQueue_reg[15][6]/NET0131  , \P2_P1_InstQueue_reg[15][7]/NET0131  , \P2_P1_InstQueue_reg[1][0]/NET0131  , \P2_P1_InstQueue_reg[1][1]/NET0131  , \P2_P1_InstQueue_reg[1][2]/NET0131  , \P2_P1_InstQueue_reg[1][3]/NET0131  , \P2_P1_InstQueue_reg[1][4]/NET0131  , \P2_P1_InstQueue_reg[1][5]/NET0131  , \P2_P1_InstQueue_reg[1][6]/NET0131  , \P2_P1_InstQueue_reg[1][7]/NET0131  , \P2_P1_InstQueue_reg[2][0]/NET0131  , \P2_P1_InstQueue_reg[2][1]/NET0131  , \P2_P1_InstQueue_reg[2][2]/NET0131  , \P2_P1_InstQueue_reg[2][3]/NET0131  , \P2_P1_InstQueue_reg[2][4]/NET0131  , \P2_P1_InstQueue_reg[2][5]/NET0131  , \P2_P1_InstQueue_reg[2][6]/NET0131  , \P2_P1_InstQueue_reg[2][7]/NET0131  , \P2_P1_InstQueue_reg[3][0]/NET0131  , \P2_P1_InstQueue_reg[3][1]/NET0131  , \P2_P1_InstQueue_reg[3][2]/NET0131  , \P2_P1_InstQueue_reg[3][3]/NET0131  , \P2_P1_InstQueue_reg[3][4]/NET0131  , \P2_P1_InstQueue_reg[3][5]/NET0131  , \P2_P1_InstQueue_reg[3][6]/NET0131  , \P2_P1_InstQueue_reg[3][7]/NET0131  , \P2_P1_InstQueue_reg[4][0]/NET0131  , \P2_P1_InstQueue_reg[4][1]/NET0131  , \P2_P1_InstQueue_reg[4][2]/NET0131  , \P2_P1_InstQueue_reg[4][3]/NET0131  , \P2_P1_InstQueue_reg[4][4]/NET0131  , \P2_P1_InstQueue_reg[4][5]/NET0131  , \P2_P1_InstQueue_reg[4][6]/NET0131  , \P2_P1_InstQueue_reg[4][7]/NET0131  , \P2_P1_InstQueue_reg[5][0]/NET0131  , \P2_P1_InstQueue_reg[5][1]/NET0131  , \P2_P1_InstQueue_reg[5][2]/NET0131  , \P2_P1_InstQueue_reg[5][3]/NET0131  , \P2_P1_InstQueue_reg[5][4]/NET0131  , \P2_P1_InstQueue_reg[5][5]/NET0131  , \P2_P1_InstQueue_reg[5][6]/NET0131  , \P2_P1_InstQueue_reg[5][7]/NET0131  , \P2_P1_InstQueue_reg[6][0]/NET0131  , \P2_P1_InstQueue_reg[6][1]/NET0131  , \P2_P1_InstQueue_reg[6][2]/NET0131  , \P2_P1_InstQueue_reg[6][3]/NET0131  , \P2_P1_InstQueue_reg[6][4]/NET0131  , \P2_P1_InstQueue_reg[6][5]/NET0131  , \P2_P1_InstQueue_reg[6][6]/NET0131  , \P2_P1_InstQueue_reg[6][7]/NET0131  , \P2_P1_InstQueue_reg[7][0]/NET0131  , \P2_P1_InstQueue_reg[7][1]/NET0131  , \P2_P1_InstQueue_reg[7][2]/NET0131  , \P2_P1_InstQueue_reg[7][3]/NET0131  , \P2_P1_InstQueue_reg[7][4]/NET0131  , \P2_P1_InstQueue_reg[7][5]/NET0131  , \P2_P1_InstQueue_reg[7][6]/NET0131  , \P2_P1_InstQueue_reg[7][7]/NET0131  , \P2_P1_InstQueue_reg[8][0]/NET0131  , \P2_P1_InstQueue_reg[8][1]/NET0131  , \P2_P1_InstQueue_reg[8][2]/NET0131  , \P2_P1_InstQueue_reg[8][3]/NET0131  , \P2_P1_InstQueue_reg[8][4]/NET0131  , \P2_P1_InstQueue_reg[8][5]/NET0131  , \P2_P1_InstQueue_reg[8][6]/NET0131  , \P2_P1_InstQueue_reg[8][7]/NET0131  , \P2_P1_InstQueue_reg[9][0]/NET0131  , \P2_P1_InstQueue_reg[9][1]/NET0131  , \P2_P1_InstQueue_reg[9][2]/NET0131  , \P2_P1_InstQueue_reg[9][3]/NET0131  , \P2_P1_InstQueue_reg[9][4]/NET0131  , \P2_P1_InstQueue_reg[9][5]/NET0131  , \P2_P1_InstQueue_reg[9][6]/NET0131  , \P2_P1_InstQueue_reg[9][7]/NET0131  , \P2_P1_M_IO_n_reg/NET0131  , \P2_P1_MemoryFetch_reg/NET0131  , \P2_P1_More_reg/NET0131  , \P2_P1_PhyAddrPointer_reg[0]/NET0131  , \P2_P1_PhyAddrPointer_reg[10]/NET0131  , \P2_P1_PhyAddrPointer_reg[11]/NET0131  , \P2_P1_PhyAddrPointer_reg[12]/NET0131  , \P2_P1_PhyAddrPointer_reg[13]/NET0131  , \P2_P1_PhyAddrPointer_reg[14]/NET0131  , \P2_P1_PhyAddrPointer_reg[15]/NET0131  , \P2_P1_PhyAddrPointer_reg[16]/NET0131  , \P2_P1_PhyAddrPointer_reg[17]/NET0131  , \P2_P1_PhyAddrPointer_reg[18]/NET0131  , \P2_P1_PhyAddrPointer_reg[19]/NET0131  , \P2_P1_PhyAddrPointer_reg[1]/NET0131  , \P2_P1_PhyAddrPointer_reg[20]/NET0131  , \P2_P1_PhyAddrPointer_reg[21]/NET0131  , \P2_P1_PhyAddrPointer_reg[22]/NET0131  , \P2_P1_PhyAddrPointer_reg[23]/NET0131  , \P2_P1_PhyAddrPointer_reg[24]/NET0131  , \P2_P1_PhyAddrPointer_reg[25]/NET0131  , \P2_P1_PhyAddrPointer_reg[26]/NET0131  , \P2_P1_PhyAddrPointer_reg[27]/NET0131  , \P2_P1_PhyAddrPointer_reg[28]/NET0131  , \P2_P1_PhyAddrPointer_reg[29]/NET0131  , \P2_P1_PhyAddrPointer_reg[2]/NET0131  , \P2_P1_PhyAddrPointer_reg[30]/NET0131  , \P2_P1_PhyAddrPointer_reg[31]/NET0131  , \P2_P1_PhyAddrPointer_reg[3]/NET0131  , \P2_P1_PhyAddrPointer_reg[4]/NET0131  , \P2_P1_PhyAddrPointer_reg[5]/NET0131  , \P2_P1_PhyAddrPointer_reg[6]/NET0131  , \P2_P1_PhyAddrPointer_reg[7]/NET0131  , \P2_P1_PhyAddrPointer_reg[8]/NET0131  , \P2_P1_PhyAddrPointer_reg[9]/NET0131  , \P2_P1_ReadRequest_reg/NET0131  , \P2_P1_RequestPending_reg/NET0131  , \P2_P1_State2_reg[0]/NET0131  , \P2_P1_State2_reg[1]/NET0131  , \P2_P1_State2_reg[2]/NET0131  , \P2_P1_State2_reg[3]/NET0131  , \P2_P1_State_reg[0]/NET0131  , \P2_P1_State_reg[1]/NET0131  , \P2_P1_State_reg[2]/NET0131  , \P2_P1_W_R_n_reg/NET0131  , \P2_P1_lWord_reg[0]/NET0131  , \P2_P1_lWord_reg[10]/NET0131  , \P2_P1_lWord_reg[11]/NET0131  , \P2_P1_lWord_reg[12]/NET0131  , \P2_P1_lWord_reg[13]/NET0131  , \P2_P1_lWord_reg[14]/NET0131  , \P2_P1_lWord_reg[15]/NET0131  , \P2_P1_lWord_reg[1]/NET0131  , \P2_P1_lWord_reg[2]/NET0131  , \P2_P1_lWord_reg[3]/NET0131  , \P2_P1_lWord_reg[4]/NET0131  , \P2_P1_lWord_reg[5]/NET0131  , \P2_P1_lWord_reg[6]/NET0131  , \P2_P1_lWord_reg[7]/NET0131  , \P2_P1_lWord_reg[8]/NET0131  , \P2_P1_lWord_reg[9]/NET0131  , \P2_P1_rEIP_reg[0]/NET0131  , \P2_P1_rEIP_reg[10]/NET0131  , \P2_P1_rEIP_reg[11]/NET0131  , \P2_P1_rEIP_reg[12]/NET0131  , \P2_P1_rEIP_reg[13]/NET0131  , \P2_P1_rEIP_reg[14]/NET0131  , \P2_P1_rEIP_reg[15]/NET0131  , \P2_P1_rEIP_reg[16]/NET0131  , \P2_P1_rEIP_reg[17]/NET0131  , \P2_P1_rEIP_reg[18]/NET0131  , \P2_P1_rEIP_reg[19]/NET0131  , \P2_P1_rEIP_reg[1]/NET0131  , \P2_P1_rEIP_reg[20]/NET0131  , \P2_P1_rEIP_reg[21]/NET0131  , \P2_P1_rEIP_reg[22]/NET0131  , \P2_P1_rEIP_reg[23]/NET0131  , \P2_P1_rEIP_reg[24]/NET0131  , \P2_P1_rEIP_reg[25]/NET0131  , \P2_P1_rEIP_reg[26]/NET0131  , \P2_P1_rEIP_reg[27]/NET0131  , \P2_P1_rEIP_reg[28]/NET0131  , \P2_P1_rEIP_reg[29]/NET0131  , \P2_P1_rEIP_reg[2]/NET0131  , \P2_P1_rEIP_reg[30]/NET0131  , \P2_P1_rEIP_reg[31]/NET0131  , \P2_P1_rEIP_reg[3]/NET0131  , \P2_P1_rEIP_reg[4]/NET0131  , \P2_P1_rEIP_reg[5]/NET0131  , \P2_P1_rEIP_reg[6]/NET0131  , \P2_P1_rEIP_reg[7]/NET0131  , \P2_P1_rEIP_reg[8]/NET0131  , \P2_P1_rEIP_reg[9]/NET0131  , \P2_P1_uWord_reg[0]/NET0131  , \P2_P1_uWord_reg[10]/NET0131  , \P2_P1_uWord_reg[11]/NET0131  , \P2_P1_uWord_reg[12]/NET0131  , \P2_P1_uWord_reg[13]/NET0131  , \P2_P1_uWord_reg[14]/NET0131  , \P2_P1_uWord_reg[1]/NET0131  , \P2_P1_uWord_reg[2]/NET0131  , \P2_P1_uWord_reg[3]/NET0131  , \P2_P1_uWord_reg[4]/NET0131  , \P2_P1_uWord_reg[5]/NET0131  , \P2_P1_uWord_reg[6]/NET0131  , \P2_P1_uWord_reg[7]/NET0131  , \P2_P1_uWord_reg[8]/NET0131  , \P2_P1_uWord_reg[9]/NET0131  , \P2_P2_ADS_n_reg/NET0131  , \P2_P2_Address_reg[0]/NET0131  , \P2_P2_Address_reg[10]/NET0131  , \P2_P2_Address_reg[11]/NET0131  , \P2_P2_Address_reg[12]/NET0131  , \P2_P2_Address_reg[13]/NET0131  , \P2_P2_Address_reg[14]/NET0131  , \P2_P2_Address_reg[15]/NET0131  , \P2_P2_Address_reg[16]/NET0131  , \P2_P2_Address_reg[17]/NET0131  , \P2_P2_Address_reg[18]/NET0131  , \P2_P2_Address_reg[19]/NET0131  , \P2_P2_Address_reg[1]/NET0131  , \P2_P2_Address_reg[20]/NET0131  , \P2_P2_Address_reg[21]/NET0131  , \P2_P2_Address_reg[22]/NET0131  , \P2_P2_Address_reg[23]/NET0131  , \P2_P2_Address_reg[24]/NET0131  , \P2_P2_Address_reg[25]/NET0131  , \P2_P2_Address_reg[26]/NET0131  , \P2_P2_Address_reg[27]/NET0131  , \P2_P2_Address_reg[28]/NET0131  , \P2_P2_Address_reg[29]/NET0131  , \P2_P2_Address_reg[2]/NET0131  , \P2_P2_Address_reg[3]/NET0131  , \P2_P2_Address_reg[4]/NET0131  , \P2_P2_Address_reg[5]/NET0131  , \P2_P2_Address_reg[6]/NET0131  , \P2_P2_Address_reg[7]/NET0131  , \P2_P2_Address_reg[8]/NET0131  , \P2_P2_Address_reg[9]/NET0131  , \P2_P2_BE_n_reg[0]/NET0131  , \P2_P2_BE_n_reg[1]/NET0131  , \P2_P2_BE_n_reg[2]/NET0131  , \P2_P2_BE_n_reg[3]/NET0131  , \P2_P2_ByteEnable_reg[0]/NET0131  , \P2_P2_ByteEnable_reg[1]/NET0131  , \P2_P2_ByteEnable_reg[2]/NET0131  , \P2_P2_ByteEnable_reg[3]/NET0131  , \P2_P2_CodeFetch_reg/NET0131  , \P2_P2_D_C_n_reg/NET0131  , \P2_P2_DataWidth_reg[0]/NET0131  , \P2_P2_DataWidth_reg[1]/NET0131  , \P2_P2_Datao_reg[0]/NET0131  , \P2_P2_Datao_reg[10]/NET0131  , \P2_P2_Datao_reg[11]/NET0131  , \P2_P2_Datao_reg[12]/NET0131  , \P2_P2_Datao_reg[13]/NET0131  , \P2_P2_Datao_reg[14]/NET0131  , \P2_P2_Datao_reg[15]/NET0131  , \P2_P2_Datao_reg[16]/NET0131  , \P2_P2_Datao_reg[17]/NET0131  , \P2_P2_Datao_reg[18]/NET0131  , \P2_P2_Datao_reg[19]/NET0131  , \P2_P2_Datao_reg[1]/NET0131  , \P2_P2_Datao_reg[20]/NET0131  , \P2_P2_Datao_reg[21]/NET0131  , \P2_P2_Datao_reg[22]/NET0131  , \P2_P2_Datao_reg[23]/NET0131  , \P2_P2_Datao_reg[24]/NET0131  , \P2_P2_Datao_reg[25]/NET0131  , \P2_P2_Datao_reg[26]/NET0131  , \P2_P2_Datao_reg[27]/NET0131  , \P2_P2_Datao_reg[28]/NET0131  , \P2_P2_Datao_reg[29]/NET0131  , \P2_P2_Datao_reg[2]/NET0131  , \P2_P2_Datao_reg[30]/NET0131  , \P2_P2_Datao_reg[3]/NET0131  , \P2_P2_Datao_reg[4]/NET0131  , \P2_P2_Datao_reg[5]/NET0131  , \P2_P2_Datao_reg[6]/NET0131  , \P2_P2_Datao_reg[7]/NET0131  , \P2_P2_Datao_reg[8]/NET0131  , \P2_P2_Datao_reg[9]/NET0131  , \P2_P2_EAX_reg[0]/NET0131  , \P2_P2_EAX_reg[10]/NET0131  , \P2_P2_EAX_reg[11]/NET0131  , \P2_P2_EAX_reg[12]/NET0131  , \P2_P2_EAX_reg[13]/NET0131  , \P2_P2_EAX_reg[14]/NET0131  , \P2_P2_EAX_reg[15]/NET0131  , \P2_P2_EAX_reg[16]/NET0131  , \P2_P2_EAX_reg[17]/NET0131  , \P2_P2_EAX_reg[18]/NET0131  , \P2_P2_EAX_reg[19]/NET0131  , \P2_P2_EAX_reg[1]/NET0131  , \P2_P2_EAX_reg[20]/NET0131  , \P2_P2_EAX_reg[21]/NET0131  , \P2_P2_EAX_reg[22]/NET0131  , \P2_P2_EAX_reg[23]/NET0131  , \P2_P2_EAX_reg[24]/NET0131  , \P2_P2_EAX_reg[25]/NET0131  , \P2_P2_EAX_reg[26]/NET0131  , \P2_P2_EAX_reg[27]/NET0131  , \P2_P2_EAX_reg[28]/NET0131  , \P2_P2_EAX_reg[29]/NET0131  , \P2_P2_EAX_reg[2]/NET0131  , \P2_P2_EAX_reg[30]/NET0131  , \P2_P2_EAX_reg[31]/NET0131  , \P2_P2_EAX_reg[3]/NET0131  , \P2_P2_EAX_reg[4]/NET0131  , \P2_P2_EAX_reg[5]/NET0131  , \P2_P2_EAX_reg[6]/NET0131  , \P2_P2_EAX_reg[7]/NET0131  , \P2_P2_EAX_reg[8]/NET0131  , \P2_P2_EAX_reg[9]/NET0131  , \P2_P2_EBX_reg[0]/NET0131  , \P2_P2_EBX_reg[10]/NET0131  , \P2_P2_EBX_reg[11]/NET0131  , \P2_P2_EBX_reg[12]/NET0131  , \P2_P2_EBX_reg[13]/NET0131  , \P2_P2_EBX_reg[14]/NET0131  , \P2_P2_EBX_reg[15]/NET0131  , \P2_P2_EBX_reg[16]/NET0131  , \P2_P2_EBX_reg[17]/NET0131  , \P2_P2_EBX_reg[18]/NET0131  , \P2_P2_EBX_reg[19]/NET0131  , \P2_P2_EBX_reg[1]/NET0131  , \P2_P2_EBX_reg[20]/NET0131  , \P2_P2_EBX_reg[21]/NET0131  , \P2_P2_EBX_reg[22]/NET0131  , \P2_P2_EBX_reg[23]/NET0131  , \P2_P2_EBX_reg[24]/NET0131  , \P2_P2_EBX_reg[25]/NET0131  , \P2_P2_EBX_reg[26]/NET0131  , \P2_P2_EBX_reg[27]/NET0131  , \P2_P2_EBX_reg[28]/NET0131  , \P2_P2_EBX_reg[29]/NET0131  , \P2_P2_EBX_reg[2]/NET0131  , \P2_P2_EBX_reg[30]/NET0131  , \P2_P2_EBX_reg[31]/NET0131  , \P2_P2_EBX_reg[3]/NET0131  , \P2_P2_EBX_reg[4]/NET0131  , \P2_P2_EBX_reg[5]/NET0131  , \P2_P2_EBX_reg[6]/NET0131  , \P2_P2_EBX_reg[7]/NET0131  , \P2_P2_EBX_reg[8]/NET0131  , \P2_P2_EBX_reg[9]/NET0131  , \P2_P2_Flush_reg/NET0131  , \P2_P2_InstAddrPointer_reg[0]/NET0131  , \P2_P2_InstAddrPointer_reg[10]/NET0131  , \P2_P2_InstAddrPointer_reg[11]/NET0131  , \P2_P2_InstAddrPointer_reg[12]/NET0131  , \P2_P2_InstAddrPointer_reg[13]/NET0131  , \P2_P2_InstAddrPointer_reg[14]/NET0131  , \P2_P2_InstAddrPointer_reg[15]/NET0131  , \P2_P2_InstAddrPointer_reg[16]/NET0131  , \P2_P2_InstAddrPointer_reg[17]/NET0131  , \P2_P2_InstAddrPointer_reg[18]/NET0131  , \P2_P2_InstAddrPointer_reg[19]/NET0131  , \P2_P2_InstAddrPointer_reg[1]/NET0131  , \P2_P2_InstAddrPointer_reg[20]/NET0131  , \P2_P2_InstAddrPointer_reg[21]/NET0131  , \P2_P2_InstAddrPointer_reg[22]/NET0131  , \P2_P2_InstAddrPointer_reg[23]/NET0131  , \P2_P2_InstAddrPointer_reg[24]/NET0131  , \P2_P2_InstAddrPointer_reg[25]/NET0131  , \P2_P2_InstAddrPointer_reg[26]/NET0131  , \P2_P2_InstAddrPointer_reg[27]/NET0131  , \P2_P2_InstAddrPointer_reg[28]/NET0131  , \P2_P2_InstAddrPointer_reg[29]/NET0131  , \P2_P2_InstAddrPointer_reg[2]/NET0131  , \P2_P2_InstAddrPointer_reg[30]/NET0131  , \P2_P2_InstAddrPointer_reg[31]/NET0131  , \P2_P2_InstAddrPointer_reg[3]/NET0131  , \P2_P2_InstAddrPointer_reg[4]/NET0131  , \P2_P2_InstAddrPointer_reg[5]/NET0131  , \P2_P2_InstAddrPointer_reg[6]/NET0131  , \P2_P2_InstAddrPointer_reg[7]/NET0131  , \P2_P2_InstAddrPointer_reg[8]/NET0131  , \P2_P2_InstAddrPointer_reg[9]/NET0131  , \P2_P2_InstQueueRd_Addr_reg[0]/NET0131  , \P2_P2_InstQueueRd_Addr_reg[1]/NET0131  , \P2_P2_InstQueueRd_Addr_reg[2]/NET0131  , \P2_P2_InstQueueRd_Addr_reg[3]/NET0131  , \P2_P2_InstQueueWr_Addr_reg[0]/NET0131  , \P2_P2_InstQueueWr_Addr_reg[1]/NET0131  , \P2_P2_InstQueueWr_Addr_reg[2]/NET0131  , \P2_P2_InstQueueWr_Addr_reg[3]/NET0131  , \P2_P2_InstQueue_reg[0][0]/NET0131  , \P2_P2_InstQueue_reg[0][1]/NET0131  , \P2_P2_InstQueue_reg[0][2]/NET0131  , \P2_P2_InstQueue_reg[0][3]/NET0131  , \P2_P2_InstQueue_reg[0][4]/NET0131  , \P2_P2_InstQueue_reg[0][5]/NET0131  , \P2_P2_InstQueue_reg[0][6]/NET0131  , \P2_P2_InstQueue_reg[0][7]/NET0131  , \P2_P2_InstQueue_reg[10][0]/NET0131  , \P2_P2_InstQueue_reg[10][1]/NET0131  , \P2_P2_InstQueue_reg[10][2]/NET0131  , \P2_P2_InstQueue_reg[10][3]/NET0131  , \P2_P2_InstQueue_reg[10][4]/NET0131  , \P2_P2_InstQueue_reg[10][5]/NET0131  , \P2_P2_InstQueue_reg[10][6]/NET0131  , \P2_P2_InstQueue_reg[10][7]/NET0131  , \P2_P2_InstQueue_reg[11][0]/NET0131  , \P2_P2_InstQueue_reg[11][1]/NET0131  , \P2_P2_InstQueue_reg[11][2]/NET0131  , \P2_P2_InstQueue_reg[11][3]/NET0131  , \P2_P2_InstQueue_reg[11][4]/NET0131  , \P2_P2_InstQueue_reg[11][5]/NET0131  , \P2_P2_InstQueue_reg[11][6]/NET0131  , \P2_P2_InstQueue_reg[11][7]/NET0131  , \P2_P2_InstQueue_reg[12][0]/NET0131  , \P2_P2_InstQueue_reg[12][1]/NET0131  , \P2_P2_InstQueue_reg[12][2]/NET0131  , \P2_P2_InstQueue_reg[12][3]/NET0131  , \P2_P2_InstQueue_reg[12][4]/NET0131  , \P2_P2_InstQueue_reg[12][5]/NET0131  , \P2_P2_InstQueue_reg[12][6]/NET0131  , \P2_P2_InstQueue_reg[12][7]/NET0131  , \P2_P2_InstQueue_reg[13][0]/NET0131  , \P2_P2_InstQueue_reg[13][1]/NET0131  , \P2_P2_InstQueue_reg[13][2]/NET0131  , \P2_P2_InstQueue_reg[13][3]/NET0131  , \P2_P2_InstQueue_reg[13][4]/NET0131  , \P2_P2_InstQueue_reg[13][5]/NET0131  , \P2_P2_InstQueue_reg[13][6]/NET0131  , \P2_P2_InstQueue_reg[13][7]/NET0131  , \P2_P2_InstQueue_reg[14][0]/NET0131  , \P2_P2_InstQueue_reg[14][1]/NET0131  , \P2_P2_InstQueue_reg[14][2]/NET0131  , \P2_P2_InstQueue_reg[14][3]/NET0131  , \P2_P2_InstQueue_reg[14][4]/NET0131  , \P2_P2_InstQueue_reg[14][5]/NET0131  , \P2_P2_InstQueue_reg[14][6]/NET0131  , \P2_P2_InstQueue_reg[14][7]/NET0131  , \P2_P2_InstQueue_reg[15][0]/NET0131  , \P2_P2_InstQueue_reg[15][1]/NET0131  , \P2_P2_InstQueue_reg[15][2]/NET0131  , \P2_P2_InstQueue_reg[15][3]/NET0131  , \P2_P2_InstQueue_reg[15][4]/NET0131  , \P2_P2_InstQueue_reg[15][5]/NET0131  , \P2_P2_InstQueue_reg[15][6]/NET0131  , \P2_P2_InstQueue_reg[15][7]/NET0131  , \P2_P2_InstQueue_reg[1][0]/NET0131  , \P2_P2_InstQueue_reg[1][1]/NET0131  , \P2_P2_InstQueue_reg[1][2]/NET0131  , \P2_P2_InstQueue_reg[1][3]/NET0131  , \P2_P2_InstQueue_reg[1][4]/NET0131  , \P2_P2_InstQueue_reg[1][5]/NET0131  , \P2_P2_InstQueue_reg[1][6]/NET0131  , \P2_P2_InstQueue_reg[1][7]/NET0131  , \P2_P2_InstQueue_reg[2][0]/NET0131  , \P2_P2_InstQueue_reg[2][1]/NET0131  , \P2_P2_InstQueue_reg[2][2]/NET0131  , \P2_P2_InstQueue_reg[2][3]/NET0131  , \P2_P2_InstQueue_reg[2][4]/NET0131  , \P2_P2_InstQueue_reg[2][5]/NET0131  , \P2_P2_InstQueue_reg[2][6]/NET0131  , \P2_P2_InstQueue_reg[2][7]/NET0131  , \P2_P2_InstQueue_reg[3][0]/NET0131  , \P2_P2_InstQueue_reg[3][1]/NET0131  , \P2_P2_InstQueue_reg[3][2]/NET0131  , \P2_P2_InstQueue_reg[3][3]/NET0131  , \P2_P2_InstQueue_reg[3][4]/NET0131  , \P2_P2_InstQueue_reg[3][5]/NET0131  , \P2_P2_InstQueue_reg[3][6]/NET0131  , \P2_P2_InstQueue_reg[3][7]/NET0131  , \P2_P2_InstQueue_reg[4][0]/NET0131  , \P2_P2_InstQueue_reg[4][1]/NET0131  , \P2_P2_InstQueue_reg[4][2]/NET0131  , \P2_P2_InstQueue_reg[4][3]/NET0131  , \P2_P2_InstQueue_reg[4][4]/NET0131  , \P2_P2_InstQueue_reg[4][5]/NET0131  , \P2_P2_InstQueue_reg[4][6]/NET0131  , \P2_P2_InstQueue_reg[4][7]/NET0131  , \P2_P2_InstQueue_reg[5][0]/NET0131  , \P2_P2_InstQueue_reg[5][1]/NET0131  , \P2_P2_InstQueue_reg[5][2]/NET0131  , \P2_P2_InstQueue_reg[5][3]/NET0131  , \P2_P2_InstQueue_reg[5][4]/NET0131  , \P2_P2_InstQueue_reg[5][5]/NET0131  , \P2_P2_InstQueue_reg[5][6]/NET0131  , \P2_P2_InstQueue_reg[5][7]/NET0131  , \P2_P2_InstQueue_reg[6][0]/NET0131  , \P2_P2_InstQueue_reg[6][1]/NET0131  , \P2_P2_InstQueue_reg[6][2]/NET0131  , \P2_P2_InstQueue_reg[6][3]/NET0131  , \P2_P2_InstQueue_reg[6][4]/NET0131  , \P2_P2_InstQueue_reg[6][5]/NET0131  , \P2_P2_InstQueue_reg[6][6]/NET0131  , \P2_P2_InstQueue_reg[6][7]/NET0131  , \P2_P2_InstQueue_reg[7][0]/NET0131  , \P2_P2_InstQueue_reg[7][1]/NET0131  , \P2_P2_InstQueue_reg[7][2]/NET0131  , \P2_P2_InstQueue_reg[7][3]/NET0131  , \P2_P2_InstQueue_reg[7][4]/NET0131  , \P2_P2_InstQueue_reg[7][5]/NET0131  , \P2_P2_InstQueue_reg[7][6]/NET0131  , \P2_P2_InstQueue_reg[7][7]/NET0131  , \P2_P2_InstQueue_reg[8][0]/NET0131  , \P2_P2_InstQueue_reg[8][1]/NET0131  , \P2_P2_InstQueue_reg[8][2]/NET0131  , \P2_P2_InstQueue_reg[8][3]/NET0131  , \P2_P2_InstQueue_reg[8][4]/NET0131  , \P2_P2_InstQueue_reg[8][5]/NET0131  , \P2_P2_InstQueue_reg[8][6]/NET0131  , \P2_P2_InstQueue_reg[8][7]/NET0131  , \P2_P2_InstQueue_reg[9][0]/NET0131  , \P2_P2_InstQueue_reg[9][1]/NET0131  , \P2_P2_InstQueue_reg[9][2]/NET0131  , \P2_P2_InstQueue_reg[9][3]/NET0131  , \P2_P2_InstQueue_reg[9][4]/NET0131  , \P2_P2_InstQueue_reg[9][5]/NET0131  , \P2_P2_InstQueue_reg[9][6]/NET0131  , \P2_P2_InstQueue_reg[9][7]/NET0131  , \P2_P2_M_IO_n_reg/NET0131  , \P2_P2_MemoryFetch_reg/NET0131  , \P2_P2_More_reg/NET0131  , \P2_P2_PhyAddrPointer_reg[0]/NET0131  , \P2_P2_PhyAddrPointer_reg[10]/NET0131  , \P2_P2_PhyAddrPointer_reg[11]/NET0131  , \P2_P2_PhyAddrPointer_reg[12]/NET0131  , \P2_P2_PhyAddrPointer_reg[13]/NET0131  , \P2_P2_PhyAddrPointer_reg[14]/NET0131  , \P2_P2_PhyAddrPointer_reg[15]/NET0131  , \P2_P2_PhyAddrPointer_reg[16]/NET0131  , \P2_P2_PhyAddrPointer_reg[17]/NET0131  , \P2_P2_PhyAddrPointer_reg[18]/NET0131  , \P2_P2_PhyAddrPointer_reg[19]/NET0131  , \P2_P2_PhyAddrPointer_reg[1]/NET0131  , \P2_P2_PhyAddrPointer_reg[20]/NET0131  , \P2_P2_PhyAddrPointer_reg[21]/NET0131  , \P2_P2_PhyAddrPointer_reg[22]/NET0131  , \P2_P2_PhyAddrPointer_reg[23]/NET0131  , \P2_P2_PhyAddrPointer_reg[24]/NET0131  , \P2_P2_PhyAddrPointer_reg[25]/NET0131  , \P2_P2_PhyAddrPointer_reg[26]/NET0131  , \P2_P2_PhyAddrPointer_reg[27]/NET0131  , \P2_P2_PhyAddrPointer_reg[28]/NET0131  , \P2_P2_PhyAddrPointer_reg[29]/NET0131  , \P2_P2_PhyAddrPointer_reg[2]/NET0131  , \P2_P2_PhyAddrPointer_reg[30]/NET0131  , \P2_P2_PhyAddrPointer_reg[31]/NET0131  , \P2_P2_PhyAddrPointer_reg[3]/NET0131  , \P2_P2_PhyAddrPointer_reg[4]/NET0131  , \P2_P2_PhyAddrPointer_reg[5]/NET0131  , \P2_P2_PhyAddrPointer_reg[6]/NET0131  , \P2_P2_PhyAddrPointer_reg[7]/NET0131  , \P2_P2_PhyAddrPointer_reg[8]/NET0131  , \P2_P2_PhyAddrPointer_reg[9]/NET0131  , \P2_P2_ReadRequest_reg/NET0131  , \P2_P2_RequestPending_reg/NET0131  , \P2_P2_State2_reg[0]/NET0131  , \P2_P2_State2_reg[1]/NET0131  , \P2_P2_State2_reg[2]/NET0131  , \P2_P2_State2_reg[3]/NET0131  , \P2_P2_State_reg[0]/NET0131  , \P2_P2_State_reg[1]/NET0131  , \P2_P2_State_reg[2]/NET0131  , \P2_P2_W_R_n_reg/NET0131  , \P2_P2_lWord_reg[0]/NET0131  , \P2_P2_lWord_reg[10]/NET0131  , \P2_P2_lWord_reg[11]/NET0131  , \P2_P2_lWord_reg[12]/NET0131  , \P2_P2_lWord_reg[13]/NET0131  , \P2_P2_lWord_reg[14]/NET0131  , \P2_P2_lWord_reg[15]/NET0131  , \P2_P2_lWord_reg[1]/NET0131  , \P2_P2_lWord_reg[2]/NET0131  , \P2_P2_lWord_reg[3]/NET0131  , \P2_P2_lWord_reg[4]/NET0131  , \P2_P2_lWord_reg[5]/NET0131  , \P2_P2_lWord_reg[6]/NET0131  , \P2_P2_lWord_reg[7]/NET0131  , \P2_P2_lWord_reg[8]/NET0131  , \P2_P2_lWord_reg[9]/NET0131  , \P2_P2_rEIP_reg[0]/NET0131  , \P2_P2_rEIP_reg[10]/NET0131  , \P2_P2_rEIP_reg[11]/NET0131  , \P2_P2_rEIP_reg[12]/NET0131  , \P2_P2_rEIP_reg[13]/NET0131  , \P2_P2_rEIP_reg[14]/NET0131  , \P2_P2_rEIP_reg[15]/NET0131  , \P2_P2_rEIP_reg[16]/NET0131  , \P2_P2_rEIP_reg[17]/NET0131  , \P2_P2_rEIP_reg[18]/NET0131  , \P2_P2_rEIP_reg[19]/NET0131  , \P2_P2_rEIP_reg[1]/NET0131  , \P2_P2_rEIP_reg[20]/NET0131  , \P2_P2_rEIP_reg[21]/NET0131  , \P2_P2_rEIP_reg[22]/NET0131  , \P2_P2_rEIP_reg[23]/NET0131  , \P2_P2_rEIP_reg[24]/NET0131  , \P2_P2_rEIP_reg[25]/NET0131  , \P2_P2_rEIP_reg[26]/NET0131  , \P2_P2_rEIP_reg[27]/NET0131  , \P2_P2_rEIP_reg[28]/NET0131  , \P2_P2_rEIP_reg[29]/NET0131  , \P2_P2_rEIP_reg[2]/NET0131  , \P2_P2_rEIP_reg[30]/NET0131  , \P2_P2_rEIP_reg[31]/NET0131  , \P2_P2_rEIP_reg[3]/NET0131  , \P2_P2_rEIP_reg[4]/NET0131  , \P2_P2_rEIP_reg[5]/NET0131  , \P2_P2_rEIP_reg[6]/NET0131  , \P2_P2_rEIP_reg[7]/NET0131  , \P2_P2_rEIP_reg[8]/NET0131  , \P2_P2_rEIP_reg[9]/NET0131  , \P2_P2_uWord_reg[0]/NET0131  , \P2_P2_uWord_reg[10]/NET0131  , \P2_P2_uWord_reg[11]/NET0131  , \P2_P2_uWord_reg[12]/NET0131  , \P2_P2_uWord_reg[13]/NET0131  , \P2_P2_uWord_reg[14]/NET0131  , \P2_P2_uWord_reg[1]/NET0131  , \P2_P2_uWord_reg[2]/NET0131  , \P2_P2_uWord_reg[3]/NET0131  , \P2_P2_uWord_reg[4]/NET0131  , \P2_P2_uWord_reg[5]/NET0131  , \P2_P2_uWord_reg[6]/NET0131  , \P2_P2_uWord_reg[7]/NET0131  , \P2_P2_uWord_reg[8]/NET0131  , \P2_P2_uWord_reg[9]/NET0131  , \P2_P3_ADS_n_reg/NET0131  , \P2_P3_Address_reg[0]/NET0131  , \P2_P3_Address_reg[10]/NET0131  , \P2_P3_Address_reg[11]/NET0131  , \P2_P3_Address_reg[12]/NET0131  , \P2_P3_Address_reg[13]/NET0131  , \P2_P3_Address_reg[14]/NET0131  , \P2_P3_Address_reg[15]/NET0131  , \P2_P3_Address_reg[16]/NET0131  , \P2_P3_Address_reg[17]/NET0131  , \P2_P3_Address_reg[18]/NET0131  , \P2_P3_Address_reg[1]/NET0131  , \P2_P3_Address_reg[2]/NET0131  , \P2_P3_Address_reg[3]/NET0131  , \P2_P3_Address_reg[4]/NET0131  , \P2_P3_Address_reg[5]/NET0131  , \P2_P3_Address_reg[6]/NET0131  , \P2_P3_Address_reg[7]/NET0131  , \P2_P3_Address_reg[8]/NET0131  , \P2_P3_Address_reg[9]/NET0131  , \P2_P3_BE_n_reg[0]/NET0131  , \P2_P3_BE_n_reg[1]/NET0131  , \P2_P3_BE_n_reg[2]/NET0131  , \P2_P3_BE_n_reg[3]/NET0131  , \P2_P3_ByteEnable_reg[0]/NET0131  , \P2_P3_ByteEnable_reg[1]/NET0131  , \P2_P3_ByteEnable_reg[2]/NET0131  , \P2_P3_ByteEnable_reg[3]/NET0131  , \P2_P3_CodeFetch_reg/NET0131  , \P2_P3_D_C_n_reg/NET0131  , \P2_P3_DataWidth_reg[0]/NET0131  , \P2_P3_DataWidth_reg[1]/NET0131  , \P2_P3_Datao_reg[0]/NET0131  , \P2_P3_Datao_reg[10]/NET0131  , \P2_P3_Datao_reg[11]/NET0131  , \P2_P3_Datao_reg[12]/NET0131  , \P2_P3_Datao_reg[13]/NET0131  , \P2_P3_Datao_reg[14]/NET0131  , \P2_P3_Datao_reg[15]/NET0131  , \P2_P3_Datao_reg[16]/NET0131  , \P2_P3_Datao_reg[17]/NET0131  , \P2_P3_Datao_reg[18]/NET0131  , \P2_P3_Datao_reg[19]/NET0131  , \P2_P3_Datao_reg[1]/NET0131  , \P2_P3_Datao_reg[20]/NET0131  , \P2_P3_Datao_reg[21]/NET0131  , \P2_P3_Datao_reg[22]/NET0131  , \P2_P3_Datao_reg[23]/NET0131  , \P2_P3_Datao_reg[24]/NET0131  , \P2_P3_Datao_reg[25]/NET0131  , \P2_P3_Datao_reg[26]/NET0131  , \P2_P3_Datao_reg[27]/NET0131  , \P2_P3_Datao_reg[28]/NET0131  , \P2_P3_Datao_reg[29]/NET0131  , \P2_P3_Datao_reg[2]/NET0131  , \P2_P3_Datao_reg[30]/NET0131  , \P2_P3_Datao_reg[3]/NET0131  , \P2_P3_Datao_reg[4]/NET0131  , \P2_P3_Datao_reg[5]/NET0131  , \P2_P3_Datao_reg[6]/NET0131  , \P2_P3_Datao_reg[7]/NET0131  , \P2_P3_Datao_reg[8]/NET0131  , \P2_P3_Datao_reg[9]/NET0131  , \P2_P3_EAX_reg[0]/NET0131  , \P2_P3_EAX_reg[10]/NET0131  , \P2_P3_EAX_reg[11]/NET0131  , \P2_P3_EAX_reg[12]/NET0131  , \P2_P3_EAX_reg[13]/NET0131  , \P2_P3_EAX_reg[14]/NET0131  , \P2_P3_EAX_reg[15]/NET0131  , \P2_P3_EAX_reg[16]/NET0131  , \P2_P3_EAX_reg[17]/NET0131  , \P2_P3_EAX_reg[18]/NET0131  , \P2_P3_EAX_reg[19]/NET0131  , \P2_P3_EAX_reg[1]/NET0131  , \P2_P3_EAX_reg[20]/NET0131  , \P2_P3_EAX_reg[21]/NET0131  , \P2_P3_EAX_reg[22]/NET0131  , \P2_P3_EAX_reg[23]/NET0131  , \P2_P3_EAX_reg[24]/NET0131  , \P2_P3_EAX_reg[25]/NET0131  , \P2_P3_EAX_reg[26]/NET0131  , \P2_P3_EAX_reg[27]/NET0131  , \P2_P3_EAX_reg[28]/NET0131  , \P2_P3_EAX_reg[29]/NET0131  , \P2_P3_EAX_reg[2]/NET0131  , \P2_P3_EAX_reg[30]/NET0131  , \P2_P3_EAX_reg[31]/NET0131  , \P2_P3_EAX_reg[3]/NET0131  , \P2_P3_EAX_reg[4]/NET0131  , \P2_P3_EAX_reg[5]/NET0131  , \P2_P3_EAX_reg[6]/NET0131  , \P2_P3_EAX_reg[7]/NET0131  , \P2_P3_EAX_reg[8]/NET0131  , \P2_P3_EAX_reg[9]/NET0131  , \P2_P3_EBX_reg[0]/NET0131  , \P2_P3_EBX_reg[10]/NET0131  , \P2_P3_EBX_reg[11]/NET0131  , \P2_P3_EBX_reg[12]/NET0131  , \P2_P3_EBX_reg[13]/NET0131  , \P2_P3_EBX_reg[14]/NET0131  , \P2_P3_EBX_reg[15]/NET0131  , \P2_P3_EBX_reg[16]/NET0131  , \P2_P3_EBX_reg[17]/NET0131  , \P2_P3_EBX_reg[18]/NET0131  , \P2_P3_EBX_reg[19]/NET0131  , \P2_P3_EBX_reg[1]/NET0131  , \P2_P3_EBX_reg[20]/NET0131  , \P2_P3_EBX_reg[21]/NET0131  , \P2_P3_EBX_reg[22]/NET0131  , \P2_P3_EBX_reg[23]/NET0131  , \P2_P3_EBX_reg[24]/NET0131  , \P2_P3_EBX_reg[25]/NET0131  , \P2_P3_EBX_reg[26]/NET0131  , \P2_P3_EBX_reg[27]/NET0131  , \P2_P3_EBX_reg[28]/NET0131  , \P2_P3_EBX_reg[29]/NET0131  , \P2_P3_EBX_reg[2]/NET0131  , \P2_P3_EBX_reg[30]/NET0131  , \P2_P3_EBX_reg[31]/NET0131  , \P2_P3_EBX_reg[3]/NET0131  , \P2_P3_EBX_reg[4]/NET0131  , \P2_P3_EBX_reg[5]/NET0131  , \P2_P3_EBX_reg[6]/NET0131  , \P2_P3_EBX_reg[7]/NET0131  , \P2_P3_EBX_reg[8]/NET0131  , \P2_P3_EBX_reg[9]/NET0131  , \P2_P3_Flush_reg/NET0131  , \P2_P3_InstAddrPointer_reg[0]/NET0131  , \P2_P3_InstAddrPointer_reg[10]/NET0131  , \P2_P3_InstAddrPointer_reg[11]/NET0131  , \P2_P3_InstAddrPointer_reg[12]/NET0131  , \P2_P3_InstAddrPointer_reg[13]/NET0131  , \P2_P3_InstAddrPointer_reg[14]/NET0131  , \P2_P3_InstAddrPointer_reg[15]/NET0131  , \P2_P3_InstAddrPointer_reg[16]/NET0131  , \P2_P3_InstAddrPointer_reg[17]/NET0131  , \P2_P3_InstAddrPointer_reg[18]/NET0131  , \P2_P3_InstAddrPointer_reg[19]/NET0131  , \P2_P3_InstAddrPointer_reg[1]/NET0131  , \P2_P3_InstAddrPointer_reg[20]/NET0131  , \P2_P3_InstAddrPointer_reg[21]/NET0131  , \P2_P3_InstAddrPointer_reg[22]/NET0131  , \P2_P3_InstAddrPointer_reg[23]/NET0131  , \P2_P3_InstAddrPointer_reg[24]/NET0131  , \P2_P3_InstAddrPointer_reg[25]/NET0131  , \P2_P3_InstAddrPointer_reg[26]/NET0131  , \P2_P3_InstAddrPointer_reg[27]/NET0131  , \P2_P3_InstAddrPointer_reg[28]/NET0131  , \P2_P3_InstAddrPointer_reg[29]/NET0131  , \P2_P3_InstAddrPointer_reg[2]/NET0131  , \P2_P3_InstAddrPointer_reg[30]/NET0131  , \P2_P3_InstAddrPointer_reg[31]/NET0131  , \P2_P3_InstAddrPointer_reg[3]/NET0131  , \P2_P3_InstAddrPointer_reg[4]/NET0131  , \P2_P3_InstAddrPointer_reg[5]/NET0131  , \P2_P3_InstAddrPointer_reg[6]/NET0131  , \P2_P3_InstAddrPointer_reg[7]/NET0131  , \P2_P3_InstAddrPointer_reg[8]/NET0131  , \P2_P3_InstAddrPointer_reg[9]/NET0131  , \P2_P3_InstQueueRd_Addr_reg[0]/NET0131  , \P2_P3_InstQueueRd_Addr_reg[1]/NET0131  , \P2_P3_InstQueueRd_Addr_reg[2]/NET0131  , \P2_P3_InstQueueRd_Addr_reg[3]/NET0131  , \P2_P3_InstQueueWr_Addr_reg[0]/NET0131  , \P2_P3_InstQueueWr_Addr_reg[1]/NET0131  , \P2_P3_InstQueueWr_Addr_reg[2]/NET0131  , \P2_P3_InstQueueWr_Addr_reg[3]/NET0131  , \P2_P3_InstQueue_reg[0][0]/NET0131  , \P2_P3_InstQueue_reg[0][1]/NET0131  , \P2_P3_InstQueue_reg[0][2]/NET0131  , \P2_P3_InstQueue_reg[0][3]/NET0131  , \P2_P3_InstQueue_reg[0][4]/NET0131  , \P2_P3_InstQueue_reg[0][5]/NET0131  , \P2_P3_InstQueue_reg[0][6]/NET0131  , \P2_P3_InstQueue_reg[0][7]/NET0131  , \P2_P3_InstQueue_reg[10][0]/NET0131  , \P2_P3_InstQueue_reg[10][1]/NET0131  , \P2_P3_InstQueue_reg[10][2]/NET0131  , \P2_P3_InstQueue_reg[10][3]/NET0131  , \P2_P3_InstQueue_reg[10][4]/NET0131  , \P2_P3_InstQueue_reg[10][5]/NET0131  , \P2_P3_InstQueue_reg[10][6]/NET0131  , \P2_P3_InstQueue_reg[10][7]/NET0131  , \P2_P3_InstQueue_reg[11][0]/NET0131  , \P2_P3_InstQueue_reg[11][1]/NET0131  , \P2_P3_InstQueue_reg[11][2]/NET0131  , \P2_P3_InstQueue_reg[11][3]/NET0131  , \P2_P3_InstQueue_reg[11][4]/NET0131  , \P2_P3_InstQueue_reg[11][5]/NET0131  , \P2_P3_InstQueue_reg[11][6]/NET0131  , \P2_P3_InstQueue_reg[11][7]/NET0131  , \P2_P3_InstQueue_reg[12][0]/NET0131  , \P2_P3_InstQueue_reg[12][1]/NET0131  , \P2_P3_InstQueue_reg[12][2]/NET0131  , \P2_P3_InstQueue_reg[12][3]/NET0131  , \P2_P3_InstQueue_reg[12][4]/NET0131  , \P2_P3_InstQueue_reg[12][5]/NET0131  , \P2_P3_InstQueue_reg[12][6]/NET0131  , \P2_P3_InstQueue_reg[12][7]/NET0131  , \P2_P3_InstQueue_reg[13][0]/NET0131  , \P2_P3_InstQueue_reg[13][1]/NET0131  , \P2_P3_InstQueue_reg[13][2]/NET0131  , \P2_P3_InstQueue_reg[13][3]/NET0131  , \P2_P3_InstQueue_reg[13][4]/NET0131  , \P2_P3_InstQueue_reg[13][5]/NET0131  , \P2_P3_InstQueue_reg[13][6]/NET0131  , \P2_P3_InstQueue_reg[13][7]/NET0131  , \P2_P3_InstQueue_reg[14][0]/NET0131  , \P2_P3_InstQueue_reg[14][1]/NET0131  , \P2_P3_InstQueue_reg[14][2]/NET0131  , \P2_P3_InstQueue_reg[14][3]/NET0131  , \P2_P3_InstQueue_reg[14][4]/NET0131  , \P2_P3_InstQueue_reg[14][5]/NET0131  , \P2_P3_InstQueue_reg[14][6]/NET0131  , \P2_P3_InstQueue_reg[14][7]/NET0131  , \P2_P3_InstQueue_reg[15][0]/NET0131  , \P2_P3_InstQueue_reg[15][1]/NET0131  , \P2_P3_InstQueue_reg[15][2]/NET0131  , \P2_P3_InstQueue_reg[15][3]/NET0131  , \P2_P3_InstQueue_reg[15][4]/NET0131  , \P2_P3_InstQueue_reg[15][5]/NET0131  , \P2_P3_InstQueue_reg[15][6]/NET0131  , \P2_P3_InstQueue_reg[15][7]/NET0131  , \P2_P3_InstQueue_reg[1][0]/NET0131  , \P2_P3_InstQueue_reg[1][1]/NET0131  , \P2_P3_InstQueue_reg[1][2]/NET0131  , \P2_P3_InstQueue_reg[1][3]/NET0131  , \P2_P3_InstQueue_reg[1][4]/NET0131  , \P2_P3_InstQueue_reg[1][5]/NET0131  , \P2_P3_InstQueue_reg[1][6]/NET0131  , \P2_P3_InstQueue_reg[1][7]/NET0131  , \P2_P3_InstQueue_reg[2][0]/NET0131  , \P2_P3_InstQueue_reg[2][1]/NET0131  , \P2_P3_InstQueue_reg[2][2]/NET0131  , \P2_P3_InstQueue_reg[2][3]/NET0131  , \P2_P3_InstQueue_reg[2][4]/NET0131  , \P2_P3_InstQueue_reg[2][5]/NET0131  , \P2_P3_InstQueue_reg[2][6]/NET0131  , \P2_P3_InstQueue_reg[2][7]/NET0131  , \P2_P3_InstQueue_reg[3][0]/NET0131  , \P2_P3_InstQueue_reg[3][1]/NET0131  , \P2_P3_InstQueue_reg[3][2]/NET0131  , \P2_P3_InstQueue_reg[3][3]/NET0131  , \P2_P3_InstQueue_reg[3][4]/NET0131  , \P2_P3_InstQueue_reg[3][5]/NET0131  , \P2_P3_InstQueue_reg[3][6]/NET0131  , \P2_P3_InstQueue_reg[3][7]/NET0131  , \P2_P3_InstQueue_reg[4][0]/NET0131  , \P2_P3_InstQueue_reg[4][1]/NET0131  , \P2_P3_InstQueue_reg[4][2]/NET0131  , \P2_P3_InstQueue_reg[4][3]/NET0131  , \P2_P3_InstQueue_reg[4][4]/NET0131  , \P2_P3_InstQueue_reg[4][5]/NET0131  , \P2_P3_InstQueue_reg[4][6]/NET0131  , \P2_P3_InstQueue_reg[4][7]/NET0131  , \P2_P3_InstQueue_reg[5][0]/NET0131  , \P2_P3_InstQueue_reg[5][1]/NET0131  , \P2_P3_InstQueue_reg[5][2]/NET0131  , \P2_P3_InstQueue_reg[5][3]/NET0131  , \P2_P3_InstQueue_reg[5][4]/NET0131  , \P2_P3_InstQueue_reg[5][5]/NET0131  , \P2_P3_InstQueue_reg[5][6]/NET0131  , \P2_P3_InstQueue_reg[5][7]/NET0131  , \P2_P3_InstQueue_reg[6][0]/NET0131  , \P2_P3_InstQueue_reg[6][1]/NET0131  , \P2_P3_InstQueue_reg[6][2]/NET0131  , \P2_P3_InstQueue_reg[6][3]/NET0131  , \P2_P3_InstQueue_reg[6][4]/NET0131  , \P2_P3_InstQueue_reg[6][5]/NET0131  , \P2_P3_InstQueue_reg[6][6]/NET0131  , \P2_P3_InstQueue_reg[6][7]/NET0131  , \P2_P3_InstQueue_reg[7][0]/NET0131  , \P2_P3_InstQueue_reg[7][1]/NET0131  , \P2_P3_InstQueue_reg[7][2]/NET0131  , \P2_P3_InstQueue_reg[7][3]/NET0131  , \P2_P3_InstQueue_reg[7][4]/NET0131  , \P2_P3_InstQueue_reg[7][5]/NET0131  , \P2_P3_InstQueue_reg[7][6]/NET0131  , \P2_P3_InstQueue_reg[7][7]/NET0131  , \P2_P3_InstQueue_reg[8][0]/NET0131  , \P2_P3_InstQueue_reg[8][1]/NET0131  , \P2_P3_InstQueue_reg[8][2]/NET0131  , \P2_P3_InstQueue_reg[8][3]/NET0131  , \P2_P3_InstQueue_reg[8][4]/NET0131  , \P2_P3_InstQueue_reg[8][5]/NET0131  , \P2_P3_InstQueue_reg[8][6]/NET0131  , \P2_P3_InstQueue_reg[8][7]/NET0131  , \P2_P3_InstQueue_reg[9][0]/NET0131  , \P2_P3_InstQueue_reg[9][1]/NET0131  , \P2_P3_InstQueue_reg[9][2]/NET0131  , \P2_P3_InstQueue_reg[9][3]/NET0131  , \P2_P3_InstQueue_reg[9][4]/NET0131  , \P2_P3_InstQueue_reg[9][5]/NET0131  , \P2_P3_InstQueue_reg[9][6]/NET0131  , \P2_P3_InstQueue_reg[9][7]/NET0131  , \P2_P3_M_IO_n_reg/NET0131  , \P2_P3_MemoryFetch_reg/NET0131  , \P2_P3_More_reg/NET0131  , \P2_P3_PhyAddrPointer_reg[0]/NET0131  , \P2_P3_PhyAddrPointer_reg[10]/NET0131  , \P2_P3_PhyAddrPointer_reg[11]/NET0131  , \P2_P3_PhyAddrPointer_reg[12]/NET0131  , \P2_P3_PhyAddrPointer_reg[13]/NET0131  , \P2_P3_PhyAddrPointer_reg[14]/NET0131  , \P2_P3_PhyAddrPointer_reg[15]/NET0131  , \P2_P3_PhyAddrPointer_reg[16]/NET0131  , \P2_P3_PhyAddrPointer_reg[17]/NET0131  , \P2_P3_PhyAddrPointer_reg[18]/NET0131  , \P2_P3_PhyAddrPointer_reg[19]/NET0131  , \P2_P3_PhyAddrPointer_reg[1]/NET0131  , \P2_P3_PhyAddrPointer_reg[20]/NET0131  , \P2_P3_PhyAddrPointer_reg[21]/NET0131  , \P2_P3_PhyAddrPointer_reg[22]/NET0131  , \P2_P3_PhyAddrPointer_reg[23]/NET0131  , \P2_P3_PhyAddrPointer_reg[24]/NET0131  , \P2_P3_PhyAddrPointer_reg[25]/NET0131  , \P2_P3_PhyAddrPointer_reg[26]/NET0131  , \P2_P3_PhyAddrPointer_reg[27]/NET0131  , \P2_P3_PhyAddrPointer_reg[28]/NET0131  , \P2_P3_PhyAddrPointer_reg[29]/NET0131  , \P2_P3_PhyAddrPointer_reg[2]/NET0131  , \P2_P3_PhyAddrPointer_reg[30]/NET0131  , \P2_P3_PhyAddrPointer_reg[31]/NET0131  , \P2_P3_PhyAddrPointer_reg[3]/NET0131  , \P2_P3_PhyAddrPointer_reg[4]/NET0131  , \P2_P3_PhyAddrPointer_reg[5]/NET0131  , \P2_P3_PhyAddrPointer_reg[6]/NET0131  , \P2_P3_PhyAddrPointer_reg[7]/NET0131  , \P2_P3_PhyAddrPointer_reg[8]/NET0131  , \P2_P3_PhyAddrPointer_reg[9]/NET0131  , \P2_P3_ReadRequest_reg/NET0131  , \P2_P3_RequestPending_reg/NET0131  , \P2_P3_State2_reg[0]/NET0131  , \P2_P3_State2_reg[1]/NET0131  , \P2_P3_State2_reg[2]/NET0131  , \P2_P3_State2_reg[3]/NET0131  , \P2_P3_State_reg[0]/NET0131  , \P2_P3_State_reg[1]/NET0131  , \P2_P3_State_reg[2]/NET0131  , \P2_P3_W_R_n_reg/NET0131  , \P2_P3_lWord_reg[0]/NET0131  , \P2_P3_lWord_reg[10]/NET0131  , \P2_P3_lWord_reg[11]/NET0131  , \P2_P3_lWord_reg[12]/NET0131  , \P2_P3_lWord_reg[13]/NET0131  , \P2_P3_lWord_reg[14]/NET0131  , \P2_P3_lWord_reg[15]/NET0131  , \P2_P3_lWord_reg[1]/NET0131  , \P2_P3_lWord_reg[2]/NET0131  , \P2_P3_lWord_reg[3]/NET0131  , \P2_P3_lWord_reg[4]/NET0131  , \P2_P3_lWord_reg[5]/NET0131  , \P2_P3_lWord_reg[6]/NET0131  , \P2_P3_lWord_reg[7]/NET0131  , \P2_P3_lWord_reg[8]/NET0131  , \P2_P3_lWord_reg[9]/NET0131  , \P2_P3_rEIP_reg[0]/NET0131  , \P2_P3_rEIP_reg[10]/NET0131  , \P2_P3_rEIP_reg[11]/NET0131  , \P2_P3_rEIP_reg[12]/NET0131  , \P2_P3_rEIP_reg[13]/NET0131  , \P2_P3_rEIP_reg[14]/NET0131  , \P2_P3_rEIP_reg[15]/NET0131  , \P2_P3_rEIP_reg[16]/NET0131  , \P2_P3_rEIP_reg[17]/NET0131  , \P2_P3_rEIP_reg[18]/NET0131  , \P2_P3_rEIP_reg[19]/NET0131  , \P2_P3_rEIP_reg[1]/NET0131  , \P2_P3_rEIP_reg[20]/NET0131  , \P2_P3_rEIP_reg[21]/NET0131  , \P2_P3_rEIP_reg[22]/NET0131  , \P2_P3_rEIP_reg[23]/NET0131  , \P2_P3_rEIP_reg[24]/NET0131  , \P2_P3_rEIP_reg[25]/NET0131  , \P2_P3_rEIP_reg[26]/NET0131  , \P2_P3_rEIP_reg[27]/NET0131  , \P2_P3_rEIP_reg[28]/NET0131  , \P2_P3_rEIP_reg[29]/NET0131  , \P2_P3_rEIP_reg[2]/NET0131  , \P2_P3_rEIP_reg[30]/NET0131  , \P2_P3_rEIP_reg[31]/NET0131  , \P2_P3_rEIP_reg[3]/NET0131  , \P2_P3_rEIP_reg[4]/NET0131  , \P2_P3_rEIP_reg[5]/NET0131  , \P2_P3_rEIP_reg[6]/NET0131  , \P2_P3_rEIP_reg[7]/NET0131  , \P2_P3_rEIP_reg[8]/NET0131  , \P2_P3_rEIP_reg[9]/NET0131  , \P2_P3_uWord_reg[0]/NET0131  , \P2_P3_uWord_reg[10]/NET0131  , \P2_P3_uWord_reg[11]/NET0131  , \P2_P3_uWord_reg[12]/NET0131  , \P2_P3_uWord_reg[13]/NET0131  , \P2_P3_uWord_reg[14]/NET0131  , \P2_P3_uWord_reg[1]/NET0131  , \P2_P3_uWord_reg[2]/NET0131  , \P2_P3_uWord_reg[3]/NET0131  , \P2_P3_uWord_reg[4]/NET0131  , \P2_P3_uWord_reg[5]/NET0131  , \P2_P3_uWord_reg[6]/NET0131  , \P2_P3_uWord_reg[7]/NET0131  , \P2_P3_uWord_reg[8]/NET0131  , \P2_P3_uWord_reg[9]/NET0131  , \P2_buf1_reg[0]/NET0131  , \P2_buf1_reg[10]/NET0131  , \P2_buf1_reg[11]/NET0131  , \P2_buf1_reg[12]/NET0131  , \P2_buf1_reg[13]/NET0131  , \P2_buf1_reg[14]/NET0131  , \P2_buf1_reg[15]/NET0131  , \P2_buf1_reg[16]/NET0131  , \P2_buf1_reg[17]/NET0131  , \P2_buf1_reg[18]/NET0131  , \P2_buf1_reg[19]/NET0131  , \P2_buf1_reg[1]/NET0131  , \P2_buf1_reg[20]/NET0131  , \P2_buf1_reg[21]/NET0131  , \P2_buf1_reg[22]/NET0131  , \P2_buf1_reg[23]/NET0131  , \P2_buf1_reg[24]/NET0131  , \P2_buf1_reg[25]/NET0131  , \P2_buf1_reg[26]/NET0131  , \P2_buf1_reg[27]/NET0131  , \P2_buf1_reg[28]/NET0131  , \P2_buf1_reg[29]/NET0131  , \P2_buf1_reg[2]/NET0131  , \P2_buf1_reg[30]/NET0131  , \P2_buf1_reg[3]/NET0131  , \P2_buf1_reg[4]/NET0131  , \P2_buf1_reg[5]/NET0131  , \P2_buf1_reg[6]/NET0131  , \P2_buf1_reg[7]/NET0131  , \P2_buf1_reg[8]/NET0131  , \P2_buf1_reg[9]/NET0131  , \P2_buf2_reg[0]/NET0131  , \P2_buf2_reg[10]/NET0131  , \P2_buf2_reg[11]/NET0131  , \P2_buf2_reg[12]/NET0131  , \P2_buf2_reg[13]/NET0131  , \P2_buf2_reg[14]/NET0131  , \P2_buf2_reg[15]/NET0131  , \P2_buf2_reg[16]/NET0131  , \P2_buf2_reg[17]/NET0131  , \P2_buf2_reg[18]/NET0131  , \P2_buf2_reg[19]/NET0131  , \P2_buf2_reg[1]/NET0131  , \P2_buf2_reg[20]/NET0131  , \P2_buf2_reg[21]/NET0131  , \P2_buf2_reg[22]/NET0131  , \P2_buf2_reg[23]/NET0131  , \P2_buf2_reg[24]/NET0131  , \P2_buf2_reg[25]/NET0131  , \P2_buf2_reg[26]/NET0131  , \P2_buf2_reg[27]/NET0131  , \P2_buf2_reg[28]/NET0131  , \P2_buf2_reg[29]/NET0131  , \P2_buf2_reg[2]/NET0131  , \P2_buf2_reg[30]/NET0131  , \P2_buf2_reg[3]/NET0131  , \P2_buf2_reg[4]/NET0131  , \P2_buf2_reg[5]/NET0131  , \P2_buf2_reg[6]/NET0131  , \P2_buf2_reg[7]/NET0131  , \P2_buf2_reg[8]/NET0131  , \P2_buf2_reg[9]/NET0131  , \P2_ready11_reg/NET0131  , \P2_ready12_reg/NET0131  , \P2_ready21_reg/NET0131  , \P2_ready22_reg/NET0131  , \P3_rd_reg/NET0131  , \P4_B_reg/NET0131  , \P4_IR_reg[0]/NET0131  , \P4_IR_reg[10]/NET0131  , \P4_IR_reg[11]/NET0131  , \P4_IR_reg[12]/NET0131  , \P4_IR_reg[13]/NET0131  , \P4_IR_reg[14]/NET0131  , \P4_IR_reg[15]/NET0131  , \P4_IR_reg[16]/NET0131  , \P4_IR_reg[17]/NET0131  , \P4_IR_reg[18]/NET0131  , \P4_IR_reg[19]/NET0131  , \P4_IR_reg[1]/NET0131  , \P4_IR_reg[20]/NET0131  , \P4_IR_reg[21]/NET0131  , \P4_IR_reg[22]/NET0131  , \P4_IR_reg[23]/NET0131  , \P4_IR_reg[24]/NET0131  , \P4_IR_reg[25]/NET0131  , \P4_IR_reg[26]/NET0131  , \P4_IR_reg[27]/NET0131  , \P4_IR_reg[28]/NET0131  , \P4_IR_reg[29]/NET0131  , \P4_IR_reg[2]/NET0131  , \P4_IR_reg[30]/NET0131  , \P4_IR_reg[3]/NET0131  , \P4_IR_reg[4]/NET0131  , \P4_IR_reg[5]/NET0131  , \P4_IR_reg[6]/NET0131  , \P4_IR_reg[7]/NET0131  , \P4_IR_reg[8]/NET0131  , \P4_IR_reg[9]/NET0131  , \P4_addr_reg[0]/NET0131  , \P4_addr_reg[10]/NET0131  , \P4_addr_reg[11]/NET0131  , \P4_addr_reg[12]/NET0131  , \P4_addr_reg[13]/NET0131  , \P4_addr_reg[14]/NET0131  , \P4_addr_reg[15]/NET0131  , \P4_addr_reg[16]/NET0131  , \P4_addr_reg[17]/NET0131  , \P4_addr_reg[18]/NET0131  , \P4_addr_reg[1]/NET0131  , \P4_addr_reg[2]/NET0131  , \P4_addr_reg[3]/NET0131  , \P4_addr_reg[4]/NET0131  , \P4_addr_reg[5]/NET0131  , \P4_addr_reg[6]/NET0131  , \P4_addr_reg[7]/NET0131  , \P4_addr_reg[8]/NET0131  , \P4_addr_reg[9]/NET0131  , \P4_d_reg[0]/NET0131  , \P4_d_reg[1]/NET0131  , \P4_datao_reg[0]/NET0131  , \P4_datao_reg[10]/NET0131  , \P4_datao_reg[11]/NET0131  , \P4_datao_reg[12]/NET0131  , \P4_datao_reg[13]/NET0131  , \P4_datao_reg[14]/NET0131  , \P4_datao_reg[15]/NET0131  , \P4_datao_reg[16]/NET0131  , \P4_datao_reg[17]/NET0131  , \P4_datao_reg[18]/NET0131  , \P4_datao_reg[19]/NET0131  , \P4_datao_reg[1]/NET0131  , \P4_datao_reg[20]/NET0131  , \P4_datao_reg[21]/NET0131  , \P4_datao_reg[22]/NET0131  , \P4_datao_reg[23]/NET0131  , \P4_datao_reg[24]/NET0131  , \P4_datao_reg[25]/NET0131  , \P4_datao_reg[26]/NET0131  , \P4_datao_reg[27]/NET0131  , \P4_datao_reg[28]/NET0131  , \P4_datao_reg[29]/NET0131  , \P4_datao_reg[2]/NET0131  , \P4_datao_reg[30]/NET0131  , \P4_datao_reg[31]/NET0131  , \P4_datao_reg[3]/NET0131  , \P4_datao_reg[4]/NET0131  , \P4_datao_reg[5]/NET0131  , \P4_datao_reg[6]/NET0131  , \P4_datao_reg[7]/NET0131  , \P4_datao_reg[8]/NET0131  , \P4_datao_reg[9]/NET0131  , \P4_rd_reg/NET0131  , \P4_reg0_reg[0]/NET0131  , \P4_reg0_reg[10]/NET0131  , \P4_reg0_reg[11]/NET0131  , \P4_reg0_reg[12]/NET0131  , \P4_reg0_reg[13]/NET0131  , \P4_reg0_reg[14]/NET0131  , \P4_reg0_reg[15]/NET0131  , \P4_reg0_reg[16]/NET0131  , \P4_reg0_reg[17]/NET0131  , \P4_reg0_reg[18]/NET0131  , \P4_reg0_reg[19]/NET0131  , \P4_reg0_reg[1]/NET0131  , \P4_reg0_reg[20]/NET0131  , \P4_reg0_reg[21]/NET0131  , \P4_reg0_reg[22]/NET0131  , \P4_reg0_reg[23]/NET0131  , \P4_reg0_reg[24]/NET0131  , \P4_reg0_reg[25]/NET0131  , \P4_reg0_reg[26]/NET0131  , \P4_reg0_reg[27]/NET0131  , \P4_reg0_reg[28]/NET0131  , \P4_reg0_reg[29]/NET0131  , \P4_reg0_reg[2]/NET0131  , \P4_reg0_reg[30]/NET0131  , \P4_reg0_reg[31]/NET0131  , \P4_reg0_reg[3]/NET0131  , \P4_reg0_reg[4]/NET0131  , \P4_reg0_reg[5]/NET0131  , \P4_reg0_reg[6]/NET0131  , \P4_reg0_reg[7]/NET0131  , \P4_reg0_reg[8]/NET0131  , \P4_reg0_reg[9]/NET0131  , \P4_reg1_reg[0]/NET0131  , \P4_reg1_reg[10]/NET0131  , \P4_reg1_reg[11]/NET0131  , \P4_reg1_reg[12]/NET0131  , \P4_reg1_reg[13]/NET0131  , \P4_reg1_reg[14]/NET0131  , \P4_reg1_reg[15]/NET0131  , \P4_reg1_reg[16]/NET0131  , \P4_reg1_reg[17]/NET0131  , \P4_reg1_reg[18]/NET0131  , \P4_reg1_reg[19]/NET0131  , \P4_reg1_reg[1]/NET0131  , \P4_reg1_reg[20]/NET0131  , \P4_reg1_reg[21]/NET0131  , \P4_reg1_reg[22]/NET0131  , \P4_reg1_reg[23]/NET0131  , \P4_reg1_reg[24]/NET0131  , \P4_reg1_reg[25]/NET0131  , \P4_reg1_reg[26]/NET0131  , \P4_reg1_reg[27]/NET0131  , \P4_reg1_reg[28]/NET0131  , \P4_reg1_reg[29]/NET0131  , \P4_reg1_reg[2]/NET0131  , \P4_reg1_reg[30]/NET0131  , \P4_reg1_reg[31]/NET0131  , \P4_reg1_reg[3]/NET0131  , \P4_reg1_reg[4]/NET0131  , \P4_reg1_reg[5]/NET0131  , \P4_reg1_reg[6]/NET0131  , \P4_reg1_reg[7]/NET0131  , \P4_reg1_reg[8]/NET0131  , \P4_reg1_reg[9]/NET0131  , \P4_reg2_reg[0]/NET0131  , \P4_reg2_reg[10]/NET0131  , \P4_reg2_reg[11]/NET0131  , \P4_reg2_reg[12]/NET0131  , \P4_reg2_reg[13]/NET0131  , \P4_reg2_reg[14]/NET0131  , \P4_reg2_reg[15]/NET0131  , \P4_reg2_reg[16]/NET0131  , \P4_reg2_reg[17]/NET0131  , \P4_reg2_reg[18]/NET0131  , \P4_reg2_reg[19]/NET0131  , \P4_reg2_reg[1]/NET0131  , \P4_reg2_reg[20]/NET0131  , \P4_reg2_reg[21]/NET0131  , \P4_reg2_reg[22]/NET0131  , \P4_reg2_reg[23]/NET0131  , \P4_reg2_reg[24]/NET0131  , \P4_reg2_reg[25]/NET0131  , \P4_reg2_reg[26]/NET0131  , \P4_reg2_reg[27]/NET0131  , \P4_reg2_reg[28]/NET0131  , \P4_reg2_reg[29]/NET0131  , \P4_reg2_reg[2]/NET0131  , \P4_reg2_reg[30]/NET0131  , \P4_reg2_reg[31]/NET0131  , \P4_reg2_reg[3]/NET0131  , \P4_reg2_reg[4]/NET0131  , \P4_reg2_reg[5]/NET0131  , \P4_reg2_reg[6]/NET0131  , \P4_reg2_reg[7]/NET0131  , \P4_reg2_reg[8]/NET0131  , \P4_reg2_reg[9]/NET0131  , \P4_reg3_reg[0]/NET0131  , \P4_reg3_reg[10]/NET0131  , \P4_reg3_reg[11]/NET0131  , \P4_reg3_reg[12]/NET0131  , \P4_reg3_reg[13]/NET0131  , \P4_reg3_reg[14]/NET0131  , \P4_reg3_reg[15]/NET0131  , \P4_reg3_reg[16]/NET0131  , \P4_reg3_reg[17]/NET0131  , \P4_reg3_reg[18]/NET0131  , \P4_reg3_reg[19]/NET0131  , \P4_reg3_reg[1]/NET0131  , \P4_reg3_reg[20]/NET0131  , \P4_reg3_reg[21]/NET0131  , \P4_reg3_reg[22]/NET0131  , \P4_reg3_reg[23]/NET0131  , \P4_reg3_reg[24]/NET0131  , \P4_reg3_reg[25]/NET0131  , \P4_reg3_reg[26]/NET0131  , \P4_reg3_reg[27]/NET0131  , \P4_reg3_reg[28]/NET0131  , \P4_reg3_reg[2]/NET0131  , \P4_reg3_reg[3]/NET0131  , \P4_reg3_reg[4]/NET0131  , \P4_reg3_reg[5]/NET0131  , \P4_reg3_reg[6]/NET0131  , \P4_reg3_reg[7]/NET0131  , \P4_reg3_reg[8]/NET0131  , \P4_reg3_reg[9]/NET0131  , \P4_wr_reg/NET0131  , bs_pad , \din[0]_pad  , \din[10]_pad  , \din[11]_pad  , \din[12]_pad  , \din[13]_pad  , \din[14]_pad  , \din[15]_pad  , \din[16]_pad  , \din[17]_pad  , \din[18]_pad  , \din[19]_pad  , \din[1]_pad  , \din[20]_pad  , \din[21]_pad  , \din[22]_pad  , \din[23]_pad  , \din[24]_pad  , \din[25]_pad  , \din[26]_pad  , \din[27]_pad  , \din[28]_pad  , \din[29]_pad  , \din[2]_pad  , \din[30]_pad  , \din[31]_pad  , \din[3]_pad  , \din[4]_pad  , \din[5]_pad  , \din[6]_pad  , \din[7]_pad  , \din[8]_pad  , \din[9]_pad  , hold_pad , na_pad , sel_pad , \P3_state_reg[0]/NET0131_syn_2  , \_al_n1  , \aux[0]_pad  , \aux[1]_pad  , \aux[2]_pad  , \dout[0]_pad  , \dout[10]_pad  , \dout[11]_pad  , \dout[12]_pad  , \dout[13]_pad  , \dout[14]_pad  , \dout[15]_pad  , \dout[16]_pad  , \dout[17]_pad  , \dout[18]_pad  , \dout[19]_pad  , \dout[1]_pad  , \dout[2]_pad  , \dout[3]_pad  , \dout[4]_pad  , \dout[5]_pad  , \dout[6]_pad  , \dout[7]_pad  , \dout[8]_pad  , \dout[9]_pad  , \g326201/_0_  , \g326202/_0_  , \g326203/_0_  , \g326204/_0_  , \g326205/_0_  , \g326206/_0_  , \g326207/_0_  , \g326208/_0_  , \g326209/_0_  , \g326210/_0_  , \g326211/_0_  , \g326212/_0_  , \g326213/_0_  , \g326214/_0_  , \g326215/_0_  , \g326216/_0_  , \g326251/_0_  , \g326255/_0_  , \g326256/_0_  , \g326271/_0_  , \g326272/_0_  , \g326273/_0_  , \g326274/_0_  , \g326275/_0_  , \g326276/_0_  , \g326277/_0_  , \g326278/_0_  , \g326279/_0_  , \g326280/_0_  , \g326281/_0_  , \g326282/_0_  , \g326283/_0_  , \g326284/_0_  , \g326285/_0_  , \g326286/_0_  , \g326287/_0_  , \g326288/_0_  , \g326289/_0_  , \g326290/_0_  , \g326291/_0_  , \g326292/_0_  , \g326293/_0_  , \g326294/_0_  , \g326295/_0_  , \g326296/_0_  , \g326297/_0_  , \g326298/_0_  , \g326299/_0_  , \g326300/_0_  , \g326301/_0_  , \g326335/_0_  , \g326369/_0_  , \g326370/_0_  , \g326371/_0_  , \g326372/_0_  , \g326373/_0_  , \g326374/_0_  , \g326375/_0_  , \g326376/_0_  , \g326377/_0_  , \g326378/_0_  , \g326379/_0_  , \g326380/_0_  , \g326381/_0_  , \g326382/_0_  , \g326383/_0_  , \g326384/_0_  , \g326385/_0_  , \g326386/_0_  , \g326387/_0_  , \g326388/_0_  , \g326389/_0_  , \g326390/_0_  , \g326391/_0_  , \g326392/_0_  , \g326393/_0_  , \g326394/_0_  , \g326395/_0_  , \g326396/_0_  , \g326397/_0_  , \g326398/_0_  , \g326399/_0_  , \g326400/_0_  , \g326401/_0_  , \g326423/_0_  , \g326438/_0_  , \g326439/_0_  , \g326440/_0_  , \g326441/_0_  , \g326442/_0_  , \g326443/_0_  , \g326444/_0_  , \g326445/_0_  , \g326446/_0_  , \g326447/_0_  , \g326448/_0_  , \g326449/_0_  , \g326450/_0_  , \g326451/_0_  , \g326452/_0_  , \g326561/_0_  , \g326571/_0_  , \g326572/_0_  , \g326597/_0_  , \g326598/_0_  , \g326599/_0_  , \g326600/_0_  , \g326601/_0_  , \g326602/_0_  , \g326603/_0_  , \g326604/_0_  , \g326605/_0_  , \g326606/_0_  , \g326607/_0_  , \g326608/_0_  , \g326609/_0_  , \g326611/_0_  , \g326612/_0_  , \g326613/_0_  , \g326614/_0_  , \g326615/_0_  , \g326616/_0_  , \g326617/_0_  , \g326618/_0_  , \g326619/_0_  , \g326620/_0_  , \g326621/_0_  , \g326622/_0_  , \g326623/_0_  , \g326624/_0_  , \g326625/_0_  , \g326626/_0_  , \g326627/_0_  , \g326628/_0_  , \g326629/_0_  , \g326630/_0_  , \g326631/_0_  , \g326632/_0_  , \g326633/_0_  , \g326634/_0_  , \g326635/_0_  , \g326636/_0_  , \g326637/_0_  , \g326638/_0_  , \g326639/_0_  , \g326640/_0_  , \g326641/_0_  , \g326798/_0_  , \g326821/_0_  , \g326822/_0_  , \g326823/_0_  , \g326824/_0_  , \g326825/_0_  , \g326826/_0_  , \g326827/_0_  , \g326828/_0_  , \g326829/_0_  , \g326830/_0_  , \g326831/_0_  , \g326832/_0_  , \g326833/_0_  , \g326834/_0_  , \g326835/_0_  , \g326868/_0_  , \g326887/_0_  , \g326926/_0_  , \g326927/_0_  , \g326928/_0_  , \g326929/_0_  , \g326930/_0_  , \g326931/_0_  , \g326932/_0_  , \g326933/_0_  , \g326934/_0_  , \g326935/_0_  , \g326936/_0_  , \g326937/_0_  , \g326938/_0_  , \g326939/_0_  , \g326940/_0_  , \g326941/_0_  , \g326942/_0_  , \g326943/_0_  , \g326944/_0_  , \g326945/_0_  , \g326946/_0_  , \g326947/_0_  , \g326948/_0_  , \g326949/_0_  , \g326950/_0_  , \g326951/_0_  , \g326952/_0_  , \g326953/_0_  , \g326954/_0_  , \g326955/_0_  , \g327192/_0_  , \g327234/_0_  , \g327237/_0_  , \g327241/_0_  , \g327242/_0_  , \g327243/_0_  , \g327247/_0_  , \g327290/_0_  , \g327311/_0_  , \g327369/_0_  , \g327370/_0_  , \g327371/_0_  , \g327373/_0_  , \g327375/_0_  , \g327377/_0_  , \g327379/_0_  , \g327380/_0_  , \g327381/_0_  , \g327382/_0_  , \g327383/_0_  , \g327384/_0_  , \g327385/_0_  , \g327386/_0_  , \g327387/_0_  , \g327388/_0_  , \g327389/_0_  , \g327390/_0_  , \g327391/_0_  , \g327392/_0_  , \g327393/_0_  , \g327394/_0_  , \g327395/_0_  , \g327396/_0_  , \g327397/_0_  , \g327398/_0_  , \g327399/_0_  , \g327400/_0_  , \g327401/_0_  , \g327402/_0_  , \g327601/_0_  , \g327602/_0_  , \g327698/_0_  , \g327781/_0_  , \g327798/_0_  , \g327799/_0_  , \g327800/_0_  , \g327801/_0_  , \g327802/_0_  , \g327803/_0_  , \g327804/_0_  , \g327805/_0_  , \g327806/_0_  , \g327807/_0_  , \g327826/_0_  , \g327828/_0_  , \g327829/_0_  , \g327830/_0_  , \g327831/_0_  , \g327832/_0_  , \g327833/_0_  , \g327834/_0_  , \g327835/_0_  , \g327836/_0_  , \g327970/_0_  , \g328019/_0_  , \g328020/_0_  , \g328021/_0_  , \g328022/_0_  , \g328023/_0_  , \g328024/_0_  , \g328027/_0_  , \g328028/_0_  , \g328029/_0_  , \g328030/_0_  , \g328031/_0_  , \g328032/_0_  , \g328033/_0_  , \g328034/_0_  , \g328035/_0_  , \g328046/_0_  , \g328048/_0_  , \g328049/_0_  , \g328052/_0_  , \g328054/_0_  , \g328056/_0_  , \g328058/_0_  , \g328059/_0_  , \g328060/_0_  , \g328061/_0_  , \g328062/_0_  , \g328063/_0_  , \g328064/_0_  , \g328065/_0_  , \g328066/_0_  , \g328067/_0_  , \g328068/_0_  , \g328069/_0_  , \g328070/_0_  , \g328071/_0_  , \g328120/_0_  , \g328152/_0_  , \g328153/_0_  , \g328154/_0_  , \g328155/_0_  , \g328156/_0_  , \g328157/_0_  , \g328158/_0_  , \g328159/_0_  , \g328160/_0_  , \g328161/_0_  , \g328257/_0_  , \g328280/_0_  , \g328302/_0_  , \g328303/_0_  , \g328332/_0_  , \g328333/_0_  , \g328334/_0_  , \g328335/_0_  , \g328336/_0_  , \g328337/_0_  , \g328338/_0_  , \g328339/_0_  , \g328340/_0_  , \g328341/_0_  , \g328342/_0_  , \g328343/_0_  , \g328344/_0_  , \g328345/_0_  , \g328346/_0_  , \g328347/_0_  , \g328348/_0_  , \g328349/_0_  , \g328350/_0_  , \g328351/_0_  , \g328352/_0_  , \g328353/_0_  , \g328354/_0_  , \g328355/_0_  , \g328356/_0_  , \g328357/_0_  , \g328358/_0_  , \g328359/_0_  , \g328360/_0_  , \g328361/_0_  , \g328372/_0_  , \g328373/_0_  , \g328374/_0_  , \g328375/_0_  , \g328376/_0_  , \g328377/_0_  , \g328378/_0_  , \g328379/_0_  , \g328380/_0_  , \g328381/_0_  , \g328382/_0_  , \g328383/_0_  , \g328384/_0_  , \g328385/_0_  , \g328569/_0_  , \g328587/_0_  , \g328658/_0_  , \g328662/_3_  , \g328664/_3_  , \g328666/_3_  , \g328669/_3_  , \g328670/_0_  , \g328671/_0_  , \g328672/_0_  , \g328674/_0_  , \g328809/_0_  , \g328810/_0_  , \g328811/_0_  , \g328812/_0_  , \g328856/_0_  , \g328887/_0_  , \g328931/_0_  , \g328945/_0_  , \g328960/_0_  , \g328991/_0_  , \g328992/_0_  , \g329022/_3_  , \g329024/_3_  , \g329025/_0_  , \g329026/_0_  , \g329027/_0_  , \g329029/_3_  , \g329030/_0_  , \g329032/_0_  , \g329033/_0_  , \g329034/_0_  , \g329182/_0_  , \g329228/_0_  , \g329281/_0_  , \g329301/_0_  , \g329302/_0_  , \g329322/_2_  , \g329324/_3_  , \g329334/_3_  , \g329336/_3_  , \g329338/_3_  , \g329340/_2_  , \g329342/_3_  , \g329343/_0_  , \g329345/_3_  , \g329347/_3_  , \g329349/_3_  , \g329351/_3_  , \g329353/_3_  , \g329355/_3_  , \g329357/_3_  , \g329359/_3_  , \g329360/_0_  , \g329362/_3_  , \g329364/_3_  , \g329366/_3_  , \g329368/_3_  , \g329370/_3_  , \g329372/_3_  , \g329374/_3_  , \g329376/_3_  , \g329378/_3_  , \g329379/_0_  , \g329380/_0_  , \g329381/_0_  , \g329388/_0_  , \g329516/_0_  , \g329517/_0_  , \g329518/_0_  , \g329587/_0_  , \g329605/_0_  , \g329687/_0_  , \g329703/_0_  , \g329709/_3_  , \g329716/_3_  , \g329718/_3_  , \g329720/_3_  , \g329722/_3_  , \g329724/_3_  , \g329725/_0_  , \g329727/_0_  , \g329805/_0_  , \g329807/_0_  , \g329809/_0_  , \g329810/_0_  , \g329811/_0_  , \g329812/_0_  , \g330065/_3_  , \g330067/_3_  , \g330069/_3_  , \g330071/_3_  , \g330073/_3_  , \g330075/_3_  , \g330077/_3_  , \g330079/_3_  , \g330081/_3_  , \g330083/_3_  , \g330085/_3_  , \g330087/_3_  , \g330089/_3_  , \g330091/_3_  , \g330093/_3_  , \g330095/_3_  , \g330097/_3_  , \g330099/_0_  , \g330188/_0_  , \g330337/_0_  , \g330388/_3_  , \g330418/_3_  , \g330420/_3_  , \g330422/_3_  , \g330424/_3_  , \g330426/_3_  , \g330428/_3_  , \g330429/_0_  , \g330431/_3_  , \g330433/_3_  , \g330435/_3_  , \g330436/_0_  , \g330438/_3_  , \g330440/_3_  , \g330441/_0_  , \g330443/_3_  , \g330444/_0_  , \g330446/_3_  , \g330448/_3_  , \g330450/_3_  , \g330451/_0_  , \g330452/_0_  , \g330453/_0_  , \g330535/_0_  , \g330762/_3_  , \g330764/_3_  , \g330766/_3_  , \g330768/_3_  , \g330770/_3_  , \g330772/_3_  , \g330774/_3_  , \g330776/_3_  , \g331141/_3_  , \g331142/_0_  , \g331144/_3_  , \g331145/_0_  , \g331147/_3_  , \g331484/_0_  , \g331485/_0_  , \g331486/_0_  , \g331497/_0_  , \g331498/_0_  , \g331502/_0_  , \g332061/_0_  , \g332062/_0_  , \g332063/_0_  , \g332064/_0_  , \g332065/_0_  , \g332066/_0_  , \g332070/_0_  , \g332071/_0_  , \g332672/_0_  , \g332673/_0_  , \g332678/_0_  , \g332679/_0_  , \g332680/_0_  , \g332681/_0_  , \g332682/_0_  , \g332700/_0_  , \g333449/_0_  , \g333453/_0_  , \g333454/_0_  , \g333462/_0_  , \g333463/_0_  , \g334369/_0_  , \g334370/_0_  , \g335243/_0_  , \g335244/_0_  , \g335965/_0_  , \g335969/_0_  , \g336538/_0_  , \g336539/_0_  , \g336540/_0_  , \g336546/_0_  , \g336551/_0_  , \g336552/_0_  , \g336557/_0_  , \g336558/_0_  , \g336654/_0_  , \g336655/_0_  , \g336656/_0_  , \g336657/_0_  , \g336660/_0_  , \g336850/_0_  , \g337247/_0_  , \g337248/_0_  , \g337249/_0_  , \g337250/_0_  , \g337251/_0_  , \g337629/_0_  , \g337635/_0_  , \g337637/_0_  , \g337879/_0_  , \g337905/_0_  , \g337906/_0_  , \g337907/_0_  , \g337916/_0_  , \g337917/_0_  , \g337946/_0_  , \g337947/_0_  , \g337948/_0_  , \g337949/_0_  , \g337950/_0_  , \g338030/_0_  , \g338034/_0_  , \g338388/_0_  , \g338442/_0_  , \g338443/_0_  , \g338513/_0_  , \g338514/_0_  , \g338750/_0_  , \g338759/_0_  , \g338800/_0_  , \g338801/_0_  , \g338802/_0_  , \g338803/_0_  , \g338804/_0_  , \g338805/_0_  , \g338806/_0_  , \g338807/_0_  , \g338808/_0_  , \g338809/_0_  , \g338810/_0_  , \g338811/_0_  , \g338812/_0_  , \g338813/_0_  , \g338814/_0_  , \g338815/_0_  , \g338816/_0_  , \g338817/_0_  , \g338818/_0_  , \g338819/_0_  , \g338820/_0_  , \g338821/_0_  , \g338822/_0_  , \g338823/_0_  , \g338824/_0_  , \g338825/_0_  , \g338826/_0_  , \g338827/_0_  , \g338828/_0_  , \g338829/_0_  , \g338869/_0_  , \g338886/_0_  , \g338887/_0_  , \g338888/_0_  , \g339020/_0_  , \g339021/_0_  , \g339022/_0_  , \g339023/_0_  , \g339024/_0_  , \g339045/_0_  , \g339060/_0_  , \g339125/_0_  , \g339142/_0_  , \g339143/_0_  , \g339144/_0_  , \g339145/_0_  , \g339146/_0_  , \g339147/_0_  , \g339148/_0_  , \g339149/_0_  , \g339150/_0_  , \g339151/_0_  , \g339152/_0_  , \g339153/_0_  , \g339154/_0_  , \g339155/_0_  , \g339156/_0_  , \g339157/_0_  , \g339158/_0_  , \g339159/_0_  , \g339160/_0_  , \g339161/_0_  , \g339162/_0_  , \g339163/_0_  , \g339164/_0_  , \g339165/_0_  , \g339166/_0_  , \g339167/_0_  , \g339168/_0_  , \g339169/_0_  , \g339170/_0_  , \g339171/_0_  , \g339254/_0_  , \g339255/_0_  , \g339257/_0_  , \g339458/_0_  , \g339459/_0_  , \g339460/_0_  , \g339461/_0_  , \g339462/_0_  , \g339463/_0_  , \g339464/_0_  , \g339466/_0_  , \g339469/_0_  , \g339470/_0_  , \g339472/_0_  , \g339504/_0_  , \g339505/_0_  , \g339535/_0_  , \g339601/_0_  , \g339614/_0_  , \g339615/_0_  , \g339616/_0_  , \g339617/_0_  , \g339618/_0_  , \g339619/_0_  , \g339620/_0_  , \g339621/_0_  , \g339622/_0_  , \g339623/_0_  , \g339624/_0_  , \g339625/_0_  , \g339626/_0_  , \g339627/_0_  , \g339628/_0_  , \g339629/_0_  , \g339630/_0_  , \g339631/_0_  , \g339632/_0_  , \g339633/_0_  , \g339634/_0_  , \g339635/_0_  , \g339636/_0_  , \g339637/_0_  , \g339638/_0_  , \g339639/_0_  , \g339640/_0_  , \g339641/_0_  , \g339642/_0_  , \g339643/_0_  , \g339644/_0_  , \g339645/_0_  , \g339646/_0_  , \g339647/_0_  , \g339648/_0_  , \g339649/_0_  , \g339650/_0_  , \g339651/_0_  , \g339652/_0_  , \g339653/_0_  , \g339654/_0_  , \g339655/_0_  , \g339656/_0_  , \g339657/_0_  , \g339658/_0_  , \g339718/_0_  , \g339719/_0_  , \g339720/_0_  , \g339721/_0_  , \g339723/_0_  , \g339725/_0_  , \g339727/_0_  , \g340058/_0_  , \g340102/_0_  , \g340103/_0_  , \g340104/_0_  , \g340106/_0_  , \g340109/_0_  , \g340244/_0_  , \g340245/_0_  , \g340246/_0_  , \g340247/_0_  , \g340464/_0_  , \g340505/_0_  , \g340612/_0_  , \g340613/_0_  , \g340614/_0_  , \g340615/_0_  , \g340616/_0_  , \g340617/_0_  , \g340618/_0_  , \g340619/_0_  , \g340620/_0_  , \g340621/_0_  , \g340622/_0_  , \g340623/_0_  , \g340624/_0_  , \g340625/_0_  , \g340626/_0_  , \g340630/_0_  , \g340631/_0_  , \g340632/_0_  , \g340633/_0_  , \g340634/_0_  , \g340635/_0_  , \g340636/_0_  , \g340637/_0_  , \g340638/_0_  , \g340640/_0_  , \g340641/_0_  , \g340642/_0_  , \g340643/_0_  , \g340644/_0_  , \g340645/_0_  , \g340701/_0_  , \g340702/_0_  , \g340703/_0_  , \g340704/_0_  , \g340714/_0_  , \g340716/_0_  , \g340717/_0_  , \g340718/_0_  , \g340728/_0_  , \g340729/_0_  , \g340730/_0_  , \g340731/_0_  , \g340747/_0_  , \g340748/_0_  , \g340749/_0_  , \g340750/_0_  , \g340751/_0_  , \g340752/_0_  , \g340753/_0_  , \g340754/_0_  , \g340792/_0_  , \g340793/_0_  , \g340794/_0_  , \g340795/_0_  , \g340796/_0_  , \g340797/_0_  , \g340988/_0_  , \g341033/_0_  , \g341191/_0_  , \g341192/_0_  , \g341193/_0_  , \g341194/_0_  , \g341195/_0_  , \g341196/_0_  , \g341197/_0_  , \g341198/_0_  , \g341199/_0_  , \g341200/_0_  , \g341201/_0_  , \g341202/_0_  , \g341203/_0_  , \g341205/_0_  , \g341206/_0_  , \g341207/_0_  , \g341208/_0_  , \g341209/_0_  , \g341210/_0_  , \g341211/_0_  , \g341212/_0_  , \g341213/_0_  , \g341214/_0_  , \g341215/_0_  , \g341216/_0_  , \g341217/_0_  , \g341218/_0_  , \g341219/_0_  , \g341220/_0_  , \g341221/_0_  , \g341241/_0_  , \g341242/_0_  , \g341245/_0_  , \g341248/_0_  , \g341250/_0_  , \g341251/_0_  , \g341339/_0_  , \g341347/_0_  , \g341349/_0_  , \g341350/_0_  , \g341352/_0_  , \g341353/_0_  , \g341354/_0_  , \g341365/_0_  , \g341366/_0_  , \g341367/_0_  , \g341368/_0_  , \g341369/_0_  , \g341370/_0_  , \g341373/_0_  , \g341388/_0_  , \g341389/_0_  , \g341390/_0_  , \g341391/_0_  , \g341392/_0_  , \g341393/_0_  , \g341394/_0_  , \g341395/_0_  , \g341396/_0_  , \g341397/_0_  , \g341398/_0_  , \g341400/_0_  , \g341401/_0_  , \g341419/_0_  , \g341435/_0_  , \g341436/_0_  , \g341455/_0_  , \g341456/_0_  , \g341457/_0_  , \g341458/_0_  , \g342136/_0_  , \g342137/_0_  , \g342141/_0_  , \g342145/_0_  , \g342148/_0_  , \g342149/_0_  , \g342308/_0_  , \g342318/_0_  , \g342322/_0_  , \g342323/_0_  , \g342327/_0_  , \g342331/_0_  , \g342333/_0_  , \g342354/_0_  , \g342355/_0_  , \g342356/_0_  , \g342357/_0_  , \g342358/_0_  , \g342359/_0_  , \g342383/_0_  , \g342384/_0_  , \g342385/_0_  , \g342386/_0_  , \g342387/_0_  , \g342388/_0_  , \g342389/_0_  , \g342390/_0_  , \g342391/_0_  , \g342392/_0_  , \g342393/_0_  , \g342394/_0_  , \g342397/_0_  , \g342398/_0_  , \g342399/_0_  , \g342400/_0_  , \g342401/_0_  , \g342454/u3_syn_4  , \g342800/_0_  , \g343406/_0_  , \g343407/_0_  , \g343408/_0_  , \g343409/_0_  , \g343410/_0_  , \g343411/_0_  , \g343412/_0_  , \g343413/_0_  , \g343414/_0_  , \g343415/_0_  , \g343416/_0_  , \g343417/_0_  , \g343418/_0_  , \g343419/_0_  , \g343420/_0_  , \g343431/_0_  , \g343432/_0_  , \g343433/_0_  , \g343434/_0_  , \g343435/_0_  , \g343436/_0_  , \g343437/_0_  , \g343439/_0_  , \g343440/_0_  , \g343441/_0_  , \g343443/_0_  , \g343444/_0_  , \g343445/_0_  , \g343446/_0_  , \g343447/_0_  , \g343452/_0_  , \g343453/_0_  , \g343454/_0_  , \g343455/_0_  , \g343456/_0_  , \g343458/_0_  , \g343459/_0_  , \g343460/_0_  , \g343461/_0_  , \g343462/_0_  , \g343463/_0_  , \g343464/_0_  , \g343465/_0_  , \g343466/_0_  , \g343467/_0_  , \g343512/_0_  , \g343514/_0_  , \g343515/_0_  , \g343517/_0_  , \g343524/_0_  , \g343531/_0_  , \g343533/_0_  , \g343534/_0_  , \g343535/_0_  , \g343536/_0_  , \g343537/_0_  , \g343555/_0_  , \g343556/_0_  , \g343557/_0_  , \g343558/_0_  , \g343559/_0_  , \g343560/_0_  , \g343561/_0_  , \g343563/_0_  , \g343564/_0_  , \g343566/_0_  , \g343567/_0_  , \g343568/_0_  , \g343569/_0_  , \g343570/_0_  , \g343699/_0_  , \g343703/_0_  , \g343944/_0_  , \g343992/_0_  , \g344429/_0_  , \g344430/_0_  , \g344431/_0_  , \g344432/_0_  , \g344433/_0_  , \g344434/_0_  , \g344435/_0_  , \g344437/_0_  , \g344438/_0_  , \g344439/_0_  , \g344440/_0_  , \g344441/_0_  , \g344442/_0_  , \g344443/_0_  , \g344444/_0_  , \g344447/_0_  , \g344448/_0_  , \g344449/_0_  , \g344450/_0_  , \g344451/_0_  , \g344452/_0_  , \g344453/_0_  , \g344454/_0_  , \g344455/_0_  , \g344456/_0_  , \g344457/_0_  , \g344458/_0_  , \g344459/_0_  , \g344460/_0_  , \g344461/_0_  , \g344495/_0_  , \g344496/_0_  , \g344497/_0_  , \g344498/_0_  , \g344499/_0_  , \g344500/_0_  , \g344501/_0_  , \g344502/_0_  , \g344503/_0_  , \g344504/_0_  , \g344505/_0_  , \g344506/_0_  , \g344507/_0_  , \g344508/_0_  , \g344511/_0_  , \g344512/_0_  , \g344513/_0_  , \g344514/_0_  , \g344515/_0_  , \g344516/_0_  , \g344517/_0_  , \g344523/_0_  , \g344524/_0_  , \g344525/_0_  , \g344526/_0_  , \g344527/_0_  , \g344528/_0_  , \g344529/_0_  , \g344536/_0_  , \g344537/_0_  , \g344538/_0_  , \g344539/_0_  , \g344540/_0_  , \g344541/_0_  , \g344542/_0_  , \g344543/_0_  , \g344545/_0_  , \g344546/_0_  , \g344547/_0_  , \g344548/_0_  , \g344549/_0_  , \g344550/_0_  , \g344711/_0_  , \g344712/_0_  , \g344729/_0_  , \g344737/_0_  , \g344738/_0_  , \g344783/_0_  , \g344784/_0_  , \g344786/_0_  , \g344791/_0_  , \g344792/_0_  , \g344816/_0_  , \g344819/_0_  , \g344823/_0_  , \g344825/_0_  , \g345116/_0_  , \g345129/_0_  , \g345149/_0_  , \g345161/_0_  , \g345170/_0_  , \g345237/_0_  , \g345313/_0_  , \g345314/_0_  , \g345316/_0_  , \g345317/_0_  , \g345318/_0_  , \g345319/_0_  , \g345320/_0_  , \g345321/_0_  , \g345322/_0_  , \g345323/_0_  , \g345324/_0_  , \g345325/_0_  , \g345326/_0_  , \g345327/_0_  , \g345328/_0_  , \g345329/_0_  , \g345333/_0_  , \g345334/_0_  , \g345335/_0_  , \g345336/_0_  , \g345337/_0_  , \g345338/_0_  , \g345339/_0_  , \g345340/_0_  , \g345349/_0_  , \g345350/_0_  , \g345351/_0_  , \g345352/_0_  , \g345353/_0_  , \g345354/_0_  , \g345355/_0_  , \g345356/_0_  , \g345365/_0_  , \g345366/_0_  , \g345367/_0_  , \g345368/_0_  , \g345369/_0_  , \g345370/_0_  , \g345371/_0_  , \g345373/_0_  , \g345374/_0_  , \g345377/_0_  , \g345378/_0_  , \g345379/_0_  , \g345380/_0_  , \g345381/_0_  , \g345382/_0_  , \g345383/_0_  , \g345488/_0_  , \g345491/_0_  , \g345524/_0_  , \g345525/_0_  , \g345545/_0_  , \g345546/_0_  , \g345574/_0_  , \g345575/_0_  , \g345638/_0_  , \g345639/_0_  , \g345690/_0_  , \g345691/_0_  , \g345692/_0_  , \g345694/_0_  , \g345695/_0_  , \g345698/_0_  , \g345699/_0_  , \g345701/_0_  , \g345703/_0_  , \g346299/_0_  , \g346326/_0_  , \g346364/_0_  , \g346707/_0_  , \g346711/_0_  , \g346721/_0_  , \g346726/_0_  , \g346729/_0_  , \g346730/_0_  , \g346731/_0_  , \g346733/_0_  , \g346735/_0_  , \g346738/_0_  , \g346740/_0_  , \g346741/_0_  , \g346746/_0_  , \g346748/_0_  , \g346750/_0_  , \g346751/_0_  , \g346758/_0_  , \g346759/_0_  , \g346761/_0_  , \g346762/_0_  , \g346763/_0_  , \g346765/_0_  , \g346766/_0_  , \g346965/_0_  , \g346971/_0_  , \g346981/_0_  , \g346986/_0_  , \g346988/_0_  , \g346989/_0_  , \g346994/_0_  , \g346998/_0_  , \g347015/_0_  , \g347016/_0_  , \g347017/_0_  , \g347018/_0_  , \g347019/_0_  , \g347020/_0_  , \g347043/_0_  , \g347050/_0_  , \g347051/_0_  , \g347052/_0_  , \g347053/_0_  , \g347054/_0_  , \g347055/_0_  , \g347056/_0_  , \g347057/_0_  , \g347058/_0_  , \g347059/_0_  , \g347061/_0_  , \g347062/_0_  , \g347063/_0_  , \g347064/_0_  , \g347065/_0_  , \g347066/_0_  , \g347067/_0_  , \g347068/_0_  , \g347069/_0_  , \g347070/_0_  , \g347071/_0_  , \g347083/_0_  , \g347085/_0_  , \g347087/_0_  , \g347089/_0_  , \g347090/_0_  , \g347091/_0_  , \g347092/_0_  , \g347093/_0_  , \g347096/_0_  , \g347097/_0_  , \g347098/_0_  , \g347099/_0_  , \g347100/_0_  , \g347101/_0_  , \g347102/_0_  , \g347104/_0_  , \g347106/_0_  , \g347108/_0_  , \g347318/_0_  , \g347400/_0_  , \g347449/_0_  , \g347477/_0_  , \g347488/_0_  , \g347531/_0_  , \g347537/_0_  , \g347544/_0_  , \g347546/_0_  , \g347553/_0_  , \g347560/_0_  , \g347569/_0_  , \g347575/_0_  , \g347581/_1_  , \g347587/_0_  , \g347592/_0_  , \g347597/_0_  , \g347603/_0_  , \g347610/_0_  , \g347611/_0_  , \g347616/_0_  , \g347624/_0_  , \g347628/_1_  , \g347632/_0_  , \g347641/_0_  , \g347645/_0_  , \g347653/_0_  , \g347661/_0_  , \g347671/_0_  , \g347678/_0_  , \g347881/_0_  , \g347883/_0_  , \g347885/_0_  , \g347886/_0_  , \g347888/_0_  , \g347889/_0_  , \g347890/_0_  , \g347891/_0_  , \g347892/_0_  , \g347893/_0_  , \g347895/_0_  , \g347896/_0_  , \g347897/_0_  , \g347898/_0_  , \g347899/_0_  , \g347902/_0_  , \g347903/_0_  , \g347904/_0_  , \g347906/_0_  , \g347907/_0_  , \g347908/_0_  , \g347909/_0_  , \g347910/_0_  , \g347911/_0_  , \g347912/_0_  , \g347913/_0_  , \g347914/_0_  , \g347915/_0_  , \g347916/_0_  , \g347917/_0_  , \g347974/_0_  , \g347977/_0_  , \g347983/_0_  , \g347999/_0_  , \g348012/_0_  , \g348015/_0_  , \g348288/_0_  , \g348291/_0_  , \g348292/_0_  , \g348293/_0_  , \g348294/_0_  , \g348295/_0_  , \g348296/_0_  , \g348300/_0_  , \g348301/_0_  , \g348302/_0_  , \g348303/_0_  , \g348304/_0_  , \g348307/_0_  , \g348308/_0_  , \g349018/_0_  , \g349020/_0_  , \g349021/_0_  , \g349025/_0_  , \g349026/_0_  , \g349027/_0_  , \g349035/_0_  , \g349036/_0_  , \g349037/_0_  , \g349049/_0_  , \g349050/_0_  , \g349051/_0_  , \g349070/_0_  , \g349071/_0_  , \g349072/_0_  , \g349076/_0_  , \g349077/_0_  , \g349078/_0_  , \g349326/_0_  , \g349333/_0_  , \g349334/_0_  , \g349335/_0_  , \g349343/_0_  , \g349345/_0_  , \g349349/_0_  , \g349350/_0_  , \g349355/_0_  , \g349357/_0_  , \g349358/_0_  , \g349873/_0_  , \g350037/_0_  , \g350042/_0_  , \g350050/_0_  , \g350051/_0_  , \g350089/_0_  , \g350090/_0_  , \g350093/_0_  , \g350094/_0_  , \g350096/_0_  , \g350097/_0_  , \g350165/_0_  , \g350166/_0_  , \g350168/_0_  , \g350170/_0_  , \g350171/_0_  , \g350172/_0_  , \g350173/_0_  , \g350174/_0_  , \g350175/_0_  , \g350176/_0_  , \g350177/_0_  , \g350178/_0_  , \g350179/_0_  , \g350180/_0_  , \g350181/_0_  , \g350183/_0_  , \g350184/_0_  , \g350185/_0_  , \g350186/_0_  , \g350187/_0_  , \g350188/_0_  , \g350189/_0_  , \g350190/_0_  , \g350191/_0_  , \g350192/_0_  , \g350193/_0_  , \g350194/_0_  , \g350195/_0_  , \g350196/_0_  , \g350197/_0_  , \g350198/_0_  , \g350199/_0_  , \g350200/_0_  , \g350201/_0_  , \g350202/_0_  , \g350203/_0_  , \g350204/_0_  , \g350205/_0_  , \g350654/_0_  , \g350655/_0_  , \g350656/_0_  , \g350658/_0_  , \g350660/_0_  , \g350661/_0_  , \g350662/_0_  , \g350663/_0_  , \g350664/_0_  , \g350665/_0_  , \g350666/_0_  , \g350667/_0_  , \g350668/_0_  , \g350669/_0_  , \g350670/_0_  , \g350671/_0_  , \g350672/_0_  , \g350673/_0_  , \g350674/_0_  , \g350675/_0_  , \g350676/_0_  , \g350677/_0_  , \g350678/_0_  , \g350679/_0_  , \g350680/_0_  , \g350681/_0_  , \g350682/_0_  , \g350683/_0_  , \g350684/_0_  , \g350685/_0_  , \g350686/_0_  , \g350687/_0_  , \g350723/_0_  , \g350724/_0_  , \g350725/_0_  , \g350726/_0_  , \g350727/_0_  , \g350728/_0_  , \g350729/_0_  , \g350730/_0_  , \g350731/_0_  , \g350814/_0_  , \g350815/_0_  , \g350816/_0_  , \g350817/_0_  , \g350818/_0_  , \g350819/_0_  , \g350820/_0_  , \g350821/_0_  , \g350822/_0_  , \g350823/_0_  , \g350824/_0_  , \g350825/_0_  , \g350826/_0_  , \g350827/_0_  , \g350828/_0_  , \g350829/_0_  , \g350830/_0_  , \g350831/_0_  , \g350832/_0_  , \g350833/_0_  , \g350834/_0_  , \g350835/_0_  , \g350836/_0_  , \g350839/_0_  , \g350840/_0_  , \g350842/_0_  , \g350843/_0_  , \g350844/_0_  , \g350845/_0_  , \g350846/_0_  , \g350847/_0_  , \g350848/_0_  , \g350849/_0_  , \g350850/_0_  , \g350852/_0_  , \g350853/_0_  , \g350854/_0_  , \g350856/_0_  , \g350857/_0_  , \g350858/_0_  , \g350859/_0_  , \g350860/_0_  , \g350861/_0_  , \g350862/_0_  , \g350863/_0_  , \g350866/_0_  , \g350867/_0_  , \g350868/_0_  , \g350869/_0_  , \g350870/_0_  , \g350871/_0_  , \g350872/_0_  , \g350873/_0_  , \g350874/_0_  , \g350952/_0_  , \g350959/_0_  , \g350961/_0_  , \g350964/_0_  , \g350974/_0_  , \g350977/_0_  , \g351003/_0_  , \g351005/_0_  , \g351037/_0_  , \g351045/_0_  , \g351048/_0_  , \g351129/_0_  , \g351147/_0_  , \g351169/_0_  , \g351171/_0_  , \g351175/_0_  , \g351195/_0_  , \g351196/_0_  , \g351197/_0_  , \g351198/_0_  , \g351201/_0_  , \g351202/_0_  , \g351203/_0_  , \g351204/_0_  , \g351205/_0_  , \g351206/_0_  , \g351207/_0_  , \g351208/_0_  , \g351209/_0_  , \g351210/_0_  , \g351211/_0_  , \g351214/_0_  , \g351215/_0_  , \g351216/_0_  , \g351217/_0_  , \g351218/_0_  , \g351219/_0_  , \g351220/_0_  , \g351221/_0_  , \g351222/_0_  , \g351223/_0_  , \g351224/_0_  , \g351225/_0_  , \g351226/_0_  , \g351227/_0_  , \g351228/_0_  , \g351229/_0_  , \g351230/_0_  , \g351231/_0_  , \g351671/_0_  , \g351699/_0_  , \g351703/_0_  , \g351704/_0_  , \g351709/_0_  , \g351711/_0_  , \g351712/_0_  , \g351715/_0_  , \g351716/_0_  , \g351717/_0_  , \g351721/_0_  , \g351722/_0_  , \g351723/_0_  , \g351724/_0_  , \g351725/_0_  , \g351726/_0_  , \g351727/_0_  , \g351728/_0_  , \g351739/_0_  , \g351741/_0_  , \g351742/_0_  , \g351750/_0_  , \g351752/_0_  , \g351753/_0_  , \g351756/_0_  , \g351757/_0_  , \g351759/_0_  , \g351760/_0_  , \g351761/_0_  , \g351766/_0_  , \g351767/_0_  , \g351768/_0_  , \g351771/_0_  , \g351772/_0_  , \g351773/_0_  , \g351775/_0_  , \g351776/_0_  , \g351779/_0_  , \g351780/_0_  , \g351782/_0_  , \g351785/_0_  , \g351786/_0_  , \g351788/_0_  , \g351789/_0_  , \g351790/_0_  , \g351791/_0_  , \g351792/_0_  , \g351793/_0_  , \g351794/_0_  , \g351795/_0_  , \g351796/_0_  , \g351797/_0_  , \g351798/_0_  , \g351799/_0_  , \g351800/_0_  , \g351801/_0_  , \g351802/_0_  , \g351803/_0_  , \g351804/_0_  , \g351805/_0_  , \g351806/_0_  , \g351807/_0_  , \g351808/_0_  , \g351809/_0_  , \g351810/_0_  , \g351811/_0_  , \g351812/_0_  , \g351814/_0_  , \g351817/_0_  , \g351818/_0_  , \g351819/_0_  , \g351821/_0_  , \g351822/_0_  , \g351823/_0_  , \g351841/_0_  , \g351842/_0_  , \g351843/_0_  , \g351844/_0_  , \g351845/_0_  , \g351846/_0_  , \g351847/_0_  , \g351848/_0_  , \g351849/_0_  , \g351850/_0_  , \g351851/_0_  , \g351852/_0_  , \g351853/_0_  , \g351854/_0_  , \g351855/_0_  , \g351856/_0_  , \g351857/_0_  , \g351858/_0_  , \g351859/_0_  , \g351860/_0_  , \g351861/_0_  , \g351862/_0_  , \g351863/_0_  , \g351864/_0_  , \g351865/_0_  , \g351866/_0_  , \g351867/_0_  , \g351868/_0_  , \g351869/_0_  , \g351870/_0_  , \g351871/_0_  , \g351872/_0_  , \g351873/_0_  , \g351874/_0_  , \g351875/_0_  , \g351876/_0_  , \g351877/_0_  , \g351878/_0_  , \g351879/_0_  , \g351880/_0_  , \g351881/_0_  , \g351882/_0_  , \g351883/_0_  , \g351884/_0_  , \g351885/_0_  , \g351889/_0_  , \g351920/_0_  , \g351921/_0_  , \g351922/_0_  , \g351923/_0_  , \g351924/_0_  , \g351925/_0_  , \g351926/_0_  , \g351927/_0_  , \g351928/_0_  , \g351929/_0_  , \g351930/_0_  , \g351954/_0_  , \g351955/_0_  , \g351956/_0_  , \g351957/_0_  , \g352167/_0_  , \g352178/_0_  , \g352211/_0_  , \g352215/_0_  , \g352219/_0_  , \g352237/_0_  , \g352238/_0_  , \g352239/_0_  , \g352240/_0_  , \g352241/_0_  , \g352242/_0_  , \g352243/_0_  , \g352244/_0_  , \g352245/_0_  , \g352246/_0_  , \g352247/_0_  , \g352248/_0_  , \g352249/_0_  , \g352250/_0_  , \g352251/_0_  , \g352252/_0_  , \g352253/_0_  , \g352254/_0_  , \g352255/_0_  , \g352256/_0_  , \g352257/_0_  , \g352258/_0_  , \g352259/_0_  , \g352260/_0_  , \g352261/_0_  , \g352262/_0_  , \g352263/_0_  , \g352264/_0_  , \g352265/_0_  , \g352266/_0_  , \g352267/_0_  , \g352268/_0_  , \g352269/_0_  , \g352271/_0_  , \g352272/_0_  , \g352273/_0_  , \g352274/_0_  , \g352275/_0_  , \g352276/_0_  , \g352277/_0_  , \g352278/_0_  , \g352279/_0_  , \g352280/_0_  , \g352281/_0_  , \g352282/_0_  , \g352283/_0_  , \g352284/_0_  , \g352285/_0_  , \g352286/_0_  , \g352287/_0_  , \g352288/_0_  , \g352289/_0_  , \g352290/_0_  , \g352291/_0_  , \g352292/_0_  , \g352293/_0_  , \g352294/_0_  , \g352295/_0_  , \g352296/_0_  , \g352297/_0_  , \g352298/_0_  , \g352299/_0_  , \g352300/_0_  , \g352301/_0_  , \g352302/_0_  , \g352303/_0_  , \g352304/_0_  , \g352305/_0_  , \g352306/_0_  , \g352307/_0_  , \g352308/_0_  , \g352309/_0_  , \g352310/_0_  , \g352311/_0_  , \g352312/_0_  , \g352313/_0_  , \g352314/_0_  , \g352315/_0_  , \g352525/_0_  , \g352527/_0_  , \g352529/_0_  , \g352547/_0_  , \g352553/_0_  , \g352554/_0_  , \g352556/_0_  , \g352558/_0_  , \g352559/_0_  , \g352560/_0_  , \g352561/_0_  , \g352563/_0_  , \g352564/_0_  , \g352565/_0_  , \g352567/_0_  , \g352568/_0_  , \g352569/_0_  , \g352570/_0_  , \g352572/_0_  , \g352574/_0_  , \g352575/_0_  , \g352577/_0_  , \g352579/_0_  , \g352581/_0_  , \g352583/_0_  , \g352584/_0_  , \g352585/_0_  , \g352586/_0_  , \g352587/_0_  , \g352588/_0_  , \g352589/_0_  , \g352590/_0_  , \g352591/_0_  , \g352592/_0_  , \g352593/_0_  , \g352594/_0_  , \g352595/_0_  , \g352596/_0_  , \g352597/_0_  , \g352598/_0_  , \g352599/_0_  , \g352600/_0_  , \g352601/_0_  , \g352602/_0_  , \g352603/_0_  , \g352605/_0_  , \g352606/_0_  , \g352607/_0_  , \g352608/_0_  , \g352609/_0_  , \g352610/_0_  , \g352611/_0_  , \g352612/_0_  , \g352613/_0_  , \g352614/_0_  , \g352615/_0_  , \g352616/_0_  , \g352617/_0_  , \g352618/_0_  , \g352619/_0_  , \g352620/_0_  , \g352621/_0_  , \g352622/_0_  , \g352623/_0_  , \g352624/_0_  , \g352625/_0_  , \g352626/_0_  , \g352627/_0_  , \g352628/_0_  , \g352629/_0_  , \g352662/_0_  , \g352663/_0_  , \g352666/_0_  , \g352667/_0_  , \g352668/_0_  , \g352676/_0_  , \g352677/_0_  , \g352678/_0_  , \g352683/_0_  , \g352684/_0_  , \g352685/_0_  , \g353014/_0_  , \g353016/_0_  , \g353035/_0_  , \g353036/_0_  , \g353065/_0_  , \g353067/_0_  , \g353071/_0_  , \g353073/_0_  , \g353085/_0_  , \g353087/_0_  , \g353116/_0_  , \g353119/_0_  , \g353120/_0_  , \g353121/_0_  , \g353122/_0_  , \g353123/_0_  , \g353124/_0_  , \g353125/_0_  , \g353126/_0_  , \g353127/_0_  , \g353128/_0_  , \g353130/_0_  , \g353131/_0_  , \g353132/_0_  , \g353133/_0_  , \g353134/_0_  , \g353135/_0_  , \g353136/_0_  , \g353137/_0_  , \g353138/_0_  , \g353142/_0_  , \g353148/_0_  , \g353149/_0_  , \g353150/_0_  , \g353151/_0_  , \g353152/_0_  , \g353153/_0_  , \g353154/_0_  , \g353155/_0_  , \g353157/_0_  , \g353158/_0_  , \g353159/_0_  , \g353160/_0_  , \g353161/_0_  , \g353162/_0_  , \g353163/_0_  , \g353164/_0_  , \g353165/_0_  , \g353166/_0_  , \g353167/_0_  , \g353168/_0_  , \g353169/_0_  , \g353170/_0_  , \g353171/_0_  , \g353172/_0_  , \g353173/_0_  , \g353174/_0_  , \g353175/_0_  , \g353176/_0_  , \g353177/_0_  , \g353178/_0_  , \g353179/_0_  , \g353180/_0_  , \g353181/_0_  , \g353184/_0_  , \g353185/_0_  , \g353186/_0_  , \g353187/_0_  , \g353188/_0_  , \g353189/_0_  , \g353190/_0_  , \g353191/_0_  , \g353192/_0_  , \g353193/_0_  , \g353194/_0_  , \g353195/_0_  , \g353196/_0_  , \g353197/_0_  , \g353198/_0_  , \g353199/_0_  , \g353200/_0_  , \g353201/_0_  , \g353202/_0_  , \g353203/_0_  , \g353204/_0_  , \g353205/_0_  , \g353206/_0_  , \g353207/_0_  , \g353208/_0_  , \g353209/_0_  , \g353210/_0_  , \g353211/_0_  , \g353212/_0_  , \g353213/_0_  , \g353214/_0_  , \g353215/_0_  , \g353216/_0_  , \g353217/_0_  , \g353218/_0_  , \g353219/_0_  , \g353220/_0_  , \g353221/_0_  , \g353222/_0_  , \g353223/_0_  , \g353224/_0_  , \g353225/_0_  , \g353226/_0_  , \g353227/_0_  , \g353228/_0_  , \g353229/_0_  , \g353230/_0_  , \g353231/_0_  , \g353232/_0_  , \g353233/_0_  , \g353234/_0_  , \g353235/_0_  , \g353236/_0_  , \g353237/_0_  , \g353238/_0_  , \g353239/_0_  , \g353240/_0_  , \g353241/_0_  , \g353242/_0_  , \g353243/_0_  , \g353244/_0_  , \g353245/_0_  , \g353246/_0_  , \g353247/_0_  , \g353248/_0_  , \g353249/_0_  , \g353250/_0_  , \g353251/_0_  , \g353252/_0_  , \g353253/_0_  , \g353254/_0_  , \g353255/_0_  , \g353256/_0_  , \g353257/_0_  , \g353258/_0_  , \g353259/_0_  , \g353260/_0_  , \g353261/_0_  , \g353262/_0_  , \g353263/_0_  , \g353264/_0_  , \g353265/_0_  , \g353266/_0_  , \g353267/_0_  , \g353268/_0_  , \g353269/_0_  , \g353270/_0_  , \g353271/_0_  , \g353272/_0_  , \g353273/_0_  , \g353274/_0_  , \g353275/_0_  , \g353276/_0_  , \g353277/_0_  , \g353278/_0_  , \g353279/_0_  , \g353280/_0_  , \g353281/_0_  , \g354206/_0_  , \g354214/_0_  , \g354216/_0_  , \g354217/_0_  , \g354222/_0_  , \g354278/_0_  , \g354282/_0_  , \g354284/_0_  , \g354289/_0_  , \g354301/_0_  , \g354330/_0_  , \g354331/_0_  , \g354332/_0_  , \g354333/_0_  , \g354335/_0_  , \g354336/_0_  , \g354337/_0_  , \g354338/_0_  , \g354339/_0_  , \g354340/_0_  , \g354341/_0_  , \g354342/_0_  , \g354343/_0_  , \g354344/_0_  , \g354345/_0_  , \g354346/_0_  , \g354358/_0_  , \g354364/_0_  , \g354442/_0_  , \g354444/_0_  , \g354445/_0_  , \g354447/_0_  , \g354448/_0_  , \g354449/_0_  , \g354450/_0_  , \g354451/_0_  , \g354452/_0_  , \g354455/_0_  , \g354456/_0_  , \g354464/_0_  , \g354465/_0_  , \g354466/_0_  , \g354468/_0_  , \g354469/_0_  , \g354470/_0_  , \g354471/_0_  , \g354472/_0_  , \g354473/_0_  , \g354474/_0_  , \g354477/_0_  , \g354478/_0_  , \g354479/_0_  , \g354480/_0_  , \g354482/_0_  , \g354483/_0_  , \g354484/_0_  , \g354485/_0_  , \g354486/_0_  , \g354487/_0_  , \g354488/_0_  , \g354490/_0_  , \g354491/_0_  , \g354492/_0_  , \g354493/_0_  , \g354494/_0_  , \g354495/_0_  , \g354504/_0_  , \g354505/_0_  , \g354506/_0_  , \g354508/_0_  , \g354509/_0_  , \g354510/_0_  , \g354511/_0_  , \g354512/_0_  , \g354513/_0_  , \g354522/_0_  , \g354524/_0_  , \g354525/_0_  , \g354526/_0_  , \g354527/_0_  , \g354920/_1_  , \g355460/_0_  , \g355461/_0_  , \g355463/_0_  , \g355464/_0_  , \g355466/_0_  , \g355467/_0_  , \g355470/_0_  , \g355471/_0_  , \g355475/_0_  , \g355476/_0_  , \g355477/_0_  , \g355479/_0_  , \g355480/_0_  , \g355481/_0_  , \g355482/_0_  , \g355483/_0_  , \g355508/_0_  , \g355509/_0_  , \g355510/_0_  , \g355511/_0_  , \g355512/_0_  , \g355513/_0_  , \g355514/_0_  , \g355515/_0_  , \g355520/_0_  , \g355521/_0_  , \g355523/_0_  , \g355525/_0_  , \g355527/_0_  , \g355530/_0_  , \g355532/_0_  , \g355534/_0_  , \g355564/_0_  , \g355565/_0_  , \g355566/_0_  , \g355567/_0_  , \g355568/_0_  , \g355569/_0_  , \g355570/_0_  , \g355571/_0_  , \g355980/_0_  , \g356052/_0_  , \g356106/_0_  , \g356111/_0_  , \g356114/_0_  , \g356117/_0_  , \g356122/_0_  , \g356126/_0_  , \g356129/_0_  , \g356133/_0_  , \g356142/_0_  , \g356148/_0_  , \g356151/_0_  , \g356155/_0_  , \g356160/_0_  , \g356162/_0_  , \g356165/_0_  , \g356167/_0_  , \g356170/_0_  , \g356174/_0_  , \g356176/_0_  , \g356179/_0_  , \g356183/_0_  , \g356185/_0_  , \g356189/_0_  , \g356193/_0_  , \g356196/_0_  , \g356199/_0_  , \g356202/_0_  , \g356205/_0_  , \g356207/_0_  , \g356210/_0_  , \g356213/_0_  , \g356215/_0_  , \g357046/_0_  , \g357047/_0_  , \g357048/_0_  , \g357051/_0_  , \g357052/_0_  , \g357053/_0_  , \g357054/_0_  , \g357055/_0_  , \g357056/_0_  , \g357057/_0_  , \g357058/_0_  , \g357059/_0_  , \g357060/_0_  , \g357061/_0_  , \g357062/_0_  , \g357063/_0_  , \g357064/_0_  , \g357065/_0_  , \g357066/_0_  , \g357067/_0_  , \g357068/_0_  , \g357069/_0_  , \g357070/_0_  , \g357071/_0_  , \g357072/_0_  , \g357073/_0_  , \g357074/_0_  , \g357099/_0_  , \g357100/_0_  , \g357101/_0_  , \g357102/_0_  , \g357103/_0_  , \g357104/_0_  , \g357105/_0_  , \g357106/_0_  , \g357107/_0_  , \g357108/_0_  , \g357109/_0_  , \g357110/_0_  , \g357111/_0_  , \g357112/_0_  , \g357113/_0_  , \g357114/_0_  , \g357116/_0_  , \g357119/_0_  , \g357121/_0_  , \g357122/_0_  , \g357123/_0_  , \g357124/_0_  , \g357125/_0_  , \g357126/_0_  , \g357128/_0_  , \g357129/_0_  , \g357130/_0_  , \g357131/_0_  , \g357132/_0_  , \g357133/_0_  , \g357134/_0_  , \g357135/_0_  , \g357142/_0_  , \g357144/_0_  , \g357145/_0_  , \g357146/_0_  , \g357147/_0_  , \g357148/_0_  , \g357149/_0_  , \g357150/_0_  , \g357151/_0_  , \g357152/_0_  , \g357153/_0_  , \g357154/_0_  , \g357155/_0_  , \g357156/_0_  , \g357157/_0_  , \g357158/_0_  , \g357160/_0_  , \g357161/_0_  , \g357163/_0_  , \g357164/_0_  , \g357165/_0_  , \g357288/_0_  , \g357289/_0_  , \g357413/_0_  , \g357414/_0_  , \g357464/_0_  , \g357510/_0_  , \g357733/_0_  , \g357769/_0_  , \g357781/_0_  , \g357828/_0_  , \g358792/_0_  , \g358802/_0_  , \g359042/_0_  , \g359043/_0_  , \g359045/_0_  , \g359048/_0_  , \g359051/_0_  , \g359053/_0_  , \g359057/_0_  , \g359060/_0_  , \g359064/_0_  , \g359070/_0_  , \g359074/_0_  , \g359077/_0_  , \g359080/_0_  , \g359086/_0_  , \g359087/_0_  , \g359088/_0_  , \g359090/_0_  , \g359092/_0_  , \g359094/_0_  , \g359096/_0_  , \g359097/_0_  , \g359099/_0_  , \g359101/_0_  , \g359102/_0_  , \g359104/_0_  , \g359106/_0_  , \g359107/_0_  , \g359108/_0_  , \g359110/_0_  , \g359111/_0_  , \g359112/_0_  , \g359113/_0_  , \g359116/_0_  , \g359118/_0_  , \g359572/_0_  , \g359573/_0_  , \g359577/_0_  , \g359585/_0_  , \g359887/_0_  , \g359888/_0_  , \g360077/_0_  , \g360083/_0_  , \g360113/_0_  , \g360124/_0_  , \g360302/_0_  , \g360303/_0_  , \g360304/_0_  , \g360305/_0_  , \g360320/_0_  , \g360325/_0_  , \g360361/_0_  , \g360371/_0_  , \g360440/_0_  , \g360441/_0_  , \g360443/_0_  , \g360445/_0_  , \g360446/_0_  , \g360448/_0_  , \g360450/_0_  , \g360453/_0_  , \g360462/_0_  , \g360469/_0_  , \g360476/_0_  , \g360478/_0_  , \g360480/_0_  , \g360485/_0_  , \g360487/_0_  , \g360489/_0_  , \g360491/_0_  , \g360492/_0_  , \g360494/_0_  , \g360497/_0_  , \g360498/_0_  , \g360504/_0_  , \g360506/_0_  , \g360514/_0_  , \g360516/_0_  , \g360518/_0_  , \g360522/_0_  , \g360524/_0_  , \g360527/_0_  , \g360528/_0_  , \g360530/_0_  , \g360533/_0_  , \g360535/_0_  , \g360538/_0_  , \g360539/_0_  , \g360542/_0_  , \g360546/_0_  , \g360593/_0_  , \g361116/_0_  , \g361128/_0_  , \g361132/_0_  , \g361137/_0_  , \g361616/_0_  , \g361624/_0_  , \g361626/_0_  , \g361627/_0_  , \g361630/_0_  , \g361631/_0_  , \g362129/_0_  , \g362558/_0_  , \g362560/_0_  , \g362564/_0_  , \g362567/_0_  , \g362575/_0_  , \g362586/_0_  , \g362598/_0_  , \g362608/_0_  , \g362627/_0_  , \g362638/_0_  , \g362648/_0_  , \g362650/_0_  , \g362653/_0_  , \g362663/_0_  , \g362664/_0_  , \g362667/_0_  , \g362671/_0_  , \g362673/_0_  , \g362676/_0_  , \g362679/_0_  , \g362686/_0_  , \g362688/_0_  , \g362693/_0_  , \g362697/_0_  , \g362703/_0_  , \g363274/_0_  , \g363290/_0_  , \g363294/_0_  , \g363303/_0_  , \g363608/_0_  , \g363609/_0_  , \g363615/_0_  , \g363616/_0_  , \g363617/_0_  , \g363627/_0_  , \g363818/_3_  , \g365385/_0_  , \g365388/_0_  , \g365391/_0_  , \g365393/_0_  , \g365394/_0_  , \g365398/_0_  , \g365474/_0_  , \g365477/_0_  , \g366167/_0_  , \g366168/_0_  , \g366169/_0_  , \g366170/_0_  , \g366171/_0_  , \g366172/_0_  , \g366173/_0_  , \g366174/_0_  , \g366523/_3_  , \g369170/_0_  , \g369171/_0_  , \g369173/_0_  , \g369177/_0_  , \g369289/_0_  , \g369290/_0_  , \g369291/_0_  , \g369292/_0_  , \g369293/_0_  , \g369294/_0_  , \g369453/_3_  , \g371379/_0_  , \g371381/_0_  , \g371384/_0_  , \g371386/_0_  , \g371387/_0_  , \g371391/_0_  , \g372221/_0_  , \g372222/_0_  , \g372232/_0_  , \g372246/_0_  , \g372249/_0_  , \g372250/_0_  , \g372251/_0_  , \g372252/_0_  , \g372253/_0_  , \g372254/_0_  , \g372454/_3_  , \g372455/_3_  , \g372456/_3_  , \g372457/_3_  , \g372458/_3_  , \g372459/_3_  , \g372460/_3_  , \g372461/_3_  , \g372462/_3_  , \g372463/_3_  , \g372464/_3_  , \g372465/_3_  , \g372466/_3_  , \g372467/_3_  , \g372468/_3_  , \g372469/_3_  , \g372470/_3_  , \g372471/_3_  , \g372472/_3_  , \g372473/_3_  , \g372474/_3_  , \g372475/_3_  , \g372476/_3_  , \g372477/_3_  , \g372478/_3_  , \g372479/_3_  , \g372480/_3_  , \g372481/_3_  , \g372482/_3_  , \g372483/_3_  , \g372484/_3_  , \g372485/_3_  , \g372487/_3_  , \g372488/_3_  , \g372489/_3_  , \g372490/_3_  , \g372491/_3_  , \g372492/_3_  , \g372493/_3_  , \g372494/_3_  , \g372495/_3_  , \g372496/_3_  , \g372497/_3_  , \g372498/_3_  , \g372499/_3_  , \g372500/_3_  , \g372501/_3_  , \g372502/_3_  , \g372503/_3_  , \g372504/_3_  , \g372506/_3_  , \g372507/_3_  , \g372508/_3_  , \g372509/_3_  , \g372510/_3_  , \g372511/_3_  , \g372512/_3_  , \g372513/_3_  , \g372514/_3_  , \g372515/_3_  , \g372516/_3_  , \g372517/_3_  , \g372531/_3_  , \g372532/_3_  , \g372533/_3_  , \g374644/_0_  , \g374645/_0_  , \g374648/_0_  , \g374697/_0_  , \g374701/_0_  , \g374749/_0_  , \g374956/_0_  , \g374961/_0_  , \g374965/_0_  , \g374982/_0_  , \g375071/_0_  , \g375073/_0_  , \g375075/_0_  , \g375078/_0_  , \g375315/_3_  , \g375316/_3_  , \g376101/_0_  , \g376479/_0_  , \g377693/_0_  , \g377694/_0_  , \g377695/_0_  , \g377720/_0_  , \g377721/_0_  , \g377722/_0_  , \g378092/_3_  , \g378093/_3_  , \g378094/_3_  , \g378523/_0_  , \g378524/_0_  , \g382190/_0_  , \g382191/_0_  , \g382192/_0_  , \g382193/_0_  , \g382194/_0_  , \g382195/_0_  , \g382279/_0_  , \g382284/_0_  , \g382292/_0_  , \g382299/_0_  , \g382534/_0_  , \g382535/_0_  , \g382555/_0_  , \g382562/_0_  , \g382563/_0_  , \g382564/_0_  , \g382565/_0_  , \g382571/_0_  , \g382773/_3_  , \g382774/_3_  , \g382775/_3_  , \g383503/_2_  , \g383932/_2_  , \g384194/_0_  , \g384195/_0_  , \g384208/_0_  , \g385644/_0_  , \g385649/_0_  , \g385654/_0_  , \g385672/_0_  , \g385812/_0_  , \g385813/_0_  , \g385816/_0_  , \g385819/_0_  , \g386657/_0_  , \g386660/_0_  , \g386710/_0_  , \g386868/_0_  , \g387282/_0_  , \g387284/_0_  , \g387287/_0_  , \g387292/_0_  , \g387559/_0_  , \g387560/_0_  , \g387561/_0_  , \g387562/_0_  , \g387563/_0_  , \g387564/_0_  , \g387735/_0_  , \g387736/_0_  , \g387738/_0_  , \g387739/_0_  , \g387740/_0_  , \g387743/_0_  , \g387788/_0_  , \g387793/_0_  , \g387796/_0_  , \g387803/_0_  , \g388323/_3_  , \g388332/_3_  , \g388543/_0_  , \g388544/_0_  , \g388545/_0_  , \g388547/_0_  , \g388585/_0_  , \g388694/_0_  , \g388830/_0_  , \g388869/_0_  , \g388998/_0_  , \g389009/_0_  , \g389221/_0_  , \g389225/_0_  , \g389226/_0_  , \g389231/_0_  , \g389234/_0_  , \g389242/_0_  , \g389368/_2_  , \g389368/_2__syn_2  , \g389369/_2_  , \g389369/_2__syn_2  , \g389746/_0_  , \g389751/_0_  , \g389774/_0_  , \g389776/_0_  , \g389777/_0_  , \g389779/_0_  , \g389781/_0_  , \g389784/_0_  , \g389787/_0_  , \g389796/_0_  , \g389797/_0_  , \g389801/_0_  , \g390034/_0_  , \g390035/_0_  , \g390037/_0_  , \g390038/_0_  , \g390039/_0_  , \g390043/_0_  , \g390303/_3_  , \g390322/_3_  , \g390323/_3_  , \g390324/_3_  , \g390706/_0_  , \g390876/_0_  , \g390894/_0_  , \g390968/_0_  , \g391050/_0_  , \g391077/_0_  , \g392543/_3_  , \g392565/_3_  , \g392566/_3_  , \g394544/_3_  , \g394545/_3_  , \g394586/_3_  , \g395723/_0_  , \g395757/_0_  , \g395821/_0_  , \g395857/_0_  , \g395858/_0_  , \g395929/_0_  , \g396850/_3_  , \g396876/_3_  , \g396877/_3_  , \g397026/_1_  , \g397035/_1_  , \g397074/_1_  , \g397144/_1_  , \g397344/_1_  , \g397418/_1_  , \g397980/_0_  , \g398209/_0_  , \g398361/_0_  , \g398409/_0_  , \g398458/_0_  , \g398728/_0_  , \g401059/_0_  , \g401066/_0_  , \g401091/_0_  , \g401127/_0_  , \g401160/_0_  , \g401368/_0_  , \g401408/_0_  , \g401455/_0_  , \g401485/_0_  , \g401487/_0_  , \g401506/_0_  , \g401515/_0_  , \g401534/_0_  , \g401549/_0_  , \g401554/_0_  , \g401555/_0_  , \g401592/_0_  , \g401616/_0_  , \g401617/_0_  , \g401618/_0_  , \g401619/_0_  , \g401635/_0_  , \g401657/_0_  , \g401671/_0_  , \g401672/_0_  , \g401684/_0_  , \g401704/_0_  , \g401794/_0_  , \g401807/_0_  , \g401919/_0_  , \g401932/_0_  , \g401935/_0_  , \g401951/_0_  , \g401959/_0_  , \g401961/_0_  , \g401962/_0_  , \g401963/_0_  , \g401998/_0_  , \g402049/_0_  , \g402057/_0_  , \g402063/_0_  , \g402165/_0_  , \g402194/_0_  , \g402298/_0_  , \g402302/_0_  , \g402336/_0_  , \g402346/_0_  , \g402398/_0_  , \g402909/_0_  , \g402910/_0_  , \g402911/_0_  , \g402912/_0_  , \g402913/_0_  , \g402914/_0_  , \g403206/_3_  , \g427842/_1_  , \g427994/_0_  , \g428519/_1_  , \g429040/_1_  , \g429357/_0_  , \g429711/_1_  , \g440733/_0_  , \g440782/_0_  , \g441022/_0_  , \g441242/_0_  , \g441305/_0_  , \g441317/_0_  , \g441329/_0_  , \g441341/_0_  , \g441370/_0_  , \g441382/_0_  , \g441394/_0_  , \g441939/_0_  );
  input \P1_P1_ADS_n_reg/NET0131  ;
  input \P1_P1_Address_reg[0]/NET0131  ;
  input \P1_P1_Address_reg[10]/NET0131  ;
  input \P1_P1_Address_reg[11]/NET0131  ;
  input \P1_P1_Address_reg[12]/NET0131  ;
  input \P1_P1_Address_reg[13]/NET0131  ;
  input \P1_P1_Address_reg[14]/NET0131  ;
  input \P1_P1_Address_reg[15]/NET0131  ;
  input \P1_P1_Address_reg[16]/NET0131  ;
  input \P1_P1_Address_reg[17]/NET0131  ;
  input \P1_P1_Address_reg[18]/NET0131  ;
  input \P1_P1_Address_reg[19]/NET0131  ;
  input \P1_P1_Address_reg[1]/NET0131  ;
  input \P1_P1_Address_reg[20]/NET0131  ;
  input \P1_P1_Address_reg[21]/NET0131  ;
  input \P1_P1_Address_reg[22]/NET0131  ;
  input \P1_P1_Address_reg[23]/NET0131  ;
  input \P1_P1_Address_reg[24]/NET0131  ;
  input \P1_P1_Address_reg[25]/NET0131  ;
  input \P1_P1_Address_reg[26]/NET0131  ;
  input \P1_P1_Address_reg[27]/NET0131  ;
  input \P1_P1_Address_reg[28]/NET0131  ;
  input \P1_P1_Address_reg[29]/NET0131  ;
  input \P1_P1_Address_reg[2]/NET0131  ;
  input \P1_P1_Address_reg[3]/NET0131  ;
  input \P1_P1_Address_reg[4]/NET0131  ;
  input \P1_P1_Address_reg[5]/NET0131  ;
  input \P1_P1_Address_reg[6]/NET0131  ;
  input \P1_P1_Address_reg[7]/NET0131  ;
  input \P1_P1_Address_reg[8]/NET0131  ;
  input \P1_P1_Address_reg[9]/NET0131  ;
  input \P1_P1_BE_n_reg[0]/NET0131  ;
  input \P1_P1_BE_n_reg[1]/NET0131  ;
  input \P1_P1_BE_n_reg[2]/NET0131  ;
  input \P1_P1_BE_n_reg[3]/NET0131  ;
  input \P1_P1_ByteEnable_reg[0]/NET0131  ;
  input \P1_P1_ByteEnable_reg[1]/NET0131  ;
  input \P1_P1_ByteEnable_reg[2]/NET0131  ;
  input \P1_P1_ByteEnable_reg[3]/NET0131  ;
  input \P1_P1_CodeFetch_reg/NET0131  ;
  input \P1_P1_D_C_n_reg/NET0131  ;
  input \P1_P1_DataWidth_reg[0]/NET0131  ;
  input \P1_P1_DataWidth_reg[1]/NET0131  ;
  input \P1_P1_Datao_reg[0]/NET0131  ;
  input \P1_P1_Datao_reg[10]/NET0131  ;
  input \P1_P1_Datao_reg[11]/NET0131  ;
  input \P1_P1_Datao_reg[12]/NET0131  ;
  input \P1_P1_Datao_reg[13]/NET0131  ;
  input \P1_P1_Datao_reg[14]/NET0131  ;
  input \P1_P1_Datao_reg[15]/NET0131  ;
  input \P1_P1_Datao_reg[16]/NET0131  ;
  input \P1_P1_Datao_reg[17]/NET0131  ;
  input \P1_P1_Datao_reg[18]/NET0131  ;
  input \P1_P1_Datao_reg[19]/NET0131  ;
  input \P1_P1_Datao_reg[1]/NET0131  ;
  input \P1_P1_Datao_reg[20]/NET0131  ;
  input \P1_P1_Datao_reg[21]/NET0131  ;
  input \P1_P1_Datao_reg[22]/NET0131  ;
  input \P1_P1_Datao_reg[23]/NET0131  ;
  input \P1_P1_Datao_reg[24]/NET0131  ;
  input \P1_P1_Datao_reg[25]/NET0131  ;
  input \P1_P1_Datao_reg[26]/NET0131  ;
  input \P1_P1_Datao_reg[27]/NET0131  ;
  input \P1_P1_Datao_reg[28]/NET0131  ;
  input \P1_P1_Datao_reg[29]/NET0131  ;
  input \P1_P1_Datao_reg[2]/NET0131  ;
  input \P1_P1_Datao_reg[30]/NET0131  ;
  input \P1_P1_Datao_reg[3]/NET0131  ;
  input \P1_P1_Datao_reg[4]/NET0131  ;
  input \P1_P1_Datao_reg[5]/NET0131  ;
  input \P1_P1_Datao_reg[6]/NET0131  ;
  input \P1_P1_Datao_reg[7]/NET0131  ;
  input \P1_P1_Datao_reg[8]/NET0131  ;
  input \P1_P1_Datao_reg[9]/NET0131  ;
  input \P1_P1_EAX_reg[0]/NET0131  ;
  input \P1_P1_EAX_reg[10]/NET0131  ;
  input \P1_P1_EAX_reg[11]/NET0131  ;
  input \P1_P1_EAX_reg[12]/NET0131  ;
  input \P1_P1_EAX_reg[13]/NET0131  ;
  input \P1_P1_EAX_reg[14]/NET0131  ;
  input \P1_P1_EAX_reg[15]/NET0131  ;
  input \P1_P1_EAX_reg[16]/NET0131  ;
  input \P1_P1_EAX_reg[17]/NET0131  ;
  input \P1_P1_EAX_reg[18]/NET0131  ;
  input \P1_P1_EAX_reg[19]/NET0131  ;
  input \P1_P1_EAX_reg[1]/NET0131  ;
  input \P1_P1_EAX_reg[20]/NET0131  ;
  input \P1_P1_EAX_reg[21]/NET0131  ;
  input \P1_P1_EAX_reg[22]/NET0131  ;
  input \P1_P1_EAX_reg[23]/NET0131  ;
  input \P1_P1_EAX_reg[24]/NET0131  ;
  input \P1_P1_EAX_reg[25]/NET0131  ;
  input \P1_P1_EAX_reg[26]/NET0131  ;
  input \P1_P1_EAX_reg[27]/NET0131  ;
  input \P1_P1_EAX_reg[28]/NET0131  ;
  input \P1_P1_EAX_reg[29]/NET0131  ;
  input \P1_P1_EAX_reg[2]/NET0131  ;
  input \P1_P1_EAX_reg[30]/NET0131  ;
  input \P1_P1_EAX_reg[31]/NET0131  ;
  input \P1_P1_EAX_reg[3]/NET0131  ;
  input \P1_P1_EAX_reg[4]/NET0131  ;
  input \P1_P1_EAX_reg[5]/NET0131  ;
  input \P1_P1_EAX_reg[6]/NET0131  ;
  input \P1_P1_EAX_reg[7]/NET0131  ;
  input \P1_P1_EAX_reg[8]/NET0131  ;
  input \P1_P1_EAX_reg[9]/NET0131  ;
  input \P1_P1_EBX_reg[0]/NET0131  ;
  input \P1_P1_EBX_reg[10]/NET0131  ;
  input \P1_P1_EBX_reg[11]/NET0131  ;
  input \P1_P1_EBX_reg[12]/NET0131  ;
  input \P1_P1_EBX_reg[13]/NET0131  ;
  input \P1_P1_EBX_reg[14]/NET0131  ;
  input \P1_P1_EBX_reg[15]/NET0131  ;
  input \P1_P1_EBX_reg[16]/NET0131  ;
  input \P1_P1_EBX_reg[17]/NET0131  ;
  input \P1_P1_EBX_reg[18]/NET0131  ;
  input \P1_P1_EBX_reg[19]/NET0131  ;
  input \P1_P1_EBX_reg[1]/NET0131  ;
  input \P1_P1_EBX_reg[20]/NET0131  ;
  input \P1_P1_EBX_reg[21]/NET0131  ;
  input \P1_P1_EBX_reg[22]/NET0131  ;
  input \P1_P1_EBX_reg[23]/NET0131  ;
  input \P1_P1_EBX_reg[24]/NET0131  ;
  input \P1_P1_EBX_reg[25]/NET0131  ;
  input \P1_P1_EBX_reg[26]/NET0131  ;
  input \P1_P1_EBX_reg[27]/NET0131  ;
  input \P1_P1_EBX_reg[28]/NET0131  ;
  input \P1_P1_EBX_reg[29]/NET0131  ;
  input \P1_P1_EBX_reg[2]/NET0131  ;
  input \P1_P1_EBX_reg[30]/NET0131  ;
  input \P1_P1_EBX_reg[31]/NET0131  ;
  input \P1_P1_EBX_reg[3]/NET0131  ;
  input \P1_P1_EBX_reg[4]/NET0131  ;
  input \P1_P1_EBX_reg[5]/NET0131  ;
  input \P1_P1_EBX_reg[6]/NET0131  ;
  input \P1_P1_EBX_reg[7]/NET0131  ;
  input \P1_P1_EBX_reg[8]/NET0131  ;
  input \P1_P1_EBX_reg[9]/NET0131  ;
  input \P1_P1_Flush_reg/NET0131  ;
  input \P1_P1_InstAddrPointer_reg[0]/NET0131  ;
  input \P1_P1_InstAddrPointer_reg[10]/NET0131  ;
  input \P1_P1_InstAddrPointer_reg[11]/NET0131  ;
  input \P1_P1_InstAddrPointer_reg[12]/NET0131  ;
  input \P1_P1_InstAddrPointer_reg[13]/NET0131  ;
  input \P1_P1_InstAddrPointer_reg[14]/NET0131  ;
  input \P1_P1_InstAddrPointer_reg[15]/NET0131  ;
  input \P1_P1_InstAddrPointer_reg[16]/NET0131  ;
  input \P1_P1_InstAddrPointer_reg[17]/NET0131  ;
  input \P1_P1_InstAddrPointer_reg[18]/NET0131  ;
  input \P1_P1_InstAddrPointer_reg[19]/NET0131  ;
  input \P1_P1_InstAddrPointer_reg[1]/NET0131  ;
  input \P1_P1_InstAddrPointer_reg[20]/NET0131  ;
  input \P1_P1_InstAddrPointer_reg[21]/NET0131  ;
  input \P1_P1_InstAddrPointer_reg[22]/NET0131  ;
  input \P1_P1_InstAddrPointer_reg[23]/NET0131  ;
  input \P1_P1_InstAddrPointer_reg[24]/NET0131  ;
  input \P1_P1_InstAddrPointer_reg[25]/NET0131  ;
  input \P1_P1_InstAddrPointer_reg[26]/NET0131  ;
  input \P1_P1_InstAddrPointer_reg[27]/NET0131  ;
  input \P1_P1_InstAddrPointer_reg[28]/NET0131  ;
  input \P1_P1_InstAddrPointer_reg[29]/NET0131  ;
  input \P1_P1_InstAddrPointer_reg[2]/NET0131  ;
  input \P1_P1_InstAddrPointer_reg[30]/NET0131  ;
  input \P1_P1_InstAddrPointer_reg[31]/NET0131  ;
  input \P1_P1_InstAddrPointer_reg[3]/NET0131  ;
  input \P1_P1_InstAddrPointer_reg[4]/NET0131  ;
  input \P1_P1_InstAddrPointer_reg[5]/NET0131  ;
  input \P1_P1_InstAddrPointer_reg[6]/NET0131  ;
  input \P1_P1_InstAddrPointer_reg[7]/NET0131  ;
  input \P1_P1_InstAddrPointer_reg[8]/NET0131  ;
  input \P1_P1_InstAddrPointer_reg[9]/NET0131  ;
  input \P1_P1_InstQueueRd_Addr_reg[0]/NET0131  ;
  input \P1_P1_InstQueueRd_Addr_reg[1]/NET0131  ;
  input \P1_P1_InstQueueRd_Addr_reg[2]/NET0131  ;
  input \P1_P1_InstQueueRd_Addr_reg[3]/NET0131  ;
  input \P1_P1_InstQueueWr_Addr_reg[0]/NET0131  ;
  input \P1_P1_InstQueueWr_Addr_reg[1]/NET0131  ;
  input \P1_P1_InstQueueWr_Addr_reg[2]/NET0131  ;
  input \P1_P1_InstQueueWr_Addr_reg[3]/NET0131  ;
  input \P1_P1_InstQueue_reg[0][0]/NET0131  ;
  input \P1_P1_InstQueue_reg[0][1]/NET0131  ;
  input \P1_P1_InstQueue_reg[0][2]/NET0131  ;
  input \P1_P1_InstQueue_reg[0][3]/NET0131  ;
  input \P1_P1_InstQueue_reg[0][4]/NET0131  ;
  input \P1_P1_InstQueue_reg[0][5]/NET0131  ;
  input \P1_P1_InstQueue_reg[0][6]/NET0131  ;
  input \P1_P1_InstQueue_reg[0][7]/NET0131  ;
  input \P1_P1_InstQueue_reg[10][0]/NET0131  ;
  input \P1_P1_InstQueue_reg[10][1]/NET0131  ;
  input \P1_P1_InstQueue_reg[10][2]/NET0131  ;
  input \P1_P1_InstQueue_reg[10][3]/NET0131  ;
  input \P1_P1_InstQueue_reg[10][4]/NET0131  ;
  input \P1_P1_InstQueue_reg[10][5]/NET0131  ;
  input \P1_P1_InstQueue_reg[10][6]/NET0131  ;
  input \P1_P1_InstQueue_reg[10][7]/NET0131  ;
  input \P1_P1_InstQueue_reg[11][0]/NET0131  ;
  input \P1_P1_InstQueue_reg[11][1]/NET0131  ;
  input \P1_P1_InstQueue_reg[11][2]/NET0131  ;
  input \P1_P1_InstQueue_reg[11][3]/NET0131  ;
  input \P1_P1_InstQueue_reg[11][4]/NET0131  ;
  input \P1_P1_InstQueue_reg[11][5]/NET0131  ;
  input \P1_P1_InstQueue_reg[11][6]/NET0131  ;
  input \P1_P1_InstQueue_reg[11][7]/NET0131  ;
  input \P1_P1_InstQueue_reg[12][0]/NET0131  ;
  input \P1_P1_InstQueue_reg[12][1]/NET0131  ;
  input \P1_P1_InstQueue_reg[12][2]/NET0131  ;
  input \P1_P1_InstQueue_reg[12][3]/NET0131  ;
  input \P1_P1_InstQueue_reg[12][4]/NET0131  ;
  input \P1_P1_InstQueue_reg[12][5]/NET0131  ;
  input \P1_P1_InstQueue_reg[12][6]/NET0131  ;
  input \P1_P1_InstQueue_reg[12][7]/NET0131  ;
  input \P1_P1_InstQueue_reg[13][0]/NET0131  ;
  input \P1_P1_InstQueue_reg[13][1]/NET0131  ;
  input \P1_P1_InstQueue_reg[13][2]/NET0131  ;
  input \P1_P1_InstQueue_reg[13][3]/NET0131  ;
  input \P1_P1_InstQueue_reg[13][4]/NET0131  ;
  input \P1_P1_InstQueue_reg[13][5]/NET0131  ;
  input \P1_P1_InstQueue_reg[13][6]/NET0131  ;
  input \P1_P1_InstQueue_reg[13][7]/NET0131  ;
  input \P1_P1_InstQueue_reg[14][0]/NET0131  ;
  input \P1_P1_InstQueue_reg[14][1]/NET0131  ;
  input \P1_P1_InstQueue_reg[14][2]/NET0131  ;
  input \P1_P1_InstQueue_reg[14][3]/NET0131  ;
  input \P1_P1_InstQueue_reg[14][4]/NET0131  ;
  input \P1_P1_InstQueue_reg[14][5]/NET0131  ;
  input \P1_P1_InstQueue_reg[14][6]/NET0131  ;
  input \P1_P1_InstQueue_reg[14][7]/NET0131  ;
  input \P1_P1_InstQueue_reg[15][0]/NET0131  ;
  input \P1_P1_InstQueue_reg[15][1]/NET0131  ;
  input \P1_P1_InstQueue_reg[15][2]/NET0131  ;
  input \P1_P1_InstQueue_reg[15][3]/NET0131  ;
  input \P1_P1_InstQueue_reg[15][4]/NET0131  ;
  input \P1_P1_InstQueue_reg[15][5]/NET0131  ;
  input \P1_P1_InstQueue_reg[15][6]/NET0131  ;
  input \P1_P1_InstQueue_reg[15][7]/NET0131  ;
  input \P1_P1_InstQueue_reg[1][0]/NET0131  ;
  input \P1_P1_InstQueue_reg[1][1]/NET0131  ;
  input \P1_P1_InstQueue_reg[1][2]/NET0131  ;
  input \P1_P1_InstQueue_reg[1][3]/NET0131  ;
  input \P1_P1_InstQueue_reg[1][4]/NET0131  ;
  input \P1_P1_InstQueue_reg[1][5]/NET0131  ;
  input \P1_P1_InstQueue_reg[1][6]/NET0131  ;
  input \P1_P1_InstQueue_reg[1][7]/NET0131  ;
  input \P1_P1_InstQueue_reg[2][0]/NET0131  ;
  input \P1_P1_InstQueue_reg[2][1]/NET0131  ;
  input \P1_P1_InstQueue_reg[2][2]/NET0131  ;
  input \P1_P1_InstQueue_reg[2][3]/NET0131  ;
  input \P1_P1_InstQueue_reg[2][4]/NET0131  ;
  input \P1_P1_InstQueue_reg[2][5]/NET0131  ;
  input \P1_P1_InstQueue_reg[2][6]/NET0131  ;
  input \P1_P1_InstQueue_reg[2][7]/NET0131  ;
  input \P1_P1_InstQueue_reg[3][0]/NET0131  ;
  input \P1_P1_InstQueue_reg[3][1]/NET0131  ;
  input \P1_P1_InstQueue_reg[3][2]/NET0131  ;
  input \P1_P1_InstQueue_reg[3][3]/NET0131  ;
  input \P1_P1_InstQueue_reg[3][4]/NET0131  ;
  input \P1_P1_InstQueue_reg[3][5]/NET0131  ;
  input \P1_P1_InstQueue_reg[3][6]/NET0131  ;
  input \P1_P1_InstQueue_reg[3][7]/NET0131  ;
  input \P1_P1_InstQueue_reg[4][0]/NET0131  ;
  input \P1_P1_InstQueue_reg[4][1]/NET0131  ;
  input \P1_P1_InstQueue_reg[4][2]/NET0131  ;
  input \P1_P1_InstQueue_reg[4][3]/NET0131  ;
  input \P1_P1_InstQueue_reg[4][4]/NET0131  ;
  input \P1_P1_InstQueue_reg[4][5]/NET0131  ;
  input \P1_P1_InstQueue_reg[4][6]/NET0131  ;
  input \P1_P1_InstQueue_reg[4][7]/NET0131  ;
  input \P1_P1_InstQueue_reg[5][0]/NET0131  ;
  input \P1_P1_InstQueue_reg[5][1]/NET0131  ;
  input \P1_P1_InstQueue_reg[5][2]/NET0131  ;
  input \P1_P1_InstQueue_reg[5][3]/NET0131  ;
  input \P1_P1_InstQueue_reg[5][4]/NET0131  ;
  input \P1_P1_InstQueue_reg[5][5]/NET0131  ;
  input \P1_P1_InstQueue_reg[5][6]/NET0131  ;
  input \P1_P1_InstQueue_reg[5][7]/NET0131  ;
  input \P1_P1_InstQueue_reg[6][0]/NET0131  ;
  input \P1_P1_InstQueue_reg[6][1]/NET0131  ;
  input \P1_P1_InstQueue_reg[6][2]/NET0131  ;
  input \P1_P1_InstQueue_reg[6][3]/NET0131  ;
  input \P1_P1_InstQueue_reg[6][4]/NET0131  ;
  input \P1_P1_InstQueue_reg[6][5]/NET0131  ;
  input \P1_P1_InstQueue_reg[6][6]/NET0131  ;
  input \P1_P1_InstQueue_reg[6][7]/NET0131  ;
  input \P1_P1_InstQueue_reg[7][0]/NET0131  ;
  input \P1_P1_InstQueue_reg[7][1]/NET0131  ;
  input \P1_P1_InstQueue_reg[7][2]/NET0131  ;
  input \P1_P1_InstQueue_reg[7][3]/NET0131  ;
  input \P1_P1_InstQueue_reg[7][4]/NET0131  ;
  input \P1_P1_InstQueue_reg[7][5]/NET0131  ;
  input \P1_P1_InstQueue_reg[7][6]/NET0131  ;
  input \P1_P1_InstQueue_reg[7][7]/NET0131  ;
  input \P1_P1_InstQueue_reg[8][0]/NET0131  ;
  input \P1_P1_InstQueue_reg[8][1]/NET0131  ;
  input \P1_P1_InstQueue_reg[8][2]/NET0131  ;
  input \P1_P1_InstQueue_reg[8][3]/NET0131  ;
  input \P1_P1_InstQueue_reg[8][4]/NET0131  ;
  input \P1_P1_InstQueue_reg[8][5]/NET0131  ;
  input \P1_P1_InstQueue_reg[8][6]/NET0131  ;
  input \P1_P1_InstQueue_reg[8][7]/NET0131  ;
  input \P1_P1_InstQueue_reg[9][0]/NET0131  ;
  input \P1_P1_InstQueue_reg[9][1]/NET0131  ;
  input \P1_P1_InstQueue_reg[9][2]/NET0131  ;
  input \P1_P1_InstQueue_reg[9][3]/NET0131  ;
  input \P1_P1_InstQueue_reg[9][4]/NET0131  ;
  input \P1_P1_InstQueue_reg[9][5]/NET0131  ;
  input \P1_P1_InstQueue_reg[9][6]/NET0131  ;
  input \P1_P1_InstQueue_reg[9][7]/NET0131  ;
  input \P1_P1_M_IO_n_reg/NET0131  ;
  input \P1_P1_MemoryFetch_reg/NET0131  ;
  input \P1_P1_More_reg/NET0131  ;
  input \P1_P1_PhyAddrPointer_reg[0]/NET0131  ;
  input \P1_P1_PhyAddrPointer_reg[10]/NET0131  ;
  input \P1_P1_PhyAddrPointer_reg[11]/NET0131  ;
  input \P1_P1_PhyAddrPointer_reg[12]/NET0131  ;
  input \P1_P1_PhyAddrPointer_reg[13]/NET0131  ;
  input \P1_P1_PhyAddrPointer_reg[14]/NET0131  ;
  input \P1_P1_PhyAddrPointer_reg[15]/NET0131  ;
  input \P1_P1_PhyAddrPointer_reg[16]/NET0131  ;
  input \P1_P1_PhyAddrPointer_reg[17]/NET0131  ;
  input \P1_P1_PhyAddrPointer_reg[18]/NET0131  ;
  input \P1_P1_PhyAddrPointer_reg[19]/NET0131  ;
  input \P1_P1_PhyAddrPointer_reg[1]/NET0131  ;
  input \P1_P1_PhyAddrPointer_reg[20]/NET0131  ;
  input \P1_P1_PhyAddrPointer_reg[21]/NET0131  ;
  input \P1_P1_PhyAddrPointer_reg[22]/NET0131  ;
  input \P1_P1_PhyAddrPointer_reg[23]/NET0131  ;
  input \P1_P1_PhyAddrPointer_reg[24]/NET0131  ;
  input \P1_P1_PhyAddrPointer_reg[25]/NET0131  ;
  input \P1_P1_PhyAddrPointer_reg[26]/NET0131  ;
  input \P1_P1_PhyAddrPointer_reg[27]/NET0131  ;
  input \P1_P1_PhyAddrPointer_reg[28]/NET0131  ;
  input \P1_P1_PhyAddrPointer_reg[29]/NET0131  ;
  input \P1_P1_PhyAddrPointer_reg[2]/NET0131  ;
  input \P1_P1_PhyAddrPointer_reg[30]/NET0131  ;
  input \P1_P1_PhyAddrPointer_reg[31]/NET0131  ;
  input \P1_P1_PhyAddrPointer_reg[3]/NET0131  ;
  input \P1_P1_PhyAddrPointer_reg[4]/NET0131  ;
  input \P1_P1_PhyAddrPointer_reg[5]/NET0131  ;
  input \P1_P1_PhyAddrPointer_reg[6]/NET0131  ;
  input \P1_P1_PhyAddrPointer_reg[7]/NET0131  ;
  input \P1_P1_PhyAddrPointer_reg[8]/NET0131  ;
  input \P1_P1_PhyAddrPointer_reg[9]/NET0131  ;
  input \P1_P1_ReadRequest_reg/NET0131  ;
  input \P1_P1_RequestPending_reg/NET0131  ;
  input \P1_P1_State2_reg[0]/NET0131  ;
  input \P1_P1_State2_reg[1]/NET0131  ;
  input \P1_P1_State2_reg[2]/NET0131  ;
  input \P1_P1_State2_reg[3]/NET0131  ;
  input \P1_P1_State_reg[0]/NET0131  ;
  input \P1_P1_State_reg[1]/NET0131  ;
  input \P1_P1_State_reg[2]/NET0131  ;
  input \P1_P1_W_R_n_reg/NET0131  ;
  input \P1_P1_lWord_reg[0]/NET0131  ;
  input \P1_P1_lWord_reg[10]/NET0131  ;
  input \P1_P1_lWord_reg[11]/NET0131  ;
  input \P1_P1_lWord_reg[12]/NET0131  ;
  input \P1_P1_lWord_reg[13]/NET0131  ;
  input \P1_P1_lWord_reg[14]/NET0131  ;
  input \P1_P1_lWord_reg[15]/NET0131  ;
  input \P1_P1_lWord_reg[1]/NET0131  ;
  input \P1_P1_lWord_reg[2]/NET0131  ;
  input \P1_P1_lWord_reg[3]/NET0131  ;
  input \P1_P1_lWord_reg[4]/NET0131  ;
  input \P1_P1_lWord_reg[5]/NET0131  ;
  input \P1_P1_lWord_reg[6]/NET0131  ;
  input \P1_P1_lWord_reg[7]/NET0131  ;
  input \P1_P1_lWord_reg[8]/NET0131  ;
  input \P1_P1_lWord_reg[9]/NET0131  ;
  input \P1_P1_rEIP_reg[0]/NET0131  ;
  input \P1_P1_rEIP_reg[10]/NET0131  ;
  input \P1_P1_rEIP_reg[11]/NET0131  ;
  input \P1_P1_rEIP_reg[12]/NET0131  ;
  input \P1_P1_rEIP_reg[13]/NET0131  ;
  input \P1_P1_rEIP_reg[14]/NET0131  ;
  input \P1_P1_rEIP_reg[15]/NET0131  ;
  input \P1_P1_rEIP_reg[16]/NET0131  ;
  input \P1_P1_rEIP_reg[17]/NET0131  ;
  input \P1_P1_rEIP_reg[18]/NET0131  ;
  input \P1_P1_rEIP_reg[19]/NET0131  ;
  input \P1_P1_rEIP_reg[1]/NET0131  ;
  input \P1_P1_rEIP_reg[20]/NET0131  ;
  input \P1_P1_rEIP_reg[21]/NET0131  ;
  input \P1_P1_rEIP_reg[22]/NET0131  ;
  input \P1_P1_rEIP_reg[23]/NET0131  ;
  input \P1_P1_rEIP_reg[24]/NET0131  ;
  input \P1_P1_rEIP_reg[25]/NET0131  ;
  input \P1_P1_rEIP_reg[26]/NET0131  ;
  input \P1_P1_rEIP_reg[27]/NET0131  ;
  input \P1_P1_rEIP_reg[28]/NET0131  ;
  input \P1_P1_rEIP_reg[29]/NET0131  ;
  input \P1_P1_rEIP_reg[2]/NET0131  ;
  input \P1_P1_rEIP_reg[30]/NET0131  ;
  input \P1_P1_rEIP_reg[31]/NET0131  ;
  input \P1_P1_rEIP_reg[3]/NET0131  ;
  input \P1_P1_rEIP_reg[4]/NET0131  ;
  input \P1_P1_rEIP_reg[5]/NET0131  ;
  input \P1_P1_rEIP_reg[6]/NET0131  ;
  input \P1_P1_rEIP_reg[7]/NET0131  ;
  input \P1_P1_rEIP_reg[8]/NET0131  ;
  input \P1_P1_rEIP_reg[9]/NET0131  ;
  input \P1_P1_uWord_reg[0]/NET0131  ;
  input \P1_P1_uWord_reg[10]/NET0131  ;
  input \P1_P1_uWord_reg[11]/NET0131  ;
  input \P1_P1_uWord_reg[12]/NET0131  ;
  input \P1_P1_uWord_reg[13]/NET0131  ;
  input \P1_P1_uWord_reg[14]/NET0131  ;
  input \P1_P1_uWord_reg[1]/NET0131  ;
  input \P1_P1_uWord_reg[2]/NET0131  ;
  input \P1_P1_uWord_reg[3]/NET0131  ;
  input \P1_P1_uWord_reg[4]/NET0131  ;
  input \P1_P1_uWord_reg[5]/NET0131  ;
  input \P1_P1_uWord_reg[6]/NET0131  ;
  input \P1_P1_uWord_reg[7]/NET0131  ;
  input \P1_P1_uWord_reg[8]/NET0131  ;
  input \P1_P1_uWord_reg[9]/NET0131  ;
  input \P1_P2_ADS_n_reg/NET0131  ;
  input \P1_P2_Address_reg[0]/NET0131  ;
  input \P1_P2_Address_reg[10]/NET0131  ;
  input \P1_P2_Address_reg[11]/NET0131  ;
  input \P1_P2_Address_reg[12]/NET0131  ;
  input \P1_P2_Address_reg[13]/NET0131  ;
  input \P1_P2_Address_reg[14]/NET0131  ;
  input \P1_P2_Address_reg[15]/NET0131  ;
  input \P1_P2_Address_reg[16]/NET0131  ;
  input \P1_P2_Address_reg[17]/NET0131  ;
  input \P1_P2_Address_reg[18]/NET0131  ;
  input \P1_P2_Address_reg[19]/NET0131  ;
  input \P1_P2_Address_reg[1]/NET0131  ;
  input \P1_P2_Address_reg[20]/NET0131  ;
  input \P1_P2_Address_reg[21]/NET0131  ;
  input \P1_P2_Address_reg[22]/NET0131  ;
  input \P1_P2_Address_reg[23]/NET0131  ;
  input \P1_P2_Address_reg[24]/NET0131  ;
  input \P1_P2_Address_reg[25]/NET0131  ;
  input \P1_P2_Address_reg[26]/NET0131  ;
  input \P1_P2_Address_reg[27]/NET0131  ;
  input \P1_P2_Address_reg[28]/NET0131  ;
  input \P1_P2_Address_reg[29]/NET0131  ;
  input \P1_P2_Address_reg[2]/NET0131  ;
  input \P1_P2_Address_reg[3]/NET0131  ;
  input \P1_P2_Address_reg[4]/NET0131  ;
  input \P1_P2_Address_reg[5]/NET0131  ;
  input \P1_P2_Address_reg[6]/NET0131  ;
  input \P1_P2_Address_reg[7]/NET0131  ;
  input \P1_P2_Address_reg[8]/NET0131  ;
  input \P1_P2_Address_reg[9]/NET0131  ;
  input \P1_P2_BE_n_reg[0]/NET0131  ;
  input \P1_P2_BE_n_reg[1]/NET0131  ;
  input \P1_P2_BE_n_reg[2]/NET0131  ;
  input \P1_P2_BE_n_reg[3]/NET0131  ;
  input \P1_P2_ByteEnable_reg[0]/NET0131  ;
  input \P1_P2_ByteEnable_reg[1]/NET0131  ;
  input \P1_P2_ByteEnable_reg[2]/NET0131  ;
  input \P1_P2_ByteEnable_reg[3]/NET0131  ;
  input \P1_P2_CodeFetch_reg/NET0131  ;
  input \P1_P2_D_C_n_reg/NET0131  ;
  input \P1_P2_DataWidth_reg[0]/NET0131  ;
  input \P1_P2_DataWidth_reg[1]/NET0131  ;
  input \P1_P2_Datao_reg[0]/NET0131  ;
  input \P1_P2_Datao_reg[10]/NET0131  ;
  input \P1_P2_Datao_reg[11]/NET0131  ;
  input \P1_P2_Datao_reg[12]/NET0131  ;
  input \P1_P2_Datao_reg[13]/NET0131  ;
  input \P1_P2_Datao_reg[14]/NET0131  ;
  input \P1_P2_Datao_reg[15]/NET0131  ;
  input \P1_P2_Datao_reg[16]/NET0131  ;
  input \P1_P2_Datao_reg[17]/NET0131  ;
  input \P1_P2_Datao_reg[18]/NET0131  ;
  input \P1_P2_Datao_reg[19]/NET0131  ;
  input \P1_P2_Datao_reg[1]/NET0131  ;
  input \P1_P2_Datao_reg[20]/NET0131  ;
  input \P1_P2_Datao_reg[21]/NET0131  ;
  input \P1_P2_Datao_reg[22]/NET0131  ;
  input \P1_P2_Datao_reg[23]/NET0131  ;
  input \P1_P2_Datao_reg[24]/NET0131  ;
  input \P1_P2_Datao_reg[25]/NET0131  ;
  input \P1_P2_Datao_reg[26]/NET0131  ;
  input \P1_P2_Datao_reg[27]/NET0131  ;
  input \P1_P2_Datao_reg[28]/NET0131  ;
  input \P1_P2_Datao_reg[29]/NET0131  ;
  input \P1_P2_Datao_reg[2]/NET0131  ;
  input \P1_P2_Datao_reg[30]/NET0131  ;
  input \P1_P2_Datao_reg[3]/NET0131  ;
  input \P1_P2_Datao_reg[4]/NET0131  ;
  input \P1_P2_Datao_reg[5]/NET0131  ;
  input \P1_P2_Datao_reg[6]/NET0131  ;
  input \P1_P2_Datao_reg[7]/NET0131  ;
  input \P1_P2_Datao_reg[8]/NET0131  ;
  input \P1_P2_Datao_reg[9]/NET0131  ;
  input \P1_P2_EAX_reg[0]/NET0131  ;
  input \P1_P2_EAX_reg[10]/NET0131  ;
  input \P1_P2_EAX_reg[11]/NET0131  ;
  input \P1_P2_EAX_reg[12]/NET0131  ;
  input \P1_P2_EAX_reg[13]/NET0131  ;
  input \P1_P2_EAX_reg[14]/NET0131  ;
  input \P1_P2_EAX_reg[15]/NET0131  ;
  input \P1_P2_EAX_reg[16]/NET0131  ;
  input \P1_P2_EAX_reg[17]/NET0131  ;
  input \P1_P2_EAX_reg[18]/NET0131  ;
  input \P1_P2_EAX_reg[19]/NET0131  ;
  input \P1_P2_EAX_reg[1]/NET0131  ;
  input \P1_P2_EAX_reg[20]/NET0131  ;
  input \P1_P2_EAX_reg[21]/NET0131  ;
  input \P1_P2_EAX_reg[22]/NET0131  ;
  input \P1_P2_EAX_reg[23]/NET0131  ;
  input \P1_P2_EAX_reg[24]/NET0131  ;
  input \P1_P2_EAX_reg[25]/NET0131  ;
  input \P1_P2_EAX_reg[26]/NET0131  ;
  input \P1_P2_EAX_reg[27]/NET0131  ;
  input \P1_P2_EAX_reg[28]/NET0131  ;
  input \P1_P2_EAX_reg[29]/NET0131  ;
  input \P1_P2_EAX_reg[2]/NET0131  ;
  input \P1_P2_EAX_reg[30]/NET0131  ;
  input \P1_P2_EAX_reg[31]/NET0131  ;
  input \P1_P2_EAX_reg[3]/NET0131  ;
  input \P1_P2_EAX_reg[4]/NET0131  ;
  input \P1_P2_EAX_reg[5]/NET0131  ;
  input \P1_P2_EAX_reg[6]/NET0131  ;
  input \P1_P2_EAX_reg[7]/NET0131  ;
  input \P1_P2_EAX_reg[8]/NET0131  ;
  input \P1_P2_EAX_reg[9]/NET0131  ;
  input \P1_P2_EBX_reg[0]/NET0131  ;
  input \P1_P2_EBX_reg[10]/NET0131  ;
  input \P1_P2_EBX_reg[11]/NET0131  ;
  input \P1_P2_EBX_reg[12]/NET0131  ;
  input \P1_P2_EBX_reg[13]/NET0131  ;
  input \P1_P2_EBX_reg[14]/NET0131  ;
  input \P1_P2_EBX_reg[15]/NET0131  ;
  input \P1_P2_EBX_reg[16]/NET0131  ;
  input \P1_P2_EBX_reg[17]/NET0131  ;
  input \P1_P2_EBX_reg[18]/NET0131  ;
  input \P1_P2_EBX_reg[19]/NET0131  ;
  input \P1_P2_EBX_reg[1]/NET0131  ;
  input \P1_P2_EBX_reg[20]/NET0131  ;
  input \P1_P2_EBX_reg[21]/NET0131  ;
  input \P1_P2_EBX_reg[22]/NET0131  ;
  input \P1_P2_EBX_reg[23]/NET0131  ;
  input \P1_P2_EBX_reg[24]/NET0131  ;
  input \P1_P2_EBX_reg[25]/NET0131  ;
  input \P1_P2_EBX_reg[26]/NET0131  ;
  input \P1_P2_EBX_reg[27]/NET0131  ;
  input \P1_P2_EBX_reg[28]/NET0131  ;
  input \P1_P2_EBX_reg[29]/NET0131  ;
  input \P1_P2_EBX_reg[2]/NET0131  ;
  input \P1_P2_EBX_reg[30]/NET0131  ;
  input \P1_P2_EBX_reg[31]/NET0131  ;
  input \P1_P2_EBX_reg[3]/NET0131  ;
  input \P1_P2_EBX_reg[4]/NET0131  ;
  input \P1_P2_EBX_reg[5]/NET0131  ;
  input \P1_P2_EBX_reg[6]/NET0131  ;
  input \P1_P2_EBX_reg[7]/NET0131  ;
  input \P1_P2_EBX_reg[8]/NET0131  ;
  input \P1_P2_EBX_reg[9]/NET0131  ;
  input \P1_P2_Flush_reg/NET0131  ;
  input \P1_P2_InstAddrPointer_reg[0]/NET0131  ;
  input \P1_P2_InstAddrPointer_reg[10]/NET0131  ;
  input \P1_P2_InstAddrPointer_reg[11]/NET0131  ;
  input \P1_P2_InstAddrPointer_reg[12]/NET0131  ;
  input \P1_P2_InstAddrPointer_reg[13]/NET0131  ;
  input \P1_P2_InstAddrPointer_reg[14]/NET0131  ;
  input \P1_P2_InstAddrPointer_reg[15]/NET0131  ;
  input \P1_P2_InstAddrPointer_reg[16]/NET0131  ;
  input \P1_P2_InstAddrPointer_reg[17]/NET0131  ;
  input \P1_P2_InstAddrPointer_reg[18]/NET0131  ;
  input \P1_P2_InstAddrPointer_reg[19]/NET0131  ;
  input \P1_P2_InstAddrPointer_reg[1]/NET0131  ;
  input \P1_P2_InstAddrPointer_reg[20]/NET0131  ;
  input \P1_P2_InstAddrPointer_reg[21]/NET0131  ;
  input \P1_P2_InstAddrPointer_reg[22]/NET0131  ;
  input \P1_P2_InstAddrPointer_reg[23]/NET0131  ;
  input \P1_P2_InstAddrPointer_reg[24]/NET0131  ;
  input \P1_P2_InstAddrPointer_reg[25]/NET0131  ;
  input \P1_P2_InstAddrPointer_reg[26]/NET0131  ;
  input \P1_P2_InstAddrPointer_reg[27]/NET0131  ;
  input \P1_P2_InstAddrPointer_reg[28]/NET0131  ;
  input \P1_P2_InstAddrPointer_reg[29]/NET0131  ;
  input \P1_P2_InstAddrPointer_reg[2]/NET0131  ;
  input \P1_P2_InstAddrPointer_reg[30]/NET0131  ;
  input \P1_P2_InstAddrPointer_reg[31]/NET0131  ;
  input \P1_P2_InstAddrPointer_reg[3]/NET0131  ;
  input \P1_P2_InstAddrPointer_reg[4]/NET0131  ;
  input \P1_P2_InstAddrPointer_reg[5]/NET0131  ;
  input \P1_P2_InstAddrPointer_reg[6]/NET0131  ;
  input \P1_P2_InstAddrPointer_reg[7]/NET0131  ;
  input \P1_P2_InstAddrPointer_reg[8]/NET0131  ;
  input \P1_P2_InstAddrPointer_reg[9]/NET0131  ;
  input \P1_P2_InstQueueRd_Addr_reg[0]/NET0131  ;
  input \P1_P2_InstQueueRd_Addr_reg[1]/NET0131  ;
  input \P1_P2_InstQueueRd_Addr_reg[2]/NET0131  ;
  input \P1_P2_InstQueueRd_Addr_reg[3]/NET0131  ;
  input \P1_P2_InstQueueWr_Addr_reg[0]/NET0131  ;
  input \P1_P2_InstQueueWr_Addr_reg[1]/NET0131  ;
  input \P1_P2_InstQueueWr_Addr_reg[2]/NET0131  ;
  input \P1_P2_InstQueueWr_Addr_reg[3]/NET0131  ;
  input \P1_P2_InstQueue_reg[0][0]/NET0131  ;
  input \P1_P2_InstQueue_reg[0][1]/NET0131  ;
  input \P1_P2_InstQueue_reg[0][2]/NET0131  ;
  input \P1_P2_InstQueue_reg[0][3]/NET0131  ;
  input \P1_P2_InstQueue_reg[0][4]/NET0131  ;
  input \P1_P2_InstQueue_reg[0][5]/NET0131  ;
  input \P1_P2_InstQueue_reg[0][6]/NET0131  ;
  input \P1_P2_InstQueue_reg[0][7]/NET0131  ;
  input \P1_P2_InstQueue_reg[10][0]/NET0131  ;
  input \P1_P2_InstQueue_reg[10][1]/NET0131  ;
  input \P1_P2_InstQueue_reg[10][2]/NET0131  ;
  input \P1_P2_InstQueue_reg[10][3]/NET0131  ;
  input \P1_P2_InstQueue_reg[10][4]/NET0131  ;
  input \P1_P2_InstQueue_reg[10][5]/NET0131  ;
  input \P1_P2_InstQueue_reg[10][6]/NET0131  ;
  input \P1_P2_InstQueue_reg[10][7]/NET0131  ;
  input \P1_P2_InstQueue_reg[11][0]/NET0131  ;
  input \P1_P2_InstQueue_reg[11][1]/NET0131  ;
  input \P1_P2_InstQueue_reg[11][2]/NET0131  ;
  input \P1_P2_InstQueue_reg[11][3]/NET0131  ;
  input \P1_P2_InstQueue_reg[11][4]/NET0131  ;
  input \P1_P2_InstQueue_reg[11][5]/NET0131  ;
  input \P1_P2_InstQueue_reg[11][6]/NET0131  ;
  input \P1_P2_InstQueue_reg[11][7]/NET0131  ;
  input \P1_P2_InstQueue_reg[12][0]/NET0131  ;
  input \P1_P2_InstQueue_reg[12][1]/NET0131  ;
  input \P1_P2_InstQueue_reg[12][2]/NET0131  ;
  input \P1_P2_InstQueue_reg[12][3]/NET0131  ;
  input \P1_P2_InstQueue_reg[12][4]/NET0131  ;
  input \P1_P2_InstQueue_reg[12][5]/NET0131  ;
  input \P1_P2_InstQueue_reg[12][6]/NET0131  ;
  input \P1_P2_InstQueue_reg[12][7]/NET0131  ;
  input \P1_P2_InstQueue_reg[13][0]/NET0131  ;
  input \P1_P2_InstQueue_reg[13][1]/NET0131  ;
  input \P1_P2_InstQueue_reg[13][2]/NET0131  ;
  input \P1_P2_InstQueue_reg[13][3]/NET0131  ;
  input \P1_P2_InstQueue_reg[13][4]/NET0131  ;
  input \P1_P2_InstQueue_reg[13][5]/NET0131  ;
  input \P1_P2_InstQueue_reg[13][6]/NET0131  ;
  input \P1_P2_InstQueue_reg[13][7]/NET0131  ;
  input \P1_P2_InstQueue_reg[14][0]/NET0131  ;
  input \P1_P2_InstQueue_reg[14][1]/NET0131  ;
  input \P1_P2_InstQueue_reg[14][2]/NET0131  ;
  input \P1_P2_InstQueue_reg[14][3]/NET0131  ;
  input \P1_P2_InstQueue_reg[14][4]/NET0131  ;
  input \P1_P2_InstQueue_reg[14][5]/NET0131  ;
  input \P1_P2_InstQueue_reg[14][6]/NET0131  ;
  input \P1_P2_InstQueue_reg[14][7]/NET0131  ;
  input \P1_P2_InstQueue_reg[15][0]/NET0131  ;
  input \P1_P2_InstQueue_reg[15][1]/NET0131  ;
  input \P1_P2_InstQueue_reg[15][2]/NET0131  ;
  input \P1_P2_InstQueue_reg[15][3]/NET0131  ;
  input \P1_P2_InstQueue_reg[15][4]/NET0131  ;
  input \P1_P2_InstQueue_reg[15][5]/NET0131  ;
  input \P1_P2_InstQueue_reg[15][6]/NET0131  ;
  input \P1_P2_InstQueue_reg[15][7]/NET0131  ;
  input \P1_P2_InstQueue_reg[1][0]/NET0131  ;
  input \P1_P2_InstQueue_reg[1][1]/NET0131  ;
  input \P1_P2_InstQueue_reg[1][2]/NET0131  ;
  input \P1_P2_InstQueue_reg[1][3]/NET0131  ;
  input \P1_P2_InstQueue_reg[1][4]/NET0131  ;
  input \P1_P2_InstQueue_reg[1][5]/NET0131  ;
  input \P1_P2_InstQueue_reg[1][6]/NET0131  ;
  input \P1_P2_InstQueue_reg[1][7]/NET0131  ;
  input \P1_P2_InstQueue_reg[2][0]/NET0131  ;
  input \P1_P2_InstQueue_reg[2][1]/NET0131  ;
  input \P1_P2_InstQueue_reg[2][2]/NET0131  ;
  input \P1_P2_InstQueue_reg[2][3]/NET0131  ;
  input \P1_P2_InstQueue_reg[2][4]/NET0131  ;
  input \P1_P2_InstQueue_reg[2][5]/NET0131  ;
  input \P1_P2_InstQueue_reg[2][6]/NET0131  ;
  input \P1_P2_InstQueue_reg[2][7]/NET0131  ;
  input \P1_P2_InstQueue_reg[3][0]/NET0131  ;
  input \P1_P2_InstQueue_reg[3][1]/NET0131  ;
  input \P1_P2_InstQueue_reg[3][2]/NET0131  ;
  input \P1_P2_InstQueue_reg[3][3]/NET0131  ;
  input \P1_P2_InstQueue_reg[3][4]/NET0131  ;
  input \P1_P2_InstQueue_reg[3][5]/NET0131  ;
  input \P1_P2_InstQueue_reg[3][6]/NET0131  ;
  input \P1_P2_InstQueue_reg[3][7]/NET0131  ;
  input \P1_P2_InstQueue_reg[4][0]/NET0131  ;
  input \P1_P2_InstQueue_reg[4][1]/NET0131  ;
  input \P1_P2_InstQueue_reg[4][2]/NET0131  ;
  input \P1_P2_InstQueue_reg[4][3]/NET0131  ;
  input \P1_P2_InstQueue_reg[4][4]/NET0131  ;
  input \P1_P2_InstQueue_reg[4][5]/NET0131  ;
  input \P1_P2_InstQueue_reg[4][6]/NET0131  ;
  input \P1_P2_InstQueue_reg[4][7]/NET0131  ;
  input \P1_P2_InstQueue_reg[5][0]/NET0131  ;
  input \P1_P2_InstQueue_reg[5][1]/NET0131  ;
  input \P1_P2_InstQueue_reg[5][2]/NET0131  ;
  input \P1_P2_InstQueue_reg[5][3]/NET0131  ;
  input \P1_P2_InstQueue_reg[5][4]/NET0131  ;
  input \P1_P2_InstQueue_reg[5][5]/NET0131  ;
  input \P1_P2_InstQueue_reg[5][6]/NET0131  ;
  input \P1_P2_InstQueue_reg[5][7]/NET0131  ;
  input \P1_P2_InstQueue_reg[6][0]/NET0131  ;
  input \P1_P2_InstQueue_reg[6][1]/NET0131  ;
  input \P1_P2_InstQueue_reg[6][2]/NET0131  ;
  input \P1_P2_InstQueue_reg[6][3]/NET0131  ;
  input \P1_P2_InstQueue_reg[6][4]/NET0131  ;
  input \P1_P2_InstQueue_reg[6][5]/NET0131  ;
  input \P1_P2_InstQueue_reg[6][6]/NET0131  ;
  input \P1_P2_InstQueue_reg[6][7]/NET0131  ;
  input \P1_P2_InstQueue_reg[7][0]/NET0131  ;
  input \P1_P2_InstQueue_reg[7][1]/NET0131  ;
  input \P1_P2_InstQueue_reg[7][2]/NET0131  ;
  input \P1_P2_InstQueue_reg[7][3]/NET0131  ;
  input \P1_P2_InstQueue_reg[7][4]/NET0131  ;
  input \P1_P2_InstQueue_reg[7][5]/NET0131  ;
  input \P1_P2_InstQueue_reg[7][6]/NET0131  ;
  input \P1_P2_InstQueue_reg[7][7]/NET0131  ;
  input \P1_P2_InstQueue_reg[8][0]/NET0131  ;
  input \P1_P2_InstQueue_reg[8][1]/NET0131  ;
  input \P1_P2_InstQueue_reg[8][2]/NET0131  ;
  input \P1_P2_InstQueue_reg[8][3]/NET0131  ;
  input \P1_P2_InstQueue_reg[8][4]/NET0131  ;
  input \P1_P2_InstQueue_reg[8][5]/NET0131  ;
  input \P1_P2_InstQueue_reg[8][6]/NET0131  ;
  input \P1_P2_InstQueue_reg[8][7]/NET0131  ;
  input \P1_P2_InstQueue_reg[9][0]/NET0131  ;
  input \P1_P2_InstQueue_reg[9][1]/NET0131  ;
  input \P1_P2_InstQueue_reg[9][2]/NET0131  ;
  input \P1_P2_InstQueue_reg[9][3]/NET0131  ;
  input \P1_P2_InstQueue_reg[9][4]/NET0131  ;
  input \P1_P2_InstQueue_reg[9][5]/NET0131  ;
  input \P1_P2_InstQueue_reg[9][6]/NET0131  ;
  input \P1_P2_InstQueue_reg[9][7]/NET0131  ;
  input \P1_P2_M_IO_n_reg/NET0131  ;
  input \P1_P2_MemoryFetch_reg/NET0131  ;
  input \P1_P2_More_reg/NET0131  ;
  input \P1_P2_PhyAddrPointer_reg[0]/NET0131  ;
  input \P1_P2_PhyAddrPointer_reg[10]/NET0131  ;
  input \P1_P2_PhyAddrPointer_reg[11]/NET0131  ;
  input \P1_P2_PhyAddrPointer_reg[12]/NET0131  ;
  input \P1_P2_PhyAddrPointer_reg[13]/NET0131  ;
  input \P1_P2_PhyAddrPointer_reg[14]/NET0131  ;
  input \P1_P2_PhyAddrPointer_reg[15]/NET0131  ;
  input \P1_P2_PhyAddrPointer_reg[16]/NET0131  ;
  input \P1_P2_PhyAddrPointer_reg[17]/NET0131  ;
  input \P1_P2_PhyAddrPointer_reg[18]/NET0131  ;
  input \P1_P2_PhyAddrPointer_reg[19]/NET0131  ;
  input \P1_P2_PhyAddrPointer_reg[1]/NET0131  ;
  input \P1_P2_PhyAddrPointer_reg[20]/NET0131  ;
  input \P1_P2_PhyAddrPointer_reg[21]/NET0131  ;
  input \P1_P2_PhyAddrPointer_reg[22]/NET0131  ;
  input \P1_P2_PhyAddrPointer_reg[23]/NET0131  ;
  input \P1_P2_PhyAddrPointer_reg[24]/NET0131  ;
  input \P1_P2_PhyAddrPointer_reg[25]/NET0131  ;
  input \P1_P2_PhyAddrPointer_reg[26]/NET0131  ;
  input \P1_P2_PhyAddrPointer_reg[27]/NET0131  ;
  input \P1_P2_PhyAddrPointer_reg[28]/NET0131  ;
  input \P1_P2_PhyAddrPointer_reg[29]/NET0131  ;
  input \P1_P2_PhyAddrPointer_reg[2]/NET0131  ;
  input \P1_P2_PhyAddrPointer_reg[30]/NET0131  ;
  input \P1_P2_PhyAddrPointer_reg[31]/NET0131  ;
  input \P1_P2_PhyAddrPointer_reg[3]/NET0131  ;
  input \P1_P2_PhyAddrPointer_reg[4]/NET0131  ;
  input \P1_P2_PhyAddrPointer_reg[5]/NET0131  ;
  input \P1_P2_PhyAddrPointer_reg[6]/NET0131  ;
  input \P1_P2_PhyAddrPointer_reg[7]/NET0131  ;
  input \P1_P2_PhyAddrPointer_reg[8]/NET0131  ;
  input \P1_P2_PhyAddrPointer_reg[9]/NET0131  ;
  input \P1_P2_ReadRequest_reg/NET0131  ;
  input \P1_P2_RequestPending_reg/NET0131  ;
  input \P1_P2_State2_reg[0]/NET0131  ;
  input \P1_P2_State2_reg[1]/NET0131  ;
  input \P1_P2_State2_reg[2]/NET0131  ;
  input \P1_P2_State2_reg[3]/NET0131  ;
  input \P1_P2_State_reg[0]/NET0131  ;
  input \P1_P2_State_reg[1]/NET0131  ;
  input \P1_P2_State_reg[2]/NET0131  ;
  input \P1_P2_W_R_n_reg/NET0131  ;
  input \P1_P2_lWord_reg[0]/NET0131  ;
  input \P1_P2_lWord_reg[10]/NET0131  ;
  input \P1_P2_lWord_reg[11]/NET0131  ;
  input \P1_P2_lWord_reg[12]/NET0131  ;
  input \P1_P2_lWord_reg[13]/NET0131  ;
  input \P1_P2_lWord_reg[14]/NET0131  ;
  input \P1_P2_lWord_reg[15]/NET0131  ;
  input \P1_P2_lWord_reg[1]/NET0131  ;
  input \P1_P2_lWord_reg[2]/NET0131  ;
  input \P1_P2_lWord_reg[3]/NET0131  ;
  input \P1_P2_lWord_reg[4]/NET0131  ;
  input \P1_P2_lWord_reg[5]/NET0131  ;
  input \P1_P2_lWord_reg[6]/NET0131  ;
  input \P1_P2_lWord_reg[7]/NET0131  ;
  input \P1_P2_lWord_reg[8]/NET0131  ;
  input \P1_P2_lWord_reg[9]/NET0131  ;
  input \P1_P2_rEIP_reg[0]/NET0131  ;
  input \P1_P2_rEIP_reg[10]/NET0131  ;
  input \P1_P2_rEIP_reg[11]/NET0131  ;
  input \P1_P2_rEIP_reg[12]/NET0131  ;
  input \P1_P2_rEIP_reg[13]/NET0131  ;
  input \P1_P2_rEIP_reg[14]/NET0131  ;
  input \P1_P2_rEIP_reg[15]/NET0131  ;
  input \P1_P2_rEIP_reg[16]/NET0131  ;
  input \P1_P2_rEIP_reg[17]/NET0131  ;
  input \P1_P2_rEIP_reg[18]/NET0131  ;
  input \P1_P2_rEIP_reg[19]/NET0131  ;
  input \P1_P2_rEIP_reg[1]/NET0131  ;
  input \P1_P2_rEIP_reg[20]/NET0131  ;
  input \P1_P2_rEIP_reg[21]/NET0131  ;
  input \P1_P2_rEIP_reg[22]/NET0131  ;
  input \P1_P2_rEIP_reg[23]/NET0131  ;
  input \P1_P2_rEIP_reg[24]/NET0131  ;
  input \P1_P2_rEIP_reg[25]/NET0131  ;
  input \P1_P2_rEIP_reg[26]/NET0131  ;
  input \P1_P2_rEIP_reg[27]/NET0131  ;
  input \P1_P2_rEIP_reg[28]/NET0131  ;
  input \P1_P2_rEIP_reg[29]/NET0131  ;
  input \P1_P2_rEIP_reg[2]/NET0131  ;
  input \P1_P2_rEIP_reg[30]/NET0131  ;
  input \P1_P2_rEIP_reg[31]/NET0131  ;
  input \P1_P2_rEIP_reg[3]/NET0131  ;
  input \P1_P2_rEIP_reg[4]/NET0131  ;
  input \P1_P2_rEIP_reg[5]/NET0131  ;
  input \P1_P2_rEIP_reg[6]/NET0131  ;
  input \P1_P2_rEIP_reg[7]/NET0131  ;
  input \P1_P2_rEIP_reg[8]/NET0131  ;
  input \P1_P2_rEIP_reg[9]/NET0131  ;
  input \P1_P2_uWord_reg[0]/NET0131  ;
  input \P1_P2_uWord_reg[10]/NET0131  ;
  input \P1_P2_uWord_reg[11]/NET0131  ;
  input \P1_P2_uWord_reg[12]/NET0131  ;
  input \P1_P2_uWord_reg[13]/NET0131  ;
  input \P1_P2_uWord_reg[14]/NET0131  ;
  input \P1_P2_uWord_reg[1]/NET0131  ;
  input \P1_P2_uWord_reg[2]/NET0131  ;
  input \P1_P2_uWord_reg[3]/NET0131  ;
  input \P1_P2_uWord_reg[4]/NET0131  ;
  input \P1_P2_uWord_reg[5]/NET0131  ;
  input \P1_P2_uWord_reg[6]/NET0131  ;
  input \P1_P2_uWord_reg[7]/NET0131  ;
  input \P1_P2_uWord_reg[8]/NET0131  ;
  input \P1_P2_uWord_reg[9]/NET0131  ;
  input \P1_P3_ADS_n_reg/NET0131  ;
  input \P1_P3_Address_reg[0]/NET0131  ;
  input \P1_P3_Address_reg[10]/NET0131  ;
  input \P1_P3_Address_reg[11]/NET0131  ;
  input \P1_P3_Address_reg[12]/NET0131  ;
  input \P1_P3_Address_reg[13]/NET0131  ;
  input \P1_P3_Address_reg[14]/NET0131  ;
  input \P1_P3_Address_reg[15]/NET0131  ;
  input \P1_P3_Address_reg[16]/NET0131  ;
  input \P1_P3_Address_reg[17]/NET0131  ;
  input \P1_P3_Address_reg[18]/NET0131  ;
  input \P1_P3_Address_reg[1]/NET0131  ;
  input \P1_P3_Address_reg[2]/NET0131  ;
  input \P1_P3_Address_reg[3]/NET0131  ;
  input \P1_P3_Address_reg[4]/NET0131  ;
  input \P1_P3_Address_reg[5]/NET0131  ;
  input \P1_P3_Address_reg[6]/NET0131  ;
  input \P1_P3_Address_reg[7]/NET0131  ;
  input \P1_P3_Address_reg[8]/NET0131  ;
  input \P1_P3_Address_reg[9]/NET0131  ;
  input \P1_P3_BE_n_reg[0]/NET0131  ;
  input \P1_P3_BE_n_reg[1]/NET0131  ;
  input \P1_P3_BE_n_reg[2]/NET0131  ;
  input \P1_P3_BE_n_reg[3]/NET0131  ;
  input \P1_P3_ByteEnable_reg[0]/NET0131  ;
  input \P1_P3_ByteEnable_reg[1]/NET0131  ;
  input \P1_P3_ByteEnable_reg[2]/NET0131  ;
  input \P1_P3_ByteEnable_reg[3]/NET0131  ;
  input \P1_P3_CodeFetch_reg/NET0131  ;
  input \P1_P3_D_C_n_reg/NET0131  ;
  input \P1_P3_DataWidth_reg[0]/NET0131  ;
  input \P1_P3_DataWidth_reg[1]/NET0131  ;
  input \P1_P3_Datao_reg[30]/NET0131  ;
  input \P1_P3_EAX_reg[0]/NET0131  ;
  input \P1_P3_EAX_reg[10]/NET0131  ;
  input \P1_P3_EAX_reg[11]/NET0131  ;
  input \P1_P3_EAX_reg[12]/NET0131  ;
  input \P1_P3_EAX_reg[13]/NET0131  ;
  input \P1_P3_EAX_reg[14]/NET0131  ;
  input \P1_P3_EAX_reg[15]/NET0131  ;
  input \P1_P3_EAX_reg[16]/NET0131  ;
  input \P1_P3_EAX_reg[17]/NET0131  ;
  input \P1_P3_EAX_reg[18]/NET0131  ;
  input \P1_P3_EAX_reg[19]/NET0131  ;
  input \P1_P3_EAX_reg[1]/NET0131  ;
  input \P1_P3_EAX_reg[20]/NET0131  ;
  input \P1_P3_EAX_reg[21]/NET0131  ;
  input \P1_P3_EAX_reg[22]/NET0131  ;
  input \P1_P3_EAX_reg[23]/NET0131  ;
  input \P1_P3_EAX_reg[24]/NET0131  ;
  input \P1_P3_EAX_reg[25]/NET0131  ;
  input \P1_P3_EAX_reg[26]/NET0131  ;
  input \P1_P3_EAX_reg[27]/NET0131  ;
  input \P1_P3_EAX_reg[28]/NET0131  ;
  input \P1_P3_EAX_reg[29]/NET0131  ;
  input \P1_P3_EAX_reg[2]/NET0131  ;
  input \P1_P3_EAX_reg[30]/NET0131  ;
  input \P1_P3_EAX_reg[31]/NET0131  ;
  input \P1_P3_EAX_reg[3]/NET0131  ;
  input \P1_P3_EAX_reg[4]/NET0131  ;
  input \P1_P3_EAX_reg[5]/NET0131  ;
  input \P1_P3_EAX_reg[6]/NET0131  ;
  input \P1_P3_EAX_reg[7]/NET0131  ;
  input \P1_P3_EAX_reg[8]/NET0131  ;
  input \P1_P3_EAX_reg[9]/NET0131  ;
  input \P1_P3_EBX_reg[0]/NET0131  ;
  input \P1_P3_EBX_reg[10]/NET0131  ;
  input \P1_P3_EBX_reg[11]/NET0131  ;
  input \P1_P3_EBX_reg[12]/NET0131  ;
  input \P1_P3_EBX_reg[13]/NET0131  ;
  input \P1_P3_EBX_reg[14]/NET0131  ;
  input \P1_P3_EBX_reg[15]/NET0131  ;
  input \P1_P3_EBX_reg[16]/NET0131  ;
  input \P1_P3_EBX_reg[17]/NET0131  ;
  input \P1_P3_EBX_reg[18]/NET0131  ;
  input \P1_P3_EBX_reg[19]/NET0131  ;
  input \P1_P3_EBX_reg[1]/NET0131  ;
  input \P1_P3_EBX_reg[20]/NET0131  ;
  input \P1_P3_EBX_reg[21]/NET0131  ;
  input \P1_P3_EBX_reg[22]/NET0131  ;
  input \P1_P3_EBX_reg[23]/NET0131  ;
  input \P1_P3_EBX_reg[24]/NET0131  ;
  input \P1_P3_EBX_reg[25]/NET0131  ;
  input \P1_P3_EBX_reg[26]/NET0131  ;
  input \P1_P3_EBX_reg[27]/NET0131  ;
  input \P1_P3_EBX_reg[28]/NET0131  ;
  input \P1_P3_EBX_reg[29]/NET0131  ;
  input \P1_P3_EBX_reg[2]/NET0131  ;
  input \P1_P3_EBX_reg[30]/NET0131  ;
  input \P1_P3_EBX_reg[31]/NET0131  ;
  input \P1_P3_EBX_reg[3]/NET0131  ;
  input \P1_P3_EBX_reg[4]/NET0131  ;
  input \P1_P3_EBX_reg[5]/NET0131  ;
  input \P1_P3_EBX_reg[6]/NET0131  ;
  input \P1_P3_EBX_reg[7]/NET0131  ;
  input \P1_P3_EBX_reg[8]/NET0131  ;
  input \P1_P3_EBX_reg[9]/NET0131  ;
  input \P1_P3_Flush_reg/NET0131  ;
  input \P1_P3_InstAddrPointer_reg[0]/NET0131  ;
  input \P1_P3_InstAddrPointer_reg[10]/NET0131  ;
  input \P1_P3_InstAddrPointer_reg[11]/NET0131  ;
  input \P1_P3_InstAddrPointer_reg[12]/NET0131  ;
  input \P1_P3_InstAddrPointer_reg[13]/NET0131  ;
  input \P1_P3_InstAddrPointer_reg[14]/NET0131  ;
  input \P1_P3_InstAddrPointer_reg[15]/NET0131  ;
  input \P1_P3_InstAddrPointer_reg[16]/NET0131  ;
  input \P1_P3_InstAddrPointer_reg[17]/NET0131  ;
  input \P1_P3_InstAddrPointer_reg[18]/NET0131  ;
  input \P1_P3_InstAddrPointer_reg[19]/NET0131  ;
  input \P1_P3_InstAddrPointer_reg[1]/NET0131  ;
  input \P1_P3_InstAddrPointer_reg[20]/NET0131  ;
  input \P1_P3_InstAddrPointer_reg[21]/NET0131  ;
  input \P1_P3_InstAddrPointer_reg[22]/NET0131  ;
  input \P1_P3_InstAddrPointer_reg[23]/NET0131  ;
  input \P1_P3_InstAddrPointer_reg[24]/NET0131  ;
  input \P1_P3_InstAddrPointer_reg[25]/NET0131  ;
  input \P1_P3_InstAddrPointer_reg[26]/NET0131  ;
  input \P1_P3_InstAddrPointer_reg[27]/NET0131  ;
  input \P1_P3_InstAddrPointer_reg[28]/NET0131  ;
  input \P1_P3_InstAddrPointer_reg[29]/NET0131  ;
  input \P1_P3_InstAddrPointer_reg[2]/NET0131  ;
  input \P1_P3_InstAddrPointer_reg[30]/NET0131  ;
  input \P1_P3_InstAddrPointer_reg[31]/NET0131  ;
  input \P1_P3_InstAddrPointer_reg[3]/NET0131  ;
  input \P1_P3_InstAddrPointer_reg[4]/NET0131  ;
  input \P1_P3_InstAddrPointer_reg[5]/NET0131  ;
  input \P1_P3_InstAddrPointer_reg[6]/NET0131  ;
  input \P1_P3_InstAddrPointer_reg[7]/NET0131  ;
  input \P1_P3_InstAddrPointer_reg[8]/NET0131  ;
  input \P1_P3_InstAddrPointer_reg[9]/NET0131  ;
  input \P1_P3_InstQueueRd_Addr_reg[0]/NET0131  ;
  input \P1_P3_InstQueueRd_Addr_reg[1]/NET0131  ;
  input \P1_P3_InstQueueRd_Addr_reg[2]/NET0131  ;
  input \P1_P3_InstQueueRd_Addr_reg[3]/NET0131  ;
  input \P1_P3_InstQueueWr_Addr_reg[0]/NET0131  ;
  input \P1_P3_InstQueueWr_Addr_reg[1]/NET0131  ;
  input \P1_P3_InstQueueWr_Addr_reg[2]/NET0131  ;
  input \P1_P3_InstQueueWr_Addr_reg[3]/NET0131  ;
  input \P1_P3_InstQueue_reg[0][0]/NET0131  ;
  input \P1_P3_InstQueue_reg[0][1]/NET0131  ;
  input \P1_P3_InstQueue_reg[0][2]/NET0131  ;
  input \P1_P3_InstQueue_reg[0][3]/NET0131  ;
  input \P1_P3_InstQueue_reg[0][4]/NET0131  ;
  input \P1_P3_InstQueue_reg[0][5]/NET0131  ;
  input \P1_P3_InstQueue_reg[0][6]/NET0131  ;
  input \P1_P3_InstQueue_reg[0][7]/NET0131  ;
  input \P1_P3_InstQueue_reg[10][0]/NET0131  ;
  input \P1_P3_InstQueue_reg[10][1]/NET0131  ;
  input \P1_P3_InstQueue_reg[10][2]/NET0131  ;
  input \P1_P3_InstQueue_reg[10][3]/NET0131  ;
  input \P1_P3_InstQueue_reg[10][4]/NET0131  ;
  input \P1_P3_InstQueue_reg[10][5]/NET0131  ;
  input \P1_P3_InstQueue_reg[10][6]/NET0131  ;
  input \P1_P3_InstQueue_reg[10][7]/NET0131  ;
  input \P1_P3_InstQueue_reg[11][0]/NET0131  ;
  input \P1_P3_InstQueue_reg[11][1]/NET0131  ;
  input \P1_P3_InstQueue_reg[11][2]/NET0131  ;
  input \P1_P3_InstQueue_reg[11][3]/NET0131  ;
  input \P1_P3_InstQueue_reg[11][4]/NET0131  ;
  input \P1_P3_InstQueue_reg[11][5]/NET0131  ;
  input \P1_P3_InstQueue_reg[11][6]/NET0131  ;
  input \P1_P3_InstQueue_reg[11][7]/NET0131  ;
  input \P1_P3_InstQueue_reg[12][0]/NET0131  ;
  input \P1_P3_InstQueue_reg[12][1]/NET0131  ;
  input \P1_P3_InstQueue_reg[12][2]/NET0131  ;
  input \P1_P3_InstQueue_reg[12][3]/NET0131  ;
  input \P1_P3_InstQueue_reg[12][4]/NET0131  ;
  input \P1_P3_InstQueue_reg[12][5]/NET0131  ;
  input \P1_P3_InstQueue_reg[12][6]/NET0131  ;
  input \P1_P3_InstQueue_reg[12][7]/NET0131  ;
  input \P1_P3_InstQueue_reg[13][0]/NET0131  ;
  input \P1_P3_InstQueue_reg[13][1]/NET0131  ;
  input \P1_P3_InstQueue_reg[13][2]/NET0131  ;
  input \P1_P3_InstQueue_reg[13][3]/NET0131  ;
  input \P1_P3_InstQueue_reg[13][4]/NET0131  ;
  input \P1_P3_InstQueue_reg[13][5]/NET0131  ;
  input \P1_P3_InstQueue_reg[13][6]/NET0131  ;
  input \P1_P3_InstQueue_reg[13][7]/NET0131  ;
  input \P1_P3_InstQueue_reg[14][0]/NET0131  ;
  input \P1_P3_InstQueue_reg[14][1]/NET0131  ;
  input \P1_P3_InstQueue_reg[14][2]/NET0131  ;
  input \P1_P3_InstQueue_reg[14][3]/NET0131  ;
  input \P1_P3_InstQueue_reg[14][4]/NET0131  ;
  input \P1_P3_InstQueue_reg[14][5]/NET0131  ;
  input \P1_P3_InstQueue_reg[14][6]/NET0131  ;
  input \P1_P3_InstQueue_reg[14][7]/NET0131  ;
  input \P1_P3_InstQueue_reg[15][0]/NET0131  ;
  input \P1_P3_InstQueue_reg[15][1]/NET0131  ;
  input \P1_P3_InstQueue_reg[15][2]/NET0131  ;
  input \P1_P3_InstQueue_reg[15][3]/NET0131  ;
  input \P1_P3_InstQueue_reg[15][4]/NET0131  ;
  input \P1_P3_InstQueue_reg[15][5]/NET0131  ;
  input \P1_P3_InstQueue_reg[15][6]/NET0131  ;
  input \P1_P3_InstQueue_reg[15][7]/NET0131  ;
  input \P1_P3_InstQueue_reg[1][0]/NET0131  ;
  input \P1_P3_InstQueue_reg[1][1]/NET0131  ;
  input \P1_P3_InstQueue_reg[1][2]/NET0131  ;
  input \P1_P3_InstQueue_reg[1][3]/NET0131  ;
  input \P1_P3_InstQueue_reg[1][4]/NET0131  ;
  input \P1_P3_InstQueue_reg[1][5]/NET0131  ;
  input \P1_P3_InstQueue_reg[1][6]/NET0131  ;
  input \P1_P3_InstQueue_reg[1][7]/NET0131  ;
  input \P1_P3_InstQueue_reg[2][0]/NET0131  ;
  input \P1_P3_InstQueue_reg[2][1]/NET0131  ;
  input \P1_P3_InstQueue_reg[2][2]/NET0131  ;
  input \P1_P3_InstQueue_reg[2][3]/NET0131  ;
  input \P1_P3_InstQueue_reg[2][4]/NET0131  ;
  input \P1_P3_InstQueue_reg[2][5]/NET0131  ;
  input \P1_P3_InstQueue_reg[2][6]/NET0131  ;
  input \P1_P3_InstQueue_reg[2][7]/NET0131  ;
  input \P1_P3_InstQueue_reg[3][0]/NET0131  ;
  input \P1_P3_InstQueue_reg[3][1]/NET0131  ;
  input \P1_P3_InstQueue_reg[3][2]/NET0131  ;
  input \P1_P3_InstQueue_reg[3][3]/NET0131  ;
  input \P1_P3_InstQueue_reg[3][4]/NET0131  ;
  input \P1_P3_InstQueue_reg[3][5]/NET0131  ;
  input \P1_P3_InstQueue_reg[3][6]/NET0131  ;
  input \P1_P3_InstQueue_reg[3][7]/NET0131  ;
  input \P1_P3_InstQueue_reg[4][0]/NET0131  ;
  input \P1_P3_InstQueue_reg[4][1]/NET0131  ;
  input \P1_P3_InstQueue_reg[4][2]/NET0131  ;
  input \P1_P3_InstQueue_reg[4][3]/NET0131  ;
  input \P1_P3_InstQueue_reg[4][4]/NET0131  ;
  input \P1_P3_InstQueue_reg[4][5]/NET0131  ;
  input \P1_P3_InstQueue_reg[4][6]/NET0131  ;
  input \P1_P3_InstQueue_reg[4][7]/NET0131  ;
  input \P1_P3_InstQueue_reg[5][0]/NET0131  ;
  input \P1_P3_InstQueue_reg[5][1]/NET0131  ;
  input \P1_P3_InstQueue_reg[5][2]/NET0131  ;
  input \P1_P3_InstQueue_reg[5][3]/NET0131  ;
  input \P1_P3_InstQueue_reg[5][4]/NET0131  ;
  input \P1_P3_InstQueue_reg[5][5]/NET0131  ;
  input \P1_P3_InstQueue_reg[5][6]/NET0131  ;
  input \P1_P3_InstQueue_reg[5][7]/NET0131  ;
  input \P1_P3_InstQueue_reg[6][0]/NET0131  ;
  input \P1_P3_InstQueue_reg[6][1]/NET0131  ;
  input \P1_P3_InstQueue_reg[6][2]/NET0131  ;
  input \P1_P3_InstQueue_reg[6][3]/NET0131  ;
  input \P1_P3_InstQueue_reg[6][4]/NET0131  ;
  input \P1_P3_InstQueue_reg[6][5]/NET0131  ;
  input \P1_P3_InstQueue_reg[6][6]/NET0131  ;
  input \P1_P3_InstQueue_reg[6][7]/NET0131  ;
  input \P1_P3_InstQueue_reg[7][0]/NET0131  ;
  input \P1_P3_InstQueue_reg[7][1]/NET0131  ;
  input \P1_P3_InstQueue_reg[7][2]/NET0131  ;
  input \P1_P3_InstQueue_reg[7][3]/NET0131  ;
  input \P1_P3_InstQueue_reg[7][4]/NET0131  ;
  input \P1_P3_InstQueue_reg[7][5]/NET0131  ;
  input \P1_P3_InstQueue_reg[7][6]/NET0131  ;
  input \P1_P3_InstQueue_reg[7][7]/NET0131  ;
  input \P1_P3_InstQueue_reg[8][0]/NET0131  ;
  input \P1_P3_InstQueue_reg[8][1]/NET0131  ;
  input \P1_P3_InstQueue_reg[8][2]/NET0131  ;
  input \P1_P3_InstQueue_reg[8][3]/NET0131  ;
  input \P1_P3_InstQueue_reg[8][4]/NET0131  ;
  input \P1_P3_InstQueue_reg[8][5]/NET0131  ;
  input \P1_P3_InstQueue_reg[8][6]/NET0131  ;
  input \P1_P3_InstQueue_reg[8][7]/NET0131  ;
  input \P1_P3_InstQueue_reg[9][0]/NET0131  ;
  input \P1_P3_InstQueue_reg[9][1]/NET0131  ;
  input \P1_P3_InstQueue_reg[9][2]/NET0131  ;
  input \P1_P3_InstQueue_reg[9][3]/NET0131  ;
  input \P1_P3_InstQueue_reg[9][4]/NET0131  ;
  input \P1_P3_InstQueue_reg[9][5]/NET0131  ;
  input \P1_P3_InstQueue_reg[9][6]/NET0131  ;
  input \P1_P3_InstQueue_reg[9][7]/NET0131  ;
  input \P1_P3_M_IO_n_reg/NET0131  ;
  input \P1_P3_MemoryFetch_reg/NET0131  ;
  input \P1_P3_More_reg/NET0131  ;
  input \P1_P3_PhyAddrPointer_reg[0]/NET0131  ;
  input \P1_P3_PhyAddrPointer_reg[10]/NET0131  ;
  input \P1_P3_PhyAddrPointer_reg[11]/NET0131  ;
  input \P1_P3_PhyAddrPointer_reg[12]/NET0131  ;
  input \P1_P3_PhyAddrPointer_reg[13]/NET0131  ;
  input \P1_P3_PhyAddrPointer_reg[14]/NET0131  ;
  input \P1_P3_PhyAddrPointer_reg[15]/NET0131  ;
  input \P1_P3_PhyAddrPointer_reg[16]/NET0131  ;
  input \P1_P3_PhyAddrPointer_reg[17]/NET0131  ;
  input \P1_P3_PhyAddrPointer_reg[18]/NET0131  ;
  input \P1_P3_PhyAddrPointer_reg[19]/NET0131  ;
  input \P1_P3_PhyAddrPointer_reg[1]/NET0131  ;
  input \P1_P3_PhyAddrPointer_reg[20]/NET0131  ;
  input \P1_P3_PhyAddrPointer_reg[21]/NET0131  ;
  input \P1_P3_PhyAddrPointer_reg[22]/NET0131  ;
  input \P1_P3_PhyAddrPointer_reg[23]/NET0131  ;
  input \P1_P3_PhyAddrPointer_reg[24]/NET0131  ;
  input \P1_P3_PhyAddrPointer_reg[25]/NET0131  ;
  input \P1_P3_PhyAddrPointer_reg[26]/NET0131  ;
  input \P1_P3_PhyAddrPointer_reg[27]/NET0131  ;
  input \P1_P3_PhyAddrPointer_reg[28]/NET0131  ;
  input \P1_P3_PhyAddrPointer_reg[29]/NET0131  ;
  input \P1_P3_PhyAddrPointer_reg[2]/NET0131  ;
  input \P1_P3_PhyAddrPointer_reg[30]/NET0131  ;
  input \P1_P3_PhyAddrPointer_reg[31]/NET0131  ;
  input \P1_P3_PhyAddrPointer_reg[3]/NET0131  ;
  input \P1_P3_PhyAddrPointer_reg[4]/NET0131  ;
  input \P1_P3_PhyAddrPointer_reg[5]/NET0131  ;
  input \P1_P3_PhyAddrPointer_reg[6]/NET0131  ;
  input \P1_P3_PhyAddrPointer_reg[7]/NET0131  ;
  input \P1_P3_PhyAddrPointer_reg[8]/NET0131  ;
  input \P1_P3_PhyAddrPointer_reg[9]/NET0131  ;
  input \P1_P3_ReadRequest_reg/NET0131  ;
  input \P1_P3_RequestPending_reg/NET0131  ;
  input \P1_P3_State2_reg[0]/NET0131  ;
  input \P1_P3_State2_reg[1]/NET0131  ;
  input \P1_P3_State2_reg[2]/NET0131  ;
  input \P1_P3_State2_reg[3]/NET0131  ;
  input \P1_P3_State_reg[0]/NET0131  ;
  input \P1_P3_State_reg[1]/NET0131  ;
  input \P1_P3_State_reg[2]/NET0131  ;
  input \P1_P3_W_R_n_reg/NET0131  ;
  input \P1_P3_rEIP_reg[0]/NET0131  ;
  input \P1_P3_rEIP_reg[10]/NET0131  ;
  input \P1_P3_rEIP_reg[11]/NET0131  ;
  input \P1_P3_rEIP_reg[12]/NET0131  ;
  input \P1_P3_rEIP_reg[13]/NET0131  ;
  input \P1_P3_rEIP_reg[14]/NET0131  ;
  input \P1_P3_rEIP_reg[15]/NET0131  ;
  input \P1_P3_rEIP_reg[16]/NET0131  ;
  input \P1_P3_rEIP_reg[17]/NET0131  ;
  input \P1_P3_rEIP_reg[18]/NET0131  ;
  input \P1_P3_rEIP_reg[19]/NET0131  ;
  input \P1_P3_rEIP_reg[1]/NET0131  ;
  input \P1_P3_rEIP_reg[20]/NET0131  ;
  input \P1_P3_rEIP_reg[21]/NET0131  ;
  input \P1_P3_rEIP_reg[22]/NET0131  ;
  input \P1_P3_rEIP_reg[23]/NET0131  ;
  input \P1_P3_rEIP_reg[24]/NET0131  ;
  input \P1_P3_rEIP_reg[25]/NET0131  ;
  input \P1_P3_rEIP_reg[26]/NET0131  ;
  input \P1_P3_rEIP_reg[27]/NET0131  ;
  input \P1_P3_rEIP_reg[28]/NET0131  ;
  input \P1_P3_rEIP_reg[29]/NET0131  ;
  input \P1_P3_rEIP_reg[2]/NET0131  ;
  input \P1_P3_rEIP_reg[30]/NET0131  ;
  input \P1_P3_rEIP_reg[31]/NET0131  ;
  input \P1_P3_rEIP_reg[3]/NET0131  ;
  input \P1_P3_rEIP_reg[4]/NET0131  ;
  input \P1_P3_rEIP_reg[5]/NET0131  ;
  input \P1_P3_rEIP_reg[6]/NET0131  ;
  input \P1_P3_rEIP_reg[7]/NET0131  ;
  input \P1_P3_rEIP_reg[8]/NET0131  ;
  input \P1_P3_rEIP_reg[9]/NET0131  ;
  input \P1_P3_uWord_reg[14]/NET0131  ;
  input \P1_buf1_reg[0]/NET0131  ;
  input \P1_buf1_reg[10]/NET0131  ;
  input \P1_buf1_reg[11]/NET0131  ;
  input \P1_buf1_reg[12]/NET0131  ;
  input \P1_buf1_reg[13]/NET0131  ;
  input \P1_buf1_reg[14]/NET0131  ;
  input \P1_buf1_reg[15]/NET0131  ;
  input \P1_buf1_reg[16]/NET0131  ;
  input \P1_buf1_reg[17]/NET0131  ;
  input \P1_buf1_reg[18]/NET0131  ;
  input \P1_buf1_reg[19]/NET0131  ;
  input \P1_buf1_reg[1]/NET0131  ;
  input \P1_buf1_reg[20]/NET0131  ;
  input \P1_buf1_reg[21]/NET0131  ;
  input \P1_buf1_reg[22]/NET0131  ;
  input \P1_buf1_reg[23]/NET0131  ;
  input \P1_buf1_reg[24]/NET0131  ;
  input \P1_buf1_reg[25]/NET0131  ;
  input \P1_buf1_reg[26]/NET0131  ;
  input \P1_buf1_reg[27]/NET0131  ;
  input \P1_buf1_reg[28]/NET0131  ;
  input \P1_buf1_reg[29]/NET0131  ;
  input \P1_buf1_reg[2]/NET0131  ;
  input \P1_buf1_reg[30]/NET0131  ;
  input \P1_buf1_reg[3]/NET0131  ;
  input \P1_buf1_reg[4]/NET0131  ;
  input \P1_buf1_reg[5]/NET0131  ;
  input \P1_buf1_reg[6]/NET0131  ;
  input \P1_buf1_reg[7]/NET0131  ;
  input \P1_buf1_reg[8]/NET0131  ;
  input \P1_buf1_reg[9]/NET0131  ;
  input \P1_buf2_reg[0]/NET0131  ;
  input \P1_buf2_reg[10]/NET0131  ;
  input \P1_buf2_reg[11]/NET0131  ;
  input \P1_buf2_reg[12]/NET0131  ;
  input \P1_buf2_reg[13]/NET0131  ;
  input \P1_buf2_reg[14]/NET0131  ;
  input \P1_buf2_reg[15]/NET0131  ;
  input \P1_buf2_reg[16]/NET0131  ;
  input \P1_buf2_reg[17]/NET0131  ;
  input \P1_buf2_reg[18]/NET0131  ;
  input \P1_buf2_reg[19]/NET0131  ;
  input \P1_buf2_reg[1]/NET0131  ;
  input \P1_buf2_reg[20]/NET0131  ;
  input \P1_buf2_reg[21]/NET0131  ;
  input \P1_buf2_reg[22]/NET0131  ;
  input \P1_buf2_reg[23]/NET0131  ;
  input \P1_buf2_reg[24]/NET0131  ;
  input \P1_buf2_reg[25]/NET0131  ;
  input \P1_buf2_reg[26]/NET0131  ;
  input \P1_buf2_reg[27]/NET0131  ;
  input \P1_buf2_reg[28]/NET0131  ;
  input \P1_buf2_reg[29]/NET0131  ;
  input \P1_buf2_reg[2]/NET0131  ;
  input \P1_buf2_reg[30]/NET0131  ;
  input \P1_buf2_reg[3]/NET0131  ;
  input \P1_buf2_reg[4]/NET0131  ;
  input \P1_buf2_reg[5]/NET0131  ;
  input \P1_buf2_reg[6]/NET0131  ;
  input \P1_buf2_reg[7]/NET0131  ;
  input \P1_buf2_reg[8]/NET0131  ;
  input \P1_buf2_reg[9]/NET0131  ;
  input \P1_ready11_reg/NET0131  ;
  input \P1_ready12_reg/NET0131  ;
  input \P1_ready21_reg/NET0131  ;
  input \P1_ready22_reg/NET0131  ;
  input \P2_P1_ADS_n_reg/NET0131  ;
  input \P2_P1_Address_reg[0]/NET0131  ;
  input \P2_P1_Address_reg[10]/NET0131  ;
  input \P2_P1_Address_reg[11]/NET0131  ;
  input \P2_P1_Address_reg[12]/NET0131  ;
  input \P2_P1_Address_reg[13]/NET0131  ;
  input \P2_P1_Address_reg[14]/NET0131  ;
  input \P2_P1_Address_reg[15]/NET0131  ;
  input \P2_P1_Address_reg[16]/NET0131  ;
  input \P2_P1_Address_reg[17]/NET0131  ;
  input \P2_P1_Address_reg[18]/NET0131  ;
  input \P2_P1_Address_reg[19]/NET0131  ;
  input \P2_P1_Address_reg[1]/NET0131  ;
  input \P2_P1_Address_reg[20]/NET0131  ;
  input \P2_P1_Address_reg[21]/NET0131  ;
  input \P2_P1_Address_reg[22]/NET0131  ;
  input \P2_P1_Address_reg[23]/NET0131  ;
  input \P2_P1_Address_reg[24]/NET0131  ;
  input \P2_P1_Address_reg[25]/NET0131  ;
  input \P2_P1_Address_reg[26]/NET0131  ;
  input \P2_P1_Address_reg[27]/NET0131  ;
  input \P2_P1_Address_reg[28]/NET0131  ;
  input \P2_P1_Address_reg[29]/NET0131  ;
  input \P2_P1_Address_reg[2]/NET0131  ;
  input \P2_P1_Address_reg[3]/NET0131  ;
  input \P2_P1_Address_reg[4]/NET0131  ;
  input \P2_P1_Address_reg[5]/NET0131  ;
  input \P2_P1_Address_reg[6]/NET0131  ;
  input \P2_P1_Address_reg[7]/NET0131  ;
  input \P2_P1_Address_reg[8]/NET0131  ;
  input \P2_P1_Address_reg[9]/NET0131  ;
  input \P2_P1_BE_n_reg[0]/NET0131  ;
  input \P2_P1_BE_n_reg[1]/NET0131  ;
  input \P2_P1_BE_n_reg[2]/NET0131  ;
  input \P2_P1_BE_n_reg[3]/NET0131  ;
  input \P2_P1_ByteEnable_reg[0]/NET0131  ;
  input \P2_P1_ByteEnable_reg[1]/NET0131  ;
  input \P2_P1_ByteEnable_reg[2]/NET0131  ;
  input \P2_P1_ByteEnable_reg[3]/NET0131  ;
  input \P2_P1_CodeFetch_reg/NET0131  ;
  input \P2_P1_D_C_n_reg/NET0131  ;
  input \P2_P1_DataWidth_reg[0]/NET0131  ;
  input \P2_P1_DataWidth_reg[1]/NET0131  ;
  input \P2_P1_Datao_reg[0]/NET0131  ;
  input \P2_P1_Datao_reg[10]/NET0131  ;
  input \P2_P1_Datao_reg[11]/NET0131  ;
  input \P2_P1_Datao_reg[12]/NET0131  ;
  input \P2_P1_Datao_reg[13]/NET0131  ;
  input \P2_P1_Datao_reg[14]/NET0131  ;
  input \P2_P1_Datao_reg[15]/NET0131  ;
  input \P2_P1_Datao_reg[16]/NET0131  ;
  input \P2_P1_Datao_reg[17]/NET0131  ;
  input \P2_P1_Datao_reg[18]/NET0131  ;
  input \P2_P1_Datao_reg[19]/NET0131  ;
  input \P2_P1_Datao_reg[1]/NET0131  ;
  input \P2_P1_Datao_reg[20]/NET0131  ;
  input \P2_P1_Datao_reg[21]/NET0131  ;
  input \P2_P1_Datao_reg[22]/NET0131  ;
  input \P2_P1_Datao_reg[23]/NET0131  ;
  input \P2_P1_Datao_reg[24]/NET0131  ;
  input \P2_P1_Datao_reg[25]/NET0131  ;
  input \P2_P1_Datao_reg[26]/NET0131  ;
  input \P2_P1_Datao_reg[27]/NET0131  ;
  input \P2_P1_Datao_reg[28]/NET0131  ;
  input \P2_P1_Datao_reg[29]/NET0131  ;
  input \P2_P1_Datao_reg[2]/NET0131  ;
  input \P2_P1_Datao_reg[30]/NET0131  ;
  input \P2_P1_Datao_reg[3]/NET0131  ;
  input \P2_P1_Datao_reg[4]/NET0131  ;
  input \P2_P1_Datao_reg[5]/NET0131  ;
  input \P2_P1_Datao_reg[6]/NET0131  ;
  input \P2_P1_Datao_reg[7]/NET0131  ;
  input \P2_P1_Datao_reg[8]/NET0131  ;
  input \P2_P1_Datao_reg[9]/NET0131  ;
  input \P2_P1_EAX_reg[0]/NET0131  ;
  input \P2_P1_EAX_reg[10]/NET0131  ;
  input \P2_P1_EAX_reg[11]/NET0131  ;
  input \P2_P1_EAX_reg[12]/NET0131  ;
  input \P2_P1_EAX_reg[13]/NET0131  ;
  input \P2_P1_EAX_reg[14]/NET0131  ;
  input \P2_P1_EAX_reg[15]/NET0131  ;
  input \P2_P1_EAX_reg[16]/NET0131  ;
  input \P2_P1_EAX_reg[17]/NET0131  ;
  input \P2_P1_EAX_reg[18]/NET0131  ;
  input \P2_P1_EAX_reg[19]/NET0131  ;
  input \P2_P1_EAX_reg[1]/NET0131  ;
  input \P2_P1_EAX_reg[20]/NET0131  ;
  input \P2_P1_EAX_reg[21]/NET0131  ;
  input \P2_P1_EAX_reg[22]/NET0131  ;
  input \P2_P1_EAX_reg[23]/NET0131  ;
  input \P2_P1_EAX_reg[24]/NET0131  ;
  input \P2_P1_EAX_reg[25]/NET0131  ;
  input \P2_P1_EAX_reg[26]/NET0131  ;
  input \P2_P1_EAX_reg[27]/NET0131  ;
  input \P2_P1_EAX_reg[28]/NET0131  ;
  input \P2_P1_EAX_reg[29]/NET0131  ;
  input \P2_P1_EAX_reg[2]/NET0131  ;
  input \P2_P1_EAX_reg[30]/NET0131  ;
  input \P2_P1_EAX_reg[31]/NET0131  ;
  input \P2_P1_EAX_reg[3]/NET0131  ;
  input \P2_P1_EAX_reg[4]/NET0131  ;
  input \P2_P1_EAX_reg[5]/NET0131  ;
  input \P2_P1_EAX_reg[6]/NET0131  ;
  input \P2_P1_EAX_reg[7]/NET0131  ;
  input \P2_P1_EAX_reg[8]/NET0131  ;
  input \P2_P1_EAX_reg[9]/NET0131  ;
  input \P2_P1_EBX_reg[0]/NET0131  ;
  input \P2_P1_EBX_reg[10]/NET0131  ;
  input \P2_P1_EBX_reg[11]/NET0131  ;
  input \P2_P1_EBX_reg[12]/NET0131  ;
  input \P2_P1_EBX_reg[13]/NET0131  ;
  input \P2_P1_EBX_reg[14]/NET0131  ;
  input \P2_P1_EBX_reg[15]/NET0131  ;
  input \P2_P1_EBX_reg[16]/NET0131  ;
  input \P2_P1_EBX_reg[17]/NET0131  ;
  input \P2_P1_EBX_reg[18]/NET0131  ;
  input \P2_P1_EBX_reg[19]/NET0131  ;
  input \P2_P1_EBX_reg[1]/NET0131  ;
  input \P2_P1_EBX_reg[20]/NET0131  ;
  input \P2_P1_EBX_reg[21]/NET0131  ;
  input \P2_P1_EBX_reg[22]/NET0131  ;
  input \P2_P1_EBX_reg[23]/NET0131  ;
  input \P2_P1_EBX_reg[24]/NET0131  ;
  input \P2_P1_EBX_reg[25]/NET0131  ;
  input \P2_P1_EBX_reg[26]/NET0131  ;
  input \P2_P1_EBX_reg[27]/NET0131  ;
  input \P2_P1_EBX_reg[28]/NET0131  ;
  input \P2_P1_EBX_reg[29]/NET0131  ;
  input \P2_P1_EBX_reg[2]/NET0131  ;
  input \P2_P1_EBX_reg[30]/NET0131  ;
  input \P2_P1_EBX_reg[31]/NET0131  ;
  input \P2_P1_EBX_reg[3]/NET0131  ;
  input \P2_P1_EBX_reg[4]/NET0131  ;
  input \P2_P1_EBX_reg[5]/NET0131  ;
  input \P2_P1_EBX_reg[6]/NET0131  ;
  input \P2_P1_EBX_reg[7]/NET0131  ;
  input \P2_P1_EBX_reg[8]/NET0131  ;
  input \P2_P1_EBX_reg[9]/NET0131  ;
  input \P2_P1_Flush_reg/NET0131  ;
  input \P2_P1_InstAddrPointer_reg[0]/NET0131  ;
  input \P2_P1_InstAddrPointer_reg[10]/NET0131  ;
  input \P2_P1_InstAddrPointer_reg[11]/NET0131  ;
  input \P2_P1_InstAddrPointer_reg[12]/NET0131  ;
  input \P2_P1_InstAddrPointer_reg[13]/NET0131  ;
  input \P2_P1_InstAddrPointer_reg[14]/NET0131  ;
  input \P2_P1_InstAddrPointer_reg[15]/NET0131  ;
  input \P2_P1_InstAddrPointer_reg[16]/NET0131  ;
  input \P2_P1_InstAddrPointer_reg[17]/NET0131  ;
  input \P2_P1_InstAddrPointer_reg[18]/NET0131  ;
  input \P2_P1_InstAddrPointer_reg[19]/NET0131  ;
  input \P2_P1_InstAddrPointer_reg[1]/NET0131  ;
  input \P2_P1_InstAddrPointer_reg[20]/NET0131  ;
  input \P2_P1_InstAddrPointer_reg[21]/NET0131  ;
  input \P2_P1_InstAddrPointer_reg[22]/NET0131  ;
  input \P2_P1_InstAddrPointer_reg[23]/NET0131  ;
  input \P2_P1_InstAddrPointer_reg[24]/NET0131  ;
  input \P2_P1_InstAddrPointer_reg[25]/NET0131  ;
  input \P2_P1_InstAddrPointer_reg[26]/NET0131  ;
  input \P2_P1_InstAddrPointer_reg[27]/NET0131  ;
  input \P2_P1_InstAddrPointer_reg[28]/NET0131  ;
  input \P2_P1_InstAddrPointer_reg[29]/NET0131  ;
  input \P2_P1_InstAddrPointer_reg[2]/NET0131  ;
  input \P2_P1_InstAddrPointer_reg[30]/NET0131  ;
  input \P2_P1_InstAddrPointer_reg[31]/NET0131  ;
  input \P2_P1_InstAddrPointer_reg[3]/NET0131  ;
  input \P2_P1_InstAddrPointer_reg[4]/NET0131  ;
  input \P2_P1_InstAddrPointer_reg[5]/NET0131  ;
  input \P2_P1_InstAddrPointer_reg[6]/NET0131  ;
  input \P2_P1_InstAddrPointer_reg[7]/NET0131  ;
  input \P2_P1_InstAddrPointer_reg[8]/NET0131  ;
  input \P2_P1_InstAddrPointer_reg[9]/NET0131  ;
  input \P2_P1_InstQueueRd_Addr_reg[0]/NET0131  ;
  input \P2_P1_InstQueueRd_Addr_reg[1]/NET0131  ;
  input \P2_P1_InstQueueRd_Addr_reg[2]/NET0131  ;
  input \P2_P1_InstQueueRd_Addr_reg[3]/NET0131  ;
  input \P2_P1_InstQueueWr_Addr_reg[0]/NET0131  ;
  input \P2_P1_InstQueueWr_Addr_reg[1]/NET0131  ;
  input \P2_P1_InstQueueWr_Addr_reg[2]/NET0131  ;
  input \P2_P1_InstQueueWr_Addr_reg[3]/NET0131  ;
  input \P2_P1_InstQueue_reg[0][0]/NET0131  ;
  input \P2_P1_InstQueue_reg[0][1]/NET0131  ;
  input \P2_P1_InstQueue_reg[0][2]/NET0131  ;
  input \P2_P1_InstQueue_reg[0][3]/NET0131  ;
  input \P2_P1_InstQueue_reg[0][4]/NET0131  ;
  input \P2_P1_InstQueue_reg[0][5]/NET0131  ;
  input \P2_P1_InstQueue_reg[0][6]/NET0131  ;
  input \P2_P1_InstQueue_reg[0][7]/NET0131  ;
  input \P2_P1_InstQueue_reg[10][0]/NET0131  ;
  input \P2_P1_InstQueue_reg[10][1]/NET0131  ;
  input \P2_P1_InstQueue_reg[10][2]/NET0131  ;
  input \P2_P1_InstQueue_reg[10][3]/NET0131  ;
  input \P2_P1_InstQueue_reg[10][4]/NET0131  ;
  input \P2_P1_InstQueue_reg[10][5]/NET0131  ;
  input \P2_P1_InstQueue_reg[10][6]/NET0131  ;
  input \P2_P1_InstQueue_reg[10][7]/NET0131  ;
  input \P2_P1_InstQueue_reg[11][0]/NET0131  ;
  input \P2_P1_InstQueue_reg[11][1]/NET0131  ;
  input \P2_P1_InstQueue_reg[11][2]/NET0131  ;
  input \P2_P1_InstQueue_reg[11][3]/NET0131  ;
  input \P2_P1_InstQueue_reg[11][4]/NET0131  ;
  input \P2_P1_InstQueue_reg[11][5]/NET0131  ;
  input \P2_P1_InstQueue_reg[11][6]/NET0131  ;
  input \P2_P1_InstQueue_reg[11][7]/NET0131  ;
  input \P2_P1_InstQueue_reg[12][0]/NET0131  ;
  input \P2_P1_InstQueue_reg[12][1]/NET0131  ;
  input \P2_P1_InstQueue_reg[12][2]/NET0131  ;
  input \P2_P1_InstQueue_reg[12][3]/NET0131  ;
  input \P2_P1_InstQueue_reg[12][4]/NET0131  ;
  input \P2_P1_InstQueue_reg[12][5]/NET0131  ;
  input \P2_P1_InstQueue_reg[12][6]/NET0131  ;
  input \P2_P1_InstQueue_reg[12][7]/NET0131  ;
  input \P2_P1_InstQueue_reg[13][0]/NET0131  ;
  input \P2_P1_InstQueue_reg[13][1]/NET0131  ;
  input \P2_P1_InstQueue_reg[13][2]/NET0131  ;
  input \P2_P1_InstQueue_reg[13][3]/NET0131  ;
  input \P2_P1_InstQueue_reg[13][4]/NET0131  ;
  input \P2_P1_InstQueue_reg[13][5]/NET0131  ;
  input \P2_P1_InstQueue_reg[13][6]/NET0131  ;
  input \P2_P1_InstQueue_reg[13][7]/NET0131  ;
  input \P2_P1_InstQueue_reg[14][0]/NET0131  ;
  input \P2_P1_InstQueue_reg[14][1]/NET0131  ;
  input \P2_P1_InstQueue_reg[14][2]/NET0131  ;
  input \P2_P1_InstQueue_reg[14][3]/NET0131  ;
  input \P2_P1_InstQueue_reg[14][4]/NET0131  ;
  input \P2_P1_InstQueue_reg[14][5]/NET0131  ;
  input \P2_P1_InstQueue_reg[14][6]/NET0131  ;
  input \P2_P1_InstQueue_reg[14][7]/NET0131  ;
  input \P2_P1_InstQueue_reg[15][0]/NET0131  ;
  input \P2_P1_InstQueue_reg[15][1]/NET0131  ;
  input \P2_P1_InstQueue_reg[15][2]/NET0131  ;
  input \P2_P1_InstQueue_reg[15][3]/NET0131  ;
  input \P2_P1_InstQueue_reg[15][4]/NET0131  ;
  input \P2_P1_InstQueue_reg[15][5]/NET0131  ;
  input \P2_P1_InstQueue_reg[15][6]/NET0131  ;
  input \P2_P1_InstQueue_reg[15][7]/NET0131  ;
  input \P2_P1_InstQueue_reg[1][0]/NET0131  ;
  input \P2_P1_InstQueue_reg[1][1]/NET0131  ;
  input \P2_P1_InstQueue_reg[1][2]/NET0131  ;
  input \P2_P1_InstQueue_reg[1][3]/NET0131  ;
  input \P2_P1_InstQueue_reg[1][4]/NET0131  ;
  input \P2_P1_InstQueue_reg[1][5]/NET0131  ;
  input \P2_P1_InstQueue_reg[1][6]/NET0131  ;
  input \P2_P1_InstQueue_reg[1][7]/NET0131  ;
  input \P2_P1_InstQueue_reg[2][0]/NET0131  ;
  input \P2_P1_InstQueue_reg[2][1]/NET0131  ;
  input \P2_P1_InstQueue_reg[2][2]/NET0131  ;
  input \P2_P1_InstQueue_reg[2][3]/NET0131  ;
  input \P2_P1_InstQueue_reg[2][4]/NET0131  ;
  input \P2_P1_InstQueue_reg[2][5]/NET0131  ;
  input \P2_P1_InstQueue_reg[2][6]/NET0131  ;
  input \P2_P1_InstQueue_reg[2][7]/NET0131  ;
  input \P2_P1_InstQueue_reg[3][0]/NET0131  ;
  input \P2_P1_InstQueue_reg[3][1]/NET0131  ;
  input \P2_P1_InstQueue_reg[3][2]/NET0131  ;
  input \P2_P1_InstQueue_reg[3][3]/NET0131  ;
  input \P2_P1_InstQueue_reg[3][4]/NET0131  ;
  input \P2_P1_InstQueue_reg[3][5]/NET0131  ;
  input \P2_P1_InstQueue_reg[3][6]/NET0131  ;
  input \P2_P1_InstQueue_reg[3][7]/NET0131  ;
  input \P2_P1_InstQueue_reg[4][0]/NET0131  ;
  input \P2_P1_InstQueue_reg[4][1]/NET0131  ;
  input \P2_P1_InstQueue_reg[4][2]/NET0131  ;
  input \P2_P1_InstQueue_reg[4][3]/NET0131  ;
  input \P2_P1_InstQueue_reg[4][4]/NET0131  ;
  input \P2_P1_InstQueue_reg[4][5]/NET0131  ;
  input \P2_P1_InstQueue_reg[4][6]/NET0131  ;
  input \P2_P1_InstQueue_reg[4][7]/NET0131  ;
  input \P2_P1_InstQueue_reg[5][0]/NET0131  ;
  input \P2_P1_InstQueue_reg[5][1]/NET0131  ;
  input \P2_P1_InstQueue_reg[5][2]/NET0131  ;
  input \P2_P1_InstQueue_reg[5][3]/NET0131  ;
  input \P2_P1_InstQueue_reg[5][4]/NET0131  ;
  input \P2_P1_InstQueue_reg[5][5]/NET0131  ;
  input \P2_P1_InstQueue_reg[5][6]/NET0131  ;
  input \P2_P1_InstQueue_reg[5][7]/NET0131  ;
  input \P2_P1_InstQueue_reg[6][0]/NET0131  ;
  input \P2_P1_InstQueue_reg[6][1]/NET0131  ;
  input \P2_P1_InstQueue_reg[6][2]/NET0131  ;
  input \P2_P1_InstQueue_reg[6][3]/NET0131  ;
  input \P2_P1_InstQueue_reg[6][4]/NET0131  ;
  input \P2_P1_InstQueue_reg[6][5]/NET0131  ;
  input \P2_P1_InstQueue_reg[6][6]/NET0131  ;
  input \P2_P1_InstQueue_reg[6][7]/NET0131  ;
  input \P2_P1_InstQueue_reg[7][0]/NET0131  ;
  input \P2_P1_InstQueue_reg[7][1]/NET0131  ;
  input \P2_P1_InstQueue_reg[7][2]/NET0131  ;
  input \P2_P1_InstQueue_reg[7][3]/NET0131  ;
  input \P2_P1_InstQueue_reg[7][4]/NET0131  ;
  input \P2_P1_InstQueue_reg[7][5]/NET0131  ;
  input \P2_P1_InstQueue_reg[7][6]/NET0131  ;
  input \P2_P1_InstQueue_reg[7][7]/NET0131  ;
  input \P2_P1_InstQueue_reg[8][0]/NET0131  ;
  input \P2_P1_InstQueue_reg[8][1]/NET0131  ;
  input \P2_P1_InstQueue_reg[8][2]/NET0131  ;
  input \P2_P1_InstQueue_reg[8][3]/NET0131  ;
  input \P2_P1_InstQueue_reg[8][4]/NET0131  ;
  input \P2_P1_InstQueue_reg[8][5]/NET0131  ;
  input \P2_P1_InstQueue_reg[8][6]/NET0131  ;
  input \P2_P1_InstQueue_reg[8][7]/NET0131  ;
  input \P2_P1_InstQueue_reg[9][0]/NET0131  ;
  input \P2_P1_InstQueue_reg[9][1]/NET0131  ;
  input \P2_P1_InstQueue_reg[9][2]/NET0131  ;
  input \P2_P1_InstQueue_reg[9][3]/NET0131  ;
  input \P2_P1_InstQueue_reg[9][4]/NET0131  ;
  input \P2_P1_InstQueue_reg[9][5]/NET0131  ;
  input \P2_P1_InstQueue_reg[9][6]/NET0131  ;
  input \P2_P1_InstQueue_reg[9][7]/NET0131  ;
  input \P2_P1_M_IO_n_reg/NET0131  ;
  input \P2_P1_MemoryFetch_reg/NET0131  ;
  input \P2_P1_More_reg/NET0131  ;
  input \P2_P1_PhyAddrPointer_reg[0]/NET0131  ;
  input \P2_P1_PhyAddrPointer_reg[10]/NET0131  ;
  input \P2_P1_PhyAddrPointer_reg[11]/NET0131  ;
  input \P2_P1_PhyAddrPointer_reg[12]/NET0131  ;
  input \P2_P1_PhyAddrPointer_reg[13]/NET0131  ;
  input \P2_P1_PhyAddrPointer_reg[14]/NET0131  ;
  input \P2_P1_PhyAddrPointer_reg[15]/NET0131  ;
  input \P2_P1_PhyAddrPointer_reg[16]/NET0131  ;
  input \P2_P1_PhyAddrPointer_reg[17]/NET0131  ;
  input \P2_P1_PhyAddrPointer_reg[18]/NET0131  ;
  input \P2_P1_PhyAddrPointer_reg[19]/NET0131  ;
  input \P2_P1_PhyAddrPointer_reg[1]/NET0131  ;
  input \P2_P1_PhyAddrPointer_reg[20]/NET0131  ;
  input \P2_P1_PhyAddrPointer_reg[21]/NET0131  ;
  input \P2_P1_PhyAddrPointer_reg[22]/NET0131  ;
  input \P2_P1_PhyAddrPointer_reg[23]/NET0131  ;
  input \P2_P1_PhyAddrPointer_reg[24]/NET0131  ;
  input \P2_P1_PhyAddrPointer_reg[25]/NET0131  ;
  input \P2_P1_PhyAddrPointer_reg[26]/NET0131  ;
  input \P2_P1_PhyAddrPointer_reg[27]/NET0131  ;
  input \P2_P1_PhyAddrPointer_reg[28]/NET0131  ;
  input \P2_P1_PhyAddrPointer_reg[29]/NET0131  ;
  input \P2_P1_PhyAddrPointer_reg[2]/NET0131  ;
  input \P2_P1_PhyAddrPointer_reg[30]/NET0131  ;
  input \P2_P1_PhyAddrPointer_reg[31]/NET0131  ;
  input \P2_P1_PhyAddrPointer_reg[3]/NET0131  ;
  input \P2_P1_PhyAddrPointer_reg[4]/NET0131  ;
  input \P2_P1_PhyAddrPointer_reg[5]/NET0131  ;
  input \P2_P1_PhyAddrPointer_reg[6]/NET0131  ;
  input \P2_P1_PhyAddrPointer_reg[7]/NET0131  ;
  input \P2_P1_PhyAddrPointer_reg[8]/NET0131  ;
  input \P2_P1_PhyAddrPointer_reg[9]/NET0131  ;
  input \P2_P1_ReadRequest_reg/NET0131  ;
  input \P2_P1_RequestPending_reg/NET0131  ;
  input \P2_P1_State2_reg[0]/NET0131  ;
  input \P2_P1_State2_reg[1]/NET0131  ;
  input \P2_P1_State2_reg[2]/NET0131  ;
  input \P2_P1_State2_reg[3]/NET0131  ;
  input \P2_P1_State_reg[0]/NET0131  ;
  input \P2_P1_State_reg[1]/NET0131  ;
  input \P2_P1_State_reg[2]/NET0131  ;
  input \P2_P1_W_R_n_reg/NET0131  ;
  input \P2_P1_lWord_reg[0]/NET0131  ;
  input \P2_P1_lWord_reg[10]/NET0131  ;
  input \P2_P1_lWord_reg[11]/NET0131  ;
  input \P2_P1_lWord_reg[12]/NET0131  ;
  input \P2_P1_lWord_reg[13]/NET0131  ;
  input \P2_P1_lWord_reg[14]/NET0131  ;
  input \P2_P1_lWord_reg[15]/NET0131  ;
  input \P2_P1_lWord_reg[1]/NET0131  ;
  input \P2_P1_lWord_reg[2]/NET0131  ;
  input \P2_P1_lWord_reg[3]/NET0131  ;
  input \P2_P1_lWord_reg[4]/NET0131  ;
  input \P2_P1_lWord_reg[5]/NET0131  ;
  input \P2_P1_lWord_reg[6]/NET0131  ;
  input \P2_P1_lWord_reg[7]/NET0131  ;
  input \P2_P1_lWord_reg[8]/NET0131  ;
  input \P2_P1_lWord_reg[9]/NET0131  ;
  input \P2_P1_rEIP_reg[0]/NET0131  ;
  input \P2_P1_rEIP_reg[10]/NET0131  ;
  input \P2_P1_rEIP_reg[11]/NET0131  ;
  input \P2_P1_rEIP_reg[12]/NET0131  ;
  input \P2_P1_rEIP_reg[13]/NET0131  ;
  input \P2_P1_rEIP_reg[14]/NET0131  ;
  input \P2_P1_rEIP_reg[15]/NET0131  ;
  input \P2_P1_rEIP_reg[16]/NET0131  ;
  input \P2_P1_rEIP_reg[17]/NET0131  ;
  input \P2_P1_rEIP_reg[18]/NET0131  ;
  input \P2_P1_rEIP_reg[19]/NET0131  ;
  input \P2_P1_rEIP_reg[1]/NET0131  ;
  input \P2_P1_rEIP_reg[20]/NET0131  ;
  input \P2_P1_rEIP_reg[21]/NET0131  ;
  input \P2_P1_rEIP_reg[22]/NET0131  ;
  input \P2_P1_rEIP_reg[23]/NET0131  ;
  input \P2_P1_rEIP_reg[24]/NET0131  ;
  input \P2_P1_rEIP_reg[25]/NET0131  ;
  input \P2_P1_rEIP_reg[26]/NET0131  ;
  input \P2_P1_rEIP_reg[27]/NET0131  ;
  input \P2_P1_rEIP_reg[28]/NET0131  ;
  input \P2_P1_rEIP_reg[29]/NET0131  ;
  input \P2_P1_rEIP_reg[2]/NET0131  ;
  input \P2_P1_rEIP_reg[30]/NET0131  ;
  input \P2_P1_rEIP_reg[31]/NET0131  ;
  input \P2_P1_rEIP_reg[3]/NET0131  ;
  input \P2_P1_rEIP_reg[4]/NET0131  ;
  input \P2_P1_rEIP_reg[5]/NET0131  ;
  input \P2_P1_rEIP_reg[6]/NET0131  ;
  input \P2_P1_rEIP_reg[7]/NET0131  ;
  input \P2_P1_rEIP_reg[8]/NET0131  ;
  input \P2_P1_rEIP_reg[9]/NET0131  ;
  input \P2_P1_uWord_reg[0]/NET0131  ;
  input \P2_P1_uWord_reg[10]/NET0131  ;
  input \P2_P1_uWord_reg[11]/NET0131  ;
  input \P2_P1_uWord_reg[12]/NET0131  ;
  input \P2_P1_uWord_reg[13]/NET0131  ;
  input \P2_P1_uWord_reg[14]/NET0131  ;
  input \P2_P1_uWord_reg[1]/NET0131  ;
  input \P2_P1_uWord_reg[2]/NET0131  ;
  input \P2_P1_uWord_reg[3]/NET0131  ;
  input \P2_P1_uWord_reg[4]/NET0131  ;
  input \P2_P1_uWord_reg[5]/NET0131  ;
  input \P2_P1_uWord_reg[6]/NET0131  ;
  input \P2_P1_uWord_reg[7]/NET0131  ;
  input \P2_P1_uWord_reg[8]/NET0131  ;
  input \P2_P1_uWord_reg[9]/NET0131  ;
  input \P2_P2_ADS_n_reg/NET0131  ;
  input \P2_P2_Address_reg[0]/NET0131  ;
  input \P2_P2_Address_reg[10]/NET0131  ;
  input \P2_P2_Address_reg[11]/NET0131  ;
  input \P2_P2_Address_reg[12]/NET0131  ;
  input \P2_P2_Address_reg[13]/NET0131  ;
  input \P2_P2_Address_reg[14]/NET0131  ;
  input \P2_P2_Address_reg[15]/NET0131  ;
  input \P2_P2_Address_reg[16]/NET0131  ;
  input \P2_P2_Address_reg[17]/NET0131  ;
  input \P2_P2_Address_reg[18]/NET0131  ;
  input \P2_P2_Address_reg[19]/NET0131  ;
  input \P2_P2_Address_reg[1]/NET0131  ;
  input \P2_P2_Address_reg[20]/NET0131  ;
  input \P2_P2_Address_reg[21]/NET0131  ;
  input \P2_P2_Address_reg[22]/NET0131  ;
  input \P2_P2_Address_reg[23]/NET0131  ;
  input \P2_P2_Address_reg[24]/NET0131  ;
  input \P2_P2_Address_reg[25]/NET0131  ;
  input \P2_P2_Address_reg[26]/NET0131  ;
  input \P2_P2_Address_reg[27]/NET0131  ;
  input \P2_P2_Address_reg[28]/NET0131  ;
  input \P2_P2_Address_reg[29]/NET0131  ;
  input \P2_P2_Address_reg[2]/NET0131  ;
  input \P2_P2_Address_reg[3]/NET0131  ;
  input \P2_P2_Address_reg[4]/NET0131  ;
  input \P2_P2_Address_reg[5]/NET0131  ;
  input \P2_P2_Address_reg[6]/NET0131  ;
  input \P2_P2_Address_reg[7]/NET0131  ;
  input \P2_P2_Address_reg[8]/NET0131  ;
  input \P2_P2_Address_reg[9]/NET0131  ;
  input \P2_P2_BE_n_reg[0]/NET0131  ;
  input \P2_P2_BE_n_reg[1]/NET0131  ;
  input \P2_P2_BE_n_reg[2]/NET0131  ;
  input \P2_P2_BE_n_reg[3]/NET0131  ;
  input \P2_P2_ByteEnable_reg[0]/NET0131  ;
  input \P2_P2_ByteEnable_reg[1]/NET0131  ;
  input \P2_P2_ByteEnable_reg[2]/NET0131  ;
  input \P2_P2_ByteEnable_reg[3]/NET0131  ;
  input \P2_P2_CodeFetch_reg/NET0131  ;
  input \P2_P2_D_C_n_reg/NET0131  ;
  input \P2_P2_DataWidth_reg[0]/NET0131  ;
  input \P2_P2_DataWidth_reg[1]/NET0131  ;
  input \P2_P2_Datao_reg[0]/NET0131  ;
  input \P2_P2_Datao_reg[10]/NET0131  ;
  input \P2_P2_Datao_reg[11]/NET0131  ;
  input \P2_P2_Datao_reg[12]/NET0131  ;
  input \P2_P2_Datao_reg[13]/NET0131  ;
  input \P2_P2_Datao_reg[14]/NET0131  ;
  input \P2_P2_Datao_reg[15]/NET0131  ;
  input \P2_P2_Datao_reg[16]/NET0131  ;
  input \P2_P2_Datao_reg[17]/NET0131  ;
  input \P2_P2_Datao_reg[18]/NET0131  ;
  input \P2_P2_Datao_reg[19]/NET0131  ;
  input \P2_P2_Datao_reg[1]/NET0131  ;
  input \P2_P2_Datao_reg[20]/NET0131  ;
  input \P2_P2_Datao_reg[21]/NET0131  ;
  input \P2_P2_Datao_reg[22]/NET0131  ;
  input \P2_P2_Datao_reg[23]/NET0131  ;
  input \P2_P2_Datao_reg[24]/NET0131  ;
  input \P2_P2_Datao_reg[25]/NET0131  ;
  input \P2_P2_Datao_reg[26]/NET0131  ;
  input \P2_P2_Datao_reg[27]/NET0131  ;
  input \P2_P2_Datao_reg[28]/NET0131  ;
  input \P2_P2_Datao_reg[29]/NET0131  ;
  input \P2_P2_Datao_reg[2]/NET0131  ;
  input \P2_P2_Datao_reg[30]/NET0131  ;
  input \P2_P2_Datao_reg[3]/NET0131  ;
  input \P2_P2_Datao_reg[4]/NET0131  ;
  input \P2_P2_Datao_reg[5]/NET0131  ;
  input \P2_P2_Datao_reg[6]/NET0131  ;
  input \P2_P2_Datao_reg[7]/NET0131  ;
  input \P2_P2_Datao_reg[8]/NET0131  ;
  input \P2_P2_Datao_reg[9]/NET0131  ;
  input \P2_P2_EAX_reg[0]/NET0131  ;
  input \P2_P2_EAX_reg[10]/NET0131  ;
  input \P2_P2_EAX_reg[11]/NET0131  ;
  input \P2_P2_EAX_reg[12]/NET0131  ;
  input \P2_P2_EAX_reg[13]/NET0131  ;
  input \P2_P2_EAX_reg[14]/NET0131  ;
  input \P2_P2_EAX_reg[15]/NET0131  ;
  input \P2_P2_EAX_reg[16]/NET0131  ;
  input \P2_P2_EAX_reg[17]/NET0131  ;
  input \P2_P2_EAX_reg[18]/NET0131  ;
  input \P2_P2_EAX_reg[19]/NET0131  ;
  input \P2_P2_EAX_reg[1]/NET0131  ;
  input \P2_P2_EAX_reg[20]/NET0131  ;
  input \P2_P2_EAX_reg[21]/NET0131  ;
  input \P2_P2_EAX_reg[22]/NET0131  ;
  input \P2_P2_EAX_reg[23]/NET0131  ;
  input \P2_P2_EAX_reg[24]/NET0131  ;
  input \P2_P2_EAX_reg[25]/NET0131  ;
  input \P2_P2_EAX_reg[26]/NET0131  ;
  input \P2_P2_EAX_reg[27]/NET0131  ;
  input \P2_P2_EAX_reg[28]/NET0131  ;
  input \P2_P2_EAX_reg[29]/NET0131  ;
  input \P2_P2_EAX_reg[2]/NET0131  ;
  input \P2_P2_EAX_reg[30]/NET0131  ;
  input \P2_P2_EAX_reg[31]/NET0131  ;
  input \P2_P2_EAX_reg[3]/NET0131  ;
  input \P2_P2_EAX_reg[4]/NET0131  ;
  input \P2_P2_EAX_reg[5]/NET0131  ;
  input \P2_P2_EAX_reg[6]/NET0131  ;
  input \P2_P2_EAX_reg[7]/NET0131  ;
  input \P2_P2_EAX_reg[8]/NET0131  ;
  input \P2_P2_EAX_reg[9]/NET0131  ;
  input \P2_P2_EBX_reg[0]/NET0131  ;
  input \P2_P2_EBX_reg[10]/NET0131  ;
  input \P2_P2_EBX_reg[11]/NET0131  ;
  input \P2_P2_EBX_reg[12]/NET0131  ;
  input \P2_P2_EBX_reg[13]/NET0131  ;
  input \P2_P2_EBX_reg[14]/NET0131  ;
  input \P2_P2_EBX_reg[15]/NET0131  ;
  input \P2_P2_EBX_reg[16]/NET0131  ;
  input \P2_P2_EBX_reg[17]/NET0131  ;
  input \P2_P2_EBX_reg[18]/NET0131  ;
  input \P2_P2_EBX_reg[19]/NET0131  ;
  input \P2_P2_EBX_reg[1]/NET0131  ;
  input \P2_P2_EBX_reg[20]/NET0131  ;
  input \P2_P2_EBX_reg[21]/NET0131  ;
  input \P2_P2_EBX_reg[22]/NET0131  ;
  input \P2_P2_EBX_reg[23]/NET0131  ;
  input \P2_P2_EBX_reg[24]/NET0131  ;
  input \P2_P2_EBX_reg[25]/NET0131  ;
  input \P2_P2_EBX_reg[26]/NET0131  ;
  input \P2_P2_EBX_reg[27]/NET0131  ;
  input \P2_P2_EBX_reg[28]/NET0131  ;
  input \P2_P2_EBX_reg[29]/NET0131  ;
  input \P2_P2_EBX_reg[2]/NET0131  ;
  input \P2_P2_EBX_reg[30]/NET0131  ;
  input \P2_P2_EBX_reg[31]/NET0131  ;
  input \P2_P2_EBX_reg[3]/NET0131  ;
  input \P2_P2_EBX_reg[4]/NET0131  ;
  input \P2_P2_EBX_reg[5]/NET0131  ;
  input \P2_P2_EBX_reg[6]/NET0131  ;
  input \P2_P2_EBX_reg[7]/NET0131  ;
  input \P2_P2_EBX_reg[8]/NET0131  ;
  input \P2_P2_EBX_reg[9]/NET0131  ;
  input \P2_P2_Flush_reg/NET0131  ;
  input \P2_P2_InstAddrPointer_reg[0]/NET0131  ;
  input \P2_P2_InstAddrPointer_reg[10]/NET0131  ;
  input \P2_P2_InstAddrPointer_reg[11]/NET0131  ;
  input \P2_P2_InstAddrPointer_reg[12]/NET0131  ;
  input \P2_P2_InstAddrPointer_reg[13]/NET0131  ;
  input \P2_P2_InstAddrPointer_reg[14]/NET0131  ;
  input \P2_P2_InstAddrPointer_reg[15]/NET0131  ;
  input \P2_P2_InstAddrPointer_reg[16]/NET0131  ;
  input \P2_P2_InstAddrPointer_reg[17]/NET0131  ;
  input \P2_P2_InstAddrPointer_reg[18]/NET0131  ;
  input \P2_P2_InstAddrPointer_reg[19]/NET0131  ;
  input \P2_P2_InstAddrPointer_reg[1]/NET0131  ;
  input \P2_P2_InstAddrPointer_reg[20]/NET0131  ;
  input \P2_P2_InstAddrPointer_reg[21]/NET0131  ;
  input \P2_P2_InstAddrPointer_reg[22]/NET0131  ;
  input \P2_P2_InstAddrPointer_reg[23]/NET0131  ;
  input \P2_P2_InstAddrPointer_reg[24]/NET0131  ;
  input \P2_P2_InstAddrPointer_reg[25]/NET0131  ;
  input \P2_P2_InstAddrPointer_reg[26]/NET0131  ;
  input \P2_P2_InstAddrPointer_reg[27]/NET0131  ;
  input \P2_P2_InstAddrPointer_reg[28]/NET0131  ;
  input \P2_P2_InstAddrPointer_reg[29]/NET0131  ;
  input \P2_P2_InstAddrPointer_reg[2]/NET0131  ;
  input \P2_P2_InstAddrPointer_reg[30]/NET0131  ;
  input \P2_P2_InstAddrPointer_reg[31]/NET0131  ;
  input \P2_P2_InstAddrPointer_reg[3]/NET0131  ;
  input \P2_P2_InstAddrPointer_reg[4]/NET0131  ;
  input \P2_P2_InstAddrPointer_reg[5]/NET0131  ;
  input \P2_P2_InstAddrPointer_reg[6]/NET0131  ;
  input \P2_P2_InstAddrPointer_reg[7]/NET0131  ;
  input \P2_P2_InstAddrPointer_reg[8]/NET0131  ;
  input \P2_P2_InstAddrPointer_reg[9]/NET0131  ;
  input \P2_P2_InstQueueRd_Addr_reg[0]/NET0131  ;
  input \P2_P2_InstQueueRd_Addr_reg[1]/NET0131  ;
  input \P2_P2_InstQueueRd_Addr_reg[2]/NET0131  ;
  input \P2_P2_InstQueueRd_Addr_reg[3]/NET0131  ;
  input \P2_P2_InstQueueWr_Addr_reg[0]/NET0131  ;
  input \P2_P2_InstQueueWr_Addr_reg[1]/NET0131  ;
  input \P2_P2_InstQueueWr_Addr_reg[2]/NET0131  ;
  input \P2_P2_InstQueueWr_Addr_reg[3]/NET0131  ;
  input \P2_P2_InstQueue_reg[0][0]/NET0131  ;
  input \P2_P2_InstQueue_reg[0][1]/NET0131  ;
  input \P2_P2_InstQueue_reg[0][2]/NET0131  ;
  input \P2_P2_InstQueue_reg[0][3]/NET0131  ;
  input \P2_P2_InstQueue_reg[0][4]/NET0131  ;
  input \P2_P2_InstQueue_reg[0][5]/NET0131  ;
  input \P2_P2_InstQueue_reg[0][6]/NET0131  ;
  input \P2_P2_InstQueue_reg[0][7]/NET0131  ;
  input \P2_P2_InstQueue_reg[10][0]/NET0131  ;
  input \P2_P2_InstQueue_reg[10][1]/NET0131  ;
  input \P2_P2_InstQueue_reg[10][2]/NET0131  ;
  input \P2_P2_InstQueue_reg[10][3]/NET0131  ;
  input \P2_P2_InstQueue_reg[10][4]/NET0131  ;
  input \P2_P2_InstQueue_reg[10][5]/NET0131  ;
  input \P2_P2_InstQueue_reg[10][6]/NET0131  ;
  input \P2_P2_InstQueue_reg[10][7]/NET0131  ;
  input \P2_P2_InstQueue_reg[11][0]/NET0131  ;
  input \P2_P2_InstQueue_reg[11][1]/NET0131  ;
  input \P2_P2_InstQueue_reg[11][2]/NET0131  ;
  input \P2_P2_InstQueue_reg[11][3]/NET0131  ;
  input \P2_P2_InstQueue_reg[11][4]/NET0131  ;
  input \P2_P2_InstQueue_reg[11][5]/NET0131  ;
  input \P2_P2_InstQueue_reg[11][6]/NET0131  ;
  input \P2_P2_InstQueue_reg[11][7]/NET0131  ;
  input \P2_P2_InstQueue_reg[12][0]/NET0131  ;
  input \P2_P2_InstQueue_reg[12][1]/NET0131  ;
  input \P2_P2_InstQueue_reg[12][2]/NET0131  ;
  input \P2_P2_InstQueue_reg[12][3]/NET0131  ;
  input \P2_P2_InstQueue_reg[12][4]/NET0131  ;
  input \P2_P2_InstQueue_reg[12][5]/NET0131  ;
  input \P2_P2_InstQueue_reg[12][6]/NET0131  ;
  input \P2_P2_InstQueue_reg[12][7]/NET0131  ;
  input \P2_P2_InstQueue_reg[13][0]/NET0131  ;
  input \P2_P2_InstQueue_reg[13][1]/NET0131  ;
  input \P2_P2_InstQueue_reg[13][2]/NET0131  ;
  input \P2_P2_InstQueue_reg[13][3]/NET0131  ;
  input \P2_P2_InstQueue_reg[13][4]/NET0131  ;
  input \P2_P2_InstQueue_reg[13][5]/NET0131  ;
  input \P2_P2_InstQueue_reg[13][6]/NET0131  ;
  input \P2_P2_InstQueue_reg[13][7]/NET0131  ;
  input \P2_P2_InstQueue_reg[14][0]/NET0131  ;
  input \P2_P2_InstQueue_reg[14][1]/NET0131  ;
  input \P2_P2_InstQueue_reg[14][2]/NET0131  ;
  input \P2_P2_InstQueue_reg[14][3]/NET0131  ;
  input \P2_P2_InstQueue_reg[14][4]/NET0131  ;
  input \P2_P2_InstQueue_reg[14][5]/NET0131  ;
  input \P2_P2_InstQueue_reg[14][6]/NET0131  ;
  input \P2_P2_InstQueue_reg[14][7]/NET0131  ;
  input \P2_P2_InstQueue_reg[15][0]/NET0131  ;
  input \P2_P2_InstQueue_reg[15][1]/NET0131  ;
  input \P2_P2_InstQueue_reg[15][2]/NET0131  ;
  input \P2_P2_InstQueue_reg[15][3]/NET0131  ;
  input \P2_P2_InstQueue_reg[15][4]/NET0131  ;
  input \P2_P2_InstQueue_reg[15][5]/NET0131  ;
  input \P2_P2_InstQueue_reg[15][6]/NET0131  ;
  input \P2_P2_InstQueue_reg[15][7]/NET0131  ;
  input \P2_P2_InstQueue_reg[1][0]/NET0131  ;
  input \P2_P2_InstQueue_reg[1][1]/NET0131  ;
  input \P2_P2_InstQueue_reg[1][2]/NET0131  ;
  input \P2_P2_InstQueue_reg[1][3]/NET0131  ;
  input \P2_P2_InstQueue_reg[1][4]/NET0131  ;
  input \P2_P2_InstQueue_reg[1][5]/NET0131  ;
  input \P2_P2_InstQueue_reg[1][6]/NET0131  ;
  input \P2_P2_InstQueue_reg[1][7]/NET0131  ;
  input \P2_P2_InstQueue_reg[2][0]/NET0131  ;
  input \P2_P2_InstQueue_reg[2][1]/NET0131  ;
  input \P2_P2_InstQueue_reg[2][2]/NET0131  ;
  input \P2_P2_InstQueue_reg[2][3]/NET0131  ;
  input \P2_P2_InstQueue_reg[2][4]/NET0131  ;
  input \P2_P2_InstQueue_reg[2][5]/NET0131  ;
  input \P2_P2_InstQueue_reg[2][6]/NET0131  ;
  input \P2_P2_InstQueue_reg[2][7]/NET0131  ;
  input \P2_P2_InstQueue_reg[3][0]/NET0131  ;
  input \P2_P2_InstQueue_reg[3][1]/NET0131  ;
  input \P2_P2_InstQueue_reg[3][2]/NET0131  ;
  input \P2_P2_InstQueue_reg[3][3]/NET0131  ;
  input \P2_P2_InstQueue_reg[3][4]/NET0131  ;
  input \P2_P2_InstQueue_reg[3][5]/NET0131  ;
  input \P2_P2_InstQueue_reg[3][6]/NET0131  ;
  input \P2_P2_InstQueue_reg[3][7]/NET0131  ;
  input \P2_P2_InstQueue_reg[4][0]/NET0131  ;
  input \P2_P2_InstQueue_reg[4][1]/NET0131  ;
  input \P2_P2_InstQueue_reg[4][2]/NET0131  ;
  input \P2_P2_InstQueue_reg[4][3]/NET0131  ;
  input \P2_P2_InstQueue_reg[4][4]/NET0131  ;
  input \P2_P2_InstQueue_reg[4][5]/NET0131  ;
  input \P2_P2_InstQueue_reg[4][6]/NET0131  ;
  input \P2_P2_InstQueue_reg[4][7]/NET0131  ;
  input \P2_P2_InstQueue_reg[5][0]/NET0131  ;
  input \P2_P2_InstQueue_reg[5][1]/NET0131  ;
  input \P2_P2_InstQueue_reg[5][2]/NET0131  ;
  input \P2_P2_InstQueue_reg[5][3]/NET0131  ;
  input \P2_P2_InstQueue_reg[5][4]/NET0131  ;
  input \P2_P2_InstQueue_reg[5][5]/NET0131  ;
  input \P2_P2_InstQueue_reg[5][6]/NET0131  ;
  input \P2_P2_InstQueue_reg[5][7]/NET0131  ;
  input \P2_P2_InstQueue_reg[6][0]/NET0131  ;
  input \P2_P2_InstQueue_reg[6][1]/NET0131  ;
  input \P2_P2_InstQueue_reg[6][2]/NET0131  ;
  input \P2_P2_InstQueue_reg[6][3]/NET0131  ;
  input \P2_P2_InstQueue_reg[6][4]/NET0131  ;
  input \P2_P2_InstQueue_reg[6][5]/NET0131  ;
  input \P2_P2_InstQueue_reg[6][6]/NET0131  ;
  input \P2_P2_InstQueue_reg[6][7]/NET0131  ;
  input \P2_P2_InstQueue_reg[7][0]/NET0131  ;
  input \P2_P2_InstQueue_reg[7][1]/NET0131  ;
  input \P2_P2_InstQueue_reg[7][2]/NET0131  ;
  input \P2_P2_InstQueue_reg[7][3]/NET0131  ;
  input \P2_P2_InstQueue_reg[7][4]/NET0131  ;
  input \P2_P2_InstQueue_reg[7][5]/NET0131  ;
  input \P2_P2_InstQueue_reg[7][6]/NET0131  ;
  input \P2_P2_InstQueue_reg[7][7]/NET0131  ;
  input \P2_P2_InstQueue_reg[8][0]/NET0131  ;
  input \P2_P2_InstQueue_reg[8][1]/NET0131  ;
  input \P2_P2_InstQueue_reg[8][2]/NET0131  ;
  input \P2_P2_InstQueue_reg[8][3]/NET0131  ;
  input \P2_P2_InstQueue_reg[8][4]/NET0131  ;
  input \P2_P2_InstQueue_reg[8][5]/NET0131  ;
  input \P2_P2_InstQueue_reg[8][6]/NET0131  ;
  input \P2_P2_InstQueue_reg[8][7]/NET0131  ;
  input \P2_P2_InstQueue_reg[9][0]/NET0131  ;
  input \P2_P2_InstQueue_reg[9][1]/NET0131  ;
  input \P2_P2_InstQueue_reg[9][2]/NET0131  ;
  input \P2_P2_InstQueue_reg[9][3]/NET0131  ;
  input \P2_P2_InstQueue_reg[9][4]/NET0131  ;
  input \P2_P2_InstQueue_reg[9][5]/NET0131  ;
  input \P2_P2_InstQueue_reg[9][6]/NET0131  ;
  input \P2_P2_InstQueue_reg[9][7]/NET0131  ;
  input \P2_P2_M_IO_n_reg/NET0131  ;
  input \P2_P2_MemoryFetch_reg/NET0131  ;
  input \P2_P2_More_reg/NET0131  ;
  input \P2_P2_PhyAddrPointer_reg[0]/NET0131  ;
  input \P2_P2_PhyAddrPointer_reg[10]/NET0131  ;
  input \P2_P2_PhyAddrPointer_reg[11]/NET0131  ;
  input \P2_P2_PhyAddrPointer_reg[12]/NET0131  ;
  input \P2_P2_PhyAddrPointer_reg[13]/NET0131  ;
  input \P2_P2_PhyAddrPointer_reg[14]/NET0131  ;
  input \P2_P2_PhyAddrPointer_reg[15]/NET0131  ;
  input \P2_P2_PhyAddrPointer_reg[16]/NET0131  ;
  input \P2_P2_PhyAddrPointer_reg[17]/NET0131  ;
  input \P2_P2_PhyAddrPointer_reg[18]/NET0131  ;
  input \P2_P2_PhyAddrPointer_reg[19]/NET0131  ;
  input \P2_P2_PhyAddrPointer_reg[1]/NET0131  ;
  input \P2_P2_PhyAddrPointer_reg[20]/NET0131  ;
  input \P2_P2_PhyAddrPointer_reg[21]/NET0131  ;
  input \P2_P2_PhyAddrPointer_reg[22]/NET0131  ;
  input \P2_P2_PhyAddrPointer_reg[23]/NET0131  ;
  input \P2_P2_PhyAddrPointer_reg[24]/NET0131  ;
  input \P2_P2_PhyAddrPointer_reg[25]/NET0131  ;
  input \P2_P2_PhyAddrPointer_reg[26]/NET0131  ;
  input \P2_P2_PhyAddrPointer_reg[27]/NET0131  ;
  input \P2_P2_PhyAddrPointer_reg[28]/NET0131  ;
  input \P2_P2_PhyAddrPointer_reg[29]/NET0131  ;
  input \P2_P2_PhyAddrPointer_reg[2]/NET0131  ;
  input \P2_P2_PhyAddrPointer_reg[30]/NET0131  ;
  input \P2_P2_PhyAddrPointer_reg[31]/NET0131  ;
  input \P2_P2_PhyAddrPointer_reg[3]/NET0131  ;
  input \P2_P2_PhyAddrPointer_reg[4]/NET0131  ;
  input \P2_P2_PhyAddrPointer_reg[5]/NET0131  ;
  input \P2_P2_PhyAddrPointer_reg[6]/NET0131  ;
  input \P2_P2_PhyAddrPointer_reg[7]/NET0131  ;
  input \P2_P2_PhyAddrPointer_reg[8]/NET0131  ;
  input \P2_P2_PhyAddrPointer_reg[9]/NET0131  ;
  input \P2_P2_ReadRequest_reg/NET0131  ;
  input \P2_P2_RequestPending_reg/NET0131  ;
  input \P2_P2_State2_reg[0]/NET0131  ;
  input \P2_P2_State2_reg[1]/NET0131  ;
  input \P2_P2_State2_reg[2]/NET0131  ;
  input \P2_P2_State2_reg[3]/NET0131  ;
  input \P2_P2_State_reg[0]/NET0131  ;
  input \P2_P2_State_reg[1]/NET0131  ;
  input \P2_P2_State_reg[2]/NET0131  ;
  input \P2_P2_W_R_n_reg/NET0131  ;
  input \P2_P2_lWord_reg[0]/NET0131  ;
  input \P2_P2_lWord_reg[10]/NET0131  ;
  input \P2_P2_lWord_reg[11]/NET0131  ;
  input \P2_P2_lWord_reg[12]/NET0131  ;
  input \P2_P2_lWord_reg[13]/NET0131  ;
  input \P2_P2_lWord_reg[14]/NET0131  ;
  input \P2_P2_lWord_reg[15]/NET0131  ;
  input \P2_P2_lWord_reg[1]/NET0131  ;
  input \P2_P2_lWord_reg[2]/NET0131  ;
  input \P2_P2_lWord_reg[3]/NET0131  ;
  input \P2_P2_lWord_reg[4]/NET0131  ;
  input \P2_P2_lWord_reg[5]/NET0131  ;
  input \P2_P2_lWord_reg[6]/NET0131  ;
  input \P2_P2_lWord_reg[7]/NET0131  ;
  input \P2_P2_lWord_reg[8]/NET0131  ;
  input \P2_P2_lWord_reg[9]/NET0131  ;
  input \P2_P2_rEIP_reg[0]/NET0131  ;
  input \P2_P2_rEIP_reg[10]/NET0131  ;
  input \P2_P2_rEIP_reg[11]/NET0131  ;
  input \P2_P2_rEIP_reg[12]/NET0131  ;
  input \P2_P2_rEIP_reg[13]/NET0131  ;
  input \P2_P2_rEIP_reg[14]/NET0131  ;
  input \P2_P2_rEIP_reg[15]/NET0131  ;
  input \P2_P2_rEIP_reg[16]/NET0131  ;
  input \P2_P2_rEIP_reg[17]/NET0131  ;
  input \P2_P2_rEIP_reg[18]/NET0131  ;
  input \P2_P2_rEIP_reg[19]/NET0131  ;
  input \P2_P2_rEIP_reg[1]/NET0131  ;
  input \P2_P2_rEIP_reg[20]/NET0131  ;
  input \P2_P2_rEIP_reg[21]/NET0131  ;
  input \P2_P2_rEIP_reg[22]/NET0131  ;
  input \P2_P2_rEIP_reg[23]/NET0131  ;
  input \P2_P2_rEIP_reg[24]/NET0131  ;
  input \P2_P2_rEIP_reg[25]/NET0131  ;
  input \P2_P2_rEIP_reg[26]/NET0131  ;
  input \P2_P2_rEIP_reg[27]/NET0131  ;
  input \P2_P2_rEIP_reg[28]/NET0131  ;
  input \P2_P2_rEIP_reg[29]/NET0131  ;
  input \P2_P2_rEIP_reg[2]/NET0131  ;
  input \P2_P2_rEIP_reg[30]/NET0131  ;
  input \P2_P2_rEIP_reg[31]/NET0131  ;
  input \P2_P2_rEIP_reg[3]/NET0131  ;
  input \P2_P2_rEIP_reg[4]/NET0131  ;
  input \P2_P2_rEIP_reg[5]/NET0131  ;
  input \P2_P2_rEIP_reg[6]/NET0131  ;
  input \P2_P2_rEIP_reg[7]/NET0131  ;
  input \P2_P2_rEIP_reg[8]/NET0131  ;
  input \P2_P2_rEIP_reg[9]/NET0131  ;
  input \P2_P2_uWord_reg[0]/NET0131  ;
  input \P2_P2_uWord_reg[10]/NET0131  ;
  input \P2_P2_uWord_reg[11]/NET0131  ;
  input \P2_P2_uWord_reg[12]/NET0131  ;
  input \P2_P2_uWord_reg[13]/NET0131  ;
  input \P2_P2_uWord_reg[14]/NET0131  ;
  input \P2_P2_uWord_reg[1]/NET0131  ;
  input \P2_P2_uWord_reg[2]/NET0131  ;
  input \P2_P2_uWord_reg[3]/NET0131  ;
  input \P2_P2_uWord_reg[4]/NET0131  ;
  input \P2_P2_uWord_reg[5]/NET0131  ;
  input \P2_P2_uWord_reg[6]/NET0131  ;
  input \P2_P2_uWord_reg[7]/NET0131  ;
  input \P2_P2_uWord_reg[8]/NET0131  ;
  input \P2_P2_uWord_reg[9]/NET0131  ;
  input \P2_P3_ADS_n_reg/NET0131  ;
  input \P2_P3_Address_reg[0]/NET0131  ;
  input \P2_P3_Address_reg[10]/NET0131  ;
  input \P2_P3_Address_reg[11]/NET0131  ;
  input \P2_P3_Address_reg[12]/NET0131  ;
  input \P2_P3_Address_reg[13]/NET0131  ;
  input \P2_P3_Address_reg[14]/NET0131  ;
  input \P2_P3_Address_reg[15]/NET0131  ;
  input \P2_P3_Address_reg[16]/NET0131  ;
  input \P2_P3_Address_reg[17]/NET0131  ;
  input \P2_P3_Address_reg[18]/NET0131  ;
  input \P2_P3_Address_reg[1]/NET0131  ;
  input \P2_P3_Address_reg[2]/NET0131  ;
  input \P2_P3_Address_reg[3]/NET0131  ;
  input \P2_P3_Address_reg[4]/NET0131  ;
  input \P2_P3_Address_reg[5]/NET0131  ;
  input \P2_P3_Address_reg[6]/NET0131  ;
  input \P2_P3_Address_reg[7]/NET0131  ;
  input \P2_P3_Address_reg[8]/NET0131  ;
  input \P2_P3_Address_reg[9]/NET0131  ;
  input \P2_P3_BE_n_reg[0]/NET0131  ;
  input \P2_P3_BE_n_reg[1]/NET0131  ;
  input \P2_P3_BE_n_reg[2]/NET0131  ;
  input \P2_P3_BE_n_reg[3]/NET0131  ;
  input \P2_P3_ByteEnable_reg[0]/NET0131  ;
  input \P2_P3_ByteEnable_reg[1]/NET0131  ;
  input \P2_P3_ByteEnable_reg[2]/NET0131  ;
  input \P2_P3_ByteEnable_reg[3]/NET0131  ;
  input \P2_P3_CodeFetch_reg/NET0131  ;
  input \P2_P3_D_C_n_reg/NET0131  ;
  input \P2_P3_DataWidth_reg[0]/NET0131  ;
  input \P2_P3_DataWidth_reg[1]/NET0131  ;
  input \P2_P3_Datao_reg[0]/NET0131  ;
  input \P2_P3_Datao_reg[10]/NET0131  ;
  input \P2_P3_Datao_reg[11]/NET0131  ;
  input \P2_P3_Datao_reg[12]/NET0131  ;
  input \P2_P3_Datao_reg[13]/NET0131  ;
  input \P2_P3_Datao_reg[14]/NET0131  ;
  input \P2_P3_Datao_reg[15]/NET0131  ;
  input \P2_P3_Datao_reg[16]/NET0131  ;
  input \P2_P3_Datao_reg[17]/NET0131  ;
  input \P2_P3_Datao_reg[18]/NET0131  ;
  input \P2_P3_Datao_reg[19]/NET0131  ;
  input \P2_P3_Datao_reg[1]/NET0131  ;
  input \P2_P3_Datao_reg[20]/NET0131  ;
  input \P2_P3_Datao_reg[21]/NET0131  ;
  input \P2_P3_Datao_reg[22]/NET0131  ;
  input \P2_P3_Datao_reg[23]/NET0131  ;
  input \P2_P3_Datao_reg[24]/NET0131  ;
  input \P2_P3_Datao_reg[25]/NET0131  ;
  input \P2_P3_Datao_reg[26]/NET0131  ;
  input \P2_P3_Datao_reg[27]/NET0131  ;
  input \P2_P3_Datao_reg[28]/NET0131  ;
  input \P2_P3_Datao_reg[29]/NET0131  ;
  input \P2_P3_Datao_reg[2]/NET0131  ;
  input \P2_P3_Datao_reg[30]/NET0131  ;
  input \P2_P3_Datao_reg[3]/NET0131  ;
  input \P2_P3_Datao_reg[4]/NET0131  ;
  input \P2_P3_Datao_reg[5]/NET0131  ;
  input \P2_P3_Datao_reg[6]/NET0131  ;
  input \P2_P3_Datao_reg[7]/NET0131  ;
  input \P2_P3_Datao_reg[8]/NET0131  ;
  input \P2_P3_Datao_reg[9]/NET0131  ;
  input \P2_P3_EAX_reg[0]/NET0131  ;
  input \P2_P3_EAX_reg[10]/NET0131  ;
  input \P2_P3_EAX_reg[11]/NET0131  ;
  input \P2_P3_EAX_reg[12]/NET0131  ;
  input \P2_P3_EAX_reg[13]/NET0131  ;
  input \P2_P3_EAX_reg[14]/NET0131  ;
  input \P2_P3_EAX_reg[15]/NET0131  ;
  input \P2_P3_EAX_reg[16]/NET0131  ;
  input \P2_P3_EAX_reg[17]/NET0131  ;
  input \P2_P3_EAX_reg[18]/NET0131  ;
  input \P2_P3_EAX_reg[19]/NET0131  ;
  input \P2_P3_EAX_reg[1]/NET0131  ;
  input \P2_P3_EAX_reg[20]/NET0131  ;
  input \P2_P3_EAX_reg[21]/NET0131  ;
  input \P2_P3_EAX_reg[22]/NET0131  ;
  input \P2_P3_EAX_reg[23]/NET0131  ;
  input \P2_P3_EAX_reg[24]/NET0131  ;
  input \P2_P3_EAX_reg[25]/NET0131  ;
  input \P2_P3_EAX_reg[26]/NET0131  ;
  input \P2_P3_EAX_reg[27]/NET0131  ;
  input \P2_P3_EAX_reg[28]/NET0131  ;
  input \P2_P3_EAX_reg[29]/NET0131  ;
  input \P2_P3_EAX_reg[2]/NET0131  ;
  input \P2_P3_EAX_reg[30]/NET0131  ;
  input \P2_P3_EAX_reg[31]/NET0131  ;
  input \P2_P3_EAX_reg[3]/NET0131  ;
  input \P2_P3_EAX_reg[4]/NET0131  ;
  input \P2_P3_EAX_reg[5]/NET0131  ;
  input \P2_P3_EAX_reg[6]/NET0131  ;
  input \P2_P3_EAX_reg[7]/NET0131  ;
  input \P2_P3_EAX_reg[8]/NET0131  ;
  input \P2_P3_EAX_reg[9]/NET0131  ;
  input \P2_P3_EBX_reg[0]/NET0131  ;
  input \P2_P3_EBX_reg[10]/NET0131  ;
  input \P2_P3_EBX_reg[11]/NET0131  ;
  input \P2_P3_EBX_reg[12]/NET0131  ;
  input \P2_P3_EBX_reg[13]/NET0131  ;
  input \P2_P3_EBX_reg[14]/NET0131  ;
  input \P2_P3_EBX_reg[15]/NET0131  ;
  input \P2_P3_EBX_reg[16]/NET0131  ;
  input \P2_P3_EBX_reg[17]/NET0131  ;
  input \P2_P3_EBX_reg[18]/NET0131  ;
  input \P2_P3_EBX_reg[19]/NET0131  ;
  input \P2_P3_EBX_reg[1]/NET0131  ;
  input \P2_P3_EBX_reg[20]/NET0131  ;
  input \P2_P3_EBX_reg[21]/NET0131  ;
  input \P2_P3_EBX_reg[22]/NET0131  ;
  input \P2_P3_EBX_reg[23]/NET0131  ;
  input \P2_P3_EBX_reg[24]/NET0131  ;
  input \P2_P3_EBX_reg[25]/NET0131  ;
  input \P2_P3_EBX_reg[26]/NET0131  ;
  input \P2_P3_EBX_reg[27]/NET0131  ;
  input \P2_P3_EBX_reg[28]/NET0131  ;
  input \P2_P3_EBX_reg[29]/NET0131  ;
  input \P2_P3_EBX_reg[2]/NET0131  ;
  input \P2_P3_EBX_reg[30]/NET0131  ;
  input \P2_P3_EBX_reg[31]/NET0131  ;
  input \P2_P3_EBX_reg[3]/NET0131  ;
  input \P2_P3_EBX_reg[4]/NET0131  ;
  input \P2_P3_EBX_reg[5]/NET0131  ;
  input \P2_P3_EBX_reg[6]/NET0131  ;
  input \P2_P3_EBX_reg[7]/NET0131  ;
  input \P2_P3_EBX_reg[8]/NET0131  ;
  input \P2_P3_EBX_reg[9]/NET0131  ;
  input \P2_P3_Flush_reg/NET0131  ;
  input \P2_P3_InstAddrPointer_reg[0]/NET0131  ;
  input \P2_P3_InstAddrPointer_reg[10]/NET0131  ;
  input \P2_P3_InstAddrPointer_reg[11]/NET0131  ;
  input \P2_P3_InstAddrPointer_reg[12]/NET0131  ;
  input \P2_P3_InstAddrPointer_reg[13]/NET0131  ;
  input \P2_P3_InstAddrPointer_reg[14]/NET0131  ;
  input \P2_P3_InstAddrPointer_reg[15]/NET0131  ;
  input \P2_P3_InstAddrPointer_reg[16]/NET0131  ;
  input \P2_P3_InstAddrPointer_reg[17]/NET0131  ;
  input \P2_P3_InstAddrPointer_reg[18]/NET0131  ;
  input \P2_P3_InstAddrPointer_reg[19]/NET0131  ;
  input \P2_P3_InstAddrPointer_reg[1]/NET0131  ;
  input \P2_P3_InstAddrPointer_reg[20]/NET0131  ;
  input \P2_P3_InstAddrPointer_reg[21]/NET0131  ;
  input \P2_P3_InstAddrPointer_reg[22]/NET0131  ;
  input \P2_P3_InstAddrPointer_reg[23]/NET0131  ;
  input \P2_P3_InstAddrPointer_reg[24]/NET0131  ;
  input \P2_P3_InstAddrPointer_reg[25]/NET0131  ;
  input \P2_P3_InstAddrPointer_reg[26]/NET0131  ;
  input \P2_P3_InstAddrPointer_reg[27]/NET0131  ;
  input \P2_P3_InstAddrPointer_reg[28]/NET0131  ;
  input \P2_P3_InstAddrPointer_reg[29]/NET0131  ;
  input \P2_P3_InstAddrPointer_reg[2]/NET0131  ;
  input \P2_P3_InstAddrPointer_reg[30]/NET0131  ;
  input \P2_P3_InstAddrPointer_reg[31]/NET0131  ;
  input \P2_P3_InstAddrPointer_reg[3]/NET0131  ;
  input \P2_P3_InstAddrPointer_reg[4]/NET0131  ;
  input \P2_P3_InstAddrPointer_reg[5]/NET0131  ;
  input \P2_P3_InstAddrPointer_reg[6]/NET0131  ;
  input \P2_P3_InstAddrPointer_reg[7]/NET0131  ;
  input \P2_P3_InstAddrPointer_reg[8]/NET0131  ;
  input \P2_P3_InstAddrPointer_reg[9]/NET0131  ;
  input \P2_P3_InstQueueRd_Addr_reg[0]/NET0131  ;
  input \P2_P3_InstQueueRd_Addr_reg[1]/NET0131  ;
  input \P2_P3_InstQueueRd_Addr_reg[2]/NET0131  ;
  input \P2_P3_InstQueueRd_Addr_reg[3]/NET0131  ;
  input \P2_P3_InstQueueWr_Addr_reg[0]/NET0131  ;
  input \P2_P3_InstQueueWr_Addr_reg[1]/NET0131  ;
  input \P2_P3_InstQueueWr_Addr_reg[2]/NET0131  ;
  input \P2_P3_InstQueueWr_Addr_reg[3]/NET0131  ;
  input \P2_P3_InstQueue_reg[0][0]/NET0131  ;
  input \P2_P3_InstQueue_reg[0][1]/NET0131  ;
  input \P2_P3_InstQueue_reg[0][2]/NET0131  ;
  input \P2_P3_InstQueue_reg[0][3]/NET0131  ;
  input \P2_P3_InstQueue_reg[0][4]/NET0131  ;
  input \P2_P3_InstQueue_reg[0][5]/NET0131  ;
  input \P2_P3_InstQueue_reg[0][6]/NET0131  ;
  input \P2_P3_InstQueue_reg[0][7]/NET0131  ;
  input \P2_P3_InstQueue_reg[10][0]/NET0131  ;
  input \P2_P3_InstQueue_reg[10][1]/NET0131  ;
  input \P2_P3_InstQueue_reg[10][2]/NET0131  ;
  input \P2_P3_InstQueue_reg[10][3]/NET0131  ;
  input \P2_P3_InstQueue_reg[10][4]/NET0131  ;
  input \P2_P3_InstQueue_reg[10][5]/NET0131  ;
  input \P2_P3_InstQueue_reg[10][6]/NET0131  ;
  input \P2_P3_InstQueue_reg[10][7]/NET0131  ;
  input \P2_P3_InstQueue_reg[11][0]/NET0131  ;
  input \P2_P3_InstQueue_reg[11][1]/NET0131  ;
  input \P2_P3_InstQueue_reg[11][2]/NET0131  ;
  input \P2_P3_InstQueue_reg[11][3]/NET0131  ;
  input \P2_P3_InstQueue_reg[11][4]/NET0131  ;
  input \P2_P3_InstQueue_reg[11][5]/NET0131  ;
  input \P2_P3_InstQueue_reg[11][6]/NET0131  ;
  input \P2_P3_InstQueue_reg[11][7]/NET0131  ;
  input \P2_P3_InstQueue_reg[12][0]/NET0131  ;
  input \P2_P3_InstQueue_reg[12][1]/NET0131  ;
  input \P2_P3_InstQueue_reg[12][2]/NET0131  ;
  input \P2_P3_InstQueue_reg[12][3]/NET0131  ;
  input \P2_P3_InstQueue_reg[12][4]/NET0131  ;
  input \P2_P3_InstQueue_reg[12][5]/NET0131  ;
  input \P2_P3_InstQueue_reg[12][6]/NET0131  ;
  input \P2_P3_InstQueue_reg[12][7]/NET0131  ;
  input \P2_P3_InstQueue_reg[13][0]/NET0131  ;
  input \P2_P3_InstQueue_reg[13][1]/NET0131  ;
  input \P2_P3_InstQueue_reg[13][2]/NET0131  ;
  input \P2_P3_InstQueue_reg[13][3]/NET0131  ;
  input \P2_P3_InstQueue_reg[13][4]/NET0131  ;
  input \P2_P3_InstQueue_reg[13][5]/NET0131  ;
  input \P2_P3_InstQueue_reg[13][6]/NET0131  ;
  input \P2_P3_InstQueue_reg[13][7]/NET0131  ;
  input \P2_P3_InstQueue_reg[14][0]/NET0131  ;
  input \P2_P3_InstQueue_reg[14][1]/NET0131  ;
  input \P2_P3_InstQueue_reg[14][2]/NET0131  ;
  input \P2_P3_InstQueue_reg[14][3]/NET0131  ;
  input \P2_P3_InstQueue_reg[14][4]/NET0131  ;
  input \P2_P3_InstQueue_reg[14][5]/NET0131  ;
  input \P2_P3_InstQueue_reg[14][6]/NET0131  ;
  input \P2_P3_InstQueue_reg[14][7]/NET0131  ;
  input \P2_P3_InstQueue_reg[15][0]/NET0131  ;
  input \P2_P3_InstQueue_reg[15][1]/NET0131  ;
  input \P2_P3_InstQueue_reg[15][2]/NET0131  ;
  input \P2_P3_InstQueue_reg[15][3]/NET0131  ;
  input \P2_P3_InstQueue_reg[15][4]/NET0131  ;
  input \P2_P3_InstQueue_reg[15][5]/NET0131  ;
  input \P2_P3_InstQueue_reg[15][6]/NET0131  ;
  input \P2_P3_InstQueue_reg[15][7]/NET0131  ;
  input \P2_P3_InstQueue_reg[1][0]/NET0131  ;
  input \P2_P3_InstQueue_reg[1][1]/NET0131  ;
  input \P2_P3_InstQueue_reg[1][2]/NET0131  ;
  input \P2_P3_InstQueue_reg[1][3]/NET0131  ;
  input \P2_P3_InstQueue_reg[1][4]/NET0131  ;
  input \P2_P3_InstQueue_reg[1][5]/NET0131  ;
  input \P2_P3_InstQueue_reg[1][6]/NET0131  ;
  input \P2_P3_InstQueue_reg[1][7]/NET0131  ;
  input \P2_P3_InstQueue_reg[2][0]/NET0131  ;
  input \P2_P3_InstQueue_reg[2][1]/NET0131  ;
  input \P2_P3_InstQueue_reg[2][2]/NET0131  ;
  input \P2_P3_InstQueue_reg[2][3]/NET0131  ;
  input \P2_P3_InstQueue_reg[2][4]/NET0131  ;
  input \P2_P3_InstQueue_reg[2][5]/NET0131  ;
  input \P2_P3_InstQueue_reg[2][6]/NET0131  ;
  input \P2_P3_InstQueue_reg[2][7]/NET0131  ;
  input \P2_P3_InstQueue_reg[3][0]/NET0131  ;
  input \P2_P3_InstQueue_reg[3][1]/NET0131  ;
  input \P2_P3_InstQueue_reg[3][2]/NET0131  ;
  input \P2_P3_InstQueue_reg[3][3]/NET0131  ;
  input \P2_P3_InstQueue_reg[3][4]/NET0131  ;
  input \P2_P3_InstQueue_reg[3][5]/NET0131  ;
  input \P2_P3_InstQueue_reg[3][6]/NET0131  ;
  input \P2_P3_InstQueue_reg[3][7]/NET0131  ;
  input \P2_P3_InstQueue_reg[4][0]/NET0131  ;
  input \P2_P3_InstQueue_reg[4][1]/NET0131  ;
  input \P2_P3_InstQueue_reg[4][2]/NET0131  ;
  input \P2_P3_InstQueue_reg[4][3]/NET0131  ;
  input \P2_P3_InstQueue_reg[4][4]/NET0131  ;
  input \P2_P3_InstQueue_reg[4][5]/NET0131  ;
  input \P2_P3_InstQueue_reg[4][6]/NET0131  ;
  input \P2_P3_InstQueue_reg[4][7]/NET0131  ;
  input \P2_P3_InstQueue_reg[5][0]/NET0131  ;
  input \P2_P3_InstQueue_reg[5][1]/NET0131  ;
  input \P2_P3_InstQueue_reg[5][2]/NET0131  ;
  input \P2_P3_InstQueue_reg[5][3]/NET0131  ;
  input \P2_P3_InstQueue_reg[5][4]/NET0131  ;
  input \P2_P3_InstQueue_reg[5][5]/NET0131  ;
  input \P2_P3_InstQueue_reg[5][6]/NET0131  ;
  input \P2_P3_InstQueue_reg[5][7]/NET0131  ;
  input \P2_P3_InstQueue_reg[6][0]/NET0131  ;
  input \P2_P3_InstQueue_reg[6][1]/NET0131  ;
  input \P2_P3_InstQueue_reg[6][2]/NET0131  ;
  input \P2_P3_InstQueue_reg[6][3]/NET0131  ;
  input \P2_P3_InstQueue_reg[6][4]/NET0131  ;
  input \P2_P3_InstQueue_reg[6][5]/NET0131  ;
  input \P2_P3_InstQueue_reg[6][6]/NET0131  ;
  input \P2_P3_InstQueue_reg[6][7]/NET0131  ;
  input \P2_P3_InstQueue_reg[7][0]/NET0131  ;
  input \P2_P3_InstQueue_reg[7][1]/NET0131  ;
  input \P2_P3_InstQueue_reg[7][2]/NET0131  ;
  input \P2_P3_InstQueue_reg[7][3]/NET0131  ;
  input \P2_P3_InstQueue_reg[7][4]/NET0131  ;
  input \P2_P3_InstQueue_reg[7][5]/NET0131  ;
  input \P2_P3_InstQueue_reg[7][6]/NET0131  ;
  input \P2_P3_InstQueue_reg[7][7]/NET0131  ;
  input \P2_P3_InstQueue_reg[8][0]/NET0131  ;
  input \P2_P3_InstQueue_reg[8][1]/NET0131  ;
  input \P2_P3_InstQueue_reg[8][2]/NET0131  ;
  input \P2_P3_InstQueue_reg[8][3]/NET0131  ;
  input \P2_P3_InstQueue_reg[8][4]/NET0131  ;
  input \P2_P3_InstQueue_reg[8][5]/NET0131  ;
  input \P2_P3_InstQueue_reg[8][6]/NET0131  ;
  input \P2_P3_InstQueue_reg[8][7]/NET0131  ;
  input \P2_P3_InstQueue_reg[9][0]/NET0131  ;
  input \P2_P3_InstQueue_reg[9][1]/NET0131  ;
  input \P2_P3_InstQueue_reg[9][2]/NET0131  ;
  input \P2_P3_InstQueue_reg[9][3]/NET0131  ;
  input \P2_P3_InstQueue_reg[9][4]/NET0131  ;
  input \P2_P3_InstQueue_reg[9][5]/NET0131  ;
  input \P2_P3_InstQueue_reg[9][6]/NET0131  ;
  input \P2_P3_InstQueue_reg[9][7]/NET0131  ;
  input \P2_P3_M_IO_n_reg/NET0131  ;
  input \P2_P3_MemoryFetch_reg/NET0131  ;
  input \P2_P3_More_reg/NET0131  ;
  input \P2_P3_PhyAddrPointer_reg[0]/NET0131  ;
  input \P2_P3_PhyAddrPointer_reg[10]/NET0131  ;
  input \P2_P3_PhyAddrPointer_reg[11]/NET0131  ;
  input \P2_P3_PhyAddrPointer_reg[12]/NET0131  ;
  input \P2_P3_PhyAddrPointer_reg[13]/NET0131  ;
  input \P2_P3_PhyAddrPointer_reg[14]/NET0131  ;
  input \P2_P3_PhyAddrPointer_reg[15]/NET0131  ;
  input \P2_P3_PhyAddrPointer_reg[16]/NET0131  ;
  input \P2_P3_PhyAddrPointer_reg[17]/NET0131  ;
  input \P2_P3_PhyAddrPointer_reg[18]/NET0131  ;
  input \P2_P3_PhyAddrPointer_reg[19]/NET0131  ;
  input \P2_P3_PhyAddrPointer_reg[1]/NET0131  ;
  input \P2_P3_PhyAddrPointer_reg[20]/NET0131  ;
  input \P2_P3_PhyAddrPointer_reg[21]/NET0131  ;
  input \P2_P3_PhyAddrPointer_reg[22]/NET0131  ;
  input \P2_P3_PhyAddrPointer_reg[23]/NET0131  ;
  input \P2_P3_PhyAddrPointer_reg[24]/NET0131  ;
  input \P2_P3_PhyAddrPointer_reg[25]/NET0131  ;
  input \P2_P3_PhyAddrPointer_reg[26]/NET0131  ;
  input \P2_P3_PhyAddrPointer_reg[27]/NET0131  ;
  input \P2_P3_PhyAddrPointer_reg[28]/NET0131  ;
  input \P2_P3_PhyAddrPointer_reg[29]/NET0131  ;
  input \P2_P3_PhyAddrPointer_reg[2]/NET0131  ;
  input \P2_P3_PhyAddrPointer_reg[30]/NET0131  ;
  input \P2_P3_PhyAddrPointer_reg[31]/NET0131  ;
  input \P2_P3_PhyAddrPointer_reg[3]/NET0131  ;
  input \P2_P3_PhyAddrPointer_reg[4]/NET0131  ;
  input \P2_P3_PhyAddrPointer_reg[5]/NET0131  ;
  input \P2_P3_PhyAddrPointer_reg[6]/NET0131  ;
  input \P2_P3_PhyAddrPointer_reg[7]/NET0131  ;
  input \P2_P3_PhyAddrPointer_reg[8]/NET0131  ;
  input \P2_P3_PhyAddrPointer_reg[9]/NET0131  ;
  input \P2_P3_ReadRequest_reg/NET0131  ;
  input \P2_P3_RequestPending_reg/NET0131  ;
  input \P2_P3_State2_reg[0]/NET0131  ;
  input \P2_P3_State2_reg[1]/NET0131  ;
  input \P2_P3_State2_reg[2]/NET0131  ;
  input \P2_P3_State2_reg[3]/NET0131  ;
  input \P2_P3_State_reg[0]/NET0131  ;
  input \P2_P3_State_reg[1]/NET0131  ;
  input \P2_P3_State_reg[2]/NET0131  ;
  input \P2_P3_W_R_n_reg/NET0131  ;
  input \P2_P3_lWord_reg[0]/NET0131  ;
  input \P2_P3_lWord_reg[10]/NET0131  ;
  input \P2_P3_lWord_reg[11]/NET0131  ;
  input \P2_P3_lWord_reg[12]/NET0131  ;
  input \P2_P3_lWord_reg[13]/NET0131  ;
  input \P2_P3_lWord_reg[14]/NET0131  ;
  input \P2_P3_lWord_reg[15]/NET0131  ;
  input \P2_P3_lWord_reg[1]/NET0131  ;
  input \P2_P3_lWord_reg[2]/NET0131  ;
  input \P2_P3_lWord_reg[3]/NET0131  ;
  input \P2_P3_lWord_reg[4]/NET0131  ;
  input \P2_P3_lWord_reg[5]/NET0131  ;
  input \P2_P3_lWord_reg[6]/NET0131  ;
  input \P2_P3_lWord_reg[7]/NET0131  ;
  input \P2_P3_lWord_reg[8]/NET0131  ;
  input \P2_P3_lWord_reg[9]/NET0131  ;
  input \P2_P3_rEIP_reg[0]/NET0131  ;
  input \P2_P3_rEIP_reg[10]/NET0131  ;
  input \P2_P3_rEIP_reg[11]/NET0131  ;
  input \P2_P3_rEIP_reg[12]/NET0131  ;
  input \P2_P3_rEIP_reg[13]/NET0131  ;
  input \P2_P3_rEIP_reg[14]/NET0131  ;
  input \P2_P3_rEIP_reg[15]/NET0131  ;
  input \P2_P3_rEIP_reg[16]/NET0131  ;
  input \P2_P3_rEIP_reg[17]/NET0131  ;
  input \P2_P3_rEIP_reg[18]/NET0131  ;
  input \P2_P3_rEIP_reg[19]/NET0131  ;
  input \P2_P3_rEIP_reg[1]/NET0131  ;
  input \P2_P3_rEIP_reg[20]/NET0131  ;
  input \P2_P3_rEIP_reg[21]/NET0131  ;
  input \P2_P3_rEIP_reg[22]/NET0131  ;
  input \P2_P3_rEIP_reg[23]/NET0131  ;
  input \P2_P3_rEIP_reg[24]/NET0131  ;
  input \P2_P3_rEIP_reg[25]/NET0131  ;
  input \P2_P3_rEIP_reg[26]/NET0131  ;
  input \P2_P3_rEIP_reg[27]/NET0131  ;
  input \P2_P3_rEIP_reg[28]/NET0131  ;
  input \P2_P3_rEIP_reg[29]/NET0131  ;
  input \P2_P3_rEIP_reg[2]/NET0131  ;
  input \P2_P3_rEIP_reg[30]/NET0131  ;
  input \P2_P3_rEIP_reg[31]/NET0131  ;
  input \P2_P3_rEIP_reg[3]/NET0131  ;
  input \P2_P3_rEIP_reg[4]/NET0131  ;
  input \P2_P3_rEIP_reg[5]/NET0131  ;
  input \P2_P3_rEIP_reg[6]/NET0131  ;
  input \P2_P3_rEIP_reg[7]/NET0131  ;
  input \P2_P3_rEIP_reg[8]/NET0131  ;
  input \P2_P3_rEIP_reg[9]/NET0131  ;
  input \P2_P3_uWord_reg[0]/NET0131  ;
  input \P2_P3_uWord_reg[10]/NET0131  ;
  input \P2_P3_uWord_reg[11]/NET0131  ;
  input \P2_P3_uWord_reg[12]/NET0131  ;
  input \P2_P3_uWord_reg[13]/NET0131  ;
  input \P2_P3_uWord_reg[14]/NET0131  ;
  input \P2_P3_uWord_reg[1]/NET0131  ;
  input \P2_P3_uWord_reg[2]/NET0131  ;
  input \P2_P3_uWord_reg[3]/NET0131  ;
  input \P2_P3_uWord_reg[4]/NET0131  ;
  input \P2_P3_uWord_reg[5]/NET0131  ;
  input \P2_P3_uWord_reg[6]/NET0131  ;
  input \P2_P3_uWord_reg[7]/NET0131  ;
  input \P2_P3_uWord_reg[8]/NET0131  ;
  input \P2_P3_uWord_reg[9]/NET0131  ;
  input \P2_buf1_reg[0]/NET0131  ;
  input \P2_buf1_reg[10]/NET0131  ;
  input \P2_buf1_reg[11]/NET0131  ;
  input \P2_buf1_reg[12]/NET0131  ;
  input \P2_buf1_reg[13]/NET0131  ;
  input \P2_buf1_reg[14]/NET0131  ;
  input \P2_buf1_reg[15]/NET0131  ;
  input \P2_buf1_reg[16]/NET0131  ;
  input \P2_buf1_reg[17]/NET0131  ;
  input \P2_buf1_reg[18]/NET0131  ;
  input \P2_buf1_reg[19]/NET0131  ;
  input \P2_buf1_reg[1]/NET0131  ;
  input \P2_buf1_reg[20]/NET0131  ;
  input \P2_buf1_reg[21]/NET0131  ;
  input \P2_buf1_reg[22]/NET0131  ;
  input \P2_buf1_reg[23]/NET0131  ;
  input \P2_buf1_reg[24]/NET0131  ;
  input \P2_buf1_reg[25]/NET0131  ;
  input \P2_buf1_reg[26]/NET0131  ;
  input \P2_buf1_reg[27]/NET0131  ;
  input \P2_buf1_reg[28]/NET0131  ;
  input \P2_buf1_reg[29]/NET0131  ;
  input \P2_buf1_reg[2]/NET0131  ;
  input \P2_buf1_reg[30]/NET0131  ;
  input \P2_buf1_reg[3]/NET0131  ;
  input \P2_buf1_reg[4]/NET0131  ;
  input \P2_buf1_reg[5]/NET0131  ;
  input \P2_buf1_reg[6]/NET0131  ;
  input \P2_buf1_reg[7]/NET0131  ;
  input \P2_buf1_reg[8]/NET0131  ;
  input \P2_buf1_reg[9]/NET0131  ;
  input \P2_buf2_reg[0]/NET0131  ;
  input \P2_buf2_reg[10]/NET0131  ;
  input \P2_buf2_reg[11]/NET0131  ;
  input \P2_buf2_reg[12]/NET0131  ;
  input \P2_buf2_reg[13]/NET0131  ;
  input \P2_buf2_reg[14]/NET0131  ;
  input \P2_buf2_reg[15]/NET0131  ;
  input \P2_buf2_reg[16]/NET0131  ;
  input \P2_buf2_reg[17]/NET0131  ;
  input \P2_buf2_reg[18]/NET0131  ;
  input \P2_buf2_reg[19]/NET0131  ;
  input \P2_buf2_reg[1]/NET0131  ;
  input \P2_buf2_reg[20]/NET0131  ;
  input \P2_buf2_reg[21]/NET0131  ;
  input \P2_buf2_reg[22]/NET0131  ;
  input \P2_buf2_reg[23]/NET0131  ;
  input \P2_buf2_reg[24]/NET0131  ;
  input \P2_buf2_reg[25]/NET0131  ;
  input \P2_buf2_reg[26]/NET0131  ;
  input \P2_buf2_reg[27]/NET0131  ;
  input \P2_buf2_reg[28]/NET0131  ;
  input \P2_buf2_reg[29]/NET0131  ;
  input \P2_buf2_reg[2]/NET0131  ;
  input \P2_buf2_reg[30]/NET0131  ;
  input \P2_buf2_reg[3]/NET0131  ;
  input \P2_buf2_reg[4]/NET0131  ;
  input \P2_buf2_reg[5]/NET0131  ;
  input \P2_buf2_reg[6]/NET0131  ;
  input \P2_buf2_reg[7]/NET0131  ;
  input \P2_buf2_reg[8]/NET0131  ;
  input \P2_buf2_reg[9]/NET0131  ;
  input \P2_ready11_reg/NET0131  ;
  input \P2_ready12_reg/NET0131  ;
  input \P2_ready21_reg/NET0131  ;
  input \P2_ready22_reg/NET0131  ;
  input \P3_rd_reg/NET0131  ;
  input \P4_B_reg/NET0131  ;
  input \P4_IR_reg[0]/NET0131  ;
  input \P4_IR_reg[10]/NET0131  ;
  input \P4_IR_reg[11]/NET0131  ;
  input \P4_IR_reg[12]/NET0131  ;
  input \P4_IR_reg[13]/NET0131  ;
  input \P4_IR_reg[14]/NET0131  ;
  input \P4_IR_reg[15]/NET0131  ;
  input \P4_IR_reg[16]/NET0131  ;
  input \P4_IR_reg[17]/NET0131  ;
  input \P4_IR_reg[18]/NET0131  ;
  input \P4_IR_reg[19]/NET0131  ;
  input \P4_IR_reg[1]/NET0131  ;
  input \P4_IR_reg[20]/NET0131  ;
  input \P4_IR_reg[21]/NET0131  ;
  input \P4_IR_reg[22]/NET0131  ;
  input \P4_IR_reg[23]/NET0131  ;
  input \P4_IR_reg[24]/NET0131  ;
  input \P4_IR_reg[25]/NET0131  ;
  input \P4_IR_reg[26]/NET0131  ;
  input \P4_IR_reg[27]/NET0131  ;
  input \P4_IR_reg[28]/NET0131  ;
  input \P4_IR_reg[29]/NET0131  ;
  input \P4_IR_reg[2]/NET0131  ;
  input \P4_IR_reg[30]/NET0131  ;
  input \P4_IR_reg[3]/NET0131  ;
  input \P4_IR_reg[4]/NET0131  ;
  input \P4_IR_reg[5]/NET0131  ;
  input \P4_IR_reg[6]/NET0131  ;
  input \P4_IR_reg[7]/NET0131  ;
  input \P4_IR_reg[8]/NET0131  ;
  input \P4_IR_reg[9]/NET0131  ;
  input \P4_addr_reg[0]/NET0131  ;
  input \P4_addr_reg[10]/NET0131  ;
  input \P4_addr_reg[11]/NET0131  ;
  input \P4_addr_reg[12]/NET0131  ;
  input \P4_addr_reg[13]/NET0131  ;
  input \P4_addr_reg[14]/NET0131  ;
  input \P4_addr_reg[15]/NET0131  ;
  input \P4_addr_reg[16]/NET0131  ;
  input \P4_addr_reg[17]/NET0131  ;
  input \P4_addr_reg[18]/NET0131  ;
  input \P4_addr_reg[1]/NET0131  ;
  input \P4_addr_reg[2]/NET0131  ;
  input \P4_addr_reg[3]/NET0131  ;
  input \P4_addr_reg[4]/NET0131  ;
  input \P4_addr_reg[5]/NET0131  ;
  input \P4_addr_reg[6]/NET0131  ;
  input \P4_addr_reg[7]/NET0131  ;
  input \P4_addr_reg[8]/NET0131  ;
  input \P4_addr_reg[9]/NET0131  ;
  input \P4_d_reg[0]/NET0131  ;
  input \P4_d_reg[1]/NET0131  ;
  input \P4_datao_reg[0]/NET0131  ;
  input \P4_datao_reg[10]/NET0131  ;
  input \P4_datao_reg[11]/NET0131  ;
  input \P4_datao_reg[12]/NET0131  ;
  input \P4_datao_reg[13]/NET0131  ;
  input \P4_datao_reg[14]/NET0131  ;
  input \P4_datao_reg[15]/NET0131  ;
  input \P4_datao_reg[16]/NET0131  ;
  input \P4_datao_reg[17]/NET0131  ;
  input \P4_datao_reg[18]/NET0131  ;
  input \P4_datao_reg[19]/NET0131  ;
  input \P4_datao_reg[1]/NET0131  ;
  input \P4_datao_reg[20]/NET0131  ;
  input \P4_datao_reg[21]/NET0131  ;
  input \P4_datao_reg[22]/NET0131  ;
  input \P4_datao_reg[23]/NET0131  ;
  input \P4_datao_reg[24]/NET0131  ;
  input \P4_datao_reg[25]/NET0131  ;
  input \P4_datao_reg[26]/NET0131  ;
  input \P4_datao_reg[27]/NET0131  ;
  input \P4_datao_reg[28]/NET0131  ;
  input \P4_datao_reg[29]/NET0131  ;
  input \P4_datao_reg[2]/NET0131  ;
  input \P4_datao_reg[30]/NET0131  ;
  input \P4_datao_reg[31]/NET0131  ;
  input \P4_datao_reg[3]/NET0131  ;
  input \P4_datao_reg[4]/NET0131  ;
  input \P4_datao_reg[5]/NET0131  ;
  input \P4_datao_reg[6]/NET0131  ;
  input \P4_datao_reg[7]/NET0131  ;
  input \P4_datao_reg[8]/NET0131  ;
  input \P4_datao_reg[9]/NET0131  ;
  input \P4_rd_reg/NET0131  ;
  input \P4_reg0_reg[0]/NET0131  ;
  input \P4_reg0_reg[10]/NET0131  ;
  input \P4_reg0_reg[11]/NET0131  ;
  input \P4_reg0_reg[12]/NET0131  ;
  input \P4_reg0_reg[13]/NET0131  ;
  input \P4_reg0_reg[14]/NET0131  ;
  input \P4_reg0_reg[15]/NET0131  ;
  input \P4_reg0_reg[16]/NET0131  ;
  input \P4_reg0_reg[17]/NET0131  ;
  input \P4_reg0_reg[18]/NET0131  ;
  input \P4_reg0_reg[19]/NET0131  ;
  input \P4_reg0_reg[1]/NET0131  ;
  input \P4_reg0_reg[20]/NET0131  ;
  input \P4_reg0_reg[21]/NET0131  ;
  input \P4_reg0_reg[22]/NET0131  ;
  input \P4_reg0_reg[23]/NET0131  ;
  input \P4_reg0_reg[24]/NET0131  ;
  input \P4_reg0_reg[25]/NET0131  ;
  input \P4_reg0_reg[26]/NET0131  ;
  input \P4_reg0_reg[27]/NET0131  ;
  input \P4_reg0_reg[28]/NET0131  ;
  input \P4_reg0_reg[29]/NET0131  ;
  input \P4_reg0_reg[2]/NET0131  ;
  input \P4_reg0_reg[30]/NET0131  ;
  input \P4_reg0_reg[31]/NET0131  ;
  input \P4_reg0_reg[3]/NET0131  ;
  input \P4_reg0_reg[4]/NET0131  ;
  input \P4_reg0_reg[5]/NET0131  ;
  input \P4_reg0_reg[6]/NET0131  ;
  input \P4_reg0_reg[7]/NET0131  ;
  input \P4_reg0_reg[8]/NET0131  ;
  input \P4_reg0_reg[9]/NET0131  ;
  input \P4_reg1_reg[0]/NET0131  ;
  input \P4_reg1_reg[10]/NET0131  ;
  input \P4_reg1_reg[11]/NET0131  ;
  input \P4_reg1_reg[12]/NET0131  ;
  input \P4_reg1_reg[13]/NET0131  ;
  input \P4_reg1_reg[14]/NET0131  ;
  input \P4_reg1_reg[15]/NET0131  ;
  input \P4_reg1_reg[16]/NET0131  ;
  input \P4_reg1_reg[17]/NET0131  ;
  input \P4_reg1_reg[18]/NET0131  ;
  input \P4_reg1_reg[19]/NET0131  ;
  input \P4_reg1_reg[1]/NET0131  ;
  input \P4_reg1_reg[20]/NET0131  ;
  input \P4_reg1_reg[21]/NET0131  ;
  input \P4_reg1_reg[22]/NET0131  ;
  input \P4_reg1_reg[23]/NET0131  ;
  input \P4_reg1_reg[24]/NET0131  ;
  input \P4_reg1_reg[25]/NET0131  ;
  input \P4_reg1_reg[26]/NET0131  ;
  input \P4_reg1_reg[27]/NET0131  ;
  input \P4_reg1_reg[28]/NET0131  ;
  input \P4_reg1_reg[29]/NET0131  ;
  input \P4_reg1_reg[2]/NET0131  ;
  input \P4_reg1_reg[30]/NET0131  ;
  input \P4_reg1_reg[31]/NET0131  ;
  input \P4_reg1_reg[3]/NET0131  ;
  input \P4_reg1_reg[4]/NET0131  ;
  input \P4_reg1_reg[5]/NET0131  ;
  input \P4_reg1_reg[6]/NET0131  ;
  input \P4_reg1_reg[7]/NET0131  ;
  input \P4_reg1_reg[8]/NET0131  ;
  input \P4_reg1_reg[9]/NET0131  ;
  input \P4_reg2_reg[0]/NET0131  ;
  input \P4_reg2_reg[10]/NET0131  ;
  input \P4_reg2_reg[11]/NET0131  ;
  input \P4_reg2_reg[12]/NET0131  ;
  input \P4_reg2_reg[13]/NET0131  ;
  input \P4_reg2_reg[14]/NET0131  ;
  input \P4_reg2_reg[15]/NET0131  ;
  input \P4_reg2_reg[16]/NET0131  ;
  input \P4_reg2_reg[17]/NET0131  ;
  input \P4_reg2_reg[18]/NET0131  ;
  input \P4_reg2_reg[19]/NET0131  ;
  input \P4_reg2_reg[1]/NET0131  ;
  input \P4_reg2_reg[20]/NET0131  ;
  input \P4_reg2_reg[21]/NET0131  ;
  input \P4_reg2_reg[22]/NET0131  ;
  input \P4_reg2_reg[23]/NET0131  ;
  input \P4_reg2_reg[24]/NET0131  ;
  input \P4_reg2_reg[25]/NET0131  ;
  input \P4_reg2_reg[26]/NET0131  ;
  input \P4_reg2_reg[27]/NET0131  ;
  input \P4_reg2_reg[28]/NET0131  ;
  input \P4_reg2_reg[29]/NET0131  ;
  input \P4_reg2_reg[2]/NET0131  ;
  input \P4_reg2_reg[30]/NET0131  ;
  input \P4_reg2_reg[31]/NET0131  ;
  input \P4_reg2_reg[3]/NET0131  ;
  input \P4_reg2_reg[4]/NET0131  ;
  input \P4_reg2_reg[5]/NET0131  ;
  input \P4_reg2_reg[6]/NET0131  ;
  input \P4_reg2_reg[7]/NET0131  ;
  input \P4_reg2_reg[8]/NET0131  ;
  input \P4_reg2_reg[9]/NET0131  ;
  input \P4_reg3_reg[0]/NET0131  ;
  input \P4_reg3_reg[10]/NET0131  ;
  input \P4_reg3_reg[11]/NET0131  ;
  input \P4_reg3_reg[12]/NET0131  ;
  input \P4_reg3_reg[13]/NET0131  ;
  input \P4_reg3_reg[14]/NET0131  ;
  input \P4_reg3_reg[15]/NET0131  ;
  input \P4_reg3_reg[16]/NET0131  ;
  input \P4_reg3_reg[17]/NET0131  ;
  input \P4_reg3_reg[18]/NET0131  ;
  input \P4_reg3_reg[19]/NET0131  ;
  input \P4_reg3_reg[1]/NET0131  ;
  input \P4_reg3_reg[20]/NET0131  ;
  input \P4_reg3_reg[21]/NET0131  ;
  input \P4_reg3_reg[22]/NET0131  ;
  input \P4_reg3_reg[23]/NET0131  ;
  input \P4_reg3_reg[24]/NET0131  ;
  input \P4_reg3_reg[25]/NET0131  ;
  input \P4_reg3_reg[26]/NET0131  ;
  input \P4_reg3_reg[27]/NET0131  ;
  input \P4_reg3_reg[28]/NET0131  ;
  input \P4_reg3_reg[2]/NET0131  ;
  input \P4_reg3_reg[3]/NET0131  ;
  input \P4_reg3_reg[4]/NET0131  ;
  input \P4_reg3_reg[5]/NET0131  ;
  input \P4_reg3_reg[6]/NET0131  ;
  input \P4_reg3_reg[7]/NET0131  ;
  input \P4_reg3_reg[8]/NET0131  ;
  input \P4_reg3_reg[9]/NET0131  ;
  input \P4_wr_reg/NET0131  ;
  input bs_pad ;
  input \din[0]_pad  ;
  input \din[10]_pad  ;
  input \din[11]_pad  ;
  input \din[12]_pad  ;
  input \din[13]_pad  ;
  input \din[14]_pad  ;
  input \din[15]_pad  ;
  input \din[16]_pad  ;
  input \din[17]_pad  ;
  input \din[18]_pad  ;
  input \din[19]_pad  ;
  input \din[1]_pad  ;
  input \din[20]_pad  ;
  input \din[21]_pad  ;
  input \din[22]_pad  ;
  input \din[23]_pad  ;
  input \din[24]_pad  ;
  input \din[25]_pad  ;
  input \din[26]_pad  ;
  input \din[27]_pad  ;
  input \din[28]_pad  ;
  input \din[29]_pad  ;
  input \din[2]_pad  ;
  input \din[30]_pad  ;
  input \din[31]_pad  ;
  input \din[3]_pad  ;
  input \din[4]_pad  ;
  input \din[5]_pad  ;
  input \din[6]_pad  ;
  input \din[7]_pad  ;
  input \din[8]_pad  ;
  input \din[9]_pad  ;
  input hold_pad ;
  input na_pad ;
  input sel_pad ;
  output \P3_state_reg[0]/NET0131_syn_2  ;
  output \_al_n1  ;
  output \aux[0]_pad  ;
  output \aux[1]_pad  ;
  output \aux[2]_pad  ;
  output \dout[0]_pad  ;
  output \dout[10]_pad  ;
  output \dout[11]_pad  ;
  output \dout[12]_pad  ;
  output \dout[13]_pad  ;
  output \dout[14]_pad  ;
  output \dout[15]_pad  ;
  output \dout[16]_pad  ;
  output \dout[17]_pad  ;
  output \dout[18]_pad  ;
  output \dout[19]_pad  ;
  output \dout[1]_pad  ;
  output \dout[2]_pad  ;
  output \dout[3]_pad  ;
  output \dout[4]_pad  ;
  output \dout[5]_pad  ;
  output \dout[6]_pad  ;
  output \dout[7]_pad  ;
  output \dout[8]_pad  ;
  output \dout[9]_pad  ;
  output \g326201/_0_  ;
  output \g326202/_0_  ;
  output \g326203/_0_  ;
  output \g326204/_0_  ;
  output \g326205/_0_  ;
  output \g326206/_0_  ;
  output \g326207/_0_  ;
  output \g326208/_0_  ;
  output \g326209/_0_  ;
  output \g326210/_0_  ;
  output \g326211/_0_  ;
  output \g326212/_0_  ;
  output \g326213/_0_  ;
  output \g326214/_0_  ;
  output \g326215/_0_  ;
  output \g326216/_0_  ;
  output \g326251/_0_  ;
  output \g326255/_0_  ;
  output \g326256/_0_  ;
  output \g326271/_0_  ;
  output \g326272/_0_  ;
  output \g326273/_0_  ;
  output \g326274/_0_  ;
  output \g326275/_0_  ;
  output \g326276/_0_  ;
  output \g326277/_0_  ;
  output \g326278/_0_  ;
  output \g326279/_0_  ;
  output \g326280/_0_  ;
  output \g326281/_0_  ;
  output \g326282/_0_  ;
  output \g326283/_0_  ;
  output \g326284/_0_  ;
  output \g326285/_0_  ;
  output \g326286/_0_  ;
  output \g326287/_0_  ;
  output \g326288/_0_  ;
  output \g326289/_0_  ;
  output \g326290/_0_  ;
  output \g326291/_0_  ;
  output \g326292/_0_  ;
  output \g326293/_0_  ;
  output \g326294/_0_  ;
  output \g326295/_0_  ;
  output \g326296/_0_  ;
  output \g326297/_0_  ;
  output \g326298/_0_  ;
  output \g326299/_0_  ;
  output \g326300/_0_  ;
  output \g326301/_0_  ;
  output \g326335/_0_  ;
  output \g326369/_0_  ;
  output \g326370/_0_  ;
  output \g326371/_0_  ;
  output \g326372/_0_  ;
  output \g326373/_0_  ;
  output \g326374/_0_  ;
  output \g326375/_0_  ;
  output \g326376/_0_  ;
  output \g326377/_0_  ;
  output \g326378/_0_  ;
  output \g326379/_0_  ;
  output \g326380/_0_  ;
  output \g326381/_0_  ;
  output \g326382/_0_  ;
  output \g326383/_0_  ;
  output \g326384/_0_  ;
  output \g326385/_0_  ;
  output \g326386/_0_  ;
  output \g326387/_0_  ;
  output \g326388/_0_  ;
  output \g326389/_0_  ;
  output \g326390/_0_  ;
  output \g326391/_0_  ;
  output \g326392/_0_  ;
  output \g326393/_0_  ;
  output \g326394/_0_  ;
  output \g326395/_0_  ;
  output \g326396/_0_  ;
  output \g326397/_0_  ;
  output \g326398/_0_  ;
  output \g326399/_0_  ;
  output \g326400/_0_  ;
  output \g326401/_0_  ;
  output \g326423/_0_  ;
  output \g326438/_0_  ;
  output \g326439/_0_  ;
  output \g326440/_0_  ;
  output \g326441/_0_  ;
  output \g326442/_0_  ;
  output \g326443/_0_  ;
  output \g326444/_0_  ;
  output \g326445/_0_  ;
  output \g326446/_0_  ;
  output \g326447/_0_  ;
  output \g326448/_0_  ;
  output \g326449/_0_  ;
  output \g326450/_0_  ;
  output \g326451/_0_  ;
  output \g326452/_0_  ;
  output \g326561/_0_  ;
  output \g326571/_0_  ;
  output \g326572/_0_  ;
  output \g326597/_0_  ;
  output \g326598/_0_  ;
  output \g326599/_0_  ;
  output \g326600/_0_  ;
  output \g326601/_0_  ;
  output \g326602/_0_  ;
  output \g326603/_0_  ;
  output \g326604/_0_  ;
  output \g326605/_0_  ;
  output \g326606/_0_  ;
  output \g326607/_0_  ;
  output \g326608/_0_  ;
  output \g326609/_0_  ;
  output \g326611/_0_  ;
  output \g326612/_0_  ;
  output \g326613/_0_  ;
  output \g326614/_0_  ;
  output \g326615/_0_  ;
  output \g326616/_0_  ;
  output \g326617/_0_  ;
  output \g326618/_0_  ;
  output \g326619/_0_  ;
  output \g326620/_0_  ;
  output \g326621/_0_  ;
  output \g326622/_0_  ;
  output \g326623/_0_  ;
  output \g326624/_0_  ;
  output \g326625/_0_  ;
  output \g326626/_0_  ;
  output \g326627/_0_  ;
  output \g326628/_0_  ;
  output \g326629/_0_  ;
  output \g326630/_0_  ;
  output \g326631/_0_  ;
  output \g326632/_0_  ;
  output \g326633/_0_  ;
  output \g326634/_0_  ;
  output \g326635/_0_  ;
  output \g326636/_0_  ;
  output \g326637/_0_  ;
  output \g326638/_0_  ;
  output \g326639/_0_  ;
  output \g326640/_0_  ;
  output \g326641/_0_  ;
  output \g326798/_0_  ;
  output \g326821/_0_  ;
  output \g326822/_0_  ;
  output \g326823/_0_  ;
  output \g326824/_0_  ;
  output \g326825/_0_  ;
  output \g326826/_0_  ;
  output \g326827/_0_  ;
  output \g326828/_0_  ;
  output \g326829/_0_  ;
  output \g326830/_0_  ;
  output \g326831/_0_  ;
  output \g326832/_0_  ;
  output \g326833/_0_  ;
  output \g326834/_0_  ;
  output \g326835/_0_  ;
  output \g326868/_0_  ;
  output \g326887/_0_  ;
  output \g326926/_0_  ;
  output \g326927/_0_  ;
  output \g326928/_0_  ;
  output \g326929/_0_  ;
  output \g326930/_0_  ;
  output \g326931/_0_  ;
  output \g326932/_0_  ;
  output \g326933/_0_  ;
  output \g326934/_0_  ;
  output \g326935/_0_  ;
  output \g326936/_0_  ;
  output \g326937/_0_  ;
  output \g326938/_0_  ;
  output \g326939/_0_  ;
  output \g326940/_0_  ;
  output \g326941/_0_  ;
  output \g326942/_0_  ;
  output \g326943/_0_  ;
  output \g326944/_0_  ;
  output \g326945/_0_  ;
  output \g326946/_0_  ;
  output \g326947/_0_  ;
  output \g326948/_0_  ;
  output \g326949/_0_  ;
  output \g326950/_0_  ;
  output \g326951/_0_  ;
  output \g326952/_0_  ;
  output \g326953/_0_  ;
  output \g326954/_0_  ;
  output \g326955/_0_  ;
  output \g327192/_0_  ;
  output \g327234/_0_  ;
  output \g327237/_0_  ;
  output \g327241/_0_  ;
  output \g327242/_0_  ;
  output \g327243/_0_  ;
  output \g327247/_0_  ;
  output \g327290/_0_  ;
  output \g327311/_0_  ;
  output \g327369/_0_  ;
  output \g327370/_0_  ;
  output \g327371/_0_  ;
  output \g327373/_0_  ;
  output \g327375/_0_  ;
  output \g327377/_0_  ;
  output \g327379/_0_  ;
  output \g327380/_0_  ;
  output \g327381/_0_  ;
  output \g327382/_0_  ;
  output \g327383/_0_  ;
  output \g327384/_0_  ;
  output \g327385/_0_  ;
  output \g327386/_0_  ;
  output \g327387/_0_  ;
  output \g327388/_0_  ;
  output \g327389/_0_  ;
  output \g327390/_0_  ;
  output \g327391/_0_  ;
  output \g327392/_0_  ;
  output \g327393/_0_  ;
  output \g327394/_0_  ;
  output \g327395/_0_  ;
  output \g327396/_0_  ;
  output \g327397/_0_  ;
  output \g327398/_0_  ;
  output \g327399/_0_  ;
  output \g327400/_0_  ;
  output \g327401/_0_  ;
  output \g327402/_0_  ;
  output \g327601/_0_  ;
  output \g327602/_0_  ;
  output \g327698/_0_  ;
  output \g327781/_0_  ;
  output \g327798/_0_  ;
  output \g327799/_0_  ;
  output \g327800/_0_  ;
  output \g327801/_0_  ;
  output \g327802/_0_  ;
  output \g327803/_0_  ;
  output \g327804/_0_  ;
  output \g327805/_0_  ;
  output \g327806/_0_  ;
  output \g327807/_0_  ;
  output \g327826/_0_  ;
  output \g327828/_0_  ;
  output \g327829/_0_  ;
  output \g327830/_0_  ;
  output \g327831/_0_  ;
  output \g327832/_0_  ;
  output \g327833/_0_  ;
  output \g327834/_0_  ;
  output \g327835/_0_  ;
  output \g327836/_0_  ;
  output \g327970/_0_  ;
  output \g328019/_0_  ;
  output \g328020/_0_  ;
  output \g328021/_0_  ;
  output \g328022/_0_  ;
  output \g328023/_0_  ;
  output \g328024/_0_  ;
  output \g328027/_0_  ;
  output \g328028/_0_  ;
  output \g328029/_0_  ;
  output \g328030/_0_  ;
  output \g328031/_0_  ;
  output \g328032/_0_  ;
  output \g328033/_0_  ;
  output \g328034/_0_  ;
  output \g328035/_0_  ;
  output \g328046/_0_  ;
  output \g328048/_0_  ;
  output \g328049/_0_  ;
  output \g328052/_0_  ;
  output \g328054/_0_  ;
  output \g328056/_0_  ;
  output \g328058/_0_  ;
  output \g328059/_0_  ;
  output \g328060/_0_  ;
  output \g328061/_0_  ;
  output \g328062/_0_  ;
  output \g328063/_0_  ;
  output \g328064/_0_  ;
  output \g328065/_0_  ;
  output \g328066/_0_  ;
  output \g328067/_0_  ;
  output \g328068/_0_  ;
  output \g328069/_0_  ;
  output \g328070/_0_  ;
  output \g328071/_0_  ;
  output \g328120/_0_  ;
  output \g328152/_0_  ;
  output \g328153/_0_  ;
  output \g328154/_0_  ;
  output \g328155/_0_  ;
  output \g328156/_0_  ;
  output \g328157/_0_  ;
  output \g328158/_0_  ;
  output \g328159/_0_  ;
  output \g328160/_0_  ;
  output \g328161/_0_  ;
  output \g328257/_0_  ;
  output \g328280/_0_  ;
  output \g328302/_0_  ;
  output \g328303/_0_  ;
  output \g328332/_0_  ;
  output \g328333/_0_  ;
  output \g328334/_0_  ;
  output \g328335/_0_  ;
  output \g328336/_0_  ;
  output \g328337/_0_  ;
  output \g328338/_0_  ;
  output \g328339/_0_  ;
  output \g328340/_0_  ;
  output \g328341/_0_  ;
  output \g328342/_0_  ;
  output \g328343/_0_  ;
  output \g328344/_0_  ;
  output \g328345/_0_  ;
  output \g328346/_0_  ;
  output \g328347/_0_  ;
  output \g328348/_0_  ;
  output \g328349/_0_  ;
  output \g328350/_0_  ;
  output \g328351/_0_  ;
  output \g328352/_0_  ;
  output \g328353/_0_  ;
  output \g328354/_0_  ;
  output \g328355/_0_  ;
  output \g328356/_0_  ;
  output \g328357/_0_  ;
  output \g328358/_0_  ;
  output \g328359/_0_  ;
  output \g328360/_0_  ;
  output \g328361/_0_  ;
  output \g328372/_0_  ;
  output \g328373/_0_  ;
  output \g328374/_0_  ;
  output \g328375/_0_  ;
  output \g328376/_0_  ;
  output \g328377/_0_  ;
  output \g328378/_0_  ;
  output \g328379/_0_  ;
  output \g328380/_0_  ;
  output \g328381/_0_  ;
  output \g328382/_0_  ;
  output \g328383/_0_  ;
  output \g328384/_0_  ;
  output \g328385/_0_  ;
  output \g328569/_0_  ;
  output \g328587/_0_  ;
  output \g328658/_0_  ;
  output \g328662/_3_  ;
  output \g328664/_3_  ;
  output \g328666/_3_  ;
  output \g328669/_3_  ;
  output \g328670/_0_  ;
  output \g328671/_0_  ;
  output \g328672/_0_  ;
  output \g328674/_0_  ;
  output \g328809/_0_  ;
  output \g328810/_0_  ;
  output \g328811/_0_  ;
  output \g328812/_0_  ;
  output \g328856/_0_  ;
  output \g328887/_0_  ;
  output \g328931/_0_  ;
  output \g328945/_0_  ;
  output \g328960/_0_  ;
  output \g328991/_0_  ;
  output \g328992/_0_  ;
  output \g329022/_3_  ;
  output \g329024/_3_  ;
  output \g329025/_0_  ;
  output \g329026/_0_  ;
  output \g329027/_0_  ;
  output \g329029/_3_  ;
  output \g329030/_0_  ;
  output \g329032/_0_  ;
  output \g329033/_0_  ;
  output \g329034/_0_  ;
  output \g329182/_0_  ;
  output \g329228/_0_  ;
  output \g329281/_0_  ;
  output \g329301/_0_  ;
  output \g329302/_0_  ;
  output \g329322/_2_  ;
  output \g329324/_3_  ;
  output \g329334/_3_  ;
  output \g329336/_3_  ;
  output \g329338/_3_  ;
  output \g329340/_2_  ;
  output \g329342/_3_  ;
  output \g329343/_0_  ;
  output \g329345/_3_  ;
  output \g329347/_3_  ;
  output \g329349/_3_  ;
  output \g329351/_3_  ;
  output \g329353/_3_  ;
  output \g329355/_3_  ;
  output \g329357/_3_  ;
  output \g329359/_3_  ;
  output \g329360/_0_  ;
  output \g329362/_3_  ;
  output \g329364/_3_  ;
  output \g329366/_3_  ;
  output \g329368/_3_  ;
  output \g329370/_3_  ;
  output \g329372/_3_  ;
  output \g329374/_3_  ;
  output \g329376/_3_  ;
  output \g329378/_3_  ;
  output \g329379/_0_  ;
  output \g329380/_0_  ;
  output \g329381/_0_  ;
  output \g329388/_0_  ;
  output \g329516/_0_  ;
  output \g329517/_0_  ;
  output \g329518/_0_  ;
  output \g329587/_0_  ;
  output \g329605/_0_  ;
  output \g329687/_0_  ;
  output \g329703/_0_  ;
  output \g329709/_3_  ;
  output \g329716/_3_  ;
  output \g329718/_3_  ;
  output \g329720/_3_  ;
  output \g329722/_3_  ;
  output \g329724/_3_  ;
  output \g329725/_0_  ;
  output \g329727/_0_  ;
  output \g329805/_0_  ;
  output \g329807/_0_  ;
  output \g329809/_0_  ;
  output \g329810/_0_  ;
  output \g329811/_0_  ;
  output \g329812/_0_  ;
  output \g330065/_3_  ;
  output \g330067/_3_  ;
  output \g330069/_3_  ;
  output \g330071/_3_  ;
  output \g330073/_3_  ;
  output \g330075/_3_  ;
  output \g330077/_3_  ;
  output \g330079/_3_  ;
  output \g330081/_3_  ;
  output \g330083/_3_  ;
  output \g330085/_3_  ;
  output \g330087/_3_  ;
  output \g330089/_3_  ;
  output \g330091/_3_  ;
  output \g330093/_3_  ;
  output \g330095/_3_  ;
  output \g330097/_3_  ;
  output \g330099/_0_  ;
  output \g330188/_0_  ;
  output \g330337/_0_  ;
  output \g330388/_3_  ;
  output \g330418/_3_  ;
  output \g330420/_3_  ;
  output \g330422/_3_  ;
  output \g330424/_3_  ;
  output \g330426/_3_  ;
  output \g330428/_3_  ;
  output \g330429/_0_  ;
  output \g330431/_3_  ;
  output \g330433/_3_  ;
  output \g330435/_3_  ;
  output \g330436/_0_  ;
  output \g330438/_3_  ;
  output \g330440/_3_  ;
  output \g330441/_0_  ;
  output \g330443/_3_  ;
  output \g330444/_0_  ;
  output \g330446/_3_  ;
  output \g330448/_3_  ;
  output \g330450/_3_  ;
  output \g330451/_0_  ;
  output \g330452/_0_  ;
  output \g330453/_0_  ;
  output \g330535/_0_  ;
  output \g330762/_3_  ;
  output \g330764/_3_  ;
  output \g330766/_3_  ;
  output \g330768/_3_  ;
  output \g330770/_3_  ;
  output \g330772/_3_  ;
  output \g330774/_3_  ;
  output \g330776/_3_  ;
  output \g331141/_3_  ;
  output \g331142/_0_  ;
  output \g331144/_3_  ;
  output \g331145/_0_  ;
  output \g331147/_3_  ;
  output \g331484/_0_  ;
  output \g331485/_0_  ;
  output \g331486/_0_  ;
  output \g331497/_0_  ;
  output \g331498/_0_  ;
  output \g331502/_0_  ;
  output \g332061/_0_  ;
  output \g332062/_0_  ;
  output \g332063/_0_  ;
  output \g332064/_0_  ;
  output \g332065/_0_  ;
  output \g332066/_0_  ;
  output \g332070/_0_  ;
  output \g332071/_0_  ;
  output \g332672/_0_  ;
  output \g332673/_0_  ;
  output \g332678/_0_  ;
  output \g332679/_0_  ;
  output \g332680/_0_  ;
  output \g332681/_0_  ;
  output \g332682/_0_  ;
  output \g332700/_0_  ;
  output \g333449/_0_  ;
  output \g333453/_0_  ;
  output \g333454/_0_  ;
  output \g333462/_0_  ;
  output \g333463/_0_  ;
  output \g334369/_0_  ;
  output \g334370/_0_  ;
  output \g335243/_0_  ;
  output \g335244/_0_  ;
  output \g335965/_0_  ;
  output \g335969/_0_  ;
  output \g336538/_0_  ;
  output \g336539/_0_  ;
  output \g336540/_0_  ;
  output \g336546/_0_  ;
  output \g336551/_0_  ;
  output \g336552/_0_  ;
  output \g336557/_0_  ;
  output \g336558/_0_  ;
  output \g336654/_0_  ;
  output \g336655/_0_  ;
  output \g336656/_0_  ;
  output \g336657/_0_  ;
  output \g336660/_0_  ;
  output \g336850/_0_  ;
  output \g337247/_0_  ;
  output \g337248/_0_  ;
  output \g337249/_0_  ;
  output \g337250/_0_  ;
  output \g337251/_0_  ;
  output \g337629/_0_  ;
  output \g337635/_0_  ;
  output \g337637/_0_  ;
  output \g337879/_0_  ;
  output \g337905/_0_  ;
  output \g337906/_0_  ;
  output \g337907/_0_  ;
  output \g337916/_0_  ;
  output \g337917/_0_  ;
  output \g337946/_0_  ;
  output \g337947/_0_  ;
  output \g337948/_0_  ;
  output \g337949/_0_  ;
  output \g337950/_0_  ;
  output \g338030/_0_  ;
  output \g338034/_0_  ;
  output \g338388/_0_  ;
  output \g338442/_0_  ;
  output \g338443/_0_  ;
  output \g338513/_0_  ;
  output \g338514/_0_  ;
  output \g338750/_0_  ;
  output \g338759/_0_  ;
  output \g338800/_0_  ;
  output \g338801/_0_  ;
  output \g338802/_0_  ;
  output \g338803/_0_  ;
  output \g338804/_0_  ;
  output \g338805/_0_  ;
  output \g338806/_0_  ;
  output \g338807/_0_  ;
  output \g338808/_0_  ;
  output \g338809/_0_  ;
  output \g338810/_0_  ;
  output \g338811/_0_  ;
  output \g338812/_0_  ;
  output \g338813/_0_  ;
  output \g338814/_0_  ;
  output \g338815/_0_  ;
  output \g338816/_0_  ;
  output \g338817/_0_  ;
  output \g338818/_0_  ;
  output \g338819/_0_  ;
  output \g338820/_0_  ;
  output \g338821/_0_  ;
  output \g338822/_0_  ;
  output \g338823/_0_  ;
  output \g338824/_0_  ;
  output \g338825/_0_  ;
  output \g338826/_0_  ;
  output \g338827/_0_  ;
  output \g338828/_0_  ;
  output \g338829/_0_  ;
  output \g338869/_0_  ;
  output \g338886/_0_  ;
  output \g338887/_0_  ;
  output \g338888/_0_  ;
  output \g339020/_0_  ;
  output \g339021/_0_  ;
  output \g339022/_0_  ;
  output \g339023/_0_  ;
  output \g339024/_0_  ;
  output \g339045/_0_  ;
  output \g339060/_0_  ;
  output \g339125/_0_  ;
  output \g339142/_0_  ;
  output \g339143/_0_  ;
  output \g339144/_0_  ;
  output \g339145/_0_  ;
  output \g339146/_0_  ;
  output \g339147/_0_  ;
  output \g339148/_0_  ;
  output \g339149/_0_  ;
  output \g339150/_0_  ;
  output \g339151/_0_  ;
  output \g339152/_0_  ;
  output \g339153/_0_  ;
  output \g339154/_0_  ;
  output \g339155/_0_  ;
  output \g339156/_0_  ;
  output \g339157/_0_  ;
  output \g339158/_0_  ;
  output \g339159/_0_  ;
  output \g339160/_0_  ;
  output \g339161/_0_  ;
  output \g339162/_0_  ;
  output \g339163/_0_  ;
  output \g339164/_0_  ;
  output \g339165/_0_  ;
  output \g339166/_0_  ;
  output \g339167/_0_  ;
  output \g339168/_0_  ;
  output \g339169/_0_  ;
  output \g339170/_0_  ;
  output \g339171/_0_  ;
  output \g339254/_0_  ;
  output \g339255/_0_  ;
  output \g339257/_0_  ;
  output \g339458/_0_  ;
  output \g339459/_0_  ;
  output \g339460/_0_  ;
  output \g339461/_0_  ;
  output \g339462/_0_  ;
  output \g339463/_0_  ;
  output \g339464/_0_  ;
  output \g339466/_0_  ;
  output \g339469/_0_  ;
  output \g339470/_0_  ;
  output \g339472/_0_  ;
  output \g339504/_0_  ;
  output \g339505/_0_  ;
  output \g339535/_0_  ;
  output \g339601/_0_  ;
  output \g339614/_0_  ;
  output \g339615/_0_  ;
  output \g339616/_0_  ;
  output \g339617/_0_  ;
  output \g339618/_0_  ;
  output \g339619/_0_  ;
  output \g339620/_0_  ;
  output \g339621/_0_  ;
  output \g339622/_0_  ;
  output \g339623/_0_  ;
  output \g339624/_0_  ;
  output \g339625/_0_  ;
  output \g339626/_0_  ;
  output \g339627/_0_  ;
  output \g339628/_0_  ;
  output \g339629/_0_  ;
  output \g339630/_0_  ;
  output \g339631/_0_  ;
  output \g339632/_0_  ;
  output \g339633/_0_  ;
  output \g339634/_0_  ;
  output \g339635/_0_  ;
  output \g339636/_0_  ;
  output \g339637/_0_  ;
  output \g339638/_0_  ;
  output \g339639/_0_  ;
  output \g339640/_0_  ;
  output \g339641/_0_  ;
  output \g339642/_0_  ;
  output \g339643/_0_  ;
  output \g339644/_0_  ;
  output \g339645/_0_  ;
  output \g339646/_0_  ;
  output \g339647/_0_  ;
  output \g339648/_0_  ;
  output \g339649/_0_  ;
  output \g339650/_0_  ;
  output \g339651/_0_  ;
  output \g339652/_0_  ;
  output \g339653/_0_  ;
  output \g339654/_0_  ;
  output \g339655/_0_  ;
  output \g339656/_0_  ;
  output \g339657/_0_  ;
  output \g339658/_0_  ;
  output \g339718/_0_  ;
  output \g339719/_0_  ;
  output \g339720/_0_  ;
  output \g339721/_0_  ;
  output \g339723/_0_  ;
  output \g339725/_0_  ;
  output \g339727/_0_  ;
  output \g340058/_0_  ;
  output \g340102/_0_  ;
  output \g340103/_0_  ;
  output \g340104/_0_  ;
  output \g340106/_0_  ;
  output \g340109/_0_  ;
  output \g340244/_0_  ;
  output \g340245/_0_  ;
  output \g340246/_0_  ;
  output \g340247/_0_  ;
  output \g340464/_0_  ;
  output \g340505/_0_  ;
  output \g340612/_0_  ;
  output \g340613/_0_  ;
  output \g340614/_0_  ;
  output \g340615/_0_  ;
  output \g340616/_0_  ;
  output \g340617/_0_  ;
  output \g340618/_0_  ;
  output \g340619/_0_  ;
  output \g340620/_0_  ;
  output \g340621/_0_  ;
  output \g340622/_0_  ;
  output \g340623/_0_  ;
  output \g340624/_0_  ;
  output \g340625/_0_  ;
  output \g340626/_0_  ;
  output \g340630/_0_  ;
  output \g340631/_0_  ;
  output \g340632/_0_  ;
  output \g340633/_0_  ;
  output \g340634/_0_  ;
  output \g340635/_0_  ;
  output \g340636/_0_  ;
  output \g340637/_0_  ;
  output \g340638/_0_  ;
  output \g340640/_0_  ;
  output \g340641/_0_  ;
  output \g340642/_0_  ;
  output \g340643/_0_  ;
  output \g340644/_0_  ;
  output \g340645/_0_  ;
  output \g340701/_0_  ;
  output \g340702/_0_  ;
  output \g340703/_0_  ;
  output \g340704/_0_  ;
  output \g340714/_0_  ;
  output \g340716/_0_  ;
  output \g340717/_0_  ;
  output \g340718/_0_  ;
  output \g340728/_0_  ;
  output \g340729/_0_  ;
  output \g340730/_0_  ;
  output \g340731/_0_  ;
  output \g340747/_0_  ;
  output \g340748/_0_  ;
  output \g340749/_0_  ;
  output \g340750/_0_  ;
  output \g340751/_0_  ;
  output \g340752/_0_  ;
  output \g340753/_0_  ;
  output \g340754/_0_  ;
  output \g340792/_0_  ;
  output \g340793/_0_  ;
  output \g340794/_0_  ;
  output \g340795/_0_  ;
  output \g340796/_0_  ;
  output \g340797/_0_  ;
  output \g340988/_0_  ;
  output \g341033/_0_  ;
  output \g341191/_0_  ;
  output \g341192/_0_  ;
  output \g341193/_0_  ;
  output \g341194/_0_  ;
  output \g341195/_0_  ;
  output \g341196/_0_  ;
  output \g341197/_0_  ;
  output \g341198/_0_  ;
  output \g341199/_0_  ;
  output \g341200/_0_  ;
  output \g341201/_0_  ;
  output \g341202/_0_  ;
  output \g341203/_0_  ;
  output \g341205/_0_  ;
  output \g341206/_0_  ;
  output \g341207/_0_  ;
  output \g341208/_0_  ;
  output \g341209/_0_  ;
  output \g341210/_0_  ;
  output \g341211/_0_  ;
  output \g341212/_0_  ;
  output \g341213/_0_  ;
  output \g341214/_0_  ;
  output \g341215/_0_  ;
  output \g341216/_0_  ;
  output \g341217/_0_  ;
  output \g341218/_0_  ;
  output \g341219/_0_  ;
  output \g341220/_0_  ;
  output \g341221/_0_  ;
  output \g341241/_0_  ;
  output \g341242/_0_  ;
  output \g341245/_0_  ;
  output \g341248/_0_  ;
  output \g341250/_0_  ;
  output \g341251/_0_  ;
  output \g341339/_0_  ;
  output \g341347/_0_  ;
  output \g341349/_0_  ;
  output \g341350/_0_  ;
  output \g341352/_0_  ;
  output \g341353/_0_  ;
  output \g341354/_0_  ;
  output \g341365/_0_  ;
  output \g341366/_0_  ;
  output \g341367/_0_  ;
  output \g341368/_0_  ;
  output \g341369/_0_  ;
  output \g341370/_0_  ;
  output \g341373/_0_  ;
  output \g341388/_0_  ;
  output \g341389/_0_  ;
  output \g341390/_0_  ;
  output \g341391/_0_  ;
  output \g341392/_0_  ;
  output \g341393/_0_  ;
  output \g341394/_0_  ;
  output \g341395/_0_  ;
  output \g341396/_0_  ;
  output \g341397/_0_  ;
  output \g341398/_0_  ;
  output \g341400/_0_  ;
  output \g341401/_0_  ;
  output \g341419/_0_  ;
  output \g341435/_0_  ;
  output \g341436/_0_  ;
  output \g341455/_0_  ;
  output \g341456/_0_  ;
  output \g341457/_0_  ;
  output \g341458/_0_  ;
  output \g342136/_0_  ;
  output \g342137/_0_  ;
  output \g342141/_0_  ;
  output \g342145/_0_  ;
  output \g342148/_0_  ;
  output \g342149/_0_  ;
  output \g342308/_0_  ;
  output \g342318/_0_  ;
  output \g342322/_0_  ;
  output \g342323/_0_  ;
  output \g342327/_0_  ;
  output \g342331/_0_  ;
  output \g342333/_0_  ;
  output \g342354/_0_  ;
  output \g342355/_0_  ;
  output \g342356/_0_  ;
  output \g342357/_0_  ;
  output \g342358/_0_  ;
  output \g342359/_0_  ;
  output \g342383/_0_  ;
  output \g342384/_0_  ;
  output \g342385/_0_  ;
  output \g342386/_0_  ;
  output \g342387/_0_  ;
  output \g342388/_0_  ;
  output \g342389/_0_  ;
  output \g342390/_0_  ;
  output \g342391/_0_  ;
  output \g342392/_0_  ;
  output \g342393/_0_  ;
  output \g342394/_0_  ;
  output \g342397/_0_  ;
  output \g342398/_0_  ;
  output \g342399/_0_  ;
  output \g342400/_0_  ;
  output \g342401/_0_  ;
  output \g342454/u3_syn_4  ;
  output \g342800/_0_  ;
  output \g343406/_0_  ;
  output \g343407/_0_  ;
  output \g343408/_0_  ;
  output \g343409/_0_  ;
  output \g343410/_0_  ;
  output \g343411/_0_  ;
  output \g343412/_0_  ;
  output \g343413/_0_  ;
  output \g343414/_0_  ;
  output \g343415/_0_  ;
  output \g343416/_0_  ;
  output \g343417/_0_  ;
  output \g343418/_0_  ;
  output \g343419/_0_  ;
  output \g343420/_0_  ;
  output \g343431/_0_  ;
  output \g343432/_0_  ;
  output \g343433/_0_  ;
  output \g343434/_0_  ;
  output \g343435/_0_  ;
  output \g343436/_0_  ;
  output \g343437/_0_  ;
  output \g343439/_0_  ;
  output \g343440/_0_  ;
  output \g343441/_0_  ;
  output \g343443/_0_  ;
  output \g343444/_0_  ;
  output \g343445/_0_  ;
  output \g343446/_0_  ;
  output \g343447/_0_  ;
  output \g343452/_0_  ;
  output \g343453/_0_  ;
  output \g343454/_0_  ;
  output \g343455/_0_  ;
  output \g343456/_0_  ;
  output \g343458/_0_  ;
  output \g343459/_0_  ;
  output \g343460/_0_  ;
  output \g343461/_0_  ;
  output \g343462/_0_  ;
  output \g343463/_0_  ;
  output \g343464/_0_  ;
  output \g343465/_0_  ;
  output \g343466/_0_  ;
  output \g343467/_0_  ;
  output \g343512/_0_  ;
  output \g343514/_0_  ;
  output \g343515/_0_  ;
  output \g343517/_0_  ;
  output \g343524/_0_  ;
  output \g343531/_0_  ;
  output \g343533/_0_  ;
  output \g343534/_0_  ;
  output \g343535/_0_  ;
  output \g343536/_0_  ;
  output \g343537/_0_  ;
  output \g343555/_0_  ;
  output \g343556/_0_  ;
  output \g343557/_0_  ;
  output \g343558/_0_  ;
  output \g343559/_0_  ;
  output \g343560/_0_  ;
  output \g343561/_0_  ;
  output \g343563/_0_  ;
  output \g343564/_0_  ;
  output \g343566/_0_  ;
  output \g343567/_0_  ;
  output \g343568/_0_  ;
  output \g343569/_0_  ;
  output \g343570/_0_  ;
  output \g343699/_0_  ;
  output \g343703/_0_  ;
  output \g343944/_0_  ;
  output \g343992/_0_  ;
  output \g344429/_0_  ;
  output \g344430/_0_  ;
  output \g344431/_0_  ;
  output \g344432/_0_  ;
  output \g344433/_0_  ;
  output \g344434/_0_  ;
  output \g344435/_0_  ;
  output \g344437/_0_  ;
  output \g344438/_0_  ;
  output \g344439/_0_  ;
  output \g344440/_0_  ;
  output \g344441/_0_  ;
  output \g344442/_0_  ;
  output \g344443/_0_  ;
  output \g344444/_0_  ;
  output \g344447/_0_  ;
  output \g344448/_0_  ;
  output \g344449/_0_  ;
  output \g344450/_0_  ;
  output \g344451/_0_  ;
  output \g344452/_0_  ;
  output \g344453/_0_  ;
  output \g344454/_0_  ;
  output \g344455/_0_  ;
  output \g344456/_0_  ;
  output \g344457/_0_  ;
  output \g344458/_0_  ;
  output \g344459/_0_  ;
  output \g344460/_0_  ;
  output \g344461/_0_  ;
  output \g344495/_0_  ;
  output \g344496/_0_  ;
  output \g344497/_0_  ;
  output \g344498/_0_  ;
  output \g344499/_0_  ;
  output \g344500/_0_  ;
  output \g344501/_0_  ;
  output \g344502/_0_  ;
  output \g344503/_0_  ;
  output \g344504/_0_  ;
  output \g344505/_0_  ;
  output \g344506/_0_  ;
  output \g344507/_0_  ;
  output \g344508/_0_  ;
  output \g344511/_0_  ;
  output \g344512/_0_  ;
  output \g344513/_0_  ;
  output \g344514/_0_  ;
  output \g344515/_0_  ;
  output \g344516/_0_  ;
  output \g344517/_0_  ;
  output \g344523/_0_  ;
  output \g344524/_0_  ;
  output \g344525/_0_  ;
  output \g344526/_0_  ;
  output \g344527/_0_  ;
  output \g344528/_0_  ;
  output \g344529/_0_  ;
  output \g344536/_0_  ;
  output \g344537/_0_  ;
  output \g344538/_0_  ;
  output \g344539/_0_  ;
  output \g344540/_0_  ;
  output \g344541/_0_  ;
  output \g344542/_0_  ;
  output \g344543/_0_  ;
  output \g344545/_0_  ;
  output \g344546/_0_  ;
  output \g344547/_0_  ;
  output \g344548/_0_  ;
  output \g344549/_0_  ;
  output \g344550/_0_  ;
  output \g344711/_0_  ;
  output \g344712/_0_  ;
  output \g344729/_0_  ;
  output \g344737/_0_  ;
  output \g344738/_0_  ;
  output \g344783/_0_  ;
  output \g344784/_0_  ;
  output \g344786/_0_  ;
  output \g344791/_0_  ;
  output \g344792/_0_  ;
  output \g344816/_0_  ;
  output \g344819/_0_  ;
  output \g344823/_0_  ;
  output \g344825/_0_  ;
  output \g345116/_0_  ;
  output \g345129/_0_  ;
  output \g345149/_0_  ;
  output \g345161/_0_  ;
  output \g345170/_0_  ;
  output \g345237/_0_  ;
  output \g345313/_0_  ;
  output \g345314/_0_  ;
  output \g345316/_0_  ;
  output \g345317/_0_  ;
  output \g345318/_0_  ;
  output \g345319/_0_  ;
  output \g345320/_0_  ;
  output \g345321/_0_  ;
  output \g345322/_0_  ;
  output \g345323/_0_  ;
  output \g345324/_0_  ;
  output \g345325/_0_  ;
  output \g345326/_0_  ;
  output \g345327/_0_  ;
  output \g345328/_0_  ;
  output \g345329/_0_  ;
  output \g345333/_0_  ;
  output \g345334/_0_  ;
  output \g345335/_0_  ;
  output \g345336/_0_  ;
  output \g345337/_0_  ;
  output \g345338/_0_  ;
  output \g345339/_0_  ;
  output \g345340/_0_  ;
  output \g345349/_0_  ;
  output \g345350/_0_  ;
  output \g345351/_0_  ;
  output \g345352/_0_  ;
  output \g345353/_0_  ;
  output \g345354/_0_  ;
  output \g345355/_0_  ;
  output \g345356/_0_  ;
  output \g345365/_0_  ;
  output \g345366/_0_  ;
  output \g345367/_0_  ;
  output \g345368/_0_  ;
  output \g345369/_0_  ;
  output \g345370/_0_  ;
  output \g345371/_0_  ;
  output \g345373/_0_  ;
  output \g345374/_0_  ;
  output \g345377/_0_  ;
  output \g345378/_0_  ;
  output \g345379/_0_  ;
  output \g345380/_0_  ;
  output \g345381/_0_  ;
  output \g345382/_0_  ;
  output \g345383/_0_  ;
  output \g345488/_0_  ;
  output \g345491/_0_  ;
  output \g345524/_0_  ;
  output \g345525/_0_  ;
  output \g345545/_0_  ;
  output \g345546/_0_  ;
  output \g345574/_0_  ;
  output \g345575/_0_  ;
  output \g345638/_0_  ;
  output \g345639/_0_  ;
  output \g345690/_0_  ;
  output \g345691/_0_  ;
  output \g345692/_0_  ;
  output \g345694/_0_  ;
  output \g345695/_0_  ;
  output \g345698/_0_  ;
  output \g345699/_0_  ;
  output \g345701/_0_  ;
  output \g345703/_0_  ;
  output \g346299/_0_  ;
  output \g346326/_0_  ;
  output \g346364/_0_  ;
  output \g346707/_0_  ;
  output \g346711/_0_  ;
  output \g346721/_0_  ;
  output \g346726/_0_  ;
  output \g346729/_0_  ;
  output \g346730/_0_  ;
  output \g346731/_0_  ;
  output \g346733/_0_  ;
  output \g346735/_0_  ;
  output \g346738/_0_  ;
  output \g346740/_0_  ;
  output \g346741/_0_  ;
  output \g346746/_0_  ;
  output \g346748/_0_  ;
  output \g346750/_0_  ;
  output \g346751/_0_  ;
  output \g346758/_0_  ;
  output \g346759/_0_  ;
  output \g346761/_0_  ;
  output \g346762/_0_  ;
  output \g346763/_0_  ;
  output \g346765/_0_  ;
  output \g346766/_0_  ;
  output \g346965/_0_  ;
  output \g346971/_0_  ;
  output \g346981/_0_  ;
  output \g346986/_0_  ;
  output \g346988/_0_  ;
  output \g346989/_0_  ;
  output \g346994/_0_  ;
  output \g346998/_0_  ;
  output \g347015/_0_  ;
  output \g347016/_0_  ;
  output \g347017/_0_  ;
  output \g347018/_0_  ;
  output \g347019/_0_  ;
  output \g347020/_0_  ;
  output \g347043/_0_  ;
  output \g347050/_0_  ;
  output \g347051/_0_  ;
  output \g347052/_0_  ;
  output \g347053/_0_  ;
  output \g347054/_0_  ;
  output \g347055/_0_  ;
  output \g347056/_0_  ;
  output \g347057/_0_  ;
  output \g347058/_0_  ;
  output \g347059/_0_  ;
  output \g347061/_0_  ;
  output \g347062/_0_  ;
  output \g347063/_0_  ;
  output \g347064/_0_  ;
  output \g347065/_0_  ;
  output \g347066/_0_  ;
  output \g347067/_0_  ;
  output \g347068/_0_  ;
  output \g347069/_0_  ;
  output \g347070/_0_  ;
  output \g347071/_0_  ;
  output \g347083/_0_  ;
  output \g347085/_0_  ;
  output \g347087/_0_  ;
  output \g347089/_0_  ;
  output \g347090/_0_  ;
  output \g347091/_0_  ;
  output \g347092/_0_  ;
  output \g347093/_0_  ;
  output \g347096/_0_  ;
  output \g347097/_0_  ;
  output \g347098/_0_  ;
  output \g347099/_0_  ;
  output \g347100/_0_  ;
  output \g347101/_0_  ;
  output \g347102/_0_  ;
  output \g347104/_0_  ;
  output \g347106/_0_  ;
  output \g347108/_0_  ;
  output \g347318/_0_  ;
  output \g347400/_0_  ;
  output \g347449/_0_  ;
  output \g347477/_0_  ;
  output \g347488/_0_  ;
  output \g347531/_0_  ;
  output \g347537/_0_  ;
  output \g347544/_0_  ;
  output \g347546/_0_  ;
  output \g347553/_0_  ;
  output \g347560/_0_  ;
  output \g347569/_0_  ;
  output \g347575/_0_  ;
  output \g347581/_1_  ;
  output \g347587/_0_  ;
  output \g347592/_0_  ;
  output \g347597/_0_  ;
  output \g347603/_0_  ;
  output \g347610/_0_  ;
  output \g347611/_0_  ;
  output \g347616/_0_  ;
  output \g347624/_0_  ;
  output \g347628/_1_  ;
  output \g347632/_0_  ;
  output \g347641/_0_  ;
  output \g347645/_0_  ;
  output \g347653/_0_  ;
  output \g347661/_0_  ;
  output \g347671/_0_  ;
  output \g347678/_0_  ;
  output \g347881/_0_  ;
  output \g347883/_0_  ;
  output \g347885/_0_  ;
  output \g347886/_0_  ;
  output \g347888/_0_  ;
  output \g347889/_0_  ;
  output \g347890/_0_  ;
  output \g347891/_0_  ;
  output \g347892/_0_  ;
  output \g347893/_0_  ;
  output \g347895/_0_  ;
  output \g347896/_0_  ;
  output \g347897/_0_  ;
  output \g347898/_0_  ;
  output \g347899/_0_  ;
  output \g347902/_0_  ;
  output \g347903/_0_  ;
  output \g347904/_0_  ;
  output \g347906/_0_  ;
  output \g347907/_0_  ;
  output \g347908/_0_  ;
  output \g347909/_0_  ;
  output \g347910/_0_  ;
  output \g347911/_0_  ;
  output \g347912/_0_  ;
  output \g347913/_0_  ;
  output \g347914/_0_  ;
  output \g347915/_0_  ;
  output \g347916/_0_  ;
  output \g347917/_0_  ;
  output \g347974/_0_  ;
  output \g347977/_0_  ;
  output \g347983/_0_  ;
  output \g347999/_0_  ;
  output \g348012/_0_  ;
  output \g348015/_0_  ;
  output \g348288/_0_  ;
  output \g348291/_0_  ;
  output \g348292/_0_  ;
  output \g348293/_0_  ;
  output \g348294/_0_  ;
  output \g348295/_0_  ;
  output \g348296/_0_  ;
  output \g348300/_0_  ;
  output \g348301/_0_  ;
  output \g348302/_0_  ;
  output \g348303/_0_  ;
  output \g348304/_0_  ;
  output \g348307/_0_  ;
  output \g348308/_0_  ;
  output \g349018/_0_  ;
  output \g349020/_0_  ;
  output \g349021/_0_  ;
  output \g349025/_0_  ;
  output \g349026/_0_  ;
  output \g349027/_0_  ;
  output \g349035/_0_  ;
  output \g349036/_0_  ;
  output \g349037/_0_  ;
  output \g349049/_0_  ;
  output \g349050/_0_  ;
  output \g349051/_0_  ;
  output \g349070/_0_  ;
  output \g349071/_0_  ;
  output \g349072/_0_  ;
  output \g349076/_0_  ;
  output \g349077/_0_  ;
  output \g349078/_0_  ;
  output \g349326/_0_  ;
  output \g349333/_0_  ;
  output \g349334/_0_  ;
  output \g349335/_0_  ;
  output \g349343/_0_  ;
  output \g349345/_0_  ;
  output \g349349/_0_  ;
  output \g349350/_0_  ;
  output \g349355/_0_  ;
  output \g349357/_0_  ;
  output \g349358/_0_  ;
  output \g349873/_0_  ;
  output \g350037/_0_  ;
  output \g350042/_0_  ;
  output \g350050/_0_  ;
  output \g350051/_0_  ;
  output \g350089/_0_  ;
  output \g350090/_0_  ;
  output \g350093/_0_  ;
  output \g350094/_0_  ;
  output \g350096/_0_  ;
  output \g350097/_0_  ;
  output \g350165/_0_  ;
  output \g350166/_0_  ;
  output \g350168/_0_  ;
  output \g350170/_0_  ;
  output \g350171/_0_  ;
  output \g350172/_0_  ;
  output \g350173/_0_  ;
  output \g350174/_0_  ;
  output \g350175/_0_  ;
  output \g350176/_0_  ;
  output \g350177/_0_  ;
  output \g350178/_0_  ;
  output \g350179/_0_  ;
  output \g350180/_0_  ;
  output \g350181/_0_  ;
  output \g350183/_0_  ;
  output \g350184/_0_  ;
  output \g350185/_0_  ;
  output \g350186/_0_  ;
  output \g350187/_0_  ;
  output \g350188/_0_  ;
  output \g350189/_0_  ;
  output \g350190/_0_  ;
  output \g350191/_0_  ;
  output \g350192/_0_  ;
  output \g350193/_0_  ;
  output \g350194/_0_  ;
  output \g350195/_0_  ;
  output \g350196/_0_  ;
  output \g350197/_0_  ;
  output \g350198/_0_  ;
  output \g350199/_0_  ;
  output \g350200/_0_  ;
  output \g350201/_0_  ;
  output \g350202/_0_  ;
  output \g350203/_0_  ;
  output \g350204/_0_  ;
  output \g350205/_0_  ;
  output \g350654/_0_  ;
  output \g350655/_0_  ;
  output \g350656/_0_  ;
  output \g350658/_0_  ;
  output \g350660/_0_  ;
  output \g350661/_0_  ;
  output \g350662/_0_  ;
  output \g350663/_0_  ;
  output \g350664/_0_  ;
  output \g350665/_0_  ;
  output \g350666/_0_  ;
  output \g350667/_0_  ;
  output \g350668/_0_  ;
  output \g350669/_0_  ;
  output \g350670/_0_  ;
  output \g350671/_0_  ;
  output \g350672/_0_  ;
  output \g350673/_0_  ;
  output \g350674/_0_  ;
  output \g350675/_0_  ;
  output \g350676/_0_  ;
  output \g350677/_0_  ;
  output \g350678/_0_  ;
  output \g350679/_0_  ;
  output \g350680/_0_  ;
  output \g350681/_0_  ;
  output \g350682/_0_  ;
  output \g350683/_0_  ;
  output \g350684/_0_  ;
  output \g350685/_0_  ;
  output \g350686/_0_  ;
  output \g350687/_0_  ;
  output \g350723/_0_  ;
  output \g350724/_0_  ;
  output \g350725/_0_  ;
  output \g350726/_0_  ;
  output \g350727/_0_  ;
  output \g350728/_0_  ;
  output \g350729/_0_  ;
  output \g350730/_0_  ;
  output \g350731/_0_  ;
  output \g350814/_0_  ;
  output \g350815/_0_  ;
  output \g350816/_0_  ;
  output \g350817/_0_  ;
  output \g350818/_0_  ;
  output \g350819/_0_  ;
  output \g350820/_0_  ;
  output \g350821/_0_  ;
  output \g350822/_0_  ;
  output \g350823/_0_  ;
  output \g350824/_0_  ;
  output \g350825/_0_  ;
  output \g350826/_0_  ;
  output \g350827/_0_  ;
  output \g350828/_0_  ;
  output \g350829/_0_  ;
  output \g350830/_0_  ;
  output \g350831/_0_  ;
  output \g350832/_0_  ;
  output \g350833/_0_  ;
  output \g350834/_0_  ;
  output \g350835/_0_  ;
  output \g350836/_0_  ;
  output \g350839/_0_  ;
  output \g350840/_0_  ;
  output \g350842/_0_  ;
  output \g350843/_0_  ;
  output \g350844/_0_  ;
  output \g350845/_0_  ;
  output \g350846/_0_  ;
  output \g350847/_0_  ;
  output \g350848/_0_  ;
  output \g350849/_0_  ;
  output \g350850/_0_  ;
  output \g350852/_0_  ;
  output \g350853/_0_  ;
  output \g350854/_0_  ;
  output \g350856/_0_  ;
  output \g350857/_0_  ;
  output \g350858/_0_  ;
  output \g350859/_0_  ;
  output \g350860/_0_  ;
  output \g350861/_0_  ;
  output \g350862/_0_  ;
  output \g350863/_0_  ;
  output \g350866/_0_  ;
  output \g350867/_0_  ;
  output \g350868/_0_  ;
  output \g350869/_0_  ;
  output \g350870/_0_  ;
  output \g350871/_0_  ;
  output \g350872/_0_  ;
  output \g350873/_0_  ;
  output \g350874/_0_  ;
  output \g350952/_0_  ;
  output \g350959/_0_  ;
  output \g350961/_0_  ;
  output \g350964/_0_  ;
  output \g350974/_0_  ;
  output \g350977/_0_  ;
  output \g351003/_0_  ;
  output \g351005/_0_  ;
  output \g351037/_0_  ;
  output \g351045/_0_  ;
  output \g351048/_0_  ;
  output \g351129/_0_  ;
  output \g351147/_0_  ;
  output \g351169/_0_  ;
  output \g351171/_0_  ;
  output \g351175/_0_  ;
  output \g351195/_0_  ;
  output \g351196/_0_  ;
  output \g351197/_0_  ;
  output \g351198/_0_  ;
  output \g351201/_0_  ;
  output \g351202/_0_  ;
  output \g351203/_0_  ;
  output \g351204/_0_  ;
  output \g351205/_0_  ;
  output \g351206/_0_  ;
  output \g351207/_0_  ;
  output \g351208/_0_  ;
  output \g351209/_0_  ;
  output \g351210/_0_  ;
  output \g351211/_0_  ;
  output \g351214/_0_  ;
  output \g351215/_0_  ;
  output \g351216/_0_  ;
  output \g351217/_0_  ;
  output \g351218/_0_  ;
  output \g351219/_0_  ;
  output \g351220/_0_  ;
  output \g351221/_0_  ;
  output \g351222/_0_  ;
  output \g351223/_0_  ;
  output \g351224/_0_  ;
  output \g351225/_0_  ;
  output \g351226/_0_  ;
  output \g351227/_0_  ;
  output \g351228/_0_  ;
  output \g351229/_0_  ;
  output \g351230/_0_  ;
  output \g351231/_0_  ;
  output \g351671/_0_  ;
  output \g351699/_0_  ;
  output \g351703/_0_  ;
  output \g351704/_0_  ;
  output \g351709/_0_  ;
  output \g351711/_0_  ;
  output \g351712/_0_  ;
  output \g351715/_0_  ;
  output \g351716/_0_  ;
  output \g351717/_0_  ;
  output \g351721/_0_  ;
  output \g351722/_0_  ;
  output \g351723/_0_  ;
  output \g351724/_0_  ;
  output \g351725/_0_  ;
  output \g351726/_0_  ;
  output \g351727/_0_  ;
  output \g351728/_0_  ;
  output \g351739/_0_  ;
  output \g351741/_0_  ;
  output \g351742/_0_  ;
  output \g351750/_0_  ;
  output \g351752/_0_  ;
  output \g351753/_0_  ;
  output \g351756/_0_  ;
  output \g351757/_0_  ;
  output \g351759/_0_  ;
  output \g351760/_0_  ;
  output \g351761/_0_  ;
  output \g351766/_0_  ;
  output \g351767/_0_  ;
  output \g351768/_0_  ;
  output \g351771/_0_  ;
  output \g351772/_0_  ;
  output \g351773/_0_  ;
  output \g351775/_0_  ;
  output \g351776/_0_  ;
  output \g351779/_0_  ;
  output \g351780/_0_  ;
  output \g351782/_0_  ;
  output \g351785/_0_  ;
  output \g351786/_0_  ;
  output \g351788/_0_  ;
  output \g351789/_0_  ;
  output \g351790/_0_  ;
  output \g351791/_0_  ;
  output \g351792/_0_  ;
  output \g351793/_0_  ;
  output \g351794/_0_  ;
  output \g351795/_0_  ;
  output \g351796/_0_  ;
  output \g351797/_0_  ;
  output \g351798/_0_  ;
  output \g351799/_0_  ;
  output \g351800/_0_  ;
  output \g351801/_0_  ;
  output \g351802/_0_  ;
  output \g351803/_0_  ;
  output \g351804/_0_  ;
  output \g351805/_0_  ;
  output \g351806/_0_  ;
  output \g351807/_0_  ;
  output \g351808/_0_  ;
  output \g351809/_0_  ;
  output \g351810/_0_  ;
  output \g351811/_0_  ;
  output \g351812/_0_  ;
  output \g351814/_0_  ;
  output \g351817/_0_  ;
  output \g351818/_0_  ;
  output \g351819/_0_  ;
  output \g351821/_0_  ;
  output \g351822/_0_  ;
  output \g351823/_0_  ;
  output \g351841/_0_  ;
  output \g351842/_0_  ;
  output \g351843/_0_  ;
  output \g351844/_0_  ;
  output \g351845/_0_  ;
  output \g351846/_0_  ;
  output \g351847/_0_  ;
  output \g351848/_0_  ;
  output \g351849/_0_  ;
  output \g351850/_0_  ;
  output \g351851/_0_  ;
  output \g351852/_0_  ;
  output \g351853/_0_  ;
  output \g351854/_0_  ;
  output \g351855/_0_  ;
  output \g351856/_0_  ;
  output \g351857/_0_  ;
  output \g351858/_0_  ;
  output \g351859/_0_  ;
  output \g351860/_0_  ;
  output \g351861/_0_  ;
  output \g351862/_0_  ;
  output \g351863/_0_  ;
  output \g351864/_0_  ;
  output \g351865/_0_  ;
  output \g351866/_0_  ;
  output \g351867/_0_  ;
  output \g351868/_0_  ;
  output \g351869/_0_  ;
  output \g351870/_0_  ;
  output \g351871/_0_  ;
  output \g351872/_0_  ;
  output \g351873/_0_  ;
  output \g351874/_0_  ;
  output \g351875/_0_  ;
  output \g351876/_0_  ;
  output \g351877/_0_  ;
  output \g351878/_0_  ;
  output \g351879/_0_  ;
  output \g351880/_0_  ;
  output \g351881/_0_  ;
  output \g351882/_0_  ;
  output \g351883/_0_  ;
  output \g351884/_0_  ;
  output \g351885/_0_  ;
  output \g351889/_0_  ;
  output \g351920/_0_  ;
  output \g351921/_0_  ;
  output \g351922/_0_  ;
  output \g351923/_0_  ;
  output \g351924/_0_  ;
  output \g351925/_0_  ;
  output \g351926/_0_  ;
  output \g351927/_0_  ;
  output \g351928/_0_  ;
  output \g351929/_0_  ;
  output \g351930/_0_  ;
  output \g351954/_0_  ;
  output \g351955/_0_  ;
  output \g351956/_0_  ;
  output \g351957/_0_  ;
  output \g352167/_0_  ;
  output \g352178/_0_  ;
  output \g352211/_0_  ;
  output \g352215/_0_  ;
  output \g352219/_0_  ;
  output \g352237/_0_  ;
  output \g352238/_0_  ;
  output \g352239/_0_  ;
  output \g352240/_0_  ;
  output \g352241/_0_  ;
  output \g352242/_0_  ;
  output \g352243/_0_  ;
  output \g352244/_0_  ;
  output \g352245/_0_  ;
  output \g352246/_0_  ;
  output \g352247/_0_  ;
  output \g352248/_0_  ;
  output \g352249/_0_  ;
  output \g352250/_0_  ;
  output \g352251/_0_  ;
  output \g352252/_0_  ;
  output \g352253/_0_  ;
  output \g352254/_0_  ;
  output \g352255/_0_  ;
  output \g352256/_0_  ;
  output \g352257/_0_  ;
  output \g352258/_0_  ;
  output \g352259/_0_  ;
  output \g352260/_0_  ;
  output \g352261/_0_  ;
  output \g352262/_0_  ;
  output \g352263/_0_  ;
  output \g352264/_0_  ;
  output \g352265/_0_  ;
  output \g352266/_0_  ;
  output \g352267/_0_  ;
  output \g352268/_0_  ;
  output \g352269/_0_  ;
  output \g352271/_0_  ;
  output \g352272/_0_  ;
  output \g352273/_0_  ;
  output \g352274/_0_  ;
  output \g352275/_0_  ;
  output \g352276/_0_  ;
  output \g352277/_0_  ;
  output \g352278/_0_  ;
  output \g352279/_0_  ;
  output \g352280/_0_  ;
  output \g352281/_0_  ;
  output \g352282/_0_  ;
  output \g352283/_0_  ;
  output \g352284/_0_  ;
  output \g352285/_0_  ;
  output \g352286/_0_  ;
  output \g352287/_0_  ;
  output \g352288/_0_  ;
  output \g352289/_0_  ;
  output \g352290/_0_  ;
  output \g352291/_0_  ;
  output \g352292/_0_  ;
  output \g352293/_0_  ;
  output \g352294/_0_  ;
  output \g352295/_0_  ;
  output \g352296/_0_  ;
  output \g352297/_0_  ;
  output \g352298/_0_  ;
  output \g352299/_0_  ;
  output \g352300/_0_  ;
  output \g352301/_0_  ;
  output \g352302/_0_  ;
  output \g352303/_0_  ;
  output \g352304/_0_  ;
  output \g352305/_0_  ;
  output \g352306/_0_  ;
  output \g352307/_0_  ;
  output \g352308/_0_  ;
  output \g352309/_0_  ;
  output \g352310/_0_  ;
  output \g352311/_0_  ;
  output \g352312/_0_  ;
  output \g352313/_0_  ;
  output \g352314/_0_  ;
  output \g352315/_0_  ;
  output \g352525/_0_  ;
  output \g352527/_0_  ;
  output \g352529/_0_  ;
  output \g352547/_0_  ;
  output \g352553/_0_  ;
  output \g352554/_0_  ;
  output \g352556/_0_  ;
  output \g352558/_0_  ;
  output \g352559/_0_  ;
  output \g352560/_0_  ;
  output \g352561/_0_  ;
  output \g352563/_0_  ;
  output \g352564/_0_  ;
  output \g352565/_0_  ;
  output \g352567/_0_  ;
  output \g352568/_0_  ;
  output \g352569/_0_  ;
  output \g352570/_0_  ;
  output \g352572/_0_  ;
  output \g352574/_0_  ;
  output \g352575/_0_  ;
  output \g352577/_0_  ;
  output \g352579/_0_  ;
  output \g352581/_0_  ;
  output \g352583/_0_  ;
  output \g352584/_0_  ;
  output \g352585/_0_  ;
  output \g352586/_0_  ;
  output \g352587/_0_  ;
  output \g352588/_0_  ;
  output \g352589/_0_  ;
  output \g352590/_0_  ;
  output \g352591/_0_  ;
  output \g352592/_0_  ;
  output \g352593/_0_  ;
  output \g352594/_0_  ;
  output \g352595/_0_  ;
  output \g352596/_0_  ;
  output \g352597/_0_  ;
  output \g352598/_0_  ;
  output \g352599/_0_  ;
  output \g352600/_0_  ;
  output \g352601/_0_  ;
  output \g352602/_0_  ;
  output \g352603/_0_  ;
  output \g352605/_0_  ;
  output \g352606/_0_  ;
  output \g352607/_0_  ;
  output \g352608/_0_  ;
  output \g352609/_0_  ;
  output \g352610/_0_  ;
  output \g352611/_0_  ;
  output \g352612/_0_  ;
  output \g352613/_0_  ;
  output \g352614/_0_  ;
  output \g352615/_0_  ;
  output \g352616/_0_  ;
  output \g352617/_0_  ;
  output \g352618/_0_  ;
  output \g352619/_0_  ;
  output \g352620/_0_  ;
  output \g352621/_0_  ;
  output \g352622/_0_  ;
  output \g352623/_0_  ;
  output \g352624/_0_  ;
  output \g352625/_0_  ;
  output \g352626/_0_  ;
  output \g352627/_0_  ;
  output \g352628/_0_  ;
  output \g352629/_0_  ;
  output \g352662/_0_  ;
  output \g352663/_0_  ;
  output \g352666/_0_  ;
  output \g352667/_0_  ;
  output \g352668/_0_  ;
  output \g352676/_0_  ;
  output \g352677/_0_  ;
  output \g352678/_0_  ;
  output \g352683/_0_  ;
  output \g352684/_0_  ;
  output \g352685/_0_  ;
  output \g353014/_0_  ;
  output \g353016/_0_  ;
  output \g353035/_0_  ;
  output \g353036/_0_  ;
  output \g353065/_0_  ;
  output \g353067/_0_  ;
  output \g353071/_0_  ;
  output \g353073/_0_  ;
  output \g353085/_0_  ;
  output \g353087/_0_  ;
  output \g353116/_0_  ;
  output \g353119/_0_  ;
  output \g353120/_0_  ;
  output \g353121/_0_  ;
  output \g353122/_0_  ;
  output \g353123/_0_  ;
  output \g353124/_0_  ;
  output \g353125/_0_  ;
  output \g353126/_0_  ;
  output \g353127/_0_  ;
  output \g353128/_0_  ;
  output \g353130/_0_  ;
  output \g353131/_0_  ;
  output \g353132/_0_  ;
  output \g353133/_0_  ;
  output \g353134/_0_  ;
  output \g353135/_0_  ;
  output \g353136/_0_  ;
  output \g353137/_0_  ;
  output \g353138/_0_  ;
  output \g353142/_0_  ;
  output \g353148/_0_  ;
  output \g353149/_0_  ;
  output \g353150/_0_  ;
  output \g353151/_0_  ;
  output \g353152/_0_  ;
  output \g353153/_0_  ;
  output \g353154/_0_  ;
  output \g353155/_0_  ;
  output \g353157/_0_  ;
  output \g353158/_0_  ;
  output \g353159/_0_  ;
  output \g353160/_0_  ;
  output \g353161/_0_  ;
  output \g353162/_0_  ;
  output \g353163/_0_  ;
  output \g353164/_0_  ;
  output \g353165/_0_  ;
  output \g353166/_0_  ;
  output \g353167/_0_  ;
  output \g353168/_0_  ;
  output \g353169/_0_  ;
  output \g353170/_0_  ;
  output \g353171/_0_  ;
  output \g353172/_0_  ;
  output \g353173/_0_  ;
  output \g353174/_0_  ;
  output \g353175/_0_  ;
  output \g353176/_0_  ;
  output \g353177/_0_  ;
  output \g353178/_0_  ;
  output \g353179/_0_  ;
  output \g353180/_0_  ;
  output \g353181/_0_  ;
  output \g353184/_0_  ;
  output \g353185/_0_  ;
  output \g353186/_0_  ;
  output \g353187/_0_  ;
  output \g353188/_0_  ;
  output \g353189/_0_  ;
  output \g353190/_0_  ;
  output \g353191/_0_  ;
  output \g353192/_0_  ;
  output \g353193/_0_  ;
  output \g353194/_0_  ;
  output \g353195/_0_  ;
  output \g353196/_0_  ;
  output \g353197/_0_  ;
  output \g353198/_0_  ;
  output \g353199/_0_  ;
  output \g353200/_0_  ;
  output \g353201/_0_  ;
  output \g353202/_0_  ;
  output \g353203/_0_  ;
  output \g353204/_0_  ;
  output \g353205/_0_  ;
  output \g353206/_0_  ;
  output \g353207/_0_  ;
  output \g353208/_0_  ;
  output \g353209/_0_  ;
  output \g353210/_0_  ;
  output \g353211/_0_  ;
  output \g353212/_0_  ;
  output \g353213/_0_  ;
  output \g353214/_0_  ;
  output \g353215/_0_  ;
  output \g353216/_0_  ;
  output \g353217/_0_  ;
  output \g353218/_0_  ;
  output \g353219/_0_  ;
  output \g353220/_0_  ;
  output \g353221/_0_  ;
  output \g353222/_0_  ;
  output \g353223/_0_  ;
  output \g353224/_0_  ;
  output \g353225/_0_  ;
  output \g353226/_0_  ;
  output \g353227/_0_  ;
  output \g353228/_0_  ;
  output \g353229/_0_  ;
  output \g353230/_0_  ;
  output \g353231/_0_  ;
  output \g353232/_0_  ;
  output \g353233/_0_  ;
  output \g353234/_0_  ;
  output \g353235/_0_  ;
  output \g353236/_0_  ;
  output \g353237/_0_  ;
  output \g353238/_0_  ;
  output \g353239/_0_  ;
  output \g353240/_0_  ;
  output \g353241/_0_  ;
  output \g353242/_0_  ;
  output \g353243/_0_  ;
  output \g353244/_0_  ;
  output \g353245/_0_  ;
  output \g353246/_0_  ;
  output \g353247/_0_  ;
  output \g353248/_0_  ;
  output \g353249/_0_  ;
  output \g353250/_0_  ;
  output \g353251/_0_  ;
  output \g353252/_0_  ;
  output \g353253/_0_  ;
  output \g353254/_0_  ;
  output \g353255/_0_  ;
  output \g353256/_0_  ;
  output \g353257/_0_  ;
  output \g353258/_0_  ;
  output \g353259/_0_  ;
  output \g353260/_0_  ;
  output \g353261/_0_  ;
  output \g353262/_0_  ;
  output \g353263/_0_  ;
  output \g353264/_0_  ;
  output \g353265/_0_  ;
  output \g353266/_0_  ;
  output \g353267/_0_  ;
  output \g353268/_0_  ;
  output \g353269/_0_  ;
  output \g353270/_0_  ;
  output \g353271/_0_  ;
  output \g353272/_0_  ;
  output \g353273/_0_  ;
  output \g353274/_0_  ;
  output \g353275/_0_  ;
  output \g353276/_0_  ;
  output \g353277/_0_  ;
  output \g353278/_0_  ;
  output \g353279/_0_  ;
  output \g353280/_0_  ;
  output \g353281/_0_  ;
  output \g354206/_0_  ;
  output \g354214/_0_  ;
  output \g354216/_0_  ;
  output \g354217/_0_  ;
  output \g354222/_0_  ;
  output \g354278/_0_  ;
  output \g354282/_0_  ;
  output \g354284/_0_  ;
  output \g354289/_0_  ;
  output \g354301/_0_  ;
  output \g354330/_0_  ;
  output \g354331/_0_  ;
  output \g354332/_0_  ;
  output \g354333/_0_  ;
  output \g354335/_0_  ;
  output \g354336/_0_  ;
  output \g354337/_0_  ;
  output \g354338/_0_  ;
  output \g354339/_0_  ;
  output \g354340/_0_  ;
  output \g354341/_0_  ;
  output \g354342/_0_  ;
  output \g354343/_0_  ;
  output \g354344/_0_  ;
  output \g354345/_0_  ;
  output \g354346/_0_  ;
  output \g354358/_0_  ;
  output \g354364/_0_  ;
  output \g354442/_0_  ;
  output \g354444/_0_  ;
  output \g354445/_0_  ;
  output \g354447/_0_  ;
  output \g354448/_0_  ;
  output \g354449/_0_  ;
  output \g354450/_0_  ;
  output \g354451/_0_  ;
  output \g354452/_0_  ;
  output \g354455/_0_  ;
  output \g354456/_0_  ;
  output \g354464/_0_  ;
  output \g354465/_0_  ;
  output \g354466/_0_  ;
  output \g354468/_0_  ;
  output \g354469/_0_  ;
  output \g354470/_0_  ;
  output \g354471/_0_  ;
  output \g354472/_0_  ;
  output \g354473/_0_  ;
  output \g354474/_0_  ;
  output \g354477/_0_  ;
  output \g354478/_0_  ;
  output \g354479/_0_  ;
  output \g354480/_0_  ;
  output \g354482/_0_  ;
  output \g354483/_0_  ;
  output \g354484/_0_  ;
  output \g354485/_0_  ;
  output \g354486/_0_  ;
  output \g354487/_0_  ;
  output \g354488/_0_  ;
  output \g354490/_0_  ;
  output \g354491/_0_  ;
  output \g354492/_0_  ;
  output \g354493/_0_  ;
  output \g354494/_0_  ;
  output \g354495/_0_  ;
  output \g354504/_0_  ;
  output \g354505/_0_  ;
  output \g354506/_0_  ;
  output \g354508/_0_  ;
  output \g354509/_0_  ;
  output \g354510/_0_  ;
  output \g354511/_0_  ;
  output \g354512/_0_  ;
  output \g354513/_0_  ;
  output \g354522/_0_  ;
  output \g354524/_0_  ;
  output \g354525/_0_  ;
  output \g354526/_0_  ;
  output \g354527/_0_  ;
  output \g354920/_1_  ;
  output \g355460/_0_  ;
  output \g355461/_0_  ;
  output \g355463/_0_  ;
  output \g355464/_0_  ;
  output \g355466/_0_  ;
  output \g355467/_0_  ;
  output \g355470/_0_  ;
  output \g355471/_0_  ;
  output \g355475/_0_  ;
  output \g355476/_0_  ;
  output \g355477/_0_  ;
  output \g355479/_0_  ;
  output \g355480/_0_  ;
  output \g355481/_0_  ;
  output \g355482/_0_  ;
  output \g355483/_0_  ;
  output \g355508/_0_  ;
  output \g355509/_0_  ;
  output \g355510/_0_  ;
  output \g355511/_0_  ;
  output \g355512/_0_  ;
  output \g355513/_0_  ;
  output \g355514/_0_  ;
  output \g355515/_0_  ;
  output \g355520/_0_  ;
  output \g355521/_0_  ;
  output \g355523/_0_  ;
  output \g355525/_0_  ;
  output \g355527/_0_  ;
  output \g355530/_0_  ;
  output \g355532/_0_  ;
  output \g355534/_0_  ;
  output \g355564/_0_  ;
  output \g355565/_0_  ;
  output \g355566/_0_  ;
  output \g355567/_0_  ;
  output \g355568/_0_  ;
  output \g355569/_0_  ;
  output \g355570/_0_  ;
  output \g355571/_0_  ;
  output \g355980/_0_  ;
  output \g356052/_0_  ;
  output \g356106/_0_  ;
  output \g356111/_0_  ;
  output \g356114/_0_  ;
  output \g356117/_0_  ;
  output \g356122/_0_  ;
  output \g356126/_0_  ;
  output \g356129/_0_  ;
  output \g356133/_0_  ;
  output \g356142/_0_  ;
  output \g356148/_0_  ;
  output \g356151/_0_  ;
  output \g356155/_0_  ;
  output \g356160/_0_  ;
  output \g356162/_0_  ;
  output \g356165/_0_  ;
  output \g356167/_0_  ;
  output \g356170/_0_  ;
  output \g356174/_0_  ;
  output \g356176/_0_  ;
  output \g356179/_0_  ;
  output \g356183/_0_  ;
  output \g356185/_0_  ;
  output \g356189/_0_  ;
  output \g356193/_0_  ;
  output \g356196/_0_  ;
  output \g356199/_0_  ;
  output \g356202/_0_  ;
  output \g356205/_0_  ;
  output \g356207/_0_  ;
  output \g356210/_0_  ;
  output \g356213/_0_  ;
  output \g356215/_0_  ;
  output \g357046/_0_  ;
  output \g357047/_0_  ;
  output \g357048/_0_  ;
  output \g357051/_0_  ;
  output \g357052/_0_  ;
  output \g357053/_0_  ;
  output \g357054/_0_  ;
  output \g357055/_0_  ;
  output \g357056/_0_  ;
  output \g357057/_0_  ;
  output \g357058/_0_  ;
  output \g357059/_0_  ;
  output \g357060/_0_  ;
  output \g357061/_0_  ;
  output \g357062/_0_  ;
  output \g357063/_0_  ;
  output \g357064/_0_  ;
  output \g357065/_0_  ;
  output \g357066/_0_  ;
  output \g357067/_0_  ;
  output \g357068/_0_  ;
  output \g357069/_0_  ;
  output \g357070/_0_  ;
  output \g357071/_0_  ;
  output \g357072/_0_  ;
  output \g357073/_0_  ;
  output \g357074/_0_  ;
  output \g357099/_0_  ;
  output \g357100/_0_  ;
  output \g357101/_0_  ;
  output \g357102/_0_  ;
  output \g357103/_0_  ;
  output \g357104/_0_  ;
  output \g357105/_0_  ;
  output \g357106/_0_  ;
  output \g357107/_0_  ;
  output \g357108/_0_  ;
  output \g357109/_0_  ;
  output \g357110/_0_  ;
  output \g357111/_0_  ;
  output \g357112/_0_  ;
  output \g357113/_0_  ;
  output \g357114/_0_  ;
  output \g357116/_0_  ;
  output \g357119/_0_  ;
  output \g357121/_0_  ;
  output \g357122/_0_  ;
  output \g357123/_0_  ;
  output \g357124/_0_  ;
  output \g357125/_0_  ;
  output \g357126/_0_  ;
  output \g357128/_0_  ;
  output \g357129/_0_  ;
  output \g357130/_0_  ;
  output \g357131/_0_  ;
  output \g357132/_0_  ;
  output \g357133/_0_  ;
  output \g357134/_0_  ;
  output \g357135/_0_  ;
  output \g357142/_0_  ;
  output \g357144/_0_  ;
  output \g357145/_0_  ;
  output \g357146/_0_  ;
  output \g357147/_0_  ;
  output \g357148/_0_  ;
  output \g357149/_0_  ;
  output \g357150/_0_  ;
  output \g357151/_0_  ;
  output \g357152/_0_  ;
  output \g357153/_0_  ;
  output \g357154/_0_  ;
  output \g357155/_0_  ;
  output \g357156/_0_  ;
  output \g357157/_0_  ;
  output \g357158/_0_  ;
  output \g357160/_0_  ;
  output \g357161/_0_  ;
  output \g357163/_0_  ;
  output \g357164/_0_  ;
  output \g357165/_0_  ;
  output \g357288/_0_  ;
  output \g357289/_0_  ;
  output \g357413/_0_  ;
  output \g357414/_0_  ;
  output \g357464/_0_  ;
  output \g357510/_0_  ;
  output \g357733/_0_  ;
  output \g357769/_0_  ;
  output \g357781/_0_  ;
  output \g357828/_0_  ;
  output \g358792/_0_  ;
  output \g358802/_0_  ;
  output \g359042/_0_  ;
  output \g359043/_0_  ;
  output \g359045/_0_  ;
  output \g359048/_0_  ;
  output \g359051/_0_  ;
  output \g359053/_0_  ;
  output \g359057/_0_  ;
  output \g359060/_0_  ;
  output \g359064/_0_  ;
  output \g359070/_0_  ;
  output \g359074/_0_  ;
  output \g359077/_0_  ;
  output \g359080/_0_  ;
  output \g359086/_0_  ;
  output \g359087/_0_  ;
  output \g359088/_0_  ;
  output \g359090/_0_  ;
  output \g359092/_0_  ;
  output \g359094/_0_  ;
  output \g359096/_0_  ;
  output \g359097/_0_  ;
  output \g359099/_0_  ;
  output \g359101/_0_  ;
  output \g359102/_0_  ;
  output \g359104/_0_  ;
  output \g359106/_0_  ;
  output \g359107/_0_  ;
  output \g359108/_0_  ;
  output \g359110/_0_  ;
  output \g359111/_0_  ;
  output \g359112/_0_  ;
  output \g359113/_0_  ;
  output \g359116/_0_  ;
  output \g359118/_0_  ;
  output \g359572/_0_  ;
  output \g359573/_0_  ;
  output \g359577/_0_  ;
  output \g359585/_0_  ;
  output \g359887/_0_  ;
  output \g359888/_0_  ;
  output \g360077/_0_  ;
  output \g360083/_0_  ;
  output \g360113/_0_  ;
  output \g360124/_0_  ;
  output \g360302/_0_  ;
  output \g360303/_0_  ;
  output \g360304/_0_  ;
  output \g360305/_0_  ;
  output \g360320/_0_  ;
  output \g360325/_0_  ;
  output \g360361/_0_  ;
  output \g360371/_0_  ;
  output \g360440/_0_  ;
  output \g360441/_0_  ;
  output \g360443/_0_  ;
  output \g360445/_0_  ;
  output \g360446/_0_  ;
  output \g360448/_0_  ;
  output \g360450/_0_  ;
  output \g360453/_0_  ;
  output \g360462/_0_  ;
  output \g360469/_0_  ;
  output \g360476/_0_  ;
  output \g360478/_0_  ;
  output \g360480/_0_  ;
  output \g360485/_0_  ;
  output \g360487/_0_  ;
  output \g360489/_0_  ;
  output \g360491/_0_  ;
  output \g360492/_0_  ;
  output \g360494/_0_  ;
  output \g360497/_0_  ;
  output \g360498/_0_  ;
  output \g360504/_0_  ;
  output \g360506/_0_  ;
  output \g360514/_0_  ;
  output \g360516/_0_  ;
  output \g360518/_0_  ;
  output \g360522/_0_  ;
  output \g360524/_0_  ;
  output \g360527/_0_  ;
  output \g360528/_0_  ;
  output \g360530/_0_  ;
  output \g360533/_0_  ;
  output \g360535/_0_  ;
  output \g360538/_0_  ;
  output \g360539/_0_  ;
  output \g360542/_0_  ;
  output \g360546/_0_  ;
  output \g360593/_0_  ;
  output \g361116/_0_  ;
  output \g361128/_0_  ;
  output \g361132/_0_  ;
  output \g361137/_0_  ;
  output \g361616/_0_  ;
  output \g361624/_0_  ;
  output \g361626/_0_  ;
  output \g361627/_0_  ;
  output \g361630/_0_  ;
  output \g361631/_0_  ;
  output \g362129/_0_  ;
  output \g362558/_0_  ;
  output \g362560/_0_  ;
  output \g362564/_0_  ;
  output \g362567/_0_  ;
  output \g362575/_0_  ;
  output \g362586/_0_  ;
  output \g362598/_0_  ;
  output \g362608/_0_  ;
  output \g362627/_0_  ;
  output \g362638/_0_  ;
  output \g362648/_0_  ;
  output \g362650/_0_  ;
  output \g362653/_0_  ;
  output \g362663/_0_  ;
  output \g362664/_0_  ;
  output \g362667/_0_  ;
  output \g362671/_0_  ;
  output \g362673/_0_  ;
  output \g362676/_0_  ;
  output \g362679/_0_  ;
  output \g362686/_0_  ;
  output \g362688/_0_  ;
  output \g362693/_0_  ;
  output \g362697/_0_  ;
  output \g362703/_0_  ;
  output \g363274/_0_  ;
  output \g363290/_0_  ;
  output \g363294/_0_  ;
  output \g363303/_0_  ;
  output \g363608/_0_  ;
  output \g363609/_0_  ;
  output \g363615/_0_  ;
  output \g363616/_0_  ;
  output \g363617/_0_  ;
  output \g363627/_0_  ;
  output \g363818/_3_  ;
  output \g365385/_0_  ;
  output \g365388/_0_  ;
  output \g365391/_0_  ;
  output \g365393/_0_  ;
  output \g365394/_0_  ;
  output \g365398/_0_  ;
  output \g365474/_0_  ;
  output \g365477/_0_  ;
  output \g366167/_0_  ;
  output \g366168/_0_  ;
  output \g366169/_0_  ;
  output \g366170/_0_  ;
  output \g366171/_0_  ;
  output \g366172/_0_  ;
  output \g366173/_0_  ;
  output \g366174/_0_  ;
  output \g366523/_3_  ;
  output \g369170/_0_  ;
  output \g369171/_0_  ;
  output \g369173/_0_  ;
  output \g369177/_0_  ;
  output \g369289/_0_  ;
  output \g369290/_0_  ;
  output \g369291/_0_  ;
  output \g369292/_0_  ;
  output \g369293/_0_  ;
  output \g369294/_0_  ;
  output \g369453/_3_  ;
  output \g371379/_0_  ;
  output \g371381/_0_  ;
  output \g371384/_0_  ;
  output \g371386/_0_  ;
  output \g371387/_0_  ;
  output \g371391/_0_  ;
  output \g372221/_0_  ;
  output \g372222/_0_  ;
  output \g372232/_0_  ;
  output \g372246/_0_  ;
  output \g372249/_0_  ;
  output \g372250/_0_  ;
  output \g372251/_0_  ;
  output \g372252/_0_  ;
  output \g372253/_0_  ;
  output \g372254/_0_  ;
  output \g372454/_3_  ;
  output \g372455/_3_  ;
  output \g372456/_3_  ;
  output \g372457/_3_  ;
  output \g372458/_3_  ;
  output \g372459/_3_  ;
  output \g372460/_3_  ;
  output \g372461/_3_  ;
  output \g372462/_3_  ;
  output \g372463/_3_  ;
  output \g372464/_3_  ;
  output \g372465/_3_  ;
  output \g372466/_3_  ;
  output \g372467/_3_  ;
  output \g372468/_3_  ;
  output \g372469/_3_  ;
  output \g372470/_3_  ;
  output \g372471/_3_  ;
  output \g372472/_3_  ;
  output \g372473/_3_  ;
  output \g372474/_3_  ;
  output \g372475/_3_  ;
  output \g372476/_3_  ;
  output \g372477/_3_  ;
  output \g372478/_3_  ;
  output \g372479/_3_  ;
  output \g372480/_3_  ;
  output \g372481/_3_  ;
  output \g372482/_3_  ;
  output \g372483/_3_  ;
  output \g372484/_3_  ;
  output \g372485/_3_  ;
  output \g372487/_3_  ;
  output \g372488/_3_  ;
  output \g372489/_3_  ;
  output \g372490/_3_  ;
  output \g372491/_3_  ;
  output \g372492/_3_  ;
  output \g372493/_3_  ;
  output \g372494/_3_  ;
  output \g372495/_3_  ;
  output \g372496/_3_  ;
  output \g372497/_3_  ;
  output \g372498/_3_  ;
  output \g372499/_3_  ;
  output \g372500/_3_  ;
  output \g372501/_3_  ;
  output \g372502/_3_  ;
  output \g372503/_3_  ;
  output \g372504/_3_  ;
  output \g372506/_3_  ;
  output \g372507/_3_  ;
  output \g372508/_3_  ;
  output \g372509/_3_  ;
  output \g372510/_3_  ;
  output \g372511/_3_  ;
  output \g372512/_3_  ;
  output \g372513/_3_  ;
  output \g372514/_3_  ;
  output \g372515/_3_  ;
  output \g372516/_3_  ;
  output \g372517/_3_  ;
  output \g372531/_3_  ;
  output \g372532/_3_  ;
  output \g372533/_3_  ;
  output \g374644/_0_  ;
  output \g374645/_0_  ;
  output \g374648/_0_  ;
  output \g374697/_0_  ;
  output \g374701/_0_  ;
  output \g374749/_0_  ;
  output \g374956/_0_  ;
  output \g374961/_0_  ;
  output \g374965/_0_  ;
  output \g374982/_0_  ;
  output \g375071/_0_  ;
  output \g375073/_0_  ;
  output \g375075/_0_  ;
  output \g375078/_0_  ;
  output \g375315/_3_  ;
  output \g375316/_3_  ;
  output \g376101/_0_  ;
  output \g376479/_0_  ;
  output \g377693/_0_  ;
  output \g377694/_0_  ;
  output \g377695/_0_  ;
  output \g377720/_0_  ;
  output \g377721/_0_  ;
  output \g377722/_0_  ;
  output \g378092/_3_  ;
  output \g378093/_3_  ;
  output \g378094/_3_  ;
  output \g378523/_0_  ;
  output \g378524/_0_  ;
  output \g382190/_0_  ;
  output \g382191/_0_  ;
  output \g382192/_0_  ;
  output \g382193/_0_  ;
  output \g382194/_0_  ;
  output \g382195/_0_  ;
  output \g382279/_0_  ;
  output \g382284/_0_  ;
  output \g382292/_0_  ;
  output \g382299/_0_  ;
  output \g382534/_0_  ;
  output \g382535/_0_  ;
  output \g382555/_0_  ;
  output \g382562/_0_  ;
  output \g382563/_0_  ;
  output \g382564/_0_  ;
  output \g382565/_0_  ;
  output \g382571/_0_  ;
  output \g382773/_3_  ;
  output \g382774/_3_  ;
  output \g382775/_3_  ;
  output \g383503/_2_  ;
  output \g383932/_2_  ;
  output \g384194/_0_  ;
  output \g384195/_0_  ;
  output \g384208/_0_  ;
  output \g385644/_0_  ;
  output \g385649/_0_  ;
  output \g385654/_0_  ;
  output \g385672/_0_  ;
  output \g385812/_0_  ;
  output \g385813/_0_  ;
  output \g385816/_0_  ;
  output \g385819/_0_  ;
  output \g386657/_0_  ;
  output \g386660/_0_  ;
  output \g386710/_0_  ;
  output \g386868/_0_  ;
  output \g387282/_0_  ;
  output \g387284/_0_  ;
  output \g387287/_0_  ;
  output \g387292/_0_  ;
  output \g387559/_0_  ;
  output \g387560/_0_  ;
  output \g387561/_0_  ;
  output \g387562/_0_  ;
  output \g387563/_0_  ;
  output \g387564/_0_  ;
  output \g387735/_0_  ;
  output \g387736/_0_  ;
  output \g387738/_0_  ;
  output \g387739/_0_  ;
  output \g387740/_0_  ;
  output \g387743/_0_  ;
  output \g387788/_0_  ;
  output \g387793/_0_  ;
  output \g387796/_0_  ;
  output \g387803/_0_  ;
  output \g388323/_3_  ;
  output \g388332/_3_  ;
  output \g388543/_0_  ;
  output \g388544/_0_  ;
  output \g388545/_0_  ;
  output \g388547/_0_  ;
  output \g388585/_0_  ;
  output \g388694/_0_  ;
  output \g388830/_0_  ;
  output \g388869/_0_  ;
  output \g388998/_0_  ;
  output \g389009/_0_  ;
  output \g389221/_0_  ;
  output \g389225/_0_  ;
  output \g389226/_0_  ;
  output \g389231/_0_  ;
  output \g389234/_0_  ;
  output \g389242/_0_  ;
  output \g389368/_2_  ;
  output \g389368/_2__syn_2  ;
  output \g389369/_2_  ;
  output \g389369/_2__syn_2  ;
  output \g389746/_0_  ;
  output \g389751/_0_  ;
  output \g389774/_0_  ;
  output \g389776/_0_  ;
  output \g389777/_0_  ;
  output \g389779/_0_  ;
  output \g389781/_0_  ;
  output \g389784/_0_  ;
  output \g389787/_0_  ;
  output \g389796/_0_  ;
  output \g389797/_0_  ;
  output \g389801/_0_  ;
  output \g390034/_0_  ;
  output \g390035/_0_  ;
  output \g390037/_0_  ;
  output \g390038/_0_  ;
  output \g390039/_0_  ;
  output \g390043/_0_  ;
  output \g390303/_3_  ;
  output \g390322/_3_  ;
  output \g390323/_3_  ;
  output \g390324/_3_  ;
  output \g390706/_0_  ;
  output \g390876/_0_  ;
  output \g390894/_0_  ;
  output \g390968/_0_  ;
  output \g391050/_0_  ;
  output \g391077/_0_  ;
  output \g392543/_3_  ;
  output \g392565/_3_  ;
  output \g392566/_3_  ;
  output \g394544/_3_  ;
  output \g394545/_3_  ;
  output \g394586/_3_  ;
  output \g395723/_0_  ;
  output \g395757/_0_  ;
  output \g395821/_0_  ;
  output \g395857/_0_  ;
  output \g395858/_0_  ;
  output \g395929/_0_  ;
  output \g396850/_3_  ;
  output \g396876/_3_  ;
  output \g396877/_3_  ;
  output \g397026/_1_  ;
  output \g397035/_1_  ;
  output \g397074/_1_  ;
  output \g397144/_1_  ;
  output \g397344/_1_  ;
  output \g397418/_1_  ;
  output \g397980/_0_  ;
  output \g398209/_0_  ;
  output \g398361/_0_  ;
  output \g398409/_0_  ;
  output \g398458/_0_  ;
  output \g398728/_0_  ;
  output \g401059/_0_  ;
  output \g401066/_0_  ;
  output \g401091/_0_  ;
  output \g401127/_0_  ;
  output \g401160/_0_  ;
  output \g401368/_0_  ;
  output \g401408/_0_  ;
  output \g401455/_0_  ;
  output \g401485/_0_  ;
  output \g401487/_0_  ;
  output \g401506/_0_  ;
  output \g401515/_0_  ;
  output \g401534/_0_  ;
  output \g401549/_0_  ;
  output \g401554/_0_  ;
  output \g401555/_0_  ;
  output \g401592/_0_  ;
  output \g401616/_0_  ;
  output \g401617/_0_  ;
  output \g401618/_0_  ;
  output \g401619/_0_  ;
  output \g401635/_0_  ;
  output \g401657/_0_  ;
  output \g401671/_0_  ;
  output \g401672/_0_  ;
  output \g401684/_0_  ;
  output \g401704/_0_  ;
  output \g401794/_0_  ;
  output \g401807/_0_  ;
  output \g401919/_0_  ;
  output \g401932/_0_  ;
  output \g401935/_0_  ;
  output \g401951/_0_  ;
  output \g401959/_0_  ;
  output \g401961/_0_  ;
  output \g401962/_0_  ;
  output \g401963/_0_  ;
  output \g401998/_0_  ;
  output \g402049/_0_  ;
  output \g402057/_0_  ;
  output \g402063/_0_  ;
  output \g402165/_0_  ;
  output \g402194/_0_  ;
  output \g402298/_0_  ;
  output \g402302/_0_  ;
  output \g402336/_0_  ;
  output \g402346/_0_  ;
  output \g402398/_0_  ;
  output \g402909/_0_  ;
  output \g402910/_0_  ;
  output \g402911/_0_  ;
  output \g402912/_0_  ;
  output \g402913/_0_  ;
  output \g402914/_0_  ;
  output \g403206/_3_  ;
  output \g427842/_1_  ;
  output \g427994/_0_  ;
  output \g428519/_1_  ;
  output \g429040/_1_  ;
  output \g429357/_0_  ;
  output \g429711/_1_  ;
  output \g440733/_0_  ;
  output \g440782/_0_  ;
  output \g441022/_0_  ;
  output \g441242/_0_  ;
  output \g441305/_0_  ;
  output \g441317/_0_  ;
  output \g441329/_0_  ;
  output \g441341/_0_  ;
  output \g441370/_0_  ;
  output \g441382/_0_  ;
  output \g441394/_0_  ;
  output \g441939/_0_  ;
  wire n2790 , n2791 , n2792 , n2793 , n2794 , n2795 , n2796 , n2797 , n2798 , n2799 , n2800 , n2801 , n2802 , n2803 , n2804 , n2805 , n2806 , n2807 , n2808 , n2809 , n2810 , n2811 , n2812 , n2813 , n2814 , n2815 , n2816 , n2817 , n2818 , n2819 , n2820 , n2821 , n2822 , n2823 , n2824 , n2825 , n2826 , n2827 , n2828 , n2829 , n2830 , n2831 , n2832 , n2833 , n2834 , n2835 , n2836 , n2837 , n2838 , n2839 , n2840 , n2841 , n2842 , n2843 , n2844 , n2845 , n2846 , n2847 , n2848 , n2849 , n2850 , n2851 , n2852 , n2853 , n2854 , n2855 , n2856 , n2857 , n2858 , n2859 , n2860 , n2861 , n2862 , n2863 , n2864 , n2865 , n2866 , n2867 , n2868 , n2869 , n2870 , n2871 , n2872 , n2873 , n2874 , n2875 , n2876 , n2877 , n2878 , n2879 , n2880 , n2881 , n2882 , n2883 , n2884 , n2885 , n2886 , n2887 , n2888 , n2889 , n2890 , n2891 , n2892 , n2893 , n2894 , n2895 , n2896 , n2897 , n2898 , n2899 , n2900 , n2901 , n2902 , n2903 , n2904 , n2905 , n2906 , n2907 , n2908 , n2909 , n2910 , n2911 , n2912 , n2913 , n2914 , n2915 , n2916 , n2917 , n2918 , n2919 , n2920 , n2921 , n2922 , n2923 , n2924 , n2925 , n2926 , n2927 , n2928 , n2929 , n2930 , n2931 , n2932 , n2933 , n2934 , n2935 , n2936 , n2937 , n2938 , n2939 , n2940 , n2941 , n2942 , n2943 , n2944 , n2945 , n2946 , n2947 , n2948 , n2949 , n2950 , n2951 , n2952 , n2953 , n2954 , n2955 , n2956 , n2957 , n2958 , n2959 , n2960 , n2961 , n2962 , n2963 , n2964 , n2965 , n2966 , n2967 , n2968 , n2969 , n2970 , n2971 , n2972 , n2973 , n2974 , n2975 , n2976 , n2977 , n2978 , n2979 , n2980 , n2981 , n2982 , n2983 , n2984 , n2985 , n2986 , n2987 , n2988 , n2989 , n2990 , n2991 , n2992 , n2993 , n2994 , n2995 , n2996 , n2997 , n2998 , n2999 , n3000 , n3001 , n3002 , n3003 , n3004 , n3005 , n3006 , n3007 , n3008 , n3009 , n3010 , n3011 , n3012 , n3013 , n3014 , n3015 , n3016 , n3017 , n3018 , n3019 , n3020 , n3021 , n3022 , n3023 , n3024 , n3025 , n3026 , n3027 , n3028 , n3029 , n3030 , n3031 , n3032 , n3033 , n3034 , n3035 , n3036 , n3037 , n3038 , n3039 , n3040 , n3041 , n3042 , n3043 , n3044 , n3045 , n3046 , n3047 , n3048 , n3049 , n3050 , n3051 , n3052 , n3053 , n3054 , n3055 , n3056 , n3057 , n3058 , n3059 , n3060 , n3061 , n3062 , n3063 , n3064 , n3065 , n3066 , n3067 , n3068 , n3069 , n3070 , n3071 , n3072 , n3073 , n3074 , n3075 , n3076 , n3077 , n3078 , n3079 , n3080 , n3081 , n3082 , n3083 , n3084 , n3085 , n3086 , n3087 , n3088 , n3089 , n3090 , n3091 , n3092 , n3093 , n3094 , n3095 , n3096 , n3097 , n3098 , n3099 , n3100 , n3101 , n3102 , n3103 , n3104 , n3105 , n3106 , n3107 , n3108 , n3109 , n3110 , n3111 , n3112 , n3113 , n3114 , n3115 , n3116 , n3117 , n3118 , n3119 , n3120 , n3121 , n3122 , n3123 , n3124 , n3125 , n3126 , n3127 , n3128 , n3129 , n3130 , n3131 , n3132 , n3133 , n3134 , n3135 , n3136 , n3137 , n3138 , n3139 , n3140 , n3141 , n3142 , n3143 , n3144 , n3145 , n3146 , n3147 , n3148 , n3149 , n3150 , n3151 , n3152 , n3153 , n3154 , n3155 , n3156 , n3157 , n3158 , n3159 , n3160 , n3161 , n3162 , n3163 , n3164 , n3165 , n3166 , n3167 , n3168 , n3169 , n3170 , n3171 , n3172 , n3173 , n3174 , n3175 , n3176 , n3177 , n3178 , n3179 , n3180 , n3181 , n3182 , n3183 , n3184 , n3185 , n3186 , n3187 , n3188 , n3189 , n3190 , n3191 , n3192 , n3193 , n3194 , n3195 , n3196 , n3197 , n3198 , n3199 , n3200 , n3201 , n3202 , n3203 , n3204 , n3205 , n3206 , n3207 , n3208 , n3209 , n3210 , n3211 , n3212 , n3213 , n3214 , n3215 , n3216 , n3217 , n3218 , n3219 , n3220 , n3221 , n3222 , n3223 , n3224 , n3225 , n3226 , n3227 , n3228 , n3229 , n3230 , n3231 , n3232 , n3233 , n3234 , n3235 , n3236 , n3237 , n3238 , n3239 , n3240 , n3241 , n3242 , n3243 , n3244 , n3245 , n3246 , n3247 , n3248 , n3249 , n3250 , n3251 , n3252 , n3253 , n3254 , n3255 , n3256 , n3257 , n3258 , n3259 , n3260 , n3261 , n3262 , n3263 , n3264 , n3265 , n3266 , n3267 , n3268 , n3269 , n3270 , n3271 , n3272 , n3273 , n3274 , n3275 , n3276 , n3277 , n3278 , n3279 , n3280 , n3281 , n3282 , n3283 , n3284 , n3285 , n3286 , n3287 , n3288 , n3289 , n3290 , n3291 , n3292 , n3293 , n3294 , n3295 , n3296 , n3297 , n3298 , n3299 , n3300 , n3301 , n3302 , n3303 , n3304 , n3305 , n3306 , n3307 , n3308 , n3309 , n3310 , n3311 , n3312 , n3313 , n3314 , n3315 , n3316 , n3317 , n3318 , n3319 , n3320 , n3321 , n3322 , n3323 , n3324 , n3325 , n3326 , n3327 , n3328 , n3329 , n3330 , n3331 , n3332 , n3333 , n3334 , n3335 , n3336 , n3337 , n3338 , n3339 , n3340 , n3341 , n3342 , n3343 , n3344 , n3345 , n3346 , n3347 , n3348 , n3349 , n3350 , n3351 , n3352 , n3353 , n3354 , n3355 , n3356 , n3357 , n3358 , n3359 , n3360 , n3361 , n3362 , n3363 , n3364 , n3365 , n3366 , n3367 , n3368 , n3369 , n3370 , n3371 , n3372 , n3373 , n3374 , n3375 , n3376 , n3377 , n3378 , n3379 , n3380 , n3381 , n3382 , n3383 , n3384 , n3385 , n3386 , n3387 , n3388 , n3389 , n3390 , n3391 , n3392 , n3393 , n3394 , n3395 , n3396 , n3397 , n3398 , n3399 , n3400 , n3401 , n3402 , n3403 , n3404 , n3405 , n3406 , n3407 , n3408 , n3409 , n3410 , n3411 , n3412 , n3413 , n3414 , n3415 , n3416 , n3417 , n3418 , n3419 , n3420 , n3421 , n3422 , n3423 , n3424 , n3425 , n3426 , n3427 , n3428 , n3429 , n3430 , n3431 , n3432 , n3433 , n3434 , n3435 , n3436 , n3437 , n3438 , n3439 , n3440 , n3441 , n3442 , n3443 , n3444 , n3445 , n3446 , n3447 , n3448 , n3449 , n3450 , n3451 , n3452 , n3453 , n3454 , n3455 , n3456 , n3457 , n3458 , n3459 , n3460 , n3461 , n3462 , n3463 , n3464 , n3465 , n3466 , n3467 , n3468 , n3469 , n3470 , n3471 , n3472 , n3473 , n3474 , n3475 , n3476 , n3477 , n3478 , n3479 , n3480 , n3481 , n3482 , n3483 , n3484 , n3485 , n3486 , n3487 , n3488 , n3489 , n3490 , n3491 , n3492 , n3493 , n3494 , n3495 , n3496 , n3497 , n3498 , n3499 , n3500 , n3501 , n3502 , n3503 , n3504 , n3505 , n3506 , n3507 , n3508 , n3509 , n3510 , n3511 , n3512 , n3513 , n3514 , n3515 , n3516 , n3517 , n3518 , n3519 , n3520 , n3521 , n3522 , n3523 , n3524 , n3525 , n3526 , n3527 , n3528 , n3529 , n3530 , n3531 , n3532 , n3533 , n3534 , n3535 , n3536 , n3537 , n3538 , n3539 , n3540 , n3541 , n3542 , n3543 , n3544 , n3545 , n3546 , n3547 , n3548 , n3549 , n3550 , n3551 , n3552 , n3553 , n3554 , n3555 , n3556 , n3557 , n3558 , n3559 , n3560 , n3561 , n3562 , n3563 , n3564 , n3565 , n3566 , n3567 , n3568 , n3569 , n3570 , n3571 , n3572 , n3573 , n3574 , n3575 , n3576 , n3577 , n3578 , n3579 , n3580 , n3581 , n3582 , n3583 , n3584 , n3585 , n3586 , n3587 , n3588 , n3589 , n3590 , n3591 , n3592 , n3593 , n3594 , n3595 , n3596 , n3597 , n3598 , n3599 , n3600 , n3601 , n3602 , n3603 , n3604 , n3605 , n3606 , n3607 , n3608 , n3609 , n3610 , n3611 , n3612 , n3613 , n3614 , n3615 , n3616 , n3617 , n3618 , n3619 , n3620 , n3621 , n3622 , n3623 , n3624 , n3625 , n3626 , n3627 , n3628 , n3629 , n3630 , n3631 , n3632 , n3633 , n3634 , n3635 , n3636 , n3637 , n3638 , n3639 , n3640 , n3641 , n3642 , n3643 , n3644 , n3645 , n3646 , n3647 , n3648 , n3649 , n3650 , n3651 , n3652 , n3653 , n3654 , n3655 , n3656 , n3657 , n3658 , n3659 , n3660 , n3661 , n3662 , n3663 , n3664 , n3665 , n3666 , n3667 , n3668 , n3669 , n3670 , n3671 , n3672 , n3673 , n3674 , n3675 , n3676 , n3677 , n3678 , n3679 , n3680 , n3681 , n3682 , n3683 , n3684 , n3685 , n3686 , n3687 , n3688 , n3689 , n3690 , n3691 , n3692 , n3693 , n3694 , n3695 , n3696 , n3697 , n3698 , n3699 , n3700 , n3701 , n3702 , n3703 , n3704 , n3705 , n3706 , n3707 , n3708 , n3709 , n3710 , n3711 , n3712 , n3713 , n3714 , n3715 , n3716 , n3717 , n3718 , n3719 , n3720 , n3721 , n3722 , n3723 , n3724 , n3725 , n3726 , n3727 , n3728 , n3729 , n3730 , n3731 , n3732 , n3733 , n3734 , n3735 , n3736 , n3737 , n3738 , n3739 , n3740 , n3741 , n3742 , n3743 , n3744 , n3745 , n3746 , n3747 , n3748 , n3749 , n3750 , n3751 , n3752 , n3753 , n3754 , n3755 , n3756 , n3757 , n3758 , n3759 , n3760 , n3761 , n3762 , n3763 , n3764 , n3765 , n3766 , n3767 , n3768 , n3769 , n3770 , n3771 , n3772 , n3773 , n3774 , n3775 , n3776 , n3777 , n3778 , n3779 , n3780 , n3781 , n3782 , n3783 , n3784 , n3785 , n3786 , n3787 , n3788 , n3789 , n3790 , n3791 , n3792 , n3793 , n3794 , n3795 , n3796 , n3797 , n3798 , n3799 , n3800 , n3801 , n3802 , n3803 , n3804 , n3805 , n3806 , n3807 , n3808 , n3809 , n3810 , n3811 , n3812 , n3813 , n3814 , n3815 , n3816 , n3817 , n3818 , n3819 , n3820 , n3821 , n3822 , n3823 , n3824 , n3825 , n3826 , n3827 , n3828 , n3829 , n3830 , n3831 , n3832 , n3833 , n3834 , n3835 , n3836 , n3837 , n3838 , n3839 , n3840 , n3841 , n3842 , n3843 , n3844 , n3845 , n3846 , n3847 , n3848 , n3849 , n3850 , n3851 , n3852 , n3853 , n3854 , n3855 , n3856 , n3857 , n3858 , n3859 , n3860 , n3861 , n3862 , n3863 , n3864 , n3865 , n3866 , n3867 , n3868 , n3869 , n3870 , n3871 , n3872 , n3873 , n3874 , n3875 , n3876 , n3877 , n3878 , n3879 , n3880 , n3881 , n3882 , n3883 , n3884 , n3885 , n3886 , n3887 , n3888 , n3889 , n3890 , n3891 , n3892 , n3893 , n3894 , n3895 , n3896 , n3897 , n3898 , n3899 , n3900 , n3901 , n3902 , n3903 , n3904 , n3905 , n3906 , n3907 , n3908 , n3909 , n3910 , n3911 , n3912 , n3913 , n3914 , n3915 , n3916 , n3917 , n3918 , n3919 , n3920 , n3921 , n3922 , n3923 , n3924 , n3925 , n3926 , n3927 , n3928 , n3929 , n3930 , n3931 , n3932 , n3933 , n3934 , n3935 , n3936 , n3937 , n3938 , n3939 , n3940 , n3941 , n3942 , n3943 , n3944 , n3945 , n3946 , n3947 , n3948 , n3949 , n3950 , n3951 , n3952 , n3953 , n3954 , n3955 , n3956 , n3957 , n3958 , n3959 , n3960 , n3961 , n3962 , n3963 , n3964 , n3965 , n3966 , n3967 , n3968 , n3969 , n3970 , n3971 , n3972 , n3973 , n3974 , n3975 , n3976 , n3977 , n3978 , n3979 , n3980 , n3981 , n3982 , n3983 , n3984 , n3985 , n3986 , n3987 , n3988 , n3989 , n3990 , n3991 , n3992 , n3993 , n3994 , n3995 , n3996 , n3997 , n3998 , n3999 , n4000 , n4001 , n4002 , n4003 , n4004 , n4005 , n4006 , n4007 , n4008 , n4009 , n4010 , n4011 , n4012 , n4013 , n4014 , n4015 , n4016 , n4017 , n4018 , n4019 , n4020 , n4021 , n4022 , n4023 , n4024 , n4025 , n4026 , n4027 , n4028 , n4029 , n4030 , n4031 , n4032 , n4033 , n4034 , n4035 , n4036 , n4037 , n4038 , n4039 , n4040 , n4041 , n4042 , n4043 , n4044 , n4045 , n4046 , n4047 , n4048 , n4049 , n4050 , n4051 , n4052 , n4053 , n4054 , n4055 , n4056 , n4057 , n4058 , n4059 , n4060 , n4061 , n4062 , n4063 , n4064 , n4065 , n4066 , n4067 , n4068 , n4069 , n4070 , n4071 , n4072 , n4073 , n4074 , n4075 , n4076 , n4077 , n4078 , n4079 , n4080 , n4081 , n4082 , n4083 , n4084 , n4085 , n4086 , n4087 , n4088 , n4089 , n4090 , n4091 , n4092 , n4093 , n4094 , n4095 , n4096 , n4097 , n4098 , n4099 , n4100 , n4101 , n4102 , n4103 , n4104 , n4105 , n4106 , n4107 , n4108 , n4109 , n4110 , n4111 , n4112 , n4113 , n4114 , n4115 , n4116 , n4117 , n4118 , n4119 , n4120 , n4121 , n4122 , n4123 , n4124 , n4125 , n4126 , n4127 , n4128 , n4129 , n4130 , n4131 , n4132 , n4133 , n4134 , n4135 , n4136 , n4137 , n4138 , n4139 , n4140 , n4141 , n4142 , n4143 , n4144 , n4145 , n4146 , n4147 , n4148 , n4149 , n4150 , n4151 , n4152 , n4153 , n4154 , n4155 , n4156 , n4157 , n4158 , n4159 , n4160 , n4161 , n4162 , n4163 , n4164 , n4165 , n4166 , n4167 , n4168 , n4169 , n4170 , n4171 , n4172 , n4173 , n4174 , n4175 , n4176 , n4177 , n4178 , n4179 , n4180 , n4181 , n4182 , n4183 , n4184 , n4185 , n4186 , n4187 , n4188 , n4189 , n4190 , n4191 , n4192 , n4193 , n4194 , n4195 , n4196 , n4197 , n4198 , n4199 , n4200 , n4201 , n4202 , n4203 , n4204 , n4205 , n4206 , n4207 , n4208 , n4209 , n4210 , n4211 , n4212 , n4213 , n4214 , n4215 , n4216 , n4217 , n4218 , n4219 , n4220 , n4221 , n4222 , n4223 , n4224 , n4225 , n4226 , n4227 , n4228 , n4229 , n4230 , n4231 , n4232 , n4233 , n4234 , n4235 , n4236 , n4237 , n4238 , n4239 , n4240 , n4241 , n4242 , n4243 , n4244 , n4245 , n4246 , n4247 , n4248 , n4249 , n4250 , n4251 , n4252 , n4253 , n4254 , n4255 , n4256 , n4257 , n4258 , n4259 , n4260 , n4261 , n4262 , n4263 , n4264 , n4265 , n4266 , n4267 , n4268 , n4269 , n4270 , n4271 , n4272 , n4273 , n4274 , n4275 , n4276 , n4277 , n4278 , n4279 , n4280 , n4281 , n4282 , n4283 , n4284 , n4285 , n4286 , n4287 , n4288 , n4289 , n4290 , n4291 , n4292 , n4293 , n4294 , n4295 , n4296 , n4297 , n4298 , n4299 , n4300 , n4301 , n4302 , n4303 , n4304 , n4305 , n4306 , n4307 , n4308 , n4309 , n4310 , n4311 , n4312 , n4313 , n4314 , n4315 , n4316 , n4317 , n4318 , n4319 , n4320 , n4321 , n4322 , n4323 , n4324 , n4325 , n4326 , n4327 , n4328 , n4329 , n4330 , n4331 , n4332 , n4333 , n4334 , n4335 , n4336 , n4337 , n4338 , n4339 , n4340 , n4341 , n4342 , n4343 , n4344 , n4345 , n4346 , n4347 , n4348 , n4349 , n4350 , n4351 , n4352 , n4353 , n4354 , n4355 , n4356 , n4357 , n4358 , n4359 , n4360 , n4361 , n4362 , n4363 , n4364 , n4365 , n4366 , n4367 , n4368 , n4369 , n4370 , n4371 , n4372 , n4373 , n4374 , n4375 , n4376 , n4377 , n4378 , n4379 , n4380 , n4381 , n4382 , n4383 , n4384 , n4385 , n4386 , n4387 , n4388 , n4389 , n4390 , n4391 , n4392 , n4393 , n4394 , n4395 , n4396 , n4397 , n4398 , n4399 , n4400 , n4401 , n4402 , n4403 , n4404 , n4405 , n4406 , n4407 , n4408 , n4409 , n4410 , n4411 , n4412 , n4413 , n4414 , n4415 , n4416 , n4417 , n4418 , n4419 , n4420 , n4421 , n4422 , n4423 , n4424 , n4425 , n4426 , n4427 , n4428 , n4429 , n4430 , n4431 , n4432 , n4433 , n4434 , n4435 , n4436 , n4437 , n4438 , n4439 , n4440 , n4441 , n4442 , n4443 , n4444 , n4445 , n4446 , n4447 , n4448 , n4449 , n4450 , n4451 , n4452 , n4453 , n4454 , n4455 , n4456 , n4457 , n4458 , n4459 , n4460 , n4461 , n4462 , n4463 , n4464 , n4465 , n4466 , n4467 , n4468 , n4469 , n4470 , n4471 , n4472 , n4473 , n4474 , n4475 , n4476 , n4477 , n4478 , n4479 , n4480 , n4481 , n4482 , n4483 , n4484 , n4485 , n4486 , n4487 , n4488 , n4489 , n4490 , n4491 , n4492 , n4493 , n4494 , n4495 , n4496 , n4497 , n4498 , n4499 , n4500 , n4501 , n4502 , n4503 , n4504 , n4505 , n4506 , n4507 , n4508 , n4509 , n4510 , n4511 , n4512 , n4513 , n4514 , n4515 , n4516 , n4517 , n4518 , n4519 , n4520 , n4521 , n4522 , n4523 , n4524 , n4525 , n4526 , n4527 , n4528 , n4529 , n4530 , n4531 , n4532 , n4533 , n4534 , n4535 , n4536 , n4537 , n4538 , n4539 , n4540 , n4541 , n4542 , n4543 , n4544 , n4545 , n4546 , n4547 , n4548 , n4549 , n4550 , n4551 , n4552 , n4553 , n4554 , n4555 , n4556 , n4557 , n4558 , n4559 , n4560 , n4561 , n4562 , n4563 , n4564 , n4565 , n4566 , n4567 , n4568 , n4569 , n4570 , n4571 , n4572 , n4573 , n4574 , n4575 , n4576 , n4577 , n4578 , n4579 , n4580 , n4581 , n4582 , n4583 , n4584 , n4585 , n4586 , n4587 , n4588 , n4589 , n4590 , n4591 , n4592 , n4593 , n4594 , n4595 , n4596 , n4597 , n4598 , n4599 , n4600 , n4601 , n4602 , n4603 , n4604 , n4605 , n4606 , n4607 , n4608 , n4609 , n4610 , n4611 , n4612 , n4613 , n4614 , n4615 , n4616 , n4617 , n4618 , n4619 , n4620 , n4621 , n4622 , n4623 , n4624 , n4625 , n4626 , n4627 , n4628 , n4629 , n4630 , n4631 , n4632 , n4633 , n4634 , n4635 , n4636 , n4637 , n4638 , n4639 , n4640 , n4641 , n4642 , n4643 , n4644 , n4645 , n4646 , n4647 , n4648 , n4649 , n4650 , n4651 , n4652 , n4653 , n4654 , n4655 , n4656 , n4657 , n4658 , n4659 , n4660 , n4661 , n4662 , n4663 , n4664 , n4665 , n4666 , n4667 , n4668 , n4669 , n4670 , n4671 , n4672 , n4673 , n4674 , n4675 , n4676 , n4677 , n4678 , n4679 , n4680 , n4681 , n4682 , n4683 , n4684 , n4685 , n4686 , n4687 , n4688 , n4689 , n4690 , n4691 , n4692 , n4693 , n4694 , n4695 , n4696 , n4697 , n4698 , n4699 , n4700 , n4701 , n4702 , n4703 , n4704 , n4705 , n4706 , n4707 , n4708 , n4709 , n4710 , n4711 , n4712 , n4713 , n4714 , n4715 , n4716 , n4717 , n4718 , n4719 , n4720 , n4721 , n4722 , n4723 , n4724 , n4725 , n4726 , n4727 , n4728 , n4729 , n4730 , n4731 , n4732 , n4733 , n4734 , n4735 , n4736 , n4737 , n4738 , n4739 , n4740 , n4741 , n4742 , n4743 , n4744 , n4745 , n4746 , n4747 , n4748 , n4749 , n4750 , n4751 , n4752 , n4753 , n4754 , n4755 , n4756 , n4757 , n4758 , n4759 , n4760 , n4761 , n4762 , n4763 , n4764 , n4765 , n4766 , n4767 , n4768 , n4769 , n4770 , n4771 , n4772 , n4773 , n4774 , n4775 , n4776 , n4777 , n4778 , n4779 , n4780 , n4781 , n4782 , n4783 , n4784 , n4785 , n4786 , n4787 , n4788 , n4789 , n4790 , n4791 , n4792 , n4793 , n4794 , n4795 , n4796 , n4797 , n4798 , n4799 , n4800 , n4801 , n4802 , n4803 , n4804 , n4805 , n4806 , n4807 , n4808 , n4809 , n4810 , n4811 , n4812 , n4813 , n4814 , n4815 , n4816 , n4817 , n4818 , n4819 , n4820 , n4821 , n4822 , n4823 , n4824 , n4825 , n4826 , n4827 , n4828 , n4829 , n4830 , n4831 , n4832 , n4833 , n4834 , n4835 , n4836 , n4837 , n4838 , n4839 , n4840 , n4841 , n4842 , n4843 , n4844 , n4845 , n4846 , n4847 , n4848 , n4849 , n4850 , n4851 , n4852 , n4853 , n4854 , n4855 , n4856 , n4857 , n4858 , n4859 , n4860 , n4861 , n4862 , n4863 , n4864 , n4865 , n4866 , n4867 , n4868 , n4869 , n4870 , n4871 , n4872 , n4873 , n4874 , n4875 , n4876 , n4877 , n4878 , n4879 , n4880 , n4881 , n4882 , n4883 , n4884 , n4885 , n4886 , n4887 , n4888 , n4889 , n4890 , n4891 , n4892 , n4893 , n4894 , n4895 , n4896 , n4897 , n4898 , n4899 , n4900 , n4901 , n4902 , n4903 , n4904 , n4905 , n4906 , n4907 , n4908 , n4909 , n4910 , n4911 , n4912 , n4913 , n4914 , n4915 , n4916 , n4917 , n4918 , n4919 , n4920 , n4921 , n4922 , n4923 , n4924 , n4925 , n4926 , n4927 , n4928 , n4929 , n4930 , n4931 , n4932 , n4933 , n4934 , n4935 , n4936 , n4937 , n4938 , n4939 , n4940 , n4941 , n4942 , n4943 , n4944 , n4945 , n4946 , n4947 , n4948 , n4949 , n4950 , n4951 , n4952 , n4953 , n4954 , n4955 , n4956 , n4957 , n4958 , n4959 , n4960 , n4961 , n4962 , n4963 , n4964 , n4965 , n4966 , n4967 , n4968 , n4969 , n4970 , n4971 , n4972 , n4973 , n4974 , n4975 , n4976 , n4977 , n4978 , n4979 , n4980 , n4981 , n4982 , n4983 , n4984 , n4985 , n4986 , n4987 , n4988 , n4989 , n4990 , n4991 , n4992 , n4993 , n4994 , n4995 , n4996 , n4997 , n4998 , n4999 , n5000 , n5001 , n5002 , n5003 , n5004 , n5005 , n5006 , n5007 , n5008 , n5009 , n5010 , n5011 , n5012 , n5013 , n5014 , n5015 , n5016 , n5017 , n5018 , n5019 , n5020 , n5021 , n5022 , n5023 , n5024 , n5025 , n5026 , n5027 , n5028 , n5029 , n5030 , n5031 , n5032 , n5033 , n5034 , n5035 , n5036 , n5037 , n5038 , n5039 , n5040 , n5041 , n5042 , n5043 , n5044 , n5045 , n5046 , n5047 , n5048 , n5049 , n5050 , n5051 , n5052 , n5053 , n5054 , n5055 , n5056 , n5057 , n5058 , n5059 , n5060 , n5061 , n5062 , n5063 , n5064 , n5065 , n5066 , n5067 , n5068 , n5069 , n5070 , n5071 , n5072 , n5073 , n5074 , n5075 , n5076 , n5077 , n5078 , n5079 , n5080 , n5081 , n5082 , n5083 , n5084 , n5085 , n5086 , n5087 , n5088 , n5089 , n5090 , n5091 , n5092 , n5093 , n5094 , n5095 , n5096 , n5097 , n5098 , n5099 , n5100 , n5101 , n5102 , n5103 , n5104 , n5105 , n5106 , n5107 , n5108 , n5109 , n5110 , n5111 , n5112 , n5113 , n5114 , n5115 , n5116 , n5117 , n5118 , n5119 , n5120 , n5121 , n5122 , n5123 , n5124 , n5125 , n5126 , n5127 , n5128 , n5129 , n5130 , n5131 , n5132 , n5133 , n5134 , n5135 , n5136 , n5137 , n5138 , n5139 , n5140 , n5141 , n5142 , n5143 , n5144 , n5145 , n5146 , n5147 , n5148 , n5149 , n5150 , n5151 , n5152 , n5153 , n5154 , n5155 , n5156 , n5157 , n5158 , n5159 , n5160 , n5161 , n5162 , n5163 , n5164 , n5165 , n5166 , n5167 , n5168 , n5169 , n5170 , n5171 , n5172 , n5173 , n5174 , n5175 , n5176 , n5177 , n5178 , n5179 , n5180 , n5181 , n5182 , n5183 , n5184 , n5185 , n5186 , n5187 , n5188 , n5189 , n5190 , n5191 , n5192 , n5193 , n5194 , n5195 , n5196 , n5197 , n5198 , n5199 , n5200 , n5201 , n5202 , n5203 , n5204 , n5205 , n5206 , n5207 , n5208 , n5209 , n5210 , n5211 , n5212 , n5213 , n5214 , n5215 , n5216 , n5217 , n5218 , n5219 , n5220 , n5221 , n5222 , n5223 , n5224 , n5225 , n5226 , n5227 , n5228 , n5229 , n5230 , n5231 , n5232 , n5233 , n5234 , n5235 , n5236 , n5237 , n5238 , n5239 , n5240 , n5241 , n5242 , n5243 , n5244 , n5245 , n5246 , n5247 , n5248 , n5249 , n5250 , n5251 , n5252 , n5253 , n5254 , n5255 , n5256 , n5257 , n5258 , n5259 , n5260 , n5261 , n5262 , n5263 , n5264 , n5265 , n5266 , n5267 , n5268 , n5269 , n5270 , n5271 , n5272 , n5273 , n5274 , n5275 , n5276 , n5277 , n5278 , n5279 , n5280 , n5281 , n5282 , n5283 , n5284 , n5285 , n5286 , n5287 , n5288 , n5289 , n5290 , n5291 , n5292 , n5293 , n5294 , n5295 , n5296 , n5297 , n5298 , n5299 , n5300 , n5301 , n5302 , n5303 , n5304 , n5305 , n5306 , n5307 , n5308 , n5309 , n5310 , n5311 , n5312 , n5313 , n5314 , n5315 , n5316 , n5317 , n5318 , n5319 , n5320 , n5321 , n5322 , n5323 , n5324 , n5325 , n5326 , n5327 , n5328 , n5329 , n5330 , n5331 , n5332 , n5333 , n5334 , n5335 , n5336 , n5337 , n5338 , n5339 , n5340 , n5341 , n5342 , n5343 , n5344 , n5345 , n5346 , n5347 , n5348 , n5349 , n5350 , n5351 , n5352 , n5353 , n5354 , n5355 , n5356 , n5357 , n5358 , n5359 , n5360 , n5361 , n5362 , n5363 , n5364 , n5365 , n5366 , n5367 , n5368 , n5369 , n5370 , n5371 , n5372 , n5373 , n5374 , n5375 , n5376 , n5377 , n5378 , n5379 , n5380 , n5381 , n5382 , n5383 , n5384 , n5385 , n5386 , n5387 , n5388 , n5389 , n5390 , n5391 , n5392 , n5393 , n5394 , n5395 , n5396 , n5397 , n5398 , n5399 , n5400 , n5401 , n5402 , n5403 , n5404 , n5405 , n5406 , n5407 , n5408 , n5409 , n5410 , n5411 , n5412 , n5413 , n5414 , n5415 , n5416 , n5417 , n5418 , n5419 , n5420 , n5421 , n5422 , n5423 , n5424 , n5425 , n5426 , n5427 , n5428 , n5429 , n5430 , n5431 , n5432 , n5433 , n5434 , n5435 , n5436 , n5437 , n5438 , n5439 , n5440 , n5441 , n5442 , n5443 , n5444 , n5445 , n5446 , n5447 , n5448 , n5449 , n5450 , n5451 , n5452 , n5453 , n5454 , n5455 , n5456 , n5457 , n5458 , n5459 , n5460 , n5461 , n5462 , n5463 , n5464 , n5465 , n5466 , n5467 , n5468 , n5469 , n5470 , n5471 , n5472 , n5473 , n5474 , n5475 , n5476 , n5477 , n5478 , n5479 , n5480 , n5481 , n5482 , n5483 , n5484 , n5485 , n5486 , n5487 , n5488 , n5489 , n5490 , n5491 , n5492 , n5493 , n5494 , n5495 , n5496 , n5497 , n5498 , n5499 , n5500 , n5501 , n5502 , n5503 , n5504 , n5505 , n5506 , n5507 , n5508 , n5509 , n5510 , n5511 , n5512 , n5513 , n5514 , n5515 , n5516 , n5517 , n5518 , n5519 , n5520 , n5521 , n5522 , n5523 , n5524 , n5525 , n5526 , n5527 , n5528 , n5529 , n5530 , n5531 , n5532 , n5533 , n5534 , n5535 , n5536 , n5537 , n5538 , n5539 , n5540 , n5541 , n5542 , n5543 , n5544 , n5545 , n5546 , n5547 , n5548 , n5549 , n5550 , n5551 , n5552 , n5553 , n5554 , n5555 , n5556 , n5557 , n5558 , n5559 , n5560 , n5561 , n5562 , n5563 , n5564 , n5565 , n5566 , n5567 , n5568 , n5569 , n5570 , n5571 , n5572 , n5573 , n5574 , n5575 , n5576 , n5577 , n5578 , n5579 , n5580 , n5581 , n5582 , n5583 , n5584 , n5585 , n5586 , n5587 , n5588 , n5589 , n5590 , n5591 , n5592 , n5593 , n5594 , n5595 , n5596 , n5597 , n5598 , n5599 , n5600 , n5601 , n5602 , n5603 , n5604 , n5605 , n5606 , n5607 , n5608 , n5609 , n5610 , n5611 , n5612 , n5613 , n5614 , n5615 , n5616 , n5617 , n5618 , n5619 , n5620 , n5621 , n5622 , n5623 , n5624 , n5625 , n5626 , n5627 , n5628 , n5629 , n5630 , n5631 , n5632 , n5633 , n5634 , n5635 , n5636 , n5637 , n5638 , n5639 , n5640 , n5641 , n5642 , n5643 , n5644 , n5645 , n5646 , n5647 , n5648 , n5649 , n5650 , n5651 , n5652 , n5653 , n5654 , n5655 , n5656 , n5657 , n5658 , n5659 , n5660 , n5661 , n5662 , n5663 , n5664 , n5665 , n5666 , n5667 , n5668 , n5669 , n5670 , n5671 , n5672 , n5673 , n5674 , n5675 , n5676 , n5677 , n5678 , n5679 , n5680 , n5681 , n5682 , n5683 , n5684 , n5685 , n5686 , n5687 , n5688 , n5689 , n5690 , n5691 , n5692 , n5693 , n5694 , n5695 , n5696 , n5697 , n5698 , n5699 , n5700 , n5701 , n5702 , n5703 , n5704 , n5705 , n5706 , n5707 , n5708 , n5709 , n5710 , n5711 , n5712 , n5713 , n5714 , n5715 , n5716 , n5717 , n5718 , n5719 , n5720 , n5721 , n5722 , n5723 , n5724 , n5725 , n5726 , n5727 , n5728 , n5729 , n5730 , n5731 , n5732 , n5733 , n5734 , n5735 , n5736 , n5737 , n5738 , n5739 , n5740 , n5741 , n5742 , n5743 , n5744 , n5745 , n5746 , n5747 , n5748 , n5749 , n5750 , n5751 , n5752 , n5753 , n5754 , n5755 , n5756 , n5757 , n5758 , n5759 , n5760 , n5761 , n5762 , n5763 , n5764 , n5765 , n5766 , n5767 , n5768 , n5769 , n5770 , n5771 , n5772 , n5773 , n5774 , n5775 , n5776 , n5777 , n5778 , n5779 , n5780 , n5781 , n5782 , n5783 , n5784 , n5785 , n5786 , n5787 , n5788 , n5789 , n5790 , n5791 , n5792 , n5793 , n5794 , n5795 , n5796 , n5797 , n5798 , n5799 , n5800 , n5801 , n5802 , n5803 , n5804 , n5805 , n5806 , n5807 , n5808 , n5809 , n5810 , n5811 , n5812 , n5813 , n5814 , n5815 , n5816 , n5817 , n5818 , n5819 , n5820 , n5821 , n5822 , n5823 , n5824 , n5825 , n5826 , n5827 , n5828 , n5829 , n5830 , n5831 , n5832 , n5833 , n5834 , n5835 , n5836 , n5837 , n5838 , n5839 , n5840 , n5841 , n5842 , n5843 , n5844 , n5845 , n5846 , n5847 , n5848 , n5849 , n5850 , n5851 , n5852 , n5853 , n5854 , n5855 , n5856 , n5857 , n5858 , n5859 , n5860 , n5861 , n5862 , n5863 , n5864 , n5865 , n5866 , n5867 , n5868 , n5869 , n5870 , n5871 , n5872 , n5873 , n5874 , n5875 , n5876 , n5877 , n5878 , n5879 , n5880 , n5881 , n5882 , n5883 , n5884 , n5885 , n5886 , n5887 , n5888 , n5889 , n5890 , n5891 , n5892 , n5893 , n5894 , n5895 , n5896 , n5897 , n5898 , n5899 , n5900 , n5901 , n5902 , n5903 , n5904 , n5905 , n5906 , n5907 , n5908 , n5909 , n5910 , n5911 , n5912 , n5913 , n5914 , n5915 , n5916 , n5917 , n5918 , n5919 , n5920 , n5921 , n5922 , n5923 , n5924 , n5925 , n5926 , n5927 , n5928 , n5929 , n5930 , n5931 , n5932 , n5933 , n5934 , n5935 , n5936 , n5937 , n5938 , n5939 , n5940 , n5941 , n5942 , n5943 , n5944 , n5945 , n5946 , n5947 , n5948 , n5949 , n5950 , n5951 , n5952 , n5953 , n5954 , n5955 , n5956 , n5957 , n5958 , n5959 , n5960 , n5961 , n5962 , n5963 , n5964 , n5965 , n5966 , n5967 , n5968 , n5969 , n5970 , n5971 , n5972 , n5973 , n5974 , n5975 , n5976 , n5977 , n5978 , n5979 , n5980 , n5981 , n5982 , n5983 , n5984 , n5985 , n5986 , n5987 , n5988 , n5989 , n5990 , n5991 , n5992 , n5993 , n5994 , n5995 , n5996 , n5997 , n5998 , n5999 , n6000 , n6001 , n6002 , n6003 , n6004 , n6005 , n6006 , n6007 , n6008 , n6009 , n6010 , n6011 , n6012 , n6013 , n6014 , n6015 , n6016 , n6017 , n6018 , n6019 , n6020 , n6021 , n6022 , n6023 , n6024 , n6025 , n6026 , n6027 , n6028 , n6029 , n6030 , n6031 , n6032 , n6033 , n6034 , n6035 , n6036 , n6037 , n6038 , n6039 , n6040 , n6041 , n6042 , n6043 , n6044 , n6045 , n6046 , n6047 , n6048 , n6049 , n6050 , n6051 , n6052 , n6053 , n6054 , n6055 , n6056 , n6057 , n6058 , n6059 , n6060 , n6061 , n6062 , n6063 , n6064 , n6065 , n6066 , n6067 , n6068 , n6069 , n6070 , n6071 , n6072 , n6073 , n6074 , n6075 , n6076 , n6077 , n6078 , n6079 , n6080 , n6081 , n6082 , n6083 , n6084 , n6085 , n6086 , n6087 , n6088 , n6089 , n6090 , n6091 , n6092 , n6093 , n6094 , n6095 , n6096 , n6097 , n6098 , n6099 , n6100 , n6101 , n6102 , n6103 , n6104 , n6105 , n6106 , n6107 , n6108 , n6109 , n6110 , n6111 , n6112 , n6113 , n6114 , n6115 , n6116 , n6117 , n6118 , n6119 , n6120 , n6121 , n6122 , n6123 , n6124 , n6125 , n6126 , n6127 , n6128 , n6129 , n6130 , n6131 , n6132 , n6133 , n6134 , n6135 , n6136 , n6137 , n6138 , n6139 , n6140 , n6141 , n6142 , n6143 , n6144 , n6145 , n6146 , n6147 , n6148 , n6149 , n6150 , n6151 , n6152 , n6153 , n6154 , n6155 , n6156 , n6157 , n6158 , n6159 , n6160 , n6161 , n6162 , n6163 , n6164 , n6165 , n6166 , n6167 , n6168 , n6169 , n6170 , n6171 , n6172 , n6173 , n6174 , n6175 , n6176 , n6177 , n6178 , n6179 , n6180 , n6181 , n6182 , n6183 , n6184 , n6185 , n6186 , n6187 , n6188 , n6189 , n6190 , n6191 , n6192 , n6193 , n6194 , n6195 , n6196 , n6197 , n6198 , n6199 , n6200 , n6201 , n6202 , n6203 , n6204 , n6205 , n6206 , n6207 , n6208 , n6209 , n6210 , n6211 , n6212 , n6213 , n6214 , n6215 , n6216 , n6217 , n6218 , n6219 , n6220 , n6221 , n6222 , n6223 , n6224 , n6225 , n6226 , n6227 , n6228 , n6229 , n6230 , n6231 , n6232 , n6233 , n6234 , n6235 , n6236 , n6237 , n6238 , n6239 , n6240 , n6241 , n6242 , n6243 , n6244 , n6245 , n6246 , n6247 , n6248 , n6249 , n6250 , n6251 , n6252 , n6253 , n6254 , n6255 , n6256 , n6257 , n6258 , n6259 , n6260 , n6261 , n6262 , n6263 , n6264 , n6265 , n6266 , n6267 , n6268 , n6269 , n6270 , n6271 , n6272 , n6273 , n6274 , n6275 , n6276 , n6277 , n6278 , n6279 , n6280 , n6281 , n6282 , n6283 , n6284 , n6285 , n6286 , n6287 , n6288 , n6289 , n6290 , n6291 , n6292 , n6293 , n6294 , n6295 , n6296 , n6297 , n6298 , n6299 , n6300 , n6301 , n6302 , n6303 , n6304 , n6305 , n6306 , n6307 , n6308 , n6309 , n6310 , n6311 , n6312 , n6313 , n6314 , n6315 , n6316 , n6317 , n6318 , n6319 , n6320 , n6321 , n6322 , n6323 , n6324 , n6325 , n6326 , n6327 , n6328 , n6329 , n6330 , n6331 , n6332 , n6333 , n6334 , n6335 , n6336 , n6337 , n6338 , n6339 , n6340 , n6341 , n6342 , n6343 , n6344 , n6345 , n6346 , n6347 , n6348 , n6349 , n6350 , n6351 , n6352 , n6353 , n6354 , n6355 , n6356 , n6357 , n6358 , n6359 , n6360 , n6361 , n6362 , n6363 , n6364 , n6365 , n6366 , n6367 , n6368 , n6369 , n6370 , n6371 , n6372 , n6373 , n6374 , n6375 , n6376 , n6377 , n6378 , n6379 , n6380 , n6381 , n6382 , n6383 , n6384 , n6385 , n6386 , n6387 , n6388 , n6389 , n6390 , n6391 , n6392 , n6393 , n6394 , n6395 , n6396 , n6397 , n6398 , n6399 , n6400 , n6401 , n6402 , n6403 , n6404 , n6405 , n6406 , n6407 , n6408 , n6409 , n6410 , n6411 , n6412 , n6413 , n6414 , n6415 , n6416 , n6417 , n6418 , n6419 , n6420 , n6421 , n6422 , n6423 , n6424 , n6425 , n6426 , n6427 , n6428 , n6429 , n6430 , n6431 , n6432 , n6433 , n6434 , n6435 , n6436 , n6437 , n6438 , n6439 , n6440 , n6441 , n6442 , n6443 , n6444 , n6445 , n6446 , n6447 , n6448 , n6449 , n6450 , n6451 , n6452 , n6453 , n6454 , n6455 , n6456 , n6457 , n6458 , n6459 , n6460 , n6461 , n6462 , n6463 , n6464 , n6465 , n6466 , n6467 , n6468 , n6469 , n6470 , n6471 , n6472 , n6473 , n6474 , n6475 , n6476 , n6477 , n6478 , n6479 , n6480 , n6481 , n6482 , n6483 , n6484 , n6485 , n6486 , n6487 , n6488 , n6489 , n6490 , n6491 , n6492 , n6493 , n6494 , n6495 , n6496 , n6497 , n6498 , n6499 , n6500 , n6501 , n6502 , n6503 , n6504 , n6505 , n6506 , n6507 , n6508 , n6509 , n6510 , n6511 , n6512 , n6513 , n6514 , n6515 , n6516 , n6517 , n6518 , n6519 , n6520 , n6521 , n6522 , n6523 , n6524 , n6525 , n6526 , n6527 , n6528 , n6529 , n6530 , n6531 , n6532 , n6533 , n6534 , n6535 , n6536 , n6537 , n6538 , n6539 , n6540 , n6541 , n6542 , n6543 , n6544 , n6545 , n6546 , n6547 , n6548 , n6549 , n6550 , n6551 , n6552 , n6553 , n6554 , n6555 , n6556 , n6557 , n6558 , n6559 , n6560 , n6561 , n6562 , n6563 , n6564 , n6565 , n6566 , n6567 , n6568 , n6569 , n6570 , n6571 , n6572 , n6573 , n6574 , n6575 , n6576 , n6577 , n6578 , n6579 , n6580 , n6581 , n6582 , n6583 , n6584 , n6585 , n6586 , n6587 , n6588 , n6589 , n6590 , n6591 , n6592 , n6593 , n6594 , n6595 , n6596 , n6597 , n6598 , n6599 , n6600 , n6601 , n6602 , n6603 , n6604 , n6605 , n6606 , n6607 , n6608 , n6609 , n6610 , n6611 , n6612 , n6613 , n6614 , n6615 , n6616 , n6617 , n6618 , n6619 , n6620 , n6621 , n6622 , n6623 , n6624 , n6625 , n6626 , n6627 , n6628 , n6629 , n6630 , n6631 , n6632 , n6633 , n6634 , n6635 , n6636 , n6637 , n6638 , n6639 , n6640 , n6641 , n6642 , n6643 , n6644 , n6645 , n6646 , n6647 , n6648 , n6649 , n6650 , n6651 , n6652 , n6653 , n6654 , n6655 , n6656 , n6657 , n6658 , n6659 , n6660 , n6661 , n6662 , n6663 , n6664 , n6665 , n6666 , n6667 , n6668 , n6669 , n6670 , n6671 , n6672 , n6673 , n6674 , n6675 , n6676 , n6677 , n6678 , n6679 , n6680 , n6681 , n6682 , n6683 , n6684 , n6685 , n6686 , n6687 , n6688 , n6689 , n6690 , n6691 , n6692 , n6693 , n6694 , n6695 , n6696 , n6697 , n6698 , n6699 , n6700 , n6701 , n6702 , n6703 , n6704 , n6705 , n6706 , n6707 , n6708 , n6709 , n6710 , n6711 , n6712 , n6713 , n6714 , n6715 , n6716 , n6717 , n6718 , n6719 , n6720 , n6721 , n6722 , n6723 , n6724 , n6725 , n6726 , n6727 , n6728 , n6729 , n6730 , n6731 , n6732 , n6733 , n6734 , n6735 , n6736 , n6737 , n6738 , n6739 , n6740 , n6741 , n6742 , n6743 , n6744 , n6745 , n6746 , n6747 , n6748 , n6749 , n6750 , n6751 , n6752 , n6753 , n6754 , n6755 , n6756 , n6757 , n6758 , n6759 , n6760 , n6761 , n6762 , n6763 , n6764 , n6765 , n6766 , n6767 , n6768 , n6769 , n6770 , n6771 , n6772 , n6773 , n6774 , n6775 , n6776 , n6777 , n6778 , n6779 , n6780 , n6781 , n6782 , n6783 , n6784 , n6785 , n6786 , n6787 , n6788 , n6789 , n6790 , n6791 , n6792 , n6793 , n6794 , n6795 , n6796 , n6797 , n6798 , n6799 , n6800 , n6801 , n6802 , n6803 , n6804 , n6805 , n6806 , n6807 , n6808 , n6809 , n6810 , n6811 , n6812 , n6813 , n6814 , n6815 , n6816 , n6817 , n6818 , n6819 , n6820 , n6821 , n6822 , n6823 , n6824 , n6825 , n6826 , n6827 , n6828 , n6829 , n6830 , n6831 , n6832 , n6833 , n6834 , n6835 , n6836 , n6837 , n6838 , n6839 , n6840 , n6841 , n6842 , n6843 , n6844 , n6845 , n6846 , n6847 , n6848 , n6849 , n6850 , n6851 , n6852 , n6853 , n6854 , n6855 , n6856 , n6857 , n6858 , n6859 , n6860 , n6861 , n6862 , n6863 , n6864 , n6865 , n6866 , n6867 , n6868 , n6869 , n6870 , n6871 , n6872 , n6873 , n6874 , n6875 , n6876 , n6877 , n6878 , n6879 , n6880 , n6881 , n6882 , n6883 , n6884 , n6885 , n6886 , n6887 , n6888 , n6889 , n6890 , n6891 , n6892 , n6893 , n6894 , n6895 , n6896 , n6897 , n6898 , n6899 , n6900 , n6901 , n6902 , n6903 , n6904 , n6905 , n6906 , n6907 , n6908 , n6909 , n6910 , n6911 , n6912 , n6913 , n6914 , n6915 , n6916 , n6917 , n6918 , n6919 , n6920 , n6921 , n6922 , n6923 , n6924 , n6925 , n6926 , n6927 , n6928 , n6929 , n6930 , n6931 , n6932 , n6933 , n6934 , n6935 , n6936 , n6937 , n6938 , n6939 , n6940 , n6941 , n6942 , n6943 , n6944 , n6945 , n6946 , n6947 , n6948 , n6949 , n6950 , n6951 , n6952 , n6953 , n6954 , n6955 , n6956 , n6957 , n6958 , n6959 , n6960 , n6961 , n6962 , n6963 , n6964 , n6965 , n6966 , n6967 , n6968 , n6969 , n6970 , n6971 , n6972 , n6973 , n6974 , n6975 , n6976 , n6977 , n6978 , n6979 , n6980 , n6981 , n6982 , n6983 , n6984 , n6985 , n6986 , n6987 , n6988 , n6989 , n6990 , n6991 , n6992 , n6993 , n6994 , n6995 , n6996 , n6997 , n6998 , n6999 , n7000 , n7001 , n7002 , n7003 , n7004 , n7005 , n7006 , n7007 , n7008 , n7009 , n7010 , n7011 , n7012 , n7013 , n7014 , n7015 , n7016 , n7017 , n7018 , n7019 , n7020 , n7021 , n7022 , n7023 , n7024 , n7025 , n7026 , n7027 , n7028 , n7029 , n7030 , n7031 , n7032 , n7033 , n7034 , n7035 , n7036 , n7037 , n7038 , n7039 , n7040 , n7041 , n7042 , n7043 , n7044 , n7045 , n7046 , n7047 , n7048 , n7049 , n7050 , n7051 , n7052 , n7053 , n7054 , n7055 , n7056 , n7057 , n7058 , n7059 , n7060 , n7061 , n7062 , n7063 , n7064 , n7065 , n7066 , n7067 , n7068 , n7069 , n7070 , n7071 , n7072 , n7073 , n7074 , n7075 , n7076 , n7077 , n7078 , n7079 , n7080 , n7081 , n7082 , n7083 , n7084 , n7085 , n7086 , n7087 , n7088 , n7089 , n7090 , n7091 , n7092 , n7093 , n7094 , n7095 , n7096 , n7097 , n7098 , n7099 , n7100 , n7101 , n7102 , n7103 , n7104 , n7105 , n7106 , n7107 , n7108 , n7109 , n7110 , n7111 , n7112 , n7113 , n7114 , n7115 , n7116 , n7117 , n7118 , n7119 , n7120 , n7121 , n7122 , n7123 , n7124 , n7125 , n7126 , n7127 , n7128 , n7129 , n7130 , n7131 , n7132 , n7133 , n7134 , n7135 , n7136 , n7137 , n7138 , n7139 , n7140 , n7141 , n7142 , n7143 , n7144 , n7145 , n7146 , n7147 , n7148 , n7149 , n7150 , n7151 , n7152 , n7153 , n7154 , n7155 , n7156 , n7157 , n7158 , n7159 , n7160 , n7161 , n7162 , n7163 , n7164 , n7165 , n7166 , n7167 , n7168 , n7169 , n7170 , n7171 , n7172 , n7173 , n7174 , n7175 , n7176 , n7177 , n7178 , n7179 , n7180 , n7181 , n7182 , n7183 , n7184 , n7185 , n7186 , n7187 , n7188 , n7189 , n7190 , n7191 , n7192 , n7193 , n7194 , n7195 , n7196 , n7197 , n7198 , n7199 , n7200 , n7201 , n7202 , n7203 , n7204 , n7205 , n7206 , n7207 , n7208 , n7209 , n7210 , n7211 , n7212 , n7213 , n7214 , n7215 , n7216 , n7217 , n7218 , n7219 , n7220 , n7221 , n7222 , n7223 , n7224 , n7225 , n7226 , n7227 , n7228 , n7229 , n7230 , n7231 , n7232 , n7233 , n7234 , n7235 , n7236 , n7237 , n7238 , n7239 , n7240 , n7241 , n7242 , n7243 , n7244 , n7245 , n7246 , n7247 , n7248 , n7249 , n7250 , n7251 , n7252 , n7253 , n7254 , n7255 , n7256 , n7257 , n7258 , n7259 , n7260 , n7261 , n7262 , n7263 , n7264 , n7265 , n7266 , n7267 , n7268 , n7269 , n7270 , n7271 , n7272 , n7273 , n7274 , n7275 , n7276 , n7277 , n7278 , n7279 , n7280 , n7281 , n7282 , n7283 , n7284 , n7285 , n7286 , n7287 , n7288 , n7289 , n7290 , n7291 , n7292 , n7293 , n7294 , n7295 , n7296 , n7297 , n7298 , n7299 , n7300 , n7301 , n7302 , n7303 , n7304 , n7305 , n7306 , n7307 , n7308 , n7309 , n7310 , n7311 , n7312 , n7313 , n7314 , n7315 , n7316 , n7317 , n7318 , n7319 , n7320 , n7321 , n7322 , n7323 , n7324 , n7325 , n7326 , n7327 , n7328 , n7329 , n7330 , n7331 , n7332 , n7333 , n7334 , n7335 , n7336 , n7337 , n7338 , n7339 , n7340 , n7341 , n7342 , n7343 , n7344 , n7345 , n7346 , n7347 , n7348 , n7349 , n7350 , n7351 , n7352 , n7353 , n7354 , n7355 , n7356 , n7357 , n7358 , n7359 , n7360 , n7361 , n7362 , n7363 , n7364 , n7365 , n7366 , n7367 , n7368 , n7369 , n7370 , n7371 , n7372 , n7373 , n7374 , n7375 , n7376 , n7377 , n7378 , n7379 , n7380 , n7381 , n7382 , n7383 , n7384 , n7385 , n7386 , n7387 , n7388 , n7389 , n7390 , n7391 , n7392 , n7393 , n7394 , n7395 , n7396 , n7397 , n7398 , n7399 , n7400 , n7401 , n7402 , n7403 , n7404 , n7405 , n7406 , n7407 , n7408 , n7409 , n7410 , n7411 , n7412 , n7413 , n7414 , n7415 , n7416 , n7417 , n7418 , n7419 , n7420 , n7421 , n7422 , n7423 , n7424 , n7425 , n7426 , n7427 , n7428 , n7429 , n7430 , n7431 , n7432 , n7433 , n7434 , n7435 , n7436 , n7437 , n7438 , n7439 , n7440 , n7441 , n7442 , n7443 , n7444 , n7445 , n7446 , n7447 , n7448 , n7449 , n7450 , n7451 , n7452 , n7453 , n7454 , n7455 , n7456 , n7457 , n7458 , n7459 , n7460 , n7461 , n7462 , n7463 , n7464 , n7465 , n7466 , n7467 , n7468 , n7469 , n7470 , n7471 , n7472 , n7473 , n7474 , n7475 , n7476 , n7477 , n7478 , n7479 , n7480 , n7481 , n7482 , n7483 , n7484 , n7485 , n7486 , n7487 , n7488 , n7489 , n7490 , n7491 , n7492 , n7493 , n7494 , n7495 , n7496 , n7497 , n7498 , n7499 , n7500 , n7501 , n7502 , n7503 , n7504 , n7505 , n7506 , n7507 , n7508 , n7509 , n7510 , n7511 , n7512 , n7513 , n7514 , n7515 , n7516 , n7517 , n7518 , n7519 , n7520 , n7521 , n7522 , n7523 , n7524 , n7525 , n7526 , n7527 , n7528 , n7529 , n7530 , n7531 , n7532 , n7533 , n7534 , n7535 , n7536 , n7537 , n7538 , n7539 , n7540 , n7541 , n7542 , n7543 , n7544 , n7545 , n7546 , n7547 , n7548 , n7549 , n7550 , n7551 , n7552 , n7553 , n7554 , n7555 , n7556 , n7557 , n7558 , n7559 , n7560 , n7561 , n7562 , n7563 , n7564 , n7565 , n7566 , n7567 , n7568 , n7569 , n7570 , n7571 , n7572 , n7573 , n7574 , n7575 , n7576 , n7577 , n7578 , n7579 , n7580 , n7581 , n7582 , n7583 , n7584 , n7585 , n7586 , n7587 , n7588 , n7589 , n7590 , n7591 , n7592 , n7593 , n7594 , n7595 , n7596 , n7597 , n7598 , n7599 , n7600 , n7601 , n7602 , n7603 , n7604 , n7605 , n7606 , n7607 , n7608 , n7609 , n7610 , n7611 , n7612 , n7613 , n7614 , n7615 , n7616 , n7617 , n7618 , n7619 , n7620 , n7621 , n7622 , n7623 , n7624 , n7625 , n7626 , n7627 , n7628 , n7629 , n7630 , n7631 , n7632 , n7633 , n7634 , n7635 , n7636 , n7637 , n7638 , n7639 , n7640 , n7641 , n7642 , n7643 , n7644 , n7645 , n7646 , n7647 , n7648 , n7649 , n7650 , n7651 , n7652 , n7653 , n7654 , n7655 , n7656 , n7657 , n7658 , n7659 , n7660 , n7661 , n7662 , n7663 , n7664 , n7665 , n7666 , n7667 , n7668 , n7669 , n7670 , n7671 , n7672 , n7673 , n7674 , n7675 , n7676 , n7677 , n7678 , n7679 , n7680 , n7681 , n7682 , n7683 , n7684 , n7685 , n7686 , n7687 , n7688 , n7689 , n7690 , n7691 , n7692 , n7693 , n7694 , n7695 , n7696 , n7697 , n7698 , n7699 , n7700 , n7701 , n7702 , n7703 , n7704 , n7705 , n7706 , n7707 , n7708 , n7709 , n7710 , n7711 , n7712 , n7713 , n7714 , n7715 , n7716 , n7717 , n7718 , n7719 , n7720 , n7721 , n7722 , n7723 , n7724 , n7725 , n7726 , n7727 , n7728 , n7729 , n7730 , n7731 , n7732 , n7733 , n7734 , n7735 , n7736 , n7737 , n7738 , n7739 , n7740 , n7741 , n7742 , n7743 , n7744 , n7745 , n7746 , n7747 , n7748 , n7749 , n7750 , n7751 , n7752 , n7753 , n7754 , n7755 , n7756 , n7757 , n7758 , n7759 , n7760 , n7761 , n7762 , n7763 , n7764 , n7765 , n7766 , n7767 , n7768 , n7769 , n7770 , n7771 , n7772 , n7773 , n7774 , n7775 , n7776 , n7777 , n7778 , n7779 , n7780 , n7781 , n7782 , n7783 , n7784 , n7785 , n7786 , n7787 , n7788 , n7789 , n7790 , n7791 , n7792 , n7793 , n7794 , n7795 , n7796 , n7797 , n7798 , n7799 , n7800 , n7801 , n7802 , n7803 , n7804 , n7805 , n7806 , n7807 , n7808 , n7809 , n7810 , n7811 , n7812 , n7813 , n7814 , n7815 , n7816 , n7817 , n7818 , n7819 , n7820 , n7821 , n7822 , n7823 , n7824 , n7825 , n7826 , n7827 , n7828 , n7829 , n7830 , n7831 , n7832 , n7833 , n7834 , n7835 , n7836 , n7837 , n7838 , n7839 , n7840 , n7841 , n7842 , n7843 , n7844 , n7845 , n7846 , n7847 , n7848 , n7849 , n7850 , n7851 , n7852 , n7853 , n7854 , n7855 , n7856 , n7857 , n7858 , n7859 , n7860 , n7861 , n7862 , n7863 , n7864 , n7865 , n7866 , n7867 , n7868 , n7869 , n7870 , n7871 , n7872 , n7873 , n7874 , n7875 , n7876 , n7877 , n7878 , n7879 , n7880 , n7881 , n7882 , n7883 , n7884 , n7885 , n7886 , n7887 , n7888 , n7889 , n7890 , n7891 , n7892 , n7893 , n7894 , n7895 , n7896 , n7897 , n7898 , n7899 , n7900 , n7901 , n7902 , n7903 , n7904 , n7905 , n7906 , n7907 , n7908 , n7909 , n7910 , n7911 , n7912 , n7913 , n7914 , n7915 , n7916 , n7917 , n7918 , n7919 , n7920 , n7921 , n7922 , n7923 , n7924 , n7925 , n7926 , n7927 , n7928 , n7929 , n7930 , n7931 , n7932 , n7933 , n7934 , n7935 , n7936 , n7937 , n7938 , n7939 , n7940 , n7941 , n7942 , n7943 , n7944 , n7945 , n7946 , n7947 , n7948 , n7949 , n7950 , n7951 , n7952 , n7953 , n7954 , n7955 , n7956 , n7957 , n7958 , n7959 , n7960 , n7961 , n7962 , n7963 , n7964 , n7965 , n7966 , n7967 , n7968 , n7969 , n7970 , n7971 , n7972 , n7973 , n7974 , n7975 , n7976 , n7977 , n7978 , n7979 , n7980 , n7981 , n7982 , n7983 , n7984 , n7985 , n7986 , n7987 , n7988 , n7989 , n7990 , n7991 , n7992 , n7993 , n7994 , n7995 , n7996 , n7997 , n7998 , n7999 , n8000 , n8001 , n8002 , n8003 , n8004 , n8005 , n8006 , n8007 , n8008 , n8009 , n8010 , n8011 , n8012 , n8013 , n8014 , n8015 , n8016 , n8017 , n8018 , n8019 , n8020 , n8021 , n8022 , n8023 , n8024 , n8025 , n8026 , n8027 , n8028 , n8029 , n8030 , n8031 , n8032 , n8033 , n8034 , n8035 , n8036 , n8037 , n8038 , n8039 , n8040 , n8041 , n8042 , n8043 , n8044 , n8045 , n8046 , n8047 , n8048 , n8049 , n8050 , n8051 , n8052 , n8053 , n8054 , n8055 , n8056 , n8057 , n8058 , n8059 , n8060 , n8061 , n8062 , n8063 , n8064 , n8065 , n8066 , n8067 , n8068 , n8069 , n8070 , n8071 , n8072 , n8073 , n8074 , n8075 , n8076 , n8077 , n8078 , n8079 , n8080 , n8081 , n8082 , n8083 , n8084 , n8085 , n8086 , n8087 , n8088 , n8089 , n8090 , n8091 , n8092 , n8093 , n8094 , n8095 , n8096 , n8097 , n8098 , n8099 , n8100 , n8101 , n8102 , n8103 , n8104 , n8105 , n8106 , n8107 , n8108 , n8109 , n8110 , n8111 , n8112 , n8113 , n8114 , n8115 , n8116 , n8117 , n8118 , n8119 , n8120 , n8121 , n8122 , n8123 , n8124 , n8125 , n8126 , n8127 , n8128 , n8129 , n8130 , n8131 , n8132 , n8133 , n8134 , n8135 , n8136 , n8137 , n8138 , n8139 , n8140 , n8141 , n8142 , n8143 , n8144 , n8145 , n8146 , n8147 , n8148 , n8149 , n8150 , n8151 , n8152 , n8153 , n8154 , n8155 , n8156 , n8157 , n8158 , n8159 , n8160 , n8161 , n8162 , n8163 , n8164 , n8165 , n8166 , n8167 , n8168 , n8169 , n8170 , n8171 , n8172 , n8173 , n8174 , n8175 , n8176 , n8177 , n8178 , n8179 , n8180 , n8181 , n8182 , n8183 , n8184 , n8185 , n8186 , n8187 , n8188 , n8189 , n8190 , n8191 , n8192 , n8193 , n8194 , n8195 , n8196 , n8197 , n8198 , n8199 , n8200 , n8201 , n8202 , n8203 , n8204 , n8205 , n8206 , n8207 , n8208 , n8209 , n8210 , n8211 , n8212 , n8213 , n8214 , n8215 , n8216 , n8217 , n8218 , n8219 , n8220 , n8221 , n8222 , n8223 , n8224 , n8225 , n8226 , n8227 , n8228 , n8229 , n8230 , n8231 , n8232 , n8233 , n8234 , n8235 , n8236 , n8237 , n8238 , n8239 , n8240 , n8241 , n8242 , n8243 , n8244 , n8245 , n8246 , n8247 , n8248 , n8249 , n8250 , n8251 , n8252 , n8253 , n8254 , n8255 , n8256 , n8257 , n8258 , n8259 , n8260 , n8261 , n8262 , n8263 , n8264 , n8265 , n8266 , n8267 , n8268 , n8269 , n8270 , n8271 , n8272 , n8273 , n8274 , n8275 , n8276 , n8277 , n8278 , n8279 , n8280 , n8281 , n8282 , n8283 , n8284 , n8285 , n8286 , n8287 , n8288 , n8289 , n8290 , n8291 , n8292 , n8293 , n8294 , n8295 , n8296 , n8297 , n8298 , n8299 , n8300 , n8301 , n8302 , n8303 , n8304 , n8305 , n8306 , n8307 , n8308 , n8309 , n8310 , n8311 , n8312 , n8313 , n8314 , n8315 , n8316 , n8317 , n8318 , n8319 , n8320 , n8321 , n8322 , n8323 , n8324 , n8325 , n8326 , n8327 , n8328 , n8329 , n8330 , n8331 , n8332 , n8333 , n8334 , n8335 , n8336 , n8337 , n8338 , n8339 , n8340 , n8341 , n8342 , n8343 , n8344 , n8345 , n8346 , n8347 , n8348 , n8349 , n8350 , n8351 , n8352 , n8353 , n8354 , n8355 , n8356 , n8357 , n8358 , n8359 , n8360 , n8361 , n8362 , n8363 , n8364 , n8365 , n8366 , n8367 , n8368 , n8369 , n8370 , n8371 , n8372 , n8373 , n8374 , n8375 , n8376 , n8377 , n8378 , n8379 , n8380 , n8381 , n8382 , n8383 , n8384 , n8385 , n8386 , n8387 , n8388 , n8389 , n8390 , n8391 , n8392 , n8393 , n8394 , n8395 , n8396 , n8397 , n8398 , n8399 , n8400 , n8401 , n8402 , n8403 , n8404 , n8405 , n8406 , n8407 , n8408 , n8409 , n8410 , n8411 , n8412 , n8413 , n8414 , n8415 , n8416 , n8417 , n8418 , n8419 , n8420 , n8421 , n8422 , n8423 , n8424 , n8425 , n8426 , n8427 , n8428 , n8429 , n8430 , n8431 , n8432 , n8433 , n8434 , n8435 , n8436 , n8437 , n8438 , n8439 , n8440 , n8441 , n8442 , n8443 , n8444 , n8445 , n8446 , n8447 , n8448 , n8449 , n8450 , n8451 , n8452 , n8453 , n8454 , n8455 , n8456 , n8457 , n8458 , n8459 , n8460 , n8461 , n8462 , n8463 , n8464 , n8465 , n8466 , n8467 , n8468 , n8469 , n8470 , n8471 , n8472 , n8473 , n8474 , n8475 , n8476 , n8477 , n8478 , n8479 , n8480 , n8481 , n8482 , n8483 , n8484 , n8485 , n8486 , n8487 , n8488 , n8489 , n8490 , n8491 , n8492 , n8493 , n8494 , n8495 , n8496 , n8497 , n8498 , n8499 , n8500 , n8501 , n8502 , n8503 , n8504 , n8505 , n8506 , n8507 , n8508 , n8509 , n8510 , n8511 , n8512 , n8513 , n8514 , n8515 , n8516 , n8517 , n8518 , n8519 , n8520 , n8521 , n8522 , n8523 , n8524 , n8525 , n8526 , n8527 , n8528 , n8529 , n8530 , n8531 , n8532 , n8533 , n8534 , n8535 , n8536 , n8537 , n8538 , n8539 , n8540 , n8541 , n8542 , n8543 , n8544 , n8545 , n8546 , n8547 , n8548 , n8549 , n8550 , n8551 , n8552 , n8553 , n8554 , n8555 , n8556 , n8557 , n8558 , n8559 , n8560 , n8561 , n8562 , n8563 , n8564 , n8565 , n8566 , n8567 , n8568 , n8569 , n8570 , n8571 , n8572 , n8573 , n8574 , n8575 , n8576 , n8577 , n8578 , n8579 , n8580 , n8581 , n8582 , n8583 , n8584 , n8585 , n8586 , n8587 , n8588 , n8589 , n8590 , n8591 , n8592 , n8593 , n8594 , n8595 , n8596 , n8597 , n8598 , n8599 , n8600 , n8601 , n8602 , n8603 , n8604 , n8605 , n8606 , n8607 , n8608 , n8609 , n8610 , n8611 , n8612 , n8613 , n8614 , n8615 , n8616 , n8617 , n8618 , n8619 , n8620 , n8621 , n8622 , n8623 , n8624 , n8625 , n8626 , n8627 , n8628 , n8629 , n8630 , n8631 , n8632 , n8633 , n8634 , n8635 , n8636 , n8637 , n8638 , n8639 , n8640 , n8641 , n8642 , n8643 , n8644 , n8645 , n8646 , n8647 , n8648 , n8649 , n8650 , n8651 , n8652 , n8653 , n8654 , n8655 , n8656 , n8657 , n8658 , n8659 , n8660 , n8661 , n8662 , n8663 , n8664 , n8665 , n8666 , n8667 , n8668 , n8669 , n8670 , n8671 , n8672 , n8673 , n8674 , n8675 , n8676 , n8677 , n8678 , n8679 , n8680 , n8681 , n8682 , n8683 , n8684 , n8685 , n8686 , n8687 , n8688 , n8689 , n8690 , n8691 , n8692 , n8693 , n8694 , n8695 , n8696 , n8697 , n8698 , n8699 , n8700 , n8701 , n8702 , n8703 , n8704 , n8705 , n8706 , n8707 , n8708 , n8709 , n8710 , n8711 , n8712 , n8713 , n8714 , n8715 , n8716 , n8717 , n8718 , n8719 , n8720 , n8721 , n8722 , n8723 , n8724 , n8725 , n8726 , n8727 , n8728 , n8729 , n8730 , n8731 , n8732 , n8733 , n8734 , n8735 , n8736 , n8737 , n8738 , n8739 , n8740 , n8741 , n8742 , n8743 , n8744 , n8745 , n8746 , n8747 , n8748 , n8749 , n8750 , n8751 , n8752 , n8753 , n8754 , n8755 , n8756 , n8757 , n8758 , n8759 , n8760 , n8761 , n8762 , n8763 , n8764 , n8765 , n8766 , n8767 , n8768 , n8769 , n8770 , n8771 , n8772 , n8773 , n8774 , n8775 , n8776 , n8777 , n8778 , n8779 , n8780 , n8781 , n8782 , n8783 , n8784 , n8785 , n8786 , n8787 , n8788 , n8789 , n8790 , n8791 , n8792 , n8793 , n8794 , n8795 , n8796 , n8797 , n8798 , n8799 , n8800 , n8801 , n8802 , n8803 , n8804 , n8805 , n8806 , n8807 , n8808 , n8809 , n8810 , n8811 , n8812 , n8813 , n8814 , n8815 , n8816 , n8817 , n8818 , n8819 , n8820 , n8821 , n8822 , n8823 , n8824 , n8825 , n8826 , n8827 , n8828 , n8829 , n8830 , n8831 , n8832 , n8833 , n8834 , n8835 , n8836 , n8837 , n8838 , n8839 , n8840 , n8841 , n8842 , n8843 , n8844 , n8845 , n8846 , n8847 , n8848 , n8849 , n8850 , n8851 , n8852 , n8853 , n8854 , n8855 , n8856 , n8857 , n8858 , n8859 , n8860 , n8861 , n8862 , n8863 , n8864 , n8865 , n8866 , n8867 , n8868 , n8869 , n8870 , n8871 , n8872 , n8873 , n8874 , n8875 , n8876 , n8877 , n8878 , n8879 , n8880 , n8881 , n8882 , n8883 , n8884 , n8885 , n8886 , n8887 , n8888 , n8889 , n8890 , n8891 , n8892 , n8893 , n8894 , n8895 , n8896 , n8897 , n8898 , n8899 , n8900 , n8901 , n8902 , n8903 , n8904 , n8905 , n8906 , n8907 , n8908 , n8909 , n8910 , n8911 , n8912 , n8913 , n8914 , n8915 , n8916 , n8917 , n8918 , n8919 , n8920 , n8921 , n8922 , n8923 , n8924 , n8925 , n8926 , n8927 , n8928 , n8929 , n8930 , n8931 , n8932 , n8933 , n8934 , n8935 , n8936 , n8937 , n8938 , n8939 , n8940 , n8941 , n8942 , n8943 , n8944 , n8945 , n8946 , n8947 , n8948 , n8949 , n8950 , n8951 , n8952 , n8953 , n8954 , n8955 , n8956 , n8957 , n8958 , n8959 , n8960 , n8961 , n8962 , n8963 , n8964 , n8965 , n8966 , n8967 , n8968 , n8969 , n8970 , n8971 , n8972 , n8973 , n8974 , n8975 , n8976 , n8977 , n8978 , n8979 , n8980 , n8981 , n8982 , n8983 , n8984 , n8985 , n8986 , n8987 , n8988 , n8989 , n8990 , n8991 , n8992 , n8993 , n8994 , n8995 , n8996 , n8997 , n8998 , n8999 , n9000 , n9001 , n9002 , n9003 , n9004 , n9005 , n9006 , n9007 , n9008 , n9009 , n9010 , n9011 , n9012 , n9013 , n9014 , n9015 , n9016 , n9017 , n9018 , n9019 , n9020 , n9021 , n9022 , n9023 , n9024 , n9025 , n9026 , n9027 , n9028 , n9029 , n9030 , n9031 , n9032 , n9033 , n9034 , n9035 , n9036 , n9037 , n9038 , n9039 , n9040 , n9041 , n9042 , n9043 , n9044 , n9045 , n9046 , n9047 , n9048 , n9049 , n9050 , n9051 , n9052 , n9053 , n9054 , n9055 , n9056 , n9057 , n9058 , n9059 , n9060 , n9061 , n9062 , n9063 , n9064 , n9065 , n9066 , n9067 , n9068 , n9069 , n9070 , n9071 , n9072 , n9073 , n9074 , n9075 , n9076 , n9077 , n9078 , n9079 , n9080 , n9081 , n9082 , n9083 , n9084 , n9085 , n9086 , n9087 , n9088 , n9089 , n9090 , n9091 , n9092 , n9093 , n9094 , n9095 , n9096 , n9097 , n9098 , n9099 , n9100 , n9101 , n9102 , n9103 , n9104 , n9105 , n9106 , n9107 , n9108 , n9109 , n9110 , n9111 , n9112 , n9113 , n9114 , n9115 , n9116 , n9117 , n9118 , n9119 , n9120 , n9121 , n9122 , n9123 , n9124 , n9125 , n9126 , n9127 , n9128 , n9129 , n9130 , n9131 , n9132 , n9133 , n9134 , n9135 , n9136 , n9137 , n9138 , n9139 , n9140 , n9141 , n9142 , n9143 , n9144 , n9145 , n9146 , n9147 , n9148 , n9149 , n9150 , n9151 , n9152 , n9153 , n9154 , n9155 , n9156 , n9157 , n9158 , n9159 , n9160 , n9161 , n9162 , n9163 , n9164 , n9165 , n9166 , n9167 , n9168 , n9169 , n9170 , n9171 , n9172 , n9173 , n9174 , n9175 , n9176 , n9177 , n9178 , n9179 , n9180 , n9181 , n9182 , n9183 , n9184 , n9185 , n9186 , n9187 , n9188 , n9189 , n9190 , n9191 , n9192 , n9193 , n9194 , n9195 , n9196 , n9197 , n9198 , n9199 , n9200 , n9201 , n9202 , n9203 , n9204 , n9205 , n9206 , n9207 , n9208 , n9209 , n9210 , n9211 , n9212 , n9213 , n9214 , n9215 , n9216 , n9217 , n9218 , n9219 , n9220 , n9221 , n9222 , n9223 , n9224 , n9225 , n9226 , n9227 , n9228 , n9229 , n9230 , n9231 , n9232 , n9233 , n9234 , n9235 , n9236 , n9237 , n9238 , n9239 , n9240 , n9241 , n9242 , n9243 , n9244 , n9245 , n9246 , n9247 , n9248 , n9249 , n9250 , n9251 , n9252 , n9253 , n9254 , n9255 , n9256 , n9257 , n9258 , n9259 , n9260 , n9261 , n9262 , n9263 , n9264 , n9265 , n9266 , n9267 , n9268 , n9269 , n9270 , n9271 , n9272 , n9273 , n9274 , n9275 , n9276 , n9277 , n9278 , n9279 , n9280 , n9281 , n9282 , n9283 , n9284 , n9285 , n9286 , n9287 , n9288 , n9289 , n9290 , n9291 , n9292 , n9293 , n9294 , n9295 , n9296 , n9297 , n9298 , n9299 , n9300 , n9301 , n9302 , n9303 , n9304 , n9305 , n9306 , n9307 , n9308 , n9309 , n9310 , n9311 , n9312 , n9313 , n9314 , n9315 , n9316 , n9317 , n9318 , n9319 , n9320 , n9321 , n9322 , n9323 , n9324 , n9325 , n9326 , n9327 , n9328 , n9329 , n9330 , n9331 , n9332 , n9333 , n9334 , n9335 , n9336 , n9337 , n9338 , n9339 , n9340 , n9341 , n9342 , n9343 , n9344 , n9345 , n9346 , n9347 , n9348 , n9349 , n9350 , n9351 , n9352 , n9353 , n9354 , n9355 , n9356 , n9357 , n9358 , n9359 , n9360 , n9361 , n9362 , n9363 , n9364 , n9365 , n9366 , n9367 , n9368 , n9369 , n9370 , n9371 , n9372 , n9373 , n9374 , n9375 , n9376 , n9377 , n9378 , n9379 , n9380 , n9381 , n9382 , n9383 , n9384 , n9385 , n9386 , n9387 , n9388 , n9389 , n9390 , n9391 , n9392 , n9393 , n9394 , n9395 , n9396 , n9397 , n9398 , n9399 , n9400 , n9401 , n9402 , n9403 , n9404 , n9405 , n9406 , n9407 , n9408 , n9409 , n9410 , n9411 , n9412 , n9413 , n9414 , n9415 , n9416 , n9417 , n9418 , n9419 , n9420 , n9421 , n9422 , n9423 , n9424 , n9425 , n9426 , n9427 , n9428 , n9429 , n9430 , n9431 , n9432 , n9433 , n9434 , n9435 , n9436 , n9437 , n9438 , n9439 , n9440 , n9441 , n9442 , n9443 , n9444 , n9445 , n9446 , n9447 , n9448 , n9449 , n9450 , n9451 , n9452 , n9453 , n9454 , n9455 , n9456 , n9457 , n9458 , n9459 , n9460 , n9461 , n9462 , n9463 , n9464 , n9465 , n9466 , n9467 , n9468 , n9469 , n9470 , n9471 , n9472 , n9473 , n9474 , n9475 , n9476 , n9477 , n9478 , n9479 , n9480 , n9481 , n9482 , n9483 , n9484 , n9485 , n9486 , n9487 , n9488 , n9489 , n9490 , n9491 , n9492 , n9493 , n9494 , n9495 , n9496 , n9497 , n9498 , n9499 , n9500 , n9501 , n9502 , n9503 , n9504 , n9505 , n9506 , n9507 , n9508 , n9509 , n9510 , n9511 , n9512 , n9513 , n9514 , n9515 , n9516 , n9517 , n9518 , n9519 , n9520 , n9521 , n9522 , n9523 , n9524 , n9525 , n9526 , n9527 , n9528 , n9529 , n9530 , n9531 , n9532 , n9533 , n9534 , n9535 , n9536 , n9537 , n9538 , n9539 , n9540 , n9541 , n9542 , n9543 , n9544 , n9545 , n9546 , n9547 , n9548 , n9549 , n9550 , n9551 , n9552 , n9553 , n9554 , n9555 , n9556 , n9557 , n9558 , n9559 , n9560 , n9561 , n9562 , n9563 , n9564 , n9565 , n9566 , n9567 , n9568 , n9569 , n9570 , n9571 , n9572 , n9573 , n9574 , n9575 , n9576 , n9577 , n9578 , n9579 , n9580 , n9581 , n9582 , n9583 , n9584 , n9585 , n9586 , n9587 , n9588 , n9589 , n9590 , n9591 , n9592 , n9593 , n9594 , n9595 , n9596 , n9597 , n9598 , n9599 , n9600 , n9601 , n9602 , n9603 , n9604 , n9605 , n9606 , n9607 , n9608 , n9609 , n9610 , n9611 , n9612 , n9613 , n9614 , n9615 , n9616 , n9617 , n9618 , n9619 , n9620 , n9621 , n9622 , n9623 , n9624 , n9625 , n9626 , n9627 , n9628 , n9629 , n9630 , n9631 , n9632 , n9633 , n9634 , n9635 , n9636 , n9637 , n9638 , n9639 , n9640 , n9641 , n9642 , n9643 , n9644 , n9645 , n9646 , n9647 , n9648 , n9649 , n9650 , n9651 , n9652 , n9653 , n9654 , n9655 , n9656 , n9657 , n9658 , n9659 , n9660 , n9661 , n9662 , n9663 , n9664 , n9665 , n9666 , n9667 , n9668 , n9669 , n9670 , n9671 , n9672 , n9673 , n9674 , n9675 , n9676 , n9677 , n9678 , n9679 , n9680 , n9681 , n9682 , n9683 , n9684 , n9685 , n9686 , n9687 , n9688 , n9689 , n9690 , n9691 , n9692 , n9693 , n9694 , n9695 , n9696 , n9697 , n9698 , n9699 , n9700 , n9701 , n9702 , n9703 , n9704 , n9705 , n9706 , n9707 , n9708 , n9709 , n9710 , n9711 , n9712 , n9713 , n9714 , n9715 , n9716 , n9717 , n9718 , n9719 , n9720 , n9721 , n9722 , n9723 , n9724 , n9725 , n9726 , n9727 , n9728 , n9729 , n9730 , n9731 , n9732 , n9733 , n9734 , n9735 , n9736 , n9737 , n9738 , n9739 , n9740 , n9741 , n9742 , n9743 , n9744 , n9745 , n9746 , n9747 , n9748 , n9749 , n9750 , n9751 , n9752 , n9753 , n9754 , n9755 , n9756 , n9757 , n9758 , n9759 , n9760 , n9761 , n9762 , n9763 , n9764 , n9765 , n9766 , n9767 , n9768 , n9769 , n9770 , n9771 , n9772 , n9773 , n9774 , n9775 , n9776 , n9777 , n9778 , n9779 , n9780 , n9781 , n9782 , n9783 , n9784 , n9785 , n9786 , n9787 , n9788 , n9789 , n9790 , n9791 , n9792 , n9793 , n9794 , n9795 , n9796 , n9797 , n9798 , n9799 , n9800 , n9801 , n9802 , n9803 , n9804 , n9805 , n9806 , n9807 , n9808 , n9809 , n9810 , n9811 , n9812 , n9813 , n9814 , n9815 , n9816 , n9817 , n9818 , n9819 , n9820 , n9821 , n9822 , n9823 , n9824 , n9825 , n9826 , n9827 , n9828 , n9829 , n9830 , n9831 , n9832 , n9833 , n9834 , n9835 , n9836 , n9837 , n9838 , n9839 , n9840 , n9841 , n9842 , n9843 , n9844 , n9845 , n9846 , n9847 , n9848 , n9849 , n9850 , n9851 , n9852 , n9853 , n9854 , n9855 , n9856 , n9857 , n9858 , n9859 , n9860 , n9861 , n9862 , n9863 , n9864 , n9865 , n9866 , n9867 , n9868 , n9869 , n9870 , n9871 , n9872 , n9873 , n9874 , n9875 , n9876 , n9877 , n9878 , n9879 , n9880 , n9881 , n9882 , n9883 , n9884 , n9885 , n9886 , n9887 , n9888 , n9889 , n9890 , n9891 , n9892 , n9893 , n9894 , n9895 , n9896 , n9897 , n9898 , n9899 , n9900 , n9901 , n9902 , n9903 , n9904 , n9905 , n9906 , n9907 , n9908 , n9909 , n9910 , n9911 , n9912 , n9913 , n9914 , n9915 , n9916 , n9917 , n9918 , n9919 , n9920 , n9921 , n9922 , n9923 , n9924 , n9925 , n9926 , n9927 , n9928 , n9929 , n9930 , n9931 , n9932 , n9933 , n9934 , n9935 , n9936 , n9937 , n9938 , n9939 , n9940 , n9941 , n9942 , n9943 , n9944 , n9945 , n9946 , n9947 , n9948 , n9949 , n9950 , n9951 , n9952 , n9953 , n9954 , n9955 , n9956 , n9957 , n9958 , n9959 , n9960 , n9961 , n9962 , n9963 , n9964 , n9965 , n9966 , n9967 , n9968 , n9969 , n9970 , n9971 , n9972 , n9973 , n9974 , n9975 , n9976 , n9977 , n9978 , n9979 , n9980 , n9981 , n9982 , n9983 , n9984 , n9985 , n9986 , n9987 , n9988 , n9989 , n9990 , n9991 , n9992 , n9993 , n9994 , n9995 , n9996 , n9997 , n9998 , n9999 , n10000 , n10001 , n10002 , n10003 , n10004 , n10005 , n10006 , n10007 , n10008 , n10009 , n10010 , n10011 , n10012 , n10013 , n10014 , n10015 , n10016 , n10017 , n10018 , n10019 , n10020 , n10021 , n10022 , n10023 , n10024 , n10025 , n10026 , n10027 , n10028 , n10029 , n10030 , n10031 , n10032 , n10033 , n10034 , n10035 , n10036 , n10037 , n10038 , n10039 , n10040 , n10041 , n10042 , n10043 , n10044 , n10045 , n10046 , n10047 , n10048 , n10049 , n10050 , n10051 , n10052 , n10053 , n10054 , n10055 , n10056 , n10057 , n10058 , n10059 , n10060 , n10061 , n10062 , n10063 , n10064 , n10065 , n10066 , n10067 , n10068 , n10069 , n10070 , n10071 , n10072 , n10073 , n10074 , n10075 , n10076 , n10077 , n10078 , n10079 , n10080 , n10081 , n10082 , n10083 , n10084 , n10085 , n10086 , n10087 , n10088 , n10089 , n10090 , n10091 , n10092 , n10093 , n10094 , n10095 , n10096 , n10097 , n10098 , n10099 , n10100 , n10101 , n10102 , n10103 , n10104 , n10105 , n10106 , n10107 , n10108 , n10109 , n10110 , n10111 , n10112 , n10113 , n10114 , n10115 , n10116 , n10117 , n10118 , n10119 , n10120 , n10121 , n10122 , n10123 , n10124 , n10125 , n10126 , n10127 , n10128 , n10129 , n10130 , n10131 , n10132 , n10133 , n10134 , n10135 , n10136 , n10137 , n10138 , n10139 , n10140 , n10141 , n10142 , n10143 , n10144 , n10145 , n10146 , n10147 , n10148 , n10149 , n10150 , n10151 , n10152 , n10153 , n10154 , n10155 , n10156 , n10157 , n10158 , n10159 , n10160 , n10161 , n10162 , n10163 , n10164 , n10165 , n10166 , n10167 , n10168 , n10169 , n10170 , n10171 , n10172 , n10173 , n10174 , n10175 , n10176 , n10177 , n10178 , n10179 , n10180 , n10181 , n10182 , n10183 , n10184 , n10185 , n10186 , n10187 , n10188 , n10189 , n10190 , n10191 , n10192 , n10193 , n10194 , n10195 , n10196 , n10197 , n10198 , n10199 , n10200 , n10201 , n10202 , n10203 , n10204 , n10205 , n10206 , n10207 , n10208 , n10209 , n10210 , n10211 , n10212 , n10213 , n10214 , n10215 , n10216 , n10217 , n10218 , n10219 , n10220 , n10221 , n10222 , n10223 , n10224 , n10225 , n10226 , n10227 , n10228 , n10229 , n10230 , n10231 , n10232 , n10233 , n10234 , n10235 , n10236 , n10237 , n10238 , n10239 , n10240 , n10241 , n10242 , n10243 , n10244 , n10245 , n10246 , n10247 , n10248 , n10249 , n10250 , n10251 , n10252 , n10253 , n10254 , n10255 , n10256 , n10257 , n10258 , n10259 , n10260 , n10261 , n10262 , n10263 , n10264 , n10265 , n10266 , n10267 , n10268 , n10269 , n10270 , n10271 , n10272 , n10273 , n10274 , n10275 , n10276 , n10277 , n10278 , n10279 , n10280 , n10281 , n10282 , n10283 , n10284 , n10285 , n10286 , n10287 , n10288 , n10289 , n10290 , n10291 , n10292 , n10293 , n10294 , n10295 , n10296 , n10297 , n10298 , n10299 , n10300 , n10301 , n10302 , n10303 , n10304 , n10305 , n10306 , n10307 , n10308 , n10309 , n10310 , n10311 , n10312 , n10313 , n10314 , n10315 , n10316 , n10317 , n10318 , n10319 , n10320 , n10321 , n10322 , n10323 , n10324 , n10325 , n10326 , n10327 , n10328 , n10329 , n10330 , n10331 , n10332 , n10333 , n10334 , n10335 , n10336 , n10337 , n10338 , n10339 , n10340 , n10341 , n10342 , n10343 , n10344 , n10345 , n10346 , n10347 , n10348 , n10349 , n10350 , n10351 , n10352 , n10353 , n10354 , n10355 , n10356 , n10357 , n10358 , n10359 , n10360 , n10361 , n10362 , n10363 , n10364 , n10365 , n10366 , n10367 , n10368 , n10369 , n10370 , n10371 , n10372 , n10373 , n10374 , n10375 , n10376 , n10377 , n10378 , n10379 , n10380 , n10381 , n10382 , n10383 , n10384 , n10385 , n10386 , n10387 , n10388 , n10389 , n10390 , n10391 , n10392 , n10393 , n10394 , n10395 , n10396 , n10397 , n10398 , n10399 , n10400 , n10401 , n10402 , n10403 , n10404 , n10405 , n10406 , n10407 , n10408 , n10409 , n10410 , n10411 , n10412 , n10413 , n10414 , n10415 , n10416 , n10417 , n10418 , n10419 , n10420 , n10421 , n10422 , n10423 , n10424 , n10425 , n10426 , n10427 , n10428 , n10429 , n10430 , n10431 , n10432 , n10433 , n10434 , n10435 , n10436 , n10437 , n10438 , n10439 , n10440 , n10441 , n10442 , n10443 , n10444 , n10445 , n10446 , n10447 , n10448 , n10449 , n10450 , n10451 , n10452 , n10453 , n10454 , n10455 , n10456 , n10457 , n10458 , n10459 , n10460 , n10461 , n10462 , n10463 , n10464 , n10465 , n10466 , n10467 , n10468 , n10469 , n10470 , n10471 , n10472 , n10473 , n10474 , n10475 , n10476 , n10477 , n10478 , n10479 , n10480 , n10481 , n10482 , n10483 , n10484 , n10485 , n10486 , n10487 , n10488 , n10489 , n10490 , n10491 , n10492 , n10493 , n10494 , n10495 , n10496 , n10497 , n10498 , n10499 , n10500 , n10501 , n10502 , n10503 , n10504 , n10505 , n10506 , n10507 , n10508 , n10509 , n10510 , n10511 , n10512 , n10513 , n10514 , n10515 , n10516 , n10517 , n10518 , n10519 , n10520 , n10521 , n10522 , n10523 , n10524 , n10525 , n10526 , n10527 , n10528 , n10529 , n10530 , n10531 , n10532 , n10533 , n10534 , n10535 , n10536 , n10537 , n10538 , n10539 , n10540 , n10541 , n10542 , n10543 , n10544 , n10545 , n10546 , n10547 , n10548 , n10549 , n10550 , n10551 , n10552 , n10553 , n10554 , n10555 , n10556 , n10557 , n10558 , n10559 , n10560 , n10561 , n10562 , n10563 , n10564 , n10565 , n10566 , n10567 , n10568 , n10569 , n10570 , n10571 , n10572 , n10573 , n10574 , n10575 , n10576 , n10577 , n10578 , n10579 , n10580 , n10581 , n10582 , n10583 , n10584 , n10585 , n10586 , n10587 , n10588 , n10589 , n10590 , n10591 , n10592 , n10593 , n10594 , n10595 , n10596 , n10597 , n10598 , n10599 , n10600 , n10601 , n10602 , n10603 , n10604 , n10605 , n10606 , n10607 , n10608 , n10609 , n10610 , n10611 , n10612 , n10613 , n10614 , n10615 , n10616 , n10617 , n10618 , n10619 , n10620 , n10621 , n10622 , n10623 , n10624 , n10625 , n10626 , n10627 , n10628 , n10629 , n10630 , n10631 , n10632 , n10633 , n10634 , n10635 , n10636 , n10637 , n10638 , n10639 , n10640 , n10641 , n10642 , n10643 , n10644 , n10645 , n10646 , n10647 , n10648 , n10649 , n10650 , n10651 , n10652 , n10653 , n10654 , n10655 , n10656 , n10657 , n10658 , n10659 , n10660 , n10661 , n10662 , n10663 , n10664 , n10665 , n10666 , n10667 , n10668 , n10669 , n10670 , n10671 , n10672 , n10673 , n10674 , n10675 , n10676 , n10677 , n10678 , n10679 , n10680 , n10681 , n10682 , n10683 , n10684 , n10685 , n10686 , n10687 , n10688 , n10689 , n10690 , n10691 , n10692 , n10693 , n10694 , n10695 , n10696 , n10697 , n10698 , n10699 , n10700 , n10701 , n10702 , n10703 , n10704 , n10705 , n10706 , n10707 , n10708 , n10709 , n10710 , n10711 , n10712 , n10713 , n10714 , n10715 , n10716 , n10717 , n10718 , n10719 , n10720 , n10721 , n10722 , n10723 , n10724 , n10725 , n10726 , n10727 , n10728 , n10729 , n10730 , n10731 , n10732 , n10733 , n10734 , n10735 , n10736 , n10737 , n10738 , n10739 , n10740 , n10741 , n10742 , n10743 , n10744 , n10745 , n10746 , n10747 , n10748 , n10749 , n10750 , n10751 , n10752 , n10753 , n10754 , n10755 , n10756 , n10757 , n10758 , n10759 , n10760 , n10761 , n10762 , n10763 , n10764 , n10765 , n10766 , n10767 , n10768 , n10769 , n10770 , n10771 , n10772 , n10773 , n10774 , n10775 , n10776 , n10777 , n10778 , n10779 , n10780 , n10781 , n10782 , n10783 , n10784 , n10785 , n10786 , n10787 , n10788 , n10789 , n10790 , n10791 , n10792 , n10793 , n10794 , n10795 , n10796 , n10797 , n10798 , n10799 , n10800 , n10801 , n10802 , n10803 , n10804 , n10805 , n10806 , n10807 , n10808 , n10809 , n10810 , n10811 , n10812 , n10813 , n10814 , n10815 , n10816 , n10817 , n10818 , n10819 , n10820 , n10821 , n10822 , n10823 , n10824 , n10825 , n10826 , n10827 , n10828 , n10829 , n10830 , n10831 , n10832 , n10833 , n10834 , n10835 , n10836 , n10837 , n10838 , n10839 , n10840 , n10841 , n10842 , n10843 , n10844 , n10845 , n10846 , n10847 , n10848 , n10849 , n10850 , n10851 , n10852 , n10853 , n10854 , n10855 , n10856 , n10857 , n10858 , n10859 , n10860 , n10861 , n10862 , n10863 , n10864 , n10865 , n10866 , n10867 , n10868 , n10869 , n10870 , n10871 , n10872 , n10873 , n10874 , n10875 , n10876 , n10877 , n10878 , n10879 , n10880 , n10881 , n10882 , n10883 , n10884 , n10885 , n10886 , n10887 , n10888 , n10889 , n10890 , n10891 , n10892 , n10893 , n10894 , n10895 , n10896 , n10897 , n10898 , n10899 , n10900 , n10901 , n10902 , n10903 , n10904 , n10905 , n10906 , n10907 , n10908 , n10909 , n10910 , n10911 , n10912 , n10913 , n10914 , n10915 , n10916 , n10917 , n10918 , n10919 , n10920 , n10921 , n10922 , n10923 , n10924 , n10925 , n10926 , n10927 , n10928 , n10929 , n10930 , n10931 , n10932 , n10933 , n10934 , n10935 , n10936 , n10937 , n10938 , n10939 , n10940 , n10941 , n10942 , n10943 , n10944 , n10945 , n10946 , n10947 , n10948 , n10949 , n10950 , n10951 , n10952 , n10953 , n10954 , n10955 , n10956 , n10957 , n10958 , n10959 , n10960 , n10961 , n10962 , n10963 , n10964 , n10965 , n10966 , n10967 , n10968 , n10969 , n10970 , n10971 , n10972 , n10973 , n10974 , n10975 , n10976 , n10977 , n10978 , n10979 , n10980 , n10981 , n10982 , n10983 , n10984 , n10985 , n10986 , n10987 , n10988 , n10989 , n10990 , n10991 , n10992 , n10993 , n10994 , n10995 , n10996 , n10997 , n10998 , n10999 , n11000 , n11001 , n11002 , n11003 , n11004 , n11005 , n11006 , n11007 , n11008 , n11009 , n11010 , n11011 , n11012 , n11013 , n11014 , n11015 , n11016 , n11017 , n11018 , n11019 , n11020 , n11021 , n11022 , n11023 , n11024 , n11025 , n11026 , n11027 , n11028 , n11029 , n11030 , n11031 , n11032 , n11033 , n11034 , n11035 , n11036 , n11037 , n11038 , n11039 , n11040 , n11041 , n11042 , n11043 , n11044 , n11045 , n11046 , n11047 , n11048 , n11049 , n11050 , n11051 , n11052 , n11053 , n11054 , n11055 , n11056 , n11057 , n11058 , n11059 , n11060 , n11061 , n11062 , n11063 , n11064 , n11065 , n11066 , n11067 , n11068 , n11069 , n11070 , n11071 , n11072 , n11073 , n11074 , n11075 , n11076 , n11077 , n11078 , n11079 , n11080 , n11081 , n11082 , n11083 , n11084 , n11085 , n11086 , n11087 , n11088 , n11089 , n11090 , n11091 , n11092 , n11093 , n11094 , n11095 , n11096 , n11097 , n11098 , n11099 , n11100 , n11101 , n11102 , n11103 , n11104 , n11105 , n11106 , n11107 , n11108 , n11109 , n11110 , n11111 , n11112 , n11113 , n11114 , n11115 , n11116 , n11117 , n11118 , n11119 , n11120 , n11121 , n11122 , n11123 , n11124 , n11125 , n11126 , n11127 , n11128 , n11129 , n11130 , n11131 , n11132 , n11133 , n11134 , n11135 , n11136 , n11137 , n11138 , n11139 , n11140 , n11141 , n11142 , n11143 , n11144 , n11145 , n11146 , n11147 , n11148 , n11149 , n11150 , n11151 , n11152 , n11153 , n11154 , n11155 , n11156 , n11157 , n11158 , n11159 , n11160 , n11161 , n11162 , n11163 , n11164 , n11165 , n11166 , n11167 , n11168 , n11169 , n11170 , n11171 , n11172 , n11173 , n11174 , n11175 , n11176 , n11177 , n11178 , n11179 , n11180 , n11181 , n11182 , n11183 , n11184 , n11185 , n11186 , n11187 , n11188 , n11189 , n11190 , n11191 , n11192 , n11193 , n11194 , n11195 , n11196 , n11197 , n11198 , n11199 , n11200 , n11201 , n11202 , n11203 , n11204 , n11205 , n11206 , n11207 , n11208 , n11209 , n11210 , n11211 , n11212 , n11213 , n11214 , n11215 , n11216 , n11217 , n11218 , n11219 , n11220 , n11221 , n11222 , n11223 , n11224 , n11225 , n11226 , n11227 , n11228 , n11229 , n11230 , n11231 , n11232 , n11233 , n11234 , n11235 , n11236 , n11237 , n11238 , n11239 , n11240 , n11241 , n11242 , n11243 , n11244 , n11245 , n11246 , n11247 , n11248 , n11249 , n11250 , n11251 , n11252 , n11253 , n11254 , n11255 , n11256 , n11257 , n11258 , n11259 , n11260 , n11261 , n11262 , n11263 , n11264 , n11265 , n11266 , n11267 , n11268 , n11269 , n11270 , n11271 , n11272 , n11273 , n11274 , n11275 , n11276 , n11277 , n11278 , n11279 , n11280 , n11281 , n11282 , n11283 , n11284 , n11285 , n11286 , n11287 , n11288 , n11289 , n11290 , n11291 , n11292 , n11293 , n11294 , n11295 , n11296 , n11297 , n11298 , n11299 , n11300 , n11301 , n11302 , n11303 , n11304 , n11305 , n11306 , n11307 , n11308 , n11309 , n11310 , n11311 , n11312 , n11313 , n11314 , n11315 , n11316 , n11317 , n11318 , n11319 , n11320 , n11321 , n11322 , n11323 , n11324 , n11325 , n11326 , n11327 , n11328 , n11329 , n11330 , n11331 , n11332 , n11333 , n11334 , n11335 , n11336 , n11337 , n11338 , n11339 , n11340 , n11341 , n11342 , n11343 , n11344 , n11345 , n11346 , n11347 , n11348 , n11349 , n11350 , n11351 , n11352 , n11353 , n11354 , n11355 , n11356 , n11357 , n11358 , n11359 , n11360 , n11361 , n11362 , n11363 , n11364 , n11365 , n11366 , n11367 , n11368 , n11369 , n11370 , n11371 , n11372 , n11373 , n11374 , n11375 , n11376 , n11377 , n11378 , n11379 , n11380 , n11381 , n11382 , n11383 , n11384 , n11385 , n11386 , n11387 , n11388 , n11389 , n11390 , n11391 , n11392 , n11393 , n11394 , n11395 , n11396 , n11397 , n11398 , n11399 , n11400 , n11401 , n11402 , n11403 , n11404 , n11405 , n11406 , n11407 , n11408 , n11409 , n11410 , n11411 , n11412 , n11413 , n11414 , n11415 , n11416 , n11417 , n11418 , n11419 , n11420 , n11421 , n11422 , n11423 , n11424 , n11425 , n11426 , n11427 , n11428 , n11429 , n11430 , n11431 , n11432 , n11433 , n11434 , n11435 , n11436 , n11437 , n11438 , n11439 , n11440 , n11441 , n11442 , n11443 , n11444 , n11445 , n11446 , n11447 , n11448 , n11449 , n11450 , n11451 , n11452 , n11453 , n11454 , n11455 , n11456 , n11457 , n11458 , n11459 , n11460 , n11461 , n11462 , n11463 , n11464 , n11465 , n11466 , n11467 , n11468 , n11469 , n11470 , n11471 , n11472 , n11473 , n11474 , n11475 , n11476 , n11477 , n11478 , n11479 , n11480 , n11481 , n11482 , n11483 , n11484 , n11485 , n11486 , n11487 , n11488 , n11489 , n11490 , n11491 , n11492 , n11493 , n11494 , n11495 , n11496 , n11497 , n11498 , n11499 , n11500 , n11501 , n11502 , n11503 , n11504 , n11505 , n11506 , n11507 , n11508 , n11509 , n11510 , n11511 , n11512 , n11513 , n11514 , n11515 , n11516 , n11517 , n11518 , n11519 , n11520 , n11521 , n11522 , n11523 , n11524 , n11525 , n11526 , n11527 , n11528 , n11529 , n11530 , n11531 , n11532 , n11533 , n11534 , n11535 , n11536 , n11537 , n11538 , n11539 , n11540 , n11541 , n11542 , n11543 , n11544 , n11545 , n11546 , n11547 , n11548 , n11549 , n11550 , n11551 , n11552 , n11553 , n11554 , n11555 , n11556 , n11557 , n11558 , n11559 , n11560 , n11561 , n11562 , n11563 , n11564 , n11565 , n11566 , n11567 , n11568 , n11569 , n11570 , n11571 , n11572 , n11573 , n11574 , n11575 , n11576 , n11577 , n11578 , n11579 , n11580 , n11581 , n11582 , n11583 , n11584 , n11585 , n11586 , n11587 , n11588 , n11589 , n11590 , n11591 , n11592 , n11593 , n11594 , n11595 , n11596 , n11597 , n11598 , n11599 , n11600 , n11601 , n11602 , n11603 , n11604 , n11605 , n11606 , n11607 , n11608 , n11609 , n11610 , n11611 , n11612 , n11613 , n11614 , n11615 , n11616 , n11617 , n11618 , n11619 , n11620 , n11621 , n11622 , n11623 , n11624 , n11625 , n11626 , n11627 , n11628 , n11629 , n11630 , n11631 , n11632 , n11633 , n11634 , n11635 , n11636 , n11637 , n11638 , n11639 , n11640 , n11641 , n11642 , n11643 , n11644 , n11645 , n11646 , n11647 , n11648 , n11649 , n11650 , n11651 , n11652 , n11653 , n11654 , n11655 , n11656 , n11657 , n11658 , n11659 , n11660 , n11661 , n11662 , n11663 , n11664 , n11665 , n11666 , n11667 , n11668 , n11669 , n11670 , n11671 , n11672 , n11673 , n11674 , n11675 , n11676 , n11677 , n11678 , n11679 , n11680 , n11681 , n11682 , n11683 , n11684 , n11685 , n11686 , n11687 , n11688 , n11689 , n11690 , n11691 , n11692 , n11693 , n11694 , n11695 , n11696 , n11697 , n11698 , n11699 , n11700 , n11701 , n11702 , n11703 , n11704 , n11705 , n11706 , n11707 , n11708 , n11709 , n11710 , n11711 , n11712 , n11713 , n11714 , n11715 , n11716 , n11717 , n11718 , n11719 , n11720 , n11721 , n11722 , n11723 , n11724 , n11725 , n11726 , n11727 , n11728 , n11729 , n11730 , n11731 , n11732 , n11733 , n11734 , n11735 , n11736 , n11737 , n11738 , n11739 , n11740 , n11741 , n11742 , n11743 , n11744 , n11745 , n11746 , n11747 , n11748 , n11749 , n11750 , n11751 , n11752 , n11753 , n11754 , n11755 , n11756 , n11757 , n11758 , n11759 , n11760 , n11761 , n11762 , n11763 , n11764 , n11765 , n11766 , n11767 , n11768 , n11769 , n11770 , n11771 , n11772 , n11773 , n11774 , n11775 , n11776 , n11777 , n11778 , n11779 , n11780 , n11781 , n11782 , n11783 , n11784 , n11785 , n11786 , n11787 , n11788 , n11789 , n11790 , n11791 , n11792 , n11793 , n11794 , n11795 , n11796 , n11797 , n11798 , n11799 , n11800 , n11801 , n11802 , n11803 , n11804 , n11805 , n11806 , n11807 , n11808 , n11809 , n11810 , n11811 , n11812 , n11813 , n11814 , n11815 , n11816 , n11817 , n11818 , n11819 , n11820 , n11821 , n11822 , n11823 , n11824 , n11825 , n11826 , n11827 , n11828 , n11829 , n11830 , n11831 , n11832 , n11833 , n11834 , n11835 , n11836 , n11837 , n11838 , n11839 , n11840 , n11841 , n11842 , n11843 , n11844 , n11845 , n11846 , n11847 , n11848 , n11849 , n11850 , n11851 , n11852 , n11853 , n11854 , n11855 , n11856 , n11857 , n11858 , n11859 , n11860 , n11861 , n11862 , n11863 , n11864 , n11865 , n11866 , n11867 , n11868 , n11869 , n11870 , n11871 , n11872 , n11873 , n11874 , n11875 , n11876 , n11877 , n11878 , n11879 , n11880 , n11881 , n11882 , n11883 , n11884 , n11885 , n11886 , n11887 , n11888 , n11889 , n11890 , n11891 , n11892 , n11893 , n11894 , n11895 , n11896 , n11897 , n11898 , n11899 , n11900 , n11901 , n11902 , n11903 , n11904 , n11905 , n11906 , n11907 , n11908 , n11909 , n11910 , n11911 , n11912 , n11913 , n11914 , n11915 , n11916 , n11917 , n11918 , n11919 , n11920 , n11921 , n11922 , n11923 , n11924 , n11925 , n11926 , n11927 , n11928 , n11929 , n11930 , n11931 , n11932 , n11933 , n11934 , n11935 , n11936 , n11937 , n11938 , n11939 , n11940 , n11941 , n11942 , n11943 , n11944 , n11945 , n11946 , n11947 , n11948 , n11949 , n11950 , n11951 , n11952 , n11953 , n11954 , n11955 , n11956 , n11957 , n11958 , n11959 , n11960 , n11961 , n11962 , n11963 , n11964 , n11965 , n11966 , n11967 , n11968 , n11969 , n11970 , n11971 , n11972 , n11973 , n11974 , n11975 , n11976 , n11977 , n11978 , n11979 , n11980 , n11981 , n11982 , n11983 , n11984 , n11985 , n11986 , n11987 , n11988 , n11989 , n11990 , n11991 , n11992 , n11993 , n11994 , n11995 , n11996 , n11997 , n11998 , n11999 , n12000 , n12001 , n12002 , n12003 , n12004 , n12005 , n12006 , n12007 , n12008 , n12009 , n12010 , n12011 , n12012 , n12013 , n12014 , n12015 , n12016 , n12017 , n12018 , n12019 , n12020 , n12021 , n12022 , n12023 , n12024 , n12025 , n12026 , n12027 , n12028 , n12029 , n12030 , n12031 , n12032 , n12033 , n12034 , n12035 , n12036 , n12037 , n12038 , n12039 , n12040 , n12041 , n12042 , n12043 , n12044 , n12045 , n12046 , n12047 , n12048 , n12049 , n12050 , n12051 , n12052 , n12053 , n12054 , n12055 , n12056 , n12057 , n12058 , n12059 , n12060 , n12061 , n12062 , n12063 , n12064 , n12065 , n12066 , n12067 , n12068 , n12069 , n12070 , n12071 , n12072 , n12073 , n12074 , n12075 , n12076 , n12077 , n12078 , n12079 , n12080 , n12081 , n12082 , n12083 , n12084 , n12085 , n12086 , n12087 , n12088 , n12089 , n12090 , n12091 , n12092 , n12093 , n12094 , n12095 , n12096 , n12097 , n12098 , n12099 , n12100 , n12101 , n12102 , n12103 , n12104 , n12105 , n12106 , n12107 , n12108 , n12109 , n12110 , n12111 , n12112 , n12113 , n12114 , n12115 , n12116 , n12117 , n12118 , n12119 , n12120 , n12121 , n12122 , n12123 , n12124 , n12125 , n12126 , n12127 , n12128 , n12129 , n12130 , n12131 , n12132 , n12133 , n12134 , n12135 , n12136 , n12137 , n12138 , n12139 , n12140 , n12141 , n12142 , n12143 , n12144 , n12145 , n12146 , n12147 , n12148 , n12149 , n12150 , n12151 , n12152 , n12153 , n12154 , n12155 , n12156 , n12157 , n12158 , n12159 , n12160 , n12161 , n12162 , n12163 , n12164 , n12165 , n12166 , n12167 , n12168 , n12169 , n12170 , n12171 , n12172 , n12173 , n12174 , n12175 , n12176 , n12177 , n12178 , n12179 , n12180 , n12181 , n12182 , n12183 , n12184 , n12185 , n12186 , n12187 , n12188 , n12189 , n12190 , n12191 , n12192 , n12193 , n12194 , n12195 , n12196 , n12197 , n12198 , n12199 , n12200 , n12201 , n12202 , n12203 , n12204 , n12205 , n12206 , n12207 , n12208 , n12209 , n12210 , n12211 , n12212 , n12213 , n12214 , n12215 , n12216 , n12217 , n12218 , n12219 , n12220 , n12221 , n12222 , n12223 , n12224 , n12225 , n12226 , n12227 , n12228 , n12229 , n12230 , n12231 , n12232 , n12233 , n12234 , n12235 , n12236 , n12237 , n12238 , n12239 , n12240 , n12241 , n12242 , n12243 , n12244 , n12245 , n12246 , n12247 , n12248 , n12249 , n12250 , n12251 , n12252 , n12253 , n12254 , n12255 , n12256 , n12257 , n12258 , n12259 , n12260 , n12261 , n12262 , n12263 , n12264 , n12265 , n12266 , n12267 , n12268 , n12269 , n12270 , n12271 , n12272 , n12273 , n12274 , n12275 , n12276 , n12277 , n12278 , n12279 , n12280 , n12281 , n12282 , n12283 , n12284 , n12285 , n12286 , n12287 , n12288 , n12289 , n12290 , n12291 , n12292 , n12293 , n12294 , n12295 , n12296 , n12297 , n12298 , n12299 , n12300 , n12301 , n12302 , n12303 , n12304 , n12305 , n12306 , n12307 , n12308 , n12309 , n12310 , n12311 , n12312 , n12313 , n12314 , n12315 , n12316 , n12317 , n12318 , n12319 , n12320 , n12321 , n12322 , n12323 , n12324 , n12325 , n12326 , n12327 , n12328 , n12329 , n12330 , n12331 , n12332 , n12333 , n12334 , n12335 , n12336 , n12337 , n12338 , n12339 , n12340 , n12341 , n12342 , n12343 , n12344 , n12345 , n12346 , n12347 , n12348 , n12349 , n12350 , n12351 , n12352 , n12353 , n12354 , n12355 , n12356 , n12357 , n12358 , n12359 , n12360 , n12361 , n12362 , n12363 , n12364 , n12365 , n12366 , n12367 , n12368 , n12369 , n12370 , n12371 , n12372 , n12373 , n12374 , n12375 , n12376 , n12377 , n12378 , n12379 , n12380 , n12381 , n12382 , n12383 , n12384 , n12385 , n12386 , n12387 , n12388 , n12389 , n12390 , n12391 , n12392 , n12393 , n12394 , n12395 , n12396 , n12397 , n12398 , n12399 , n12400 , n12401 , n12402 , n12403 , n12404 , n12405 , n12406 , n12407 , n12408 , n12409 , n12410 , n12411 , n12412 , n12413 , n12414 , n12415 , n12416 , n12417 , n12418 , n12419 , n12420 , n12421 , n12422 , n12423 , n12424 , n12425 , n12426 , n12427 , n12428 , n12429 , n12430 , n12431 , n12432 , n12433 , n12434 , n12435 , n12436 , n12437 , n12438 , n12439 , n12440 , n12441 , n12442 , n12443 , n12444 , n12445 , n12446 , n12447 , n12448 , n12449 , n12450 , n12451 , n12452 , n12453 , n12454 , n12455 , n12456 , n12457 , n12458 , n12459 , n12460 , n12461 , n12462 , n12463 , n12464 , n12465 , n12466 , n12467 , n12468 , n12469 , n12470 , n12471 , n12472 , n12473 , n12474 , n12475 , n12476 , n12477 , n12478 , n12479 , n12480 , n12481 , n12482 , n12483 , n12484 , n12485 , n12486 , n12487 , n12488 , n12489 , n12490 , n12491 , n12492 , n12493 , n12494 , n12495 , n12496 , n12497 , n12498 , n12499 , n12500 , n12501 , n12502 , n12503 , n12504 , n12505 , n12506 , n12507 , n12508 , n12509 , n12510 , n12511 , n12512 , n12513 , n12514 , n12515 , n12516 , n12517 , n12518 , n12519 , n12520 , n12521 , n12522 , n12523 , n12524 , n12525 , n12526 , n12527 , n12528 , n12529 , n12530 , n12531 , n12532 , n12533 , n12534 , n12535 , n12536 , n12537 , n12538 , n12539 , n12540 , n12541 , n12542 , n12543 , n12544 , n12545 , n12546 , n12547 , n12548 , n12549 , n12550 , n12551 , n12552 , n12553 , n12554 , n12555 , n12556 , n12557 , n12558 , n12559 , n12560 , n12561 , n12562 , n12563 , n12564 , n12565 , n12566 , n12567 , n12568 , n12569 , n12570 , n12571 , n12572 , n12573 , n12574 , n12575 , n12576 , n12577 , n12578 , n12579 , n12580 , n12581 , n12582 , n12583 , n12584 , n12585 , n12586 , n12587 , n12588 , n12589 , n12590 , n12591 , n12592 , n12593 , n12594 , n12595 , n12596 , n12597 , n12598 , n12599 , n12600 , n12601 , n12602 , n12603 , n12604 , n12605 , n12606 , n12607 , n12608 , n12609 , n12610 , n12611 , n12612 , n12613 , n12614 , n12615 , n12616 , n12617 , n12618 , n12619 , n12620 , n12621 , n12622 , n12623 , n12624 , n12625 , n12626 , n12627 , n12628 , n12629 , n12630 , n12631 , n12632 , n12633 , n12634 , n12635 , n12636 , n12637 , n12638 , n12639 , n12640 , n12641 , n12642 , n12643 , n12644 , n12645 , n12646 , n12647 , n12648 , n12649 , n12650 , n12651 , n12652 , n12653 , n12654 , n12655 , n12656 , n12657 , n12658 , n12659 , n12660 , n12661 , n12662 , n12663 , n12664 , n12665 , n12666 , n12667 , n12668 , n12669 , n12670 , n12671 , n12672 , n12673 , n12674 , n12675 , n12676 , n12677 , n12678 , n12679 , n12680 , n12681 , n12682 , n12683 , n12684 , n12685 , n12686 , n12687 , n12688 , n12689 , n12690 , n12691 , n12692 , n12693 , n12694 , n12695 , n12696 , n12697 , n12698 , n12699 , n12700 , n12701 , n12702 , n12703 , n12704 , n12705 , n12706 , n12707 , n12708 , n12709 , n12710 , n12711 , n12712 , n12713 , n12714 , n12715 , n12716 , n12717 , n12718 , n12719 , n12720 , n12721 , n12722 , n12723 , n12724 , n12725 , n12726 , n12727 , n12728 , n12729 , n12730 , n12731 , n12732 , n12733 , n12734 , n12735 , n12736 , n12737 , n12738 , n12739 , n12740 , n12741 , n12742 , n12743 , n12744 , n12745 , n12746 , n12747 , n12748 , n12749 , n12750 , n12751 , n12752 , n12753 , n12754 , n12755 , n12756 , n12757 , n12758 , n12759 , n12760 , n12761 , n12762 , n12763 , n12764 , n12765 , n12766 , n12767 , n12768 , n12769 , n12770 , n12771 , n12772 , n12773 , n12774 , n12775 , n12776 , n12777 , n12778 , n12779 , n12780 , n12781 , n12782 , n12783 , n12784 , n12785 , n12786 , n12787 , n12788 , n12789 , n12790 , n12791 , n12792 , n12793 , n12794 , n12795 , n12796 , n12797 , n12798 , n12799 , n12800 , n12801 , n12802 , n12803 , n12804 , n12805 , n12806 , n12807 , n12808 , n12809 , n12810 , n12811 , n12812 , n12813 , n12814 , n12815 , n12816 , n12817 , n12818 , n12819 , n12820 , n12821 , n12822 , n12823 , n12824 , n12825 , n12826 , n12827 , n12828 , n12829 , n12830 , n12831 , n12832 , n12833 , n12834 , n12835 , n12836 , n12837 , n12838 , n12839 , n12840 , n12841 , n12842 , n12843 , n12844 , n12845 , n12846 , n12847 , n12848 , n12849 , n12850 , n12851 , n12852 , n12853 , n12854 , n12855 , n12856 , n12857 , n12858 , n12859 , n12860 , n12861 , n12862 , n12863 , n12864 , n12865 , n12866 , n12867 , n12868 , n12869 , n12870 , n12871 , n12872 , n12873 , n12874 , n12875 , n12876 , n12877 , n12878 , n12879 , n12880 , n12881 , n12882 , n12883 , n12884 , n12885 , n12886 , n12887 , n12888 , n12889 , n12890 , n12891 , n12892 , n12893 , n12894 , n12895 , n12896 , n12897 , n12898 , n12899 , n12900 , n12901 , n12902 , n12903 , n12904 , n12905 , n12906 , n12907 , n12908 , n12909 , n12910 , n12911 , n12912 , n12913 , n12914 , n12915 , n12916 , n12917 , n12918 , n12919 , n12920 , n12921 , n12922 , n12923 , n12924 , n12925 , n12926 , n12927 , n12928 , n12929 , n12930 , n12931 , n12932 , n12933 , n12934 , n12935 , n12936 , n12937 , n12938 , n12939 , n12940 , n12941 , n12942 , n12943 , n12944 , n12945 , n12946 , n12947 , n12948 , n12949 , n12950 , n12951 , n12952 , n12953 , n12954 , n12955 , n12956 , n12957 , n12958 , n12959 , n12960 , n12961 , n12962 , n12963 , n12964 , n12965 , n12966 , n12967 , n12968 , n12969 , n12970 , n12971 , n12972 , n12973 , n12974 , n12975 , n12976 , n12977 , n12978 , n12979 , n12980 , n12981 , n12982 , n12983 , n12984 , n12985 , n12986 , n12987 , n12988 , n12989 , n12990 , n12991 , n12992 , n12993 , n12994 , n12995 , n12996 , n12997 , n12998 , n12999 , n13000 , n13001 , n13002 , n13003 , n13004 , n13005 , n13006 , n13007 , n13008 , n13009 , n13010 , n13011 , n13012 , n13013 , n13014 , n13015 , n13016 , n13017 , n13018 , n13019 , n13020 , n13021 , n13022 , n13023 , n13024 , n13025 , n13026 , n13027 , n13028 , n13029 , n13030 , n13031 , n13032 , n13033 , n13034 , n13035 , n13036 , n13037 , n13038 , n13039 , n13040 , n13041 , n13042 , n13043 , n13044 , n13045 , n13046 , n13047 , n13048 , n13049 , n13050 , n13051 , n13052 , n13053 , n13054 , n13055 , n13056 , n13057 , n13058 , n13059 , n13060 , n13061 , n13062 , n13063 , n13064 , n13065 , n13066 , n13067 , n13068 , n13069 , n13070 , n13071 , n13072 , n13073 , n13074 , n13075 , n13076 , n13077 , n13078 , n13079 , n13080 , n13081 , n13082 , n13083 , n13084 , n13085 , n13086 , n13087 , n13088 , n13089 , n13090 , n13091 , n13092 , n13093 , n13094 , n13095 , n13096 , n13097 , n13098 , n13099 , n13100 , n13101 , n13102 , n13103 , n13104 , n13105 , n13106 , n13107 , n13108 , n13109 , n13110 , n13111 , n13112 , n13113 , n13114 , n13115 , n13116 , n13117 , n13118 , n13119 , n13120 , n13121 , n13122 , n13123 , n13124 , n13125 , n13126 , n13127 , n13128 , n13129 , n13130 , n13131 , n13132 , n13133 , n13134 , n13135 , n13136 , n13137 , n13138 , n13139 , n13140 , n13141 , n13142 , n13143 , n13144 , n13145 , n13146 , n13147 , n13148 , n13149 , n13150 , n13151 , n13152 , n13153 , n13154 , n13155 , n13156 , n13157 , n13158 , n13159 , n13160 , n13161 , n13162 , n13163 , n13164 , n13165 , n13166 , n13167 , n13168 , n13169 , n13170 , n13171 , n13172 , n13173 , n13174 , n13175 , n13176 , n13177 , n13178 , n13179 , n13180 , n13181 , n13182 , n13183 , n13184 , n13185 , n13186 , n13187 , n13188 , n13189 , n13190 , n13191 , n13192 , n13193 , n13194 , n13195 , n13196 , n13197 , n13198 , n13199 , n13200 , n13201 , n13202 , n13203 , n13204 , n13205 , n13206 , n13207 , n13208 , n13209 , n13210 , n13211 , n13212 , n13213 , n13214 , n13215 , n13216 , n13217 , n13218 , n13219 , n13220 , n13221 , n13222 , n13223 , n13224 , n13225 , n13226 , n13227 , n13228 , n13229 , n13230 , n13231 , n13232 , n13233 , n13234 , n13235 , n13236 , n13237 , n13238 , n13239 , n13240 , n13241 , n13242 , n13243 , n13244 , n13245 , n13246 , n13247 , n13248 , n13249 , n13250 , n13251 , n13252 , n13253 , n13254 , n13255 , n13256 , n13257 , n13258 , n13259 , n13260 , n13261 , n13262 , n13263 , n13264 , n13265 , n13266 , n13267 , n13268 , n13269 , n13270 , n13271 , n13272 , n13273 , n13274 , n13275 , n13276 , n13277 , n13278 , n13279 , n13280 , n13281 , n13282 , n13283 , n13284 , n13285 , n13286 , n13287 , n13288 , n13289 , n13290 , n13291 , n13292 , n13293 , n13294 , n13295 , n13296 , n13297 , n13298 , n13299 , n13300 , n13301 , n13302 , n13303 , n13304 , n13305 , n13306 , n13307 , n13308 , n13309 , n13310 , n13311 , n13312 , n13313 , n13314 , n13315 , n13316 , n13317 , n13318 , n13319 , n13320 , n13321 , n13322 , n13323 , n13324 , n13325 , n13326 , n13327 , n13328 , n13329 , n13330 , n13331 , n13332 , n13333 , n13334 , n13335 , n13336 , n13337 , n13338 , n13339 , n13340 , n13341 , n13342 , n13343 , n13344 , n13345 , n13346 , n13347 , n13348 , n13349 , n13350 , n13351 , n13352 , n13353 , n13354 , n13355 , n13356 , n13357 , n13358 , n13359 , n13360 , n13361 , n13362 , n13363 , n13364 , n13365 , n13366 , n13367 , n13368 , n13369 , n13370 , n13371 , n13372 , n13373 , n13374 , n13375 , n13376 , n13377 , n13378 , n13379 , n13380 , n13381 , n13382 , n13383 , n13384 , n13385 , n13386 , n13387 , n13388 , n13389 , n13390 , n13391 , n13392 , n13393 , n13394 , n13395 , n13396 , n13397 , n13398 , n13399 , n13400 , n13401 , n13402 , n13403 , n13404 , n13405 , n13406 , n13407 , n13408 , n13409 , n13410 , n13411 , n13412 , n13413 , n13414 , n13415 , n13416 , n13417 , n13418 , n13419 , n13420 , n13421 , n13422 , n13423 , n13424 , n13425 , n13426 , n13427 , n13428 , n13429 , n13430 , n13431 , n13432 , n13433 , n13434 , n13435 , n13436 , n13437 , n13438 , n13439 , n13440 , n13441 , n13442 , n13443 , n13444 , n13445 , n13446 , n13447 , n13448 , n13449 , n13450 , n13451 , n13452 , n13453 , n13454 , n13455 , n13456 , n13457 , n13458 , n13459 , n13460 , n13461 , n13462 , n13463 , n13464 , n13465 , n13466 , n13467 , n13468 , n13469 , n13470 , n13471 , n13472 , n13473 , n13474 , n13475 , n13476 , n13477 , n13478 , n13479 , n13480 , n13481 , n13482 , n13483 , n13484 , n13485 , n13486 , n13487 , n13488 , n13489 , n13490 , n13491 , n13492 , n13493 , n13494 , n13495 , n13496 , n13497 , n13498 , n13499 , n13500 , n13501 , n13502 , n13503 , n13504 , n13505 , n13506 , n13507 , n13508 , n13509 , n13510 , n13511 , n13512 , n13513 , n13514 , n13515 , n13516 , n13517 , n13518 , n13519 , n13520 , n13521 , n13522 , n13523 , n13524 , n13525 , n13526 , n13527 , n13528 , n13529 , n13530 , n13531 , n13532 , n13533 , n13534 , n13535 , n13536 , n13537 , n13538 , n13539 , n13540 , n13541 , n13542 , n13543 , n13544 , n13545 , n13546 , n13547 , n13548 , n13549 , n13550 , n13551 , n13552 , n13553 , n13554 , n13555 , n13556 , n13557 , n13558 , n13559 , n13560 , n13561 , n13562 , n13563 , n13564 , n13565 , n13566 , n13567 , n13568 , n13569 , n13570 , n13571 , n13572 , n13573 , n13574 , n13575 , n13576 , n13577 , n13578 , n13579 , n13580 , n13581 , n13582 , n13583 , n13584 , n13585 , n13586 , n13587 , n13588 , n13589 , n13590 , n13591 , n13592 , n13593 , n13594 , n13595 , n13596 , n13597 , n13598 , n13599 , n13600 , n13601 , n13602 , n13603 , n13604 , n13605 , n13606 , n13607 , n13608 , n13609 , n13610 , n13611 , n13612 , n13613 , n13614 , n13615 , n13616 , n13617 , n13618 , n13619 , n13620 , n13621 , n13622 , n13623 , n13624 , n13625 , n13626 , n13627 , n13628 , n13629 , n13630 , n13631 , n13632 , n13633 , n13634 , n13635 , n13636 , n13637 , n13638 , n13639 , n13640 , n13641 , n13642 , n13643 , n13644 , n13645 , n13646 , n13647 , n13648 , n13649 , n13650 , n13651 , n13652 , n13653 , n13654 , n13655 , n13656 , n13657 , n13658 , n13659 , n13660 , n13661 , n13662 , n13663 , n13664 , n13665 , n13666 , n13667 , n13668 , n13669 , n13670 , n13671 , n13672 , n13673 , n13674 , n13675 , n13676 , n13677 , n13678 , n13679 , n13680 , n13681 , n13682 , n13683 , n13684 , n13685 , n13686 , n13687 , n13688 , n13689 , n13690 , n13691 , n13692 , n13693 , n13694 , n13695 , n13696 , n13697 , n13698 , n13699 , n13700 , n13701 , n13702 , n13703 , n13704 , n13705 , n13706 , n13707 , n13708 , n13709 , n13710 , n13711 , n13712 , n13713 , n13714 , n13715 , n13716 , n13717 , n13718 , n13719 , n13720 , n13721 , n13722 , n13723 , n13724 , n13725 , n13726 , n13727 , n13728 , n13729 , n13730 , n13731 , n13732 , n13733 , n13734 , n13735 , n13736 , n13737 , n13738 , n13739 , n13740 , n13741 , n13742 , n13743 , n13744 , n13745 , n13746 , n13747 , n13748 , n13749 , n13750 , n13751 , n13752 , n13753 , n13754 , n13755 , n13756 , n13757 , n13758 , n13759 , n13760 , n13761 , n13762 , n13763 , n13764 , n13765 , n13766 , n13767 , n13768 , n13769 , n13770 , n13771 , n13772 , n13773 , n13774 , n13775 , n13776 , n13777 , n13778 , n13779 , n13780 , n13781 , n13782 , n13783 , n13784 , n13785 , n13786 , n13787 , n13788 , n13789 , n13790 , n13791 , n13792 , n13793 , n13794 , n13795 , n13796 , n13797 , n13798 , n13799 , n13800 , n13801 , n13802 , n13803 , n13804 , n13805 , n13806 , n13807 , n13808 , n13809 , n13810 , n13811 , n13812 , n13813 , n13814 , n13815 , n13816 , n13817 , n13818 , n13819 , n13820 , n13821 , n13822 , n13823 , n13824 , n13825 , n13826 , n13827 , n13828 , n13829 , n13830 , n13831 , n13832 , n13833 , n13834 , n13835 , n13836 , n13837 , n13838 , n13839 , n13840 , n13841 , n13842 , n13843 , n13844 , n13845 , n13846 , n13847 , n13848 , n13849 , n13850 , n13851 , n13852 , n13853 , n13854 , n13855 , n13856 , n13857 , n13858 , n13859 , n13860 , n13861 , n13862 , n13863 , n13864 , n13865 , n13866 , n13867 , n13868 , n13869 , n13870 , n13871 , n13872 , n13873 , n13874 , n13875 , n13876 , n13877 , n13878 , n13879 , n13880 , n13881 , n13882 , n13883 , n13884 , n13885 , n13886 , n13887 , n13888 , n13889 , n13890 , n13891 , n13892 , n13893 , n13894 , n13895 , n13896 , n13897 , n13898 , n13899 , n13900 , n13901 , n13902 , n13903 , n13904 , n13905 , n13906 , n13907 , n13908 , n13909 , n13910 , n13911 , n13912 , n13913 , n13914 , n13915 , n13916 , n13917 , n13918 , n13919 , n13920 , n13921 , n13922 , n13923 , n13924 , n13925 , n13926 , n13927 , n13928 , n13929 , n13930 , n13931 , n13932 , n13933 , n13934 , n13935 , n13936 , n13937 , n13938 , n13939 , n13940 , n13941 , n13942 , n13943 , n13944 , n13945 , n13946 , n13947 , n13948 , n13949 , n13950 , n13951 , n13952 , n13953 , n13954 , n13955 , n13956 , n13957 , n13958 , n13959 , n13960 , n13961 , n13962 , n13963 , n13964 , n13965 , n13966 , n13967 , n13968 , n13969 , n13970 , n13971 , n13972 , n13973 , n13974 , n13975 , n13976 , n13977 , n13978 , n13979 , n13980 , n13981 , n13982 , n13983 , n13984 , n13985 , n13986 , n13987 , n13988 , n13989 , n13990 , n13991 , n13992 , n13993 , n13994 , n13995 , n13996 , n13997 , n13998 , n13999 , n14000 , n14001 , n14002 , n14003 , n14004 , n14005 , n14006 , n14007 , n14008 , n14009 , n14010 , n14011 , n14012 , n14013 , n14014 , n14015 , n14016 , n14017 , n14018 , n14019 , n14020 , n14021 , n14022 , n14023 , n14024 , n14025 , n14026 , n14027 , n14028 , n14029 , n14030 , n14031 , n14032 , n14033 , n14034 , n14035 , n14036 , n14037 , n14038 , n14039 , n14040 , n14041 , n14042 , n14043 , n14044 , n14045 , n14046 , n14047 , n14048 , n14049 , n14050 , n14051 , n14052 , n14053 , n14054 , n14055 , n14056 , n14057 , n14058 , n14059 , n14060 , n14061 , n14062 , n14063 , n14064 , n14065 , n14066 , n14067 , n14068 , n14069 , n14070 , n14071 , n14072 , n14073 , n14074 , n14075 , n14076 , n14077 , n14078 , n14079 , n14080 , n14081 , n14082 , n14083 , n14084 , n14085 , n14086 , n14087 , n14088 , n14089 , n14090 , n14091 , n14092 , n14093 , n14094 , n14095 , n14096 , n14097 , n14098 , n14099 , n14100 , n14101 , n14102 , n14103 , n14104 , n14105 , n14106 , n14107 , n14108 , n14109 , n14110 , n14111 , n14112 , n14113 , n14114 , n14115 , n14116 , n14117 , n14118 , n14119 , n14120 , n14121 , n14122 , n14123 , n14124 , n14125 , n14126 , n14127 , n14128 , n14129 , n14130 , n14131 , n14132 , n14133 , n14134 , n14135 , n14136 , n14137 , n14138 , n14139 , n14140 , n14141 , n14142 , n14143 , n14144 , n14145 , n14146 , n14147 , n14148 , n14149 , n14150 , n14151 , n14152 , n14153 , n14154 , n14155 , n14156 , n14157 , n14158 , n14159 , n14160 , n14161 , n14162 , n14163 , n14164 , n14165 , n14166 , n14167 , n14168 , n14169 , n14170 , n14171 , n14172 , n14173 , n14174 , n14175 , n14176 , n14177 , n14178 , n14179 , n14180 , n14181 , n14182 , n14183 , n14184 , n14185 , n14186 , n14187 , n14188 , n14189 , n14190 , n14191 , n14192 , n14193 , n14194 , n14195 , n14196 , n14197 , n14198 , n14199 , n14200 , n14201 , n14202 , n14203 , n14204 , n14205 , n14206 , n14207 , n14208 , n14209 , n14210 , n14211 , n14212 , n14213 , n14214 , n14215 , n14216 , n14217 , n14218 , n14219 , n14220 , n14221 , n14222 , n14223 , n14224 , n14225 , n14226 , n14227 , n14228 , n14229 , n14230 , n14231 , n14232 , n14233 , n14234 , n14235 , n14236 , n14237 , n14238 , n14239 , n14240 , n14241 , n14242 , n14243 , n14244 , n14245 , n14246 , n14247 , n14248 , n14249 , n14250 , n14251 , n14252 , n14253 , n14254 , n14255 , n14256 , n14257 , n14258 , n14259 , n14260 , n14261 , n14262 , n14263 , n14264 , n14265 , n14266 , n14267 , n14268 , n14269 , n14270 , n14271 , n14272 , n14273 , n14274 , n14275 , n14276 , n14277 , n14278 , n14279 , n14280 , n14281 , n14282 , n14283 , n14284 , n14285 , n14286 , n14287 , n14288 , n14289 , n14290 , n14291 , n14292 , n14293 , n14294 , n14295 , n14296 , n14297 , n14298 , n14299 , n14300 , n14301 , n14302 , n14303 , n14304 , n14305 , n14306 , n14307 , n14308 , n14309 , n14310 , n14311 , n14312 , n14313 , n14314 , n14315 , n14316 , n14317 , n14318 , n14319 , n14320 , n14321 , n14322 , n14323 , n14324 , n14325 , n14326 , n14327 , n14328 , n14329 , n14330 , n14331 , n14332 , n14333 , n14334 , n14335 , n14336 , n14337 , n14338 , n14339 , n14340 , n14341 , n14342 , n14343 , n14344 , n14345 , n14346 , n14347 , n14348 , n14349 , n14350 , n14351 , n14352 , n14353 , n14354 , n14355 , n14356 , n14357 , n14358 , n14359 , n14360 , n14361 , n14362 , n14363 , n14364 , n14365 , n14366 , n14367 , n14368 , n14369 , n14370 , n14371 , n14372 , n14373 , n14374 , n14375 , n14376 , n14377 , n14378 , n14379 , n14380 , n14381 , n14382 , n14383 , n14384 , n14385 , n14386 , n14387 , n14388 , n14389 , n14390 , n14391 , n14392 , n14393 , n14394 , n14395 , n14396 , n14397 , n14398 , n14399 , n14400 , n14401 , n14402 , n14403 , n14404 , n14405 , n14406 , n14407 , n14408 , n14409 , n14410 , n14411 , n14412 , n14413 , n14414 , n14415 , n14416 , n14417 , n14418 , n14419 , n14420 , n14421 , n14422 , n14423 , n14424 , n14425 , n14426 , n14427 , n14428 , n14429 , n14430 , n14431 , n14432 , n14433 , n14434 , n14435 , n14436 , n14437 , n14438 , n14439 , n14440 , n14441 , n14442 , n14443 , n14444 , n14445 , n14446 , n14447 , n14448 , n14449 , n14450 , n14451 , n14452 , n14453 , n14454 , n14455 , n14456 , n14457 , n14458 , n14459 , n14460 , n14461 , n14462 , n14463 , n14464 , n14465 , n14466 , n14467 , n14468 , n14469 , n14470 , n14471 , n14472 , n14473 , n14474 , n14475 , n14476 , n14477 , n14478 , n14479 , n14480 , n14481 , n14482 , n14483 , n14484 , n14485 , n14486 , n14487 , n14488 , n14489 , n14490 , n14491 , n14492 , n14493 , n14494 , n14495 , n14496 , n14497 , n14498 , n14499 , n14500 , n14501 , n14502 , n14503 , n14504 , n14505 , n14506 , n14507 , n14508 , n14509 , n14510 , n14511 , n14512 , n14513 , n14514 , n14515 , n14516 , n14517 , n14518 , n14519 , n14520 , n14521 , n14522 , n14523 , n14524 , n14525 , n14526 , n14527 , n14528 , n14529 , n14530 , n14531 , n14532 , n14533 , n14534 , n14535 , n14536 , n14537 , n14538 , n14539 , n14540 , n14541 , n14542 , n14543 , n14544 , n14545 , n14546 , n14547 , n14548 , n14549 , n14550 , n14551 , n14552 , n14553 , n14554 , n14555 , n14556 , n14557 , n14558 , n14559 , n14560 , n14561 , n14562 , n14563 , n14564 , n14565 , n14566 , n14567 , n14568 , n14569 , n14570 , n14571 , n14572 , n14573 , n14574 , n14575 , n14576 , n14577 , n14578 , n14579 , n14580 , n14581 , n14582 , n14583 , n14584 , n14585 , n14586 , n14587 , n14588 , n14589 , n14590 , n14591 , n14592 , n14593 , n14594 , n14595 , n14596 , n14597 , n14598 , n14599 , n14600 , n14601 , n14602 , n14603 , n14604 , n14605 , n14606 , n14607 , n14608 , n14609 , n14610 , n14611 , n14612 , n14613 , n14614 , n14615 , n14616 , n14617 , n14618 , n14619 , n14620 , n14621 , n14622 , n14623 , n14624 , n14625 , n14626 , n14627 , n14628 , n14629 , n14630 , n14631 , n14632 , n14633 , n14634 , n14635 , n14636 , n14637 , n14638 , n14639 , n14640 , n14641 , n14642 , n14643 , n14644 , n14645 , n14646 , n14647 , n14648 , n14649 , n14650 , n14651 , n14652 , n14653 , n14654 , n14655 , n14656 , n14657 , n14658 , n14659 , n14660 , n14661 , n14662 , n14663 , n14664 , n14665 , n14666 , n14667 , n14668 , n14669 , n14670 , n14671 , n14672 , n14673 , n14674 , n14675 , n14676 , n14677 , n14678 , n14679 , n14680 , n14681 , n14682 , n14683 , n14684 , n14685 , n14686 , n14687 , n14688 , n14689 , n14690 , n14691 , n14692 , n14693 , n14694 , n14695 , n14696 , n14697 , n14698 , n14699 , n14700 , n14701 , n14702 , n14703 , n14704 , n14705 , n14706 , n14707 , n14708 , n14709 , n14710 , n14711 , n14712 , n14713 , n14714 , n14715 , n14716 , n14717 , n14718 , n14719 , n14720 , n14721 , n14722 , n14723 , n14724 , n14725 , n14726 , n14727 , n14728 , n14729 , n14730 , n14731 , n14732 , n14733 , n14734 , n14735 , n14736 , n14737 , n14738 , n14739 , n14740 , n14741 , n14742 , n14743 , n14744 , n14745 , n14746 , n14747 , n14748 , n14749 , n14750 , n14751 , n14752 , n14753 , n14754 , n14755 , n14756 , n14757 , n14758 , n14759 , n14760 , n14761 , n14762 , n14763 , n14764 , n14765 , n14766 , n14767 , n14768 , n14769 , n14770 , n14771 , n14772 , n14773 , n14774 , n14775 , n14776 , n14777 , n14778 , n14779 , n14780 , n14781 , n14782 , n14783 , n14784 , n14785 , n14786 , n14787 , n14788 , n14789 , n14790 , n14791 , n14792 , n14793 , n14794 , n14795 , n14796 , n14797 , n14798 , n14799 , n14800 , n14801 , n14802 , n14803 , n14804 , n14805 , n14806 , n14807 , n14808 , n14809 , n14810 , n14811 , n14812 , n14813 , n14814 , n14815 , n14816 , n14817 , n14818 , n14819 , n14820 , n14821 , n14822 , n14823 , n14824 , n14825 , n14826 , n14827 , n14828 , n14829 , n14830 , n14831 , n14832 , n14833 , n14834 , n14835 , n14836 , n14837 , n14838 , n14839 , n14840 , n14841 , n14842 , n14843 , n14844 , n14845 , n14846 , n14847 , n14848 , n14849 , n14850 , n14851 , n14852 , n14853 , n14854 , n14855 , n14856 , n14857 , n14858 , n14859 , n14860 , n14861 , n14862 , n14863 , n14864 , n14865 , n14866 , n14867 , n14868 , n14869 , n14870 , n14871 , n14872 , n14873 , n14874 , n14875 , n14876 , n14877 , n14878 , n14879 , n14880 , n14881 , n14882 , n14883 , n14884 , n14885 , n14886 , n14887 , n14888 , n14889 , n14890 , n14891 , n14892 , n14893 , n14894 , n14895 , n14896 , n14897 , n14898 , n14899 , n14900 , n14901 , n14902 , n14903 , n14904 , n14905 , n14906 , n14907 , n14908 , n14909 , n14910 , n14911 , n14912 , n14913 , n14914 , n14915 , n14916 , n14917 , n14918 , n14919 , n14920 , n14921 , n14922 , n14923 , n14924 , n14925 , n14926 , n14927 , n14928 , n14929 , n14930 , n14931 , n14932 , n14933 , n14934 , n14935 , n14936 , n14937 , n14938 , n14939 , n14940 , n14941 , n14942 , n14943 , n14944 , n14945 , n14946 , n14947 , n14948 , n14949 , n14950 , n14951 , n14952 , n14953 , n14954 , n14955 , n14956 , n14957 , n14958 , n14959 , n14960 , n14961 , n14962 , n14963 , n14964 , n14965 , n14966 , n14967 , n14968 , n14969 , n14970 , n14971 , n14972 , n14973 , n14974 , n14975 , n14976 , n14977 , n14978 , n14979 , n14980 , n14981 , n14982 , n14983 , n14984 , n14985 , n14986 , n14987 , n14988 , n14989 , n14990 , n14991 , n14992 , n14993 , n14994 , n14995 , n14996 , n14997 , n14998 , n14999 , n15000 , n15001 , n15002 , n15003 , n15004 , n15005 , n15006 , n15007 , n15008 , n15009 , n15010 , n15011 , n15012 , n15013 , n15014 , n15015 , n15016 , n15017 , n15018 , n15019 , n15020 , n15021 , n15022 , n15023 , n15024 , n15025 , n15026 , n15027 , n15028 , n15029 , n15030 , n15031 , n15032 , n15033 , n15034 , n15035 , n15036 , n15037 , n15038 , n15039 , n15040 , n15041 , n15042 , n15043 , n15044 , n15045 , n15046 , n15047 , n15048 , n15049 , n15050 , n15051 , n15052 , n15053 , n15054 , n15055 , n15056 , n15057 , n15058 , n15059 , n15060 , n15061 , n15062 , n15063 , n15064 , n15065 , n15066 , n15067 , n15068 , n15069 , n15070 , n15071 , n15072 , n15073 , n15074 , n15075 , n15076 , n15077 , n15078 , n15079 , n15080 , n15081 , n15082 , n15083 , n15084 , n15085 , n15086 , n15087 , n15088 , n15089 , n15090 , n15091 , n15092 , n15093 , n15094 , n15095 , n15096 , n15097 , n15098 , n15099 , n15100 , n15101 , n15102 , n15103 , n15104 , n15105 , n15106 , n15107 , n15108 , n15109 , n15110 , n15111 , n15112 , n15113 , n15114 , n15115 , n15116 , n15117 , n15118 , n15119 , n15120 , n15121 , n15122 , n15123 , n15124 , n15125 , n15126 , n15127 , n15128 , n15129 , n15130 , n15131 , n15132 , n15133 , n15134 , n15135 , n15136 , n15137 , n15138 , n15139 , n15140 , n15141 , n15142 , n15143 , n15144 , n15145 , n15146 , n15147 , n15148 , n15149 , n15150 , n15151 , n15152 , n15153 , n15154 , n15155 , n15156 , n15157 , n15158 , n15159 , n15160 , n15161 , n15162 , n15163 , n15164 , n15165 , n15166 , n15167 , n15168 , n15169 , n15170 , n15171 , n15172 , n15173 , n15174 , n15175 , n15176 , n15177 , n15178 , n15179 , n15180 , n15181 , n15182 , n15183 , n15184 , n15185 , n15186 , n15187 , n15188 , n15189 , n15190 , n15191 , n15192 , n15193 , n15194 , n15195 , n15196 , n15197 , n15198 , n15199 , n15200 , n15201 , n15202 , n15203 , n15204 , n15205 , n15206 , n15207 , n15208 , n15209 , n15210 , n15211 , n15212 , n15213 , n15214 , n15215 , n15216 , n15217 , n15218 , n15219 , n15220 , n15221 , n15222 , n15223 , n15224 , n15225 , n15226 , n15227 , n15228 , n15229 , n15230 , n15231 , n15232 , n15233 , n15234 , n15235 , n15236 , n15237 , n15238 , n15239 , n15240 , n15241 , n15242 , n15243 , n15244 , n15245 , n15246 , n15247 , n15248 , n15249 , n15250 , n15251 , n15252 , n15253 , n15254 , n15255 , n15256 , n15257 , n15258 , n15259 , n15260 , n15261 , n15262 , n15263 , n15264 , n15265 , n15266 , n15267 , n15268 , n15269 , n15270 , n15271 , n15272 , n15273 , n15274 , n15275 , n15276 , n15277 , n15278 , n15279 , n15280 , n15281 , n15282 , n15283 , n15284 , n15285 , n15286 , n15287 , n15288 , n15289 , n15290 , n15291 , n15292 , n15293 , n15294 , n15295 , n15296 , n15297 , n15298 , n15299 , n15300 , n15301 , n15302 , n15303 , n15304 , n15305 , n15306 , n15307 , n15308 , n15309 , n15310 , n15311 , n15312 , n15313 , n15314 , n15315 , n15316 , n15317 , n15318 , n15319 , n15320 , n15321 , n15322 , n15323 , n15324 , n15325 , n15326 , n15327 , n15328 , n15329 , n15330 , n15331 , n15332 , n15333 , n15334 , n15335 , n15336 , n15337 , n15338 , n15339 , n15340 , n15341 , n15342 , n15343 , n15344 , n15345 , n15346 , n15347 , n15348 , n15349 , n15350 , n15351 , n15352 , n15353 , n15354 , n15355 , n15356 , n15357 , n15358 , n15359 , n15360 , n15361 , n15362 , n15363 , n15364 , n15365 , n15366 , n15367 , n15368 , n15369 , n15370 , n15371 , n15372 , n15373 , n15374 , n15375 , n15376 , n15377 , n15378 , n15379 , n15380 , n15381 , n15382 , n15383 , n15384 , n15385 , n15386 , n15387 , n15388 , n15389 , n15390 , n15391 , n15392 , n15393 , n15394 , n15395 , n15396 , n15397 , n15398 , n15399 , n15400 , n15401 , n15402 , n15403 , n15404 , n15405 , n15406 , n15407 , n15408 , n15409 , n15410 , n15411 , n15412 , n15413 , n15414 , n15415 , n15416 , n15417 , n15418 , n15419 , n15420 , n15421 , n15422 , n15423 , n15424 , n15425 , n15426 , n15427 , n15428 , n15429 , n15430 , n15431 , n15432 , n15433 , n15434 , n15435 , n15436 , n15437 , n15438 , n15439 , n15440 , n15441 , n15442 , n15443 , n15444 , n15445 , n15446 , n15447 , n15448 , n15449 , n15450 , n15451 , n15452 , n15453 , n15454 , n15455 , n15456 , n15457 , n15458 , n15459 , n15460 , n15461 , n15462 , n15463 , n15464 , n15465 , n15466 , n15467 , n15468 , n15469 , n15470 , n15471 , n15472 , n15473 , n15474 , n15475 , n15476 , n15477 , n15478 , n15479 , n15480 , n15481 , n15482 , n15483 , n15484 , n15485 , n15486 , n15487 , n15488 , n15489 , n15490 , n15491 , n15492 , n15493 , n15494 , n15495 , n15496 , n15497 , n15498 , n15499 , n15500 , n15501 , n15502 , n15503 , n15504 , n15505 , n15506 , n15507 , n15508 , n15509 , n15510 , n15511 , n15512 , n15513 , n15514 , n15515 , n15516 , n15517 , n15518 , n15519 , n15520 , n15521 , n15522 , n15523 , n15524 , n15525 , n15526 , n15527 , n15528 , n15529 , n15530 , n15531 , n15532 , n15533 , n15534 , n15535 , n15536 , n15537 , n15538 , n15539 , n15540 , n15541 , n15542 , n15543 , n15544 , n15545 , n15546 , n15547 , n15548 , n15549 , n15550 , n15551 , n15552 , n15553 , n15554 , n15555 , n15556 , n15557 , n15558 , n15559 , n15560 , n15561 , n15562 , n15563 , n15564 , n15565 , n15566 , n15567 , n15568 , n15569 , n15570 , n15571 , n15572 , n15573 , n15574 , n15575 , n15576 , n15577 , n15578 , n15579 , n15580 , n15581 , n15582 , n15583 , n15584 , n15585 , n15586 , n15587 , n15588 , n15589 , n15590 , n15591 , n15592 , n15593 , n15594 , n15595 , n15596 , n15597 , n15598 , n15599 , n15600 , n15601 , n15602 , n15603 , n15604 , n15605 , n15606 , n15607 , n15608 , n15609 , n15610 , n15611 , n15612 , n15613 , n15614 , n15615 , n15616 , n15617 , n15618 , n15619 , n15620 , n15621 , n15622 , n15623 , n15624 , n15625 , n15626 , n15627 , n15628 , n15629 , n15630 , n15631 , n15632 , n15633 , n15634 , n15635 , n15636 , n15637 , n15638 , n15639 , n15640 , n15641 , n15642 , n15643 , n15644 , n15645 , n15646 , n15647 , n15648 , n15649 , n15650 , n15651 , n15652 , n15653 , n15654 , n15655 , n15656 , n15657 , n15658 , n15659 , n15660 , n15661 , n15662 , n15663 , n15664 , n15665 , n15666 , n15667 , n15668 , n15669 , n15670 , n15671 , n15672 , n15673 , n15674 , n15675 , n15676 , n15677 , n15678 , n15679 , n15680 , n15681 , n15682 , n15683 , n15684 , n15685 , n15686 , n15687 , n15688 , n15689 , n15690 , n15691 , n15692 , n15693 , n15694 , n15695 , n15696 , n15697 , n15698 , n15699 , n15700 , n15701 , n15702 , n15703 , n15704 , n15705 , n15706 , n15707 , n15708 , n15709 , n15710 , n15711 , n15712 , n15713 , n15714 , n15715 , n15716 , n15717 , n15718 , n15719 , n15720 , n15721 , n15722 , n15723 , n15724 , n15725 , n15726 , n15727 , n15728 , n15729 , n15730 , n15731 , n15732 , n15733 , n15734 , n15735 , n15736 , n15737 , n15738 , n15739 , n15740 , n15741 , n15742 , n15743 , n15744 , n15745 , n15746 , n15747 , n15748 , n15749 , n15750 , n15751 , n15752 , n15753 , n15754 , n15755 , n15756 , n15757 , n15758 , n15759 , n15760 , n15761 , n15762 , n15763 , n15764 , n15765 , n15766 , n15767 , n15768 , n15769 , n15770 , n15771 , n15772 , n15773 , n15774 , n15775 , n15776 , n15777 , n15778 , n15779 , n15780 , n15781 , n15782 , n15783 , n15784 , n15785 , n15786 , n15787 , n15788 , n15789 , n15790 , n15791 , n15792 , n15793 , n15794 , n15795 , n15796 , n15797 , n15798 , n15799 , n15800 , n15801 , n15802 , n15803 , n15804 , n15805 , n15806 , n15807 , n15808 , n15809 , n15810 , n15811 , n15812 , n15813 , n15814 , n15815 , n15816 , n15817 , n15818 , n15819 , n15820 , n15821 , n15822 , n15823 , n15824 , n15825 , n15826 , n15827 , n15828 , n15829 , n15830 , n15831 , n15832 , n15833 , n15834 , n15835 , n15836 , n15837 , n15838 , n15839 , n15840 , n15841 , n15842 , n15843 , n15844 , n15845 , n15846 , n15847 , n15848 , n15849 , n15850 , n15851 , n15852 , n15853 , n15854 , n15855 , n15856 , n15857 , n15858 , n15859 , n15860 , n15861 , n15862 , n15863 , n15864 , n15865 , n15866 , n15867 , n15868 , n15869 , n15870 , n15871 , n15872 , n15873 , n15874 , n15875 , n15876 , n15877 , n15878 , n15879 , n15880 , n15881 , n15882 , n15883 , n15884 , n15885 , n15886 , n15887 , n15888 , n15889 , n15890 , n15891 , n15892 , n15893 , n15894 , n15895 , n15896 , n15897 , n15898 , n15899 , n15900 , n15901 , n15902 , n15903 , n15904 , n15905 , n15906 , n15907 , n15908 , n15909 , n15910 , n15911 , n15912 , n15913 , n15914 , n15915 , n15916 , n15917 , n15918 , n15919 , n15920 , n15921 , n15922 , n15923 , n15924 , n15925 , n15926 , n15927 , n15928 , n15929 , n15930 , n15931 , n15932 , n15933 , n15934 , n15935 , n15936 , n15937 , n15938 , n15939 , n15940 , n15941 , n15942 , n15943 , n15944 , n15945 , n15946 , n15947 , n15948 , n15949 , n15950 , n15951 , n15952 , n15953 , n15954 , n15955 , n15956 , n15957 , n15958 , n15959 , n15960 , n15961 , n15962 , n15963 , n15964 , n15965 , n15966 , n15967 , n15968 , n15969 , n15970 , n15971 , n15972 , n15973 , n15974 , n15975 , n15976 , n15977 , n15978 , n15979 , n15980 , n15981 , n15982 , n15983 , n15984 , n15985 , n15986 , n15987 , n15988 , n15989 , n15990 , n15991 , n15992 , n15993 , n15994 , n15995 , n15996 , n15997 , n15998 , n15999 , n16000 , n16001 , n16002 , n16003 , n16004 , n16005 , n16006 , n16007 , n16008 , n16009 , n16010 , n16011 , n16012 , n16013 , n16014 , n16015 , n16016 , n16017 , n16018 , n16019 , n16020 , n16021 , n16022 , n16023 , n16024 , n16025 , n16026 , n16027 , n16028 , n16029 , n16030 , n16031 , n16032 , n16033 , n16034 , n16035 , n16036 , n16037 , n16038 , n16039 , n16040 , n16041 , n16042 , n16043 , n16044 , n16045 , n16046 , n16047 , n16048 , n16049 , n16050 , n16051 , n16052 , n16053 , n16054 , n16055 , n16056 , n16057 , n16058 , n16059 , n16060 , n16061 , n16062 , n16063 , n16064 , n16065 , n16066 , n16067 , n16068 , n16069 , n16070 , n16071 , n16072 , n16073 , n16074 , n16075 , n16076 , n16077 , n16078 , n16079 , n16080 , n16081 , n16082 , n16083 , n16084 , n16085 , n16086 , n16087 , n16088 , n16089 , n16090 , n16091 , n16092 , n16093 , n16094 , n16095 , n16096 , n16097 , n16098 , n16099 , n16100 , n16101 , n16102 , n16103 , n16104 , n16105 , n16106 , n16107 , n16108 , n16109 , n16110 , n16111 , n16112 , n16113 , n16114 , n16115 , n16116 , n16117 , n16118 , n16119 , n16120 , n16121 , n16122 , n16123 , n16124 , n16125 , n16126 , n16127 , n16128 , n16129 , n16130 , n16131 , n16132 , n16133 , n16134 , n16135 , n16136 , n16137 , n16138 , n16139 , n16140 , n16141 , n16142 , n16143 , n16144 , n16145 , n16146 , n16147 , n16148 , n16149 , n16150 , n16151 , n16152 , n16153 , n16154 , n16155 , n16156 , n16157 , n16158 , n16159 , n16160 , n16161 , n16162 , n16163 , n16164 , n16165 , n16166 , n16167 , n16168 , n16169 , n16170 , n16171 , n16172 , n16173 , n16174 , n16175 , n16176 , n16177 , n16178 , n16179 , n16180 , n16181 , n16182 , n16183 , n16184 , n16185 , n16186 , n16187 , n16188 , n16189 , n16190 , n16191 , n16192 , n16193 , n16194 , n16195 , n16196 , n16197 , n16198 , n16199 , n16200 , n16201 , n16202 , n16203 , n16204 , n16205 , n16206 , n16207 , n16208 , n16209 , n16210 , n16211 , n16212 , n16213 , n16214 , n16215 , n16216 , n16217 , n16218 , n16219 , n16220 , n16221 , n16222 , n16223 , n16224 , n16225 , n16226 , n16227 , n16228 , n16229 , n16230 , n16231 , n16232 , n16233 , n16234 , n16235 , n16236 , n16237 , n16238 , n16239 , n16240 , n16241 , n16242 , n16243 , n16244 , n16245 , n16246 , n16247 , n16248 , n16249 , n16250 , n16251 , n16252 , n16253 , n16254 , n16255 , n16256 , n16257 , n16258 , n16259 , n16260 , n16261 , n16262 , n16263 , n16264 , n16265 , n16266 , n16267 , n16268 , n16269 , n16270 , n16271 , n16272 , n16273 , n16274 , n16275 , n16276 , n16277 , n16278 , n16279 , n16280 , n16281 , n16282 , n16283 , n16284 , n16285 , n16286 , n16287 , n16288 , n16289 , n16290 , n16291 , n16292 , n16293 , n16294 , n16295 , n16296 , n16297 , n16298 , n16299 , n16300 , n16301 , n16302 , n16303 , n16304 , n16305 , n16306 , n16307 , n16308 , n16309 , n16310 , n16311 , n16312 , n16313 , n16314 , n16315 , n16316 , n16317 , n16318 , n16319 , n16320 , n16321 , n16322 , n16323 , n16324 , n16325 , n16326 , n16327 , n16328 , n16329 , n16330 , n16331 , n16332 , n16333 , n16334 , n16335 , n16336 , n16337 , n16338 , n16339 , n16340 , n16341 , n16342 , n16343 , n16344 , n16345 , n16346 , n16347 , n16348 , n16349 , n16350 , n16351 , n16352 , n16353 , n16354 , n16355 , n16356 , n16357 , n16358 , n16359 , n16360 , n16361 , n16362 , n16363 , n16364 , n16365 , n16366 , n16367 , n16368 , n16369 , n16370 , n16371 , n16372 , n16373 , n16374 , n16375 , n16376 , n16377 , n16378 , n16379 , n16380 , n16381 , n16382 , n16383 , n16384 , n16385 , n16386 , n16387 , n16388 , n16389 , n16390 , n16391 , n16392 , n16393 , n16394 , n16395 , n16396 , n16397 , n16398 , n16399 , n16400 , n16401 , n16402 , n16403 , n16404 , n16405 , n16406 , n16407 , n16408 , n16409 , n16410 , n16411 , n16412 , n16413 , n16414 , n16415 , n16416 , n16417 , n16418 , n16419 , n16420 , n16421 , n16422 , n16423 , n16424 , n16425 , n16426 , n16427 , n16428 , n16429 , n16430 , n16431 , n16432 , n16433 , n16434 , n16435 , n16436 , n16437 , n16438 , n16439 , n16440 , n16441 , n16442 , n16443 , n16444 , n16445 , n16446 , n16447 , n16448 , n16449 , n16450 , n16451 , n16452 , n16453 , n16454 , n16455 , n16456 , n16457 , n16458 , n16459 , n16460 , n16461 , n16462 , n16463 , n16464 , n16465 , n16466 , n16467 , n16468 , n16469 , n16470 , n16471 , n16472 , n16473 , n16474 , n16475 , n16476 , n16477 , n16478 , n16479 , n16480 , n16481 , n16482 , n16483 , n16484 , n16485 , n16486 , n16487 , n16488 , n16489 , n16490 , n16491 , n16492 , n16493 , n16494 , n16495 , n16496 , n16497 , n16498 , n16499 , n16500 , n16501 , n16502 , n16503 , n16504 , n16505 , n16506 , n16507 , n16508 , n16509 , n16510 , n16511 , n16512 , n16513 , n16514 , n16515 , n16516 , n16517 , n16518 , n16519 , n16520 , n16521 , n16522 , n16523 , n16524 , n16525 , n16526 , n16527 , n16528 , n16529 , n16530 , n16531 , n16532 , n16533 , n16534 , n16535 , n16536 , n16537 , n16538 , n16539 , n16540 , n16541 , n16542 , n16543 , n16544 , n16545 , n16546 , n16547 , n16548 , n16549 , n16550 , n16551 , n16552 , n16553 , n16554 , n16555 , n16556 , n16557 , n16558 , n16559 , n16560 , n16561 , n16562 , n16563 , n16564 , n16565 , n16566 , n16567 , n16568 , n16569 , n16570 , n16571 , n16572 , n16573 , n16574 , n16575 , n16576 , n16577 , n16578 , n16579 , n16580 , n16581 , n16582 , n16583 , n16584 , n16585 , n16586 , n16587 , n16588 , n16589 , n16590 , n16591 , n16592 , n16593 , n16594 , n16595 , n16596 , n16597 , n16598 , n16599 , n16600 , n16601 , n16602 , n16603 , n16604 , n16605 , n16606 , n16607 , n16608 , n16609 , n16610 , n16611 , n16612 , n16613 , n16614 , n16615 , n16616 , n16617 , n16618 , n16619 , n16620 , n16621 , n16622 , n16623 , n16624 , n16625 , n16626 , n16627 , n16628 , n16629 , n16630 , n16631 , n16632 , n16633 , n16634 , n16635 , n16636 , n16637 , n16638 , n16639 , n16640 , n16641 , n16642 , n16643 , n16644 , n16645 , n16646 , n16647 , n16648 , n16649 , n16650 , n16651 , n16652 , n16653 , n16654 , n16655 , n16656 , n16657 , n16658 , n16659 , n16660 , n16661 , n16662 , n16663 , n16664 , n16665 , n16666 , n16667 , n16668 , n16669 , n16670 , n16671 , n16672 , n16673 , n16674 , n16675 , n16676 , n16677 , n16678 , n16679 , n16680 , n16681 , n16682 , n16683 , n16684 , n16685 , n16686 , n16687 , n16688 , n16689 , n16690 , n16691 , n16692 , n16693 , n16694 , n16695 , n16696 , n16697 , n16698 , n16699 , n16700 , n16701 , n16702 , n16703 , n16704 , n16705 , n16706 , n16707 , n16708 , n16709 , n16710 , n16711 , n16712 , n16713 , n16714 , n16715 , n16716 , n16717 , n16718 , n16719 , n16720 , n16721 , n16722 , n16723 , n16724 , n16725 , n16726 , n16727 , n16728 , n16729 , n16730 , n16731 , n16732 , n16733 , n16734 , n16735 , n16736 , n16737 , n16738 , n16739 , n16740 , n16741 , n16742 , n16743 , n16744 , n16745 , n16746 , n16747 , n16748 , n16749 , n16750 , n16751 , n16752 , n16753 , n16754 , n16755 , n16756 , n16757 , n16758 , n16759 , n16760 , n16761 , n16762 , n16763 , n16764 , n16765 , n16766 , n16767 , n16768 , n16769 , n16770 , n16771 , n16772 , n16773 , n16774 , n16775 , n16776 , n16777 , n16778 , n16779 , n16780 , n16781 , n16782 , n16783 , n16784 , n16785 , n16786 , n16787 , n16788 , n16789 , n16790 , n16791 , n16792 , n16793 , n16794 , n16795 , n16796 , n16797 , n16798 , n16799 , n16800 , n16801 , n16802 , n16803 , n16804 , n16805 , n16806 , n16807 , n16808 , n16809 , n16810 , n16811 , n16812 , n16813 , n16814 , n16815 , n16816 , n16817 , n16818 , n16819 , n16820 , n16821 , n16822 , n16823 , n16824 , n16825 , n16826 , n16827 , n16828 , n16829 , n16830 , n16831 , n16832 , n16833 , n16834 , n16835 , n16836 , n16837 , n16838 , n16839 , n16840 , n16841 , n16842 , n16843 , n16844 , n16845 , n16846 , n16847 , n16848 , n16849 , n16850 , n16851 , n16852 , n16853 , n16854 , n16855 , n16856 , n16857 , n16858 , n16859 , n16860 , n16861 , n16862 , n16863 , n16864 , n16865 , n16866 , n16867 , n16868 , n16869 , n16870 , n16871 , n16872 , n16873 , n16874 , n16875 , n16876 , n16877 , n16878 , n16879 , n16880 , n16881 , n16882 , n16883 , n16884 , n16885 , n16886 , n16887 , n16888 , n16889 , n16890 , n16891 , n16892 , n16893 , n16894 , n16895 , n16896 , n16897 , n16898 , n16899 , n16900 , n16901 , n16902 , n16903 , n16904 , n16905 , n16906 , n16907 , n16908 , n16909 , n16910 , n16911 , n16912 , n16913 , n16914 , n16915 , n16916 , n16917 , n16918 , n16919 , n16920 , n16921 , n16922 , n16923 , n16924 , n16925 , n16926 , n16927 , n16928 , n16929 , n16930 , n16931 , n16932 , n16933 , n16934 , n16935 , n16936 , n16937 , n16938 , n16939 , n16940 , n16941 , n16942 , n16943 , n16944 , n16945 , n16946 , n16947 , n16948 , n16949 , n16950 , n16951 , n16952 , n16953 , n16954 , n16955 , n16956 , n16957 , n16958 , n16959 , n16960 , n16961 , n16962 , n16963 , n16964 , n16965 , n16966 , n16967 , n16968 , n16969 , n16970 , n16971 , n16972 , n16973 , n16974 , n16975 , n16976 , n16977 , n16978 , n16979 , n16980 , n16981 , n16982 , n16983 , n16984 , n16985 , n16986 , n16987 , n16988 , n16989 , n16990 , n16991 , n16992 , n16993 , n16994 , n16995 , n16996 , n16997 , n16998 , n16999 , n17000 , n17001 , n17002 , n17003 , n17004 , n17005 , n17006 , n17007 , n17008 , n17009 , n17010 , n17011 , n17012 , n17013 , n17014 , n17015 , n17016 , n17017 , n17018 , n17019 , n17020 , n17021 , n17022 , n17023 , n17024 , n17025 , n17026 , n17027 , n17028 , n17029 , n17030 , n17031 , n17032 , n17033 , n17034 , n17035 , n17036 , n17037 , n17038 , n17039 , n17040 , n17041 , n17042 , n17043 , n17044 , n17045 , n17046 , n17047 , n17048 , n17049 , n17050 , n17051 , n17052 , n17053 , n17054 , n17055 , n17056 , n17057 , n17058 , n17059 , n17060 , n17061 , n17062 , n17063 , n17064 , n17065 , n17066 , n17067 , n17068 , n17069 , n17070 , n17071 , n17072 , n17073 , n17074 , n17075 , n17076 , n17077 , n17078 , n17079 , n17080 , n17081 , n17082 , n17083 , n17084 , n17085 , n17086 , n17087 , n17088 , n17089 , n17090 , n17091 , n17092 , n17093 , n17094 , n17095 , n17096 , n17097 , n17098 , n17099 , n17100 , n17101 , n17102 , n17103 , n17104 , n17105 , n17106 , n17107 , n17108 , n17109 , n17110 , n17111 , n17112 , n17113 , n17114 , n17115 , n17116 , n17117 , n17118 , n17119 , n17120 , n17121 , n17122 , n17123 , n17124 , n17125 , n17126 , n17127 , n17128 , n17129 , n17130 , n17131 , n17132 , n17133 , n17134 , n17135 , n17136 , n17137 , n17138 , n17139 , n17140 , n17141 , n17142 , n17143 , n17144 , n17145 , n17146 , n17147 , n17148 , n17149 , n17150 , n17151 , n17152 , n17153 , n17154 , n17155 , n17156 , n17157 , n17158 , n17159 , n17160 , n17161 , n17162 , n17163 , n17164 , n17165 , n17166 , n17167 , n17168 , n17169 , n17170 , n17171 , n17172 , n17173 , n17174 , n17175 , n17176 , n17177 , n17178 , n17179 , n17180 , n17181 , n17182 , n17183 , n17184 , n17185 , n17186 , n17187 , n17188 , n17189 , n17190 , n17191 , n17192 , n17193 , n17194 , n17195 , n17196 , n17197 , n17198 , n17199 , n17200 , n17201 , n17202 , n17203 , n17204 , n17205 , n17206 , n17207 , n17208 , n17209 , n17210 , n17211 , n17212 , n17213 , n17214 , n17215 , n17216 , n17217 , n17218 , n17219 , n17220 , n17221 , n17222 , n17223 , n17224 , n17225 , n17226 , n17227 , n17228 , n17229 , n17230 , n17231 , n17232 , n17233 , n17234 , n17235 , n17236 , n17237 , n17238 , n17239 , n17240 , n17241 , n17242 , n17243 , n17244 , n17245 , n17246 , n17247 , n17248 , n17249 , n17250 , n17251 , n17252 , n17253 , n17254 , n17255 , n17256 , n17257 , n17258 , n17259 , n17260 , n17261 , n17262 , n17263 , n17264 , n17265 , n17266 , n17267 , n17268 , n17269 , n17270 , n17271 , n17272 , n17273 , n17274 , n17275 , n17276 , n17277 , n17278 , n17279 , n17280 , n17281 , n17282 , n17283 , n17284 , n17285 , n17286 , n17287 , n17288 , n17289 , n17290 , n17291 , n17292 , n17293 , n17294 , n17295 , n17296 , n17297 , n17298 , n17299 , n17300 , n17301 , n17302 , n17303 , n17304 , n17305 , n17306 , n17307 , n17308 , n17309 , n17310 , n17311 , n17312 , n17313 , n17314 , n17315 , n17316 , n17317 , n17318 , n17319 , n17320 , n17321 , n17322 , n17323 , n17324 , n17325 , n17326 , n17327 , n17328 , n17329 , n17330 , n17331 , n17332 , n17333 , n17334 , n17335 , n17336 , n17337 , n17338 , n17339 , n17340 , n17341 , n17342 , n17343 , n17344 , n17345 , n17346 , n17347 , n17348 , n17349 , n17350 , n17351 , n17352 , n17353 , n17354 , n17355 , n17356 , n17357 , n17358 , n17359 , n17360 , n17361 , n17362 , n17363 , n17364 , n17365 , n17366 , n17367 , n17368 , n17369 , n17370 , n17371 , n17372 , n17373 , n17374 , n17375 , n17376 , n17377 , n17378 , n17379 , n17380 , n17381 , n17382 , n17383 , n17384 , n17385 , n17386 , n17387 , n17388 , n17389 , n17390 , n17391 , n17392 , n17393 , n17394 , n17395 , n17396 , n17397 , n17398 , n17399 , n17400 , n17401 , n17402 , n17403 , n17404 , n17405 , n17406 , n17407 , n17408 , n17409 , n17410 , n17411 , n17412 , n17413 , n17414 , n17415 , n17416 , n17417 , n17418 , n17419 , n17420 , n17421 , n17422 , n17423 , n17424 , n17425 , n17426 , n17427 , n17428 , n17429 , n17430 , n17431 , n17432 , n17433 , n17434 , n17435 , n17436 , n17437 , n17438 , n17439 , n17440 , n17441 , n17442 , n17443 , n17444 , n17445 , n17446 , n17447 , n17448 , n17449 , n17450 , n17451 , n17452 , n17453 , n17454 , n17455 , n17456 , n17457 , n17458 , n17459 , n17460 , n17461 , n17462 , n17463 , n17464 , n17465 , n17466 , n17467 , n17468 , n17469 , n17470 , n17471 , n17472 , n17473 , n17474 , n17475 , n17476 , n17477 , n17478 , n17479 , n17480 , n17481 , n17482 , n17483 , n17484 , n17485 , n17486 , n17487 , n17488 , n17489 , n17490 , n17491 , n17492 , n17493 , n17494 , n17495 , n17496 , n17497 , n17498 , n17499 , n17500 , n17501 , n17502 , n17503 , n17504 , n17505 , n17506 , n17507 , n17508 , n17509 , n17510 , n17511 , n17512 , n17513 , n17514 , n17515 , n17516 , n17517 , n17518 , n17519 , n17520 , n17521 , n17522 , n17523 , n17524 , n17525 , n17526 , n17527 , n17528 , n17529 , n17530 , n17531 , n17532 , n17533 , n17534 , n17535 , n17536 , n17537 , n17538 , n17539 , n17540 , n17541 , n17542 , n17543 , n17544 , n17545 , n17546 , n17547 , n17548 , n17549 , n17550 , n17551 , n17552 , n17553 , n17554 , n17555 , n17556 , n17557 , n17558 , n17559 , n17560 , n17561 , n17562 , n17563 , n17564 , n17565 , n17566 , n17567 , n17568 , n17569 , n17570 , n17571 , n17572 , n17573 , n17574 , n17575 , n17576 , n17577 , n17578 , n17579 , n17580 , n17581 , n17582 , n17583 , n17584 , n17585 , n17586 , n17587 , n17588 , n17589 , n17590 , n17591 , n17592 , n17593 , n17594 , n17595 , n17596 , n17597 , n17598 , n17599 , n17600 , n17601 , n17602 , n17603 , n17604 , n17605 , n17606 , n17607 , n17608 , n17609 , n17610 , n17611 , n17612 , n17613 , n17614 , n17615 , n17616 , n17617 , n17618 , n17619 , n17620 , n17621 , n17622 , n17623 , n17624 , n17625 , n17626 , n17627 , n17628 , n17629 , n17630 , n17631 , n17632 , n17633 , n17634 , n17635 , n17636 , n17637 , n17638 , n17639 , n17640 , n17641 , n17642 , n17643 , n17644 , n17645 , n17646 , n17647 , n17648 , n17649 , n17650 , n17651 , n17652 , n17653 , n17654 , n17655 , n17656 , n17657 , n17658 , n17659 , n17660 , n17661 , n17662 , n17663 , n17664 , n17665 , n17666 , n17667 , n17668 , n17669 , n17670 , n17671 , n17672 , n17673 , n17674 , n17675 , n17676 , n17677 , n17678 , n17679 , n17680 , n17681 , n17682 , n17683 , n17684 , n17685 , n17686 , n17687 , n17688 , n17689 , n17690 , n17691 , n17692 , n17693 , n17694 , n17695 , n17696 , n17697 , n17698 , n17699 , n17700 , n17701 , n17702 , n17703 , n17704 , n17705 , n17706 , n17707 , n17708 , n17709 , n17710 , n17711 , n17712 , n17713 , n17714 , n17715 , n17716 , n17717 , n17718 , n17719 , n17720 , n17721 , n17722 , n17723 , n17724 , n17725 , n17726 , n17727 , n17728 , n17729 , n17730 , n17731 , n17732 , n17733 , n17734 , n17735 , n17736 , n17737 , n17738 , n17739 , n17740 , n17741 , n17742 , n17743 , n17744 , n17745 , n17746 , n17747 , n17748 , n17749 , n17750 , n17751 , n17752 , n17753 , n17754 , n17755 , n17756 , n17757 , n17758 , n17759 , n17760 , n17761 , n17762 , n17763 , n17764 , n17765 , n17766 , n17767 , n17768 , n17769 , n17770 , n17771 , n17772 , n17773 , n17774 , n17775 , n17776 , n17777 , n17778 , n17779 , n17780 , n17781 , n17782 , n17783 , n17784 , n17785 , n17786 , n17787 , n17788 , n17789 , n17790 , n17791 , n17792 , n17793 , n17794 , n17795 , n17796 , n17797 , n17798 , n17799 , n17800 , n17801 , n17802 , n17803 , n17804 , n17805 , n17806 , n17807 , n17808 , n17809 , n17810 , n17811 , n17812 , n17813 , n17814 , n17815 , n17816 , n17817 , n17818 , n17819 , n17820 , n17821 , n17822 , n17823 , n17824 , n17825 , n17826 , n17827 , n17828 , n17829 , n17830 , n17831 , n17832 , n17833 , n17834 , n17835 , n17836 , n17837 , n17838 , n17839 , n17840 , n17841 , n17842 , n17843 , n17844 , n17845 , n17846 , n17847 , n17848 , n17849 , n17850 , n17851 , n17852 , n17853 , n17854 , n17855 , n17856 , n17857 , n17858 , n17859 , n17860 , n17861 , n17862 , n17863 , n17864 , n17865 , n17866 , n17867 , n17868 , n17869 , n17870 , n17871 , n17872 , n17873 , n17874 , n17875 , n17876 , n17877 , n17878 , n17879 , n17880 , n17881 , n17882 , n17883 , n17884 , n17885 , n17886 , n17887 , n17888 , n17889 , n17890 , n17891 , n17892 , n17893 , n17894 , n17895 , n17896 , n17897 , n17898 , n17899 , n17900 , n17901 , n17902 , n17903 , n17904 , n17905 , n17906 , n17907 , n17908 , n17909 , n17910 , n17911 , n17912 , n17913 , n17914 , n17915 , n17916 , n17917 , n17918 , n17919 , n17920 , n17921 , n17922 , n17923 , n17924 , n17925 , n17926 , n17927 , n17928 , n17929 , n17930 , n17931 , n17932 , n17933 , n17934 , n17935 , n17936 , n17937 , n17938 , n17939 , n17940 , n17941 , n17942 , n17943 , n17944 , n17945 , n17946 , n17947 , n17948 , n17949 , n17950 , n17951 , n17952 , n17953 , n17954 , n17955 , n17956 , n17957 , n17958 , n17959 , n17960 , n17961 , n17962 , n17963 , n17964 , n17965 , n17966 , n17967 , n17968 , n17969 , n17970 , n17971 , n17972 , n17973 , n17974 , n17975 , n17976 , n17977 , n17978 , n17979 , n17980 , n17981 , n17982 , n17983 , n17984 , n17985 , n17986 , n17987 , n17988 , n17989 , n17990 , n17991 , n17992 , n17993 , n17994 , n17995 , n17996 , n17997 , n17998 , n17999 , n18000 , n18001 , n18002 , n18003 , n18004 , n18005 , n18006 , n18007 , n18008 , n18009 , n18010 , n18011 , n18012 , n18013 , n18014 , n18015 , n18016 , n18017 , n18018 , n18019 , n18020 , n18021 , n18022 , n18023 , n18024 , n18025 , n18026 , n18027 , n18028 , n18029 , n18030 , n18031 , n18032 , n18033 , n18034 , n18035 , n18036 , n18037 , n18038 , n18039 , n18040 , n18041 , n18042 , n18043 , n18044 , n18045 , n18046 , n18047 , n18048 , n18049 , n18050 , n18051 , n18052 , n18053 , n18054 , n18055 , n18056 , n18057 , n18058 , n18059 , n18060 , n18061 , n18062 , n18063 , n18064 , n18065 , n18066 , n18067 , n18068 , n18069 , n18070 , n18071 , n18072 , n18073 , n18074 , n18075 , n18076 , n18077 , n18078 , n18079 , n18080 , n18081 , n18082 , n18083 , n18084 , n18085 , n18086 , n18087 , n18088 , n18089 , n18090 , n18091 , n18092 , n18093 , n18094 , n18095 , n18096 , n18097 , n18098 , n18099 , n18100 , n18101 , n18102 , n18103 , n18104 , n18105 , n18106 , n18107 , n18108 , n18109 , n18110 , n18111 , n18112 , n18113 , n18114 , n18115 , n18116 , n18117 , n18118 , n18119 , n18120 , n18121 , n18122 , n18123 , n18124 , n18125 , n18126 , n18127 , n18128 , n18129 , n18130 , n18131 , n18132 , n18133 , n18134 , n18135 , n18136 , n18137 , n18138 , n18139 , n18140 , n18141 , n18142 , n18143 , n18144 , n18145 , n18146 , n18147 , n18148 , n18149 , n18150 , n18151 , n18152 , n18153 , n18154 , n18155 , n18156 , n18157 , n18158 , n18159 , n18160 , n18161 , n18162 , n18163 , n18164 , n18165 , n18166 , n18167 , n18168 , n18169 , n18170 , n18171 , n18172 , n18173 , n18174 , n18175 , n18176 , n18177 , n18178 , n18179 , n18180 , n18181 , n18182 , n18183 , n18184 , n18185 , n18186 , n18187 , n18188 , n18189 , n18190 , n18191 , n18192 , n18193 , n18194 , n18195 , n18196 , n18197 , n18198 , n18199 , n18200 , n18201 , n18202 , n18203 , n18204 , n18205 , n18206 , n18207 , n18208 , n18209 , n18210 , n18211 , n18212 , n18213 , n18214 , n18215 , n18216 , n18217 , n18218 , n18219 , n18220 , n18221 , n18222 , n18223 , n18224 , n18225 , n18226 , n18227 , n18228 , n18229 , n18230 , n18231 , n18232 , n18233 , n18234 , n18235 , n18236 , n18237 , n18238 , n18239 , n18240 , n18241 , n18242 , n18243 , n18244 , n18245 , n18246 , n18247 , n18248 , n18249 , n18250 , n18251 , n18252 , n18253 , n18254 , n18255 , n18256 , n18257 , n18258 , n18259 , n18260 , n18261 , n18262 , n18263 , n18264 , n18265 , n18266 , n18267 , n18268 , n18269 , n18270 , n18271 , n18272 , n18273 , n18274 , n18275 , n18276 , n18277 , n18278 , n18279 , n18280 , n18281 , n18282 , n18283 , n18284 , n18285 , n18286 , n18287 , n18288 , n18289 , n18290 , n18291 , n18292 , n18293 , n18294 , n18295 , n18296 , n18297 , n18298 , n18299 , n18300 , n18301 , n18302 , n18303 , n18304 , n18305 , n18306 , n18307 , n18308 , n18309 , n18310 , n18311 , n18312 , n18313 , n18314 , n18315 , n18316 , n18317 , n18318 , n18319 , n18320 , n18321 , n18322 , n18323 , n18324 , n18325 , n18326 , n18327 , n18328 , n18329 , n18330 , n18331 , n18332 , n18333 , n18334 , n18335 , n18336 , n18337 , n18338 , n18339 , n18340 , n18341 , n18342 , n18343 , n18344 , n18345 , n18346 , n18347 , n18348 , n18349 , n18350 , n18351 , n18352 , n18353 , n18354 , n18355 , n18356 , n18357 , n18358 , n18359 , n18360 , n18361 , n18362 , n18363 , n18364 , n18365 , n18366 , n18367 , n18368 , n18369 , n18370 , n18371 , n18372 , n18373 , n18374 , n18375 , n18376 , n18377 , n18378 , n18379 , n18380 , n18381 , n18382 , n18383 , n18384 , n18385 , n18386 , n18387 , n18388 , n18389 , n18390 , n18391 , n18392 , n18393 , n18394 , n18395 , n18396 , n18397 , n18398 , n18399 , n18400 , n18401 , n18402 , n18403 , n18404 , n18405 , n18406 , n18407 , n18408 , n18409 , n18410 , n18411 , n18412 , n18413 , n18414 , n18415 , n18416 , n18417 , n18418 , n18419 , n18420 , n18421 , n18422 , n18423 , n18424 , n18425 , n18426 , n18427 , n18428 , n18429 , n18430 , n18431 , n18432 , n18433 , n18434 , n18435 , n18436 , n18437 , n18438 , n18439 , n18440 , n18441 , n18442 , n18443 , n18444 , n18445 , n18446 , n18447 , n18448 , n18449 , n18450 , n18451 , n18452 , n18453 , n18454 , n18455 , n18456 , n18457 , n18458 , n18459 , n18460 , n18461 , n18462 , n18463 , n18464 , n18465 , n18466 , n18467 , n18468 , n18469 , n18470 , n18471 , n18472 , n18473 , n18474 , n18475 , n18476 , n18477 , n18478 , n18479 , n18480 , n18481 , n18482 , n18483 , n18484 , n18485 , n18486 , n18487 , n18488 , n18489 , n18490 , n18491 , n18492 , n18493 , n18494 , n18495 , n18496 , n18497 , n18498 , n18499 , n18500 , n18501 , n18502 , n18503 , n18504 , n18505 , n18506 , n18507 , n18508 , n18509 , n18510 , n18511 , n18512 , n18513 , n18514 , n18515 , n18516 , n18517 , n18518 , n18519 , n18520 , n18521 , n18522 , n18523 , n18524 , n18525 , n18526 , n18527 , n18528 , n18529 , n18530 , n18531 , n18532 , n18533 , n18534 , n18535 , n18536 , n18537 , n18538 , n18539 , n18540 , n18541 , n18542 , n18543 , n18544 , n18545 , n18546 , n18547 , n18548 , n18549 , n18550 , n18551 , n18552 , n18553 , n18554 , n18555 , n18556 , n18557 , n18558 , n18559 , n18560 , n18561 , n18562 , n18563 , n18564 , n18565 , n18566 , n18567 , n18568 , n18569 , n18570 , n18571 , n18572 , n18573 , n18574 , n18575 , n18576 , n18577 , n18578 , n18579 , n18580 , n18581 , n18582 , n18583 , n18584 , n18585 , n18586 , n18587 , n18588 , n18589 , n18590 , n18591 , n18592 , n18593 , n18594 , n18595 , n18596 , n18597 , n18598 , n18599 , n18600 , n18601 , n18602 , n18603 , n18604 , n18605 , n18606 , n18607 , n18608 , n18609 , n18610 , n18611 , n18612 , n18613 , n18614 , n18615 , n18616 , n18617 , n18618 , n18619 , n18620 , n18621 , n18622 , n18623 , n18624 , n18625 , n18626 , n18627 , n18628 , n18629 , n18630 , n18631 , n18632 , n18633 , n18634 , n18635 , n18636 , n18637 , n18638 , n18639 , n18640 , n18641 , n18642 , n18643 , n18644 , n18645 , n18646 , n18647 , n18648 , n18649 , n18650 , n18651 , n18652 , n18653 , n18654 , n18655 , n18656 , n18657 , n18658 , n18659 , n18660 , n18661 , n18662 , n18663 , n18664 , n18665 , n18666 , n18667 , n18668 , n18669 , n18670 , n18671 , n18672 , n18673 , n18674 , n18675 , n18676 , n18677 , n18678 , n18679 , n18680 , n18681 , n18682 , n18683 , n18684 , n18685 , n18686 , n18687 , n18688 , n18689 , n18690 , n18691 , n18692 , n18693 , n18694 , n18695 , n18696 , n18697 , n18698 , n18699 , n18700 , n18701 , n18702 , n18703 , n18704 , n18705 , n18706 , n18707 , n18708 , n18709 , n18710 , n18711 , n18712 , n18713 , n18714 , n18715 , n18716 , n18717 , n18718 , n18719 , n18720 , n18721 , n18722 , n18723 , n18724 , n18725 , n18726 , n18727 , n18728 , n18729 , n18730 , n18731 , n18732 , n18733 , n18734 , n18735 , n18736 , n18737 , n18738 , n18739 , n18740 , n18741 , n18742 , n18743 , n18744 , n18745 , n18746 , n18747 , n18748 , n18749 , n18750 , n18751 , n18752 , n18753 , n18754 , n18755 , n18756 , n18757 , n18758 , n18759 , n18760 , n18761 , n18762 , n18763 , n18764 , n18765 , n18766 , n18767 , n18768 , n18769 , n18770 , n18771 , n18772 , n18773 , n18774 , n18775 , n18776 , n18777 , n18778 , n18779 , n18780 , n18781 , n18782 , n18783 , n18784 , n18785 , n18786 , n18787 , n18788 , n18789 , n18790 , n18791 , n18792 , n18793 , n18794 , n18795 , n18796 , n18797 , n18798 , n18799 , n18800 , n18801 , n18802 , n18803 , n18804 , n18805 , n18806 , n18807 , n18808 , n18809 , n18810 , n18811 , n18812 , n18813 , n18814 , n18815 , n18816 , n18817 , n18818 , n18819 , n18820 , n18821 , n18822 , n18823 , n18824 , n18825 , n18826 , n18827 , n18828 , n18829 , n18830 , n18831 , n18832 , n18833 , n18834 , n18835 , n18836 , n18837 , n18838 , n18839 , n18840 , n18841 , n18842 , n18843 , n18844 , n18845 , n18846 , n18847 , n18848 , n18849 , n18850 , n18851 , n18852 , n18853 , n18854 , n18855 , n18856 , n18857 , n18858 , n18859 , n18860 , n18861 , n18862 , n18863 , n18864 , n18865 , n18866 , n18867 , n18868 , n18869 , n18870 , n18871 , n18872 , n18873 , n18874 , n18875 , n18876 , n18877 , n18878 , n18879 , n18880 , n18881 , n18882 , n18883 , n18884 , n18885 , n18886 , n18887 , n18888 , n18889 , n18890 , n18891 , n18892 , n18893 , n18894 , n18895 , n18896 , n18897 , n18898 , n18899 , n18900 , n18901 , n18902 , n18903 , n18904 , n18905 , n18906 , n18907 , n18908 , n18909 , n18910 , n18911 , n18912 , n18913 , n18914 , n18915 , n18916 , n18917 , n18918 , n18919 , n18920 , n18921 , n18922 , n18923 , n18924 , n18925 , n18926 , n18927 , n18928 , n18929 , n18930 , n18931 , n18932 , n18933 , n18934 , n18935 , n18936 , n18937 , n18938 , n18939 , n18940 , n18941 , n18942 , n18943 , n18944 , n18945 , n18946 , n18947 , n18948 , n18949 , n18950 , n18951 , n18952 , n18953 , n18954 , n18955 , n18956 , n18957 , n18958 , n18959 , n18960 , n18961 , n18962 , n18963 , n18964 , n18965 , n18966 , n18967 , n18968 , n18969 , n18970 , n18971 , n18972 , n18973 , n18974 , n18975 , n18976 , n18977 , n18978 , n18979 , n18980 , n18981 , n18982 , n18983 , n18984 , n18985 , n18986 , n18987 , n18988 , n18989 , n18990 , n18991 , n18992 , n18993 , n18994 , n18995 , n18996 , n18997 , n18998 , n18999 , n19000 , n19001 , n19002 , n19003 , n19004 , n19005 , n19006 , n19007 , n19008 , n19009 , n19010 , n19011 , n19012 , n19013 , n19014 , n19015 , n19016 , n19017 , n19018 , n19019 , n19020 , n19021 , n19022 , n19023 , n19024 , n19025 , n19026 , n19027 , n19028 , n19029 , n19030 , n19031 , n19032 , n19033 , n19034 , n19035 , n19036 , n19037 , n19038 , n19039 , n19040 , n19041 , n19042 , n19043 , n19044 , n19045 , n19046 , n19047 , n19048 , n19049 , n19050 , n19051 , n19052 , n19053 , n19054 , n19055 , n19056 , n19057 , n19058 , n19059 , n19060 , n19061 , n19062 , n19063 , n19064 , n19065 , n19066 , n19067 , n19068 , n19069 , n19070 , n19071 , n19072 , n19073 , n19074 , n19075 , n19076 , n19077 , n19078 , n19079 , n19080 , n19081 , n19082 , n19083 , n19084 , n19085 , n19086 , n19087 , n19088 , n19089 , n19090 , n19091 , n19092 , n19093 , n19094 , n19095 , n19096 , n19097 , n19098 , n19099 , n19100 , n19101 , n19102 , n19103 , n19104 , n19105 , n19106 , n19107 , n19108 , n19109 , n19110 , n19111 , n19112 , n19113 , n19114 , n19115 , n19116 , n19117 , n19118 , n19119 , n19120 , n19121 , n19122 , n19123 , n19124 , n19125 , n19126 , n19127 , n19128 , n19129 , n19130 , n19131 , n19132 , n19133 , n19134 , n19135 , n19136 , n19137 , n19138 , n19139 , n19140 , n19141 , n19142 , n19143 , n19144 , n19145 , n19146 , n19147 , n19148 , n19149 , n19150 , n19151 , n19152 , n19153 , n19154 , n19155 , n19156 , n19157 , n19158 , n19159 , n19160 , n19161 , n19162 , n19163 , n19164 , n19165 , n19166 , n19167 , n19168 , n19169 , n19170 , n19171 , n19172 , n19173 , n19174 , n19175 , n19176 , n19177 , n19178 , n19179 , n19180 , n19181 , n19182 , n19183 , n19184 , n19185 , n19186 , n19187 , n19188 , n19189 , n19190 , n19191 , n19192 , n19193 , n19194 , n19195 , n19196 , n19197 , n19198 , n19199 , n19200 , n19201 , n19202 , n19203 , n19204 , n19205 , n19206 , n19207 , n19208 , n19209 , n19210 , n19211 , n19212 , n19213 , n19214 , n19215 , n19216 , n19217 , n19218 , n19219 , n19220 , n19221 , n19222 , n19223 , n19224 , n19225 , n19226 , n19227 , n19228 , n19229 , n19230 , n19231 , n19232 , n19233 , n19234 , n19235 , n19236 , n19237 , n19238 , n19239 , n19240 , n19241 , n19242 , n19243 , n19244 , n19245 , n19246 , n19247 , n19248 , n19249 , n19250 , n19251 , n19252 , n19253 , n19254 , n19255 , n19256 , n19257 , n19258 , n19259 , n19260 , n19261 , n19262 , n19263 , n19264 , n19265 , n19266 , n19267 , n19268 , n19269 , n19270 , n19271 , n19272 , n19273 , n19274 , n19275 , n19276 , n19277 , n19278 , n19279 , n19280 , n19281 , n19282 , n19283 , n19284 , n19285 , n19286 , n19287 , n19288 , n19289 , n19290 , n19291 , n19292 , n19293 , n19294 , n19295 , n19296 , n19297 , n19298 , n19299 , n19300 , n19301 , n19302 , n19303 , n19304 , n19305 , n19306 , n19307 , n19308 , n19309 , n19310 , n19311 , n19312 , n19313 , n19314 , n19315 , n19316 , n19317 , n19318 , n19319 , n19320 , n19321 , n19322 , n19323 , n19324 , n19325 , n19326 , n19327 , n19328 , n19329 , n19330 , n19331 , n19332 , n19333 , n19334 , n19335 , n19336 , n19337 , n19338 , n19339 , n19340 , n19341 , n19342 , n19343 , n19344 , n19345 , n19346 , n19347 , n19348 , n19349 , n19350 , n19351 , n19352 , n19353 , n19354 , n19355 , n19356 , n19357 , n19358 , n19359 , n19360 , n19361 , n19362 , n19363 , n19364 , n19365 , n19366 , n19367 , n19368 , n19369 , n19370 , n19371 , n19372 , n19373 , n19374 , n19375 , n19376 , n19377 , n19378 , n19379 , n19380 , n19381 , n19382 , n19383 , n19384 , n19385 , n19386 , n19387 , n19388 , n19389 , n19390 , n19391 , n19392 , n19393 , n19394 , n19395 , n19396 , n19397 , n19398 , n19399 , n19400 , n19401 , n19402 , n19403 , n19404 , n19405 , n19406 , n19407 , n19408 , n19409 , n19410 , n19411 , n19412 , n19413 , n19414 , n19415 , n19416 , n19417 , n19418 , n19419 , n19420 , n19421 , n19422 , n19423 , n19424 , n19425 , n19426 , n19427 , n19428 , n19429 , n19430 , n19431 , n19432 , n19433 , n19434 , n19435 , n19436 , n19437 , n19438 , n19439 , n19440 , n19441 , n19442 , n19443 , n19444 , n19445 , n19446 , n19447 , n19448 , n19449 , n19450 , n19451 , n19452 , n19453 , n19454 , n19455 , n19456 , n19457 , n19458 , n19459 , n19460 , n19461 , n19462 , n19463 , n19464 , n19465 , n19466 , n19467 , n19468 , n19469 , n19470 , n19471 , n19472 , n19473 , n19474 , n19475 , n19476 , n19477 , n19478 , n19479 , n19480 , n19481 , n19482 , n19483 , n19484 , n19485 , n19486 , n19487 , n19488 , n19489 , n19490 , n19491 , n19492 , n19493 , n19494 , n19495 , n19496 , n19497 , n19498 , n19499 , n19500 , n19501 , n19502 , n19503 , n19504 , n19505 , n19506 , n19507 , n19508 , n19509 , n19510 , n19511 , n19512 , n19513 , n19514 , n19515 , n19516 , n19517 , n19518 , n19519 , n19520 , n19521 , n19522 , n19523 , n19524 , n19525 , n19526 , n19527 , n19528 , n19529 , n19530 , n19531 , n19532 , n19533 , n19534 , n19535 , n19536 , n19537 , n19538 , n19539 , n19540 , n19541 , n19542 , n19543 , n19544 , n19545 , n19546 , n19547 , n19548 , n19549 , n19550 , n19551 , n19552 , n19553 , n19554 , n19555 , n19556 , n19557 , n19558 , n19559 , n19560 , n19561 , n19562 , n19563 , n19564 , n19565 , n19566 , n19567 , n19568 , n19569 , n19570 , n19571 , n19572 , n19573 , n19574 , n19575 , n19576 , n19577 , n19578 , n19579 , n19580 , n19581 , n19582 , n19583 , n19584 , n19585 , n19586 , n19587 , n19588 , n19589 , n19590 , n19591 , n19592 , n19593 , n19594 , n19595 , n19596 , n19597 , n19598 , n19599 , n19600 , n19601 , n19602 , n19603 , n19604 , n19605 , n19606 , n19607 , n19608 , n19609 , n19610 , n19611 , n19612 , n19613 , n19614 , n19615 , n19616 , n19617 , n19618 , n19619 , n19620 , n19621 , n19622 , n19623 , n19624 , n19625 , n19626 , n19627 , n19628 , n19629 , n19630 , n19631 , n19632 , n19633 , n19634 , n19635 , n19636 , n19637 , n19638 , n19639 , n19640 , n19641 , n19642 , n19643 , n19644 , n19645 , n19646 , n19647 , n19648 , n19649 , n19650 , n19651 , n19652 , n19653 , n19654 , n19655 , n19656 , n19657 , n19658 , n19659 , n19660 , n19661 , n19662 , n19663 , n19664 , n19665 , n19666 , n19667 , n19668 , n19669 , n19670 , n19671 , n19672 , n19673 , n19674 , n19675 , n19676 , n19677 , n19678 , n19679 , n19680 , n19681 , n19682 , n19683 , n19684 , n19685 , n19686 , n19687 , n19688 , n19689 , n19690 , n19691 , n19692 , n19693 , n19694 , n19695 , n19696 , n19697 , n19698 , n19699 , n19700 , n19701 , n19702 , n19703 , n19704 , n19705 , n19706 , n19707 , n19708 , n19709 , n19710 , n19711 , n19712 , n19713 , n19714 , n19715 , n19716 , n19717 , n19718 , n19719 , n19720 , n19721 , n19722 , n19723 , n19724 , n19725 , n19726 , n19727 , n19728 , n19729 , n19730 , n19731 , n19732 , n19733 , n19734 , n19735 , n19736 , n19737 , n19738 , n19739 , n19740 , n19741 , n19742 , n19743 , n19744 , n19745 , n19746 , n19747 , n19748 , n19749 , n19750 , n19751 , n19752 , n19753 , n19754 , n19755 , n19756 , n19757 , n19758 , n19759 , n19760 , n19761 , n19762 , n19763 , n19764 , n19765 , n19766 , n19767 , n19768 , n19769 , n19770 , n19771 , n19772 , n19773 , n19774 , n19775 , n19776 , n19777 , n19778 , n19779 , n19780 , n19781 , n19782 , n19783 , n19784 , n19785 , n19786 , n19787 , n19788 , n19789 , n19790 , n19791 , n19792 , n19793 , n19794 , n19795 , n19796 , n19797 , n19798 , n19799 , n19800 , n19801 , n19802 , n19803 , n19804 , n19805 , n19806 , n19807 , n19808 , n19809 , n19810 , n19811 , n19812 , n19813 , n19814 , n19815 , n19816 , n19817 , n19818 , n19819 , n19820 , n19821 , n19822 , n19823 , n19824 , n19825 , n19826 , n19827 , n19828 , n19829 , n19830 , n19831 , n19832 , n19833 , n19834 , n19835 , n19836 , n19837 , n19838 , n19839 , n19840 , n19841 , n19842 , n19843 , n19844 , n19845 , n19846 , n19847 , n19848 , n19849 , n19850 , n19851 , n19852 , n19853 , n19854 , n19855 , n19856 , n19857 , n19858 , n19859 , n19860 , n19861 , n19862 , n19863 , n19864 , n19865 , n19866 , n19867 , n19868 , n19869 , n19870 , n19871 , n19872 , n19873 , n19874 , n19875 , n19876 , n19877 , n19878 , n19879 , n19880 , n19881 , n19882 , n19883 , n19884 , n19885 , n19886 , n19887 , n19888 , n19889 , n19890 , n19891 , n19892 , n19893 , n19894 , n19895 , n19896 , n19897 , n19898 , n19899 , n19900 , n19901 , n19902 , n19903 , n19904 , n19905 , n19906 , n19907 , n19908 , n19909 , n19910 , n19911 , n19912 , n19913 , n19914 , n19915 , n19916 , n19917 , n19918 , n19919 , n19920 , n19921 , n19922 , n19923 , n19924 , n19925 , n19926 , n19927 , n19928 , n19929 , n19930 , n19931 , n19932 , n19933 , n19934 , n19935 , n19936 , n19937 , n19938 , n19939 , n19940 , n19941 , n19942 , n19943 , n19944 , n19945 , n19946 , n19947 , n19948 , n19949 , n19950 , n19951 , n19952 , n19953 , n19954 , n19955 , n19956 , n19957 , n19958 , n19959 , n19960 , n19961 , n19962 , n19963 , n19964 , n19965 , n19966 , n19967 , n19968 , n19969 , n19970 , n19971 , n19972 , n19973 , n19974 , n19975 , n19976 , n19977 , n19978 , n19979 , n19980 , n19981 , n19982 , n19983 , n19984 , n19985 , n19986 , n19987 , n19988 , n19989 , n19990 , n19991 , n19992 , n19993 , n19994 , n19995 , n19996 , n19997 , n19998 , n19999 , n20000 , n20001 , n20002 , n20003 , n20004 , n20005 , n20006 , n20007 , n20008 , n20009 , n20010 , n20011 , n20012 , n20013 , n20014 , n20015 , n20016 , n20017 , n20018 , n20019 , n20020 , n20021 , n20022 , n20023 , n20024 , n20025 , n20026 , n20027 , n20028 , n20029 , n20030 , n20031 , n20032 , n20033 , n20034 , n20035 , n20036 , n20037 , n20038 , n20039 , n20040 , n20041 , n20042 , n20043 , n20044 , n20045 , n20046 , n20047 , n20048 , n20049 , n20050 , n20051 , n20052 , n20053 , n20054 , n20055 , n20056 , n20057 , n20058 , n20059 , n20060 , n20061 , n20062 , n20063 , n20064 , n20065 , n20066 , n20067 , n20068 , n20069 , n20070 , n20071 , n20072 , n20073 , n20074 , n20075 , n20076 , n20077 , n20078 , n20079 , n20080 , n20081 , n20082 , n20083 , n20084 , n20085 , n20086 , n20087 , n20088 , n20089 , n20090 , n20091 , n20092 , n20093 , n20094 , n20095 , n20096 , n20097 , n20098 , n20099 , n20100 , n20101 , n20102 , n20103 , n20104 , n20105 , n20106 , n20107 , n20108 , n20109 , n20110 , n20111 , n20112 , n20113 , n20114 , n20115 , n20116 , n20117 , n20118 , n20119 , n20120 , n20121 , n20122 , n20123 , n20124 , n20125 , n20126 , n20127 , n20128 , n20129 , n20130 , n20131 , n20132 , n20133 , n20134 , n20135 , n20136 , n20137 , n20138 , n20139 , n20140 , n20141 , n20142 , n20143 , n20144 , n20145 , n20146 , n20147 , n20148 , n20149 , n20150 , n20151 , n20152 , n20153 , n20154 , n20155 , n20156 , n20157 , n20158 , n20159 , n20160 , n20161 , n20162 , n20163 , n20164 , n20165 , n20166 , n20167 , n20168 , n20169 , n20170 , n20171 , n20172 , n20173 , n20174 , n20175 , n20176 , n20177 , n20178 , n20179 , n20180 , n20181 , n20182 , n20183 , n20184 , n20185 , n20186 , n20187 , n20188 , n20189 , n20190 , n20191 , n20192 , n20193 , n20194 , n20195 , n20196 , n20197 , n20198 , n20199 , n20200 , n20201 , n20202 , n20203 , n20204 , n20205 , n20206 , n20207 , n20208 , n20209 , n20210 , n20211 , n20212 , n20213 , n20214 , n20215 , n20216 , n20217 , n20218 , n20219 , n20220 , n20221 , n20222 , n20223 , n20224 , n20225 , n20226 , n20227 , n20228 , n20229 , n20230 , n20231 , n20232 , n20233 , n20234 , n20235 , n20236 , n20237 , n20238 , n20239 , n20240 , n20241 , n20242 , n20243 , n20244 , n20245 , n20246 , n20247 , n20248 , n20249 , n20250 , n20251 , n20252 , n20253 , n20254 , n20255 , n20256 , n20257 , n20258 , n20259 , n20260 , n20261 , n20262 , n20263 , n20264 , n20265 , n20266 , n20267 , n20268 , n20269 , n20270 , n20271 , n20272 , n20273 , n20274 , n20275 , n20276 , n20277 , n20278 , n20279 , n20280 , n20281 , n20282 , n20283 , n20284 , n20285 , n20286 , n20287 , n20288 , n20289 , n20290 , n20291 , n20292 , n20293 , n20294 , n20295 , n20296 , n20297 , n20298 , n20299 , n20300 , n20301 , n20302 , n20303 , n20304 , n20305 , n20306 , n20307 , n20308 , n20309 , n20310 , n20311 , n20312 , n20313 , n20314 , n20315 , n20316 , n20317 , n20318 , n20319 , n20320 , n20321 , n20322 , n20323 , n20324 , n20325 , n20326 , n20327 , n20328 , n20329 , n20330 , n20331 , n20332 , n20333 , n20334 , n20335 , n20336 , n20337 , n20338 , n20339 , n20340 , n20341 , n20342 , n20343 , n20344 , n20345 , n20346 , n20347 , n20348 , n20349 , n20350 , n20351 , n20352 , n20353 , n20354 , n20355 , n20356 , n20357 , n20358 , n20359 , n20360 , n20361 , n20362 , n20363 , n20364 , n20365 , n20366 , n20367 , n20368 , n20369 , n20370 , n20371 , n20372 , n20373 , n20374 , n20375 , n20376 , n20377 , n20378 , n20379 , n20380 , n20381 , n20382 , n20383 , n20384 , n20385 , n20386 , n20387 , n20388 , n20389 , n20390 , n20391 , n20392 , n20393 , n20394 , n20395 , n20396 , n20397 , n20398 , n20399 , n20400 , n20401 , n20402 , n20403 , n20404 , n20405 , n20406 , n20407 , n20408 , n20409 , n20410 , n20411 , n20412 , n20413 , n20414 , n20415 , n20416 , n20417 , n20418 , n20419 , n20420 , n20421 , n20422 , n20423 , n20424 , n20425 , n20426 , n20427 , n20428 , n20429 , n20430 , n20431 , n20432 , n20433 , n20434 , n20435 , n20436 , n20437 , n20438 , n20439 , n20440 , n20441 , n20442 , n20443 , n20444 , n20445 , n20446 , n20447 , n20448 , n20449 , n20450 , n20451 , n20452 , n20453 , n20454 , n20455 , n20456 , n20457 , n20458 , n20459 , n20460 , n20461 , n20462 , n20463 , n20464 , n20465 , n20466 , n20467 , n20468 , n20469 , n20470 , n20471 , n20472 , n20473 , n20474 , n20475 , n20476 , n20477 , n20478 , n20479 , n20480 , n20481 , n20482 , n20483 , n20484 , n20485 , n20486 , n20487 , n20488 , n20489 , n20490 , n20491 , n20492 , n20493 , n20494 , n20495 , n20496 , n20497 , n20498 , n20499 , n20500 , n20501 , n20502 , n20503 , n20504 , n20505 , n20506 , n20507 , n20508 , n20509 , n20510 , n20511 , n20512 , n20513 , n20514 , n20515 , n20516 , n20517 , n20518 , n20519 , n20520 , n20521 , n20522 , n20523 , n20524 , n20525 , n20526 , n20527 , n20528 , n20529 , n20530 , n20531 , n20532 , n20533 , n20534 , n20535 , n20536 , n20537 , n20538 , n20539 , n20540 , n20541 , n20542 , n20543 , n20544 , n20545 , n20546 , n20547 , n20548 , n20549 , n20550 , n20551 , n20552 , n20553 , n20554 , n20555 , n20556 , n20557 , n20558 , n20559 , n20560 , n20561 , n20562 , n20563 , n20564 , n20565 , n20566 , n20567 , n20568 , n20569 , n20570 , n20571 , n20572 , n20573 , n20574 , n20575 , n20576 , n20577 , n20578 , n20579 , n20580 , n20581 , n20582 , n20583 , n20584 , n20585 , n20586 , n20587 , n20588 , n20589 , n20590 , n20591 , n20592 , n20593 , n20594 , n20595 , n20596 , n20597 , n20598 , n20599 , n20600 , n20601 , n20602 , n20603 , n20604 , n20605 , n20606 , n20607 , n20608 , n20609 , n20610 , n20611 , n20612 , n20613 , n20614 , n20615 , n20616 , n20617 , n20618 , n20619 , n20620 , n20621 , n20622 , n20623 , n20624 , n20625 , n20626 , n20627 , n20628 , n20629 , n20630 , n20631 , n20632 , n20633 , n20634 , n20635 , n20636 , n20637 , n20638 , n20639 , n20640 , n20641 , n20642 , n20643 , n20644 , n20645 , n20646 , n20647 , n20648 , n20649 , n20650 , n20651 , n20652 , n20653 , n20654 , n20655 , n20656 , n20657 , n20658 , n20659 , n20660 , n20661 , n20662 , n20663 , n20664 , n20665 , n20666 , n20667 , n20668 , n20669 , n20670 , n20671 , n20672 , n20673 , n20674 , n20675 , n20676 , n20677 , n20678 , n20679 , n20680 , n20681 , n20682 , n20683 , n20684 , n20685 , n20686 , n20687 , n20688 , n20689 , n20690 , n20691 , n20692 , n20693 , n20694 , n20695 , n20696 , n20697 , n20698 , n20699 , n20700 , n20701 , n20702 , n20703 , n20704 , n20705 , n20706 , n20707 , n20708 , n20709 , n20710 , n20711 , n20712 , n20713 , n20714 , n20715 , n20716 , n20717 , n20718 , n20719 , n20720 , n20721 , n20722 , n20723 , n20724 , n20725 , n20726 , n20727 , n20728 , n20729 , n20730 , n20731 , n20732 , n20733 , n20734 , n20735 , n20736 , n20737 , n20738 , n20739 , n20740 , n20741 , n20742 , n20743 , n20744 , n20745 , n20746 , n20747 , n20748 , n20749 , n20750 , n20751 , n20752 , n20753 , n20754 , n20755 , n20756 , n20757 , n20758 , n20759 , n20760 , n20761 , n20762 , n20763 , n20764 , n20765 , n20766 , n20767 , n20768 , n20769 , n20770 , n20771 , n20772 , n20773 , n20774 , n20775 , n20776 , n20777 , n20778 , n20779 , n20780 , n20781 , n20782 , n20783 , n20784 , n20785 , n20786 , n20787 , n20788 , n20789 , n20790 , n20791 , n20792 , n20793 , n20794 , n20795 , n20796 , n20797 , n20798 , n20799 , n20800 , n20801 , n20802 , n20803 , n20804 , n20805 , n20806 , n20807 , n20808 , n20809 , n20810 , n20811 , n20812 , n20813 , n20814 , n20815 , n20816 , n20817 , n20818 , n20819 , n20820 , n20821 , n20822 , n20823 , n20824 , n20825 , n20826 , n20827 , n20828 , n20829 , n20830 , n20831 , n20832 , n20833 , n20834 , n20835 , n20836 , n20837 , n20838 , n20839 , n20840 , n20841 , n20842 , n20843 , n20844 , n20845 , n20846 , n20847 , n20848 , n20849 , n20850 , n20851 , n20852 , n20853 , n20854 , n20855 , n20856 , n20857 , n20858 , n20859 , n20860 , n20861 , n20862 , n20863 , n20864 , n20865 , n20866 , n20867 , n20868 , n20869 , n20870 , n20871 , n20872 , n20873 , n20874 , n20875 , n20876 , n20877 , n20878 , n20879 , n20880 , n20881 , n20882 , n20883 , n20884 , n20885 , n20886 , n20887 , n20888 , n20889 , n20890 , n20891 , n20892 , n20893 , n20894 , n20895 , n20896 , n20897 , n20898 , n20899 , n20900 , n20901 , n20902 , n20903 , n20904 , n20905 , n20906 , n20907 , n20908 , n20909 , n20910 , n20911 , n20912 , n20913 , n20914 , n20915 , n20916 , n20917 , n20918 , n20919 , n20920 , n20921 , n20922 , n20923 , n20924 , n20925 , n20926 , n20927 , n20928 , n20929 , n20930 , n20931 , n20932 , n20933 , n20934 , n20935 , n20936 , n20937 , n20938 , n20939 , n20940 , n20941 , n20942 , n20943 , n20944 , n20945 , n20946 , n20947 , n20948 , n20949 , n20950 , n20951 , n20952 , n20953 , n20954 , n20955 , n20956 , n20957 , n20958 , n20959 , n20960 , n20961 , n20962 , n20963 , n20964 , n20965 , n20966 , n20967 , n20968 , n20969 , n20970 , n20971 , n20972 , n20973 , n20974 , n20975 , n20976 , n20977 , n20978 , n20979 , n20980 , n20981 , n20982 , n20983 , n20984 , n20985 , n20986 , n20987 , n20988 , n20989 , n20990 , n20991 , n20992 , n20993 , n20994 , n20995 , n20996 , n20997 , n20998 , n20999 , n21000 , n21001 , n21002 , n21003 , n21004 , n21005 , n21006 , n21007 , n21008 , n21009 , n21010 , n21011 , n21012 , n21013 , n21014 , n21015 , n21016 , n21017 , n21018 , n21019 , n21020 , n21021 , n21022 , n21023 , n21024 , n21025 , n21026 , n21027 , n21028 , n21029 , n21030 , n21031 , n21032 , n21033 , n21034 , n21035 , n21036 , n21037 , n21038 , n21039 , n21040 , n21041 , n21042 , n21043 , n21044 , n21045 , n21046 , n21047 , n21048 , n21049 , n21050 , n21051 , n21052 , n21053 , n21054 , n21055 , n21056 , n21057 , n21058 , n21059 , n21060 , n21061 , n21062 , n21063 , n21064 , n21065 , n21066 , n21067 , n21068 , n21069 , n21070 , n21071 , n21072 , n21073 , n21074 , n21075 , n21076 , n21077 , n21078 , n21079 , n21080 , n21081 , n21082 , n21083 , n21084 , n21085 , n21086 , n21087 , n21088 , n21089 , n21090 , n21091 , n21092 , n21093 , n21094 , n21095 , n21096 , n21097 , n21098 , n21099 , n21100 , n21101 , n21102 , n21103 , n21104 , n21105 , n21106 , n21107 , n21108 , n21109 , n21110 , n21111 , n21112 , n21113 , n21114 , n21115 , n21116 , n21117 , n21118 , n21119 , n21120 , n21121 , n21122 , n21123 , n21124 , n21125 , n21126 , n21127 , n21128 , n21129 , n21130 , n21131 , n21132 , n21133 , n21134 , n21135 , n21136 , n21137 , n21138 , n21139 , n21140 , n21141 , n21142 , n21143 , n21144 , n21145 , n21146 , n21147 , n21148 , n21149 , n21150 , n21151 , n21152 , n21153 , n21154 , n21155 , n21156 , n21157 , n21158 , n21159 , n21160 , n21161 , n21162 , n21163 , n21164 , n21165 , n21166 , n21167 , n21168 , n21169 , n21170 , n21171 , n21172 , n21173 , n21174 , n21175 , n21176 , n21177 , n21178 , n21179 , n21180 , n21181 , n21182 , n21183 , n21184 , n21185 , n21186 , n21187 , n21188 , n21189 , n21190 , n21191 , n21192 , n21193 , n21194 , n21195 , n21196 , n21197 , n21198 , n21199 , n21200 , n21201 , n21202 , n21203 , n21204 , n21205 , n21206 , n21207 , n21208 , n21209 , n21210 , n21211 , n21212 , n21213 , n21214 , n21215 , n21216 , n21217 , n21218 , n21219 , n21220 , n21221 , n21222 , n21223 , n21224 , n21225 , n21226 , n21227 , n21228 , n21229 , n21230 , n21231 , n21232 , n21233 , n21234 , n21235 , n21236 , n21237 , n21238 , n21239 , n21240 , n21241 , n21242 , n21243 , n21244 , n21245 , n21246 , n21247 , n21248 , n21249 , n21250 , n21251 , n21252 , n21253 , n21254 , n21255 , n21256 , n21257 , n21258 , n21259 , n21260 , n21261 , n21262 , n21263 , n21264 , n21265 , n21266 , n21267 , n21268 , n21269 , n21270 , n21271 , n21272 , n21273 , n21274 , n21275 , n21276 , n21277 , n21278 , n21279 , n21280 , n21281 , n21282 , n21283 , n21284 , n21285 , n21286 , n21287 , n21288 , n21289 , n21290 , n21291 , n21292 , n21293 , n21294 , n21295 , n21296 , n21297 , n21298 , n21299 , n21300 , n21301 , n21302 , n21303 , n21304 , n21305 , n21306 , n21307 , n21308 , n21309 , n21310 , n21311 , n21312 , n21313 , n21314 , n21315 , n21316 , n21317 , n21318 , n21319 , n21320 , n21321 , n21322 , n21323 , n21324 , n21325 , n21326 , n21327 , n21328 , n21329 , n21330 , n21331 , n21332 , n21333 , n21334 , n21335 , n21336 , n21337 , n21338 , n21339 , n21340 , n21341 , n21342 , n21343 , n21344 , n21345 , n21346 , n21347 , n21348 , n21349 , n21350 , n21351 , n21352 , n21353 , n21354 , n21355 , n21356 , n21357 , n21358 , n21359 , n21360 , n21361 , n21362 , n21363 , n21364 , n21365 , n21366 , n21367 , n21368 , n21369 , n21370 , n21371 , n21372 , n21373 , n21374 , n21375 , n21376 , n21377 , n21378 , n21379 , n21380 , n21381 , n21382 , n21383 , n21384 , n21385 , n21386 , n21387 , n21388 , n21389 , n21390 , n21391 , n21392 , n21393 , n21394 , n21395 , n21396 , n21397 , n21398 , n21399 , n21400 , n21401 , n21402 , n21403 , n21404 , n21405 , n21406 , n21407 , n21408 , n21409 , n21410 , n21411 , n21412 , n21413 , n21414 , n21415 , n21416 , n21417 , n21418 , n21419 , n21420 , n21421 , n21422 , n21423 , n21424 , n21425 , n21426 , n21427 , n21428 , n21429 , n21430 , n21431 , n21432 , n21433 , n21434 , n21435 , n21436 , n21437 , n21438 , n21439 , n21440 , n21441 , n21442 , n21443 , n21444 , n21445 , n21446 , n21447 , n21448 , n21449 , n21450 , n21451 , n21452 , n21453 , n21454 , n21455 , n21456 , n21457 , n21458 , n21459 , n21460 , n21461 , n21462 , n21463 , n21464 , n21465 , n21466 , n21467 , n21468 , n21469 , n21470 , n21471 , n21472 , n21473 , n21474 , n21475 , n21476 , n21477 , n21478 , n21479 , n21480 , n21481 , n21482 , n21483 , n21484 , n21485 , n21486 , n21487 , n21488 , n21489 , n21490 , n21491 , n21492 , n21493 , n21494 , n21495 , n21496 , n21497 , n21498 , n21499 , n21500 , n21501 , n21502 , n21503 , n21504 , n21505 , n21506 , n21507 , n21508 , n21509 , n21510 , n21511 , n21512 , n21513 , n21514 , n21515 , n21516 , n21517 , n21518 , n21519 , n21520 , n21521 , n21522 , n21523 , n21524 , n21525 , n21526 , n21527 , n21528 , n21529 , n21530 , n21531 , n21532 , n21533 , n21534 , n21535 , n21536 , n21537 , n21538 , n21539 , n21540 , n21541 , n21542 , n21543 , n21544 , n21545 , n21546 , n21547 , n21548 , n21549 , n21550 , n21551 , n21552 , n21553 , n21554 , n21555 , n21556 , n21557 , n21558 , n21559 , n21560 , n21561 , n21562 , n21563 , n21564 , n21565 , n21566 , n21567 , n21568 , n21569 , n21570 , n21571 , n21572 , n21573 , n21574 , n21575 , n21576 , n21577 , n21578 , n21579 , n21580 , n21581 , n21582 , n21583 , n21584 , n21585 , n21586 , n21587 , n21588 , n21589 , n21590 , n21591 , n21592 , n21593 , n21594 , n21595 , n21596 , n21597 , n21598 , n21599 , n21600 , n21601 , n21602 , n21603 , n21604 , n21605 , n21606 , n21607 , n21608 , n21609 , n21610 , n21611 , n21612 , n21613 , n21614 , n21615 , n21616 , n21617 , n21618 , n21619 , n21620 , n21621 , n21622 , n21623 , n21624 , n21625 , n21626 , n21627 , n21628 , n21629 , n21630 , n21631 , n21632 , n21633 , n21634 , n21635 , n21636 , n21637 , n21638 , n21639 , n21640 , n21641 , n21642 , n21643 , n21644 , n21645 , n21646 , n21647 , n21648 , n21649 , n21650 , n21651 , n21652 , n21653 , n21654 , n21655 , n21656 , n21657 , n21658 , n21659 , n21660 , n21661 , n21662 , n21663 , n21664 , n21665 , n21666 , n21667 , n21668 , n21669 , n21670 , n21671 , n21672 , n21673 , n21674 , n21675 , n21676 , n21677 , n21678 , n21679 , n21680 , n21681 , n21682 , n21683 , n21684 , n21685 , n21686 , n21687 , n21688 , n21689 , n21690 , n21691 , n21692 , n21693 , n21694 , n21695 , n21696 , n21697 , n21698 , n21699 , n21700 , n21701 , n21702 , n21703 , n21704 , n21705 , n21706 , n21707 , n21708 , n21709 , n21710 , n21711 , n21712 , n21713 , n21714 , n21715 , n21716 , n21717 , n21718 , n21719 , n21720 , n21721 , n21722 , n21723 , n21724 , n21725 , n21726 , n21727 , n21728 , n21729 , n21730 , n21731 , n21732 , n21733 , n21734 , n21735 , n21736 , n21737 , n21738 , n21739 , n21740 , n21741 , n21742 , n21743 , n21744 , n21745 , n21746 , n21747 , n21748 , n21749 , n21750 , n21751 , n21752 , n21753 , n21754 , n21755 , n21756 , n21757 , n21758 , n21759 , n21760 , n21761 , n21762 , n21763 , n21764 , n21765 , n21766 , n21767 , n21768 , n21769 , n21770 , n21771 , n21772 , n21773 , n21774 , n21775 , n21776 , n21777 , n21778 , n21779 , n21780 , n21781 , n21782 , n21783 , n21784 , n21785 , n21786 , n21787 , n21788 , n21789 , n21790 , n21791 , n21792 , n21793 , n21794 , n21795 , n21796 , n21797 , n21798 , n21799 , n21800 , n21801 , n21802 , n21803 , n21804 , n21805 , n21806 , n21807 , n21808 , n21809 , n21810 , n21811 , n21812 , n21813 , n21814 , n21815 , n21816 , n21817 , n21818 , n21819 , n21820 , n21821 , n21822 , n21823 , n21824 , n21825 , n21826 , n21827 , n21828 , n21829 , n21830 , n21831 , n21832 , n21833 , n21834 , n21835 , n21836 , n21837 , n21838 , n21839 , n21840 , n21841 , n21842 , n21843 , n21844 , n21845 , n21846 , n21847 , n21848 , n21849 , n21850 , n21851 , n21852 , n21853 , n21854 , n21855 , n21856 , n21857 , n21858 , n21859 , n21860 , n21861 , n21862 , n21863 , n21864 , n21865 , n21866 , n21867 , n21868 , n21869 , n21870 , n21871 , n21872 , n21873 , n21874 , n21875 , n21876 , n21877 , n21878 , n21879 , n21880 , n21881 , n21882 , n21883 , n21884 , n21885 , n21886 , n21887 , n21888 , n21889 , n21890 , n21891 , n21892 , n21893 , n21894 , n21895 , n21896 , n21897 , n21898 , n21899 , n21900 , n21901 , n21902 , n21903 , n21904 , n21905 , n21906 , n21907 , n21908 , n21909 , n21910 , n21911 , n21912 , n21913 , n21914 , n21915 , n21916 , n21917 , n21918 , n21919 , n21920 , n21921 , n21922 , n21923 , n21924 , n21925 , n21926 , n21927 , n21928 , n21929 , n21930 , n21931 , n21932 , n21933 , n21934 , n21935 , n21936 , n21937 , n21938 , n21939 , n21940 , n21941 , n21942 , n21943 , n21944 , n21945 , n21946 , n21947 , n21948 , n21949 , n21950 , n21951 , n21952 , n21953 , n21954 , n21955 , n21956 , n21957 , n21958 , n21959 , n21960 , n21961 , n21962 , n21963 , n21964 , n21965 , n21966 , n21967 , n21968 , n21969 , n21970 , n21971 , n21972 , n21973 , n21974 , n21975 , n21976 , n21977 , n21978 , n21979 , n21980 , n21981 , n21982 , n21983 , n21984 , n21985 , n21986 , n21987 , n21988 , n21989 , n21990 , n21991 , n21992 , n21993 , n21994 , n21995 , n21996 , n21997 , n21998 , n21999 , n22000 , n22001 , n22002 , n22003 , n22004 , n22005 , n22006 , n22007 , n22008 , n22009 , n22010 , n22011 , n22012 , n22013 , n22014 , n22015 , n22016 , n22017 , n22018 , n22019 , n22020 , n22021 , n22022 , n22023 , n22024 , n22025 , n22026 , n22027 , n22028 , n22029 , n22030 , n22031 , n22032 , n22033 , n22034 , n22035 , n22036 , n22037 , n22038 , n22039 , n22040 , n22041 , n22042 , n22043 , n22044 , n22045 , n22046 , n22047 , n22048 , n22049 , n22050 , n22051 , n22052 , n22053 , n22054 , n22055 , n22056 , n22057 , n22058 , n22059 , n22060 , n22061 , n22062 , n22063 , n22064 , n22065 , n22066 , n22067 , n22068 , n22069 , n22070 , n22071 , n22072 , n22073 , n22074 , n22075 , n22076 , n22077 , n22078 , n22079 , n22080 , n22081 , n22082 , n22083 , n22084 , n22085 , n22086 , n22087 , n22088 , n22089 , n22090 , n22091 , n22092 , n22093 , n22094 , n22095 , n22096 , n22097 , n22098 , n22099 , n22100 , n22101 , n22102 , n22103 , n22104 , n22105 , n22106 , n22107 , n22108 , n22109 , n22110 , n22111 , n22112 , n22113 , n22114 , n22115 , n22116 , n22117 , n22118 , n22119 , n22120 , n22121 , n22122 , n22123 , n22124 , n22125 , n22126 , n22127 , n22128 , n22129 , n22130 , n22131 , n22132 , n22133 , n22134 , n22135 , n22136 , n22137 , n22138 , n22139 , n22140 , n22141 , n22142 , n22143 , n22144 , n22145 , n22146 , n22147 , n22148 , n22149 , n22150 , n22151 , n22152 , n22153 , n22154 , n22155 , n22156 , n22157 , n22158 , n22159 , n22160 , n22161 , n22162 , n22163 , n22164 , n22165 , n22166 , n22167 , n22168 , n22169 , n22170 , n22171 , n22172 , n22173 , n22174 , n22175 , n22176 , n22177 , n22178 , n22179 , n22180 , n22181 , n22182 , n22183 , n22184 , n22185 , n22186 , n22187 , n22188 , n22189 , n22190 , n22191 , n22192 , n22193 , n22194 , n22195 , n22196 , n22197 , n22198 , n22199 , n22200 , n22201 , n22202 , n22203 , n22204 , n22205 , n22206 , n22207 , n22208 , n22209 , n22210 , n22211 , n22212 , n22213 , n22214 , n22215 , n22216 , n22217 , n22218 , n22219 , n22220 , n22221 , n22222 , n22223 , n22224 , n22225 , n22226 , n22227 , n22228 , n22229 , n22230 , n22231 , n22232 , n22233 , n22234 , n22235 , n22236 , n22237 , n22238 , n22239 , n22240 , n22241 , n22242 , n22243 , n22244 , n22245 , n22246 , n22247 , n22248 , n22249 , n22250 , n22251 , n22252 , n22253 , n22254 , n22255 , n22256 , n22257 , n22258 , n22259 , n22260 , n22261 , n22262 , n22263 , n22264 , n22265 , n22266 , n22267 , n22268 , n22269 , n22270 , n22271 , n22272 , n22273 , n22274 , n22275 , n22276 , n22277 , n22278 , n22279 , n22280 , n22281 , n22282 , n22283 , n22284 , n22285 , n22286 , n22287 , n22288 , n22289 , n22290 , n22291 , n22292 , n22293 , n22294 , n22295 , n22296 , n22297 , n22298 , n22299 , n22300 , n22301 , n22302 , n22303 , n22304 , n22305 , n22306 , n22307 , n22308 , n22309 , n22310 , n22311 , n22312 , n22313 , n22314 , n22315 , n22316 , n22317 , n22318 , n22319 , n22320 , n22321 , n22322 , n22323 , n22324 , n22325 , n22326 , n22327 , n22328 , n22329 , n22330 , n22331 , n22332 , n22333 , n22334 , n22335 , n22336 , n22337 , n22338 , n22339 , n22340 , n22341 , n22342 , n22343 , n22344 , n22345 , n22346 , n22347 , n22348 , n22349 , n22350 , n22351 , n22352 , n22353 , n22354 , n22355 , n22356 , n22357 , n22358 , n22359 , n22360 , n22361 , n22362 , n22363 , n22364 , n22365 , n22366 , n22367 , n22368 , n22369 , n22370 , n22371 , n22372 , n22373 , n22374 , n22375 , n22376 , n22377 , n22378 , n22379 , n22380 , n22381 , n22382 , n22383 , n22384 , n22385 , n22386 , n22387 , n22388 , n22389 , n22390 , n22391 , n22392 , n22393 , n22394 , n22395 , n22396 , n22397 , n22398 , n22399 , n22400 , n22401 , n22402 , n22403 , n22404 , n22405 , n22406 , n22407 , n22408 , n22409 , n22410 , n22411 , n22412 , n22413 , n22414 , n22415 , n22416 , n22417 , n22418 , n22419 , n22420 , n22421 , n22422 , n22423 , n22424 , n22425 , n22426 , n22427 , n22428 , n22429 , n22430 , n22431 , n22432 , n22433 , n22434 , n22435 , n22436 , n22437 , n22438 , n22439 , n22440 , n22441 , n22442 , n22443 , n22444 , n22445 , n22446 , n22447 , n22448 , n22449 , n22450 , n22451 , n22452 , n22453 , n22454 , n22455 , n22456 , n22457 , n22458 , n22459 , n22460 , n22461 , n22462 , n22463 , n22464 , n22465 , n22466 , n22467 , n22468 , n22469 , n22470 , n22471 , n22472 , n22473 , n22474 , n22475 , n22476 , n22477 , n22478 , n22479 , n22480 , n22481 , n22482 , n22483 , n22484 , n22485 , n22486 , n22487 , n22488 , n22489 , n22490 , n22491 , n22492 , n22493 , n22494 , n22495 , n22496 , n22497 , n22498 , n22499 , n22500 , n22501 , n22502 , n22503 , n22504 , n22505 , n22506 , n22507 , n22508 , n22509 , n22510 , n22511 , n22512 , n22513 , n22514 , n22515 , n22516 , n22517 , n22518 , n22519 , n22520 , n22521 , n22522 , n22523 , n22524 , n22525 , n22526 , n22527 , n22528 , n22529 , n22530 , n22531 , n22532 , n22533 , n22534 , n22535 , n22536 , n22537 , n22538 , n22539 , n22540 , n22541 , n22542 , n22543 , n22544 , n22545 , n22546 , n22547 , n22548 , n22549 , n22550 , n22551 , n22552 , n22553 , n22554 , n22555 , n22556 , n22557 , n22558 , n22559 , n22560 , n22561 , n22562 , n22563 , n22564 , n22565 , n22566 , n22567 , n22568 , n22569 , n22570 , n22571 , n22572 , n22573 , n22574 , n22575 , n22576 , n22577 , n22578 , n22579 , n22580 , n22581 , n22582 , n22583 , n22584 , n22585 , n22586 , n22587 , n22588 , n22589 , n22590 , n22591 , n22592 , n22593 , n22594 , n22595 , n22596 , n22597 , n22598 , n22599 , n22600 , n22601 , n22602 , n22603 , n22604 , n22605 , n22606 , n22607 , n22608 , n22609 , n22610 , n22611 , n22612 , n22613 , n22614 , n22615 , n22616 , n22617 , n22618 , n22619 , n22620 , n22621 , n22622 , n22623 , n22624 , n22625 , n22626 , n22627 , n22628 , n22629 , n22630 , n22631 , n22632 , n22633 , n22634 , n22635 , n22636 , n22637 , n22638 , n22639 , n22640 , n22641 , n22642 , n22643 , n22644 , n22645 , n22646 , n22647 , n22648 , n22649 , n22650 , n22651 , n22652 , n22653 , n22654 , n22655 , n22656 , n22657 , n22658 , n22659 , n22660 , n22661 , n22662 , n22663 , n22664 , n22665 , n22666 , n22667 , n22668 , n22669 , n22670 , n22671 , n22672 , n22673 , n22674 , n22675 , n22676 , n22677 , n22678 , n22679 , n22680 , n22681 , n22682 , n22683 , n22684 , n22685 , n22686 , n22687 , n22688 , n22689 , n22690 , n22691 , n22692 , n22693 , n22694 , n22695 , n22696 , n22697 , n22698 , n22699 , n22700 , n22701 , n22702 , n22703 , n22704 , n22705 , n22706 , n22707 , n22708 , n22709 , n22710 , n22711 , n22712 , n22713 , n22714 , n22715 , n22716 , n22717 , n22718 , n22719 , n22720 , n22721 , n22722 , n22723 , n22724 , n22725 , n22726 , n22727 , n22728 , n22729 , n22730 , n22731 , n22732 , n22733 , n22734 , n22735 , n22736 , n22737 , n22738 , n22739 , n22740 , n22741 , n22742 , n22743 , n22744 , n22745 , n22746 , n22747 , n22748 , n22749 , n22750 , n22751 , n22752 , n22753 , n22754 , n22755 , n22756 , n22757 , n22758 , n22759 , n22760 , n22761 , n22762 , n22763 , n22764 , n22765 , n22766 , n22767 , n22768 , n22769 , n22770 , n22771 , n22772 , n22773 , n22774 , n22775 , n22776 , n22777 , n22778 , n22779 , n22780 , n22781 , n22782 , n22783 , n22784 , n22785 , n22786 , n22787 , n22788 , n22789 , n22790 , n22791 , n22792 , n22793 , n22794 , n22795 , n22796 , n22797 , n22798 , n22799 , n22800 , n22801 , n22802 , n22803 , n22804 , n22805 , n22806 , n22807 , n22808 , n22809 , n22810 , n22811 , n22812 , n22813 , n22814 , n22815 , n22816 , n22817 , n22818 , n22819 , n22820 , n22821 , n22822 , n22823 , n22824 , n22825 , n22826 , n22827 , n22828 , n22829 , n22830 , n22831 , n22832 , n22833 , n22834 , n22835 , n22836 , n22837 , n22838 , n22839 , n22840 , n22841 , n22842 , n22843 , n22844 , n22845 , n22846 , n22847 , n22848 , n22849 , n22850 , n22851 , n22852 , n22853 , n22854 , n22855 , n22856 , n22857 , n22858 , n22859 , n22860 , n22861 , n22862 , n22863 , n22864 , n22865 , n22866 , n22867 , n22868 , n22869 , n22870 , n22871 , n22872 , n22873 , n22874 , n22875 , n22876 , n22877 , n22878 , n22879 , n22880 , n22881 , n22882 , n22883 , n22884 , n22885 , n22886 , n22887 , n22888 , n22889 , n22890 , n22891 , n22892 , n22893 , n22894 , n22895 , n22896 , n22897 , n22898 , n22899 , n22900 , n22901 , n22902 , n22903 , n22904 , n22905 , n22906 , n22907 , n22908 , n22909 , n22910 , n22911 , n22912 , n22913 , n22914 , n22915 , n22916 , n22917 , n22918 , n22919 , n22920 , n22921 , n22922 , n22923 , n22924 , n22925 , n22926 , n22927 , n22928 , n22929 , n22930 , n22931 , n22932 , n22933 , n22934 , n22935 , n22936 , n22937 , n22938 , n22939 , n22940 , n22941 , n22942 , n22943 , n22944 , n22945 , n22946 , n22947 , n22948 , n22949 , n22950 , n22951 , n22952 , n22953 , n22954 , n22955 , n22956 , n22957 , n22958 , n22959 , n22960 , n22961 , n22962 , n22963 , n22964 , n22965 , n22966 , n22967 , n22968 , n22969 , n22970 , n22971 , n22972 , n22973 , n22974 , n22975 , n22976 , n22977 , n22978 , n22979 , n22980 , n22981 , n22982 , n22983 , n22984 , n22985 , n22986 , n22987 , n22988 , n22989 , n22990 , n22991 , n22992 , n22993 , n22994 , n22995 , n22996 , n22997 , n22998 , n22999 , n23000 , n23001 , n23002 , n23003 , n23004 , n23005 , n23006 , n23007 , n23008 , n23009 , n23010 , n23011 , n23012 , n23013 , n23014 , n23015 , n23016 , n23017 , n23018 , n23019 , n23020 , n23021 , n23022 , n23023 , n23024 , n23025 , n23026 , n23027 , n23028 , n23029 , n23030 , n23031 , n23032 , n23033 , n23034 , n23035 , n23036 , n23037 , n23038 , n23039 , n23040 , n23041 , n23042 , n23043 , n23044 , n23045 , n23046 , n23047 , n23048 , n23049 , n23050 , n23051 , n23052 , n23053 , n23054 , n23055 , n23056 , n23057 , n23058 , n23059 , n23060 , n23061 , n23062 , n23063 , n23064 , n23065 , n23066 , n23067 , n23068 , n23069 , n23070 , n23071 , n23072 , n23073 , n23074 , n23075 , n23076 , n23077 , n23078 , n23079 , n23080 , n23081 , n23082 , n23083 , n23084 , n23085 , n23086 , n23087 , n23088 , n23089 , n23090 , n23091 , n23092 , n23093 , n23094 , n23095 , n23096 , n23097 , n23098 , n23099 , n23100 , n23101 , n23102 , n23103 , n23104 , n23105 , n23106 , n23107 , n23108 , n23109 , n23110 , n23111 , n23112 , n23113 , n23114 , n23115 , n23116 , n23117 , n23118 , n23119 , n23120 , n23121 , n23122 , n23123 , n23124 , n23125 , n23126 , n23127 , n23128 , n23129 , n23130 , n23131 , n23132 , n23133 , n23134 , n23135 , n23136 , n23137 , n23138 , n23139 , n23140 , n23141 , n23142 , n23143 , n23144 , n23145 , n23146 , n23147 , n23148 , n23149 , n23150 , n23151 , n23152 , n23153 , n23154 , n23155 , n23156 , n23157 , n23158 , n23159 , n23160 , n23161 , n23162 , n23163 , n23164 , n23165 , n23166 , n23167 , n23168 , n23169 , n23170 , n23171 , n23172 , n23173 , n23174 , n23175 , n23176 , n23177 , n23178 , n23179 , n23180 , n23181 , n23182 , n23183 , n23184 , n23185 , n23186 , n23187 , n23188 , n23189 , n23190 , n23191 , n23192 , n23193 , n23194 , n23195 , n23196 , n23197 , n23198 , n23199 , n23200 , n23201 , n23202 , n23203 , n23204 , n23205 , n23206 , n23207 , n23208 , n23209 , n23210 , n23211 , n23212 , n23213 , n23214 , n23215 , n23216 , n23217 , n23218 , n23219 , n23220 , n23221 , n23222 , n23223 , n23224 , n23225 , n23226 , n23227 , n23228 , n23229 , n23230 , n23231 , n23232 , n23233 , n23234 , n23235 , n23236 , n23237 , n23238 , n23239 , n23240 , n23241 , n23242 , n23243 , n23244 , n23245 , n23246 , n23247 , n23248 , n23249 , n23250 , n23251 , n23252 , n23253 , n23254 , n23255 , n23256 , n23257 , n23258 , n23259 , n23260 , n23261 , n23262 , n23263 , n23264 , n23265 , n23266 , n23267 , n23268 , n23269 , n23270 , n23271 , n23272 , n23273 , n23274 , n23275 , n23276 , n23277 , n23278 , n23279 , n23280 , n23281 , n23282 , n23283 , n23284 , n23285 , n23286 , n23287 , n23288 , n23289 , n23290 , n23291 , n23292 , n23293 , n23294 , n23295 , n23296 , n23297 , n23298 , n23299 , n23300 , n23301 , n23302 , n23303 , n23304 , n23305 , n23306 , n23307 , n23308 , n23309 , n23310 , n23311 , n23312 , n23313 , n23314 , n23315 , n23316 , n23317 , n23318 , n23319 , n23320 , n23321 , n23322 , n23323 , n23324 , n23325 , n23326 , n23327 , n23328 , n23329 , n23330 , n23331 , n23332 , n23333 , n23334 , n23335 , n23336 , n23337 , n23338 , n23339 , n23340 , n23341 , n23342 , n23343 , n23344 , n23345 , n23346 , n23347 , n23348 , n23349 , n23350 , n23351 , n23352 , n23353 , n23354 , n23355 , n23356 , n23357 , n23358 , n23359 , n23360 , n23361 , n23362 , n23363 , n23364 , n23365 , n23366 , n23367 , n23368 , n23369 , n23370 , n23371 , n23372 , n23373 , n23374 , n23375 , n23376 , n23377 , n23378 , n23379 , n23380 , n23381 , n23382 , n23383 , n23384 , n23385 , n23386 , n23387 , n23388 , n23389 , n23390 , n23391 , n23392 , n23393 , n23394 , n23395 , n23396 , n23397 , n23398 , n23399 , n23400 , n23401 , n23402 , n23403 , n23404 , n23405 , n23406 , n23407 , n23408 , n23409 , n23410 , n23411 , n23412 , n23413 , n23414 , n23415 , n23416 , n23417 , n23418 , n23419 , n23420 , n23421 , n23422 , n23423 , n23424 , n23425 , n23426 , n23427 , n23428 , n23429 , n23430 , n23431 , n23432 , n23433 , n23434 , n23435 , n23436 , n23437 , n23438 , n23439 , n23440 , n23441 , n23442 , n23443 , n23444 , n23445 , n23446 , n23447 , n23448 , n23449 , n23450 , n23451 , n23452 , n23453 , n23454 , n23455 , n23456 , n23457 , n23458 , n23459 , n23460 , n23461 , n23462 , n23463 , n23464 , n23465 , n23466 , n23467 , n23468 , n23469 , n23470 , n23471 , n23472 , n23473 , n23474 , n23475 , n23476 , n23477 , n23478 , n23479 , n23480 , n23481 , n23482 , n23483 , n23484 , n23485 , n23486 , n23487 , n23488 , n23489 , n23490 , n23491 , n23492 , n23493 , n23494 , n23495 , n23496 , n23497 , n23498 , n23499 , n23500 , n23501 , n23502 , n23503 , n23504 , n23505 , n23506 , n23507 , n23508 , n23509 , n23510 , n23511 , n23512 , n23513 , n23514 , n23515 , n23516 , n23517 , n23518 , n23519 , n23520 , n23521 , n23522 , n23523 , n23524 , n23525 , n23526 , n23527 , n23528 , n23529 , n23530 , n23531 , n23532 , n23533 , n23534 , n23535 , n23536 , n23537 , n23538 , n23539 , n23540 , n23541 , n23542 , n23543 , n23544 , n23545 , n23546 , n23547 , n23548 , n23549 , n23550 , n23551 , n23552 , n23553 , n23554 , n23555 , n23556 , n23557 , n23558 , n23559 , n23560 , n23561 , n23562 , n23563 , n23564 , n23565 , n23566 , n23567 , n23568 , n23569 , n23570 , n23571 , n23572 , n23573 , n23574 , n23575 , n23576 , n23577 , n23578 , n23579 , n23580 , n23581 , n23582 , n23583 , n23584 , n23585 , n23586 , n23587 , n23588 , n23589 , n23590 , n23591 , n23592 , n23593 , n23594 , n23595 , n23596 , n23597 , n23598 , n23599 , n23600 , n23601 , n23602 , n23603 , n23604 , n23605 , n23606 , n23607 , n23608 , n23609 , n23610 , n23611 , n23612 , n23613 , n23614 , n23615 , n23616 , n23617 , n23618 , n23619 , n23620 , n23621 , n23622 , n23623 , n23624 , n23625 , n23626 , n23627 , n23628 , n23629 , n23630 , n23631 , n23632 , n23633 , n23634 , n23635 , n23636 , n23637 , n23638 , n23639 , n23640 , n23641 , n23642 , n23643 , n23644 , n23645 , n23646 , n23647 , n23648 , n23649 , n23650 , n23651 , n23652 , n23653 , n23654 , n23655 , n23656 , n23657 , n23658 , n23659 , n23660 , n23661 , n23662 , n23663 , n23664 , n23665 , n23666 , n23667 , n23668 , n23669 , n23670 , n23671 , n23672 , n23673 , n23674 , n23675 , n23676 , n23677 , n23678 , n23679 , n23680 , n23681 , n23682 , n23683 , n23684 , n23685 , n23686 , n23687 , n23688 , n23689 , n23690 , n23691 , n23692 , n23693 , n23694 , n23695 , n23696 , n23697 , n23698 , n23699 , n23700 , n23701 , n23702 , n23703 , n23704 , n23705 , n23706 , n23707 , n23708 , n23709 , n23710 , n23711 , n23712 , n23713 , n23714 , n23715 , n23716 , n23717 , n23718 , n23719 , n23720 , n23721 , n23722 , n23723 , n23724 , n23725 , n23726 , n23727 , n23728 , n23729 , n23730 , n23731 , n23732 , n23733 , n23734 , n23735 , n23736 , n23737 , n23738 , n23739 , n23740 , n23741 , n23742 , n23743 , n23744 , n23745 , n23746 , n23747 , n23748 , n23749 , n23750 , n23751 , n23752 , n23753 , n23754 , n23755 , n23756 , n23757 , n23758 , n23759 , n23760 , n23761 , n23762 , n23763 , n23764 , n23765 , n23766 , n23767 , n23768 , n23769 , n23770 , n23771 , n23772 , n23773 , n23774 , n23775 , n23776 , n23777 , n23778 , n23779 , n23780 , n23781 , n23782 , n23783 , n23784 , n23785 , n23786 , n23787 , n23788 , n23789 , n23790 , n23791 , n23792 , n23793 , n23794 , n23795 , n23796 , n23797 , n23798 , n23799 , n23800 , n23801 , n23802 , n23803 , n23804 , n23805 , n23806 , n23807 , n23808 , n23809 , n23810 , n23811 , n23812 , n23813 , n23814 , n23815 , n23816 , n23817 , n23818 , n23819 , n23820 , n23821 , n23822 , n23823 , n23824 , n23825 , n23826 , n23827 , n23828 , n23829 , n23830 , n23831 , n23832 , n23833 , n23834 , n23835 , n23836 , n23837 , n23838 , n23839 , n23840 , n23841 , n23842 , n23843 , n23844 , n23845 , n23846 , n23847 , n23848 , n23849 , n23850 , n23851 , n23852 , n23853 , n23854 , n23855 , n23856 , n23857 , n23858 , n23859 , n23860 , n23861 , n23862 , n23863 , n23864 , n23865 , n23866 , n23867 , n23868 , n23869 , n23870 , n23871 , n23872 , n23873 , n23874 , n23875 , n23876 , n23877 , n23878 , n23879 , n23880 , n23881 , n23882 , n23883 , n23884 , n23885 , n23886 , n23887 , n23888 , n23889 , n23890 , n23891 , n23892 , n23893 , n23894 , n23895 , n23896 , n23897 , n23898 , n23899 , n23900 , n23901 , n23902 , n23903 , n23904 , n23905 , n23906 , n23907 , n23908 , n23909 , n23910 , n23911 , n23912 , n23913 , n23914 , n23915 , n23916 , n23917 , n23918 , n23919 , n23920 , n23921 , n23922 , n23923 , n23924 , n23925 , n23926 , n23927 , n23928 , n23929 , n23930 , n23931 , n23932 , n23933 , n23934 , n23935 , n23936 , n23937 , n23938 , n23939 , n23940 , n23941 , n23942 , n23943 , n23944 , n23945 , n23946 , n23947 , n23948 , n23949 , n23950 , n23951 , n23952 , n23953 , n23954 , n23955 , n23956 , n23957 , n23958 , n23959 , n23960 , n23961 , n23962 , n23963 , n23964 , n23965 , n23966 , n23967 , n23968 , n23969 , n23970 , n23971 , n23972 , n23973 , n23974 , n23975 , n23976 , n23977 , n23978 , n23979 , n23980 , n23981 , n23982 , n23983 , n23984 , n23985 , n23986 , n23987 , n23988 , n23989 , n23990 , n23991 , n23992 , n23993 , n23994 , n23995 , n23996 , n23997 , n23998 , n23999 , n24000 , n24001 , n24002 , n24003 , n24004 , n24005 , n24006 , n24007 , n24008 , n24009 , n24010 , n24011 , n24012 , n24013 , n24014 , n24015 , n24016 , n24017 , n24018 , n24019 , n24020 , n24021 , n24022 , n24023 , n24024 , n24025 , n24026 , n24027 , n24028 , n24029 , n24030 , n24031 , n24032 , n24033 , n24034 , n24035 , n24036 , n24037 , n24038 , n24039 , n24040 , n24041 , n24042 , n24043 , n24044 , n24045 , n24046 , n24047 , n24048 , n24049 , n24050 , n24051 , n24052 , n24053 , n24054 , n24055 , n24056 , n24057 , n24058 , n24059 , n24060 , n24061 , n24062 , n24063 , n24064 , n24065 , n24066 , n24067 , n24068 , n24069 , n24070 , n24071 , n24072 , n24073 , n24074 , n24075 , n24076 , n24077 , n24078 , n24079 , n24080 , n24081 , n24082 , n24083 , n24084 , n24085 , n24086 , n24087 , n24088 , n24089 , n24090 , n24091 , n24092 , n24093 , n24094 , n24095 , n24096 , n24097 , n24098 , n24099 , n24100 , n24101 , n24102 , n24103 , n24104 , n24105 , n24106 , n24107 , n24108 , n24109 , n24110 , n24111 , n24112 , n24113 , n24114 , n24115 , n24116 , n24117 , n24118 , n24119 , n24120 , n24121 , n24122 , n24123 , n24124 , n24125 , n24126 , n24127 , n24128 , n24129 , n24130 , n24131 , n24132 , n24133 , n24134 , n24135 , n24136 , n24137 , n24138 , n24139 , n24140 , n24141 , n24142 , n24143 , n24144 , n24145 , n24146 , n24147 , n24148 , n24149 , n24150 , n24151 , n24152 , n24153 , n24154 , n24155 , n24156 , n24157 , n24158 , n24159 , n24160 , n24161 , n24162 , n24163 , n24164 , n24165 , n24166 , n24167 , n24168 , n24169 , n24170 , n24171 , n24172 , n24173 , n24174 , n24175 , n24176 , n24177 , n24178 , n24179 , n24180 , n24181 , n24182 , n24183 , n24184 , n24185 , n24186 , n24187 , n24188 , n24189 , n24190 , n24191 , n24192 , n24193 , n24194 , n24195 , n24196 , n24197 , n24198 , n24199 , n24200 , n24201 , n24202 , n24203 , n24204 , n24205 , n24206 , n24207 , n24208 , n24209 , n24210 , n24211 , n24212 , n24213 , n24214 , n24215 , n24216 , n24217 , n24218 , n24219 , n24220 , n24221 , n24222 , n24223 , n24224 , n24225 , n24226 , n24227 , n24228 , n24229 , n24230 , n24231 , n24232 , n24233 , n24234 , n24235 , n24236 , n24237 , n24238 , n24239 , n24240 , n24241 , n24242 , n24243 , n24244 , n24245 , n24246 , n24247 , n24248 , n24249 , n24250 , n24251 , n24252 , n24253 , n24254 , n24255 , n24256 , n24257 , n24258 , n24259 , n24260 , n24261 , n24262 , n24263 , n24264 , n24265 , n24266 , n24267 , n24268 , n24269 , n24270 , n24271 , n24272 , n24273 , n24274 , n24275 , n24276 , n24277 , n24278 , n24279 , n24280 , n24281 , n24282 , n24283 , n24284 , n24285 , n24286 , n24287 , n24288 , n24289 , n24290 , n24291 , n24292 , n24293 , n24294 , n24295 , n24296 , n24297 , n24298 , n24299 , n24300 , n24301 , n24302 , n24303 , n24304 , n24305 , n24306 , n24307 , n24308 , n24309 , n24310 , n24311 , n24312 , n24313 , n24314 , n24315 , n24316 , n24317 , n24318 , n24319 , n24320 , n24321 , n24322 , n24323 , n24324 , n24325 , n24326 , n24327 , n24328 , n24329 , n24330 , n24331 , n24332 , n24333 , n24334 , n24335 , n24336 , n24337 , n24338 , n24339 , n24340 , n24341 , n24342 , n24343 , n24344 , n24345 , n24346 , n24347 , n24348 , n24349 , n24350 , n24351 , n24352 , n24353 , n24354 , n24355 , n24356 , n24357 , n24358 , n24359 , n24360 , n24361 , n24362 , n24363 , n24364 , n24365 , n24366 , n24367 , n24368 , n24369 , n24370 , n24371 , n24372 , n24373 , n24374 , n24375 , n24376 , n24377 , n24378 , n24379 , n24380 , n24381 , n24382 , n24383 , n24384 , n24385 , n24386 , n24387 , n24388 , n24389 , n24390 , n24391 , n24392 , n24393 , n24394 , n24395 , n24396 , n24397 , n24398 , n24399 , n24400 , n24401 , n24402 , n24403 , n24404 , n24405 , n24406 , n24407 , n24408 , n24409 , n24410 , n24411 , n24412 , n24413 , n24414 , n24415 , n24416 , n24417 , n24418 , n24419 , n24420 , n24421 , n24422 , n24423 , n24424 , n24425 , n24426 , n24427 , n24428 , n24429 , n24430 , n24431 , n24432 , n24433 , n24434 , n24435 , n24436 , n24437 , n24438 , n24439 , n24440 , n24441 , n24442 , n24443 , n24444 , n24445 , n24446 , n24447 , n24448 , n24449 , n24450 , n24451 , n24452 , n24453 , n24454 , n24455 , n24456 , n24457 , n24458 , n24459 , n24460 , n24461 , n24462 , n24463 , n24464 , n24465 , n24466 , n24467 , n24468 , n24469 , n24470 , n24471 , n24472 , n24473 , n24474 , n24475 , n24476 , n24477 , n24478 , n24479 , n24480 , n24481 , n24482 , n24483 , n24484 , n24485 , n24486 , n24487 , n24488 , n24489 , n24490 , n24491 , n24492 , n24493 , n24494 , n24495 , n24496 , n24497 , n24498 , n24499 , n24500 , n24501 , n24502 , n24503 , n24504 , n24505 , n24506 , n24507 , n24508 , n24509 , n24510 , n24511 , n24512 , n24513 , n24514 , n24515 , n24516 , n24517 , n24518 , n24519 , n24520 , n24521 , n24522 , n24523 , n24524 , n24525 , n24526 , n24527 , n24528 , n24529 , n24530 , n24531 , n24532 , n24533 , n24534 , n24535 , n24536 , n24537 , n24538 , n24539 , n24540 , n24541 , n24542 , n24543 , n24544 , n24545 , n24546 , n24547 , n24548 , n24549 , n24550 , n24551 , n24552 , n24553 , n24554 , n24555 , n24556 , n24557 , n24558 , n24559 , n24560 , n24561 , n24562 , n24563 , n24564 , n24565 , n24566 , n24567 , n24568 , n24569 , n24570 , n24571 , n24572 , n24573 , n24574 , n24575 , n24576 , n24577 , n24578 , n24579 , n24580 , n24581 , n24582 , n24583 , n24584 , n24585 , n24586 , n24587 , n24588 , n24589 , n24590 , n24591 , n24592 , n24593 , n24594 , n24595 , n24596 , n24597 , n24598 , n24599 , n24600 , n24601 , n24602 , n24603 , n24604 , n24605 , n24606 , n24607 , n24608 , n24609 , n24610 , n24611 , n24612 , n24613 , n24614 , n24615 , n24616 , n24617 , n24618 , n24619 , n24620 , n24621 , n24622 , n24623 , n24624 , n24625 , n24626 , n24627 , n24628 , n24629 , n24630 , n24631 , n24632 , n24633 , n24634 , n24635 , n24636 , n24637 , n24638 , n24639 , n24640 , n24641 , n24642 , n24643 , n24644 , n24645 , n24646 , n24647 , n24648 , n24649 , n24650 , n24651 , n24652 , n24653 , n24654 , n24655 , n24656 , n24657 , n24658 , n24659 , n24660 , n24661 , n24662 , n24663 , n24664 , n24665 , n24666 , n24667 , n24668 , n24669 , n24670 , n24671 , n24672 , n24673 , n24674 , n24675 , n24676 , n24677 , n24678 , n24679 , n24680 , n24681 , n24682 , n24683 , n24684 , n24685 , n24686 , n24687 , n24688 , n24689 , n24690 , n24691 , n24692 , n24693 , n24694 , n24695 , n24696 , n24697 , n24698 , n24699 , n24700 , n24701 , n24702 , n24703 , n24704 , n24705 , n24706 , n24707 , n24708 , n24709 , n24710 , n24711 , n24712 , n24713 , n24714 , n24715 , n24716 , n24717 , n24718 , n24719 , n24720 , n24721 , n24722 , n24723 , n24724 , n24725 , n24726 , n24727 , n24728 , n24729 , n24730 , n24731 , n24732 , n24733 , n24734 , n24735 , n24736 , n24737 , n24738 , n24739 , n24740 , n24741 , n24742 , n24743 , n24744 , n24745 , n24746 , n24747 , n24748 , n24749 , n24750 , n24751 , n24752 , n24753 , n24754 , n24755 , n24756 , n24757 , n24758 , n24759 , n24760 , n24761 , n24762 , n24763 , n24764 , n24765 , n24766 , n24767 , n24768 , n24769 , n24770 , n24771 , n24772 , n24773 , n24774 , n24775 , n24776 , n24777 , n24778 , n24779 , n24780 , n24781 , n24782 , n24783 , n24784 , n24785 , n24786 , n24787 , n24788 , n24789 , n24790 , n24791 , n24792 , n24793 , n24794 , n24795 , n24796 , n24797 , n24798 , n24799 , n24800 , n24801 , n24802 , n24803 , n24804 , n24805 , n24806 , n24807 , n24808 , n24809 , n24810 , n24811 , n24812 , n24813 , n24814 , n24815 , n24816 , n24817 , n24818 , n24819 , n24820 , n24821 , n24822 , n24823 , n24824 , n24825 , n24826 , n24827 , n24828 , n24829 , n24830 , n24831 , n24832 , n24833 , n24834 , n24835 , n24836 , n24837 , n24838 , n24839 , n24840 , n24841 , n24842 , n24843 , n24844 , n24845 , n24846 , n24847 , n24848 , n24849 , n24850 , n24851 , n24852 , n24853 , n24854 , n24855 , n24856 , n24857 , n24858 , n24859 , n24860 , n24861 , n24862 , n24863 , n24864 , n24865 , n24866 , n24867 , n24868 , n24869 , n24870 , n24871 , n24872 , n24873 , n24874 , n24875 , n24876 , n24877 , n24878 , n24879 , n24880 , n24881 , n24882 , n24883 , n24884 , n24885 , n24886 , n24887 , n24888 , n24889 , n24890 , n24891 , n24892 , n24893 , n24894 , n24895 , n24896 , n24897 , n24898 , n24899 , n24900 , n24901 , n24902 , n24903 , n24904 , n24905 , n24906 , n24907 , n24908 , n24909 , n24910 , n24911 , n24912 , n24913 , n24914 , n24915 , n24916 , n24917 , n24918 , n24919 , n24920 , n24921 , n24922 , n24923 , n24924 , n24925 , n24926 , n24927 , n24928 , n24929 , n24930 , n24931 , n24932 , n24933 , n24934 , n24935 , n24936 , n24937 , n24938 , n24939 , n24940 , n24941 , n24942 , n24943 , n24944 , n24945 , n24946 , n24947 , n24948 , n24949 , n24950 , n24951 , n24952 , n24953 , n24954 , n24955 , n24956 , n24957 , n24958 , n24959 , n24960 , n24961 , n24962 , n24963 , n24964 , n24965 , n24966 , n24967 , n24968 , n24969 , n24970 , n24971 , n24972 , n24973 , n24974 , n24975 , n24976 , n24977 , n24978 , n24979 , n24980 , n24981 , n24982 , n24983 , n24984 , n24985 , n24986 , n24987 , n24988 , n24989 , n24990 , n24991 , n24992 , n24993 , n24994 , n24995 , n24996 , n24997 , n24998 , n24999 , n25000 , n25001 , n25002 , n25003 , n25004 , n25005 , n25006 , n25007 , n25008 , n25009 , n25010 , n25011 , n25012 , n25013 , n25014 , n25015 , n25016 , n25017 , n25018 , n25019 , n25020 , n25021 , n25022 , n25023 , n25024 , n25025 , n25026 , n25027 , n25028 , n25029 , n25030 , n25031 , n25032 , n25033 , n25034 , n25035 , n25036 , n25037 , n25038 , n25039 , n25040 , n25041 , n25042 , n25043 , n25044 , n25045 , n25046 , n25047 , n25048 , n25049 , n25050 , n25051 , n25052 , n25053 , n25054 , n25055 , n25056 , n25057 , n25058 , n25059 , n25060 , n25061 , n25062 , n25063 , n25064 , n25065 , n25066 , n25067 , n25068 , n25069 , n25070 , n25071 , n25072 , n25073 , n25074 , n25075 , n25076 , n25077 , n25078 , n25079 , n25080 , n25081 , n25082 , n25083 , n25084 , n25085 , n25086 , n25087 , n25088 , n25089 , n25090 , n25091 , n25092 , n25093 , n25094 , n25095 , n25096 , n25097 , n25098 , n25099 , n25100 , n25101 , n25102 , n25103 , n25104 , n25105 , n25106 , n25107 , n25108 , n25109 , n25110 , n25111 , n25112 , n25113 , n25114 , n25115 , n25116 , n25117 , n25118 , n25119 , n25120 , n25121 , n25122 , n25123 , n25124 , n25125 , n25126 , n25127 , n25128 , n25129 , n25130 , n25131 , n25132 , n25133 , n25134 , n25135 , n25136 , n25137 , n25138 , n25139 , n25140 , n25141 , n25142 , n25143 , n25144 , n25145 , n25146 , n25147 , n25148 , n25149 , n25150 , n25151 , n25152 , n25153 , n25154 , n25155 , n25156 , n25157 , n25158 , n25159 , n25160 , n25161 , n25162 , n25163 , n25164 , n25165 , n25166 , n25167 , n25168 , n25169 , n25170 , n25171 , n25172 , n25173 , n25174 , n25175 , n25176 , n25177 , n25178 , n25179 , n25180 , n25181 , n25182 , n25183 , n25184 , n25185 , n25186 , n25187 , n25188 , n25189 , n25190 , n25191 , n25192 , n25193 , n25194 , n25195 , n25196 , n25197 , n25198 , n25199 , n25200 , n25201 , n25202 , n25203 , n25204 , n25205 , n25206 , n25207 , n25208 , n25209 , n25210 , n25211 , n25212 , n25213 , n25214 , n25215 , n25216 , n25217 , n25218 , n25219 , n25220 , n25221 , n25222 , n25223 , n25224 , n25225 , n25226 , n25227 , n25228 , n25229 , n25230 , n25231 , n25232 , n25233 , n25234 , n25235 , n25236 , n25237 , n25238 , n25239 , n25240 , n25241 , n25242 , n25243 , n25244 , n25245 , n25246 , n25247 , n25248 , n25249 , n25250 , n25251 , n25252 , n25253 , n25254 , n25255 , n25256 , n25257 , n25258 , n25259 , n25260 , n25261 , n25262 , n25263 , n25264 , n25265 , n25266 , n25267 , n25268 , n25269 , n25270 , n25271 , n25272 , n25273 , n25274 , n25275 , n25276 , n25277 , n25278 , n25279 , n25280 , n25281 , n25282 , n25283 , n25284 , n25285 , n25286 , n25287 , n25288 , n25289 , n25290 , n25291 , n25292 , n25293 , n25294 , n25295 , n25296 , n25297 , n25298 , n25299 , n25300 , n25301 , n25302 , n25303 , n25304 , n25305 , n25306 , n25307 , n25308 , n25309 , n25310 , n25311 , n25312 , n25313 , n25314 , n25315 , n25316 , n25317 , n25318 , n25319 , n25320 , n25321 , n25322 , n25323 , n25324 , n25325 , n25326 , n25327 , n25328 , n25329 , n25330 , n25331 , n25332 , n25333 , n25334 , n25335 , n25336 , n25337 , n25338 , n25339 , n25340 , n25341 , n25342 , n25343 , n25344 , n25345 , n25346 , n25347 , n25348 , n25349 , n25350 , n25351 , n25352 , n25353 , n25354 , n25355 , n25356 , n25357 , n25358 , n25359 , n25360 , n25361 , n25362 , n25363 , n25364 , n25365 , n25366 , n25367 , n25368 , n25369 , n25370 , n25371 , n25372 , n25373 , n25374 , n25375 , n25376 , n25377 , n25378 , n25379 , n25380 , n25381 , n25382 , n25383 , n25384 , n25385 , n25386 , n25387 , n25388 , n25389 , n25390 , n25391 , n25392 , n25393 , n25394 , n25395 , n25396 , n25397 , n25398 , n25399 , n25400 , n25401 , n25402 , n25403 , n25404 , n25405 , n25406 , n25407 , n25408 , n25409 , n25410 , n25411 , n25412 , n25413 , n25414 , n25415 , n25416 , n25417 , n25418 , n25419 , n25420 , n25421 , n25422 , n25423 , n25424 , n25425 , n25426 , n25427 , n25428 , n25429 , n25430 , n25431 , n25432 , n25433 , n25434 , n25435 , n25436 , n25437 , n25438 , n25439 , n25440 , n25441 , n25442 , n25443 , n25444 , n25445 , n25446 , n25447 , n25448 , n25449 , n25450 , n25451 , n25452 , n25453 , n25454 , n25455 , n25456 , n25457 , n25458 , n25459 , n25460 , n25461 , n25462 , n25463 , n25464 , n25465 , n25466 , n25467 , n25468 , n25469 , n25470 , n25471 , n25472 , n25473 , n25474 , n25475 , n25476 , n25477 , n25478 , n25479 , n25480 , n25481 , n25482 , n25483 , n25484 , n25485 , n25486 , n25487 , n25488 , n25489 , n25490 , n25491 , n25492 , n25493 , n25494 , n25495 , n25496 , n25497 , n25498 , n25499 , n25500 , n25501 , n25502 , n25503 , n25504 , n25505 , n25506 , n25507 , n25508 , n25509 , n25510 , n25511 , n25512 , n25513 , n25514 , n25515 , n25516 , n25517 , n25518 , n25519 , n25520 , n25521 , n25522 , n25523 , n25524 , n25525 , n25526 , n25527 , n25528 , n25529 , n25530 , n25531 , n25532 , n25533 , n25534 , n25535 , n25536 , n25537 , n25538 , n25539 , n25540 , n25541 , n25542 , n25543 , n25544 , n25545 , n25546 , n25547 , n25548 , n25549 , n25550 , n25551 , n25552 , n25553 , n25554 , n25555 , n25556 , n25557 , n25558 , n25559 , n25560 , n25561 , n25562 , n25563 , n25564 , n25565 , n25566 , n25567 , n25568 , n25569 , n25570 , n25571 , n25572 , n25573 , n25574 , n25575 , n25576 , n25577 , n25578 , n25579 , n25580 , n25581 , n25582 , n25583 , n25584 , n25585 , n25586 , n25587 , n25588 , n25589 , n25590 , n25591 , n25592 , n25593 , n25594 , n25595 , n25596 , n25597 , n25598 , n25599 , n25600 , n25601 , n25602 , n25603 , n25604 , n25605 , n25606 , n25607 , n25608 , n25609 , n25610 , n25611 , n25612 , n25613 , n25614 , n25615 , n25616 , n25617 , n25618 , n25619 , n25620 , n25621 , n25622 , n25623 , n25624 , n25625 , n25626 , n25627 , n25628 , n25629 , n25630 , n25631 , n25632 , n25633 , n25634 , n25635 , n25636 , n25637 , n25638 , n25639 , n25640 , n25641 , n25642 , n25643 , n25644 , n25645 , n25646 , n25647 , n25648 , n25649 , n25650 , n25651 , n25652 , n25653 , n25654 , n25655 , n25656 , n25657 , n25658 , n25659 , n25660 , n25661 , n25662 , n25663 , n25664 , n25665 , n25666 , n25667 , n25668 , n25669 , n25670 , n25671 , n25672 , n25673 , n25674 , n25675 , n25676 , n25677 , n25678 , n25679 , n25680 , n25681 , n25682 , n25683 , n25684 , n25685 , n25686 , n25687 , n25688 , n25689 , n25690 , n25691 , n25692 , n25693 , n25694 , n25695 , n25696 , n25697 , n25698 , n25699 , n25700 , n25701 , n25702 , n25703 , n25704 , n25705 , n25706 , n25707 , n25708 , n25709 , n25710 , n25711 , n25712 , n25713 , n25714 , n25715 , n25716 , n25717 , n25718 , n25719 , n25720 , n25721 , n25722 , n25723 , n25724 , n25725 , n25726 , n25727 , n25728 , n25729 , n25730 , n25731 , n25732 , n25733 , n25734 , n25735 , n25736 , n25737 , n25738 , n25739 , n25740 , n25741 , n25742 , n25743 , n25744 , n25745 , n25746 , n25747 , n25748 , n25749 , n25750 , n25751 , n25752 , n25753 , n25754 , n25755 , n25756 , n25757 , n25758 , n25759 , n25760 , n25761 , n25762 , n25763 , n25764 , n25765 , n25766 , n25767 , n25768 , n25769 , n25770 , n25771 , n25772 , n25773 , n25774 , n25775 , n25776 , n25777 , n25778 , n25779 , n25780 , n25781 , n25782 , n25783 , n25784 , n25785 , n25786 , n25787 , n25788 , n25789 , n25790 , n25791 , n25792 , n25793 , n25794 , n25795 , n25796 , n25797 , n25798 , n25799 , n25800 , n25801 , n25802 , n25803 , n25804 , n25805 , n25806 , n25807 , n25808 , n25809 , n25810 , n25811 , n25812 , n25813 , n25814 , n25815 , n25816 , n25817 , n25818 , n25819 , n25820 , n25821 , n25822 , n25823 , n25824 , n25825 , n25826 , n25827 , n25828 , n25829 , n25830 , n25831 , n25832 , n25833 , n25834 , n25835 , n25836 , n25837 , n25838 , n25839 , n25840 , n25841 , n25842 , n25843 , n25844 , n25845 , n25846 , n25847 , n25848 , n25849 , n25850 , n25851 , n25852 , n25853 , n25854 , n25855 , n25856 , n25857 , n25858 , n25859 , n25860 , n25861 , n25862 , n25863 , n25864 , n25865 , n25866 , n25867 , n25868 , n25869 , n25870 , n25871 , n25872 , n25873 , n25874 , n25875 , n25876 , n25877 , n25878 , n25879 , n25880 , n25881 , n25882 , n25883 , n25884 , n25885 , n25886 , n25887 , n25888 , n25889 , n25890 , n25891 , n25892 , n25893 , n25894 , n25895 , n25896 , n25897 , n25898 , n25899 , n25900 , n25901 , n25902 , n25903 , n25904 , n25905 , n25906 , n25907 , n25908 , n25909 , n25910 , n25911 , n25912 , n25913 , n25914 , n25915 , n25916 , n25917 , n25918 , n25919 , n25920 , n25921 , n25922 , n25923 , n25924 , n25925 , n25926 , n25927 , n25928 , n25929 , n25930 , n25931 , n25932 , n25933 , n25934 , n25935 , n25936 , n25937 , n25938 , n25939 , n25940 , n25941 , n25942 , n25943 , n25944 , n25945 , n25946 , n25947 , n25948 , n25949 , n25950 , n25951 , n25952 , n25953 , n25954 , n25955 , n25956 , n25957 , n25958 , n25959 , n25960 , n25961 , n25962 , n25963 , n25964 , n25965 , n25966 , n25967 , n25968 , n25969 , n25970 , n25971 , n25972 , n25973 , n25974 , n25975 , n25976 , n25977 , n25978 , n25979 , n25980 , n25981 , n25982 , n25983 , n25984 , n25985 , n25986 , n25987 , n25988 , n25989 , n25990 , n25991 , n25992 , n25993 , n25994 , n25995 , n25996 , n25997 , n25998 , n25999 , n26000 , n26001 , n26002 , n26003 , n26004 , n26005 , n26006 , n26007 , n26008 , n26009 , n26010 , n26011 , n26012 , n26013 , n26014 , n26015 , n26016 , n26017 , n26018 , n26019 , n26020 , n26021 , n26022 , n26023 , n26024 , n26025 , n26026 , n26027 , n26028 , n26029 , n26030 , n26031 , n26032 , n26033 , n26034 , n26035 , n26036 , n26037 , n26038 , n26039 , n26040 , n26041 , n26042 , n26043 , n26044 , n26045 , n26046 , n26047 , n26048 , n26049 , n26050 , n26051 , n26052 , n26053 , n26054 , n26055 , n26056 , n26057 , n26058 , n26059 , n26060 , n26061 , n26062 , n26063 , n26064 , n26065 , n26066 , n26067 , n26068 , n26069 , n26070 , n26071 , n26072 , n26073 , n26074 , n26075 , n26076 , n26077 , n26078 , n26079 , n26080 , n26081 , n26082 , n26083 , n26084 , n26085 , n26086 , n26087 , n26088 , n26089 , n26090 , n26091 , n26092 , n26093 , n26094 , n26095 , n26096 , n26097 , n26098 , n26099 , n26100 , n26101 , n26102 , n26103 , n26104 , n26105 , n26106 , n26107 , n26108 , n26109 , n26110 , n26111 , n26112 , n26113 , n26114 , n26115 , n26116 , n26117 , n26118 , n26119 , n26120 , n26121 , n26122 , n26123 , n26124 , n26125 , n26126 , n26127 , n26128 , n26129 , n26130 , n26131 , n26132 , n26133 , n26134 , n26135 , n26136 , n26137 , n26138 , n26139 , n26140 , n26141 , n26142 , n26143 , n26144 , n26145 , n26146 , n26147 , n26148 , n26149 , n26150 , n26151 , n26152 , n26153 , n26154 , n26155 , n26156 , n26157 , n26158 , n26159 , n26160 , n26161 , n26162 , n26163 , n26164 , n26165 , n26166 , n26167 , n26168 , n26169 , n26170 , n26171 , n26172 , n26173 , n26174 , n26175 , n26176 , n26177 , n26178 , n26179 , n26180 , n26181 , n26182 , n26183 , n26184 , n26185 , n26186 , n26187 , n26188 , n26189 , n26190 , n26191 , n26192 , n26193 , n26194 , n26195 , n26196 , n26197 , n26198 , n26199 , n26200 , n26201 , n26202 , n26203 , n26204 , n26205 , n26206 , n26207 , n26208 , n26209 , n26210 , n26211 , n26212 , n26213 , n26214 , n26215 , n26216 , n26217 , n26218 , n26219 , n26220 , n26221 , n26222 , n26223 , n26224 , n26225 , n26226 , n26227 , n26228 , n26229 , n26230 , n26231 , n26232 , n26233 , n26234 , n26235 , n26236 , n26237 , n26238 , n26239 , n26240 , n26241 , n26242 , n26243 , n26244 , n26245 , n26246 , n26247 , n26248 , n26249 , n26250 , n26251 , n26252 , n26253 , n26254 , n26255 , n26256 , n26257 , n26258 , n26259 , n26260 , n26261 , n26262 , n26263 , n26264 , n26265 , n26266 , n26267 , n26268 , n26269 , n26270 , n26271 , n26272 , n26273 , n26274 , n26275 , n26276 , n26277 , n26278 , n26279 , n26280 , n26281 , n26282 , n26283 , n26284 , n26285 , n26286 , n26287 , n26288 , n26289 , n26290 , n26291 , n26292 , n26293 , n26294 , n26295 , n26296 , n26297 , n26298 , n26299 , n26300 , n26301 , n26302 , n26303 , n26304 , n26305 , n26306 , n26307 , n26308 , n26309 , n26310 , n26311 , n26312 , n26313 , n26314 , n26315 , n26316 , n26317 , n26318 , n26319 , n26320 , n26321 , n26322 , n26323 , n26324 , n26325 , n26326 , n26327 , n26328 , n26329 , n26330 , n26331 , n26332 , n26333 , n26334 , n26335 , n26336 , n26337 , n26338 , n26339 , n26340 , n26341 , n26342 , n26343 , n26344 , n26345 , n26346 , n26347 , n26348 , n26349 , n26350 , n26351 , n26352 , n26353 , n26354 , n26355 , n26356 , n26357 , n26358 , n26359 , n26360 , n26361 , n26362 , n26363 , n26364 , n26365 , n26366 , n26367 , n26368 , n26369 , n26370 , n26371 , n26372 , n26373 , n26374 , n26375 , n26376 , n26377 , n26378 , n26379 , n26380 , n26381 , n26382 , n26383 , n26384 , n26385 , n26386 , n26387 , n26388 , n26389 , n26390 , n26391 , n26392 , n26393 , n26394 , n26395 , n26396 , n26397 , n26398 , n26399 , n26400 , n26401 , n26402 , n26403 , n26404 , n26405 , n26406 , n26407 , n26408 , n26409 , n26410 , n26411 , n26412 , n26413 , n26414 , n26415 , n26416 , n26417 , n26418 , n26419 , n26420 , n26421 , n26422 , n26423 , n26424 , n26425 , n26426 , n26427 , n26428 , n26429 , n26430 , n26431 , n26432 , n26433 , n26434 , n26435 , n26436 , n26437 , n26438 , n26439 , n26440 , n26441 , n26442 , n26443 , n26444 , n26445 , n26446 , n26447 , n26448 , n26449 , n26450 , n26451 , n26452 , n26453 , n26454 , n26455 , n26456 , n26457 , n26458 , n26459 , n26460 , n26461 , n26462 , n26463 , n26464 , n26465 , n26466 , n26467 , n26468 , n26469 , n26470 , n26471 , n26472 , n26473 , n26474 , n26475 , n26476 , n26477 , n26478 , n26479 , n26480 , n26481 , n26482 , n26483 , n26484 , n26485 , n26486 , n26487 , n26488 , n26489 , n26490 , n26491 , n26492 , n26493 , n26494 , n26495 , n26496 , n26497 , n26498 , n26499 , n26500 , n26501 , n26502 , n26503 , n26504 , n26505 , n26506 , n26507 , n26508 , n26509 , n26510 , n26511 , n26512 , n26513 , n26514 , n26515 , n26516 , n26517 , n26518 , n26519 , n26520 , n26521 , n26522 , n26523 , n26524 , n26525 , n26526 , n26527 , n26528 , n26529 , n26530 , n26531 , n26532 , n26533 , n26534 , n26535 , n26536 , n26537 , n26538 , n26539 , n26540 , n26541 , n26542 , n26543 , n26544 , n26545 , n26546 , n26547 , n26548 , n26549 , n26550 , n26551 , n26552 , n26553 , n26554 , n26555 , n26556 , n26557 , n26558 , n26559 , n26560 , n26561 , n26562 , n26563 , n26564 , n26565 , n26566 , n26567 , n26568 , n26569 , n26570 , n26571 , n26572 , n26573 , n26574 , n26575 , n26576 , n26577 , n26578 , n26579 , n26580 , n26581 , n26582 , n26583 , n26584 , n26585 , n26586 , n26587 , n26588 , n26589 , n26590 , n26591 , n26592 , n26593 , n26594 , n26595 , n26596 , n26597 , n26598 , n26599 , n26600 , n26601 , n26602 , n26603 , n26604 , n26605 , n26606 , n26607 , n26608 , n26609 , n26610 , n26611 , n26612 , n26613 , n26614 , n26615 , n26616 , n26617 , n26618 , n26619 , n26620 , n26621 , n26622 , n26623 , n26624 , n26625 , n26626 , n26627 , n26628 , n26629 , n26630 , n26631 , n26632 , n26633 , n26634 , n26635 , n26636 , n26637 , n26638 , n26639 , n26640 , n26641 , n26642 , n26643 , n26644 , n26645 , n26646 , n26647 , n26648 , n26649 , n26650 , n26651 , n26652 , n26653 , n26654 , n26655 , n26656 , n26657 , n26658 , n26659 , n26660 , n26661 , n26662 , n26663 , n26664 , n26665 , n26666 , n26667 , n26668 , n26669 , n26670 , n26671 , n26672 , n26673 , n26674 , n26675 , n26676 , n26677 , n26678 , n26679 , n26680 , n26681 , n26682 , n26683 , n26684 , n26685 , n26686 , n26687 , n26688 , n26689 , n26690 , n26691 , n26692 , n26693 , n26694 , n26695 , n26696 , n26697 , n26698 , n26699 , n26700 , n26701 , n26702 , n26703 , n26704 , n26705 , n26706 , n26707 , n26708 , n26709 , n26710 , n26711 , n26712 , n26713 , n26714 , n26715 , n26716 , n26717 , n26718 , n26719 , n26720 , n26721 , n26722 , n26723 , n26724 , n26725 , n26726 , n26727 , n26728 , n26729 , n26730 , n26731 , n26732 , n26733 , n26734 , n26735 , n26736 , n26737 , n26738 , n26739 , n26740 , n26741 , n26742 , n26743 , n26744 , n26745 , n26746 , n26747 , n26748 , n26749 , n26750 , n26751 , n26752 , n26753 , n26754 , n26755 , n26756 , n26757 , n26758 , n26759 , n26760 , n26761 , n26762 , n26763 , n26764 , n26765 , n26766 , n26767 , n26768 , n26769 , n26770 , n26771 , n26772 , n26773 , n26774 , n26775 , n26776 , n26777 , n26778 , n26779 , n26780 , n26781 , n26782 , n26783 , n26784 , n26785 , n26786 , n26787 , n26788 , n26789 , n26790 , n26791 , n26792 , n26793 , n26794 , n26795 , n26796 , n26797 , n26798 , n26799 , n26800 , n26801 , n26802 , n26803 , n26804 , n26805 , n26806 , n26807 , n26808 , n26809 , n26810 , n26811 , n26812 , n26813 , n26814 , n26815 , n26816 , n26817 , n26818 , n26819 , n26820 , n26821 , n26822 , n26823 , n26824 , n26825 , n26826 , n26827 , n26828 , n26829 , n26830 , n26831 , n26832 , n26833 , n26834 , n26835 , n26836 , n26837 , n26838 , n26839 , n26840 , n26841 , n26842 , n26843 , n26844 , n26845 , n26846 , n26847 , n26848 , n26849 , n26850 , n26851 , n26852 , n26853 , n26854 , n26855 , n26856 , n26857 , n26858 , n26859 , n26860 , n26861 , n26862 , n26863 , n26864 , n26865 , n26866 , n26867 , n26868 , n26869 , n26870 , n26871 , n26872 , n26873 , n26874 , n26875 , n26876 , n26877 , n26878 , n26879 , n26880 , n26881 , n26882 , n26883 , n26884 , n26885 , n26886 , n26887 , n26888 , n26889 , n26890 , n26891 , n26892 , n26893 , n26894 , n26895 , n26896 , n26897 , n26898 , n26899 , n26900 , n26901 , n26902 , n26903 , n26904 , n26905 , n26906 , n26907 , n26908 , n26909 , n26910 , n26911 , n26912 , n26913 , n26914 , n26915 , n26916 , n26917 , n26918 , n26919 , n26920 , n26921 , n26922 , n26923 , n26924 , n26925 , n26926 , n26927 , n26928 , n26929 , n26930 , n26931 , n26932 , n26933 , n26934 , n26935 , n26936 , n26937 , n26938 , n26939 , n26940 , n26941 , n26942 , n26943 , n26944 , n26945 , n26946 , n26947 , n26948 , n26949 , n26950 , n26951 , n26952 , n26953 , n26954 , n26955 , n26956 , n26957 , n26958 , n26959 , n26960 , n26961 , n26962 , n26963 , n26964 , n26965 , n26966 , n26967 , n26968 , n26969 , n26970 , n26971 , n26972 , n26973 , n26974 , n26975 , n26976 , n26977 , n26978 , n26979 , n26980 , n26981 , n26982 , n26983 , n26984 , n26985 , n26986 , n26987 , n26988 , n26989 , n26990 , n26991 , n26992 , n26993 , n26994 , n26995 , n26996 , n26997 , n26998 , n26999 , n27000 , n27001 , n27002 , n27003 , n27004 , n27005 , n27006 , n27007 , n27008 , n27009 , n27010 , n27011 , n27012 , n27013 , n27014 , n27015 , n27016 , n27017 , n27018 , n27019 , n27020 , n27021 , n27022 , n27023 , n27024 , n27025 , n27026 , n27027 , n27028 , n27029 , n27030 , n27031 , n27032 , n27033 , n27034 , n27035 , n27036 , n27037 , n27038 , n27039 , n27040 , n27041 , n27042 , n27043 , n27044 , n27045 , n27046 , n27047 , n27048 , n27049 , n27050 , n27051 , n27052 , n27053 , n27054 , n27055 , n27056 , n27057 , n27058 , n27059 , n27060 , n27061 , n27062 , n27063 , n27064 , n27065 , n27066 , n27067 , n27068 , n27069 , n27070 , n27071 , n27072 , n27073 , n27074 , n27075 , n27076 , n27077 , n27078 , n27079 , n27080 , n27081 , n27082 , n27083 , n27084 , n27085 , n27086 , n27087 , n27088 , n27089 , n27090 , n27091 , n27092 , n27093 , n27094 , n27095 , n27096 , n27097 , n27098 , n27099 , n27100 , n27101 , n27102 , n27103 , n27104 , n27105 , n27106 , n27107 , n27108 , n27109 , n27110 , n27111 , n27112 , n27113 , n27114 , n27115 , n27116 , n27117 , n27118 , n27119 , n27120 , n27121 , n27122 , n27123 , n27124 , n27125 , n27126 , n27127 , n27128 , n27129 , n27130 , n27131 , n27132 , n27133 , n27134 , n27135 , n27136 , n27137 , n27138 , n27139 , n27140 , n27141 , n27142 , n27143 , n27144 , n27145 , n27146 , n27147 , n27148 , n27149 , n27150 , n27151 , n27152 , n27153 , n27154 , n27155 , n27156 , n27157 , n27158 , n27159 , n27160 , n27161 , n27162 , n27163 , n27164 , n27165 , n27166 , n27167 , n27168 , n27169 , n27170 , n27171 , n27172 , n27173 , n27174 , n27175 , n27176 , n27177 , n27178 , n27179 , n27180 , n27181 , n27182 , n27183 , n27184 , n27185 , n27186 , n27187 , n27188 , n27189 , n27190 , n27191 , n27192 , n27193 , n27194 , n27195 , n27196 , n27197 , n27198 , n27199 , n27200 , n27201 , n27202 , n27203 , n27204 , n27205 , n27206 , n27207 , n27208 , n27209 , n27210 , n27211 , n27212 , n27213 , n27214 , n27215 , n27216 , n27217 , n27218 , n27219 , n27220 , n27221 , n27222 , n27223 , n27224 , n27225 , n27226 , n27227 , n27228 , n27229 , n27230 , n27231 , n27232 , n27233 , n27234 , n27235 , n27236 , n27237 , n27238 , n27239 , n27240 , n27241 , n27242 , n27243 , n27244 , n27245 , n27246 , n27247 , n27248 , n27249 , n27250 , n27251 , n27252 , n27253 , n27254 , n27255 , n27256 , n27257 , n27258 , n27259 , n27260 , n27261 , n27262 , n27263 , n27264 , n27265 , n27266 , n27267 , n27268 , n27269 , n27270 , n27271 , n27272 , n27273 , n27274 , n27275 , n27276 , n27277 , n27278 , n27279 , n27280 , n27281 , n27282 , n27283 , n27284 , n27285 , n27286 , n27287 , n27288 , n27289 , n27290 , n27291 , n27292 , n27293 , n27294 , n27295 , n27296 , n27297 , n27298 , n27299 , n27300 , n27301 , n27302 , n27303 , n27304 , n27305 , n27306 , n27307 , n27308 , n27309 , n27310 , n27311 , n27312 , n27313 , n27314 , n27315 , n27316 , n27317 , n27318 , n27319 , n27320 , n27321 , n27322 , n27323 , n27324 , n27325 , n27326 , n27327 , n27328 , n27329 , n27330 , n27331 , n27332 , n27333 , n27334 , n27335 , n27336 , n27337 , n27338 , n27339 , n27340 , n27341 , n27342 , n27343 , n27344 , n27345 , n27346 , n27347 , n27348 , n27349 , n27350 , n27351 , n27352 , n27353 , n27354 , n27355 , n27356 , n27357 , n27358 , n27359 , n27360 , n27361 , n27362 , n27363 , n27364 , n27365 , n27366 , n27367 , n27368 , n27369 , n27370 , n27371 , n27372 , n27373 , n27374 , n27375 , n27376 , n27377 , n27378 , n27379 , n27380 , n27381 , n27382 , n27383 , n27384 , n27385 , n27386 , n27387 , n27388 , n27389 , n27390 , n27391 , n27392 , n27393 , n27394 , n27395 , n27396 , n27397 , n27398 , n27399 , n27400 , n27401 , n27402 , n27403 , n27404 , n27405 , n27406 , n27407 , n27408 , n27409 , n27410 , n27411 , n27412 , n27413 , n27414 , n27415 , n27416 , n27417 , n27418 , n27419 , n27420 , n27421 , n27422 , n27423 , n27424 , n27425 , n27426 , n27427 , n27428 , n27429 , n27430 , n27431 , n27432 , n27433 , n27434 , n27435 , n27436 , n27437 , n27438 , n27439 , n27440 , n27441 , n27442 , n27443 , n27444 , n27445 , n27446 , n27447 , n27448 , n27449 , n27450 , n27451 , n27452 , n27453 , n27454 , n27455 , n27456 , n27457 , n27458 , n27459 , n27460 , n27461 , n27462 , n27463 , n27464 , n27465 , n27466 , n27467 , n27468 , n27469 , n27470 , n27471 , n27472 , n27473 , n27474 , n27475 , n27476 , n27477 , n27478 , n27479 , n27480 , n27481 , n27482 , n27483 , n27484 , n27485 , n27486 , n27487 , n27488 , n27489 , n27490 , n27491 , n27492 , n27493 , n27494 , n27495 , n27496 , n27497 , n27498 , n27499 , n27500 , n27501 , n27502 , n27503 , n27504 , n27505 , n27506 , n27507 , n27508 , n27509 , n27510 , n27511 , n27512 , n27513 , n27514 , n27515 , n27516 , n27517 , n27518 , n27519 , n27520 , n27521 , n27522 , n27523 , n27524 , n27525 , n27526 , n27527 , n27528 , n27529 , n27530 , n27531 , n27532 , n27533 , n27534 , n27535 , n27536 , n27537 , n27538 , n27539 , n27540 , n27541 , n27542 , n27543 , n27544 , n27545 , n27546 , n27547 , n27548 , n27549 , n27550 , n27551 , n27552 , n27553 , n27554 , n27555 , n27556 , n27557 , n27558 , n27559 , n27560 , n27561 , n27562 , n27563 , n27564 , n27565 , n27566 , n27567 , n27568 , n27569 , n27570 , n27571 , n27572 , n27573 , n27574 , n27575 , n27576 , n27577 , n27578 , n27579 , n27580 , n27581 , n27582 , n27583 , n27584 , n27585 , n27586 , n27587 , n27588 , n27589 , n27590 , n27591 , n27592 , n27593 , n27594 , n27595 , n27596 , n27597 , n27598 , n27599 , n27600 , n27601 , n27602 , n27603 , n27604 , n27605 , n27606 , n27607 , n27608 , n27609 , n27610 , n27611 , n27612 , n27613 , n27614 , n27615 , n27616 , n27617 , n27618 , n27619 , n27620 , n27621 , n27622 , n27623 , n27624 , n27625 , n27626 , n27627 , n27628 , n27629 , n27630 , n27631 , n27632 , n27633 , n27634 , n27635 , n27636 , n27637 , n27638 , n27639 , n27640 , n27641 , n27642 , n27643 , n27644 , n27645 , n27646 , n27647 , n27648 , n27649 , n27650 , n27651 , n27652 , n27653 , n27654 , n27655 , n27656 , n27657 , n27658 , n27659 , n27660 , n27661 , n27662 , n27663 , n27664 , n27665 , n27666 , n27667 , n27668 , n27669 , n27670 , n27671 , n27672 , n27673 , n27674 , n27675 , n27676 , n27677 , n27678 , n27679 , n27680 , n27681 , n27682 , n27683 , n27684 , n27685 , n27686 , n27687 , n27688 , n27689 , n27690 , n27691 , n27692 , n27693 , n27694 , n27695 , n27696 , n27697 , n27698 , n27699 , n27700 , n27701 , n27702 , n27703 , n27704 , n27705 , n27706 , n27707 , n27708 , n27709 , n27710 , n27711 , n27712 , n27713 , n27714 , n27715 , n27716 , n27717 , n27718 , n27719 , n27720 , n27721 , n27722 , n27723 , n27724 , n27725 , n27726 , n27727 , n27728 , n27729 , n27730 , n27731 , n27732 , n27733 , n27734 , n27735 , n27736 , n27737 , n27738 , n27739 , n27740 , n27741 , n27742 , n27743 , n27744 , n27745 , n27746 , n27747 , n27748 , n27749 , n27750 , n27751 , n27752 , n27753 , n27754 , n27755 , n27756 , n27757 , n27758 , n27759 , n27760 , n27761 , n27762 , n27763 , n27764 , n27765 , n27766 , n27767 , n27768 , n27769 , n27770 , n27771 , n27772 , n27773 , n27774 , n27775 , n27776 , n27777 , n27778 , n27779 , n27780 , n27781 , n27782 , n27783 , n27784 , n27785 , n27786 , n27787 , n27788 , n27789 , n27790 , n27791 , n27792 , n27793 , n27794 , n27795 , n27796 , n27797 , n27798 , n27799 , n27800 , n27801 , n27802 , n27803 , n27804 , n27805 , n27806 , n27807 , n27808 , n27809 , n27810 , n27811 , n27812 , n27813 , n27814 , n27815 , n27816 , n27817 , n27818 , n27819 , n27820 , n27821 , n27822 , n27823 , n27824 , n27825 , n27826 , n27827 , n27828 , n27829 , n27830 , n27831 , n27832 , n27833 , n27834 , n27835 , n27836 , n27837 , n27838 , n27839 , n27840 , n27841 , n27842 , n27843 , n27844 , n27845 , n27846 , n27847 , n27848 , n27849 , n27850 , n27851 , n27852 , n27853 , n27854 , n27855 , n27856 , n27857 , n27858 , n27859 , n27860 , n27861 , n27862 , n27863 , n27864 , n27865 , n27866 , n27867 , n27868 , n27869 , n27870 , n27871 , n27872 , n27873 , n27874 , n27875 , n27876 , n27877 , n27878 , n27879 , n27880 , n27881 , n27882 , n27883 , n27884 , n27885 , n27886 , n27887 , n27888 , n27889 , n27890 , n27891 , n27892 , n27893 , n27894 , n27895 , n27896 , n27897 , n27898 , n27899 , n27900 , n27901 , n27902 , n27903 , n27904 , n27905 , n27906 , n27907 , n27908 , n27909 , n27910 , n27911 , n27912 , n27913 , n27914 , n27915 , n27916 , n27917 , n27918 , n27919 , n27920 , n27921 , n27922 , n27923 , n27924 , n27925 , n27926 , n27927 , n27928 , n27929 , n27930 , n27931 , n27932 , n27933 , n27934 , n27935 , n27936 , n27937 , n27938 , n27939 , n27940 , n27941 , n27942 , n27943 , n27944 , n27945 , n27946 , n27947 , n27948 , n27949 , n27950 , n27951 , n27952 , n27953 , n27954 , n27955 , n27956 , n27957 , n27958 , n27959 , n27960 , n27961 , n27962 , n27963 , n27964 , n27965 , n27966 , n27967 , n27968 , n27969 , n27970 , n27971 , n27972 , n27973 , n27974 , n27975 , n27976 , n27977 , n27978 , n27979 , n27980 , n27981 , n27982 , n27983 , n27984 , n27985 , n27986 , n27987 , n27988 , n27989 , n27990 , n27991 , n27992 , n27993 , n27994 , n27995 , n27996 , n27997 , n27998 , n27999 , n28000 , n28001 , n28002 , n28003 , n28004 , n28005 , n28006 , n28007 , n28008 , n28009 , n28010 , n28011 , n28012 , n28013 , n28014 , n28015 , n28016 , n28017 , n28018 , n28019 , n28020 , n28021 , n28022 , n28023 , n28024 , n28025 , n28026 , n28027 , n28028 , n28029 , n28030 , n28031 , n28032 , n28033 , n28034 , n28035 , n28036 , n28037 , n28038 , n28039 , n28040 , n28041 , n28042 , n28043 , n28044 , n28045 , n28046 , n28047 , n28048 , n28049 , n28050 , n28051 , n28052 , n28053 , n28054 , n28055 , n28056 , n28057 , n28058 , n28059 , n28060 , n28061 , n28062 , n28063 , n28064 , n28065 , n28066 , n28067 , n28068 , n28069 , n28070 , n28071 , n28072 , n28073 , n28074 , n28075 , n28076 , n28077 , n28078 , n28079 , n28080 , n28081 , n28082 , n28083 , n28084 , n28085 , n28086 , n28087 , n28088 , n28089 , n28090 , n28091 , n28092 , n28093 , n28094 , n28095 , n28096 , n28097 , n28098 , n28099 , n28100 , n28101 , n28102 , n28103 , n28104 , n28105 , n28106 , n28107 , n28108 , n28109 , n28110 , n28111 , n28112 , n28113 , n28114 , n28115 , n28116 , n28117 , n28118 , n28119 , n28120 , n28121 , n28122 , n28123 , n28124 , n28125 , n28126 , n28127 , n28128 , n28129 , n28130 , n28131 , n28132 , n28133 , n28134 , n28135 , n28136 , n28137 , n28138 , n28139 , n28140 , n28141 , n28142 , n28143 , n28144 , n28145 , n28146 , n28147 , n28148 , n28149 , n28150 , n28151 , n28152 , n28153 , n28154 , n28155 , n28156 , n28157 , n28158 , n28159 , n28160 , n28161 , n28162 , n28163 , n28164 , n28165 , n28166 , n28167 , n28168 , n28169 , n28170 , n28171 , n28172 , n28173 , n28174 , n28175 , n28176 , n28177 , n28178 , n28179 , n28180 , n28181 , n28182 , n28183 , n28184 , n28185 , n28186 , n28187 , n28188 , n28189 , n28190 , n28191 , n28192 , n28193 , n28194 , n28195 , n28196 , n28197 , n28198 , n28199 , n28200 , n28201 , n28202 , n28203 , n28204 , n28205 , n28206 , n28207 , n28208 , n28209 , n28210 , n28211 , n28212 , n28213 , n28214 , n28215 , n28216 , n28217 , n28218 , n28219 , n28220 , n28221 , n28222 , n28223 , n28224 , n28225 , n28226 , n28227 , n28228 , n28229 , n28230 , n28231 , n28232 , n28233 , n28234 , n28235 , n28236 , n28237 , n28238 , n28239 , n28240 , n28241 , n28242 , n28243 , n28244 , n28245 , n28246 , n28247 , n28248 , n28249 , n28250 , n28251 , n28252 , n28253 , n28254 , n28255 , n28256 , n28257 , n28258 , n28259 , n28260 , n28261 , n28262 , n28263 , n28264 , n28265 , n28266 , n28267 , n28268 , n28269 , n28270 , n28271 , n28272 , n28273 , n28274 , n28275 , n28276 , n28277 , n28278 , n28279 , n28280 , n28281 , n28282 , n28283 , n28284 , n28285 , n28286 , n28287 , n28288 , n28289 , n28290 , n28291 , n28292 , n28293 , n28294 , n28295 , n28296 , n28297 , n28298 , n28299 , n28300 , n28301 , n28302 , n28303 , n28304 , n28305 , n28306 , n28307 , n28308 , n28309 , n28310 , n28311 , n28312 , n28313 , n28314 , n28315 , n28316 , n28317 , n28318 , n28319 , n28320 , n28321 , n28322 , n28323 , n28324 , n28325 , n28326 , n28327 , n28328 , n28329 , n28330 , n28331 , n28332 , n28333 , n28334 , n28335 , n28336 , n28337 , n28338 , n28339 , n28340 , n28341 , n28342 , n28343 , n28344 , n28345 , n28346 , n28347 , n28348 , n28349 , n28350 , n28351 , n28352 , n28353 , n28354 , n28355 , n28356 , n28357 , n28358 , n28359 , n28360 , n28361 , n28362 , n28363 , n28364 , n28365 , n28366 , n28367 , n28368 , n28369 , n28370 , n28371 , n28372 , n28373 , n28374 , n28375 , n28376 , n28377 , n28378 , n28379 , n28380 , n28381 , n28382 , n28383 , n28384 , n28385 , n28386 , n28387 , n28388 , n28389 , n28390 , n28391 , n28392 , n28393 , n28394 , n28395 , n28396 , n28397 , n28398 , n28399 , n28400 , n28401 , n28402 , n28403 , n28404 , n28405 , n28406 , n28407 , n28408 , n28409 , n28410 , n28411 , n28412 , n28413 , n28414 , n28415 , n28416 , n28417 , n28418 , n28419 , n28420 , n28421 , n28422 , n28423 , n28424 , n28425 , n28426 , n28427 , n28428 , n28429 , n28430 , n28431 , n28432 , n28433 , n28434 , n28435 , n28436 , n28437 , n28438 , n28439 , n28440 , n28441 , n28442 , n28443 , n28444 , n28445 , n28446 , n28447 , n28448 , n28449 , n28450 , n28451 , n28452 , n28453 , n28454 , n28455 , n28456 , n28457 , n28458 , n28459 , n28460 , n28461 , n28462 , n28463 , n28464 , n28465 , n28466 , n28467 , n28468 , n28469 , n28470 , n28471 , n28472 , n28473 , n28474 , n28475 , n28476 , n28477 , n28478 , n28479 , n28480 , n28481 , n28482 , n28483 , n28484 , n28485 , n28486 , n28487 , n28488 , n28489 , n28490 , n28491 , n28492 , n28493 , n28494 , n28495 , n28496 , n28497 , n28498 , n28499 , n28500 , n28501 , n28502 , n28503 , n28504 , n28505 , n28506 , n28507 , n28508 , n28509 , n28510 , n28511 , n28512 , n28513 , n28514 , n28515 , n28516 , n28517 , n28518 , n28519 , n28520 , n28521 , n28522 , n28523 , n28524 , n28525 , n28526 , n28527 , n28528 , n28529 , n28530 , n28531 , n28532 , n28533 , n28534 , n28535 , n28536 , n28537 , n28538 , n28539 , n28540 , n28541 , n28542 , n28543 , n28544 , n28545 , n28546 , n28547 , n28548 , n28549 , n28550 , n28551 , n28552 , n28553 , n28554 , n28555 , n28556 , n28557 , n28558 , n28559 , n28560 , n28561 , n28562 , n28563 , n28564 , n28565 , n28566 , n28567 , n28568 , n28569 , n28570 , n28571 , n28572 , n28573 , n28574 , n28575 , n28576 , n28577 , n28578 , n28579 , n28580 , n28581 , n28582 , n28583 , n28584 , n28585 , n28586 , n28587 , n28588 , n28589 , n28590 , n28591 , n28592 , n28593 , n28594 , n28595 , n28596 , n28597 , n28598 , n28599 , n28600 , n28601 , n28602 , n28603 , n28604 , n28605 , n28606 , n28607 , n28608 , n28609 , n28610 , n28611 , n28612 , n28613 , n28614 , n28615 , n28616 , n28617 , n28618 , n28619 , n28620 , n28621 , n28622 , n28623 , n28624 , n28625 , n28626 , n28627 , n28628 , n28629 , n28630 , n28631 , n28632 , n28633 , n28634 , n28635 , n28636 , n28637 , n28638 , n28639 , n28640 , n28641 , n28642 , n28643 , n28644 , n28645 , n28646 , n28647 , n28648 , n28649 , n28650 , n28651 , n28652 , n28653 , n28654 , n28655 , n28656 , n28657 , n28658 , n28659 , n28660 , n28661 , n28662 , n28663 , n28664 , n28665 , n28666 , n28667 , n28668 , n28669 , n28670 , n28671 , n28672 , n28673 , n28674 , n28675 , n28676 , n28677 , n28678 , n28679 , n28680 , n28681 , n28682 , n28683 , n28684 , n28685 , n28686 , n28687 , n28688 , n28689 , n28690 , n28691 , n28692 , n28693 , n28694 , n28695 , n28696 , n28697 , n28698 , n28699 , n28700 , n28701 , n28702 , n28703 , n28704 , n28705 , n28706 , n28707 , n28708 , n28709 , n28710 , n28711 , n28712 , n28713 , n28714 , n28715 , n28716 , n28717 , n28718 , n28719 , n28720 , n28721 , n28722 , n28723 , n28724 , n28725 , n28726 , n28727 , n28728 , n28729 , n28730 , n28731 , n28732 , n28733 , n28734 , n28735 , n28736 , n28737 , n28738 , n28739 , n28740 , n28741 , n28742 , n28743 , n28744 , n28745 , n28746 , n28747 , n28748 , n28749 , n28750 , n28751 , n28752 , n28753 , n28754 , n28755 , n28756 , n28757 , n28758 , n28759 , n28760 , n28761 , n28762 , n28763 , n28764 , n28765 , n28766 , n28767 , n28768 , n28769 , n28770 , n28771 , n28772 , n28773 , n28774 , n28775 , n28776 , n28777 , n28778 , n28779 , n28780 , n28781 , n28782 , n28783 , n28784 , n28785 , n28786 , n28787 , n28788 , n28789 , n28790 , n28791 , n28792 , n28793 , n28794 , n28795 , n28796 , n28797 , n28798 , n28799 , n28800 , n28801 , n28802 , n28803 , n28804 , n28805 , n28806 , n28807 , n28808 , n28809 , n28810 , n28811 , n28812 , n28813 , n28814 , n28815 , n28816 , n28817 , n28818 , n28819 , n28820 , n28821 , n28822 , n28823 , n28824 , n28825 , n28826 , n28827 , n28828 , n28829 , n28830 , n28831 , n28832 , n28833 , n28834 , n28835 , n28836 , n28837 , n28838 , n28839 , n28840 , n28841 , n28842 , n28843 , n28844 , n28845 , n28846 , n28847 , n28848 , n28849 , n28850 , n28851 , n28852 , n28853 , n28854 , n28855 , n28856 , n28857 , n28858 , n28859 , n28860 , n28861 , n28862 , n28863 , n28864 , n28865 , n28866 , n28867 , n28868 , n28869 , n28870 , n28871 , n28872 , n28873 , n28874 , n28875 , n28876 , n28877 , n28878 , n28879 , n28880 , n28881 , n28882 , n28883 , n28884 , n28885 , n28886 , n28887 , n28888 , n28889 , n28890 , n28891 , n28892 , n28893 , n28894 , n28895 , n28896 , n28897 , n28898 , n28899 , n28900 , n28901 , n28902 , n28903 , n28904 , n28905 , n28906 , n28907 , n28908 , n28909 , n28910 , n28911 , n28912 , n28913 , n28914 , n28915 , n28916 , n28917 , n28918 , n28919 , n28920 , n28921 , n28922 , n28923 , n28924 , n28925 , n28926 , n28927 , n28928 , n28929 , n28930 , n28931 , n28932 , n28933 , n28934 , n28935 , n28936 , n28937 , n28938 , n28939 , n28940 , n28941 , n28942 , n28943 , n28944 , n28945 , n28946 , n28947 , n28948 , n28949 , n28950 , n28951 , n28952 , n28953 , n28954 , n28955 , n28956 , n28957 , n28958 , n28959 , n28960 , n28961 , n28962 , n28963 , n28964 , n28965 , n28966 , n28967 , n28968 , n28969 , n28970 , n28971 , n28972 , n28973 , n28974 , n28975 , n28976 , n28977 , n28978 , n28979 , n28980 , n28981 , n28982 , n28983 , n28984 , n28985 , n28986 , n28987 , n28988 , n28989 , n28990 , n28991 , n28992 , n28993 , n28994 , n28995 , n28996 , n28997 , n28998 , n28999 , n29000 , n29001 , n29002 , n29003 , n29004 , n29005 , n29006 , n29007 , n29008 , n29009 , n29010 , n29011 , n29012 , n29013 , n29014 , n29015 , n29016 , n29017 , n29018 , n29019 , n29020 , n29021 , n29022 , n29023 , n29024 , n29025 , n29026 , n29027 , n29028 , n29029 , n29030 , n29031 , n29032 , n29033 , n29034 , n29035 , n29036 , n29037 , n29038 , n29039 , n29040 , n29041 , n29042 , n29043 , n29044 , n29045 , n29046 , n29047 , n29048 , n29049 , n29050 , n29051 , n29052 , n29053 , n29054 , n29055 , n29056 , n29057 , n29058 , n29059 , n29060 , n29061 , n29062 , n29063 , n29064 , n29065 , n29066 , n29067 , n29068 , n29069 , n29070 , n29071 , n29072 , n29073 , n29074 , n29075 , n29076 , n29077 , n29078 , n29079 , n29080 , n29081 , n29082 , n29083 , n29084 , n29085 , n29086 , n29087 , n29088 , n29089 , n29090 , n29091 , n29092 , n29093 , n29094 , n29095 , n29096 , n29097 , n29098 , n29099 , n29100 , n29101 , n29102 , n29103 , n29104 , n29105 , n29106 , n29107 , n29108 , n29109 , n29110 , n29111 , n29112 , n29113 , n29114 , n29115 , n29116 , n29117 , n29118 , n29119 , n29120 , n29121 , n29122 , n29123 , n29124 , n29125 , n29126 , n29127 , n29128 , n29129 , n29130 , n29131 , n29132 , n29133 , n29134 , n29135 , n29136 , n29137 , n29138 , n29139 , n29140 , n29141 , n29142 , n29143 , n29144 , n29145 , n29146 , n29147 , n29148 , n29149 , n29150 , n29151 , n29152 , n29153 , n29154 , n29155 , n29156 , n29157 , n29158 , n29159 , n29160 , n29161 , n29162 , n29163 , n29164 , n29165 , n29166 , n29167 , n29168 , n29169 , n29170 , n29171 , n29172 , n29173 , n29174 , n29175 , n29176 , n29177 , n29178 , n29179 , n29180 , n29181 , n29182 , n29183 , n29184 , n29185 , n29186 , n29187 , n29188 , n29189 , n29190 , n29191 , n29192 , n29193 , n29194 , n29195 , n29196 , n29197 , n29198 , n29199 , n29200 , n29201 , n29202 , n29203 , n29204 , n29205 , n29206 , n29207 , n29208 , n29209 , n29210 , n29211 , n29212 , n29213 , n29214 , n29215 , n29216 , n29217 , n29218 , n29219 , n29220 , n29221 , n29222 , n29223 , n29224 , n29225 , n29226 , n29227 , n29228 , n29229 , n29230 , n29231 , n29232 , n29233 , n29234 , n29235 , n29236 , n29237 , n29238 , n29239 , n29240 , n29241 , n29242 , n29243 , n29244 , n29245 , n29246 , n29247 , n29248 , n29249 , n29250 , n29251 , n29252 , n29253 , n29254 , n29255 , n29256 , n29257 , n29258 , n29259 , n29260 , n29261 , n29262 , n29263 , n29264 , n29265 , n29266 , n29267 , n29268 , n29269 , n29270 , n29271 , n29272 , n29273 , n29274 , n29275 , n29276 , n29277 , n29278 , n29279 , n29280 , n29281 , n29282 , n29283 , n29284 , n29285 , n29286 , n29287 , n29288 , n29289 , n29290 , n29291 , n29292 , n29293 , n29294 , n29295 , n29296 , n29297 , n29298 , n29299 , n29300 , n29301 , n29302 , n29303 , n29304 , n29305 , n29306 , n29307 , n29308 , n29309 , n29310 , n29311 , n29312 , n29313 , n29314 , n29315 , n29316 , n29317 , n29318 , n29319 , n29320 , n29321 , n29322 , n29323 , n29324 , n29325 , n29326 , n29327 , n29328 , n29329 , n29330 , n29331 , n29332 , n29333 , n29334 , n29335 , n29336 , n29337 , n29338 , n29339 , n29340 , n29341 , n29342 , n29343 , n29344 , n29345 , n29346 , n29347 , n29348 , n29349 , n29350 , n29351 , n29352 , n29353 , n29354 , n29355 , n29356 , n29357 , n29358 , n29359 , n29360 , n29361 , n29362 , n29363 , n29364 , n29365 , n29366 , n29367 , n29368 , n29369 , n29370 , n29371 , n29372 , n29373 , n29374 , n29375 , n29376 , n29377 , n29378 , n29379 , n29380 , n29381 , n29382 , n29383 , n29384 , n29385 , n29386 , n29387 , n29388 , n29389 , n29390 , n29391 , n29392 , n29393 , n29394 , n29395 , n29396 , n29397 , n29398 , n29399 , n29400 , n29401 , n29402 , n29403 , n29404 , n29405 , n29406 , n29407 , n29408 , n29409 , n29410 , n29411 , n29412 , n29413 , n29414 , n29415 , n29416 , n29417 , n29418 , n29419 , n29420 , n29421 , n29422 , n29423 , n29424 , n29425 , n29426 , n29427 , n29428 , n29429 , n29430 , n29431 , n29432 , n29433 , n29434 , n29435 , n29436 , n29437 , n29438 , n29439 , n29440 , n29441 , n29442 , n29443 , n29444 , n29445 , n29446 , n29447 , n29448 , n29449 , n29450 , n29451 , n29452 , n29453 , n29454 , n29455 , n29456 , n29457 , n29458 , n29459 , n29460 , n29461 , n29462 , n29463 , n29464 , n29465 , n29466 , n29467 , n29468 , n29469 , n29470 , n29471 , n29472 , n29473 , n29474 , n29475 , n29476 , n29477 , n29478 , n29479 , n29480 , n29481 , n29482 , n29483 , n29484 , n29485 , n29486 , n29487 , n29488 , n29489 , n29490 , n29491 , n29492 , n29493 , n29494 , n29495 , n29496 , n29497 , n29498 , n29499 , n29500 , n29501 , n29502 , n29503 , n29504 , n29505 , n29506 , n29507 , n29508 , n29509 , n29510 , n29511 , n29512 , n29513 , n29514 , n29515 , n29516 , n29517 , n29518 , n29519 , n29520 , n29521 , n29522 , n29523 , n29524 , n29525 , n29526 , n29527 , n29528 , n29529 , n29530 , n29531 , n29532 , n29533 , n29534 , n29535 , n29536 , n29537 , n29538 , n29539 , n29540 , n29541 , n29542 , n29543 , n29544 , n29545 , n29546 , n29547 , n29548 , n29549 , n29550 , n29551 , n29552 , n29553 , n29554 , n29555 , n29556 , n29557 , n29558 , n29559 , n29560 , n29561 , n29562 , n29563 , n29564 , n29565 , n29566 , n29567 , n29568 , n29569 , n29570 , n29571 , n29572 , n29573 , n29574 , n29575 , n29576 , n29577 , n29578 , n29579 , n29580 , n29581 , n29582 , n29583 , n29584 , n29585 , n29586 , n29587 , n29588 , n29589 , n29590 , n29591 , n29592 , n29593 , n29594 , n29595 , n29596 , n29597 , n29598 , n29599 , n29600 , n29601 , n29602 , n29603 , n29604 , n29605 , n29606 , n29607 , n29608 , n29609 , n29610 , n29611 , n29612 , n29613 , n29614 , n29615 , n29616 , n29617 , n29618 , n29619 , n29620 , n29621 , n29622 , n29623 , n29624 , n29625 , n29626 , n29627 , n29628 , n29629 , n29630 , n29631 , n29632 , n29633 , n29634 , n29635 , n29636 , n29637 , n29638 , n29639 , n29640 , n29641 , n29642 , n29643 , n29644 , n29645 , n29646 , n29647 , n29648 , n29649 , n29650 , n29651 , n29652 , n29653 , n29654 , n29655 , n29656 , n29657 , n29658 , n29659 , n29660 , n29661 , n29662 , n29663 , n29664 , n29665 , n29666 , n29667 , n29668 , n29669 , n29670 , n29671 , n29672 , n29673 , n29674 , n29675 , n29676 , n29677 , n29678 , n29679 , n29680 , n29681 , n29682 , n29683 , n29684 , n29685 , n29686 , n29687 , n29688 , n29689 , n29690 , n29691 , n29692 , n29693 , n29694 , n29695 , n29696 , n29697 , n29698 , n29699 , n29700 , n29701 , n29702 , n29703 , n29704 , n29705 , n29706 , n29707 , n29708 , n29709 , n29710 , n29711 , n29712 , n29713 , n29714 , n29715 , n29716 , n29717 , n29718 , n29719 , n29720 , n29721 , n29722 , n29723 , n29724 , n29725 , n29726 , n29727 , n29728 , n29729 , n29730 , n29731 , n29732 , n29733 , n29734 , n29735 , n29736 , n29737 , n29738 , n29739 , n29740 , n29741 , n29742 , n29743 , n29744 , n29745 , n29746 , n29747 , n29748 , n29749 , n29750 , n29751 , n29752 , n29753 , n29754 , n29755 , n29756 , n29757 , n29758 , n29759 , n29760 , n29761 , n29762 , n29763 , n29764 , n29765 , n29766 , n29767 , n29768 , n29769 , n29770 , n29771 , n29772 , n29773 , n29774 , n29775 , n29776 , n29777 , n29778 , n29779 , n29780 , n29781 , n29782 , n29783 , n29784 , n29785 , n29786 , n29787 , n29788 , n29789 , n29790 , n29791 , n29792 , n29793 , n29794 , n29795 , n29796 , n29797 , n29798 , n29799 , n29800 , n29801 , n29802 , n29803 , n29804 , n29805 , n29806 , n29807 , n29808 , n29809 , n29810 , n29811 , n29812 , n29813 , n29814 , n29815 , n29816 , n29817 , n29818 , n29819 , n29820 , n29821 , n29822 , n29823 , n29824 , n29825 , n29826 , n29827 , n29828 , n29829 , n29830 , n29831 , n29832 , n29833 , n29834 , n29835 , n29836 , n29837 , n29838 , n29839 , n29840 , n29841 , n29842 , n29843 , n29844 , n29845 , n29846 , n29847 , n29848 , n29849 , n29850 , n29851 , n29852 , n29853 , n29854 , n29855 , n29856 , n29857 , n29858 , n29859 , n29860 , n29861 , n29862 , n29863 , n29864 , n29865 , n29866 , n29867 , n29868 , n29869 , n29870 , n29871 , n29872 , n29873 , n29874 , n29875 , n29876 , n29877 , n29878 , n29879 , n29880 , n29881 , n29882 , n29883 , n29884 , n29885 , n29886 , n29887 , n29888 , n29889 , n29890 , n29891 , n29892 , n29893 , n29894 , n29895 , n29896 , n29897 , n29898 , n29899 , n29900 , n29901 , n29902 , n29903 , n29904 , n29905 , n29906 , n29907 , n29908 , n29909 , n29910 , n29911 , n29912 , n29913 , n29914 , n29915 , n29916 , n29917 , n29918 , n29919 , n29920 , n29921 , n29922 , n29923 , n29924 , n29925 , n29926 , n29927 , n29928 , n29929 , n29930 , n29931 , n29932 , n29933 , n29934 , n29935 , n29936 , n29937 , n29938 , n29939 , n29940 , n29941 , n29942 , n29943 , n29944 , n29945 , n29946 , n29947 , n29948 , n29949 , n29950 , n29951 , n29952 , n29953 , n29954 , n29955 , n29956 , n29957 , n29958 , n29959 , n29960 , n29961 , n29962 , n29963 , n29964 , n29965 , n29966 , n29967 , n29968 , n29969 , n29970 , n29971 , n29972 , n29973 , n29974 , n29975 , n29976 , n29977 , n29978 , n29979 , n29980 , n29981 , n29982 , n29983 , n29984 , n29985 , n29986 , n29987 , n29988 , n29989 , n29990 , n29991 , n29992 , n29993 , n29994 , n29995 , n29996 , n29997 , n29998 , n29999 , n30000 , n30001 , n30002 , n30003 , n30004 , n30005 , n30006 , n30007 , n30008 , n30009 , n30010 , n30011 , n30012 , n30013 , n30014 , n30015 , n30016 , n30017 , n30018 , n30019 , n30020 , n30021 , n30022 , n30023 , n30024 , n30025 , n30026 , n30027 , n30028 , n30029 , n30030 , n30031 , n30032 , n30033 , n30034 , n30035 , n30036 , n30037 , n30038 , n30039 , n30040 , n30041 , n30042 , n30043 , n30044 , n30045 , n30046 , n30047 , n30048 , n30049 , n30050 , n30051 , n30052 , n30053 , n30054 , n30055 , n30056 , n30057 , n30058 , n30059 , n30060 , n30061 , n30062 , n30063 , n30064 , n30065 , n30066 , n30067 , n30068 , n30069 , n30070 , n30071 , n30072 , n30073 , n30074 , n30075 , n30076 , n30077 , n30078 , n30079 , n30080 , n30081 , n30082 , n30083 , n30084 , n30085 , n30086 , n30087 , n30088 , n30089 , n30090 , n30091 , n30092 , n30093 , n30094 , n30095 , n30096 , n30097 , n30098 , n30099 , n30100 , n30101 , n30102 , n30103 , n30104 , n30105 , n30106 , n30107 , n30108 , n30109 , n30110 , n30111 , n30112 , n30113 , n30114 , n30115 , n30116 , n30117 , n30118 , n30119 , n30120 , n30121 , n30122 , n30123 , n30124 , n30125 , n30126 , n30127 , n30128 , n30129 , n30130 , n30131 , n30132 , n30133 , n30134 , n30135 , n30136 , n30137 , n30138 , n30139 , n30140 , n30141 , n30142 , n30143 , n30144 , n30145 , n30146 , n30147 , n30148 , n30149 , n30150 , n30151 , n30152 , n30153 , n30154 , n30155 , n30156 , n30157 , n30158 , n30159 , n30160 , n30161 , n30162 , n30163 , n30164 , n30165 , n30166 , n30167 , n30168 , n30169 , n30170 , n30171 , n30172 , n30173 , n30174 , n30175 , n30176 , n30177 , n30178 , n30179 , n30180 , n30181 , n30182 , n30183 , n30184 , n30185 , n30186 , n30187 , n30188 , n30189 , n30190 , n30191 , n30192 , n30193 , n30194 , n30195 , n30196 , n30197 , n30198 , n30199 , n30200 , n30201 , n30202 , n30203 , n30204 , n30205 , n30206 , n30207 , n30208 , n30209 , n30210 , n30211 , n30212 , n30213 , n30214 , n30215 , n30216 , n30217 , n30218 , n30219 , n30220 , n30221 , n30222 , n30223 , n30224 , n30225 , n30226 , n30227 , n30228 , n30229 , n30230 , n30231 , n30232 , n30233 , n30234 , n30235 , n30236 , n30237 , n30238 , n30239 , n30240 , n30241 , n30242 , n30243 , n30244 , n30245 , n30246 , n30247 , n30248 , n30249 , n30250 , n30251 , n30252 , n30253 , n30254 , n30255 , n30256 , n30257 , n30258 , n30259 , n30260 , n30261 , n30262 , n30263 , n30264 , n30265 , n30266 , n30267 , n30268 , n30269 , n30270 , n30271 , n30272 , n30273 , n30274 , n30275 , n30276 , n30277 , n30278 , n30279 , n30280 , n30281 , n30282 , n30283 , n30284 , n30285 , n30286 , n30287 , n30288 , n30289 , n30290 , n30291 , n30292 , n30293 , n30294 , n30295 , n30296 , n30297 , n30298 , n30299 , n30300 , n30301 , n30302 , n30303 , n30304 , n30305 , n30306 , n30307 , n30308 , n30309 , n30310 , n30311 , n30312 , n30313 , n30314 , n30315 , n30316 , n30317 , n30318 , n30319 , n30320 , n30321 , n30322 , n30323 , n30324 , n30325 , n30326 , n30327 , n30328 , n30329 , n30330 , n30331 , n30332 , n30333 , n30334 , n30335 , n30336 , n30337 , n30338 , n30339 , n30340 , n30341 , n30342 , n30343 , n30344 , n30345 , n30346 , n30347 , n30348 , n30349 , n30350 , n30351 , n30352 , n30353 , n30354 , n30355 , n30356 , n30357 , n30358 , n30359 , n30360 , n30361 , n30362 , n30363 , n30364 , n30365 , n30366 , n30367 , n30368 , n30369 , n30370 , n30371 , n30372 , n30373 , n30374 , n30375 , n30376 , n30377 , n30378 , n30379 , n30380 , n30381 , n30382 , n30383 , n30384 , n30385 , n30386 , n30387 , n30388 , n30389 , n30390 , n30391 , n30392 , n30393 , n30394 , n30395 , n30396 , n30397 , n30398 , n30399 , n30400 , n30401 , n30402 , n30403 , n30404 , n30405 , n30406 , n30407 , n30408 , n30409 , n30410 , n30411 , n30412 , n30413 , n30414 , n30415 , n30416 , n30417 , n30418 , n30419 , n30420 , n30421 , n30422 , n30423 , n30424 , n30425 , n30426 , n30427 , n30428 , n30429 , n30430 , n30431 , n30432 , n30433 , n30434 , n30435 , n30436 , n30437 , n30438 , n30439 , n30440 , n30441 , n30442 , n30443 , n30444 , n30445 , n30446 , n30447 , n30448 , n30449 , n30450 , n30451 , n30452 , n30453 , n30454 , n30455 , n30456 , n30457 , n30458 , n30459 , n30460 , n30461 , n30462 , n30463 , n30464 , n30465 , n30466 , n30467 , n30468 , n30469 , n30470 , n30471 , n30472 , n30473 , n30474 , n30475 , n30476 , n30477 , n30478 , n30479 , n30480 , n30481 , n30482 , n30483 , n30484 , n30485 , n30486 , n30487 , n30488 , n30489 , n30490 , n30491 , n30492 , n30493 , n30494 , n30495 , n30496 , n30497 , n30498 , n30499 , n30500 , n30501 , n30502 , n30503 , n30504 , n30505 , n30506 , n30507 , n30508 , n30509 , n30510 , n30511 , n30512 , n30513 , n30514 , n30515 , n30516 , n30517 , n30518 , n30519 , n30520 , n30521 , n30522 , n30523 , n30524 , n30525 , n30526 , n30527 , n30528 , n30529 , n30530 , n30531 , n30532 , n30533 , n30534 , n30535 , n30536 , n30537 , n30538 , n30539 , n30540 , n30541 , n30542 , n30543 , n30544 , n30545 , n30546 , n30547 , n30548 , n30549 , n30550 , n30551 , n30552 , n30553 , n30554 , n30555 , n30556 , n30557 , n30558 , n30559 , n30560 , n30561 , n30562 , n30563 , n30564 , n30565 , n30566 , n30567 , n30568 , n30569 , n30570 , n30571 , n30572 , n30573 , n30574 , n30575 , n30576 , n30577 , n30578 , n30579 , n30580 , n30581 , n30582 , n30583 , n30584 , n30585 , n30586 , n30587 , n30588 , n30589 , n30590 , n30591 , n30592 , n30593 , n30594 , n30595 , n30596 , n30597 , n30598 , n30599 , n30600 , n30601 , n30602 , n30603 , n30604 , n30605 , n30606 , n30607 , n30608 , n30609 , n30610 , n30611 , n30612 , n30613 , n30614 , n30615 , n30616 , n30617 , n30618 , n30619 , n30620 , n30621 , n30622 , n30623 , n30624 , n30625 , n30626 , n30627 , n30628 , n30629 , n30630 , n30631 , n30632 , n30633 , n30634 , n30635 , n30636 , n30637 , n30638 , n30639 , n30640 , n30641 , n30642 , n30643 , n30644 , n30645 , n30646 , n30647 , n30648 , n30649 , n30650 , n30651 , n30652 , n30653 , n30654 , n30655 , n30656 , n30657 , n30658 , n30659 , n30660 , n30661 , n30662 , n30663 , n30664 , n30665 , n30666 , n30667 , n30668 , n30669 , n30670 , n30671 , n30672 , n30673 , n30674 , n30675 , n30676 , n30677 , n30678 , n30679 , n30680 , n30681 , n30682 , n30683 , n30684 , n30685 , n30686 , n30687 , n30688 , n30689 , n30690 , n30691 , n30692 , n30693 , n30694 , n30695 , n30696 , n30697 , n30698 , n30699 , n30700 , n30701 , n30702 , n30703 , n30704 , n30705 , n30706 , n30707 , n30708 , n30709 , n30710 , n30711 , n30712 , n30713 , n30714 , n30715 , n30716 , n30717 , n30718 , n30719 , n30720 , n30721 , n30722 , n30723 , n30724 , n30725 , n30726 , n30727 , n30728 , n30729 , n30730 , n30731 , n30732 , n30733 , n30734 , n30735 , n30736 , n30737 , n30738 , n30739 , n30740 , n30741 , n30742 , n30743 , n30744 , n30745 , n30746 , n30747 , n30748 , n30749 , n30750 , n30751 , n30752 , n30753 , n30754 , n30755 , n30756 , n30757 , n30758 , n30759 , n30760 , n30761 , n30762 , n30763 , n30764 , n30765 , n30766 , n30767 , n30768 , n30769 , n30770 , n30771 , n30772 , n30773 , n30774 , n30775 , n30776 , n30777 , n30778 , n30779 , n30780 , n30781 , n30782 , n30783 , n30784 , n30785 , n30786 , n30787 , n30788 , n30789 , n30790 , n30791 , n30792 , n30793 , n30794 , n30795 , n30796 , n30797 , n30798 , n30799 , n30800 , n30801 , n30802 , n30803 , n30804 , n30805 , n30806 , n30807 , n30808 , n30809 , n30810 , n30811 , n30812 , n30813 , n30814 , n30815 , n30816 , n30817 , n30818 , n30819 , n30820 , n30821 , n30822 , n30823 , n30824 , n30825 , n30826 , n30827 , n30828 , n30829 , n30830 , n30831 , n30832 , n30833 , n30834 , n30835 , n30836 , n30837 , n30838 , n30839 , n30840 , n30841 , n30842 , n30843 , n30844 , n30845 , n30846 , n30847 , n30848 , n30849 , n30850 , n30851 , n30852 , n30853 , n30854 , n30855 , n30856 , n30857 , n30858 , n30859 , n30860 , n30861 , n30862 , n30863 , n30864 , n30865 , n30866 , n30867 , n30868 , n30869 , n30870 , n30871 , n30872 , n30873 , n30874 , n30875 , n30876 , n30877 , n30878 , n30879 , n30880 , n30881 , n30882 , n30883 , n30884 , n30885 , n30886 , n30887 , n30888 , n30889 , n30890 , n30891 , n30892 , n30893 , n30894 , n30895 , n30896 , n30897 , n30898 , n30899 , n30900 , n30901 , n30902 , n30903 , n30904 , n30905 , n30906 , n30907 , n30908 , n30909 , n30910 , n30911 , n30912 , n30913 , n30914 , n30915 , n30916 , n30917 , n30918 , n30919 , n30920 , n30921 , n30922 , n30923 , n30924 , n30925 , n30926 , n30927 , n30928 , n30929 , n30930 , n30931 , n30932 , n30933 , n30934 , n30935 , n30936 , n30937 , n30938 , n30939 , n30940 , n30941 , n30942 , n30943 , n30944 , n30945 , n30946 , n30947 , n30948 , n30949 , n30950 , n30951 , n30952 , n30953 , n30954 , n30955 , n30956 , n30957 , n30958 , n30959 , n30960 , n30961 , n30962 , n30963 , n30964 , n30965 , n30966 , n30967 , n30968 , n30969 , n30970 , n30971 , n30972 , n30973 , n30974 , n30975 , n30976 , n30977 , n30978 , n30979 , n30980 , n30981 , n30982 , n30983 , n30984 , n30985 , n30986 , n30987 , n30988 , n30989 , n30990 , n30991 , n30992 , n30993 , n30994 , n30995 , n30996 , n30997 , n30998 , n30999 , n31000 , n31001 , n31002 , n31003 , n31004 , n31005 , n31006 , n31007 , n31008 , n31009 , n31010 , n31011 , n31012 , n31013 , n31014 , n31015 , n31016 , n31017 , n31018 , n31019 , n31020 , n31021 , n31022 , n31023 , n31024 , n31025 , n31026 , n31027 , n31028 , n31029 , n31030 , n31031 , n31032 , n31033 , n31034 , n31035 , n31036 , n31037 , n31038 , n31039 , n31040 , n31041 , n31042 , n31043 , n31044 , n31045 , n31046 , n31047 , n31048 , n31049 , n31050 , n31051 , n31052 , n31053 , n31054 , n31055 , n31056 , n31057 , n31058 , n31059 , n31060 , n31061 , n31062 , n31063 , n31064 , n31065 , n31066 , n31067 , n31068 , n31069 , n31070 , n31071 , n31072 , n31073 , n31074 , n31075 , n31076 , n31077 , n31078 , n31079 , n31080 , n31081 , n31082 , n31083 , n31084 , n31085 , n31086 , n31087 , n31088 , n31089 , n31090 , n31091 , n31092 , n31093 , n31094 , n31095 , n31096 , n31097 , n31098 , n31099 , n31100 , n31101 , n31102 , n31103 , n31104 , n31105 , n31106 , n31107 , n31108 , n31109 , n31110 , n31111 , n31112 , n31113 , n31114 , n31115 , n31116 , n31117 , n31118 , n31119 , n31120 , n31121 , n31122 , n31123 , n31124 , n31125 , n31126 , n31127 , n31128 , n31129 , n31130 , n31131 , n31132 , n31133 , n31134 , n31135 , n31136 , n31137 , n31138 , n31139 , n31140 , n31141 , n31142 , n31143 , n31144 , n31145 , n31146 , n31147 , n31148 , n31149 , n31150 , n31151 , n31152 , n31153 , n31154 , n31155 , n31156 , n31157 , n31158 , n31159 , n31160 , n31161 , n31162 , n31163 , n31164 , n31165 , n31166 , n31167 , n31168 , n31169 , n31170 , n31171 , n31172 , n31173 , n31174 , n31175 , n31176 , n31177 , n31178 , n31179 , n31180 , n31181 , n31182 , n31183 , n31184 , n31185 , n31186 , n31187 , n31188 , n31189 , n31190 , n31191 , n31192 , n31193 , n31194 , n31195 , n31196 , n31197 , n31198 , n31199 , n31200 , n31201 , n31202 , n31203 , n31204 , n31205 , n31206 , n31207 , n31208 , n31209 , n31210 , n31211 , n31212 , n31213 , n31214 , n31215 , n31216 , n31217 , n31218 , n31219 , n31220 , n31221 , n31222 , n31223 , n31224 , n31225 , n31226 , n31227 , n31228 , n31229 , n31230 , n31231 , n31232 , n31233 , n31234 , n31235 , n31236 , n31237 , n31238 , n31239 , n31240 , n31241 , n31242 , n31243 , n31244 , n31245 , n31246 , n31247 , n31248 , n31249 , n31250 , n31251 , n31252 , n31253 , n31254 , n31255 , n31256 , n31257 , n31258 , n31259 , n31260 , n31261 , n31262 , n31263 , n31264 , n31265 , n31266 , n31267 , n31268 , n31269 , n31270 , n31271 , n31272 , n31273 , n31274 , n31275 , n31276 , n31277 , n31278 , n31279 , n31280 , n31281 , n31282 , n31283 , n31284 , n31285 , n31286 , n31287 , n31288 , n31289 , n31290 , n31291 , n31292 , n31293 , n31294 , n31295 , n31296 , n31297 , n31298 , n31299 , n31300 , n31301 , n31302 , n31303 , n31304 , n31305 , n31306 , n31307 , n31308 , n31309 , n31310 , n31311 , n31312 , n31313 , n31314 , n31315 , n31316 , n31317 , n31318 , n31319 , n31320 , n31321 , n31322 , n31323 , n31324 , n31325 , n31326 , n31327 , n31328 , n31329 , n31330 , n31331 , n31332 , n31333 , n31334 , n31335 , n31336 , n31337 , n31338 , n31339 , n31340 , n31341 , n31342 , n31343 , n31344 , n31345 , n31346 , n31347 , n31348 , n31349 , n31350 , n31351 , n31352 , n31353 , n31354 , n31355 , n31356 , n31357 , n31358 , n31359 , n31360 , n31361 , n31362 , n31363 , n31364 , n31365 , n31366 , n31367 , n31368 , n31369 , n31370 , n31371 , n31372 , n31373 , n31374 , n31375 , n31376 , n31377 , n31378 , n31379 , n31380 , n31381 , n31382 , n31383 , n31384 , n31385 , n31386 , n31387 , n31388 , n31389 , n31390 , n31391 , n31392 , n31393 , n31394 , n31395 , n31396 , n31397 , n31398 , n31399 , n31400 , n31401 , n31402 , n31403 , n31404 , n31405 , n31406 , n31407 , n31408 , n31409 , n31410 , n31411 , n31412 , n31413 , n31414 , n31415 , n31416 , n31417 , n31418 , n31419 , n31420 , n31421 , n31422 , n31423 , n31424 , n31425 , n31426 , n31427 , n31428 , n31429 , n31430 , n31431 , n31432 , n31433 , n31434 , n31435 , n31436 , n31437 , n31438 , n31439 , n31440 , n31441 , n31442 , n31443 , n31444 , n31445 , n31446 , n31447 , n31448 , n31449 , n31450 , n31451 , n31452 , n31453 , n31454 , n31455 , n31456 , n31457 , n31458 , n31459 , n31460 , n31461 , n31462 , n31463 , n31464 , n31465 , n31466 , n31467 , n31468 , n31469 , n31470 , n31471 , n31472 , n31473 , n31474 , n31475 , n31476 , n31477 , n31478 , n31479 , n31480 , n31481 , n31482 , n31483 , n31484 , n31485 , n31486 , n31487 , n31488 , n31489 , n31490 , n31491 , n31492 , n31493 , n31494 , n31495 , n31496 , n31497 , n31498 , n31499 , n31500 , n31501 , n31502 , n31503 , n31504 , n31505 , n31506 , n31507 , n31508 , n31509 , n31510 , n31511 , n31512 , n31513 , n31514 , n31515 , n31516 , n31517 , n31518 , n31519 , n31520 , n31521 , n31522 , n31523 , n31524 , n31525 , n31526 , n31527 , n31528 , n31529 , n31530 , n31531 , n31532 , n31533 , n31534 , n31535 , n31536 , n31537 , n31538 , n31539 , n31540 , n31541 , n31542 , n31543 , n31544 , n31545 , n31546 , n31547 , n31548 , n31549 , n31550 , n31551 , n31552 , n31553 , n31554 , n31555 , n31556 , n31557 , n31558 , n31559 , n31560 , n31561 , n31562 , n31563 , n31564 , n31565 , n31566 , n31567 , n31568 , n31569 , n31570 , n31571 , n31572 , n31573 , n31574 , n31575 , n31576 , n31577 , n31578 , n31579 , n31580 , n31581 , n31582 , n31583 , n31584 , n31585 , n31586 , n31587 , n31588 , n31589 , n31590 , n31591 , n31592 , n31593 , n31594 , n31595 , n31596 , n31597 , n31598 , n31599 , n31600 , n31601 , n31602 , n31603 , n31604 , n31605 , n31606 , n31607 , n31608 , n31609 , n31610 , n31611 , n31612 , n31613 , n31614 , n31615 , n31616 , n31617 , n31618 , n31619 , n31620 , n31621 , n31622 , n31623 , n31624 , n31625 , n31626 , n31627 , n31628 , n31629 , n31630 , n31631 , n31632 , n31633 , n31634 , n31635 , n31636 , n31637 , n31638 , n31639 , n31640 , n31641 , n31642 , n31643 , n31644 , n31645 , n31646 , n31647 , n31648 , n31649 , n31650 , n31651 , n31652 , n31653 , n31654 , n31655 , n31656 , n31657 , n31658 , n31659 , n31660 , n31661 , n31662 , n31663 , n31664 , n31665 , n31666 , n31667 , n31668 , n31669 , n31670 , n31671 , n31672 , n31673 , n31674 , n31675 , n31676 , n31677 , n31678 , n31679 , n31680 , n31681 , n31682 , n31683 , n31684 , n31685 , n31686 , n31687 , n31688 , n31689 , n31690 , n31691 , n31692 , n31693 , n31694 , n31695 , n31696 , n31697 , n31698 , n31699 , n31700 , n31701 , n31702 , n31703 , n31704 , n31705 , n31706 , n31707 , n31708 , n31709 , n31710 , n31711 , n31712 , n31713 , n31714 , n31715 , n31716 , n31717 , n31718 , n31719 , n31720 , n31721 , n31722 , n31723 , n31724 , n31725 , n31726 , n31727 , n31728 , n31729 , n31730 , n31731 , n31732 , n31733 , n31734 , n31735 , n31736 , n31737 , n31738 , n31739 , n31740 , n31741 , n31742 , n31743 , n31744 , n31745 , n31746 , n31747 , n31748 , n31749 , n31750 , n31751 , n31752 , n31753 , n31754 , n31755 , n31756 , n31757 , n31758 , n31759 , n31760 , n31761 , n31762 , n31763 , n31764 , n31765 , n31766 , n31767 , n31768 , n31769 , n31770 , n31771 , n31772 , n31773 , n31774 , n31775 , n31776 , n31777 , n31778 , n31779 , n31780 , n31781 , n31782 , n31783 , n31784 , n31785 , n31786 , n31787 , n31788 , n31789 , n31790 , n31791 , n31792 , n31793 , n31794 , n31795 , n31796 , n31797 , n31798 , n31799 , n31800 , n31801 , n31802 , n31803 , n31804 , n31805 , n31806 , n31807 , n31808 , n31809 , n31810 , n31811 , n31812 , n31813 , n31814 , n31815 , n31816 , n31817 , n31818 , n31819 , n31820 , n31821 , n31822 , n31823 , n31824 , n31825 , n31826 , n31827 , n31828 , n31829 , n31830 , n31831 , n31832 , n31833 , n31834 , n31835 , n31836 , n31837 , n31838 , n31839 , n31840 , n31841 , n31842 , n31843 , n31844 , n31845 , n31846 , n31847 , n31848 , n31849 , n31850 , n31851 , n31852 , n31853 , n31854 , n31855 , n31856 , n31857 , n31858 , n31859 , n31860 , n31861 , n31862 , n31863 , n31864 , n31865 , n31866 , n31867 , n31868 , n31869 , n31870 , n31871 , n31872 , n31873 , n31874 , n31875 , n31876 , n31877 , n31878 , n31879 , n31880 , n31881 , n31882 , n31883 , n31884 , n31885 , n31886 , n31887 , n31888 , n31889 , n31890 , n31891 , n31892 , n31893 , n31894 , n31895 , n31896 , n31897 , n31898 , n31899 , n31900 , n31901 , n31902 , n31903 , n31904 , n31905 , n31906 , n31907 , n31908 , n31909 , n31910 , n31911 , n31912 , n31913 , n31914 , n31915 , n31916 , n31917 , n31918 , n31919 , n31920 , n31921 , n31922 , n31923 , n31924 , n31925 , n31926 , n31927 , n31928 , n31929 , n31930 , n31931 , n31932 , n31933 , n31934 , n31935 , n31936 , n31937 , n31938 , n31939 , n31940 , n31941 , n31942 , n31943 , n31944 , n31945 , n31946 , n31947 , n31948 , n31949 , n31950 , n31951 , n31952 , n31953 , n31954 , n31955 , n31956 , n31957 , n31958 , n31959 , n31960 , n31961 , n31962 , n31963 , n31964 , n31965 , n31966 , n31967 , n31968 , n31969 , n31970 , n31971 , n31972 , n31973 , n31974 , n31975 , n31976 , n31977 , n31978 , n31979 , n31980 , n31981 , n31982 , n31983 , n31984 , n31985 , n31986 , n31987 , n31988 , n31989 , n31990 , n31991 , n31992 , n31993 , n31994 , n31995 , n31996 , n31997 , n31998 , n31999 , n32000 , n32001 , n32002 , n32003 , n32004 , n32005 , n32006 , n32007 , n32008 , n32009 , n32010 , n32011 , n32012 , n32013 , n32014 , n32015 , n32016 , n32017 , n32018 , n32019 , n32020 , n32021 , n32022 , n32023 , n32024 , n32025 , n32026 , n32027 , n32028 , n32029 , n32030 , n32031 , n32032 , n32033 , n32034 , n32035 , n32036 , n32037 , n32038 , n32039 , n32040 , n32041 , n32042 , n32043 , n32044 , n32045 , n32046 , n32047 , n32048 , n32049 , n32050 , n32051 , n32052 , n32053 , n32054 , n32055 , n32056 , n32057 , n32058 , n32059 , n32060 , n32061 , n32062 , n32063 , n32064 , n32065 , n32066 , n32067 , n32068 , n32069 , n32070 , n32071 , n32072 , n32073 , n32074 , n32075 , n32076 , n32077 , n32078 , n32079 , n32080 , n32081 , n32082 , n32083 , n32084 , n32085 , n32086 , n32087 , n32088 , n32089 , n32090 , n32091 , n32092 , n32093 , n32094 , n32095 , n32096 , n32097 , n32098 , n32099 , n32100 , n32101 , n32102 , n32103 , n32104 , n32105 , n32106 , n32107 , n32108 , n32109 , n32110 , n32111 , n32112 , n32113 , n32114 , n32115 , n32116 , n32117 , n32118 , n32119 , n32120 , n32121 , n32122 , n32123 , n32124 , n32125 , n32126 , n32127 , n32128 , n32129 , n32130 , n32131 , n32132 , n32133 , n32134 , n32135 , n32136 , n32137 , n32138 , n32139 , n32140 , n32141 , n32142 , n32143 , n32144 , n32145 , n32146 , n32147 , n32148 , n32149 , n32150 , n32151 , n32152 , n32153 , n32154 , n32155 , n32156 , n32157 , n32158 , n32159 , n32160 , n32161 , n32162 , n32163 , n32164 , n32165 , n32166 , n32167 , n32168 , n32169 , n32170 , n32171 , n32172 , n32173 , n32174 , n32175 , n32176 , n32177 , n32178 , n32179 , n32180 , n32181 , n32182 , n32183 , n32184 , n32185 , n32186 , n32187 , n32188 , n32189 , n32190 , n32191 , n32192 , n32193 , n32194 , n32195 , n32196 , n32197 , n32198 , n32199 , n32200 , n32201 , n32202 , n32203 , n32204 , n32205 , n32206 , n32207 , n32208 , n32209 , n32210 , n32211 , n32212 , n32213 , n32214 , n32215 , n32216 , n32217 , n32218 , n32219 , n32220 , n32221 , n32222 , n32223 , n32224 , n32225 , n32226 , n32227 , n32228 , n32229 , n32230 , n32231 , n32232 , n32233 , n32234 , n32235 , n32236 , n32237 , n32238 , n32239 , n32240 , n32241 , n32242 , n32243 , n32244 , n32245 , n32246 , n32247 , n32248 , n32249 , n32250 , n32251 , n32252 , n32253 , n32254 , n32255 , n32256 , n32257 , n32258 , n32259 , n32260 , n32261 , n32262 , n32263 , n32264 , n32265 , n32266 , n32267 , n32268 , n32269 , n32270 , n32271 , n32272 , n32273 , n32274 , n32275 , n32276 , n32277 , n32278 , n32279 , n32280 , n32281 , n32282 , n32283 , n32284 , n32285 , n32286 , n32287 , n32288 , n32289 , n32290 , n32291 , n32292 , n32293 , n32294 , n32295 , n32296 , n32297 , n32298 , n32299 , n32300 , n32301 , n32302 , n32303 , n32304 , n32305 , n32306 , n32307 , n32308 , n32309 , n32310 , n32311 , n32312 , n32313 , n32314 , n32315 , n32316 , n32317 , n32318 , n32319 , n32320 , n32321 , n32322 , n32323 , n32324 , n32325 , n32326 , n32327 , n32328 , n32329 , n32330 , n32331 , n32332 , n32333 , n32334 , n32335 , n32336 , n32337 , n32338 , n32339 , n32340 , n32341 , n32342 , n32343 , n32344 , n32345 , n32346 , n32347 , n32348 , n32349 , n32350 , n32351 , n32352 , n32353 , n32354 , n32355 , n32356 , n32357 , n32358 , n32359 , n32360 , n32361 , n32362 , n32363 , n32364 , n32365 , n32366 , n32367 , n32368 , n32369 , n32370 , n32371 , n32372 , n32373 , n32374 , n32375 , n32376 , n32377 , n32378 , n32379 , n32380 , n32381 , n32382 , n32383 , n32384 , n32385 , n32386 , n32387 , n32388 , n32389 , n32390 , n32391 , n32392 , n32393 , n32394 , n32395 , n32396 , n32397 , n32398 , n32399 , n32400 , n32401 , n32402 , n32403 , n32404 , n32405 , n32406 , n32407 , n32408 , n32409 , n32410 , n32411 , n32412 , n32413 , n32414 , n32415 , n32416 , n32417 , n32418 , n32419 , n32420 , n32421 , n32422 , n32423 , n32424 , n32425 , n32426 , n32427 , n32428 , n32429 , n32430 , n32431 , n32432 , n32433 , n32434 , n32435 , n32436 , n32437 , n32438 , n32439 , n32440 , n32441 , n32442 , n32443 , n32444 , n32445 , n32446 , n32447 , n32448 , n32449 , n32450 , n32451 , n32452 , n32453 , n32454 , n32455 , n32456 , n32457 , n32458 , n32459 , n32460 , n32461 , n32462 , n32463 , n32464 , n32465 , n32466 , n32467 , n32468 , n32469 , n32470 , n32471 , n32472 , n32473 , n32474 , n32475 , n32476 , n32477 , n32478 , n32479 , n32480 , n32481 , n32482 , n32483 , n32484 , n32485 , n32486 , n32487 , n32488 , n32489 , n32490 , n32491 , n32492 , n32493 , n32494 , n32495 , n32496 , n32497 , n32498 , n32499 , n32500 , n32501 , n32502 , n32503 , n32504 , n32505 , n32506 , n32507 , n32508 , n32509 , n32510 , n32511 , n32512 , n32513 , n32514 , n32515 , n32516 , n32517 , n32518 , n32519 , n32520 , n32521 , n32522 , n32523 , n32524 , n32525 , n32526 , n32527 , n32528 , n32529 , n32530 , n32531 , n32532 , n32533 , n32534 , n32535 , n32536 , n32537 , n32538 , n32539 , n32540 , n32541 , n32542 , n32543 , n32544 , n32545 , n32546 , n32547 , n32548 , n32549 , n32550 , n32551 , n32552 , n32553 , n32554 , n32555 , n32556 , n32557 , n32558 , n32559 , n32560 , n32561 , n32562 , n32563 , n32564 , n32565 , n32566 , n32567 , n32568 , n32569 , n32570 , n32571 , n32572 , n32573 , n32574 , n32575 , n32576 , n32577 , n32578 , n32579 , n32580 , n32581 , n32582 , n32583 , n32584 , n32585 , n32586 , n32587 , n32588 , n32589 , n32590 , n32591 , n32592 , n32593 , n32594 , n32595 , n32596 , n32597 , n32598 , n32599 , n32600 , n32601 , n32602 , n32603 , n32604 , n32605 , n32606 , n32607 , n32608 , n32609 , n32610 , n32611 , n32612 , n32613 , n32614 , n32615 , n32616 , n32617 , n32618 , n32619 , n32620 , n32621 , n32622 , n32623 , n32624 , n32625 , n32626 , n32627 , n32628 , n32629 , n32630 , n32631 , n32632 , n32633 , n32634 , n32635 , n32636 , n32637 , n32638 , n32639 , n32640 , n32641 , n32642 , n32643 , n32644 , n32645 , n32646 , n32647 , n32648 , n32649 , n32650 , n32651 , n32652 , n32653 , n32654 , n32655 , n32656 , n32657 , n32658 , n32659 , n32660 , n32661 , n32662 , n32663 , n32664 , n32665 , n32666 , n32667 , n32668 , n32669 , n32670 , n32671 , n32672 , n32673 , n32674 , n32675 , n32676 , n32677 , n32678 , n32679 , n32680 , n32681 , n32682 , n32683 , n32684 , n32685 , n32686 , n32687 , n32688 , n32689 , n32690 , n32691 , n32692 , n32693 , n32694 , n32695 , n32696 , n32697 , n32698 , n32699 , n32700 , n32701 , n32702 , n32703 , n32704 , n32705 , n32706 , n32707 , n32708 , n32709 , n32710 , n32711 , n32712 , n32713 , n32714 , n32715 , n32716 , n32717 , n32718 , n32719 , n32720 , n32721 , n32722 , n32723 , n32724 , n32725 , n32726 , n32727 , n32728 , n32729 , n32730 , n32731 , n32732 , n32733 , n32734 , n32735 , n32736 , n32737 , n32738 , n32739 , n32740 , n32741 , n32742 , n32743 , n32744 , n32745 , n32746 , n32747 , n32748 , n32749 , n32750 , n32751 , n32752 , n32753 , n32754 , n32755 , n32756 , n32757 , n32758 , n32759 , n32760 , n32761 , n32762 , n32763 , n32764 , n32765 , n32766 , n32767 , n32768 , n32769 , n32770 , n32771 , n32772 , n32773 , n32774 , n32775 , n32776 , n32777 , n32778 , n32779 , n32780 , n32781 , n32782 , n32783 , n32784 , n32785 , n32786 , n32787 , n32788 , n32789 , n32790 , n32791 , n32792 , n32793 , n32794 , n32795 , n32796 , n32797 , n32798 , n32799 , n32800 , n32801 , n32802 , n32803 , n32804 , n32805 , n32806 , n32807 , n32808 , n32809 , n32810 , n32811 , n32812 , n32813 , n32814 , n32815 , n32816 , n32817 , n32818 , n32819 , n32820 , n32821 , n32822 , n32823 , n32824 , n32825 , n32826 , n32827 , n32828 , n32829 , n32830 , n32831 , n32832 , n32833 , n32834 , n32835 , n32836 , n32837 , n32838 , n32839 , n32840 , n32841 , n32842 , n32843 , n32844 , n32845 , n32846 , n32847 , n32848 , n32849 , n32850 , n32851 , n32852 , n32853 , n32854 , n32855 , n32856 , n32857 , n32858 , n32859 , n32860 , n32861 , n32862 , n32863 , n32864 , n32865 , n32866 , n32867 , n32868 , n32869 , n32870 , n32871 , n32872 , n32873 , n32874 , n32875 , n32876 , n32877 , n32878 , n32879 , n32880 , n32881 , n32882 , n32883 , n32884 , n32885 , n32886 , n32887 , n32888 , n32889 , n32890 , n32891 , n32892 , n32893 , n32894 , n32895 , n32896 , n32897 , n32898 , n32899 , n32900 , n32901 , n32902 , n32903 , n32904 , n32905 , n32906 , n32907 , n32908 , n32909 , n32910 , n32911 , n32912 , n32913 , n32914 , n32915 , n32916 , n32917 , n32918 , n32919 , n32920 , n32921 , n32922 , n32923 , n32924 , n32925 , n32926 , n32927 , n32928 , n32929 , n32930 , n32931 , n32932 , n32933 , n32934 , n32935 , n32936 , n32937 , n32938 , n32939 , n32940 , n32941 , n32942 , n32943 , n32944 , n32945 , n32946 , n32947 , n32948 , n32949 , n32950 , n32951 , n32952 , n32953 , n32954 , n32955 , n32956 , n32957 , n32958 , n32959 , n32960 , n32961 , n32962 , n32963 , n32964 , n32965 , n32966 , n32967 , n32968 , n32969 , n32970 , n32971 , n32972 , n32973 , n32974 , n32975 , n32976 , n32977 , n32978 , n32979 , n32980 , n32981 , n32982 , n32983 , n32984 , n32985 , n32986 , n32987 , n32988 , n32989 , n32990 , n32991 , n32992 , n32993 , n32994 , n32995 , n32996 , n32997 , n32998 , n32999 , n33000 , n33001 , n33002 , n33003 , n33004 , n33005 , n33006 , n33007 , n33008 , n33009 , n33010 , n33011 , n33012 , n33013 , n33014 , n33015 , n33016 , n33017 , n33018 , n33019 , n33020 , n33021 , n33022 , n33023 , n33024 , n33025 , n33026 , n33027 , n33028 , n33029 , n33030 , n33031 , n33032 , n33033 , n33034 , n33035 , n33036 , n33037 , n33038 , n33039 , n33040 , n33041 , n33042 , n33043 , n33044 , n33045 , n33046 , n33047 , n33048 , n33049 , n33050 , n33051 , n33052 , n33053 , n33054 , n33055 , n33056 , n33057 , n33058 , n33059 , n33060 , n33061 , n33062 , n33063 , n33064 , n33065 , n33066 , n33067 , n33068 , n33069 , n33070 , n33071 , n33072 , n33073 , n33074 , n33075 , n33076 , n33077 , n33078 , n33079 , n33080 , n33081 , n33082 , n33083 , n33084 , n33085 , n33086 , n33087 , n33088 , n33089 , n33090 , n33091 , n33092 , n33093 , n33094 , n33095 , n33096 , n33097 , n33098 , n33099 , n33100 , n33101 , n33102 , n33103 , n33104 , n33105 , n33106 , n33107 , n33108 , n33109 , n33110 , n33111 , n33112 , n33113 , n33114 , n33115 , n33116 , n33117 , n33118 , n33119 , n33120 , n33121 , n33122 , n33123 , n33124 , n33125 , n33126 , n33127 , n33128 , n33129 , n33130 , n33131 , n33132 , n33133 , n33134 , n33135 , n33136 , n33137 , n33138 , n33139 , n33140 , n33141 , n33142 , n33143 , n33144 , n33145 , n33146 , n33147 , n33148 , n33149 , n33150 , n33151 , n33152 , n33153 , n33154 , n33155 , n33156 , n33157 , n33158 , n33159 , n33160 , n33161 , n33162 , n33163 , n33164 , n33165 , n33166 , n33167 , n33168 , n33169 , n33170 , n33171 , n33172 , n33173 , n33174 , n33175 , n33176 , n33177 , n33178 , n33179 , n33180 , n33181 , n33182 , n33183 , n33184 , n33185 , n33186 , n33187 , n33188 , n33189 , n33190 , n33191 , n33192 , n33193 , n33194 , n33195 , n33196 , n33197 , n33198 , n33199 , n33200 , n33201 , n33202 , n33203 , n33204 , n33205 , n33206 , n33207 , n33208 , n33209 , n33210 , n33211 , n33212 , n33213 , n33214 , n33215 , n33216 , n33217 , n33218 , n33219 , n33220 , n33221 , n33222 , n33223 , n33224 , n33225 , n33226 , n33227 , n33228 , n33229 , n33230 , n33231 , n33232 , n33233 , n33234 , n33235 , n33236 , n33237 , n33238 , n33239 , n33240 , n33241 , n33242 , n33243 , n33244 , n33245 , n33246 , n33247 , n33248 , n33249 , n33250 , n33251 , n33252 , n33253 , n33254 , n33255 , n33256 , n33257 , n33258 , n33259 , n33260 , n33261 , n33262 , n33263 , n33264 , n33265 , n33266 , n33267 , n33268 , n33269 , n33270 , n33271 , n33272 , n33273 , n33274 , n33275 , n33276 , n33277 , n33278 , n33279 , n33280 , n33281 , n33282 , n33283 , n33284 , n33285 , n33286 , n33287 , n33288 , n33289 , n33290 , n33291 , n33292 , n33293 , n33294 , n33295 , n33296 , n33297 , n33298 , n33299 , n33300 , n33301 , n33302 , n33303 , n33304 , n33305 , n33306 , n33307 , n33308 , n33309 , n33310 , n33311 , n33312 , n33313 , n33314 , n33315 , n33316 , n33317 , n33318 , n33319 , n33320 , n33321 , n33322 , n33323 , n33324 , n33325 , n33326 , n33327 , n33328 , n33329 , n33330 , n33331 , n33332 , n33333 , n33334 , n33335 , n33336 , n33337 , n33338 , n33339 , n33340 , n33341 , n33342 , n33343 , n33344 , n33345 , n33346 , n33347 , n33348 , n33349 , n33350 , n33351 , n33352 , n33353 , n33354 , n33355 , n33356 , n33357 , n33358 , n33359 , n33360 , n33361 , n33362 , n33363 , n33364 , n33365 , n33366 , n33367 , n33368 , n33369 , n33370 , n33371 , n33372 , n33373 , n33374 , n33375 , n33376 , n33377 , n33378 , n33379 , n33380 , n33381 , n33382 , n33383 , n33384 , n33385 , n33386 , n33387 , n33388 , n33389 , n33390 , n33391 , n33392 , n33393 , n33394 , n33395 , n33396 , n33397 , n33398 , n33399 , n33400 , n33401 , n33402 , n33403 , n33404 , n33405 , n33406 , n33407 , n33408 , n33409 , n33410 , n33411 , n33412 , n33413 , n33414 , n33415 , n33416 , n33417 , n33418 , n33419 , n33420 , n33421 , n33422 , n33423 , n33424 , n33425 , n33426 , n33427 , n33428 , n33429 , n33430 , n33431 , n33432 , n33433 , n33434 , n33435 , n33436 , n33437 , n33438 , n33439 , n33440 , n33441 , n33442 , n33443 , n33444 , n33445 , n33446 , n33447 , n33448 , n33449 , n33450 , n33451 , n33452 , n33453 , n33454 , n33455 , n33456 , n33457 , n33458 , n33459 , n33460 , n33461 , n33462 , n33463 , n33464 , n33465 , n33466 , n33467 , n33468 , n33469 , n33470 , n33471 , n33472 , n33473 , n33474 , n33475 , n33476 , n33477 , n33478 , n33479 , n33480 , n33481 , n33482 , n33483 , n33484 , n33485 , n33486 , n33487 , n33488 , n33489 , n33490 , n33491 , n33492 , n33493 , n33494 , n33495 , n33496 , n33497 , n33498 , n33499 , n33500 , n33501 , n33502 , n33503 , n33504 , n33505 , n33506 , n33507 , n33508 , n33509 , n33510 , n33511 , n33512 , n33513 , n33514 , n33515 , n33516 , n33517 , n33518 , n33519 , n33520 , n33521 , n33522 , n33523 , n33524 , n33525 , n33526 , n33527 , n33528 , n33529 , n33530 , n33531 , n33532 , n33533 , n33534 , n33535 , n33536 , n33537 , n33538 , n33539 , n33540 , n33541 , n33542 , n33543 , n33544 , n33545 , n33546 , n33547 , n33548 , n33549 , n33550 , n33551 , n33552 , n33553 , n33554 , n33555 , n33556 , n33557 , n33558 , n33559 , n33560 , n33561 , n33562 , n33563 , n33564 , n33565 , n33566 , n33567 , n33568 , n33569 , n33570 , n33571 , n33572 , n33573 , n33574 , n33575 , n33576 , n33577 , n33578 , n33579 , n33580 , n33581 , n33582 , n33583 , n33584 , n33585 , n33586 , n33587 , n33588 , n33589 , n33590 , n33591 , n33592 , n33593 , n33594 , n33595 , n33596 , n33597 , n33598 , n33599 , n33600 , n33601 , n33602 , n33603 , n33604 , n33605 , n33606 , n33607 , n33608 , n33609 , n33610 , n33611 , n33612 , n33613 , n33614 , n33615 , n33616 , n33617 , n33618 , n33619 , n33620 , n33621 , n33622 , n33623 , n33624 , n33625 , n33626 , n33627 , n33628 , n33629 , n33630 , n33631 , n33632 , n33633 , n33634 , n33635 , n33636 , n33637 , n33638 , n33639 , n33640 , n33641 , n33642 , n33643 , n33644 , n33645 , n33646 , n33647 , n33648 , n33649 , n33650 , n33651 , n33652 , n33653 , n33654 , n33655 , n33656 , n33657 , n33658 , n33659 , n33660 , n33661 , n33662 , n33663 , n33664 , n33665 , n33666 , n33667 , n33668 , n33669 , n33670 , n33671 , n33672 , n33673 , n33674 , n33675 , n33676 , n33677 , n33678 , n33679 , n33680 , n33681 , n33682 , n33683 , n33684 , n33685 , n33686 , n33687 , n33688 , n33689 , n33690 , n33691 , n33692 , n33693 , n33694 , n33695 , n33696 , n33697 , n33698 , n33699 , n33700 , n33701 , n33702 , n33703 , n33704 , n33705 , n33706 , n33707 , n33708 , n33709 , n33710 , n33711 , n33712 , n33713 , n33714 , n33715 , n33716 , n33717 , n33718 , n33719 , n33720 , n33721 , n33722 , n33723 , n33724 , n33725 , n33726 , n33727 , n33728 , n33729 , n33730 , n33731 , n33732 , n33733 , n33734 , n33735 , n33736 , n33737 , n33738 , n33739 , n33740 , n33741 , n33742 , n33743 , n33744 , n33745 , n33746 , n33747 , n33748 , n33749 , n33750 , n33751 , n33752 , n33753 , n33754 , n33755 , n33756 , n33757 , n33758 , n33759 , n33760 , n33761 , n33762 , n33763 , n33764 , n33765 , n33766 , n33767 , n33768 , n33769 , n33770 , n33771 , n33772 , n33773 , n33774 , n33775 , n33776 , n33777 , n33778 , n33779 , n33780 , n33781 , n33782 , n33783 , n33784 , n33785 , n33786 , n33787 , n33788 , n33789 , n33790 , n33791 , n33792 , n33793 , n33794 , n33795 , n33796 , n33797 , n33798 , n33799 , n33800 , n33801 , n33802 , n33803 , n33804 , n33805 , n33806 , n33807 , n33808 , n33809 , n33810 , n33811 , n33812 , n33813 , n33814 , n33815 , n33816 , n33817 , n33818 , n33819 , n33820 , n33821 , n33822 , n33823 , n33824 , n33825 , n33826 , n33827 , n33828 , n33829 , n33830 , n33831 , n33832 , n33833 , n33834 , n33835 , n33836 , n33837 , n33838 , n33839 , n33840 , n33841 , n33842 , n33843 , n33844 , n33845 , n33846 , n33847 , n33848 , n33849 , n33850 , n33851 , n33852 , n33853 , n33854 , n33855 , n33856 , n33857 , n33858 , n33859 , n33860 , n33861 , n33862 , n33863 , n33864 , n33865 , n33866 , n33867 , n33868 , n33869 , n33870 , n33871 , n33872 , n33873 , n33874 , n33875 , n33876 , n33877 , n33878 , n33879 , n33880 , n33881 , n33882 , n33883 , n33884 , n33885 , n33886 , n33887 , n33888 , n33889 , n33890 , n33891 , n33892 , n33893 , n33894 , n33895 , n33896 , n33897 , n33898 , n33899 , n33900 , n33901 , n33902 , n33903 , n33904 , n33905 , n33906 , n33907 , n33908 , n33909 , n33910 , n33911 , n33912 , n33913 , n33914 , n33915 , n33916 , n33917 , n33918 , n33919 , n33920 , n33921 , n33922 , n33923 , n33924 , n33925 , n33926 , n33927 , n33928 , n33929 , n33930 , n33931 , n33932 , n33933 , n33934 , n33935 , n33936 , n33937 , n33938 , n33939 , n33940 , n33941 , n33942 , n33943 , n33944 , n33945 , n33946 , n33947 , n33948 , n33949 , n33950 , n33951 , n33952 , n33953 , n33954 , n33955 , n33956 , n33957 , n33958 , n33959 , n33960 , n33961 , n33962 , n33963 , n33964 , n33965 , n33966 , n33967 , n33968 , n33969 , n33970 , n33971 , n33972 , n33973 , n33974 , n33975 , n33976 , n33977 , n33978 , n33979 , n33980 , n33981 , n33982 , n33983 , n33984 , n33985 , n33986 , n33987 , n33988 , n33989 , n33990 , n33991 , n33992 , n33993 , n33994 , n33995 , n33996 , n33997 , n33998 , n33999 , n34000 , n34001 , n34002 , n34003 , n34004 , n34005 , n34006 , n34007 , n34008 , n34009 , n34010 , n34011 , n34012 , n34013 , n34014 , n34015 , n34016 , n34017 , n34018 , n34019 , n34020 , n34021 , n34022 , n34023 , n34024 , n34025 , n34026 , n34027 , n34028 , n34029 , n34030 , n34031 , n34032 , n34033 , n34034 , n34035 , n34036 , n34037 , n34038 , n34039 , n34040 , n34041 , n34042 , n34043 , n34044 , n34045 , n34046 , n34047 , n34048 , n34049 , n34050 , n34051 , n34052 , n34053 , n34054 , n34055 , n34056 , n34057 , n34058 , n34059 , n34060 , n34061 , n34062 , n34063 , n34064 , n34065 , n34066 , n34067 , n34068 , n34069 , n34070 , n34071 , n34072 , n34073 , n34074 , n34075 , n34076 , n34077 , n34078 , n34079 , n34080 , n34081 , n34082 , n34083 , n34084 , n34085 , n34086 , n34087 , n34088 , n34089 , n34090 , n34091 , n34092 , n34093 , n34094 , n34095 , n34096 , n34097 , n34098 , n34099 , n34100 , n34101 , n34102 , n34103 , n34104 , n34105 , n34106 , n34107 , n34108 , n34109 , n34110 , n34111 , n34112 , n34113 , n34114 , n34115 , n34116 , n34117 , n34118 , n34119 , n34120 , n34121 , n34122 , n34123 , n34124 , n34125 , n34126 , n34127 , n34128 , n34129 , n34130 , n34131 , n34132 , n34133 , n34134 , n34135 , n34136 , n34137 , n34138 , n34139 , n34140 , n34141 , n34142 , n34143 , n34144 , n34145 , n34146 , n34147 , n34148 , n34149 , n34150 , n34151 , n34152 , n34153 , n34154 , n34155 , n34156 , n34157 , n34158 , n34159 , n34160 , n34161 , n34162 , n34163 , n34164 , n34165 , n34166 , n34167 , n34168 , n34169 , n34170 , n34171 , n34172 , n34173 , n34174 , n34175 , n34176 , n34177 , n34178 , n34179 , n34180 , n34181 , n34182 , n34183 , n34184 , n34185 , n34186 , n34187 , n34188 , n34189 , n34190 , n34191 , n34192 , n34193 , n34194 , n34195 , n34196 , n34197 , n34198 , n34199 , n34200 , n34201 , n34202 , n34203 , n34204 , n34205 , n34206 , n34207 , n34208 , n34209 , n34210 , n34211 , n34212 , n34213 , n34214 , n34215 , n34216 , n34217 , n34218 , n34219 , n34220 , n34221 , n34222 , n34223 , n34224 , n34225 , n34226 , n34227 , n34228 , n34229 , n34230 , n34231 , n34232 , n34233 , n34234 , n34235 , n34236 , n34237 , n34238 , n34239 , n34240 , n34241 , n34242 , n34243 , n34244 , n34245 , n34246 , n34247 , n34248 , n34249 , n34250 , n34251 , n34252 , n34253 , n34254 , n34255 , n34256 , n34257 , n34258 , n34259 , n34260 , n34261 , n34262 , n34263 , n34264 , n34265 , n34266 , n34267 , n34268 , n34269 , n34270 , n34271 , n34272 , n34273 , n34274 , n34275 , n34276 , n34277 , n34278 , n34279 , n34280 , n34281 , n34282 , n34283 , n34284 , n34285 , n34286 , n34287 , n34288 , n34289 , n34290 , n34291 , n34292 , n34293 , n34294 , n34295 , n34296 , n34297 , n34298 , n34299 , n34300 , n34301 , n34302 , n34303 , n34304 , n34305 , n34306 , n34307 , n34308 , n34309 , n34310 , n34311 , n34312 , n34313 , n34314 , n34315 , n34316 , n34317 , n34318 , n34319 , n34320 , n34321 , n34322 , n34323 , n34324 , n34325 , n34326 , n34327 , n34328 , n34329 , n34330 , n34331 , n34332 , n34333 , n34334 , n34335 , n34336 , n34337 , n34338 , n34339 , n34340 , n34341 , n34342 , n34343 , n34344 , n34345 , n34346 , n34347 , n34348 , n34349 , n34350 , n34351 , n34352 , n34353 , n34354 , n34355 , n34356 , n34357 , n34358 , n34359 , n34360 , n34361 , n34362 , n34363 , n34364 , n34365 , n34366 , n34367 , n34368 , n34369 , n34370 , n34371 , n34372 , n34373 , n34374 , n34375 , n34376 , n34377 , n34378 , n34379 , n34380 , n34381 , n34382 , n34383 , n34384 , n34385 , n34386 , n34387 , n34388 , n34389 , n34390 , n34391 , n34392 , n34393 , n34394 , n34395 , n34396 , n34397 , n34398 , n34399 , n34400 , n34401 , n34402 , n34403 , n34404 , n34405 , n34406 , n34407 , n34408 , n34409 , n34410 , n34411 , n34412 , n34413 , n34414 , n34415 , n34416 , n34417 , n34418 , n34419 , n34420 , n34421 , n34422 , n34423 , n34424 , n34425 , n34426 , n34427 , n34428 , n34429 , n34430 , n34431 , n34432 , n34433 , n34434 , n34435 , n34436 , n34437 , n34438 , n34439 , n34440 , n34441 , n34442 , n34443 , n34444 , n34445 , n34446 , n34447 , n34448 , n34449 , n34450 , n34451 , n34452 , n34453 , n34454 , n34455 , n34456 , n34457 , n34458 , n34459 , n34460 , n34461 , n34462 , n34463 , n34464 , n34465 , n34466 , n34467 , n34468 , n34469 , n34470 , n34471 , n34472 , n34473 , n34474 , n34475 , n34476 , n34477 , n34478 , n34479 , n34480 , n34481 , n34482 , n34483 , n34484 , n34485 , n34486 , n34487 , n34488 , n34489 , n34490 , n34491 , n34492 , n34493 , n34494 , n34495 , n34496 , n34497 , n34498 , n34499 , n34500 , n34501 , n34502 , n34503 , n34504 , n34505 , n34506 , n34507 , n34508 , n34509 , n34510 , n34511 , n34512 , n34513 , n34514 , n34515 , n34516 , n34517 , n34518 , n34519 , n34520 , n34521 , n34522 , n34523 , n34524 , n34525 , n34526 , n34527 , n34528 , n34529 , n34530 , n34531 , n34532 , n34533 , n34534 , n34535 , n34536 , n34537 , n34538 , n34539 , n34540 , n34541 , n34542 , n34543 , n34544 , n34545 , n34546 , n34547 , n34548 , n34549 , n34550 , n34551 , n34552 , n34553 , n34554 , n34555 , n34556 , n34557 , n34558 , n34559 , n34560 , n34561 , n34562 , n34563 , n34564 , n34565 , n34566 , n34567 , n34568 , n34569 , n34570 , n34571 , n34572 , n34573 , n34574 , n34575 , n34576 , n34577 , n34578 , n34579 , n34580 , n34581 , n34582 , n34583 , n34584 , n34585 , n34586 , n34587 , n34588 , n34589 , n34590 , n34591 , n34592 , n34593 , n34594 , n34595 , n34596 , n34597 , n34598 , n34599 , n34600 , n34601 , n34602 , n34603 , n34604 , n34605 , n34606 , n34607 , n34608 , n34609 , n34610 , n34611 , n34612 , n34613 , n34614 , n34615 , n34616 , n34617 , n34618 , n34619 , n34620 , n34621 , n34622 , n34623 , n34624 , n34625 , n34626 , n34627 , n34628 , n34629 , n34630 , n34631 , n34632 , n34633 , n34634 , n34635 , n34636 , n34637 , n34638 , n34639 , n34640 , n34641 , n34642 , n34643 , n34644 , n34645 , n34646 , n34647 , n34648 , n34649 , n34650 , n34651 , n34652 , n34653 , n34654 , n34655 , n34656 , n34657 , n34658 , n34659 , n34660 , n34661 , n34662 , n34663 , n34664 , n34665 , n34666 , n34667 , n34668 , n34669 , n34670 , n34671 , n34672 , n34673 , n34674 , n34675 , n34676 , n34677 , n34678 , n34679 , n34680 , n34681 , n34682 , n34683 , n34684 , n34685 , n34686 , n34687 , n34688 , n34689 , n34690 , n34691 , n34692 , n34693 , n34694 , n34695 , n34696 , n34697 , n34698 , n34699 , n34700 , n34701 , n34702 , n34703 , n34704 , n34705 , n34706 , n34707 , n34708 , n34709 , n34710 , n34711 , n34712 , n34713 , n34714 , n34715 , n34716 , n34717 , n34718 , n34719 , n34720 , n34721 , n34722 , n34723 , n34724 , n34725 , n34726 , n34727 , n34728 , n34729 , n34730 , n34731 , n34732 , n34733 , n34734 , n34735 , n34736 , n34737 , n34738 , n34739 , n34740 , n34741 , n34742 , n34743 , n34744 , n34745 , n34746 , n34747 , n34748 , n34749 , n34750 , n34751 , n34752 , n34753 , n34754 , n34755 , n34756 , n34757 , n34758 , n34759 , n34760 , n34761 , n34762 , n34763 , n34764 , n34765 , n34766 , n34767 , n34768 , n34769 , n34770 , n34771 , n34772 , n34773 , n34774 , n34775 , n34776 , n34777 , n34778 , n34779 , n34780 , n34781 , n34782 , n34783 , n34784 , n34785 , n34786 , n34787 , n34788 , n34789 , n34790 , n34791 , n34792 , n34793 , n34794 , n34795 , n34796 , n34797 , n34798 , n34799 , n34800 , n34801 , n34802 , n34803 , n34804 , n34805 , n34806 , n34807 , n34808 , n34809 , n34810 , n34811 , n34812 , n34813 , n34814 , n34815 , n34816 , n34817 , n34818 , n34819 , n34820 , n34821 , n34822 , n34823 , n34824 , n34825 , n34826 , n34827 , n34828 , n34829 , n34830 , n34831 , n34832 , n34833 , n34834 , n34835 , n34836 , n34837 , n34838 , n34839 , n34840 , n34841 , n34842 , n34843 , n34844 , n34845 , n34846 , n34847 , n34848 , n34849 , n34850 , n34851 , n34852 , n34853 , n34854 , n34855 , n34856 , n34857 , n34858 , n34859 , n34860 , n34861 , n34862 , n34863 , n34864 , n34865 , n34866 , n34867 , n34868 , n34869 , n34870 , n34871 , n34872 , n34873 , n34874 , n34875 , n34876 , n34877 , n34878 , n34879 , n34880 , n34881 , n34882 , n34883 , n34884 , n34885 , n34886 , n34887 , n34888 , n34889 , n34890 , n34891 , n34892 , n34893 , n34894 , n34895 , n34896 , n34897 , n34898 , n34899 , n34900 , n34901 , n34902 , n34903 , n34904 , n34905 , n34906 , n34907 , n34908 , n34909 , n34910 , n34911 , n34912 , n34913 , n34914 , n34915 , n34916 , n34917 , n34918 , n34919 , n34920 , n34921 , n34922 , n34923 , n34924 , n34925 , n34926 , n34927 , n34928 , n34929 , n34930 , n34931 , n34932 , n34933 , n34934 , n34935 , n34936 , n34937 , n34938 , n34939 , n34940 , n34941 , n34942 , n34943 , n34944 , n34945 , n34946 , n34947 , n34948 , n34949 , n34950 , n34951 , n34952 , n34953 , n34954 , n34955 , n34956 , n34957 , n34958 , n34959 , n34960 , n34961 , n34962 , n34963 , n34964 , n34965 , n34966 , n34967 , n34968 , n34969 , n34970 , n34971 , n34972 , n34973 , n34974 , n34975 , n34976 , n34977 , n34978 , n34979 , n34980 , n34981 , n34982 , n34983 , n34984 , n34985 , n34986 , n34987 , n34988 , n34989 , n34990 , n34991 , n34992 , n34993 , n34994 , n34995 , n34996 , n34997 , n34998 , n34999 , n35000 , n35001 , n35002 , n35003 , n35004 , n35005 , n35006 , n35007 , n35008 , n35009 , n35010 , n35011 , n35012 , n35013 , n35014 , n35015 , n35016 , n35017 , n35018 , n35019 , n35020 , n35021 , n35022 , n35023 , n35024 , n35025 , n35026 , n35027 , n35028 , n35029 , n35030 , n35031 , n35032 , n35033 , n35034 , n35035 , n35036 , n35037 , n35038 , n35039 , n35040 , n35041 , n35042 , n35043 , n35044 , n35045 , n35046 , n35047 , n35048 , n35049 , n35050 , n35051 , n35052 , n35053 , n35054 , n35055 , n35056 , n35057 , n35058 , n35059 , n35060 , n35061 , n35062 , n35063 , n35064 , n35065 , n35066 , n35067 , n35068 , n35069 , n35070 , n35071 , n35072 , n35073 , n35074 , n35075 , n35076 , n35077 , n35078 , n35079 , n35080 , n35081 , n35082 , n35083 , n35084 , n35085 , n35086 , n35087 , n35088 , n35089 , n35090 , n35091 , n35092 , n35093 , n35094 , n35095 , n35096 , n35097 , n35098 , n35099 , n35100 , n35101 , n35102 , n35103 , n35104 , n35105 , n35106 , n35107 , n35108 , n35109 , n35110 , n35111 , n35112 , n35113 , n35114 , n35115 , n35116 , n35117 , n35118 , n35119 , n35120 , n35121 , n35122 , n35123 , n35124 , n35125 , n35126 , n35127 , n35128 , n35129 , n35130 , n35131 , n35132 , n35133 , n35134 , n35135 , n35136 , n35137 , n35138 , n35139 , n35140 , n35141 , n35142 , n35143 , n35144 , n35145 , n35146 , n35147 , n35148 , n35149 , n35150 , n35151 , n35152 , n35153 , n35154 , n35155 , n35156 , n35157 , n35158 , n35159 , n35160 , n35161 , n35162 , n35163 , n35164 , n35165 , n35166 , n35167 , n35168 , n35169 , n35170 , n35171 , n35172 , n35173 , n35174 , n35175 , n35176 , n35177 , n35178 , n35179 , n35180 , n35181 , n35182 , n35183 , n35184 , n35185 , n35186 , n35187 , n35188 , n35189 , n35190 , n35191 , n35192 , n35193 , n35194 , n35195 , n35196 , n35197 , n35198 , n35199 , n35200 , n35201 , n35202 , n35203 , n35204 , n35205 , n35206 , n35207 , n35208 , n35209 , n35210 , n35211 , n35212 , n35213 , n35214 , n35215 , n35216 , n35217 , n35218 , n35219 , n35220 , n35221 , n35222 , n35223 , n35224 , n35225 , n35226 , n35227 , n35228 , n35229 , n35230 , n35231 , n35232 , n35233 , n35234 , n35235 , n35236 , n35237 , n35238 , n35239 , n35240 , n35241 , n35242 , n35243 , n35244 , n35245 , n35246 , n35247 , n35248 , n35249 , n35250 , n35251 , n35252 , n35253 , n35254 , n35255 , n35256 , n35257 , n35258 , n35259 , n35260 , n35261 , n35262 , n35263 , n35264 , n35265 , n35266 , n35267 , n35268 , n35269 , n35270 , n35271 , n35272 , n35273 , n35274 , n35275 , n35276 , n35277 , n35278 , n35279 , n35280 , n35281 , n35282 , n35283 , n35284 , n35285 , n35286 , n35287 , n35288 , n35289 , n35290 , n35291 , n35292 , n35293 , n35294 , n35295 , n35296 , n35297 , n35298 , n35299 , n35300 , n35301 , n35302 , n35303 , n35304 , n35305 , n35306 , n35307 , n35308 , n35309 , n35310 , n35311 , n35312 , n35313 , n35314 , n35315 , n35316 , n35317 , n35318 , n35319 , n35320 , n35321 , n35322 , n35323 , n35324 , n35325 , n35326 , n35327 , n35328 , n35329 , n35330 , n35331 , n35332 , n35333 , n35334 , n35335 , n35336 , n35337 , n35338 , n35339 , n35340 , n35341 , n35342 , n35343 , n35344 , n35345 , n35346 , n35347 , n35348 , n35349 , n35350 , n35351 , n35352 , n35353 , n35354 , n35355 , n35356 , n35357 , n35358 , n35359 , n35360 , n35361 , n35362 , n35363 , n35364 , n35365 , n35366 , n35367 , n35368 , n35369 , n35370 , n35371 , n35372 , n35373 , n35374 , n35375 , n35376 , n35377 , n35378 , n35379 , n35380 , n35381 , n35382 , n35383 , n35384 , n35385 , n35386 , n35387 , n35388 , n35389 , n35390 , n35391 , n35392 , n35393 , n35394 , n35395 , n35396 , n35397 , n35398 , n35399 , n35400 , n35401 , n35402 , n35403 , n35404 , n35405 , n35406 , n35407 , n35408 , n35409 , n35410 , n35411 , n35412 , n35413 , n35414 , n35415 , n35416 , n35417 , n35418 , n35419 , n35420 , n35421 , n35422 , n35423 , n35424 , n35425 , n35426 , n35427 , n35428 , n35429 , n35430 , n35431 , n35432 , n35433 , n35434 , n35435 , n35436 , n35437 , n35438 , n35439 , n35440 , n35441 , n35442 , n35443 , n35444 , n35445 , n35446 , n35447 , n35448 , n35449 , n35450 , n35451 , n35452 , n35453 , n35454 , n35455 , n35456 , n35457 , n35458 , n35459 , n35460 , n35461 , n35462 , n35463 , n35464 , n35465 , n35466 , n35467 , n35468 , n35469 , n35470 , n35471 , n35472 , n35473 , n35474 , n35475 , n35476 , n35477 , n35478 , n35479 , n35480 , n35481 , n35482 , n35483 , n35484 , n35485 , n35486 , n35487 , n35488 , n35489 , n35490 , n35491 , n35492 , n35493 , n35494 , n35495 , n35496 , n35497 , n35498 , n35499 , n35500 , n35501 , n35502 , n35503 , n35504 , n35505 , n35506 , n35507 , n35508 , n35509 , n35510 , n35511 , n35512 , n35513 , n35514 , n35515 , n35516 , n35517 , n35518 , n35519 , n35520 , n35521 , n35522 , n35523 , n35524 , n35525 , n35526 , n35527 , n35528 , n35529 , n35530 , n35531 , n35532 , n35533 , n35534 , n35535 , n35536 , n35537 , n35538 , n35539 , n35540 , n35541 , n35542 , n35543 , n35544 , n35545 , n35546 , n35547 , n35548 , n35549 , n35550 , n35551 , n35552 , n35553 , n35554 , n35555 , n35556 , n35557 , n35558 , n35559 , n35560 , n35561 , n35562 , n35563 , n35564 , n35565 , n35566 , n35567 , n35568 , n35569 , n35570 , n35571 , n35572 , n35573 , n35574 , n35575 , n35576 , n35577 , n35578 , n35579 , n35580 , n35581 , n35582 , n35583 , n35584 , n35585 , n35586 , n35587 , n35588 , n35589 , n35590 , n35591 , n35592 , n35593 , n35594 , n35595 , n35596 , n35597 , n35598 , n35599 , n35600 , n35601 , n35602 , n35603 , n35604 , n35605 , n35606 , n35607 , n35608 , n35609 , n35610 , n35611 , n35612 , n35613 , n35614 , n35615 , n35616 , n35617 , n35618 , n35619 , n35620 , n35621 , n35622 , n35623 , n35624 , n35625 , n35626 , n35627 , n35628 , n35629 , n35630 , n35631 , n35632 , n35633 , n35634 , n35635 , n35636 , n35637 , n35638 , n35639 , n35640 , n35641 , n35642 , n35643 , n35644 , n35645 , n35646 , n35647 , n35648 , n35649 , n35650 , n35651 , n35652 , n35653 , n35654 , n35655 , n35656 , n35657 , n35658 , n35659 , n35660 , n35661 , n35662 , n35663 , n35664 , n35665 , n35666 , n35667 , n35668 , n35669 , n35670 , n35671 , n35672 , n35673 , n35674 , n35675 , n35676 , n35677 , n35678 , n35679 , n35680 , n35681 , n35682 , n35683 , n35684 , n35685 , n35686 , n35687 , n35688 , n35689 , n35690 , n35691 , n35692 , n35693 , n35694 , n35695 , n35696 , n35697 , n35698 , n35699 , n35700 , n35701 , n35702 , n35703 , n35704 , n35705 , n35706 , n35707 , n35708 , n35709 , n35710 , n35711 , n35712 , n35713 , n35714 , n35715 , n35716 , n35717 , n35718 , n35719 , n35720 , n35721 , n35722 , n35723 , n35724 , n35725 , n35726 , n35727 , n35728 , n35729 , n35730 , n35731 , n35732 , n35733 , n35734 , n35735 , n35736 , n35737 , n35738 , n35739 , n35740 , n35741 , n35742 , n35743 , n35744 , n35745 , n35746 , n35747 , n35748 , n35749 , n35750 , n35751 , n35752 , n35753 , n35754 , n35755 , n35756 , n35757 , n35758 , n35759 , n35760 , n35761 , n35762 , n35763 , n35764 , n35765 , n35766 , n35767 , n35768 , n35769 , n35770 , n35771 , n35772 , n35773 , n35774 , n35775 , n35776 , n35777 , n35778 , n35779 , n35780 , n35781 , n35782 , n35783 , n35784 , n35785 , n35786 , n35787 , n35788 , n35789 , n35790 , n35791 , n35792 , n35793 , n35794 , n35795 , n35796 , n35797 , n35798 , n35799 , n35800 , n35801 , n35802 , n35803 , n35804 , n35805 , n35806 , n35807 , n35808 , n35809 , n35810 , n35811 , n35812 , n35813 , n35814 , n35815 , n35816 , n35817 , n35818 , n35819 , n35820 , n35821 , n35822 , n35823 , n35824 , n35825 , n35826 , n35827 , n35828 , n35829 , n35830 , n35831 , n35832 , n35833 , n35834 , n35835 , n35836 , n35837 , n35838 , n35839 , n35840 , n35841 , n35842 , n35843 , n35844 , n35845 , n35846 , n35847 , n35848 , n35849 , n35850 , n35851 , n35852 , n35853 , n35854 , n35855 , n35856 , n35857 , n35858 , n35859 , n35860 , n35861 , n35862 , n35863 , n35864 , n35865 , n35866 , n35867 , n35868 , n35869 , n35870 , n35871 , n35872 , n35873 , n35874 , n35875 , n35876 , n35877 , n35878 , n35879 , n35880 , n35881 , n35882 , n35883 , n35884 , n35885 , n35886 , n35887 , n35888 , n35889 , n35890 , n35891 , n35892 , n35893 , n35894 , n35895 , n35896 , n35897 , n35898 , n35899 , n35900 , n35901 , n35902 , n35903 , n35904 , n35905 , n35906 , n35907 , n35908 , n35909 , n35910 , n35911 , n35912 , n35913 , n35914 , n35915 , n35916 , n35917 , n35918 , n35919 , n35920 , n35921 , n35922 , n35923 , n35924 , n35925 , n35926 , n35927 , n35928 , n35929 , n35930 , n35931 , n35932 , n35933 , n35934 , n35935 , n35936 , n35937 , n35938 , n35939 , n35940 , n35941 , n35942 , n35943 , n35944 , n35945 , n35946 , n35947 , n35948 , n35949 , n35950 , n35951 , n35952 , n35953 , n35954 , n35955 , n35956 , n35957 , n35958 , n35959 , n35960 , n35961 , n35962 , n35963 , n35964 , n35965 , n35966 , n35967 , n35968 , n35969 , n35970 , n35971 , n35972 , n35973 , n35974 , n35975 , n35976 , n35977 , n35978 , n35979 , n35980 , n35981 , n35982 , n35983 , n35984 , n35985 , n35986 , n35987 , n35988 , n35989 , n35990 , n35991 , n35992 , n35993 , n35994 , n35995 , n35996 , n35997 , n35998 , n35999 , n36000 , n36001 , n36002 , n36003 , n36004 , n36005 , n36006 , n36007 , n36008 , n36009 , n36010 , n36011 , n36012 , n36013 , n36014 , n36015 , n36016 , n36017 , n36018 , n36019 , n36020 , n36021 , n36022 , n36023 , n36024 , n36025 , n36026 , n36027 , n36028 , n36029 , n36030 , n36031 , n36032 , n36033 , n36034 , n36035 , n36036 , n36037 , n36038 , n36039 , n36040 , n36041 , n36042 , n36043 , n36044 , n36045 , n36046 , n36047 , n36048 , n36049 , n36050 , n36051 , n36052 , n36053 , n36054 , n36055 , n36056 , n36057 , n36058 , n36059 , n36060 , n36061 , n36062 , n36063 , n36064 , n36065 , n36066 , n36067 , n36068 , n36069 , n36070 , n36071 , n36072 , n36073 , n36074 , n36075 , n36076 , n36077 , n36078 , n36079 , n36080 , n36081 , n36082 , n36083 , n36084 , n36085 , n36086 , n36087 , n36088 , n36089 , n36090 , n36091 , n36092 , n36093 , n36094 , n36095 , n36096 , n36097 , n36098 , n36099 , n36100 , n36101 , n36102 , n36103 , n36104 , n36105 , n36106 , n36107 , n36108 , n36109 , n36110 , n36111 , n36112 , n36113 , n36114 , n36115 , n36116 , n36117 , n36118 , n36119 , n36120 , n36121 , n36122 , n36123 , n36124 , n36125 , n36126 , n36127 , n36128 , n36129 , n36130 , n36131 , n36132 , n36133 , n36134 , n36135 , n36136 , n36137 , n36138 , n36139 , n36140 , n36141 , n36142 , n36143 , n36144 , n36145 , n36146 , n36147 , n36148 , n36149 , n36150 , n36151 , n36152 , n36153 , n36154 , n36155 , n36156 , n36157 , n36158 , n36159 , n36160 , n36161 , n36162 , n36163 , n36164 , n36165 , n36166 , n36167 , n36168 , n36169 , n36170 , n36171 , n36172 , n36173 , n36174 , n36175 , n36176 , n36177 , n36178 , n36179 , n36180 , n36181 , n36182 , n36183 , n36184 , n36185 , n36186 , n36187 , n36188 , n36189 , n36190 , n36191 , n36192 , n36193 , n36194 , n36195 , n36196 , n36197 , n36198 , n36199 , n36200 , n36201 , n36202 , n36203 , n36204 , n36205 , n36206 , n36207 , n36208 , n36209 , n36210 , n36211 , n36212 , n36213 , n36214 , n36215 , n36216 , n36217 , n36218 , n36219 , n36220 , n36221 , n36222 , n36223 , n36224 , n36225 , n36226 , n36227 , n36228 , n36229 , n36230 , n36231 , n36232 , n36233 , n36234 , n36235 , n36236 , n36237 , n36238 , n36239 , n36240 , n36241 , n36242 , n36243 , n36244 , n36245 , n36246 , n36247 , n36248 , n36249 , n36250 , n36251 , n36252 , n36253 , n36254 , n36255 , n36256 , n36257 , n36258 , n36259 , n36260 , n36261 , n36262 , n36263 , n36264 , n36265 , n36266 , n36267 , n36268 , n36269 , n36270 , n36271 , n36272 , n36273 , n36274 , n36275 , n36276 , n36277 , n36278 , n36279 , n36280 , n36281 , n36282 , n36283 , n36284 , n36285 , n36286 , n36287 , n36288 , n36289 , n36290 , n36291 , n36292 , n36293 , n36294 , n36295 , n36296 , n36297 , n36298 , n36299 , n36300 , n36301 , n36302 , n36303 , n36304 , n36305 , n36306 , n36307 , n36308 , n36309 , n36310 , n36311 , n36312 , n36313 , n36314 , n36315 , n36316 , n36317 , n36318 , n36319 , n36320 , n36321 , n36322 , n36323 , n36324 , n36325 , n36326 , n36327 , n36328 , n36329 , n36330 , n36331 , n36332 , n36333 , n36334 , n36335 , n36336 , n36337 , n36338 , n36339 , n36340 , n36341 , n36342 , n36343 , n36344 , n36345 , n36346 , n36347 , n36348 , n36349 , n36350 , n36351 , n36352 , n36353 , n36354 , n36355 , n36356 , n36357 , n36358 , n36359 , n36360 , n36361 , n36362 , n36363 , n36364 , n36365 , n36366 , n36367 , n36368 , n36369 , n36370 , n36371 , n36372 , n36373 , n36374 , n36375 , n36376 , n36377 , n36378 , n36379 , n36380 , n36381 , n36382 , n36383 , n36384 , n36385 , n36386 , n36387 , n36388 , n36389 , n36390 , n36391 , n36392 , n36393 , n36394 , n36395 , n36396 , n36397 , n36398 , n36399 , n36400 , n36401 , n36402 , n36403 , n36404 , n36405 , n36406 , n36407 , n36408 , n36409 , n36410 , n36411 , n36412 , n36413 , n36414 , n36415 , n36416 , n36417 , n36418 , n36419 , n36420 , n36421 , n36422 , n36423 , n36424 , n36425 , n36426 , n36427 , n36428 , n36429 , n36430 , n36431 , n36432 , n36433 , n36434 , n36435 , n36436 , n36437 , n36438 , n36439 , n36440 , n36441 , n36442 , n36443 , n36444 , n36445 , n36446 , n36447 , n36448 , n36449 , n36450 , n36451 , n36452 , n36453 , n36454 , n36455 , n36456 , n36457 , n36458 , n36459 , n36460 , n36461 , n36462 , n36463 , n36464 , n36465 , n36466 , n36467 , n36468 , n36469 , n36470 , n36471 , n36472 , n36473 , n36474 , n36475 , n36476 , n36477 , n36478 , n36479 , n36480 , n36481 , n36482 , n36483 , n36484 , n36485 , n36486 , n36487 , n36488 , n36489 , n36490 , n36491 , n36492 , n36493 , n36494 , n36495 , n36496 , n36497 , n36498 , n36499 , n36500 , n36501 , n36502 , n36503 , n36504 , n36505 , n36506 , n36507 , n36508 , n36509 , n36510 , n36511 , n36512 , n36513 , n36514 , n36515 , n36516 , n36517 , n36518 , n36519 , n36520 , n36521 , n36522 , n36523 , n36524 , n36525 , n36526 , n36527 , n36528 , n36529 , n36530 , n36531 , n36532 , n36533 , n36534 , n36535 , n36536 , n36537 , n36538 , n36539 , n36540 , n36541 , n36542 , n36543 , n36544 , n36545 , n36546 , n36547 , n36548 , n36549 , n36550 , n36551 , n36552 , n36553 , n36554 , n36555 , n36556 , n36557 , n36558 , n36559 , n36560 , n36561 , n36562 , n36563 , n36564 , n36565 , n36566 , n36567 , n36568 , n36569 , n36570 , n36571 , n36572 , n36573 , n36574 , n36575 , n36576 , n36577 , n36578 , n36579 , n36580 , n36581 , n36582 , n36583 , n36584 , n36585 , n36586 , n36587 , n36588 , n36589 , n36590 , n36591 , n36592 , n36593 , n36594 , n36595 , n36596 , n36597 , n36598 , n36599 , n36600 , n36601 , n36602 , n36603 , n36604 , n36605 , n36606 , n36607 , n36608 , n36609 , n36610 , n36611 , n36612 , n36613 , n36614 , n36615 , n36616 , n36617 , n36618 , n36619 , n36620 , n36621 , n36622 , n36623 , n36624 , n36625 , n36626 , n36627 , n36628 , n36629 , n36630 , n36631 , n36632 , n36633 , n36634 , n36635 , n36636 , n36637 , n36638 , n36639 , n36640 , n36641 , n36642 , n36643 , n36644 , n36645 , n36646 , n36647 , n36648 , n36649 , n36650 , n36651 , n36652 , n36653 , n36654 , n36655 , n36656 , n36657 , n36658 , n36659 , n36660 , n36661 , n36662 , n36663 , n36664 , n36665 , n36666 , n36667 , n36668 , n36669 , n36670 , n36671 , n36672 , n36673 , n36674 , n36675 , n36676 , n36677 , n36678 , n36679 , n36680 , n36681 , n36682 , n36683 , n36684 , n36685 , n36686 , n36687 , n36688 , n36689 , n36690 , n36691 , n36692 , n36693 , n36694 , n36695 , n36696 , n36697 , n36698 , n36699 , n36700 , n36701 , n36702 , n36703 , n36704 , n36705 , n36706 , n36707 , n36708 , n36709 , n36710 , n36711 , n36712 , n36713 , n36714 , n36715 , n36716 , n36717 , n36718 , n36719 , n36720 , n36721 , n36722 , n36723 , n36724 , n36725 , n36726 , n36727 , n36728 , n36729 , n36730 , n36731 , n36732 , n36733 , n36734 , n36735 , n36736 , n36737 , n36738 , n36739 , n36740 , n36741 , n36742 , n36743 , n36744 , n36745 , n36746 , n36747 , n36748 , n36749 , n36750 , n36751 , n36752 , n36753 , n36754 , n36755 , n36756 , n36757 , n36758 , n36759 , n36760 , n36761 , n36762 , n36763 , n36764 , n36765 , n36766 , n36767 , n36768 , n36769 , n36770 , n36771 , n36772 , n36773 , n36774 , n36775 , n36776 , n36777 , n36778 , n36779 , n36780 , n36781 , n36782 , n36783 , n36784 , n36785 , n36786 , n36787 , n36788 , n36789 , n36790 , n36791 , n36792 , n36793 , n36794 , n36795 , n36796 , n36797 , n36798 , n36799 , n36800 , n36801 , n36802 , n36803 , n36804 , n36805 , n36806 , n36807 , n36808 , n36809 , n36810 , n36811 , n36812 , n36813 , n36814 , n36815 , n36816 , n36817 , n36818 , n36819 , n36820 , n36821 , n36822 , n36823 , n36824 , n36825 , n36826 , n36827 , n36828 , n36829 , n36830 , n36831 , n36832 , n36833 , n36834 , n36835 , n36836 , n36837 , n36838 , n36839 , n36840 , n36841 , n36842 , n36843 , n36844 , n36845 , n36846 , n36847 , n36848 , n36849 , n36850 , n36851 , n36852 , n36853 , n36854 , n36855 , n36856 , n36857 , n36858 , n36859 , n36860 , n36861 , n36862 , n36863 , n36864 , n36865 , n36866 , n36867 , n36868 , n36869 , n36870 , n36871 , n36872 , n36873 , n36874 , n36875 , n36876 , n36877 , n36878 , n36879 , n36880 , n36881 , n36882 , n36883 , n36884 , n36885 , n36886 , n36887 , n36888 , n36889 , n36890 , n36891 , n36892 , n36893 , n36894 , n36895 , n36896 , n36897 , n36898 , n36899 , n36900 , n36901 , n36902 , n36903 , n36904 , n36905 , n36906 , n36907 , n36908 , n36909 , n36910 , n36911 , n36912 , n36913 , n36914 , n36915 , n36916 , n36917 , n36918 , n36919 , n36920 , n36921 , n36922 , n36923 , n36924 , n36925 , n36926 , n36927 , n36928 , n36929 , n36930 , n36931 , n36932 , n36933 , n36934 , n36935 , n36936 , n36937 , n36938 , n36939 , n36940 , n36941 , n36942 , n36943 , n36944 , n36945 , n36946 , n36947 , n36948 , n36949 , n36950 , n36951 , n36952 , n36953 , n36954 , n36955 , n36956 , n36957 , n36958 , n36959 , n36960 , n36961 , n36962 , n36963 , n36964 , n36965 , n36966 , n36967 , n36968 , n36969 , n36970 , n36971 , n36972 , n36973 , n36974 , n36975 , n36976 , n36977 , n36978 , n36979 , n36980 , n36981 , n36982 , n36983 , n36984 , n36985 , n36986 , n36987 , n36988 , n36989 , n36990 , n36991 , n36992 , n36993 , n36994 , n36995 , n36996 , n36997 , n36998 , n36999 , n37000 , n37001 , n37002 , n37003 , n37004 , n37005 , n37006 , n37007 , n37008 , n37009 , n37010 , n37011 , n37012 , n37013 , n37014 , n37015 , n37016 , n37017 , n37018 , n37019 , n37020 , n37021 , n37022 , n37023 , n37024 , n37025 , n37026 , n37027 , n37028 , n37029 , n37030 , n37031 , n37032 , n37033 , n37034 , n37035 , n37036 , n37037 , n37038 , n37039 , n37040 , n37041 , n37042 , n37043 , n37044 , n37045 , n37046 , n37047 , n37048 , n37049 , n37050 , n37051 , n37052 , n37053 , n37054 , n37055 , n37056 , n37057 , n37058 , n37059 , n37060 , n37061 , n37062 , n37063 , n37064 , n37065 , n37066 , n37067 , n37068 , n37069 , n37070 , n37071 , n37072 , n37073 , n37074 , n37075 , n37076 , n37077 , n37078 , n37079 , n37080 , n37081 , n37082 , n37083 , n37084 , n37085 , n37086 , n37087 , n37088 , n37089 , n37090 , n37091 , n37092 , n37093 , n37094 , n37095 , n37096 , n37097 , n37098 , n37099 , n37100 , n37101 , n37102 , n37103 , n37104 , n37105 , n37106 , n37107 , n37108 , n37109 , n37110 , n37111 , n37112 , n37113 , n37114 , n37115 , n37116 , n37117 , n37118 , n37119 , n37120 , n37121 , n37122 , n37123 , n37124 , n37125 , n37126 , n37127 , n37128 , n37129 , n37130 , n37131 , n37132 , n37133 , n37134 , n37135 , n37136 , n37137 , n37138 , n37139 , n37140 , n37141 , n37142 , n37143 , n37144 , n37145 , n37146 , n37147 , n37148 , n37149 , n37150 , n37151 , n37152 , n37153 , n37154 , n37155 , n37156 , n37157 , n37158 , n37159 , n37160 , n37161 , n37162 , n37163 , n37164 , n37165 , n37166 , n37167 , n37168 , n37169 , n37170 , n37171 , n37172 , n37173 , n37174 , n37175 , n37176 , n37177 , n37178 , n37179 , n37180 , n37181 , n37182 , n37183 , n37184 , n37185 , n37186 , n37187 , n37188 , n37189 , n37190 , n37191 , n37192 , n37193 , n37194 , n37195 , n37196 , n37197 , n37198 , n37199 , n37200 , n37201 , n37202 , n37203 , n37204 , n37205 , n37206 , n37207 , n37208 , n37209 , n37210 , n37211 , n37212 , n37213 , n37214 , n37215 , n37216 , n37217 , n37218 , n37219 , n37220 , n37221 , n37222 , n37223 , n37224 , n37225 , n37226 , n37227 , n37228 , n37229 , n37230 , n37231 , n37232 , n37233 , n37234 , n37235 , n37236 , n37237 , n37238 , n37239 , n37240 , n37241 , n37242 , n37243 , n37244 , n37245 , n37246 , n37247 , n37248 , n37249 , n37250 , n37251 , n37252 , n37253 , n37254 , n37255 , n37256 , n37257 , n37258 , n37259 , n37260 , n37261 , n37262 , n37263 , n37264 , n37265 , n37266 , n37267 , n37268 , n37269 , n37270 , n37271 , n37272 , n37273 , n37274 , n37275 , n37276 , n37277 , n37278 , n37279 , n37280 , n37281 , n37282 , n37283 , n37284 , n37285 , n37286 , n37287 , n37288 , n37289 , n37290 , n37291 , n37292 , n37293 , n37294 , n37295 , n37296 , n37297 , n37298 , n37299 , n37300 , n37301 , n37302 , n37303 , n37304 , n37305 , n37306 , n37307 , n37308 , n37309 , n37310 , n37311 , n37312 , n37313 , n37314 , n37315 , n37316 , n37317 , n37318 , n37319 , n37320 , n37321 , n37322 , n37323 , n37324 , n37325 , n37326 , n37327 , n37328 , n37329 , n37330 , n37331 , n37332 , n37333 , n37334 , n37335 , n37336 , n37337 , n37338 , n37339 , n37340 , n37341 , n37342 , n37343 , n37344 , n37345 , n37346 , n37347 , n37348 , n37349 , n37350 , n37351 , n37352 , n37353 , n37354 , n37355 , n37356 , n37357 , n37358 , n37359 , n37360 , n37361 , n37362 , n37363 , n37364 , n37365 , n37366 , n37367 , n37368 , n37369 , n37370 , n37371 , n37372 , n37373 , n37374 , n37375 , n37376 , n37377 , n37378 , n37379 , n37380 , n37381 , n37382 , n37383 , n37384 , n37385 , n37386 , n37387 , n37388 , n37389 , n37390 , n37391 , n37392 , n37393 , n37394 , n37395 , n37396 , n37397 , n37398 , n37399 , n37400 , n37401 , n37402 , n37403 , n37404 , n37405 , n37406 , n37407 , n37408 , n37409 , n37410 , n37411 , n37412 , n37413 , n37414 , n37415 , n37416 , n37417 , n37418 , n37419 , n37420 , n37421 , n37422 , n37423 , n37424 , n37425 , n37426 , n37427 , n37428 , n37429 , n37430 , n37431 , n37432 , n37433 , n37434 , n37435 , n37436 , n37437 , n37438 , n37439 , n37440 , n37441 , n37442 , n37443 , n37444 , n37445 , n37446 , n37447 , n37448 , n37449 , n37450 , n37451 , n37452 , n37453 , n37454 , n37455 , n37456 , n37457 , n37458 , n37459 , n37460 , n37461 , n37462 , n37463 , n37464 , n37465 , n37466 , n37467 , n37468 , n37469 , n37470 , n37471 , n37472 , n37473 , n37474 , n37475 , n37476 , n37477 , n37478 , n37479 , n37480 , n37481 , n37482 , n37483 , n37484 , n37485 , n37486 , n37487 , n37488 , n37489 , n37490 , n37491 , n37492 , n37493 , n37494 , n37495 , n37496 , n37497 , n37498 , n37499 , n37500 , n37501 , n37502 , n37503 , n37504 , n37505 , n37506 , n37507 , n37508 , n37509 , n37510 , n37511 , n37512 , n37513 , n37514 , n37515 , n37516 , n37517 , n37518 , n37519 , n37520 , n37521 , n37522 , n37523 , n37524 , n37525 , n37526 , n37527 , n37528 , n37529 , n37530 , n37531 , n37532 , n37533 , n37534 , n37535 , n37536 , n37537 , n37538 , n37539 , n37540 , n37541 , n37542 , n37543 , n37544 , n37545 , n37546 , n37547 , n37548 , n37549 , n37550 , n37551 , n37552 , n37553 , n37554 , n37555 , n37556 , n37557 , n37558 , n37559 , n37560 , n37561 , n37562 , n37563 , n37564 , n37565 , n37566 , n37567 , n37568 , n37569 , n37570 , n37571 , n37572 , n37573 , n37574 , n37575 , n37576 , n37577 , n37578 , n37579 , n37580 , n37581 , n37582 , n37583 , n37584 , n37585 , n37586 , n37587 , n37588 , n37589 , n37590 , n37591 , n37592 , n37593 , n37594 , n37595 , n37596 , n37597 , n37598 , n37599 , n37600 , n37601 , n37602 , n37603 , n37604 , n37605 , n37606 , n37607 , n37608 , n37609 , n37610 , n37611 , n37612 , n37613 , n37614 , n37615 , n37616 , n37617 , n37618 , n37619 , n37620 , n37621 , n37622 , n37623 , n37624 , n37625 , n37626 , n37627 , n37628 , n37629 , n37630 , n37631 , n37632 , n37633 , n37634 , n37635 , n37636 , n37637 , n37638 , n37639 , n37640 , n37641 , n37642 , n37643 , n37644 , n37645 , n37646 , n37647 , n37648 , n37649 , n37650 , n37651 , n37652 , n37653 , n37654 , n37655 , n37656 , n37657 , n37658 , n37659 , n37660 , n37661 , n37662 , n37663 , n37664 , n37665 , n37666 , n37667 , n37668 , n37669 , n37670 , n37671 , n37672 , n37673 , n37674 , n37675 , n37676 , n37677 , n37678 , n37679 , n37680 , n37681 , n37682 , n37683 , n37684 , n37685 , n37686 , n37687 , n37688 , n37689 , n37690 , n37691 , n37692 , n37693 , n37694 , n37695 , n37696 , n37697 , n37698 , n37699 , n37700 , n37701 , n37702 , n37703 , n37704 , n37705 , n37706 , n37707 , n37708 , n37709 , n37710 , n37711 , n37712 , n37713 , n37714 , n37715 , n37716 , n37717 , n37718 , n37719 , n37720 , n37721 , n37722 , n37723 , n37724 , n37725 , n37726 , n37727 , n37728 , n37729 , n37730 , n37731 , n37732 , n37733 , n37734 , n37735 , n37736 , n37737 , n37738 , n37739 , n37740 , n37741 , n37742 , n37743 , n37744 , n37745 , n37746 , n37747 , n37748 , n37749 , n37750 , n37751 , n37752 , n37753 , n37754 , n37755 , n37756 , n37757 , n37758 , n37759 , n37760 , n37761 , n37762 , n37763 , n37764 , n37765 , n37766 , n37767 , n37768 , n37769 , n37770 , n37771 , n37772 , n37773 , n37774 , n37775 , n37776 , n37777 , n37778 , n37779 , n37780 , n37781 , n37782 , n37783 , n37784 , n37785 , n37786 , n37787 , n37788 , n37789 , n37790 , n37791 , n37792 , n37793 , n37794 , n37795 , n37796 , n37797 , n37798 , n37799 , n37800 , n37801 , n37802 , n37803 , n37804 , n37805 , n37806 , n37807 , n37808 , n37809 , n37810 , n37811 , n37812 , n37813 , n37814 , n37815 , n37816 , n37817 , n37818 , n37819 , n37820 , n37821 , n37822 , n37823 , n37824 , n37825 , n37826 , n37827 , n37828 , n37829 , n37830 , n37831 , n37832 , n37833 , n37834 , n37835 , n37836 , n37837 , n37838 , n37839 , n37840 , n37841 , n37842 , n37843 , n37844 , n37845 , n37846 , n37847 , n37848 , n37849 , n37850 , n37851 , n37852 , n37853 , n37854 , n37855 , n37856 , n37857 , n37858 , n37859 , n37860 , n37861 , n37862 , n37863 , n37864 , n37865 , n37866 , n37867 , n37868 , n37869 , n37870 , n37871 , n37872 , n37873 , n37874 , n37875 , n37876 , n37877 , n37878 , n37879 , n37880 , n37881 , n37882 , n37883 , n37884 , n37885 , n37886 , n37887 , n37888 , n37889 , n37890 , n37891 , n37892 , n37893 , n37894 , n37895 , n37896 , n37897 , n37898 , n37899 , n37900 , n37901 , n37902 , n37903 , n37904 , n37905 , n37906 , n37907 , n37908 , n37909 , n37910 , n37911 , n37912 , n37913 , n37914 , n37915 , n37916 , n37917 , n37918 , n37919 , n37920 , n37921 , n37922 , n37923 , n37924 , n37925 , n37926 , n37927 , n37928 , n37929 , n37930 , n37931 , n37932 , n37933 , n37934 , n37935 , n37936 , n37937 , n37938 , n37939 , n37940 , n37941 , n37942 , n37943 , n37944 , n37945 , n37946 , n37947 , n37948 , n37949 , n37950 , n37951 , n37952 , n37953 , n37954 , n37955 , n37956 , n37957 , n37958 , n37959 , n37960 , n37961 , n37962 , n37963 , n37964 , n37965 , n37966 , n37967 , n37968 , n37969 , n37970 , n37971 , n37972 , n37973 , n37974 , n37975 , n37976 , n37977 , n37978 , n37979 , n37980 , n37981 , n37982 , n37983 , n37984 , n37985 , n37986 , n37987 , n37988 , n37989 , n37990 , n37991 , n37992 , n37993 , n37994 , n37995 , n37996 , n37997 , n37998 , n37999 , n38000 , n38001 , n38002 , n38003 , n38004 , n38005 , n38006 , n38007 , n38008 , n38009 , n38010 , n38011 , n38012 , n38013 , n38014 , n38015 , n38016 , n38017 , n38018 , n38019 , n38020 , n38021 , n38022 , n38023 , n38024 , n38025 , n38026 , n38027 , n38028 , n38029 , n38030 , n38031 , n38032 , n38033 , n38034 , n38035 , n38036 , n38037 , n38038 , n38039 , n38040 , n38041 , n38042 , n38043 , n38044 , n38045 , n38046 , n38047 , n38048 , n38049 , n38050 , n38051 , n38052 , n38053 , n38054 , n38055 , n38056 , n38057 , n38058 , n38059 , n38060 , n38061 , n38062 , n38063 , n38064 , n38065 , n38066 , n38067 , n38068 , n38069 , n38070 , n38071 , n38072 , n38073 , n38074 , n38075 , n38076 , n38077 , n38078 , n38079 , n38080 , n38081 , n38082 , n38083 , n38084 , n38085 , n38086 , n38087 , n38088 , n38089 , n38090 , n38091 , n38092 , n38093 , n38094 , n38095 , n38096 , n38097 , n38098 , n38099 , n38100 , n38101 , n38102 , n38103 , n38104 , n38105 , n38106 , n38107 , n38108 , n38109 , n38110 , n38111 , n38112 , n38113 , n38114 , n38115 , n38116 , n38117 , n38118 , n38119 , n38120 , n38121 , n38122 , n38123 , n38124 , n38125 , n38126 , n38127 , n38128 , n38129 , n38130 , n38131 , n38132 , n38133 , n38134 , n38135 , n38136 , n38137 , n38138 , n38139 , n38140 , n38141 , n38142 , n38143 , n38144 , n38145 , n38146 , n38147 , n38148 , n38149 , n38150 , n38151 , n38152 , n38153 , n38154 , n38155 , n38156 , n38157 , n38158 , n38159 , n38160 , n38161 , n38162 , n38163 , n38164 , n38165 , n38166 , n38167 , n38168 , n38169 , n38170 , n38171 , n38172 , n38173 , n38174 , n38175 , n38176 , n38177 , n38178 , n38179 , n38180 , n38181 , n38182 , n38183 , n38184 , n38185 , n38186 , n38187 , n38188 , n38189 , n38190 , n38191 , n38192 , n38193 , n38194 , n38195 , n38196 , n38197 , n38198 , n38199 , n38200 , n38201 , n38202 , n38203 , n38204 , n38205 , n38206 , n38207 , n38208 , n38209 , n38210 , n38211 , n38212 , n38213 , n38214 , n38215 , n38216 , n38217 , n38218 , n38219 , n38220 , n38221 , n38222 , n38223 , n38224 , n38225 , n38226 , n38227 , n38228 , n38229 , n38230 , n38231 , n38232 , n38233 , n38234 , n38235 , n38236 , n38237 , n38238 , n38239 , n38240 , n38241 , n38242 , n38243 , n38244 , n38245 , n38246 , n38247 , n38248 , n38249 , n38250 , n38251 , n38252 , n38253 , n38254 , n38255 , n38256 , n38257 , n38258 , n38259 , n38260 , n38261 , n38262 , n38263 , n38264 , n38265 , n38266 , n38267 , n38268 , n38269 , n38270 , n38271 , n38272 , n38273 , n38274 , n38275 , n38276 , n38277 , n38278 , n38279 , n38280 , n38281 , n38282 , n38283 , n38284 , n38285 , n38286 , n38287 , n38288 , n38289 , n38290 , n38291 , n38292 , n38293 , n38294 , n38295 , n38296 , n38297 , n38298 , n38299 , n38300 , n38301 , n38302 , n38303 , n38304 , n38305 , n38306 , n38307 , n38308 , n38309 , n38310 , n38311 , n38312 , n38313 , n38314 , n38315 , n38316 , n38317 , n38318 , n38319 , n38320 , n38321 , n38322 , n38323 , n38324 , n38325 , n38326 , n38327 , n38328 , n38329 , n38330 , n38331 , n38332 , n38333 , n38334 , n38335 , n38336 , n38337 , n38338 , n38339 , n38340 , n38341 , n38342 , n38343 , n38344 , n38345 , n38346 , n38347 , n38348 , n38349 , n38350 , n38351 , n38352 , n38353 , n38354 , n38355 , n38356 , n38357 , n38358 , n38359 , n38360 , n38361 , n38362 , n38363 , n38364 , n38365 , n38366 , n38367 , n38368 , n38369 , n38370 , n38371 , n38372 , n38373 , n38374 , n38375 , n38376 , n38377 , n38378 , n38379 , n38380 , n38381 , n38382 , n38383 , n38384 , n38385 , n38386 , n38387 , n38388 , n38389 , n38390 , n38391 , n38392 , n38393 , n38394 , n38395 , n38396 , n38397 , n38398 , n38399 , n38400 , n38401 , n38402 , n38403 , n38404 , n38405 , n38406 , n38407 , n38408 , n38409 , n38410 , n38411 , n38412 , n38413 , n38414 , n38415 , n38416 , n38417 , n38418 , n38419 , n38420 , n38421 , n38422 , n38423 , n38424 , n38425 , n38426 , n38427 , n38428 , n38429 , n38430 , n38431 , n38432 , n38433 , n38434 , n38435 , n38436 , n38437 , n38438 , n38439 , n38440 , n38441 , n38442 , n38443 , n38444 , n38445 , n38446 , n38447 , n38448 , n38449 , n38450 , n38451 , n38452 , n38453 , n38454 , n38455 , n38456 , n38457 , n38458 , n38459 , n38460 , n38461 , n38462 , n38463 , n38464 , n38465 , n38466 , n38467 , n38468 , n38469 , n38470 , n38471 , n38472 , n38473 , n38474 , n38475 , n38476 , n38477 , n38478 , n38479 , n38480 , n38481 , n38482 , n38483 , n38484 , n38485 , n38486 , n38487 , n38488 , n38489 , n38490 , n38491 , n38492 , n38493 , n38494 , n38495 , n38496 , n38497 , n38498 , n38499 , n38500 , n38501 , n38502 , n38503 , n38504 , n38505 , n38506 , n38507 , n38508 , n38509 , n38510 , n38511 , n38512 , n38513 , n38514 , n38515 , n38516 , n38517 , n38518 , n38519 , n38520 , n38521 , n38522 , n38523 , n38524 , n38525 , n38526 , n38527 , n38528 , n38529 , n38530 , n38531 , n38532 , n38533 , n38534 , n38535 , n38536 , n38537 , n38538 , n38539 , n38540 , n38541 , n38542 , n38543 , n38544 , n38545 , n38546 , n38547 , n38548 , n38549 , n38550 , n38551 , n38552 , n38553 , n38554 , n38555 , n38556 , n38557 , n38558 , n38559 , n38560 , n38561 , n38562 , n38563 , n38564 , n38565 , n38566 , n38567 , n38568 , n38569 , n38570 , n38571 , n38572 , n38573 , n38574 , n38575 , n38576 , n38577 , n38578 , n38579 , n38580 , n38581 , n38582 , n38583 , n38584 , n38585 , n38586 , n38587 , n38588 , n38589 , n38590 , n38591 , n38592 , n38593 , n38594 , n38595 , n38596 , n38597 , n38598 , n38599 , n38600 , n38601 , n38602 , n38603 , n38604 , n38605 , n38606 , n38607 , n38608 , n38609 , n38610 , n38611 , n38612 , n38613 , n38614 , n38615 , n38616 , n38617 , n38618 , n38619 , n38620 , n38621 , n38622 , n38623 , n38624 , n38625 , n38626 , n38627 , n38628 , n38629 , n38630 , n38631 , n38632 , n38633 , n38634 , n38635 , n38636 , n38637 , n38638 , n38639 , n38640 , n38641 , n38642 , n38643 , n38644 , n38645 , n38646 , n38647 , n38648 , n38649 , n38650 , n38651 , n38652 , n38653 , n38654 , n38655 , n38656 , n38657 , n38658 , n38659 , n38660 , n38661 , n38662 , n38663 , n38664 , n38665 , n38666 , n38667 , n38668 , n38669 , n38670 , n38671 , n38672 , n38673 , n38674 , n38675 , n38676 , n38677 , n38678 , n38679 , n38680 , n38681 , n38682 , n38683 , n38684 , n38685 , n38686 , n38687 , n38688 , n38689 , n38690 , n38691 , n38692 , n38693 , n38694 , n38695 , n38696 , n38697 , n38698 , n38699 , n38700 , n38701 , n38702 , n38703 , n38704 , n38705 , n38706 , n38707 , n38708 , n38709 , n38710 , n38711 , n38712 , n38713 , n38714 , n38715 , n38716 , n38717 , n38718 , n38719 , n38720 , n38721 , n38722 , n38723 , n38724 , n38725 , n38726 , n38727 , n38728 , n38729 , n38730 , n38731 , n38732 , n38733 , n38734 , n38735 , n38736 , n38737 , n38738 , n38739 , n38740 , n38741 , n38742 , n38743 , n38744 , n38745 , n38746 , n38747 , n38748 , n38749 , n38750 , n38751 , n38752 , n38753 , n38754 , n38755 , n38756 , n38757 , n38758 , n38759 , n38760 , n38761 , n38762 , n38763 , n38764 , n38765 , n38766 , n38767 , n38768 , n38769 , n38770 , n38771 , n38772 , n38773 , n38774 , n38775 , n38776 , n38777 , n38778 , n38779 , n38780 , n38781 , n38782 , n38783 , n38784 , n38785 , n38786 , n38787 , n38788 , n38789 , n38790 , n38791 , n38792 , n38793 , n38794 , n38795 , n38796 , n38797 , n38798 , n38799 , n38800 , n38801 , n38802 , n38803 , n38804 , n38805 , n38806 , n38807 , n38808 , n38809 , n38810 , n38811 , n38812 , n38813 , n38814 , n38815 , n38816 , n38817 , n38818 , n38819 , n38820 , n38821 , n38822 , n38823 , n38824 , n38825 , n38826 , n38827 , n38828 , n38829 , n38830 , n38831 , n38832 , n38833 , n38834 , n38835 , n38836 , n38837 , n38838 , n38839 , n38840 , n38841 , n38842 , n38843 , n38844 , n38845 , n38846 , n38847 , n38848 , n38849 , n38850 , n38851 , n38852 , n38853 , n38854 , n38855 , n38856 , n38857 , n38858 , n38859 , n38860 , n38861 , n38862 , n38863 , n38864 , n38865 , n38866 , n38867 , n38868 , n38869 , n38870 , n38871 , n38872 , n38873 , n38874 , n38875 , n38876 , n38877 , n38878 , n38879 , n38880 , n38881 , n38882 , n38883 , n38884 , n38885 , n38886 , n38887 , n38888 , n38889 , n38890 , n38891 , n38892 , n38893 , n38894 , n38895 , n38896 , n38897 , n38898 , n38899 , n38900 , n38901 , n38902 , n38903 , n38904 , n38905 , n38906 , n38907 , n38908 , n38909 , n38910 , n38911 , n38912 , n38913 , n38914 , n38915 , n38916 , n38917 , n38918 , n38919 , n38920 , n38921 , n38922 , n38923 , n38924 , n38925 , n38926 , n38927 , n38928 , n38929 , n38930 , n38931 , n38932 , n38933 , n38934 , n38935 , n38936 , n38937 , n38938 , n38939 , n38940 , n38941 , n38942 , n38943 , n38944 , n38945 , n38946 , n38947 , n38948 , n38949 , n38950 , n38951 , n38952 , n38953 , n38954 , n38955 , n38956 , n38957 , n38958 , n38959 , n38960 , n38961 , n38962 , n38963 , n38964 , n38965 , n38966 , n38967 , n38968 , n38969 , n38970 , n38971 , n38972 , n38973 , n38974 , n38975 , n38976 , n38977 , n38978 , n38979 , n38980 , n38981 , n38982 , n38983 , n38984 , n38985 , n38986 , n38987 , n38988 , n38989 , n38990 , n38991 , n38992 , n38993 , n38994 , n38995 , n38996 , n38997 , n38998 , n38999 , n39000 , n39001 , n39002 , n39003 , n39004 , n39005 , n39006 , n39007 , n39008 , n39009 , n39010 , n39011 , n39012 , n39013 , n39014 , n39015 , n39016 , n39017 , n39018 , n39019 , n39020 , n39021 , n39022 , n39023 , n39024 , n39025 , n39026 , n39027 , n39028 , n39029 , n39030 , n39031 , n39032 , n39033 , n39034 , n39035 , n39036 , n39037 , n39038 , n39039 , n39040 , n39041 , n39042 , n39043 , n39044 , n39045 , n39046 , n39047 , n39048 , n39049 , n39050 , n39051 , n39052 , n39053 , n39054 , n39055 , n39056 , n39057 , n39058 , n39059 , n39060 , n39061 , n39062 , n39063 , n39064 , n39065 , n39066 , n39067 , n39068 , n39069 , n39070 , n39071 , n39072 , n39073 , n39074 , n39075 , n39076 , n39077 , n39078 , n39079 , n39080 , n39081 , n39082 , n39083 , n39084 , n39085 , n39086 , n39087 , n39088 , n39089 , n39090 , n39091 , n39092 , n39093 , n39094 , n39095 , n39096 , n39097 , n39098 , n39099 , n39100 , n39101 , n39102 , n39103 , n39104 , n39105 , n39106 , n39107 , n39108 , n39109 , n39110 , n39111 , n39112 , n39113 , n39114 , n39115 , n39116 , n39117 , n39118 , n39119 , n39120 , n39121 , n39122 , n39123 , n39124 , n39125 , n39126 , n39127 , n39128 , n39129 , n39130 , n39131 , n39132 , n39133 , n39134 , n39135 , n39136 , n39137 , n39138 , n39139 , n39140 , n39141 , n39142 , n39143 , n39144 , n39145 , n39146 , n39147 , n39148 , n39149 , n39150 , n39151 , n39152 , n39153 , n39154 , n39155 , n39156 , n39157 , n39158 , n39159 , n39160 , n39161 , n39162 , n39163 , n39164 , n39165 , n39166 , n39167 , n39168 , n39169 , n39170 , n39171 , n39172 , n39173 , n39174 , n39175 , n39176 , n39177 , n39178 , n39179 , n39180 , n39181 , n39182 , n39183 , n39184 , n39185 , n39186 , n39187 , n39188 , n39189 , n39190 , n39191 , n39192 , n39193 , n39194 , n39195 , n39196 , n39197 , n39198 , n39199 , n39200 , n39201 , n39202 , n39203 , n39204 , n39205 , n39206 , n39207 , n39208 , n39209 , n39210 , n39211 , n39212 , n39213 , n39214 , n39215 , n39216 , n39217 , n39218 , n39219 , n39220 , n39221 , n39222 , n39223 , n39224 , n39225 , n39226 , n39227 , n39228 , n39229 , n39230 , n39231 , n39232 , n39233 , n39234 , n39235 , n39236 , n39237 , n39238 , n39239 , n39240 , n39241 , n39242 , n39243 , n39244 , n39245 , n39246 , n39247 , n39248 , n39249 , n39250 , n39251 , n39252 , n39253 , n39254 , n39255 , n39256 , n39257 , n39258 , n39259 , n39260 , n39261 , n39262 , n39263 , n39264 , n39265 , n39266 , n39267 , n39268 , n39269 , n39270 , n39271 , n39272 , n39273 , n39274 , n39275 , n39276 , n39277 , n39278 , n39279 , n39280 , n39281 , n39282 , n39283 , n39284 , n39285 , n39286 , n39287 , n39288 , n39289 , n39290 , n39291 , n39292 , n39293 , n39294 , n39295 , n39296 , n39297 , n39298 , n39299 , n39300 , n39301 , n39302 , n39303 , n39304 , n39305 , n39306 , n39307 , n39308 , n39309 , n39310 , n39311 , n39312 , n39313 , n39314 , n39315 , n39316 , n39317 , n39318 , n39319 , n39320 , n39321 , n39322 , n39323 , n39324 , n39325 , n39326 , n39327 , n39328 , n39329 , n39330 , n39331 , n39332 , n39333 , n39334 , n39335 , n39336 , n39337 , n39338 , n39339 , n39340 , n39341 , n39342 , n39343 , n39344 , n39345 , n39346 , n39347 , n39348 , n39349 , n39350 , n39351 , n39352 , n39353 , n39354 , n39355 , n39356 , n39357 , n39358 , n39359 , n39360 , n39361 , n39362 , n39363 , n39364 , n39365 , n39366 , n39367 , n39368 , n39369 , n39370 , n39371 , n39372 , n39373 , n39374 , n39375 , n39376 , n39377 , n39378 , n39379 , n39380 , n39381 , n39382 , n39383 , n39384 , n39385 , n39386 , n39387 , n39388 , n39389 , n39390 , n39391 , n39392 , n39393 , n39394 , n39395 , n39396 , n39397 , n39398 , n39399 , n39400 , n39401 , n39402 , n39403 , n39404 , n39405 , n39406 , n39407 , n39408 , n39409 , n39410 , n39411 , n39412 , n39413 , n39414 , n39415 , n39416 , n39417 , n39418 , n39419 , n39420 , n39421 , n39422 , n39423 , n39424 , n39425 , n39426 , n39427 , n39428 , n39429 , n39430 , n39431 , n39432 , n39433 , n39434 , n39435 , n39436 , n39437 , n39438 , n39439 , n39440 , n39441 , n39442 , n39443 , n39444 , n39445 , n39446 , n39447 , n39448 , n39449 , n39450 , n39451 , n39452 , n39453 , n39454 , n39455 , n39456 , n39457 , n39458 , n39459 , n39460 , n39461 , n39462 , n39463 , n39464 , n39465 , n39466 , n39467 , n39468 , n39469 , n39470 , n39471 , n39472 , n39473 , n39474 , n39475 , n39476 , n39477 , n39478 , n39479 , n39480 , n39481 , n39482 , n39483 , n39484 , n39485 , n39486 , n39487 , n39488 , n39489 , n39490 , n39491 , n39492 , n39493 , n39494 , n39495 , n39496 , n39497 , n39498 , n39499 , n39500 , n39501 , n39502 , n39503 , n39504 , n39505 , n39506 , n39507 , n39508 , n39509 , n39510 , n39511 , n39512 , n39513 , n39514 , n39515 , n39516 , n39517 , n39518 , n39519 , n39520 , n39521 , n39522 , n39523 , n39524 , n39525 , n39526 , n39527 , n39528 , n39529 , n39530 , n39531 , n39532 , n39533 , n39534 , n39535 , n39536 , n39537 , n39538 , n39539 , n39540 , n39541 , n39542 , n39543 , n39544 , n39545 , n39546 , n39547 , n39548 , n39549 , n39550 , n39551 , n39552 , n39553 , n39554 , n39555 , n39556 , n39557 , n39558 , n39559 , n39560 , n39561 , n39562 , n39563 , n39564 , n39565 , n39566 , n39567 , n39568 , n39569 , n39570 , n39571 , n39572 , n39573 , n39574 , n39575 , n39576 , n39577 , n39578 , n39579 , n39580 , n39581 , n39582 , n39583 , n39584 , n39585 , n39586 , n39587 , n39588 , n39589 , n39590 , n39591 , n39592 , n39593 , n39594 , n39595 , n39596 , n39597 , n39598 , n39599 , n39600 , n39601 , n39602 , n39603 , n39604 , n39605 , n39606 , n39607 , n39608 , n39609 , n39610 , n39611 , n39612 , n39613 , n39614 , n39615 , n39616 , n39617 , n39618 , n39619 , n39620 , n39621 , n39622 , n39623 , n39624 , n39625 , n39626 , n39627 , n39628 , n39629 , n39630 , n39631 , n39632 , n39633 , n39634 , n39635 , n39636 , n39637 , n39638 , n39639 , n39640 , n39641 , n39642 , n39643 , n39644 , n39645 , n39646 , n39647 , n39648 , n39649 , n39650 , n39651 , n39652 , n39653 , n39654 , n39655 , n39656 , n39657 , n39658 , n39659 , n39660 , n39661 , n39662 , n39663 , n39664 , n39665 , n39666 , n39667 , n39668 , n39669 , n39670 , n39671 , n39672 , n39673 , n39674 , n39675 , n39676 , n39677 , n39678 , n39679 , n39680 , n39681 , n39682 , n39683 , n39684 , n39685 , n39686 , n39687 , n39688 , n39689 , n39690 , n39691 , n39692 , n39693 , n39694 , n39695 , n39696 , n39697 , n39698 , n39699 , n39700 , n39701 , n39702 , n39703 , n39704 , n39705 , n39706 , n39707 , n39708 , n39709 , n39710 , n39711 , n39712 , n39713 , n39714 , n39715 , n39716 , n39717 , n39718 , n39719 , n39720 , n39721 , n39722 , n39723 , n39724 , n39725 , n39726 , n39727 , n39728 , n39729 , n39730 , n39731 , n39732 , n39733 , n39734 , n39735 , n39736 , n39737 , n39738 , n39739 , n39740 , n39741 , n39742 , n39743 , n39744 , n39745 , n39746 , n39747 , n39748 , n39749 , n39750 , n39751 , n39752 , n39753 , n39754 , n39755 , n39756 , n39757 , n39758 , n39759 , n39760 , n39761 , n39762 , n39763 , n39764 , n39765 , n39766 , n39767 , n39768 , n39769 , n39770 , n39771 , n39772 , n39773 , n39774 , n39775 , n39776 , n39777 , n39778 , n39779 , n39780 , n39781 , n39782 , n39783 , n39784 , n39785 , n39786 , n39787 , n39788 , n39789 , n39790 , n39791 , n39792 , n39793 , n39794 , n39795 , n39796 , n39797 , n39798 , n39799 , n39800 , n39801 , n39802 , n39803 , n39804 , n39805 , n39806 , n39807 , n39808 , n39809 , n39810 , n39811 , n39812 , n39813 , n39814 , n39815 , n39816 , n39817 , n39818 , n39819 , n39820 , n39821 , n39822 , n39823 , n39824 , n39825 , n39826 , n39827 , n39828 , n39829 , n39830 , n39831 , n39832 , n39833 , n39834 , n39835 , n39836 , n39837 , n39838 , n39839 , n39840 , n39841 , n39842 , n39843 , n39844 , n39845 , n39846 , n39847 , n39848 , n39849 , n39850 , n39851 , n39852 , n39853 , n39854 , n39855 , n39856 , n39857 , n39858 , n39859 , n39860 , n39861 , n39862 , n39863 , n39864 , n39865 , n39866 , n39867 , n39868 , n39869 , n39870 , n39871 , n39872 , n39873 , n39874 , n39875 , n39876 , n39877 , n39878 , n39879 , n39880 , n39881 , n39882 , n39883 , n39884 , n39885 , n39886 , n39887 , n39888 , n39889 , n39890 , n39891 , n39892 , n39893 , n39894 , n39895 , n39896 , n39897 , n39898 , n39899 , n39900 , n39901 , n39902 , n39903 , n39904 , n39905 , n39906 , n39907 , n39908 , n39909 , n39910 , n39911 , n39912 , n39913 , n39914 , n39915 , n39916 , n39917 , n39918 , n39919 , n39920 , n39921 , n39922 , n39923 , n39924 , n39925 , n39926 , n39927 , n39928 , n39929 , n39930 , n39931 , n39932 , n39933 , n39934 , n39935 , n39936 , n39937 , n39938 , n39939 , n39940 , n39941 , n39942 , n39943 , n39944 , n39945 , n39946 , n39947 , n39948 , n39949 , n39950 , n39951 , n39952 , n39953 , n39954 , n39955 , n39956 , n39957 , n39958 , n39959 , n39960 , n39961 , n39962 , n39963 , n39964 , n39965 , n39966 , n39967 , n39968 , n39969 , n39970 , n39971 , n39972 , n39973 , n39974 , n39975 , n39976 , n39977 , n39978 , n39979 , n39980 , n39981 , n39982 , n39983 , n39984 , n39985 , n39986 , n39987 , n39988 , n39989 , n39990 , n39991 , n39992 , n39993 , n39994 , n39995 , n39996 , n39997 , n39998 , n39999 , n40000 , n40001 , n40002 , n40003 , n40004 , n40005 , n40006 , n40007 , n40008 , n40009 , n40010 , n40011 , n40012 , n40013 , n40014 , n40015 , n40016 , n40017 , n40018 , n40019 , n40020 , n40021 , n40022 , n40023 , n40024 , n40025 , n40026 , n40027 , n40028 , n40029 , n40030 , n40031 , n40032 , n40033 , n40034 , n40035 , n40036 , n40037 , n40038 , n40039 , n40040 , n40041 , n40042 , n40043 , n40044 , n40045 , n40046 , n40047 , n40048 , n40049 , n40050 , n40051 , n40052 , n40053 , n40054 , n40055 , n40056 , n40057 , n40058 , n40059 , n40060 , n40061 , n40062 , n40063 , n40064 , n40065 , n40066 , n40067 , n40068 , n40069 , n40070 , n40071 , n40072 , n40073 , n40074 , n40075 , n40076 , n40077 , n40078 , n40079 , n40080 , n40081 , n40082 , n40083 , n40084 , n40085 , n40086 , n40087 , n40088 , n40089 , n40090 , n40091 , n40092 , n40093 , n40094 , n40095 , n40096 , n40097 , n40098 , n40099 , n40100 , n40101 , n40102 , n40103 , n40104 , n40105 , n40106 , n40107 , n40108 , n40109 , n40110 , n40111 , n40112 , n40113 , n40114 , n40115 , n40116 , n40117 , n40118 , n40119 , n40120 , n40121 , n40122 , n40123 , n40124 , n40125 , n40126 , n40127 , n40128 , n40129 , n40130 , n40131 , n40132 , n40133 , n40134 , n40135 , n40136 , n40137 , n40138 , n40139 , n40140 , n40141 , n40142 , n40143 , n40144 , n40145 , n40146 , n40147 , n40148 , n40149 , n40150 , n40151 , n40152 , n40153 , n40154 , n40155 , n40156 , n40157 , n40158 , n40159 , n40160 , n40161 , n40162 , n40163 , n40164 , n40165 , n40166 , n40167 , n40168 , n40169 , n40170 , n40171 , n40172 , n40173 , n40174 , n40175 , n40176 , n40177 , n40178 , n40179 , n40180 , n40181 , n40182 , n40183 , n40184 , n40185 , n40186 , n40187 , n40188 , n40189 , n40190 , n40191 , n40192 , n40193 , n40194 , n40195 , n40196 , n40197 , n40198 , n40199 , n40200 , n40201 , n40202 , n40203 , n40204 , n40205 , n40206 , n40207 , n40208 , n40209 , n40210 , n40211 , n40212 , n40213 , n40214 , n40215 , n40216 , n40217 , n40218 , n40219 , n40220 , n40221 , n40222 , n40223 , n40224 , n40225 , n40226 , n40227 , n40228 , n40229 , n40230 , n40231 , n40232 , n40233 , n40234 , n40235 , n40236 , n40237 , n40238 , n40239 , n40240 , n40241 , n40242 , n40243 , n40244 , n40245 , n40246 , n40247 , n40248 , n40249 , n40250 , n40251 , n40252 , n40253 , n40254 , n40255 , n40256 , n40257 , n40258 , n40259 , n40260 , n40261 , n40262 , n40263 , n40264 , n40265 , n40266 , n40267 , n40268 , n40269 , n40270 , n40271 , n40272 , n40273 , n40274 , n40275 , n40276 , n40277 , n40278 , n40279 , n40280 , n40281 , n40282 , n40283 , n40284 , n40285 , n40286 , n40287 , n40288 , n40289 , n40290 , n40291 , n40292 , n40293 , n40294 , n40295 , n40296 , n40297 , n40298 , n40299 , n40300 , n40301 , n40302 , n40303 , n40304 , n40305 , n40306 , n40307 , n40308 , n40309 , n40310 , n40311 , n40312 , n40313 , n40314 , n40315 , n40316 , n40317 , n40318 , n40319 , n40320 , n40321 , n40322 , n40323 , n40324 , n40325 , n40326 , n40327 , n40328 , n40329 , n40330 , n40331 , n40332 , n40333 , n40334 , n40335 , n40336 , n40337 , n40338 , n40339 , n40340 , n40341 , n40342 , n40343 , n40344 , n40345 , n40346 , n40347 , n40348 , n40349 , n40350 , n40351 , n40352 , n40353 , n40354 , n40355 , n40356 , n40357 , n40358 , n40359 , n40360 , n40361 , n40362 , n40363 , n40364 , n40365 , n40366 , n40367 , n40368 , n40369 , n40370 , n40371 , n40372 , n40373 , n40374 , n40375 , n40376 , n40377 , n40378 , n40379 , n40380 , n40381 , n40382 , n40383 , n40384 , n40385 , n40386 , n40387 , n40388 , n40389 , n40390 , n40391 , n40392 , n40393 , n40394 , n40395 , n40396 , n40397 , n40398 , n40399 , n40400 , n40401 , n40402 , n40403 , n40404 , n40405 , n40406 , n40407 , n40408 , n40409 , n40410 , n40411 , n40412 , n40413 , n40414 , n40415 , n40416 , n40417 , n40418 , n40419 , n40420 , n40421 , n40422 , n40423 , n40424 , n40425 , n40426 , n40427 , n40428 , n40429 , n40430 , n40431 , n40432 , n40433 , n40434 , n40435 , n40436 , n40437 , n40438 , n40439 , n40440 , n40441 , n40442 , n40443 , n40444 , n40445 , n40446 , n40447 , n40448 , n40449 , n40450 , n40451 , n40452 , n40453 , n40454 , n40455 , n40456 , n40457 , n40458 , n40459 , n40460 , n40461 , n40462 , n40463 , n40464 , n40465 , n40466 , n40467 , n40468 , n40469 , n40470 , n40471 , n40472 , n40473 , n40474 , n40475 , n40476 , n40477 , n40478 , n40479 , n40480 , n40481 , n40482 , n40483 , n40484 , n40485 , n40486 , n40487 , n40488 , n40489 , n40490 , n40491 , n40492 , n40493 , n40494 , n40495 , n40496 , n40497 , n40498 , n40499 , n40500 , n40501 , n40502 , n40503 , n40504 , n40505 , n40506 , n40507 , n40508 , n40509 , n40510 , n40511 , n40512 , n40513 , n40514 , n40515 , n40516 , n40517 , n40518 , n40519 , n40520 , n40521 , n40522 , n40523 , n40524 , n40525 , n40526 , n40527 , n40528 , n40529 , n40530 , n40531 , n40532 , n40533 , n40534 , n40535 , n40536 , n40537 , n40538 , n40539 , n40540 , n40541 , n40542 , n40543 , n40544 , n40545 , n40546 , n40547 , n40548 , n40549 , n40550 , n40551 , n40552 , n40553 , n40554 , n40555 , n40556 , n40557 , n40558 , n40559 , n40560 , n40561 , n40562 , n40563 , n40564 , n40565 , n40566 , n40567 , n40568 , n40569 , n40570 , n40571 , n40572 , n40573 , n40574 , n40575 , n40576 , n40577 , n40578 , n40579 , n40580 , n40581 , n40582 , n40583 , n40584 , n40585 , n40586 , n40587 , n40588 , n40589 , n40590 , n40591 , n40592 , n40593 , n40594 , n40595 , n40596 , n40597 , n40598 , n40599 , n40600 , n40601 , n40602 , n40603 , n40604 , n40605 , n40606 , n40607 , n40608 , n40609 , n40610 , n40611 , n40612 , n40613 , n40614 , n40615 , n40616 , n40617 , n40618 , n40619 , n40620 , n40621 , n40622 , n40623 , n40624 , n40625 , n40626 , n40627 , n40628 , n40629 , n40630 , n40631 , n40632 , n40633 , n40634 , n40635 , n40636 , n40637 , n40638 , n40639 , n40640 , n40641 , n40642 , n40643 , n40644 , n40645 , n40646 , n40647 , n40648 , n40649 , n40650 , n40651 , n40652 , n40653 , n40654 , n40655 , n40656 , n40657 , n40658 , n40659 , n40660 , n40661 , n40662 , n40663 , n40664 , n40665 , n40666 , n40667 , n40668 , n40669 , n40670 , n40671 , n40672 , n40673 , n40674 , n40675 , n40676 , n40677 , n40678 , n40679 , n40680 , n40681 , n40682 , n40683 , n40684 , n40685 , n40686 , n40687 , n40688 , n40689 , n40690 , n40691 , n40692 , n40693 , n40694 , n40695 , n40696 , n40697 , n40698 , n40699 , n40700 , n40701 , n40702 , n40703 , n40704 , n40705 , n40706 , n40707 , n40708 , n40709 , n40710 , n40711 , n40712 , n40713 , n40714 , n40715 , n40716 , n40717 , n40718 , n40719 , n40720 , n40721 , n40722 , n40723 , n40724 , n40725 , n40726 , n40727 , n40728 , n40729 , n40730 , n40731 , n40732 , n40733 , n40734 , n40735 , n40736 , n40737 , n40738 , n40739 , n40740 , n40741 , n40742 , n40743 , n40744 , n40745 , n40746 , n40747 , n40748 , n40749 , n40750 , n40751 , n40752 , n40753 , n40754 , n40755 , n40756 , n40757 , n40758 , n40759 , n40760 , n40761 , n40762 , n40763 , n40764 , n40765 , n40766 , n40767 , n40768 , n40769 , n40770 , n40771 , n40772 , n40773 , n40774 , n40775 , n40776 , n40777 , n40778 , n40779 , n40780 , n40781 , n40782 , n40783 , n40784 , n40785 , n40786 , n40787 , n40788 , n40789 , n40790 , n40791 , n40792 , n40793 , n40794 , n40795 , n40796 , n40797 , n40798 , n40799 , n40800 , n40801 , n40802 , n40803 , n40804 , n40805 , n40806 , n40807 , n40808 , n40809 , n40810 , n40811 , n40812 , n40813 , n40814 , n40815 , n40816 , n40817 , n40818 , n40819 , n40820 , n40821 , n40822 , n40823 , n40824 , n40825 , n40826 , n40827 , n40828 , n40829 , n40830 , n40831 , n40832 , n40833 , n40834 , n40835 , n40836 , n40837 , n40838 , n40839 , n40840 , n40841 , n40842 , n40843 , n40844 , n40845 , n40846 , n40847 , n40848 , n40849 , n40850 , n40851 , n40852 , n40853 , n40854 , n40855 , n40856 , n40857 , n40858 , n40859 , n40860 , n40861 , n40862 , n40863 , n40864 , n40865 , n40866 , n40867 , n40868 , n40869 , n40870 , n40871 , n40872 , n40873 , n40874 , n40875 , n40876 , n40877 , n40878 , n40879 , n40880 , n40881 , n40882 , n40883 , n40884 , n40885 , n40886 , n40887 , n40888 , n40889 , n40890 , n40891 , n40892 , n40893 , n40894 , n40895 , n40896 , n40897 , n40898 , n40899 , n40900 , n40901 , n40902 , n40903 , n40904 , n40905 , n40906 , n40907 , n40908 , n40909 , n40910 , n40911 , n40912 , n40913 , n40914 , n40915 , n40916 , n40917 , n40918 , n40919 , n40920 , n40921 , n40922 , n40923 , n40924 , n40925 , n40926 , n40927 , n40928 , n40929 , n40930 , n40931 , n40932 , n40933 , n40934 , n40935 , n40936 , n40937 , n40938 , n40939 , n40940 , n40941 , n40942 , n40943 , n40944 , n40945 , n40946 , n40947 , n40948 , n40949 , n40950 , n40951 , n40952 , n40953 , n40954 , n40955 , n40956 , n40957 , n40958 , n40959 , n40960 , n40961 , n40962 , n40963 , n40964 , n40965 , n40966 , n40967 , n40968 , n40969 , n40970 , n40971 , n40972 , n40973 , n40974 , n40975 , n40976 , n40977 , n40978 , n40979 , n40980 , n40981 , n40982 , n40983 , n40984 , n40985 , n40986 , n40987 , n40988 , n40989 , n40990 , n40991 , n40992 , n40993 , n40994 , n40995 , n40996 , n40997 , n40998 , n40999 , n41000 , n41001 , n41002 , n41003 , n41004 , n41005 , n41006 , n41007 , n41008 , n41009 , n41010 , n41011 , n41012 , n41013 , n41014 , n41015 , n41016 , n41017 , n41018 , n41019 , n41020 , n41021 , n41022 , n41023 , n41024 , n41025 , n41026 , n41027 , n41028 , n41029 , n41030 , n41031 , n41032 , n41033 , n41034 , n41035 , n41036 , n41037 , n41038 , n41039 , n41040 , n41041 , n41042 , n41043 , n41044 , n41045 , n41046 , n41047 , n41048 , n41049 , n41050 , n41051 , n41052 , n41053 , n41054 , n41055 , n41056 , n41057 , n41058 , n41059 , n41060 , n41061 , n41062 , n41063 , n41064 , n41065 , n41066 , n41067 , n41068 , n41069 , n41070 , n41071 , n41072 , n41073 , n41074 , n41075 , n41076 , n41077 , n41078 , n41079 , n41080 , n41081 , n41082 , n41083 , n41084 , n41085 , n41086 , n41087 , n41088 , n41089 , n41090 , n41091 , n41092 , n41093 , n41094 , n41095 , n41096 , n41097 , n41098 , n41099 , n41100 , n41101 , n41102 , n41103 , n41104 , n41105 , n41106 , n41107 , n41108 , n41109 , n41110 , n41111 , n41112 , n41113 , n41114 , n41115 , n41116 , n41117 , n41118 , n41119 , n41120 , n41121 , n41122 , n41123 , n41124 , n41125 , n41126 , n41127 , n41128 , n41129 , n41130 , n41131 , n41132 , n41133 , n41134 , n41135 , n41136 , n41137 , n41138 , n41139 , n41140 , n41141 , n41142 , n41143 , n41144 , n41145 , n41146 , n41147 , n41148 , n41149 , n41150 , n41151 , n41152 , n41153 , n41154 , n41155 , n41156 , n41157 , n41158 , n41159 , n41160 , n41161 , n41162 , n41163 , n41164 , n41165 , n41166 , n41167 , n41168 , n41169 , n41170 , n41171 , n41172 , n41173 , n41174 , n41175 , n41176 , n41177 , n41178 , n41179 , n41180 , n41181 , n41182 , n41183 , n41184 , n41185 , n41186 , n41187 , n41188 , n41189 , n41190 , n41191 , n41192 , n41193 , n41194 , n41195 , n41196 , n41197 , n41198 , n41199 , n41200 , n41201 , n41202 , n41203 , n41204 , n41205 , n41206 , n41207 , n41208 , n41209 , n41210 , n41211 , n41212 , n41213 , n41214 , n41215 , n41216 , n41217 , n41218 , n41219 , n41220 , n41221 , n41222 , n41223 , n41224 , n41225 , n41226 , n41227 , n41228 , n41229 , n41230 , n41231 , n41232 , n41233 , n41234 , n41235 , n41236 , n41237 , n41238 , n41239 , n41240 , n41241 , n41242 , n41243 , n41244 , n41245 , n41246 , n41247 , n41248 , n41249 , n41250 , n41251 , n41252 , n41253 , n41254 , n41255 , n41256 , n41257 , n41258 , n41259 , n41260 , n41261 , n41262 , n41263 , n41264 , n41265 , n41266 , n41267 , n41268 , n41269 , n41270 , n41271 , n41272 , n41273 , n41274 , n41275 , n41276 , n41277 , n41278 , n41279 , n41280 , n41281 , n41282 , n41283 , n41284 , n41285 , n41286 , n41287 , n41288 , n41289 , n41290 , n41291 , n41292 , n41293 , n41294 , n41295 , n41296 , n41297 , n41298 , n41299 , n41300 , n41301 , n41302 , n41303 , n41304 , n41305 , n41306 , n41307 , n41308 , n41309 , n41310 , n41311 , n41312 , n41313 , n41314 , n41315 , n41316 , n41317 , n41318 , n41319 , n41320 , n41321 , n41322 , n41323 , n41324 , n41325 , n41326 , n41327 , n41328 , n41329 , n41330 , n41331 , n41332 , n41333 , n41334 , n41335 , n41336 , n41337 , n41338 , n41339 , n41340 , n41341 , n41342 , n41343 , n41344 , n41345 , n41346 , n41347 , n41348 , n41349 , n41350 , n41351 , n41352 , n41353 , n41354 , n41355 , n41356 , n41357 , n41358 , n41359 , n41360 , n41361 , n41362 , n41363 , n41364 , n41365 , n41366 , n41367 , n41368 , n41369 , n41370 , n41371 , n41372 , n41373 , n41374 , n41375 , n41376 , n41377 , n41378 , n41379 , n41380 , n41381 , n41382 , n41383 , n41384 , n41385 , n41386 , n41387 , n41388 , n41389 , n41390 , n41391 , n41392 , n41393 , n41394 , n41395 , n41396 , n41397 , n41398 , n41399 , n41400 , n41401 , n41402 , n41403 , n41404 , n41405 , n41406 , n41407 , n41408 , n41409 , n41410 , n41411 , n41412 , n41413 , n41414 , n41415 , n41416 , n41417 , n41418 , n41419 , n41420 , n41421 , n41422 , n41423 , n41424 , n41425 , n41426 , n41427 , n41428 , n41429 , n41430 , n41431 , n41432 , n41433 , n41434 , n41435 , n41436 , n41437 , n41438 , n41439 , n41440 , n41441 , n41442 , n41443 , n41444 , n41445 , n41446 , n41447 , n41448 , n41449 , n41450 , n41451 , n41452 , n41453 , n41454 , n41455 , n41456 , n41457 , n41458 , n41459 , n41460 , n41461 , n41462 , n41463 , n41464 , n41465 , n41466 , n41467 , n41468 , n41469 , n41470 , n41471 , n41472 , n41473 , n41474 , n41475 , n41476 , n41477 , n41478 , n41479 , n41480 , n41481 , n41482 , n41483 , n41484 , n41485 , n41486 , n41487 , n41488 , n41489 , n41490 , n41491 , n41492 , n41493 , n41494 , n41495 , n41496 , n41497 , n41498 , n41499 , n41500 , n41501 , n41502 , n41503 , n41504 , n41505 , n41506 , n41507 , n41508 , n41509 , n41510 , n41511 , n41512 , n41513 , n41514 , n41515 , n41516 , n41517 , n41518 , n41519 , n41520 , n41521 , n41522 , n41523 , n41524 , n41525 , n41526 , n41527 , n41528 , n41529 , n41530 , n41531 , n41532 , n41533 , n41534 , n41535 , n41536 , n41537 , n41538 , n41539 , n41540 , n41541 , n41542 , n41543 , n41544 , n41545 , n41546 , n41547 , n41548 , n41549 , n41550 , n41551 , n41552 , n41553 , n41554 , n41555 , n41556 , n41557 , n41558 , n41559 , n41560 , n41561 , n41562 , n41563 , n41564 , n41565 , n41566 , n41567 , n41568 , n41569 , n41570 , n41571 , n41572 , n41573 , n41574 , n41575 , n41576 , n41577 , n41578 , n41579 , n41580 , n41581 , n41582 , n41583 , n41584 , n41585 , n41586 , n41587 , n41588 , n41589 , n41590 , n41591 , n41592 , n41593 , n41594 , n41595 , n41596 , n41597 , n41598 , n41599 , n41600 , n41601 , n41602 , n41603 , n41604 , n41605 , n41606 , n41607 , n41608 , n41609 , n41610 , n41611 , n41612 , n41613 , n41614 , n41615 , n41616 , n41617 , n41618 , n41619 , n41620 , n41621 , n41622 , n41623 , n41624 , n41625 , n41626 , n41627 , n41628 , n41629 , n41630 , n41631 , n41632 , n41633 , n41634 , n41635 , n41636 , n41637 , n41638 , n41639 , n41640 , n41641 , n41642 , n41643 , n41644 , n41645 , n41646 , n41647 , n41648 , n41649 , n41650 , n41651 , n41652 , n41653 , n41654 , n41655 , n41656 , n41657 , n41658 , n41659 , n41660 , n41661 , n41662 , n41663 , n41664 , n41665 , n41666 , n41667 , n41668 , n41669 , n41670 , n41671 , n41672 , n41673 , n41674 , n41675 , n41676 , n41677 , n41678 , n41679 , n41680 , n41681 , n41682 , n41683 , n41684 , n41685 , n41686 , n41687 , n41688 , n41689 , n41690 , n41691 , n41692 , n41693 , n41694 , n41695 , n41696 , n41697 , n41698 , n41699 , n41700 , n41701 , n41702 , n41703 , n41704 , n41705 , n41706 , n41707 , n41708 , n41709 , n41710 , n41711 , n41712 , n41713 , n41714 , n41715 , n41716 , n41717 , n41718 , n41719 , n41720 , n41721 , n41722 , n41723 , n41724 , n41725 , n41726 , n41727 , n41728 , n41729 , n41730 , n41731 , n41732 , n41733 , n41734 , n41735 , n41736 , n41737 , n41738 , n41739 , n41740 , n41741 , n41742 , n41743 , n41744 , n41745 , n41746 , n41747 , n41748 , n41749 , n41750 , n41751 , n41752 , n41753 , n41754 , n41755 , n41756 , n41757 , n41758 , n41759 , n41760 , n41761 , n41762 , n41763 , n41764 , n41765 , n41766 , n41767 , n41768 , n41769 , n41770 , n41771 , n41772 , n41773 , n41774 , n41775 , n41776 , n41777 , n41778 , n41779 , n41780 , n41781 , n41782 , n41783 , n41784 , n41785 , n41786 , n41787 , n41788 , n41789 , n41790 , n41791 , n41792 , n41793 , n41794 , n41795 , n41796 , n41797 , n41798 , n41799 , n41800 , n41801 , n41802 , n41803 , n41804 , n41805 , n41806 , n41807 , n41808 , n41809 , n41810 , n41811 , n41812 , n41813 , n41814 , n41815 , n41816 , n41817 , n41818 , n41819 , n41820 , n41821 , n41822 , n41823 , n41824 , n41825 , n41826 , n41827 , n41828 , n41829 , n41830 , n41831 , n41832 , n41833 , n41834 , n41835 , n41836 , n41837 , n41838 , n41839 , n41840 , n41841 , n41842 , n41843 , n41844 , n41845 , n41846 , n41847 , n41848 , n41849 , n41850 , n41851 , n41852 , n41853 , n41854 , n41855 , n41856 , n41857 , n41858 , n41859 , n41860 , n41861 , n41862 , n41863 , n41864 , n41865 , n41866 , n41867 , n41868 , n41869 , n41870 , n41871 , n41872 , n41873 , n41874 , n41875 , n41876 , n41877 , n41878 , n41879 , n41880 , n41881 , n41882 , n41883 , n41884 , n41885 , n41886 , n41887 , n41888 , n41889 , n41890 , n41891 , n41892 , n41893 , n41894 , n41895 , n41896 , n41897 , n41898 , n41899 , n41900 , n41901 , n41902 , n41903 , n41904 , n41905 , n41906 , n41907 , n41908 , n41909 , n41910 , n41911 , n41912 , n41913 , n41914 , n41915 , n41916 , n41917 , n41918 , n41919 , n41920 , n41921 , n41922 , n41923 , n41924 , n41925 , n41926 , n41927 , n41928 , n41929 , n41930 , n41931 , n41932 , n41933 , n41934 , n41935 , n41936 , n41937 , n41938 , n41939 , n41940 , n41941 , n41942 , n41943 , n41944 , n41945 , n41946 , n41947 , n41948 , n41949 , n41950 , n41951 , n41952 , n41953 , n41954 , n41955 , n41956 , n41957 , n41958 , n41959 , n41960 , n41961 , n41962 , n41963 , n41964 , n41965 , n41966 , n41967 , n41968 , n41969 , n41970 , n41971 , n41972 , n41973 , n41974 , n41975 , n41976 , n41977 , n41978 , n41979 , n41980 , n41981 , n41982 , n41983 , n41984 , n41985 , n41986 , n41987 , n41988 , n41989 , n41990 , n41991 , n41992 , n41993 , n41994 , n41995 , n41996 , n41997 , n41998 , n41999 , n42000 , n42001 , n42002 , n42003 , n42004 , n42005 , n42006 , n42007 , n42008 , n42009 , n42010 , n42011 , n42012 , n42013 , n42014 , n42015 , n42016 , n42017 , n42018 , n42019 , n42020 , n42021 , n42022 , n42023 , n42024 , n42025 , n42026 , n42027 , n42028 , n42029 , n42030 , n42031 , n42032 , n42033 , n42034 , n42035 , n42036 , n42037 , n42038 , n42039 , n42040 , n42041 , n42042 , n42043 , n42044 , n42045 , n42046 , n42047 , n42048 , n42049 , n42050 , n42051 , n42052 , n42053 , n42054 , n42055 , n42056 , n42057 , n42058 , n42059 , n42060 , n42061 , n42062 , n42063 , n42064 , n42065 , n42066 , n42067 , n42068 , n42069 , n42070 , n42071 , n42072 , n42073 , n42074 , n42075 , n42076 , n42077 , n42078 , n42079 , n42080 , n42081 , n42082 , n42083 , n42084 , n42085 , n42086 , n42087 , n42088 , n42089 , n42090 , n42091 , n42092 , n42093 , n42094 , n42095 , n42096 , n42097 , n42098 , n42099 , n42100 , n42101 , n42102 , n42103 , n42104 , n42105 , n42106 , n42107 , n42108 , n42109 , n42110 , n42111 , n42112 , n42113 , n42114 , n42115 , n42116 , n42117 , n42118 , n42119 , n42120 , n42121 , n42122 , n42123 , n42124 , n42125 , n42126 , n42127 , n42128 , n42129 , n42130 , n42131 , n42132 , n42133 , n42134 , n42135 , n42136 , n42137 , n42138 , n42139 , n42140 , n42141 , n42142 , n42143 , n42144 , n42145 , n42146 , n42147 , n42148 , n42149 , n42150 , n42151 , n42152 , n42153 , n42154 , n42155 , n42156 , n42157 , n42158 , n42159 , n42160 , n42161 , n42162 , n42163 , n42164 , n42165 , n42166 , n42167 , n42168 , n42169 , n42170 , n42171 , n42172 , n42173 , n42174 , n42175 , n42176 , n42177 , n42178 , n42179 , n42180 , n42181 , n42182 , n42183 , n42184 , n42185 , n42186 , n42187 , n42188 , n42189 , n42190 , n42191 , n42192 , n42193 , n42194 , n42195 , n42196 , n42197 , n42198 , n42199 , n42200 , n42201 , n42202 , n42203 , n42204 , n42205 , n42206 , n42207 , n42208 , n42209 , n42210 , n42211 , n42212 , n42213 , n42214 , n42215 , n42216 , n42217 , n42218 , n42219 , n42220 , n42221 , n42222 , n42223 , n42224 , n42225 , n42226 , n42227 , n42228 , n42229 , n42230 , n42231 , n42232 , n42233 , n42234 , n42235 , n42236 , n42237 , n42238 , n42239 , n42240 , n42241 , n42242 , n42243 , n42244 , n42245 , n42246 , n42247 , n42248 , n42249 , n42250 , n42251 , n42252 , n42253 , n42254 , n42255 , n42256 , n42257 , n42258 , n42259 , n42260 , n42261 , n42262 , n42263 , n42264 , n42265 , n42266 , n42267 , n42268 , n42269 , n42270 , n42271 , n42272 , n42273 , n42274 , n42275 , n42276 , n42277 , n42278 , n42279 , n42280 , n42281 , n42282 , n42283 , n42284 , n42285 , n42286 , n42287 , n42288 , n42289 , n42290 , n42291 , n42292 , n42293 , n42294 , n42295 , n42296 , n42297 , n42298 , n42299 , n42300 , n42301 , n42302 , n42303 , n42304 , n42305 , n42306 , n42307 , n42308 , n42309 , n42310 , n42311 , n42312 , n42313 , n42314 , n42315 , n42316 , n42317 , n42318 , n42319 , n42320 , n42321 , n42322 , n42323 , n42324 , n42325 , n42326 , n42327 , n42328 , n42329 , n42330 , n42331 , n42332 , n42333 , n42334 , n42335 , n42336 , n42337 , n42338 , n42339 , n42340 , n42341 , n42342 , n42343 , n42344 , n42345 , n42346 , n42347 , n42348 , n42349 , n42350 , n42351 , n42352 , n42353 , n42354 , n42355 , n42356 , n42357 , n42358 , n42359 , n42360 , n42361 , n42362 , n42363 , n42364 , n42365 , n42366 , n42367 , n42368 , n42369 , n42370 , n42371 , n42372 , n42373 , n42374 , n42375 , n42376 , n42377 , n42378 , n42379 , n42380 , n42381 , n42382 , n42383 , n42384 , n42385 , n42386 , n42387 , n42388 , n42389 , n42390 , n42391 , n42392 , n42393 , n42394 , n42395 , n42396 , n42397 , n42398 , n42399 , n42400 , n42401 , n42402 , n42403 , n42404 , n42405 , n42406 , n42407 , n42408 , n42409 , n42410 , n42411 , n42412 , n42413 , n42414 , n42415 , n42416 , n42417 , n42418 , n42419 , n42420 , n42421 , n42422 , n42423 , n42424 , n42425 , n42426 , n42427 , n42428 , n42429 , n42430 , n42431 , n42432 , n42433 , n42434 , n42435 , n42436 , n42437 , n42438 , n42439 , n42440 , n42441 , n42442 , n42443 , n42444 , n42445 , n42446 , n42447 , n42448 , n42449 , n42450 , n42451 , n42452 , n42453 , n42454 , n42455 , n42456 , n42457 , n42458 , n42459 , n42460 , n42461 , n42462 , n42463 , n42464 , n42465 , n42466 , n42467 , n42468 , n42469 , n42470 , n42471 , n42472 , n42473 , n42474 , n42475 , n42476 , n42477 , n42478 , n42479 , n42480 , n42481 , n42482 , n42483 , n42484 , n42485 , n42486 , n42487 , n42488 , n42489 , n42490 , n42491 , n42492 , n42493 , n42494 , n42495 , n42496 , n42497 , n42498 , n42499 , n42500 , n42501 , n42502 , n42503 , n42504 , n42505 , n42506 , n42507 , n42508 , n42509 , n42510 , n42511 , n42512 , n42513 , n42514 , n42515 , n42516 , n42517 , n42518 , n42519 , n42520 , n42521 , n42522 , n42523 , n42524 , n42525 , n42526 , n42527 , n42528 , n42529 , n42530 , n42531 , n42532 , n42533 , n42534 , n42535 , n42536 , n42537 , n42538 , n42539 , n42540 , n42541 , n42542 , n42543 , n42544 , n42545 , n42546 , n42547 , n42548 , n42549 , n42550 , n42551 , n42552 , n42553 , n42554 , n42555 , n42556 , n42557 , n42558 , n42559 , n42560 , n42561 , n42562 , n42563 , n42564 , n42565 , n42566 , n42567 , n42568 , n42569 , n42570 , n42571 , n42572 , n42573 , n42574 , n42575 , n42576 , n42577 , n42578 , n42579 , n42580 , n42581 , n42582 , n42583 , n42584 , n42585 , n42586 , n42587 , n42588 , n42589 , n42590 , n42591 , n42592 , n42593 , n42594 , n42595 , n42596 , n42597 , n42598 , n42599 , n42600 , n42601 , n42602 , n42603 , n42604 , n42605 , n42606 , n42607 , n42608 , n42609 , n42610 , n42611 , n42612 , n42613 , n42614 , n42615 , n42616 , n42617 , n42618 , n42619 , n42620 , n42621 , n42622 , n42623 , n42624 , n42625 , n42626 , n42627 , n42628 , n42629 , n42630 , n42631 , n42632 , n42633 , n42634 , n42635 , n42636 , n42637 , n42638 , n42639 , n42640 , n42641 , n42642 , n42643 , n42644 , n42645 , n42646 , n42647 , n42648 , n42649 , n42650 , n42651 , n42652 , n42653 , n42654 , n42655 , n42656 , n42657 , n42658 , n42659 , n42660 , n42661 , n42662 , n42663 , n42664 , n42665 , n42666 , n42667 , n42668 , n42669 , n42670 , n42671 , n42672 , n42673 , n42674 , n42675 , n42676 , n42677 , n42678 , n42679 , n42680 , n42681 , n42682 , n42683 , n42684 , n42685 , n42686 , n42687 , n42688 , n42689 , n42690 , n42691 , n42692 , n42693 , n42694 , n42695 , n42696 , n42697 , n42698 , n42699 , n42700 , n42701 , n42702 , n42703 , n42704 , n42705 , n42706 , n42707 , n42708 , n42709 , n42710 , n42711 , n42712 , n42713 , n42714 , n42715 , n42716 , n42717 , n42718 , n42719 , n42720 , n42721 , n42722 , n42723 , n42724 , n42725 , n42726 , n42727 , n42728 , n42729 , n42730 , n42731 , n42732 , n42733 , n42734 , n42735 , n42736 , n42737 , n42738 , n42739 , n42740 , n42741 , n42742 , n42743 , n42744 , n42745 , n42746 , n42747 , n42748 , n42749 , n42750 , n42751 , n42752 , n42753 , n42754 , n42755 , n42756 , n42757 , n42758 , n42759 , n42760 , n42761 , n42762 , n42763 , n42764 , n42765 , n42766 , n42767 , n42768 , n42769 , n42770 , n42771 , n42772 , n42773 , n42774 , n42775 , n42776 , n42777 , n42778 , n42779 , n42780 , n42781 , n42782 , n42783 , n42784 , n42785 , n42786 , n42787 , n42788 , n42789 , n42790 , n42791 , n42792 , n42793 , n42794 , n42795 , n42796 , n42797 , n42798 , n42799 , n42800 , n42801 , n42802 , n42803 , n42804 , n42805 , n42806 , n42807 , n42808 , n42809 , n42810 , n42811 , n42812 , n42813 , n42814 , n42815 , n42816 , n42817 , n42818 , n42819 , n42820 , n42821 , n42822 , n42823 , n42824 , n42825 , n42826 , n42827 , n42828 , n42829 , n42830 , n42831 , n42832 , n42833 , n42834 , n42835 , n42836 , n42837 , n42838 , n42839 , n42840 , n42841 , n42842 , n42843 , n42844 , n42845 , n42846 , n42847 , n42848 , n42849 , n42850 , n42851 , n42852 , n42853 , n42854 , n42855 , n42856 , n42857 , n42858 , n42859 , n42860 , n42861 , n42862 , n42863 , n42864 , n42865 , n42866 , n42867 , n42868 , n42869 , n42870 , n42871 , n42872 , n42873 , n42874 , n42875 , n42876 , n42877 , n42878 , n42879 , n42880 , n42881 , n42882 , n42883 , n42884 , n42885 , n42886 , n42887 , n42888 , n42889 , n42890 , n42891 , n42892 , n42893 , n42894 , n42895 , n42896 , n42897 , n42898 , n42899 , n42900 , n42901 , n42902 , n42903 , n42904 , n42905 , n42906 , n42907 , n42908 , n42909 , n42910 , n42911 , n42912 , n42913 , n42914 , n42915 , n42916 , n42917 , n42918 , n42919 , n42920 , n42921 , n42922 , n42923 , n42924 , n42925 , n42926 , n42927 , n42928 , n42929 , n42930 , n42931 , n42932 , n42933 , n42934 , n42935 , n42936 , n42937 , n42938 , n42939 , n42940 , n42941 , n42942 , n42943 , n42944 , n42945 , n42946 , n42947 , n42948 , n42949 , n42950 , n42951 , n42952 , n42953 , n42954 , n42955 , n42956 , n42957 , n42958 , n42959 , n42960 , n42961 , n42962 , n42963 , n42964 , n42965 , n42966 , n42967 , n42968 , n42969 , n42970 , n42971 , n42972 , n42973 , n42974 , n42975 , n42976 , n42977 , n42978 , n42979 , n42980 , n42981 , n42982 , n42983 , n42984 , n42985 , n42986 , n42987 , n42988 , n42989 , n42990 , n42991 , n42992 , n42993 , n42994 , n42995 , n42996 , n42997 , n42998 , n42999 , n43000 , n43001 , n43002 , n43003 , n43004 , n43005 , n43006 , n43007 , n43008 , n43009 , n43010 , n43011 , n43012 , n43013 , n43014 , n43015 , n43016 , n43017 , n43018 , n43019 , n43020 , n43021 , n43022 , n43023 , n43024 , n43025 , n43026 , n43027 , n43028 , n43029 , n43030 , n43031 , n43032 , n43033 , n43034 , n43035 , n43036 , n43037 , n43038 , n43039 , n43040 , n43041 , n43042 , n43043 , n43044 , n43045 , n43046 , n43047 , n43048 , n43049 , n43050 , n43051 , n43052 , n43053 , n43054 , n43055 , n43056 , n43057 , n43058 , n43059 , n43060 , n43061 , n43062 , n43063 , n43064 , n43065 , n43066 , n43067 , n43068 , n43069 , n43070 , n43071 , n43072 , n43073 , n43074 , n43075 , n43076 , n43077 , n43078 , n43079 , n43080 , n43081 , n43082 , n43083 , n43084 , n43085 , n43086 , n43087 , n43088 , n43089 , n43090 , n43091 , n43092 , n43093 , n43094 , n43095 , n43096 , n43097 , n43098 , n43099 , n43100 , n43101 , n43102 , n43103 , n43104 , n43105 , n43106 , n43107 , n43108 , n43109 , n43110 , n43111 , n43112 , n43113 , n43114 , n43115 , n43116 , n43117 , n43118 , n43119 , n43120 , n43121 , n43122 , n43123 , n43124 , n43125 , n43126 , n43127 , n43128 , n43129 , n43130 , n43131 , n43132 , n43133 , n43134 , n43135 , n43136 , n43137 , n43138 , n43139 , n43140 , n43141 , n43142 , n43143 , n43144 , n43145 , n43146 , n43147 , n43148 , n43149 , n43150 , n43151 , n43152 , n43153 , n43154 , n43155 , n43156 , n43157 , n43158 , n43159 , n43160 , n43161 , n43162 , n43163 , n43164 , n43165 , n43166 , n43167 , n43168 , n43169 , n43170 , n43171 , n43172 , n43173 , n43174 , n43175 , n43176 , n43177 , n43178 , n43179 , n43180 , n43181 , n43182 , n43183 , n43184 , n43185 , n43186 , n43187 , n43188 , n43189 , n43190 , n43191 , n43192 , n43193 , n43194 , n43195 , n43196 , n43197 , n43198 , n43199 , n43200 , n43201 , n43202 , n43203 , n43204 , n43205 , n43206 , n43207 , n43208 , n43209 , n43210 , n43211 , n43212 , n43213 , n43214 , n43215 , n43216 , n43217 , n43218 , n43219 , n43220 , n43221 , n43222 , n43223 , n43224 , n43225 , n43226 , n43227 , n43228 , n43229 , n43230 , n43231 , n43232 , n43233 , n43234 , n43235 , n43236 , n43237 , n43238 , n43239 , n43240 , n43241 , n43242 , n43243 , n43244 , n43245 , n43246 , n43247 , n43248 , n43249 , n43250 , n43251 , n43252 , n43253 , n43254 , n43255 , n43256 , n43257 , n43258 , n43259 , n43260 , n43261 , n43262 , n43263 , n43264 , n43265 , n43266 , n43267 , n43268 , n43269 , n43270 , n43271 , n43272 , n43273 , n43274 , n43275 , n43276 , n43277 , n43278 , n43279 , n43280 , n43281 , n43282 , n43283 , n43284 , n43285 , n43286 , n43287 , n43288 , n43289 , n43290 , n43291 , n43292 , n43293 , n43294 , n43295 , n43296 , n43297 , n43298 , n43299 , n43300 , n43301 , n43302 , n43303 , n43304 , n43305 , n43306 , n43307 , n43308 , n43309 , n43310 , n43311 , n43312 , n43313 , n43314 , n43315 , n43316 , n43317 , n43318 , n43319 , n43320 , n43321 , n43322 , n43323 , n43324 , n43325 , n43326 , n43327 , n43328 , n43329 , n43330 , n43331 , n43332 , n43333 , n43334 , n43335 , n43336 , n43337 , n43338 , n43339 , n43340 , n43341 , n43342 , n43343 , n43344 , n43345 , n43346 , n43347 , n43348 , n43349 , n43350 , n43351 , n43352 , n43353 , n43354 , n43355 , n43356 , n43357 , n43358 , n43359 , n43360 , n43361 , n43362 , n43363 , n43364 , n43365 , n43366 , n43367 , n43368 , n43369 , n43370 , n43371 , n43372 , n43373 , n43374 , n43375 , n43376 , n43377 , n43378 , n43379 , n43380 , n43381 , n43382 , n43383 , n43384 , n43385 , n43386 , n43387 , n43388 , n43389 , n43390 , n43391 , n43392 , n43393 , n43394 , n43395 , n43396 , n43397 , n43398 , n43399 , n43400 , n43401 , n43402 , n43403 , n43404 , n43405 , n43406 , n43407 , n43408 , n43409 , n43410 , n43411 , n43412 , n43413 , n43414 , n43415 , n43416 , n43417 , n43418 , n43419 , n43420 , n43421 , n43422 , n43423 , n43424 , n43425 , n43426 , n43427 , n43428 , n43429 , n43430 , n43431 , n43432 , n43433 , n43434 , n43435 , n43436 , n43437 , n43438 , n43439 , n43440 , n43441 , n43442 , n43443 , n43444 , n43445 , n43446 , n43447 , n43448 , n43449 , n43450 , n43451 , n43452 , n43453 , n43454 , n43455 , n43456 , n43457 , n43458 , n43459 , n43460 , n43461 , n43462 , n43463 , n43464 , n43465 , n43466 , n43467 , n43468 , n43469 , n43470 , n43471 , n43472 , n43473 , n43474 , n43475 , n43476 , n43477 , n43478 , n43479 , n43480 , n43481 , n43482 , n43483 , n43484 , n43485 , n43486 , n43487 , n43488 , n43489 , n43490 , n43491 , n43492 , n43493 , n43494 , n43495 , n43496 , n43497 , n43498 , n43499 , n43500 , n43501 , n43502 , n43503 , n43504 , n43505 , n43506 , n43507 , n43508 , n43509 , n43510 , n43511 , n43512 , n43513 , n43514 , n43515 , n43516 , n43517 , n43518 , n43519 , n43520 , n43521 , n43522 , n43523 , n43524 , n43525 , n43526 , n43527 , n43528 , n43529 , n43530 , n43531 , n43532 , n43533 , n43534 , n43535 , n43536 , n43537 , n43538 , n43539 , n43540 , n43541 , n43542 , n43543 , n43544 , n43545 , n43546 , n43547 , n43548 , n43549 , n43550 , n43551 , n43552 , n43553 , n43554 , n43555 , n43556 , n43557 , n43558 , n43559 , n43560 , n43561 , n43562 , n43563 , n43564 , n43565 , n43566 , n43567 , n43568 , n43569 , n43570 , n43571 , n43572 , n43573 , n43574 , n43575 , n43576 , n43577 , n43578 , n43579 , n43580 , n43581 , n43582 , n43583 , n43584 , n43585 , n43586 , n43587 , n43588 , n43589 , n43590 , n43591 , n43592 , n43593 , n43594 , n43595 , n43596 , n43597 , n43598 , n43599 , n43600 , n43601 , n43602 , n43603 , n43604 , n43605 , n43606 , n43607 , n43608 , n43609 , n43610 , n43611 , n43612 , n43613 , n43614 , n43615 , n43616 , n43617 , n43618 , n43619 , n43620 , n43621 , n43622 , n43623 , n43624 , n43625 , n43626 , n43627 , n43628 , n43629 , n43630 , n43631 , n43632 , n43633 , n43634 , n43635 , n43636 , n43637 , n43638 , n43639 , n43640 , n43641 , n43642 , n43643 , n43644 , n43645 , n43646 , n43647 , n43648 , n43649 , n43650 , n43651 , n43652 , n43653 , n43654 , n43655 , n43656 , n43657 , n43658 , n43659 , n43660 , n43661 , n43662 , n43663 , n43664 , n43665 , n43666 , n43667 , n43668 , n43669 , n43670 , n43671 , n43672 , n43673 , n43674 , n43675 , n43676 , n43677 , n43678 , n43679 , n43680 , n43681 , n43682 , n43683 , n43684 , n43685 , n43686 , n43687 , n43688 , n43689 , n43690 , n43691 , n43692 , n43693 , n43694 , n43695 , n43696 , n43697 , n43698 , n43699 , n43700 , n43701 , n43702 , n43703 , n43704 , n43705 , n43706 , n43707 , n43708 , n43709 , n43710 , n43711 , n43712 , n43713 , n43714 , n43715 , n43716 , n43717 , n43718 , n43719 , n43720 , n43721 , n43722 , n43723 , n43724 , n43725 , n43726 , n43727 , n43728 , n43729 , n43730 , n43731 , n43732 , n43733 , n43734 , n43735 , n43736 , n43737 , n43738 , n43739 , n43740 , n43741 , n43742 , n43743 , n43744 , n43745 , n43746 , n43747 , n43748 , n43749 , n43750 , n43751 , n43752 , n43753 , n43754 , n43755 , n43756 , n43757 , n43758 , n43759 , n43760 , n43761 , n43762 , n43763 , n43764 , n43765 , n43766 , n43767 , n43768 , n43769 , n43770 , n43771 , n43772 , n43773 , n43774 , n43775 , n43776 , n43777 , n43778 , n43779 , n43780 , n43781 , n43782 , n43783 , n43784 , n43785 , n43786 , n43787 , n43788 , n43789 , n43790 , n43791 , n43792 , n43793 , n43794 , n43795 , n43796 , n43797 , n43798 , n43799 , n43800 , n43801 , n43802 , n43803 , n43804 , n43805 , n43806 , n43807 , n43808 , n43809 , n43810 , n43811 , n43812 , n43813 , n43814 , n43815 , n43816 , n43817 , n43818 , n43819 , n43820 , n43821 , n43822 , n43823 , n43824 , n43825 , n43826 , n43827 , n43828 , n43829 , n43830 , n43831 , n43832 , n43833 , n43834 , n43835 , n43836 , n43837 , n43838 , n43839 , n43840 , n43841 , n43842 , n43843 , n43844 , n43845 , n43846 , n43847 , n43848 , n43849 , n43850 , n43851 , n43852 , n43853 , n43854 , n43855 , n43856 , n43857 , n43858 , n43859 , n43860 , n43861 , n43862 , n43863 , n43864 , n43865 , n43866 , n43867 , n43868 , n43869 , n43870 , n43871 , n43872 , n43873 , n43874 , n43875 , n43876 , n43877 , n43878 , n43879 , n43880 , n43881 , n43882 , n43883 , n43884 , n43885 , n43886 , n43887 , n43888 , n43889 , n43890 , n43891 , n43892 , n43893 , n43894 , n43895 , n43896 , n43897 , n43898 , n43899 , n43900 , n43901 , n43902 , n43903 , n43904 , n43905 , n43906 , n43907 , n43908 , n43909 , n43910 , n43911 , n43912 , n43913 , n43914 , n43915 , n43916 , n43917 , n43918 , n43919 , n43920 , n43921 , n43922 , n43923 , n43924 , n43925 , n43926 , n43927 , n43928 , n43929 , n43930 , n43931 , n43932 , n43933 , n43934 , n43935 , n43936 , n43937 , n43938 , n43939 , n43940 , n43941 , n43942 , n43943 , n43944 , n43945 , n43946 , n43947 , n43948 , n43949 , n43950 , n43951 , n43952 , n43953 , n43954 , n43955 , n43956 , n43957 , n43958 , n43959 , n43960 , n43961 , n43962 , n43963 , n43964 , n43965 , n43966 , n43967 , n43968 , n43969 , n43970 , n43971 , n43972 , n43973 , n43974 , n43975 , n43976 , n43977 , n43978 , n43979 , n43980 , n43981 , n43982 , n43983 , n43984 , n43985 , n43986 , n43987 , n43988 , n43989 , n43990 , n43991 , n43992 , n43993 , n43994 , n43995 , n43996 , n43997 , n43998 , n43999 , n44000 , n44001 , n44002 , n44003 , n44004 , n44005 , n44006 , n44007 , n44008 , n44009 , n44010 , n44011 , n44012 , n44013 , n44014 , n44015 , n44016 , n44017 , n44018 , n44019 , n44020 , n44021 , n44022 , n44023 , n44024 , n44025 , n44026 , n44027 , n44028 , n44029 , n44030 , n44031 , n44032 , n44033 , n44034 , n44035 , n44036 , n44037 , n44038 , n44039 , n44040 , n44041 , n44042 , n44043 , n44044 , n44045 , n44046 , n44047 , n44048 , n44049 , n44050 , n44051 , n44052 , n44053 , n44054 , n44055 , n44056 , n44057 , n44058 , n44059 , n44060 , n44061 , n44062 , n44063 , n44064 , n44065 , n44066 , n44067 , n44068 , n44069 , n44070 , n44071 , n44072 , n44073 , n44074 , n44075 , n44076 , n44077 , n44078 , n44079 , n44080 , n44081 , n44082 , n44083 , n44084 , n44085 , n44086 , n44087 , n44088 , n44089 , n44090 , n44091 , n44092 , n44093 , n44094 , n44095 , n44096 , n44097 , n44098 , n44099 , n44100 , n44101 , n44102 , n44103 , n44104 , n44105 , n44106 , n44107 , n44108 , n44109 , n44110 , n44111 , n44112 , n44113 , n44114 , n44115 , n44116 , n44117 , n44118 , n44119 , n44120 , n44121 , n44122 , n44123 , n44124 , n44125 , n44126 , n44127 , n44128 , n44129 , n44130 , n44131 , n44132 , n44133 , n44134 , n44135 , n44136 , n44137 , n44138 , n44139 , n44140 , n44141 , n44142 , n44143 , n44144 , n44145 , n44146 , n44147 , n44148 , n44149 , n44150 , n44151 , n44152 , n44153 , n44154 , n44155 , n44156 , n44157 , n44158 , n44159 , n44160 , n44161 , n44162 , n44163 , n44164 , n44165 , n44166 , n44167 , n44168 , n44169 , n44170 , n44171 , n44172 , n44173 , n44174 , n44175 , n44176 , n44177 , n44178 , n44179 , n44180 , n44181 , n44182 , n44183 , n44184 , n44185 , n44186 , n44187 , n44188 , n44189 , n44190 , n44191 , n44192 , n44193 , n44194 , n44195 , n44196 , n44197 , n44198 , n44199 , n44200 , n44201 , n44202 , n44203 , n44204 , n44205 , n44206 , n44207 , n44208 , n44209 , n44210 , n44211 , n44212 , n44213 , n44214 , n44215 , n44216 , n44217 , n44218 , n44219 , n44220 , n44221 , n44222 , n44223 , n44224 , n44225 , n44226 , n44227 , n44228 , n44229 , n44230 , n44231 , n44232 , n44233 , n44234 , n44235 , n44236 , n44237 , n44238 , n44239 , n44240 , n44241 , n44242 , n44243 , n44244 , n44245 , n44246 , n44247 , n44248 , n44249 , n44250 , n44251 , n44252 , n44253 , n44254 , n44255 , n44256 , n44257 , n44258 , n44259 , n44260 , n44261 , n44262 , n44263 , n44264 , n44265 , n44266 , n44267 , n44268 , n44269 , n44270 , n44271 , n44272 , n44273 , n44274 , n44275 , n44276 , n44277 , n44278 , n44279 , n44280 , n44281 , n44282 , n44283 , n44284 , n44285 , n44286 , n44287 , n44288 , n44289 , n44290 , n44291 , n44292 , n44293 , n44294 , n44295 , n44296 , n44297 , n44298 , n44299 , n44300 , n44301 , n44302 , n44303 , n44304 , n44305 , n44306 , n44307 , n44308 , n44309 , n44310 , n44311 , n44312 , n44313 , n44314 , n44315 , n44316 , n44317 , n44318 , n44319 , n44320 , n44321 , n44322 , n44323 , n44324 , n44325 , n44326 , n44327 , n44328 , n44329 , n44330 , n44331 , n44332 , n44333 , n44334 , n44335 , n44336 , n44337 , n44338 , n44339 , n44340 , n44341 , n44342 , n44343 , n44344 , n44345 , n44346 , n44347 , n44348 , n44349 , n44350 , n44351 , n44352 , n44353 , n44354 , n44355 , n44356 , n44357 , n44358 , n44359 , n44360 , n44361 , n44362 , n44363 , n44364 , n44365 , n44366 , n44367 , n44368 , n44369 , n44370 , n44371 , n44372 , n44373 , n44374 , n44375 , n44376 , n44377 , n44378 , n44379 , n44380 , n44381 , n44382 , n44383 , n44384 , n44385 , n44386 , n44387 , n44388 , n44389 , n44390 , n44391 , n44392 , n44393 , n44394 , n44395 , n44396 , n44397 , n44398 , n44399 , n44400 , n44401 , n44402 , n44403 , n44404 , n44405 , n44406 , n44407 , n44408 , n44409 , n44410 , n44411 , n44412 , n44413 , n44414 , n44415 , n44416 , n44417 , n44418 , n44419 , n44420 , n44421 , n44422 , n44423 , n44424 , n44425 , n44426 , n44427 , n44428 , n44429 , n44430 , n44431 , n44432 , n44433 , n44434 , n44435 , n44436 , n44437 , n44438 , n44439 , n44440 , n44441 , n44442 , n44443 , n44444 , n44445 , n44446 , n44447 , n44448 , n44449 , n44450 , n44451 , n44452 , n44453 , n44454 , n44455 , n44456 , n44457 , n44458 , n44459 , n44460 , n44461 , n44462 , n44463 , n44464 , n44465 , n44466 , n44467 , n44468 , n44469 , n44470 , n44471 , n44472 , n44473 , n44474 , n44475 , n44476 , n44477 , n44478 , n44479 , n44480 , n44481 , n44482 , n44483 , n44484 , n44485 , n44486 , n44487 , n44488 , n44489 , n44490 , n44491 , n44492 , n44493 , n44494 , n44495 , n44496 , n44497 , n44498 , n44499 , n44500 , n44501 , n44502 , n44503 , n44504 , n44505 , n44506 , n44507 , n44508 , n44509 , n44510 , n44511 , n44512 , n44513 , n44514 , n44515 , n44516 , n44517 , n44518 , n44519 , n44520 , n44521 , n44522 , n44523 , n44524 , n44525 , n44526 , n44527 , n44528 , n44529 , n44530 , n44531 , n44532 , n44533 , n44534 , n44535 , n44536 , n44537 , n44538 , n44539 , n44540 , n44541 , n44542 , n44543 , n44544 , n44545 , n44546 , n44547 , n44548 , n44549 , n44550 , n44551 , n44552 , n44553 , n44554 , n44555 , n44556 , n44557 , n44558 , n44559 , n44560 , n44561 , n44562 , n44563 , n44564 , n44565 , n44566 , n44567 , n44568 , n44569 , n44570 , n44571 , n44572 , n44573 , n44574 , n44575 , n44576 , n44577 , n44578 , n44579 , n44580 , n44581 , n44582 , n44583 , n44584 , n44585 , n44586 , n44587 , n44588 , n44589 , n44590 , n44591 , n44592 , n44593 , n44594 , n44595 , n44596 , n44597 , n44598 , n44599 , n44600 , n44601 , n44602 , n44603 , n44604 , n44605 , n44606 , n44607 , n44608 , n44609 , n44610 , n44611 , n44612 , n44613 , n44614 , n44615 , n44616 , n44617 , n44618 , n44619 , n44620 , n44621 , n44622 , n44623 , n44624 , n44625 , n44626 , n44627 , n44628 , n44629 , n44630 , n44631 , n44632 , n44633 , n44634 , n44635 , n44636 , n44637 , n44638 , n44639 , n44640 , n44641 , n44642 , n44643 , n44644 , n44645 , n44646 , n44647 , n44648 , n44649 , n44650 , n44651 , n44652 , n44653 , n44654 , n44655 , n44656 , n44657 , n44658 , n44659 , n44660 , n44661 , n44662 , n44663 , n44664 , n44665 , n44666 , n44667 , n44668 , n44669 , n44670 , n44671 , n44672 , n44673 , n44674 , n44675 , n44676 , n44677 , n44678 , n44679 , n44680 , n44681 , n44682 , n44683 , n44684 , n44685 , n44686 , n44687 , n44688 , n44689 , n44690 , n44691 , n44692 , n44693 , n44694 , n44695 , n44696 , n44697 , n44698 , n44699 , n44700 , n44701 , n44702 , n44703 , n44704 , n44705 , n44706 , n44707 , n44708 , n44709 , n44710 , n44711 , n44712 , n44713 , n44714 , n44715 , n44716 , n44717 , n44718 , n44719 , n44720 , n44721 , n44722 , n44723 , n44724 , n44725 , n44726 , n44727 , n44728 , n44729 , n44730 , n44731 , n44732 , n44733 , n44734 , n44735 , n44736 , n44737 , n44738 , n44739 , n44740 , n44741 , n44742 , n44743 , n44744 , n44745 , n44746 , n44747 , n44748 , n44749 , n44750 , n44751 , n44752 , n44753 , n44754 , n44755 , n44756 , n44757 , n44758 , n44759 , n44760 , n44761 , n44762 , n44763 , n44764 , n44765 , n44766 , n44767 , n44768 , n44769 , n44770 , n44771 , n44772 , n44773 , n44774 , n44775 , n44776 , n44777 , n44778 , n44779 , n44780 , n44781 , n44782 , n44783 , n44784 , n44785 , n44786 , n44787 , n44788 , n44789 , n44790 , n44791 , n44792 , n44793 , n44794 , n44795 , n44796 , n44797 , n44798 , n44799 , n44800 , n44801 , n44802 , n44803 , n44804 , n44805 , n44806 , n44807 , n44808 , n44809 , n44810 , n44811 , n44812 , n44813 , n44814 , n44815 , n44816 , n44817 , n44818 , n44819 , n44820 , n44821 , n44822 , n44823 , n44824 , n44825 , n44826 , n44827 , n44828 , n44829 , n44830 , n44831 , n44832 , n44833 , n44834 , n44835 , n44836 , n44837 , n44838 , n44839 , n44840 , n44841 , n44842 , n44843 , n44844 , n44845 , n44846 , n44847 , n44848 , n44849 , n44850 , n44851 , n44852 , n44853 , n44854 , n44855 , n44856 , n44857 , n44858 , n44859 , n44860 , n44861 , n44862 , n44863 , n44864 , n44865 , n44866 , n44867 , n44868 , n44869 , n44870 , n44871 , n44872 , n44873 , n44874 , n44875 , n44876 , n44877 , n44878 , n44879 , n44880 , n44881 , n44882 , n44883 , n44884 , n44885 , n44886 , n44887 , n44888 , n44889 , n44890 , n44891 , n44892 , n44893 , n44894 , n44895 , n44896 , n44897 , n44898 , n44899 , n44900 , n44901 , n44902 , n44903 , n44904 , n44905 , n44906 , n44907 , n44908 , n44909 , n44910 , n44911 , n44912 , n44913 , n44914 , n44915 , n44916 , n44917 , n44918 , n44919 , n44920 , n44921 , n44922 , n44923 , n44924 , n44925 , n44926 , n44927 , n44928 , n44929 , n44930 , n44931 , n44932 , n44933 , n44934 , n44935 , n44936 , n44937 , n44938 , n44939 , n44940 , n44941 , n44942 , n44943 , n44944 , n44945 , n44946 , n44947 , n44948 , n44949 , n44950 , n44951 , n44952 , n44953 , n44954 , n44955 , n44956 , n44957 , n44958 , n44959 , n44960 , n44961 , n44962 , n44963 , n44964 , n44965 , n44966 , n44967 , n44968 , n44969 , n44970 , n44971 , n44972 , n44973 , n44974 , n44975 , n44976 , n44977 , n44978 , n44979 , n44980 , n44981 , n44982 , n44983 , n44984 , n44985 , n44986 , n44987 , n44988 , n44989 , n44990 , n44991 , n44992 , n44993 , n44994 , n44995 , n44996 , n44997 , n44998 , n44999 , n45000 , n45001 , n45002 , n45003 , n45004 , n45005 , n45006 , n45007 , n45008 , n45009 , n45010 , n45011 , n45012 , n45013 , n45014 , n45015 , n45016 , n45017 , n45018 , n45019 , n45020 , n45021 , n45022 , n45023 , n45024 , n45025 , n45026 , n45027 , n45028 , n45029 , n45030 , n45031 , n45032 , n45033 , n45034 , n45035 , n45036 , n45037 , n45038 , n45039 , n45040 , n45041 , n45042 , n45043 , n45044 , n45045 , n45046 , n45047 , n45048 , n45049 , n45050 , n45051 , n45052 , n45053 , n45054 , n45055 , n45056 , n45057 , n45058 , n45059 , n45060 , n45061 , n45062 , n45063 , n45064 , n45065 , n45066 , n45067 , n45068 , n45069 , n45070 , n45071 , n45072 , n45073 , n45074 , n45075 , n45076 , n45077 , n45078 , n45079 , n45080 , n45081 , n45082 , n45083 , n45084 , n45085 , n45086 , n45087 , n45088 , n45089 , n45090 , n45091 , n45092 , n45093 , n45094 , n45095 , n45096 , n45097 , n45098 , n45099 , n45100 , n45101 , n45102 , n45103 , n45104 , n45105 , n45106 , n45107 , n45108 , n45109 , n45110 , n45111 , n45112 , n45113 , n45114 , n45115 , n45116 , n45117 , n45118 , n45119 , n45120 , n45121 , n45122 , n45123 , n45124 , n45125 , n45126 , n45127 , n45128 , n45129 , n45130 , n45131 , n45132 , n45133 , n45134 , n45135 , n45136 , n45137 , n45138 , n45139 , n45140 , n45141 , n45142 , n45143 , n45144 , n45145 , n45146 , n45147 , n45148 , n45149 , n45150 , n45151 , n45152 , n45153 , n45154 , n45155 , n45156 , n45157 , n45158 , n45159 , n45160 , n45161 , n45162 , n45163 , n45164 , n45165 , n45166 , n45167 , n45168 , n45169 , n45170 , n45171 , n45172 , n45173 , n45174 , n45175 , n45176 , n45177 , n45178 , n45179 , n45180 , n45181 , n45182 , n45183 , n45184 , n45185 , n45186 , n45187 , n45188 , n45189 , n45190 , n45191 , n45192 , n45193 , n45194 , n45195 , n45196 , n45197 , n45198 , n45199 , n45200 , n45201 , n45202 , n45203 , n45204 , n45205 , n45206 , n45207 , n45208 , n45209 , n45210 , n45211 , n45212 , n45213 , n45214 , n45215 , n45216 , n45217 , n45218 , n45219 , n45220 , n45221 , n45222 , n45223 , n45224 , n45225 , n45226 , n45227 , n45228 , n45229 , n45230 , n45231 , n45232 , n45233 , n45234 , n45235 , n45236 , n45237 , n45238 , n45239 , n45240 , n45241 , n45242 , n45243 , n45244 , n45245 , n45246 , n45247 , n45248 , n45249 , n45250 , n45251 , n45252 , n45253 , n45254 , n45255 , n45256 , n45257 , n45258 , n45259 , n45260 , n45261 , n45262 , n45263 , n45264 , n45265 , n45266 , n45267 , n45268 , n45269 , n45270 , n45271 , n45272 , n45273 , n45274 , n45275 , n45276 , n45277 , n45278 , n45279 , n45280 , n45281 , n45282 , n45283 , n45284 , n45285 , n45286 , n45287 , n45288 , n45289 , n45290 , n45291 , n45292 , n45293 , n45294 , n45295 , n45296 , n45297 , n45298 , n45299 , n45300 , n45301 , n45302 , n45303 , n45304 , n45305 , n45306 , n45307 , n45308 , n45309 , n45310 , n45311 , n45312 , n45313 , n45314 , n45315 , n45316 , n45317 , n45318 , n45319 , n45320 , n45321 , n45322 , n45323 , n45324 , n45325 , n45326 , n45327 , n45328 , n45329 , n45330 , n45331 , n45332 , n45333 , n45334 , n45335 , n45336 , n45337 , n45338 , n45339 , n45340 , n45341 , n45342 , n45343 , n45344 , n45345 , n45346 , n45347 , n45348 , n45349 , n45350 , n45351 , n45352 , n45353 , n45354 , n45355 , n45356 , n45357 , n45358 , n45359 , n45360 , n45361 , n45362 , n45363 , n45364 , n45365 , n45366 , n45367 , n45368 , n45369 , n45370 , n45371 , n45372 , n45373 , n45374 , n45375 , n45376 , n45377 , n45378 , n45379 , n45380 , n45381 , n45382 , n45383 , n45384 , n45385 , n45386 , n45387 , n45388 , n45389 , n45390 , n45391 , n45392 , n45393 , n45394 , n45395 , n45396 , n45397 , n45398 , n45399 , n45400 , n45401 , n45402 , n45403 , n45404 , n45405 , n45406 , n45407 , n45408 , n45409 , n45410 , n45411 , n45412 , n45413 , n45414 , n45415 , n45416 , n45417 , n45418 , n45419 , n45420 , n45421 , n45422 , n45423 , n45424 , n45425 , n45426 , n45427 , n45428 , n45429 , n45430 , n45431 , n45432 , n45433 , n45434 , n45435 , n45436 , n45437 , n45438 , n45439 , n45440 , n45441 , n45442 , n45443 , n45444 , n45445 , n45446 , n45447 , n45448 , n45449 , n45450 , n45451 , n45452 , n45453 , n45454 , n45455 , n45456 , n45457 , n45458 , n45459 , n45460 , n45461 , n45462 , n45463 , n45464 , n45465 , n45466 , n45467 , n45468 , n45469 , n45470 , n45471 , n45472 , n45473 , n45474 , n45475 , n45476 , n45477 , n45478 , n45479 , n45480 , n45481 , n45482 , n45483 , n45484 , n45485 , n45486 , n45487 , n45488 , n45489 , n45490 , n45491 , n45492 , n45493 , n45494 , n45495 , n45496 , n45497 , n45498 , n45499 , n45500 , n45501 , n45502 , n45503 , n45504 , n45505 , n45506 , n45507 , n45508 , n45509 , n45510 , n45511 , n45512 , n45513 , n45514 , n45515 , n45516 , n45517 , n45518 , n45519 , n45520 , n45521 , n45522 , n45523 , n45524 , n45525 , n45526 , n45527 , n45528 , n45529 , n45530 , n45531 , n45532 , n45533 , n45534 , n45535 , n45536 , n45537 , n45538 , n45539 , n45540 , n45541 , n45542 , n45543 , n45544 , n45545 , n45546 , n45547 , n45548 , n45549 , n45550 , n45551 , n45552 , n45553 , n45554 , n45555 , n45556 , n45557 , n45558 , n45559 , n45560 , n45561 , n45562 , n45563 , n45564 , n45565 , n45566 , n45567 , n45568 , n45569 , n45570 , n45571 , n45572 , n45573 , n45574 , n45575 , n45576 , n45577 , n45578 , n45579 , n45580 , n45581 , n45582 , n45583 , n45584 , n45585 , n45586 , n45587 , n45588 , n45589 , n45590 , n45591 , n45592 , n45593 , n45594 , n45595 , n45596 , n45597 , n45598 , n45599 , n45600 , n45601 , n45602 , n45603 , n45604 , n45605 , n45606 , n45607 , n45608 , n45609 , n45610 , n45611 , n45612 , n45613 , n45614 , n45615 , n45616 , n45617 , n45618 , n45619 , n45620 , n45621 , n45622 , n45623 , n45624 , n45625 , n45626 , n45627 , n45628 , n45629 , n45630 , n45631 , n45632 , n45633 , n45634 , n45635 , n45636 , n45637 , n45638 , n45639 , n45640 , n45641 , n45642 , n45643 , n45644 , n45645 , n45646 , n45647 , n45648 , n45649 , n45650 , n45651 , n45652 , n45653 , n45654 , n45655 , n45656 , n45657 , n45658 , n45659 , n45660 , n45661 , n45662 , n45663 , n45664 , n45665 , n45666 , n45667 , n45668 , n45669 , n45670 , n45671 , n45672 , n45673 , n45674 , n45675 , n45676 , n45677 , n45678 , n45679 , n45680 , n45681 , n45682 , n45683 , n45684 , n45685 , n45686 , n45687 , n45688 , n45689 , n45690 , n45691 , n45692 , n45693 , n45694 , n45695 , n45696 , n45697 , n45698 , n45699 , n45700 , n45701 , n45702 , n45703 , n45704 , n45705 , n45706 , n45707 , n45708 , n45709 , n45710 , n45711 , n45712 , n45713 , n45714 , n45715 , n45716 , n45717 , n45718 , n45719 , n45720 , n45721 , n45722 , n45723 , n45724 , n45725 , n45726 , n45727 , n45728 , n45729 , n45730 , n45731 , n45732 , n45733 , n45734 , n45735 , n45736 , n45737 , n45738 , n45739 , n45740 , n45741 , n45742 , n45743 , n45744 , n45745 , n45746 , n45747 , n45748 , n45749 , n45750 , n45751 , n45752 , n45753 , n45754 , n45755 , n45756 , n45757 , n45758 , n45759 , n45760 , n45761 , n45762 , n45763 , n45764 , n45765 , n45766 , n45767 , n45768 , n45769 , n45770 , n45771 , n45772 , n45773 , n45774 , n45775 , n45776 , n45777 , n45778 , n45779 , n45780 , n45781 , n45782 , n45783 , n45784 , n45785 , n45786 , n45787 , n45788 , n45789 , n45790 , n45791 , n45792 , n45793 , n45794 , n45795 , n45796 , n45797 , n45798 , n45799 , n45800 , n45801 , n45802 , n45803 , n45804 , n45805 , n45806 , n45807 , n45808 , n45809 , n45810 , n45811 , n45812 , n45813 , n45814 , n45815 , n45816 , n45817 , n45818 , n45819 , n45820 , n45821 , n45822 , n45823 , n45824 , n45825 , n45826 , n45827 , n45828 , n45829 , n45830 , n45831 , n45832 , n45833 , n45834 , n45835 , n45836 , n45837 , n45838 , n45839 , n45840 , n45841 , n45842 , n45843 , n45844 , n45845 , n45846 , n45847 , n45848 , n45849 , n45850 , n45851 , n45852 , n45853 , n45854 , n45855 , n45856 , n45857 , n45858 , n45859 , n45860 , n45861 , n45862 , n45863 , n45864 , n45865 , n45866 , n45867 , n45868 , n45869 , n45870 , n45871 , n45872 , n45873 , n45874 , n45875 , n45876 , n45877 , n45878 , n45879 , n45880 , n45881 , n45882 , n45883 , n45884 , n45885 , n45886 , n45887 , n45888 , n45889 , n45890 , n45891 , n45892 , n45893 , n45894 , n45895 , n45896 , n45897 , n45898 , n45899 , n45900 , n45901 , n45902 , n45903 , n45904 , n45905 , n45906 , n45907 , n45908 , n45909 , n45910 , n45911 , n45912 , n45913 , n45914 , n45915 , n45916 , n45917 , n45918 , n45919 , n45920 , n45921 , n45922 , n45923 , n45924 , n45925 , n45926 , n45927 , n45928 , n45929 , n45930 , n45931 , n45932 , n45933 , n45934 , n45935 , n45936 , n45937 , n45938 , n45939 , n45940 , n45941 , n45942 , n45943 , n45944 , n45945 , n45946 , n45947 , n45948 , n45949 , n45950 , n45951 , n45952 , n45953 , n45954 , n45955 , n45956 , n45957 , n45958 , n45959 , n45960 , n45961 , n45962 , n45963 , n45964 , n45965 , n45966 , n45967 , n45968 , n45969 , n45970 , n45971 , n45972 , n45973 , n45974 , n45975 , n45976 , n45977 , n45978 , n45979 , n45980 , n45981 , n45982 , n45983 , n45984 , n45985 , n45986 , n45987 , n45988 , n45989 , n45990 , n45991 , n45992 , n45993 , n45994 , n45995 , n45996 , n45997 , n45998 , n45999 , n46000 , n46001 , n46002 , n46003 , n46004 , n46005 , n46006 , n46007 , n46008 , n46009 , n46010 , n46011 , n46012 , n46013 , n46014 , n46015 , n46016 , n46017 , n46018 , n46019 , n46020 , n46021 , n46022 , n46023 , n46024 , n46025 , n46026 , n46027 , n46028 , n46029 , n46030 , n46031 , n46032 , n46033 , n46034 , n46035 , n46036 , n46037 , n46038 , n46039 , n46040 , n46041 , n46042 , n46043 , n46044 , n46045 , n46046 , n46047 , n46048 , n46049 , n46050 , n46051 , n46052 , n46053 , n46054 , n46055 , n46056 , n46057 , n46058 , n46059 , n46060 , n46061 , n46062 , n46063 , n46064 , n46065 , n46066 , n46067 , n46068 , n46069 , n46070 , n46071 , n46072 , n46073 , n46074 , n46075 , n46076 , n46077 , n46078 , n46079 , n46080 , n46081 , n46082 , n46083 , n46084 , n46085 , n46086 , n46087 , n46088 , n46089 , n46090 , n46091 , n46092 , n46093 , n46094 , n46095 , n46096 , n46097 , n46098 , n46099 , n46100 , n46101 , n46102 , n46103 , n46104 , n46105 , n46106 , n46107 , n46108 , n46109 , n46110 , n46111 , n46112 , n46113 , n46114 , n46115 , n46116 , n46117 , n46118 , n46119 , n46120 , n46121 , n46122 , n46123 , n46124 , n46125 , n46126 , n46127 , n46128 , n46129 , n46130 , n46131 , n46132 , n46133 , n46134 , n46135 , n46136 , n46137 , n46138 , n46139 , n46140 , n46141 , n46142 , n46143 , n46144 , n46145 , n46146 , n46147 , n46148 , n46149 , n46150 , n46151 , n46152 , n46153 , n46154 , n46155 , n46156 , n46157 , n46158 , n46159 , n46160 , n46161 , n46162 , n46163 , n46164 , n46165 , n46166 , n46167 , n46168 , n46169 , n46170 , n46171 , n46172 , n46173 , n46174 , n46175 , n46176 , n46177 , n46178 , n46179 , n46180 , n46181 , n46182 , n46183 , n46184 , n46185 , n46186 , n46187 , n46188 , n46189 , n46190 , n46191 , n46192 , n46193 , n46194 , n46195 , n46196 , n46197 , n46198 , n46199 , n46200 , n46201 , n46202 , n46203 , n46204 , n46205 , n46206 , n46207 , n46208 , n46209 , n46210 , n46211 , n46212 , n46213 , n46214 , n46215 , n46216 , n46217 , n46218 , n46219 , n46220 , n46221 , n46222 , n46223 , n46224 , n46225 , n46226 , n46227 , n46228 , n46229 , n46230 , n46231 , n46232 , n46233 , n46234 , n46235 , n46236 , n46237 , n46238 , n46239 , n46240 , n46241 , n46242 , n46243 , n46244 , n46245 , n46246 , n46247 , n46248 , n46249 , n46250 , n46251 , n46252 , n46253 , n46254 , n46255 , n46256 , n46257 , n46258 , n46259 , n46260 , n46261 , n46262 , n46263 , n46264 , n46265 , n46266 , n46267 , n46268 , n46269 , n46270 , n46271 , n46272 , n46273 , n46274 , n46275 , n46276 , n46277 , n46278 , n46279 , n46280 , n46281 , n46282 , n46283 , n46284 , n46285 , n46286 , n46287 , n46288 , n46289 , n46290 , n46291 , n46292 , n46293 , n46294 , n46295 , n46296 , n46297 , n46298 , n46299 , n46300 , n46301 , n46302 , n46303 , n46304 , n46305 , n46306 , n46307 , n46308 , n46309 , n46310 , n46311 , n46312 , n46313 , n46314 , n46315 , n46316 , n46317 , n46318 , n46319 , n46320 , n46321 , n46322 , n46323 , n46324 , n46325 , n46326 , n46327 , n46328 , n46329 , n46330 , n46331 , n46332 , n46333 , n46334 , n46335 , n46336 , n46337 , n46338 , n46339 , n46340 , n46341 , n46342 , n46343 , n46344 , n46345 , n46346 , n46347 , n46348 , n46349 , n46350 , n46351 , n46352 , n46353 , n46354 , n46355 , n46356 , n46357 , n46358 , n46359 , n46360 , n46361 , n46362 , n46363 , n46364 , n46365 , n46366 , n46367 , n46368 , n46369 , n46370 , n46371 , n46372 , n46373 , n46374 , n46375 , n46376 , n46377 , n46378 , n46379 , n46380 , n46381 , n46382 , n46383 , n46384 , n46385 , n46386 , n46387 , n46388 , n46389 , n46390 , n46391 , n46392 , n46393 , n46394 , n46395 , n46396 , n46397 , n46398 , n46399 , n46400 , n46401 , n46402 , n46403 , n46404 , n46405 , n46406 , n46407 , n46408 , n46409 , n46410 , n46411 , n46412 , n46413 , n46414 , n46415 , n46416 , n46417 , n46418 , n46419 , n46420 , n46421 , n46422 , n46423 , n46424 , n46425 , n46426 , n46427 , n46428 , n46429 , n46430 , n46431 , n46432 , n46433 , n46434 , n46435 , n46436 , n46437 , n46438 , n46439 , n46440 , n46441 , n46442 , n46443 , n46444 , n46445 , n46446 , n46447 , n46448 , n46449 , n46450 , n46451 , n46452 , n46453 , n46454 , n46455 , n46456 , n46457 , n46458 , n46459 , n46460 , n46461 , n46462 , n46463 , n46464 , n46465 , n46466 , n46467 , n46468 , n46469 , n46470 , n46471 , n46472 , n46473 , n46474 , n46475 , n46476 , n46477 , n46478 , n46479 , n46480 , n46481 , n46482 , n46483 , n46484 , n46485 , n46486 , n46487 , n46488 , n46489 , n46490 , n46491 , n46492 , n46493 , n46494 , n46495 , n46496 , n46497 , n46498 , n46499 , n46500 , n46501 , n46502 , n46503 , n46504 , n46505 , n46506 , n46507 , n46508 , n46509 , n46510 , n46511 , n46512 , n46513 , n46514 , n46515 , n46516 , n46517 , n46518 , n46519 , n46520 , n46521 , n46522 , n46523 , n46524 , n46525 , n46526 , n46527 , n46528 , n46529 , n46530 , n46531 , n46532 , n46533 , n46534 , n46535 , n46536 , n46537 , n46538 , n46539 , n46540 , n46541 , n46542 , n46543 , n46544 , n46545 , n46546 , n46547 , n46548 , n46549 , n46550 , n46551 , n46552 , n46553 , n46554 , n46555 , n46556 , n46557 , n46558 , n46559 , n46560 , n46561 , n46562 , n46563 , n46564 , n46565 , n46566 , n46567 , n46568 , n46569 , n46570 , n46571 , n46572 , n46573 , n46574 , n46575 , n46576 , n46577 , n46578 , n46579 , n46580 , n46581 , n46582 , n46583 , n46584 , n46585 , n46586 , n46587 , n46588 , n46589 , n46590 , n46591 , n46592 , n46593 , n46594 , n46595 , n46596 , n46597 , n46598 , n46599 , n46600 , n46601 , n46602 , n46603 , n46604 , n46605 , n46606 , n46607 , n46608 , n46609 , n46610 , n46611 , n46612 , n46613 , n46614 , n46615 , n46616 , n46617 , n46618 , n46619 , n46620 , n46621 , n46622 , n46623 , n46624 , n46625 , n46626 , n46627 , n46628 , n46629 , n46630 , n46631 , n46632 , n46633 , n46634 , n46635 , n46636 , n46637 , n46638 , n46639 , n46640 , n46641 , n46642 , n46643 , n46644 , n46645 , n46646 , n46647 , n46648 , n46649 , n46650 , n46651 , n46652 , n46653 , n46654 , n46655 , n46656 , n46657 , n46658 , n46659 , n46660 , n46661 , n46662 , n46663 , n46664 , n46665 , n46666 , n46667 , n46668 , n46669 , n46670 , n46671 , n46672 , n46673 , n46674 , n46675 , n46676 , n46677 , n46678 , n46679 , n46680 , n46681 , n46682 , n46683 , n46684 , n46685 , n46686 , n46687 , n46688 , n46689 , n46690 , n46691 , n46692 , n46693 , n46694 , n46695 , n46696 , n46697 , n46698 , n46699 , n46700 , n46701 , n46702 , n46703 , n46704 , n46705 , n46706 , n46707 , n46708 , n46709 , n46710 , n46711 , n46712 , n46713 , n46714 , n46715 , n46716 , n46717 , n46718 , n46719 , n46720 , n46721 , n46722 , n46723 , n46724 , n46725 , n46726 , n46727 , n46728 , n46729 , n46730 , n46731 , n46732 , n46733 , n46734 , n46735 , n46736 , n46737 , n46738 , n46739 , n46740 , n46741 , n46742 , n46743 , n46744 , n46745 , n46746 , n46747 , n46748 , n46749 , n46750 , n46751 , n46752 , n46753 , n46754 , n46755 , n46756 , n46757 , n46758 , n46759 , n46760 , n46761 , n46762 , n46763 , n46764 , n46765 , n46766 , n46767 , n46768 , n46769 , n46770 , n46771 , n46772 , n46773 , n46774 , n46775 , n46776 , n46777 , n46778 , n46779 , n46780 , n46781 , n46782 , n46783 , n46784 , n46785 , n46786 , n46787 , n46788 , n46789 , n46790 , n46791 , n46792 , n46793 , n46794 , n46795 , n46796 , n46797 , n46798 , n46799 , n46800 , n46801 , n46802 , n46803 , n46804 , n46805 , n46806 , n46807 , n46808 , n46809 , n46810 , n46811 , n46812 , n46813 , n46814 , n46815 , n46816 , n46817 , n46818 , n46819 , n46820 , n46821 , n46822 , n46823 , n46824 , n46825 , n46826 , n46827 , n46828 , n46829 , n46830 , n46831 , n46832 , n46833 , n46834 , n46835 , n46836 , n46837 , n46838 , n46839 , n46840 , n46841 , n46842 , n46843 , n46844 , n46845 , n46846 , n46847 , n46848 , n46849 , n46850 , n46851 , n46852 , n46853 , n46854 , n46855 , n46856 , n46857 , n46858 , n46859 , n46860 , n46861 , n46862 , n46863 , n46864 , n46865 , n46866 , n46867 , n46868 , n46869 , n46870 , n46871 , n46872 , n46873 , n46874 , n46875 , n46876 , n46877 , n46878 , n46879 , n46880 , n46881 , n46882 , n46883 , n46884 , n46885 , n46886 , n46887 , n46888 , n46889 , n46890 , n46891 , n46892 , n46893 , n46894 , n46895 , n46896 , n46897 , n46898 , n46899 , n46900 , n46901 , n46902 , n46903 , n46904 , n46905 , n46906 , n46907 , n46908 , n46909 , n46910 , n46911 , n46912 , n46913 , n46914 , n46915 , n46916 , n46917 , n46918 , n46919 , n46920 , n46921 , n46922 , n46923 , n46924 , n46925 , n46926 , n46927 , n46928 , n46929 , n46930 , n46931 , n46932 , n46933 , n46934 , n46935 , n46936 , n46937 , n46938 , n46939 , n46940 , n46941 , n46942 , n46943 , n46944 , n46945 , n46946 , n46947 , n46948 , n46949 , n46950 , n46951 , n46952 , n46953 , n46954 , n46955 , n46956 , n46957 , n46958 , n46959 , n46960 , n46961 , n46962 , n46963 , n46964 , n46965 , n46966 , n46967 , n46968 , n46969 , n46970 , n46971 , n46972 , n46973 , n46974 , n46975 , n46976 , n46977 , n46978 , n46979 , n46980 , n46981 , n46982 , n46983 , n46984 , n46985 , n46986 , n46987 , n46988 , n46989 , n46990 , n46991 , n46992 , n46993 , n46994 , n46995 , n46996 , n46997 , n46998 , n46999 , n47000 , n47001 , n47002 , n47003 , n47004 , n47005 , n47006 , n47007 , n47008 , n47009 , n47010 , n47011 , n47012 , n47013 , n47014 , n47015 , n47016 , n47017 , n47018 , n47019 , n47020 , n47021 , n47022 , n47023 , n47024 , n47025 , n47026 , n47027 , n47028 , n47029 , n47030 , n47031 , n47032 , n47033 , n47034 , n47035 , n47036 , n47037 , n47038 , n47039 , n47040 , n47041 , n47042 , n47043 , n47044 , n47045 , n47046 , n47047 , n47048 , n47049 , n47050 , n47051 , n47052 , n47053 , n47054 , n47055 , n47056 , n47057 , n47058 , n47059 , n47060 , n47061 , n47062 , n47063 , n47064 , n47065 , n47066 , n47067 , n47068 , n47069 , n47070 , n47071 , n47072 , n47073 , n47074 , n47075 , n47076 , n47077 , n47078 , n47079 , n47080 , n47081 , n47082 , n47083 , n47084 , n47085 , n47086 , n47087 , n47088 , n47089 , n47090 , n47091 , n47092 , n47093 , n47094 , n47095 , n47096 , n47097 , n47098 , n47099 , n47100 , n47101 , n47102 , n47103 , n47104 , n47105 , n47106 , n47107 , n47108 , n47109 , n47110 , n47111 , n47112 , n47113 , n47114 , n47115 , n47116 , n47117 , n47118 , n47119 , n47120 , n47121 , n47122 , n47123 , n47124 , n47125 , n47126 , n47127 , n47128 , n47129 , n47130 , n47131 , n47132 , n47133 , n47134 , n47135 , n47136 , n47137 , n47138 , n47139 , n47140 , n47141 , n47142 , n47143 , n47144 , n47145 , n47146 , n47147 , n47148 , n47149 , n47150 , n47151 , n47152 , n47153 , n47154 , n47155 , n47156 , n47157 , n47158 , n47159 , n47160 , n47161 , n47162 , n47163 , n47164 , n47165 , n47166 , n47167 , n47168 , n47169 , n47170 , n47171 , n47172 , n47173 , n47174 , n47175 , n47176 , n47177 , n47178 , n47179 , n47180 , n47181 , n47182 , n47183 , n47184 , n47185 , n47186 , n47187 , n47188 , n47189 , n47190 , n47191 , n47192 , n47193 , n47194 , n47195 , n47196 , n47197 , n47198 , n47199 , n47200 , n47201 , n47202 , n47203 , n47204 , n47205 , n47206 , n47207 , n47208 , n47209 , n47210 , n47211 , n47212 , n47213 , n47214 , n47215 , n47216 , n47217 , n47218 , n47219 , n47220 , n47221 , n47222 , n47223 , n47224 , n47225 , n47226 , n47227 , n47228 , n47229 , n47230 , n47231 , n47232 , n47233 , n47234 , n47235 , n47236 , n47237 , n47238 , n47239 , n47240 , n47241 , n47242 , n47243 , n47244 , n47245 , n47246 , n47247 , n47248 , n47249 , n47250 , n47251 , n47252 , n47253 , n47254 , n47255 , n47256 , n47257 , n47258 , n47259 , n47260 , n47261 , n47262 , n47263 , n47264 , n47265 , n47266 , n47267 , n47268 , n47269 , n47270 , n47271 , n47272 , n47273 , n47274 , n47275 , n47276 , n47277 , n47278 , n47279 , n47280 , n47281 , n47282 , n47283 , n47284 , n47285 , n47286 , n47287 , n47288 , n47289 , n47290 , n47291 , n47292 , n47293 , n47294 , n47295 , n47296 , n47297 , n47298 , n47299 , n47300 , n47301 , n47302 , n47303 , n47304 , n47305 , n47306 , n47307 , n47308 , n47309 , n47310 , n47311 , n47312 , n47313 , n47314 , n47315 , n47316 , n47317 , n47318 , n47319 , n47320 , n47321 , n47322 , n47323 , n47324 , n47325 , n47326 , n47327 , n47328 , n47329 , n47330 , n47331 , n47332 , n47333 , n47334 , n47335 , n47336 , n47337 , n47338 , n47339 , n47340 , n47341 , n47342 , n47343 , n47344 , n47345 , n47346 , n47347 , n47348 , n47349 , n47350 , n47351 , n47352 , n47353 , n47354 , n47355 , n47356 , n47357 , n47358 , n47359 , n47360 , n47361 , n47362 , n47363 , n47364 , n47365 , n47366 , n47367 , n47368 , n47369 , n47370 , n47371 , n47372 , n47373 , n47374 , n47375 , n47376 , n47377 , n47378 , n47379 , n47380 , n47381 , n47382 , n47383 , n47384 , n47385 , n47386 , n47387 , n47388 , n47389 , n47390 , n47391 , n47392 , n47393 , n47394 , n47395 , n47396 , n47397 , n47398 , n47399 , n47400 , n47401 , n47402 , n47403 , n47404 , n47405 , n47406 , n47407 , n47408 , n47409 , n47410 , n47411 , n47412 , n47413 , n47414 , n47415 , n47416 , n47417 , n47418 , n47419 , n47420 , n47421 , n47422 , n47423 , n47424 , n47425 , n47426 , n47427 , n47428 , n47429 , n47430 , n47431 , n47432 , n47433 , n47434 , n47435 , n47436 , n47437 , n47438 , n47439 , n47440 , n47441 , n47442 , n47443 , n47444 , n47445 , n47446 , n47447 , n47448 , n47449 , n47450 , n47451 , n47452 , n47453 , n47454 , n47455 , n47456 , n47457 , n47458 , n47459 , n47460 , n47461 , n47462 , n47463 , n47464 , n47465 , n47466 , n47467 , n47468 , n47469 , n47470 , n47471 , n47472 , n47473 , n47474 , n47475 , n47476 , n47477 , n47478 , n47479 , n47480 , n47481 , n47482 , n47483 , n47484 , n47485 , n47486 , n47487 , n47488 , n47489 , n47490 , n47491 , n47492 , n47493 , n47494 , n47495 , n47496 , n47497 , n47498 , n47499 , n47500 , n47501 , n47502 , n47503 , n47504 , n47505 , n47506 , n47507 , n47508 , n47509 , n47510 , n47511 , n47512 , n47513 , n47514 , n47515 , n47516 , n47517 , n47518 , n47519 , n47520 , n47521 , n47522 , n47523 , n47524 , n47525 , n47526 , n47527 , n47528 , n47529 , n47530 , n47531 , n47532 , n47533 , n47534 , n47535 , n47536 , n47537 , n47538 , n47539 , n47540 , n47541 , n47542 , n47543 , n47544 , n47545 , n47546 , n47547 , n47548 , n47549 , n47550 , n47551 , n47552 , n47553 , n47554 , n47555 , n47556 , n47557 , n47558 , n47559 , n47560 , n47561 , n47562 , n47563 , n47564 , n47565 , n47566 , n47567 , n47568 , n47569 , n47570 , n47571 , n47572 , n47573 , n47574 , n47575 , n47576 , n47577 , n47578 , n47579 , n47580 , n47581 , n47582 , n47583 , n47584 , n47585 , n47586 , n47587 , n47588 , n47589 , n47590 , n47591 , n47592 , n47593 , n47594 , n47595 , n47596 , n47597 , n47598 , n47599 , n47600 , n47601 , n47602 , n47603 , n47604 , n47605 , n47606 , n47607 , n47608 , n47609 , n47610 , n47611 , n47612 , n47613 , n47614 , n47615 , n47616 , n47617 , n47618 , n47619 , n47620 , n47621 , n47622 , n47623 , n47624 , n47625 , n47626 , n47627 , n47628 , n47629 , n47630 , n47631 , n47632 , n47633 , n47634 , n47635 , n47636 , n47637 , n47638 , n47639 , n47640 , n47641 , n47642 , n47643 , n47644 , n47645 , n47646 , n47647 , n47648 , n47649 , n47650 , n47651 , n47652 , n47653 , n47654 , n47655 , n47656 , n47657 , n47658 , n47659 , n47660 , n47661 , n47662 , n47663 , n47664 , n47665 , n47666 , n47667 , n47668 , n47669 , n47670 , n47671 , n47672 , n47673 , n47674 , n47675 , n47676 , n47677 , n47678 , n47679 , n47680 , n47681 , n47682 , n47683 , n47684 , n47685 , n47686 , n47687 , n47688 , n47689 , n47690 , n47691 , n47692 , n47693 , n47694 , n47695 , n47696 , n47697 , n47698 , n47699 , n47700 , n47701 , n47702 , n47703 , n47704 , n47705 , n47706 , n47707 , n47708 , n47709 , n47710 , n47711 , n47712 , n47713 , n47714 , n47715 , n47716 , n47717 , n47718 , n47719 , n47720 , n47721 , n47722 , n47723 , n47724 , n47725 , n47726 , n47727 , n47728 , n47729 , n47730 , n47731 , n47732 , n47733 , n47734 , n47735 , n47736 , n47737 , n47738 , n47739 , n47740 , n47741 , n47742 , n47743 , n47744 , n47745 , n47746 , n47747 , n47748 , n47749 , n47750 , n47751 , n47752 , n47753 , n47754 , n47755 , n47756 , n47757 , n47758 , n47759 , n47760 , n47761 , n47762 , n47763 , n47764 , n47765 , n47766 , n47767 , n47768 , n47769 , n47770 , n47771 , n47772 , n47773 , n47774 , n47775 , n47776 , n47777 , n47778 , n47779 , n47780 , n47781 , n47782 , n47783 , n47784 , n47785 , n47786 , n47787 , n47788 , n47789 , n47790 , n47791 , n47792 , n47793 , n47794 , n47795 , n47796 , n47797 , n47798 , n47799 , n47800 , n47801 , n47802 , n47803 , n47804 , n47805 , n47806 , n47807 , n47808 , n47809 , n47810 , n47811 , n47812 , n47813 , n47814 , n47815 , n47816 , n47817 , n47818 , n47819 , n47820 , n47821 , n47822 , n47823 , n47824 , n47825 , n47826 , n47827 , n47828 , n47829 , n47830 , n47831 , n47832 , n47833 , n47834 , n47835 , n47836 , n47837 , n47838 , n47839 , n47840 , n47841 , n47842 , n47843 , n47844 , n47845 , n47846 , n47847 , n47848 , n47849 , n47850 , n47851 , n47852 , n47853 , n47854 , n47855 , n47856 , n47857 , n47858 , n47859 , n47860 , n47861 , n47862 , n47863 , n47864 , n47865 , n47866 , n47867 , n47868 , n47869 , n47870 , n47871 , n47872 , n47873 , n47874 , n47875 , n47876 , n47877 , n47878 , n47879 , n47880 , n47881 , n47882 , n47883 , n47884 , n47885 , n47886 , n47887 , n47888 , n47889 , n47890 , n47891 , n47892 , n47893 , n47894 , n47895 , n47896 , n47897 , n47898 , n47899 , n47900 , n47901 , n47902 , n47903 , n47904 , n47905 , n47906 , n47907 , n47908 , n47909 , n47910 , n47911 , n47912 , n47913 , n47914 , n47915 , n47916 , n47917 , n47918 , n47919 , n47920 , n47921 , n47922 , n47923 , n47924 , n47925 , n47926 , n47927 , n47928 , n47929 , n47930 , n47931 , n47932 , n47933 , n47934 , n47935 , n47936 , n47937 , n47938 , n47939 , n47940 , n47941 , n47942 , n47943 , n47944 , n47945 , n47946 , n47947 , n47948 , n47949 , n47950 , n47951 , n47952 , n47953 , n47954 , n47955 , n47956 , n47957 , n47958 , n47959 , n47960 , n47961 , n47962 , n47963 , n47964 , n47965 , n47966 , n47967 , n47968 , n47969 , n47970 , n47971 , n47972 , n47973 , n47974 , n47975 , n47976 , n47977 , n47978 , n47979 , n47980 , n47981 , n47982 , n47983 , n47984 , n47985 , n47986 , n47987 , n47988 , n47989 , n47990 , n47991 , n47992 , n47993 , n47994 , n47995 , n47996 , n47997 , n47998 , n47999 , n48000 , n48001 , n48002 , n48003 , n48004 , n48005 , n48006 , n48007 , n48008 , n48009 , n48010 , n48011 , n48012 , n48013 , n48014 , n48015 , n48016 , n48017 , n48018 , n48019 , n48020 , n48021 , n48022 , n48023 , n48024 , n48025 , n48026 , n48027 , n48028 , n48029 , n48030 , n48031 , n48032 , n48033 , n48034 , n48035 , n48036 , n48037 , n48038 , n48039 , n48040 , n48041 , n48042 , n48043 , n48044 , n48045 , n48046 , n48047 , n48048 , n48049 , n48050 , n48051 , n48052 , n48053 , n48054 , n48055 , n48056 , n48057 , n48058 , n48059 , n48060 , n48061 , n48062 , n48063 , n48064 , n48065 , n48066 , n48067 , n48068 , n48069 , n48070 , n48071 , n48072 , n48073 , n48074 , n48075 , n48076 , n48077 , n48078 , n48079 , n48080 , n48081 , n48082 , n48083 , n48084 , n48085 , n48086 , n48087 , n48088 , n48089 , n48090 , n48091 , n48092 , n48093 , n48094 , n48095 , n48096 , n48097 , n48098 , n48099 , n48100 , n48101 , n48102 , n48103 , n48104 , n48105 , n48106 , n48107 , n48108 , n48109 , n48110 , n48111 , n48112 , n48113 , n48114 , n48115 , n48116 , n48117 , n48118 , n48119 , n48120 , n48121 , n48122 , n48123 , n48124 , n48125 , n48126 , n48127 , n48128 , n48129 , n48130 , n48131 , n48132 , n48133 , n48134 , n48135 , n48136 , n48137 , n48138 , n48139 , n48140 , n48141 , n48142 , n48143 , n48144 , n48145 , n48146 , n48147 , n48148 , n48149 , n48150 , n48151 , n48152 , n48153 , n48154 , n48155 , n48156 , n48157 , n48158 , n48159 , n48160 , n48161 , n48162 , n48163 , n48164 , n48165 , n48166 , n48167 , n48168 , n48169 , n48170 , n48171 , n48172 , n48173 , n48174 , n48175 , n48176 , n48177 , n48178 , n48179 , n48180 , n48181 , n48182 , n48183 , n48184 , n48185 , n48186 , n48187 , n48188 , n48189 , n48190 , n48191 , n48192 , n48193 , n48194 , n48195 , n48196 , n48197 , n48198 , n48199 , n48200 , n48201 , n48202 , n48203 , n48204 , n48205 , n48206 , n48207 , n48208 , n48209 , n48210 , n48211 , n48212 , n48213 , n48214 , n48215 , n48216 , n48217 , n48218 , n48219 , n48220 , n48221 , n48222 , n48223 , n48224 , n48225 , n48226 , n48227 , n48228 , n48229 , n48230 , n48231 , n48232 , n48233 , n48234 , n48235 , n48236 , n48237 , n48238 , n48239 , n48240 , n48241 , n48242 , n48243 , n48244 , n48245 , n48246 , n48247 , n48248 , n48249 , n48250 , n48251 , n48252 , n48253 , n48254 , n48255 , n48256 , n48257 , n48258 , n48259 , n48260 , n48261 , n48262 , n48263 , n48264 , n48265 , n48266 , n48267 , n48268 , n48269 , n48270 , n48271 , n48272 , n48273 , n48274 , n48275 , n48276 , n48277 , n48278 , n48279 , n48280 , n48281 , n48282 , n48283 , n48284 , n48285 , n48286 , n48287 , n48288 , n48289 , n48290 , n48291 , n48292 , n48293 , n48294 , n48295 , n48296 , n48297 , n48298 , n48299 , n48300 , n48301 , n48302 , n48303 , n48304 , n48305 , n48306 , n48307 , n48308 , n48309 , n48310 , n48311 , n48312 , n48313 , n48314 , n48315 , n48316 , n48317 , n48318 , n48319 , n48320 , n48321 , n48322 , n48323 , n48324 , n48325 , n48326 , n48327 , n48328 , n48329 , n48330 , n48331 , n48332 , n48333 , n48334 , n48335 , n48336 , n48337 , n48338 , n48339 , n48340 , n48341 , n48342 , n48343 , n48344 , n48345 , n48346 , n48347 , n48348 , n48349 , n48350 , n48351 , n48352 , n48353 , n48354 , n48355 , n48356 , n48357 , n48358 , n48359 , n48360 , n48361 , n48362 , n48363 , n48364 , n48365 , n48366 , n48367 , n48368 , n48369 , n48370 , n48371 , n48372 , n48373 , n48374 , n48375 , n48376 , n48377 , n48378 , n48379 , n48380 , n48381 , n48382 , n48383 , n48384 , n48385 , n48386 , n48387 , n48388 , n48389 , n48390 , n48391 , n48392 , n48393 , n48394 , n48395 , n48396 , n48397 , n48398 , n48399 , n48400 , n48401 , n48402 , n48403 , n48404 , n48405 , n48406 , n48407 , n48408 , n48409 , n48410 , n48411 , n48412 , n48413 , n48414 , n48415 , n48416 , n48417 , n48418 , n48419 , n48420 , n48421 , n48422 , n48423 , n48424 , n48425 , n48426 , n48427 , n48428 , n48429 , n48430 , n48431 , n48432 , n48433 , n48434 , n48435 , n48436 , n48437 , n48438 , n48439 , n48440 , n48441 , n48442 , n48443 , n48444 , n48445 , n48446 , n48447 , n48448 , n48449 , n48450 , n48451 , n48452 , n48453 , n48454 , n48455 , n48456 , n48457 , n48458 , n48459 , n48460 , n48461 , n48462 , n48463 , n48464 , n48465 , n48466 , n48467 , n48468 , n48469 , n48470 , n48471 , n48472 , n48473 , n48474 , n48475 , n48476 , n48477 , n48478 , n48479 , n48480 , n48481 , n48482 , n48483 , n48484 , n48485 , n48486 , n48487 , n48488 , n48489 , n48490 , n48491 , n48492 , n48493 , n48494 , n48495 , n48496 , n48497 , n48498 , n48499 , n48500 , n48501 , n48502 , n48503 , n48504 , n48505 , n48506 , n48507 , n48508 , n48509 , n48510 , n48511 , n48512 , n48513 , n48514 , n48515 , n48516 , n48517 , n48518 , n48519 , n48520 , n48521 , n48522 , n48523 , n48524 , n48525 , n48526 , n48527 , n48528 , n48529 , n48530 , n48531 , n48532 , n48533 , n48534 , n48535 , n48536 , n48537 , n48538 , n48539 , n48540 , n48541 , n48542 , n48543 , n48544 , n48545 , n48546 , n48547 , n48548 , n48549 , n48550 , n48551 , n48552 , n48553 , n48554 , n48555 , n48556 , n48557 , n48558 , n48559 , n48560 , n48561 , n48562 , n48563 , n48564 , n48565 , n48566 , n48567 , n48568 , n48569 , n48570 , n48571 , n48572 , n48573 , n48574 , n48575 , n48576 , n48577 , n48578 , n48579 , n48580 , n48581 , n48582 , n48583 , n48584 , n48585 , n48586 , n48587 , n48588 , n48589 , n48590 , n48591 , n48592 , n48593 , n48594 , n48595 , n48596 , n48597 , n48598 , n48599 , n48600 , n48601 , n48602 , n48603 , n48604 , n48605 , n48606 , n48607 , n48608 , n48609 , n48610 , n48611 , n48612 , n48613 , n48614 , n48615 , n48616 , n48617 , n48618 , n48619 , n48620 , n48621 , n48622 , n48623 , n48624 , n48625 , n48626 , n48627 , n48628 , n48629 , n48630 , n48631 , n48632 , n48633 , n48634 , n48635 , n48636 , n48637 , n48638 , n48639 , n48640 , n48641 , n48642 , n48643 , n48644 , n48645 , n48646 , n48647 , n48648 , n48649 , n48650 , n48651 , n48652 , n48653 , n48654 , n48655 , n48656 , n48657 , n48658 , n48659 , n48660 , n48661 , n48662 , n48663 , n48664 , n48665 , n48666 , n48667 , n48668 , n48669 , n48670 , n48671 , n48672 , n48673 , n48674 , n48675 , n48676 , n48677 , n48678 , n48679 , n48680 , n48681 , n48682 , n48683 , n48684 , n48685 , n48686 , n48687 , n48688 , n48689 , n48690 , n48691 , n48692 , n48693 , n48694 , n48695 , n48696 , n48697 , n48698 , n48699 , n48700 , n48701 , n48702 , n48703 , n48704 , n48705 , n48706 , n48707 , n48708 , n48709 , n48710 , n48711 , n48712 , n48713 , n48714 , n48715 , n48716 , n48717 , n48718 , n48719 , n48720 , n48721 , n48722 , n48723 , n48724 , n48725 , n48726 , n48727 , n48728 , n48729 , n48730 , n48731 , n48732 , n48733 , n48734 , n48735 , n48736 , n48737 , n48738 , n48739 , n48740 , n48741 , n48742 , n48743 , n48744 , n48745 , n48746 , n48747 , n48748 , n48749 , n48750 , n48751 , n48752 , n48753 , n48754 , n48755 , n48756 , n48757 , n48758 , n48759 , n48760 , n48761 , n48762 , n48763 , n48764 , n48765 , n48766 , n48767 , n48768 , n48769 , n48770 , n48771 , n48772 , n48773 , n48774 , n48775 , n48776 , n48777 , n48778 , n48779 , n48780 , n48781 , n48782 , n48783 , n48784 , n48785 , n48786 , n48787 , n48788 , n48789 , n48790 , n48791 , n48792 , n48793 , n48794 , n48795 , n48796 , n48797 , n48798 , n48799 , n48800 , n48801 , n48802 , n48803 , n48804 , n48805 , n48806 , n48807 , n48808 , n48809 , n48810 , n48811 , n48812 , n48813 , n48814 , n48815 , n48816 , n48817 , n48818 , n48819 , n48820 , n48821 , n48822 , n48823 , n48824 , n48825 , n48826 , n48827 , n48828 , n48829 , n48830 , n48831 , n48832 , n48833 , n48834 , n48835 , n48836 , n48837 , n48838 , n48839 , n48840 , n48841 , n48842 , n48843 , n48844 , n48845 , n48846 , n48847 , n48848 , n48849 , n48850 , n48851 , n48852 , n48853 , n48854 , n48855 , n48856 , n48857 , n48858 , n48859 , n48860 , n48861 , n48862 , n48863 , n48864 , n48865 , n48866 , n48867 , n48868 , n48869 , n48870 , n48871 , n48872 , n48873 , n48874 , n48875 , n48876 , n48877 , n48878 , n48879 , n48880 , n48881 , n48882 , n48883 , n48884 , n48885 , n48886 , n48887 , n48888 , n48889 , n48890 , n48891 , n48892 , n48893 , n48894 , n48895 , n48896 , n48897 , n48898 , n48899 , n48900 , n48901 , n48902 , n48903 , n48904 , n48905 , n48906 , n48907 , n48908 , n48909 , n48910 , n48911 , n48912 , n48913 , n48914 , n48915 , n48916 , n48917 , n48918 , n48919 , n48920 , n48921 , n48922 , n48923 , n48924 , n48925 , n48926 , n48927 , n48928 , n48929 , n48930 , n48931 , n48932 , n48933 , n48934 , n48935 , n48936 , n48937 , n48938 , n48939 , n48940 , n48941 , n48942 , n48943 , n48944 , n48945 , n48946 , n48947 , n48948 , n48949 , n48950 , n48951 , n48952 , n48953 , n48954 , n48955 , n48956 , n48957 , n48958 , n48959 , n48960 , n48961 , n48962 , n48963 , n48964 , n48965 , n48966 , n48967 , n48968 , n48969 , n48970 , n48971 , n48972 , n48973 , n48974 , n48975 , n48976 , n48977 , n48978 , n48979 , n48980 , n48981 , n48982 , n48983 , n48984 , n48985 , n48986 , n48987 , n48988 , n48989 , n48990 , n48991 , n48992 , n48993 , n48994 , n48995 , n48996 , n48997 , n48998 , n48999 , n49000 , n49001 , n49002 , n49003 , n49004 , n49005 , n49006 , n49007 , n49008 , n49009 , n49010 , n49011 , n49012 , n49013 , n49014 , n49015 , n49016 , n49017 , n49018 , n49019 , n49020 , n49021 , n49022 , n49023 , n49024 , n49025 , n49026 , n49027 , n49028 , n49029 , n49030 , n49031 , n49032 , n49033 , n49034 , n49035 , n49036 , n49037 , n49038 , n49039 , n49040 , n49041 , n49042 , n49043 , n49044 , n49045 , n49046 , n49047 , n49048 , n49049 , n49050 , n49051 , n49052 , n49053 , n49054 , n49055 , n49056 , n49057 , n49058 , n49059 , n49060 , n49061 , n49062 , n49063 , n49064 , n49065 , n49066 , n49067 , n49068 , n49069 , n49070 , n49071 , n49072 , n49073 , n49074 , n49075 , n49076 , n49077 , n49078 , n49079 , n49080 , n49081 , n49082 , n49083 , n49084 , n49085 , n49086 , n49087 , n49088 , n49089 , n49090 , n49091 , n49092 , n49093 , n49094 , n49095 , n49096 , n49097 , n49098 , n49099 , n49100 , n49101 , n49102 , n49103 , n49104 , n49105 , n49106 , n49107 , n49108 , n49109 , n49110 , n49111 , n49112 , n49113 , n49114 , n49115 , n49116 , n49117 , n49118 , n49119 , n49120 , n49121 , n49122 , n49123 , n49124 , n49125 , n49126 , n49127 , n49128 , n49129 , n49130 , n49131 , n49132 , n49133 , n49134 , n49135 , n49136 , n49137 , n49138 , n49139 , n49140 , n49141 , n49142 , n49143 , n49144 , n49145 , n49146 , n49147 , n49148 , n49149 , n49150 , n49151 , n49152 , n49153 , n49154 , n49155 , n49156 , n49157 , n49158 , n49159 , n49160 , n49161 , n49162 , n49163 , n49164 , n49165 , n49166 , n49167 , n49168 , n49169 , n49170 , n49171 , n49172 , n49173 , n49174 , n49175 , n49176 , n49177 , n49178 , n49179 , n49180 , n49181 , n49182 , n49183 , n49184 , n49185 , n49186 , n49187 , n49188 , n49189 , n49190 , n49191 , n49192 , n49193 , n49194 , n49195 , n49196 , n49197 , n49198 , n49199 , n49200 , n49201 , n49202 , n49203 , n49204 , n49205 , n49206 , n49207 , n49208 , n49209 , n49210 , n49211 , n49212 , n49213 , n49214 , n49215 , n49216 , n49217 , n49218 , n49219 , n49220 , n49221 , n49222 , n49223 , n49224 , n49225 , n49226 , n49227 , n49228 , n49229 , n49230 , n49231 , n49232 , n49233 , n49234 , n49235 , n49236 , n49237 , n49238 , n49239 , n49240 , n49241 , n49242 , n49243 , n49244 , n49245 , n49246 , n49247 , n49248 , n49249 , n49250 , n49251 , n49252 , n49253 , n49254 , n49255 , n49256 , n49257 , n49258 , n49259 , n49260 , n49261 , n49262 , n49263 , n49264 , n49265 , n49266 , n49267 , n49268 , n49269 , n49270 , n49271 , n49272 , n49273 , n49274 , n49275 , n49276 , n49277 , n49278 , n49279 , n49280 , n49281 , n49282 , n49283 , n49284 , n49285 , n49286 , n49287 , n49288 , n49289 , n49290 , n49291 , n49292 , n49293 , n49294 , n49295 , n49296 , n49297 , n49298 , n49299 , n49300 , n49301 , n49302 , n49303 , n49304 , n49305 , n49306 , n49307 , n49308 , n49309 , n49310 , n49311 , n49312 , n49313 , n49314 , n49315 , n49316 , n49317 , n49318 , n49319 , n49320 , n49321 , n49322 , n49323 , n49324 , n49325 , n49326 , n49327 , n49328 , n49329 , n49330 , n49331 , n49332 , n49333 , n49334 , n49335 , n49336 , n49337 , n49338 , n49339 , n49340 , n49341 , n49342 , n49343 , n49344 , n49345 , n49346 , n49347 , n49348 , n49349 , n49350 , n49351 , n49352 , n49353 , n49354 , n49355 , n49356 , n49357 , n49358 , n49359 , n49360 , n49361 , n49362 , n49363 , n49364 , n49365 , n49366 , n49367 , n49368 , n49369 , n49370 , n49371 , n49372 , n49373 , n49374 , n49375 , n49376 , n49377 , n49378 , n49379 , n49380 , n49381 , n49382 , n49383 , n49384 , n49385 , n49386 , n49387 , n49388 , n49389 , n49390 , n49391 , n49392 , n49393 , n49394 , n49395 , n49396 , n49397 , n49398 , n49399 , n49400 , n49401 , n49402 , n49403 , n49404 , n49405 , n49406 , n49407 , n49408 , n49409 , n49410 , n49411 , n49412 , n49413 , n49414 , n49415 , n49416 , n49417 , n49418 , n49419 , n49420 , n49421 , n49422 , n49423 , n49424 , n49425 , n49426 , n49427 , n49428 , n49429 , n49430 , n49431 , n49432 , n49433 , n49434 , n49435 , n49436 , n49437 , n49438 , n49439 , n49440 , n49441 , n49442 , n49443 , n49444 , n49445 , n49446 , n49447 , n49448 , n49449 , n49450 , n49451 , n49452 , n49453 , n49454 , n49455 , n49456 , n49457 , n49458 , n49459 , n49460 , n49461 , n49462 , n49463 , n49464 , n49465 , n49466 , n49467 , n49468 , n49469 , n49470 , n49471 , n49472 , n49473 , n49474 , n49475 , n49476 , n49477 , n49478 , n49479 , n49480 , n49481 , n49482 , n49483 , n49484 , n49485 , n49486 , n49487 , n49488 , n49489 , n49490 , n49491 , n49492 , n49493 , n49494 , n49495 , n49496 , n49497 , n49498 , n49499 , n49500 , n49501 , n49502 , n49503 , n49504 , n49505 , n49506 , n49507 , n49508 , n49509 , n49510 , n49511 , n49512 , n49513 , n49514 , n49515 , n49516 , n49517 , n49518 , n49519 , n49520 , n49521 , n49522 , n49523 , n49524 , n49525 , n49526 , n49527 , n49528 , n49529 , n49530 , n49531 , n49532 , n49533 , n49534 , n49535 , n49536 , n49537 , n49538 , n49539 , n49540 , n49541 , n49542 , n49543 , n49544 , n49545 , n49546 , n49547 , n49548 , n49549 , n49550 , n49551 , n49552 , n49553 , n49554 , n49555 , n49556 , n49557 , n49558 , n49559 , n49560 , n49561 , n49562 , n49563 , n49564 , n49565 , n49566 , n49567 , n49568 , n49569 , n49570 , n49571 , n49572 , n49573 , n49574 , n49575 , n49576 , n49577 , n49578 , n49579 , n49580 , n49581 , n49582 , n49583 , n49584 , n49585 , n49586 , n49587 , n49588 , n49589 , n49590 , n49591 , n49592 , n49593 , n49594 , n49595 , n49596 , n49597 , n49598 , n49599 , n49600 , n49601 , n49602 , n49603 , n49604 , n49605 , n49606 , n49607 , n49608 , n49609 , n49610 , n49611 , n49612 , n49613 , n49614 , n49615 , n49616 , n49617 , n49618 , n49619 , n49620 , n49621 , n49622 , n49623 , n49624 , n49625 , n49626 , n49627 , n49628 , n49629 , n49630 , n49631 , n49632 , n49633 , n49634 , n49635 , n49636 , n49637 , n49638 , n49639 , n49640 , n49641 , n49642 , n49643 , n49644 , n49645 , n49646 , n49647 , n49648 , n49649 , n49650 , n49651 , n49652 , n49653 , n49654 , n49655 , n49656 , n49657 , n49658 , n49659 , n49660 , n49661 , n49662 , n49663 , n49664 , n49665 , n49666 , n49667 , n49668 , n49669 , n49670 , n49671 , n49672 , n49673 , n49674 , n49675 , n49676 , n49677 , n49678 , n49679 , n49680 , n49681 , n49682 , n49683 , n49684 , n49685 , n49686 , n49687 , n49688 , n49689 , n49690 , n49691 , n49692 , n49693 , n49694 , n49695 , n49696 , n49697 , n49698 , n49699 , n49700 , n49701 , n49702 , n49703 , n49704 , n49705 , n49706 , n49707 , n49708 , n49709 , n49710 , n49711 , n49712 , n49713 , n49714 , n49715 , n49716 , n49717 , n49718 , n49719 , n49720 , n49721 , n49722 , n49723 , n49724 , n49725 , n49726 , n49727 , n49728 , n49729 , n49730 , n49731 , n49732 , n49733 , n49734 , n49735 , n49736 , n49737 , n49738 , n49739 , n49740 , n49741 , n49742 , n49743 , n49744 , n49745 , n49746 , n49747 , n49748 , n49749 , n49750 , n49751 , n49752 , n49753 , n49754 , n49755 , n49756 , n49757 , n49758 , n49759 , n49760 , n49761 , n49762 , n49763 , n49764 , n49765 , n49766 , n49767 , n49768 , n49769 , n49770 , n49771 , n49772 , n49773 , n49774 , n49775 , n49776 , n49777 , n49778 , n49779 , n49780 , n49781 , n49782 , n49783 , n49784 , n49785 , n49786 , n49787 , n49788 , n49789 , n49790 , n49791 , n49792 , n49793 , n49794 , n49795 , n49796 , n49797 , n49798 , n49799 , n49800 , n49801 , n49802 , n49803 , n49804 , n49805 , n49806 , n49807 , n49808 , n49809 , n49810 , n49811 , n49812 , n49813 , n49814 , n49815 , n49816 , n49817 , n49818 , n49819 , n49820 , n49821 , n49822 , n49823 , n49824 , n49825 , n49826 , n49827 , n49828 , n49829 , n49830 , n49831 , n49832 , n49833 , n49834 , n49835 , n49836 , n49837 , n49838 , n49839 , n49840 , n49841 , n49842 , n49843 , n49844 , n49845 , n49846 , n49847 , n49848 , n49849 , n49850 , n49851 , n49852 , n49853 , n49854 , n49855 , n49856 , n49857 , n49858 , n49859 , n49860 , n49861 , n49862 , n49863 , n49864 , n49865 , n49866 , n49867 , n49868 , n49869 , n49870 , n49871 , n49872 , n49873 , n49874 , n49875 , n49876 , n49877 , n49878 , n49879 , n49880 , n49881 , n49882 , n49883 , n49884 , n49885 , n49886 , n49887 , n49888 , n49889 , n49890 , n49891 , n49892 , n49893 , n49894 , n49895 , n49896 , n49897 , n49898 , n49899 , n49900 , n49901 , n49902 , n49903 , n49904 , n49905 , n49906 , n49907 , n49908 , n49909 , n49910 , n49911 , n49912 , n49913 , n49914 , n49915 , n49916 , n49917 , n49918 , n49919 , n49920 , n49921 , n49922 , n49923 , n49924 , n49925 , n49926 , n49927 , n49928 , n49929 , n49930 , n49931 , n49932 , n49933 , n49934 , n49935 , n49936 , n49937 , n49938 , n49939 , n49940 , n49941 , n49942 , n49943 , n49944 , n49945 , n49946 , n49947 , n49948 , n49949 , n49950 , n49951 , n49952 , n49953 , n49954 , n49955 , n49956 , n49957 , n49958 , n49959 , n49960 , n49961 , n49962 , n49963 , n49964 , n49965 , n49966 , n49967 , n49968 , n49969 , n49970 , n49971 , n49972 , n49973 , n49974 , n49975 , n49976 , n49977 , n49978 , n49979 , n49980 , n49981 , n49982 , n49983 , n49984 , n49985 , n49986 , n49987 , n49988 , n49989 , n49990 , n49991 , n49992 , n49993 , n49994 , n49995 , n49996 , n49997 , n49998 , n49999 , n50000 , n50001 , n50002 , n50003 , n50004 , n50005 , n50006 , n50007 , n50008 , n50009 , n50010 , n50011 , n50012 , n50013 , n50014 , n50015 , n50016 , n50017 , n50018 , n50019 , n50020 , n50021 , n50022 , n50023 , n50024 , n50025 , n50026 , n50027 , n50028 , n50029 , n50030 , n50031 , n50032 , n50033 , n50034 , n50035 , n50036 , n50037 , n50038 , n50039 , n50040 , n50041 , n50042 , n50043 , n50044 , n50045 , n50046 , n50047 , n50048 , n50049 , n50050 , n50051 , n50052 , n50053 , n50054 , n50055 , n50056 , n50057 , n50058 , n50059 , n50060 , n50061 , n50062 , n50063 , n50064 , n50065 , n50066 , n50067 , n50068 , n50069 , n50070 , n50071 , n50072 , n50073 , n50074 , n50075 , n50076 , n50077 , n50078 , n50079 , n50080 , n50081 , n50082 , n50083 , n50084 , n50085 , n50086 , n50087 , n50088 , n50089 , n50090 , n50091 , n50092 , n50093 , n50094 , n50095 , n50096 , n50097 , n50098 , n50099 , n50100 , n50101 , n50102 , n50103 , n50104 , n50105 , n50106 , n50107 , n50108 , n50109 , n50110 , n50111 , n50112 , n50113 , n50114 , n50115 , n50116 , n50117 , n50118 , n50119 , n50120 , n50121 , n50122 , n50123 , n50124 , n50125 , n50126 , n50127 , n50128 , n50129 , n50130 , n50131 , n50132 , n50133 , n50134 , n50135 , n50136 , n50137 , n50138 , n50139 , n50140 , n50141 , n50142 , n50143 , n50144 , n50145 , n50146 , n50147 , n50148 , n50149 , n50150 , n50151 , n50152 , n50153 , n50154 , n50155 , n50156 , n50157 , n50158 , n50159 , n50160 , n50161 , n50162 , n50163 , n50164 , n50165 , n50166 , n50167 , n50168 , n50169 , n50170 , n50171 , n50172 , n50173 , n50174 , n50175 , n50176 , n50177 , n50178 , n50179 , n50180 , n50181 , n50182 , n50183 , n50184 , n50185 , n50186 , n50187 , n50188 , n50189 , n50190 , n50191 , n50192 , n50193 , n50194 , n50195 , n50196 , n50197 , n50198 , n50199 , n50200 , n50201 , n50202 , n50203 , n50204 , n50205 , n50206 , n50207 , n50208 , n50209 , n50210 , n50211 , n50212 , n50213 , n50214 , n50215 , n50216 , n50217 , n50218 , n50219 , n50220 , n50221 , n50222 , n50223 , n50224 , n50225 , n50226 , n50227 , n50228 , n50229 , n50230 , n50231 , n50232 , n50233 , n50234 , n50235 , n50236 , n50237 , n50238 , n50239 , n50240 , n50241 , n50242 , n50243 , n50244 , n50245 , n50246 , n50247 , n50248 , n50249 , n50250 , n50251 , n50252 , n50253 , n50254 , n50255 , n50256 , n50257 , n50258 , n50259 , n50260 , n50261 , n50262 , n50263 , n50264 , n50265 , n50266 , n50267 , n50268 , n50269 , n50270 , n50271 , n50272 , n50273 , n50274 , n50275 , n50276 , n50277 , n50278 , n50279 , n50280 , n50281 , n50282 , n50283 , n50284 , n50285 , n50286 , n50287 , n50288 , n50289 , n50290 , n50291 , n50292 , n50293 , n50294 , n50295 , n50296 , n50297 , n50298 , n50299 , n50300 , n50301 , n50302 , n50303 , n50304 , n50305 , n50306 , n50307 , n50308 , n50309 , n50310 , n50311 , n50312 , n50313 , n50314 , n50315 , n50316 , n50317 , n50318 , n50319 , n50320 , n50321 , n50322 , n50323 , n50324 , n50325 , n50326 , n50327 , n50328 , n50329 , n50330 , n50331 , n50332 , n50333 , n50334 , n50335 , n50336 , n50337 , n50338 , n50339 , n50340 , n50341 , n50342 , n50343 , n50344 , n50345 , n50346 , n50347 , n50348 , n50349 , n50350 , n50351 , n50352 , n50353 , n50354 , n50355 , n50356 , n50357 , n50358 , n50359 , n50360 , n50361 , n50362 , n50363 , n50364 , n50365 , n50366 , n50367 , n50368 , n50369 , n50370 , n50371 , n50372 , n50373 , n50374 , n50375 , n50376 , n50377 , n50378 , n50379 , n50380 , n50381 , n50382 , n50383 , n50384 , n50385 , n50386 , n50387 , n50388 , n50389 , n50390 , n50391 , n50392 , n50393 , n50394 , n50395 , n50396 , n50397 , n50398 , n50399 , n50400 , n50401 , n50402 , n50403 , n50404 , n50405 , n50406 , n50407 , n50408 , n50409 , n50410 , n50411 , n50412 , n50413 , n50414 , n50415 , n50416 , n50417 , n50418 , n50419 , n50420 , n50421 , n50422 , n50423 , n50424 , n50425 , n50426 , n50427 , n50428 , n50429 , n50430 , n50431 , n50432 , n50433 , n50434 , n50435 , n50436 , n50437 , n50438 , n50439 , n50440 , n50441 , n50442 , n50443 , n50444 , n50445 , n50446 , n50447 , n50448 , n50449 , n50450 , n50451 , n50452 , n50453 , n50454 , n50455 , n50456 , n50457 , n50458 , n50459 , n50460 , n50461 , n50462 , n50463 , n50464 , n50465 , n50466 , n50467 , n50468 , n50469 , n50470 , n50471 , n50472 , n50473 , n50474 , n50475 , n50476 , n50477 , n50478 , n50479 , n50480 , n50481 , n50482 , n50483 , n50484 , n50485 , n50486 , n50487 , n50488 , n50489 , n50490 , n50491 , n50492 , n50493 , n50494 , n50495 , n50496 , n50497 , n50498 , n50499 , n50500 , n50501 , n50502 , n50503 , n50504 , n50505 , n50506 , n50507 , n50508 , n50509 , n50510 , n50511 , n50512 , n50513 , n50514 , n50515 , n50516 , n50517 , n50518 , n50519 , n50520 , n50521 , n50522 , n50523 , n50524 , n50525 , n50526 , n50527 , n50528 , n50529 , n50530 , n50531 , n50532 , n50533 , n50534 , n50535 , n50536 , n50537 , n50538 , n50539 , n50540 , n50541 , n50542 , n50543 , n50544 , n50545 , n50546 , n50547 , n50548 , n50549 , n50550 , n50551 , n50552 , n50553 , n50554 , n50555 , n50556 , n50557 , n50558 , n50559 , n50560 , n50561 , n50562 , n50563 , n50564 , n50565 , n50566 , n50567 , n50568 , n50569 , n50570 , n50571 , n50572 , n50573 , n50574 , n50575 , n50576 , n50577 , n50578 , n50579 , n50580 , n50581 , n50582 , n50583 , n50584 , n50585 , n50586 , n50587 , n50588 , n50589 , n50590 , n50591 , n50592 , n50593 , n50594 , n50595 , n50596 , n50597 , n50598 , n50599 , n50600 , n50601 , n50602 , n50603 , n50604 , n50605 , n50606 , n50607 , n50608 , n50609 , n50610 , n50611 , n50612 , n50613 , n50614 , n50615 , n50616 , n50617 , n50618 , n50619 , n50620 , n50621 , n50622 , n50623 , n50624 , n50625 , n50626 , n50627 , n50628 , n50629 , n50630 , n50631 , n50632 , n50633 , n50634 , n50635 , n50636 , n50637 , n50638 , n50639 , n50640 , n50641 , n50642 , n50643 , n50644 , n50645 , n50646 , n50647 , n50648 , n50649 , n50650 , n50651 , n50652 , n50653 , n50654 , n50655 , n50656 , n50657 , n50658 , n50659 , n50660 , n50661 , n50662 , n50663 , n50664 , n50665 , n50666 , n50667 , n50668 , n50669 , n50670 , n50671 , n50672 , n50673 , n50674 , n50675 , n50676 , n50677 , n50678 , n50679 , n50680 , n50681 , n50682 , n50683 , n50684 , n50685 , n50686 , n50687 , n50688 , n50689 , n50690 , n50691 , n50692 , n50693 , n50694 , n50695 , n50696 , n50697 , n50698 , n50699 , n50700 , n50701 , n50702 , n50703 , n50704 , n50705 , n50706 , n50707 , n50708 , n50709 , n50710 , n50711 , n50712 , n50713 , n50714 , n50715 , n50716 , n50717 , n50718 , n50719 , n50720 , n50721 , n50722 , n50723 , n50724 , n50725 , n50726 , n50727 , n50728 , n50729 , n50730 , n50731 , n50732 , n50733 , n50734 , n50735 , n50736 , n50737 , n50738 , n50739 , n50740 , n50741 , n50742 , n50743 , n50744 , n50745 , n50746 , n50747 , n50748 , n50749 , n50750 , n50751 , n50752 , n50753 , n50754 , n50755 , n50756 , n50757 , n50758 , n50759 , n50760 , n50761 , n50762 , n50763 , n50764 , n50765 , n50766 , n50767 , n50768 , n50769 , n50770 , n50771 , n50772 , n50773 , n50774 , n50775 , n50776 , n50777 , n50778 , n50779 , n50780 , n50781 , n50782 , n50783 , n50784 , n50785 , n50786 , n50787 , n50788 , n50789 , n50790 , n50791 , n50792 , n50793 , n50794 , n50795 , n50796 , n50797 , n50798 , n50799 , n50800 , n50801 , n50802 , n50803 , n50804 , n50805 , n50806 , n50807 , n50808 , n50809 , n50810 , n50811 , n50812 , n50813 , n50814 , n50815 , n50816 , n50817 , n50818 , n50819 , n50820 , n50821 , n50822 , n50823 , n50824 , n50825 , n50826 , n50827 , n50828 , n50829 , n50830 , n50831 , n50832 , n50833 , n50834 , n50835 , n50836 , n50837 , n50838 , n50839 , n50840 , n50841 , n50842 , n50843 , n50844 , n50845 , n50846 , n50847 , n50848 , n50849 , n50850 , n50851 , n50852 , n50853 , n50854 , n50855 , n50856 , n50857 , n50858 , n50859 , n50860 , n50861 , n50862 , n50863 , n50864 , n50865 , n50866 , n50867 , n50868 , n50869 , n50870 , n50871 , n50872 , n50873 , n50874 , n50875 , n50876 , n50877 , n50878 , n50879 , n50880 , n50881 , n50882 , n50883 , n50884 , n50885 , n50886 , n50887 , n50888 , n50889 , n50890 , n50891 , n50892 , n50893 , n50894 , n50895 , n50896 , n50897 , n50898 , n50899 , n50900 , n50901 , n50902 , n50903 , n50904 , n50905 , n50906 , n50907 , n50908 , n50909 , n50910 , n50911 , n50912 , n50913 , n50914 , n50915 , n50916 , n50917 , n50918 , n50919 , n50920 , n50921 , n50922 , n50923 , n50924 , n50925 , n50926 , n50927 , n50928 , n50929 , n50930 , n50931 , n50932 , n50933 , n50934 , n50935 , n50936 , n50937 , n50938 , n50939 , n50940 , n50941 , n50942 , n50943 , n50944 , n50945 , n50946 , n50947 , n50948 , n50949 , n50950 , n50951 , n50952 , n50953 , n50954 , n50955 , n50956 , n50957 , n50958 , n50959 , n50960 , n50961 , n50962 , n50963 , n50964 , n50965 , n50966 , n50967 , n50968 , n50969 , n50970 , n50971 , n50972 , n50973 , n50974 , n50975 , n50976 , n50977 , n50978 , n50979 , n50980 , n50981 , n50982 , n50983 , n50984 , n50985 , n50986 , n50987 , n50988 , n50989 , n50990 , n50991 , n50992 , n50993 , n50994 , n50995 , n50996 , n50997 , n50998 , n50999 , n51000 , n51001 , n51002 , n51003 , n51004 , n51005 , n51006 , n51007 , n51008 , n51009 , n51010 , n51011 , n51012 , n51013 , n51014 , n51015 , n51016 , n51017 , n51018 , n51019 , n51020 , n51021 , n51022 , n51023 , n51024 , n51025 , n51026 , n51027 , n51028 , n51029 , n51030 , n51031 , n51032 , n51033 , n51034 , n51035 , n51036 , n51037 , n51038 , n51039 , n51040 , n51041 , n51042 , n51043 , n51044 , n51045 , n51046 , n51047 , n51048 , n51049 , n51050 , n51051 , n51052 , n51053 , n51054 , n51055 , n51056 , n51057 , n51058 , n51059 , n51060 , n51061 , n51062 , n51063 , n51064 , n51065 , n51066 , n51067 , n51068 , n51069 , n51070 , n51071 , n51072 , n51073 , n51074 , n51075 , n51076 , n51077 , n51078 , n51079 , n51080 , n51081 , n51082 , n51083 , n51084 , n51085 , n51086 , n51087 , n51088 , n51089 , n51090 , n51091 , n51092 , n51093 , n51094 , n51095 , n51096 , n51097 , n51098 , n51099 , n51100 , n51101 , n51102 , n51103 , n51104 , n51105 , n51106 , n51107 , n51108 , n51109 , n51110 , n51111 , n51112 , n51113 , n51114 , n51115 , n51116 , n51117 , n51118 , n51119 , n51120 , n51121 , n51122 , n51123 , n51124 , n51125 , n51126 , n51127 , n51128 , n51129 , n51130 , n51131 , n51132 , n51133 , n51134 , n51135 , n51136 , n51137 , n51138 , n51139 , n51140 , n51141 , n51142 , n51143 , n51144 , n51145 , n51146 , n51147 , n51148 , n51149 , n51150 , n51151 , n51152 , n51153 , n51154 , n51155 , n51156 , n51157 , n51158 , n51159 , n51160 , n51161 , n51162 , n51163 , n51164 , n51165 , n51166 , n51167 , n51168 , n51169 , n51170 , n51171 , n51172 , n51173 , n51174 , n51175 , n51176 , n51177 , n51178 , n51179 , n51180 , n51181 , n51182 , n51183 , n51184 , n51185 , n51186 , n51187 , n51188 , n51189 , n51190 , n51191 , n51192 , n51193 , n51194 , n51195 , n51196 , n51197 , n51198 , n51199 , n51200 , n51201 , n51202 , n51203 , n51204 , n51205 , n51206 , n51207 , n51208 , n51209 , n51210 , n51211 , n51212 , n51213 , n51214 , n51215 , n51216 , n51217 , n51218 , n51219 , n51220 , n51221 , n51222 , n51223 , n51224 , n51225 , n51226 , n51227 , n51228 , n51229 , n51230 , n51231 , n51232 , n51233 , n51234 , n51235 , n51236 , n51237 , n51238 , n51239 , n51240 , n51241 , n51242 , n51243 , n51244 , n51245 , n51246 , n51247 , n51248 , n51249 , n51250 , n51251 , n51252 , n51253 , n51254 , n51255 , n51256 , n51257 , n51258 , n51259 , n51260 , n51261 , n51262 , n51263 , n51264 , n51265 , n51266 , n51267 , n51268 , n51269 , n51270 , n51271 , n51272 , n51273 , n51274 , n51275 , n51276 , n51277 , n51278 , n51279 , n51280 , n51281 , n51282 , n51283 , n51284 , n51285 , n51286 , n51287 , n51288 , n51289 , n51290 , n51291 , n51292 , n51293 , n51294 , n51295 , n51296 , n51297 , n51298 , n51299 , n51300 , n51301 , n51302 , n51303 , n51304 , n51305 , n51306 , n51307 , n51308 , n51309 , n51310 , n51311 , n51312 , n51313 , n51314 , n51315 , n51316 , n51317 , n51318 , n51319 , n51320 , n51321 , n51322 , n51323 , n51324 , n51325 , n51326 , n51327 , n51328 , n51329 , n51330 , n51331 , n51332 , n51333 , n51334 , n51335 , n51336 , n51337 , n51338 , n51339 , n51340 , n51341 , n51342 , n51343 , n51344 , n51345 , n51346 , n51347 , n51348 , n51349 , n51350 , n51351 , n51352 , n51353 , n51354 , n51355 , n51356 , n51357 , n51358 , n51359 , n51360 , n51361 , n51362 , n51363 , n51364 , n51365 , n51366 , n51367 , n51368 , n51369 , n51370 , n51371 , n51372 , n51373 , n51374 , n51375 , n51376 , n51377 , n51378 , n51379 , n51380 , n51381 , n51382 , n51383 , n51384 , n51385 , n51386 , n51387 , n51388 , n51389 , n51390 , n51391 , n51392 , n51393 , n51394 , n51395 , n51396 , n51397 , n51398 , n51399 , n51400 , n51401 , n51402 , n51403 , n51404 , n51405 , n51406 , n51407 , n51408 , n51409 , n51410 , n51411 , n51412 , n51413 , n51414 , n51415 , n51416 , n51417 , n51418 , n51419 , n51420 , n51421 , n51422 , n51423 , n51424 , n51425 , n51426 , n51427 , n51428 , n51429 , n51430 , n51431 , n51432 , n51433 , n51434 , n51435 , n51436 , n51437 , n51438 , n51439 , n51440 , n51441 , n51442 , n51443 , n51444 , n51445 , n51446 , n51447 , n51448 , n51449 , n51450 , n51451 , n51452 , n51453 , n51454 , n51455 , n51456 , n51457 , n51458 , n51459 , n51460 , n51461 , n51462 , n51463 , n51464 , n51465 , n51466 , n51467 , n51468 , n51469 , n51470 , n51471 , n51472 , n51473 , n51474 , n51475 , n51476 , n51477 , n51478 , n51479 , n51480 , n51481 , n51482 , n51483 , n51484 , n51485 , n51486 , n51487 , n51488 , n51489 , n51490 , n51491 , n51492 , n51493 , n51494 , n51495 , n51496 , n51497 , n51498 , n51499 , n51500 , n51501 , n51502 , n51503 , n51504 , n51505 , n51506 , n51507 , n51508 , n51509 , n51510 , n51511 , n51512 , n51513 , n51514 , n51515 , n51516 , n51517 , n51518 , n51519 , n51520 , n51521 , n51522 , n51523 , n51524 , n51525 , n51526 , n51527 , n51528 , n51529 , n51530 , n51531 , n51532 , n51533 , n51534 , n51535 , n51536 , n51537 , n51538 , n51539 , n51540 , n51541 , n51542 , n51543 , n51544 , n51545 , n51546 , n51547 , n51548 , n51549 , n51550 , n51551 , n51552 , n51553 , n51554 , n51555 , n51556 , n51557 , n51558 , n51559 , n51560 , n51561 , n51562 , n51563 , n51564 , n51565 , n51566 , n51567 , n51568 , n51569 , n51570 , n51571 , n51572 , n51573 , n51574 , n51575 , n51576 , n51577 , n51578 , n51579 , n51580 , n51581 , n51582 , n51583 , n51584 , n51585 , n51586 , n51587 , n51588 , n51589 , n51590 , n51591 , n51592 , n51593 , n51594 , n51595 , n51596 , n51597 , n51598 , n51599 , n51600 , n51601 , n51602 , n51603 , n51604 , n51605 , n51606 , n51607 , n51608 , n51609 , n51610 , n51611 , n51612 , n51613 , n51614 , n51615 , n51616 , n51617 , n51618 , n51619 , n51620 , n51621 , n51622 , n51623 , n51624 , n51625 , n51626 , n51627 , n51628 , n51629 , n51630 , n51631 , n51632 , n51633 , n51634 , n51635 , n51636 , n51637 , n51638 , n51639 , n51640 , n51641 , n51642 , n51643 , n51644 , n51645 , n51646 , n51647 , n51648 , n51649 , n51650 , n51651 , n51652 , n51653 , n51654 , n51655 , n51656 , n51657 , n51658 , n51659 , n51660 , n51661 , n51662 , n51663 , n51664 , n51665 , n51666 , n51667 , n51668 , n51669 , n51670 , n51671 , n51672 , n51673 , n51674 , n51675 , n51676 , n51677 , n51678 , n51679 , n51680 , n51681 , n51682 , n51683 , n51684 , n51685 , n51686 , n51687 , n51688 , n51689 , n51690 , n51691 , n51692 , n51693 , n51694 , n51695 , n51696 , n51697 , n51698 , n51699 , n51700 , n51701 , n51702 , n51703 , n51704 , n51705 , n51706 , n51707 , n51708 , n51709 , n51710 , n51711 , n51712 , n51713 , n51714 , n51715 , n51716 , n51717 , n51718 , n51719 , n51720 , n51721 , n51722 , n51723 , n51724 , n51725 , n51726 , n51727 , n51728 , n51729 , n51730 , n51731 , n51732 , n51733 , n51734 , n51735 , n51736 , n51737 , n51738 , n51739 , n51740 , n51741 , n51742 , n51743 , n51744 , n51745 , n51746 , n51747 , n51748 , n51749 , n51750 , n51751 , n51752 , n51753 , n51754 , n51755 , n51756 , n51757 , n51758 , n51759 , n51760 , n51761 , n51762 , n51763 , n51764 , n51765 , n51766 , n51767 , n51768 , n51769 , n51770 , n51771 , n51772 , n51773 , n51774 , n51775 , n51776 , n51777 , n51778 , n51779 , n51780 , n51781 , n51782 , n51783 , n51784 , n51785 , n51786 , n51787 , n51788 , n51789 , n51790 , n51791 , n51792 , n51793 , n51794 , n51795 , n51796 , n51797 , n51798 , n51799 , n51800 , n51801 , n51802 , n51803 , n51804 , n51805 , n51806 , n51807 , n51808 , n51809 , n51810 , n51811 , n51812 , n51813 , n51814 , n51815 , n51816 , n51817 , n51818 , n51819 , n51820 , n51821 , n51822 , n51823 , n51824 , n51825 , n51826 , n51827 , n51828 , n51829 , n51830 , n51831 , n51832 , n51833 , n51834 , n51835 , n51836 , n51837 , n51838 , n51839 , n51840 , n51841 , n51842 , n51843 , n51844 , n51845 , n51846 , n51847 , n51848 , n51849 , n51850 , n51851 , n51852 , n51853 , n51854 , n51855 , n51856 , n51857 , n51858 , n51859 , n51860 , n51861 , n51862 , n51863 , n51864 , n51865 , n51866 , n51867 , n51868 , n51869 , n51870 , n51871 , n51872 , n51873 , n51874 , n51875 , n51876 , n51877 , n51878 , n51879 , n51880 , n51881 , n51882 , n51883 , n51884 , n51885 , n51886 , n51887 , n51888 , n51889 , n51890 , n51891 , n51892 , n51893 , n51894 , n51895 , n51896 , n51897 , n51898 , n51899 , n51900 , n51901 , n51902 , n51903 , n51904 , n51905 , n51906 , n51907 , n51908 , n51909 , n51910 , n51911 , n51912 , n51913 , n51914 , n51915 , n51916 , n51917 , n51918 , n51919 , n51920 , n51921 , n51922 , n51923 , n51924 , n51925 , n51926 , n51927 , n51928 , n51929 , n51930 , n51931 , n51932 , n51933 , n51934 , n51935 , n51936 , n51937 , n51938 , n51939 , n51940 , n51941 , n51942 , n51943 , n51944 , n51945 , n51946 , n51947 , n51948 , n51949 , n51950 , n51951 , n51952 , n51953 , n51954 , n51955 , n51956 , n51957 , n51958 , n51959 , n51960 , n51961 , n51962 , n51963 , n51964 , n51965 , n51966 , n51967 , n51968 , n51969 , n51970 , n51971 , n51972 , n51973 , n51974 , n51975 , n51976 , n51977 , n51978 , n51979 , n51980 , n51981 , n51982 , n51983 , n51984 , n51985 , n51986 , n51987 , n51988 , n51989 , n51990 , n51991 , n51992 , n51993 , n51994 , n51995 , n51996 , n51997 , n51998 , n51999 , n52000 , n52001 , n52002 , n52003 , n52004 , n52005 , n52006 , n52007 , n52008 , n52009 , n52010 , n52011 , n52012 , n52013 , n52014 , n52015 , n52016 , n52017 , n52018 , n52019 , n52020 , n52021 , n52022 , n52023 , n52024 , n52025 , n52026 , n52027 , n52028 , n52029 , n52030 , n52031 , n52032 , n52033 , n52034 , n52035 , n52036 , n52037 , n52038 , n52039 , n52040 , n52041 , n52042 , n52043 , n52044 , n52045 , n52046 , n52047 , n52048 , n52049 , n52050 , n52051 , n52052 , n52053 , n52054 , n52055 , n52056 , n52057 , n52058 , n52059 , n52060 , n52061 , n52062 , n52063 , n52064 , n52065 , n52066 , n52067 , n52068 , n52069 , n52070 , n52071 , n52072 , n52073 , n52074 , n52075 , n52076 , n52077 , n52078 , n52079 , n52080 , n52081 , n52082 , n52083 , n52084 , n52085 , n52086 , n52087 , n52088 , n52089 , n52090 , n52091 , n52092 , n52093 , n52094 , n52095 , n52096 , n52097 , n52098 , n52099 , n52100 , n52101 , n52102 , n52103 , n52104 , n52105 , n52106 , n52107 , n52108 , n52109 , n52110 , n52111 , n52112 , n52113 , n52114 , n52115 , n52116 , n52117 , n52118 , n52119 , n52120 , n52121 , n52122 , n52123 , n52124 , n52125 , n52126 , n52127 , n52128 , n52129 , n52130 , n52131 , n52132 , n52133 , n52134 , n52135 , n52136 , n52137 , n52138 , n52139 , n52140 , n52141 , n52142 , n52143 , n52144 , n52145 , n52146 , n52147 , n52148 , n52149 , n52150 , n52151 , n52152 , n52153 , n52154 , n52155 , n52156 , n52157 , n52158 , n52159 , n52160 , n52161 , n52162 , n52163 , n52164 , n52165 , n52166 , n52167 , n52168 , n52169 , n52170 , n52171 , n52172 , n52173 , n52174 , n52175 , n52176 , n52177 , n52178 , n52179 , n52180 , n52181 , n52182 , n52183 , n52184 , n52185 , n52186 , n52187 , n52188 , n52189 , n52190 , n52191 , n52192 , n52193 , n52194 , n52195 , n52196 , n52197 , n52198 , n52199 , n52200 , n52201 , n52202 , n52203 , n52204 , n52205 , n52206 , n52207 , n52208 , n52209 , n52210 , n52211 , n52212 , n52213 , n52214 , n52215 , n52216 , n52217 , n52218 , n52219 , n52220 , n52221 , n52222 , n52223 , n52224 , n52225 , n52226 , n52227 , n52228 , n52229 , n52230 , n52231 , n52232 , n52233 , n52234 , n52235 , n52236 , n52237 , n52238 , n52239 , n52240 , n52241 , n52242 , n52243 , n52244 , n52245 , n52246 , n52247 , n52248 , n52249 , n52250 , n52251 , n52252 , n52253 , n52254 , n52255 , n52256 , n52257 , n52258 , n52259 , n52260 , n52261 , n52262 , n52263 , n52264 , n52265 , n52266 , n52267 , n52268 , n52269 , n52270 , n52271 , n52272 , n52273 , n52274 , n52275 , n52276 , n52277 , n52278 , n52279 , n52280 , n52281 , n52282 , n52283 , n52284 , n52285 , n52286 , n52287 , n52288 , n52289 , n52290 , n52291 , n52292 , n52293 , n52294 , n52295 , n52296 , n52297 , n52298 , n52299 , n52300 , n52301 , n52302 , n52303 , n52304 , n52305 , n52306 , n52307 , n52308 , n52309 , n52310 , n52311 , n52312 , n52313 , n52314 , n52315 , n52316 , n52317 , n52318 , n52319 , n52320 , n52321 , n52322 , n52323 , n52324 , n52325 , n52326 , n52327 , n52328 , n52329 , n52330 , n52331 , n52332 , n52333 , n52334 , n52335 , n52336 , n52337 , n52338 , n52339 , n52340 , n52341 , n52342 , n52343 , n52344 , n52345 , n52346 , n52347 , n52348 , n52349 , n52350 , n52351 , n52352 , n52353 , n52354 , n52355 , n52356 , n52357 , n52358 , n52359 , n52360 , n52361 , n52362 , n52363 , n52364 , n52365 , n52366 , n52367 , n52368 , n52369 , n52370 , n52371 , n52372 , n52373 , n52374 , n52375 , n52376 , n52377 , n52378 , n52379 , n52380 , n52381 , n52382 , n52383 , n52384 , n52385 , n52386 , n52387 , n52388 , n52389 , n52390 , n52391 , n52392 , n52393 , n52394 , n52395 , n52396 , n52397 , n52398 , n52399 , n52400 , n52401 , n52402 , n52403 , n52404 , n52405 , n52406 , n52407 , n52408 , n52409 , n52410 , n52411 , n52412 , n52413 , n52414 , n52415 , n52416 , n52417 , n52418 , n52419 , n52420 , n52421 , n52422 , n52423 , n52424 , n52425 , n52426 , n52427 , n52428 , n52429 , n52430 , n52431 , n52432 , n52433 , n52434 , n52435 , n52436 , n52437 , n52438 , n52439 , n52440 , n52441 , n52442 , n52443 , n52444 , n52445 , n52446 , n52447 , n52448 , n52449 , n52450 , n52451 , n52452 , n52453 , n52454 , n52455 , n52456 , n52457 , n52458 , n52459 , n52460 , n52461 , n52462 , n52463 , n52464 , n52465 , n52466 , n52467 , n52468 , n52469 , n52470 , n52471 , n52472 , n52473 , n52474 , n52475 , n52476 , n52477 , n52478 , n52479 , n52480 , n52481 , n52482 , n52483 , n52484 , n52485 , n52486 , n52487 , n52488 , n52489 , n52490 , n52491 , n52492 , n52493 , n52494 , n52495 , n52496 , n52497 , n52498 , n52499 , n52500 , n52501 , n52502 , n52503 , n52504 , n52505 , n52506 , n52507 , n52508 , n52509 , n52510 , n52511 , n52512 , n52513 , n52514 , n52515 , n52516 , n52517 , n52518 , n52519 , n52520 , n52521 , n52522 , n52523 , n52524 , n52525 , n52526 , n52527 , n52528 , n52529 , n52530 , n52531 , n52532 , n52533 , n52534 , n52535 , n52536 , n52537 , n52538 , n52539 , n52540 , n52541 , n52542 , n52543 , n52544 , n52545 , n52546 , n52547 , n52548 , n52549 , n52550 , n52551 , n52552 , n52553 , n52554 , n52555 , n52556 , n52557 , n52558 , n52559 , n52560 , n52561 , n52562 , n52563 , n52564 , n52565 , n52566 , n52567 , n52568 , n52569 , n52570 , n52571 , n52572 , n52573 , n52574 , n52575 , n52576 , n52577 , n52578 , n52579 , n52580 , n52581 , n52582 , n52583 , n52584 , n52585 , n52586 , n52587 , n52588 , n52589 , n52590 , n52591 , n52592 , n52593 , n52594 , n52595 , n52596 , n52597 , n52598 , n52599 , n52600 , n52601 , n52602 , n52603 , n52604 , n52605 , n52606 , n52607 , n52608 , n52609 , n52610 , n52611 , n52612 , n52613 , n52614 , n52615 , n52616 , n52617 , n52618 , n52619 , n52620 , n52621 , n52622 , n52623 , n52624 , n52625 , n52626 , n52627 , n52628 , n52629 , n52630 , n52631 , n52632 , n52633 , n52634 , n52635 , n52636 , n52637 , n52638 , n52639 , n52640 , n52641 , n52642 , n52643 , n52644 , n52645 , n52646 , n52647 , n52648 , n52649 , n52650 , n52651 , n52652 , n52653 , n52654 , n52655 , n52656 , n52657 , n52658 , n52659 , n52660 , n52661 , n52662 , n52663 , n52664 , n52665 , n52666 , n52667 , n52668 , n52669 , n52670 , n52671 , n52672 , n52673 , n52674 , n52675 , n52676 , n52677 , n52678 , n52679 , n52680 , n52681 , n52682 , n52683 , n52684 , n52685 , n52686 , n52687 , n52688 , n52689 , n52690 , n52691 , n52692 , n52693 , n52694 , n52695 , n52696 , n52697 , n52698 , n52699 , n52700 , n52701 , n52702 , n52703 , n52704 , n52705 , n52706 , n52707 , n52708 , n52709 , n52710 , n52711 , n52712 , n52713 , n52714 , n52715 , n52716 , n52717 , n52718 , n52719 , n52720 , n52721 , n52722 , n52723 , n52724 , n52725 , n52726 , n52727 , n52728 , n52729 , n52730 , n52731 , n52732 , n52733 , n52734 , n52735 , n52736 , n52737 , n52738 , n52739 , n52740 , n52741 , n52742 , n52743 , n52744 , n52745 , n52746 , n52747 , n52748 , n52749 , n52750 , n52751 , n52752 , n52753 , n52754 , n52755 , n52756 , n52757 , n52758 , n52759 , n52760 , n52761 , n52762 , n52763 , n52764 , n52765 , n52766 , n52767 , n52768 , n52769 , n52770 , n52771 , n52772 , n52773 , n52774 , n52775 , n52776 , n52777 , n52778 , n52779 , n52780 , n52781 , n52782 , n52783 , n52784 , n52785 , n52786 , n52787 , n52788 , n52789 , n52790 , n52791 , n52792 , n52793 , n52794 , n52795 , n52796 , n52797 , n52798 , n52799 , n52800 , n52801 , n52802 , n52803 , n52804 , n52805 , n52806 , n52807 , n52808 , n52809 , n52810 , n52811 , n52812 , n52813 , n52814 , n52815 , n52816 , n52817 , n52818 , n52819 , n52820 , n52821 , n52822 , n52823 , n52824 , n52825 , n52826 , n52827 , n52828 , n52829 , n52830 , n52831 , n52832 , n52833 , n52834 , n52835 , n52836 , n52837 , n52838 , n52839 , n52840 , n52841 , n52842 , n52843 , n52844 , n52845 , n52846 , n52847 , n52848 , n52849 , n52850 , n52851 , n52852 , n52853 , n52854 , n52855 , n52856 , n52857 , n52858 , n52859 , n52860 , n52861 , n52862 , n52863 , n52864 , n52865 , n52866 , n52867 , n52868 , n52869 , n52870 , n52871 , n52872 , n52873 , n52874 , n52875 , n52876 , n52877 , n52878 , n52879 , n52880 , n52881 , n52882 , n52883 , n52884 , n52885 , n52886 , n52887 , n52888 , n52889 , n52890 , n52891 , n52892 , n52893 , n52894 , n52895 , n52896 , n52897 , n52898 , n52899 , n52900 , n52901 , n52902 , n52903 , n52904 , n52905 , n52906 , n52907 , n52908 , n52909 , n52910 , n52911 , n52912 , n52913 , n52914 , n52915 , n52916 , n52917 , n52918 , n52919 , n52920 , n52921 , n52922 , n52923 , n52924 , n52925 , n52926 , n52927 , n52928 , n52929 , n52930 , n52931 , n52932 , n52933 , n52934 , n52935 , n52936 , n52937 , n52938 , n52939 , n52940 , n52941 , n52942 , n52943 , n52944 , n52945 , n52946 , n52947 , n52948 , n52949 , n52950 , n52951 , n52952 , n52953 , n52954 , n52955 , n52956 , n52957 , n52958 , n52959 , n52960 , n52961 , n52962 , n52963 , n52964 , n52965 , n52966 , n52967 , n52968 , n52969 , n52970 , n52971 , n52972 , n52973 , n52974 , n52975 , n52976 , n52977 , n52978 , n52979 , n52980 , n52981 , n52982 , n52983 , n52984 , n52985 , n52986 , n52987 , n52988 , n52989 , n52990 , n52991 , n52992 , n52993 , n52994 , n52995 , n52996 , n52997 , n52998 , n52999 , n53000 , n53001 , n53002 , n53003 , n53004 , n53005 , n53006 , n53007 , n53008 , n53009 , n53010 , n53011 , n53012 , n53013 , n53014 , n53015 , n53016 , n53017 , n53018 , n53019 , n53020 , n53021 , n53022 , n53023 , n53024 , n53025 , n53026 , n53027 , n53028 , n53029 , n53030 , n53031 , n53032 , n53033 , n53034 , n53035 , n53036 , n53037 , n53038 , n53039 , n53040 , n53041 , n53042 , n53043 , n53044 , n53045 , n53046 , n53047 , n53048 , n53049 , n53050 , n53051 , n53052 , n53053 , n53054 , n53055 , n53056 , n53057 , n53058 , n53059 , n53060 , n53061 , n53062 , n53063 , n53064 , n53065 , n53066 , n53067 , n53068 , n53069 , n53070 , n53071 , n53072 , n53073 , n53074 , n53075 , n53076 , n53077 , n53078 , n53079 , n53080 , n53081 , n53082 , n53083 , n53084 , n53085 , n53086 , n53087 , n53088 , n53089 , n53090 , n53091 , n53092 , n53093 , n53094 , n53095 , n53096 , n53097 , n53098 , n53099 , n53100 , n53101 , n53102 , n53103 , n53104 , n53105 , n53106 , n53107 , n53108 , n53109 , n53110 , n53111 , n53112 , n53113 , n53114 , n53115 , n53116 , n53117 , n53118 , n53119 , n53120 , n53121 , n53122 , n53123 , n53124 , n53125 , n53126 , n53127 , n53128 , n53129 , n53130 , n53131 , n53132 , n53133 , n53134 , n53135 , n53136 , n53137 , n53138 , n53139 , n53140 , n53141 , n53142 , n53143 , n53144 , n53145 , n53146 , n53147 , n53148 , n53149 , n53150 , n53151 , n53152 , n53153 , n53154 , n53155 , n53156 , n53157 , n53158 , n53159 , n53160 , n53161 , n53162 , n53163 , n53164 , n53165 , n53166 , n53167 , n53168 , n53169 , n53170 , n53171 , n53172 , n53173 , n53174 , n53175 , n53176 , n53177 , n53178 , n53179 , n53180 , n53181 , n53182 , n53183 , n53184 , n53185 , n53186 , n53187 , n53188 , n53189 , n53190 , n53191 , n53192 , n53193 , n53194 , n53195 , n53196 , n53197 , n53198 , n53199 , n53200 , n53201 , n53202 , n53203 , n53204 , n53205 , n53206 , n53207 , n53208 , n53209 , n53210 , n53211 , n53212 , n53213 , n53214 , n53215 , n53216 , n53217 , n53218 , n53219 , n53220 , n53221 , n53222 , n53223 , n53224 , n53225 , n53226 , n53227 , n53228 , n53229 , n53230 , n53231 , n53232 , n53233 , n53234 , n53235 , n53236 , n53237 , n53238 , n53239 , n53240 , n53241 , n53242 , n53243 , n53244 , n53245 , n53246 , n53247 , n53248 , n53249 , n53250 , n53251 , n53252 , n53253 , n53254 , n53255 , n53256 , n53257 , n53258 , n53259 , n53260 , n53261 , n53262 , n53263 , n53264 , n53265 , n53266 , n53267 , n53268 , n53269 , n53270 , n53271 , n53272 , n53273 , n53274 , n53275 , n53276 , n53277 , n53278 , n53279 , n53280 , n53281 , n53282 , n53283 , n53284 , n53285 , n53286 , n53287 , n53288 , n53289 , n53290 , n53291 , n53292 , n53293 , n53294 , n53295 , n53296 , n53297 , n53298 , n53299 , n53300 , n53301 , n53302 , n53303 , n53304 , n53305 , n53306 , n53307 , n53308 , n53309 , n53310 , n53311 , n53312 , n53313 , n53314 , n53315 , n53316 , n53317 , n53318 , n53319 , n53320 , n53321 , n53322 , n53323 , n53324 , n53325 , n53326 , n53327 , n53328 , n53329 , n53330 , n53331 , n53332 , n53333 , n53334 , n53335 , n53336 , n53337 , n53338 , n53339 , n53340 , n53341 , n53342 , n53343 , n53344 , n53345 , n53346 , n53347 , n53348 , n53349 , n53350 , n53351 , n53352 , n53353 , n53354 , n53355 , n53356 , n53357 , n53358 , n53359 , n53360 , n53361 , n53362 , n53363 , n53364 , n53365 , n53366 , n53367 , n53368 , n53369 , n53370 , n53371 , n53372 , n53373 , n53374 , n53375 , n53376 , n53377 , n53378 , n53379 , n53380 , n53381 , n53382 , n53383 , n53384 , n53385 , n53386 , n53387 , n53388 , n53389 , n53390 , n53391 , n53392 , n53393 , n53394 , n53395 , n53396 , n53397 , n53398 , n53399 , n53400 , n53401 , n53402 , n53403 , n53404 , n53405 , n53406 , n53407 , n53408 , n53409 , n53410 , n53411 , n53412 , n53413 , n53414 , n53415 , n53416 , n53417 , n53418 , n53419 , n53420 , n53421 , n53422 , n53423 , n53424 , n53425 , n53426 , n53427 , n53428 , n53429 , n53430 , n53431 , n53432 , n53433 , n53434 , n53435 , n53436 , n53437 , n53438 , n53439 , n53440 , n53441 , n53442 , n53443 , n53444 , n53445 , n53446 , n53447 , n53448 , n53449 , n53450 , n53451 , n53452 , n53453 , n53454 , n53455 , n53456 , n53457 , n53458 , n53459 , n53460 , n53461 , n53462 , n53463 , n53464 , n53465 , n53466 , n53467 , n53468 , n53469 , n53470 , n53471 , n53472 , n53473 , n53474 , n53475 , n53476 , n53477 , n53478 , n53479 , n53480 , n53481 , n53482 , n53483 , n53484 , n53485 , n53486 , n53487 , n53488 , n53489 , n53490 , n53491 , n53492 , n53493 , n53494 , n53495 , n53496 , n53497 , n53498 , n53499 , n53500 , n53501 , n53502 , n53503 , n53504 , n53505 , n53506 , n53507 , n53508 , n53509 , n53510 , n53511 , n53512 , n53513 , n53514 , n53515 , n53516 , n53517 , n53518 , n53519 , n53520 , n53521 , n53522 , n53523 , n53524 , n53525 , n53526 , n53527 , n53528 , n53529 , n53530 , n53531 , n53532 , n53533 , n53534 , n53535 , n53536 , n53537 , n53538 , n53539 , n53540 , n53541 , n53542 , n53543 , n53544 , n53545 , n53546 , n53547 , n53548 , n53549 , n53550 , n53551 , n53552 , n53553 , n53554 , n53555 , n53556 , n53557 , n53558 , n53559 , n53560 , n53561 , n53562 , n53563 , n53564 , n53565 , n53566 , n53567 , n53568 , n53569 , n53570 , n53571 , n53572 , n53573 , n53574 , n53575 , n53576 , n53577 , n53578 , n53579 , n53580 , n53581 , n53582 , n53583 , n53584 , n53585 , n53586 , n53587 , n53588 , n53589 , n53590 , n53591 , n53592 , n53593 , n53594 , n53595 , n53596 , n53597 , n53598 , n53599 , n53600 , n53601 , n53602 , n53603 , n53604 , n53605 , n53606 , n53607 , n53608 , n53609 , n53610 , n53611 , n53612 , n53613 , n53614 , n53615 , n53616 , n53617 , n53618 , n53619 , n53620 , n53621 , n53622 , n53623 , n53624 , n53625 , n53626 , n53627 , n53628 , n53629 , n53630 , n53631 , n53632 , n53633 , n53634 , n53635 , n53636 , n53637 , n53638 , n53639 , n53640 , n53641 , n53642 , n53643 , n53644 , n53645 , n53646 , n53647 , n53648 , n53649 , n53650 , n53651 , n53652 , n53653 , n53654 , n53655 , n53656 , n53657 , n53658 , n53659 , n53660 , n53661 , n53662 , n53663 , n53664 , n53665 , n53666 , n53667 , n53668 , n53669 , n53670 , n53671 , n53672 , n53673 , n53674 , n53675 , n53676 , n53677 , n53678 , n53679 , n53680 , n53681 , n53682 , n53683 , n53684 , n53685 , n53686 , n53687 , n53688 , n53689 , n53690 , n53691 , n53692 , n53693 , n53694 , n53695 , n53696 , n53697 , n53698 , n53699 , n53700 , n53701 , n53702 , n53703 , n53704 , n53705 , n53706 , n53707 , n53708 , n53709 , n53710 , n53711 , n53712 , n53713 , n53714 , n53715 , n53716 , n53717 , n53718 , n53719 , n53720 , n53721 , n53722 , n53723 , n53724 , n53725 , n53726 , n53727 , n53728 , n53729 , n53730 , n53731 , n53732 , n53733 , n53734 , n53735 , n53736 , n53737 , n53738 , n53739 , n53740 , n53741 , n53742 , n53743 , n53744 , n53745 , n53746 , n53747 , n53748 , n53749 , n53750 , n53751 , n53752 , n53753 , n53754 , n53755 , n53756 , n53757 , n53758 , n53759 , n53760 , n53761 , n53762 , n53763 , n53764 , n53765 , n53766 , n53767 , n53768 , n53769 , n53770 , n53771 , n53772 , n53773 , n53774 , n53775 , n53776 , n53777 , n53778 , n53779 , n53780 , n53781 , n53782 , n53783 , n53784 , n53785 , n53786 , n53787 , n53788 , n53789 , n53790 , n53791 , n53792 , n53793 , n53794 , n53795 , n53796 , n53797 , n53798 , n53799 , n53800 , n53801 , n53802 , n53803 , n53804 , n53805 , n53806 , n53807 , n53808 , n53809 , n53810 , n53811 , n53812 , n53813 , n53814 , n53815 , n53816 , n53817 , n53818 , n53819 , n53820 , n53821 , n53822 , n53823 , n53824 , n53825 , n53826 , n53827 , n53828 , n53829 , n53830 , n53831 , n53832 , n53833 , n53834 , n53835 , n53836 , n53837 , n53838 , n53839 , n53840 , n53841 , n53842 , n53843 , n53844 , n53845 , n53846 , n53847 , n53848 , n53849 , n53850 , n53851 , n53852 , n53853 , n53854 , n53855 , n53856 , n53857 , n53858 , n53859 , n53860 , n53861 , n53862 , n53863 , n53864 , n53865 , n53866 , n53867 , n53868 , n53869 , n53870 , n53871 , n53872 , n53873 , n53874 , n53875 , n53876 , n53877 , n53878 , n53879 , n53880 , n53881 , n53882 , n53883 , n53884 , n53885 , n53886 , n53887 , n53888 , n53889 , n53890 , n53891 , n53892 , n53893 , n53894 , n53895 , n53896 , n53897 , n53898 , n53899 , n53900 , n53901 , n53902 , n53903 , n53904 , n53905 , n53906 , n53907 , n53908 , n53909 , n53910 , n53911 , n53912 , n53913 , n53914 , n53915 , n53916 , n53917 , n53918 , n53919 , n53920 , n53921 , n53922 , n53923 , n53924 , n53925 , n53926 , n53927 , n53928 , n53929 , n53930 , n53931 , n53932 , n53933 , n53934 , n53935 , n53936 , n53937 , n53938 , n53939 , n53940 , n53941 , n53942 , n53943 , n53944 , n53945 , n53946 , n53947 , n53948 , n53949 , n53950 , n53951 , n53952 , n53953 , n53954 , n53955 , n53956 , n53957 , n53958 , n53959 , n53960 , n53961 , n53962 , n53963 , n53964 , n53965 , n53966 , n53967 , n53968 , n53969 , n53970 , n53971 , n53972 , n53973 , n53974 , n53975 , n53976 , n53977 , n53978 , n53979 , n53980 , n53981 , n53982 , n53983 , n53984 , n53985 , n53986 , n53987 , n53988 , n53989 , n53990 , n53991 , n53992 , n53993 , n53994 , n53995 , n53996 , n53997 , n53998 , n53999 , n54000 , n54001 , n54002 , n54003 , n54004 , n54005 , n54006 , n54007 , n54008 , n54009 , n54010 , n54011 , n54012 , n54013 , n54014 , n54015 , n54016 , n54017 , n54018 , n54019 , n54020 , n54021 , n54022 , n54023 , n54024 , n54025 , n54026 , n54027 , n54028 , n54029 , n54030 , n54031 , n54032 , n54033 , n54034 , n54035 , n54036 , n54037 , n54038 , n54039 , n54040 , n54041 , n54042 , n54043 , n54044 , n54045 , n54046 , n54047 , n54048 , n54049 , n54050 , n54051 , n54052 , n54053 , n54054 , n54055 , n54056 , n54057 , n54058 , n54059 , n54060 , n54061 , n54062 , n54063 , n54064 , n54065 , n54066 , n54067 , n54068 , n54069 , n54070 , n54071 , n54072 , n54073 , n54074 , n54075 , n54076 , n54077 , n54078 , n54079 , n54080 , n54081 , n54082 , n54083 , n54084 , n54085 , n54086 , n54087 , n54088 , n54089 , n54090 , n54091 , n54092 , n54093 , n54094 , n54095 , n54096 , n54097 , n54098 , n54099 , n54100 , n54101 , n54102 , n54103 , n54104 , n54105 , n54106 , n54107 , n54108 , n54109 , n54110 , n54111 , n54112 , n54113 , n54114 , n54115 , n54116 , n54117 , n54118 , n54119 , n54120 , n54121 , n54122 , n54123 , n54124 , n54125 , n54126 , n54127 , n54128 , n54129 , n54130 , n54131 , n54132 , n54133 , n54134 , n54135 , n54136 , n54137 , n54138 , n54139 , n54140 , n54141 , n54142 , n54143 , n54144 , n54145 , n54146 , n54147 , n54148 , n54149 , n54150 , n54151 , n54152 , n54153 , n54154 , n54155 , n54156 , n54157 , n54158 , n54159 , n54160 , n54161 , n54162 , n54163 , n54164 , n54165 , n54166 , n54167 , n54168 , n54169 , n54170 , n54171 , n54172 , n54173 , n54174 , n54175 , n54176 , n54177 , n54178 , n54179 , n54180 , n54181 , n54182 , n54183 , n54184 , n54185 , n54186 , n54187 , n54188 , n54189 , n54190 , n54191 , n54192 , n54193 , n54194 , n54195 , n54196 , n54197 , n54198 , n54199 , n54200 , n54201 , n54202 , n54203 , n54204 , n54205 , n54206 , n54207 , n54208 , n54209 , n54210 , n54211 , n54212 , n54213 , n54214 , n54215 , n54216 , n54217 , n54218 , n54219 , n54220 , n54221 , n54222 , n54223 , n54224 , n54225 , n54226 , n54227 , n54228 , n54229 , n54230 , n54231 , n54232 , n54233 , n54234 , n54235 , n54236 , n54237 , n54238 , n54239 , n54240 , n54241 , n54242 , n54243 , n54244 , n54245 , n54246 , n54247 , n54248 , n54249 , n54250 , n54251 , n54252 , n54253 , n54254 , n54255 , n54256 , n54257 , n54258 , n54259 , n54260 , n54261 , n54262 , n54263 , n54264 , n54265 , n54266 , n54267 , n54268 , n54269 , n54270 , n54271 , n54272 , n54273 , n54274 , n54275 , n54276 , n54277 , n54278 , n54279 , n54280 , n54281 , n54282 , n54283 , n54284 , n54285 , n54286 , n54287 , n54288 , n54289 , n54290 , n54291 , n54292 , n54293 , n54294 , n54295 , n54296 , n54297 , n54298 , n54299 , n54300 , n54301 , n54302 , n54303 , n54304 , n54305 , n54306 , n54307 , n54308 , n54309 , n54310 , n54311 , n54312 , n54313 , n54314 , n54315 , n54316 , n54317 , n54318 , n54319 , n54320 , n54321 , n54322 , n54323 , n54324 , n54325 , n54326 , n54327 , n54328 , n54329 , n54330 , n54331 , n54332 , n54333 , n54334 , n54335 , n54336 , n54337 , n54338 , n54339 , n54340 , n54341 , n54342 , n54343 , n54344 , n54345 , n54346 , n54347 , n54348 , n54349 , n54350 , n54351 , n54352 , n54353 , n54354 , n54355 , n54356 , n54357 , n54358 , n54359 , n54360 , n54361 , n54362 , n54363 , n54364 , n54365 , n54366 , n54367 , n54368 , n54369 , n54370 , n54371 , n54372 , n54373 , n54374 , n54375 , n54376 , n54377 , n54378 , n54379 , n54380 , n54381 , n54382 , n54383 , n54384 , n54385 , n54386 , n54387 , n54388 , n54389 , n54390 , n54391 , n54392 , n54393 , n54394 , n54395 , n54396 , n54397 , n54398 , n54399 , n54400 , n54401 , n54402 , n54403 , n54404 , n54405 , n54406 , n54407 , n54408 , n54409 , n54410 , n54411 , n54412 , n54413 , n54414 , n54415 , n54416 , n54417 , n54418 , n54419 , n54420 , n54421 , n54422 , n54423 , n54424 , n54425 , n54426 , n54427 , n54428 , n54429 , n54430 , n54431 , n54432 , n54433 , n54434 , n54435 , n54436 , n54437 , n54438 , n54439 , n54440 , n54441 , n54442 , n54443 , n54444 , n54445 , n54446 , n54447 , n54448 , n54449 , n54450 , n54451 , n54452 , n54453 , n54454 , n54455 , n54456 , n54457 , n54458 , n54459 , n54460 , n54461 , n54462 , n54463 , n54464 , n54465 , n54466 , n54467 , n54468 , n54469 , n54470 , n54471 , n54472 , n54473 , n54474 , n54475 , n54476 , n54477 , n54478 , n54479 , n54480 , n54481 , n54482 , n54483 , n54484 , n54485 , n54486 , n54487 , n54488 , n54489 , n54490 , n54491 , n54492 , n54493 , n54494 , n54495 , n54496 , n54497 , n54498 , n54499 , n54500 , n54501 , n54502 , n54503 , n54504 , n54505 , n54506 , n54507 , n54508 , n54509 , n54510 , n54511 , n54512 , n54513 , n54514 , n54515 , n54516 , n54517 , n54518 , n54519 , n54520 , n54521 , n54522 , n54523 , n54524 , n54525 , n54526 , n54527 , n54528 , n54529 , n54530 , n54531 , n54532 , n54533 , n54534 , n54535 , n54536 , n54537 , n54538 , n54539 , n54540 , n54541 , n54542 , n54543 , n54544 , n54545 , n54546 , n54547 , n54548 , n54549 , n54550 , n54551 , n54552 , n54553 , n54554 , n54555 , n54556 , n54557 , n54558 , n54559 , n54560 , n54561 , n54562 , n54563 , n54564 , n54565 , n54566 , n54567 , n54568 , n54569 , n54570 , n54571 , n54572 , n54573 , n54574 , n54575 , n54576 , n54577 , n54578 , n54579 , n54580 , n54581 , n54582 , n54583 , n54584 , n54585 , n54586 , n54587 , n54588 , n54589 , n54590 , n54591 , n54592 , n54593 , n54594 , n54595 , n54596 , n54597 , n54598 , n54599 , n54600 , n54601 , n54602 , n54603 , n54604 , n54605 , n54606 , n54607 , n54608 , n54609 , n54610 , n54611 , n54612 , n54613 , n54614 , n54615 , n54616 , n54617 , n54618 , n54619 , n54620 , n54621 , n54622 , n54623 , n54624 , n54625 , n54626 , n54627 , n54628 , n54629 , n54630 , n54631 , n54632 , n54633 , n54634 , n54635 , n54636 , n54637 , n54638 , n54639 , n54640 , n54641 , n54642 , n54643 , n54644 , n54645 , n54646 , n54647 , n54648 , n54649 , n54650 , n54651 , n54652 , n54653 , n54654 , n54655 , n54656 , n54657 , n54658 , n54659 , n54660 , n54661 , n54662 , n54663 , n54664 , n54665 , n54666 , n54667 , n54668 , n54669 , n54670 , n54671 , n54672 , n54673 , n54674 , n54675 , n54676 , n54677 , n54678 , n54679 , n54680 , n54681 , n54682 , n54683 , n54684 , n54685 , n54686 , n54687 , n54688 , n54689 , n54690 , n54691 , n54692 , n54693 , n54694 , n54695 , n54696 , n54697 , n54698 , n54699 , n54700 , n54701 , n54702 , n54703 , n54704 , n54705 , n54706 , n54707 , n54708 , n54709 , n54710 , n54711 , n54712 , n54713 , n54714 , n54715 , n54716 , n54717 , n54718 , n54719 , n54720 , n54721 , n54722 , n54723 , n54724 , n54725 , n54726 , n54727 , n54728 , n54729 , n54730 , n54731 , n54732 , n54733 , n54734 , n54735 , n54736 , n54737 , n54738 , n54739 , n54740 , n54741 , n54742 , n54743 , n54744 , n54745 , n54746 , n54747 , n54748 , n54749 , n54750 , n54751 , n54752 , n54753 , n54754 , n54755 , n54756 , n54757 , n54758 , n54759 , n54760 , n54761 , n54762 , n54763 , n54764 , n54765 , n54766 , n54767 , n54768 , n54769 , n54770 , n54771 , n54772 , n54773 , n54774 , n54775 , n54776 , n54777 , n54778 , n54779 , n54780 , n54781 , n54782 , n54783 , n54784 , n54785 , n54786 , n54787 , n54788 , n54789 , n54790 , n54791 , n54792 , n54793 , n54794 , n54795 , n54796 , n54797 , n54798 , n54799 , n54800 , n54801 , n54802 , n54803 , n54804 , n54805 , n54806 , n54807 , n54808 , n54809 , n54810 , n54811 , n54812 , n54813 , n54814 , n54815 , n54816 , n54817 , n54818 , n54819 , n54820 , n54821 , n54822 , n54823 , n54824 , n54825 , n54826 , n54827 , n54828 , n54829 , n54830 , n54831 , n54832 , n54833 , n54834 , n54835 , n54836 , n54837 , n54838 , n54839 , n54840 , n54841 , n54842 , n54843 , n54844 , n54845 , n54846 , n54847 , n54848 , n54849 , n54850 , n54851 , n54852 , n54853 , n54854 , n54855 , n54856 , n54857 , n54858 , n54859 , n54860 , n54861 , n54862 , n54863 , n54864 , n54865 , n54866 , n54867 , n54868 , n54869 , n54870 , n54871 , n54872 , n54873 , n54874 , n54875 , n54876 , n54877 , n54878 , n54879 , n54880 , n54881 , n54882 , n54883 , n54884 , n54885 , n54886 , n54887 , n54888 , n54889 , n54890 , n54891 , n54892 , n54893 , n54894 , n54895 , n54896 , n54897 , n54898 , n54899 , n54900 , n54901 , n54902 , n54903 , n54904 , n54905 , n54906 , n54907 , n54908 , n54909 , n54910 , n54911 , n54912 , n54913 , n54914 , n54915 , n54916 , n54917 , n54918 , n54919 , n54920 , n54921 , n54922 , n54923 , n54924 , n54925 , n54926 , n54927 , n54928 , n54929 , n54930 , n54931 , n54932 , n54933 , n54934 , n54935 , n54936 , n54937 , n54938 , n54939 , n54940 , n54941 , n54942 , n54943 , n54944 , n54945 , n54946 , n54947 , n54948 , n54949 , n54950 , n54951 , n54952 , n54953 , n54954 , n54955 , n54956 , n54957 , n54958 , n54959 , n54960 , n54961 , n54962 , n54963 , n54964 , n54965 , n54966 , n54967 , n54968 , n54969 , n54970 , n54971 , n54972 , n54973 , n54974 , n54975 , n54976 , n54977 , n54978 , n54979 , n54980 , n54981 , n54982 , n54983 , n54984 , n54985 , n54986 , n54987 , n54988 , n54989 , n54990 , n54991 , n54992 , n54993 , n54994 , n54995 , n54996 , n54997 , n54998 , n54999 , n55000 , n55001 , n55002 , n55003 , n55004 , n55005 , n55006 , n55007 , n55008 , n55009 , n55010 , n55011 , n55012 , n55013 , n55014 , n55015 , n55016 , n55017 , n55018 , n55019 , n55020 , n55021 , n55022 , n55023 , n55024 , n55025 , n55026 , n55027 , n55028 , n55029 , n55030 , n55031 , n55032 , n55033 , n55034 , n55035 , n55036 , n55037 , n55038 , n55039 , n55040 , n55041 , n55042 , n55043 , n55044 , n55045 , n55046 , n55047 , n55048 , n55049 , n55050 , n55051 , n55052 , n55053 , n55054 , n55055 , n55056 , n55057 , n55058 , n55059 , n55060 , n55061 , n55062 , n55063 , n55064 , n55065 , n55066 , n55067 , n55068 , n55069 , n55070 , n55071 , n55072 , n55073 , n55074 , n55075 , n55076 , n55077 , n55078 , n55079 , n55080 , n55081 , n55082 , n55083 , n55084 , n55085 , n55086 , n55087 , n55088 , n55089 , n55090 , n55091 , n55092 , n55093 , n55094 , n55095 , n55096 , n55097 , n55098 , n55099 , n55100 , n55101 , n55102 , n55103 , n55104 , n55105 , n55106 , n55107 , n55108 , n55109 , n55110 , n55111 , n55112 , n55113 , n55114 , n55115 , n55116 , n55117 , n55118 , n55119 , n55120 , n55121 , n55122 , n55123 , n55124 , n55125 , n55126 , n55127 , n55128 , n55129 , n55130 , n55131 , n55132 , n55133 , n55134 , n55135 , n55136 , n55137 , n55138 , n55139 , n55140 , n55141 , n55142 , n55143 , n55144 , n55145 , n55146 , n55147 , n55148 , n55149 , n55150 , n55151 , n55152 , n55153 , n55154 , n55155 , n55156 , n55157 , n55158 , n55159 , n55160 , n55161 , n55162 , n55163 , n55164 , n55165 , n55166 , n55167 , n55168 , n55169 , n55170 , n55171 , n55172 , n55173 , n55174 , n55175 , n55176 , n55177 , n55178 , n55179 , n55180 , n55181 , n55182 , n55183 , n55184 , n55185 , n55186 , n55187 , n55188 , n55189 , n55190 , n55191 , n55192 , n55193 , n55194 , n55195 , n55196 , n55197 , n55198 , n55199 , n55200 , n55201 , n55202 , n55203 , n55204 , n55205 , n55206 , n55207 , n55208 , n55209 , n55210 , n55211 , n55212 , n55213 , n55214 , n55215 , n55216 , n55217 , n55218 , n55219 , n55220 , n55221 , n55222 , n55223 , n55224 , n55225 , n55226 , n55227 , n55228 , n55229 , n55230 , n55231 , n55232 , n55233 , n55234 , n55235 , n55236 , n55237 , n55238 , n55239 , n55240 , n55241 , n55242 , n55243 , n55244 , n55245 , n55246 , n55247 , n55248 , n55249 , n55250 , n55251 , n55252 , n55253 , n55254 , n55255 , n55256 , n55257 , n55258 , n55259 , n55260 , n55261 , n55262 , n55263 , n55264 , n55265 , n55266 , n55267 , n55268 , n55269 , n55270 , n55271 , n55272 , n55273 , n55274 , n55275 , n55276 , n55277 , n55278 , n55279 , n55280 , n55281 , n55282 , n55283 , n55284 , n55285 , n55286 , n55287 , n55288 , n55289 , n55290 , n55291 , n55292 , n55293 , n55294 , n55295 , n55296 , n55297 , n55298 , n55299 , n55300 , n55301 , n55302 , n55303 , n55304 , n55305 , n55306 , n55307 , n55308 , n55309 , n55310 , n55311 , n55312 , n55313 , n55314 , n55315 , n55316 , n55317 , n55318 , n55319 , n55320 , n55321 , n55322 , n55323 , n55324 , n55325 , n55326 , n55327 , n55328 , n55329 , n55330 , n55331 , n55332 , n55333 , n55334 , n55335 , n55336 , n55337 , n55338 , n55339 , n55340 , n55341 , n55342 , n55343 , n55344 , n55345 , n55346 , n55347 , n55348 , n55349 , n55350 , n55351 , n55352 , n55353 , n55354 , n55355 , n55356 , n55357 , n55358 , n55359 , n55360 , n55361 , n55362 , n55363 , n55364 , n55365 , n55366 , n55367 , n55368 , n55369 , n55370 , n55371 , n55372 , n55373 , n55374 , n55375 , n55376 , n55377 , n55378 , n55379 , n55380 , n55381 , n55382 , n55383 , n55384 , n55385 , n55386 , n55387 , n55388 , n55389 , n55390 , n55391 , n55392 , n55393 , n55394 , n55395 , n55396 , n55397 , n55398 , n55399 , n55400 , n55401 , n55402 , n55403 , n55404 , n55405 , n55406 , n55407 , n55408 , n55409 , n55410 , n55411 , n55412 , n55413 , n55414 , n55415 , n55416 , n55417 , n55418 , n55419 , n55420 , n55421 , n55422 , n55423 , n55424 , n55425 , n55426 , n55427 , n55428 , n55429 , n55430 , n55431 , n55432 , n55433 , n55434 , n55435 , n55436 , n55437 , n55438 , n55439 , n55440 , n55441 , n55442 , n55443 , n55444 , n55445 , n55446 , n55447 , n55448 , n55449 , n55450 , n55451 , n55452 , n55453 , n55454 , n55455 , n55456 , n55457 , n55458 , n55459 , n55460 , n55461 , n55462 , n55463 , n55464 , n55465 , n55466 , n55467 , n55468 , n55469 , n55470 , n55471 , n55472 , n55473 , n55474 , n55475 , n55476 , n55477 , n55478 , n55479 , n55480 , n55481 , n55482 , n55483 , n55484 , n55485 , n55486 , n55487 , n55488 , n55489 , n55490 , n55491 , n55492 , n55493 , n55494 , n55495 , n55496 , n55497 , n55498 , n55499 , n55500 , n55501 , n55502 , n55503 , n55504 , n55505 , n55506 , n55507 , n55508 , n55509 , n55510 , n55511 , n55512 , n55513 , n55514 , n55515 , n55516 , n55517 , n55518 , n55519 , n55520 , n55521 , n55522 , n55523 , n55524 , n55525 , n55526 , n55527 , n55528 , n55529 , n55530 , n55531 , n55532 , n55533 , n55534 , n55535 , n55536 , n55537 , n55538 , n55539 , n55540 , n55541 , n55542 , n55543 , n55544 , n55545 , n55546 , n55547 , n55548 , n55549 , n55550 , n55551 , n55552 , n55553 , n55554 , n55555 , n55556 , n55557 , n55558 , n55559 , n55560 , n55561 , n55562 , n55563 , n55564 , n55565 , n55566 , n55567 , n55568 , n55569 , n55570 , n55571 , n55572 , n55573 , n55574 , n55575 , n55576 , n55577 , n55578 , n55579 , n55580 , n55581 , n55582 , n55583 , n55584 , n55585 , n55586 , n55587 , n55588 , n55589 , n55590 , n55591 , n55592 , n55593 , n55594 , n55595 , n55596 , n55597 , n55598 , n55599 , n55600 , n55601 , n55602 , n55603 , n55604 , n55605 , n55606 , n55607 , n55608 , n55609 , n55610 , n55611 , n55612 , n55613 , n55614 , n55615 , n55616 , n55617 , n55618 , n55619 , n55620 , n55621 , n55622 , n55623 , n55624 , n55625 , n55626 , n55627 , n55628 , n55629 , n55630 , n55631 , n55632 , n55633 , n55634 , n55635 , n55636 , n55637 , n55638 , n55639 , n55640 , n55641 , n55642 , n55643 , n55644 , n55645 , n55646 , n55647 , n55648 , n55649 , n55650 , n55651 , n55652 , n55653 , n55654 , n55655 , n55656 , n55657 , n55658 , n55659 , n55660 , n55661 , n55662 , n55663 , n55664 , n55665 , n55666 , n55667 , n55668 , n55669 , n55670 , n55671 , n55672 , n55673 , n55674 , n55675 , n55676 , n55677 , n55678 , n55679 , n55680 , n55681 , n55682 , n55683 , n55684 , n55685 , n55686 , n55687 , n55688 , n55689 , n55690 , n55691 , n55692 , n55693 , n55694 , n55695 , n55696 , n55697 , n55698 , n55699 , n55700 , n55701 , n55702 , n55703 , n55704 , n55705 , n55706 , n55707 , n55708 , n55709 , n55710 , n55711 , n55712 , n55713 , n55714 , n55715 , n55716 , n55717 , n55718 , n55719 , n55720 , n55721 , n55722 , n55723 , n55724 , n55725 , n55726 , n55727 , n55728 , n55729 , n55730 , n55731 , n55732 , n55733 , n55734 , n55735 , n55736 , n55737 , n55738 , n55739 , n55740 , n55741 , n55742 , n55743 , n55744 , n55745 , n55746 , n55747 , n55748 , n55749 , n55750 , n55751 , n55752 , n55753 , n55754 , n55755 , n55756 , n55757 , n55758 , n55759 , n55760 , n55761 , n55762 , n55763 , n55764 , n55765 , n55766 , n55767 , n55768 , n55769 , n55770 , n55771 , n55772 , n55773 , n55774 , n55775 , n55776 , n55777 , n55778 , n55779 , n55780 , n55781 , n55782 , n55783 , n55784 , n55785 , n55786 , n55787 , n55788 , n55789 , n55790 , n55791 , n55792 , n55793 , n55794 , n55795 , n55796 , n55797 , n55798 , n55799 , n55800 , n55801 , n55802 , n55803 , n55804 , n55805 , n55806 , n55807 , n55808 , n55809 , n55810 , n55811 , n55812 , n55813 , n55814 , n55815 , n55816 , n55817 , n55818 , n55819 , n55820 , n55821 , n55822 , n55823 , n55824 , n55825 , n55826 , n55827 , n55828 , n55829 , n55830 , n55831 , n55832 , n55833 , n55834 , n55835 , n55836 , n55837 , n55838 , n55839 , n55840 , n55841 , n55842 , n55843 , n55844 , n55845 , n55846 , n55847 , n55848 , n55849 , n55850 , n55851 , n55852 , n55853 , n55854 , n55855 , n55856 , n55857 , n55858 , n55859 , n55860 , n55861 , n55862 , n55863 , n55864 , n55865 , n55866 , n55867 , n55868 , n55869 , n55870 , n55871 , n55872 , n55873 , n55874 , n55875 , n55876 , n55877 , n55878 , n55879 , n55880 , n55881 , n55882 , n55883 , n55884 , n55885 , n55886 , n55887 , n55888 , n55889 , n55890 , n55891 , n55892 , n55893 , n55894 , n55895 , n55896 , n55897 , n55898 , n55899 , n55900 , n55901 , n55902 , n55903 , n55904 , n55905 , n55906 , n55907 , n55908 , n55909 , n55910 , n55911 , n55912 , n55913 , n55914 , n55915 , n55916 , n55917 , n55918 , n55919 , n55920 , n55921 , n55922 , n55923 , n55924 , n55925 , n55926 , n55927 , n55928 , n55929 , n55930 , n55931 , n55932 , n55933 , n55934 , n55935 , n55936 , n55937 , n55938 , n55939 , n55940 , n55941 , n55942 , n55943 , n55944 , n55945 , n55946 , n55947 , n55948 , n55949 , n55950 , n55951 , n55952 , n55953 , n55954 , n55955 , n55956 , n55957 , n55958 , n55959 , n55960 , n55961 , n55962 , n55963 , n55964 , n55965 , n55966 , n55967 , n55968 , n55969 , n55970 , n55971 , n55972 , n55973 , n55974 , n55975 , n55976 , n55977 , n55978 , n55979 , n55980 , n55981 , n55982 , n55983 , n55984 , n55985 , n55986 , n55987 , n55988 , n55989 , n55990 , n55991 , n55992 , n55993 , n55994 , n55995 , n55996 , n55997 , n55998 , n55999 , n56000 , n56001 , n56002 , n56003 , n56004 , n56005 , n56006 , n56007 , n56008 , n56009 , n56010 , n56011 , n56012 , n56013 , n56014 , n56015 , n56016 , n56017 , n56018 , n56019 , n56020 , n56021 , n56022 , n56023 , n56024 , n56025 , n56026 , n56027 , n56028 , n56029 , n56030 , n56031 , n56032 , n56033 , n56034 , n56035 , n56036 , n56037 , n56038 , n56039 , n56040 , n56041 , n56042 , n56043 , n56044 , n56045 , n56046 , n56047 , n56048 , n56049 , n56050 , n56051 , n56052 , n56053 , n56054 , n56055 , n56056 , n56057 , n56058 , n56059 , n56060 , n56061 , n56062 , n56063 , n56064 , n56065 , n56066 , n56067 , n56068 , n56069 , n56070 , n56071 , n56072 , n56073 , n56074 , n56075 , n56076 , n56077 , n56078 , n56079 , n56080 , n56081 , n56082 , n56083 , n56084 , n56085 , n56086 , n56087 , n56088 , n56089 , n56090 , n56091 , n56092 , n56093 , n56094 , n56095 , n56096 , n56097 , n56098 , n56099 , n56100 , n56101 , n56102 , n56103 , n56104 , n56105 , n56106 , n56107 , n56108 , n56109 , n56110 , n56111 , n56112 , n56113 , n56114 , n56115 , n56116 , n56117 , n56118 , n56119 , n56120 , n56121 , n56122 , n56123 , n56124 , n56125 , n56126 , n56127 , n56128 , n56129 , n56130 , n56131 , n56132 , n56133 , n56134 , n56135 , n56136 , n56137 , n56138 , n56139 , n56140 , n56141 , n56142 , n56143 , n56144 , n56145 , n56146 , n56147 , n56148 , n56149 , n56150 , n56151 , n56152 , n56153 , n56154 , n56155 , n56156 , n56157 , n56158 , n56159 , n56160 , n56161 , n56162 , n56163 , n56164 , n56165 , n56166 , n56167 , n56168 , n56169 , n56170 , n56171 , n56172 , n56173 , n56174 , n56175 , n56176 , n56177 , n56178 , n56179 , n56180 , n56181 , n56182 , n56183 , n56184 , n56185 , n56186 , n56187 , n56188 , n56189 , n56190 , n56191 , n56192 , n56193 , n56194 , n56195 , n56196 , n56197 , n56198 , n56199 , n56200 , n56201 , n56202 , n56203 , n56204 , n56205 , n56206 , n56207 , n56208 , n56209 , n56210 , n56211 , n56212 , n56213 , n56214 , n56215 , n56216 , n56217 , n56218 , n56219 , n56220 , n56221 , n56222 , n56223 , n56224 , n56225 , n56226 , n56227 , n56228 , n56229 , n56230 , n56231 , n56232 , n56233 , n56234 , n56235 , n56236 , n56237 , n56238 , n56239 , n56240 , n56241 , n56242 , n56243 , n56244 , n56245 , n56246 , n56247 , n56248 , n56249 , n56250 , n56251 , n56252 , n56253 , n56254 , n56255 , n56256 , n56257 , n56258 , n56259 , n56260 , n56261 , n56262 , n56263 , n56264 , n56265 , n56266 , n56267 , n56268 , n56269 , n56270 , n56271 , n56272 , n56273 , n56274 , n56275 , n56276 , n56277 , n56278 , n56279 , n56280 , n56281 , n56282 , n56283 , n56284 , n56285 , n56286 , n56287 , n56288 , n56289 , n56290 , n56291 , n56292 , n56293 , n56294 , n56295 , n56296 , n56297 , n56298 , n56299 , n56300 , n56301 , n56302 , n56303 , n56304 , n56305 , n56306 , n56307 , n56308 , n56309 , n56310 , n56311 , n56312 , n56313 , n56314 , n56315 , n56316 , n56317 , n56318 , n56319 , n56320 , n56321 , n56322 , n56323 , n56324 , n56325 , n56326 , n56327 , n56328 , n56329 , n56330 , n56331 , n56332 , n56333 , n56334 , n56335 , n56336 , n56337 , n56338 , n56339 , n56340 , n56341 , n56342 , n56343 , n56344 , n56345 , n56346 , n56347 , n56348 , n56349 , n56350 , n56351 , n56352 , n56353 , n56354 , n56355 , n56356 , n56357 , n56358 , n56359 , n56360 , n56361 , n56362 , n56363 , n56364 , n56365 , n56366 , n56367 , n56368 , n56369 , n56370 , n56371 , n56372 , n56373 , n56374 , n56375 , n56376 , n56377 , n56378 , n56379 , n56380 , n56381 , n56382 , n56383 , n56384 , n56385 , n56386 , n56387 , n56388 , n56389 , n56390 , n56391 , n56392 , n56393 , n56394 , n56395 , n56396 , n56397 , n56398 , n56399 , n56400 , n56401 , n56402 , n56403 , n56404 , n56405 , n56406 , n56407 , n56408 , n56409 , n56410 , n56411 , n56412 , n56413 , n56414 , n56415 , n56416 , n56417 , n56418 , n56419 , n56420 , n56421 , n56422 , n56423 , n56424 , n56425 , n56426 , n56427 , n56428 , n56429 , n56430 , n56431 , n56432 , n56433 , n56434 , n56435 , n56436 , n56437 , n56438 , n56439 , n56440 , n56441 , n56442 , n56443 , n56444 , n56445 , n56446 , n56447 , n56448 , n56449 , n56450 , n56451 , n56452 , n56453 , n56454 , n56455 , n56456 , n56457 , n56458 , n56459 , n56460 , n56461 , n56462 , n56463 , n56464 , n56465 , n56466 , n56467 , n56468 , n56469 , n56470 , n56471 , n56472 , n56473 , n56474 , n56475 , n56476 , n56477 , n56478 , n56479 , n56480 , n56481 , n56482 , n56483 , n56484 , n56485 , n56486 , n56487 , n56488 , n56489 , n56490 , n56491 , n56492 , n56493 , n56494 , n56495 , n56496 , n56497 , n56498 , n56499 , n56500 , n56501 , n56502 , n56503 , n56504 , n56505 , n56506 , n56507 , n56508 , n56509 , n56510 , n56511 , n56512 , n56513 , n56514 , n56515 , n56516 , n56517 , n56518 , n56519 , n56520 , n56521 , n56522 , n56523 , n56524 , n56525 , n56526 , n56527 , n56528 , n56529 , n56530 , n56531 , n56532 , n56533 , n56534 , n56535 , n56536 , n56537 , n56538 , n56539 , n56540 , n56541 , n56542 , n56543 , n56544 , n56545 , n56546 , n56547 , n56548 , n56549 , n56550 , n56551 , n56552 , n56553 , n56554 , n56555 , n56556 , n56557 , n56558 , n56559 , n56560 , n56561 , n56562 , n56563 , n56564 , n56565 , n56566 , n56567 , n56568 , n56569 , n56570 , n56571 , n56572 , n56573 , n56574 , n56575 , n56576 , n56577 , n56578 , n56579 , n56580 , n56581 , n56582 , n56583 , n56584 , n56585 , n56586 , n56587 , n56588 , n56589 , n56590 , n56591 , n56592 , n56593 , n56594 , n56595 , n56596 , n56597 , n56598 , n56599 , n56600 , n56601 , n56602 , n56603 , n56604 , n56605 , n56606 , n56607 , n56608 , n56609 , n56610 , n56611 , n56612 , n56613 , n56614 , n56615 , n56616 , n56617 , n56618 , n56619 , n56620 , n56621 , n56622 , n56623 , n56624 , n56625 , n56626 , n56627 , n56628 , n56629 , n56630 , n56631 , n56632 , n56633 , n56634 , n56635 , n56636 , n56637 , n56638 , n56639 , n56640 , n56641 , n56642 , n56643 , n56644 , n56645 , n56646 , n56647 , n56648 , n56649 , n56650 , n56651 , n56652 , n56653 , n56654 , n56655 , n56656 , n56657 , n56658 , n56659 , n56660 , n56661 , n56662 , n56663 , n56664 , n56665 , n56666 , n56667 , n56668 , n56669 , n56670 , n56671 , n56672 , n56673 , n56674 , n56675 , n56676 , n56677 , n56678 , n56679 , n56680 , n56681 , n56682 , n56683 , n56684 , n56685 , n56686 , n56687 , n56688 , n56689 , n56690 , n56691 , n56692 , n56693 , n56694 , n56695 , n56696 , n56697 , n56698 , n56699 , n56700 , n56701 , n56702 , n56703 , n56704 , n56705 , n56706 , n56707 , n56708 , n56709 , n56710 , n56711 , n56712 , n56713 , n56714 , n56715 , n56716 , n56717 , n56718 , n56719 , n56720 , n56721 , n56722 , n56723 , n56724 , n56725 , n56726 , n56727 , n56728 , n56729 , n56730 , n56731 , n56732 , n56733 , n56734 , n56735 , n56736 , n56737 , n56738 , n56739 , n56740 , n56741 , n56742 , n56743 , n56744 , n56745 , n56746 , n56747 , n56748 , n56749 , n56750 , n56751 , n56752 , n56753 , n56754 , n56755 , n56756 , n56757 , n56758 , n56759 , n56760 , n56761 , n56762 , n56763 , n56764 , n56765 , n56766 , n56767 , n56768 , n56769 , n56770 , n56771 , n56772 , n56773 , n56774 , n56775 , n56776 , n56777 , n56778 , n56779 , n56780 , n56781 , n56782 , n56783 , n56784 , n56785 , n56786 , n56787 , n56788 , n56789 , n56790 , n56791 , n56792 , n56793 , n56794 , n56795 , n56796 , n56797 , n56798 , n56799 , n56800 , n56801 , n56802 , n56803 , n56804 , n56805 , n56806 , n56807 , n56808 , n56809 , n56810 , n56811 , n56812 , n56813 , n56814 , n56815 , n56816 , n56817 , n56818 , n56819 , n56820 , n56821 , n56822 , n56823 , n56824 , n56825 , n56826 , n56827 , n56828 , n56829 , n56830 , n56831 , n56832 , n56833 , n56834 , n56835 , n56836 , n56837 , n56838 , n56839 , n56840 , n56841 , n56842 , n56843 , n56844 , n56845 , n56846 , n56847 , n56848 , n56849 , n56850 , n56851 , n56852 , n56853 , n56854 , n56855 , n56856 , n56857 , n56858 , n56859 , n56860 , n56861 , n56862 , n56863 , n56864 , n56865 , n56866 , n56867 , n56868 , n56869 , n56870 , n56871 , n56872 , n56873 , n56874 , n56875 , n56876 , n56877 , n56878 , n56879 , n56880 , n56881 , n56882 , n56883 , n56884 , n56885 , n56886 , n56887 , n56888 , n56889 , n56890 , n56891 , n56892 , n56893 , n56894 , n56895 , n56896 , n56897 , n56898 , n56899 , n56900 , n56901 , n56902 , n56903 , n56904 , n56905 , n56906 , n56907 , n56908 , n56909 , n56910 , n56911 , n56912 , n56913 , n56914 , n56915 , n56916 , n56917 , n56918 , n56919 , n56920 , n56921 , n56922 , n56923 , n56924 , n56925 , n56926 , n56927 , n56928 , n56929 , n56930 , n56931 , n56932 , n56933 , n56934 , n56935 , n56936 , n56937 , n56938 , n56939 , n56940 , n56941 , n56942 , n56943 , n56944 , n56945 , n56946 , n56947 , n56948 , n56949 , n56950 , n56951 , n56952 , n56953 , n56954 , n56955 , n56956 , n56957 , n56958 , n56959 , n56960 , n56961 , n56962 , n56963 , n56964 , n56965 , n56966 , n56967 , n56968 , n56969 , n56970 , n56971 , n56972 , n56973 , n56974 , n56975 , n56976 , n56977 , n56978 , n56979 , n56980 , n56981 , n56982 , n56983 , n56984 , n56985 , n56986 , n56987 , n56988 , n56989 , n56990 , n56991 , n56992 , n56993 , n56994 , n56995 , n56996 , n56997 , n56998 , n56999 , n57000 , n57001 , n57002 , n57003 , n57004 , n57005 , n57006 , n57007 , n57008 , n57009 , n57010 , n57011 , n57012 , n57013 , n57014 , n57015 , n57016 , n57017 , n57018 , n57019 , n57020 , n57021 , n57022 , n57023 , n57024 , n57025 , n57026 , n57027 , n57028 , n57029 , n57030 , n57031 , n57032 , n57033 , n57034 , n57035 , n57036 , n57037 , n57038 , n57039 , n57040 , n57041 , n57042 , n57043 , n57044 , n57045 , n57046 , n57047 , n57048 , n57049 , n57050 , n57051 , n57052 , n57053 , n57054 , n57055 , n57056 , n57057 , n57058 , n57059 , n57060 , n57061 , n57062 , n57063 , n57064 , n57065 , n57066 , n57067 , n57068 , n57069 , n57070 , n57071 , n57072 , n57073 , n57074 , n57075 , n57076 , n57077 , n57078 , n57079 , n57080 , n57081 , n57082 , n57083 , n57084 , n57085 , n57086 , n57087 , n57088 , n57089 , n57090 , n57091 , n57092 , n57093 , n57094 , n57095 , n57096 , n57097 , n57098 , n57099 , n57100 , n57101 , n57102 , n57103 , n57104 , n57105 , n57106 , n57107 , n57108 , n57109 , n57110 , n57111 , n57112 , n57113 , n57114 , n57115 , n57116 , n57117 , n57118 , n57119 , n57120 , n57121 , n57122 , n57123 , n57124 , n57125 , n57126 , n57127 , n57128 , n57129 , n57130 , n57131 , n57132 , n57133 , n57134 , n57135 , n57136 , n57137 , n57138 , n57139 , n57140 , n57141 , n57142 , n57143 , n57144 , n57145 , n57146 , n57147 , n57148 , n57149 , n57150 , n57151 , n57152 , n57153 , n57154 , n57155 , n57156 , n57157 , n57158 , n57159 , n57160 , n57161 , n57162 , n57163 , n57164 , n57165 , n57166 , n57167 , n57168 , n57169 , n57170 , n57171 , n57172 , n57173 , n57174 , n57175 , n57176 , n57177 , n57178 , n57179 , n57180 , n57181 , n57182 , n57183 , n57184 , n57185 , n57186 , n57187 , n57188 , n57189 , n57190 , n57191 , n57192 , n57193 , n57194 , n57195 , n57196 , n57197 , n57198 , n57199 , n57200 , n57201 , n57202 , n57203 , n57204 , n57205 , n57206 , n57207 , n57208 , n57209 , n57210 , n57211 , n57212 , n57213 , n57214 , n57215 , n57216 , n57217 , n57218 , n57219 , n57220 , n57221 , n57222 , n57223 , n57224 , n57225 , n57226 , n57227 , n57228 , n57229 , n57230 , n57231 , n57232 , n57233 , n57234 , n57235 , n57236 , n57237 , n57238 , n57239 , n57240 , n57241 , n57242 , n57243 , n57244 , n57245 , n57246 , n57247 , n57248 , n57249 , n57250 , n57251 , n57252 , n57253 , n57254 , n57255 , n57256 , n57257 , n57258 , n57259 , n57260 , n57261 , n57262 , n57263 , n57264 , n57265 , n57266 , n57267 , n57268 , n57269 , n57270 , n57271 , n57272 , n57273 , n57274 , n57275 , n57276 , n57277 , n57278 , n57279 , n57280 , n57281 , n57282 , n57283 , n57284 , n57285 , n57286 , n57287 , n57288 , n57289 , n57290 , n57291 , n57292 , n57293 , n57294 , n57295 , n57296 , n57297 , n57298 , n57299 , n57300 , n57301 , n57302 , n57303 , n57304 , n57305 , n57306 , n57307 , n57308 , n57309 , n57310 , n57311 , n57312 , n57313 , n57314 , n57315 , n57316 , n57317 , n57318 , n57319 , n57320 , n57321 , n57322 , n57323 , n57324 , n57325 , n57326 , n57327 , n57328 , n57329 , n57330 , n57331 , n57332 , n57333 , n57334 , n57335 , n57336 , n57337 , n57338 , n57339 , n57340 , n57341 , n57342 , n57343 , n57344 , n57345 , n57346 , n57347 , n57348 , n57349 , n57350 , n57351 , n57352 , n57353 , n57354 , n57355 , n57356 , n57357 , n57358 , n57359 , n57360 , n57361 , n57362 , n57363 , n57364 , n57365 , n57366 , n57367 , n57368 , n57369 , n57370 , n57371 , n57372 , n57373 , n57374 , n57375 , n57376 , n57377 , n57378 , n57379 , n57380 , n57381 , n57382 , n57383 , n57384 , n57385 , n57386 , n57387 , n57388 , n57389 , n57390 , n57391 , n57392 , n57393 , n57394 , n57395 , n57396 , n57397 , n57398 , n57399 , n57400 , n57401 , n57402 , n57403 , n57404 , n57405 , n57406 , n57407 , n57408 , n57409 , n57410 , n57411 , n57412 , n57413 , n57414 , n57415 , n57416 , n57417 , n57418 , n57419 , n57420 , n57421 , n57422 , n57423 , n57424 , n57425 , n57426 , n57427 , n57428 , n57429 , n57430 , n57431 , n57432 , n57433 , n57434 , n57435 , n57436 , n57437 , n57438 , n57439 , n57440 , n57441 , n57442 , n57443 , n57444 , n57445 , n57446 , n57447 , n57448 , n57449 , n57450 , n57451 , n57452 , n57453 , n57454 , n57455 , n57456 , n57457 , n57458 , n57459 , n57460 , n57461 , n57462 , n57463 , n57464 , n57465 , n57466 , n57467 , n57468 , n57469 , n57470 , n57471 , n57472 , n57473 , n57474 , n57475 , n57476 , n57477 , n57478 , n57479 , n57480 , n57481 , n57482 , n57483 , n57484 , n57485 , n57486 , n57487 , n57488 , n57489 , n57490 , n57491 , n57492 , n57493 , n57494 , n57495 , n57496 , n57497 , n57498 , n57499 , n57500 , n57501 , n57502 , n57503 , n57504 , n57505 , n57506 , n57507 , n57508 , n57509 , n57510 , n57511 , n57512 , n57513 , n57514 , n57515 , n57516 , n57517 , n57518 , n57519 , n57520 , n57521 , n57522 , n57523 , n57524 , n57525 , n57526 , n57527 , n57528 , n57529 , n57530 , n57531 , n57532 , n57533 , n57534 , n57535 , n57536 , n57537 , n57538 , n57539 , n57540 , n57541 , n57542 , n57543 , n57544 , n57545 , n57546 , n57547 , n57548 , n57549 , n57550 , n57551 , n57552 , n57553 , n57554 , n57555 , n57556 , n57557 , n57558 , n57559 , n57560 , n57561 , n57562 , n57563 , n57564 , n57565 , n57566 , n57567 , n57568 , n57569 , n57570 , n57571 , n57572 , n57573 , n57574 , n57575 , n57576 , n57577 , n57578 , n57579 , n57580 , n57581 , n57582 , n57583 , n57584 , n57585 , n57586 , n57587 , n57588 , n57589 , n57590 , n57591 , n57592 , n57593 , n57594 , n57595 , n57596 , n57597 , n57598 , n57599 , n57600 , n57601 , n57602 , n57603 , n57604 , n57605 , n57606 , n57607 , n57608 , n57609 , n57610 , n57611 , n57612 , n57613 , n57614 , n57615 , n57616 , n57617 , n57618 , n57619 , n57620 , n57621 , n57622 , n57623 , n57624 , n57625 , n57626 , n57627 , n57628 , n57629 , n57630 , n57631 , n57632 , n57633 , n57634 , n57635 , n57636 , n57637 , n57638 , n57639 , n57640 , n57641 , n57642 , n57643 , n57644 , n57645 , n57646 , n57647 , n57648 , n57649 , n57650 , n57651 , n57652 , n57653 , n57654 , n57655 , n57656 , n57657 , n57658 , n57659 , n57660 , n57661 , n57662 , n57663 , n57664 , n57665 , n57666 , n57667 , n57668 , n57669 , n57670 , n57671 , n57672 , n57673 , n57674 , n57675 , n57676 , n57677 , n57678 , n57679 , n57680 , n57681 , n57682 , n57683 , n57684 , n57685 , n57686 , n57687 , n57688 , n57689 , n57690 , n57691 , n57692 , n57693 , n57694 , n57695 , n57696 , n57697 , n57698 , n57699 , n57700 , n57701 , n57702 , n57703 , n57704 , n57705 , n57706 , n57707 , n57708 , n57709 , n57710 , n57711 , n57712 , n57713 , n57714 , n57715 , n57716 , n57717 , n57718 , n57719 , n57720 , n57721 , n57722 , n57723 , n57724 , n57725 , n57726 , n57727 , n57728 , n57729 , n57730 , n57731 , n57732 , n57733 , n57734 , n57735 , n57736 , n57737 , n57738 , n57739 , n57740 , n57741 , n57742 , n57743 , n57744 , n57745 , n57746 , n57747 , n57748 , n57749 , n57750 , n57751 , n57752 , n57753 , n57754 , n57755 , n57756 , n57757 , n57758 , n57759 , n57760 , n57761 , n57762 , n57763 , n57764 , n57765 , n57766 , n57767 , n57768 , n57769 , n57770 , n57771 , n57772 , n57773 , n57774 , n57775 , n57776 , n57777 , n57778 , n57779 , n57780 , n57781 , n57782 , n57783 , n57784 , n57785 , n57786 , n57787 , n57788 , n57789 , n57790 , n57791 , n57792 , n57793 , n57794 , n57795 , n57796 , n57797 , n57798 , n57799 , n57800 , n57801 , n57802 , n57803 , n57804 , n57805 , n57806 , n57807 , n57808 , n57809 , n57810 , n57811 , n57812 , n57813 , n57814 , n57815 , n57816 , n57817 , n57818 , n57819 , n57820 , n57821 , n57822 , n57823 , n57824 , n57825 , n57826 , n57827 , n57828 , n57829 , n57830 , n57831 , n57832 , n57833 , n57834 , n57835 , n57836 , n57837 , n57838 , n57839 , n57840 , n57841 , n57842 , n57843 , n57844 , n57845 , n57846 , n57847 , n57848 , n57849 , n57850 , n57851 , n57852 , n57853 , n57854 , n57855 , n57856 , n57857 , n57858 , n57859 , n57860 , n57861 , n57862 , n57863 , n57864 , n57865 , n57866 , n57867 , n57868 , n57869 , n57870 , n57871 , n57872 , n57873 , n57874 , n57875 , n57876 , n57877 , n57878 , n57879 , n57880 , n57881 , n57882 , n57883 , n57884 , n57885 , n57886 , n57887 , n57888 , n57889 , n57890 , n57891 , n57892 , n57893 , n57894 , n57895 , n57896 , n57897 , n57898 , n57899 , n57900 , n57901 , n57902 , n57903 , n57904 , n57905 , n57906 , n57907 , n57908 , n57909 , n57910 , n57911 , n57912 , n57913 , n57914 , n57915 , n57916 , n57917 , n57918 , n57919 , n57920 , n57921 , n57922 , n57923 , n57924 , n57925 , n57926 , n57927 , n57928 , n57929 , n57930 , n57931 , n57932 , n57933 , n57934 , n57935 , n57936 , n57937 , n57938 , n57939 , n57940 , n57941 , n57942 , n57943 , n57944 , n57945 , n57946 , n57947 , n57948 , n57949 , n57950 , n57951 , n57952 , n57953 , n57954 , n57955 , n57956 , n57957 , n57958 , n57959 , n57960 , n57961 , n57962 , n57963 , n57964 , n57965 , n57966 , n57967 , n57968 , n57969 , n57970 , n57971 , n57972 , n57973 , n57974 , n57975 , n57976 , n57977 , n57978 , n57979 , n57980 , n57981 , n57982 , n57983 , n57984 , n57985 , n57986 , n57987 , n57988 , n57989 , n57990 , n57991 , n57992 , n57993 , n57994 , n57995 , n57996 , n57997 , n57998 , n57999 , n58000 , n58001 , n58002 , n58003 , n58004 , n58005 , n58006 , n58007 , n58008 , n58009 , n58010 , n58011 , n58012 , n58013 , n58014 , n58015 , n58016 , n58017 , n58018 , n58019 , n58020 , n58021 , n58022 , n58023 , n58024 , n58025 , n58026 , n58027 , n58028 , n58029 , n58030 , n58031 , n58032 , n58033 , n58034 , n58035 , n58036 , n58037 , n58038 , n58039 , n58040 , n58041 , n58042 , n58043 , n58044 , n58045 , n58046 , n58047 , n58048 , n58049 , n58050 , n58051 , n58052 , n58053 , n58054 , n58055 , n58056 , n58057 , n58058 , n58059 , n58060 , n58061 , n58062 , n58063 , n58064 , n58065 , n58066 , n58067 , n58068 , n58069 , n58070 , n58071 , n58072 , n58073 , n58074 , n58075 , n58076 , n58077 , n58078 , n58079 , n58080 , n58081 , n58082 , n58083 , n58084 , n58085 , n58086 , n58087 , n58088 , n58089 , n58090 , n58091 , n58092 , n58093 , n58094 , n58095 , n58096 , n58097 , n58098 , n58099 , n58100 , n58101 , n58102 , n58103 , n58104 , n58105 , n58106 , n58107 , n58108 , n58109 , n58110 , n58111 , n58112 , n58113 , n58114 , n58115 , n58116 , n58117 , n58118 , n58119 , n58120 , n58121 , n58122 , n58123 , n58124 , n58125 , n58126 , n58127 , n58128 , n58129 , n58130 , n58131 , n58132 , n58133 , n58134 , n58135 , n58136 , n58137 , n58138 , n58139 , n58140 , n58141 , n58142 , n58143 , n58144 , n58145 , n58146 , n58147 , n58148 , n58149 , n58150 , n58151 , n58152 , n58153 , n58154 , n58155 , n58156 , n58157 , n58158 , n58159 , n58160 , n58161 , n58162 , n58163 , n58164 , n58165 , n58166 , n58167 , n58168 , n58169 , n58170 , n58171 , n58172 , n58173 , n58174 , n58175 , n58176 , n58177 , n58178 , n58179 , n58180 , n58181 , n58182 , n58183 , n58184 , n58185 , n58186 , n58187 , n58188 , n58189 , n58190 , n58191 , n58192 , n58193 , n58194 , n58195 , n58196 , n58197 , n58198 , n58199 , n58200 , n58201 , n58202 , n58203 , n58204 , n58205 , n58206 , n58207 , n58208 , n58209 , n58210 , n58211 , n58212 , n58213 , n58214 , n58215 , n58216 , n58217 , n58218 , n58219 , n58220 , n58221 , n58222 , n58223 , n58224 , n58225 , n58226 , n58227 , n58228 , n58229 , n58230 , n58231 , n58232 , n58233 , n58234 , n58235 , n58236 , n58237 , n58238 , n58239 , n58240 , n58241 , n58242 , n58243 , n58244 , n58245 , n58246 , n58247 , n58248 , n58249 , n58250 , n58251 , n58252 , n58253 , n58254 , n58255 , n58256 , n58257 , n58258 , n58259 , n58260 , n58261 , n58262 , n58263 , n58264 , n58265 , n58266 , n58267 , n58268 , n58269 , n58270 , n58271 , n58272 , n58273 , n58274 , n58275 , n58276 , n58277 , n58278 , n58279 , n58280 , n58281 , n58282 , n58283 , n58284 , n58285 , n58286 , n58287 , n58288 , n58289 , n58290 , n58291 , n58292 , n58293 , n58294 , n58295 , n58296 , n58297 , n58298 , n58299 , n58300 , n58301 , n58302 , n58303 , n58304 , n58305 , n58306 , n58307 , n58308 , n58309 , n58310 , n58311 , n58312 , n58313 , n58314 , n58315 , n58316 , n58317 , n58318 , n58319 , n58320 , n58321 , n58322 , n58323 , n58324 , n58325 , n58326 , n58327 , n58328 , n58329 , n58330 , n58331 , n58332 , n58333 , n58334 , n58335 , n58336 , n58337 , n58338 , n58339 , n58340 , n58341 , n58342 , n58343 , n58344 , n58345 , n58346 , n58347 , n58348 , n58349 , n58350 , n58351 , n58352 , n58353 , n58354 , n58355 , n58356 , n58357 , n58358 , n58359 , n58360 , n58361 , n58362 , n58363 , n58364 , n58365 , n58366 , n58367 , n58368 , n58369 , n58370 , n58371 , n58372 , n58373 , n58374 , n58375 , n58376 , n58377 , n58378 , n58379 , n58380 , n58381 , n58382 , n58383 , n58384 , n58385 , n58386 , n58387 , n58388 , n58389 , n58390 , n58391 , n58392 , n58393 , n58394 , n58395 , n58396 , n58397 , n58398 , n58399 , n58400 , n58401 , n58402 , n58403 , n58404 , n58405 , n58406 , n58407 , n58408 , n58409 , n58410 , n58411 , n58412 , n58413 , n58414 , n58415 , n58416 , n58417 , n58418 , n58419 , n58420 , n58421 , n58422 , n58423 , n58424 , n58425 , n58426 , n58427 , n58428 , n58429 , n58430 , n58431 , n58432 , n58433 , n58434 , n58435 , n58436 , n58437 , n58438 , n58439 , n58440 , n58441 , n58442 , n58443 , n58444 , n58445 , n58446 , n58447 , n58448 , n58449 , n58450 , n58451 , n58452 , n58453 , n58454 , n58455 , n58456 , n58457 , n58458 , n58459 , n58460 , n58461 , n58462 , n58463 , n58464 , n58465 , n58466 , n58467 , n58468 , n58469 , n58470 , n58471 , n58472 , n58473 , n58474 , n58475 , n58476 , n58477 , n58478 , n58479 , n58480 , n58481 , n58482 , n58483 , n58484 , n58485 , n58486 , n58487 , n58488 , n58489 , n58490 , n58491 , n58492 , n58493 , n58494 , n58495 , n58496 , n58497 , n58498 , n58499 , n58500 , n58501 , n58502 , n58503 , n58504 , n58505 , n58506 , n58507 , n58508 , n58509 , n58510 , n58511 , n58512 , n58513 , n58514 , n58515 , n58516 , n58517 , n58518 , n58519 , n58520 , n58521 , n58522 , n58523 , n58524 , n58525 , n58526 , n58527 , n58528 , n58529 , n58530 , n58531 , n58532 , n58533 , n58534 , n58535 , n58536 , n58537 , n58538 , n58539 , n58540 , n58541 , n58542 , n58543 , n58544 , n58545 , n58546 , n58547 , n58548 , n58549 , n58550 , n58551 , n58552 , n58553 , n58554 , n58555 , n58556 , n58557 , n58558 , n58559 , n58560 , n58561 , n58562 , n58563 , n58564 , n58565 , n58566 , n58567 , n58568 , n58569 , n58570 , n58571 , n58572 , n58573 , n58574 , n58575 , n58576 , n58577 , n58578 , n58579 , n58580 , n58581 , n58582 , n58583 , n58584 , n58585 , n58586 , n58587 , n58588 , n58589 , n58590 , n58591 , n58592 , n58593 , n58594 , n58595 , n58596 , n58597 , n58598 , n58599 , n58600 , n58601 , n58602 , n58603 , n58604 , n58605 , n58606 , n58607 , n58608 , n58609 , n58610 , n58611 , n58612 , n58613 , n58614 , n58615 , n58616 , n58617 , n58618 , n58619 , n58620 , n58621 , n58622 , n58623 , n58624 , n58625 , n58626 , n58627 , n58628 , n58629 , n58630 , n58631 , n58632 , n58633 , n58634 , n58635 , n58636 , n58637 , n58638 , n58639 , n58640 , n58641 , n58642 , n58643 , n58644 , n58645 , n58646 , n58647 , n58648 , n58649 , n58650 , n58651 , n58652 , n58653 , n58654 , n58655 , n58656 , n58657 , n58658 , n58659 , n58660 , n58661 , n58662 , n58663 , n58664 , n58665 , n58666 , n58667 , n58668 , n58669 , n58670 , n58671 , n58672 , n58673 , n58674 , n58675 , n58676 , n58677 , n58678 , n58679 , n58680 , n58681 , n58682 , n58683 , n58684 , n58685 , n58686 , n58687 , n58688 , n58689 , n58690 , n58691 , n58692 , n58693 , n58694 , n58695 , n58696 , n58697 , n58698 , n58699 , n58700 , n58701 , n58702 , n58703 , n58704 , n58705 , n58706 , n58707 , n58708 , n58709 , n58710 , n58711 , n58712 , n58713 , n58714 , n58715 , n58716 , n58717 , n58718 , n58719 , n58720 , n58721 , n58722 , n58723 , n58724 , n58725 , n58726 , n58727 , n58728 , n58729 , n58730 , n58731 , n58732 , n58733 , n58734 , n58735 , n58736 , n58737 , n58738 , n58739 , n58740 , n58741 , n58742 , n58743 , n58744 , n58745 , n58746 , n58747 , n58748 , n58749 , n58750 , n58751 , n58752 , n58753 , n58754 , n58755 , n58756 , n58757 , n58758 , n58759 , n58760 , n58761 , n58762 , n58763 , n58764 , n58765 , n58766 , n58767 , n58768 , n58769 , n58770 , n58771 , n58772 , n58773 , n58774 , n58775 , n58776 , n58777 , n58778 , n58779 , n58780 , n58781 , n58782 , n58783 , n58784 , n58785 , n58786 , n58787 , n58788 , n58789 , n58790 , n58791 , n58792 , n58793 , n58794 , n58795 , n58796 , n58797 , n58798 , n58799 , n58800 , n58801 , n58802 , n58803 , n58804 , n58805 , n58806 , n58807 , n58808 , n58809 , n58810 , n58811 , n58812 , n58813 , n58814 , n58815 , n58816 , n58817 , n58818 , n58819 , n58820 , n58821 , n58822 , n58823 , n58824 , n58825 , n58826 , n58827 , n58828 , n58829 , n58830 , n58831 , n58832 , n58833 , n58834 , n58835 , n58836 , n58837 , n58838 , n58839 , n58840 , n58841 , n58842 , n58843 , n58844 , n58845 , n58846 , n58847 , n58848 , n58849 , n58850 , n58851 , n58852 , n58853 , n58854 , n58855 , n58856 , n58857 , n58858 , n58859 , n58860 , n58861 , n58862 , n58863 , n58864 , n58865 , n58866 , n58867 , n58868 , n58869 , n58870 , n58871 , n58872 , n58873 , n58874 , n58875 , n58876 , n58877 , n58878 , n58879 , n58880 , n58881 , n58882 , n58883 , n58884 , n58885 , n58886 , n58887 , n58888 , n58889 , n58890 , n58891 , n58892 , n58893 , n58894 , n58895 , n58896 , n58897 , n58898 , n58899 , n58900 , n58901 , n58902 , n58903 , n58904 , n58905 , n58906 , n58907 , n58908 , n58909 , n58910 , n58911 , n58912 , n58913 , n58914 , n58915 , n58916 , n58917 , n58918 , n58919 , n58920 , n58921 , n58922 , n58923 , n58924 , n58925 , n58926 , n58927 , n58928 , n58929 , n58930 , n58931 , n58932 , n58933 , n58934 , n58935 , n58936 , n58937 , n58938 , n58939 , n58940 , n58941 , n58942 , n58943 , n58944 , n58945 , n58946 , n58947 , n58948 , n58949 , n58950 , n58951 , n58952 , n58953 , n58954 , n58955 , n58956 , n58957 , n58958 , n58959 , n58960 , n58961 , n58962 , n58963 , n58964 , n58965 , n58966 , n58967 , n58968 , n58969 , n58970 , n58971 , n58972 , n58973 , n58974 , n58975 , n58976 , n58977 , n58978 , n58979 , n58980 , n58981 , n58982 , n58983 , n58984 , n58985 , n58986 , n58987 , n58988 , n58989 , n58990 , n58991 , n58992 , n58993 , n58994 , n58995 , n58996 , n58997 , n58998 , n58999 , n59000 , n59001 , n59002 , n59003 , n59004 , n59005 , n59006 , n59007 , n59008 , n59009 , n59010 , n59011 , n59012 , n59013 , n59014 , n59015 , n59016 , n59017 , n59018 , n59019 , n59020 , n59021 , n59022 , n59023 , n59024 , n59025 , n59026 , n59027 , n59028 , n59029 , n59030 , n59031 , n59032 , n59033 , n59034 , n59035 , n59036 , n59037 , n59038 , n59039 , n59040 , n59041 , n59042 , n59043 , n59044 , n59045 , n59046 , n59047 , n59048 , n59049 , n59050 , n59051 , n59052 , n59053 , n59054 , n59055 , n59056 , n59057 , n59058 , n59059 , n59060 , n59061 , n59062 , n59063 , n59064 , n59065 , n59066 , n59067 , n59068 , n59069 , n59070 , n59071 , n59072 , n59073 , n59074 , n59075 , n59076 , n59077 , n59078 , n59079 , n59080 , n59081 , n59082 , n59083 , n59084 , n59085 , n59086 , n59087 , n59088 , n59089 , n59090 , n59091 , n59092 , n59093 , n59094 , n59095 , n59096 , n59097 , n59098 , n59099 , n59100 , n59101 , n59102 , n59103 , n59104 , n59105 , n59106 , n59107 , n59108 , n59109 , n59110 , n59111 , n59112 , n59113 , n59114 , n59115 , n59116 , n59117 , n59118 , n59119 , n59120 , n59121 , n59122 , n59123 , n59124 , n59125 , n59126 , n59127 , n59128 , n59129 , n59130 , n59131 , n59132 , n59133 , n59134 , n59135 , n59136 , n59137 , n59138 , n59139 , n59140 , n59141 , n59142 , n59143 , n59144 , n59145 , n59146 , n59147 , n59148 , n59149 , n59150 , n59151 , n59152 , n59153 , n59154 , n59155 , n59156 , n59157 , n59158 , n59159 , n59160 , n59161 , n59162 , n59163 , n59164 , n59165 , n59166 , n59167 , n59168 , n59169 , n59170 , n59171 , n59172 , n59173 , n59174 , n59175 , n59176 , n59177 , n59178 , n59179 , n59180 , n59181 , n59182 , n59183 , n59184 , n59185 , n59186 , n59187 , n59188 , n59189 , n59190 , n59191 , n59192 , n59193 , n59194 , n59195 , n59196 , n59197 , n59198 , n59199 , n59200 , n59201 , n59202 , n59203 , n59204 , n59205 , n59206 , n59207 , n59208 , n59209 , n59210 , n59211 , n59212 , n59213 , n59214 , n59215 , n59216 , n59217 , n59218 , n59219 , n59220 , n59221 , n59222 , n59223 , n59224 , n59225 , n59226 , n59227 , n59228 , n59229 , n59230 , n59231 , n59232 , n59233 , n59234 , n59235 , n59236 , n59237 , n59238 , n59239 , n59240 , n59241 , n59242 , n59243 , n59244 , n59245 , n59246 , n59247 , n59248 , n59249 , n59250 , n59251 , n59252 , n59253 , n59254 , n59255 , n59256 , n59257 , n59258 , n59259 , n59260 , n59261 , n59262 , n59263 , n59264 , n59265 , n59266 , n59267 , n59268 , n59269 , n59270 , n59271 , n59272 , n59273 , n59274 , n59275 , n59276 , n59277 , n59278 , n59279 , n59280 , n59281 , n59282 , n59283 , n59284 , n59285 , n59286 , n59287 , n59288 , n59289 , n59290 , n59291 , n59292 , n59293 , n59294 , n59295 , n59296 , n59297 , n59298 , n59299 , n59300 , n59301 , n59302 , n59303 , n59304 , n59305 , n59306 , n59307 , n59308 , n59309 , n59310 , n59311 , n59312 , n59313 , n59314 , n59315 , n59316 , n59317 , n59318 , n59319 , n59320 , n59321 , n59322 , n59323 , n59324 , n59325 , n59326 , n59327 , n59328 , n59329 , n59330 , n59331 , n59332 , n59333 , n59334 , n59335 , n59336 , n59337 , n59338 , n59339 , n59340 , n59341 , n59342 , n59343 , n59344 , n59345 , n59346 , n59347 , n59348 , n59349 , n59350 , n59351 , n59352 , n59353 , n59354 , n59355 , n59356 , n59357 , n59358 , n59359 , n59360 , n59361 , n59362 , n59363 , n59364 , n59365 , n59366 , n59367 , n59368 , n59369 , n59370 , n59371 , n59372 , n59373 , n59374 , n59375 , n59376 , n59377 , n59378 , n59379 , n59380 , n59381 , n59382 , n59383 , n59384 , n59385 , n59386 , n59387 , n59388 , n59389 , n59390 , n59391 , n59392 , n59393 , n59394 , n59395 , n59396 , n59397 , n59398 , n59399 , n59400 , n59401 , n59402 , n59403 , n59404 , n59405 , n59406 , n59407 , n59408 , n59409 , n59410 , n59411 , n59412 , n59413 , n59414 , n59415 , n59416 , n59417 , n59418 , n59419 , n59420 , n59421 , n59422 , n59423 , n59424 , n59425 , n59426 , n59427 , n59428 , n59429 , n59430 , n59431 , n59432 , n59433 , n59434 , n59435 , n59436 , n59437 , n59438 , n59439 , n59440 , n59441 , n59442 , n59443 , n59444 , n59445 , n59446 , n59447 , n59448 , n59449 , n59450 , n59451 , n59452 , n59453 , n59454 , n59455 , n59456 , n59457 , n59458 , n59459 , n59460 , n59461 , n59462 , n59463 , n59464 , n59465 , n59466 , n59467 , n59468 , n59469 , n59470 , n59471 , n59472 , n59473 , n59474 , n59475 , n59476 , n59477 , n59478 , n59479 , n59480 , n59481 , n59482 , n59483 , n59484 , n59485 , n59486 , n59487 , n59488 , n59489 , n59490 , n59491 , n59492 , n59493 , n59494 , n59495 , n59496 , n59497 , n59498 , n59499 , n59500 , n59501 , n59502 , n59503 , n59504 , n59505 , n59506 , n59507 , n59508 , n59509 , n59510 , n59511 , n59512 , n59513 , n59514 , n59515 , n59516 , n59517 , n59518 , n59519 , n59520 , n59521 , n59522 , n59523 , n59524 , n59525 , n59526 , n59527 , n59528 , n59529 , n59530 , n59531 , n59532 , n59533 , n59534 , n59535 , n59536 , n59537 , n59538 , n59539 , n59540 , n59541 , n59542 , n59543 , n59544 , n59545 , n59546 , n59547 , n59548 , n59549 , n59550 , n59551 , n59552 , n59553 , n59554 , n59555 , n59556 , n59557 , n59558 , n59559 , n59560 , n59561 , n59562 , n59563 , n59564 , n59565 , n59566 , n59567 , n59568 , n59569 , n59570 , n59571 , n59572 , n59573 , n59574 , n59575 , n59576 , n59577 , n59578 , n59579 , n59580 , n59581 , n59582 , n59583 , n59584 , n59585 , n59586 , n59587 , n59588 , n59589 , n59590 , n59591 , n59592 , n59593 , n59594 , n59595 , n59596 , n59597 , n59598 , n59599 , n59600 , n59601 , n59602 , n59603 , n59604 , n59605 , n59606 , n59607 , n59608 , n59609 , n59610 , n59611 , n59612 , n59613 , n59614 , n59615 , n59616 , n59617 , n59618 , n59619 , n59620 , n59621 , n59622 , n59623 , n59624 , n59625 , n59626 , n59627 , n59628 , n59629 , n59630 , n59631 , n59632 , n59633 , n59634 , n59635 , n59636 , n59637 , n59638 , n59639 , n59640 , n59641 , n59642 , n59643 , n59644 , n59645 , n59646 , n59647 , n59648 , n59649 , n59650 , n59651 , n59652 , n59653 , n59654 , n59655 , n59656 , n59657 , n59658 , n59659 , n59660 , n59661 , n59662 , n59663 , n59664 , n59665 , n59666 , n59667 , n59668 , n59669 , n59670 , n59671 , n59672 , n59673 , n59674 , n59675 , n59676 , n59677 , n59678 , n59679 , n59680 , n59681 , n59682 , n59683 , n59684 , n59685 , n59686 , n59687 , n59688 , n59689 , n59690 , n59691 , n59692 , n59693 , n59694 , n59695 , n59696 , n59697 , n59698 , n59699 , n59700 , n59701 , n59702 , n59703 , n59704 , n59705 , n59706 , n59707 , n59708 , n59709 , n59710 , n59711 , n59712 , n59713 , n59714 , n59715 , n59716 , n59717 , n59718 , n59719 , n59720 , n59721 , n59722 , n59723 , n59724 , n59725 , n59726 , n59727 , n59728 , n59729 , n59730 , n59731 , n59732 , n59733 , n59734 , n59735 , n59736 , n59737 , n59738 , n59739 , n59740 , n59741 , n59742 , n59743 , n59744 , n59745 , n59746 , n59747 , n59748 , n59749 , n59750 , n59751 , n59752 , n59753 , n59754 , n59755 , n59756 , n59757 , n59758 , n59759 , n59760 , n59761 , n59762 , n59763 , n59764 , n59765 , n59766 , n59767 , n59768 , n59769 , n59770 , n59771 , n59772 , n59773 , n59774 , n59775 , n59776 , n59777 , n59778 , n59779 , n59780 , n59781 , n59782 , n59783 , n59784 , n59785 , n59786 , n59787 , n59788 , n59789 , n59790 , n59791 , n59792 , n59793 , n59794 , n59795 , n59796 , n59797 , n59798 , n59799 , n59800 , n59801 , n59802 , n59803 , n59804 , n59805 , n59806 , n59807 , n59808 , n59809 , n59810 , n59811 , n59812 , n59813 , n59814 , n59815 , n59816 , n59817 , n59818 , n59819 , n59820 , n59821 , n59822 , n59823 , n59824 , n59825 , n59826 , n59827 , n59828 , n59829 , n59830 , n59831 , n59832 , n59833 , n59834 , n59835 , n59836 , n59837 , n59838 , n59839 , n59840 , n59841 , n59842 , n59843 , n59844 , n59845 , n59846 , n59847 , n59848 , n59849 , n59850 , n59851 , n59852 , n59853 , n59854 , n59855 , n59856 , n59857 , n59858 , n59859 , n59860 , n59861 , n59862 , n59863 , n59864 , n59865 , n59866 , n59867 , n59868 , n59869 , n59870 , n59871 , n59872 , n59873 , n59874 , n59875 , n59876 , n59877 , n59878 , n59879 , n59880 , n59881 , n59882 , n59883 , n59884 , n59885 , n59886 , n59887 , n59888 , n59889 , n59890 , n59891 , n59892 , n59893 , n59894 , n59895 , n59896 , n59897 , n59898 , n59899 , n59900 , n59901 , n59902 , n59903 , n59904 , n59905 , n59906 , n59907 , n59908 , n59909 , n59910 , n59911 , n59912 , n59913 , n59914 , n59915 , n59916 , n59917 , n59918 , n59919 , n59920 , n59921 , n59922 , n59923 , n59924 , n59925 , n59926 , n59927 , n59928 , n59929 , n59930 , n59931 , n59932 , n59933 , n59934 , n59935 , n59936 , n59937 , n59938 , n59939 , n59940 , n59941 , n59942 , n59943 , n59944 , n59945 , n59946 , n59947 , n59948 , n59949 , n59950 , n59951 , n59952 , n59953 , n59954 , n59955 , n59956 , n59957 , n59958 , n59959 , n59960 , n59961 , n59962 , n59963 , n59964 , n59965 , n59966 , n59967 , n59968 , n59969 , n59970 , n59971 , n59972 , n59973 , n59974 , n59975 , n59976 , n59977 , n59978 , n59979 , n59980 , n59981 , n59982 , n59983 , n59984 , n59985 , n59986 , n59987 , n59988 , n59989 , n59990 , n59991 , n59992 , n59993 , n59994 , n59995 , n59996 , n59997 , n59998 , n59999 , n60000 , n60001 , n60002 , n60003 , n60004 , n60005 , n60006 , n60007 , n60008 , n60009 , n60010 , n60011 , n60012 , n60013 , n60014 , n60015 , n60016 , n60017 , n60018 , n60019 , n60020 , n60021 , n60022 , n60023 , n60024 , n60025 , n60026 , n60027 , n60028 , n60029 , n60030 , n60031 , n60032 , n60033 , n60034 , n60035 , n60036 , n60037 , n60038 , n60039 , n60040 , n60041 , n60042 , n60043 , n60044 , n60045 , n60046 , n60047 , n60048 , n60049 , n60050 , n60051 , n60052 , n60053 , n60054 , n60055 , n60056 , n60057 , n60058 , n60059 , n60060 , n60061 , n60062 , n60063 , n60064 , n60065 , n60066 , n60067 , n60068 , n60069 , n60070 , n60071 , n60072 , n60073 , n60074 , n60075 , n60076 , n60077 , n60078 , n60079 , n60080 , n60081 , n60082 , n60083 , n60084 , n60085 , n60086 , n60087 , n60088 , n60089 , n60090 , n60091 , n60092 , n60093 , n60094 , n60095 , n60096 , n60097 , n60098 , n60099 , n60100 , n60101 , n60102 , n60103 , n60104 , n60105 , n60106 , n60107 , n60108 , n60109 , n60110 , n60111 , n60112 , n60113 , n60114 , n60115 , n60116 , n60117 , n60118 , n60119 , n60120 , n60121 , n60122 , n60123 , n60124 , n60125 , n60126 , n60127 , n60128 , n60129 , n60130 , n60131 , n60132 , n60133 , n60134 , n60135 , n60136 , n60137 , n60138 , n60139 , n60140 , n60141 , n60142 , n60143 , n60144 , n60145 , n60146 , n60147 , n60148 , n60149 , n60150 , n60151 , n60152 , n60153 , n60154 , n60155 , n60156 , n60157 , n60158 , n60159 , n60160 , n60161 , n60162 , n60163 , n60164 , n60165 , n60166 , n60167 , n60168 , n60169 , n60170 , n60171 , n60172 , n60173 , n60174 , n60175 , n60176 , n60177 , n60178 , n60179 , n60180 , n60181 , n60182 , n60183 , n60184 , n60185 , n60186 , n60187 , n60188 , n60189 , n60190 , n60191 , n60192 , n60193 , n60194 , n60195 , n60196 , n60197 , n60198 , n60199 , n60200 , n60201 , n60202 , n60203 , n60204 , n60205 , n60206 , n60207 , n60208 , n60209 , n60210 , n60211 , n60212 , n60213 , n60214 , n60215 , n60216 , n60217 , n60218 , n60219 , n60220 , n60221 , n60222 , n60223 , n60224 , n60225 , n60226 , n60227 , n60228 , n60229 , n60230 , n60231 , n60232 , n60233 , n60234 , n60235 , n60236 , n60237 , n60238 , n60239 , n60240 , n60241 , n60242 , n60243 , n60244 , n60245 , n60246 , n60247 , n60248 , n60249 , n60250 , n60251 , n60252 , n60253 , n60254 , n60255 , n60256 , n60257 , n60258 , n60259 , n60260 , n60261 , n60262 , n60263 , n60264 , n60265 , n60266 , n60267 , n60268 , n60269 , n60270 , n60271 , n60272 , n60273 , n60274 , n60275 , n60276 , n60277 , n60278 , n60279 , n60280 , n60281 , n60282 , n60283 , n60284 , n60285 , n60286 , n60287 , n60288 , n60289 , n60290 , n60291 , n60292 , n60293 , n60294 , n60295 , n60296 , n60297 , n60298 , n60299 , n60300 , n60301 , n60302 , n60303 , n60304 , n60305 , n60306 , n60307 , n60308 , n60309 , n60310 , n60311 , n60312 , n60313 , n60314 , n60315 , n60316 , n60317 , n60318 , n60319 , n60320 , n60321 , n60322 , n60323 , n60324 , n60325 , n60326 , n60327 , n60328 , n60329 , n60330 , n60331 , n60332 , n60333 , n60334 , n60335 , n60336 , n60337 , n60338 , n60339 , n60340 , n60341 , n60342 , n60343 , n60344 , n60345 , n60346 , n60347 , n60348 , n60349 , n60350 , n60351 , n60352 , n60353 , n60354 , n60355 , n60356 , n60357 , n60358 , n60359 , n60360 , n60361 , n60362 , n60363 , n60364 , n60365 , n60366 , n60367 , n60368 , n60369 , n60370 , n60371 , n60372 , n60373 , n60374 , n60375 , n60376 , n60377 , n60378 , n60379 , n60380 , n60381 , n60382 , n60383 , n60384 , n60385 , n60386 , n60387 , n60388 , n60389 , n60390 , n60391 , n60392 , n60393 , n60394 , n60395 , n60396 , n60397 , n60398 , n60399 , n60400 , n60401 , n60402 , n60403 , n60404 , n60405 , n60406 , n60407 , n60408 , n60409 , n60410 , n60411 , n60412 , n60413 , n60414 , n60415 , n60416 , n60417 , n60418 , n60419 , n60420 , n60421 , n60422 , n60423 , n60424 , n60425 , n60426 , n60427 , n60428 , n60429 , n60430 , n60431 , n60432 , n60433 , n60434 , n60435 , n60436 , n60437 , n60438 , n60439 , n60440 , n60441 , n60442 , n60443 , n60444 , n60445 , n60446 , n60447 , n60448 , n60449 , n60450 , n60451 , n60452 , n60453 , n60454 , n60455 , n60456 , n60457 , n60458 , n60459 , n60460 , n60461 , n60462 , n60463 , n60464 , n60465 , n60466 , n60467 , n60468 , n60469 , n60470 , n60471 , n60472 , n60473 , n60474 , n60475 , n60476 , n60477 , n60478 , n60479 , n60480 , n60481 , n60482 , n60483 , n60484 , n60485 , n60486 , n60487 , n60488 , n60489 , n60490 , n60491 , n60492 , n60493 , n60494 , n60495 , n60496 , n60497 , n60498 , n60499 , n60500 , n60501 , n60502 , n60503 , n60504 , n60505 , n60506 , n60507 , n60508 , n60509 , n60510 , n60511 , n60512 , n60513 , n60514 , n60515 , n60516 , n60517 , n60518 , n60519 , n60520 , n60521 , n60522 , n60523 , n60524 , n60525 , n60526 , n60527 , n60528 , n60529 , n60530 , n60531 , n60532 , n60533 , n60534 , n60535 , n60536 , n60537 , n60538 , n60539 , n60540 , n60541 , n60542 , n60543 , n60544 , n60545 , n60546 , n60547 , n60548 , n60549 , n60550 , n60551 , n60552 , n60553 , n60554 , n60555 , n60556 , n60557 , n60558 , n60559 , n60560 , n60561 , n60562 , n60563 , n60564 , n60565 , n60566 , n60567 , n60568 , n60569 , n60570 , n60571 , n60572 , n60573 , n60574 , n60575 , n60576 , n60577 , n60578 , n60579 , n60580 , n60581 , n60582 , n60583 , n60584 , n60585 , n60586 , n60587 , n60588 , n60589 , n60590 , n60591 , n60592 , n60593 , n60594 , n60595 , n60596 , n60597 , n60598 , n60599 , n60600 , n60601 , n60602 , n60603 , n60604 , n60605 , n60606 , n60607 , n60608 , n60609 , n60610 , n60611 , n60612 , n60613 , n60614 , n60615 , n60616 , n60617 , n60618 , n60619 , n60620 , n60621 , n60622 , n60623 , n60624 , n60625 , n60626 , n60627 , n60628 , n60629 , n60630 , n60631 , n60632 , n60633 , n60634 , n60635 , n60636 , n60637 , n60638 , n60639 , n60640 , n60641 , n60642 , n60643 , n60644 , n60645 , n60646 , n60647 , n60648 , n60649 , n60650 , n60651 , n60652 , n60653 , n60654 , n60655 , n60656 , n60657 , n60658 , n60659 , n60660 , n60661 , n60662 , n60663 , n60664 , n60665 , n60666 , n60667 , n60668 , n60669 , n60670 , n60671 , n60672 , n60673 , n60674 , n60675 , n60676 , n60677 , n60678 , n60679 , n60680 , n60681 , n60682 , n60683 , n60684 , n60685 , n60686 , n60687 , n60688 , n60689 , n60690 , n60691 , n60692 , n60693 , n60694 , n60695 , n60696 , n60697 , n60698 , n60699 , n60700 , n60701 , n60702 , n60703 , n60704 , n60705 , n60706 , n60707 , n60708 , n60709 , n60710 , n60711 , n60712 , n60713 , n60714 , n60715 , n60716 , n60717 , n60718 , n60719 , n60720 , n60721 , n60722 , n60723 , n60724 , n60725 , n60726 , n60727 , n60728 , n60729 , n60730 , n60731 , n60732 , n60733 , n60734 , n60735 , n60736 , n60737 , n60738 , n60739 , n60740 , n60741 , n60742 , n60743 , n60744 , n60745 , n60746 , n60747 , n60748 , n60749 , n60750 , n60751 , n60752 , n60753 , n60754 , n60755 , n60756 , n60757 , n60758 , n60759 , n60760 , n60761 , n60762 , n60763 , n60764 , n60765 , n60766 , n60767 , n60768 , n60769 , n60770 , n60771 , n60772 , n60773 , n60774 , n60775 , n60776 , n60777 , n60778 , n60779 , n60780 , n60781 , n60782 , n60783 , n60784 , n60785 , n60786 , n60787 , n60788 , n60789 , n60790 , n60791 , n60792 , n60793 , n60794 , n60795 , n60796 , n60797 , n60798 , n60799 , n60800 , n60801 , n60802 , n60803 , n60804 , n60805 , n60806 , n60807 , n60808 , n60809 , n60810 , n60811 , n60812 , n60813 , n60814 , n60815 , n60816 , n60817 , n60818 , n60819 , n60820 , n60821 , n60822 , n60823 , n60824 , n60825 , n60826 , n60827 , n60828 , n60829 , n60830 , n60831 , n60832 , n60833 , n60834 , n60835 , n60836 , n60837 , n60838 , n60839 , n60840 , n60841 , n60842 , n60843 , n60844 , n60845 , n60846 , n60847 , n60848 , n60849 , n60850 , n60851 , n60852 , n60853 , n60854 , n60855 , n60856 , n60857 , n60858 , n60859 , n60860 , n60861 , n60862 , n60863 , n60864 , n60865 , n60866 , n60867 , n60868 , n60869 , n60870 , n60871 , n60872 , n60873 , n60874 , n60875 , n60876 , n60877 , n60878 , n60879 , n60880 , n60881 , n60882 , n60883 , n60884 , n60885 , n60886 , n60887 , n60888 , n60889 , n60890 , n60891 , n60892 , n60893 , n60894 , n60895 , n60896 , n60897 , n60898 , n60899 , n60900 , n60901 , n60902 , n60903 , n60904 , n60905 , n60906 , n60907 , n60908 , n60909 , n60910 , n60911 , n60912 , n60913 , n60914 , n60915 , n60916 , n60917 , n60918 , n60919 , n60920 , n60921 , n60922 , n60923 , n60924 , n60925 , n60926 , n60927 , n60928 , n60929 , n60930 , n60931 , n60932 , n60933 , n60934 , n60935 , n60936 , n60937 , n60938 , n60939 , n60940 , n60941 , n60942 , n60943 , n60944 , n60945 , n60946 , n60947 , n60948 , n60949 , n60950 , n60951 , n60952 , n60953 , n60954 , n60955 , n60956 , n60957 , n60958 , n60959 , n60960 , n60961 , n60962 , n60963 , n60964 , n60965 , n60966 , n60967 , n60968 , n60969 , n60970 , n60971 , n60972 , n60973 , n60974 , n60975 , n60976 , n60977 , n60978 , n60979 , n60980 , n60981 , n60982 , n60983 , n60984 , n60985 , n60986 , n60987 , n60988 , n60989 , n60990 , n60991 , n60992 , n60993 , n60994 , n60995 , n60996 , n60997 , n60998 , n60999 , n61000 , n61001 , n61002 , n61003 , n61004 , n61005 , n61006 , n61007 , n61008 , n61009 , n61010 , n61011 , n61012 , n61013 , n61014 , n61015 , n61016 , n61017 , n61018 , n61019 , n61020 , n61021 , n61022 , n61023 , n61024 , n61025 , n61026 , n61027 , n61028 , n61029 , n61030 , n61031 , n61032 , n61033 , n61034 , n61035 , n61036 , n61037 , n61038 , n61039 , n61040 , n61041 , n61042 , n61043 , n61044 , n61045 , n61046 , n61047 , n61048 , n61049 , n61050 , n61051 , n61052 , n61053 , n61054 , n61055 , n61056 , n61057 , n61058 , n61059 , n61060 , n61061 , n61062 , n61063 , n61064 , n61065 , n61066 , n61067 , n61068 , n61069 , n61070 , n61071 , n61072 , n61073 , n61074 , n61075 , n61076 , n61077 , n61078 , n61079 , n61080 , n61081 , n61082 , n61083 , n61084 , n61085 , n61086 , n61087 , n61088 , n61089 , n61090 , n61091 , n61092 , n61093 , n61094 , n61095 , n61096 , n61097 , n61098 , n61099 , n61100 , n61101 , n61102 , n61103 , n61104 , n61105 , n61106 , n61107 , n61108 , n61109 , n61110 , n61111 , n61112 , n61113 , n61114 , n61115 , n61116 , n61117 , n61118 , n61119 , n61120 , n61121 , n61122 , n61123 , n61124 , n61125 , n61126 , n61127 , n61128 , n61129 , n61130 , n61131 , n61132 , n61133 , n61134 , n61135 , n61136 , n61137 , n61138 , n61139 , n61140 , n61141 , n61142 , n61143 , n61144 , n61145 , n61146 , n61147 , n61148 , n61149 , n61150 , n61151 , n61152 , n61153 , n61154 , n61155 , n61156 , n61157 , n61158 , n61159 , n61160 , n61161 , n61162 , n61163 , n61164 , n61165 , n61166 , n61167 , n61168 , n61169 , n61170 , n61171 , n61172 , n61173 , n61174 , n61175 , n61176 , n61177 , n61178 , n61179 , n61180 , n61181 , n61182 , n61183 , n61184 , n61185 , n61186 , n61187 , n61188 , n61189 , n61190 , n61191 , n61192 , n61193 , n61194 , n61195 , n61196 , n61197 , n61198 , n61199 , n61200 , n61201 , n61202 , n61203 , n61204 , n61205 , n61206 , n61207 , n61208 , n61209 , n61210 , n61211 , n61212 , n61213 , n61214 , n61215 , n61216 , n61217 , n61218 , n61219 , n61220 , n61221 , n61222 , n61223 , n61224 , n61225 , n61226 , n61227 , n61228 , n61229 , n61230 , n61231 , n61232 , n61233 , n61234 , n61235 , n61236 , n61237 , n61238 , n61239 , n61240 , n61241 , n61242 , n61243 , n61244 , n61245 , n61246 , n61247 , n61248 , n61249 , n61250 , n61251 , n61252 , n61253 , n61254 , n61255 , n61256 , n61257 , n61258 , n61259 , n61260 , n61261 , n61262 , n61263 , n61264 , n61265 , n61266 , n61267 , n61268 , n61269 , n61270 , n61271 , n61272 , n61273 , n61274 , n61275 , n61276 , n61277 , n61278 , n61279 , n61280 , n61281 , n61282 , n61283 , n61284 , n61285 , n61286 , n61287 , n61288 , n61289 , n61290 , n61291 , n61292 , n61293 , n61294 , n61295 , n61296 , n61297 , n61298 , n61299 , n61300 , n61301 , n61302 , n61303 , n61304 , n61305 , n61306 , n61307 , n61308 , n61309 , n61310 , n61311 , n61312 , n61313 , n61314 , n61315 , n61316 , n61317 , n61318 , n61319 , n61320 , n61321 , n61322 , n61323 , n61324 , n61325 , n61326 , n61327 , n61328 , n61329 , n61330 , n61331 , n61332 , n61333 , n61334 , n61335 , n61336 , n61337 , n61338 , n61339 , n61340 , n61341 , n61342 , n61343 , n61344 , n61345 , n61346 , n61347 , n61348 , n61349 , n61350 , n61351 , n61352 , n61353 , n61354 , n61355 , n61356 , n61357 , n61358 , n61359 , n61360 , n61361 , n61362 , n61363 , n61364 , n61365 , n61366 , n61367 , n61368 , n61369 , n61370 , n61371 , n61372 , n61373 , n61374 , n61375 , n61376 , n61377 , n61378 , n61379 , n61380 , n61381 , n61382 , n61383 , n61384 , n61385 , n61386 , n61387 , n61388 , n61389 , n61390 , n61391 , n61392 , n61393 , n61394 , n61395 , n61396 , n61397 , n61398 , n61399 , n61400 , n61401 , n61402 , n61403 , n61404 , n61405 , n61406 , n61407 , n61408 , n61409 , n61410 , n61411 , n61412 , n61413 , n61414 , n61415 , n61416 , n61417 , n61418 , n61419 , n61420 , n61421 , n61422 , n61423 , n61424 , n61425 , n61426 , n61427 , n61428 , n61429 , n61430 , n61431 , n61432 , n61433 , n61434 , n61435 , n61436 , n61437 , n61438 , n61439 , n61440 , n61441 , n61442 , n61443 , n61444 , n61445 , n61446 , n61447 , n61448 , n61449 , n61450 , n61451 , n61452 , n61453 , n61454 , n61455 , n61456 , n61457 , n61458 , n61459 , n61460 , n61461 , n61462 , n61463 , n61464 , n61465 , n61466 , n61467 , n61468 , n61469 , n61470 , n61471 , n61472 , n61473 , n61474 , n61475 , n61476 , n61477 , n61478 , n61479 , n61480 , n61481 , n61482 , n61483 , n61484 , n61485 , n61486 , n61487 , n61488 , n61489 , n61490 , n61491 , n61492 , n61493 , n61494 , n61495 , n61496 , n61497 , n61498 , n61499 , n61500 , n61501 , n61502 , n61503 , n61504 , n61505 , n61506 , n61507 , n61508 , n61509 , n61510 , n61511 , n61512 , n61513 , n61514 , n61515 , n61516 , n61517 , n61518 , n61519 , n61520 , n61521 , n61522 , n61523 , n61524 , n61525 , n61526 , n61527 , n61528 , n61529 , n61530 , n61531 , n61532 , n61533 , n61534 , n61535 , n61536 , n61537 , n61538 , n61539 , n61540 , n61541 , n61542 , n61543 , n61544 , n61545 , n61546 , n61547 , n61548 , n61549 , n61550 , n61551 , n61552 , n61553 , n61554 , n61555 , n61556 , n61557 , n61558 , n61559 , n61560 , n61561 , n61562 , n61563 , n61564 , n61565 , n61566 , n61567 , n61568 , n61569 , n61570 , n61571 , n61572 , n61573 , n61574 , n61575 , n61576 , n61577 , n61578 , n61579 , n61580 , n61581 , n61582 , n61583 , n61584 , n61585 , n61586 , n61587 , n61588 , n61589 , n61590 , n61591 , n61592 , n61593 , n61594 , n61595 , n61596 , n61597 , n61598 , n61599 , n61600 , n61601 , n61602 , n61603 , n61604 , n61605 , n61606 , n61607 , n61608 , n61609 , n61610 , n61611 , n61612 , n61613 , n61614 , n61615 , n61616 , n61617 , n61618 , n61619 , n61620 , n61621 , n61622 , n61623 , n61624 , n61625 , n61626 , n61627 , n61628 , n61629 , n61630 , n61631 , n61632 , n61633 , n61634 , n61635 , n61636 , n61637 , n61638 , n61639 , n61640 , n61641 , n61642 , n61643 , n61644 , n61645 , n61646 , n61647 , n61648 , n61649 , n61650 , n61651 , n61652 , n61653 , n61654 , n61655 , n61656 , n61657 , n61658 , n61659 , n61660 , n61661 , n61662 , n61663 , n61664 , n61665 , n61666 , n61667 , n61668 , n61669 , n61670 , n61671 , n61672 , n61673 , n61674 , n61675 , n61676 , n61677 , n61678 , n61679 , n61680 , n61681 , n61682 , n61683 , n61684 , n61685 , n61686 , n61687 , n61688 , n61689 , n61690 , n61691 , n61692 , n61693 , n61694 , n61695 , n61696 , n61697 , n61698 , n61699 , n61700 , n61701 , n61702 , n61703 , n61704 , n61705 , n61706 , n61707 , n61708 , n61709 , n61710 , n61711 , n61712 , n61713 , n61714 , n61715 , n61716 , n61717 , n61718 , n61719 , n61720 , n61721 , n61722 , n61723 , n61724 , n61725 , n61726 , n61727 , n61728 , n61729 , n61730 , n61731 , n61732 , n61733 , n61734 , n61735 , n61736 , n61737 , n61738 , n61739 , n61740 , n61741 , n61742 , n61743 , n61744 , n61745 , n61746 , n61747 , n61748 , n61749 , n61750 , n61751 , n61752 , n61753 , n61754 , n61755 , n61756 , n61757 , n61758 , n61759 , n61760 , n61761 , n61762 , n61763 , n61764 , n61765 , n61766 , n61767 , n61768 , n61769 , n61770 , n61771 , n61772 , n61773 , n61774 , n61775 , n61776 , n61777 , n61778 , n61779 , n61780 , n61781 , n61782 , n61783 , n61784 , n61785 , n61786 , n61787 , n61788 , n61789 , n61790 , n61791 , n61792 , n61793 , n61794 , n61795 , n61796 , n61797 , n61798 , n61799 , n61800 , n61801 , n61802 , n61803 , n61804 , n61805 , n61806 , n61807 , n61808 , n61809 , n61810 , n61811 , n61812 , n61813 , n61814 , n61815 , n61816 , n61817 , n61818 , n61819 , n61820 , n61821 , n61822 , n61823 , n61824 , n61825 , n61826 , n61827 , n61828 , n61829 , n61830 , n61831 , n61832 , n61833 , n61834 , n61835 , n61836 , n61837 , n61838 , n61839 , n61840 , n61841 , n61842 , n61843 , n61844 , n61845 , n61846 , n61847 , n61848 , n61849 , n61850 , n61851 , n61852 , n61853 , n61854 , n61855 , n61856 , n61857 , n61858 , n61859 , n61860 , n61861 , n61862 , n61863 , n61864 , n61865 , n61866 , n61867 , n61868 , n61869 , n61870 , n61871 , n61872 , n61873 , n61874 , n61875 , n61876 , n61877 , n61878 , n61879 , n61880 , n61881 , n61882 , n61883 , n61884 , n61885 , n61886 , n61887 , n61888 , n61889 , n61890 , n61891 , n61892 , n61893 , n61894 , n61895 , n61896 , n61897 , n61898 , n61899 , n61900 , n61901 , n61902 , n61903 , n61904 , n61905 , n61906 , n61907 , n61908 , n61909 , n61910 , n61911 , n61912 , n61913 , n61914 , n61915 , n61916 , n61917 , n61918 , n61919 , n61920 , n61921 , n61922 , n61923 , n61924 , n61925 , n61926 , n61927 , n61928 , n61929 , n61930 , n61931 , n61932 , n61933 , n61934 , n61935 , n61936 , n61937 , n61938 , n61939 , n61940 , n61941 , n61942 , n61943 , n61944 , n61945 , n61946 , n61947 , n61948 , n61949 , n61950 , n61951 , n61952 , n61953 , n61954 , n61955 , n61956 , n61957 , n61958 , n61959 , n61960 , n61961 , n61962 , n61963 , n61964 , n61965 , n61966 , n61967 , n61968 , n61969 , n61970 , n61971 , n61972 , n61973 , n61974 , n61975 , n61976 , n61977 , n61978 , n61979 , n61980 , n61981 , n61982 , n61983 , n61984 , n61985 , n61986 , n61987 , n61988 , n61989 , n61990 , n61991 , n61992 , n61993 , n61994 , n61995 , n61996 , n61997 , n61998 , n61999 , n62000 , n62001 , n62002 , n62003 , n62004 , n62005 , n62006 , n62007 , n62008 , n62009 , n62010 , n62011 , n62012 , n62013 , n62014 , n62015 , n62016 , n62017 , n62018 , n62019 , n62020 , n62021 , n62022 , n62023 , n62024 , n62025 , n62026 , n62027 , n62028 , n62029 , n62030 , n62031 , n62032 , n62033 , n62034 , n62035 , n62036 , n62037 , n62038 , n62039 , n62040 , n62041 , n62042 , n62043 , n62044 , n62045 , n62046 , n62047 , n62048 , n62049 , n62050 , n62051 , n62052 , n62053 , n62054 , n62055 , n62056 , n62057 , n62058 , n62059 , n62060 , n62061 , n62062 , n62063 , n62064 , n62065 , n62066 , n62067 , n62068 , n62069 , n62070 , n62071 , n62072 , n62073 , n62074 , n62075 , n62076 , n62077 , n62078 , n62079 , n62080 , n62081 , n62082 , n62083 , n62084 , n62085 , n62086 , n62087 , n62088 , n62089 , n62090 , n62091 , n62092 , n62093 , n62094 , n62095 , n62096 , n62097 , n62098 , n62099 , n62100 , n62101 , n62102 , n62103 , n62104 , n62105 , n62106 , n62107 , n62108 , n62109 , n62110 , n62111 , n62112 , n62113 , n62114 , n62115 , n62116 , n62117 , n62118 , n62119 , n62120 , n62121 , n62122 , n62123 , n62124 , n62125 , n62126 , n62127 , n62128 , n62129 , n62130 , n62131 , n62132 , n62133 , n62134 , n62135 , n62136 , n62137 , n62138 , n62139 , n62140 , n62141 , n62142 , n62143 , n62144 , n62145 , n62146 , n62147 , n62148 , n62149 , n62150 , n62151 , n62152 , n62153 , n62154 , n62155 , n62156 , n62157 , n62158 , n62159 , n62160 , n62161 , n62162 , n62163 , n62164 , n62165 , n62166 , n62167 , n62168 , n62169 , n62170 , n62171 , n62172 , n62173 , n62174 , n62175 , n62176 , n62177 , n62178 , n62179 , n62180 , n62181 , n62182 , n62183 , n62184 , n62185 , n62186 , n62187 , n62188 , n62189 , n62190 , n62191 , n62192 , n62193 , n62194 , n62195 , n62196 , n62197 , n62198 , n62199 , n62200 , n62201 , n62202 , n62203 , n62204 , n62205 , n62206 , n62207 , n62208 , n62209 , n62210 , n62211 , n62212 , n62213 , n62214 , n62215 , n62216 , n62217 , n62218 , n62219 , n62220 , n62221 , n62222 , n62223 , n62224 , n62225 , n62226 , n62227 , n62228 , n62229 , n62230 , n62231 , n62232 , n62233 , n62234 , n62235 , n62236 , n62237 , n62238 , n62239 , n62240 , n62241 , n62242 , n62243 , n62244 , n62245 , n62246 , n62247 , n62248 , n62249 , n62250 , n62251 , n62252 , n62253 , n62254 , n62255 , n62256 , n62257 , n62258 , n62259 , n62260 , n62261 , n62262 , n62263 , n62264 , n62265 , n62266 , n62267 , n62268 , n62269 , n62270 , n62271 , n62272 , n62273 , n62274 , n62275 , n62276 , n62277 , n62278 , n62279 , n62280 , n62281 , n62282 , n62283 , n62284 , n62285 , n62286 , n62287 , n62288 , n62289 , n62290 , n62291 , n62292 , n62293 , n62294 , n62295 , n62296 , n62297 , n62298 , n62299 , n62300 , n62301 , n62302 , n62303 , n62304 , n62305 , n62306 , n62307 , n62308 , n62309 , n62310 , n62311 , n62312 , n62313 , n62314 , n62315 , n62316 , n62317 , n62318 , n62319 , n62320 , n62321 , n62322 , n62323 , n62324 , n62325 , n62326 , n62327 , n62328 , n62329 , n62330 , n62331 , n62332 , n62333 , n62334 , n62335 , n62336 , n62337 , n62338 , n62339 , n62340 , n62341 , n62342 , n62343 , n62344 , n62345 , n62346 , n62347 , n62348 , n62349 , n62350 , n62351 , n62352 , n62353 , n62354 , n62355 , n62356 , n62357 , n62358 , n62359 , n62360 , n62361 , n62362 , n62363 , n62364 , n62365 , n62366 , n62367 , n62368 , n62369 , n62370 , n62371 , n62372 , n62373 , n62374 , n62375 , n62376 , n62377 , n62378 , n62379 , n62380 , n62381 , n62382 , n62383 , n62384 , n62385 , n62386 , n62387 , n62388 , n62389 , n62390 , n62391 , n62392 , n62393 , n62394 , n62395 , n62396 , n62397 , n62398 , n62399 , n62400 , n62401 , n62402 , n62403 , n62404 , n62405 , n62406 , n62407 , n62408 , n62409 , n62410 , n62411 , n62412 , n62413 , n62414 , n62415 , n62416 , n62417 , n62418 , n62419 , n62420 , n62421 , n62422 , n62423 , n62424 , n62425 , n62426 , n62427 , n62428 , n62429 , n62430 , n62431 , n62432 , n62433 , n62434 , n62435 , n62436 , n62437 , n62438 , n62439 , n62440 , n62441 , n62442 , n62443 , n62444 , n62445 , n62446 , n62447 , n62448 , n62449 , n62450 , n62451 , n62452 , n62453 , n62454 , n62455 , n62456 , n62457 , n62458 , n62459 , n62460 , n62461 , n62462 , n62463 , n62464 , n62465 , n62466 , n62467 , n62468 , n62469 , n62470 , n62471 , n62472 , n62473 , n62474 , n62475 , n62476 , n62477 , n62478 , n62479 , n62480 , n62481 , n62482 , n62483 , n62484 , n62485 , n62486 , n62487 , n62488 , n62489 , n62490 , n62491 , n62492 , n62493 , n62494 , n62495 , n62496 , n62497 , n62498 , n62499 , n62500 , n62501 , n62502 , n62503 , n62504 , n62505 , n62506 , n62507 , n62508 , n62509 , n62510 , n62511 , n62512 , n62513 , n62514 , n62515 , n62516 , n62517 , n62518 , n62519 , n62520 , n62521 , n62522 , n62523 , n62524 , n62525 , n62526 , n62527 , n62528 , n62529 , n62530 , n62531 , n62532 , n62533 , n62534 , n62535 , n62536 , n62537 , n62538 , n62539 , n62540 , n62541 , n62542 , n62543 , n62544 , n62545 , n62546 , n62547 , n62548 , n62549 , n62550 , n62551 , n62552 , n62553 , n62554 , n62555 , n62556 , n62557 , n62558 , n62559 , n62560 , n62561 , n62562 , n62563 , n62564 , n62565 , n62566 , n62567 , n62568 , n62569 , n62570 , n62571 , n62572 , n62573 , n62574 , n62575 , n62576 , n62577 , n62578 , n62579 , n62580 , n62581 , n62582 , n62583 , n62584 , n62585 , n62586 , n62587 , n62588 , n62589 , n62590 , n62591 , n62592 , n62593 , n62594 , n62595 , n62596 , n62597 , n62598 , n62599 , n62600 , n62601 , n62602 , n62603 , n62604 , n62605 , n62606 , n62607 , n62608 , n62609 , n62610 , n62611 , n62612 , n62613 , n62614 , n62615 , n62616 , n62617 , n62618 , n62619 , n62620 , n62621 , n62622 , n62623 , n62624 , n62625 , n62626 , n62627 , n62628 , n62629 , n62630 , n62631 , n62632 , n62633 , n62634 , n62635 , n62636 , n62637 , n62638 , n62639 , n62640 , n62641 , n62642 , n62643 , n62644 , n62645 , n62646 , n62647 , n62648 , n62649 , n62650 , n62651 , n62652 , n62653 , n62654 , n62655 , n62656 , n62657 , n62658 , n62659 , n62660 , n62661 , n62662 , n62663 , n62664 , n62665 , n62666 , n62667 , n62668 , n62669 , n62670 , n62671 , n62672 , n62673 , n62674 , n62675 , n62676 , n62677 , n62678 , n62679 , n62680 , n62681 , n62682 , n62683 , n62684 , n62685 , n62686 , n62687 , n62688 , n62689 , n62690 , n62691 , n62692 , n62693 , n62694 , n62695 , n62696 , n62697 , n62698 , n62699 , n62700 , n62701 , n62702 , n62703 , n62704 , n62705 , n62706 , n62707 , n62708 , n62709 , n62710 , n62711 , n62712 , n62713 , n62714 , n62715 , n62716 , n62717 , n62718 , n62719 , n62720 , n62721 , n62722 , n62723 , n62724 , n62725 , n62726 , n62727 , n62728 , n62729 , n62730 , n62731 , n62732 , n62733 , n62734 , n62735 , n62736 , n62737 , n62738 , n62739 , n62740 , n62741 , n62742 , n62743 , n62744 , n62745 , n62746 , n62747 , n62748 , n62749 , n62750 , n62751 , n62752 , n62753 , n62754 , n62755 , n62756 , n62757 , n62758 , n62759 , n62760 , n62761 , n62762 , n62763 , n62764 , n62765 , n62766 , n62767 , n62768 , n62769 , n62770 , n62771 , n62772 , n62773 , n62774 , n62775 , n62776 , n62777 , n62778 , n62779 , n62780 , n62781 , n62782 , n62783 , n62784 , n62785 , n62786 , n62787 , n62788 , n62789 , n62790 , n62791 , n62792 , n62793 , n62794 , n62795 , n62796 , n62797 , n62798 , n62799 , n62800 , n62801 , n62802 , n62803 , n62804 , n62805 , n62806 , n62807 , n62808 , n62809 , n62810 , n62811 , n62812 , n62813 , n62814 , n62815 , n62816 , n62817 , n62818 , n62819 , n62820 , n62821 , n62822 , n62823 , n62824 , n62825 , n62826 , n62827 , n62828 , n62829 , n62830 , n62831 , n62832 , n62833 , n62834 , n62835 , n62836 , n62837 , n62838 , n62839 , n62840 , n62841 , n62842 , n62843 , n62844 , n62845 , n62846 , n62847 , n62848 , n62849 , n62850 , n62851 , n62852 , n62853 , n62854 , n62855 , n62856 , n62857 , n62858 , n62859 , n62860 , n62861 , n62862 , n62863 , n62864 , n62865 , n62866 , n62867 , n62868 , n62869 , n62870 , n62871 , n62872 , n62873 , n62874 , n62875 , n62876 , n62877 , n62878 , n62879 , n62880 , n62881 , n62882 , n62883 , n62884 , n62885 , n62886 , n62887 , n62888 , n62889 , n62890 , n62891 , n62892 , n62893 , n62894 , n62895 , n62896 , n62897 , n62898 , n62899 , n62900 , n62901 , n62902 , n62903 , n62904 , n62905 , n62906 , n62907 , n62908 , n62909 , n62910 , n62911 , n62912 , n62913 , n62914 , n62915 , n62916 , n62917 , n62918 , n62919 , n62920 , n62921 , n62922 , n62923 , n62924 , n62925 , n62926 , n62927 , n62928 , n62929 , n62930 , n62931 , n62932 , n62933 , n62934 , n62935 , n62936 , n62937 , n62938 , n62939 , n62940 , n62941 , n62942 , n62943 , n62944 , n62945 , n62946 , n62947 , n62948 , n62949 , n62950 , n62951 , n62952 , n62953 , n62954 , n62955 , n62956 , n62957 , n62958 , n62959 , n62960 , n62961 , n62962 , n62963 , n62964 , n62965 , n62966 , n62967 , n62968 , n62969 , n62970 , n62971 , n62972 , n62973 , n62974 , n62975 , n62976 , n62977 , n62978 , n62979 , n62980 , n62981 , n62982 , n62983 , n62984 , n62985 , n62986 , n62987 , n62988 , n62989 , n62990 , n62991 , n62992 , n62993 , n62994 , n62995 , n62996 , n62997 , n62998 , n62999 , n63000 , n63001 , n63002 , n63003 , n63004 , n63005 , n63006 , n63007 , n63008 , n63009 , n63010 , n63011 , n63012 , n63013 , n63014 , n63015 , n63016 , n63017 , n63018 , n63019 , n63020 , n63021 , n63022 , n63023 , n63024 , n63025 , n63026 , n63027 , n63028 , n63029 , n63030 , n63031 , n63032 , n63033 , n63034 , n63035 , n63036 , n63037 , n63038 , n63039 , n63040 , n63041 , n63042 , n63043 , n63044 , n63045 , n63046 , n63047 , n63048 , n63049 , n63050 , n63051 , n63052 , n63053 , n63054 , n63055 , n63056 , n63057 , n63058 , n63059 , n63060 , n63061 , n63062 , n63063 , n63064 , n63065 , n63066 , n63067 , n63068 , n63069 , n63070 , n63071 , n63072 , n63073 , n63074 , n63075 , n63076 , n63077 , n63078 , n63079 , n63080 , n63081 , n63082 , n63083 , n63084 , n63085 , n63086 , n63087 , n63088 , n63089 , n63090 , n63091 , n63092 , n63093 , n63094 , n63095 , n63096 , n63097 , n63098 , n63099 , n63100 , n63101 , n63102 , n63103 , n63104 , n63105 , n63106 , n63107 , n63108 , n63109 , n63110 , n63111 , n63112 , n63113 , n63114 , n63115 , n63116 , n63117 , n63118 , n63119 , n63120 , n63121 , n63122 , n63123 , n63124 , n63125 , n63126 , n63127 , n63128 , n63129 , n63130 , n63131 , n63132 , n63133 , n63134 , n63135 , n63136 , n63137 , n63138 , n63139 , n63140 , n63141 , n63142 , n63143 , n63144 , n63145 , n63146 , n63147 , n63148 , n63149 , n63150 , n63151 , n63152 , n63153 , n63154 , n63155 , n63156 , n63157 , n63158 , n63159 , n63160 , n63161 , n63162 , n63163 , n63164 , n63165 , n63166 , n63167 , n63168 , n63169 , n63170 , n63171 , n63172 , n63173 , n63174 , n63175 , n63176 , n63177 , n63178 , n63179 , n63180 , n63181 , n63182 , n63183 , n63184 , n63185 , n63186 , n63187 , n63188 , n63189 , n63190 , n63191 , n63192 , n63193 , n63194 , n63195 , n63196 , n63197 , n63198 , n63199 , n63200 , n63201 , n63202 , n63203 , n63204 , n63205 , n63206 , n63207 , n63208 , n63209 , n63210 , n63211 , n63212 , n63213 , n63214 , n63215 , n63216 , n63217 , n63218 , n63219 , n63220 , n63221 , n63222 , n63223 , n63224 , n63225 , n63226 , n63227 , n63228 , n63229 , n63230 , n63231 , n63232 , n63233 , n63234 , n63235 , n63236 , n63237 , n63238 , n63239 , n63240 , n63241 , n63242 , n63243 , n63244 , n63245 , n63246 , n63247 , n63248 , n63249 , n63250 , n63251 , n63252 , n63253 , n63254 , n63255 , n63256 , n63257 , n63258 , n63259 , n63260 , n63261 , n63262 , n63263 , n63264 , n63265 , n63266 , n63267 , n63268 , n63269 , n63270 , n63271 , n63272 , n63273 , n63274 , n63275 , n63276 , n63277 , n63278 , n63279 , n63280 , n63281 , n63282 , n63283 , n63284 , n63285 , n63286 , n63287 , n63288 , n63289 , n63290 , n63291 , n63292 , n63293 , n63294 , n63295 , n63296 , n63297 , n63298 , n63299 , n63300 , n63301 , n63302 , n63303 , n63304 , n63305 , n63306 , n63307 , n63308 , n63309 , n63310 , n63311 , n63312 , n63313 , n63314 , n63315 , n63316 , n63317 , n63318 , n63319 , n63320 , n63321 , n63322 , n63323 , n63324 , n63325 , n63326 , n63327 , n63328 , n63329 , n63330 , n63331 , n63332 , n63333 , n63334 , n63335 , n63336 , n63337 , n63338 , n63339 , n63340 , n63341 , n63342 , n63343 , n63344 , n63345 , n63346 , n63347 , n63348 , n63349 , n63350 , n63351 , n63352 , n63353 , n63354 , n63355 , n63356 , n63357 , n63358 , n63359 , n63360 , n63361 , n63362 , n63363 , n63364 , n63365 , n63366 , n63367 , n63368 , n63369 , n63370 , n63371 , n63372 , n63373 , n63374 , n63375 , n63376 , n63377 , n63378 , n63379 , n63380 , n63381 , n63382 , n63383 , n63384 , n63385 , n63386 , n63387 , n63388 , n63389 , n63390 , n63391 , n63392 , n63393 , n63394 , n63395 , n63396 , n63397 , n63398 , n63399 , n63400 , n63401 , n63402 , n63403 , n63404 , n63405 , n63406 , n63407 , n63408 , n63409 , n63410 , n63411 , n63412 , n63413 , n63414 , n63415 , n63416 , n63417 , n63418 , n63419 , n63420 , n63421 , n63422 , n63423 , n63424 , n63425 , n63426 , n63427 , n63428 , n63429 , n63430 , n63431 , n63432 , n63433 , n63434 , n63435 , n63436 , n63437 , n63438 , n63439 , n63440 , n63441 , n63442 , n63443 , n63444 , n63445 , n63446 , n63447 , n63448 , n63449 , n63450 , n63451 , n63452 , n63453 , n63454 , n63455 , n63456 , n63457 , n63458 , n63459 , n63460 , n63461 , n63462 , n63463 , n63464 , n63465 , n63466 , n63467 , n63468 , n63469 , n63470 , n63471 , n63472 , n63473 , n63474 , n63475 , n63476 , n63477 , n63478 , n63479 , n63480 , n63481 , n63482 , n63483 , n63484 , n63485 , n63486 , n63487 , n63488 , n63489 , n63490 , n63491 , n63492 , n63493 , n63494 , n63495 , n63496 , n63497 , n63498 , n63499 , n63500 , n63501 , n63502 , n63503 , n63504 , n63505 , n63506 , n63507 , n63508 , n63509 , n63510 , n63511 , n63512 , n63513 , n63514 , n63515 , n63516 , n63517 , n63518 , n63519 , n63520 , n63521 , n63522 , n63523 , n63524 , n63525 , n63526 , n63527 , n63528 , n63529 , n63530 , n63531 , n63532 , n63533 , n63534 , n63535 , n63536 , n63537 , n63538 , n63539 , n63540 , n63541 , n63542 , n63543 , n63544 , n63545 , n63546 , n63547 , n63548 , n63549 , n63550 , n63551 , n63552 , n63553 , n63554 , n63555 , n63556 , n63557 , n63558 , n63559 , n63560 , n63561 , n63562 , n63563 , n63564 , n63565 , n63566 , n63567 , n63568 , n63569 , n63570 , n63571 , n63572 , n63573 , n63574 , n63575 , n63576 , n63577 , n63578 , n63579 , n63580 , n63581 , n63582 , n63583 , n63584 , n63585 , n63586 , n63587 , n63588 , n63589 , n63590 , n63591 , n63592 , n63593 , n63594 , n63595 , n63596 , n63597 , n63598 , n63599 , n63600 , n63601 , n63602 , n63603 , n63604 , n63605 , n63606 , n63607 , n63608 , n63609 , n63610 , n63611 , n63612 , n63613 , n63614 , n63615 , n63616 , n63617 , n63618 , n63619 , n63620 , n63621 , n63622 , n63623 , n63624 , n63625 , n63626 , n63627 , n63628 , n63629 , n63630 , n63631 , n63632 , n63633 , n63634 , n63635 , n63636 , n63637 , n63638 , n63639 , n63640 , n63641 , n63642 , n63643 , n63644 , n63645 , n63646 , n63647 , n63648 , n63649 , n63650 , n63651 , n63652 , n63653 , n63654 , n63655 , n63656 , n63657 , n63658 , n63659 , n63660 , n63661 , n63662 , n63663 , n63664 , n63665 , n63666 , n63667 , n63668 , n63669 , n63670 , n63671 , n63672 , n63673 , n63674 , n63675 , n63676 , n63677 , n63678 , n63679 , n63680 , n63681 , n63682 , n63683 , n63684 , n63685 , n63686 , n63687 , n63688 , n63689 , n63690 , n63691 , n63692 , n63693 , n63694 , n63695 , n63696 , n63697 , n63698 , n63699 , n63700 , n63701 , n63702 , n63703 , n63704 , n63705 , n63706 , n63707 , n63708 , n63709 , n63710 , n63711 , n63712 , n63713 , n63714 , n63715 , n63716 , n63717 , n63718 , n63719 , n63720 , n63721 , n63722 , n63723 , n63724 , n63725 , n63726 , n63727 , n63728 , n63729 , n63730 , n63731 , n63732 , n63733 , n63734 , n63735 , n63736 , n63737 , n63738 , n63739 , n63740 , n63741 , n63742 , n63743 , n63744 , n63745 , n63746 , n63747 , n63748 , n63749 , n63750 , n63751 , n63752 , n63753 , n63754 , n63755 , n63756 , n63757 , n63758 , n63759 , n63760 , n63761 , n63762 , n63763 , n63764 , n63765 , n63766 , n63767 , n63768 , n63769 , n63770 , n63771 , n63772 , n63773 , n63774 , n63775 , n63776 , n63777 , n63778 , n63779 , n63780 , n63781 , n63782 , n63783 , n63784 , n63785 , n63786 , n63787 , n63788 , n63789 , n63790 , n63791 , n63792 , n63793 , n63794 , n63795 , n63796 , n63797 , n63798 , n63799 , n63800 , n63801 , n63802 , n63803 , n63804 , n63805 , n63806 , n63807 , n63808 , n63809 , n63810 , n63811 , n63812 , n63813 , n63814 , n63815 , n63816 , n63817 , n63818 , n63819 , n63820 , n63821 , n63822 , n63823 , n63824 , n63825 , n63826 , n63827 , n63828 , n63829 , n63830 , n63831 , n63832 , n63833 , n63834 , n63835 , n63836 , n63837 , n63838 , n63839 , n63840 , n63841 , n63842 , n63843 , n63844 , n63845 , n63846 , n63847 , n63848 , n63849 , n63850 , n63851 , n63852 , n63853 , n63854 , n63855 , n63856 , n63857 , n63858 , n63859 , n63860 , n63861 , n63862 , n63863 , n63864 , n63865 , n63866 , n63867 , n63868 , n63869 , n63870 , n63871 , n63872 , n63873 , n63874 , n63875 , n63876 , n63877 , n63878 , n63879 , n63880 , n63881 , n63882 , n63883 , n63884 , n63885 , n63886 , n63887 , n63888 , n63889 , n63890 , n63891 , n63892 , n63893 , n63894 , n63895 , n63896 , n63897 , n63898 , n63899 , n63900 , n63901 , n63902 , n63903 , n63904 , n63905 , n63906 , n63907 , n63908 , n63909 , n63910 , n63911 , n63912 , n63913 , n63914 , n63915 , n63916 , n63917 , n63918 , n63919 , n63920 , n63921 , n63922 , n63923 , n63924 , n63925 , n63926 , n63927 , n63928 , n63929 , n63930 , n63931 , n63932 , n63933 , n63934 , n63935 , n63936 , n63937 , n63938 , n63939 , n63940 , n63941 , n63942 , n63943 , n63944 , n63945 , n63946 , n63947 , n63948 , n63949 , n63950 , n63951 , n63952 , n63953 , n63954 , n63955 , n63956 , n63957 , n63958 , n63959 , n63960 , n63961 , n63962 , n63963 , n63964 , n63965 , n63966 , n63967 , n63968 , n63969 , n63970 , n63971 , n63972 , n63973 , n63974 , n63975 , n63976 , n63977 , n63978 , n63979 , n63980 , n63981 , n63982 , n63983 , n63984 , n63985 , n63986 , n63987 , n63988 , n63989 , n63990 , n63991 , n63992 , n63993 , n63994 , n63995 , n63996 , n63997 , n63998 , n63999 , n64000 , n64001 , n64002 , n64003 , n64004 , n64005 , n64006 , n64007 , n64008 , n64009 , n64010 , n64011 , n64012 , n64013 , n64014 , n64015 , n64016 , n64017 , n64018 , n64019 , n64020 , n64021 , n64022 , n64023 , n64024 , n64025 , n64026 , n64027 , n64028 , n64029 , n64030 , n64031 , n64032 , n64033 , n64034 , n64035 , n64036 , n64037 , n64038 , n64039 , n64040 , n64041 , n64042 , n64043 , n64044 , n64045 , n64046 , n64047 , n64048 , n64049 , n64050 , n64051 , n64052 , n64053 , n64054 , n64055 , n64056 , n64057 , n64058 , n64059 , n64060 , n64061 , n64062 , n64063 , n64064 , n64065 , n64066 , n64067 , n64068 , n64069 , n64070 , n64071 , n64072 , n64073 , n64074 , n64075 , n64076 , n64077 , n64078 , n64079 , n64080 , n64081 , n64082 , n64083 , n64084 , n64085 , n64086 , n64087 , n64088 , n64089 , n64090 , n64091 , n64092 , n64093 , n64094 , n64095 , n64096 , n64097 , n64098 , n64099 , n64100 , n64101 , n64102 , n64103 , n64104 , n64105 , n64106 , n64107 , n64108 , n64109 , n64110 , n64111 , n64112 , n64113 , n64114 , n64115 , n64116 , n64117 , n64118 , n64119 , n64120 , n64121 , n64122 , n64123 , n64124 , n64125 , n64126 , n64127 , n64128 , n64129 , n64130 , n64131 , n64132 , n64133 , n64134 , n64135 , n64136 , n64137 , n64138 , n64139 , n64140 , n64141 , n64142 , n64143 , n64144 , n64145 , n64146 , n64147 , n64148 , n64149 , n64150 , n64151 , n64152 , n64153 , n64154 , n64155 , n64156 , n64157 , n64158 , n64159 , n64160 , n64161 , n64162 , n64163 , n64164 , n64165 , n64166 , n64167 , n64168 , n64169 , n64170 , n64171 , n64172 , n64173 , n64174 , n64175 , n64176 , n64177 , n64178 , n64179 , n64180 , n64181 , n64182 , n64183 , n64184 , n64185 , n64186 , n64187 , n64188 , n64189 , n64190 , n64191 , n64192 , n64193 , n64194 , n64195 , n64196 , n64197 , n64198 , n64199 , n64200 , n64201 , n64202 , n64203 , n64204 , n64205 , n64206 , n64207 , n64208 , n64209 , n64210 , n64211 , n64212 , n64213 , n64214 , n64215 , n64216 , n64217 , n64218 , n64219 , n64220 , n64221 , n64222 , n64223 , n64224 , n64225 , n64226 , n64227 , n64228 , n64229 , n64230 , n64231 , n64232 , n64233 , n64234 , n64235 , n64236 , n64237 , n64238 , n64239 , n64240 , n64241 , n64242 , n64243 , n64244 , n64245 , n64246 , n64247 , n64248 , n64249 , n64250 , n64251 , n64252 , n64253 , n64254 , n64255 , n64256 , n64257 , n64258 , n64259 , n64260 , n64261 , n64262 , n64263 , n64264 , n64265 , n64266 , n64267 , n64268 , n64269 , n64270 , n64271 , n64272 , n64273 , n64274 , n64275 , n64276 , n64277 , n64278 , n64279 , n64280 , n64281 , n64282 , n64283 , n64284 , n64285 , n64286 , n64287 , n64288 , n64289 , n64290 , n64291 , n64292 , n64293 , n64294 , n64295 , n64296 , n64297 , n64298 , n64299 , n64300 , n64301 , n64302 , n64303 , n64304 , n64305 , n64306 , n64307 , n64308 , n64309 , n64310 , n64311 , n64312 , n64313 , n64314 , n64315 , n64316 , n64317 , n64318 , n64319 , n64320 , n64321 , n64322 , n64323 , n64324 , n64325 , n64326 , n64327 , n64328 , n64329 , n64330 , n64331 , n64332 , n64333 , n64334 , n64335 , n64336 , n64337 , n64338 , n64339 , n64340 , n64341 , n64342 , n64343 , n64344 , n64345 , n64346 , n64347 , n64348 , n64349 , n64350 , n64351 , n64352 , n64353 , n64354 , n64355 , n64356 , n64357 , n64358 , n64359 , n64360 , n64361 , n64362 , n64363 , n64364 , n64365 , n64366 , n64367 , n64368 , n64369 , n64370 , n64371 , n64372 , n64373 , n64374 , n64375 , n64376 , n64377 , n64378 , n64379 , n64380 , n64381 , n64382 , n64383 , n64384 , n64385 , n64386 , n64387 , n64388 , n64389 , n64390 , n64391 , n64392 , n64393 , n64394 , n64395 , n64396 , n64397 , n64398 , n64399 , n64400 , n64401 , n64402 , n64403 , n64404 , n64405 , n64406 , n64407 , n64408 , n64409 , n64410 , n64411 , n64412 , n64413 , n64414 , n64415 , n64416 , n64417 , n64418 , n64419 , n64420 , n64421 , n64422 , n64423 , n64424 , n64425 , n64426 , n64427 , n64428 , n64429 , n64430 , n64431 , n64432 , n64433 , n64434 , n64435 , n64436 , n64437 , n64438 , n64439 , n64440 , n64441 , n64442 , n64443 , n64444 , n64445 , n64446 , n64447 , n64448 , n64449 , n64450 , n64451 , n64452 , n64453 , n64454 , n64455 , n64456 , n64457 , n64458 , n64459 , n64460 , n64461 , n64462 , n64463 , n64464 , n64465 , n64466 , n64467 , n64468 , n64469 , n64470 , n64471 , n64472 , n64473 , n64474 , n64475 , n64476 , n64477 , n64478 , n64479 , n64480 , n64481 , n64482 , n64483 , n64484 , n64485 , n64486 , n64487 , n64488 , n64489 , n64490 , n64491 , n64492 , n64493 , n64494 , n64495 , n64496 , n64497 , n64498 , n64499 , n64500 , n64501 , n64502 , n64503 , n64504 , n64505 , n64506 , n64507 , n64508 , n64509 , n64510 , n64511 , n64512 , n64513 , n64514 , n64515 , n64516 , n64517 , n64518 , n64519 , n64520 , n64521 , n64522 , n64523 , n64524 , n64525 , n64526 , n64527 , n64528 , n64529 , n64530 , n64531 , n64532 , n64533 , n64534 , n64535 , n64536 , n64537 , n64538 , n64539 , n64540 , n64541 , n64542 , n64543 , n64544 , n64545 , n64546 , n64547 , n64548 , n64549 , n64550 , n64551 , n64552 , n64553 , n64554 , n64555 , n64556 , n64557 , n64558 , n64559 , n64560 , n64561 , n64562 , n64563 , n64564 , n64565 , n64566 , n64567 , n64568 , n64569 , n64570 , n64571 , n64572 , n64573 , n64574 , n64575 , n64576 , n64577 , n64578 , n64579 , n64580 , n64581 , n64582 , n64583 , n64584 , n64585 , n64586 , n64587 , n64588 , n64589 , n64590 , n64591 , n64592 , n64593 , n64594 , n64595 , n64596 , n64597 , n64598 , n64599 , n64600 , n64601 , n64602 , n64603 , n64604 , n64605 , n64606 , n64607 , n64608 , n64609 , n64610 , n64611 , n64612 , n64613 , n64614 , n64615 , n64616 , n64617 , n64618 , n64619 , n64620 , n64621 , n64622 , n64623 , n64624 , n64625 , n64626 , n64627 , n64628 , n64629 , n64630 , n64631 , n64632 , n64633 , n64634 , n64635 , n64636 , n64637 , n64638 , n64639 , n64640 , n64641 , n64642 , n64643 , n64644 , n64645 , n64646 , n64647 , n64648 , n64649 , n64650 , n64651 , n64652 , n64653 , n64654 , n64655 , n64656 , n64657 , n64658 , n64659 , n64660 , n64661 , n64662 , n64663 , n64664 , n64665 , n64666 , n64667 , n64668 , n64669 , n64670 , n64671 , n64672 , n64673 , n64674 , n64675 , n64676 , n64677 , n64678 , n64679 , n64680 , n64681 , n64682 , n64683 , n64684 , n64685 , n64686 , n64687 , n64688 , n64689 , n64690 , n64691 , n64692 , n64693 , n64694 , n64695 , n64696 , n64697 , n64698 , n64699 , n64700 , n64701 , n64702 , n64703 , n64704 , n64705 , n64706 , n64707 , n64708 , n64709 , n64710 , n64711 , n64712 , n64713 , n64714 , n64715 , n64716 , n64717 , n64718 , n64719 , n64720 , n64721 , n64722 , n64723 , n64724 , n64725 , n64726 , n64727 , n64728 , n64729 , n64730 , n64731 , n64732 , n64733 , n64734 , n64735 , n64736 , n64737 , n64738 , n64739 , n64740 , n64741 , n64742 , n64743 , n64744 , n64745 , n64746 , n64747 , n64748 , n64749 , n64750 , n64751 , n64752 , n64753 , n64754 , n64755 , n64756 , n64757 , n64758 , n64759 , n64760 , n64761 , n64762 , n64763 , n64764 , n64765 , n64766 , n64767 , n64768 , n64769 , n64770 , n64771 , n64772 , n64773 , n64774 , n64775 , n64776 , n64777 , n64778 , n64779 , n64780 , n64781 , n64782 , n64783 , n64784 , n64785 , n64786 , n64787 , n64788 , n64789 , n64790 , n64791 , n64792 , n64793 , n64794 , n64795 , n64796 , n64797 , n64798 , n64799 , n64800 , n64801 , n64802 , n64803 , n64804 , n64805 , n64806 , n64807 , n64808 , n64809 , n64810 , n64811 , n64812 , n64813 , n64814 , n64815 , n64816 , n64817 , n64818 , n64819 , n64820 , n64821 , n64822 , n64823 , n64824 , n64825 , n64826 , n64827 , n64828 , n64829 , n64830 , n64831 , n64832 , n64833 , n64834 , n64835 , n64836 , n64837 , n64838 , n64839 , n64840 , n64841 , n64842 , n64843 , n64844 , n64845 , n64846 , n64847 , n64848 , n64849 , n64850 , n64851 , n64852 , n64853 , n64854 , n64855 , n64856 , n64857 , n64858 , n64859 , n64860 , n64861 , n64862 , n64863 , n64864 , n64865 , n64866 , n64867 , n64868 , n64869 , n64870 , n64871 , n64872 , n64873 , n64874 , n64875 , n64876 , n64877 , n64878 , n64879 , n64880 , n64881 , n64882 , n64883 , n64884 , n64885 , n64886 , n64887 , n64888 , n64889 , n64890 , n64891 , n64892 , n64893 , n64894 , n64895 , n64896 , n64897 , n64898 , n64899 , n64900 , n64901 , n64902 , n64903 , n64904 , n64905 , n64906 , n64907 , n64908 , n64909 , n64910 , n64911 , n64912 , n64913 , n64914 , n64915 , n64916 , n64917 , n64918 , n64919 , n64920 , n64921 , n64922 , n64923 , n64924 , n64925 , n64926 , n64927 , n64928 , n64929 , n64930 , n64931 , n64932 , n64933 , n64934 , n64935 , n64936 , n64937 , n64938 , n64939 , n64940 , n64941 , n64942 , n64943 , n64944 , n64945 , n64946 , n64947 , n64948 , n64949 , n64950 , n64951 , n64952 , n64953 , n64954 , n64955 , n64956 , n64957 , n64958 , n64959 , n64960 , n64961 , n64962 , n64963 , n64964 , n64965 , n64966 , n64967 , n64968 , n64969 , n64970 , n64971 , n64972 , n64973 , n64974 , n64975 , n64976 , n64977 , n64978 , n64979 , n64980 , n64981 , n64982 , n64983 , n64984 , n64985 , n64986 , n64987 , n64988 , n64989 , n64990 , n64991 , n64992 , n64993 , n64994 , n64995 , n64996 , n64997 , n64998 , n64999 , n65000 , n65001 , n65002 , n65003 , n65004 , n65005 , n65006 , n65007 , n65008 , n65009 , n65010 , n65011 , n65012 , n65013 , n65014 , n65015 , n65016 , n65017 , n65018 , n65019 , n65020 , n65021 , n65022 , n65023 , n65024 , n65025 , n65026 , n65027 , n65028 , n65029 , n65030 , n65031 , n65032 , n65033 , n65034 , n65035 , n65036 , n65037 , n65038 , n65039 , n65040 , n65041 , n65042 , n65043 , n65044 , n65045 , n65046 , n65047 , n65048 , n65049 , n65050 , n65051 , n65052 , n65053 , n65054 , n65055 , n65056 , n65057 , n65058 , n65059 , n65060 , n65061 , n65062 , n65063 , n65064 , n65065 , n65066 , n65067 , n65068 , n65069 , n65070 , n65071 , n65072 , n65073 , n65074 , n65075 , n65076 , n65077 , n65078 , n65079 , n65080 , n65081 , n65082 , n65083 , n65084 , n65085 , n65086 , n65087 , n65088 , n65089 , n65090 , n65091 , n65092 , n65093 , n65094 , n65095 , n65096 , n65097 , n65098 , n65099 , n65100 , n65101 , n65102 , n65103 , n65104 , n65105 , n65106 , n65107 , n65108 , n65109 , n65110 , n65111 , n65112 , n65113 , n65114 , n65115 , n65116 , n65117 , n65118 , n65119 , n65120 , n65121 , n65122 , n65123 , n65124 , n65125 , n65126 , n65127 , n65128 , n65129 , n65130 , n65131 , n65132 , n65133 , n65134 , n65135 , n65136 , n65137 , n65138 , n65139 , n65140 , n65141 , n65142 , n65143 , n65144 , n65145 , n65146 , n65147 , n65148 , n65149 , n65150 , n65151 , n65152 , n65153 , n65154 , n65155 , n65156 , n65157 , n65158 , n65159 , n65160 , n65161 , n65162 , n65163 , n65164 , n65165 , n65166 , n65167 , n65168 , n65169 , n65170 , n65171 , n65172 , n65173 , n65174 , n65175 , n65176 , n65177 , n65178 , n65179 , n65180 , n65181 , n65182 , n65183 , n65184 , n65185 , n65186 , n65187 , n65188 , n65189 , n65190 , n65191 , n65192 , n65193 , n65194 , n65195 , n65196 , n65197 , n65198 , n65199 , n65200 , n65201 , n65202 , n65203 , n65204 , n65205 , n65206 , n65207 , n65208 , n65209 , n65210 , n65211 , n65212 , n65213 , n65214 , n65215 , n65216 , n65217 , n65218 , n65219 , n65220 , n65221 , n65222 , n65223 , n65224 , n65225 , n65226 , n65227 , n65228 , n65229 , n65230 , n65231 , n65232 , n65233 , n65234 , n65235 , n65236 , n65237 , n65238 , n65239 , n65240 , n65241 , n65242 , n65243 , n65244 , n65245 , n65246 , n65247 , n65248 , n65249 , n65250 , n65251 , n65252 , n65253 , n65254 , n65255 , n65256 , n65257 , n65258 , n65259 , n65260 , n65261 , n65262 , n65263 , n65264 , n65265 , n65266 , n65267 , n65268 , n65269 , n65270 , n65271 , n65272 , n65273 , n65274 , n65275 , n65276 , n65277 , n65278 , n65279 , n65280 , n65281 , n65282 , n65283 , n65284 , n65285 , n65286 , n65287 , n65288 , n65289 , n65290 , n65291 , n65292 , n65293 , n65294 , n65295 , n65296 , n65297 , n65298 , n65299 , n65300 , n65301 , n65302 , n65303 , n65304 , n65305 , n65306 , n65307 , n65308 , n65309 , n65310 , n65311 , n65312 , n65313 , n65314 , n65315 , n65316 , n65317 , n65318 , n65319 , n65320 , n65321 , n65322 , n65323 , n65324 , n65325 , n65326 , n65327 , n65328 , n65329 , n65330 , n65331 , n65332 , n65333 , n65334 , n65335 , n65336 , n65337 , n65338 , n65339 , n65340 , n65341 , n65342 , n65343 , n65344 , n65345 , n65346 , n65347 , n65348 , n65349 , n65350 , n65351 , n65352 , n65353 , n65354 , n65355 , n65356 , n65357 , n65358 , n65359 , n65360 , n65361 , n65362 , n65363 , n65364 , n65365 , n65366 , n65367 , n65368 , n65369 , n65370 , n65371 , n65372 , n65373 , n65374 , n65375 , n65376 , n65377 , n65378 , n65379 , n65380 , n65381 , n65382 , n65383 , n65384 , n65385 , n65386 , n65387 , n65388 , n65389 , n65390 , n65391 , n65392 , n65393 , n65394 , n65395 , n65396 , n65397 , n65398 , n65399 , n65400 , n65401 , n65402 , n65403 , n65404 , n65405 , n65406 , n65407 , n65408 , n65409 , n65410 , n65411 , n65412 , n65413 , n65414 , n65415 , n65416 , n65417 , n65418 , n65419 , n65420 , n65421 , n65422 , n65423 , n65424 , n65425 , n65426 , n65427 , n65428 , n65429 , n65430 , n65431 , n65432 , n65433 , n65434 , n65435 , n65436 , n65437 , n65438 , n65439 , n65440 , n65441 , n65442 , n65443 , n65444 , n65445 , n65446 , n65447 , n65448 , n65449 , n65450 , n65451 , n65452 , n65453 , n65454 , n65455 , n65456 , n65457 , n65458 , n65459 , n65460 , n65461 , n65462 , n65463 , n65464 , n65465 , n65466 , n65467 , n65468 , n65469 , n65470 , n65471 , n65472 , n65473 , n65474 , n65475 , n65476 , n65477 , n65478 , n65479 , n65480 , n65481 , n65482 , n65483 , n65484 , n65485 , n65486 , n65487 , n65488 , n65489 , n65490 , n65491 , n65492 , n65493 , n65494 , n65495 , n65496 , n65497 , n65498 , n65499 , n65500 , n65501 , n65502 , n65503 , n65504 , n65505 , n65506 , n65507 , n65508 , n65509 , n65510 , n65511 , n65512 , n65513 , n65514 , n65515 , n65516 , n65517 , n65518 , n65519 , n65520 , n65521 , n65522 , n65523 , n65524 , n65525 , n65526 , n65527 , n65528 , n65529 , n65530 , n65531 , n65532 , n65533 , n65534 , n65535 , n65536 , n65537 , n65538 , n65539 , n65540 , n65541 , n65542 , n65543 , n65544 , n65545 , n65546 , n65547 , n65548 , n65549 , n65550 , n65551 , n65552 , n65553 , n65554 , n65555 , n65556 , n65557 , n65558 , n65559 , n65560 , n65561 , n65562 , n65563 , n65564 , n65565 , n65566 , n65567 , n65568 , n65569 , n65570 , n65571 , n65572 , n65573 , n65574 , n65575 , n65576 , n65577 , n65578 , n65579 , n65580 , n65581 , n65582 , n65583 , n65584 , n65585 , n65586 , n65587 , n65588 , n65589 , n65590 , n65591 , n65592 , n65593 , n65594 , n65595 , n65596 , n65597 , n65598 , n65599 , n65600 , n65601 , n65602 , n65603 , n65604 , n65605 , n65606 , n65607 , n65608 , n65609 , n65610 , n65611 , n65612 , n65613 , n65614 , n65615 , n65616 , n65617 , n65618 , n65619 , n65620 , n65621 , n65622 , n65623 , n65624 , n65625 , n65626 , n65627 , n65628 , n65629 , n65630 , n65631 , n65632 , n65633 , n65634 , n65635 , n65636 , n65637 , n65638 , n65639 , n65640 , n65641 , n65642 , n65643 , n65644 , n65645 , n65646 , n65647 , n65648 , n65649 , n65650 , n65651 , n65652 , n65653 , n65654 , n65655 , n65656 , n65657 , n65658 , n65659 , n65660 , n65661 , n65662 , n65663 , n65664 , n65665 , n65666 , n65667 , n65668 , n65669 , n65670 , n65671 , n65672 , n65673 , n65674 , n65675 , n65676 , n65677 , n65678 , n65679 , n65680 , n65681 , n65682 , n65683 , n65684 , n65685 , n65686 , n65687 , n65688 , n65689 , n65690 , n65691 , n65692 , n65693 , n65694 , n65695 , n65696 , n65697 , n65698 , n65699 , n65700 , n65701 , n65702 , n65703 , n65704 , n65705 , n65706 , n65707 , n65708 , n65709 , n65710 , n65711 , n65712 , n65713 , n65714 , n65715 , n65716 , n65717 , n65718 , n65719 , n65720 , n65721 , n65722 , n65723 , n65724 , n65725 , n65726 , n65727 , n65728 , n65729 , n65730 , n65731 , n65732 , n65733 , n65734 , n65735 , n65736 , n65737 , n65738 , n65739 , n65740 , n65741 , n65742 , n65743 , n65744 , n65745 , n65746 , n65747 , n65748 , n65749 , n65750 , n65751 , n65752 , n65753 , n65754 , n65755 , n65756 , n65757 , n65758 , n65759 , n65760 , n65761 , n65762 , n65763 , n65764 , n65765 , n65766 , n65767 , n65768 , n65769 , n65770 , n65771 , n65772 , n65773 , n65774 , n65775 , n65776 , n65777 , n65778 , n65779 , n65780 , n65781 , n65782 , n65783 , n65784 , n65785 , n65786 , n65787 , n65788 , n65789 , n65790 , n65791 , n65792 , n65793 , n65794 , n65795 , n65796 , n65797 , n65798 , n65799 , n65800 , n65801 , n65802 , n65803 , n65804 , n65805 , n65806 , n65807 , n65808 , n65809 , n65810 , n65811 , n65812 , n65813 , n65814 , n65815 , n65816 , n65817 , n65818 , n65819 , n65820 , n65821 , n65822 , n65823 , n65824 , n65825 , n65826 , n65827 , n65828 , n65829 , n65830 , n65831 , n65832 , n65833 , n65834 , n65835 , n65836 , n65837 , n65838 , n65839 , n65840 , n65841 , n65842 , n65843 , n65844 , n65845 , n65846 , n65847 , n65848 , n65849 , n65850 , n65851 , n65852 , n65853 , n65854 , n65855 , n65856 , n65857 , n65858 , n65859 , n65860 , n65861 , n65862 , n65863 , n65864 , n65865 , n65866 , n65867 , n65868 , n65869 , n65870 , n65871 , n65872 , n65873 , n65874 , n65875 , n65876 , n65877 , n65878 , n65879 , n65880 , n65881 , n65882 , n65883 , n65884 , n65885 , n65886 , n65887 , n65888 , n65889 , n65890 , n65891 , n65892 , n65893 , n65894 , n65895 , n65896 , n65897 , n65898 , n65899 , n65900 , n65901 , n65902 , n65903 , n65904 , n65905 , n65906 , n65907 , n65908 , n65909 , n65910 , n65911 , n65912 , n65913 , n65914 , n65915 , n65916 , n65917 , n65918 , n65919 , n65920 , n65921 , n65922 , n65923 , n65924 , n65925 , n65926 , n65927 , n65928 , n65929 , n65930 , n65931 , n65932 , n65933 , n65934 , n65935 , n65936 , n65937 , n65938 , n65939 , n65940 , n65941 , n65942 , n65943 , n65944 , n65945 , n65946 , n65947 , n65948 , n65949 , n65950 , n65951 , n65952 , n65953 , n65954 , n65955 , n65956 , n65957 , n65958 , n65959 , n65960 , n65961 , n65962 , n65963 , n65964 , n65965 , n65966 , n65967 , n65968 , n65969 , n65970 , n65971 , n65972 , n65973 , n65974 , n65975 , n65976 , n65977 , n65978 , n65979 , n65980 , n65981 , n65982 , n65983 , n65984 , n65985 , n65986 , n65987 , n65988 , n65989 , n65990 , n65991 , n65992 , n65993 , n65994 , n65995 , n65996 , n65997 , n65998 , n65999 , n66000 , n66001 , n66002 , n66003 , n66004 , n66005 , n66006 , n66007 , n66008 , n66009 , n66010 , n66011 , n66012 , n66013 , n66014 , n66015 , n66016 , n66017 , n66018 , n66019 , n66020 , n66021 , n66022 , n66023 , n66024 , n66025 , n66026 , n66027 , n66028 , n66029 , n66030 , n66031 , n66032 , n66033 , n66034 , n66035 , n66036 , n66037 , n66038 , n66039 , n66040 , n66041 , n66042 , n66043 , n66044 , n66045 , n66046 , n66047 , n66048 , n66049 , n66050 , n66051 , n66052 , n66053 , n66054 , n66055 , n66056 , n66057 , n66058 , n66059 , n66060 , n66061 , n66062 , n66063 , n66064 , n66065 , n66066 , n66067 , n66068 , n66069 , n66070 , n66071 , n66072 , n66073 , n66074 , n66075 , n66076 , n66077 , n66078 , n66079 , n66080 , n66081 , n66082 , n66083 , n66084 , n66085 , n66086 , n66087 , n66088 , n66089 , n66090 , n66091 , n66092 , n66093 , n66094 , n66095 , n66096 , n66097 , n66098 , n66099 , n66100 , n66101 , n66102 , n66103 , n66104 , n66105 , n66106 , n66107 , n66108 , n66109 , n66110 , n66111 , n66112 , n66113 , n66114 , n66115 , n66116 , n66117 , n66118 , n66119 , n66120 , n66121 , n66122 , n66123 , n66124 , n66125 , n66126 , n66127 , n66128 , n66129 , n66130 , n66131 , n66132 , n66133 , n66134 , n66135 , n66136 , n66137 , n66138 , n66139 , n66140 , n66141 , n66142 , n66143 , n66144 , n66145 , n66146 , n66147 , n66148 , n66149 , n66150 , n66151 , n66152 , n66153 , n66154 , n66155 , n66156 , n66157 , n66158 , n66159 , n66160 , n66161 , n66162 , n66163 , n66164 , n66165 , n66166 , n66167 , n66168 , n66169 , n66170 , n66171 , n66172 , n66173 , n66174 , n66175 , n66176 , n66177 , n66178 , n66179 , n66180 , n66181 , n66182 , n66183 , n66184 , n66185 , n66186 , n66187 , n66188 , n66189 , n66190 , n66191 , n66192 , n66193 , n66194 , n66195 , n66196 , n66197 , n66198 , n66199 , n66200 , n66201 , n66202 , n66203 , n66204 , n66205 , n66206 , n66207 , n66208 , n66209 , n66210 , n66211 , n66212 , n66213 , n66214 , n66215 , n66216 , n66217 , n66218 , n66219 , n66220 , n66221 , n66222 , n66223 , n66224 , n66225 , n66226 , n66227 , n66228 , n66229 , n66230 , n66231 , n66232 , n66233 , n66234 , n66235 , n66236 , n66237 , n66238 , n66239 , n66240 , n66241 , n66242 , n66243 , n66244 , n66245 , n66246 , n66247 , n66248 , n66249 , n66250 , n66251 , n66252 , n66253 , n66254 , n66255 , n66256 , n66257 , n66258 , n66259 , n66260 , n66261 , n66262 , n66263 , n66264 , n66265 , n66266 , n66267 , n66268 , n66269 , n66270 , n66271 , n66272 , n66273 , n66274 , n66275 , n66276 , n66277 , n66278 , n66279 , n66280 , n66281 , n66282 , n66283 , n66284 , n66285 , n66286 , n66287 , n66288 , n66289 , n66290 , n66291 , n66292 , n66293 , n66294 , n66295 , n66296 , n66297 , n66298 , n66299 , n66300 , n66301 , n66302 , n66303 , n66304 , n66305 , n66306 , n66307 , n66308 , n66309 , n66310 , n66311 , n66312 , n66313 , n66314 , n66315 , n66316 , n66317 , n66318 , n66319 , n66320 , n66321 , n66322 , n66323 , n66324 , n66325 , n66326 , n66327 , n66328 , n66329 , n66330 , n66331 , n66332 , n66333 , n66334 , n66335 , n66336 , n66337 , n66338 , n66339 , n66340 , n66341 , n66342 , n66343 , n66344 , n66345 , n66346 , n66347 , n66348 , n66349 , n66350 , n66351 , n66352 , n66353 , n66354 , n66355 , n66356 , n66357 , n66358 , n66359 , n66360 , n66361 , n66362 , n66363 , n66364 , n66365 , n66366 , n66367 , n66368 , n66369 , n66370 , n66371 , n66372 , n66373 , n66374 , n66375 , n66376 , n66377 , n66378 , n66379 , n66380 , n66381 , n66382 , n66383 , n66384 , n66385 , n66386 , n66387 , n66388 , n66389 , n66390 , n66391 , n66392 , n66393 , n66394 , n66395 , n66396 , n66397 , n66398 , n66399 , n66400 , n66401 , n66402 , n66403 , n66404 , n66405 , n66406 , n66407 , n66408 , n66409 , n66410 , n66411 , n66412 , n66413 , n66414 , n66415 , n66416 , n66417 , n66418 , n66419 , n66420 , n66421 , n66422 , n66423 , n66424 , n66425 , n66426 , n66427 , n66428 , n66429 , n66430 , n66431 , n66432 , n66433 , n66434 , n66435 , n66436 , n66437 , n66438 , n66439 , n66440 , n66441 , n66442 , n66443 , n66444 , n66445 , n66446 , n66447 , n66448 , n66449 , n66450 , n66451 , n66452 , n66453 , n66454 , n66455 , n66456 , n66457 , n66458 , n66459 , n66460 , n66461 , n66462 , n66463 , n66464 , n66465 , n66466 , n66467 , n66468 , n66469 , n66470 , n66471 , n66472 , n66473 , n66474 , n66475 , n66476 , n66477 , n66478 , n66479 , n66480 , n66481 , n66482 , n66483 , n66484 , n66485 , n66486 , n66487 , n66488 , n66489 , n66490 , n66491 , n66492 , n66493 , n66494 , n66495 , n66496 , n66497 , n66498 , n66499 , n66500 , n66501 , n66502 , n66503 , n66504 , n66505 , n66506 , n66507 , n66508 , n66509 , n66510 , n66511 , n66512 , n66513 , n66514 , n66515 , n66516 , n66517 , n66518 , n66519 , n66520 , n66521 , n66522 , n66523 , n66524 , n66525 , n66526 , n66527 , n66528 , n66529 , n66530 , n66531 , n66532 , n66533 , n66534 , n66535 , n66536 , n66537 , n66538 , n66539 , n66540 , n66541 , n66542 , n66543 , n66544 , n66545 , n66546 , n66547 , n66548 , n66549 , n66550 , n66551 , n66552 , n66553 , n66554 , n66555 , n66556 , n66557 , n66558 , n66559 , n66560 , n66561 , n66562 , n66563 , n66564 , n66565 , n66566 , n66567 , n66568 , n66569 , n66570 , n66571 , n66572 , n66573 , n66574 , n66575 , n66576 , n66577 , n66578 , n66579 , n66580 , n66581 , n66582 , n66583 , n66584 , n66585 , n66586 , n66587 , n66588 , n66589 , n66590 , n66591 , n66592 , n66593 , n66594 , n66595 , n66596 , n66597 , n66598 , n66599 , n66600 , n66601 , n66602 , n66603 , n66604 , n66605 , n66606 , n66607 , n66608 , n66609 , n66610 , n66611 , n66612 , n66613 , n66614 , n66615 , n66616 , n66617 , n66618 , n66619 , n66620 , n66621 , n66622 , n66623 , n66624 , n66625 , n66626 , n66627 , n66628 , n66629 , n66630 , n66631 , n66632 , n66633 , n66634 , n66635 , n66636 , n66637 , n66638 , n66639 , n66640 , n66641 , n66642 , n66643 , n66644 , n66645 , n66646 , n66647 , n66648 , n66649 , n66650 , n66651 , n66652 , n66653 , n66654 , n66655 , n66656 , n66657 , n66658 , n66659 , n66660 , n66661 , n66662 , n66663 , n66664 , n66665 , n66666 , n66667 , n66668 , n66669 , n66670 , n66671 , n66672 , n66673 , n66674 , n66675 , n66676 , n66677 , n66678 , n66679 , n66680 , n66681 , n66682 , n66683 , n66684 , n66685 , n66686 , n66687 , n66688 , n66689 , n66690 , n66691 , n66692 , n66693 , n66694 , n66695 , n66696 , n66697 , n66698 , n66699 , n66700 , n66701 , n66702 , n66703 , n66704 , n66705 , n66706 , n66707 , n66708 , n66709 , n66710 , n66711 , n66712 , n66713 , n66714 , n66715 , n66716 , n66717 , n66718 , n66719 , n66720 , n66721 , n66722 , n66723 , n66724 , n66725 , n66726 , n66727 , n66728 , n66729 , n66730 , n66731 , n66732 , n66733 , n66734 , n66735 , n66736 , n66737 , n66738 , n66739 , n66740 , n66741 , n66742 , n66743 , n66744 , n66745 , n66746 , n66747 , n66748 , n66749 , n66750 , n66751 , n66752 , n66753 , n66754 , n66755 , n66756 , n66757 , n66758 , n66759 , n66760 , n66761 , n66762 , n66763 , n66764 , n66765 , n66766 , n66767 , n66768 , n66769 , n66770 , n66771 , n66772 , n66773 , n66774 , n66775 , n66776 , n66777 , n66778 , n66779 , n66780 , n66781 , n66782 , n66783 , n66784 , n66785 , n66786 , n66787 , n66788 , n66789 , n66790 , n66791 , n66792 , n66793 , n66794 , n66795 , n66796 , n66797 , n66798 , n66799 , n66800 , n66801 , n66802 , n66803 , n66804 , n66805 , n66806 , n66807 , n66808 , n66809 , n66810 , n66811 , n66812 , n66813 , n66814 , n66815 , n66816 , n66817 , n66818 , n66819 , n66820 , n66821 , n66822 , n66823 , n66824 , n66825 , n66826 , n66827 , n66828 , n66829 , n66830 , n66831 , n66832 , n66833 , n66834 , n66835 , n66836 , n66837 , n66838 , n66839 , n66840 , n66841 , n66842 , n66843 , n66844 , n66845 , n66846 , n66847 , n66848 , n66849 , n66850 , n66851 , n66852 , n66853 , n66854 , n66855 , n66856 , n66857 , n66858 , n66859 , n66860 , n66861 , n66862 , n66863 , n66864 , n66865 , n66866 , n66867 , n66868 , n66869 , n66870 , n66871 , n66872 , n66873 , n66874 , n66875 , n66876 , n66877 , n66878 , n66879 , n66880 , n66881 , n66882 , n66883 , n66884 , n66885 , n66886 , n66887 , n66888 , n66889 , n66890 , n66891 , n66892 , n66893 , n66894 , n66895 , n66896 , n66897 , n66898 , n66899 , n66900 , n66901 , n66902 , n66903 , n66904 , n66905 , n66906 , n66907 , n66908 , n66909 , n66910 , n66911 , n66912 , n66913 , n66914 , n66915 , n66916 , n66917 , n66918 , n66919 , n66920 , n66921 , n66922 , n66923 , n66924 , n66925 , n66926 , n66927 , n66928 , n66929 , n66930 , n66931 , n66932 , n66933 , n66934 , n66935 , n66936 , n66937 , n66938 , n66939 , n66940 , n66941 , n66942 , n66943 , n66944 , n66945 , n66946 , n66947 , n66948 , n66949 , n66950 , n66951 , n66952 , n66953 , n66954 , n66955 , n66956 , n66957 , n66958 , n66959 , n66960 , n66961 , n66962 , n66963 , n66964 , n66965 , n66966 , n66967 , n66968 , n66969 , n66970 , n66971 , n66972 , n66973 , n66974 , n66975 , n66976 , n66977 , n66978 , n66979 , n66980 , n66981 , n66982 , n66983 , n66984 , n66985 , n66986 , n66987 , n66988 , n66989 , n66990 , n66991 , n66992 , n66993 , n66994 , n66995 , n66996 , n66997 , n66998 , n66999 , n67000 , n67001 , n67002 , n67003 , n67004 , n67005 , n67006 , n67007 , n67008 , n67009 , n67010 , n67011 , n67012 , n67013 , n67014 , n67015 , n67016 , n67017 , n67018 , n67019 , n67020 , n67021 , n67022 , n67023 , n67024 , n67025 , n67026 , n67027 , n67028 , n67029 , n67030 , n67031 , n67032 , n67033 , n67034 , n67035 , n67036 , n67037 , n67038 , n67039 , n67040 , n67041 , n67042 , n67043 , n67044 , n67045 , n67046 , n67047 , n67048 , n67049 , n67050 , n67051 , n67052 , n67053 , n67054 , n67055 , n67056 , n67057 , n67058 , n67059 , n67060 , n67061 , n67062 , n67063 , n67064 , n67065 , n67066 , n67067 , n67068 , n67069 , n67070 , n67071 , n67072 , n67073 , n67074 , n67075 , n67076 , n67077 , n67078 , n67079 , n67080 , n67081 , n67082 , n67083 , n67084 , n67085 , n67086 , n67087 , n67088 , n67089 , n67090 , n67091 , n67092 , n67093 , n67094 , n67095 , n67096 , n67097 , n67098 , n67099 , n67100 , n67101 , n67102 , n67103 , n67104 , n67105 , n67106 , n67107 , n67108 , n67109 , n67110 , n67111 , n67112 , n67113 , n67114 , n67115 , n67116 , n67117 , n67118 , n67119 , n67120 , n67121 , n67122 , n67123 , n67124 , n67125 , n67126 , n67127 , n67128 , n67129 , n67130 , n67131 , n67132 , n67133 , n67134 , n67135 , n67136 , n67137 , n67138 , n67139 , n67140 , n67141 , n67142 , n67143 , n67144 , n67145 , n67146 , n67147 , n67148 , n67149 , n67150 , n67151 , n67152 , n67153 , n67154 , n67155 , n67156 , n67157 , n67158 , n67159 , n67160 , n67161 , n67162 , n67163 , n67164 , n67165 , n67166 , n67167 , n67168 , n67169 , n67170 , n67171 , n67172 , n67173 , n67174 , n67175 , n67176 , n67177 , n67178 , n67179 , n67180 , n67181 , n67182 , n67183 , n67184 , n67185 , n67186 , n67187 , n67188 , n67189 , n67190 , n67191 , n67192 , n67193 , n67194 , n67195 , n67196 , n67197 , n67198 , n67199 , n67200 , n67201 , n67202 , n67203 , n67204 , n67205 , n67206 , n67207 , n67208 , n67209 , n67210 , n67211 , n67212 , n67213 , n67214 , n67215 , n67216 , n67217 , n67218 , n67219 , n67220 , n67221 , n67222 , n67223 , n67224 , n67225 , n67226 , n67227 , n67228 , n67229 , n67230 , n67231 , n67232 , n67233 , n67234 , n67235 , n67236 , n67237 , n67238 , n67239 , n67240 , n67241 , n67242 , n67243 , n67244 , n67245 , n67246 , n67247 , n67248 , n67249 , n67250 , n67251 , n67252 , n67253 , n67254 , n67255 , n67256 , n67257 , n67258 , n67259 , n67260 , n67261 , n67262 , n67263 , n67264 , n67265 , n67266 , n67267 , n67268 , n67269 , n67270 , n67271 , n67272 , n67273 , n67274 , n67275 , n67276 , n67277 , n67278 , n67279 , n67280 , n67281 , n67282 , n67283 , n67284 , n67285 , n67286 , n67287 , n67288 , n67289 , n67290 , n67291 , n67292 , n67293 , n67294 , n67295 , n67296 , n67297 , n67298 , n67299 , n67300 , n67301 , n67302 , n67303 , n67304 , n67305 , n67306 , n67307 , n67308 , n67309 , n67310 , n67311 , n67312 , n67313 , n67314 , n67315 , n67316 , n67317 , n67318 , n67319 , n67320 , n67321 , n67322 , n67323 , n67324 , n67325 , n67326 , n67327 , n67328 , n67329 , n67330 , n67331 , n67332 , n67333 , n67334 , n67335 , n67336 , n67337 , n67338 , n67339 , n67340 , n67341 , n67342 , n67343 , n67344 , n67345 , n67346 , n67347 , n67348 , n67349 , n67350 , n67351 , n67352 , n67353 , n67354 , n67355 , n67356 , n67357 , n67358 , n67359 , n67360 , n67361 , n67362 , n67363 , n67364 , n67365 , n67366 , n67367 , n67368 , n67369 , n67370 , n67371 , n67372 , n67373 , n67374 , n67375 , n67376 , n67377 , n67378 , n67379 , n67380 , n67381 , n67382 , n67383 , n67384 , n67385 , n67386 , n67387 , n67388 , n67389 , n67390 , n67391 , n67392 , n67393 , n67394 , n67395 , n67396 , n67397 , n67398 , n67399 , n67400 , n67401 , n67402 , n67403 , n67404 , n67405 , n67406 , n67407 , n67408 , n67409 , n67410 , n67411 , n67412 , n67413 , n67414 , n67415 , n67416 , n67417 , n67418 , n67419 , n67420 , n67421 , n67422 , n67423 , n67424 , n67425 , n67426 , n67427 , n67428 , n67429 , n67430 , n67431 , n67432 , n67433 , n67434 , n67435 , n67436 , n67437 , n67438 , n67439 , n67440 , n67441 , n67442 , n67443 , n67444 , n67445 , n67446 , n67447 , n67448 , n67449 , n67450 , n67451 , n67452 , n67453 , n67454 , n67455 , n67456 , n67457 , n67458 , n67459 , n67460 , n67461 , n67462 , n67463 , n67464 , n67465 , n67466 , n67467 , n67468 , n67469 , n67470 , n67471 , n67472 , n67473 , n67474 , n67475 , n67476 , n67477 , n67478 , n67479 , n67480 , n67481 , n67482 , n67483 , n67484 , n67485 , n67486 , n67487 , n67488 , n67489 , n67490 , n67491 , n67492 , n67493 , n67494 , n67495 , n67496 , n67497 , n67498 , n67499 , n67500 , n67501 , n67502 , n67503 , n67504 , n67505 , n67506 , n67507 , n67508 , n67509 , n67510 , n67511 , n67512 , n67513 , n67514 , n67515 , n67516 , n67517 , n67518 , n67519 , n67520 , n67521 , n67522 , n67523 , n67524 , n67525 , n67526 , n67527 , n67528 , n67529 , n67530 , n67531 , n67532 , n67533 , n67534 , n67535 , n67536 , n67537 , n67538 , n67539 , n67540 , n67541 , n67542 , n67543 , n67544 , n67545 , n67546 , n67547 , n67548 , n67549 , n67550 , n67551 , n67552 , n67553 , n67554 , n67555 , n67556 , n67557 , n67558 , n67559 , n67560 , n67561 , n67562 , n67563 , n67564 , n67565 , n67566 , n67567 , n67568 , n67569 , n67570 , n67571 , n67572 , n67573 , n67574 , n67575 , n67576 , n67577 , n67578 , n67579 , n67580 , n67581 , n67582 , n67583 , n67584 , n67585 , n67586 , n67587 , n67588 , n67589 , n67590 , n67591 , n67592 , n67593 , n67594 , n67595 , n67596 , n67597 , n67598 , n67599 , n67600 , n67601 , n67602 , n67603 , n67604 , n67605 , n67606 , n67607 , n67608 , n67609 , n67610 , n67611 , n67612 , n67613 , n67614 , n67615 , n67616 , n67617 , n67618 , n67619 , n67620 , n67621 , n67622 , n67623 , n67624 , n67625 , n67626 , n67627 , n67628 , n67629 , n67630 , n67631 , n67632 , n67633 , n67634 , n67635 , n67636 , n67637 , n67638 , n67639 , n67640 , n67641 , n67642 , n67643 , n67644 , n67645 , n67646 , n67647 , n67648 , n67649 , n67650 , n67651 , n67652 , n67653 , n67654 , n67655 , n67656 , n67657 , n67658 , n67659 , n67660 , n67661 , n67662 , n67663 , n67664 , n67665 , n67666 , n67667 , n67668 , n67669 , n67670 , n67671 , n67672 , n67673 , n67674 , n67675 , n67676 , n67677 , n67678 , n67679 , n67680 , n67681 , n67682 , n67683 , n67684 , n67685 , n67686 , n67687 , n67688 , n67689 , n67690 , n67691 , n67692 , n67693 , n67694 , n67695 , n67696 , n67697 , n67698 , n67699 , n67700 , n67701 , n67702 , n67703 , n67704 , n67705 , n67706 , n67707 , n67708 , n67709 , n67710 , n67711 , n67712 , n67713 , n67714 , n67715 , n67716 , n67717 , n67718 , n67719 , n67720 , n67721 , n67722 , n67723 , n67724 , n67725 , n67726 , n67727 , n67728 , n67729 , n67730 , n67731 , n67732 , n67733 , n67734 , n67735 , n67736 , n67737 , n67738 , n67739 , n67740 , n67741 , n67742 , n67743 , n67744 , n67745 , n67746 , n67747 , n67748 , n67749 , n67750 , n67751 , n67752 , n67753 , n67754 , n67755 , n67756 , n67757 , n67758 , n67759 , n67760 , n67761 , n67762 , n67763 , n67764 , n67765 , n67766 , n67767 , n67768 , n67769 , n67770 , n67771 , n67772 , n67773 , n67774 , n67775 , n67776 , n67777 , n67778 , n67779 , n67780 , n67781 , n67782 , n67783 , n67784 , n67785 , n67786 , n67787 , n67788 , n67789 , n67790 , n67791 , n67792 , n67793 , n67794 , n67795 , n67796 , n67797 , n67798 , n67799 , n67800 , n67801 , n67802 , n67803 , n67804 , n67805 , n67806 , n67807 , n67808 , n67809 ;
  assign n2790 = ~\P1_P1_Datao_reg[30]/NET0131  & ~\P1_P2_Datao_reg[30]/NET0131  ;
  assign n2791 = ~\P1_P3_Datao_reg[30]/NET0131  & n2790 ;
  assign n2792 = \P1_P2_Address_reg[0]/NET0131  & ~n2791 ;
  assign n2793 = \P1_P3_Address_reg[0]/NET0131  & n2791 ;
  assign n2794 = ~n2792 & ~n2793 ;
  assign n2805 = ~\P4_datao_reg[26]/NET0131  & ~\P4_datao_reg[27]/NET0131  ;
  assign n2806 = ~\P4_datao_reg[28]/NET0131  & ~\P4_datao_reg[2]/NET0131  ;
  assign n2813 = n2805 & n2806 ;
  assign n2803 = ~\P4_datao_reg[22]/NET0131  & ~\P4_datao_reg[23]/NET0131  ;
  assign n2804 = ~\P4_datao_reg[24]/NET0131  & ~\P4_datao_reg[25]/NET0131  ;
  assign n2814 = n2803 & n2804 ;
  assign n2820 = n2813 & n2814 ;
  assign n2809 = ~\P4_datao_reg[6]/NET0131  & ~\P4_datao_reg[7]/NET0131  ;
  assign n2810 = ~\P4_datao_reg[8]/NET0131  & ~\P4_datao_reg[9]/NET0131  ;
  assign n2811 = n2809 & n2810 ;
  assign n2807 = ~\P4_datao_reg[30]/NET0131  & ~\P4_datao_reg[3]/NET0131  ;
  assign n2808 = ~\P4_datao_reg[4]/NET0131  & ~\P4_datao_reg[5]/NET0131  ;
  assign n2812 = n2807 & n2808 ;
  assign n2821 = n2811 & n2812 ;
  assign n2822 = n2820 & n2821 ;
  assign n2796 = ~\P4_datao_reg[0]/NET0131  & ~\P4_datao_reg[10]/NET0131  ;
  assign n2797 = ~\P4_datao_reg[11]/NET0131  & ~\P4_datao_reg[12]/NET0131  ;
  assign n2798 = ~\P4_datao_reg[13]/NET0131  & ~\P4_datao_reg[14]/NET0131  ;
  assign n2817 = n2797 & n2798 ;
  assign n2818 = n2796 & n2817 ;
  assign n2801 = ~\P4_datao_reg[19]/NET0131  & ~\P4_datao_reg[1]/NET0131  ;
  assign n2802 = ~\P4_datao_reg[20]/NET0131  & ~\P4_datao_reg[21]/NET0131  ;
  assign n2815 = n2801 & n2802 ;
  assign n2799 = ~\P4_datao_reg[15]/NET0131  & ~\P4_datao_reg[16]/NET0131  ;
  assign n2800 = ~\P4_datao_reg[17]/NET0131  & ~\P4_datao_reg[18]/NET0131  ;
  assign n2816 = n2799 & n2800 ;
  assign n2819 = n2815 & n2816 ;
  assign n2823 = n2818 & n2819 ;
  assign n2824 = n2822 & n2823 ;
  assign n2795 = ~\P4_datao_reg[29]/NET0131  & ~\P4_datao_reg[30]/NET0131  ;
  assign n2825 = ~\P4_datao_reg[31]/NET0131  & ~n2795 ;
  assign n2826 = ~n2824 & n2825 ;
  assign n2827 = ~\P2_P1_Datao_reg[30]/NET0131  & ~\P2_P2_Datao_reg[30]/NET0131  ;
  assign n2828 = ~\P2_P3_Datao_reg[30]/NET0131  & n2827 ;
  assign n2829 = \P2_P2_Address_reg[0]/NET0131  & ~n2828 ;
  assign n2830 = \P2_P3_Address_reg[0]/NET0131  & n2828 ;
  assign n2831 = ~n2829 & ~n2830 ;
  assign n2832 = ~n2826 & ~n2831 ;
  assign n2833 = \P2_P1_Address_reg[0]/NET0131  & n2826 ;
  assign n2834 = ~n2832 & ~n2833 ;
  assign n2835 = ~n2794 & ~n2834 ;
  assign n2836 = \P1_P2_Address_reg[1]/NET0131  & ~n2791 ;
  assign n2837 = \P1_P3_Address_reg[1]/NET0131  & n2791 ;
  assign n2838 = ~n2836 & ~n2837 ;
  assign n2839 = ~n2834 & ~n2838 ;
  assign n2840 = ~\P2_P3_Address_reg[1]/NET0131  & n2828 ;
  assign n2841 = ~\P2_P2_Address_reg[1]/NET0131  & ~n2828 ;
  assign n2842 = ~n2840 & ~n2841 ;
  assign n2843 = ~n2826 & ~n2842 ;
  assign n2844 = ~\P2_P1_Address_reg[1]/NET0131  & n2826 ;
  assign n2845 = ~n2843 & ~n2844 ;
  assign n2846 = ~n2794 & n2845 ;
  assign n2847 = n2839 & ~n2846 ;
  assign n2848 = ~n2839 & n2846 ;
  assign n2849 = ~n2847 & ~n2848 ;
  assign n2850 = \P1_P2_Address_reg[2]/NET0131  & ~n2791 ;
  assign n2851 = \P1_P3_Address_reg[2]/NET0131  & n2791 ;
  assign n2852 = ~n2850 & ~n2851 ;
  assign n2853 = ~n2834 & ~n2852 ;
  assign n2854 = ~n2838 & n2845 ;
  assign n2855 = n2834 & n2854 ;
  assign n2856 = ~n2853 & ~n2855 ;
  assign n2857 = ~n2834 & n2854 ;
  assign n2858 = n2794 & ~n2857 ;
  assign n2859 = ~\P2_P3_Address_reg[2]/NET0131  & n2828 ;
  assign n2860 = ~\P2_P2_Address_reg[2]/NET0131  & ~n2828 ;
  assign n2861 = ~n2859 & ~n2860 ;
  assign n2862 = ~n2826 & ~n2861 ;
  assign n2863 = ~\P2_P1_Address_reg[2]/NET0131  & n2826 ;
  assign n2864 = ~n2862 & ~n2863 ;
  assign n2865 = ~n2794 & ~n2864 ;
  assign n2866 = ~n2858 & ~n2865 ;
  assign n2867 = n2856 & ~n2866 ;
  assign n2868 = ~n2856 & n2866 ;
  assign n2869 = ~n2867 & ~n2868 ;
  assign n2870 = ~\P4_wr_reg/NET0131  & ~n2794 ;
  assign n2871 = \P4_addr_reg[0]/NET0131  & \P4_wr_reg/NET0131  ;
  assign n2872 = ~n2870 & ~n2871 ;
  assign n2873 = ~n2834 & ~n2872 ;
  assign n2874 = \P1_P2_Address_reg[7]/NET0131  & ~n2791 ;
  assign n2875 = \P1_P3_Address_reg[7]/NET0131  & n2791 ;
  assign n2876 = ~n2874 & ~n2875 ;
  assign n2877 = ~\P4_wr_reg/NET0131  & ~n2876 ;
  assign n2878 = \P4_addr_reg[7]/NET0131  & \P4_wr_reg/NET0131  ;
  assign n2879 = ~n2877 & ~n2878 ;
  assign n2880 = ~\P1_P2_Address_reg[8]/NET0131  & ~n2791 ;
  assign n2881 = ~\P1_P3_Address_reg[8]/NET0131  & n2791 ;
  assign n2882 = ~n2880 & ~n2881 ;
  assign n2883 = ~\P4_wr_reg/NET0131  & ~n2882 ;
  assign n2884 = ~\P4_addr_reg[8]/NET0131  & \P4_wr_reg/NET0131  ;
  assign n2885 = ~n2883 & ~n2884 ;
  assign n2886 = n2879 & ~n2885 ;
  assign n2887 = ~n2879 & n2885 ;
  assign n2888 = ~n2886 & ~n2887 ;
  assign n2889 = ~n2834 & n2888 ;
  assign n2890 = \P1_P2_Address_reg[6]/NET0131  & ~n2791 ;
  assign n2891 = \P1_P3_Address_reg[6]/NET0131  & n2791 ;
  assign n2892 = ~n2890 & ~n2891 ;
  assign n2893 = ~\P4_wr_reg/NET0131  & ~n2892 ;
  assign n2894 = \P4_addr_reg[6]/NET0131  & \P4_wr_reg/NET0131  ;
  assign n2895 = ~n2893 & ~n2894 ;
  assign n2896 = \P1_P2_Address_reg[5]/NET0131  & ~n2791 ;
  assign n2897 = \P1_P3_Address_reg[5]/NET0131  & n2791 ;
  assign n2898 = ~n2896 & ~n2897 ;
  assign n2899 = ~\P4_wr_reg/NET0131  & ~n2898 ;
  assign n2900 = \P4_addr_reg[5]/NET0131  & \P4_wr_reg/NET0131  ;
  assign n2901 = ~n2899 & ~n2900 ;
  assign n2902 = ~n2895 & ~n2901 ;
  assign n2903 = n2879 & ~n2902 ;
  assign n2904 = n2895 & n2901 ;
  assign n2905 = ~n2879 & ~n2904 ;
  assign n2906 = ~n2903 & ~n2905 ;
  assign n2907 = n2845 & n2906 ;
  assign n2908 = ~n2902 & ~n2904 ;
  assign n2909 = n2864 & n2908 ;
  assign n2910 = ~n2907 & ~n2909 ;
  assign n2911 = ~n2879 & ~n2910 ;
  assign n2912 = n2879 & n2910 ;
  assign n2913 = ~n2911 & ~n2912 ;
  assign n2914 = ~n2889 & ~n2913 ;
  assign n2915 = n2889 & n2913 ;
  assign n2923 = \P2_P2_Address_reg[8]/NET0131  & ~n2828 ;
  assign n2924 = \P2_P3_Address_reg[8]/NET0131  & n2828 ;
  assign n2925 = ~n2923 & ~n2924 ;
  assign n2926 = ~n2826 & ~n2925 ;
  assign n2927 = \P2_P1_Address_reg[8]/NET0131  & n2826 ;
  assign n2928 = ~n2926 & ~n2927 ;
  assign n2929 = ~n2872 & ~n2928 ;
  assign n2930 = ~\P4_wr_reg/NET0131  & ~n2838 ;
  assign n2931 = \P4_addr_reg[1]/NET0131  & \P4_wr_reg/NET0131  ;
  assign n2932 = ~n2930 & ~n2931 ;
  assign n2934 = ~n2929 & n2932 ;
  assign n2916 = \P2_P2_Address_reg[7]/NET0131  & ~n2828 ;
  assign n2917 = \P2_P3_Address_reg[7]/NET0131  & n2828 ;
  assign n2918 = ~n2916 & ~n2917 ;
  assign n2919 = ~n2826 & ~n2918 ;
  assign n2920 = \P2_P1_Address_reg[7]/NET0131  & n2826 ;
  assign n2921 = ~n2919 & ~n2920 ;
  assign n2922 = n2872 & ~n2921 ;
  assign n2933 = n2929 & ~n2932 ;
  assign n2935 = ~n2922 & ~n2933 ;
  assign n2936 = ~n2934 & n2935 ;
  assign n2937 = ~n2915 & ~n2936 ;
  assign n2938 = ~n2914 & ~n2937 ;
  assign n2939 = \P1_P2_Address_reg[3]/NET0131  & ~n2791 ;
  assign n2940 = \P1_P3_Address_reg[3]/NET0131  & n2791 ;
  assign n2941 = ~n2939 & ~n2940 ;
  assign n2942 = ~\P4_wr_reg/NET0131  & ~n2941 ;
  assign n2943 = \P4_addr_reg[3]/NET0131  & \P4_wr_reg/NET0131  ;
  assign n2944 = ~n2942 & ~n2943 ;
  assign n2945 = ~\P4_wr_reg/NET0131  & ~n2852 ;
  assign n2946 = \P4_addr_reg[2]/NET0131  & \P4_wr_reg/NET0131  ;
  assign n2947 = ~n2945 & ~n2946 ;
  assign n2948 = n2932 & n2947 ;
  assign n2949 = ~n2932 & ~n2947 ;
  assign n2950 = ~n2948 & ~n2949 ;
  assign n2951 = ~n2921 & n2950 ;
  assign n2952 = n2944 & ~n2949 ;
  assign n2953 = ~n2944 & ~n2948 ;
  assign n2954 = ~n2952 & ~n2953 ;
  assign n2955 = \P2_P2_Address_reg[6]/NET0131  & ~n2828 ;
  assign n2956 = \P2_P3_Address_reg[6]/NET0131  & n2828 ;
  assign n2957 = ~n2955 & ~n2956 ;
  assign n2958 = ~n2826 & ~n2957 ;
  assign n2959 = \P2_P1_Address_reg[6]/NET0131  & n2826 ;
  assign n2960 = ~n2958 & ~n2959 ;
  assign n2961 = n2954 & ~n2960 ;
  assign n2962 = ~n2951 & ~n2961 ;
  assign n2963 = n2944 & n2962 ;
  assign n2964 = ~n2944 & ~n2962 ;
  assign n2965 = ~n2963 & ~n2964 ;
  assign n2967 = \P2_P2_Address_reg[9]/NET0131  & ~n2828 ;
  assign n2968 = \P2_P3_Address_reg[9]/NET0131  & n2828 ;
  assign n2969 = ~n2967 & ~n2968 ;
  assign n2970 = ~n2826 & ~n2969 ;
  assign n2971 = \P2_P1_Address_reg[9]/NET0131  & n2826 ;
  assign n2972 = ~n2970 & ~n2971 ;
  assign n2973 = ~n2872 & ~n2972 ;
  assign n2975 = n2932 & ~n2973 ;
  assign n2966 = n2872 & ~n2928 ;
  assign n2974 = ~n2932 & n2973 ;
  assign n2976 = ~n2966 & ~n2974 ;
  assign n2977 = ~n2975 & n2976 ;
  assign n2978 = n2965 & n2977 ;
  assign n2979 = ~n2965 & ~n2977 ;
  assign n2980 = ~n2978 & ~n2979 ;
  assign n2981 = \P1_P2_Address_reg[9]/NET0131  & ~n2791 ;
  assign n2982 = \P1_P3_Address_reg[9]/NET0131  & n2791 ;
  assign n2983 = ~n2981 & ~n2982 ;
  assign n2984 = ~\P4_wr_reg/NET0131  & ~n2983 ;
  assign n2985 = \P4_addr_reg[9]/NET0131  & \P4_wr_reg/NET0131  ;
  assign n2986 = ~n2984 & ~n2985 ;
  assign n2987 = ~n2889 & ~n2986 ;
  assign n2988 = ~n2980 & ~n2987 ;
  assign n2989 = n2980 & n2987 ;
  assign n2990 = ~n2988 & ~n2989 ;
  assign n2991 = n2938 & ~n2990 ;
  assign n2992 = ~n2938 & n2990 ;
  assign n2993 = ~n2991 & ~n2992 ;
  assign n2994 = \P2_P2_Address_reg[5]/NET0131  & ~n2828 ;
  assign n2995 = \P2_P3_Address_reg[5]/NET0131  & n2828 ;
  assign n2996 = ~n2994 & ~n2995 ;
  assign n2997 = ~n2826 & ~n2996 ;
  assign n2998 = \P2_P1_Address_reg[5]/NET0131  & n2826 ;
  assign n2999 = ~n2997 & ~n2998 ;
  assign n3000 = n2950 & ~n2999 ;
  assign n3001 = ~\P2_P2_Address_reg[4]/NET0131  & ~n2828 ;
  assign n3002 = ~\P2_P3_Address_reg[4]/NET0131  & n2828 ;
  assign n3003 = ~n3001 & ~n3002 ;
  assign n3004 = ~n2826 & ~n3003 ;
  assign n3005 = ~\P2_P1_Address_reg[4]/NET0131  & n2826 ;
  assign n3006 = ~n3004 & ~n3005 ;
  assign n3007 = n2954 & n3006 ;
  assign n3008 = ~n3000 & ~n3007 ;
  assign n3009 = n2944 & n3008 ;
  assign n3010 = ~n2944 & ~n3008 ;
  assign n3011 = ~n3009 & ~n3010 ;
  assign n3013 = ~n2872 & ~n2921 ;
  assign n3015 = n2932 & ~n3013 ;
  assign n3012 = n2872 & ~n2960 ;
  assign n3014 = ~n2932 & n3013 ;
  assign n3016 = ~n3012 & ~n3014 ;
  assign n3017 = ~n3015 & n3016 ;
  assign n3018 = n3011 & n3017 ;
  assign n3019 = ~\P1_P2_Address_reg[4]/NET0131  & ~n2791 ;
  assign n3020 = ~\P1_P3_Address_reg[4]/NET0131  & n2791 ;
  assign n3021 = ~n3019 & ~n3020 ;
  assign n3022 = ~\P4_wr_reg/NET0131  & ~n3021 ;
  assign n3023 = ~\P4_addr_reg[4]/NET0131  & \P4_wr_reg/NET0131  ;
  assign n3024 = ~n3022 & ~n3023 ;
  assign n3025 = n2944 & ~n3024 ;
  assign n3026 = ~n2944 & n3024 ;
  assign n3027 = ~n3025 & ~n3026 ;
  assign n3028 = n3006 & n3027 ;
  assign n3029 = ~n2901 & n3025 ;
  assign n3030 = n2901 & n3026 ;
  assign n3031 = ~n3029 & ~n3030 ;
  assign n3032 = ~\P2_P3_Address_reg[3]/NET0131  & n2828 ;
  assign n3033 = ~\P2_P2_Address_reg[3]/NET0131  & ~n2828 ;
  assign n3034 = ~n3032 & ~n3033 ;
  assign n3035 = ~n2826 & ~n3034 ;
  assign n3036 = ~\P2_P1_Address_reg[3]/NET0131  & n2826 ;
  assign n3037 = ~n3035 & ~n3036 ;
  assign n3038 = ~n3031 & n3037 ;
  assign n3039 = ~n3028 & ~n3038 ;
  assign n3040 = ~n2901 & ~n3039 ;
  assign n3041 = n2901 & n3039 ;
  assign n3042 = ~n3040 & ~n3041 ;
  assign n3043 = n3018 & n3042 ;
  assign n3044 = ~n3018 & ~n3042 ;
  assign n3045 = n2954 & ~n2999 ;
  assign n3046 = n2950 & ~n2960 ;
  assign n3047 = ~n3045 & ~n3046 ;
  assign n3048 = ~n2944 & ~n3047 ;
  assign n3049 = n2944 & n3047 ;
  assign n3050 = ~n3048 & ~n3049 ;
  assign n3051 = ~n3044 & n3050 ;
  assign n3052 = ~n3043 & ~n3051 ;
  assign n3053 = ~n2993 & ~n3052 ;
  assign n3054 = n2993 & n3052 ;
  assign n3055 = n2908 & n3037 ;
  assign n3056 = n2864 & n2906 ;
  assign n3057 = ~n3055 & ~n3056 ;
  assign n3058 = n2879 & n3057 ;
  assign n3059 = ~n2879 & ~n3057 ;
  assign n3060 = ~n3058 & ~n3059 ;
  assign n3061 = ~n2999 & n3027 ;
  assign n3062 = n3006 & ~n3031 ;
  assign n3063 = ~n3061 & ~n3062 ;
  assign n3064 = n2901 & n3063 ;
  assign n3065 = ~n2901 & ~n3063 ;
  assign n3066 = ~n3064 & ~n3065 ;
  assign n3067 = n2845 & n2888 ;
  assign n3068 = n2886 & ~n2986 ;
  assign n3069 = n2887 & n2986 ;
  assign n3070 = ~n3068 & ~n3069 ;
  assign n3071 = ~n2834 & ~n3070 ;
  assign n3072 = ~n3067 & ~n3071 ;
  assign n3073 = n2986 & n3072 ;
  assign n3074 = ~n2986 & ~n3072 ;
  assign n3075 = ~n3073 & ~n3074 ;
  assign n3076 = n3066 & n3075 ;
  assign n3077 = ~n3066 & ~n3075 ;
  assign n3078 = ~n3076 & ~n3077 ;
  assign n3079 = n3060 & ~n3078 ;
  assign n3080 = ~n3060 & n3078 ;
  assign n3081 = ~n3079 & ~n3080 ;
  assign n3082 = ~n3054 & ~n3081 ;
  assign n3083 = ~n3053 & ~n3082 ;
  assign n3084 = n2864 & n2888 ;
  assign n3085 = n2845 & ~n3070 ;
  assign n3086 = ~n3084 & ~n3085 ;
  assign n3087 = n2986 & n3086 ;
  assign n3088 = ~n2986 & ~n3086 ;
  assign n3089 = ~n3087 & ~n3088 ;
  assign n3090 = ~n2960 & n3027 ;
  assign n3091 = ~n2999 & ~n3031 ;
  assign n3092 = ~n3090 & ~n3091 ;
  assign n3093 = n2901 & n3092 ;
  assign n3094 = ~n2901 & ~n3092 ;
  assign n3095 = ~n3093 & ~n3094 ;
  assign n3097 = \P2_P2_Address_reg[10]/NET0131  & ~n2828 ;
  assign n3098 = \P2_P3_Address_reg[10]/NET0131  & n2828 ;
  assign n3099 = ~n3097 & ~n3098 ;
  assign n3100 = ~n2826 & ~n3099 ;
  assign n3101 = \P2_P1_Address_reg[10]/NET0131  & n2826 ;
  assign n3102 = ~n3100 & ~n3101 ;
  assign n3103 = ~n2872 & ~n3102 ;
  assign n3105 = n2932 & ~n3103 ;
  assign n3096 = n2872 & ~n2972 ;
  assign n3104 = ~n2932 & n3103 ;
  assign n3106 = ~n3096 & ~n3104 ;
  assign n3107 = ~n3105 & n3106 ;
  assign n3108 = n3095 & n3107 ;
  assign n3109 = ~n3095 & ~n3107 ;
  assign n3110 = ~n3108 & ~n3109 ;
  assign n3111 = n3089 & ~n3110 ;
  assign n3112 = ~n3089 & n3110 ;
  assign n3113 = ~n3111 & ~n3112 ;
  assign n3114 = ~\P1_P2_Address_reg[10]/NET0131  & ~n2791 ;
  assign n3115 = ~\P1_P3_Address_reg[10]/NET0131  & n2791 ;
  assign n3116 = ~n3114 & ~n3115 ;
  assign n3117 = ~\P4_wr_reg/NET0131  & ~n3116 ;
  assign n3118 = ~\P4_addr_reg[10]/NET0131  & \P4_wr_reg/NET0131  ;
  assign n3119 = ~n3117 & ~n3118 ;
  assign n3120 = n2986 & ~n3119 ;
  assign n3121 = ~n2986 & n3119 ;
  assign n3122 = ~n3120 & ~n3121 ;
  assign n3123 = ~n2834 & n3122 ;
  assign n3124 = n2908 & n3006 ;
  assign n3125 = n2906 & n3037 ;
  assign n3126 = ~n3124 & ~n3125 ;
  assign n3127 = n2879 & n3126 ;
  assign n3128 = ~n2879 & ~n3126 ;
  assign n3129 = ~n3127 & ~n3128 ;
  assign n3130 = n3123 & n3129 ;
  assign n3131 = ~n3123 & ~n3129 ;
  assign n3132 = ~n3130 & ~n3131 ;
  assign n3133 = ~n2928 & n2950 ;
  assign n3134 = ~n2921 & n2954 ;
  assign n3135 = ~n3133 & ~n3134 ;
  assign n3136 = n2944 & n3135 ;
  assign n3137 = ~n2944 & ~n3135 ;
  assign n3138 = ~n3136 & ~n3137 ;
  assign n3139 = ~n3132 & n3138 ;
  assign n3140 = n3132 & ~n3138 ;
  assign n3141 = ~n3139 & ~n3140 ;
  assign n3142 = n3060 & ~n3077 ;
  assign n3143 = ~n3076 & ~n3142 ;
  assign n3144 = n3141 & n3143 ;
  assign n3145 = ~n3141 & ~n3143 ;
  assign n3146 = ~n3144 & ~n3145 ;
  assign n3147 = n2978 & ~n3146 ;
  assign n3148 = ~n2978 & n3146 ;
  assign n3149 = ~n3147 & ~n3148 ;
  assign n3150 = n3113 & n3149 ;
  assign n3151 = ~n3113 & ~n3149 ;
  assign n3152 = ~n3150 & ~n3151 ;
  assign n3153 = ~n2938 & ~n2989 ;
  assign n3154 = ~n2988 & ~n3153 ;
  assign n3155 = n3152 & ~n3154 ;
  assign n3156 = ~n3152 & n3154 ;
  assign n3157 = ~n3155 & ~n3156 ;
  assign n3158 = ~n3083 & ~n3157 ;
  assign n3159 = n3083 & n3157 ;
  assign n3160 = ~n3158 & ~n3159 ;
  assign n3161 = ~n2914 & ~n2915 ;
  assign n3162 = n2936 & ~n3161 ;
  assign n3163 = ~n2936 & n3161 ;
  assign n3164 = ~n3162 & ~n3163 ;
  assign n3165 = n3027 & n3037 ;
  assign n3166 = n2864 & ~n3031 ;
  assign n3167 = ~n3165 & ~n3166 ;
  assign n3168 = n2901 & n3167 ;
  assign n3169 = ~n2901 & ~n3167 ;
  assign n3170 = ~n3168 & ~n3169 ;
  assign n3171 = ~n2834 & n2908 ;
  assign n3172 = ~n2879 & ~n3171 ;
  assign n3173 = n3170 & n3172 ;
  assign n3174 = ~n3170 & ~n3172 ;
  assign n3175 = n2845 & n2908 ;
  assign n3176 = ~n2834 & n2906 ;
  assign n3177 = ~n3175 & ~n3176 ;
  assign n3178 = n2879 & n3177 ;
  assign n3179 = ~n2879 & ~n3177 ;
  assign n3180 = ~n3178 & ~n3179 ;
  assign n3181 = ~n3174 & n3180 ;
  assign n3182 = ~n3173 & ~n3181 ;
  assign n3183 = ~n3164 & ~n3182 ;
  assign n3184 = n3164 & n3182 ;
  assign n3185 = ~n3043 & ~n3044 ;
  assign n3186 = ~n3050 & n3185 ;
  assign n3187 = n3050 & ~n3185 ;
  assign n3188 = ~n3186 & ~n3187 ;
  assign n3189 = ~n3184 & ~n3188 ;
  assign n3190 = ~n3183 & ~n3189 ;
  assign n3191 = ~n3053 & ~n3054 ;
  assign n3192 = ~n3081 & n3191 ;
  assign n3193 = n3081 & ~n3191 ;
  assign n3194 = ~n3192 & ~n3193 ;
  assign n3195 = ~n3190 & n3194 ;
  assign n3196 = n3190 & ~n3194 ;
  assign n3197 = n2954 & n3037 ;
  assign n3198 = n2950 & n3006 ;
  assign n3199 = ~n3197 & ~n3198 ;
  assign n3200 = ~n2944 & ~n3199 ;
  assign n3201 = n2944 & n3199 ;
  assign n3202 = ~n3200 & ~n3201 ;
  assign n3204 = ~n2872 & ~n2960 ;
  assign n3206 = n2932 & ~n3204 ;
  assign n3203 = n2872 & ~n2999 ;
  assign n3205 = ~n2932 & n3204 ;
  assign n3207 = ~n3203 & ~n3205 ;
  assign n3208 = ~n3206 & n3207 ;
  assign n3209 = n3202 & n3208 ;
  assign n3210 = ~n3171 & ~n3209 ;
  assign n3211 = ~n3202 & ~n3208 ;
  assign n3212 = ~n3210 & ~n3211 ;
  assign n3213 = ~n3173 & ~n3174 ;
  assign n3214 = ~n3180 & n3213 ;
  assign n3215 = n3180 & ~n3213 ;
  assign n3216 = ~n3214 & ~n3215 ;
  assign n3217 = ~n3212 & n3216 ;
  assign n3218 = n3212 & ~n3216 ;
  assign n3219 = ~n3011 & ~n3017 ;
  assign n3220 = ~n3018 & ~n3219 ;
  assign n3221 = ~n3218 & ~n3220 ;
  assign n3222 = ~n3217 & ~n3221 ;
  assign n3223 = ~n3183 & ~n3184 ;
  assign n3224 = ~n3188 & n3223 ;
  assign n3225 = n3188 & ~n3223 ;
  assign n3226 = ~n3224 & ~n3225 ;
  assign n3227 = n3222 & n3226 ;
  assign n3228 = ~n3222 & ~n3226 ;
  assign n3229 = n2950 & n3037 ;
  assign n3230 = n2864 & n2954 ;
  assign n3231 = ~n3229 & ~n3230 ;
  assign n3232 = n2944 & n3231 ;
  assign n3233 = ~n2944 & ~n3231 ;
  assign n3234 = ~n3232 & ~n3233 ;
  assign n3236 = ~n2872 & ~n2999 ;
  assign n3238 = n2932 & ~n3236 ;
  assign n3235 = n2872 & n3006 ;
  assign n3237 = ~n2932 & n3236 ;
  assign n3239 = ~n3235 & ~n3237 ;
  assign n3240 = ~n3238 & n3239 ;
  assign n3241 = n3234 & n3240 ;
  assign n3242 = n2864 & n3027 ;
  assign n3243 = n2845 & ~n3031 ;
  assign n3244 = ~n3242 & ~n3243 ;
  assign n3245 = n2901 & n3244 ;
  assign n3246 = ~n2901 & ~n3244 ;
  assign n3247 = ~n3245 & ~n3246 ;
  assign n3248 = n3241 & n3247 ;
  assign n3249 = ~n3241 & ~n3247 ;
  assign n3250 = ~n3209 & ~n3211 ;
  assign n3251 = n3171 & ~n3250 ;
  assign n3252 = ~n3171 & n3250 ;
  assign n3253 = ~n3251 & ~n3252 ;
  assign n3254 = ~n3249 & ~n3253 ;
  assign n3255 = ~n3248 & ~n3254 ;
  assign n3256 = ~n3217 & ~n3218 ;
  assign n3257 = ~n3220 & n3256 ;
  assign n3258 = n3220 & ~n3256 ;
  assign n3259 = ~n3257 & ~n3258 ;
  assign n3260 = ~n3255 & ~n3259 ;
  assign n3261 = n3255 & n3259 ;
  assign n3262 = ~n3234 & ~n3240 ;
  assign n3263 = ~n3241 & ~n3262 ;
  assign n3264 = n2845 & n3027 ;
  assign n3265 = ~n2834 & ~n3031 ;
  assign n3266 = ~n3264 & ~n3265 ;
  assign n3267 = ~n2901 & n3266 ;
  assign n3268 = ~n2834 & n3027 ;
  assign n3269 = ~n2901 & n3268 ;
  assign n3270 = ~n3266 & ~n3269 ;
  assign n3271 = ~n3267 & ~n3270 ;
  assign n3272 = n3263 & ~n3271 ;
  assign n3273 = n3267 & ~n3268 ;
  assign n3274 = ~n3272 & ~n3273 ;
  assign n3275 = ~n3248 & ~n3249 ;
  assign n3276 = ~n3253 & n3275 ;
  assign n3277 = n3253 & ~n3275 ;
  assign n3278 = ~n3276 & ~n3277 ;
  assign n3279 = n3274 & ~n3278 ;
  assign n3280 = ~n3274 & n3278 ;
  assign n3281 = n2845 & n2954 ;
  assign n3282 = n2864 & n2950 ;
  assign n3283 = ~n3281 & ~n3282 ;
  assign n3284 = ~n2944 & ~n3283 ;
  assign n3285 = n2944 & n3283 ;
  assign n3286 = ~n3284 & ~n3285 ;
  assign n3288 = ~n2872 & n3006 ;
  assign n3290 = n2932 & ~n3288 ;
  assign n3287 = n2872 & n3037 ;
  assign n3289 = ~n2932 & n3288 ;
  assign n3291 = ~n3287 & ~n3289 ;
  assign n3292 = ~n3290 & n3291 ;
  assign n3293 = n3286 & n3292 ;
  assign n3294 = ~n3268 & ~n3293 ;
  assign n3295 = ~n3286 & ~n3292 ;
  assign n3296 = ~n3294 & ~n3295 ;
  assign n3297 = ~n3271 & ~n3273 ;
  assign n3298 = n3263 & ~n3297 ;
  assign n3299 = ~n3263 & n3297 ;
  assign n3300 = ~n3298 & ~n3299 ;
  assign n3301 = ~n3296 & n3300 ;
  assign n3302 = n3296 & ~n3300 ;
  assign n3303 = ~n2834 & n2950 ;
  assign n3304 = ~n2944 & ~n3303 ;
  assign n3306 = ~n2872 & n3037 ;
  assign n3308 = n2932 & ~n3306 ;
  assign n3305 = n2864 & n2872 ;
  assign n3307 = ~n2932 & n3306 ;
  assign n3309 = ~n3305 & ~n3307 ;
  assign n3310 = ~n3308 & n3309 ;
  assign n3311 = n3304 & n3310 ;
  assign n3312 = ~n3293 & ~n3295 ;
  assign n3313 = n3268 & ~n3312 ;
  assign n3314 = ~n3268 & n3312 ;
  assign n3315 = ~n3313 & ~n3314 ;
  assign n3316 = ~n3311 & n3315 ;
  assign n3317 = n3311 & ~n3315 ;
  assign n3318 = ~n3304 & ~n3310 ;
  assign n3319 = ~n3311 & ~n3318 ;
  assign n3320 = ~n2834 & n2954 ;
  assign n3321 = n2845 & n2950 ;
  assign n3322 = ~n3320 & ~n3321 ;
  assign n3323 = ~n2944 & ~n3322 ;
  assign n3324 = n2944 & n3322 ;
  assign n3325 = ~n3323 & ~n3324 ;
  assign n3326 = ~n3319 & ~n3325 ;
  assign n3327 = n3319 & n3325 ;
  assign n3328 = n2845 & ~n2872 ;
  assign n3329 = n2834 & ~n2932 ;
  assign n3330 = ~n3328 & n3329 ;
  assign n3331 = ~n3303 & ~n3330 ;
  assign n3333 = n2864 & ~n2872 ;
  assign n3335 = n2932 & ~n3333 ;
  assign n3332 = n2845 & n2872 ;
  assign n3334 = ~n2932 & n3333 ;
  assign n3336 = ~n3332 & ~n3334 ;
  assign n3337 = ~n3335 & n3336 ;
  assign n3338 = ~n3331 & n3337 ;
  assign n3339 = ~n3327 & ~n3338 ;
  assign n3340 = ~n3326 & ~n3339 ;
  assign n3341 = ~n3317 & ~n3340 ;
  assign n3342 = ~n3316 & ~n3341 ;
  assign n3343 = ~n3302 & ~n3342 ;
  assign n3344 = ~n3301 & ~n3343 ;
  assign n3345 = ~n3280 & ~n3344 ;
  assign n3346 = ~n3279 & ~n3345 ;
  assign n3347 = ~n3261 & n3346 ;
  assign n3348 = ~n3260 & ~n3347 ;
  assign n3349 = ~n3228 & ~n3348 ;
  assign n3350 = ~n3227 & ~n3349 ;
  assign n3351 = ~n3196 & ~n3350 ;
  assign n3352 = ~n3195 & ~n3351 ;
  assign n3353 = n3160 & ~n3352 ;
  assign n3354 = ~n3160 & n3352 ;
  assign n3355 = ~n3353 & ~n3354 ;
  assign n3356 = ~n3150 & n3154 ;
  assign n3357 = ~n3151 & ~n3356 ;
  assign n3358 = \P1_P2_Address_reg[11]/NET0131  & ~n2791 ;
  assign n3359 = \P1_P3_Address_reg[11]/NET0131  & n2791 ;
  assign n3360 = ~n3358 & ~n3359 ;
  assign n3361 = ~\P4_wr_reg/NET0131  & ~n3360 ;
  assign n3362 = \P4_addr_reg[11]/NET0131  & \P4_wr_reg/NET0131  ;
  assign n3363 = ~n3361 & ~n3362 ;
  assign n3364 = n2845 & n3122 ;
  assign n3365 = n3120 & ~n3363 ;
  assign n3366 = n3121 & n3363 ;
  assign n3367 = ~n3365 & ~n3366 ;
  assign n3368 = ~n2834 & ~n3367 ;
  assign n3369 = ~n3364 & ~n3368 ;
  assign n3370 = ~n3363 & ~n3369 ;
  assign n3371 = n3363 & n3369 ;
  assign n3372 = ~n3370 & ~n3371 ;
  assign n3373 = n2950 & ~n2972 ;
  assign n3374 = ~n2928 & n2954 ;
  assign n3375 = ~n3373 & ~n3374 ;
  assign n3376 = n2944 & n3375 ;
  assign n3377 = ~n2944 & ~n3375 ;
  assign n3378 = ~n3376 & ~n3377 ;
  assign n3380 = \P2_P2_Address_reg[11]/NET0131  & ~n2828 ;
  assign n3381 = \P2_P3_Address_reg[11]/NET0131  & n2828 ;
  assign n3382 = ~n3380 & ~n3381 ;
  assign n3383 = ~n2826 & ~n3382 ;
  assign n3384 = \P2_P1_Address_reg[11]/NET0131  & n2826 ;
  assign n3385 = ~n3383 & ~n3384 ;
  assign n3386 = ~n2872 & ~n3385 ;
  assign n3388 = n2932 & ~n3386 ;
  assign n3379 = n2872 & ~n3102 ;
  assign n3387 = ~n2932 & n3386 ;
  assign n3389 = ~n3379 & ~n3387 ;
  assign n3390 = ~n3388 & n3389 ;
  assign n3391 = n3378 & n3390 ;
  assign n3392 = ~n3378 & ~n3390 ;
  assign n3393 = ~n3391 & ~n3392 ;
  assign n3394 = ~n3123 & ~n3363 ;
  assign n3395 = ~n3393 & ~n3394 ;
  assign n3396 = n3393 & n3394 ;
  assign n3397 = ~n3395 & ~n3396 ;
  assign n3398 = n3372 & ~n3397 ;
  assign n3399 = ~n3372 & n3397 ;
  assign n3400 = ~n3398 & ~n3399 ;
  assign n3401 = n2978 & ~n3144 ;
  assign n3402 = ~n3145 & ~n3401 ;
  assign n3403 = n3400 & n3402 ;
  assign n3404 = ~n3400 & ~n3402 ;
  assign n3405 = ~n3403 & ~n3404 ;
  assign n3406 = n2908 & ~n2999 ;
  assign n3407 = n2906 & n3006 ;
  assign n3408 = ~n3406 & ~n3407 ;
  assign n3409 = n2879 & n3408 ;
  assign n3410 = ~n2879 & ~n3408 ;
  assign n3411 = ~n3409 & ~n3410 ;
  assign n3412 = ~n2921 & n3027 ;
  assign n3413 = ~n2960 & ~n3031 ;
  assign n3414 = ~n3412 & ~n3413 ;
  assign n3415 = n2901 & n3414 ;
  assign n3416 = ~n2901 & ~n3414 ;
  assign n3417 = ~n3415 & ~n3416 ;
  assign n3418 = n2888 & n3037 ;
  assign n3419 = n2864 & ~n3070 ;
  assign n3420 = ~n3418 & ~n3419 ;
  assign n3421 = n2986 & n3420 ;
  assign n3422 = ~n2986 & ~n3420 ;
  assign n3423 = ~n3421 & ~n3422 ;
  assign n3424 = n3417 & n3423 ;
  assign n3425 = ~n3417 & ~n3423 ;
  assign n3426 = ~n3424 & ~n3425 ;
  assign n3427 = n3411 & ~n3426 ;
  assign n3428 = ~n3411 & n3426 ;
  assign n3429 = ~n3427 & ~n3428 ;
  assign n3430 = n3089 & ~n3109 ;
  assign n3431 = ~n3108 & ~n3430 ;
  assign n3432 = n3429 & n3431 ;
  assign n3433 = ~n3429 & ~n3431 ;
  assign n3434 = ~n3432 & ~n3433 ;
  assign n3435 = ~n3131 & n3138 ;
  assign n3436 = ~n3130 & ~n3435 ;
  assign n3437 = n3434 & ~n3436 ;
  assign n3438 = ~n3434 & n3436 ;
  assign n3439 = ~n3437 & ~n3438 ;
  assign n3440 = n3405 & n3439 ;
  assign n3441 = ~n3405 & ~n3439 ;
  assign n3442 = ~n3440 & ~n3441 ;
  assign n3443 = ~n3357 & n3442 ;
  assign n3444 = n3357 & ~n3442 ;
  assign n3445 = ~n3443 & ~n3444 ;
  assign n3446 = ~n3159 & ~n3352 ;
  assign n3447 = ~n3158 & ~n3446 ;
  assign n3448 = n3445 & n3447 ;
  assign n3449 = ~n3445 & ~n3447 ;
  assign n3450 = ~n3448 & ~n3449 ;
  assign n3451 = ~n3404 & ~n3439 ;
  assign n3452 = ~n3403 & ~n3451 ;
  assign n3453 = ~n2928 & n3027 ;
  assign n3454 = ~n2921 & ~n3031 ;
  assign n3455 = ~n3453 & ~n3454 ;
  assign n3456 = ~n2901 & ~n3455 ;
  assign n3457 = n2901 & n3455 ;
  assign n3458 = ~n3456 & ~n3457 ;
  assign n3459 = n3411 & ~n3425 ;
  assign n3460 = ~n3424 & ~n3459 ;
  assign n3461 = ~n3391 & n3460 ;
  assign n3462 = n3391 & ~n3460 ;
  assign n3463 = ~n3461 & ~n3462 ;
  assign n3464 = n3458 & n3463 ;
  assign n3465 = ~n3458 & ~n3463 ;
  assign n3466 = ~n3464 & ~n3465 ;
  assign n3467 = n2864 & n3122 ;
  assign n3468 = n2845 & ~n3367 ;
  assign n3469 = ~n3467 & ~n3468 ;
  assign n3470 = n3363 & n3469 ;
  assign n3471 = ~n3363 & ~n3469 ;
  assign n3472 = ~n3470 & ~n3471 ;
  assign n3473 = n2888 & n3006 ;
  assign n3474 = n3037 & ~n3070 ;
  assign n3475 = ~n3473 & ~n3474 ;
  assign n3476 = n2986 & n3475 ;
  assign n3477 = ~n2986 & ~n3475 ;
  assign n3478 = ~n3476 & ~n3477 ;
  assign n3480 = \P2_P2_Address_reg[12]/NET0131  & ~n2828 ;
  assign n3481 = \P2_P3_Address_reg[12]/NET0131  & n2828 ;
  assign n3482 = ~n3480 & ~n3481 ;
  assign n3483 = ~n2826 & ~n3482 ;
  assign n3484 = \P2_P1_Address_reg[12]/NET0131  & n2826 ;
  assign n3485 = ~n3483 & ~n3484 ;
  assign n3486 = ~n2872 & ~n3485 ;
  assign n3488 = n2932 & ~n3486 ;
  assign n3479 = n2872 & ~n3385 ;
  assign n3487 = ~n2932 & n3486 ;
  assign n3489 = ~n3479 & ~n3487 ;
  assign n3490 = ~n3488 & n3489 ;
  assign n3491 = n3478 & n3490 ;
  assign n3492 = ~n3478 & ~n3490 ;
  assign n3493 = ~n3491 & ~n3492 ;
  assign n3494 = n3472 & ~n3493 ;
  assign n3495 = ~n3472 & n3493 ;
  assign n3496 = ~n3494 & ~n3495 ;
  assign n3497 = ~n3372 & ~n3396 ;
  assign n3498 = ~n3395 & ~n3497 ;
  assign n3499 = n3496 & ~n3498 ;
  assign n3500 = ~n3496 & n3498 ;
  assign n3501 = ~n3499 & ~n3500 ;
  assign n3502 = ~\P1_P2_Address_reg[12]/NET0131  & ~n2791 ;
  assign n3503 = ~\P1_P3_Address_reg[12]/NET0131  & n2791 ;
  assign n3504 = ~n3502 & ~n3503 ;
  assign n3505 = ~\P4_wr_reg/NET0131  & ~n3504 ;
  assign n3506 = ~\P4_addr_reg[12]/NET0131  & \P4_wr_reg/NET0131  ;
  assign n3507 = ~n3505 & ~n3506 ;
  assign n3508 = n3363 & ~n3507 ;
  assign n3509 = ~n3363 & n3507 ;
  assign n3510 = ~n3508 & ~n3509 ;
  assign n3511 = ~n2834 & n3510 ;
  assign n3512 = n2908 & ~n2960 ;
  assign n3513 = n2906 & ~n2999 ;
  assign n3514 = ~n3512 & ~n3513 ;
  assign n3515 = n2879 & n3514 ;
  assign n3516 = ~n2879 & ~n3514 ;
  assign n3517 = ~n3515 & ~n3516 ;
  assign n3518 = n3511 & n3517 ;
  assign n3519 = ~n3511 & ~n3517 ;
  assign n3520 = ~n3518 & ~n3519 ;
  assign n3521 = n2950 & ~n3102 ;
  assign n3522 = n2954 & ~n2972 ;
  assign n3523 = ~n3521 & ~n3522 ;
  assign n3524 = n2944 & n3523 ;
  assign n3525 = ~n2944 & ~n3523 ;
  assign n3526 = ~n3524 & ~n3525 ;
  assign n3527 = ~n3520 & n3526 ;
  assign n3528 = n3520 & ~n3526 ;
  assign n3529 = ~n3527 & ~n3528 ;
  assign n3530 = n3501 & ~n3529 ;
  assign n3531 = ~n3501 & n3529 ;
  assign n3532 = ~n3530 & ~n3531 ;
  assign n3533 = ~n3466 & ~n3532 ;
  assign n3534 = n3466 & n3532 ;
  assign n3535 = ~n3533 & ~n3534 ;
  assign n3536 = ~n3432 & ~n3436 ;
  assign n3537 = ~n3433 & ~n3536 ;
  assign n3538 = n3535 & n3537 ;
  assign n3539 = ~n3535 & ~n3537 ;
  assign n3540 = ~n3538 & ~n3539 ;
  assign n3541 = n3452 & ~n3540 ;
  assign n3542 = ~n3452 & n3540 ;
  assign n3543 = ~n3541 & ~n3542 ;
  assign n3544 = ~n3444 & ~n3447 ;
  assign n3545 = ~n3443 & ~n3544 ;
  assign n3546 = n3543 & n3545 ;
  assign n3547 = ~n3543 & ~n3545 ;
  assign n3548 = ~n3546 & ~n3547 ;
  assign n3549 = ~n3533 & ~n3537 ;
  assign n3550 = ~n3534 & ~n3549 ;
  assign n3551 = n2950 & ~n3385 ;
  assign n3552 = n2954 & ~n3102 ;
  assign n3553 = ~n3551 & ~n3552 ;
  assign n3554 = n2944 & n3553 ;
  assign n3555 = ~n2944 & ~n3553 ;
  assign n3556 = ~n3554 & ~n3555 ;
  assign n3558 = \P2_P2_Address_reg[13]/NET0131  & ~n2828 ;
  assign n3559 = \P2_P3_Address_reg[13]/NET0131  & n2828 ;
  assign n3560 = ~n3558 & ~n3559 ;
  assign n3561 = ~n2826 & ~n3560 ;
  assign n3562 = \P2_P1_Address_reg[13]/NET0131  & n2826 ;
  assign n3563 = ~n3561 & ~n3562 ;
  assign n3564 = ~n2872 & ~n3563 ;
  assign n3566 = n2932 & ~n3564 ;
  assign n3557 = n2872 & ~n3485 ;
  assign n3565 = ~n2932 & n3564 ;
  assign n3567 = ~n3557 & ~n3565 ;
  assign n3568 = ~n3566 & n3567 ;
  assign n3569 = n3556 & n3568 ;
  assign n3570 = ~n3556 & ~n3568 ;
  assign n3571 = ~n3569 & ~n3570 ;
  assign n3572 = ~n3519 & n3526 ;
  assign n3573 = ~n3518 & ~n3572 ;
  assign n3574 = ~n3571 & n3573 ;
  assign n3575 = n3571 & ~n3573 ;
  assign n3576 = ~n3574 & ~n3575 ;
  assign n3577 = n3472 & ~n3492 ;
  assign n3578 = ~n3491 & ~n3577 ;
  assign n3579 = n3576 & ~n3578 ;
  assign n3580 = ~n3576 & n3578 ;
  assign n3581 = ~n3579 & ~n3580 ;
  assign n3582 = \P1_P2_Address_reg[13]/NET0131  & ~n2791 ;
  assign n3583 = \P1_P3_Address_reg[13]/NET0131  & n2791 ;
  assign n3584 = ~n3582 & ~n3583 ;
  assign n3585 = ~\P4_wr_reg/NET0131  & ~n3584 ;
  assign n3586 = \P4_addr_reg[13]/NET0131  & \P4_wr_reg/NET0131  ;
  assign n3587 = ~n3585 & ~n3586 ;
  assign n3588 = ~n3511 & ~n3587 ;
  assign n3589 = n2888 & ~n2999 ;
  assign n3590 = n3006 & ~n3070 ;
  assign n3591 = ~n3589 & ~n3590 ;
  assign n3592 = n2986 & n3591 ;
  assign n3593 = ~n2986 & ~n3591 ;
  assign n3594 = ~n3592 & ~n3593 ;
  assign n3595 = n3588 & n3594 ;
  assign n3596 = ~n3588 & ~n3594 ;
  assign n3597 = ~n3595 & ~n3596 ;
  assign n3598 = n2908 & ~n2921 ;
  assign n3599 = n2906 & ~n2960 ;
  assign n3600 = ~n3598 & ~n3599 ;
  assign n3601 = n2879 & n3600 ;
  assign n3602 = ~n2879 & ~n3600 ;
  assign n3603 = ~n3601 & ~n3602 ;
  assign n3604 = ~n3597 & n3603 ;
  assign n3605 = n3597 & ~n3603 ;
  assign n3606 = ~n3604 & ~n3605 ;
  assign n3607 = ~n3458 & ~n3462 ;
  assign n3608 = ~n3461 & ~n3607 ;
  assign n3609 = n3606 & ~n3608 ;
  assign n3610 = ~n3606 & n3608 ;
  assign n3611 = ~n3609 & ~n3610 ;
  assign n3612 = ~n2972 & n3027 ;
  assign n3613 = ~n2928 & ~n3031 ;
  assign n3614 = ~n3612 & ~n3613 ;
  assign n3615 = n2901 & n3614 ;
  assign n3616 = ~n2901 & ~n3614 ;
  assign n3617 = ~n3615 & ~n3616 ;
  assign n3618 = n2845 & n3510 ;
  assign n3619 = n3363 & n3587 ;
  assign n3620 = ~n3363 & ~n3587 ;
  assign n3621 = ~n3619 & ~n3620 ;
  assign n3622 = ~n3510 & n3621 ;
  assign n3623 = ~n2834 & n3622 ;
  assign n3624 = ~n3618 & ~n3623 ;
  assign n3625 = n3587 & n3624 ;
  assign n3626 = ~n3587 & ~n3624 ;
  assign n3627 = ~n3625 & ~n3626 ;
  assign n3628 = n3037 & n3122 ;
  assign n3629 = n2864 & ~n3367 ;
  assign n3630 = ~n3628 & ~n3629 ;
  assign n3631 = n3363 & n3630 ;
  assign n3632 = ~n3363 & ~n3630 ;
  assign n3633 = ~n3631 & ~n3632 ;
  assign n3634 = n3627 & n3633 ;
  assign n3635 = ~n3627 & ~n3633 ;
  assign n3636 = ~n3634 & ~n3635 ;
  assign n3637 = n3617 & ~n3636 ;
  assign n3638 = ~n3617 & n3636 ;
  assign n3639 = ~n3637 & ~n3638 ;
  assign n3640 = n3611 & ~n3639 ;
  assign n3641 = ~n3611 & n3639 ;
  assign n3642 = ~n3640 & ~n3641 ;
  assign n3643 = ~n3581 & ~n3642 ;
  assign n3644 = n3581 & n3642 ;
  assign n3645 = ~n3643 & ~n3644 ;
  assign n3646 = ~n3500 & n3529 ;
  assign n3647 = ~n3499 & ~n3646 ;
  assign n3648 = n3645 & ~n3647 ;
  assign n3649 = ~n3645 & n3647 ;
  assign n3650 = ~n3648 & ~n3649 ;
  assign n3651 = ~n3550 & ~n3650 ;
  assign n3652 = n3550 & n3650 ;
  assign n3653 = ~n3651 & ~n3652 ;
  assign n3654 = ~n3542 & ~n3545 ;
  assign n3655 = ~n3541 & ~n3654 ;
  assign n3656 = n3653 & n3655 ;
  assign n3657 = ~n3653 & ~n3655 ;
  assign n3658 = ~n3656 & ~n3657 ;
  assign n3659 = ~n3644 & ~n3647 ;
  assign n3660 = ~n3643 & ~n3659 ;
  assign n3661 = n2864 & n3510 ;
  assign n3662 = n2845 & n3622 ;
  assign n3663 = ~n3661 & ~n3662 ;
  assign n3664 = ~n3587 & ~n3663 ;
  assign n3665 = n3587 & n3663 ;
  assign n3666 = ~n3664 & ~n3665 ;
  assign n3667 = n3006 & n3122 ;
  assign n3668 = n3037 & ~n3367 ;
  assign n3669 = ~n3667 & ~n3668 ;
  assign n3670 = ~n3363 & ~n3669 ;
  assign n3671 = n3363 & n3669 ;
  assign n3672 = ~n3670 & ~n3671 ;
  assign n3673 = n3569 & n3672 ;
  assign n3674 = ~n3569 & ~n3672 ;
  assign n3675 = ~n3673 & ~n3674 ;
  assign n3676 = n3666 & ~n3675 ;
  assign n3677 = ~n3666 & n3675 ;
  assign n3678 = ~n3676 & ~n3677 ;
  assign n3679 = ~n3574 & ~n3578 ;
  assign n3680 = ~n3575 & ~n3679 ;
  assign n3681 = n3678 & n3680 ;
  assign n3682 = ~n3678 & ~n3680 ;
  assign n3683 = ~n3681 & ~n3682 ;
  assign n3684 = n2950 & ~n3485 ;
  assign n3685 = n2954 & ~n3385 ;
  assign n3686 = ~n3684 & ~n3685 ;
  assign n3687 = n2944 & n3686 ;
  assign n3688 = ~n2944 & ~n3686 ;
  assign n3689 = ~n3687 & ~n3688 ;
  assign n3690 = n2888 & ~n2960 ;
  assign n3691 = ~n2999 & ~n3070 ;
  assign n3692 = ~n3690 & ~n3691 ;
  assign n3693 = n2986 & n3692 ;
  assign n3694 = ~n2986 & ~n3692 ;
  assign n3695 = ~n3693 & ~n3694 ;
  assign n3696 = n3689 & n3695 ;
  assign n3697 = ~n3689 & ~n3695 ;
  assign n3698 = ~n3696 & ~n3697 ;
  assign n3699 = n3027 & ~n3102 ;
  assign n3700 = ~n2972 & ~n3031 ;
  assign n3701 = ~n3699 & ~n3700 ;
  assign n3702 = n2901 & n3701 ;
  assign n3703 = ~n2901 & ~n3701 ;
  assign n3704 = ~n3702 & ~n3703 ;
  assign n3705 = ~n3698 & n3704 ;
  assign n3706 = n3698 & ~n3704 ;
  assign n3707 = ~n3705 & ~n3706 ;
  assign n3708 = n3683 & n3707 ;
  assign n3709 = ~n3683 & ~n3707 ;
  assign n3710 = ~n3708 & ~n3709 ;
  assign n3711 = ~\P1_P2_Address_reg[14]/NET0131  & ~n2791 ;
  assign n3712 = ~\P1_P3_Address_reg[14]/NET0131  & n2791 ;
  assign n3713 = ~n3711 & ~n3712 ;
  assign n3714 = ~\P4_wr_reg/NET0131  & ~n3713 ;
  assign n3715 = ~\P4_addr_reg[14]/NET0131  & \P4_wr_reg/NET0131  ;
  assign n3716 = ~n3714 & ~n3715 ;
  assign n3717 = n3587 & ~n3716 ;
  assign n3718 = ~n3587 & n3716 ;
  assign n3719 = ~n3717 & ~n3718 ;
  assign n3720 = ~n2834 & n3719 ;
  assign n3721 = n2906 & ~n2921 ;
  assign n3722 = n2908 & ~n2928 ;
  assign n3723 = ~n3721 & ~n3722 ;
  assign n3724 = ~n2879 & ~n3723 ;
  assign n3725 = n2879 & n3723 ;
  assign n3726 = ~n3724 & ~n3725 ;
  assign n3727 = n3720 & n3726 ;
  assign n3728 = ~n3720 & ~n3726 ;
  assign n3729 = ~n3727 & ~n3728 ;
  assign n3731 = \P2_P2_Address_reg[14]/NET0131  & ~n2828 ;
  assign n3732 = \P2_P3_Address_reg[14]/NET0131  & n2828 ;
  assign n3733 = ~n3731 & ~n3732 ;
  assign n3734 = ~n2826 & ~n3733 ;
  assign n3735 = \P2_P1_Address_reg[14]/NET0131  & n2826 ;
  assign n3736 = ~n3734 & ~n3735 ;
  assign n3737 = ~n2872 & ~n3736 ;
  assign n3739 = n2932 & ~n3737 ;
  assign n3730 = n2872 & ~n3563 ;
  assign n3738 = ~n2932 & n3737 ;
  assign n3740 = ~n3730 & ~n3738 ;
  assign n3741 = ~n3739 & n3740 ;
  assign n3742 = ~n3729 & n3741 ;
  assign n3743 = n3729 & ~n3741 ;
  assign n3744 = ~n3742 & ~n3743 ;
  assign n3745 = ~n3596 & n3603 ;
  assign n3746 = ~n3595 & ~n3745 ;
  assign n3747 = n3744 & n3746 ;
  assign n3748 = ~n3744 & ~n3746 ;
  assign n3749 = ~n3747 & ~n3748 ;
  assign n3750 = n3617 & ~n3635 ;
  assign n3751 = ~n3634 & ~n3750 ;
  assign n3752 = n3749 & ~n3751 ;
  assign n3753 = ~n3749 & n3751 ;
  assign n3754 = ~n3752 & ~n3753 ;
  assign n3755 = n3710 & ~n3754 ;
  assign n3756 = ~n3710 & n3754 ;
  assign n3757 = ~n3755 & ~n3756 ;
  assign n3758 = ~n3610 & n3639 ;
  assign n3759 = ~n3609 & ~n3758 ;
  assign n3760 = n3757 & n3759 ;
  assign n3761 = ~n3757 & ~n3759 ;
  assign n3762 = ~n3760 & ~n3761 ;
  assign n3763 = n3660 & n3762 ;
  assign n3764 = ~n3660 & ~n3762 ;
  assign n3765 = ~n3763 & ~n3764 ;
  assign n3766 = ~n3652 & ~n3655 ;
  assign n3767 = ~n3651 & ~n3766 ;
  assign n3768 = n3765 & ~n3767 ;
  assign n3769 = ~n3765 & n3767 ;
  assign n3770 = ~n3768 & ~n3769 ;
  assign n3771 = ~n3681 & ~n3707 ;
  assign n3772 = ~n3682 & ~n3771 ;
  assign n3773 = n2888 & ~n2921 ;
  assign n3774 = ~n2960 & ~n3070 ;
  assign n3775 = ~n3773 & ~n3774 ;
  assign n3776 = n2986 & n3775 ;
  assign n3777 = ~n2986 & ~n3775 ;
  assign n3778 = ~n3776 & ~n3777 ;
  assign n3779 = ~n2999 & n3122 ;
  assign n3780 = n3006 & ~n3367 ;
  assign n3781 = ~n3779 & ~n3780 ;
  assign n3782 = n3363 & n3781 ;
  assign n3783 = ~n3363 & ~n3781 ;
  assign n3784 = ~n3782 & ~n3783 ;
  assign n3785 = n3027 & ~n3385 ;
  assign n3786 = ~n3031 & ~n3102 ;
  assign n3787 = ~n3785 & ~n3786 ;
  assign n3788 = n2901 & n3787 ;
  assign n3789 = ~n2901 & ~n3787 ;
  assign n3790 = ~n3788 & ~n3789 ;
  assign n3791 = n3784 & n3790 ;
  assign n3792 = ~n3784 & ~n3790 ;
  assign n3793 = ~n3791 & ~n3792 ;
  assign n3794 = n3778 & ~n3793 ;
  assign n3795 = ~n3778 & n3793 ;
  assign n3796 = ~n3794 & ~n3795 ;
  assign n3797 = ~n3697 & n3704 ;
  assign n3798 = ~n3696 & ~n3797 ;
  assign n3799 = ~n3796 & ~n3798 ;
  assign n3800 = n3796 & n3798 ;
  assign n3801 = ~n3799 & ~n3800 ;
  assign n3802 = \P1_P2_Address_reg[15]/NET0131  & ~n2791 ;
  assign n3803 = \P1_P3_Address_reg[15]/NET0131  & n2791 ;
  assign n3804 = ~n3802 & ~n3803 ;
  assign n3805 = ~\P4_wr_reg/NET0131  & ~n3804 ;
  assign n3806 = \P4_addr_reg[15]/NET0131  & \P4_wr_reg/NET0131  ;
  assign n3807 = ~n3805 & ~n3806 ;
  assign n3808 = n2845 & n3719 ;
  assign n3809 = n3717 & ~n3807 ;
  assign n3810 = n3718 & n3807 ;
  assign n3811 = ~n3809 & ~n3810 ;
  assign n3812 = ~n2834 & ~n3811 ;
  assign n3813 = ~n3808 & ~n3812 ;
  assign n3814 = ~n3807 & n3813 ;
  assign n3815 = ~n3720 & n3814 ;
  assign n3816 = n3720 & ~n3807 ;
  assign n3817 = ~n3813 & ~n3816 ;
  assign n3818 = ~n3814 & ~n3817 ;
  assign n3819 = ~n3815 & ~n3818 ;
  assign n3820 = n2908 & ~n2972 ;
  assign n3821 = n2906 & ~n2928 ;
  assign n3822 = ~n3820 & ~n3821 ;
  assign n3823 = n2879 & n3822 ;
  assign n3824 = ~n2879 & ~n3822 ;
  assign n3825 = ~n3823 & ~n3824 ;
  assign n3826 = n3819 & ~n3825 ;
  assign n3827 = ~n3819 & n3825 ;
  assign n3828 = ~n3826 & ~n3827 ;
  assign n3829 = n3801 & n3828 ;
  assign n3830 = ~n3801 & ~n3828 ;
  assign n3831 = ~n3829 & ~n3830 ;
  assign n3832 = n3772 & n3831 ;
  assign n3833 = ~n3772 & ~n3831 ;
  assign n3834 = ~n3832 & ~n3833 ;
  assign n3835 = ~n3666 & ~n3673 ;
  assign n3836 = ~n3674 & ~n3835 ;
  assign n3837 = ~n3747 & ~n3751 ;
  assign n3838 = ~n3748 & ~n3837 ;
  assign n3839 = ~n3836 & n3838 ;
  assign n3840 = n3836 & ~n3838 ;
  assign n3841 = ~n3839 & ~n3840 ;
  assign n3842 = ~n3727 & ~n3741 ;
  assign n3843 = ~n3728 & ~n3842 ;
  assign n3844 = n2950 & ~n3563 ;
  assign n3845 = n2954 & ~n3485 ;
  assign n3846 = ~n3844 & ~n3845 ;
  assign n3847 = n2944 & n3846 ;
  assign n3848 = ~n2944 & ~n3846 ;
  assign n3849 = ~n3847 & ~n3848 ;
  assign n3851 = \P2_P2_Address_reg[15]/NET0131  & ~n2828 ;
  assign n3852 = \P2_P3_Address_reg[15]/NET0131  & n2828 ;
  assign n3853 = ~n3851 & ~n3852 ;
  assign n3854 = ~n2826 & ~n3853 ;
  assign n3855 = \P2_P1_Address_reg[15]/NET0131  & n2826 ;
  assign n3856 = ~n3854 & ~n3855 ;
  assign n3857 = ~n2872 & ~n3856 ;
  assign n3859 = n2932 & ~n3857 ;
  assign n3850 = n2872 & ~n3736 ;
  assign n3858 = ~n2932 & n3857 ;
  assign n3860 = ~n3850 & ~n3858 ;
  assign n3861 = ~n3859 & n3860 ;
  assign n3862 = n3849 & n3861 ;
  assign n3863 = ~n3849 & ~n3861 ;
  assign n3864 = ~n3862 & ~n3863 ;
  assign n3865 = n3037 & n3510 ;
  assign n3866 = n2864 & n3622 ;
  assign n3867 = ~n3865 & ~n3866 ;
  assign n3868 = ~n3587 & ~n3867 ;
  assign n3869 = n3587 & n3867 ;
  assign n3870 = ~n3868 & ~n3869 ;
  assign n3871 = n3864 & n3870 ;
  assign n3872 = ~n3864 & ~n3870 ;
  assign n3873 = ~n3871 & ~n3872 ;
  assign n3874 = n3843 & ~n3873 ;
  assign n3875 = ~n3843 & n3873 ;
  assign n3876 = ~n3874 & ~n3875 ;
  assign n3877 = n3841 & n3876 ;
  assign n3878 = ~n3841 & ~n3876 ;
  assign n3879 = ~n3877 & ~n3878 ;
  assign n3880 = n3834 & n3879 ;
  assign n3881 = ~n3834 & ~n3879 ;
  assign n3882 = ~n3880 & ~n3881 ;
  assign n3883 = ~n3756 & ~n3759 ;
  assign n3884 = ~n3755 & ~n3883 ;
  assign n3885 = ~n3882 & n3884 ;
  assign n3886 = n3882 & ~n3884 ;
  assign n3887 = ~n3885 & ~n3886 ;
  assign n3888 = ~n3763 & n3767 ;
  assign n3889 = ~n3764 & ~n3888 ;
  assign n3890 = n3887 & ~n3889 ;
  assign n3891 = ~n3887 & n3889 ;
  assign n3892 = ~n3890 & ~n3891 ;
  assign n3893 = ~n3832 & ~n3879 ;
  assign n3894 = ~n3833 & ~n3893 ;
  assign n3895 = ~n3839 & ~n3876 ;
  assign n3896 = ~n3840 & ~n3895 ;
  assign n3897 = ~\P1_P2_Address_reg[16]/NET0131  & ~n2791 ;
  assign n3898 = ~\P1_P3_Address_reg[16]/NET0131  & n2791 ;
  assign n3899 = ~n3897 & ~n3898 ;
  assign n3900 = ~\P4_wr_reg/NET0131  & ~n3899 ;
  assign n3901 = ~\P4_addr_reg[16]/NET0131  & \P4_wr_reg/NET0131  ;
  assign n3902 = ~n3900 & ~n3901 ;
  assign n3903 = n3807 & ~n3902 ;
  assign n3904 = ~n3807 & n3902 ;
  assign n3905 = ~n3903 & ~n3904 ;
  assign n3906 = ~n2834 & n3905 ;
  assign n3908 = \P2_P2_Address_reg[16]/NET0131  & ~n2828 ;
  assign n3909 = \P2_P3_Address_reg[16]/NET0131  & n2828 ;
  assign n3910 = ~n3908 & ~n3909 ;
  assign n3911 = ~n2826 & ~n3910 ;
  assign n3912 = \P2_P1_Address_reg[16]/NET0131  & n2826 ;
  assign n3913 = ~n3911 & ~n3912 ;
  assign n3914 = ~n2872 & ~n3913 ;
  assign n3916 = n2932 & ~n3914 ;
  assign n3907 = n2872 & ~n3856 ;
  assign n3915 = ~n2932 & n3914 ;
  assign n3917 = ~n3907 & ~n3915 ;
  assign n3918 = ~n3916 & n3917 ;
  assign n3919 = n3906 & n3918 ;
  assign n3920 = ~n3906 & ~n3918 ;
  assign n3921 = ~n3919 & ~n3920 ;
  assign n3922 = n2888 & ~n2928 ;
  assign n3923 = ~n2921 & ~n3070 ;
  assign n3924 = ~n3922 & ~n3923 ;
  assign n3925 = n2986 & n3924 ;
  assign n3926 = ~n2986 & ~n3924 ;
  assign n3927 = ~n3925 & ~n3926 ;
  assign n3928 = ~n3921 & n3927 ;
  assign n3929 = n3921 & ~n3927 ;
  assign n3930 = ~n3928 & ~n3929 ;
  assign n3931 = n2950 & ~n3736 ;
  assign n3932 = n2954 & ~n3563 ;
  assign n3933 = ~n3931 & ~n3932 ;
  assign n3934 = n2944 & n3933 ;
  assign n3935 = ~n2944 & ~n3933 ;
  assign n3936 = ~n3934 & ~n3935 ;
  assign n3937 = n2908 & ~n3102 ;
  assign n3938 = n2906 & ~n2972 ;
  assign n3939 = ~n3937 & ~n3938 ;
  assign n3940 = n2879 & n3939 ;
  assign n3941 = ~n2879 & ~n3939 ;
  assign n3942 = ~n3940 & ~n3941 ;
  assign n3943 = n2864 & n3719 ;
  assign n3944 = n2845 & ~n3811 ;
  assign n3945 = ~n3943 & ~n3944 ;
  assign n3946 = n3807 & n3945 ;
  assign n3947 = ~n3807 & ~n3945 ;
  assign n3948 = ~n3946 & ~n3947 ;
  assign n3949 = n3942 & n3948 ;
  assign n3950 = ~n3942 & ~n3948 ;
  assign n3951 = ~n3949 & ~n3950 ;
  assign n3952 = n3936 & ~n3951 ;
  assign n3953 = ~n3936 & n3951 ;
  assign n3954 = ~n3952 & ~n3953 ;
  assign n3955 = ~n3930 & ~n3954 ;
  assign n3956 = n3930 & n3954 ;
  assign n3957 = ~n3955 & ~n3956 ;
  assign n3958 = n3027 & ~n3485 ;
  assign n3959 = ~n3031 & ~n3385 ;
  assign n3960 = ~n3958 & ~n3959 ;
  assign n3961 = n2901 & n3960 ;
  assign n3962 = ~n2901 & ~n3960 ;
  assign n3963 = ~n3961 & ~n3962 ;
  assign n3964 = n3006 & n3510 ;
  assign n3965 = n3037 & n3622 ;
  assign n3966 = ~n3964 & ~n3965 ;
  assign n3967 = n3587 & n3966 ;
  assign n3968 = ~n3587 & ~n3966 ;
  assign n3969 = ~n3967 & ~n3968 ;
  assign n3970 = ~n2960 & n3122 ;
  assign n3971 = ~n2999 & ~n3367 ;
  assign n3972 = ~n3970 & ~n3971 ;
  assign n3973 = n3363 & n3972 ;
  assign n3974 = ~n3363 & ~n3972 ;
  assign n3975 = ~n3973 & ~n3974 ;
  assign n3976 = n3969 & n3975 ;
  assign n3977 = ~n3969 & ~n3975 ;
  assign n3978 = ~n3976 & ~n3977 ;
  assign n3979 = n3963 & ~n3978 ;
  assign n3980 = ~n3963 & n3978 ;
  assign n3981 = ~n3979 & ~n3980 ;
  assign n3982 = ~n3957 & n3981 ;
  assign n3983 = n3957 & ~n3981 ;
  assign n3984 = ~n3982 & ~n3983 ;
  assign n3985 = ~n3896 & n3984 ;
  assign n3986 = n3896 & ~n3984 ;
  assign n3987 = ~n3985 & ~n3986 ;
  assign n3988 = ~n3843 & ~n3871 ;
  assign n3989 = ~n3872 & ~n3988 ;
  assign n3990 = ~n3800 & ~n3828 ;
  assign n3991 = ~n3799 & ~n3990 ;
  assign n3992 = ~n3989 & n3991 ;
  assign n3993 = n3989 & ~n3991 ;
  assign n3994 = ~n3992 & ~n3993 ;
  assign n3995 = ~n3818 & n3825 ;
  assign n3996 = ~n3815 & ~n3995 ;
  assign n3997 = n3778 & ~n3792 ;
  assign n3998 = ~n3791 & ~n3997 ;
  assign n3999 = ~n3862 & n3998 ;
  assign n4000 = n3862 & ~n3998 ;
  assign n4001 = ~n3999 & ~n4000 ;
  assign n4002 = n3996 & n4001 ;
  assign n4003 = ~n3996 & ~n4001 ;
  assign n4004 = ~n4002 & ~n4003 ;
  assign n4005 = n3994 & ~n4004 ;
  assign n4006 = ~n3994 & n4004 ;
  assign n4007 = ~n4005 & ~n4006 ;
  assign n4008 = n3987 & ~n4007 ;
  assign n4009 = ~n3987 & n4007 ;
  assign n4010 = ~n4008 & ~n4009 ;
  assign n4011 = ~n3894 & ~n4010 ;
  assign n4012 = n3894 & n4010 ;
  assign n4013 = ~n4011 & ~n4012 ;
  assign n4014 = ~n3885 & ~n3889 ;
  assign n4015 = ~n3886 & ~n4014 ;
  assign n4016 = n4013 & n4015 ;
  assign n4017 = ~n4013 & ~n4015 ;
  assign n4018 = ~n4016 & ~n4017 ;
  assign n4019 = ~n3986 & n4007 ;
  assign n4020 = ~n3985 & ~n4019 ;
  assign n4021 = \P1_P2_Address_reg[17]/NET0131  & ~n2791 ;
  assign n4022 = \P1_P3_Address_reg[17]/NET0131  & n2791 ;
  assign n4023 = ~n4021 & ~n4022 ;
  assign n4024 = ~\P4_wr_reg/NET0131  & ~n4023 ;
  assign n4025 = \P4_addr_reg[17]/NET0131  & \P4_wr_reg/NET0131  ;
  assign n4026 = ~n4024 & ~n4025 ;
  assign n4027 = ~n3906 & ~n4026 ;
  assign n4028 = n3027 & ~n3563 ;
  assign n4029 = ~n3031 & ~n3485 ;
  assign n4030 = ~n4028 & ~n4029 ;
  assign n4031 = n2901 & n4030 ;
  assign n4032 = ~n2901 & ~n4030 ;
  assign n4033 = ~n4031 & ~n4032 ;
  assign n4034 = n4027 & n4033 ;
  assign n4035 = ~n4027 & ~n4033 ;
  assign n4036 = ~n4034 & ~n4035 ;
  assign n4037 = n2888 & ~n2972 ;
  assign n4038 = ~n2928 & ~n3070 ;
  assign n4039 = ~n4037 & ~n4038 ;
  assign n4040 = n2986 & n4039 ;
  assign n4041 = ~n2986 & ~n4039 ;
  assign n4042 = ~n4040 & ~n4041 ;
  assign n4043 = ~n4036 & n4042 ;
  assign n4044 = n4036 & ~n4042 ;
  assign n4045 = ~n4043 & ~n4044 ;
  assign n4046 = n2908 & ~n3385 ;
  assign n4047 = n2906 & ~n3102 ;
  assign n4048 = ~n4046 & ~n4047 ;
  assign n4049 = n2879 & n4048 ;
  assign n4050 = ~n2879 & ~n4048 ;
  assign n4051 = ~n4049 & ~n4050 ;
  assign n4052 = n3037 & n3719 ;
  assign n4053 = n2864 & ~n3811 ;
  assign n4054 = ~n4052 & ~n4053 ;
  assign n4055 = n3807 & n4054 ;
  assign n4056 = ~n3807 & ~n4054 ;
  assign n4057 = ~n4055 & ~n4056 ;
  assign n4058 = n2845 & n3905 ;
  assign n4059 = n3807 & n4026 ;
  assign n4060 = ~n3807 & ~n4026 ;
  assign n4061 = ~n4059 & ~n4060 ;
  assign n4062 = ~n2834 & ~n3905 ;
  assign n4063 = n4061 & n4062 ;
  assign n4064 = ~n4058 & ~n4063 ;
  assign n4065 = n4026 & n4064 ;
  assign n4066 = ~n4026 & ~n4064 ;
  assign n4067 = ~n4065 & ~n4066 ;
  assign n4068 = n4057 & n4067 ;
  assign n4069 = ~n4057 & ~n4067 ;
  assign n4070 = ~n4068 & ~n4069 ;
  assign n4071 = n4051 & ~n4070 ;
  assign n4072 = ~n4051 & n4070 ;
  assign n4073 = ~n4071 & ~n4072 ;
  assign n4074 = n4045 & n4073 ;
  assign n4075 = ~n4045 & ~n4073 ;
  assign n4076 = ~n4074 & ~n4075 ;
  assign n4077 = n2950 & ~n3856 ;
  assign n4078 = n2954 & ~n3736 ;
  assign n4079 = ~n4077 & ~n4078 ;
  assign n4080 = n2944 & n4079 ;
  assign n4081 = ~n2944 & ~n4079 ;
  assign n4082 = ~n4080 & ~n4081 ;
  assign n4084 = \P2_P2_Address_reg[17]/NET0131  & ~n2828 ;
  assign n4085 = \P2_P3_Address_reg[17]/NET0131  & n2828 ;
  assign n4086 = ~n4084 & ~n4085 ;
  assign n4087 = ~n2826 & ~n4086 ;
  assign n4088 = \P2_P1_Address_reg[17]/NET0131  & n2826 ;
  assign n4089 = ~n4087 & ~n4088 ;
  assign n4090 = ~n2872 & ~n4089 ;
  assign n4092 = n2932 & ~n4090 ;
  assign n4083 = n2872 & ~n3913 ;
  assign n4091 = ~n2932 & n4090 ;
  assign n4093 = ~n4083 & ~n4091 ;
  assign n4094 = ~n4092 & n4093 ;
  assign n4095 = n4082 & n4094 ;
  assign n4096 = ~n4082 & ~n4094 ;
  assign n4097 = ~n4095 & ~n4096 ;
  assign n4098 = ~n2999 & n3510 ;
  assign n4099 = n3006 & n3622 ;
  assign n4100 = ~n4098 & ~n4099 ;
  assign n4101 = n3587 & n4100 ;
  assign n4102 = ~n3587 & ~n4100 ;
  assign n4103 = ~n4101 & ~n4102 ;
  assign n4104 = ~n2921 & n3122 ;
  assign n4105 = ~n2960 & ~n3367 ;
  assign n4106 = ~n4104 & ~n4105 ;
  assign n4107 = n3363 & n4106 ;
  assign n4108 = ~n3363 & ~n4106 ;
  assign n4109 = ~n4107 & ~n4108 ;
  assign n4110 = n4103 & n4109 ;
  assign n4111 = ~n4103 & ~n4109 ;
  assign n4112 = ~n4110 & ~n4111 ;
  assign n4113 = n4097 & n4112 ;
  assign n4114 = ~n4097 & ~n4112 ;
  assign n4115 = ~n4113 & ~n4114 ;
  assign n4116 = n4076 & ~n4115 ;
  assign n4117 = ~n4076 & n4115 ;
  assign n4118 = ~n4116 & ~n4117 ;
  assign n4119 = ~n3956 & ~n3981 ;
  assign n4120 = ~n3955 & ~n4119 ;
  assign n4121 = n3936 & ~n3950 ;
  assign n4122 = ~n3949 & ~n4121 ;
  assign n4123 = n3963 & ~n3977 ;
  assign n4124 = ~n3976 & ~n4123 ;
  assign n4125 = ~n4122 & ~n4124 ;
  assign n4126 = n4122 & n4124 ;
  assign n4127 = ~n4125 & ~n4126 ;
  assign n4128 = ~n3920 & n3927 ;
  assign n4129 = ~n3919 & ~n4128 ;
  assign n4130 = n4127 & ~n4129 ;
  assign n4131 = ~n4127 & n4129 ;
  assign n4132 = ~n4130 & ~n4131 ;
  assign n4133 = n4120 & ~n4132 ;
  assign n4134 = ~n4120 & n4132 ;
  assign n4135 = ~n4133 & ~n4134 ;
  assign n4136 = n3996 & ~n4000 ;
  assign n4137 = ~n3999 & ~n4136 ;
  assign n4138 = n4135 & n4137 ;
  assign n4139 = ~n4135 & ~n4137 ;
  assign n4140 = ~n4138 & ~n4139 ;
  assign n4141 = n4118 & ~n4140 ;
  assign n4142 = ~n4118 & n4140 ;
  assign n4143 = ~n4141 & ~n4142 ;
  assign n4144 = ~n3992 & ~n4004 ;
  assign n4145 = ~n3993 & ~n4144 ;
  assign n4146 = n4143 & ~n4145 ;
  assign n4147 = ~n4143 & n4145 ;
  assign n4148 = ~n4146 & ~n4147 ;
  assign n4149 = ~n4020 & n4148 ;
  assign n4150 = n4020 & ~n4148 ;
  assign n4151 = ~n4149 & ~n4150 ;
  assign n4152 = ~n4012 & n4015 ;
  assign n4153 = ~n4011 & ~n4152 ;
  assign n4154 = n4151 & n4153 ;
  assign n4155 = ~n4151 & ~n4153 ;
  assign n4156 = ~n4154 & ~n4155 ;
  assign n4157 = n2888 & ~n3102 ;
  assign n4158 = ~n2972 & ~n3070 ;
  assign n4159 = ~n4157 & ~n4158 ;
  assign n4160 = ~n2901 & n4159 ;
  assign n4161 = n2901 & ~n4159 ;
  assign n4162 = ~n4160 & ~n4161 ;
  assign n4163 = n2950 & ~n3913 ;
  assign n4164 = n2954 & ~n3856 ;
  assign n4165 = ~n4163 & ~n4164 ;
  assign n4166 = ~n4141 & ~n4145 ;
  assign n4167 = ~n4142 & ~n4166 ;
  assign n4168 = n4165 & ~n4167 ;
  assign n4169 = ~n4165 & n4167 ;
  assign n4170 = ~n4168 & ~n4169 ;
  assign n4171 = n4162 & ~n4170 ;
  assign n4172 = ~n4162 & n4170 ;
  assign n4173 = ~n4171 & ~n4172 ;
  assign n4174 = n2986 & n4173 ;
  assign n4175 = ~n2986 & ~n4173 ;
  assign n4176 = ~n4174 & ~n4175 ;
  assign n4177 = ~n4074 & n4115 ;
  assign n4178 = ~n4075 & ~n4177 ;
  assign n4179 = n4176 & ~n4178 ;
  assign n4180 = ~n4176 & n4178 ;
  assign n4181 = ~n4179 & ~n4180 ;
  assign n4182 = ~\P1_P2_Address_reg[18]/NET0131  & ~n2791 ;
  assign n4183 = ~\P1_P3_Address_reg[18]/NET0131  & n2791 ;
  assign n4184 = ~n4182 & ~n4183 ;
  assign n4185 = ~\P4_wr_reg/NET0131  & ~n4184 ;
  assign n4186 = ~\P4_addr_reg[18]/NET0131  & \P4_wr_reg/NET0131  ;
  assign n4187 = ~n4185 & ~n4186 ;
  assign n4188 = ~n4026 & ~n4187 ;
  assign n4189 = n4026 & n4187 ;
  assign n4190 = ~n4188 & ~n4189 ;
  assign n4191 = ~n2834 & ~n4190 ;
  assign n4194 = ~\P2_P2_Address_reg[18]/NET0131  & ~n2828 ;
  assign n4195 = ~\P2_P3_Address_reg[18]/NET0131  & n2828 ;
  assign n4196 = ~n4194 & ~n4195 ;
  assign n4197 = ~n2826 & ~n4196 ;
  assign n4193 = ~\P2_P1_Address_reg[18]/NET0131  & n2826 ;
  assign n4198 = ~n2872 & ~n4193 ;
  assign n4199 = ~n4197 & n4198 ;
  assign n4192 = n2872 & ~n4089 ;
  assign n4200 = ~n2932 & ~n4192 ;
  assign n4201 = ~n4199 & n4200 ;
  assign n4202 = n2932 & n4199 ;
  assign n4203 = ~n4201 & ~n4202 ;
  assign n4204 = n4191 & ~n4203 ;
  assign n4205 = ~n4191 & n4203 ;
  assign n4206 = ~n4204 & ~n4205 ;
  assign n4207 = n3027 & ~n3736 ;
  assign n4208 = ~n3031 & ~n3563 ;
  assign n4209 = ~n4207 & ~n4208 ;
  assign n4210 = ~n2944 & n4209 ;
  assign n4211 = n2944 & ~n4209 ;
  assign n4212 = ~n4210 & ~n4211 ;
  assign n4213 = ~n4134 & ~n4137 ;
  assign n4214 = ~n4133 & ~n4213 ;
  assign n4215 = n4212 & ~n4214 ;
  assign n4216 = ~n4212 & n4214 ;
  assign n4217 = ~n4215 & ~n4216 ;
  assign n4218 = n4206 & ~n4217 ;
  assign n4219 = ~n4206 & n4217 ;
  assign n4220 = ~n4218 & ~n4219 ;
  assign n4221 = n4181 & ~n4220 ;
  assign n4222 = ~n4181 & n4220 ;
  assign n4223 = ~n4221 & ~n4222 ;
  assign n4224 = ~n4011 & ~n4149 ;
  assign n4225 = ~n4152 & n4224 ;
  assign n4226 = ~n4150 & ~n4225 ;
  assign n4227 = ~n4035 & n4042 ;
  assign n4228 = ~n4034 & ~n4227 ;
  assign n4229 = ~n2960 & n3510 ;
  assign n4230 = ~n2999 & n3622 ;
  assign n4231 = ~n4229 & ~n4230 ;
  assign n4232 = n4051 & ~n4069 ;
  assign n4233 = ~n4068 & ~n4232 ;
  assign n4234 = n4231 & ~n4233 ;
  assign n4235 = ~n4231 & n4233 ;
  assign n4236 = ~n4234 & ~n4235 ;
  assign n4237 = n4228 & n4236 ;
  assign n4238 = ~n4228 & ~n4236 ;
  assign n4239 = ~n4237 & ~n4238 ;
  assign n4240 = n4095 & ~n4110 ;
  assign n4241 = ~n4095 & n4110 ;
  assign n4242 = ~n4240 & ~n4241 ;
  assign n4243 = ~n4113 & n4242 ;
  assign n4244 = n4239 & ~n4243 ;
  assign n4245 = ~n4239 & n4243 ;
  assign n4246 = ~n4244 & ~n4245 ;
  assign n4247 = ~n4126 & ~n4129 ;
  assign n4248 = ~n4125 & ~n4247 ;
  assign n4249 = n3621 & ~n4248 ;
  assign n4250 = ~n3621 & n4248 ;
  assign n4251 = ~n4249 & ~n4250 ;
  assign n4253 = n2845 & ~n3905 ;
  assign n4252 = n2864 & n3905 ;
  assign n4254 = n4061 & ~n4252 ;
  assign n4255 = ~n4253 & n4254 ;
  assign n4256 = ~n4061 & n4252 ;
  assign n4257 = ~n4255 & ~n4256 ;
  assign n4258 = ~n2928 & n3122 ;
  assign n4259 = ~n2921 & ~n3367 ;
  assign n4260 = ~n4258 & ~n4259 ;
  assign n4261 = n3006 & n3719 ;
  assign n4262 = n3037 & ~n3811 ;
  assign n4263 = ~n4261 & ~n4262 ;
  assign n4264 = n4260 & ~n4263 ;
  assign n4265 = ~n4260 & n4263 ;
  assign n4266 = ~n4264 & ~n4265 ;
  assign n4267 = n4257 & ~n4266 ;
  assign n4268 = ~n4257 & n4266 ;
  assign n4269 = ~n4267 & ~n4268 ;
  assign n4270 = n4251 & n4269 ;
  assign n4271 = ~n4251 & ~n4269 ;
  assign n4272 = ~n4270 & ~n4271 ;
  assign n4273 = n2908 & ~n3485 ;
  assign n4274 = n2906 & ~n3385 ;
  assign n4275 = ~n4273 & ~n4274 ;
  assign n4276 = ~n2879 & n4275 ;
  assign n4277 = n2879 & ~n4275 ;
  assign n4278 = ~n4276 & ~n4277 ;
  assign n4279 = n4272 & ~n4278 ;
  assign n4280 = ~n4272 & n4278 ;
  assign n4281 = ~n4279 & ~n4280 ;
  assign n4282 = n4246 & n4281 ;
  assign n4283 = ~n4246 & ~n4281 ;
  assign n4284 = ~n4282 & ~n4283 ;
  assign n4285 = n4226 & ~n4284 ;
  assign n4286 = ~n4226 & n4284 ;
  assign n4287 = ~n4285 & ~n4286 ;
  assign n4288 = n4223 & n4287 ;
  assign n4289 = ~n4223 & ~n4287 ;
  assign n4290 = ~n4288 & ~n4289 ;
  assign n4291 = ~n2834 & ~n2932 ;
  assign n4292 = n3328 & ~n4291 ;
  assign n4293 = ~n3328 & n4291 ;
  assign n4294 = ~n4292 & ~n4293 ;
  assign n4295 = n3331 & ~n3337 ;
  assign n4296 = ~n3338 & ~n4295 ;
  assign n4297 = ~n3326 & ~n3327 ;
  assign n4298 = n3338 & ~n4297 ;
  assign n4299 = ~n3338 & n4297 ;
  assign n4300 = ~n4298 & ~n4299 ;
  assign n4301 = ~n3316 & ~n3317 ;
  assign n4302 = ~n3340 & n4301 ;
  assign n4303 = n3340 & ~n4301 ;
  assign n4304 = ~n4302 & ~n4303 ;
  assign n4305 = ~n3301 & ~n3302 ;
  assign n4306 = ~n3342 & n4305 ;
  assign n4307 = n3342 & ~n4305 ;
  assign n4308 = ~n4306 & ~n4307 ;
  assign n4309 = ~n3279 & ~n3280 ;
  assign n4310 = ~n3344 & n4309 ;
  assign n4311 = n3344 & ~n4309 ;
  assign n4312 = ~n4310 & ~n4311 ;
  assign n4313 = ~n3260 & ~n3261 ;
  assign n4314 = ~n3346 & n4313 ;
  assign n4315 = n3346 & ~n4313 ;
  assign n4316 = ~n4314 & ~n4315 ;
  assign n4317 = ~n3227 & ~n3228 ;
  assign n4318 = ~n3348 & n4317 ;
  assign n4319 = n3348 & ~n4317 ;
  assign n4320 = ~n4318 & ~n4319 ;
  assign n4321 = ~n3195 & ~n3196 ;
  assign n4322 = ~n3350 & n4321 ;
  assign n4323 = n3350 & ~n4321 ;
  assign n4324 = ~n4322 & ~n4323 ;
  assign n4325 = \P1_P1_InstQueueWr_Addr_reg[0]/NET0131  & ~\P1_P1_InstQueueWr_Addr_reg[1]/NET0131  ;
  assign n4326 = ~\P1_P1_InstQueueWr_Addr_reg[2]/NET0131  & n4325 ;
  assign n4327 = \P1_P1_InstQueueWr_Addr_reg[3]/NET0131  & n4326 ;
  assign n4328 = \din[3]_pad  & sel_pad ;
  assign n4329 = \din[1]_pad  & sel_pad ;
  assign n4330 = \din[2]_pad  & n4329 ;
  assign n4331 = ~n4328 & ~n4330 ;
  assign n4332 = ~\din[1]_pad  & ~\din[2]_pad  ;
  assign n4333 = sel_pad & ~n4332 ;
  assign n4334 = \din[3]_pad  & n4333 ;
  assign n4335 = ~n4331 & ~n4334 ;
  assign n4336 = \P4_datao_reg[20]/NET0131  & n4335 ;
  assign n4337 = ~n4330 & n4333 ;
  assign n4338 = \P4_datao_reg[21]/NET0131  & n4337 ;
  assign n4339 = ~n4336 & ~n4338 ;
  assign n4340 = ~n4328 & n4339 ;
  assign n4341 = n4328 & ~n4339 ;
  assign n4342 = ~n4340 & ~n4341 ;
  assign n4343 = \din[0]_pad  & sel_pad ;
  assign n4344 = \P4_datao_reg[23]/NET0131  & n4343 ;
  assign n4345 = ~\din[1]_pad  & n4344 ;
  assign n4346 = \P4_datao_reg[22]/NET0131  & ~n4343 ;
  assign n4347 = n4329 & ~n4344 ;
  assign n4348 = ~n4346 & n4347 ;
  assign n4349 = ~n4345 & ~n4348 ;
  assign n4350 = n4342 & ~n4349 ;
  assign n4351 = \din[13]_pad  & sel_pad ;
  assign n4352 = \din[11]_pad  & sel_pad ;
  assign n4353 = \din[12]_pad  & n4352 ;
  assign n4354 = ~\din[11]_pad  & ~\din[12]_pad  ;
  assign n4355 = sel_pad & ~n4354 ;
  assign n4356 = ~n4353 & n4355 ;
  assign n4357 = \P4_datao_reg[12]/NET0131  & n4356 ;
  assign n4358 = ~n4351 & ~n4353 ;
  assign n4359 = \din[13]_pad  & n4355 ;
  assign n4360 = ~n4358 & ~n4359 ;
  assign n4361 = \P4_datao_reg[11]/NET0131  & n4360 ;
  assign n4362 = ~n4357 & ~n4361 ;
  assign n4363 = n4351 & ~n4362 ;
  assign n4364 = ~n4351 & n4362 ;
  assign n4365 = ~n4363 & ~n4364 ;
  assign n4366 = ~n4350 & ~n4365 ;
  assign n4367 = n4350 & n4365 ;
  assign n4368 = \din[15]_pad  & sel_pad ;
  assign n4369 = \din[14]_pad  & n4351 ;
  assign n4370 = ~n4368 & ~n4369 ;
  assign n4371 = ~\din[13]_pad  & ~\din[14]_pad  ;
  assign n4372 = sel_pad & ~n4371 ;
  assign n4373 = \din[15]_pad  & n4372 ;
  assign n4374 = ~n4370 & ~n4373 ;
  assign n4375 = \P4_datao_reg[8]/NET0131  & n4374 ;
  assign n4376 = ~n4369 & n4372 ;
  assign n4377 = \P4_datao_reg[9]/NET0131  & n4376 ;
  assign n4378 = ~n4375 & ~n4377 ;
  assign n4379 = ~n4368 & n4378 ;
  assign n4380 = n4368 & ~n4378 ;
  assign n4381 = ~n4379 & ~n4380 ;
  assign n4382 = \din[17]_pad  & sel_pad ;
  assign n4383 = \din[16]_pad  & n4368 ;
  assign n4384 = ~n4382 & ~n4383 ;
  assign n4385 = ~\din[15]_pad  & ~\din[16]_pad  ;
  assign n4386 = sel_pad & ~n4385 ;
  assign n4387 = \din[17]_pad  & n4386 ;
  assign n4388 = ~n4384 & ~n4387 ;
  assign n4389 = \P4_datao_reg[6]/NET0131  & n4388 ;
  assign n4390 = ~n4383 & n4386 ;
  assign n4391 = \P4_datao_reg[7]/NET0131  & n4390 ;
  assign n4392 = ~n4389 & ~n4391 ;
  assign n4393 = n4382 & ~n4392 ;
  assign n4394 = ~n4382 & n4392 ;
  assign n4395 = ~n4393 & ~n4394 ;
  assign n4396 = ~n4381 & ~n4395 ;
  assign n4397 = n4381 & n4395 ;
  assign n4398 = \din[7]_pad  & sel_pad ;
  assign n4399 = \din[5]_pad  & sel_pad ;
  assign n4400 = \din[6]_pad  & n4399 ;
  assign n4401 = ~n4398 & ~n4400 ;
  assign n4402 = ~\din[5]_pad  & ~\din[6]_pad  ;
  assign n4403 = sel_pad & ~n4402 ;
  assign n4404 = \din[7]_pad  & n4403 ;
  assign n4405 = ~n4401 & ~n4404 ;
  assign n4406 = \P4_datao_reg[16]/NET0131  & n4405 ;
  assign n4407 = ~n4400 & n4403 ;
  assign n4408 = \P4_datao_reg[17]/NET0131  & n4407 ;
  assign n4409 = ~n4406 & ~n4408 ;
  assign n4410 = ~n4398 & n4409 ;
  assign n4411 = n4398 & ~n4409 ;
  assign n4412 = ~n4410 & ~n4411 ;
  assign n4413 = ~n4397 & ~n4412 ;
  assign n4414 = ~n4396 & ~n4413 ;
  assign n4415 = ~n4367 & ~n4414 ;
  assign n4416 = ~n4366 & ~n4415 ;
  assign n4417 = \din[23]_pad  & sel_pad ;
  assign n4418 = \din[24]_pad  & n4417 ;
  assign n4419 = ~\din[23]_pad  & ~\din[24]_pad  ;
  assign n4420 = sel_pad & ~n4419 ;
  assign n4421 = ~n4418 & n4420 ;
  assign n4422 = \P4_datao_reg[0]/NET0131  & n4421 ;
  assign n4423 = \P4_datao_reg[24]/NET0131  & n4343 ;
  assign n4424 = ~\din[1]_pad  & n4423 ;
  assign n4425 = \P4_datao_reg[23]/NET0131  & ~n4343 ;
  assign n4426 = n4329 & ~n4423 ;
  assign n4427 = ~n4425 & n4426 ;
  assign n4428 = ~n4424 & ~n4427 ;
  assign n4429 = n4422 & ~n4428 ;
  assign n4430 = ~n4422 & n4428 ;
  assign n4431 = \din[9]_pad  & sel_pad ;
  assign n4432 = \din[10]_pad  & n4431 ;
  assign n4433 = ~\din[10]_pad  & ~\din[9]_pad  ;
  assign n4434 = sel_pad & ~n4433 ;
  assign n4435 = ~n4432 & n4434 ;
  assign n4436 = \P4_datao_reg[14]/NET0131  & n4435 ;
  assign n4437 = ~n4352 & ~n4432 ;
  assign n4438 = \din[11]_pad  & n4434 ;
  assign n4439 = ~n4437 & ~n4438 ;
  assign n4440 = \P4_datao_reg[13]/NET0131  & n4439 ;
  assign n4441 = ~n4436 & ~n4440 ;
  assign n4442 = n4352 & ~n4441 ;
  assign n4443 = ~n4352 & n4441 ;
  assign n4444 = ~n4442 & ~n4443 ;
  assign n4445 = ~n4430 & n4444 ;
  assign n4446 = ~n4429 & ~n4445 ;
  assign n4447 = \din[25]_pad  & sel_pad ;
  assign n4448 = ~n4422 & n4447 ;
  assign n4449 = \P4_datao_reg[12]/NET0131  & n4360 ;
  assign n4450 = \P4_datao_reg[13]/NET0131  & n4356 ;
  assign n4451 = ~n4449 & ~n4450 ;
  assign n4452 = n4351 & ~n4451 ;
  assign n4453 = ~n4351 & n4451 ;
  assign n4454 = ~n4452 & ~n4453 ;
  assign n4455 = n4448 & n4454 ;
  assign n4456 = ~n4448 & ~n4454 ;
  assign n4457 = ~n4455 & ~n4456 ;
  assign n4458 = ~n4418 & ~n4447 ;
  assign n4459 = \din[25]_pad  & n4420 ;
  assign n4460 = ~n4458 & ~n4459 ;
  assign n4461 = \P4_datao_reg[0]/NET0131  & n4460 ;
  assign n4462 = \P4_datao_reg[1]/NET0131  & n4421 ;
  assign n4463 = ~n4461 & ~n4462 ;
  assign n4464 = n4447 & ~n4463 ;
  assign n4465 = ~n4447 & n4463 ;
  assign n4466 = ~n4464 & ~n4465 ;
  assign n4467 = n4457 & ~n4466 ;
  assign n4468 = ~n4457 & n4466 ;
  assign n4469 = ~n4467 & ~n4468 ;
  assign n4470 = ~n4446 & ~n4469 ;
  assign n4471 = n4446 & n4469 ;
  assign n4472 = ~n4470 & ~n4471 ;
  assign n4473 = \P4_datao_reg[17]/NET0131  & n4405 ;
  assign n4474 = \P4_datao_reg[18]/NET0131  & n4407 ;
  assign n4475 = ~n4473 & ~n4474 ;
  assign n4476 = ~n4398 & n4475 ;
  assign n4477 = n4398 & ~n4475 ;
  assign n4478 = ~n4476 & ~n4477 ;
  assign n4479 = \P4_datao_reg[9]/NET0131  & n4374 ;
  assign n4480 = \P4_datao_reg[10]/NET0131  & n4376 ;
  assign n4481 = ~n4479 & ~n4480 ;
  assign n4482 = ~n4368 & n4481 ;
  assign n4483 = n4368 & ~n4481 ;
  assign n4484 = ~n4482 & ~n4483 ;
  assign n4485 = n4478 & n4484 ;
  assign n4486 = ~n4478 & ~n4484 ;
  assign n4487 = \P4_datao_reg[22]/NET0131  & n4337 ;
  assign n4488 = \P4_datao_reg[21]/NET0131  & n4335 ;
  assign n4489 = ~n4487 & ~n4488 ;
  assign n4490 = n4328 & ~n4489 ;
  assign n4491 = ~n4328 & n4489 ;
  assign n4492 = ~n4490 & ~n4491 ;
  assign n4493 = ~n4486 & n4492 ;
  assign n4494 = ~n4485 & ~n4493 ;
  assign n4495 = n4472 & ~n4494 ;
  assign n4496 = ~n4472 & n4494 ;
  assign n4497 = ~n4495 & ~n4496 ;
  assign n4498 = ~n4416 & ~n4497 ;
  assign n4499 = n4416 & n4497 ;
  assign n4500 = ~n4485 & ~n4486 ;
  assign n4501 = ~n4492 & n4500 ;
  assign n4502 = n4492 & ~n4500 ;
  assign n4503 = ~n4501 & ~n4502 ;
  assign n4504 = \din[8]_pad  & n4398 ;
  assign n4505 = ~\din[7]_pad  & ~\din[8]_pad  ;
  assign n4506 = sel_pad & ~n4505 ;
  assign n4507 = ~n4504 & n4506 ;
  assign n4508 = \P4_datao_reg[16]/NET0131  & n4507 ;
  assign n4509 = ~n4431 & ~n4504 ;
  assign n4510 = \din[9]_pad  & n4506 ;
  assign n4511 = ~n4509 & ~n4510 ;
  assign n4512 = \P4_datao_reg[15]/NET0131  & n4511 ;
  assign n4513 = ~n4508 & ~n4512 ;
  assign n4514 = n4431 & ~n4513 ;
  assign n4515 = ~n4431 & n4513 ;
  assign n4516 = ~n4514 & ~n4515 ;
  assign n4517 = \din[19]_pad  & sel_pad ;
  assign n4518 = \din[18]_pad  & n4382 ;
  assign n4519 = ~n4517 & ~n4518 ;
  assign n4520 = ~\din[17]_pad  & ~\din[18]_pad  ;
  assign n4521 = sel_pad & ~n4520 ;
  assign n4522 = \din[19]_pad  & n4521 ;
  assign n4523 = ~n4519 & ~n4522 ;
  assign n4524 = \P4_datao_reg[5]/NET0131  & n4523 ;
  assign n4525 = ~n4518 & n4521 ;
  assign n4526 = \P4_datao_reg[6]/NET0131  & n4525 ;
  assign n4527 = ~n4524 & ~n4526 ;
  assign n4528 = n4517 & ~n4527 ;
  assign n4529 = ~n4517 & n4527 ;
  assign n4530 = ~n4528 & ~n4529 ;
  assign n4531 = \P4_datao_reg[8]/NET0131  & n4390 ;
  assign n4532 = \P4_datao_reg[7]/NET0131  & n4388 ;
  assign n4533 = ~n4531 & ~n4532 ;
  assign n4534 = n4382 & ~n4533 ;
  assign n4535 = ~n4382 & n4533 ;
  assign n4536 = ~n4534 & ~n4535 ;
  assign n4537 = ~n4530 & ~n4536 ;
  assign n4538 = n4530 & n4536 ;
  assign n4539 = ~n4537 & ~n4538 ;
  assign n4540 = n4516 & n4539 ;
  assign n4541 = ~n4516 & ~n4539 ;
  assign n4542 = ~n4540 & ~n4541 ;
  assign n4543 = n4503 & ~n4542 ;
  assign n4544 = ~n4503 & n4542 ;
  assign n4545 = \din[4]_pad  & n4328 ;
  assign n4546 = ~\din[3]_pad  & ~\din[4]_pad  ;
  assign n4547 = sel_pad & ~n4546 ;
  assign n4548 = ~n4545 & n4547 ;
  assign n4549 = \P4_datao_reg[20]/NET0131  & n4548 ;
  assign n4550 = ~n4399 & ~n4545 ;
  assign n4551 = \din[5]_pad  & n4547 ;
  assign n4552 = ~n4550 & ~n4551 ;
  assign n4553 = \P4_datao_reg[19]/NET0131  & n4552 ;
  assign n4554 = ~n4549 & ~n4553 ;
  assign n4555 = n4399 & ~n4554 ;
  assign n4556 = ~n4399 & n4554 ;
  assign n4557 = ~n4555 & ~n4556 ;
  assign n4558 = \din[21]_pad  & sel_pad ;
  assign n4559 = \din[22]_pad  & n4558 ;
  assign n4560 = ~\din[21]_pad  & ~\din[22]_pad  ;
  assign n4561 = sel_pad & ~n4560 ;
  assign n4562 = ~n4559 & n4561 ;
  assign n4563 = \P4_datao_reg[2]/NET0131  & n4562 ;
  assign n4564 = ~n4417 & ~n4559 ;
  assign n4565 = \din[23]_pad  & n4561 ;
  assign n4566 = ~n4564 & ~n4565 ;
  assign n4567 = \P4_datao_reg[1]/NET0131  & n4566 ;
  assign n4568 = ~n4563 & ~n4567 ;
  assign n4569 = n4417 & ~n4568 ;
  assign n4570 = ~n4417 & n4568 ;
  assign n4571 = ~n4569 & ~n4570 ;
  assign n4572 = \din[19]_pad  & ~\din[20]_pad  ;
  assign n4573 = ~\din[19]_pad  & \din[20]_pad  ;
  assign n4574 = ~n4572 & ~n4573 ;
  assign n4575 = sel_pad & ~n4574 ;
  assign n4576 = \P4_datao_reg[4]/NET0131  & n4575 ;
  assign n4577 = n4517 & ~n4558 ;
  assign n4578 = ~n4517 & n4558 ;
  assign n4579 = ~n4577 & ~n4578 ;
  assign n4580 = ~n4575 & ~n4579 ;
  assign n4581 = \P4_datao_reg[3]/NET0131  & n4580 ;
  assign n4582 = ~n4576 & ~n4581 ;
  assign n4583 = n4558 & ~n4582 ;
  assign n4584 = ~n4558 & n4582 ;
  assign n4585 = ~n4583 & ~n4584 ;
  assign n4586 = ~n4571 & ~n4585 ;
  assign n4587 = n4571 & n4585 ;
  assign n4588 = ~n4586 & ~n4587 ;
  assign n4589 = n4557 & n4588 ;
  assign n4590 = ~n4557 & ~n4588 ;
  assign n4591 = ~n4589 & ~n4590 ;
  assign n4592 = ~n4544 & ~n4591 ;
  assign n4593 = ~n4543 & ~n4592 ;
  assign n4594 = ~n4499 & ~n4593 ;
  assign n4595 = ~n4498 & ~n4594 ;
  assign n4596 = ~n4471 & ~n4494 ;
  assign n4597 = ~n4470 & ~n4596 ;
  assign n4598 = ~n4557 & ~n4587 ;
  assign n4599 = ~n4586 & ~n4598 ;
  assign n4600 = ~n4516 & ~n4538 ;
  assign n4601 = ~n4537 & ~n4600 ;
  assign n4602 = ~n4599 & ~n4601 ;
  assign n4603 = n4599 & n4601 ;
  assign n4604 = \P4_datao_reg[22]/NET0131  & n4335 ;
  assign n4605 = \P4_datao_reg[23]/NET0131  & n4337 ;
  assign n4606 = ~n4604 & ~n4605 ;
  assign n4607 = ~n4328 & n4606 ;
  assign n4608 = n4328 & ~n4606 ;
  assign n4609 = ~n4607 & ~n4608 ;
  assign n4610 = \P4_datao_reg[25]/NET0131  & n4343 ;
  assign n4611 = ~\din[1]_pad  & n4610 ;
  assign n4612 = \P4_datao_reg[24]/NET0131  & ~n4343 ;
  assign n4613 = n4329 & ~n4610 ;
  assign n4614 = ~n4612 & n4613 ;
  assign n4615 = ~n4611 & ~n4614 ;
  assign n4616 = n4609 & ~n4615 ;
  assign n4617 = ~n4609 & n4615 ;
  assign n4618 = ~n4616 & ~n4617 ;
  assign n4619 = ~n4603 & ~n4618 ;
  assign n4620 = ~n4602 & ~n4619 ;
  assign n4621 = n4597 & ~n4620 ;
  assign n4622 = ~n4597 & n4620 ;
  assign n4623 = ~n4621 & ~n4622 ;
  assign n4624 = \P4_datao_reg[16]/NET0131  & n4511 ;
  assign n4625 = \P4_datao_reg[17]/NET0131  & n4507 ;
  assign n4626 = ~n4624 & ~n4625 ;
  assign n4627 = ~n4431 & n4626 ;
  assign n4628 = n4431 & ~n4626 ;
  assign n4629 = ~n4627 & ~n4628 ;
  assign n4630 = \P4_datao_reg[5]/NET0131  & n4575 ;
  assign n4631 = \P4_datao_reg[4]/NET0131  & n4580 ;
  assign n4632 = ~n4630 & ~n4631 ;
  assign n4633 = n4558 & ~n4632 ;
  assign n4634 = ~n4558 & n4632 ;
  assign n4635 = ~n4633 & ~n4634 ;
  assign n4636 = \P4_datao_reg[7]/NET0131  & n4525 ;
  assign n4637 = \P4_datao_reg[6]/NET0131  & n4523 ;
  assign n4638 = ~n4636 & ~n4637 ;
  assign n4639 = n4517 & ~n4638 ;
  assign n4640 = ~n4517 & n4638 ;
  assign n4641 = ~n4639 & ~n4640 ;
  assign n4642 = ~n4635 & ~n4641 ;
  assign n4643 = n4635 & n4641 ;
  assign n4644 = ~n4642 & ~n4643 ;
  assign n4645 = n4629 & n4644 ;
  assign n4646 = ~n4629 & ~n4644 ;
  assign n4647 = ~n4645 & ~n4646 ;
  assign n4648 = \P4_datao_reg[20]/NET0131  & n4552 ;
  assign n4649 = \P4_datao_reg[21]/NET0131  & n4548 ;
  assign n4650 = ~n4648 & ~n4649 ;
  assign n4651 = ~n4399 & n4650 ;
  assign n4652 = n4399 & ~n4650 ;
  assign n4653 = ~n4651 & ~n4652 ;
  assign n4654 = \P4_datao_reg[14]/NET0131  & n4439 ;
  assign n4655 = \P4_datao_reg[15]/NET0131  & n4435 ;
  assign n4656 = ~n4654 & ~n4655 ;
  assign n4657 = ~n4352 & n4656 ;
  assign n4658 = n4352 & ~n4656 ;
  assign n4659 = ~n4657 & ~n4658 ;
  assign n4660 = \P4_datao_reg[2]/NET0131  & n4566 ;
  assign n4661 = \P4_datao_reg[3]/NET0131  & n4562 ;
  assign n4662 = ~n4660 & ~n4661 ;
  assign n4663 = ~n4417 & n4662 ;
  assign n4664 = n4417 & ~n4662 ;
  assign n4665 = ~n4663 & ~n4664 ;
  assign n4666 = ~n4659 & ~n4665 ;
  assign n4667 = n4659 & n4665 ;
  assign n4668 = ~n4666 & ~n4667 ;
  assign n4669 = n4653 & n4668 ;
  assign n4670 = ~n4653 & ~n4668 ;
  assign n4671 = ~n4669 & ~n4670 ;
  assign n4672 = n4647 & n4671 ;
  assign n4673 = ~n4647 & ~n4671 ;
  assign n4674 = \P4_datao_reg[18]/NET0131  & n4405 ;
  assign n4675 = \P4_datao_reg[19]/NET0131  & n4407 ;
  assign n4676 = ~n4674 & ~n4675 ;
  assign n4677 = ~n4398 & n4676 ;
  assign n4678 = n4398 & ~n4676 ;
  assign n4679 = ~n4677 & ~n4678 ;
  assign n4680 = \P4_datao_reg[10]/NET0131  & n4374 ;
  assign n4681 = \P4_datao_reg[11]/NET0131  & n4376 ;
  assign n4682 = ~n4680 & ~n4681 ;
  assign n4683 = n4368 & ~n4682 ;
  assign n4684 = ~n4368 & n4682 ;
  assign n4685 = ~n4683 & ~n4684 ;
  assign n4686 = \P4_datao_reg[9]/NET0131  & n4390 ;
  assign n4687 = \P4_datao_reg[8]/NET0131  & n4388 ;
  assign n4688 = ~n4686 & ~n4687 ;
  assign n4689 = n4382 & ~n4688 ;
  assign n4690 = ~n4382 & n4688 ;
  assign n4691 = ~n4689 & ~n4690 ;
  assign n4692 = n4685 & n4691 ;
  assign n4693 = ~n4685 & ~n4691 ;
  assign n4694 = ~n4692 & ~n4693 ;
  assign n4695 = n4679 & ~n4694 ;
  assign n4696 = ~n4679 & n4694 ;
  assign n4697 = ~n4695 & ~n4696 ;
  assign n4698 = ~n4673 & ~n4697 ;
  assign n4699 = ~n4672 & ~n4698 ;
  assign n4700 = n4623 & ~n4699 ;
  assign n4701 = ~n4623 & n4699 ;
  assign n4702 = ~n4700 & ~n4701 ;
  assign n4703 = n4595 & n4702 ;
  assign n4704 = ~n4595 & ~n4702 ;
  assign n4705 = \P4_datao_reg[12]/NET0131  & n4439 ;
  assign n4706 = \P4_datao_reg[13]/NET0131  & n4435 ;
  assign n4707 = ~n4705 & ~n4706 ;
  assign n4708 = n4352 & ~n4707 ;
  assign n4709 = ~n4352 & n4707 ;
  assign n4710 = ~n4708 & ~n4709 ;
  assign n4711 = \P4_datao_reg[1]/NET0131  & n4562 ;
  assign n4712 = \P4_datao_reg[0]/NET0131  & n4566 ;
  assign n4713 = ~n4711 & ~n4712 ;
  assign n4714 = n4417 & ~n4713 ;
  assign n4715 = ~n4417 & n4713 ;
  assign n4716 = ~n4714 & ~n4715 ;
  assign n4717 = ~n4710 & ~n4716 ;
  assign n4718 = n4710 & n4716 ;
  assign n4719 = \P4_datao_reg[18]/NET0131  & n4552 ;
  assign n4720 = \P4_datao_reg[19]/NET0131  & n4548 ;
  assign n4721 = ~n4719 & ~n4720 ;
  assign n4722 = ~n4399 & n4721 ;
  assign n4723 = n4399 & ~n4721 ;
  assign n4724 = ~n4722 & ~n4723 ;
  assign n4725 = ~n4718 & ~n4724 ;
  assign n4726 = ~n4717 & ~n4725 ;
  assign n4727 = ~n4429 & ~n4430 ;
  assign n4728 = n4444 & n4727 ;
  assign n4729 = ~n4444 & ~n4727 ;
  assign n4730 = ~n4728 & ~n4729 ;
  assign n4731 = ~n4726 & ~n4730 ;
  assign n4732 = n4726 & n4730 ;
  assign n4733 = \P4_datao_reg[4]/NET0131  & n4523 ;
  assign n4734 = \P4_datao_reg[5]/NET0131  & n4525 ;
  assign n4735 = ~n4733 & ~n4734 ;
  assign n4736 = ~n4517 & n4735 ;
  assign n4737 = n4517 & ~n4735 ;
  assign n4738 = ~n4736 & ~n4737 ;
  assign n4739 = \P4_datao_reg[3]/NET0131  & n4575 ;
  assign n4740 = \P4_datao_reg[2]/NET0131  & n4580 ;
  assign n4741 = ~n4739 & ~n4740 ;
  assign n4742 = n4558 & ~n4741 ;
  assign n4743 = ~n4558 & n4741 ;
  assign n4744 = ~n4742 & ~n4743 ;
  assign n4745 = ~n4738 & ~n4744 ;
  assign n4746 = n4738 & n4744 ;
  assign n4747 = \P4_datao_reg[14]/NET0131  & n4511 ;
  assign n4748 = \P4_datao_reg[15]/NET0131  & n4507 ;
  assign n4749 = ~n4747 & ~n4748 ;
  assign n4750 = n4431 & ~n4749 ;
  assign n4751 = ~n4431 & n4749 ;
  assign n4752 = ~n4750 & ~n4751 ;
  assign n4753 = ~n4746 & ~n4752 ;
  assign n4754 = ~n4745 & ~n4753 ;
  assign n4755 = ~n4732 & ~n4754 ;
  assign n4756 = ~n4731 & ~n4755 ;
  assign n4757 = ~n4602 & ~n4603 ;
  assign n4758 = ~n4618 & n4757 ;
  assign n4759 = n4618 & ~n4757 ;
  assign n4760 = ~n4758 & ~n4759 ;
  assign n4761 = n4756 & ~n4760 ;
  assign n4762 = ~n4756 & n4760 ;
  assign n4763 = ~n4672 & ~n4673 ;
  assign n4764 = ~n4697 & n4763 ;
  assign n4765 = n4697 & ~n4763 ;
  assign n4766 = ~n4764 & ~n4765 ;
  assign n4767 = ~n4762 & n4766 ;
  assign n4768 = ~n4761 & ~n4767 ;
  assign n4769 = ~n4704 & ~n4768 ;
  assign n4770 = ~n4703 & ~n4769 ;
  assign n4771 = \P4_datao_reg[21]/NET0131  & n4407 ;
  assign n4772 = \P4_datao_reg[20]/NET0131  & n4405 ;
  assign n4773 = ~n4771 & ~n4772 ;
  assign n4774 = n4398 & ~n4773 ;
  assign n4775 = ~n4398 & n4773 ;
  assign n4776 = ~n4774 & ~n4775 ;
  assign n4777 = \P4_datao_reg[13]/NET0131  & n4376 ;
  assign n4778 = \P4_datao_reg[12]/NET0131  & n4374 ;
  assign n4779 = ~n4777 & ~n4778 ;
  assign n4780 = n4368 & ~n4779 ;
  assign n4781 = ~n4368 & n4779 ;
  assign n4782 = ~n4780 & ~n4781 ;
  assign n4783 = \P4_datao_reg[11]/NET0131  & n4390 ;
  assign n4784 = \P4_datao_reg[10]/NET0131  & n4388 ;
  assign n4785 = ~n4783 & ~n4784 ;
  assign n4786 = n4382 & ~n4785 ;
  assign n4787 = ~n4382 & n4785 ;
  assign n4788 = ~n4786 & ~n4787 ;
  assign n4789 = n4782 & n4788 ;
  assign n4790 = ~n4782 & ~n4788 ;
  assign n4791 = ~n4789 & ~n4790 ;
  assign n4792 = n4776 & ~n4791 ;
  assign n4793 = ~n4776 & n4791 ;
  assign n4794 = ~n4792 & ~n4793 ;
  assign n4795 = \P4_datao_reg[15]/NET0131  & n4356 ;
  assign n4796 = \P4_datao_reg[14]/NET0131  & n4360 ;
  assign n4797 = ~n4795 & ~n4796 ;
  assign n4798 = n4351 & ~n4797 ;
  assign n4799 = ~n4351 & n4797 ;
  assign n4800 = ~n4798 & ~n4799 ;
  assign n4801 = \P4_datao_reg[2]/NET0131  & n4460 ;
  assign n4802 = \P4_datao_reg[3]/NET0131  & n4421 ;
  assign n4803 = ~n4801 & ~n4802 ;
  assign n4804 = ~n4447 & n4803 ;
  assign n4805 = n4447 & ~n4803 ;
  assign n4806 = ~n4804 & ~n4805 ;
  assign n4807 = \din[27]_pad  & sel_pad ;
  assign n4808 = \din[26]_pad  & n4447 ;
  assign n4809 = ~n4807 & ~n4808 ;
  assign n4810 = ~\din[25]_pad  & ~\din[26]_pad  ;
  assign n4811 = sel_pad & ~n4810 ;
  assign n4812 = \din[27]_pad  & n4811 ;
  assign n4813 = ~n4809 & ~n4812 ;
  assign n4814 = \P4_datao_reg[0]/NET0131  & n4813 ;
  assign n4815 = ~n4808 & n4811 ;
  assign n4816 = \P4_datao_reg[1]/NET0131  & n4815 ;
  assign n4817 = ~n4814 & ~n4816 ;
  assign n4818 = ~n4807 & n4817 ;
  assign n4819 = n4807 & ~n4817 ;
  assign n4820 = ~n4818 & ~n4819 ;
  assign n4821 = n4806 & n4820 ;
  assign n4822 = ~n4806 & ~n4820 ;
  assign n4823 = ~n4821 & ~n4822 ;
  assign n4824 = n4800 & ~n4823 ;
  assign n4825 = ~n4800 & n4823 ;
  assign n4826 = ~n4824 & ~n4825 ;
  assign n4827 = n4794 & n4826 ;
  assign n4828 = ~n4794 & ~n4826 ;
  assign n4829 = ~n4827 & ~n4828 ;
  assign n4830 = \P4_datao_reg[22]/NET0131  & n4552 ;
  assign n4831 = \P4_datao_reg[23]/NET0131  & n4548 ;
  assign n4832 = ~n4830 & ~n4831 ;
  assign n4833 = n4399 & ~n4832 ;
  assign n4834 = ~n4399 & n4832 ;
  assign n4835 = ~n4833 & ~n4834 ;
  assign n4836 = \P4_datao_reg[16]/NET0131  & n4439 ;
  assign n4837 = \P4_datao_reg[17]/NET0131  & n4435 ;
  assign n4838 = ~n4836 & ~n4837 ;
  assign n4839 = ~n4352 & n4838 ;
  assign n4840 = n4352 & ~n4838 ;
  assign n4841 = ~n4839 & ~n4840 ;
  assign n4842 = \P4_datao_reg[4]/NET0131  & n4566 ;
  assign n4843 = \P4_datao_reg[5]/NET0131  & n4562 ;
  assign n4844 = ~n4842 & ~n4843 ;
  assign n4845 = ~n4417 & n4844 ;
  assign n4846 = n4417 & ~n4844 ;
  assign n4847 = ~n4845 & ~n4846 ;
  assign n4848 = n4841 & n4847 ;
  assign n4849 = ~n4841 & ~n4847 ;
  assign n4850 = ~n4848 & ~n4849 ;
  assign n4851 = n4835 & ~n4850 ;
  assign n4852 = ~n4835 & n4850 ;
  assign n4853 = ~n4851 & ~n4852 ;
  assign n4854 = n4829 & n4853 ;
  assign n4855 = ~n4829 & ~n4853 ;
  assign n4856 = ~n4854 & ~n4855 ;
  assign n4857 = \P4_datao_reg[22]/NET0131  & n4548 ;
  assign n4858 = \P4_datao_reg[21]/NET0131  & n4552 ;
  assign n4859 = ~n4857 & ~n4858 ;
  assign n4860 = n4399 & ~n4859 ;
  assign n4861 = ~n4399 & n4859 ;
  assign n4862 = ~n4860 & ~n4861 ;
  assign n4863 = \P4_datao_reg[14]/NET0131  & n4356 ;
  assign n4864 = \P4_datao_reg[13]/NET0131  & n4360 ;
  assign n4865 = ~n4863 & ~n4864 ;
  assign n4866 = n4351 & ~n4865 ;
  assign n4867 = ~n4351 & n4865 ;
  assign n4868 = ~n4866 & ~n4867 ;
  assign n4869 = n4862 & n4868 ;
  assign n4870 = ~n4862 & ~n4868 ;
  assign n4871 = ~n4869 & ~n4870 ;
  assign n4872 = ~n4616 & n4871 ;
  assign n4873 = n4616 & ~n4871 ;
  assign n4874 = ~n4872 & ~n4873 ;
  assign n4875 = \P4_datao_reg[0]/NET0131  & n4815 ;
  assign n4876 = \P4_datao_reg[20]/NET0131  & n4407 ;
  assign n4877 = \P4_datao_reg[19]/NET0131  & n4405 ;
  assign n4878 = ~n4876 & ~n4877 ;
  assign n4879 = n4398 & ~n4878 ;
  assign n4880 = ~n4398 & n4878 ;
  assign n4881 = ~n4879 & ~n4880 ;
  assign n4882 = ~n4875 & ~n4881 ;
  assign n4883 = n4875 & n4881 ;
  assign n4884 = ~n4882 & ~n4883 ;
  assign n4885 = \P4_datao_reg[23]/NET0131  & n4335 ;
  assign n4886 = \P4_datao_reg[24]/NET0131  & n4337 ;
  assign n4887 = ~n4885 & ~n4886 ;
  assign n4888 = n4328 & ~n4887 ;
  assign n4889 = ~n4328 & n4887 ;
  assign n4890 = ~n4888 & ~n4889 ;
  assign n4891 = n4884 & ~n4890 ;
  assign n4892 = ~n4884 & n4890 ;
  assign n4893 = ~n4891 & ~n4892 ;
  assign n4894 = ~n4874 & ~n4893 ;
  assign n4895 = n4874 & n4893 ;
  assign n4896 = \P4_datao_reg[4]/NET0131  & n4562 ;
  assign n4897 = \P4_datao_reg[3]/NET0131  & n4566 ;
  assign n4898 = ~n4896 & ~n4897 ;
  assign n4899 = n4417 & ~n4898 ;
  assign n4900 = ~n4417 & n4898 ;
  assign n4901 = ~n4899 & ~n4900 ;
  assign n4902 = \P4_datao_reg[2]/NET0131  & n4421 ;
  assign n4903 = \P4_datao_reg[1]/NET0131  & n4460 ;
  assign n4904 = ~n4902 & ~n4903 ;
  assign n4905 = n4447 & ~n4904 ;
  assign n4906 = ~n4447 & n4904 ;
  assign n4907 = ~n4905 & ~n4906 ;
  assign n4908 = \P4_datao_reg[26]/NET0131  & n4343 ;
  assign n4909 = ~\din[1]_pad  & n4908 ;
  assign n4910 = \P4_datao_reg[25]/NET0131  & ~n4343 ;
  assign n4911 = n4329 & ~n4908 ;
  assign n4912 = ~n4910 & n4911 ;
  assign n4913 = ~n4909 & ~n4912 ;
  assign n4914 = n4907 & ~n4913 ;
  assign n4915 = ~n4907 & n4913 ;
  assign n4916 = ~n4914 & ~n4915 ;
  assign n4917 = n4901 & ~n4916 ;
  assign n4918 = ~n4901 & n4916 ;
  assign n4919 = ~n4917 & ~n4918 ;
  assign n4920 = ~n4895 & ~n4919 ;
  assign n4921 = ~n4894 & ~n4920 ;
  assign n4922 = n4856 & n4921 ;
  assign n4923 = ~n4856 & ~n4921 ;
  assign n4924 = ~n4922 & ~n4923 ;
  assign n4925 = ~n4616 & ~n4869 ;
  assign n4926 = ~n4870 & ~n4925 ;
  assign n4927 = \P4_datao_reg[18]/NET0131  & n4511 ;
  assign n4928 = \P4_datao_reg[19]/NET0131  & n4507 ;
  assign n4929 = ~n4927 & ~n4928 ;
  assign n4930 = ~n4431 & n4929 ;
  assign n4931 = n4431 & ~n4929 ;
  assign n4932 = ~n4930 & ~n4931 ;
  assign n4933 = \P4_datao_reg[9]/NET0131  & n4525 ;
  assign n4934 = \P4_datao_reg[8]/NET0131  & n4523 ;
  assign n4935 = ~n4933 & ~n4934 ;
  assign n4936 = n4517 & ~n4935 ;
  assign n4937 = ~n4517 & n4935 ;
  assign n4938 = ~n4936 & ~n4937 ;
  assign n4939 = \P4_datao_reg[6]/NET0131  & n4580 ;
  assign n4940 = \P4_datao_reg[7]/NET0131  & n4575 ;
  assign n4941 = ~n4939 & ~n4940 ;
  assign n4942 = n4558 & ~n4941 ;
  assign n4943 = ~n4558 & n4941 ;
  assign n4944 = ~n4942 & ~n4943 ;
  assign n4945 = n4938 & n4944 ;
  assign n4946 = ~n4938 & ~n4944 ;
  assign n4947 = ~n4945 & ~n4946 ;
  assign n4948 = n4932 & ~n4947 ;
  assign n4949 = ~n4932 & n4947 ;
  assign n4950 = ~n4948 & ~n4949 ;
  assign n4951 = n4926 & ~n4950 ;
  assign n4952 = ~n4926 & n4950 ;
  assign n4953 = ~n4951 & ~n4952 ;
  assign n4954 = n4807 & ~n4875 ;
  assign n4955 = \P4_datao_reg[24]/NET0131  & n4335 ;
  assign n4956 = \P4_datao_reg[25]/NET0131  & n4337 ;
  assign n4957 = ~n4955 & ~n4956 ;
  assign n4958 = n4328 & ~n4957 ;
  assign n4959 = ~n4328 & n4957 ;
  assign n4960 = ~n4958 & ~n4959 ;
  assign n4961 = \P4_datao_reg[27]/NET0131  & n4343 ;
  assign n4962 = ~\din[1]_pad  & n4961 ;
  assign n4963 = \P4_datao_reg[26]/NET0131  & ~n4343 ;
  assign n4964 = n4329 & ~n4961 ;
  assign n4965 = ~n4963 & n4964 ;
  assign n4966 = ~n4962 & ~n4965 ;
  assign n4967 = n4960 & ~n4966 ;
  assign n4968 = ~n4960 & n4966 ;
  assign n4969 = ~n4967 & ~n4968 ;
  assign n4970 = n4954 & n4969 ;
  assign n4971 = ~n4954 & ~n4969 ;
  assign n4972 = ~n4970 & ~n4971 ;
  assign n4973 = ~n4882 & n4890 ;
  assign n4974 = ~n4883 & ~n4973 ;
  assign n4975 = n4972 & ~n4974 ;
  assign n4976 = ~n4972 & n4974 ;
  assign n4977 = ~n4975 & ~n4976 ;
  assign n4978 = n4953 & ~n4977 ;
  assign n4979 = ~n4953 & n4977 ;
  assign n4980 = ~n4978 & ~n4979 ;
  assign n4981 = n4924 & n4980 ;
  assign n4982 = ~n4924 & ~n4980 ;
  assign n4983 = ~n4981 & ~n4982 ;
  assign n4984 = ~n4770 & ~n4983 ;
  assign n4985 = n4770 & n4983 ;
  assign n4986 = ~n4984 & ~n4985 ;
  assign n4987 = ~n4622 & n4699 ;
  assign n4988 = ~n4621 & ~n4987 ;
  assign n4989 = ~n4653 & ~n4667 ;
  assign n4990 = ~n4666 & ~n4989 ;
  assign n4991 = \P4_datao_reg[12]/NET0131  & n4376 ;
  assign n4992 = \P4_datao_reg[11]/NET0131  & n4374 ;
  assign n4993 = ~n4991 & ~n4992 ;
  assign n4994 = n4368 & ~n4993 ;
  assign n4995 = ~n4368 & n4993 ;
  assign n4996 = ~n4994 & ~n4995 ;
  assign n4997 = \P4_datao_reg[10]/NET0131  & n4390 ;
  assign n4998 = \P4_datao_reg[9]/NET0131  & n4388 ;
  assign n4999 = ~n4997 & ~n4998 ;
  assign n5000 = n4382 & ~n4999 ;
  assign n5001 = ~n4382 & n4999 ;
  assign n5002 = ~n5000 & ~n5001 ;
  assign n5003 = n4996 & n5002 ;
  assign n5004 = ~n4996 & ~n5002 ;
  assign n5005 = ~n5003 & ~n5004 ;
  assign n5006 = \P4_datao_reg[18]/NET0131  & n4507 ;
  assign n5007 = \P4_datao_reg[17]/NET0131  & n4511 ;
  assign n5008 = ~n5006 & ~n5007 ;
  assign n5009 = n4431 & ~n5008 ;
  assign n5010 = ~n4431 & n5008 ;
  assign n5011 = ~n5009 & ~n5010 ;
  assign n5012 = n5005 & ~n5011 ;
  assign n5013 = ~n5005 & n5011 ;
  assign n5014 = ~n5012 & ~n5013 ;
  assign n5015 = n4990 & ~n5014 ;
  assign n5016 = ~n4990 & n5014 ;
  assign n5017 = \P4_datao_reg[7]/NET0131  & n4523 ;
  assign n5018 = \P4_datao_reg[8]/NET0131  & n4525 ;
  assign n5019 = ~n5017 & ~n5018 ;
  assign n5020 = ~n4517 & n5019 ;
  assign n5021 = n4517 & ~n5019 ;
  assign n5022 = ~n5020 & ~n5021 ;
  assign n5023 = \P4_datao_reg[6]/NET0131  & n4575 ;
  assign n5024 = \P4_datao_reg[5]/NET0131  & n4580 ;
  assign n5025 = ~n5023 & ~n5024 ;
  assign n5026 = n4558 & ~n5025 ;
  assign n5027 = ~n4558 & n5025 ;
  assign n5028 = ~n5026 & ~n5027 ;
  assign n5029 = ~n5022 & ~n5028 ;
  assign n5030 = n5022 & n5028 ;
  assign n5031 = ~n5029 & ~n5030 ;
  assign n5032 = \P4_datao_reg[16]/NET0131  & n4435 ;
  assign n5033 = \P4_datao_reg[15]/NET0131  & n4439 ;
  assign n5034 = ~n5032 & ~n5033 ;
  assign n5035 = n4352 & ~n5034 ;
  assign n5036 = ~n4352 & n5034 ;
  assign n5037 = ~n5035 & ~n5036 ;
  assign n5038 = n5031 & ~n5037 ;
  assign n5039 = ~n5031 & n5037 ;
  assign n5040 = ~n5038 & ~n5039 ;
  assign n5041 = ~n5016 & ~n5040 ;
  assign n5042 = ~n5015 & ~n5041 ;
  assign n5043 = n4901 & ~n4915 ;
  assign n5044 = ~n4914 & ~n5043 ;
  assign n5045 = ~n5029 & n5037 ;
  assign n5046 = ~n5030 & ~n5045 ;
  assign n5047 = ~n5004 & n5011 ;
  assign n5048 = ~n5003 & ~n5047 ;
  assign n5049 = n5046 & ~n5048 ;
  assign n5050 = ~n5046 & n5048 ;
  assign n5051 = ~n5049 & ~n5050 ;
  assign n5052 = n5044 & n5051 ;
  assign n5053 = ~n5044 & ~n5051 ;
  assign n5054 = ~n5052 & ~n5053 ;
  assign n5055 = ~n5042 & n5054 ;
  assign n5056 = n5042 & ~n5054 ;
  assign n5057 = ~n5055 & ~n5056 ;
  assign n5058 = ~n4629 & ~n4643 ;
  assign n5059 = ~n4642 & ~n5058 ;
  assign n5060 = ~n4456 & n4466 ;
  assign n5061 = ~n4455 & ~n5060 ;
  assign n5062 = n5059 & ~n5061 ;
  assign n5063 = ~n5059 & n5061 ;
  assign n5064 = ~n4679 & ~n4692 ;
  assign n5065 = ~n4693 & ~n5064 ;
  assign n5066 = ~n5063 & n5065 ;
  assign n5067 = ~n5062 & ~n5066 ;
  assign n5068 = n5057 & n5067 ;
  assign n5069 = ~n5057 & ~n5067 ;
  assign n5070 = ~n5068 & ~n5069 ;
  assign n5071 = n4988 & ~n5070 ;
  assign n5072 = ~n4988 & n5070 ;
  assign n5073 = ~n5071 & ~n5072 ;
  assign n5074 = ~n5062 & ~n5063 ;
  assign n5075 = n5065 & n5074 ;
  assign n5076 = ~n5065 & ~n5074 ;
  assign n5077 = ~n5075 & ~n5076 ;
  assign n5078 = ~n5015 & ~n5016 ;
  assign n5079 = ~n5040 & n5078 ;
  assign n5080 = n5040 & ~n5078 ;
  assign n5081 = ~n5079 & ~n5080 ;
  assign n5082 = ~n5077 & ~n5081 ;
  assign n5083 = n5077 & n5081 ;
  assign n5084 = ~n4894 & ~n4895 ;
  assign n5085 = ~n4919 & n5084 ;
  assign n5086 = n4919 & ~n5084 ;
  assign n5087 = ~n5085 & ~n5086 ;
  assign n5088 = ~n5083 & ~n5087 ;
  assign n5089 = ~n5082 & ~n5088 ;
  assign n5090 = n5073 & ~n5089 ;
  assign n5091 = ~n5073 & n5089 ;
  assign n5092 = ~n5090 & ~n5091 ;
  assign n5093 = n4986 & n5092 ;
  assign n5094 = ~n4986 & ~n5092 ;
  assign n5095 = ~n5093 & ~n5094 ;
  assign n5096 = \P4_datao_reg[15]/NET0131  & n4405 ;
  assign n5097 = \P4_datao_reg[16]/NET0131  & n4407 ;
  assign n5098 = ~n5096 & ~n5097 ;
  assign n5099 = ~n4398 & n5098 ;
  assign n5100 = n4398 & ~n5098 ;
  assign n5101 = ~n5099 & ~n5100 ;
  assign n5102 = \P4_datao_reg[0]/NET0131  & n4562 ;
  assign n5103 = ~n5101 & ~n5102 ;
  assign n5104 = n5101 & n5102 ;
  assign n5105 = \P4_datao_reg[19]/NET0131  & n4335 ;
  assign n5106 = \P4_datao_reg[20]/NET0131  & n4337 ;
  assign n5107 = ~n5105 & ~n5106 ;
  assign n5108 = ~n4328 & n5107 ;
  assign n5109 = n4328 & ~n5107 ;
  assign n5110 = ~n5108 & ~n5109 ;
  assign n5111 = ~n5104 & ~n5110 ;
  assign n5112 = ~n5103 & ~n5111 ;
  assign n5113 = \P4_datao_reg[9]/NET0131  & n4360 ;
  assign n5114 = \P4_datao_reg[10]/NET0131  & n4356 ;
  assign n5115 = ~n5113 & ~n5114 ;
  assign n5116 = ~n4351 & n5115 ;
  assign n5117 = n4351 & ~n5115 ;
  assign n5118 = ~n5116 & ~n5117 ;
  assign n5119 = \P4_datao_reg[12]/NET0131  & n4435 ;
  assign n5120 = \P4_datao_reg[11]/NET0131  & n4439 ;
  assign n5121 = ~n5119 & ~n5120 ;
  assign n5122 = n4352 & ~n5121 ;
  assign n5123 = ~n4352 & n5121 ;
  assign n5124 = ~n5122 & ~n5123 ;
  assign n5125 = ~n5118 & ~n5124 ;
  assign n5126 = n5118 & n5124 ;
  assign n5127 = \P4_datao_reg[17]/NET0131  & n4552 ;
  assign n5128 = \P4_datao_reg[18]/NET0131  & n4548 ;
  assign n5129 = ~n5127 & ~n5128 ;
  assign n5130 = ~n4399 & n5129 ;
  assign n5131 = n4399 & ~n5129 ;
  assign n5132 = ~n5130 & ~n5131 ;
  assign n5133 = ~n5126 & ~n5132 ;
  assign n5134 = ~n5125 & ~n5133 ;
  assign n5135 = n5112 & n5134 ;
  assign n5136 = ~n5112 & ~n5134 ;
  assign n5137 = \P4_datao_reg[1]/NET0131  & n4580 ;
  assign n5138 = \P4_datao_reg[2]/NET0131  & n4575 ;
  assign n5139 = ~n5137 & ~n5138 ;
  assign n5140 = n4558 & ~n5139 ;
  assign n5141 = ~n4558 & n5139 ;
  assign n5142 = ~n5140 & ~n5141 ;
  assign n5143 = \P4_datao_reg[3]/NET0131  & n4523 ;
  assign n5144 = \P4_datao_reg[4]/NET0131  & n4525 ;
  assign n5145 = ~n5143 & ~n5144 ;
  assign n5146 = n4517 & ~n5145 ;
  assign n5147 = ~n4517 & n5145 ;
  assign n5148 = ~n5146 & ~n5147 ;
  assign n5149 = n5142 & n5148 ;
  assign n5150 = ~n5142 & ~n5148 ;
  assign n5151 = \P4_datao_reg[22]/NET0131  & n4343 ;
  assign n5152 = ~\din[1]_pad  & n5151 ;
  assign n5153 = \P4_datao_reg[21]/NET0131  & ~n4343 ;
  assign n5154 = n4329 & ~n5151 ;
  assign n5155 = ~n5153 & n5154 ;
  assign n5156 = ~n5152 & ~n5155 ;
  assign n5157 = ~n5150 & ~n5156 ;
  assign n5158 = ~n5149 & ~n5157 ;
  assign n5159 = ~n5136 & ~n5158 ;
  assign n5160 = ~n5135 & ~n5159 ;
  assign n5161 = \P4_datao_reg[10]/NET0131  & n4360 ;
  assign n5162 = \P4_datao_reg[11]/NET0131  & n4356 ;
  assign n5163 = ~n5161 & ~n5162 ;
  assign n5164 = ~n4351 & n5163 ;
  assign n5165 = n4351 & ~n5163 ;
  assign n5166 = ~n5164 & ~n5165 ;
  assign n5167 = n4417 & ~n5102 ;
  assign n5168 = n5166 & n5167 ;
  assign n5169 = ~n5166 & ~n5167 ;
  assign n5170 = ~n4342 & n4349 ;
  assign n5171 = ~n4350 & ~n5170 ;
  assign n5172 = ~n5169 & n5171 ;
  assign n5173 = ~n5168 & ~n5172 ;
  assign n5174 = ~n5160 & ~n5173 ;
  assign n5175 = n5160 & n5173 ;
  assign n5176 = ~n4366 & ~n4367 ;
  assign n5177 = ~n4414 & n5176 ;
  assign n5178 = n4414 & ~n5176 ;
  assign n5179 = ~n5177 & ~n5178 ;
  assign n5180 = ~n5175 & ~n5179 ;
  assign n5181 = ~n5174 & ~n5180 ;
  assign n5182 = ~n4731 & ~n4732 ;
  assign n5183 = ~n4754 & n5182 ;
  assign n5184 = n4754 & ~n5182 ;
  assign n5185 = ~n5183 & ~n5184 ;
  assign n5186 = \P4_datao_reg[7]/NET0131  & n4374 ;
  assign n5187 = \P4_datao_reg[8]/NET0131  & n4376 ;
  assign n5188 = ~n5186 & ~n5187 ;
  assign n5189 = n4368 & ~n5188 ;
  assign n5190 = ~n4368 & n5188 ;
  assign n5191 = ~n5189 & ~n5190 ;
  assign n5192 = \P4_datao_reg[13]/NET0131  & n4511 ;
  assign n5193 = \P4_datao_reg[14]/NET0131  & n4507 ;
  assign n5194 = ~n5192 & ~n5193 ;
  assign n5195 = n4431 & ~n5194 ;
  assign n5196 = ~n4431 & n5194 ;
  assign n5197 = ~n5195 & ~n5196 ;
  assign n5198 = ~n5191 & ~n5197 ;
  assign n5199 = n5191 & n5197 ;
  assign n5200 = \P4_datao_reg[5]/NET0131  & n4388 ;
  assign n5201 = \P4_datao_reg[6]/NET0131  & n4390 ;
  assign n5202 = ~n5200 & ~n5201 ;
  assign n5203 = n4382 & ~n5202 ;
  assign n5204 = ~n4382 & n5202 ;
  assign n5205 = ~n5203 & ~n5204 ;
  assign n5206 = ~n5199 & ~n5205 ;
  assign n5207 = ~n5198 & ~n5206 ;
  assign n5208 = ~n4717 & ~n4718 ;
  assign n5209 = ~n4724 & n5208 ;
  assign n5210 = n4724 & ~n5208 ;
  assign n5211 = ~n5209 & ~n5210 ;
  assign n5212 = n5207 & ~n5211 ;
  assign n5213 = ~n5207 & n5211 ;
  assign n5214 = ~n4745 & ~n4746 ;
  assign n5215 = n4752 & n5214 ;
  assign n5216 = ~n4752 & ~n5214 ;
  assign n5217 = ~n5215 & ~n5216 ;
  assign n5218 = ~n5213 & n5217 ;
  assign n5219 = ~n5212 & ~n5218 ;
  assign n5220 = ~n5185 & ~n5219 ;
  assign n5221 = n5185 & n5219 ;
  assign n5222 = ~n4543 & ~n4544 ;
  assign n5223 = ~n4591 & n5222 ;
  assign n5224 = n4591 & ~n5222 ;
  assign n5225 = ~n5223 & ~n5224 ;
  assign n5226 = ~n5221 & ~n5225 ;
  assign n5227 = ~n5220 & ~n5226 ;
  assign n5228 = ~n5181 & ~n5227 ;
  assign n5229 = n5181 & n5227 ;
  assign n5230 = ~n4498 & ~n4499 ;
  assign n5231 = ~n4593 & n5230 ;
  assign n5232 = n4593 & ~n5230 ;
  assign n5233 = ~n5231 & ~n5232 ;
  assign n5234 = ~n5229 & ~n5233 ;
  assign n5235 = ~n5228 & ~n5234 ;
  assign n5236 = ~n5082 & ~n5083 ;
  assign n5237 = ~n5087 & n5236 ;
  assign n5238 = n5087 & ~n5236 ;
  assign n5239 = ~n5237 & ~n5238 ;
  assign n5240 = ~n5235 & ~n5239 ;
  assign n5241 = n5235 & n5239 ;
  assign n5242 = ~n4703 & ~n4704 ;
  assign n5243 = ~n4768 & n5242 ;
  assign n5244 = n4768 & ~n5242 ;
  assign n5245 = ~n5243 & ~n5244 ;
  assign n5246 = ~n5241 & n5245 ;
  assign n5247 = ~n5240 & ~n5246 ;
  assign n5248 = n5095 & n5247 ;
  assign n5249 = ~n5072 & n5089 ;
  assign n5250 = ~n5071 & ~n5249 ;
  assign n5251 = \P4_datao_reg[10]/NET0131  & n4525 ;
  assign n5252 = \P4_datao_reg[9]/NET0131  & n4523 ;
  assign n5253 = ~n5251 & ~n5252 ;
  assign n5254 = n4517 & ~n5253 ;
  assign n5255 = ~n4517 & n5253 ;
  assign n5256 = ~n5254 & ~n5255 ;
  assign n5257 = \P4_datao_reg[7]/NET0131  & n4580 ;
  assign n5258 = \P4_datao_reg[8]/NET0131  & n4575 ;
  assign n5259 = ~n5257 & ~n5258 ;
  assign n5260 = n4558 & ~n5259 ;
  assign n5261 = ~n4558 & n5259 ;
  assign n5262 = ~n5260 & ~n5261 ;
  assign n5263 = n5256 & n5262 ;
  assign n5264 = ~n5256 & ~n5262 ;
  assign n5265 = ~n5263 & ~n5264 ;
  assign n5266 = \P4_datao_reg[28]/NET0131  & n4343 ;
  assign n5267 = ~\din[1]_pad  & n5266 ;
  assign n5268 = \P4_datao_reg[27]/NET0131  & ~n4343 ;
  assign n5269 = n4329 & ~n5266 ;
  assign n5270 = ~n5268 & n5269 ;
  assign n5271 = ~n5267 & ~n5270 ;
  assign n5272 = n5265 & n5271 ;
  assign n5273 = ~n5265 & ~n5271 ;
  assign n5274 = ~n5272 & ~n5273 ;
  assign n5275 = \P4_datao_reg[23]/NET0131  & n4552 ;
  assign n5276 = \P4_datao_reg[24]/NET0131  & n4548 ;
  assign n5277 = ~n5275 & ~n5276 ;
  assign n5278 = ~n4399 & n5277 ;
  assign n5279 = n4399 & ~n5277 ;
  assign n5280 = ~n5278 & ~n5279 ;
  assign n5281 = \P4_datao_reg[2]/NET0131  & n4815 ;
  assign n5282 = \P4_datao_reg[1]/NET0131  & n4813 ;
  assign n5283 = ~n5281 & ~n5282 ;
  assign n5284 = ~n4807 & n5283 ;
  assign n5285 = n4807 & ~n5283 ;
  assign n5286 = ~n5284 & ~n5285 ;
  assign n5287 = \P4_datao_reg[16]/NET0131  & n4356 ;
  assign n5288 = \P4_datao_reg[15]/NET0131  & n4360 ;
  assign n5289 = ~n5287 & ~n5288 ;
  assign n5290 = n4351 & ~n5289 ;
  assign n5291 = ~n4351 & n5289 ;
  assign n5292 = ~n5290 & ~n5291 ;
  assign n5293 = n5286 & n5292 ;
  assign n5294 = ~n5286 & ~n5292 ;
  assign n5295 = ~n5293 & ~n5294 ;
  assign n5296 = n5280 & n5295 ;
  assign n5297 = ~n5280 & ~n5295 ;
  assign n5298 = ~n5296 & ~n5297 ;
  assign n5299 = n5274 & ~n5298 ;
  assign n5300 = ~n5274 & n5298 ;
  assign n5301 = ~n5299 & ~n5300 ;
  assign n5302 = \P4_datao_reg[14]/NET0131  & n4376 ;
  assign n5303 = \P4_datao_reg[13]/NET0131  & n4374 ;
  assign n5304 = ~n5302 & ~n5303 ;
  assign n5305 = n4368 & ~n5304 ;
  assign n5306 = ~n4368 & n5304 ;
  assign n5307 = ~n5305 & ~n5306 ;
  assign n5308 = \P4_datao_reg[12]/NET0131  & n4390 ;
  assign n5309 = \P4_datao_reg[11]/NET0131  & n4388 ;
  assign n5310 = ~n5308 & ~n5309 ;
  assign n5311 = n4382 & ~n5310 ;
  assign n5312 = ~n4382 & n5310 ;
  assign n5313 = ~n5311 & ~n5312 ;
  assign n5314 = n5307 & n5313 ;
  assign n5315 = ~n5307 & ~n5313 ;
  assign n5316 = ~n5314 & ~n5315 ;
  assign n5317 = \P4_datao_reg[20]/NET0131  & n4507 ;
  assign n5318 = \P4_datao_reg[19]/NET0131  & n4511 ;
  assign n5319 = ~n5317 & ~n5318 ;
  assign n5320 = n4431 & ~n5319 ;
  assign n5321 = ~n4431 & n5319 ;
  assign n5322 = ~n5320 & ~n5321 ;
  assign n5323 = n5316 & ~n5322 ;
  assign n5324 = ~n5316 & n5322 ;
  assign n5325 = ~n5323 & ~n5324 ;
  assign n5326 = n5301 & ~n5325 ;
  assign n5327 = ~n5301 & n5325 ;
  assign n5328 = ~n5326 & ~n5327 ;
  assign n5329 = ~n5056 & ~n5067 ;
  assign n5330 = ~n5055 & ~n5329 ;
  assign n5331 = n5328 & ~n5330 ;
  assign n5332 = ~n5328 & n5330 ;
  assign n5333 = ~n5331 & ~n5332 ;
  assign n5334 = ~n4952 & n4977 ;
  assign n5335 = ~n4951 & ~n5334 ;
  assign n5336 = n5333 & n5335 ;
  assign n5337 = ~n5333 & ~n5335 ;
  assign n5338 = ~n5336 & ~n5337 ;
  assign n5339 = ~n5250 & ~n5338 ;
  assign n5340 = n5250 & n5338 ;
  assign n5341 = ~n5339 & ~n5340 ;
  assign n5342 = ~n4932 & ~n4945 ;
  assign n5343 = ~n4946 & ~n5342 ;
  assign n5344 = n4967 & n5343 ;
  assign n5345 = ~n4967 & ~n5343 ;
  assign n5346 = ~n5344 & ~n5345 ;
  assign n5347 = ~n4776 & ~n4789 ;
  assign n5348 = ~n4790 & ~n5347 ;
  assign n5349 = ~n5346 & n5348 ;
  assign n5350 = ~n5344 & ~n5348 ;
  assign n5351 = ~n5345 & n5350 ;
  assign n5352 = ~n5349 & ~n5351 ;
  assign n5353 = ~n4835 & ~n4848 ;
  assign n5354 = ~n4849 & ~n5353 ;
  assign n5355 = ~n4800 & ~n4821 ;
  assign n5356 = ~n4822 & ~n5355 ;
  assign n5357 = n5354 & n5356 ;
  assign n5358 = ~n5354 & ~n5356 ;
  assign n5359 = ~n5357 & ~n5358 ;
  assign n5360 = \din[28]_pad  & n4807 ;
  assign n5361 = ~\din[27]_pad  & ~\din[28]_pad  ;
  assign n5362 = sel_pad & ~n5361 ;
  assign n5363 = ~n5360 & n5362 ;
  assign n5364 = \P4_datao_reg[0]/NET0131  & n5363 ;
  assign n5365 = \P4_datao_reg[21]/NET0131  & n4405 ;
  assign n5366 = \P4_datao_reg[22]/NET0131  & n4407 ;
  assign n5367 = ~n5365 & ~n5366 ;
  assign n5368 = n4398 & ~n5367 ;
  assign n5369 = ~n4398 & n5367 ;
  assign n5370 = ~n5368 & ~n5369 ;
  assign n5371 = n5364 & n5370 ;
  assign n5372 = ~n5364 & ~n5370 ;
  assign n5373 = ~n5371 & ~n5372 ;
  assign n5374 = \P4_datao_reg[26]/NET0131  & n4337 ;
  assign n5375 = \P4_datao_reg[25]/NET0131  & n4335 ;
  assign n5376 = ~n5374 & ~n5375 ;
  assign n5377 = n4328 & ~n5376 ;
  assign n5378 = ~n4328 & n5376 ;
  assign n5379 = ~n5377 & ~n5378 ;
  assign n5380 = n5373 & ~n5379 ;
  assign n5381 = ~n5373 & n5379 ;
  assign n5382 = ~n5380 & ~n5381 ;
  assign n5383 = n5359 & ~n5382 ;
  assign n5384 = ~n5359 & n5382 ;
  assign n5385 = ~n5383 & ~n5384 ;
  assign n5386 = n5352 & ~n5385 ;
  assign n5387 = ~n5352 & n5385 ;
  assign n5388 = ~n5386 & ~n5387 ;
  assign n5389 = ~n4827 & ~n4853 ;
  assign n5390 = ~n4828 & ~n5389 ;
  assign n5391 = n5388 & n5390 ;
  assign n5392 = ~n5388 & ~n5390 ;
  assign n5393 = ~n5391 & ~n5392 ;
  assign n5394 = ~n4971 & ~n4974 ;
  assign n5395 = ~n4970 & ~n5394 ;
  assign n5396 = \P4_datao_reg[17]/NET0131  & n4439 ;
  assign n5397 = \P4_datao_reg[18]/NET0131  & n4435 ;
  assign n5398 = ~n5396 & ~n5397 ;
  assign n5399 = ~n4352 & n5398 ;
  assign n5400 = n4352 & ~n5398 ;
  assign n5401 = ~n5399 & ~n5400 ;
  assign n5402 = \P4_datao_reg[3]/NET0131  & n4460 ;
  assign n5403 = \P4_datao_reg[4]/NET0131  & n4421 ;
  assign n5404 = ~n5402 & ~n5403 ;
  assign n5405 = n4447 & ~n5404 ;
  assign n5406 = ~n4447 & n5404 ;
  assign n5407 = ~n5405 & ~n5406 ;
  assign n5408 = \P4_datao_reg[6]/NET0131  & n4562 ;
  assign n5409 = \P4_datao_reg[5]/NET0131  & n4566 ;
  assign n5410 = ~n5408 & ~n5409 ;
  assign n5411 = n4417 & ~n5410 ;
  assign n5412 = ~n4417 & n5410 ;
  assign n5413 = ~n5411 & ~n5412 ;
  assign n5414 = ~n5407 & ~n5413 ;
  assign n5415 = n5407 & n5413 ;
  assign n5416 = ~n5414 & ~n5415 ;
  assign n5417 = n5401 & n5416 ;
  assign n5418 = ~n5401 & ~n5416 ;
  assign n5419 = ~n5417 & ~n5418 ;
  assign n5420 = ~n5395 & n5419 ;
  assign n5421 = n5395 & ~n5419 ;
  assign n5422 = ~n5420 & ~n5421 ;
  assign n5423 = n5044 & n5046 ;
  assign n5424 = ~n5048 & ~n5423 ;
  assign n5425 = ~n5044 & ~n5046 ;
  assign n5426 = ~n5424 & ~n5425 ;
  assign n5427 = n5422 & n5426 ;
  assign n5428 = ~n5422 & ~n5426 ;
  assign n5429 = ~n5427 & ~n5428 ;
  assign n5430 = n5393 & n5429 ;
  assign n5431 = ~n5393 & ~n5429 ;
  assign n5432 = ~n5430 & ~n5431 ;
  assign n5433 = ~n4922 & ~n4980 ;
  assign n5434 = ~n4923 & ~n5433 ;
  assign n5435 = n5432 & ~n5434 ;
  assign n5436 = ~n5432 & n5434 ;
  assign n5437 = ~n5435 & ~n5436 ;
  assign n5438 = n5341 & ~n5437 ;
  assign n5439 = ~n5341 & n5437 ;
  assign n5440 = ~n5438 & ~n5439 ;
  assign n5441 = ~n4985 & ~n5092 ;
  assign n5442 = ~n4984 & ~n5441 ;
  assign n5443 = n5440 & n5442 ;
  assign n5444 = ~n5248 & ~n5443 ;
  assign n5445 = ~n5430 & ~n5434 ;
  assign n5446 = ~n5431 & ~n5445 ;
  assign n5447 = ~n5332 & ~n5335 ;
  assign n5448 = ~n5331 & ~n5447 ;
  assign n5449 = n5446 & n5448 ;
  assign n5450 = ~n5446 & ~n5448 ;
  assign n5451 = ~n5449 & ~n5450 ;
  assign n5452 = ~n5372 & n5379 ;
  assign n5453 = ~n5371 & ~n5452 ;
  assign n5454 = ~n5264 & ~n5271 ;
  assign n5455 = ~n5263 & ~n5454 ;
  assign n5456 = ~n5453 & ~n5455 ;
  assign n5457 = n5453 & n5455 ;
  assign n5458 = ~n5456 & ~n5457 ;
  assign n5459 = ~n5315 & n5322 ;
  assign n5460 = ~n5314 & ~n5459 ;
  assign n5461 = n5458 & ~n5460 ;
  assign n5462 = ~n5458 & n5460 ;
  assign n5463 = ~n5461 & ~n5462 ;
  assign n5464 = ~n5280 & ~n5293 ;
  assign n5465 = ~n5294 & ~n5464 ;
  assign n5466 = ~n5401 & ~n5415 ;
  assign n5467 = ~n5414 & ~n5466 ;
  assign n5468 = ~n5465 & ~n5467 ;
  assign n5469 = n5465 & n5467 ;
  assign n5470 = ~n5468 & ~n5469 ;
  assign n5471 = \P4_datao_reg[22]/NET0131  & n4405 ;
  assign n5472 = \P4_datao_reg[23]/NET0131  & n4407 ;
  assign n5473 = ~n5471 & ~n5472 ;
  assign n5474 = ~n4398 & n5473 ;
  assign n5475 = n4398 & ~n5473 ;
  assign n5476 = ~n5474 & ~n5475 ;
  assign n5477 = \P4_datao_reg[14]/NET0131  & n4374 ;
  assign n5478 = \P4_datao_reg[15]/NET0131  & n4376 ;
  assign n5479 = ~n5477 & ~n5478 ;
  assign n5480 = ~n4368 & n5479 ;
  assign n5481 = n4368 & ~n5479 ;
  assign n5482 = ~n5480 & ~n5481 ;
  assign n5483 = \din[29]_pad  & sel_pad ;
  assign n5484 = ~n5364 & n5483 ;
  assign n5485 = ~n5482 & ~n5484 ;
  assign n5486 = n5482 & n5484 ;
  assign n5487 = ~n5485 & ~n5486 ;
  assign n5488 = n5476 & n5487 ;
  assign n5489 = ~n5476 & ~n5487 ;
  assign n5490 = ~n5488 & ~n5489 ;
  assign n5491 = n5470 & ~n5490 ;
  assign n5492 = ~n5470 & n5490 ;
  assign n5493 = ~n5491 & ~n5492 ;
  assign n5494 = n5463 & ~n5493 ;
  assign n5495 = ~n5463 & n5493 ;
  assign n5496 = ~n5494 & ~n5495 ;
  assign n5497 = ~n5358 & ~n5382 ;
  assign n5498 = ~n5357 & ~n5497 ;
  assign n5499 = n5496 & ~n5498 ;
  assign n5500 = ~n5496 & n5498 ;
  assign n5501 = ~n5499 & ~n5500 ;
  assign n5502 = ~n5345 & ~n5350 ;
  assign n5503 = \P4_datao_reg[27]/NET0131  & n4337 ;
  assign n5504 = \P4_datao_reg[26]/NET0131  & n4335 ;
  assign n5505 = ~n5503 & ~n5504 ;
  assign n5506 = n4328 & ~n5505 ;
  assign n5507 = ~n4328 & n5505 ;
  assign n5508 = ~n5506 & ~n5507 ;
  assign n5509 = \P4_datao_reg[29]/NET0131  & n4343 ;
  assign n5510 = ~\din[1]_pad  & n5509 ;
  assign n5511 = \P4_datao_reg[28]/NET0131  & ~n4343 ;
  assign n5512 = n4329 & ~n5509 ;
  assign n5513 = ~n5511 & n5512 ;
  assign n5514 = ~n5510 & ~n5513 ;
  assign n5515 = n5508 & ~n5514 ;
  assign n5516 = ~n5508 & n5514 ;
  assign n5517 = ~n5515 & ~n5516 ;
  assign n5518 = \P4_datao_reg[2]/NET0131  & n4813 ;
  assign n5519 = \P4_datao_reg[3]/NET0131  & n4815 ;
  assign n5520 = ~n5518 & ~n5519 ;
  assign n5521 = n4807 & ~n5520 ;
  assign n5522 = ~n4807 & n5520 ;
  assign n5523 = ~n5521 & ~n5522 ;
  assign n5524 = \P4_datao_reg[1]/NET0131  & n5363 ;
  assign n5525 = ~n5360 & ~n5483 ;
  assign n5526 = \din[29]_pad  & n5362 ;
  assign n5527 = ~n5525 & ~n5526 ;
  assign n5528 = \P4_datao_reg[0]/NET0131  & n5527 ;
  assign n5529 = ~n5524 & ~n5528 ;
  assign n5530 = n5483 & ~n5529 ;
  assign n5531 = ~n5483 & n5529 ;
  assign n5532 = ~n5530 & ~n5531 ;
  assign n5533 = n5523 & n5532 ;
  assign n5534 = ~n5523 & ~n5532 ;
  assign n5535 = ~n5533 & ~n5534 ;
  assign n5536 = n5517 & ~n5535 ;
  assign n5537 = ~n5517 & n5535 ;
  assign n5538 = ~n5536 & ~n5537 ;
  assign n5539 = n5502 & ~n5538 ;
  assign n5540 = ~n5502 & n5538 ;
  assign n5541 = ~n5539 & ~n5540 ;
  assign n5542 = ~n5300 & n5325 ;
  assign n5543 = ~n5299 & ~n5542 ;
  assign n5544 = n5541 & ~n5543 ;
  assign n5545 = ~n5541 & n5543 ;
  assign n5546 = ~n5544 & ~n5545 ;
  assign n5547 = ~n5501 & n5546 ;
  assign n5548 = n5501 & ~n5546 ;
  assign n5549 = ~n5547 & ~n5548 ;
  assign n5550 = \P4_datao_reg[10]/NET0131  & n4523 ;
  assign n5551 = \P4_datao_reg[11]/NET0131  & n4525 ;
  assign n5552 = ~n5550 & ~n5551 ;
  assign n5553 = n4517 & ~n5552 ;
  assign n5554 = ~n4517 & n5552 ;
  assign n5555 = ~n5553 & ~n5554 ;
  assign n5556 = \P4_datao_reg[20]/NET0131  & n4511 ;
  assign n5557 = \P4_datao_reg[21]/NET0131  & n4507 ;
  assign n5558 = ~n5556 & ~n5557 ;
  assign n5559 = n4431 & ~n5558 ;
  assign n5560 = ~n4431 & n5558 ;
  assign n5561 = ~n5559 & ~n5560 ;
  assign n5562 = \P4_datao_reg[12]/NET0131  & n4388 ;
  assign n5563 = \P4_datao_reg[13]/NET0131  & n4390 ;
  assign n5564 = ~n5562 & ~n5563 ;
  assign n5565 = n4382 & ~n5564 ;
  assign n5566 = ~n4382 & n5564 ;
  assign n5567 = ~n5565 & ~n5566 ;
  assign n5568 = n5561 & n5567 ;
  assign n5569 = ~n5561 & ~n5567 ;
  assign n5570 = ~n5568 & ~n5569 ;
  assign n5571 = n5555 & ~n5570 ;
  assign n5572 = ~n5555 & n5570 ;
  assign n5573 = ~n5571 & ~n5572 ;
  assign n5574 = \P4_datao_reg[16]/NET0131  & n4360 ;
  assign n5575 = \P4_datao_reg[17]/NET0131  & n4356 ;
  assign n5576 = ~n5574 & ~n5575 ;
  assign n5577 = n4351 & ~n5576 ;
  assign n5578 = ~n4351 & n5576 ;
  assign n5579 = ~n5577 & ~n5578 ;
  assign n5580 = \P4_datao_reg[6]/NET0131  & n4566 ;
  assign n5581 = \P4_datao_reg[7]/NET0131  & n4562 ;
  assign n5582 = ~n5580 & ~n5581 ;
  assign n5583 = n4417 & ~n5582 ;
  assign n5584 = ~n4417 & n5582 ;
  assign n5585 = ~n5583 & ~n5584 ;
  assign n5586 = \P4_datao_reg[4]/NET0131  & n4460 ;
  assign n5587 = \P4_datao_reg[5]/NET0131  & n4421 ;
  assign n5588 = ~n5586 & ~n5587 ;
  assign n5589 = n4447 & ~n5588 ;
  assign n5590 = ~n4447 & n5588 ;
  assign n5591 = ~n5589 & ~n5590 ;
  assign n5592 = n5585 & n5591 ;
  assign n5593 = ~n5585 & ~n5591 ;
  assign n5594 = ~n5592 & ~n5593 ;
  assign n5595 = n5579 & ~n5594 ;
  assign n5596 = ~n5579 & n5594 ;
  assign n5597 = ~n5595 & ~n5596 ;
  assign n5598 = ~n5573 & ~n5597 ;
  assign n5599 = n5573 & n5597 ;
  assign n5600 = ~n5598 & ~n5599 ;
  assign n5601 = \P4_datao_reg[24]/NET0131  & n4552 ;
  assign n5602 = \P4_datao_reg[25]/NET0131  & n4548 ;
  assign n5603 = ~n5601 & ~n5602 ;
  assign n5604 = ~n4399 & n5603 ;
  assign n5605 = n4399 & ~n5603 ;
  assign n5606 = ~n5604 & ~n5605 ;
  assign n5607 = \P4_datao_reg[9]/NET0131  & n4575 ;
  assign n5608 = \P4_datao_reg[8]/NET0131  & n4580 ;
  assign n5609 = ~n5607 & ~n5608 ;
  assign n5610 = n4558 & ~n5609 ;
  assign n5611 = ~n4558 & n5609 ;
  assign n5612 = ~n5610 & ~n5611 ;
  assign n5613 = \P4_datao_reg[19]/NET0131  & n4435 ;
  assign n5614 = \P4_datao_reg[18]/NET0131  & n4439 ;
  assign n5615 = ~n5613 & ~n5614 ;
  assign n5616 = n4352 & ~n5615 ;
  assign n5617 = ~n4352 & n5615 ;
  assign n5618 = ~n5616 & ~n5617 ;
  assign n5619 = n5612 & n5618 ;
  assign n5620 = ~n5612 & ~n5618 ;
  assign n5621 = ~n5619 & ~n5620 ;
  assign n5622 = n5606 & ~n5621 ;
  assign n5623 = ~n5606 & n5621 ;
  assign n5624 = ~n5622 & ~n5623 ;
  assign n5625 = n5600 & n5624 ;
  assign n5626 = ~n5600 & ~n5624 ;
  assign n5627 = ~n5625 & ~n5626 ;
  assign n5628 = ~n5421 & ~n5426 ;
  assign n5629 = ~n5420 & ~n5628 ;
  assign n5630 = n5627 & n5629 ;
  assign n5631 = ~n5627 & ~n5629 ;
  assign n5632 = ~n5630 & ~n5631 ;
  assign n5633 = ~n5386 & ~n5390 ;
  assign n5634 = ~n5387 & ~n5633 ;
  assign n5635 = n5632 & ~n5634 ;
  assign n5636 = ~n5632 & n5634 ;
  assign n5637 = ~n5635 & ~n5636 ;
  assign n5638 = n5549 & ~n5637 ;
  assign n5639 = ~n5549 & n5637 ;
  assign n5640 = ~n5638 & ~n5639 ;
  assign n5641 = n5451 & ~n5640 ;
  assign n5642 = ~n5451 & n5640 ;
  assign n5643 = ~n5641 & ~n5642 ;
  assign n5644 = ~n5340 & n5437 ;
  assign n5645 = ~n5339 & ~n5644 ;
  assign n5646 = ~n5643 & n5645 ;
  assign n5647 = ~n5449 & ~n5640 ;
  assign n5648 = ~n5450 & ~n5647 ;
  assign n5649 = ~n5547 & n5637 ;
  assign n5650 = ~n5548 & ~n5649 ;
  assign n5651 = ~n5540 & n5543 ;
  assign n5652 = ~n5539 & ~n5651 ;
  assign n5653 = \P4_datao_reg[24]/NET0131  & n4407 ;
  assign n5654 = \P4_datao_reg[23]/NET0131  & n4405 ;
  assign n5655 = ~n5653 & ~n5654 ;
  assign n5656 = ~n4398 & n5655 ;
  assign n5657 = n4398 & ~n5655 ;
  assign n5658 = ~n5656 & ~n5657 ;
  assign n5659 = \P4_datao_reg[16]/NET0131  & n4376 ;
  assign n5660 = \P4_datao_reg[15]/NET0131  & n4374 ;
  assign n5661 = ~n5659 & ~n5660 ;
  assign n5662 = ~n4368 & n5661 ;
  assign n5663 = n4368 & ~n5661 ;
  assign n5664 = ~n5662 & ~n5663 ;
  assign n5665 = \P4_datao_reg[14]/NET0131  & n4390 ;
  assign n5666 = \P4_datao_reg[13]/NET0131  & n4388 ;
  assign n5667 = ~n5665 & ~n5666 ;
  assign n5668 = ~n4382 & n5667 ;
  assign n5669 = n4382 & ~n5667 ;
  assign n5670 = ~n5668 & ~n5669 ;
  assign n5671 = ~n5664 & ~n5670 ;
  assign n5672 = n5664 & n5670 ;
  assign n5673 = ~n5671 & ~n5672 ;
  assign n5674 = n5658 & n5673 ;
  assign n5675 = ~n5658 & ~n5673 ;
  assign n5676 = ~n5674 & ~n5675 ;
  assign n5677 = \P4_datao_reg[21]/NET0131  & n4511 ;
  assign n5678 = \P4_datao_reg[22]/NET0131  & n4507 ;
  assign n5679 = ~n5677 & ~n5678 ;
  assign n5680 = n4431 & ~n5679 ;
  assign n5681 = ~n4431 & n5679 ;
  assign n5682 = ~n5680 & ~n5681 ;
  assign n5683 = \P4_datao_reg[12]/NET0131  & n4525 ;
  assign n5684 = \P4_datao_reg[11]/NET0131  & n4523 ;
  assign n5685 = ~n5683 & ~n5684 ;
  assign n5686 = n4517 & ~n5685 ;
  assign n5687 = ~n4517 & n5685 ;
  assign n5688 = ~n5686 & ~n5687 ;
  assign n5689 = \P4_datao_reg[10]/NET0131  & n4575 ;
  assign n5690 = \P4_datao_reg[9]/NET0131  & n4580 ;
  assign n5691 = ~n5689 & ~n5690 ;
  assign n5692 = n4558 & ~n5691 ;
  assign n5693 = ~n4558 & n5691 ;
  assign n5694 = ~n5692 & ~n5693 ;
  assign n5695 = n5688 & n5694 ;
  assign n5696 = ~n5688 & ~n5694 ;
  assign n5697 = ~n5695 & ~n5696 ;
  assign n5698 = n5682 & ~n5697 ;
  assign n5699 = ~n5682 & n5697 ;
  assign n5700 = ~n5698 & ~n5699 ;
  assign n5701 = n5676 & ~n5700 ;
  assign n5702 = ~n5676 & n5700 ;
  assign n5703 = ~n5701 & ~n5702 ;
  assign n5704 = n5517 & ~n5534 ;
  assign n5705 = ~n5533 & ~n5704 ;
  assign n5706 = n5703 & n5705 ;
  assign n5707 = ~n5703 & ~n5705 ;
  assign n5708 = ~n5706 & ~n5707 ;
  assign n5709 = ~n5652 & ~n5708 ;
  assign n5710 = n5652 & n5708 ;
  assign n5711 = ~n5709 & ~n5710 ;
  assign n5712 = ~n5495 & ~n5498 ;
  assign n5713 = ~n5494 & ~n5712 ;
  assign n5714 = n5711 & ~n5713 ;
  assign n5715 = ~n5711 & n5713 ;
  assign n5716 = ~n5714 & ~n5715 ;
  assign n5717 = n5650 & ~n5716 ;
  assign n5718 = ~n5650 & n5716 ;
  assign n5719 = ~n5717 & ~n5718 ;
  assign n5720 = ~n5599 & ~n5624 ;
  assign n5721 = ~n5598 & ~n5720 ;
  assign n5722 = ~n5468 & n5490 ;
  assign n5723 = ~n5469 & ~n5722 ;
  assign n5724 = n5721 & n5723 ;
  assign n5725 = ~n5721 & ~n5723 ;
  assign n5726 = ~n5724 & ~n5725 ;
  assign n5728 = \din[30]_pad  & n5483 ;
  assign n5727 = ~\din[29]_pad  & ~\din[30]_pad  ;
  assign n5729 = sel_pad & ~n5727 ;
  assign n5730 = ~n5728 & n5729 ;
  assign n5731 = \P4_datao_reg[0]/NET0131  & n5730 ;
  assign n5732 = \P4_datao_reg[30]/NET0131  & n4343 ;
  assign n5733 = ~\din[1]_pad  & n5732 ;
  assign n5734 = \P4_datao_reg[29]/NET0131  & ~n4343 ;
  assign n5735 = n4329 & ~n5732 ;
  assign n5736 = ~n5734 & n5735 ;
  assign n5737 = ~n5733 & ~n5736 ;
  assign n5738 = n5731 & ~n5737 ;
  assign n5739 = ~n5731 & n5737 ;
  assign n5740 = ~n5738 & ~n5739 ;
  assign n5741 = \P4_datao_reg[28]/NET0131  & n4337 ;
  assign n5742 = \P4_datao_reg[27]/NET0131  & n4335 ;
  assign n5743 = ~n5741 & ~n5742 ;
  assign n5744 = n4328 & ~n5743 ;
  assign n5745 = ~n4328 & n5743 ;
  assign n5746 = ~n5744 & ~n5745 ;
  assign n5747 = ~n5740 & n5746 ;
  assign n5748 = n5740 & ~n5746 ;
  assign n5749 = ~n5747 & ~n5748 ;
  assign n5750 = \P4_datao_reg[17]/NET0131  & n4360 ;
  assign n5751 = \P4_datao_reg[18]/NET0131  & n4356 ;
  assign n5752 = ~n5750 & ~n5751 ;
  assign n5753 = ~n4351 & n5752 ;
  assign n5754 = n4351 & ~n5752 ;
  assign n5755 = ~n5753 & ~n5754 ;
  assign n5756 = \P4_datao_reg[5]/NET0131  & n4460 ;
  assign n5757 = \P4_datao_reg[6]/NET0131  & n4421 ;
  assign n5758 = ~n5756 & ~n5757 ;
  assign n5759 = n4447 & ~n5758 ;
  assign n5760 = ~n4447 & n5758 ;
  assign n5761 = ~n5759 & ~n5760 ;
  assign n5762 = \P4_datao_reg[4]/NET0131  & n4815 ;
  assign n5763 = \P4_datao_reg[3]/NET0131  & n4813 ;
  assign n5764 = ~n5762 & ~n5763 ;
  assign n5765 = n4807 & ~n5764 ;
  assign n5766 = ~n4807 & n5764 ;
  assign n5767 = ~n5765 & ~n5766 ;
  assign n5768 = n5761 & n5767 ;
  assign n5769 = ~n5761 & ~n5767 ;
  assign n5770 = ~n5768 & ~n5769 ;
  assign n5771 = n5755 & ~n5770 ;
  assign n5772 = ~n5755 & n5770 ;
  assign n5773 = ~n5771 & ~n5772 ;
  assign n5774 = n5749 & n5773 ;
  assign n5775 = ~n5749 & ~n5773 ;
  assign n5776 = ~n5774 & ~n5775 ;
  assign n5777 = \P4_datao_reg[8]/NET0131  & n4562 ;
  assign n5778 = \P4_datao_reg[7]/NET0131  & n4566 ;
  assign n5779 = ~n5777 & ~n5778 ;
  assign n5780 = ~n4417 & n5779 ;
  assign n5781 = n4417 & ~n5779 ;
  assign n5782 = ~n5780 & ~n5781 ;
  assign n5783 = \P4_datao_reg[20]/NET0131  & n4435 ;
  assign n5784 = \P4_datao_reg[19]/NET0131  & n4439 ;
  assign n5785 = ~n5783 & ~n5784 ;
  assign n5786 = n4352 & ~n5785 ;
  assign n5787 = ~n4352 & n5785 ;
  assign n5788 = ~n5786 & ~n5787 ;
  assign n5789 = n5782 & n5788 ;
  assign n5790 = ~n5782 & ~n5788 ;
  assign n5791 = ~n5789 & ~n5790 ;
  assign n5792 = \P4_datao_reg[25]/NET0131  & n4552 ;
  assign n5793 = \P4_datao_reg[26]/NET0131  & n4548 ;
  assign n5794 = ~n5792 & ~n5793 ;
  assign n5795 = n4399 & ~n5794 ;
  assign n5796 = ~n4399 & n5794 ;
  assign n5797 = ~n5795 & ~n5796 ;
  assign n5798 = n5791 & n5797 ;
  assign n5799 = ~n5791 & ~n5797 ;
  assign n5800 = ~n5798 & ~n5799 ;
  assign n5801 = n5776 & ~n5800 ;
  assign n5802 = ~n5776 & n5800 ;
  assign n5803 = ~n5801 & ~n5802 ;
  assign n5804 = n5726 & ~n5803 ;
  assign n5805 = ~n5726 & n5803 ;
  assign n5806 = ~n5804 & ~n5805 ;
  assign n5807 = \P4_datao_reg[1]/NET0131  & n5527 ;
  assign n5808 = \P4_datao_reg[2]/NET0131  & n5363 ;
  assign n5809 = ~n5807 & ~n5808 ;
  assign n5810 = ~n5483 & n5809 ;
  assign n5811 = n5483 & ~n5809 ;
  assign n5812 = ~n5810 & ~n5811 ;
  assign n5813 = ~n5515 & ~n5812 ;
  assign n5814 = n5515 & n5812 ;
  assign n5815 = ~n5813 & ~n5814 ;
  assign n5816 = ~n5476 & ~n5486 ;
  assign n5817 = ~n5485 & ~n5816 ;
  assign n5818 = n5815 & ~n5817 ;
  assign n5819 = ~n5815 & n5817 ;
  assign n5820 = ~n5818 & ~n5819 ;
  assign n5821 = ~n5457 & ~n5460 ;
  assign n5822 = ~n5456 & ~n5821 ;
  assign n5823 = ~n5820 & ~n5822 ;
  assign n5824 = n5820 & n5822 ;
  assign n5825 = ~n5823 & ~n5824 ;
  assign n5826 = ~n5579 & ~n5592 ;
  assign n5827 = ~n5593 & ~n5826 ;
  assign n5828 = ~n5606 & ~n5619 ;
  assign n5829 = ~n5620 & ~n5828 ;
  assign n5830 = ~n5555 & ~n5568 ;
  assign n5831 = ~n5569 & ~n5830 ;
  assign n5832 = n5829 & n5831 ;
  assign n5833 = ~n5829 & ~n5831 ;
  assign n5834 = ~n5832 & ~n5833 ;
  assign n5835 = n5827 & ~n5834 ;
  assign n5836 = ~n5827 & n5834 ;
  assign n5837 = ~n5835 & ~n5836 ;
  assign n5838 = n5825 & n5837 ;
  assign n5839 = ~n5825 & ~n5837 ;
  assign n5840 = ~n5838 & ~n5839 ;
  assign n5841 = n5806 & ~n5840 ;
  assign n5842 = ~n5806 & n5840 ;
  assign n5843 = ~n5841 & ~n5842 ;
  assign n5844 = ~n5630 & ~n5634 ;
  assign n5845 = ~n5631 & ~n5844 ;
  assign n5846 = n5843 & ~n5845 ;
  assign n5847 = ~n5843 & n5845 ;
  assign n5848 = ~n5846 & ~n5847 ;
  assign n5849 = n5719 & n5848 ;
  assign n5850 = ~n5719 & ~n5848 ;
  assign n5851 = ~n5849 & ~n5850 ;
  assign n5852 = n5648 & ~n5851 ;
  assign n5853 = ~n5646 & ~n5852 ;
  assign n5854 = n5444 & n5853 ;
  assign n5855 = ~n5103 & ~n5104 ;
  assign n5856 = n5110 & n5855 ;
  assign n5857 = ~n5110 & ~n5855 ;
  assign n5858 = ~n5856 & ~n5857 ;
  assign n5859 = ~n5125 & ~n5126 ;
  assign n5860 = n5132 & n5859 ;
  assign n5861 = ~n5132 & ~n5859 ;
  assign n5862 = ~n5860 & ~n5861 ;
  assign n5863 = n5858 & n5862 ;
  assign n5864 = ~n5858 & ~n5862 ;
  assign n5865 = ~n5863 & ~n5864 ;
  assign n5866 = \P4_datao_reg[18]/NET0131  & n4335 ;
  assign n5867 = \P4_datao_reg[19]/NET0131  & n4337 ;
  assign n5868 = ~n5866 & ~n5867 ;
  assign n5869 = ~n4328 & n5868 ;
  assign n5870 = n4328 & ~n5868 ;
  assign n5871 = ~n5869 & ~n5870 ;
  assign n5872 = \P4_datao_reg[21]/NET0131  & n4343 ;
  assign n5873 = ~\din[1]_pad  & n5872 ;
  assign n5874 = \P4_datao_reg[20]/NET0131  & ~n4343 ;
  assign n5875 = n4329 & ~n5872 ;
  assign n5876 = ~n5874 & n5875 ;
  assign n5877 = ~n5873 & ~n5876 ;
  assign n5878 = n5871 & ~n5877 ;
  assign n5879 = ~n5871 & n5877 ;
  assign n5880 = ~n5878 & ~n5879 ;
  assign n5881 = \P4_datao_reg[9]/NET0131  & n4356 ;
  assign n5882 = \P4_datao_reg[8]/NET0131  & n4360 ;
  assign n5883 = ~n5881 & ~n5882 ;
  assign n5884 = n4351 & ~n5883 ;
  assign n5885 = ~n4351 & n5883 ;
  assign n5886 = ~n5884 & ~n5885 ;
  assign n5887 = ~n5880 & ~n5886 ;
  assign n5888 = n5880 & n5886 ;
  assign n5889 = \P4_datao_reg[5]/NET0131  & n4374 ;
  assign n5890 = \P4_datao_reg[6]/NET0131  & n4376 ;
  assign n5891 = ~n5889 & ~n5890 ;
  assign n5892 = n4368 & ~n5891 ;
  assign n5893 = ~n4368 & n5891 ;
  assign n5894 = ~n5892 & ~n5893 ;
  assign n5895 = \P4_datao_reg[3]/NET0131  & n4388 ;
  assign n5896 = \P4_datao_reg[4]/NET0131  & n4390 ;
  assign n5897 = ~n5895 & ~n5896 ;
  assign n5898 = n4382 & ~n5897 ;
  assign n5899 = ~n4382 & n5897 ;
  assign n5900 = ~n5898 & ~n5899 ;
  assign n5901 = ~n5894 & ~n5900 ;
  assign n5902 = n5894 & n5900 ;
  assign n5903 = \P4_datao_reg[18]/NET0131  & n4337 ;
  assign n5904 = \P4_datao_reg[17]/NET0131  & n4335 ;
  assign n5905 = ~n5903 & ~n5904 ;
  assign n5906 = n4328 & ~n5905 ;
  assign n5907 = ~n4328 & n5905 ;
  assign n5908 = ~n5906 & ~n5907 ;
  assign n5909 = ~n5902 & ~n5908 ;
  assign n5910 = ~n5901 & ~n5909 ;
  assign n5911 = ~n5888 & ~n5910 ;
  assign n5912 = ~n5887 & ~n5911 ;
  assign n5913 = n5865 & ~n5912 ;
  assign n5914 = ~n5865 & n5912 ;
  assign n5915 = ~n5913 & ~n5914 ;
  assign n5916 = \P4_datao_reg[6]/NET0131  & n4374 ;
  assign n5917 = \P4_datao_reg[7]/NET0131  & n4376 ;
  assign n5918 = ~n5916 & ~n5917 ;
  assign n5919 = ~n4368 & n5918 ;
  assign n5920 = n4368 & ~n5918 ;
  assign n5921 = ~n5919 & ~n5920 ;
  assign n5922 = \P4_datao_reg[5]/NET0131  & n4390 ;
  assign n5923 = \P4_datao_reg[4]/NET0131  & n4388 ;
  assign n5924 = ~n5922 & ~n5923 ;
  assign n5925 = n4382 & ~n5924 ;
  assign n5926 = ~n4382 & n5924 ;
  assign n5927 = ~n5925 & ~n5926 ;
  assign n5928 = ~n5921 & ~n5927 ;
  assign n5929 = n5921 & n5927 ;
  assign n5930 = \P4_datao_reg[14]/NET0131  & n4405 ;
  assign n5931 = \P4_datao_reg[15]/NET0131  & n4407 ;
  assign n5932 = ~n5930 & ~n5931 ;
  assign n5933 = ~n4398 & n5932 ;
  assign n5934 = n4398 & ~n5932 ;
  assign n5935 = ~n5933 & ~n5934 ;
  assign n5936 = ~n5929 & ~n5935 ;
  assign n5937 = ~n5928 & ~n5936 ;
  assign n5938 = ~n5198 & ~n5199 ;
  assign n5939 = ~n5205 & n5938 ;
  assign n5940 = n5205 & ~n5938 ;
  assign n5941 = ~n5939 & ~n5940 ;
  assign n5942 = ~n5937 & n5941 ;
  assign n5943 = n5937 & ~n5941 ;
  assign n5944 = ~n5942 & ~n5943 ;
  assign n5945 = ~n5149 & ~n5150 ;
  assign n5946 = ~n5156 & n5945 ;
  assign n5947 = n5156 & ~n5945 ;
  assign n5948 = ~n5946 & ~n5947 ;
  assign n5949 = n5944 & ~n5948 ;
  assign n5950 = ~n5944 & n5948 ;
  assign n5951 = ~n5949 & ~n5950 ;
  assign n5952 = ~n5915 & ~n5951 ;
  assign n5953 = n5915 & n5951 ;
  assign n5954 = ~n5952 & ~n5953 ;
  assign n5955 = \P4_datao_reg[0]/NET0131  & n4525 ;
  assign n5956 = \P4_datao_reg[0]/NET0131  & n4523 ;
  assign n5957 = \P4_datao_reg[1]/NET0131  & n4525 ;
  assign n5958 = ~n5956 & ~n5957 ;
  assign n5959 = n4517 & n5958 ;
  assign n5960 = ~n5955 & n5959 ;
  assign n5961 = \P4_datao_reg[11]/NET0131  & n4507 ;
  assign n5962 = \P4_datao_reg[10]/NET0131  & n4511 ;
  assign n5963 = ~n5961 & ~n5962 ;
  assign n5964 = n4431 & ~n5963 ;
  assign n5965 = ~n4431 & n5963 ;
  assign n5966 = ~n5964 & ~n5965 ;
  assign n5967 = n4517 & n5955 ;
  assign n5968 = ~n5958 & ~n5967 ;
  assign n5969 = ~n5959 & ~n5968 ;
  assign n5970 = n5966 & ~n5969 ;
  assign n5971 = ~n5960 & ~n5970 ;
  assign n5972 = \P4_datao_reg[4]/NET0131  & n4374 ;
  assign n5973 = \P4_datao_reg[5]/NET0131  & n4376 ;
  assign n5974 = ~n5972 & ~n5973 ;
  assign n5975 = n4368 & ~n5974 ;
  assign n5976 = ~n4368 & n5974 ;
  assign n5977 = ~n5975 & ~n5976 ;
  assign n5978 = \P4_datao_reg[3]/NET0131  & n4390 ;
  assign n5979 = \P4_datao_reg[2]/NET0131  & n4388 ;
  assign n5980 = ~n5978 & ~n5979 ;
  assign n5981 = n4382 & ~n5980 ;
  assign n5982 = ~n4382 & n5980 ;
  assign n5983 = ~n5981 & ~n5982 ;
  assign n5984 = ~n5977 & ~n5983 ;
  assign n5985 = n5977 & n5983 ;
  assign n5986 = \P4_datao_reg[13]/NET0131  & n4407 ;
  assign n5987 = \P4_datao_reg[12]/NET0131  & n4405 ;
  assign n5988 = ~n5986 & ~n5987 ;
  assign n5989 = n4398 & ~n5988 ;
  assign n5990 = ~n4398 & n5988 ;
  assign n5991 = ~n5989 & ~n5990 ;
  assign n5992 = ~n5985 & ~n5991 ;
  assign n5993 = ~n5984 & ~n5992 ;
  assign n5994 = n5971 & ~n5993 ;
  assign n5995 = ~n5971 & n5993 ;
  assign n5996 = \P4_datao_reg[14]/NET0131  & n4552 ;
  assign n5997 = \P4_datao_reg[15]/NET0131  & n4548 ;
  assign n5998 = ~n5996 & ~n5997 ;
  assign n5999 = ~n4399 & n5998 ;
  assign n6000 = n4399 & ~n5998 ;
  assign n6001 = ~n5999 & ~n6000 ;
  assign n6002 = \P4_datao_reg[6]/NET0131  & n4360 ;
  assign n6003 = \P4_datao_reg[7]/NET0131  & n4356 ;
  assign n6004 = ~n6002 & ~n6003 ;
  assign n6005 = ~n4351 & n6004 ;
  assign n6006 = n4351 & ~n6004 ;
  assign n6007 = ~n6005 & ~n6006 ;
  assign n6008 = ~n6001 & ~n6007 ;
  assign n6009 = n6001 & n6007 ;
  assign n6010 = \P4_datao_reg[8]/NET0131  & n4439 ;
  assign n6011 = \P4_datao_reg[9]/NET0131  & n4435 ;
  assign n6012 = ~n6010 & ~n6011 ;
  assign n6013 = n4352 & ~n6012 ;
  assign n6014 = ~n4352 & n6012 ;
  assign n6015 = ~n6013 & ~n6014 ;
  assign n6016 = ~n6009 & ~n6015 ;
  assign n6017 = ~n6008 & ~n6016 ;
  assign n6018 = ~n5995 & ~n6017 ;
  assign n6019 = ~n5994 & ~n6018 ;
  assign n6020 = ~n5887 & ~n5888 ;
  assign n6021 = ~n5910 & n6020 ;
  assign n6022 = n5910 & ~n6020 ;
  assign n6023 = ~n6021 & ~n6022 ;
  assign n6024 = n6019 & ~n6023 ;
  assign n6025 = ~n6019 & n6023 ;
  assign n6026 = \P4_datao_reg[0]/NET0131  & n4575 ;
  assign n6027 = \P4_datao_reg[20]/NET0131  & n4343 ;
  assign n6028 = ~\din[1]_pad  & n6027 ;
  assign n6029 = \P4_datao_reg[19]/NET0131  & ~n4343 ;
  assign n6030 = n4329 & ~n6027 ;
  assign n6031 = ~n6029 & n6030 ;
  assign n6032 = ~n6028 & ~n6031 ;
  assign n6033 = n6026 & ~n6032 ;
  assign n6034 = ~n6026 & n6032 ;
  assign n6035 = \P4_datao_reg[14]/NET0131  & n4407 ;
  assign n6036 = \P4_datao_reg[13]/NET0131  & n4405 ;
  assign n6037 = ~n6035 & ~n6036 ;
  assign n6038 = n4398 & ~n6037 ;
  assign n6039 = ~n4398 & n6037 ;
  assign n6040 = ~n6038 & ~n6039 ;
  assign n6041 = ~n6034 & n6040 ;
  assign n6042 = ~n6033 & ~n6041 ;
  assign n6043 = \P4_datao_reg[16]/NET0131  & n4552 ;
  assign n6044 = \P4_datao_reg[17]/NET0131  & n4548 ;
  assign n6045 = ~n6043 & ~n6044 ;
  assign n6046 = ~n4399 & n6045 ;
  assign n6047 = n4399 & ~n6045 ;
  assign n6048 = ~n6046 & ~n6047 ;
  assign n6049 = n4558 & ~n6026 ;
  assign n6050 = \P4_datao_reg[11]/NET0131  & n4435 ;
  assign n6051 = \P4_datao_reg[10]/NET0131  & n4439 ;
  assign n6052 = ~n6050 & ~n6051 ;
  assign n6053 = n4352 & ~n6052 ;
  assign n6054 = ~n4352 & n6052 ;
  assign n6055 = ~n6053 & ~n6054 ;
  assign n6056 = n6049 & n6055 ;
  assign n6057 = ~n6049 & ~n6055 ;
  assign n6058 = ~n6056 & ~n6057 ;
  assign n6059 = n6048 & n6058 ;
  assign n6060 = ~n6048 & ~n6058 ;
  assign n6061 = ~n6059 & ~n6060 ;
  assign n6062 = n6042 & ~n6061 ;
  assign n6063 = ~n6042 & n6061 ;
  assign n6064 = ~n6062 & ~n6063 ;
  assign n6065 = \P4_datao_reg[1]/NET0131  & n4523 ;
  assign n6066 = \P4_datao_reg[2]/NET0131  & n4525 ;
  assign n6067 = ~n6065 & ~n6066 ;
  assign n6068 = ~n4517 & n6067 ;
  assign n6069 = n4517 & ~n6067 ;
  assign n6070 = ~n6068 & ~n6069 ;
  assign n6071 = \P4_datao_reg[15]/NET0131  & n4552 ;
  assign n6072 = \P4_datao_reg[16]/NET0131  & n4548 ;
  assign n6073 = ~n6071 & ~n6072 ;
  assign n6074 = ~n4399 & n6073 ;
  assign n6075 = n4399 & ~n6073 ;
  assign n6076 = ~n6074 & ~n6075 ;
  assign n6077 = n6070 & n6076 ;
  assign n6078 = ~n6070 & ~n6076 ;
  assign n6079 = \P4_datao_reg[12]/NET0131  & n4507 ;
  assign n6080 = \P4_datao_reg[11]/NET0131  & n4511 ;
  assign n6081 = ~n6079 & ~n6080 ;
  assign n6082 = n4431 & ~n6081 ;
  assign n6083 = ~n4431 & n6081 ;
  assign n6084 = ~n6082 & ~n6083 ;
  assign n6085 = ~n6078 & n6084 ;
  assign n6086 = ~n6077 & ~n6085 ;
  assign n6087 = n6064 & ~n6086 ;
  assign n6088 = ~n6064 & n6086 ;
  assign n6089 = ~n6087 & ~n6088 ;
  assign n6090 = ~n6025 & n6089 ;
  assign n6091 = ~n6024 & ~n6090 ;
  assign n6092 = n5954 & ~n6091 ;
  assign n6093 = ~n5954 & n6091 ;
  assign n6094 = ~n6092 & ~n6093 ;
  assign n6095 = ~n6048 & ~n6056 ;
  assign n6096 = ~n6057 & ~n6095 ;
  assign n6097 = n5878 & n6096 ;
  assign n6098 = ~n5878 & ~n6096 ;
  assign n6099 = ~n6097 & ~n6098 ;
  assign n6100 = \P4_datao_reg[2]/NET0131  & n4523 ;
  assign n6101 = \P4_datao_reg[3]/NET0131  & n4525 ;
  assign n6102 = ~n6100 & ~n6101 ;
  assign n6103 = ~n4517 & n6102 ;
  assign n6104 = n4517 & ~n6102 ;
  assign n6105 = ~n6103 & ~n6104 ;
  assign n6106 = \P4_datao_reg[1]/NET0131  & n4575 ;
  assign n6107 = \P4_datao_reg[0]/NET0131  & n4580 ;
  assign n6108 = ~n6106 & ~n6107 ;
  assign n6109 = n4558 & ~n6108 ;
  assign n6110 = ~n4558 & n6108 ;
  assign n6111 = ~n6109 & ~n6110 ;
  assign n6112 = n6105 & n6111 ;
  assign n6113 = ~n6105 & ~n6111 ;
  assign n6114 = \P4_datao_reg[12]/NET0131  & n4511 ;
  assign n6115 = \P4_datao_reg[13]/NET0131  & n4507 ;
  assign n6116 = ~n6114 & ~n6115 ;
  assign n6117 = ~n4431 & n6116 ;
  assign n6118 = n4431 & ~n6116 ;
  assign n6119 = ~n6117 & ~n6118 ;
  assign n6120 = ~n6113 & n6119 ;
  assign n6121 = ~n6112 & ~n6120 ;
  assign n6122 = n6099 & ~n6121 ;
  assign n6123 = ~n6099 & n6121 ;
  assign n6124 = ~n6122 & ~n6123 ;
  assign n6125 = ~n6063 & n6086 ;
  assign n6126 = ~n6062 & ~n6125 ;
  assign n6127 = ~n6124 & ~n6126 ;
  assign n6128 = n6124 & n6126 ;
  assign n6129 = ~n6127 & ~n6128 ;
  assign n6130 = \P4_datao_reg[9]/NET0131  & n4439 ;
  assign n6131 = \P4_datao_reg[10]/NET0131  & n4435 ;
  assign n6132 = ~n6130 & ~n6131 ;
  assign n6133 = n4352 & ~n6132 ;
  assign n6134 = ~n4352 & n6132 ;
  assign n6135 = ~n6133 & ~n6134 ;
  assign n6136 = \P4_datao_reg[7]/NET0131  & n4360 ;
  assign n6137 = \P4_datao_reg[8]/NET0131  & n4356 ;
  assign n6138 = ~n6136 & ~n6137 ;
  assign n6139 = n4351 & ~n6138 ;
  assign n6140 = ~n4351 & n6138 ;
  assign n6141 = ~n6139 & ~n6140 ;
  assign n6142 = ~n6135 & ~n6141 ;
  assign n6143 = \P4_datao_reg[17]/NET0131  & n4337 ;
  assign n6144 = \P4_datao_reg[16]/NET0131  & n4335 ;
  assign n6145 = ~n6143 & ~n6144 ;
  assign n6146 = n4328 & ~n6145 ;
  assign n6147 = ~n4328 & n6145 ;
  assign n6148 = ~n6146 & ~n6147 ;
  assign n6149 = \P4_datao_reg[19]/NET0131  & n4343 ;
  assign n6150 = ~\din[1]_pad  & n6149 ;
  assign n6151 = \P4_datao_reg[18]/NET0131  & ~n4343 ;
  assign n6152 = n4329 & ~n6149 ;
  assign n6153 = ~n6151 & n6152 ;
  assign n6154 = ~n6150 & ~n6153 ;
  assign n6155 = n6148 & ~n6154 ;
  assign n6156 = n6135 & n6141 ;
  assign n6157 = ~n6155 & ~n6156 ;
  assign n6158 = ~n6142 & ~n6157 ;
  assign n6159 = ~n6112 & ~n6113 ;
  assign n6160 = n6119 & n6159 ;
  assign n6161 = ~n6119 & ~n6159 ;
  assign n6162 = ~n6160 & ~n6161 ;
  assign n6163 = ~n6158 & ~n6162 ;
  assign n6164 = n6158 & n6162 ;
  assign n6165 = ~n5928 & ~n5929 ;
  assign n6166 = n5935 & n6165 ;
  assign n6167 = ~n5935 & ~n6165 ;
  assign n6168 = ~n6166 & ~n6167 ;
  assign n6169 = ~n6164 & ~n6168 ;
  assign n6170 = ~n6163 & ~n6169 ;
  assign n6171 = n6129 & ~n6170 ;
  assign n6172 = ~n6129 & n6170 ;
  assign n6173 = ~n6171 & ~n6172 ;
  assign n6174 = n6094 & ~n6173 ;
  assign n6175 = ~n6094 & n6173 ;
  assign n6176 = ~n6033 & ~n6034 ;
  assign n6177 = n6040 & n6176 ;
  assign n6178 = ~n6040 & ~n6176 ;
  assign n6179 = ~n6177 & ~n6178 ;
  assign n6180 = ~n5901 & ~n5902 ;
  assign n6181 = n5908 & n6180 ;
  assign n6182 = ~n5908 & ~n6180 ;
  assign n6183 = ~n6181 & ~n6182 ;
  assign n6184 = ~n6179 & ~n6183 ;
  assign n6185 = n6179 & n6183 ;
  assign n6186 = ~n6077 & ~n6078 ;
  assign n6187 = ~n6084 & n6186 ;
  assign n6188 = n6084 & ~n6186 ;
  assign n6189 = ~n6187 & ~n6188 ;
  assign n6190 = ~n6185 & n6189 ;
  assign n6191 = ~n6184 & ~n6190 ;
  assign n6192 = ~n6163 & ~n6164 ;
  assign n6193 = ~n6168 & n6192 ;
  assign n6194 = n6168 & ~n6192 ;
  assign n6195 = ~n6193 & ~n6194 ;
  assign n6196 = n6191 & ~n6195 ;
  assign n6197 = ~n6191 & n6195 ;
  assign n6198 = ~n6024 & ~n6025 ;
  assign n6199 = n6089 & n6198 ;
  assign n6200 = ~n6089 & ~n6198 ;
  assign n6201 = ~n6199 & ~n6200 ;
  assign n6202 = ~n6197 & n6201 ;
  assign n6203 = ~n6196 & ~n6202 ;
  assign n6204 = ~n6175 & ~n6203 ;
  assign n6205 = ~n6174 & ~n6204 ;
  assign n6206 = ~n5953 & ~n6091 ;
  assign n6207 = ~n5952 & ~n6206 ;
  assign n6208 = ~n6128 & ~n6170 ;
  assign n6209 = ~n6127 & ~n6208 ;
  assign n6210 = ~n6207 & n6209 ;
  assign n6211 = n6207 & ~n6209 ;
  assign n6212 = ~n6210 & ~n6211 ;
  assign n6213 = ~n5863 & ~n5912 ;
  assign n6214 = ~n5864 & ~n6213 ;
  assign n6215 = ~n5168 & ~n5169 ;
  assign n6216 = n5171 & n6215 ;
  assign n6217 = ~n5171 & ~n6215 ;
  assign n6218 = ~n6216 & ~n6217 ;
  assign n6219 = ~n4396 & ~n4397 ;
  assign n6220 = n4412 & n6219 ;
  assign n6221 = ~n4412 & ~n6219 ;
  assign n6222 = ~n6220 & ~n6221 ;
  assign n6223 = n6218 & n6222 ;
  assign n6224 = ~n6218 & ~n6222 ;
  assign n6225 = ~n6223 & ~n6224 ;
  assign n6226 = ~n6098 & ~n6121 ;
  assign n6227 = ~n6097 & ~n6226 ;
  assign n6228 = n6225 & ~n6227 ;
  assign n6229 = ~n6225 & n6227 ;
  assign n6230 = ~n6228 & ~n6229 ;
  assign n6231 = n6214 & n6230 ;
  assign n6232 = ~n6214 & ~n6230 ;
  assign n6233 = ~n6231 & ~n6232 ;
  assign n6234 = ~n5942 & n5948 ;
  assign n6235 = ~n5943 & ~n6234 ;
  assign n6236 = ~n5135 & ~n5136 ;
  assign n6237 = ~n5158 & n6236 ;
  assign n6238 = n5158 & ~n6236 ;
  assign n6239 = ~n6237 & ~n6238 ;
  assign n6240 = n6235 & ~n6239 ;
  assign n6241 = ~n6235 & n6239 ;
  assign n6242 = ~n6240 & ~n6241 ;
  assign n6243 = ~n5212 & ~n5213 ;
  assign n6244 = ~n5217 & n6243 ;
  assign n6245 = n5217 & ~n6243 ;
  assign n6246 = ~n6244 & ~n6245 ;
  assign n6247 = n6242 & n6246 ;
  assign n6248 = ~n6242 & ~n6246 ;
  assign n6249 = ~n6247 & ~n6248 ;
  assign n6250 = n6233 & n6249 ;
  assign n6251 = ~n6233 & ~n6249 ;
  assign n6252 = ~n6250 & ~n6251 ;
  assign n6253 = n6212 & ~n6252 ;
  assign n6254 = ~n6212 & n6252 ;
  assign n6255 = ~n6253 & ~n6254 ;
  assign n6256 = n6205 & ~n6255 ;
  assign n6257 = ~n6211 & ~n6252 ;
  assign n6258 = ~n6210 & ~n6257 ;
  assign n6259 = ~n5174 & ~n5175 ;
  assign n6260 = ~n5179 & n6259 ;
  assign n6261 = n5179 & ~n6259 ;
  assign n6262 = ~n6260 & ~n6261 ;
  assign n6263 = ~n6223 & n6227 ;
  assign n6264 = ~n6224 & ~n6263 ;
  assign n6265 = n6262 & n6264 ;
  assign n6266 = ~n6262 & ~n6264 ;
  assign n6267 = ~n6265 & ~n6266 ;
  assign n6268 = ~n6240 & ~n6246 ;
  assign n6269 = ~n6241 & ~n6268 ;
  assign n6270 = n6267 & ~n6269 ;
  assign n6271 = ~n6267 & n6269 ;
  assign n6272 = ~n6270 & ~n6271 ;
  assign n6273 = ~n5220 & ~n5221 ;
  assign n6274 = ~n5225 & n6273 ;
  assign n6275 = n5225 & ~n6273 ;
  assign n6276 = ~n6274 & ~n6275 ;
  assign n6277 = n6272 & n6276 ;
  assign n6278 = ~n6272 & ~n6276 ;
  assign n6279 = ~n6277 & ~n6278 ;
  assign n6280 = ~n6232 & ~n6249 ;
  assign n6281 = ~n6231 & ~n6280 ;
  assign n6282 = n6279 & n6281 ;
  assign n6283 = ~n6279 & ~n6281 ;
  assign n6284 = ~n6282 & ~n6283 ;
  assign n6285 = n6258 & n6284 ;
  assign n6286 = ~n6256 & ~n6285 ;
  assign n6287 = ~n6265 & n6269 ;
  assign n6288 = ~n6266 & ~n6287 ;
  assign n6289 = ~n4761 & ~n4762 ;
  assign n6290 = n4766 & n6289 ;
  assign n6291 = ~n4766 & ~n6289 ;
  assign n6292 = ~n6290 & ~n6291 ;
  assign n6293 = n6288 & n6292 ;
  assign n6294 = ~n6288 & ~n6292 ;
  assign n6295 = ~n6293 & ~n6294 ;
  assign n6296 = ~n5228 & ~n5229 ;
  assign n6297 = ~n5233 & n6296 ;
  assign n6298 = n5233 & ~n6296 ;
  assign n6299 = ~n6297 & ~n6298 ;
  assign n6300 = n6295 & ~n6299 ;
  assign n6301 = ~n6295 & n6299 ;
  assign n6302 = ~n6300 & ~n6301 ;
  assign n6303 = ~n6278 & ~n6281 ;
  assign n6304 = ~n6277 & ~n6303 ;
  assign n6305 = n6302 & n6304 ;
  assign n6306 = ~n6293 & ~n6299 ;
  assign n6307 = ~n6294 & ~n6306 ;
  assign n6308 = ~n5240 & ~n5241 ;
  assign n6309 = n5245 & n6308 ;
  assign n6310 = ~n5245 & ~n6308 ;
  assign n6311 = ~n6309 & ~n6310 ;
  assign n6312 = ~n6307 & ~n6311 ;
  assign n6313 = ~n6305 & ~n6312 ;
  assign n6314 = n6286 & n6313 ;
  assign n6315 = \P4_datao_reg[6]/NET0131  & n4439 ;
  assign n6316 = \P4_datao_reg[7]/NET0131  & n4435 ;
  assign n6317 = ~n6315 & ~n6316 ;
  assign n6318 = ~n4352 & n6317 ;
  assign n6319 = n4352 & ~n6317 ;
  assign n6320 = ~n6318 & ~n6319 ;
  assign n6321 = \P4_datao_reg[5]/NET0131  & n4356 ;
  assign n6322 = \P4_datao_reg[4]/NET0131  & n4360 ;
  assign n6323 = ~n6321 & ~n6322 ;
  assign n6324 = n4351 & ~n6323 ;
  assign n6325 = ~n4351 & n6323 ;
  assign n6326 = ~n6324 & ~n6325 ;
  assign n6327 = n6320 & n6326 ;
  assign n6328 = ~n6320 & ~n6326 ;
  assign n6329 = \P4_datao_reg[14]/NET0131  & n4335 ;
  assign n6330 = \P4_datao_reg[15]/NET0131  & n4337 ;
  assign n6331 = ~n6329 & ~n6330 ;
  assign n6332 = ~n4328 & n6331 ;
  assign n6333 = n4328 & ~n6331 ;
  assign n6334 = ~n6332 & ~n6333 ;
  assign n6335 = \P4_datao_reg[17]/NET0131  & n4343 ;
  assign n6336 = ~\din[1]_pad  & n6335 ;
  assign n6337 = \P4_datao_reg[16]/NET0131  & ~n4343 ;
  assign n6338 = n4329 & ~n6335 ;
  assign n6339 = ~n6337 & n6338 ;
  assign n6340 = ~n6336 & ~n6339 ;
  assign n6341 = n6334 & ~n6340 ;
  assign n6342 = ~n6334 & n6340 ;
  assign n6343 = ~n6341 & ~n6342 ;
  assign n6344 = ~n6328 & n6343 ;
  assign n6345 = ~n6327 & ~n6344 ;
  assign n6346 = \P4_datao_reg[15]/NET0131  & n4335 ;
  assign n6347 = \P4_datao_reg[16]/NET0131  & n4337 ;
  assign n6348 = ~n6346 & ~n6347 ;
  assign n6349 = ~n4328 & n6348 ;
  assign n6350 = n4328 & ~n6348 ;
  assign n6351 = ~n6349 & ~n6350 ;
  assign n6352 = \P4_datao_reg[14]/NET0131  & n4548 ;
  assign n6353 = \P4_datao_reg[13]/NET0131  & n4552 ;
  assign n6354 = ~n6352 & ~n6353 ;
  assign n6355 = n4399 & ~n6354 ;
  assign n6356 = ~n4399 & n6354 ;
  assign n6357 = ~n6355 & ~n6356 ;
  assign n6358 = \P4_datao_reg[8]/NET0131  & n4435 ;
  assign n6359 = \P4_datao_reg[7]/NET0131  & n4439 ;
  assign n6360 = ~n6358 & ~n6359 ;
  assign n6361 = n4352 & ~n6360 ;
  assign n6362 = ~n4352 & n6360 ;
  assign n6363 = ~n6361 & ~n6362 ;
  assign n6364 = ~n6357 & ~n6363 ;
  assign n6365 = n6357 & n6363 ;
  assign n6366 = ~n6364 & ~n6365 ;
  assign n6367 = n6351 & ~n6366 ;
  assign n6368 = ~n6351 & n6366 ;
  assign n6369 = ~n6367 & ~n6368 ;
  assign n6370 = ~n6345 & ~n6369 ;
  assign n6371 = n6345 & n6369 ;
  assign n6372 = \P4_datao_reg[4]/NET0131  & n4356 ;
  assign n6373 = \P4_datao_reg[3]/NET0131  & n4360 ;
  assign n6374 = ~n6372 & ~n6373 ;
  assign n6375 = n4351 & ~n6374 ;
  assign n6376 = ~n4351 & n6374 ;
  assign n6377 = ~n6375 & ~n6376 ;
  assign n6378 = \P4_datao_reg[6]/NET0131  & n4435 ;
  assign n6379 = \P4_datao_reg[5]/NET0131  & n4439 ;
  assign n6380 = ~n6378 & ~n6379 ;
  assign n6381 = n4352 & ~n6380 ;
  assign n6382 = ~n4352 & n6380 ;
  assign n6383 = ~n6381 & ~n6382 ;
  assign n6384 = \P4_datao_reg[12]/NET0131  & n4548 ;
  assign n6385 = \P4_datao_reg[11]/NET0131  & n4552 ;
  assign n6386 = ~n6384 & ~n6385 ;
  assign n6387 = n4399 & ~n6386 ;
  assign n6388 = ~n4399 & n6386 ;
  assign n6389 = ~n6387 & ~n6388 ;
  assign n6390 = n6383 & n6389 ;
  assign n6391 = ~n6377 & ~n6390 ;
  assign n6392 = ~n6383 & ~n6389 ;
  assign n6393 = ~n6391 & ~n6392 ;
  assign n6394 = \P4_datao_reg[2]/NET0131  & n4376 ;
  assign n6395 = \P4_datao_reg[1]/NET0131  & n4374 ;
  assign n6396 = ~n6394 & ~n6395 ;
  assign n6397 = n4368 & ~n6396 ;
  assign n6398 = ~n4368 & n6396 ;
  assign n6399 = ~n6397 & ~n6398 ;
  assign n6400 = \P4_datao_reg[10]/NET0131  & n4407 ;
  assign n6401 = \P4_datao_reg[9]/NET0131  & n4405 ;
  assign n6402 = ~n6400 & ~n6401 ;
  assign n6403 = n4398 & ~n6402 ;
  assign n6404 = ~n4398 & n6402 ;
  assign n6405 = ~n6403 & ~n6404 ;
  assign n6406 = n6399 & n6405 ;
  assign n6407 = ~n6399 & ~n6405 ;
  assign n6408 = \P4_datao_reg[14]/NET0131  & n4337 ;
  assign n6409 = \P4_datao_reg[13]/NET0131  & n4335 ;
  assign n6410 = ~n6408 & ~n6409 ;
  assign n6411 = n4328 & ~n6410 ;
  assign n6412 = ~n4328 & n6410 ;
  assign n6413 = ~n6411 & ~n6412 ;
  assign n6414 = ~n6407 & n6413 ;
  assign n6415 = ~n6406 & ~n6414 ;
  assign n6416 = n6393 & ~n6415 ;
  assign n6417 = ~n6393 & n6415 ;
  assign n6418 = \P4_datao_reg[0]/NET0131  & n4390 ;
  assign n6419 = \P4_datao_reg[16]/NET0131  & n4343 ;
  assign n6420 = ~\din[1]_pad  & n6419 ;
  assign n6421 = \P4_datao_reg[15]/NET0131  & ~n4343 ;
  assign n6422 = n4329 & ~n6419 ;
  assign n6423 = ~n6421 & n6422 ;
  assign n6424 = ~n6420 & ~n6423 ;
  assign n6425 = n6418 & ~n6424 ;
  assign n6426 = ~n6418 & n6424 ;
  assign n6427 = \P4_datao_reg[8]/NET0131  & n4507 ;
  assign n6428 = \P4_datao_reg[7]/NET0131  & n4511 ;
  assign n6429 = ~n6427 & ~n6428 ;
  assign n6430 = n4431 & ~n6429 ;
  assign n6431 = ~n4431 & n6429 ;
  assign n6432 = ~n6430 & ~n6431 ;
  assign n6433 = ~n6426 & n6432 ;
  assign n6434 = ~n6425 & ~n6433 ;
  assign n6435 = ~n6417 & ~n6434 ;
  assign n6436 = ~n6416 & ~n6435 ;
  assign n6437 = ~n6371 & ~n6436 ;
  assign n6438 = ~n6370 & ~n6437 ;
  assign n6439 = \P4_datao_reg[2]/NET0131  & n4374 ;
  assign n6440 = \P4_datao_reg[3]/NET0131  & n4376 ;
  assign n6441 = ~n6439 & ~n6440 ;
  assign n6442 = ~n4368 & n6441 ;
  assign n6443 = n4368 & ~n6441 ;
  assign n6444 = ~n6442 & ~n6443 ;
  assign n6445 = \P4_datao_reg[0]/NET0131  & n4388 ;
  assign n6446 = \P4_datao_reg[1]/NET0131  & n4390 ;
  assign n6447 = ~n6445 & ~n6446 ;
  assign n6448 = ~n4382 & n6447 ;
  assign n6449 = n4382 & ~n6447 ;
  assign n6450 = ~n6448 & ~n6449 ;
  assign n6451 = n6444 & n6450 ;
  assign n6452 = ~n6444 & ~n6450 ;
  assign n6453 = \P4_datao_reg[11]/NET0131  & n4407 ;
  assign n6454 = \P4_datao_reg[10]/NET0131  & n4405 ;
  assign n6455 = ~n6453 & ~n6454 ;
  assign n6456 = n4398 & ~n6455 ;
  assign n6457 = ~n4398 & n6455 ;
  assign n6458 = ~n6456 & ~n6457 ;
  assign n6459 = ~n6452 & n6458 ;
  assign n6460 = ~n6451 & ~n6459 ;
  assign n6461 = \P4_datao_reg[10]/NET0131  & n4507 ;
  assign n6462 = \P4_datao_reg[9]/NET0131  & n4511 ;
  assign n6463 = ~n6461 & ~n6462 ;
  assign n6464 = n4431 & ~n6463 ;
  assign n6465 = ~n4431 & n6463 ;
  assign n6466 = ~n6464 & ~n6465 ;
  assign n6467 = \P4_datao_reg[18]/NET0131  & n4343 ;
  assign n6468 = ~\din[1]_pad  & n6467 ;
  assign n6469 = \P4_datao_reg[17]/NET0131  & ~n4343 ;
  assign n6470 = n4329 & ~n6467 ;
  assign n6471 = ~n6469 & n6470 ;
  assign n6472 = ~n6468 & ~n6471 ;
  assign n6473 = n5955 & ~n6472 ;
  assign n6474 = ~n5955 & n6472 ;
  assign n6475 = ~n6473 & ~n6474 ;
  assign n6476 = n6466 & ~n6475 ;
  assign n6477 = ~n6466 & n6475 ;
  assign n6478 = ~n6476 & ~n6477 ;
  assign n6479 = ~n6460 & ~n6478 ;
  assign n6480 = n6460 & n6478 ;
  assign n6481 = \P4_datao_reg[11]/NET0131  & n4405 ;
  assign n6482 = \P4_datao_reg[12]/NET0131  & n4407 ;
  assign n6483 = ~n6481 & ~n6482 ;
  assign n6484 = ~n4398 & n6483 ;
  assign n6485 = n4398 & ~n6483 ;
  assign n6486 = ~n6484 & ~n6485 ;
  assign n6487 = \P4_datao_reg[1]/NET0131  & n4388 ;
  assign n6488 = \P4_datao_reg[2]/NET0131  & n4390 ;
  assign n6489 = ~n6487 & ~n6488 ;
  assign n6490 = ~n4382 & n6489 ;
  assign n6491 = n4382 & ~n6489 ;
  assign n6492 = ~n6490 & ~n6491 ;
  assign n6493 = \P4_datao_reg[4]/NET0131  & n4376 ;
  assign n6494 = \P4_datao_reg[3]/NET0131  & n4374 ;
  assign n6495 = ~n6493 & ~n6494 ;
  assign n6496 = n4368 & ~n6495 ;
  assign n6497 = ~n4368 & n6495 ;
  assign n6498 = ~n6496 & ~n6497 ;
  assign n6499 = ~n6492 & ~n6498 ;
  assign n6500 = n6492 & n6498 ;
  assign n6501 = ~n6499 & ~n6500 ;
  assign n6502 = n6486 & n6501 ;
  assign n6503 = ~n6486 & ~n6501 ;
  assign n6504 = ~n6502 & ~n6503 ;
  assign n6505 = ~n6480 & n6504 ;
  assign n6506 = ~n6479 & ~n6505 ;
  assign n6507 = ~n6438 & ~n6506 ;
  assign n6508 = n6438 & n6506 ;
  assign n6509 = ~n6351 & ~n6365 ;
  assign n6510 = ~n6364 & ~n6509 ;
  assign n6511 = ~n6008 & ~n6009 ;
  assign n6512 = ~n6015 & n6511 ;
  assign n6513 = n6015 & ~n6511 ;
  assign n6514 = ~n6512 & ~n6513 ;
  assign n6515 = n6510 & ~n6514 ;
  assign n6516 = ~n6510 & n6514 ;
  assign n6517 = ~n6515 & ~n6516 ;
  assign n6518 = ~n5984 & ~n5985 ;
  assign n6519 = ~n5991 & n6518 ;
  assign n6520 = n5991 & ~n6518 ;
  assign n6521 = ~n6519 & ~n6520 ;
  assign n6522 = n6517 & ~n6521 ;
  assign n6523 = ~n6517 & n6521 ;
  assign n6524 = ~n6522 & ~n6523 ;
  assign n6525 = ~n6508 & n6524 ;
  assign n6526 = ~n6507 & ~n6525 ;
  assign n6527 = \P4_datao_reg[6]/NET0131  & n4356 ;
  assign n6528 = \P4_datao_reg[5]/NET0131  & n4360 ;
  assign n6529 = ~n6527 & ~n6528 ;
  assign n6530 = n4351 & ~n6529 ;
  assign n6531 = ~n4351 & n6529 ;
  assign n6532 = ~n6530 & ~n6531 ;
  assign n6533 = n6341 & n6532 ;
  assign n6534 = ~n6341 & ~n6532 ;
  assign n6535 = \P4_datao_reg[12]/NET0131  & n4552 ;
  assign n6536 = \P4_datao_reg[13]/NET0131  & n4548 ;
  assign n6537 = ~n6535 & ~n6536 ;
  assign n6538 = ~n4399 & n6537 ;
  assign n6539 = n4399 & ~n6537 ;
  assign n6540 = ~n6538 & ~n6539 ;
  assign n6541 = n4382 & ~n6418 ;
  assign n6542 = n6540 & n6541 ;
  assign n6543 = ~n6540 & ~n6541 ;
  assign n6544 = \P4_datao_reg[9]/NET0131  & n4507 ;
  assign n6545 = \P4_datao_reg[8]/NET0131  & n4511 ;
  assign n6546 = ~n6544 & ~n6545 ;
  assign n6547 = n4431 & ~n6546 ;
  assign n6548 = ~n4431 & n6546 ;
  assign n6549 = ~n6547 & ~n6548 ;
  assign n6550 = ~n6543 & n6549 ;
  assign n6551 = ~n6542 & ~n6550 ;
  assign n6552 = ~n6534 & ~n6551 ;
  assign n6553 = ~n6533 & ~n6552 ;
  assign n6554 = ~n5960 & ~n5969 ;
  assign n6555 = n5966 & ~n6554 ;
  assign n6556 = ~n5966 & n6554 ;
  assign n6557 = ~n6555 & ~n6556 ;
  assign n6558 = ~n6553 & ~n6557 ;
  assign n6559 = n6553 & n6557 ;
  assign n6560 = ~n6148 & n6154 ;
  assign n6561 = ~n6155 & ~n6560 ;
  assign n6562 = ~n6486 & ~n6500 ;
  assign n6563 = ~n6499 & ~n6562 ;
  assign n6564 = n6561 & n6563 ;
  assign n6565 = ~n6561 & ~n6563 ;
  assign n6566 = ~n6564 & ~n6565 ;
  assign n6567 = n6466 & ~n6474 ;
  assign n6568 = ~n6473 & ~n6567 ;
  assign n6569 = n6566 & ~n6568 ;
  assign n6570 = ~n6566 & n6568 ;
  assign n6571 = ~n6569 & ~n6570 ;
  assign n6572 = ~n6559 & n6571 ;
  assign n6573 = ~n6558 & ~n6572 ;
  assign n6574 = ~n6526 & ~n6573 ;
  assign n6575 = n6526 & n6573 ;
  assign n6576 = ~n6184 & ~n6185 ;
  assign n6577 = n6189 & n6576 ;
  assign n6578 = ~n6189 & ~n6576 ;
  assign n6579 = ~n6577 & ~n6578 ;
  assign n6580 = ~n6516 & ~n6521 ;
  assign n6581 = ~n6515 & ~n6580 ;
  assign n6582 = n6579 & n6581 ;
  assign n6583 = ~n6579 & ~n6581 ;
  assign n6584 = ~n6582 & ~n6583 ;
  assign n6585 = ~n6565 & ~n6568 ;
  assign n6586 = ~n6564 & ~n6585 ;
  assign n6587 = ~n6142 & ~n6156 ;
  assign n6588 = ~n6155 & n6587 ;
  assign n6589 = n6155 & ~n6587 ;
  assign n6590 = ~n6588 & ~n6589 ;
  assign n6591 = ~n6586 & ~n6590 ;
  assign n6592 = n6586 & n6590 ;
  assign n6593 = ~n6591 & ~n6592 ;
  assign n6594 = ~n5994 & ~n5995 ;
  assign n6595 = ~n6017 & n6594 ;
  assign n6596 = n6017 & ~n6594 ;
  assign n6597 = ~n6595 & ~n6596 ;
  assign n6598 = n6593 & n6597 ;
  assign n6599 = ~n6593 & ~n6597 ;
  assign n6600 = ~n6598 & ~n6599 ;
  assign n6601 = n6584 & n6600 ;
  assign n6602 = ~n6584 & ~n6600 ;
  assign n6603 = ~n6601 & ~n6602 ;
  assign n6604 = ~n6575 & ~n6603 ;
  assign n6605 = ~n6574 & ~n6604 ;
  assign n6606 = ~n6592 & ~n6597 ;
  assign n6607 = ~n6591 & ~n6606 ;
  assign n6608 = ~n6196 & ~n6197 ;
  assign n6609 = n6201 & n6608 ;
  assign n6610 = ~n6201 & ~n6608 ;
  assign n6611 = ~n6609 & ~n6610 ;
  assign n6612 = ~n6607 & n6611 ;
  assign n6613 = n6607 & ~n6611 ;
  assign n6614 = ~n6612 & ~n6613 ;
  assign n6615 = ~n6582 & ~n6600 ;
  assign n6616 = ~n6583 & ~n6615 ;
  assign n6617 = n6614 & n6616 ;
  assign n6618 = ~n6614 & ~n6616 ;
  assign n6619 = ~n6617 & ~n6618 ;
  assign n6620 = n6605 & n6619 ;
  assign n6621 = ~n6174 & ~n6175 ;
  assign n6622 = ~n6203 & n6621 ;
  assign n6623 = n6203 & ~n6621 ;
  assign n6624 = ~n6622 & ~n6623 ;
  assign n6625 = ~n6613 & ~n6616 ;
  assign n6626 = ~n6612 & ~n6625 ;
  assign n6627 = ~n6624 & n6626 ;
  assign n6628 = ~n6620 & ~n6627 ;
  assign n6629 = ~n6574 & ~n6575 ;
  assign n6630 = ~n6603 & n6629 ;
  assign n6631 = n6603 & ~n6629 ;
  assign n6632 = ~n6630 & ~n6631 ;
  assign n6633 = ~n6327 & ~n6328 ;
  assign n6634 = ~n6343 & n6633 ;
  assign n6635 = n6343 & ~n6633 ;
  assign n6636 = ~n6634 & ~n6635 ;
  assign n6637 = ~n6542 & ~n6543 ;
  assign n6638 = ~n6549 & n6637 ;
  assign n6639 = n6549 & ~n6637 ;
  assign n6640 = ~n6638 & ~n6639 ;
  assign n6641 = ~n6636 & ~n6640 ;
  assign n6642 = n6636 & n6640 ;
  assign n6643 = ~n6451 & ~n6452 ;
  assign n6644 = ~n6458 & n6643 ;
  assign n6645 = n6458 & ~n6643 ;
  assign n6646 = ~n6644 & ~n6645 ;
  assign n6647 = ~n6642 & ~n6646 ;
  assign n6648 = ~n6641 & ~n6647 ;
  assign n6649 = ~n6533 & ~n6534 ;
  assign n6650 = ~n6551 & n6649 ;
  assign n6651 = n6551 & ~n6649 ;
  assign n6652 = ~n6650 & ~n6651 ;
  assign n6653 = ~n6648 & n6652 ;
  assign n6654 = n6648 & ~n6652 ;
  assign n6655 = ~n6479 & ~n6480 ;
  assign n6656 = ~n6504 & n6655 ;
  assign n6657 = n6504 & ~n6655 ;
  assign n6658 = ~n6656 & ~n6657 ;
  assign n6659 = ~n6654 & ~n6658 ;
  assign n6660 = ~n6653 & ~n6659 ;
  assign n6661 = ~n6507 & ~n6508 ;
  assign n6662 = n6524 & n6661 ;
  assign n6663 = ~n6524 & ~n6661 ;
  assign n6664 = ~n6662 & ~n6663 ;
  assign n6665 = n6660 & ~n6664 ;
  assign n6666 = ~n6660 & n6664 ;
  assign n6667 = ~n6558 & ~n6559 ;
  assign n6668 = ~n6571 & n6667 ;
  assign n6669 = n6571 & ~n6667 ;
  assign n6670 = ~n6668 & ~n6669 ;
  assign n6671 = ~n6666 & n6670 ;
  assign n6672 = ~n6665 & ~n6671 ;
  assign n6673 = ~n6632 & ~n6672 ;
  assign n6674 = n6632 & n6672 ;
  assign n6675 = ~n6370 & ~n6371 ;
  assign n6676 = ~n6436 & n6675 ;
  assign n6677 = n6436 & ~n6675 ;
  assign n6678 = ~n6676 & ~n6677 ;
  assign n6679 = ~n6653 & ~n6654 ;
  assign n6680 = ~n6658 & n6679 ;
  assign n6681 = n6658 & ~n6679 ;
  assign n6682 = ~n6680 & ~n6681 ;
  assign n6683 = ~n6678 & ~n6682 ;
  assign n6684 = n6678 & n6682 ;
  assign n6685 = \P4_datao_reg[8]/NET0131  & n4405 ;
  assign n6686 = \P4_datao_reg[9]/NET0131  & n4407 ;
  assign n6687 = ~n6685 & ~n6686 ;
  assign n6688 = ~n4398 & n6687 ;
  assign n6689 = n4398 & ~n6687 ;
  assign n6690 = ~n6688 & ~n6689 ;
  assign n6691 = \P4_datao_reg[1]/NET0131  & n4376 ;
  assign n6692 = \P4_datao_reg[0]/NET0131  & n4374 ;
  assign n6693 = ~n6691 & ~n6692 ;
  assign n6694 = n4368 & n6693 ;
  assign n6695 = \P4_datao_reg[0]/NET0131  & n4376 ;
  assign n6696 = n4368 & n6695 ;
  assign n6697 = ~n6693 & ~n6696 ;
  assign n6698 = ~n6694 & ~n6697 ;
  assign n6699 = n6690 & ~n6698 ;
  assign n6700 = n6694 & ~n6695 ;
  assign n6701 = ~n6699 & ~n6700 ;
  assign n6702 = \P4_datao_reg[12]/NET0131  & n4335 ;
  assign n6703 = \P4_datao_reg[13]/NET0131  & n4337 ;
  assign n6704 = ~n6702 & ~n6703 ;
  assign n6705 = ~n4328 & n6704 ;
  assign n6706 = n4328 & ~n6704 ;
  assign n6707 = ~n6705 & ~n6706 ;
  assign n6708 = \P4_datao_reg[15]/NET0131  & n4343 ;
  assign n6709 = ~\din[1]_pad  & n6708 ;
  assign n6710 = \P4_datao_reg[14]/NET0131  & ~n4343 ;
  assign n6711 = n4329 & ~n6708 ;
  assign n6712 = ~n6710 & n6711 ;
  assign n6713 = ~n6709 & ~n6712 ;
  assign n6714 = n6707 & ~n6713 ;
  assign n6715 = ~n6701 & n6714 ;
  assign n6716 = n6701 & ~n6714 ;
  assign n6717 = \P4_datao_reg[7]/NET0131  & n4507 ;
  assign n6718 = \P4_datao_reg[6]/NET0131  & n4511 ;
  assign n6719 = ~n6717 & ~n6718 ;
  assign n6720 = n4431 & ~n6719 ;
  assign n6721 = ~n4431 & n6719 ;
  assign n6722 = ~n6720 & ~n6721 ;
  assign n6723 = \P4_datao_reg[5]/NET0131  & n4435 ;
  assign n6724 = \P4_datao_reg[4]/NET0131  & n4439 ;
  assign n6725 = ~n6723 & ~n6724 ;
  assign n6726 = n4352 & ~n6725 ;
  assign n6727 = ~n4352 & n6725 ;
  assign n6728 = ~n6726 & ~n6727 ;
  assign n6729 = n6722 & n6728 ;
  assign n6730 = ~n6722 & ~n6728 ;
  assign n6731 = \P4_datao_reg[10]/NET0131  & n4552 ;
  assign n6732 = \P4_datao_reg[11]/NET0131  & n4548 ;
  assign n6733 = ~n6731 & ~n6732 ;
  assign n6734 = n4399 & ~n6733 ;
  assign n6735 = ~n4399 & n6733 ;
  assign n6736 = ~n6734 & ~n6735 ;
  assign n6737 = ~n6730 & n6736 ;
  assign n6738 = ~n6729 & ~n6737 ;
  assign n6739 = ~n6716 & ~n6738 ;
  assign n6740 = ~n6715 & ~n6739 ;
  assign n6741 = ~n6416 & ~n6417 ;
  assign n6742 = ~n6434 & n6741 ;
  assign n6743 = n6434 & ~n6741 ;
  assign n6744 = ~n6742 & ~n6743 ;
  assign n6745 = ~n6740 & n6744 ;
  assign n6746 = n6740 & ~n6744 ;
  assign n6747 = ~n6390 & ~n6392 ;
  assign n6748 = n6377 & n6747 ;
  assign n6749 = ~n6377 & ~n6747 ;
  assign n6750 = ~n6748 & ~n6749 ;
  assign n6751 = ~n6425 & ~n6426 ;
  assign n6752 = n6432 & n6751 ;
  assign n6753 = ~n6432 & ~n6751 ;
  assign n6754 = ~n6752 & ~n6753 ;
  assign n6755 = n6750 & n6754 ;
  assign n6756 = ~n6750 & ~n6754 ;
  assign n6757 = ~n6406 & ~n6407 ;
  assign n6758 = ~n6413 & n6757 ;
  assign n6759 = n6413 & ~n6757 ;
  assign n6760 = ~n6758 & ~n6759 ;
  assign n6761 = ~n6756 & ~n6760 ;
  assign n6762 = ~n6755 & ~n6761 ;
  assign n6763 = ~n6746 & ~n6762 ;
  assign n6764 = ~n6745 & ~n6763 ;
  assign n6765 = ~n6684 & n6764 ;
  assign n6766 = ~n6683 & ~n6765 ;
  assign n6767 = ~n6665 & ~n6666 ;
  assign n6768 = n6670 & n6767 ;
  assign n6769 = ~n6670 & ~n6767 ;
  assign n6770 = ~n6768 & ~n6769 ;
  assign n6771 = n6766 & ~n6770 ;
  assign n6772 = ~n6674 & ~n6771 ;
  assign n6773 = ~n6673 & ~n6772 ;
  assign n6774 = n6628 & n6773 ;
  assign n6775 = n6624 & ~n6626 ;
  assign n6776 = ~n6605 & ~n6619 ;
  assign n6777 = ~n6627 & n6776 ;
  assign n6778 = ~n6775 & ~n6777 ;
  assign n6779 = ~n6774 & n6778 ;
  assign n6780 = ~n6766 & n6770 ;
  assign n6781 = ~n6673 & ~n6780 ;
  assign n6782 = n6628 & n6781 ;
  assign n6783 = ~n6707 & n6713 ;
  assign n6784 = ~n6714 & ~n6783 ;
  assign n6785 = \P4_datao_reg[3]/NET0131  & n4356 ;
  assign n6786 = \P4_datao_reg[2]/NET0131  & n4360 ;
  assign n6787 = ~n6785 & ~n6786 ;
  assign n6788 = n4351 & ~n6787 ;
  assign n6789 = ~n4351 & n6787 ;
  assign n6790 = ~n6788 & ~n6789 ;
  assign n6791 = n6784 & n6790 ;
  assign n6792 = ~n6784 & ~n6790 ;
  assign n6793 = \P4_datao_reg[14]/NET0131  & n4343 ;
  assign n6794 = ~\din[1]_pad  & n6793 ;
  assign n6795 = \P4_datao_reg[13]/NET0131  & ~n4343 ;
  assign n6796 = n4329 & ~n6793 ;
  assign n6797 = ~n6795 & n6796 ;
  assign n6798 = ~n6794 & ~n6797 ;
  assign n6799 = n6695 & ~n6798 ;
  assign n6800 = ~n6695 & n6798 ;
  assign n6801 = \P4_datao_reg[8]/NET0131  & n4407 ;
  assign n6802 = \P4_datao_reg[7]/NET0131  & n4405 ;
  assign n6803 = ~n6801 & ~n6802 ;
  assign n6804 = n4398 & ~n6803 ;
  assign n6805 = ~n4398 & n6803 ;
  assign n6806 = ~n6804 & ~n6805 ;
  assign n6807 = ~n6800 & n6806 ;
  assign n6808 = ~n6799 & ~n6807 ;
  assign n6809 = ~n6792 & ~n6808 ;
  assign n6810 = ~n6791 & ~n6809 ;
  assign n6811 = ~n6715 & ~n6716 ;
  assign n6812 = ~n6738 & n6811 ;
  assign n6813 = n6738 & ~n6811 ;
  assign n6814 = ~n6812 & ~n6813 ;
  assign n6815 = ~n6810 & n6814 ;
  assign n6816 = n6810 & ~n6814 ;
  assign n6817 = \P4_datao_reg[10]/NET0131  & n4548 ;
  assign n6818 = \P4_datao_reg[9]/NET0131  & n4552 ;
  assign n6819 = ~n6817 & ~n6818 ;
  assign n6820 = n4399 & ~n6819 ;
  assign n6821 = ~n4399 & n6819 ;
  assign n6822 = ~n6820 & ~n6821 ;
  assign n6823 = \P4_datao_reg[5]/NET0131  & n4511 ;
  assign n6824 = \P4_datao_reg[6]/NET0131  & n4507 ;
  assign n6825 = ~n6823 & ~n6824 ;
  assign n6826 = n4431 & ~n6825 ;
  assign n6827 = ~n4431 & n6825 ;
  assign n6828 = ~n6826 & ~n6827 ;
  assign n6829 = \P4_datao_reg[12]/NET0131  & n4337 ;
  assign n6830 = \P4_datao_reg[11]/NET0131  & n4335 ;
  assign n6831 = ~n6829 & ~n6830 ;
  assign n6832 = n4328 & ~n6831 ;
  assign n6833 = ~n4328 & n6831 ;
  assign n6834 = ~n6832 & ~n6833 ;
  assign n6835 = n6828 & n6834 ;
  assign n6836 = ~n6822 & ~n6835 ;
  assign n6837 = ~n6828 & ~n6834 ;
  assign n6838 = ~n6836 & ~n6837 ;
  assign n6839 = ~n6698 & ~n6700 ;
  assign n6840 = n6690 & n6839 ;
  assign n6841 = ~n6690 & ~n6839 ;
  assign n6842 = ~n6840 & ~n6841 ;
  assign n6843 = n6838 & n6842 ;
  assign n6844 = ~n6838 & ~n6842 ;
  assign n6845 = ~n6729 & ~n6730 ;
  assign n6846 = ~n6736 & n6845 ;
  assign n6847 = n6736 & ~n6845 ;
  assign n6848 = ~n6846 & ~n6847 ;
  assign n6849 = ~n6844 & ~n6848 ;
  assign n6850 = ~n6843 & ~n6849 ;
  assign n6851 = ~n6816 & ~n6850 ;
  assign n6852 = ~n6815 & ~n6851 ;
  assign n6853 = ~n6641 & ~n6642 ;
  assign n6854 = ~n6646 & n6853 ;
  assign n6855 = n6646 & ~n6853 ;
  assign n6856 = ~n6854 & ~n6855 ;
  assign n6857 = ~n6852 & n6856 ;
  assign n6858 = n6852 & ~n6856 ;
  assign n6859 = ~n6745 & ~n6746 ;
  assign n6860 = ~n6762 & n6859 ;
  assign n6861 = n6762 & ~n6859 ;
  assign n6862 = ~n6860 & ~n6861 ;
  assign n6863 = ~n6858 & n6862 ;
  assign n6864 = ~n6857 & ~n6863 ;
  assign n6865 = ~n6683 & ~n6684 ;
  assign n6866 = n6764 & n6865 ;
  assign n6867 = ~n6764 & ~n6865 ;
  assign n6868 = ~n6866 & ~n6867 ;
  assign n6869 = n6864 & n6868 ;
  assign n6870 = \P4_datao_reg[3]/NET0131  & n4439 ;
  assign n6871 = \P4_datao_reg[4]/NET0131  & n4435 ;
  assign n6872 = ~n6870 & ~n6871 ;
  assign n6873 = ~n4352 & n6872 ;
  assign n6874 = n4352 & ~n6872 ;
  assign n6875 = ~n6873 & ~n6874 ;
  assign n6876 = \P4_datao_reg[2]/NET0131  & n4356 ;
  assign n6877 = \P4_datao_reg[1]/NET0131  & n4360 ;
  assign n6878 = ~n6876 & ~n6877 ;
  assign n6879 = n4351 & ~n6878 ;
  assign n6880 = ~n4351 & n6878 ;
  assign n6881 = ~n6879 & ~n6880 ;
  assign n6882 = ~n6875 & ~n6881 ;
  assign n6883 = n6875 & n6881 ;
  assign n6884 = \P4_datao_reg[11]/NET0131  & n4337 ;
  assign n6885 = \P4_datao_reg[10]/NET0131  & n4335 ;
  assign n6886 = ~n6884 & ~n6885 ;
  assign n6887 = n4328 & ~n6886 ;
  assign n6888 = ~n4328 & n6886 ;
  assign n6889 = ~n6887 & ~n6888 ;
  assign n6890 = \P4_datao_reg[13]/NET0131  & n4343 ;
  assign n6891 = ~\din[1]_pad  & n6890 ;
  assign n6892 = \P4_datao_reg[12]/NET0131  & ~n4343 ;
  assign n6893 = n4329 & ~n6890 ;
  assign n6894 = ~n6892 & n6893 ;
  assign n6895 = ~n6891 & ~n6894 ;
  assign n6896 = n6889 & ~n6895 ;
  assign n6897 = ~n6883 & ~n6896 ;
  assign n6898 = ~n6882 & ~n6897 ;
  assign n6899 = ~n6791 & ~n6792 ;
  assign n6900 = ~n6808 & n6899 ;
  assign n6901 = n6808 & ~n6899 ;
  assign n6902 = ~n6900 & ~n6901 ;
  assign n6903 = ~n6898 & ~n6902 ;
  assign n6904 = n6898 & n6902 ;
  assign n6905 = \P4_datao_reg[0]/NET0131  & n4360 ;
  assign n6906 = \P4_datao_reg[1]/NET0131  & n4356 ;
  assign n6907 = ~n6905 & ~n6906 ;
  assign n6908 = n4351 & ~n6907 ;
  assign n6909 = ~n4351 & n6907 ;
  assign n6910 = ~n6908 & ~n6909 ;
  assign n6911 = \P4_datao_reg[9]/NET0131  & n4548 ;
  assign n6912 = \P4_datao_reg[8]/NET0131  & n4552 ;
  assign n6913 = ~n6911 & ~n6912 ;
  assign n6914 = n4399 & ~n6913 ;
  assign n6915 = ~n4399 & n6913 ;
  assign n6916 = ~n6914 & ~n6915 ;
  assign n6917 = n6910 & n6916 ;
  assign n6918 = ~n6910 & ~n6916 ;
  assign n6919 = \P4_datao_reg[2]/NET0131  & n4439 ;
  assign n6920 = \P4_datao_reg[3]/NET0131  & n4435 ;
  assign n6921 = ~n6919 & ~n6920 ;
  assign n6922 = n4352 & ~n6921 ;
  assign n6923 = ~n4352 & n6921 ;
  assign n6924 = ~n6922 & ~n6923 ;
  assign n6925 = ~n6918 & n6924 ;
  assign n6926 = ~n6917 & ~n6925 ;
  assign n6927 = \P4_datao_reg[0]/NET0131  & n4356 ;
  assign n6928 = n4351 & ~n6927 ;
  assign n6929 = \P4_datao_reg[6]/NET0131  & n4405 ;
  assign n6930 = \P4_datao_reg[7]/NET0131  & n4407 ;
  assign n6931 = ~n6929 & ~n6930 ;
  assign n6932 = ~n4398 & n6931 ;
  assign n6933 = n4398 & ~n6931 ;
  assign n6934 = ~n6932 & ~n6933 ;
  assign n6935 = ~n6928 & ~n6934 ;
  assign n6936 = n6928 & n6934 ;
  assign n6937 = \P4_datao_reg[4]/NET0131  & n4511 ;
  assign n6938 = \P4_datao_reg[5]/NET0131  & n4507 ;
  assign n6939 = ~n6937 & ~n6938 ;
  assign n6940 = n4431 & ~n6939 ;
  assign n6941 = ~n4431 & n6939 ;
  assign n6942 = ~n6940 & ~n6941 ;
  assign n6943 = ~n6936 & ~n6942 ;
  assign n6944 = ~n6935 & ~n6943 ;
  assign n6945 = n6926 & ~n6944 ;
  assign n6946 = ~n6926 & n6944 ;
  assign n6947 = ~n6799 & ~n6800 ;
  assign n6948 = n6806 & n6947 ;
  assign n6949 = ~n6806 & ~n6947 ;
  assign n6950 = ~n6948 & ~n6949 ;
  assign n6951 = ~n6946 & ~n6950 ;
  assign n6952 = ~n6945 & ~n6951 ;
  assign n6953 = ~n6904 & ~n6952 ;
  assign n6954 = ~n6903 & ~n6953 ;
  assign n6955 = ~n6755 & ~n6756 ;
  assign n6956 = ~n6760 & n6955 ;
  assign n6957 = n6760 & ~n6955 ;
  assign n6958 = ~n6956 & ~n6957 ;
  assign n6959 = ~n6954 & ~n6958 ;
  assign n6960 = n6954 & n6958 ;
  assign n6961 = ~n6815 & ~n6816 ;
  assign n6962 = ~n6850 & n6961 ;
  assign n6963 = n6850 & ~n6961 ;
  assign n6964 = ~n6962 & ~n6963 ;
  assign n6965 = ~n6960 & ~n6964 ;
  assign n6966 = ~n6959 & ~n6965 ;
  assign n6967 = ~n6857 & ~n6858 ;
  assign n6968 = ~n6862 & n6967 ;
  assign n6969 = n6862 & ~n6967 ;
  assign n6970 = ~n6968 & ~n6969 ;
  assign n6971 = ~n6966 & n6970 ;
  assign n6972 = ~n6869 & ~n6971 ;
  assign n6973 = ~n6835 & ~n6837 ;
  assign n6974 = n6822 & n6973 ;
  assign n6975 = ~n6822 & ~n6973 ;
  assign n6976 = ~n6974 & ~n6975 ;
  assign n6977 = ~n6882 & ~n6883 ;
  assign n6978 = n6896 & n6977 ;
  assign n6979 = ~n6896 & ~n6977 ;
  assign n6980 = ~n6978 & ~n6979 ;
  assign n6981 = n6976 & n6980 ;
  assign n6982 = ~n6976 & ~n6980 ;
  assign n6983 = ~n6889 & n6895 ;
  assign n6984 = ~n6896 & ~n6983 ;
  assign n6985 = \P4_datao_reg[10]/NET0131  & n4337 ;
  assign n6986 = \P4_datao_reg[9]/NET0131  & n4335 ;
  assign n6987 = ~n6985 & ~n6986 ;
  assign n6988 = n4328 & ~n6987 ;
  assign n6989 = ~n4328 & n6987 ;
  assign n6990 = ~n6988 & ~n6989 ;
  assign n6991 = n6927 & n6990 ;
  assign n6992 = ~n6927 & ~n6990 ;
  assign n6993 = \P4_datao_reg[6]/NET0131  & n4407 ;
  assign n6994 = \P4_datao_reg[5]/NET0131  & n4405 ;
  assign n6995 = ~n6993 & ~n6994 ;
  assign n6996 = n4398 & ~n6995 ;
  assign n6997 = ~n4398 & n6995 ;
  assign n6998 = ~n6996 & ~n6997 ;
  assign n6999 = ~n6992 & n6998 ;
  assign n7000 = ~n6991 & ~n6999 ;
  assign n7001 = n6984 & ~n7000 ;
  assign n7002 = ~n6984 & n7000 ;
  assign n7003 = \P4_datao_reg[2]/NET0131  & n4435 ;
  assign n7004 = \P4_datao_reg[1]/NET0131  & n4439 ;
  assign n7005 = ~n7003 & ~n7004 ;
  assign n7006 = n4352 & ~n7005 ;
  assign n7007 = ~n4352 & n7005 ;
  assign n7008 = ~n7006 & ~n7007 ;
  assign n7009 = \P4_datao_reg[12]/NET0131  & n4343 ;
  assign n7010 = ~\din[1]_pad  & n7009 ;
  assign n7011 = n4329 & ~n4343 ;
  assign n7012 = \P4_datao_reg[11]/NET0131  & n7011 ;
  assign n7013 = n4329 & ~n7009 ;
  assign n7014 = ~n7012 & n7013 ;
  assign n7015 = ~n7010 & ~n7014 ;
  assign n7016 = n7008 & ~n7015 ;
  assign n7017 = ~n7008 & n7015 ;
  assign n7018 = \P4_datao_reg[3]/NET0131  & n4511 ;
  assign n7019 = \P4_datao_reg[4]/NET0131  & n4507 ;
  assign n7020 = ~n7018 & ~n7019 ;
  assign n7021 = n4431 & ~n7020 ;
  assign n7022 = ~n4431 & n7020 ;
  assign n7023 = ~n7021 & ~n7022 ;
  assign n7024 = ~n7017 & n7023 ;
  assign n7025 = ~n7016 & ~n7024 ;
  assign n7026 = ~n7002 & ~n7025 ;
  assign n7027 = ~n7001 & ~n7026 ;
  assign n7028 = ~n6982 & ~n7027 ;
  assign n7029 = ~n6981 & ~n7028 ;
  assign n7030 = ~n6843 & ~n6844 ;
  assign n7031 = ~n6848 & n7030 ;
  assign n7032 = n6848 & ~n7030 ;
  assign n7033 = ~n7031 & ~n7032 ;
  assign n7034 = n7029 & ~n7033 ;
  assign n7035 = ~n7029 & n7033 ;
  assign n7036 = ~n6903 & ~n6904 ;
  assign n7037 = ~n6952 & n7036 ;
  assign n7038 = n6952 & ~n7036 ;
  assign n7039 = ~n7037 & ~n7038 ;
  assign n7040 = ~n7035 & n7039 ;
  assign n7041 = ~n7034 & ~n7040 ;
  assign n7042 = ~n6959 & ~n6960 ;
  assign n7043 = ~n6964 & n7042 ;
  assign n7044 = n6964 & ~n7042 ;
  assign n7045 = ~n7043 & ~n7044 ;
  assign n7046 = n7041 & ~n7045 ;
  assign n7047 = ~n7041 & n7045 ;
  assign n7048 = ~n6917 & ~n6918 ;
  assign n7049 = ~n6924 & n7048 ;
  assign n7050 = n6924 & ~n7048 ;
  assign n7051 = ~n7049 & ~n7050 ;
  assign n7052 = ~n6935 & ~n6936 ;
  assign n7053 = ~n6942 & n7052 ;
  assign n7054 = n6942 & ~n7052 ;
  assign n7055 = ~n7053 & ~n7054 ;
  assign n7056 = ~n7051 & ~n7055 ;
  assign n7057 = n7051 & n7055 ;
  assign n7058 = \P4_datao_reg[9]/NET0131  & n4337 ;
  assign n7059 = \P4_datao_reg[8]/NET0131  & n4335 ;
  assign n7060 = ~n7058 & ~n7059 ;
  assign n7061 = ~n4328 & n7060 ;
  assign n7062 = n4328 & ~n7060 ;
  assign n7063 = ~n7061 & ~n7062 ;
  assign n7064 = \P4_datao_reg[11]/NET0131  & n4343 ;
  assign n7065 = ~\din[1]_pad  & n7064 ;
  assign n7066 = \P4_datao_reg[10]/NET0131  & n7011 ;
  assign n7067 = n4329 & ~n7064 ;
  assign n7068 = ~n7066 & n7067 ;
  assign n7069 = ~n7065 & ~n7068 ;
  assign n7070 = n7063 & ~n7069 ;
  assign n7071 = \P4_datao_reg[8]/NET0131  & n4548 ;
  assign n7072 = \P4_datao_reg[7]/NET0131  & n4552 ;
  assign n7073 = ~n7071 & ~n7072 ;
  assign n7074 = n4399 & ~n7073 ;
  assign n7075 = ~n4399 & n7073 ;
  assign n7076 = ~n7074 & ~n7075 ;
  assign n7077 = n7070 & n7076 ;
  assign n7078 = ~n7070 & ~n7076 ;
  assign n7079 = \P4_datao_reg[7]/NET0131  & n4548 ;
  assign n7080 = \P4_datao_reg[6]/NET0131  & n4552 ;
  assign n7081 = ~n7079 & ~n7080 ;
  assign n7082 = n4399 & ~n7081 ;
  assign n7083 = ~n4399 & n7081 ;
  assign n7084 = ~n7082 & ~n7083 ;
  assign n7085 = \P4_datao_reg[5]/NET0131  & n4407 ;
  assign n7086 = \P4_datao_reg[4]/NET0131  & n4405 ;
  assign n7087 = ~n7085 & ~n7086 ;
  assign n7088 = n4398 & ~n7087 ;
  assign n7089 = ~n4398 & n7087 ;
  assign n7090 = ~n7088 & ~n7089 ;
  assign n7091 = n7084 & n7090 ;
  assign n7092 = ~n7084 & ~n7090 ;
  assign n7093 = \P4_datao_reg[3]/NET0131  & n4507 ;
  assign n7094 = \P4_datao_reg[2]/NET0131  & n4511 ;
  assign n7095 = ~n7093 & ~n7094 ;
  assign n7096 = n4431 & ~n7095 ;
  assign n7097 = ~n4431 & n7095 ;
  assign n7098 = ~n7096 & ~n7097 ;
  assign n7099 = ~n7092 & n7098 ;
  assign n7100 = ~n7091 & ~n7099 ;
  assign n7101 = ~n7078 & ~n7100 ;
  assign n7102 = ~n7077 & ~n7101 ;
  assign n7103 = ~n7057 & ~n7102 ;
  assign n7104 = ~n7056 & ~n7103 ;
  assign n7105 = ~n6981 & ~n6982 ;
  assign n7106 = ~n7027 & n7105 ;
  assign n7107 = n7027 & ~n7105 ;
  assign n7108 = ~n7106 & ~n7107 ;
  assign n7109 = n7104 & ~n7108 ;
  assign n7110 = ~n7104 & n7108 ;
  assign n7111 = ~n6945 & ~n6946 ;
  assign n7112 = ~n6950 & n7111 ;
  assign n7113 = n6950 & ~n7111 ;
  assign n7114 = ~n7112 & ~n7113 ;
  assign n7115 = ~n7110 & n7114 ;
  assign n7116 = ~n7109 & ~n7115 ;
  assign n7117 = ~n7034 & ~n7035 ;
  assign n7118 = n7039 & n7117 ;
  assign n7119 = ~n7039 & ~n7117 ;
  assign n7120 = ~n7118 & ~n7119 ;
  assign n7121 = n7116 & ~n7120 ;
  assign n7122 = ~n7047 & n7121 ;
  assign n7123 = ~n7046 & ~n7122 ;
  assign n7124 = n6972 & ~n7123 ;
  assign n7125 = ~n6864 & ~n6868 ;
  assign n7126 = n6966 & ~n6970 ;
  assign n7127 = ~n6869 & n7126 ;
  assign n7128 = ~n7125 & ~n7127 ;
  assign n7129 = ~n7124 & n7128 ;
  assign n7130 = n6782 & ~n7129 ;
  assign n7131 = n6779 & ~n7130 ;
  assign n7132 = n6314 & ~n7131 ;
  assign n7133 = ~n6258 & ~n6284 ;
  assign n7134 = ~n6205 & n6255 ;
  assign n7135 = ~n6285 & n7134 ;
  assign n7136 = ~n7133 & ~n7135 ;
  assign n7137 = n6313 & ~n7136 ;
  assign n7138 = n6307 & n6311 ;
  assign n7139 = ~n6302 & ~n6304 ;
  assign n7140 = ~n7138 & ~n7139 ;
  assign n7141 = ~n6312 & ~n7140 ;
  assign n7142 = ~n7137 & ~n7141 ;
  assign n7143 = ~n7132 & n7142 ;
  assign n7144 = n5854 & ~n7143 ;
  assign n7147 = \P4_datao_reg[6]/NET0131  & n4548 ;
  assign n7148 = \P4_datao_reg[5]/NET0131  & n4552 ;
  assign n7149 = ~n7147 & ~n7148 ;
  assign n7150 = n4399 & ~n7149 ;
  assign n7151 = ~n4399 & n7149 ;
  assign n7152 = ~n7150 & ~n7151 ;
  assign n7153 = \P4_datao_reg[10]/NET0131  & n4343 ;
  assign n7154 = ~\din[1]_pad  & n7153 ;
  assign n7155 = \P4_datao_reg[9]/NET0131  & ~n4343 ;
  assign n7156 = n4329 & ~n7153 ;
  assign n7157 = ~n7155 & n7156 ;
  assign n7158 = ~n7154 & ~n7157 ;
  assign n7159 = n7152 & ~n7158 ;
  assign n7160 = ~n7152 & n7158 ;
  assign n7161 = \P4_datao_reg[2]/NET0131  & n4507 ;
  assign n7162 = \P4_datao_reg[1]/NET0131  & n4511 ;
  assign n7163 = ~n7161 & ~n7162 ;
  assign n7164 = n4431 & ~n7163 ;
  assign n7165 = ~n4431 & n7163 ;
  assign n7166 = ~n7164 & ~n7165 ;
  assign n7167 = ~n7160 & n7166 ;
  assign n7168 = ~n7159 & ~n7167 ;
  assign n7169 = \P4_datao_reg[0]/NET0131  & n4435 ;
  assign n7170 = \P4_datao_reg[7]/NET0131  & n4335 ;
  assign n7171 = \P4_datao_reg[8]/NET0131  & n4337 ;
  assign n7172 = ~n7170 & ~n7171 ;
  assign n7173 = ~n4328 & n7172 ;
  assign n7174 = n4328 & ~n7172 ;
  assign n7175 = ~n7173 & ~n7174 ;
  assign n7176 = n7169 & n7175 ;
  assign n7177 = ~n7169 & ~n7175 ;
  assign n7178 = \P4_datao_reg[4]/NET0131  & n4407 ;
  assign n7179 = \P4_datao_reg[3]/NET0131  & n4405 ;
  assign n7180 = ~n7178 & ~n7179 ;
  assign n7181 = n4398 & ~n7180 ;
  assign n7182 = ~n4398 & n7180 ;
  assign n7183 = ~n7181 & ~n7182 ;
  assign n7184 = ~n7177 & n7183 ;
  assign n7185 = ~n7176 & ~n7184 ;
  assign n7186 = ~n7168 & ~n7185 ;
  assign n7187 = n7168 & n7185 ;
  assign n7188 = ~n7186 & ~n7187 ;
  assign n7189 = ~n7091 & ~n7092 ;
  assign n7190 = ~n7098 & n7189 ;
  assign n7191 = n7098 & ~n7189 ;
  assign n7192 = ~n7190 & ~n7191 ;
  assign n7193 = n7188 & ~n7192 ;
  assign n7194 = ~n7188 & n7192 ;
  assign n7195 = ~n7193 & ~n7194 ;
  assign n7196 = ~n7063 & n7069 ;
  assign n7197 = ~n7070 & ~n7196 ;
  assign n7198 = \P4_datao_reg[1]/NET0131  & n4435 ;
  assign n7199 = \P4_datao_reg[0]/NET0131  & n4439 ;
  assign n7200 = ~n7198 & ~n7199 ;
  assign n7201 = n4352 & n7200 ;
  assign n7202 = ~n7169 & n7201 ;
  assign n7203 = n4352 & n7169 ;
  assign n7204 = ~n7200 & ~n7203 ;
  assign n7205 = ~n7201 & ~n7204 ;
  assign n7206 = ~n7202 & ~n7205 ;
  assign n7207 = n7197 & ~n7206 ;
  assign n7208 = ~n7197 & n7206 ;
  assign n7209 = ~n7207 & ~n7208 ;
  assign n7210 = n7195 & ~n7209 ;
  assign n7211 = ~n7195 & n7209 ;
  assign n7212 = \P4_datao_reg[7]/NET0131  & n4337 ;
  assign n7213 = \P4_datao_reg[6]/NET0131  & n4335 ;
  assign n7214 = ~n7212 & ~n7213 ;
  assign n7215 = n4328 & ~n7214 ;
  assign n7216 = ~n4328 & n7214 ;
  assign n7217 = ~n7215 & ~n7216 ;
  assign n7218 = \P4_datao_reg[9]/NET0131  & n4343 ;
  assign n7219 = ~\din[1]_pad  & n7218 ;
  assign n7220 = \P4_datao_reg[8]/NET0131  & ~n4343 ;
  assign n7221 = n4329 & ~n7218 ;
  assign n7222 = ~n7220 & n7221 ;
  assign n7223 = ~n7219 & ~n7222 ;
  assign n7224 = n7217 & ~n7223 ;
  assign n7225 = \P4_datao_reg[0]/NET0131  & n4511 ;
  assign n7226 = \P4_datao_reg[1]/NET0131  & n4507 ;
  assign n7227 = ~n7225 & ~n7226 ;
  assign n7228 = n4431 & ~n7227 ;
  assign n7229 = ~n4431 & n7227 ;
  assign n7230 = ~n7228 & ~n7229 ;
  assign n7231 = \P4_datao_reg[3]/NET0131  & n4407 ;
  assign n7232 = \P4_datao_reg[2]/NET0131  & n4405 ;
  assign n7233 = ~n7231 & ~n7232 ;
  assign n7234 = n4398 & ~n7233 ;
  assign n7235 = ~n4398 & n7233 ;
  assign n7236 = ~n7234 & ~n7235 ;
  assign n7237 = n7230 & n7236 ;
  assign n7238 = ~n7230 & ~n7236 ;
  assign n7239 = \P4_datao_reg[5]/NET0131  & n4548 ;
  assign n7240 = \P4_datao_reg[4]/NET0131  & n4552 ;
  assign n7241 = ~n7239 & ~n7240 ;
  assign n7242 = n4399 & ~n7241 ;
  assign n7243 = ~n4399 & n7241 ;
  assign n7244 = ~n7242 & ~n7243 ;
  assign n7245 = ~n7238 & n7244 ;
  assign n7246 = ~n7237 & ~n7245 ;
  assign n7247 = n7224 & ~n7246 ;
  assign n7248 = ~n7224 & n7246 ;
  assign n7249 = ~n7176 & ~n7177 ;
  assign n7250 = n7183 & n7249 ;
  assign n7251 = ~n7183 & ~n7249 ;
  assign n7252 = ~n7250 & ~n7251 ;
  assign n7253 = ~n7248 & n7252 ;
  assign n7254 = ~n7247 & ~n7253 ;
  assign n7255 = ~n7211 & ~n7254 ;
  assign n7256 = ~n7210 & ~n7255 ;
  assign n7257 = ~n7187 & ~n7192 ;
  assign n7258 = ~n7186 & ~n7257 ;
  assign n7259 = ~n7077 & ~n7078 ;
  assign n7260 = ~n7100 & n7259 ;
  assign n7261 = n7100 & ~n7259 ;
  assign n7262 = ~n7260 & ~n7261 ;
  assign n7263 = n7258 & ~n7262 ;
  assign n7264 = ~n7258 & n7262 ;
  assign n7265 = ~n7263 & ~n7264 ;
  assign n7266 = n7197 & ~n7205 ;
  assign n7267 = ~n7202 & ~n7266 ;
  assign n7268 = ~n6991 & ~n6992 ;
  assign n7269 = n6998 & n7268 ;
  assign n7270 = ~n6998 & ~n7268 ;
  assign n7271 = ~n7269 & ~n7270 ;
  assign n7272 = ~n7016 & ~n7017 ;
  assign n7273 = n7023 & n7272 ;
  assign n7274 = ~n7023 & ~n7272 ;
  assign n7275 = ~n7273 & ~n7274 ;
  assign n7276 = ~n7271 & ~n7275 ;
  assign n7277 = n7271 & n7275 ;
  assign n7278 = ~n7276 & ~n7277 ;
  assign n7279 = n7267 & ~n7278 ;
  assign n7280 = ~n7267 & n7278 ;
  assign n7281 = ~n7279 & ~n7280 ;
  assign n7282 = n7265 & ~n7281 ;
  assign n7283 = ~n7265 & n7281 ;
  assign n7284 = ~n7282 & ~n7283 ;
  assign n7285 = n7256 & n7284 ;
  assign n7286 = \P4_datao_reg[0]/NET0131  & n4507 ;
  assign n7287 = n4431 & ~n7286 ;
  assign n7288 = ~n7217 & n7223 ;
  assign n7289 = ~n7224 & ~n7288 ;
  assign n7290 = n7287 & n7289 ;
  assign n7291 = ~n7287 & ~n7289 ;
  assign n7292 = \P4_datao_reg[8]/NET0131  & n4343 ;
  assign n7293 = ~\din[1]_pad  & n7292 ;
  assign n7294 = \P4_datao_reg[7]/NET0131  & ~n4343 ;
  assign n7295 = n4329 & ~n7292 ;
  assign n7296 = ~n7294 & n7295 ;
  assign n7297 = ~n7293 & ~n7296 ;
  assign n7298 = n7286 & ~n7297 ;
  assign n7299 = ~n7286 & n7297 ;
  assign n7300 = \P4_datao_reg[2]/NET0131  & n4407 ;
  assign n7301 = \P4_datao_reg[1]/NET0131  & n4405 ;
  assign n7302 = ~n7300 & ~n7301 ;
  assign n7303 = n4398 & ~n7302 ;
  assign n7304 = ~n4398 & n7302 ;
  assign n7305 = ~n7303 & ~n7304 ;
  assign n7306 = ~n7299 & n7305 ;
  assign n7307 = ~n7298 & ~n7306 ;
  assign n7308 = ~n7291 & ~n7307 ;
  assign n7309 = ~n7290 & ~n7308 ;
  assign n7310 = ~n7159 & ~n7160 ;
  assign n7311 = n7166 & n7310 ;
  assign n7312 = ~n7166 & ~n7310 ;
  assign n7313 = ~n7311 & ~n7312 ;
  assign n7314 = n7309 & ~n7313 ;
  assign n7315 = ~n7309 & n7313 ;
  assign n7316 = ~n7314 & ~n7315 ;
  assign n7317 = ~n7247 & ~n7248 ;
  assign n7318 = ~n7252 & n7317 ;
  assign n7319 = n7252 & ~n7317 ;
  assign n7320 = ~n7318 & ~n7319 ;
  assign n7321 = n7316 & ~n7320 ;
  assign n7322 = ~n7316 & n7320 ;
  assign n7323 = ~n7321 & ~n7322 ;
  assign n7324 = \P4_datao_reg[6]/NET0131  & n4337 ;
  assign n7325 = \P4_datao_reg[5]/NET0131  & n4335 ;
  assign n7326 = ~n7324 & ~n7325 ;
  assign n7327 = n4328 & ~n7326 ;
  assign n7328 = ~n4328 & n7326 ;
  assign n7329 = ~n7327 & ~n7328 ;
  assign n7330 = \P4_datao_reg[4]/NET0131  & n4548 ;
  assign n7331 = \P4_datao_reg[3]/NET0131  & n4552 ;
  assign n7332 = ~n7330 & ~n7331 ;
  assign n7333 = n4399 & ~n7332 ;
  assign n7334 = ~n4399 & n7332 ;
  assign n7335 = ~n7333 & ~n7334 ;
  assign n7336 = ~n7329 & ~n7335 ;
  assign n7337 = \P4_datao_reg[5]/NET0131  & n4337 ;
  assign n7338 = \P4_datao_reg[4]/NET0131  & n4335 ;
  assign n7339 = ~n7337 & ~n7338 ;
  assign n7340 = n4328 & ~n7339 ;
  assign n7341 = ~n4328 & n7339 ;
  assign n7342 = ~n7340 & ~n7341 ;
  assign n7343 = \P4_datao_reg[7]/NET0131  & n4343 ;
  assign n7344 = ~\din[1]_pad  & n7343 ;
  assign n7345 = \P4_datao_reg[6]/NET0131  & ~n4343 ;
  assign n7346 = n4329 & ~n7343 ;
  assign n7347 = ~n7345 & n7346 ;
  assign n7348 = ~n7344 & ~n7347 ;
  assign n7349 = n7342 & ~n7348 ;
  assign n7350 = n7329 & n7335 ;
  assign n7351 = ~n7349 & ~n7350 ;
  assign n7352 = ~n7336 & ~n7351 ;
  assign n7353 = ~n7237 & ~n7238 ;
  assign n7354 = ~n7244 & n7353 ;
  assign n7355 = n7244 & ~n7353 ;
  assign n7356 = ~n7354 & ~n7355 ;
  assign n7357 = n7352 & ~n7356 ;
  assign n7358 = ~n7352 & n7356 ;
  assign n7359 = ~n7290 & ~n7291 ;
  assign n7360 = ~n7307 & n7359 ;
  assign n7361 = n7307 & ~n7359 ;
  assign n7362 = ~n7360 & ~n7361 ;
  assign n7363 = ~n7358 & n7362 ;
  assign n7364 = ~n7357 & ~n7363 ;
  assign n7365 = ~n7323 & n7364 ;
  assign n7366 = ~n7314 & ~n7320 ;
  assign n7367 = ~n7315 & ~n7366 ;
  assign n7368 = ~n7210 & ~n7211 ;
  assign n7369 = ~n7254 & n7368 ;
  assign n7370 = n7254 & ~n7368 ;
  assign n7371 = ~n7369 & ~n7370 ;
  assign n7372 = n7367 & ~n7371 ;
  assign n7373 = ~n7365 & ~n7372 ;
  assign n7374 = \P4_datao_reg[0]/NET0131  & n4407 ;
  assign n7375 = \P4_datao_reg[1]/NET0131  & n4407 ;
  assign n7376 = \P4_datao_reg[0]/NET0131  & n4405 ;
  assign n7377 = ~n7375 & ~n7376 ;
  assign n7378 = n4398 & n7377 ;
  assign n7379 = ~n7374 & n7378 ;
  assign n7380 = n4398 & n7374 ;
  assign n7381 = ~n7377 & ~n7380 ;
  assign n7382 = ~n7378 & ~n7381 ;
  assign n7383 = \P4_datao_reg[3]/NET0131  & n4548 ;
  assign n7384 = \P4_datao_reg[2]/NET0131  & n4552 ;
  assign n7385 = ~n7383 & ~n7384 ;
  assign n7386 = n4399 & ~n7385 ;
  assign n7387 = ~n4399 & n7385 ;
  assign n7388 = ~n7386 & ~n7387 ;
  assign n7389 = ~n7382 & n7388 ;
  assign n7390 = ~n7379 & ~n7389 ;
  assign n7391 = ~n7298 & ~n7299 ;
  assign n7392 = n7305 & n7391 ;
  assign n7393 = ~n7305 & ~n7391 ;
  assign n7394 = ~n7392 & ~n7393 ;
  assign n7395 = n7390 & ~n7394 ;
  assign n7396 = ~n7390 & n7394 ;
  assign n7397 = ~n7395 & ~n7396 ;
  assign n7398 = ~n7336 & ~n7350 ;
  assign n7399 = ~n7349 & n7398 ;
  assign n7400 = n7349 & ~n7398 ;
  assign n7401 = ~n7399 & ~n7400 ;
  assign n7402 = n7397 & ~n7401 ;
  assign n7403 = ~n7397 & n7401 ;
  assign n7404 = ~n7402 & ~n7403 ;
  assign n7405 = ~n7342 & n7348 ;
  assign n7406 = ~n7349 & ~n7405 ;
  assign n7407 = \P4_datao_reg[4]/NET0131  & n4337 ;
  assign n7408 = \P4_datao_reg[3]/NET0131  & n4335 ;
  assign n7409 = ~n7407 & ~n7408 ;
  assign n7410 = n4328 & ~n7409 ;
  assign n7411 = ~n4328 & n7409 ;
  assign n7412 = ~n7410 & ~n7411 ;
  assign n7413 = n7374 & n7412 ;
  assign n7414 = ~n7374 & ~n7412 ;
  assign n7415 = \P4_datao_reg[6]/NET0131  & n4343 ;
  assign n7416 = ~\din[1]_pad  & n7415 ;
  assign n7417 = \P4_datao_reg[5]/NET0131  & ~n4343 ;
  assign n7418 = n4329 & ~n7415 ;
  assign n7419 = ~n7417 & n7418 ;
  assign n7420 = ~n7416 & ~n7419 ;
  assign n7421 = ~n7414 & ~n7420 ;
  assign n7422 = ~n7413 & ~n7421 ;
  assign n7423 = n7406 & ~n7422 ;
  assign n7424 = ~n7406 & n7422 ;
  assign n7425 = ~n7379 & ~n7382 ;
  assign n7426 = n7388 & ~n7425 ;
  assign n7427 = ~n7388 & n7425 ;
  assign n7428 = ~n7426 & ~n7427 ;
  assign n7429 = ~n7424 & ~n7428 ;
  assign n7430 = ~n7423 & ~n7429 ;
  assign n7431 = ~n7404 & n7430 ;
  assign n7432 = ~n7395 & ~n7401 ;
  assign n7433 = ~n7396 & ~n7432 ;
  assign n7434 = ~n7357 & ~n7358 ;
  assign n7435 = ~n7362 & n7434 ;
  assign n7436 = n7362 & ~n7434 ;
  assign n7437 = ~n7435 & ~n7436 ;
  assign n7438 = n7433 & n7437 ;
  assign n7439 = ~n7431 & ~n7438 ;
  assign n7472 = \P4_datao_reg[0]/NET0131  & n4548 ;
  assign n7473 = \P4_datao_reg[1]/NET0131  & n4548 ;
  assign n7474 = \P4_datao_reg[0]/NET0131  & n4552 ;
  assign n7475 = ~n7473 & ~n7474 ;
  assign n7476 = n4399 & n7475 ;
  assign n7477 = ~n7472 & n7476 ;
  assign n7440 = \P4_datao_reg[3]/NET0131  & n4337 ;
  assign n7441 = \P4_datao_reg[2]/NET0131  & n4335 ;
  assign n7442 = ~n7440 & ~n7441 ;
  assign n7443 = n4328 & ~n7442 ;
  assign n7444 = ~n4328 & n7442 ;
  assign n7445 = ~n7443 & ~n7444 ;
  assign n7446 = \P4_datao_reg[5]/NET0131  & n4343 ;
  assign n7447 = ~\din[1]_pad  & n7446 ;
  assign n7448 = \P4_datao_reg[4]/NET0131  & ~n4343 ;
  assign n7449 = n4329 & ~n7446 ;
  assign n7450 = ~n7448 & n7449 ;
  assign n7451 = ~n7447 & ~n7450 ;
  assign n7452 = n7445 & ~n7451 ;
  assign n7478 = ~n7445 & n7451 ;
  assign n7479 = ~n7452 & ~n7478 ;
  assign n7480 = n4399 & n7472 ;
  assign n7481 = ~n7475 & ~n7480 ;
  assign n7482 = ~n7476 & ~n7481 ;
  assign n7483 = n7479 & ~n7482 ;
  assign n7484 = ~n7477 & ~n7483 ;
  assign n7461 = ~n7413 & ~n7414 ;
  assign n7462 = ~n7420 & n7461 ;
  assign n7463 = n7420 & ~n7461 ;
  assign n7464 = ~n7462 & ~n7463 ;
  assign n7453 = \P4_datao_reg[2]/NET0131  & n4548 ;
  assign n7454 = \P4_datao_reg[1]/NET0131  & n4552 ;
  assign n7455 = ~n7453 & ~n7454 ;
  assign n7456 = n4399 & ~n7455 ;
  assign n7457 = ~n4399 & n7455 ;
  assign n7458 = ~n7456 & ~n7457 ;
  assign n7459 = n7452 & n7458 ;
  assign n7460 = ~n7452 & ~n7458 ;
  assign n7485 = ~n7459 & ~n7460 ;
  assign n7486 = ~n7464 & n7485 ;
  assign n7487 = n7464 & ~n7485 ;
  assign n7488 = ~n7486 & ~n7487 ;
  assign n7555 = ~n7484 & ~n7488 ;
  assign n7490 = \P4_datao_reg[2]/NET0131  & n4337 ;
  assign n7491 = \P4_datao_reg[1]/NET0131  & n4335 ;
  assign n7492 = ~n7490 & ~n7491 ;
  assign n7493 = n4328 & ~n7492 ;
  assign n7494 = ~n4328 & n7492 ;
  assign n7495 = ~n7493 & ~n7494 ;
  assign n7496 = n7472 & n7495 ;
  assign n7497 = ~n7472 & ~n7495 ;
  assign n7498 = \P4_datao_reg[4]/NET0131  & n4343 ;
  assign n7499 = ~\din[1]_pad  & n7498 ;
  assign n7500 = \P4_datao_reg[3]/NET0131  & ~n4343 ;
  assign n7501 = n4329 & ~n7498 ;
  assign n7502 = ~n7500 & n7501 ;
  assign n7503 = ~n7499 & ~n7502 ;
  assign n7504 = ~n7497 & ~n7503 ;
  assign n7505 = ~n7496 & ~n7504 ;
  assign n7506 = ~n7477 & ~n7482 ;
  assign n7507 = n7479 & ~n7506 ;
  assign n7508 = ~n7479 & n7506 ;
  assign n7509 = ~n7507 & ~n7508 ;
  assign n7510 = ~n7505 & ~n7509 ;
  assign n7511 = n7505 & n7509 ;
  assign n7512 = ~n7496 & ~n7497 ;
  assign n7513 = ~n7503 & n7512 ;
  assign n7514 = n7503 & ~n7512 ;
  assign n7515 = ~n7513 & ~n7514 ;
  assign n7516 = \P4_datao_reg[0]/NET0131  & n4337 ;
  assign n7517 = n4328 & ~n7516 ;
  assign n7518 = \P4_datao_reg[3]/NET0131  & n4343 ;
  assign n7519 = ~\din[1]_pad  & n7518 ;
  assign n7520 = \P4_datao_reg[2]/NET0131  & ~n4343 ;
  assign n7521 = n4329 & ~n7518 ;
  assign n7522 = ~n7520 & n7521 ;
  assign n7523 = ~n7519 & ~n7522 ;
  assign n7524 = n7517 & ~n7523 ;
  assign n7525 = ~n7517 & n7523 ;
  assign n7526 = ~n7524 & ~n7525 ;
  assign n7527 = \P4_datao_reg[1]/NET0131  & n4337 ;
  assign n7528 = \P4_datao_reg[0]/NET0131  & n4335 ;
  assign n7529 = ~n7527 & ~n7528 ;
  assign n7530 = n4328 & ~n7529 ;
  assign n7531 = ~n4328 & n7529 ;
  assign n7532 = ~n7530 & ~n7531 ;
  assign n7533 = ~n7526 & ~n7532 ;
  assign n7534 = \P4_datao_reg[2]/NET0131  & n4343 ;
  assign n7535 = ~\din[1]_pad  & n7534 ;
  assign n7536 = \P4_datao_reg[1]/NET0131  & ~n4343 ;
  assign n7537 = n4329 & ~n7534 ;
  assign n7538 = ~n7536 & n7537 ;
  assign n7539 = ~n7535 & ~n7538 ;
  assign n7540 = n7516 & ~n7539 ;
  assign n7541 = ~n7516 & n7539 ;
  assign n7542 = \P4_datao_reg[1]/NET0131  & n4343 ;
  assign n7543 = ~\P4_datao_reg[0]/NET0131  & n4329 ;
  assign n7544 = ~n7542 & n7543 ;
  assign n7545 = ~n7541 & n7544 ;
  assign n7546 = ~n7540 & ~n7545 ;
  assign n7547 = ~n7533 & ~n7546 ;
  assign n7548 = n7526 & n7532 ;
  assign n7549 = ~n7547 & ~n7548 ;
  assign n7550 = ~n7524 & n7549 ;
  assign n7551 = n7515 & ~n7550 ;
  assign n7552 = n7524 & n7547 ;
  assign n7553 = ~n7551 & ~n7552 ;
  assign n7554 = ~n7511 & ~n7553 ;
  assign n7556 = ~n7510 & ~n7554 ;
  assign n7557 = ~n7555 & n7556 ;
  assign n7465 = ~n7460 & n7464 ;
  assign n7466 = ~n7459 & ~n7465 ;
  assign n7467 = ~n7423 & ~n7424 ;
  assign n7468 = ~n7428 & n7467 ;
  assign n7469 = n7428 & ~n7467 ;
  assign n7470 = ~n7468 & ~n7469 ;
  assign n7471 = n7466 & ~n7470 ;
  assign n7489 = n7484 & n7488 ;
  assign n7558 = ~n7471 & ~n7489 ;
  assign n7559 = ~n7557 & n7558 ;
  assign n7560 = ~n7466 & n7470 ;
  assign n7561 = n7404 & ~n7430 ;
  assign n7562 = ~n7560 & ~n7561 ;
  assign n7563 = ~n7559 & n7562 ;
  assign n7564 = n7439 & ~n7563 ;
  assign n7565 = n7323 & ~n7364 ;
  assign n7566 = ~n7433 & ~n7437 ;
  assign n7567 = ~n7565 & ~n7566 ;
  assign n7568 = ~n7564 & n7567 ;
  assign n7569 = n7373 & ~n7568 ;
  assign n7570 = ~n7256 & ~n7284 ;
  assign n7571 = ~n7367 & n7371 ;
  assign n7572 = ~n7570 & ~n7571 ;
  assign n7573 = ~n7569 & n7572 ;
  assign n7574 = ~n7285 & ~n7573 ;
  assign n7575 = n7267 & ~n7277 ;
  assign n7576 = ~n7276 & ~n7575 ;
  assign n7577 = ~n7001 & ~n7002 ;
  assign n7578 = ~n7025 & n7577 ;
  assign n7579 = n7025 & ~n7577 ;
  assign n7580 = ~n7578 & ~n7579 ;
  assign n7581 = ~n7576 & ~n7580 ;
  assign n7582 = n7576 & n7580 ;
  assign n7583 = ~n7056 & ~n7057 ;
  assign n7584 = ~n7102 & n7583 ;
  assign n7585 = n7102 & ~n7583 ;
  assign n7586 = ~n7584 & ~n7585 ;
  assign n7587 = ~n7582 & ~n7586 ;
  assign n7588 = ~n7581 & ~n7587 ;
  assign n7589 = ~n7109 & ~n7110 ;
  assign n7590 = n7114 & n7589 ;
  assign n7591 = ~n7114 & ~n7589 ;
  assign n7592 = ~n7590 & ~n7591 ;
  assign n7593 = ~n7588 & n7592 ;
  assign n7594 = ~n7264 & ~n7281 ;
  assign n7595 = ~n7263 & ~n7594 ;
  assign n7596 = ~n7581 & ~n7582 ;
  assign n7597 = ~n7586 & n7596 ;
  assign n7598 = n7586 & ~n7596 ;
  assign n7599 = ~n7597 & ~n7598 ;
  assign n7600 = ~n7595 & n7599 ;
  assign n7601 = ~n7593 & ~n7600 ;
  assign n7602 = n7574 & n7601 ;
  assign n7603 = n7588 & ~n7592 ;
  assign n7604 = n7595 & ~n7599 ;
  assign n7605 = ~n7593 & n7604 ;
  assign n7606 = ~n7603 & ~n7605 ;
  assign n7607 = ~n7602 & n7606 ;
  assign n7608 = ~n7116 & n7120 ;
  assign n7609 = ~n7047 & ~n7608 ;
  assign n7610 = n6972 & n7609 ;
  assign n7611 = ~n7607 & n7610 ;
  assign n7612 = n6782 & n7611 ;
  assign n7613 = n5854 & n7612 ;
  assign n7614 = n6314 & n7613 ;
  assign n7615 = ~n5440 & ~n5442 ;
  assign n7616 = ~n5095 & ~n5247 ;
  assign n7617 = ~n5443 & n7616 ;
  assign n7618 = ~n7615 & ~n7617 ;
  assign n7619 = n5853 & ~n7618 ;
  assign n7145 = n5643 & ~n5645 ;
  assign n7146 = ~n5852 & n7145 ;
  assign n7620 = ~n5648 & n5851 ;
  assign n7621 = ~n7146 & ~n7620 ;
  assign n7622 = ~n7619 & n7621 ;
  assign n7623 = ~n7614 & n7622 ;
  assign n7624 = ~n7144 & n7623 ;
  assign n7634 = ~\P1_P1_Address_reg[26]/NET0131  & ~\P1_P1_Address_reg[27]/NET0131  ;
  assign n7635 = ~\P1_P1_Address_reg[28]/NET0131  & ~\P1_P1_Address_reg[2]/NET0131  ;
  assign n7641 = n7634 & n7635 ;
  assign n7632 = ~\P1_P1_Address_reg[22]/NET0131  & ~\P1_P1_Address_reg[23]/NET0131  ;
  assign n7633 = ~\P1_P1_Address_reg[24]/NET0131  & ~\P1_P1_Address_reg[25]/NET0131  ;
  assign n7642 = n7632 & n7633 ;
  assign n7648 = n7641 & n7642 ;
  assign n7638 = ~\P1_P1_Address_reg[7]/NET0131  & ~\P1_P1_Address_reg[8]/NET0131  ;
  assign n7639 = ~\P1_P1_Address_reg[9]/NET0131  & n7638 ;
  assign n7636 = ~\P1_P1_Address_reg[3]/NET0131  & ~\P1_P1_Address_reg[4]/NET0131  ;
  assign n7637 = ~\P1_P1_Address_reg[5]/NET0131  & ~\P1_P1_Address_reg[6]/NET0131  ;
  assign n7640 = n7636 & n7637 ;
  assign n7649 = n7639 & n7640 ;
  assign n7650 = n7648 & n7649 ;
  assign n7625 = ~\P1_P1_Address_reg[0]/NET0131  & ~\P1_P1_Address_reg[10]/NET0131  ;
  assign n7626 = ~\P1_P1_Address_reg[11]/NET0131  & ~\P1_P1_Address_reg[12]/NET0131  ;
  assign n7627 = ~\P1_P1_Address_reg[13]/NET0131  & ~\P1_P1_Address_reg[14]/NET0131  ;
  assign n7645 = n7626 & n7627 ;
  assign n7646 = n7625 & n7645 ;
  assign n7630 = ~\P1_P1_Address_reg[19]/NET0131  & ~\P1_P1_Address_reg[1]/NET0131  ;
  assign n7631 = ~\P1_P1_Address_reg[20]/NET0131  & ~\P1_P1_Address_reg[21]/NET0131  ;
  assign n7643 = n7630 & n7631 ;
  assign n7628 = ~\P1_P1_Address_reg[15]/NET0131  & ~\P1_P1_Address_reg[16]/NET0131  ;
  assign n7629 = ~\P1_P1_Address_reg[17]/NET0131  & ~\P1_P1_Address_reg[18]/NET0131  ;
  assign n7644 = n7628 & n7629 ;
  assign n7647 = n7643 & n7644 ;
  assign n7651 = n7646 & n7647 ;
  assign n7652 = n7650 & n7651 ;
  assign n7653 = \P1_P1_Address_reg[29]/NET0131  & ~n7652 ;
  assign n7654 = \P4_datao_reg[19]/NET0131  & n4356 ;
  assign n7655 = \P4_datao_reg[18]/NET0131  & n4360 ;
  assign n7656 = ~n7654 & ~n7655 ;
  assign n7657 = \P4_datao_reg[15]/NET0131  & n4390 ;
  assign n7658 = \P4_datao_reg[14]/NET0131  & n4388 ;
  assign n7659 = ~n7657 & ~n7658 ;
  assign n7660 = n7656 & ~n7659 ;
  assign n7661 = ~n7656 & n7659 ;
  assign n7662 = ~n7660 & ~n7661 ;
  assign n7663 = \P4_datao_reg[27]/NET0131  & n4548 ;
  assign n7664 = \P4_datao_reg[26]/NET0131  & n4552 ;
  assign n7665 = ~n7663 & ~n7664 ;
  assign n7666 = \P4_datao_reg[25]/NET0131  & n4407 ;
  assign n7667 = \P4_datao_reg[24]/NET0131  & n4405 ;
  assign n7668 = ~n7666 & ~n7667 ;
  assign n7669 = n4417 & ~n7668 ;
  assign n7670 = ~n4417 & n7668 ;
  assign n7671 = ~n7669 & ~n7670 ;
  assign n7672 = \P4_datao_reg[11]/NET0131  & n4575 ;
  assign n7673 = \P4_datao_reg[10]/NET0131  & n4580 ;
  assign n7674 = ~n7672 & ~n7673 ;
  assign n7675 = n7671 & ~n7674 ;
  assign n7676 = ~n7671 & n7674 ;
  assign n7677 = ~n7675 & ~n7676 ;
  assign n7678 = n7665 & n7677 ;
  assign n7679 = ~n7665 & ~n7677 ;
  assign n7680 = ~n7678 & ~n7679 ;
  assign n7681 = n7662 & ~n7680 ;
  assign n7682 = ~n7662 & n7680 ;
  assign n7683 = ~n7681 & ~n7682 ;
  assign n7684 = \P4_datao_reg[21]/NET0131  & n4435 ;
  assign n7685 = \P4_datao_reg[20]/NET0131  & n4439 ;
  assign n7686 = ~n7684 & ~n7685 ;
  assign n7687 = \P4_datao_reg[9]/NET0131  & n4562 ;
  assign n7688 = \P4_datao_reg[8]/NET0131  & n4566 ;
  assign n7689 = ~n7687 & ~n7688 ;
  assign n7690 = \P4_datao_reg[17]/NET0131  & n4376 ;
  assign n7691 = \P4_datao_reg[16]/NET0131  & n4374 ;
  assign n7692 = ~n7690 & ~n7691 ;
  assign n7693 = n7689 & ~n7692 ;
  assign n7694 = ~n7689 & n7692 ;
  assign n7695 = ~n7693 & ~n7694 ;
  assign n7696 = ~n4447 & ~n4807 ;
  assign n7697 = n4447 & n4807 ;
  assign n7698 = ~n7696 & ~n7697 ;
  assign n7699 = n7695 & ~n7698 ;
  assign n7700 = ~n7695 & n7698 ;
  assign n7701 = ~n7699 & ~n7700 ;
  assign n7702 = n7686 & n7701 ;
  assign n7703 = ~n7686 & ~n7701 ;
  assign n7704 = ~n7702 & ~n7703 ;
  assign n7705 = \din[31]_pad  & sel_pad ;
  assign n7706 = \P4_datao_reg[1]/NET0131  & n5730 ;
  assign n7707 = ~n5727 & n7705 ;
  assign n7708 = \P4_datao_reg[0]/NET0131  & ~n7707 ;
  assign n7709 = ~n7706 & ~n7708 ;
  assign n7710 = n7705 & ~n7709 ;
  assign n7711 = n5728 & n7708 ;
  assign n7712 = ~n7705 & ~n7706 ;
  assign n7713 = ~n7711 & n7712 ;
  assign n7714 = ~n7710 & ~n7713 ;
  assign n7715 = n7704 & ~n7714 ;
  assign n7716 = ~n7704 & n7714 ;
  assign n7717 = ~n7715 & ~n7716 ;
  assign n7718 = n7683 & ~n7717 ;
  assign n7719 = ~n7683 & n7717 ;
  assign n7720 = ~n7718 & ~n7719 ;
  assign n7721 = ~n5718 & ~n5848 ;
  assign n7722 = ~n5717 & ~n7721 ;
  assign n7723 = ~n5775 & ~n5800 ;
  assign n7724 = ~n5774 & ~n7723 ;
  assign n7725 = ~n7722 & n7724 ;
  assign n7726 = n7722 & ~n7724 ;
  assign n7727 = ~n7725 & ~n7726 ;
  assign n7728 = ~n5710 & ~n5713 ;
  assign n7729 = ~n5709 & ~n7728 ;
  assign n7730 = n4431 & ~n7729 ;
  assign n7731 = ~n4431 & n7729 ;
  assign n7732 = ~n7730 & ~n7731 ;
  assign n7733 = \P4_datao_reg[3]/NET0131  & n5363 ;
  assign n7734 = \P4_datao_reg[2]/NET0131  & n5527 ;
  assign n7735 = ~n7733 & ~n7734 ;
  assign n7736 = \P4_datao_reg[5]/NET0131  & n4815 ;
  assign n7737 = \P4_datao_reg[4]/NET0131  & n4813 ;
  assign n7738 = ~n7736 & ~n7737 ;
  assign n7739 = n4351 & ~n5483 ;
  assign n7740 = ~n4351 & n5483 ;
  assign n7741 = ~n7739 & ~n7740 ;
  assign n7742 = n7738 & n7741 ;
  assign n7743 = ~n7738 & ~n7741 ;
  assign n7744 = ~n7742 & ~n7743 ;
  assign n7745 = n7735 & ~n7744 ;
  assign n7746 = ~n7735 & n7744 ;
  assign n7747 = ~n7745 & ~n7746 ;
  assign n7748 = n7732 & n7747 ;
  assign n7749 = ~n7732 & ~n7747 ;
  assign n7750 = ~n7748 & ~n7749 ;
  assign n7751 = n7727 & ~n7750 ;
  assign n7752 = ~n7727 & n7750 ;
  assign n7753 = ~n7751 & ~n7752 ;
  assign n7754 = n7720 & n7753 ;
  assign n7755 = ~n7720 & ~n7753 ;
  assign n7756 = ~n7754 & ~n7755 ;
  assign n7757 = ~n5658 & ~n5672 ;
  assign n7758 = ~n5671 & ~n7757 ;
  assign n7759 = ~n5789 & ~n5797 ;
  assign n7760 = ~n5790 & ~n7759 ;
  assign n7761 = ~n5814 & ~n5817 ;
  assign n7762 = ~n5813 & ~n7761 ;
  assign n7763 = n4352 & ~n7762 ;
  assign n7764 = ~n4352 & n7762 ;
  assign n7765 = ~n7763 & ~n7764 ;
  assign n7766 = \P4_datao_reg[13]/NET0131  & n4525 ;
  assign n7767 = \P4_datao_reg[12]/NET0131  & n4523 ;
  assign n7768 = ~n7766 & ~n7767 ;
  assign n7769 = n4398 & ~n7768 ;
  assign n7770 = ~n4398 & n7768 ;
  assign n7771 = ~n7769 & ~n7770 ;
  assign n7772 = n7765 & ~n7771 ;
  assign n7773 = ~n7765 & n7771 ;
  assign n7774 = ~n7772 & ~n7773 ;
  assign n7775 = n7760 & ~n7774 ;
  assign n7776 = ~n7760 & n7774 ;
  assign n7777 = ~n7775 & ~n7776 ;
  assign n7778 = \P4_datao_reg[29]/NET0131  & n4337 ;
  assign n7779 = \P4_datao_reg[28]/NET0131  & n4335 ;
  assign n7780 = ~n7778 & ~n7779 ;
  assign n7781 = n4328 & ~n7780 ;
  assign n7782 = ~n4328 & n7780 ;
  assign n7783 = ~n7781 & ~n7782 ;
  assign n7784 = n4399 & ~n7783 ;
  assign n7785 = ~n4399 & n7783 ;
  assign n7786 = ~n7784 & ~n7785 ;
  assign n7787 = ~n5755 & ~n5768 ;
  assign n7788 = ~n5769 & ~n7787 ;
  assign n7789 = ~n5827 & ~n5832 ;
  assign n7790 = ~n5833 & ~n7789 ;
  assign n7791 = n4368 & ~n7790 ;
  assign n7792 = ~n4368 & n7790 ;
  assign n7793 = ~n7791 & ~n7792 ;
  assign n7794 = n7788 & ~n7793 ;
  assign n7795 = ~n7788 & n7793 ;
  assign n7796 = ~n7794 & ~n7795 ;
  assign n7797 = n7786 & n7796 ;
  assign n7798 = ~n7786 & ~n7796 ;
  assign n7799 = ~n7797 & ~n7798 ;
  assign n7800 = ~n5824 & ~n5837 ;
  assign n7801 = ~n5823 & ~n7800 ;
  assign n7802 = ~n5702 & ~n5705 ;
  assign n7803 = ~n5701 & ~n7802 ;
  assign n7804 = n7801 & ~n7803 ;
  assign n7805 = ~n7801 & n7803 ;
  assign n7806 = ~n7804 & ~n7805 ;
  assign n7807 = \P4_datao_reg[23]/NET0131  & n4507 ;
  assign n7808 = \P4_datao_reg[22]/NET0131  & n4511 ;
  assign n7809 = ~n7807 & ~n7808 ;
  assign n7810 = n4579 & ~n7809 ;
  assign n7811 = ~n4579 & n7809 ;
  assign n7812 = ~n7810 & ~n7811 ;
  assign n7813 = ~n5682 & ~n5695 ;
  assign n7814 = ~n5696 & ~n7813 ;
  assign n7815 = \P4_datao_reg[31]/NET0131  & n4343 ;
  assign n7816 = ~\din[1]_pad  & n7815 ;
  assign n7817 = \P4_datao_reg[30]/NET0131  & n7011 ;
  assign n7818 = n4329 & ~n7815 ;
  assign n7819 = ~n7817 & n7818 ;
  assign n7820 = ~n7816 & ~n7819 ;
  assign n7821 = n7814 & ~n7820 ;
  assign n7822 = ~n7814 & n7820 ;
  assign n7823 = ~n7821 & ~n7822 ;
  assign n7824 = n7812 & n7823 ;
  assign n7825 = ~n7812 & ~n7823 ;
  assign n7826 = ~n7824 & ~n7825 ;
  assign n7827 = ~n5731 & n7705 ;
  assign n7828 = ~\din[17]_pad  & n7827 ;
  assign n7829 = n4382 & ~n7827 ;
  assign n7830 = ~n7828 & ~n7829 ;
  assign n7831 = n7826 & ~n7830 ;
  assign n7832 = ~n7826 & n7830 ;
  assign n7833 = ~n7831 & ~n7832 ;
  assign n7834 = n7806 & ~n7833 ;
  assign n7835 = ~n7806 & n7833 ;
  assign n7836 = ~n7834 & ~n7835 ;
  assign n7837 = n7799 & ~n7836 ;
  assign n7838 = ~n7799 & n7836 ;
  assign n7839 = ~n7837 & ~n7838 ;
  assign n7840 = n7777 & n7839 ;
  assign n7841 = ~n7777 & ~n7839 ;
  assign n7842 = ~n7840 & ~n7841 ;
  assign n7843 = n7758 & ~n7842 ;
  assign n7844 = ~n7758 & n7842 ;
  assign n7845 = ~n7843 & ~n7844 ;
  assign n7846 = \P4_datao_reg[7]/NET0131  & n4421 ;
  assign n7847 = \P4_datao_reg[6]/NET0131  & n4460 ;
  assign n7848 = ~n7846 & ~n7847 ;
  assign n7849 = ~n5724 & ~n5803 ;
  assign n7850 = ~n5725 & ~n7849 ;
  assign n7851 = n7848 & ~n7850 ;
  assign n7852 = ~n7848 & n7850 ;
  assign n7853 = ~n7851 & ~n7852 ;
  assign n7854 = ~n5738 & ~n5746 ;
  assign n7855 = ~n5739 & ~n7854 ;
  assign n7856 = n7853 & ~n7855 ;
  assign n7857 = ~n7853 & n7855 ;
  assign n7858 = ~n7856 & ~n7857 ;
  assign n7859 = ~n5842 & ~n5845 ;
  assign n7860 = ~n5841 & ~n7859 ;
  assign n7861 = n7858 & ~n7860 ;
  assign n7862 = ~n7858 & n7860 ;
  assign n7863 = ~n7861 & ~n7862 ;
  assign n7864 = n7845 & ~n7863 ;
  assign n7865 = ~n7845 & n7863 ;
  assign n7866 = ~n7864 & ~n7865 ;
  assign n7867 = n7756 & n7866 ;
  assign n7868 = ~n7756 & ~n7866 ;
  assign n7869 = ~n7867 & ~n7868 ;
  assign n7870 = ~n7653 & ~n7869 ;
  assign n7871 = ~n7624 & n7870 ;
  assign n7872 = ~n7653 & n7869 ;
  assign n7873 = n7624 & n7872 ;
  assign n7874 = ~n7871 & ~n7873 ;
  assign n7996 = ~n7121 & ~n7608 ;
  assign n7997 = ~n7607 & ~n7996 ;
  assign n7998 = n7607 & n7996 ;
  assign n7999 = ~n7997 & ~n7998 ;
  assign n8000 = ~n7653 & ~n7999 ;
  assign n8001 = \P1_buf1_reg[13]/NET0131  & n7653 ;
  assign n8002 = ~n7600 & ~n7604 ;
  assign n8004 = n7574 & n8002 ;
  assign n8003 = ~n7574 & ~n8002 ;
  assign n8005 = ~n7653 & ~n8003 ;
  assign n8006 = ~n8004 & n8005 ;
  assign n8007 = ~n8001 & ~n8006 ;
  assign n7876 = n7515 & n7524 ;
  assign n7877 = n7549 & ~n7876 ;
  assign n7878 = ~n7515 & ~n7524 ;
  assign n7879 = ~n7511 & ~n7878 ;
  assign n7880 = ~n7877 & n7879 ;
  assign n7881 = ~n7510 & ~n7880 ;
  assign n7882 = ~n7489 & ~n7881 ;
  assign n7883 = ~n7555 & ~n7560 ;
  assign n7884 = ~n7882 & n7883 ;
  assign n7885 = ~n7471 & ~n7884 ;
  assign n7958 = n7439 & n7885 ;
  assign n7959 = ~n7561 & ~n7566 ;
  assign n7960 = ~n7438 & ~n7959 ;
  assign n7961 = ~n7958 & ~n7960 ;
  assign n7976 = n7373 & ~n7961 ;
  assign n7977 = ~n7372 & n7565 ;
  assign n7978 = ~n7571 & ~n7977 ;
  assign n7979 = ~n7976 & n7978 ;
  assign n7986 = ~n7285 & ~n7600 ;
  assign n7987 = ~n7979 & n7986 ;
  assign n7988 = ~n7570 & ~n7604 ;
  assign n7989 = ~n7600 & ~n7988 ;
  assign n7990 = ~n7987 & ~n7989 ;
  assign n7991 = ~n7593 & ~n7603 ;
  assign n7992 = ~n7990 & ~n7991 ;
  assign n7993 = n7990 & n7991 ;
  assign n7994 = ~n7992 & ~n7993 ;
  assign n7995 = ~n7653 & ~n7994 ;
  assign n7975 = ~\P1_buf1_reg[12]/NET0131  & n7653 ;
  assign n7980 = ~n7285 & ~n7570 ;
  assign n7982 = n7979 & n7980 ;
  assign n7981 = ~n7979 & ~n7980 ;
  assign n7983 = ~n7653 & ~n7981 ;
  assign n7984 = ~n7982 & n7983 ;
  assign n7985 = ~n7975 & ~n7984 ;
  assign n7967 = ~\P1_buf1_reg[11]/NET0131  & n7653 ;
  assign n7968 = ~n7372 & ~n7571 ;
  assign n7969 = ~n7365 & ~n7568 ;
  assign n7971 = ~n7968 & n7969 ;
  assign n7970 = n7968 & ~n7969 ;
  assign n7972 = ~n7653 & ~n7970 ;
  assign n7973 = ~n7971 & n7972 ;
  assign n7974 = ~n7967 & ~n7973 ;
  assign n7956 = \P1_buf1_reg[10]/NET0131  & n7653 ;
  assign n7957 = ~n7365 & ~n7565 ;
  assign n7963 = ~n7957 & n7961 ;
  assign n7962 = n7957 & ~n7961 ;
  assign n7964 = ~n7653 & ~n7962 ;
  assign n7965 = ~n7963 & n7964 ;
  assign n7966 = ~n7956 & ~n7965 ;
  assign n7948 = ~\P1_buf1_reg[9]/NET0131  & n7653 ;
  assign n7949 = ~n7438 & ~n7566 ;
  assign n7950 = ~n7431 & ~n7563 ;
  assign n7952 = ~n7949 & n7950 ;
  assign n7951 = n7949 & ~n7950 ;
  assign n7953 = ~n7653 & ~n7951 ;
  assign n7954 = ~n7952 & n7953 ;
  assign n7955 = ~n7948 & ~n7954 ;
  assign n7875 = \P1_buf1_reg[8]/NET0131  & n7653 ;
  assign n7886 = ~n7431 & ~n7561 ;
  assign n7888 = n7885 & n7886 ;
  assign n7887 = ~n7885 & ~n7886 ;
  assign n7889 = ~n7653 & ~n7887 ;
  assign n7890 = ~n7888 & n7889 ;
  assign n7891 = ~n7875 & ~n7890 ;
  assign n7892 = ~\P1_buf1_reg[7]/NET0131  & n7653 ;
  assign n7893 = ~n7471 & ~n7560 ;
  assign n7894 = ~n7489 & ~n7557 ;
  assign n7896 = ~n7893 & n7894 ;
  assign n7895 = n7893 & ~n7894 ;
  assign n7897 = ~n7653 & ~n7895 ;
  assign n7898 = ~n7896 & n7897 ;
  assign n7899 = ~n7892 & ~n7898 ;
  assign n7900 = ~\P1_buf1_reg[6]/NET0131  & n7653 ;
  assign n7901 = ~n7489 & ~n7555 ;
  assign n7903 = n7881 & n7901 ;
  assign n7902 = ~n7881 & ~n7901 ;
  assign n7904 = ~n7653 & ~n7902 ;
  assign n7905 = ~n7903 & n7904 ;
  assign n7906 = ~n7900 & ~n7905 ;
  assign n7934 = \P1_buf1_reg[4]/NET0131  & n7653 ;
  assign n7935 = ~n7876 & ~n7878 ;
  assign n7937 = ~n7549 & n7935 ;
  assign n7936 = n7549 & ~n7935 ;
  assign n7938 = ~n7653 & ~n7936 ;
  assign n7939 = ~n7937 & n7938 ;
  assign n7940 = ~n7934 & ~n7939 ;
  assign n7927 = \P1_buf1_reg[5]/NET0131  & n7653 ;
  assign n7928 = ~n7510 & ~n7511 ;
  assign n7930 = n7553 & ~n7928 ;
  assign n7929 = ~n7553 & n7928 ;
  assign n7931 = ~n7653 & ~n7929 ;
  assign n7932 = ~n7930 & n7931 ;
  assign n7933 = ~n7927 & ~n7932 ;
  assign n7907 = \P1_buf1_reg[3]/NET0131  & n7653 ;
  assign n7908 = ~n7533 & ~n7548 ;
  assign n7910 = ~n7546 & n7908 ;
  assign n7909 = n7546 & ~n7908 ;
  assign n7911 = ~n7653 & ~n7909 ;
  assign n7912 = ~n7910 & n7911 ;
  assign n7913 = ~n7907 & ~n7912 ;
  assign n7941 = ~\P1_buf1_reg[2]/NET0131  & n7653 ;
  assign n7942 = ~n7540 & ~n7541 ;
  assign n7944 = n7544 & ~n7942 ;
  assign n7943 = ~n7544 & n7942 ;
  assign n7945 = ~n7653 & ~n7943 ;
  assign n7946 = ~n7944 & n7945 ;
  assign n7947 = ~n7941 & ~n7946 ;
  assign n7921 = \P1_buf1_reg[0]/NET0131  & n7653 ;
  assign n7922 = \P4_datao_reg[0]/NET0131  & n4343 ;
  assign n7923 = ~n7653 & n7922 ;
  assign n7924 = ~n7921 & ~n7923 ;
  assign n7914 = ~\P1_buf1_reg[1]/NET0131  & n7653 ;
  assign n7915 = \P4_datao_reg[0]/NET0131  & n4329 ;
  assign n7916 = n7542 & ~n7915 ;
  assign n7917 = ~n7542 & n7915 ;
  assign n7918 = ~n7916 & ~n7917 ;
  assign n7919 = ~n7653 & n7918 ;
  assign n7920 = ~n7914 & ~n7919 ;
  assign n7925 = \P1_buf1_reg[14]/NET0131  & n7653 ;
  assign n7926 = \P1_buf1_reg[15]/NET0131  & n7653 ;
  assign n8008 = ~n7925 & ~n7926 ;
  assign n8009 = ~n7920 & n8008 ;
  assign n8010 = n7924 & n8009 ;
  assign n8011 = ~n7947 & n8010 ;
  assign n8012 = n7913 & n8011 ;
  assign n8013 = n7933 & n8012 ;
  assign n8014 = n7940 & n8013 ;
  assign n8015 = ~n7906 & n8014 ;
  assign n8016 = ~n7899 & n8015 ;
  assign n8017 = n7891 & n8016 ;
  assign n8018 = ~n7955 & n8017 ;
  assign n8019 = n7966 & n8018 ;
  assign n8020 = ~n7974 & n8019 ;
  assign n8021 = ~n7985 & n8020 ;
  assign n8022 = ~n7995 & n8021 ;
  assign n8023 = n8007 & n8022 ;
  assign n8024 = ~n8000 & n8023 ;
  assign n8025 = ~n7874 & ~n8024 ;
  assign n8026 = \P1_buf1_reg[16]/NET0131  & n7653 ;
  assign n8027 = ~n7593 & ~n7608 ;
  assign n8028 = n7987 & n8027 ;
  assign n8029 = n7989 & n8027 ;
  assign n8030 = n7603 & ~n7608 ;
  assign n8031 = ~n7121 & ~n8030 ;
  assign n8032 = ~n8029 & n8031 ;
  assign n8033 = ~n8028 & n8032 ;
  assign n8034 = ~n7046 & ~n7047 ;
  assign n8036 = ~n8033 & n8034 ;
  assign n8035 = n8033 & ~n8034 ;
  assign n8037 = ~n7653 & ~n8035 ;
  assign n8038 = ~n8036 & n8037 ;
  assign n8039 = ~n8026 & ~n8038 ;
  assign n8040 = n8025 & ~n8039 ;
  assign n8041 = \P1_buf1_reg[17]/NET0131  & n7653 ;
  assign n8042 = n7601 & n7609 ;
  assign n8043 = n7574 & n8042 ;
  assign n8044 = ~n7606 & n7609 ;
  assign n8045 = n7123 & ~n8044 ;
  assign n8046 = ~n8043 & n8045 ;
  assign n8047 = ~n6971 & ~n7126 ;
  assign n8049 = ~n8046 & n8047 ;
  assign n8048 = n8046 & ~n8047 ;
  assign n8050 = ~n7653 & ~n8048 ;
  assign n8051 = ~n8049 & n8050 ;
  assign n8052 = ~n8041 & ~n8051 ;
  assign n8053 = n8040 & ~n8052 ;
  assign n8054 = \P1_buf1_reg[18]/NET0131  & n7653 ;
  assign n8055 = ~n6971 & ~n7047 ;
  assign n8056 = ~n8031 & n8055 ;
  assign n8057 = ~n6971 & n7046 ;
  assign n8058 = ~n7126 & ~n8057 ;
  assign n8059 = ~n8056 & n8058 ;
  assign n8060 = n8027 & n8055 ;
  assign n8061 = ~n7990 & n8060 ;
  assign n8062 = n8059 & ~n8061 ;
  assign n8063 = ~n6869 & ~n7125 ;
  assign n8065 = ~n8062 & n8063 ;
  assign n8064 = n8062 & ~n8063 ;
  assign n8066 = ~n7653 & ~n8064 ;
  assign n8067 = ~n8065 & n8066 ;
  assign n8068 = ~n8054 & ~n8067 ;
  assign n8069 = n8053 & ~n8068 ;
  assign n8070 = \P1_buf1_reg[19]/NET0131  & n7653 ;
  assign n8071 = n7129 & ~n7611 ;
  assign n8072 = ~n6771 & ~n6780 ;
  assign n8074 = ~n8071 & n8072 ;
  assign n8073 = n8071 & ~n8072 ;
  assign n8075 = ~n7653 & ~n8073 ;
  assign n8076 = ~n8074 & n8075 ;
  assign n8077 = ~n8070 & ~n8076 ;
  assign n8078 = \P1_buf1_reg[20]/NET0131  & n7653 ;
  assign n8079 = ~n6673 & ~n6674 ;
  assign n8080 = ~n6780 & ~n6869 ;
  assign n8084 = ~n8033 & n8055 ;
  assign n8085 = n8080 & n8084 ;
  assign n8081 = ~n8058 & n8080 ;
  assign n8082 = ~n6780 & n7125 ;
  assign n8083 = ~n6771 & ~n8082 ;
  assign n8086 = ~n8081 & n8083 ;
  assign n8087 = ~n8085 & n8086 ;
  assign n8089 = ~n8079 & n8087 ;
  assign n8088 = n8079 & ~n8087 ;
  assign n8090 = ~n7653 & ~n8088 ;
  assign n8091 = ~n8089 & n8090 ;
  assign n8092 = ~n8078 & ~n8091 ;
  assign n8093 = ~n8077 & ~n8092 ;
  assign n8094 = n8069 & n8093 ;
  assign n8095 = \P1_buf1_reg[21]/NET0131  & n7653 ;
  assign n8096 = ~n6620 & ~n6776 ;
  assign n8098 = n6781 & n6972 ;
  assign n8099 = ~n8046 & n8098 ;
  assign n8097 = n6781 & ~n7128 ;
  assign n8100 = ~n6773 & ~n8097 ;
  assign n8101 = ~n8099 & n8100 ;
  assign n8103 = ~n8096 & n8101 ;
  assign n8102 = n8096 & ~n8101 ;
  assign n8104 = ~n7653 & ~n8102 ;
  assign n8105 = ~n8103 & n8104 ;
  assign n8106 = ~n8095 & ~n8105 ;
  assign n8107 = \P1_buf1_reg[22]/NET0131  & n7653 ;
  assign n8108 = ~n6627 & ~n6775 ;
  assign n8109 = ~n6620 & ~n6673 ;
  assign n8110 = ~n8083 & n8109 ;
  assign n8111 = ~n6620 & n6674 ;
  assign n8112 = ~n6776 & ~n8111 ;
  assign n8113 = ~n8110 & n8112 ;
  assign n8114 = n8080 & n8109 ;
  assign n8115 = ~n8062 & n8114 ;
  assign n8116 = n8113 & ~n8115 ;
  assign n8118 = ~n8108 & n8116 ;
  assign n8117 = n8108 & ~n8116 ;
  assign n8119 = ~n7653 & ~n8117 ;
  assign n8120 = ~n8118 & n8119 ;
  assign n8121 = ~n8107 & ~n8120 ;
  assign n8122 = ~n8106 & ~n8121 ;
  assign n8123 = n8094 & n8122 ;
  assign n8124 = \P1_buf1_reg[23]/NET0131  & n7653 ;
  assign n8125 = ~n6256 & ~n7134 ;
  assign n8126 = n6782 & ~n8071 ;
  assign n8127 = n6779 & ~n8126 ;
  assign n8129 = ~n8125 & n8127 ;
  assign n8128 = n8125 & ~n8127 ;
  assign n8130 = ~n7653 & ~n8128 ;
  assign n8131 = ~n8129 & n8130 ;
  assign n8132 = ~n8124 & ~n8131 ;
  assign n8133 = n8123 & ~n8132 ;
  assign n8134 = ~n8123 & n8132 ;
  assign n8135 = ~n8133 & ~n8134 ;
  assign n8136 = n4327 & ~n8135 ;
  assign n8137 = ~\P1_P1_InstQueueWr_Addr_reg[0]/NET0131  & ~\P1_P1_InstQueueWr_Addr_reg[1]/NET0131  ;
  assign n8138 = ~\P1_P1_InstQueueWr_Addr_reg[2]/NET0131  & n8137 ;
  assign n8139 = \P1_P1_InstQueueWr_Addr_reg[3]/NET0131  & n8138 ;
  assign n8140 = \P1_P1_InstQueueWr_Addr_reg[0]/NET0131  & \P1_P1_InstQueueWr_Addr_reg[1]/NET0131  ;
  assign n8141 = ~\P1_P1_InstQueueWr_Addr_reg[2]/NET0131  & n8140 ;
  assign n8142 = \P1_P1_InstQueueWr_Addr_reg[3]/NET0131  & n8141 ;
  assign n8143 = ~\P1_P1_InstQueueWr_Addr_reg[0]/NET0131  & \P1_P1_InstQueueWr_Addr_reg[1]/NET0131  ;
  assign n8144 = ~\P1_P1_InstQueueWr_Addr_reg[2]/NET0131  & n8143 ;
  assign n8145 = \P1_P1_InstQueueWr_Addr_reg[3]/NET0131  & n8144 ;
  assign n8146 = ~n8142 & ~n8145 ;
  assign n8147 = n7899 & ~n8146 ;
  assign n8148 = \P1_P1_InstQueue_reg[11][7]/NET0131  & ~n8142 ;
  assign n8149 = ~n8145 & n8148 ;
  assign n8150 = ~n8147 & ~n8149 ;
  assign n8151 = ~n4327 & n8150 ;
  assign n8152 = ~n8139 & ~n8151 ;
  assign n8153 = ~n8136 & n8152 ;
  assign n8154 = n8039 & n8052 ;
  assign n8155 = n8024 & n8154 ;
  assign n8156 = n8068 & n8155 ;
  assign n8157 = n8077 & n8156 ;
  assign n8158 = n8092 & n8106 ;
  assign n8159 = n8157 & n8158 ;
  assign n8160 = n8121 & n8132 ;
  assign n8161 = n8159 & n8160 ;
  assign n8162 = ~n7874 & ~n8161 ;
  assign n8163 = \P1_buf1_reg[24]/NET0131  & n7653 ;
  assign n8164 = ~n6285 & ~n7133 ;
  assign n8165 = ~n6256 & ~n6627 ;
  assign n8166 = ~n8112 & n8165 ;
  assign n8167 = ~n6256 & n6775 ;
  assign n8168 = ~n7134 & ~n8167 ;
  assign n8169 = ~n8166 & n8168 ;
  assign n8170 = ~n8087 & n8109 ;
  assign n8171 = n8165 & n8170 ;
  assign n8172 = n8169 & ~n8171 ;
  assign n8174 = ~n8164 & n8172 ;
  assign n8173 = n8164 & ~n8172 ;
  assign n8175 = ~n7653 & ~n8173 ;
  assign n8176 = ~n8174 & n8175 ;
  assign n8177 = ~n8163 & ~n8176 ;
  assign n8178 = n8162 & ~n8177 ;
  assign n8179 = \P1_buf1_reg[25]/NET0131  & n7653 ;
  assign n8180 = ~n6305 & ~n7139 ;
  assign n8181 = n6286 & ~n6778 ;
  assign n8182 = n7136 & ~n8181 ;
  assign n8183 = n6628 & ~n8101 ;
  assign n8184 = n6286 & n8183 ;
  assign n8185 = n8182 & ~n8184 ;
  assign n8187 = ~n8180 & n8185 ;
  assign n8186 = n8180 & ~n8185 ;
  assign n8188 = ~n7653 & ~n8186 ;
  assign n8189 = ~n8187 & n8188 ;
  assign n8190 = ~n8179 & ~n8189 ;
  assign n8191 = n8178 & ~n8190 ;
  assign n8192 = \P1_buf1_reg[26]/NET0131  & n7653 ;
  assign n8193 = ~n6312 & ~n7138 ;
  assign n8194 = ~n6285 & ~n6305 ;
  assign n8195 = ~n8168 & n8194 ;
  assign n8196 = ~n6305 & n7133 ;
  assign n8197 = ~n7139 & ~n8196 ;
  assign n8198 = ~n8195 & n8197 ;
  assign n8199 = n8165 & n8194 ;
  assign n8200 = ~n8116 & n8199 ;
  assign n8201 = n8198 & ~n8200 ;
  assign n8203 = ~n8193 & n8201 ;
  assign n8202 = n8193 & ~n8201 ;
  assign n8204 = ~n7653 & ~n8202 ;
  assign n8205 = ~n8203 & n8204 ;
  assign n8206 = ~n8192 & ~n8205 ;
  assign n8207 = n8191 & ~n8206 ;
  assign n8208 = \P1_buf1_reg[28]/NET0131  & n7653 ;
  assign n8209 = ~n5248 & n7138 ;
  assign n8210 = ~n7616 & ~n8209 ;
  assign n8211 = ~n5248 & ~n6312 ;
  assign n8213 = n8170 & n8199 ;
  assign n8212 = ~n8169 & n8194 ;
  assign n8214 = n8197 & ~n8212 ;
  assign n8215 = ~n8213 & n8214 ;
  assign n8216 = n8211 & ~n8215 ;
  assign n8217 = n8210 & ~n8216 ;
  assign n8218 = ~n5443 & ~n7615 ;
  assign n8220 = ~n8217 & n8218 ;
  assign n8219 = n8217 & ~n8218 ;
  assign n8221 = ~n7653 & ~n8219 ;
  assign n8222 = ~n8220 & n8221 ;
  assign n8223 = ~n8208 & ~n8222 ;
  assign n8224 = \P1_buf1_reg[27]/NET0131  & n7653 ;
  assign n8225 = ~n5248 & ~n7616 ;
  assign n8226 = n6314 & ~n8127 ;
  assign n8227 = n7142 & ~n8226 ;
  assign n8229 = ~n8225 & n8227 ;
  assign n8228 = n8225 & ~n8227 ;
  assign n8230 = ~n7653 & ~n8228 ;
  assign n8231 = ~n8229 & n8230 ;
  assign n8232 = ~n8224 & ~n8231 ;
  assign n8233 = ~n8223 & ~n8232 ;
  assign n8234 = n8207 & n8233 ;
  assign n8235 = \P1_buf1_reg[29]/NET0131  & n7653 ;
  assign n8236 = ~n5646 & ~n7145 ;
  assign n8239 = n6313 & ~n8182 ;
  assign n8240 = ~n7141 & ~n8239 ;
  assign n8241 = n5444 & ~n8240 ;
  assign n8237 = n5444 & n6314 ;
  assign n8238 = n8183 & n8237 ;
  assign n8242 = n7618 & ~n8238 ;
  assign n8243 = ~n8241 & n8242 ;
  assign n8245 = ~n8236 & n8243 ;
  assign n8244 = n8236 & ~n8243 ;
  assign n8246 = ~n7653 & ~n8244 ;
  assign n8247 = ~n8245 & n8246 ;
  assign n8248 = ~n8235 & ~n8247 ;
  assign n8249 = \P1_buf1_reg[30]/NET0131  & n7653 ;
  assign n8250 = ~n5852 & ~n7620 ;
  assign n8251 = ~n8059 & n8114 ;
  assign n8252 = n8113 & ~n8251 ;
  assign n8253 = n8199 & ~n8252 ;
  assign n8254 = n8198 & ~n8253 ;
  assign n8255 = ~n5443 & ~n5646 ;
  assign n8256 = n8211 & n8255 ;
  assign n8257 = ~n8254 & n8256 ;
  assign n8260 = n8061 & n8114 ;
  assign n8261 = n8199 & n8260 ;
  assign n8262 = n8256 & n8261 ;
  assign n8258 = ~n7615 & n8210 ;
  assign n8259 = n8255 & ~n8258 ;
  assign n8263 = ~n7145 & ~n8259 ;
  assign n8264 = ~n8262 & n8263 ;
  assign n8265 = ~n8257 & n8264 ;
  assign n8267 = ~n8250 & n8265 ;
  assign n8266 = n8250 & ~n8265 ;
  assign n8268 = ~n7653 & ~n8266 ;
  assign n8269 = ~n8267 & n8268 ;
  assign n8270 = ~n8249 & ~n8269 ;
  assign n8271 = ~n8248 & ~n8270 ;
  assign n8272 = n8234 & n8271 ;
  assign n8273 = ~n7874 & ~n8272 ;
  assign n8274 = n7874 & n8272 ;
  assign n8275 = ~n8273 & ~n8274 ;
  assign n8276 = n8139 & ~n8275 ;
  assign n8277 = \P1_P1_DataWidth_reg[1]/NET0131  & ~n8276 ;
  assign n8278 = ~n8153 & n8277 ;
  assign n8279 = ~\P1_P1_DataWidth_reg[1]/NET0131  & n8150 ;
  assign n8280 = \P1_P1_State2_reg[1]/NET0131  & ~\P1_P1_State2_reg[2]/NET0131  ;
  assign n8281 = ~\P1_P1_State2_reg[3]/NET0131  & n8280 ;
  assign n8282 = ~\P1_P1_State2_reg[0]/NET0131  & n8281 ;
  assign n8283 = ~n8279 & n8282 ;
  assign n8284 = ~n8278 & n8283 ;
  assign n8285 = ~\P1_P1_State2_reg[1]/NET0131  & \P1_P1_State2_reg[2]/NET0131  ;
  assign n8286 = ~\P1_P1_State2_reg[3]/NET0131  & n8285 ;
  assign n8287 = ~\P1_P1_State2_reg[0]/NET0131  & n8286 ;
  assign n8288 = ~n8150 & n8287 ;
  assign n8289 = \P1_P1_InstQueueRd_Addr_reg[1]/NET0131  & \P1_P1_InstQueueRd_Addr_reg[2]/NET0131  ;
  assign n8290 = \P1_P1_InstQueueRd_Addr_reg[3]/NET0131  & n8289 ;
  assign n8291 = ~\P1_P1_InstQueueRd_Addr_reg[0]/NET0131  & n8290 ;
  assign n8292 = \P1_P1_InstQueue_reg[14][7]/NET0131  & n8291 ;
  assign n8293 = ~\P1_P1_InstQueueRd_Addr_reg[0]/NET0131  & ~\P1_P1_InstQueueRd_Addr_reg[1]/NET0131  ;
  assign n8294 = \P1_P1_InstQueueRd_Addr_reg[2]/NET0131  & ~\P1_P1_InstQueueRd_Addr_reg[3]/NET0131  ;
  assign n8295 = n8293 & n8294 ;
  assign n8296 = \P1_P1_InstQueue_reg[4][7]/NET0131  & n8295 ;
  assign n8297 = \P1_P1_InstQueueRd_Addr_reg[0]/NET0131  & ~\P1_P1_InstQueueRd_Addr_reg[1]/NET0131  ;
  assign n8298 = ~\P1_P1_InstQueueRd_Addr_reg[2]/NET0131  & ~\P1_P1_InstQueueRd_Addr_reg[3]/NET0131  ;
  assign n8299 = n8297 & n8298 ;
  assign n8300 = \P1_P1_InstQueue_reg[1][7]/NET0131  & n8299 ;
  assign n8331 = ~n8296 & ~n8300 ;
  assign n8301 = ~\P1_P1_InstQueueRd_Addr_reg[0]/NET0131  & \P1_P1_InstQueueRd_Addr_reg[1]/NET0131  ;
  assign n8302 = ~\P1_P1_InstQueueRd_Addr_reg[2]/NET0131  & \P1_P1_InstQueueRd_Addr_reg[3]/NET0131  ;
  assign n8303 = n8301 & n8302 ;
  assign n8304 = \P1_P1_InstQueue_reg[10][7]/NET0131  & n8303 ;
  assign n8305 = n8293 & n8302 ;
  assign n8306 = \P1_P1_InstQueue_reg[8][7]/NET0131  & n8305 ;
  assign n8332 = ~n8304 & ~n8306 ;
  assign n8341 = n8331 & n8332 ;
  assign n8342 = ~n8292 & n8341 ;
  assign n8320 = \P1_P1_InstQueueRd_Addr_reg[2]/NET0131  & \P1_P1_InstQueueRd_Addr_reg[3]/NET0131  ;
  assign n8329 = n8293 & n8320 ;
  assign n8330 = \P1_P1_InstQueue_reg[12][7]/NET0131  & n8329 ;
  assign n8325 = n8297 & n8302 ;
  assign n8326 = \P1_P1_InstQueue_reg[9][7]/NET0131  & n8325 ;
  assign n8327 = n8297 & n8320 ;
  assign n8328 = \P1_P1_InstQueue_reg[13][7]/NET0131  & n8327 ;
  assign n8337 = ~n8326 & ~n8328 ;
  assign n8338 = ~n8330 & n8337 ;
  assign n8316 = n8294 & n8301 ;
  assign n8317 = \P1_P1_InstQueue_reg[6][7]/NET0131  & n8316 ;
  assign n8311 = \P1_P1_InstQueueRd_Addr_reg[0]/NET0131  & \P1_P1_InstQueueRd_Addr_reg[1]/NET0131  ;
  assign n8318 = n8294 & n8311 ;
  assign n8319 = \P1_P1_InstQueue_reg[7][7]/NET0131  & n8318 ;
  assign n8335 = ~n8317 & ~n8319 ;
  assign n8321 = n8311 & n8320 ;
  assign n8322 = \P1_P1_InstQueue_reg[15][7]/NET0131  & n8321 ;
  assign n8323 = n8298 & n8311 ;
  assign n8324 = \P1_P1_InstQueue_reg[3][7]/NET0131  & n8323 ;
  assign n8336 = ~n8322 & ~n8324 ;
  assign n8339 = n8335 & n8336 ;
  assign n8307 = n8294 & n8297 ;
  assign n8308 = \P1_P1_InstQueue_reg[5][7]/NET0131  & n8307 ;
  assign n8309 = n8293 & n8298 ;
  assign n8310 = \P1_P1_InstQueue_reg[0][7]/NET0131  & n8309 ;
  assign n8333 = ~n8308 & ~n8310 ;
  assign n8312 = n8302 & n8311 ;
  assign n8313 = \P1_P1_InstQueue_reg[11][7]/NET0131  & n8312 ;
  assign n8314 = n8298 & n8301 ;
  assign n8315 = \P1_P1_InstQueue_reg[2][7]/NET0131  & n8314 ;
  assign n8334 = ~n8313 & ~n8315 ;
  assign n8340 = n8333 & n8334 ;
  assign n8343 = n8339 & n8340 ;
  assign n8344 = n8338 & n8343 ;
  assign n8345 = n8342 & n8344 ;
  assign n8346 = n8142 & ~n8345 ;
  assign n8347 = ~n8148 & ~n8346 ;
  assign n8348 = ~\P1_P1_State2_reg[1]/NET0131  & ~\P1_P1_State2_reg[2]/NET0131  ;
  assign n8349 = \P1_P1_State2_reg[3]/NET0131  & n8348 ;
  assign n8350 = ~\P1_P1_State2_reg[0]/NET0131  & n8349 ;
  assign n8351 = ~n8347 & n8350 ;
  assign n8356 = ~\P1_P1_State2_reg[0]/NET0131  & ~\P1_P1_State2_reg[3]/NET0131  ;
  assign n8357 = n8348 & n8356 ;
  assign n8358 = \P1_P1_State2_reg[0]/NET0131  & n8348 ;
  assign n8359 = ~\P1_P1_State2_reg[3]/NET0131  & n8358 ;
  assign n8360 = ~n8357 & ~n8359 ;
  assign n8361 = \P1_P1_State2_reg[0]/NET0131  & n8349 ;
  assign n8362 = n8360 & ~n8361 ;
  assign n8354 = \P1_P1_State2_reg[0]/NET0131  & ~\P1_P1_State2_reg[3]/NET0131  ;
  assign n8363 = n8280 & n8354 ;
  assign n8352 = \P1_P1_State2_reg[1]/NET0131  & \P1_P1_State2_reg[2]/NET0131  ;
  assign n8353 = ~\P1_P1_State2_reg[3]/NET0131  & n8352 ;
  assign n8355 = n8285 & n8354 ;
  assign n8364 = ~n8353 & ~n8355 ;
  assign n8365 = ~n8363 & n8364 ;
  assign n8366 = n8362 & n8365 ;
  assign n8367 = \P1_P1_InstQueue_reg[11][7]/NET0131  & ~n8366 ;
  assign n8368 = ~n8351 & ~n8367 ;
  assign n8369 = ~n8288 & n8368 ;
  assign n8370 = ~n8284 & n8369 ;
  assign n8371 = \P1_P1_InstQueueWr_Addr_reg[2]/NET0131  & n8143 ;
  assign n8372 = \P1_P1_InstQueueWr_Addr_reg[3]/NET0131  & n8371 ;
  assign n8373 = ~n8135 & n8372 ;
  assign n8374 = \P1_P1_InstQueueWr_Addr_reg[2]/NET0131  & n4325 ;
  assign n8375 = \P1_P1_InstQueueWr_Addr_reg[3]/NET0131  & n8374 ;
  assign n8376 = ~\P1_P1_InstQueueWr_Addr_reg[3]/NET0131  & n8138 ;
  assign n8377 = \P1_P1_InstQueueWr_Addr_reg[2]/NET0131  & n8140 ;
  assign n8378 = \P1_P1_InstQueueWr_Addr_reg[3]/NET0131  & n8377 ;
  assign n8379 = ~n8376 & ~n8378 ;
  assign n8380 = n7899 & ~n8379 ;
  assign n8381 = \P1_P1_InstQueue_reg[0][7]/NET0131  & ~n8376 ;
  assign n8382 = ~n8378 & n8381 ;
  assign n8383 = ~n8380 & ~n8382 ;
  assign n8384 = ~n8372 & n8383 ;
  assign n8385 = ~n8375 & ~n8384 ;
  assign n8386 = ~n8373 & n8385 ;
  assign n8387 = ~n8275 & n8375 ;
  assign n8388 = \P1_P1_DataWidth_reg[1]/NET0131  & ~n8387 ;
  assign n8389 = ~n8386 & n8388 ;
  assign n8390 = ~\P1_P1_DataWidth_reg[1]/NET0131  & n8383 ;
  assign n8391 = n8282 & ~n8390 ;
  assign n8392 = ~n8389 & n8391 ;
  assign n8393 = n8287 & ~n8383 ;
  assign n8394 = ~n8345 & n8376 ;
  assign n8395 = ~n8381 & ~n8394 ;
  assign n8396 = n8350 & ~n8395 ;
  assign n8397 = \P1_P1_InstQueue_reg[0][7]/NET0131  & ~n8366 ;
  assign n8398 = ~n8396 & ~n8397 ;
  assign n8399 = ~n8393 & n8398 ;
  assign n8400 = ~n8392 & n8399 ;
  assign n8409 = n8135 & n8139 ;
  assign n8407 = ~\P1_P1_InstQueueWr_Addr_reg[3]/NET0131  & n8377 ;
  assign n8408 = ~n8275 & n8407 ;
  assign n8401 = ~n4327 & ~n8145 ;
  assign n8402 = n7899 & ~n8401 ;
  assign n8403 = \P1_P1_InstQueue_reg[10][7]/NET0131  & ~n8145 ;
  assign n8404 = ~n4327 & n8403 ;
  assign n8405 = ~n8402 & ~n8404 ;
  assign n8410 = ~n8139 & ~n8407 ;
  assign n8411 = ~n8405 & n8410 ;
  assign n8412 = \P1_P1_DataWidth_reg[1]/NET0131  & ~n8411 ;
  assign n8413 = ~n8408 & n8412 ;
  assign n8414 = ~n8409 & n8413 ;
  assign n8406 = ~\P1_P1_DataWidth_reg[1]/NET0131  & n8405 ;
  assign n8415 = n8282 & ~n8406 ;
  assign n8416 = ~n8414 & n8415 ;
  assign n8417 = n8287 & ~n8405 ;
  assign n8418 = n8145 & ~n8345 ;
  assign n8419 = ~n8403 & ~n8418 ;
  assign n8420 = n8350 & ~n8419 ;
  assign n8421 = \P1_P1_InstQueue_reg[10][7]/NET0131  & ~n8366 ;
  assign n8422 = ~n8420 & ~n8421 ;
  assign n8423 = ~n8417 & n8422 ;
  assign n8424 = ~n8416 & n8423 ;
  assign n8425 = ~n8135 & n8145 ;
  assign n8426 = \P1_P1_InstQueueWr_Addr_reg[2]/NET0131  & n8137 ;
  assign n8427 = \P1_P1_InstQueueWr_Addr_reg[3]/NET0131  & n8426 ;
  assign n8428 = ~n8142 & ~n8427 ;
  assign n8429 = n7899 & ~n8428 ;
  assign n8430 = \P1_P1_InstQueue_reg[12][7]/NET0131  & ~n8427 ;
  assign n8431 = ~n8142 & n8430 ;
  assign n8432 = ~n8429 & ~n8431 ;
  assign n8433 = ~n8145 & n8432 ;
  assign n8434 = ~n4327 & ~n8433 ;
  assign n8435 = ~n8425 & n8434 ;
  assign n8436 = n4327 & ~n8275 ;
  assign n8437 = \P1_P1_DataWidth_reg[1]/NET0131  & ~n8436 ;
  assign n8438 = ~n8435 & n8437 ;
  assign n8439 = ~\P1_P1_DataWidth_reg[1]/NET0131  & n8432 ;
  assign n8440 = n8282 & ~n8439 ;
  assign n8441 = ~n8438 & n8440 ;
  assign n8442 = n8287 & ~n8432 ;
  assign n8443 = ~n8345 & n8427 ;
  assign n8444 = ~n8430 & ~n8443 ;
  assign n8445 = n8350 & ~n8444 ;
  assign n8446 = \P1_P1_InstQueue_reg[12][7]/NET0131  & ~n8366 ;
  assign n8447 = ~n8445 & ~n8446 ;
  assign n8448 = ~n8442 & n8447 ;
  assign n8449 = ~n8441 & n8448 ;
  assign n8450 = ~n8135 & n8142 ;
  assign n8451 = ~n8375 & ~n8427 ;
  assign n8452 = n7899 & ~n8451 ;
  assign n8453 = \P1_P1_InstQueue_reg[13][7]/NET0131  & ~n8375 ;
  assign n8454 = ~n8427 & n8453 ;
  assign n8455 = ~n8452 & ~n8454 ;
  assign n8456 = ~n8142 & n8455 ;
  assign n8457 = ~n8145 & ~n8456 ;
  assign n8458 = ~n8450 & n8457 ;
  assign n8459 = n8145 & ~n8275 ;
  assign n8460 = \P1_P1_DataWidth_reg[1]/NET0131  & ~n8459 ;
  assign n8461 = ~n8458 & n8460 ;
  assign n8462 = ~\P1_P1_DataWidth_reg[1]/NET0131  & n8455 ;
  assign n8463 = n8282 & ~n8462 ;
  assign n8464 = ~n8461 & n8463 ;
  assign n8465 = n8287 & ~n8455 ;
  assign n8466 = ~n8345 & n8375 ;
  assign n8467 = ~n8453 & ~n8466 ;
  assign n8468 = n8350 & ~n8467 ;
  assign n8469 = \P1_P1_InstQueue_reg[13][7]/NET0131  & ~n8366 ;
  assign n8470 = ~n8468 & ~n8469 ;
  assign n8471 = ~n8465 & n8470 ;
  assign n8472 = ~n8464 & n8471 ;
  assign n8473 = ~n8135 & n8427 ;
  assign n8474 = ~n8372 & ~n8375 ;
  assign n8475 = n7899 & ~n8474 ;
  assign n8476 = \P1_P1_InstQueue_reg[14][7]/NET0131  & ~n8372 ;
  assign n8477 = ~n8375 & n8476 ;
  assign n8478 = ~n8475 & ~n8477 ;
  assign n8479 = ~n8427 & n8478 ;
  assign n8480 = ~n8142 & ~n8479 ;
  assign n8481 = ~n8473 & n8480 ;
  assign n8482 = n8142 & ~n8275 ;
  assign n8483 = \P1_P1_DataWidth_reg[1]/NET0131  & ~n8482 ;
  assign n8484 = ~n8481 & n8483 ;
  assign n8485 = ~\P1_P1_DataWidth_reg[1]/NET0131  & n8478 ;
  assign n8486 = n8282 & ~n8485 ;
  assign n8487 = ~n8484 & n8486 ;
  assign n8488 = n8287 & ~n8478 ;
  assign n8489 = ~n8345 & n8372 ;
  assign n8490 = ~n8476 & ~n8489 ;
  assign n8491 = n8350 & ~n8490 ;
  assign n8492 = \P1_P1_InstQueue_reg[14][7]/NET0131  & ~n8366 ;
  assign n8493 = ~n8491 & ~n8492 ;
  assign n8494 = ~n8488 & n8493 ;
  assign n8495 = ~n8487 & n8494 ;
  assign n8496 = ~n8135 & n8375 ;
  assign n8497 = ~n8372 & ~n8378 ;
  assign n8498 = n7899 & ~n8497 ;
  assign n8499 = \P1_P1_InstQueue_reg[15][7]/NET0131  & ~n8378 ;
  assign n8500 = ~n8372 & n8499 ;
  assign n8501 = ~n8498 & ~n8500 ;
  assign n8502 = ~n8375 & n8501 ;
  assign n8503 = ~n8427 & ~n8502 ;
  assign n8504 = ~n8496 & n8503 ;
  assign n8505 = ~n8275 & n8427 ;
  assign n8506 = \P1_P1_DataWidth_reg[1]/NET0131  & ~n8505 ;
  assign n8507 = ~n8504 & n8506 ;
  assign n8508 = ~\P1_P1_DataWidth_reg[1]/NET0131  & n8501 ;
  assign n8509 = n8282 & ~n8508 ;
  assign n8510 = ~n8507 & n8509 ;
  assign n8511 = n8287 & ~n8501 ;
  assign n8512 = ~n8345 & n8378 ;
  assign n8513 = ~n8499 & ~n8512 ;
  assign n8514 = n8350 & ~n8513 ;
  assign n8515 = \P1_P1_InstQueue_reg[15][7]/NET0131  & ~n8366 ;
  assign n8516 = ~n8514 & ~n8515 ;
  assign n8517 = ~n8511 & n8516 ;
  assign n8518 = ~n8510 & n8517 ;
  assign n8519 = ~n8135 & n8378 ;
  assign n8520 = ~\P1_P1_InstQueueWr_Addr_reg[3]/NET0131  & n4326 ;
  assign n8521 = ~n8376 & ~n8520 ;
  assign n8522 = n7899 & ~n8521 ;
  assign n8523 = \P1_P1_InstQueue_reg[1][7]/NET0131  & ~n8520 ;
  assign n8524 = ~n8376 & n8523 ;
  assign n8525 = ~n8522 & ~n8524 ;
  assign n8526 = ~n8378 & n8525 ;
  assign n8527 = ~n8372 & ~n8526 ;
  assign n8528 = ~n8519 & n8527 ;
  assign n8529 = ~n8275 & n8372 ;
  assign n8530 = \P1_P1_DataWidth_reg[1]/NET0131  & ~n8529 ;
  assign n8531 = ~n8528 & n8530 ;
  assign n8532 = ~\P1_P1_DataWidth_reg[1]/NET0131  & n8525 ;
  assign n8533 = n8282 & ~n8532 ;
  assign n8534 = ~n8531 & n8533 ;
  assign n8535 = n8287 & ~n8525 ;
  assign n8536 = ~n8345 & n8520 ;
  assign n8537 = ~n8523 & ~n8536 ;
  assign n8538 = n8350 & ~n8537 ;
  assign n8539 = \P1_P1_InstQueue_reg[1][7]/NET0131  & ~n8366 ;
  assign n8540 = ~n8538 & ~n8539 ;
  assign n8541 = ~n8535 & n8540 ;
  assign n8542 = ~n8534 & n8541 ;
  assign n8543 = ~n8135 & n8376 ;
  assign n8544 = ~\P1_P1_InstQueueWr_Addr_reg[3]/NET0131  & n8144 ;
  assign n8545 = ~n8520 & ~n8544 ;
  assign n8546 = n7899 & ~n8545 ;
  assign n8547 = \P1_P1_InstQueue_reg[2][7]/NET0131  & ~n8544 ;
  assign n8548 = ~n8520 & n8547 ;
  assign n8549 = ~n8546 & ~n8548 ;
  assign n8550 = ~n8376 & n8549 ;
  assign n8551 = ~n8378 & ~n8550 ;
  assign n8552 = ~n8543 & n8551 ;
  assign n8553 = ~n8275 & n8378 ;
  assign n8554 = \P1_P1_DataWidth_reg[1]/NET0131  & ~n8553 ;
  assign n8555 = ~n8552 & n8554 ;
  assign n8556 = ~\P1_P1_DataWidth_reg[1]/NET0131  & n8549 ;
  assign n8557 = n8282 & ~n8556 ;
  assign n8558 = ~n8555 & n8557 ;
  assign n8559 = n8287 & ~n8549 ;
  assign n8560 = ~n8345 & n8544 ;
  assign n8561 = ~n8547 & ~n8560 ;
  assign n8562 = n8350 & ~n8561 ;
  assign n8563 = \P1_P1_InstQueue_reg[2][7]/NET0131  & ~n8366 ;
  assign n8564 = ~n8562 & ~n8563 ;
  assign n8565 = ~n8559 & n8564 ;
  assign n8566 = ~n8558 & n8565 ;
  assign n8567 = ~n8135 & n8520 ;
  assign n8568 = ~\P1_P1_InstQueueWr_Addr_reg[3]/NET0131  & n8141 ;
  assign n8569 = ~n8544 & ~n8568 ;
  assign n8570 = n7899 & ~n8569 ;
  assign n8571 = \P1_P1_InstQueue_reg[3][7]/NET0131  & ~n8568 ;
  assign n8572 = ~n8544 & n8571 ;
  assign n8573 = ~n8570 & ~n8572 ;
  assign n8574 = ~n8520 & n8573 ;
  assign n8575 = ~n8376 & ~n8574 ;
  assign n8576 = ~n8567 & n8575 ;
  assign n8577 = ~n8275 & n8376 ;
  assign n8578 = \P1_P1_DataWidth_reg[1]/NET0131  & ~n8577 ;
  assign n8579 = ~n8576 & n8578 ;
  assign n8580 = ~\P1_P1_DataWidth_reg[1]/NET0131  & n8573 ;
  assign n8581 = n8282 & ~n8580 ;
  assign n8582 = ~n8579 & n8581 ;
  assign n8583 = n8287 & ~n8573 ;
  assign n8584 = ~n8345 & n8568 ;
  assign n8585 = ~n8571 & ~n8584 ;
  assign n8586 = n8350 & ~n8585 ;
  assign n8587 = \P1_P1_InstQueue_reg[3][7]/NET0131  & ~n8366 ;
  assign n8588 = ~n8586 & ~n8587 ;
  assign n8589 = ~n8583 & n8588 ;
  assign n8590 = ~n8582 & n8589 ;
  assign n8591 = ~n8135 & n8544 ;
  assign n8592 = ~\P1_P1_InstQueueWr_Addr_reg[3]/NET0131  & n8426 ;
  assign n8593 = ~n8568 & ~n8592 ;
  assign n8594 = n7899 & ~n8593 ;
  assign n8595 = \P1_P1_InstQueue_reg[4][7]/NET0131  & ~n8592 ;
  assign n8596 = ~n8568 & n8595 ;
  assign n8597 = ~n8594 & ~n8596 ;
  assign n8598 = ~n8544 & n8597 ;
  assign n8599 = ~n8520 & ~n8598 ;
  assign n8600 = ~n8591 & n8599 ;
  assign n8601 = ~n8275 & n8520 ;
  assign n8602 = \P1_P1_DataWidth_reg[1]/NET0131  & ~n8601 ;
  assign n8603 = ~n8600 & n8602 ;
  assign n8604 = ~\P1_P1_DataWidth_reg[1]/NET0131  & n8597 ;
  assign n8605 = n8282 & ~n8604 ;
  assign n8606 = ~n8603 & n8605 ;
  assign n8607 = n8287 & ~n8597 ;
  assign n8608 = ~n8345 & n8592 ;
  assign n8609 = ~n8595 & ~n8608 ;
  assign n8610 = n8350 & ~n8609 ;
  assign n8611 = \P1_P1_InstQueue_reg[4][7]/NET0131  & ~n8366 ;
  assign n8612 = ~n8610 & ~n8611 ;
  assign n8613 = ~n8607 & n8612 ;
  assign n8614 = ~n8606 & n8613 ;
  assign n8615 = ~n8135 & n8568 ;
  assign n8616 = ~\P1_P1_InstQueueWr_Addr_reg[3]/NET0131  & n8374 ;
  assign n8617 = ~n8592 & ~n8616 ;
  assign n8618 = n7899 & ~n8617 ;
  assign n8619 = \P1_P1_InstQueue_reg[5][7]/NET0131  & ~n8616 ;
  assign n8620 = ~n8592 & n8619 ;
  assign n8621 = ~n8618 & ~n8620 ;
  assign n8622 = ~n8568 & n8621 ;
  assign n8623 = ~n8544 & ~n8622 ;
  assign n8624 = ~n8615 & n8623 ;
  assign n8625 = ~n8275 & n8544 ;
  assign n8626 = \P1_P1_DataWidth_reg[1]/NET0131  & ~n8625 ;
  assign n8627 = ~n8624 & n8626 ;
  assign n8628 = ~\P1_P1_DataWidth_reg[1]/NET0131  & n8621 ;
  assign n8629 = n8282 & ~n8628 ;
  assign n8630 = ~n8627 & n8629 ;
  assign n8631 = n8287 & ~n8621 ;
  assign n8632 = ~n8345 & n8616 ;
  assign n8633 = ~n8619 & ~n8632 ;
  assign n8634 = n8350 & ~n8633 ;
  assign n8635 = \P1_P1_InstQueue_reg[5][7]/NET0131  & ~n8366 ;
  assign n8636 = ~n8634 & ~n8635 ;
  assign n8637 = ~n8631 & n8636 ;
  assign n8638 = ~n8630 & n8637 ;
  assign n8639 = ~n8135 & n8592 ;
  assign n8640 = ~\P1_P1_InstQueueWr_Addr_reg[3]/NET0131  & n8371 ;
  assign n8641 = ~n8616 & ~n8640 ;
  assign n8642 = n7899 & ~n8641 ;
  assign n8643 = \P1_P1_InstQueue_reg[6][7]/NET0131  & ~n8640 ;
  assign n8644 = ~n8616 & n8643 ;
  assign n8645 = ~n8642 & ~n8644 ;
  assign n8646 = ~n8592 & n8645 ;
  assign n8647 = ~n8568 & ~n8646 ;
  assign n8648 = ~n8639 & n8647 ;
  assign n8649 = ~n8275 & n8568 ;
  assign n8650 = \P1_P1_DataWidth_reg[1]/NET0131  & ~n8649 ;
  assign n8651 = ~n8648 & n8650 ;
  assign n8652 = ~\P1_P1_DataWidth_reg[1]/NET0131  & n8645 ;
  assign n8653 = n8282 & ~n8652 ;
  assign n8654 = ~n8651 & n8653 ;
  assign n8655 = n8287 & ~n8645 ;
  assign n8656 = ~n8345 & n8640 ;
  assign n8657 = ~n8643 & ~n8656 ;
  assign n8658 = n8350 & ~n8657 ;
  assign n8659 = \P1_P1_InstQueue_reg[6][7]/NET0131  & ~n8366 ;
  assign n8660 = ~n8658 & ~n8659 ;
  assign n8661 = ~n8655 & n8660 ;
  assign n8662 = ~n8654 & n8661 ;
  assign n8663 = ~n8135 & n8616 ;
  assign n8664 = ~n8407 & ~n8640 ;
  assign n8665 = n7899 & ~n8664 ;
  assign n8666 = \P1_P1_InstQueue_reg[7][7]/NET0131  & ~n8407 ;
  assign n8667 = ~n8640 & n8666 ;
  assign n8668 = ~n8665 & ~n8667 ;
  assign n8669 = ~n8616 & n8668 ;
  assign n8670 = ~n8592 & ~n8669 ;
  assign n8671 = ~n8663 & n8670 ;
  assign n8672 = ~n8275 & n8592 ;
  assign n8673 = \P1_P1_DataWidth_reg[1]/NET0131  & ~n8672 ;
  assign n8674 = ~n8671 & n8673 ;
  assign n8675 = ~\P1_P1_DataWidth_reg[1]/NET0131  & n8668 ;
  assign n8676 = n8282 & ~n8675 ;
  assign n8677 = ~n8674 & n8676 ;
  assign n8678 = n8287 & ~n8668 ;
  assign n8679 = ~n8345 & n8407 ;
  assign n8680 = ~n8666 & ~n8679 ;
  assign n8681 = n8350 & ~n8680 ;
  assign n8682 = \P1_P1_InstQueue_reg[7][7]/NET0131  & ~n8366 ;
  assign n8683 = ~n8681 & ~n8682 ;
  assign n8684 = ~n8678 & n8683 ;
  assign n8685 = ~n8677 & n8684 ;
  assign n8686 = ~n8135 & n8640 ;
  assign n8687 = n7899 & ~n8410 ;
  assign n8688 = \P1_P1_InstQueue_reg[8][7]/NET0131  & ~n8139 ;
  assign n8689 = ~n8407 & n8688 ;
  assign n8690 = ~n8687 & ~n8689 ;
  assign n8691 = ~n8640 & n8690 ;
  assign n8692 = ~n8616 & ~n8691 ;
  assign n8693 = ~n8686 & n8692 ;
  assign n8694 = ~n8275 & n8616 ;
  assign n8695 = \P1_P1_DataWidth_reg[1]/NET0131  & ~n8694 ;
  assign n8696 = ~n8693 & n8695 ;
  assign n8697 = ~\P1_P1_DataWidth_reg[1]/NET0131  & n8690 ;
  assign n8698 = n8282 & ~n8697 ;
  assign n8699 = ~n8696 & n8698 ;
  assign n8700 = n8287 & ~n8690 ;
  assign n8701 = n8139 & ~n8345 ;
  assign n8702 = ~n8688 & ~n8701 ;
  assign n8703 = n8350 & ~n8702 ;
  assign n8704 = \P1_P1_InstQueue_reg[8][7]/NET0131  & ~n8366 ;
  assign n8705 = ~n8703 & ~n8704 ;
  assign n8706 = ~n8700 & n8705 ;
  assign n8707 = ~n8699 & n8706 ;
  assign n8708 = ~n8135 & n8407 ;
  assign n8709 = ~n4327 & ~n8139 ;
  assign n8710 = n7899 & ~n8709 ;
  assign n8711 = \P1_P1_InstQueue_reg[9][7]/NET0131  & ~n4327 ;
  assign n8712 = ~n8139 & n8711 ;
  assign n8713 = ~n8710 & ~n8712 ;
  assign n8714 = ~n8407 & n8713 ;
  assign n8715 = ~n8640 & ~n8714 ;
  assign n8716 = ~n8708 & n8715 ;
  assign n8717 = ~n8275 & n8640 ;
  assign n8718 = \P1_P1_DataWidth_reg[1]/NET0131  & ~n8717 ;
  assign n8719 = ~n8716 & n8718 ;
  assign n8720 = ~\P1_P1_DataWidth_reg[1]/NET0131  & n8713 ;
  assign n8721 = n8282 & ~n8720 ;
  assign n8722 = ~n8719 & n8721 ;
  assign n8723 = n8287 & ~n8713 ;
  assign n8724 = n4327 & ~n8345 ;
  assign n8725 = ~n8711 & ~n8724 ;
  assign n8726 = n8350 & ~n8725 ;
  assign n8727 = \P1_P1_InstQueue_reg[9][7]/NET0131  & ~n8366 ;
  assign n8728 = ~n8726 & ~n8727 ;
  assign n8729 = ~n8723 & n8728 ;
  assign n8730 = ~n8722 & n8729 ;
  assign n8756 = ~\P1_P3_InstQueueRd_Addr_reg[2]/NET0131  & \P1_P3_InstQueueRd_Addr_reg[3]/NET0131  ;
  assign n8762 = \P1_P3_InstQueueRd_Addr_reg[0]/NET0131  & ~\P1_P3_InstQueueRd_Addr_reg[1]/NET0131  ;
  assign n8763 = n8756 & n8762 ;
  assign n8834 = \P1_P3_InstQueue_reg[9][5]/NET0131  & n8763 ;
  assign n8759 = \P1_P3_InstQueueRd_Addr_reg[2]/NET0131  & \P1_P3_InstQueueRd_Addr_reg[3]/NET0131  ;
  assign n8775 = n8759 & n8762 ;
  assign n8835 = \P1_P3_InstQueue_reg[13][5]/NET0131  & n8775 ;
  assign n8848 = ~n8834 & ~n8835 ;
  assign n8744 = ~\P1_P3_InstQueueRd_Addr_reg[0]/NET0131  & ~\P1_P3_InstQueueRd_Addr_reg[1]/NET0131  ;
  assign n8769 = n8744 & n8756 ;
  assign n8836 = \P1_P3_InstQueue_reg[8][5]/NET0131  & n8769 ;
  assign n8747 = \P1_P3_InstQueueRd_Addr_reg[0]/NET0131  & \P1_P3_InstQueueRd_Addr_reg[1]/NET0131  ;
  assign n8765 = n8747 & n8756 ;
  assign n8837 = \P1_P3_InstQueue_reg[11][5]/NET0131  & n8765 ;
  assign n8849 = ~n8836 & ~n8837 ;
  assign n8856 = n8848 & n8849 ;
  assign n8760 = n8744 & n8759 ;
  assign n8830 = \P1_P3_InstQueue_reg[12][5]/NET0131  & n8760 ;
  assign n8743 = \P1_P3_InstQueueRd_Addr_reg[2]/NET0131  & ~\P1_P3_InstQueueRd_Addr_reg[3]/NET0131  ;
  assign n8748 = n8743 & n8747 ;
  assign n8831 = \P1_P3_InstQueue_reg[7][5]/NET0131  & n8748 ;
  assign n8846 = ~n8830 & ~n8831 ;
  assign n8751 = ~\P1_P3_InstQueueRd_Addr_reg[0]/NET0131  & \P1_P3_InstQueueRd_Addr_reg[1]/NET0131  ;
  assign n8757 = n8751 & n8756 ;
  assign n8832 = \P1_P3_InstQueue_reg[10][5]/NET0131  & n8757 ;
  assign n8750 = ~\P1_P3_InstQueueRd_Addr_reg[2]/NET0131  & ~\P1_P3_InstQueueRd_Addr_reg[3]/NET0131  ;
  assign n8777 = n8750 & n8762 ;
  assign n8833 = \P1_P3_InstQueue_reg[1][5]/NET0131  & n8777 ;
  assign n8847 = ~n8832 & ~n8833 ;
  assign n8857 = n8846 & n8847 ;
  assign n8858 = n8856 & n8857 ;
  assign n8767 = n8744 & n8750 ;
  assign n8842 = \P1_P3_InstQueue_reg[0][5]/NET0131  & n8767 ;
  assign n8745 = n8743 & n8744 ;
  assign n8843 = \P1_P3_InstQueue_reg[4][5]/NET0131  & n8745 ;
  assign n8852 = ~n8842 & ~n8843 ;
  assign n8752 = n8750 & n8751 ;
  assign n8844 = \P1_P3_InstQueue_reg[2][5]/NET0131  & n8752 ;
  assign n8781 = n8751 & n8759 ;
  assign n8845 = \P1_P3_InstQueue_reg[14][5]/NET0131  & n8781 ;
  assign n8853 = ~n8844 & ~n8845 ;
  assign n8854 = n8852 & n8853 ;
  assign n8754 = n8743 & n8751 ;
  assign n8838 = \P1_P3_InstQueue_reg[6][5]/NET0131  & n8754 ;
  assign n8771 = n8747 & n8750 ;
  assign n8839 = \P1_P3_InstQueue_reg[3][5]/NET0131  & n8771 ;
  assign n8850 = ~n8838 & ~n8839 ;
  assign n8779 = n8743 & n8762 ;
  assign n8840 = \P1_P3_InstQueue_reg[5][5]/NET0131  & n8779 ;
  assign n8773 = n8747 & n8759 ;
  assign n8841 = \P1_P3_InstQueue_reg[15][5]/NET0131  & n8773 ;
  assign n8851 = ~n8840 & ~n8841 ;
  assign n8855 = n8850 & n8851 ;
  assign n8859 = n8854 & n8855 ;
  assign n8860 = n8858 & n8859 ;
  assign n8865 = \P1_P3_InstQueue_reg[13][4]/NET0131  & n8775 ;
  assign n8866 = \P1_P3_InstQueue_reg[1][4]/NET0131  & n8777 ;
  assign n8879 = ~n8865 & ~n8866 ;
  assign n8867 = \P1_P3_InstQueue_reg[5][4]/NET0131  & n8779 ;
  assign n8868 = \P1_P3_InstQueue_reg[6][4]/NET0131  & n8754 ;
  assign n8880 = ~n8867 & ~n8868 ;
  assign n8887 = n8879 & n8880 ;
  assign n8861 = \P1_P3_InstQueue_reg[4][4]/NET0131  & n8745 ;
  assign n8862 = \P1_P3_InstQueue_reg[7][4]/NET0131  & n8748 ;
  assign n8877 = ~n8861 & ~n8862 ;
  assign n8863 = \P1_P3_InstQueue_reg[10][4]/NET0131  & n8757 ;
  assign n8864 = \P1_P3_InstQueue_reg[3][4]/NET0131  & n8771 ;
  assign n8878 = ~n8863 & ~n8864 ;
  assign n8888 = n8877 & n8878 ;
  assign n8889 = n8887 & n8888 ;
  assign n8873 = \P1_P3_InstQueue_reg[0][4]/NET0131  & n8767 ;
  assign n8874 = \P1_P3_InstQueue_reg[9][4]/NET0131  & n8763 ;
  assign n8883 = ~n8873 & ~n8874 ;
  assign n8875 = \P1_P3_InstQueue_reg[2][4]/NET0131  & n8752 ;
  assign n8876 = \P1_P3_InstQueue_reg[14][4]/NET0131  & n8781 ;
  assign n8884 = ~n8875 & ~n8876 ;
  assign n8885 = n8883 & n8884 ;
  assign n8869 = \P1_P3_InstQueue_reg[12][4]/NET0131  & n8760 ;
  assign n8870 = \P1_P3_InstQueue_reg[11][4]/NET0131  & n8765 ;
  assign n8881 = ~n8869 & ~n8870 ;
  assign n8871 = \P1_P3_InstQueue_reg[8][4]/NET0131  & n8769 ;
  assign n8872 = \P1_P3_InstQueue_reg[15][4]/NET0131  & n8773 ;
  assign n8882 = ~n8871 & ~n8872 ;
  assign n8886 = n8881 & n8882 ;
  assign n8890 = n8885 & n8886 ;
  assign n8891 = n8889 & n8890 ;
  assign n8758 = \P1_P3_InstQueue_reg[10][7]/NET0131  & n8757 ;
  assign n8761 = \P1_P3_InstQueue_reg[12][7]/NET0131  & n8760 ;
  assign n8785 = ~n8758 & ~n8761 ;
  assign n8764 = \P1_P3_InstQueue_reg[9][7]/NET0131  & n8763 ;
  assign n8766 = \P1_P3_InstQueue_reg[11][7]/NET0131  & n8765 ;
  assign n8786 = ~n8764 & ~n8766 ;
  assign n8793 = n8785 & n8786 ;
  assign n8746 = \P1_P3_InstQueue_reg[4][7]/NET0131  & n8745 ;
  assign n8749 = \P1_P3_InstQueue_reg[7][7]/NET0131  & n8748 ;
  assign n8783 = ~n8746 & ~n8749 ;
  assign n8753 = \P1_P3_InstQueue_reg[2][7]/NET0131  & n8752 ;
  assign n8755 = \P1_P3_InstQueue_reg[6][7]/NET0131  & n8754 ;
  assign n8784 = ~n8753 & ~n8755 ;
  assign n8794 = n8783 & n8784 ;
  assign n8795 = n8793 & n8794 ;
  assign n8776 = \P1_P3_InstQueue_reg[13][7]/NET0131  & n8775 ;
  assign n8778 = \P1_P3_InstQueue_reg[1][7]/NET0131  & n8777 ;
  assign n8789 = ~n8776 & ~n8778 ;
  assign n8780 = \P1_P3_InstQueue_reg[5][7]/NET0131  & n8779 ;
  assign n8782 = \P1_P3_InstQueue_reg[14][7]/NET0131  & n8781 ;
  assign n8790 = ~n8780 & ~n8782 ;
  assign n8791 = n8789 & n8790 ;
  assign n8768 = \P1_P3_InstQueue_reg[0][7]/NET0131  & n8767 ;
  assign n8770 = \P1_P3_InstQueue_reg[8][7]/NET0131  & n8769 ;
  assign n8787 = ~n8768 & ~n8770 ;
  assign n8772 = \P1_P3_InstQueue_reg[3][7]/NET0131  & n8771 ;
  assign n8774 = \P1_P3_InstQueue_reg[15][7]/NET0131  & n8773 ;
  assign n8788 = ~n8772 & ~n8774 ;
  assign n8792 = n8787 & n8788 ;
  assign n8796 = n8791 & n8792 ;
  assign n8797 = n8795 & n8796 ;
  assign n8802 = \P1_P3_InstQueue_reg[13][6]/NET0131  & n8775 ;
  assign n8803 = \P1_P3_InstQueue_reg[1][6]/NET0131  & n8777 ;
  assign n8816 = ~n8802 & ~n8803 ;
  assign n8804 = \P1_P3_InstQueue_reg[5][6]/NET0131  & n8779 ;
  assign n8805 = \P1_P3_InstQueue_reg[6][6]/NET0131  & n8754 ;
  assign n8817 = ~n8804 & ~n8805 ;
  assign n8824 = n8816 & n8817 ;
  assign n8798 = \P1_P3_InstQueue_reg[4][6]/NET0131  & n8745 ;
  assign n8799 = \P1_P3_InstQueue_reg[7][6]/NET0131  & n8748 ;
  assign n8814 = ~n8798 & ~n8799 ;
  assign n8800 = \P1_P3_InstQueue_reg[10][6]/NET0131  & n8757 ;
  assign n8801 = \P1_P3_InstQueue_reg[3][6]/NET0131  & n8771 ;
  assign n8815 = ~n8800 & ~n8801 ;
  assign n8825 = n8814 & n8815 ;
  assign n8826 = n8824 & n8825 ;
  assign n8810 = \P1_P3_InstQueue_reg[0][6]/NET0131  & n8767 ;
  assign n8811 = \P1_P3_InstQueue_reg[9][6]/NET0131  & n8763 ;
  assign n8820 = ~n8810 & ~n8811 ;
  assign n8812 = \P1_P3_InstQueue_reg[2][6]/NET0131  & n8752 ;
  assign n8813 = \P1_P3_InstQueue_reg[14][6]/NET0131  & n8781 ;
  assign n8821 = ~n8812 & ~n8813 ;
  assign n8822 = n8820 & n8821 ;
  assign n8806 = \P1_P3_InstQueue_reg[12][6]/NET0131  & n8760 ;
  assign n8807 = \P1_P3_InstQueue_reg[11][6]/NET0131  & n8765 ;
  assign n8818 = ~n8806 & ~n8807 ;
  assign n8808 = \P1_P3_InstQueue_reg[8][6]/NET0131  & n8769 ;
  assign n8809 = \P1_P3_InstQueue_reg[15][6]/NET0131  & n8773 ;
  assign n8819 = ~n8808 & ~n8809 ;
  assign n8823 = n8818 & n8819 ;
  assign n8827 = n8822 & n8823 ;
  assign n8828 = n8826 & n8827 ;
  assign n9051 = ~n8797 & n8828 ;
  assign n9052 = ~n8891 & n9051 ;
  assign n9053 = ~n8860 & n9052 ;
  assign n8929 = \P1_P3_InstQueue_reg[9][3]/NET0131  & n8763 ;
  assign n8930 = \P1_P3_InstQueue_reg[1][3]/NET0131  & n8777 ;
  assign n8943 = ~n8929 & ~n8930 ;
  assign n8931 = \P1_P3_InstQueue_reg[8][3]/NET0131  & n8769 ;
  assign n8932 = \P1_P3_InstQueue_reg[11][3]/NET0131  & n8765 ;
  assign n8944 = ~n8931 & ~n8932 ;
  assign n8951 = n8943 & n8944 ;
  assign n8925 = \P1_P3_InstQueue_reg[12][3]/NET0131  & n8760 ;
  assign n8926 = \P1_P3_InstQueue_reg[7][3]/NET0131  & n8748 ;
  assign n8941 = ~n8925 & ~n8926 ;
  assign n8927 = \P1_P3_InstQueue_reg[10][3]/NET0131  & n8757 ;
  assign n8928 = \P1_P3_InstQueue_reg[6][3]/NET0131  & n8754 ;
  assign n8942 = ~n8927 & ~n8928 ;
  assign n8952 = n8941 & n8942 ;
  assign n8953 = n8951 & n8952 ;
  assign n8937 = \P1_P3_InstQueue_reg[4][3]/NET0131  & n8745 ;
  assign n8938 = \P1_P3_InstQueue_reg[0][3]/NET0131  & n8767 ;
  assign n8947 = ~n8937 & ~n8938 ;
  assign n8939 = \P1_P3_InstQueue_reg[2][3]/NET0131  & n8752 ;
  assign n8940 = \P1_P3_InstQueue_reg[14][3]/NET0131  & n8781 ;
  assign n8948 = ~n8939 & ~n8940 ;
  assign n8949 = n8947 & n8948 ;
  assign n8933 = \P1_P3_InstQueue_reg[13][3]/NET0131  & n8775 ;
  assign n8934 = \P1_P3_InstQueue_reg[3][3]/NET0131  & n8771 ;
  assign n8945 = ~n8933 & ~n8934 ;
  assign n8935 = \P1_P3_InstQueue_reg[5][3]/NET0131  & n8779 ;
  assign n8936 = \P1_P3_InstQueue_reg[15][3]/NET0131  & n8773 ;
  assign n8946 = ~n8935 & ~n8936 ;
  assign n8950 = n8945 & n8946 ;
  assign n8954 = n8949 & n8950 ;
  assign n8955 = n8953 & n8954 ;
  assign n8898 = \P1_P3_InstQueue_reg[10][0]/NET0131  & n8757 ;
  assign n8899 = \P1_P3_InstQueue_reg[12][0]/NET0131  & n8760 ;
  assign n8912 = ~n8898 & ~n8899 ;
  assign n8900 = \P1_P3_InstQueue_reg[9][0]/NET0131  & n8763 ;
  assign n8901 = \P1_P3_InstQueue_reg[11][0]/NET0131  & n8765 ;
  assign n8913 = ~n8900 & ~n8901 ;
  assign n8920 = n8912 & n8913 ;
  assign n8894 = \P1_P3_InstQueue_reg[4][0]/NET0131  & n8745 ;
  assign n8895 = \P1_P3_InstQueue_reg[7][0]/NET0131  & n8748 ;
  assign n8910 = ~n8894 & ~n8895 ;
  assign n8896 = \P1_P3_InstQueue_reg[8][0]/NET0131  & n8769 ;
  assign n8897 = \P1_P3_InstQueue_reg[6][0]/NET0131  & n8754 ;
  assign n8911 = ~n8896 & ~n8897 ;
  assign n8921 = n8910 & n8911 ;
  assign n8922 = n8920 & n8921 ;
  assign n8906 = \P1_P3_InstQueue_reg[13][0]/NET0131  & n8775 ;
  assign n8907 = \P1_P3_InstQueue_reg[1][0]/NET0131  & n8777 ;
  assign n8916 = ~n8906 & ~n8907 ;
  assign n8908 = \P1_P3_InstQueue_reg[2][0]/NET0131  & n8752 ;
  assign n8909 = \P1_P3_InstQueue_reg[14][0]/NET0131  & n8781 ;
  assign n8917 = ~n8908 & ~n8909 ;
  assign n8918 = n8916 & n8917 ;
  assign n8902 = \P1_P3_InstQueue_reg[0][0]/NET0131  & n8767 ;
  assign n8903 = \P1_P3_InstQueue_reg[5][0]/NET0131  & n8779 ;
  assign n8914 = ~n8902 & ~n8903 ;
  assign n8904 = \P1_P3_InstQueue_reg[3][0]/NET0131  & n8771 ;
  assign n8905 = \P1_P3_InstQueue_reg[15][0]/NET0131  & n8773 ;
  assign n8915 = ~n8904 & ~n8905 ;
  assign n8919 = n8914 & n8915 ;
  assign n8923 = n8918 & n8919 ;
  assign n8924 = n8922 & n8923 ;
  assign n8961 = \P1_P3_InstQueue_reg[9][2]/NET0131  & n8763 ;
  assign n8962 = \P1_P3_InstQueue_reg[13][2]/NET0131  & n8775 ;
  assign n8975 = ~n8961 & ~n8962 ;
  assign n8963 = \P1_P3_InstQueue_reg[8][2]/NET0131  & n8769 ;
  assign n8964 = \P1_P3_InstQueue_reg[11][2]/NET0131  & n8765 ;
  assign n8976 = ~n8963 & ~n8964 ;
  assign n8983 = n8975 & n8976 ;
  assign n8957 = \P1_P3_InstQueue_reg[12][2]/NET0131  & n8760 ;
  assign n8958 = \P1_P3_InstQueue_reg[7][2]/NET0131  & n8748 ;
  assign n8973 = ~n8957 & ~n8958 ;
  assign n8959 = \P1_P3_InstQueue_reg[10][2]/NET0131  & n8757 ;
  assign n8960 = \P1_P3_InstQueue_reg[1][2]/NET0131  & n8777 ;
  assign n8974 = ~n8959 & ~n8960 ;
  assign n8984 = n8973 & n8974 ;
  assign n8985 = n8983 & n8984 ;
  assign n8969 = \P1_P3_InstQueue_reg[0][2]/NET0131  & n8767 ;
  assign n8970 = \P1_P3_InstQueue_reg[4][2]/NET0131  & n8745 ;
  assign n8979 = ~n8969 & ~n8970 ;
  assign n8971 = \P1_P3_InstQueue_reg[2][2]/NET0131  & n8752 ;
  assign n8972 = \P1_P3_InstQueue_reg[14][2]/NET0131  & n8781 ;
  assign n8980 = ~n8971 & ~n8972 ;
  assign n8981 = n8979 & n8980 ;
  assign n8965 = \P1_P3_InstQueue_reg[6][2]/NET0131  & n8754 ;
  assign n8966 = \P1_P3_InstQueue_reg[3][2]/NET0131  & n8771 ;
  assign n8977 = ~n8965 & ~n8966 ;
  assign n8967 = \P1_P3_InstQueue_reg[5][2]/NET0131  & n8779 ;
  assign n8968 = \P1_P3_InstQueue_reg[15][2]/NET0131  & n8773 ;
  assign n8978 = ~n8967 & ~n8968 ;
  assign n8982 = n8977 & n8978 ;
  assign n8986 = n8981 & n8982 ;
  assign n8987 = n8985 & n8986 ;
  assign n8992 = \P1_P3_InstQueue_reg[13][1]/NET0131  & n8775 ;
  assign n8993 = \P1_P3_InstQueue_reg[1][1]/NET0131  & n8777 ;
  assign n9006 = ~n8992 & ~n8993 ;
  assign n8994 = \P1_P3_InstQueue_reg[8][1]/NET0131  & n8769 ;
  assign n8995 = \P1_P3_InstQueue_reg[6][1]/NET0131  & n8754 ;
  assign n9007 = ~n8994 & ~n8995 ;
  assign n9014 = n9006 & n9007 ;
  assign n8988 = \P1_P3_InstQueue_reg[4][1]/NET0131  & n8745 ;
  assign n8989 = \P1_P3_InstQueue_reg[7][1]/NET0131  & n8748 ;
  assign n9004 = ~n8988 & ~n8989 ;
  assign n8990 = \P1_P3_InstQueue_reg[10][1]/NET0131  & n8757 ;
  assign n8991 = \P1_P3_InstQueue_reg[3][1]/NET0131  & n8771 ;
  assign n9005 = ~n8990 & ~n8991 ;
  assign n9015 = n9004 & n9005 ;
  assign n9016 = n9014 & n9015 ;
  assign n9000 = \P1_P3_InstQueue_reg[0][1]/NET0131  & n8767 ;
  assign n9001 = \P1_P3_InstQueue_reg[9][1]/NET0131  & n8763 ;
  assign n9010 = ~n9000 & ~n9001 ;
  assign n9002 = \P1_P3_InstQueue_reg[2][1]/NET0131  & n8752 ;
  assign n9003 = \P1_P3_InstQueue_reg[14][1]/NET0131  & n8781 ;
  assign n9011 = ~n9002 & ~n9003 ;
  assign n9012 = n9010 & n9011 ;
  assign n8996 = \P1_P3_InstQueue_reg[12][1]/NET0131  & n8760 ;
  assign n8997 = \P1_P3_InstQueue_reg[11][1]/NET0131  & n8765 ;
  assign n9008 = ~n8996 & ~n8997 ;
  assign n8998 = \P1_P3_InstQueue_reg[5][1]/NET0131  & n8779 ;
  assign n8999 = \P1_P3_InstQueue_reg[15][1]/NET0131  & n8773 ;
  assign n9009 = ~n8998 & ~n8999 ;
  assign n9013 = n9008 & n9009 ;
  assign n9017 = n9012 & n9013 ;
  assign n9018 = n9016 & n9017 ;
  assign n9054 = n8987 & ~n9018 ;
  assign n9055 = ~n8924 & n9054 ;
  assign n9056 = ~n8955 & n9055 ;
  assign n9057 = n9053 & n9056 ;
  assign n9019 = n8987 & n9018 ;
  assign n9058 = n8924 & ~n8955 ;
  assign n9059 = n9019 & n9058 ;
  assign n9060 = n9053 & n9059 ;
  assign n9061 = ~n9057 & ~n9060 ;
  assign n8829 = ~n8797 & ~n8828 ;
  assign n8892 = ~n8860 & n8891 ;
  assign n8893 = n8829 & n8892 ;
  assign n8956 = ~n8924 & ~n8955 ;
  assign n9020 = n8956 & n9019 ;
  assign n9021 = n8893 & n9020 ;
  assign n9063 = n8893 & n9054 ;
  assign n9064 = n8956 & n9063 ;
  assign n9114 = ~n9021 & ~n9064 ;
  assign n9077 = n8860 & n8891 ;
  assign n9078 = n9051 & n9077 ;
  assign n9079 = n9020 & n9078 ;
  assign n9080 = n8955 & ~n8987 ;
  assign n9081 = n8924 & n9080 ;
  assign n9082 = n8893 & n9081 ;
  assign n9085 = n9056 & n9078 ;
  assign n9115 = ~n9082 & ~n9085 ;
  assign n9116 = ~n9079 & n9115 ;
  assign n9110 = n8924 & n8955 ;
  assign n9111 = n9019 & n9110 ;
  assign n9117 = n8829 & n8860 ;
  assign n9118 = n9111 & n9117 ;
  assign n9119 = n9116 & ~n9118 ;
  assign n9120 = n9114 & n9119 ;
  assign n9121 = n9061 & n9120 ;
  assign n9105 = n8797 & ~n8828 ;
  assign n9106 = n9077 & n9105 ;
  assign n9107 = n8955 & n9055 ;
  assign n9108 = n9106 & n9107 ;
  assign n9125 = n8797 & n8828 ;
  assign n9126 = n9018 & n9125 ;
  assign n9127 = n9077 & n9080 ;
  assign n9128 = n9126 & n9127 ;
  assign n9129 = ~n9108 & ~n9128 ;
  assign n9122 = n8892 & ~n9018 ;
  assign n9123 = n9105 & n9122 ;
  assign n9124 = n9081 & n9123 ;
  assign n9109 = ~n9052 & ~n9106 ;
  assign n9112 = ~n9109 & n9111 ;
  assign n9113 = n9058 & n9063 ;
  assign n9130 = ~n9112 & ~n9113 ;
  assign n9131 = ~n9124 & n9130 ;
  assign n9132 = n9129 & n9131 ;
  assign n9133 = ~n9121 & n9132 ;
  assign n9022 = ~\P1_P3_InstQueueRd_Addr_reg[3]/NET0131  & \P1_P3_InstQueueWr_Addr_reg[3]/NET0131  ;
  assign n9023 = \P1_P3_InstQueueRd_Addr_reg[3]/NET0131  & ~\P1_P3_InstQueueWr_Addr_reg[3]/NET0131  ;
  assign n9024 = ~n9022 & ~n9023 ;
  assign n9025 = ~\P1_P3_InstQueueRd_Addr_reg[2]/NET0131  & \P1_P3_InstQueueWr_Addr_reg[2]/NET0131  ;
  assign n9026 = \P1_P3_InstQueueRd_Addr_reg[2]/NET0131  & ~\P1_P3_InstQueueWr_Addr_reg[2]/NET0131  ;
  assign n9027 = ~\P1_P3_InstQueueRd_Addr_reg[1]/NET0131  & \P1_P3_InstQueueWr_Addr_reg[1]/NET0131  ;
  assign n9028 = \P1_P3_InstQueueRd_Addr_reg[1]/NET0131  & ~\P1_P3_InstQueueWr_Addr_reg[1]/NET0131  ;
  assign n9029 = \P1_P3_InstQueueRd_Addr_reg[0]/NET0131  & ~\P1_P3_InstQueueWr_Addr_reg[0]/NET0131  ;
  assign n9030 = ~n9028 & ~n9029 ;
  assign n9031 = ~n9027 & ~n9030 ;
  assign n9032 = ~n9026 & ~n9031 ;
  assign n9033 = ~n9025 & ~n9032 ;
  assign n9034 = n9024 & n9033 ;
  assign n9035 = ~n9024 & ~n9033 ;
  assign n9036 = ~n9034 & ~n9035 ;
  assign n9037 = ~n9025 & ~n9026 ;
  assign n9038 = n9031 & ~n9037 ;
  assign n9039 = ~n9031 & n9037 ;
  assign n9040 = ~n9038 & ~n9039 ;
  assign n9041 = ~n9027 & ~n9028 ;
  assign n9042 = ~\P1_P3_InstQueueRd_Addr_reg[0]/NET0131  & \P1_P3_InstQueueWr_Addr_reg[0]/NET0131  ;
  assign n9043 = ~n9029 & ~n9042 ;
  assign n9044 = n9041 & n9043 ;
  assign n9045 = n9040 & ~n9044 ;
  assign n9046 = n9036 & ~n9045 ;
  assign n9047 = ~n9023 & ~n9033 ;
  assign n9048 = ~n9022 & ~n9047 ;
  assign n9049 = ~n9046 & ~n9048 ;
  assign n9220 = n9049 & ~n9061 ;
  assign n9221 = n9133 & ~n9220 ;
  assign n9222 = ~\P1_P3_InstQueueRd_Addr_reg[0]/NET0131  & n9221 ;
  assign n9062 = ~n9049 & ~n9061 ;
  assign n9223 = \P1_P3_InstQueueRd_Addr_reg[0]/NET0131  & ~n9062 ;
  assign n9224 = n9120 & n9223 ;
  assign n9225 = ~n9222 & ~n9224 ;
  assign n9207 = ~n8751 & ~n8762 ;
  assign n9208 = ~n9133 & ~n9207 ;
  assign n9065 = n9036 & ~n9040 ;
  assign n9066 = ~n9048 & ~n9065 ;
  assign n9067 = n9029 & ~n9041 ;
  assign n9068 = ~n9029 & n9041 ;
  assign n9069 = ~n9067 & ~n9068 ;
  assign n9070 = ~n9048 & n9069 ;
  assign n9075 = ~n9066 & ~n9070 ;
  assign n9086 = n9018 & n9082 ;
  assign n9087 = ~n9085 & ~n9086 ;
  assign n9135 = n9075 & ~n9087 ;
  assign n9136 = n9114 & ~n9135 ;
  assign n9083 = ~n9018 & n9082 ;
  assign n9084 = ~n9079 & ~n9083 ;
  assign n9091 = ~\P1_P3_State_reg[0]/NET0131  & \P1_P3_State_reg[1]/NET0131  ;
  assign n9092 = ~\P1_P3_State_reg[2]/NET0131  & n9091 ;
  assign n9093 = ~\P1_P3_State_reg[0]/NET0131  & ~\P1_P3_State_reg[1]/NET0131  ;
  assign n9094 = \P1_P3_State_reg[2]/NET0131  & n9093 ;
  assign n9095 = ~n9092 & ~n9094 ;
  assign n9162 = ~n9075 & ~n9095 ;
  assign n9163 = ~n9084 & ~n9162 ;
  assign n9164 = n9136 & ~n9163 ;
  assign n9209 = \P1_P3_InstQueueRd_Addr_reg[1]/NET0131  & ~n9164 ;
  assign n9147 = ~n9075 & ~n9087 ;
  assign n9165 = ~n9084 & n9162 ;
  assign n9166 = ~n9147 & ~n9165 ;
  assign n8737 = ~\P1_P3_ADS_n_reg/NET0131  & \P1_P3_D_C_n_reg/NET0131  ;
  assign n8738 = \P1_P3_M_IO_n_reg/NET0131  & \P1_P3_W_R_n_reg/NET0131  ;
  assign n8739 = \P3_rd_reg/NET0131  & n8738 ;
  assign n8740 = n8737 & n8739 ;
  assign n8741 = \P1_ready22_reg/NET0131  & ~n8740 ;
  assign n9148 = \P1_P3_InstQueueRd_Addr_reg[1]/NET0131  & ~n8741 ;
  assign n9204 = ~\P1_P3_InstQueueRd_Addr_reg[1]/NET0131  & n8741 ;
  assign n9205 = ~n9148 & ~n9204 ;
  assign n9206 = ~n9166 & n9205 ;
  assign n9210 = ~\P1_P3_InstQueueRd_Addr_reg[1]/NET0131  & n9118 ;
  assign n9211 = ~\P1_P3_InstQueueRd_Addr_reg[1]/NET0131  & ~n9049 ;
  assign n9212 = n9049 & n9207 ;
  assign n9213 = ~n9211 & ~n9212 ;
  assign n9214 = ~n9061 & n9213 ;
  assign n9215 = ~n9210 & ~n9214 ;
  assign n9216 = ~n9206 & n9215 ;
  assign n9217 = ~n9209 & n9216 ;
  assign n9218 = ~n9208 & n9217 ;
  assign n9219 = ~\P1_P3_InstQueueWr_Addr_reg[1]/NET0131  & ~n9218 ;
  assign n9226 = \P1_P3_InstQueueWr_Addr_reg[0]/NET0131  & ~n9219 ;
  assign n9227 = ~n9225 & n9226 ;
  assign n9103 = \P1_P3_InstQueueRd_Addr_reg[2]/NET0131  & n8747 ;
  assign n9179 = \P1_P3_InstQueueRd_Addr_reg[3]/NET0131  & ~n9103 ;
  assign n9180 = ~n8748 & ~n9179 ;
  assign n9181 = ~n9133 & ~n9180 ;
  assign n9144 = \P1_P3_InstQueueRd_Addr_reg[1]/NET0131  & \P1_P3_InstQueueRd_Addr_reg[2]/NET0131  ;
  assign n9168 = ~n9118 & n9166 ;
  assign n9169 = ~n9144 & ~n9168 ;
  assign n9167 = n8741 & ~n9166 ;
  assign n9170 = n9164 & ~n9167 ;
  assign n9171 = ~n9169 & n9170 ;
  assign n9172 = \P1_P3_InstQueueRd_Addr_reg[3]/NET0131  & ~n9171 ;
  assign n9096 = ~n8741 & ~n9095 ;
  assign n9097 = ~n9075 & n9096 ;
  assign n9173 = ~n9084 & n9097 ;
  assign n9174 = ~n9118 & ~n9173 ;
  assign n9088 = ~n8741 & ~n9075 ;
  assign n9175 = ~n9087 & n9088 ;
  assign n9176 = n9174 & ~n9175 ;
  assign n9177 = \P1_P3_InstQueueRd_Addr_reg[1]/NET0131  & n8743 ;
  assign n9178 = ~n9176 & n9177 ;
  assign n9102 = ~\P1_P3_InstQueueRd_Addr_reg[2]/NET0131  & ~n8747 ;
  assign n9182 = n9049 & ~n9102 ;
  assign n9183 = \P1_P3_InstQueueRd_Addr_reg[3]/NET0131  & n9182 ;
  assign n9184 = ~\P1_P3_InstQueueRd_Addr_reg[3]/NET0131  & ~n9182 ;
  assign n9185 = ~n9183 & ~n9184 ;
  assign n9186 = ~n9061 & n9185 ;
  assign n9187 = ~n9178 & ~n9186 ;
  assign n9188 = ~n9172 & n9187 ;
  assign n9189 = ~n9181 & n9188 ;
  assign n9200 = \P1_P3_InstQueueWr_Addr_reg[3]/NET0131  & n9189 ;
  assign n9104 = ~n9102 & ~n9103 ;
  assign n9134 = n9104 & ~n9133 ;
  assign n9137 = ~n9084 & ~n9097 ;
  assign n9138 = n9136 & ~n9137 ;
  assign n9139 = \P1_P3_InstQueueRd_Addr_reg[2]/NET0131  & ~n9138 ;
  assign n9141 = ~\P1_P3_InstQueueRd_Addr_reg[2]/NET0131  & ~n9097 ;
  assign n9142 = ~n9084 & ~n9141 ;
  assign n9143 = ~n9118 & ~n9142 ;
  assign n9140 = ~\P1_P3_InstQueueRd_Addr_reg[1]/NET0131  & ~\P1_P3_InstQueueRd_Addr_reg[2]/NET0131  ;
  assign n9145 = ~n9140 & ~n9144 ;
  assign n9146 = ~n9143 & n9145 ;
  assign n9149 = ~\P1_P3_InstQueueRd_Addr_reg[2]/NET0131  & ~n9148 ;
  assign n9150 = \P1_P3_InstQueueRd_Addr_reg[2]/NET0131  & n9148 ;
  assign n9151 = ~n9149 & ~n9150 ;
  assign n9152 = n9147 & n9151 ;
  assign n9153 = ~\P1_P3_InstQueueRd_Addr_reg[2]/NET0131  & ~n9049 ;
  assign n9154 = n9049 & n9104 ;
  assign n9155 = ~n9153 & ~n9154 ;
  assign n9156 = ~n9061 & n9155 ;
  assign n9157 = ~n9152 & ~n9156 ;
  assign n9158 = ~n9146 & n9157 ;
  assign n9159 = ~n9139 & n9158 ;
  assign n9160 = ~n9134 & n9159 ;
  assign n9203 = \P1_P3_InstQueueWr_Addr_reg[2]/NET0131  & n9160 ;
  assign n9228 = \P1_P3_InstQueueWr_Addr_reg[1]/NET0131  & n9218 ;
  assign n9229 = ~n9203 & ~n9228 ;
  assign n9230 = ~n9200 & n9229 ;
  assign n9231 = ~n9227 & n9230 ;
  assign n9201 = ~\P1_P3_InstQueueWr_Addr_reg[2]/NET0131  & ~n9160 ;
  assign n9202 = ~n9200 & n9201 ;
  assign n9161 = \P1_P3_InstQueueWr_Addr_reg[3]/NET0131  & n9160 ;
  assign n9190 = ~n9161 & ~n9189 ;
  assign n9089 = ~n9087 & ~n9088 ;
  assign n9090 = n9084 & ~n9089 ;
  assign n9076 = ~\P1_P3_More_reg/NET0131  & ~n9075 ;
  assign n9098 = ~n9076 & ~n9097 ;
  assign n9099 = ~n9090 & n9098 ;
  assign n9050 = n9021 & ~n9049 ;
  assign n9071 = ~n9043 & n9070 ;
  assign n9072 = ~n9066 & ~n9071 ;
  assign n9073 = n9064 & n9072 ;
  assign n9074 = ~n9062 & ~n9073 ;
  assign n9100 = ~n9050 & n9074 ;
  assign n9101 = ~n9099 & n9100 ;
  assign n9195 = ~n9075 & ~n9116 ;
  assign n9193 = ~n9084 & n9095 ;
  assign n9194 = ~n8741 & ~n9193 ;
  assign n9196 = \P1_P3_Flush_reg/NET0131  & ~n9194 ;
  assign n9197 = n9195 & n9196 ;
  assign n9191 = n9021 & n9049 ;
  assign n9192 = n9064 & ~n9072 ;
  assign n9198 = ~n9191 & ~n9192 ;
  assign n9199 = ~n9197 & n9198 ;
  assign n9232 = n9101 & n9199 ;
  assign n9233 = ~n9190 & n9232 ;
  assign n9234 = ~n9202 & n9233 ;
  assign n9235 = ~n9231 & n9234 ;
  assign n9236 = ~n9075 & n9079 ;
  assign n9237 = ~\P1_P3_DataWidth_reg[1]/NET0131  & n9236 ;
  assign n9238 = n9096 & n9237 ;
  assign n9239 = n9235 & ~n9238 ;
  assign n8731 = \P1_P3_State2_reg[0]/NET0131  & ~\P1_P3_State2_reg[3]/NET0131  ;
  assign n9240 = ~\P1_P3_State2_reg[1]/NET0131  & \P1_P3_State2_reg[2]/NET0131  ;
  assign n9241 = n8731 & n9240 ;
  assign n9242 = ~n9239 & n9241 ;
  assign n8732 = ~\P1_P3_State2_reg[2]/NET0131  & n8731 ;
  assign n9247 = ~\P1_P3_State2_reg[1]/NET0131  & n8732 ;
  assign n9248 = ~n8741 & n9247 ;
  assign n8733 = ~\P1_P3_State2_reg[0]/NET0131  & ~\P1_P3_State2_reg[3]/NET0131  ;
  assign n8734 = \P1_P3_State2_reg[2]/NET0131  & n8733 ;
  assign n8735 = ~n8732 & ~n8734 ;
  assign n8736 = \P1_P3_State2_reg[1]/NET0131  & ~n8735 ;
  assign n8742 = n8736 & n8741 ;
  assign n9243 = ~\P1_P3_State2_reg[2]/NET0131  & ~\P1_P3_State2_reg[3]/NET0131  ;
  assign n9244 = \P1_P3_State2_reg[1]/NET0131  & n9243 ;
  assign n9245 = ~\P1_P3_State2_reg[0]/NET0131  & n9244 ;
  assign n9246 = ~\P1_P3_DataWidth_reg[1]/NET0131  & n9245 ;
  assign n9249 = ~n8742 & ~n9246 ;
  assign n9250 = ~n9248 & n9249 ;
  assign n9251 = ~n9242 & n9250 ;
  assign n9261 = n8069 & ~n8077 ;
  assign n9262 = n8092 & ~n9261 ;
  assign n9263 = ~n8094 & ~n9262 ;
  assign n9264 = n4327 & ~n9263 ;
  assign n9256 = ~n7940 & ~n8146 ;
  assign n9257 = \P1_P1_InstQueue_reg[11][4]/NET0131  & ~n8142 ;
  assign n9258 = ~n8145 & n9257 ;
  assign n9259 = ~n9256 & ~n9258 ;
  assign n9260 = ~n4327 & n9259 ;
  assign n9265 = ~n8139 & ~n9260 ;
  assign n9266 = ~n9264 & n9265 ;
  assign n9252 = n8207 & ~n8232 ;
  assign n9253 = n8223 & ~n9252 ;
  assign n9254 = ~n8234 & ~n9253 ;
  assign n9255 = n8139 & n9254 ;
  assign n9267 = \P1_P1_DataWidth_reg[1]/NET0131  & ~n9255 ;
  assign n9268 = ~n9266 & n9267 ;
  assign n9269 = ~\P1_P1_DataWidth_reg[1]/NET0131  & n9259 ;
  assign n9270 = n8282 & ~n9269 ;
  assign n9271 = ~n9268 & n9270 ;
  assign n9272 = n8287 & ~n9259 ;
  assign n9273 = \P1_P1_InstQueue_reg[14][4]/NET0131  & n8291 ;
  assign n9274 = \P1_P1_InstQueue_reg[2][4]/NET0131  & n8314 ;
  assign n9275 = \P1_P1_InstQueue_reg[8][4]/NET0131  & n8305 ;
  assign n9289 = ~n9274 & ~n9275 ;
  assign n9276 = \P1_P1_InstQueue_reg[11][4]/NET0131  & n8312 ;
  assign n9277 = \P1_P1_InstQueue_reg[3][4]/NET0131  & n8323 ;
  assign n9290 = ~n9276 & ~n9277 ;
  assign n9299 = n9289 & n9290 ;
  assign n9300 = ~n9273 & n9299 ;
  assign n9288 = \P1_P1_InstQueue_reg[0][4]/NET0131  & n8309 ;
  assign n9286 = \P1_P1_InstQueue_reg[9][4]/NET0131  & n8325 ;
  assign n9287 = \P1_P1_InstQueue_reg[4][4]/NET0131  & n8295 ;
  assign n9295 = ~n9286 & ~n9287 ;
  assign n9296 = ~n9288 & n9295 ;
  assign n9282 = \P1_P1_InstQueue_reg[6][4]/NET0131  & n8316 ;
  assign n9283 = \P1_P1_InstQueue_reg[15][4]/NET0131  & n8321 ;
  assign n9293 = ~n9282 & ~n9283 ;
  assign n9284 = \P1_P1_InstQueue_reg[7][4]/NET0131  & n8318 ;
  assign n9285 = \P1_P1_InstQueue_reg[13][4]/NET0131  & n8327 ;
  assign n9294 = ~n9284 & ~n9285 ;
  assign n9297 = n9293 & n9294 ;
  assign n9278 = \P1_P1_InstQueue_reg[12][4]/NET0131  & n8329 ;
  assign n9279 = \P1_P1_InstQueue_reg[10][4]/NET0131  & n8303 ;
  assign n9291 = ~n9278 & ~n9279 ;
  assign n9280 = \P1_P1_InstQueue_reg[1][4]/NET0131  & n8299 ;
  assign n9281 = \P1_P1_InstQueue_reg[5][4]/NET0131  & n8307 ;
  assign n9292 = ~n9280 & ~n9281 ;
  assign n9298 = n9291 & n9292 ;
  assign n9301 = n9297 & n9298 ;
  assign n9302 = n9296 & n9301 ;
  assign n9303 = n9300 & n9302 ;
  assign n9304 = n8142 & ~n9303 ;
  assign n9305 = ~n9257 & ~n9304 ;
  assign n9306 = n8350 & ~n9305 ;
  assign n9307 = \P1_P1_InstQueue_reg[11][4]/NET0131  & ~n8366 ;
  assign n9308 = ~n9306 & ~n9307 ;
  assign n9309 = ~n9272 & n9308 ;
  assign n9310 = ~n9271 & n9309 ;
  assign n9311 = n8094 & ~n8106 ;
  assign n9312 = n8121 & ~n9311 ;
  assign n9313 = ~n8123 & ~n9312 ;
  assign n9314 = n4327 & ~n9313 ;
  assign n9315 = n7906 & ~n8146 ;
  assign n9316 = \P1_P1_InstQueue_reg[11][6]/NET0131  & ~n8142 ;
  assign n9317 = ~n8145 & n9316 ;
  assign n9318 = ~n9315 & ~n9317 ;
  assign n9319 = ~n4327 & n9318 ;
  assign n9320 = ~n8139 & ~n9319 ;
  assign n9321 = ~n9314 & n9320 ;
  assign n9322 = n8234 & ~n8248 ;
  assign n9323 = n8270 & ~n9322 ;
  assign n9324 = ~n8272 & ~n9323 ;
  assign n9325 = n8139 & n9324 ;
  assign n9326 = \P1_P1_DataWidth_reg[1]/NET0131  & ~n9325 ;
  assign n9327 = ~n9321 & n9326 ;
  assign n9328 = ~\P1_P1_DataWidth_reg[1]/NET0131  & n9318 ;
  assign n9329 = n8282 & ~n9328 ;
  assign n9330 = ~n9327 & n9329 ;
  assign n9331 = n8287 & ~n9318 ;
  assign n9332 = \P1_P1_InstQueue_reg[14][6]/NET0131  & n8291 ;
  assign n9333 = \P1_P1_InstQueue_reg[13][6]/NET0131  & n8327 ;
  assign n9334 = \P1_P1_InstQueue_reg[4][6]/NET0131  & n8295 ;
  assign n9348 = ~n9333 & ~n9334 ;
  assign n9335 = \P1_P1_InstQueue_reg[12][6]/NET0131  & n8329 ;
  assign n9336 = \P1_P1_InstQueue_reg[11][6]/NET0131  & n8312 ;
  assign n9349 = ~n9335 & ~n9336 ;
  assign n9358 = n9348 & n9349 ;
  assign n9359 = ~n9332 & n9358 ;
  assign n9347 = \P1_P1_InstQueue_reg[10][6]/NET0131  & n8303 ;
  assign n9345 = \P1_P1_InstQueue_reg[1][6]/NET0131  & n8299 ;
  assign n9346 = \P1_P1_InstQueue_reg[5][6]/NET0131  & n8307 ;
  assign n9354 = ~n9345 & ~n9346 ;
  assign n9355 = ~n9347 & n9354 ;
  assign n9341 = \P1_P1_InstQueue_reg[6][6]/NET0131  & n8316 ;
  assign n9342 = \P1_P1_InstQueue_reg[15][6]/NET0131  & n8321 ;
  assign n9352 = ~n9341 & ~n9342 ;
  assign n9343 = \P1_P1_InstQueue_reg[7][6]/NET0131  & n8318 ;
  assign n9344 = \P1_P1_InstQueue_reg[9][6]/NET0131  & n8325 ;
  assign n9353 = ~n9343 & ~n9344 ;
  assign n9356 = n9352 & n9353 ;
  assign n9337 = \P1_P1_InstQueue_reg[8][6]/NET0131  & n8305 ;
  assign n9338 = \P1_P1_InstQueue_reg[2][6]/NET0131  & n8314 ;
  assign n9350 = ~n9337 & ~n9338 ;
  assign n9339 = \P1_P1_InstQueue_reg[3][6]/NET0131  & n8323 ;
  assign n9340 = \P1_P1_InstQueue_reg[0][6]/NET0131  & n8309 ;
  assign n9351 = ~n9339 & ~n9340 ;
  assign n9357 = n9350 & n9351 ;
  assign n9360 = n9356 & n9357 ;
  assign n9361 = n9355 & n9360 ;
  assign n9362 = n9359 & n9361 ;
  assign n9363 = n8142 & ~n9362 ;
  assign n9364 = ~n9316 & ~n9363 ;
  assign n9365 = n8350 & ~n9364 ;
  assign n9366 = \P1_P1_InstQueue_reg[11][6]/NET0131  & ~n8366 ;
  assign n9367 = ~n9365 & ~n9366 ;
  assign n9368 = ~n9331 & n9367 ;
  assign n9369 = ~n9330 & n9368 ;
  assign n9376 = n8372 & ~n9263 ;
  assign n9371 = ~n7940 & ~n8379 ;
  assign n9372 = \P1_P1_InstQueue_reg[0][4]/NET0131  & ~n8376 ;
  assign n9373 = ~n8378 & n9372 ;
  assign n9374 = ~n9371 & ~n9373 ;
  assign n9375 = ~n8372 & n9374 ;
  assign n9377 = ~n8375 & ~n9375 ;
  assign n9378 = ~n9376 & n9377 ;
  assign n9370 = n8375 & n9254 ;
  assign n9379 = \P1_P1_DataWidth_reg[1]/NET0131  & ~n9370 ;
  assign n9380 = ~n9378 & n9379 ;
  assign n9381 = ~\P1_P1_DataWidth_reg[1]/NET0131  & n9374 ;
  assign n9382 = n8282 & ~n9381 ;
  assign n9383 = ~n9380 & n9382 ;
  assign n9384 = n8287 & ~n9374 ;
  assign n9385 = n8376 & ~n9303 ;
  assign n9386 = ~n9372 & ~n9385 ;
  assign n9387 = n8350 & ~n9386 ;
  assign n9388 = \P1_P1_InstQueue_reg[0][4]/NET0131  & ~n8366 ;
  assign n9389 = ~n9387 & ~n9388 ;
  assign n9390 = ~n9384 & n9389 ;
  assign n9391 = ~n9383 & n9390 ;
  assign n9392 = n8372 & ~n9313 ;
  assign n9393 = n7906 & ~n8379 ;
  assign n9394 = \P1_P1_InstQueue_reg[0][6]/NET0131  & ~n8376 ;
  assign n9395 = ~n8378 & n9394 ;
  assign n9396 = ~n9393 & ~n9395 ;
  assign n9397 = ~n8372 & n9396 ;
  assign n9398 = ~n8375 & ~n9397 ;
  assign n9399 = ~n9392 & n9398 ;
  assign n9400 = n8375 & n9324 ;
  assign n9401 = \P1_P1_DataWidth_reg[1]/NET0131  & ~n9400 ;
  assign n9402 = ~n9399 & n9401 ;
  assign n9403 = ~\P1_P1_DataWidth_reg[1]/NET0131  & n9396 ;
  assign n9404 = n8282 & ~n9403 ;
  assign n9405 = ~n9402 & n9404 ;
  assign n9406 = n8287 & ~n9396 ;
  assign n9407 = n8376 & ~n9362 ;
  assign n9408 = ~n9394 & ~n9407 ;
  assign n9409 = n8350 & ~n9408 ;
  assign n9410 = \P1_P1_InstQueue_reg[0][6]/NET0131  & ~n8366 ;
  assign n9411 = ~n9409 & ~n9410 ;
  assign n9412 = ~n9406 & n9411 ;
  assign n9413 = ~n9405 & n9412 ;
  assign n9414 = n8407 & n9254 ;
  assign n9415 = n8139 & n9263 ;
  assign n9416 = ~n9414 & ~n9415 ;
  assign n9417 = \P1_P1_DataWidth_reg[1]/NET0131  & ~n9416 ;
  assign n9418 = \P1_P1_DataWidth_reg[1]/NET0131  & ~n8410 ;
  assign n9419 = ~n7940 & ~n8401 ;
  assign n9420 = \P1_P1_InstQueue_reg[10][4]/NET0131  & ~n8145 ;
  assign n9421 = ~n4327 & n9420 ;
  assign n9422 = ~n9419 & ~n9421 ;
  assign n9423 = ~n9418 & ~n9422 ;
  assign n9424 = ~n9417 & ~n9423 ;
  assign n9425 = n8282 & ~n9424 ;
  assign n9427 = n8287 & ~n9422 ;
  assign n9426 = \P1_P1_InstQueue_reg[10][4]/NET0131  & ~n8366 ;
  assign n9428 = n8145 & ~n9303 ;
  assign n9429 = ~n9420 & ~n9428 ;
  assign n9430 = n8350 & ~n9429 ;
  assign n9431 = ~n9426 & ~n9430 ;
  assign n9432 = ~n9427 & n9431 ;
  assign n9433 = ~n9425 & n9432 ;
  assign n9440 = n8139 & n9313 ;
  assign n9439 = n8407 & n9324 ;
  assign n9434 = n7906 & ~n8401 ;
  assign n9435 = \P1_P1_InstQueue_reg[10][6]/NET0131  & ~n8145 ;
  assign n9436 = ~n4327 & n9435 ;
  assign n9437 = ~n9434 & ~n9436 ;
  assign n9441 = n8410 & ~n9437 ;
  assign n9442 = \P1_P1_DataWidth_reg[1]/NET0131  & ~n9441 ;
  assign n9443 = ~n9439 & n9442 ;
  assign n9444 = ~n9440 & n9443 ;
  assign n9438 = ~\P1_P1_DataWidth_reg[1]/NET0131  & n9437 ;
  assign n9445 = n8282 & ~n9438 ;
  assign n9446 = ~n9444 & n9445 ;
  assign n9447 = n8287 & ~n9437 ;
  assign n9448 = n8145 & ~n9362 ;
  assign n9449 = ~n9435 & ~n9448 ;
  assign n9450 = n8350 & ~n9449 ;
  assign n9451 = \P1_P1_InstQueue_reg[10][6]/NET0131  & ~n8366 ;
  assign n9452 = ~n9450 & ~n9451 ;
  assign n9453 = ~n9447 & n9452 ;
  assign n9454 = ~n9446 & n9453 ;
  assign n9461 = n8145 & ~n9263 ;
  assign n9456 = ~n7940 & ~n8428 ;
  assign n9457 = \P1_P1_InstQueue_reg[12][4]/NET0131  & ~n8427 ;
  assign n9458 = ~n8142 & n9457 ;
  assign n9459 = ~n9456 & ~n9458 ;
  assign n9460 = ~n8145 & n9459 ;
  assign n9462 = ~n4327 & ~n9460 ;
  assign n9463 = ~n9461 & n9462 ;
  assign n9455 = n4327 & n9254 ;
  assign n9464 = \P1_P1_DataWidth_reg[1]/NET0131  & ~n9455 ;
  assign n9465 = ~n9463 & n9464 ;
  assign n9466 = ~\P1_P1_DataWidth_reg[1]/NET0131  & n9459 ;
  assign n9467 = n8282 & ~n9466 ;
  assign n9468 = ~n9465 & n9467 ;
  assign n9469 = n8287 & ~n9459 ;
  assign n9470 = n8427 & ~n9303 ;
  assign n9471 = ~n9457 & ~n9470 ;
  assign n9472 = n8350 & ~n9471 ;
  assign n9473 = \P1_P1_InstQueue_reg[12][4]/NET0131  & ~n8366 ;
  assign n9474 = ~n9472 & ~n9473 ;
  assign n9475 = ~n9469 & n9474 ;
  assign n9476 = ~n9468 & n9475 ;
  assign n9477 = n8145 & ~n9313 ;
  assign n9478 = n7906 & ~n8428 ;
  assign n9479 = \P1_P1_InstQueue_reg[12][6]/NET0131  & ~n8427 ;
  assign n9480 = ~n8142 & n9479 ;
  assign n9481 = ~n9478 & ~n9480 ;
  assign n9482 = ~n8145 & n9481 ;
  assign n9483 = ~n4327 & ~n9482 ;
  assign n9484 = ~n9477 & n9483 ;
  assign n9485 = n4327 & n9324 ;
  assign n9486 = \P1_P1_DataWidth_reg[1]/NET0131  & ~n9485 ;
  assign n9487 = ~n9484 & n9486 ;
  assign n9488 = ~\P1_P1_DataWidth_reg[1]/NET0131  & n9481 ;
  assign n9489 = n8282 & ~n9488 ;
  assign n9490 = ~n9487 & n9489 ;
  assign n9491 = n8287 & ~n9481 ;
  assign n9492 = n8427 & ~n9362 ;
  assign n9493 = ~n9479 & ~n9492 ;
  assign n9494 = n8350 & ~n9493 ;
  assign n9495 = \P1_P1_InstQueue_reg[12][6]/NET0131  & ~n8366 ;
  assign n9496 = ~n9494 & ~n9495 ;
  assign n9497 = ~n9491 & n9496 ;
  assign n9498 = ~n9490 & n9497 ;
  assign n9499 = n8142 & ~n9313 ;
  assign n9500 = n7906 & ~n8451 ;
  assign n9501 = \P1_P1_InstQueue_reg[13][6]/NET0131  & ~n8375 ;
  assign n9502 = ~n8427 & n9501 ;
  assign n9503 = ~n9500 & ~n9502 ;
  assign n9504 = ~n8142 & n9503 ;
  assign n9505 = ~n8145 & ~n9504 ;
  assign n9506 = ~n9499 & n9505 ;
  assign n9507 = n8145 & n9324 ;
  assign n9508 = \P1_P1_DataWidth_reg[1]/NET0131  & ~n9507 ;
  assign n9509 = ~n9506 & n9508 ;
  assign n9510 = ~\P1_P1_DataWidth_reg[1]/NET0131  & n9503 ;
  assign n9511 = n8282 & ~n9510 ;
  assign n9512 = ~n9509 & n9511 ;
  assign n9513 = n8287 & ~n9503 ;
  assign n9514 = n8375 & ~n9362 ;
  assign n9515 = ~n9501 & ~n9514 ;
  assign n9516 = n8350 & ~n9515 ;
  assign n9517 = \P1_P1_InstQueue_reg[13][6]/NET0131  & ~n8366 ;
  assign n9518 = ~n9516 & ~n9517 ;
  assign n9519 = ~n9513 & n9518 ;
  assign n9520 = ~n9512 & n9519 ;
  assign n9527 = n8142 & ~n9263 ;
  assign n9522 = ~n7940 & ~n8451 ;
  assign n9523 = \P1_P1_InstQueue_reg[13][4]/NET0131  & ~n8375 ;
  assign n9524 = ~n8427 & n9523 ;
  assign n9525 = ~n9522 & ~n9524 ;
  assign n9526 = ~n8142 & n9525 ;
  assign n9528 = ~n8145 & ~n9526 ;
  assign n9529 = ~n9527 & n9528 ;
  assign n9521 = n8145 & n9254 ;
  assign n9530 = \P1_P1_DataWidth_reg[1]/NET0131  & ~n9521 ;
  assign n9531 = ~n9529 & n9530 ;
  assign n9532 = ~\P1_P1_DataWidth_reg[1]/NET0131  & n9525 ;
  assign n9533 = n8282 & ~n9532 ;
  assign n9534 = ~n9531 & n9533 ;
  assign n9535 = n8287 & ~n9525 ;
  assign n9536 = n8375 & ~n9303 ;
  assign n9537 = ~n9523 & ~n9536 ;
  assign n9538 = n8350 & ~n9537 ;
  assign n9539 = \P1_P1_InstQueue_reg[13][4]/NET0131  & ~n8366 ;
  assign n9540 = ~n9538 & ~n9539 ;
  assign n9541 = ~n9535 & n9540 ;
  assign n9542 = ~n9534 & n9541 ;
  assign n9549 = n8427 & ~n9263 ;
  assign n9544 = ~n7940 & ~n8474 ;
  assign n9545 = \P1_P1_InstQueue_reg[14][4]/NET0131  & ~n8372 ;
  assign n9546 = ~n8375 & n9545 ;
  assign n9547 = ~n9544 & ~n9546 ;
  assign n9548 = ~n8427 & n9547 ;
  assign n9550 = ~n8142 & ~n9548 ;
  assign n9551 = ~n9549 & n9550 ;
  assign n9543 = n8142 & n9254 ;
  assign n9552 = \P1_P1_DataWidth_reg[1]/NET0131  & ~n9543 ;
  assign n9553 = ~n9551 & n9552 ;
  assign n9554 = ~\P1_P1_DataWidth_reg[1]/NET0131  & n9547 ;
  assign n9555 = n8282 & ~n9554 ;
  assign n9556 = ~n9553 & n9555 ;
  assign n9557 = n8287 & ~n9547 ;
  assign n9558 = n8372 & ~n9303 ;
  assign n9559 = ~n9545 & ~n9558 ;
  assign n9560 = n8350 & ~n9559 ;
  assign n9561 = \P1_P1_InstQueue_reg[14][4]/NET0131  & ~n8366 ;
  assign n9562 = ~n9560 & ~n9561 ;
  assign n9563 = ~n9557 & n9562 ;
  assign n9564 = ~n9556 & n9563 ;
  assign n9565 = n8427 & ~n9313 ;
  assign n9566 = n7906 & ~n8474 ;
  assign n9567 = \P1_P1_InstQueue_reg[14][6]/NET0131  & ~n8372 ;
  assign n9568 = ~n8375 & n9567 ;
  assign n9569 = ~n9566 & ~n9568 ;
  assign n9570 = ~n8427 & n9569 ;
  assign n9571 = ~n8142 & ~n9570 ;
  assign n9572 = ~n9565 & n9571 ;
  assign n9573 = n8142 & n9324 ;
  assign n9574 = \P1_P1_DataWidth_reg[1]/NET0131  & ~n9573 ;
  assign n9575 = ~n9572 & n9574 ;
  assign n9576 = ~\P1_P1_DataWidth_reg[1]/NET0131  & n9569 ;
  assign n9577 = n8282 & ~n9576 ;
  assign n9578 = ~n9575 & n9577 ;
  assign n9579 = n8287 & ~n9569 ;
  assign n9580 = n8372 & ~n9362 ;
  assign n9581 = ~n9567 & ~n9580 ;
  assign n9582 = n8350 & ~n9581 ;
  assign n9583 = \P1_P1_InstQueue_reg[14][6]/NET0131  & ~n8366 ;
  assign n9584 = ~n9582 & ~n9583 ;
  assign n9585 = ~n9579 & n9584 ;
  assign n9586 = ~n9578 & n9585 ;
  assign n9593 = n8375 & ~n9263 ;
  assign n9588 = ~n7940 & ~n8497 ;
  assign n9589 = \P1_P1_InstQueue_reg[15][4]/NET0131  & ~n8378 ;
  assign n9590 = ~n8372 & n9589 ;
  assign n9591 = ~n9588 & ~n9590 ;
  assign n9592 = ~n8375 & n9591 ;
  assign n9594 = ~n8427 & ~n9592 ;
  assign n9595 = ~n9593 & n9594 ;
  assign n9587 = n8427 & n9254 ;
  assign n9596 = \P1_P1_DataWidth_reg[1]/NET0131  & ~n9587 ;
  assign n9597 = ~n9595 & n9596 ;
  assign n9598 = ~\P1_P1_DataWidth_reg[1]/NET0131  & n9591 ;
  assign n9599 = n8282 & ~n9598 ;
  assign n9600 = ~n9597 & n9599 ;
  assign n9601 = n8287 & ~n9591 ;
  assign n9602 = n8378 & ~n9303 ;
  assign n9603 = ~n9589 & ~n9602 ;
  assign n9604 = n8350 & ~n9603 ;
  assign n9605 = \P1_P1_InstQueue_reg[15][4]/NET0131  & ~n8366 ;
  assign n9606 = ~n9604 & ~n9605 ;
  assign n9607 = ~n9601 & n9606 ;
  assign n9608 = ~n9600 & n9607 ;
  assign n9609 = n8375 & ~n9313 ;
  assign n9610 = n7906 & ~n8497 ;
  assign n9611 = \P1_P1_InstQueue_reg[15][6]/NET0131  & ~n8378 ;
  assign n9612 = ~n8372 & n9611 ;
  assign n9613 = ~n9610 & ~n9612 ;
  assign n9614 = ~n8375 & n9613 ;
  assign n9615 = ~n8427 & ~n9614 ;
  assign n9616 = ~n9609 & n9615 ;
  assign n9617 = n8427 & n9324 ;
  assign n9618 = \P1_P1_DataWidth_reg[1]/NET0131  & ~n9617 ;
  assign n9619 = ~n9616 & n9618 ;
  assign n9620 = ~\P1_P1_DataWidth_reg[1]/NET0131  & n9613 ;
  assign n9621 = n8282 & ~n9620 ;
  assign n9622 = ~n9619 & n9621 ;
  assign n9623 = n8287 & ~n9613 ;
  assign n9624 = n8378 & ~n9362 ;
  assign n9625 = ~n9611 & ~n9624 ;
  assign n9626 = n8350 & ~n9625 ;
  assign n9627 = \P1_P1_InstQueue_reg[15][6]/NET0131  & ~n8366 ;
  assign n9628 = ~n9626 & ~n9627 ;
  assign n9629 = ~n9623 & n9628 ;
  assign n9630 = ~n9622 & n9629 ;
  assign n9637 = n8378 & ~n9263 ;
  assign n9632 = ~n7940 & ~n8521 ;
  assign n9633 = \P1_P1_InstQueue_reg[1][4]/NET0131  & ~n8520 ;
  assign n9634 = ~n8376 & n9633 ;
  assign n9635 = ~n9632 & ~n9634 ;
  assign n9636 = ~n8378 & n9635 ;
  assign n9638 = ~n8372 & ~n9636 ;
  assign n9639 = ~n9637 & n9638 ;
  assign n9631 = n8372 & n9254 ;
  assign n9640 = \P1_P1_DataWidth_reg[1]/NET0131  & ~n9631 ;
  assign n9641 = ~n9639 & n9640 ;
  assign n9642 = ~\P1_P1_DataWidth_reg[1]/NET0131  & n9635 ;
  assign n9643 = n8282 & ~n9642 ;
  assign n9644 = ~n9641 & n9643 ;
  assign n9645 = n8287 & ~n9635 ;
  assign n9646 = n8520 & ~n9303 ;
  assign n9647 = ~n9633 & ~n9646 ;
  assign n9648 = n8350 & ~n9647 ;
  assign n9649 = \P1_P1_InstQueue_reg[1][4]/NET0131  & ~n8366 ;
  assign n9650 = ~n9648 & ~n9649 ;
  assign n9651 = ~n9645 & n9650 ;
  assign n9652 = ~n9644 & n9651 ;
  assign n9653 = n8378 & ~n9313 ;
  assign n9654 = n7906 & ~n8521 ;
  assign n9655 = \P1_P1_InstQueue_reg[1][6]/NET0131  & ~n8520 ;
  assign n9656 = ~n8376 & n9655 ;
  assign n9657 = ~n9654 & ~n9656 ;
  assign n9658 = ~n8378 & n9657 ;
  assign n9659 = ~n8372 & ~n9658 ;
  assign n9660 = ~n9653 & n9659 ;
  assign n9661 = n8372 & n9324 ;
  assign n9662 = \P1_P1_DataWidth_reg[1]/NET0131  & ~n9661 ;
  assign n9663 = ~n9660 & n9662 ;
  assign n9664 = ~\P1_P1_DataWidth_reg[1]/NET0131  & n9657 ;
  assign n9665 = n8282 & ~n9664 ;
  assign n9666 = ~n9663 & n9665 ;
  assign n9667 = n8287 & ~n9657 ;
  assign n9668 = n8520 & ~n9362 ;
  assign n9669 = ~n9655 & ~n9668 ;
  assign n9670 = n8350 & ~n9669 ;
  assign n9671 = \P1_P1_InstQueue_reg[1][6]/NET0131  & ~n8366 ;
  assign n9672 = ~n9670 & ~n9671 ;
  assign n9673 = ~n9667 & n9672 ;
  assign n9674 = ~n9666 & n9673 ;
  assign n9675 = n8376 & ~n9313 ;
  assign n9676 = n7906 & ~n8545 ;
  assign n9677 = \P1_P1_InstQueue_reg[2][6]/NET0131  & ~n8544 ;
  assign n9678 = ~n8520 & n9677 ;
  assign n9679 = ~n9676 & ~n9678 ;
  assign n9680 = ~n8376 & n9679 ;
  assign n9681 = ~n8378 & ~n9680 ;
  assign n9682 = ~n9675 & n9681 ;
  assign n9683 = n8378 & n9324 ;
  assign n9684 = \P1_P1_DataWidth_reg[1]/NET0131  & ~n9683 ;
  assign n9685 = ~n9682 & n9684 ;
  assign n9686 = ~\P1_P1_DataWidth_reg[1]/NET0131  & n9679 ;
  assign n9687 = n8282 & ~n9686 ;
  assign n9688 = ~n9685 & n9687 ;
  assign n9689 = n8287 & ~n9679 ;
  assign n9690 = n8544 & ~n9362 ;
  assign n9691 = ~n9677 & ~n9690 ;
  assign n9692 = n8350 & ~n9691 ;
  assign n9693 = \P1_P1_InstQueue_reg[2][6]/NET0131  & ~n8366 ;
  assign n9694 = ~n9692 & ~n9693 ;
  assign n9695 = ~n9689 & n9694 ;
  assign n9696 = ~n9688 & n9695 ;
  assign n9703 = n8376 & ~n9263 ;
  assign n9698 = ~n7940 & ~n8545 ;
  assign n9699 = \P1_P1_InstQueue_reg[2][4]/NET0131  & ~n8544 ;
  assign n9700 = ~n8520 & n9699 ;
  assign n9701 = ~n9698 & ~n9700 ;
  assign n9702 = ~n8376 & n9701 ;
  assign n9704 = ~n8378 & ~n9702 ;
  assign n9705 = ~n9703 & n9704 ;
  assign n9697 = n8378 & n9254 ;
  assign n9706 = \P1_P1_DataWidth_reg[1]/NET0131  & ~n9697 ;
  assign n9707 = ~n9705 & n9706 ;
  assign n9708 = ~\P1_P1_DataWidth_reg[1]/NET0131  & n9701 ;
  assign n9709 = n8282 & ~n9708 ;
  assign n9710 = ~n9707 & n9709 ;
  assign n9711 = n8287 & ~n9701 ;
  assign n9712 = n8544 & ~n9303 ;
  assign n9713 = ~n9699 & ~n9712 ;
  assign n9714 = n8350 & ~n9713 ;
  assign n9715 = \P1_P1_InstQueue_reg[2][4]/NET0131  & ~n8366 ;
  assign n9716 = ~n9714 & ~n9715 ;
  assign n9717 = ~n9711 & n9716 ;
  assign n9718 = ~n9710 & n9717 ;
  assign n9719 = n8520 & ~n9313 ;
  assign n9720 = n7906 & ~n8569 ;
  assign n9721 = \P1_P1_InstQueue_reg[3][6]/NET0131  & ~n8568 ;
  assign n9722 = ~n8544 & n9721 ;
  assign n9723 = ~n9720 & ~n9722 ;
  assign n9724 = ~n8520 & n9723 ;
  assign n9725 = ~n8376 & ~n9724 ;
  assign n9726 = ~n9719 & n9725 ;
  assign n9727 = n8376 & n9324 ;
  assign n9728 = \P1_P1_DataWidth_reg[1]/NET0131  & ~n9727 ;
  assign n9729 = ~n9726 & n9728 ;
  assign n9730 = ~\P1_P1_DataWidth_reg[1]/NET0131  & n9723 ;
  assign n9731 = n8282 & ~n9730 ;
  assign n9732 = ~n9729 & n9731 ;
  assign n9733 = n8287 & ~n9723 ;
  assign n9734 = n8568 & ~n9362 ;
  assign n9735 = ~n9721 & ~n9734 ;
  assign n9736 = n8350 & ~n9735 ;
  assign n9737 = \P1_P1_InstQueue_reg[3][6]/NET0131  & ~n8366 ;
  assign n9738 = ~n9736 & ~n9737 ;
  assign n9739 = ~n9733 & n9738 ;
  assign n9740 = ~n9732 & n9739 ;
  assign n9747 = n8520 & ~n9263 ;
  assign n9742 = ~n7940 & ~n8569 ;
  assign n9743 = \P1_P1_InstQueue_reg[3][4]/NET0131  & ~n8568 ;
  assign n9744 = ~n8544 & n9743 ;
  assign n9745 = ~n9742 & ~n9744 ;
  assign n9746 = ~n8520 & n9745 ;
  assign n9748 = ~n8376 & ~n9746 ;
  assign n9749 = ~n9747 & n9748 ;
  assign n9741 = n8376 & n9254 ;
  assign n9750 = \P1_P1_DataWidth_reg[1]/NET0131  & ~n9741 ;
  assign n9751 = ~n9749 & n9750 ;
  assign n9752 = ~\P1_P1_DataWidth_reg[1]/NET0131  & n9745 ;
  assign n9753 = n8282 & ~n9752 ;
  assign n9754 = ~n9751 & n9753 ;
  assign n9755 = n8287 & ~n9745 ;
  assign n9756 = n8568 & ~n9303 ;
  assign n9757 = ~n9743 & ~n9756 ;
  assign n9758 = n8350 & ~n9757 ;
  assign n9759 = \P1_P1_InstQueue_reg[3][4]/NET0131  & ~n8366 ;
  assign n9760 = ~n9758 & ~n9759 ;
  assign n9761 = ~n9755 & n9760 ;
  assign n9762 = ~n9754 & n9761 ;
  assign n9769 = n8544 & ~n9263 ;
  assign n9764 = ~n7940 & ~n8593 ;
  assign n9765 = \P1_P1_InstQueue_reg[4][4]/NET0131  & ~n8592 ;
  assign n9766 = ~n8568 & n9765 ;
  assign n9767 = ~n9764 & ~n9766 ;
  assign n9768 = ~n8544 & n9767 ;
  assign n9770 = ~n8520 & ~n9768 ;
  assign n9771 = ~n9769 & n9770 ;
  assign n9763 = n8520 & n9254 ;
  assign n9772 = \P1_P1_DataWidth_reg[1]/NET0131  & ~n9763 ;
  assign n9773 = ~n9771 & n9772 ;
  assign n9774 = ~\P1_P1_DataWidth_reg[1]/NET0131  & n9767 ;
  assign n9775 = n8282 & ~n9774 ;
  assign n9776 = ~n9773 & n9775 ;
  assign n9777 = n8287 & ~n9767 ;
  assign n9778 = n8592 & ~n9303 ;
  assign n9779 = ~n9765 & ~n9778 ;
  assign n9780 = n8350 & ~n9779 ;
  assign n9781 = \P1_P1_InstQueue_reg[4][4]/NET0131  & ~n8366 ;
  assign n9782 = ~n9780 & ~n9781 ;
  assign n9783 = ~n9777 & n9782 ;
  assign n9784 = ~n9776 & n9783 ;
  assign n9785 = n8544 & ~n9313 ;
  assign n9786 = n7906 & ~n8593 ;
  assign n9787 = \P1_P1_InstQueue_reg[4][6]/NET0131  & ~n8592 ;
  assign n9788 = ~n8568 & n9787 ;
  assign n9789 = ~n9786 & ~n9788 ;
  assign n9790 = ~n8544 & n9789 ;
  assign n9791 = ~n8520 & ~n9790 ;
  assign n9792 = ~n9785 & n9791 ;
  assign n9793 = n8520 & n9324 ;
  assign n9794 = \P1_P1_DataWidth_reg[1]/NET0131  & ~n9793 ;
  assign n9795 = ~n9792 & n9794 ;
  assign n9796 = ~\P1_P1_DataWidth_reg[1]/NET0131  & n9789 ;
  assign n9797 = n8282 & ~n9796 ;
  assign n9798 = ~n9795 & n9797 ;
  assign n9799 = n8287 & ~n9789 ;
  assign n9800 = n8592 & ~n9362 ;
  assign n9801 = ~n9787 & ~n9800 ;
  assign n9802 = n8350 & ~n9801 ;
  assign n9803 = \P1_P1_InstQueue_reg[4][6]/NET0131  & ~n8366 ;
  assign n9804 = ~n9802 & ~n9803 ;
  assign n9805 = ~n9799 & n9804 ;
  assign n9806 = ~n9798 & n9805 ;
  assign n9813 = n8568 & ~n9263 ;
  assign n9808 = ~n7940 & ~n8617 ;
  assign n9809 = \P1_P1_InstQueue_reg[5][4]/NET0131  & ~n8616 ;
  assign n9810 = ~n8592 & n9809 ;
  assign n9811 = ~n9808 & ~n9810 ;
  assign n9812 = ~n8568 & n9811 ;
  assign n9814 = ~n8544 & ~n9812 ;
  assign n9815 = ~n9813 & n9814 ;
  assign n9807 = n8544 & n9254 ;
  assign n9816 = \P1_P1_DataWidth_reg[1]/NET0131  & ~n9807 ;
  assign n9817 = ~n9815 & n9816 ;
  assign n9818 = ~\P1_P1_DataWidth_reg[1]/NET0131  & n9811 ;
  assign n9819 = n8282 & ~n9818 ;
  assign n9820 = ~n9817 & n9819 ;
  assign n9821 = n8287 & ~n9811 ;
  assign n9822 = n8616 & ~n9303 ;
  assign n9823 = ~n9809 & ~n9822 ;
  assign n9824 = n8350 & ~n9823 ;
  assign n9825 = \P1_P1_InstQueue_reg[5][4]/NET0131  & ~n8366 ;
  assign n9826 = ~n9824 & ~n9825 ;
  assign n9827 = ~n9821 & n9826 ;
  assign n9828 = ~n9820 & n9827 ;
  assign n9829 = n8568 & ~n9313 ;
  assign n9830 = n7906 & ~n8617 ;
  assign n9831 = \P1_P1_InstQueue_reg[5][6]/NET0131  & ~n8616 ;
  assign n9832 = ~n8592 & n9831 ;
  assign n9833 = ~n9830 & ~n9832 ;
  assign n9834 = ~n8568 & n9833 ;
  assign n9835 = ~n8544 & ~n9834 ;
  assign n9836 = ~n9829 & n9835 ;
  assign n9837 = n8544 & n9324 ;
  assign n9838 = \P1_P1_DataWidth_reg[1]/NET0131  & ~n9837 ;
  assign n9839 = ~n9836 & n9838 ;
  assign n9840 = ~\P1_P1_DataWidth_reg[1]/NET0131  & n9833 ;
  assign n9841 = n8282 & ~n9840 ;
  assign n9842 = ~n9839 & n9841 ;
  assign n9843 = n8287 & ~n9833 ;
  assign n9844 = n8616 & ~n9362 ;
  assign n9845 = ~n9831 & ~n9844 ;
  assign n9846 = n8350 & ~n9845 ;
  assign n9847 = \P1_P1_InstQueue_reg[5][6]/NET0131  & ~n8366 ;
  assign n9848 = ~n9846 & ~n9847 ;
  assign n9849 = ~n9843 & n9848 ;
  assign n9850 = ~n9842 & n9849 ;
  assign n9857 = n8592 & ~n9263 ;
  assign n9852 = ~n7940 & ~n8641 ;
  assign n9853 = \P1_P1_InstQueue_reg[6][4]/NET0131  & ~n8640 ;
  assign n9854 = ~n8616 & n9853 ;
  assign n9855 = ~n9852 & ~n9854 ;
  assign n9856 = ~n8592 & n9855 ;
  assign n9858 = ~n8568 & ~n9856 ;
  assign n9859 = ~n9857 & n9858 ;
  assign n9851 = n8568 & n9254 ;
  assign n9860 = \P1_P1_DataWidth_reg[1]/NET0131  & ~n9851 ;
  assign n9861 = ~n9859 & n9860 ;
  assign n9862 = ~\P1_P1_DataWidth_reg[1]/NET0131  & n9855 ;
  assign n9863 = n8282 & ~n9862 ;
  assign n9864 = ~n9861 & n9863 ;
  assign n9865 = n8287 & ~n9855 ;
  assign n9866 = n8640 & ~n9303 ;
  assign n9867 = ~n9853 & ~n9866 ;
  assign n9868 = n8350 & ~n9867 ;
  assign n9869 = \P1_P1_InstQueue_reg[6][4]/NET0131  & ~n8366 ;
  assign n9870 = ~n9868 & ~n9869 ;
  assign n9871 = ~n9865 & n9870 ;
  assign n9872 = ~n9864 & n9871 ;
  assign n9873 = n8592 & ~n9313 ;
  assign n9874 = n7906 & ~n8641 ;
  assign n9875 = \P1_P1_InstQueue_reg[6][6]/NET0131  & ~n8640 ;
  assign n9876 = ~n8616 & n9875 ;
  assign n9877 = ~n9874 & ~n9876 ;
  assign n9878 = ~n8592 & n9877 ;
  assign n9879 = ~n8568 & ~n9878 ;
  assign n9880 = ~n9873 & n9879 ;
  assign n9881 = n8568 & n9324 ;
  assign n9882 = \P1_P1_DataWidth_reg[1]/NET0131  & ~n9881 ;
  assign n9883 = ~n9880 & n9882 ;
  assign n9884 = ~\P1_P1_DataWidth_reg[1]/NET0131  & n9877 ;
  assign n9885 = n8282 & ~n9884 ;
  assign n9886 = ~n9883 & n9885 ;
  assign n9887 = n8287 & ~n9877 ;
  assign n9888 = n8640 & ~n9362 ;
  assign n9889 = ~n9875 & ~n9888 ;
  assign n9890 = n8350 & ~n9889 ;
  assign n9891 = \P1_P1_InstQueue_reg[6][6]/NET0131  & ~n8366 ;
  assign n9892 = ~n9890 & ~n9891 ;
  assign n9893 = ~n9887 & n9892 ;
  assign n9894 = ~n9886 & n9893 ;
  assign n9901 = n8616 & ~n9263 ;
  assign n9896 = ~n7940 & ~n8664 ;
  assign n9897 = \P1_P1_InstQueue_reg[7][4]/NET0131  & ~n8407 ;
  assign n9898 = ~n8640 & n9897 ;
  assign n9899 = ~n9896 & ~n9898 ;
  assign n9900 = ~n8616 & n9899 ;
  assign n9902 = ~n8592 & ~n9900 ;
  assign n9903 = ~n9901 & n9902 ;
  assign n9895 = n8592 & n9254 ;
  assign n9904 = \P1_P1_DataWidth_reg[1]/NET0131  & ~n9895 ;
  assign n9905 = ~n9903 & n9904 ;
  assign n9906 = ~\P1_P1_DataWidth_reg[1]/NET0131  & n9899 ;
  assign n9907 = n8282 & ~n9906 ;
  assign n9908 = ~n9905 & n9907 ;
  assign n9909 = n8287 & ~n9899 ;
  assign n9910 = n8407 & ~n9303 ;
  assign n9911 = ~n9897 & ~n9910 ;
  assign n9912 = n8350 & ~n9911 ;
  assign n9913 = \P1_P1_InstQueue_reg[7][4]/NET0131  & ~n8366 ;
  assign n9914 = ~n9912 & ~n9913 ;
  assign n9915 = ~n9909 & n9914 ;
  assign n9916 = ~n9908 & n9915 ;
  assign n9917 = n8616 & ~n9313 ;
  assign n9918 = n7906 & ~n8664 ;
  assign n9919 = \P1_P1_InstQueue_reg[7][6]/NET0131  & ~n8407 ;
  assign n9920 = ~n8640 & n9919 ;
  assign n9921 = ~n9918 & ~n9920 ;
  assign n9922 = ~n8616 & n9921 ;
  assign n9923 = ~n8592 & ~n9922 ;
  assign n9924 = ~n9917 & n9923 ;
  assign n9925 = n8592 & n9324 ;
  assign n9926 = \P1_P1_DataWidth_reg[1]/NET0131  & ~n9925 ;
  assign n9927 = ~n9924 & n9926 ;
  assign n9928 = ~\P1_P1_DataWidth_reg[1]/NET0131  & n9921 ;
  assign n9929 = n8282 & ~n9928 ;
  assign n9930 = ~n9927 & n9929 ;
  assign n9931 = n8287 & ~n9921 ;
  assign n9932 = n8407 & ~n9362 ;
  assign n9933 = ~n9919 & ~n9932 ;
  assign n9934 = n8350 & ~n9933 ;
  assign n9935 = \P1_P1_InstQueue_reg[7][6]/NET0131  & ~n8366 ;
  assign n9936 = ~n9934 & ~n9935 ;
  assign n9937 = ~n9931 & n9936 ;
  assign n9938 = ~n9930 & n9937 ;
  assign n9945 = n8640 & ~n9263 ;
  assign n9940 = ~n7940 & ~n8410 ;
  assign n9941 = \P1_P1_InstQueue_reg[8][4]/NET0131  & ~n8139 ;
  assign n9942 = ~n8407 & n9941 ;
  assign n9943 = ~n9940 & ~n9942 ;
  assign n9944 = ~n8640 & n9943 ;
  assign n9946 = ~n8616 & ~n9944 ;
  assign n9947 = ~n9945 & n9946 ;
  assign n9939 = n8616 & n9254 ;
  assign n9948 = \P1_P1_DataWidth_reg[1]/NET0131  & ~n9939 ;
  assign n9949 = ~n9947 & n9948 ;
  assign n9950 = ~\P1_P1_DataWidth_reg[1]/NET0131  & n9943 ;
  assign n9951 = n8282 & ~n9950 ;
  assign n9952 = ~n9949 & n9951 ;
  assign n9953 = n8287 & ~n9943 ;
  assign n9954 = n8139 & ~n9303 ;
  assign n9955 = ~n9941 & ~n9954 ;
  assign n9956 = n8350 & ~n9955 ;
  assign n9957 = \P1_P1_InstQueue_reg[8][4]/NET0131  & ~n8366 ;
  assign n9958 = ~n9956 & ~n9957 ;
  assign n9959 = ~n9953 & n9958 ;
  assign n9960 = ~n9952 & n9959 ;
  assign n9961 = n8640 & ~n9313 ;
  assign n9962 = n7906 & ~n8410 ;
  assign n9963 = \P1_P1_InstQueue_reg[8][6]/NET0131  & ~n8139 ;
  assign n9964 = ~n8407 & n9963 ;
  assign n9965 = ~n9962 & ~n9964 ;
  assign n9966 = ~n8640 & n9965 ;
  assign n9967 = ~n8616 & ~n9966 ;
  assign n9968 = ~n9961 & n9967 ;
  assign n9969 = n8616 & n9324 ;
  assign n9970 = \P1_P1_DataWidth_reg[1]/NET0131  & ~n9969 ;
  assign n9971 = ~n9968 & n9970 ;
  assign n9972 = ~\P1_P1_DataWidth_reg[1]/NET0131  & n9965 ;
  assign n9973 = n8282 & ~n9972 ;
  assign n9974 = ~n9971 & n9973 ;
  assign n9975 = n8287 & ~n9965 ;
  assign n9976 = n8139 & ~n9362 ;
  assign n9977 = ~n9963 & ~n9976 ;
  assign n9978 = n8350 & ~n9977 ;
  assign n9979 = \P1_P1_InstQueue_reg[8][6]/NET0131  & ~n8366 ;
  assign n9980 = ~n9978 & ~n9979 ;
  assign n9981 = ~n9975 & n9980 ;
  assign n9982 = ~n9974 & n9981 ;
  assign n9989 = n8407 & ~n9263 ;
  assign n9984 = ~n7940 & ~n8709 ;
  assign n9985 = \P1_P1_InstQueue_reg[9][4]/NET0131  & ~n4327 ;
  assign n9986 = ~n8139 & n9985 ;
  assign n9987 = ~n9984 & ~n9986 ;
  assign n9988 = ~n8407 & n9987 ;
  assign n9990 = ~n8640 & ~n9988 ;
  assign n9991 = ~n9989 & n9990 ;
  assign n9983 = n8640 & n9254 ;
  assign n9992 = \P1_P1_DataWidth_reg[1]/NET0131  & ~n9983 ;
  assign n9993 = ~n9991 & n9992 ;
  assign n9994 = ~\P1_P1_DataWidth_reg[1]/NET0131  & n9987 ;
  assign n9995 = n8282 & ~n9994 ;
  assign n9996 = ~n9993 & n9995 ;
  assign n9997 = n8287 & ~n9987 ;
  assign n9998 = n4327 & ~n9303 ;
  assign n9999 = ~n9985 & ~n9998 ;
  assign n10000 = n8350 & ~n9999 ;
  assign n10001 = \P1_P1_InstQueue_reg[9][4]/NET0131  & ~n8366 ;
  assign n10002 = ~n10000 & ~n10001 ;
  assign n10003 = ~n9997 & n10002 ;
  assign n10004 = ~n9996 & n10003 ;
  assign n10005 = n8407 & ~n9313 ;
  assign n10006 = n7906 & ~n8709 ;
  assign n10007 = \P1_P1_InstQueue_reg[9][6]/NET0131  & ~n4327 ;
  assign n10008 = ~n8139 & n10007 ;
  assign n10009 = ~n10006 & ~n10008 ;
  assign n10010 = ~n8407 & n10009 ;
  assign n10011 = ~n8640 & ~n10010 ;
  assign n10012 = ~n10005 & n10011 ;
  assign n10013 = n8640 & n9324 ;
  assign n10014 = \P1_P1_DataWidth_reg[1]/NET0131  & ~n10013 ;
  assign n10015 = ~n10012 & n10014 ;
  assign n10016 = ~\P1_P1_DataWidth_reg[1]/NET0131  & n10009 ;
  assign n10017 = n8282 & ~n10016 ;
  assign n10018 = ~n10015 & n10017 ;
  assign n10019 = n8287 & ~n10009 ;
  assign n10020 = n4327 & ~n9362 ;
  assign n10021 = ~n10007 & ~n10020 ;
  assign n10022 = n8350 & ~n10021 ;
  assign n10023 = \P1_P1_InstQueue_reg[9][6]/NET0131  & ~n8366 ;
  assign n10024 = ~n10022 & ~n10023 ;
  assign n10025 = ~n10019 & n10024 ;
  assign n10026 = ~n10018 & n10025 ;
  assign n10027 = n9235 & n9238 ;
  assign n10028 = n9241 & ~n10027 ;
  assign n10033 = \P1_P3_State2_reg[1]/NET0131  & \P1_P3_State2_reg[2]/NET0131  ;
  assign n10034 = n8741 & n10033 ;
  assign n10035 = n8733 & ~n10034 ;
  assign n10032 = n8732 & n8741 ;
  assign n10029 = ~\P1_P3_State2_reg[1]/NET0131  & ~\P1_P3_State2_reg[2]/NET0131  ;
  assign n10030 = \P1_P3_State2_reg[3]/NET0131  & n10029 ;
  assign n10031 = \P1_P3_State2_reg[0]/NET0131  & n10030 ;
  assign n10036 = ~\P1_P3_State2_reg[3]/NET0131  & n10033 ;
  assign n10037 = \P1_P3_State2_reg[0]/NET0131  & n10036 ;
  assign n10038 = ~\P1_P3_Flush_reg/NET0131  & \P1_P3_InstQueueRd_Addr_reg[2]/NET0131  ;
  assign n10039 = \P1_P3_InstQueueRd_Addr_reg[3]/NET0131  & ~n8744 ;
  assign n10040 = n10038 & n10039 ;
  assign n10041 = n10037 & ~n10040 ;
  assign n10042 = ~n10031 & ~n10041 ;
  assign n10043 = ~n10032 & n10042 ;
  assign n10044 = ~n10035 & n10043 ;
  assign n10045 = ~n10028 & n10044 ;
  assign n10046 = ~\P1_P3_State2_reg[0]/NET0131  & n10030 ;
  assign n10047 = ~n10037 & ~n10046 ;
  assign n10049 = ~n8207 & n8232 ;
  assign n10050 = ~n9252 & ~n10049 ;
  assign n10051 = n8139 & n10050 ;
  assign n10052 = ~n8069 & n8077 ;
  assign n10053 = ~n9261 & ~n10052 ;
  assign n10054 = n4327 & n10053 ;
  assign n10055 = ~n10051 & ~n10054 ;
  assign n10056 = \P1_P1_DataWidth_reg[1]/NET0131  & ~n10055 ;
  assign n10057 = \P1_P1_DataWidth_reg[1]/NET0131  & ~n8709 ;
  assign n10058 = ~n7913 & ~n8146 ;
  assign n10059 = \P1_P1_InstQueue_reg[11][3]/NET0131  & ~n8142 ;
  assign n10060 = ~n8145 & n10059 ;
  assign n10061 = ~n10058 & ~n10060 ;
  assign n10062 = ~n10057 & ~n10061 ;
  assign n10063 = ~n10056 & ~n10062 ;
  assign n10064 = n8282 & ~n10063 ;
  assign n10065 = n8287 & ~n10061 ;
  assign n10048 = \P1_P1_InstQueue_reg[11][3]/NET0131  & ~n8366 ;
  assign n10066 = \P1_P1_InstQueue_reg[14][3]/NET0131  & n8291 ;
  assign n10067 = \P1_P1_InstQueue_reg[4][3]/NET0131  & n8295 ;
  assign n10068 = \P1_P1_InstQueue_reg[8][3]/NET0131  & n8305 ;
  assign n10082 = ~n10067 & ~n10068 ;
  assign n10069 = \P1_P1_InstQueue_reg[11][3]/NET0131  & n8312 ;
  assign n10070 = \P1_P1_InstQueue_reg[3][3]/NET0131  & n8323 ;
  assign n10083 = ~n10069 & ~n10070 ;
  assign n10092 = n10082 & n10083 ;
  assign n10093 = ~n10066 & n10092 ;
  assign n10081 = \P1_P1_InstQueue_reg[13][3]/NET0131  & n8327 ;
  assign n10079 = \P1_P1_InstQueue_reg[2][3]/NET0131  & n8314 ;
  assign n10080 = \P1_P1_InstQueue_reg[5][3]/NET0131  & n8307 ;
  assign n10088 = ~n10079 & ~n10080 ;
  assign n10089 = ~n10081 & n10088 ;
  assign n10075 = \P1_P1_InstQueue_reg[6][3]/NET0131  & n8316 ;
  assign n10076 = \P1_P1_InstQueue_reg[15][3]/NET0131  & n8321 ;
  assign n10086 = ~n10075 & ~n10076 ;
  assign n10077 = \P1_P1_InstQueue_reg[7][3]/NET0131  & n8318 ;
  assign n10078 = \P1_P1_InstQueue_reg[0][3]/NET0131  & n8309 ;
  assign n10087 = ~n10077 & ~n10078 ;
  assign n10090 = n10086 & n10087 ;
  assign n10071 = \P1_P1_InstQueue_reg[12][3]/NET0131  & n8329 ;
  assign n10072 = \P1_P1_InstQueue_reg[10][3]/NET0131  & n8303 ;
  assign n10084 = ~n10071 & ~n10072 ;
  assign n10073 = \P1_P1_InstQueue_reg[1][3]/NET0131  & n8299 ;
  assign n10074 = \P1_P1_InstQueue_reg[9][3]/NET0131  & n8325 ;
  assign n10085 = ~n10073 & ~n10074 ;
  assign n10091 = n10084 & n10085 ;
  assign n10094 = n10090 & n10091 ;
  assign n10095 = n10089 & n10094 ;
  assign n10096 = n10093 & n10095 ;
  assign n10097 = n8142 & ~n10096 ;
  assign n10098 = ~n10059 & ~n10097 ;
  assign n10099 = n8350 & ~n10098 ;
  assign n10100 = ~n10048 & ~n10099 ;
  assign n10101 = ~n10065 & n10100 ;
  assign n10102 = ~n10064 & n10101 ;
  assign n10103 = ~\P2_P1_InstQueueWr_Addr_reg[0]/NET0131  & ~\P2_P1_InstQueueWr_Addr_reg[1]/NET0131  ;
  assign n10104 = ~\P2_P1_InstQueueWr_Addr_reg[2]/NET0131  & n10103 ;
  assign n10105 = \P2_P1_InstQueueWr_Addr_reg[3]/NET0131  & n10104 ;
  assign n10115 = ~\P2_P1_Address_reg[26]/NET0131  & ~\P2_P1_Address_reg[27]/NET0131  ;
  assign n10116 = ~\P2_P1_Address_reg[28]/NET0131  & ~\P2_P1_Address_reg[2]/NET0131  ;
  assign n10122 = n10115 & n10116 ;
  assign n10113 = ~\P2_P1_Address_reg[22]/NET0131  & ~\P2_P1_Address_reg[23]/NET0131  ;
  assign n10114 = ~\P2_P1_Address_reg[24]/NET0131  & ~\P2_P1_Address_reg[25]/NET0131  ;
  assign n10123 = n10113 & n10114 ;
  assign n10129 = n10122 & n10123 ;
  assign n10119 = ~\P2_P1_Address_reg[7]/NET0131  & ~\P2_P1_Address_reg[8]/NET0131  ;
  assign n10120 = ~\P2_P1_Address_reg[9]/NET0131  & n10119 ;
  assign n10117 = ~\P2_P1_Address_reg[3]/NET0131  & ~\P2_P1_Address_reg[4]/NET0131  ;
  assign n10118 = ~\P2_P1_Address_reg[5]/NET0131  & ~\P2_P1_Address_reg[6]/NET0131  ;
  assign n10121 = n10117 & n10118 ;
  assign n10130 = n10120 & n10121 ;
  assign n10131 = n10129 & n10130 ;
  assign n10106 = ~\P2_P1_Address_reg[0]/NET0131  & ~\P2_P1_Address_reg[10]/NET0131  ;
  assign n10107 = ~\P2_P1_Address_reg[11]/NET0131  & ~\P2_P1_Address_reg[12]/NET0131  ;
  assign n10108 = ~\P2_P1_Address_reg[13]/NET0131  & ~\P2_P1_Address_reg[14]/NET0131  ;
  assign n10126 = n10107 & n10108 ;
  assign n10127 = n10106 & n10126 ;
  assign n10111 = ~\P2_P1_Address_reg[19]/NET0131  & ~\P2_P1_Address_reg[1]/NET0131  ;
  assign n10112 = ~\P2_P1_Address_reg[20]/NET0131  & ~\P2_P1_Address_reg[21]/NET0131  ;
  assign n10124 = n10111 & n10112 ;
  assign n10109 = ~\P2_P1_Address_reg[15]/NET0131  & ~\P2_P1_Address_reg[16]/NET0131  ;
  assign n10110 = ~\P2_P1_Address_reg[17]/NET0131  & ~\P2_P1_Address_reg[18]/NET0131  ;
  assign n10125 = n10109 & n10110 ;
  assign n10128 = n10124 & n10125 ;
  assign n10132 = n10127 & n10128 ;
  assign n10133 = n10131 & n10132 ;
  assign n10134 = \P2_P1_Address_reg[29]/NET0131  & ~n10133 ;
  assign n10135 = \din[3]_pad  & ~sel_pad ;
  assign n10136 = \din[1]_pad  & ~sel_pad ;
  assign n10137 = n10135 & n10136 ;
  assign n10138 = ~n10135 & ~n10136 ;
  assign n10139 = ~n10137 & ~n10138 ;
  assign n10140 = \din[5]_pad  & ~sel_pad ;
  assign n10141 = \din[21]_pad  & n10140 ;
  assign n10142 = \din[21]_pad  & ~sel_pad ;
  assign n10143 = ~n10140 & ~n10142 ;
  assign n10144 = \din[23]_pad  & ~n10143 ;
  assign n10145 = ~n10141 & ~n10144 ;
  assign n10146 = n10139 & ~n10145 ;
  assign n10147 = ~n10139 & n10145 ;
  assign n10148 = \din[9]_pad  & ~sel_pad ;
  assign n10149 = \din[17]_pad  & n10148 ;
  assign n10150 = \din[17]_pad  & ~sel_pad ;
  assign n10151 = ~n10148 & ~n10150 ;
  assign n10152 = \din[19]_pad  & ~n10151 ;
  assign n10153 = ~n10149 & ~n10152 ;
  assign n10154 = ~n10147 & ~n10153 ;
  assign n10155 = ~n10146 & ~n10154 ;
  assign n10156 = \din[15]_pad  & ~sel_pad ;
  assign n10157 = \din[7]_pad  & ~sel_pad ;
  assign n10158 = ~n10156 & ~n10157 ;
  assign n10159 = n10156 & n10157 ;
  assign n10160 = ~n10135 & ~n10159 ;
  assign n10161 = ~n10158 & ~n10160 ;
  assign n10162 = \din[11]_pad  & ~sel_pad ;
  assign n10163 = n10136 & n10162 ;
  assign n10164 = ~n10161 & ~n10163 ;
  assign n10165 = n10161 & n10163 ;
  assign n10166 = \din[13]_pad  & ~sel_pad ;
  assign n10167 = ~n10165 & ~n10166 ;
  assign n10168 = ~n10164 & ~n10167 ;
  assign n10169 = ~n10155 & n10168 ;
  assign n10170 = n10155 & ~n10168 ;
  assign n10171 = ~n10169 & ~n10170 ;
  assign n10172 = ~n10158 & ~n10159 ;
  assign n10173 = ~n10150 & n10172 ;
  assign n10174 = n10150 & ~n10172 ;
  assign n10175 = ~n10173 & ~n10174 ;
  assign n10176 = \din[19]_pad  & ~sel_pad ;
  assign n10177 = n10148 & ~n10176 ;
  assign n10178 = ~n10148 & n10176 ;
  assign n10179 = ~n10177 & ~n10178 ;
  assign n10180 = n10142 & n10179 ;
  assign n10181 = ~n10142 & ~n10179 ;
  assign n10182 = ~n10180 & ~n10181 ;
  assign n10183 = ~n10175 & ~n10182 ;
  assign n10184 = n10175 & n10182 ;
  assign n10185 = \din[23]_pad  & ~sel_pad ;
  assign n10186 = ~n10140 & ~n10162 ;
  assign n10187 = n10140 & n10162 ;
  assign n10188 = ~n10186 & ~n10187 ;
  assign n10189 = ~n10185 & n10188 ;
  assign n10190 = n10185 & ~n10188 ;
  assign n10191 = ~n10189 & ~n10190 ;
  assign n10192 = ~n10184 & ~n10191 ;
  assign n10193 = ~n10183 & ~n10192 ;
  assign n10194 = n10171 & n10193 ;
  assign n10195 = ~n10171 & ~n10193 ;
  assign n10196 = ~n10194 & ~n10195 ;
  assign n10197 = \din[13]_pad  & n10137 ;
  assign n10198 = ~n10137 & ~n10166 ;
  assign n10199 = ~n10150 & ~n10159 ;
  assign n10200 = ~n10158 & ~n10199 ;
  assign n10201 = ~n10198 & n10200 ;
  assign n10202 = ~n10197 & ~n10201 ;
  assign n10203 = ~n10164 & ~n10165 ;
  assign n10204 = n10166 & ~n10203 ;
  assign n10205 = ~n10166 & n10203 ;
  assign n10206 = ~n10204 & ~n10205 ;
  assign n10207 = ~n10202 & ~n10206 ;
  assign n10208 = n10202 & n10206 ;
  assign n10209 = n10140 & n10142 ;
  assign n10210 = ~n10143 & ~n10209 ;
  assign n10211 = ~n10185 & n10210 ;
  assign n10212 = n10185 & ~n10210 ;
  assign n10213 = ~n10211 & ~n10212 ;
  assign n10214 = n10150 & n10179 ;
  assign n10215 = ~n10150 & ~n10179 ;
  assign n10216 = ~n10214 & ~n10215 ;
  assign n10217 = ~n10213 & ~n10216 ;
  assign n10218 = n10213 & n10216 ;
  assign n10219 = n10135 & ~n10157 ;
  assign n10220 = ~n10135 & n10157 ;
  assign n10221 = ~n10219 & ~n10220 ;
  assign n10222 = n10156 & n10221 ;
  assign n10223 = ~n10156 & ~n10221 ;
  assign n10224 = ~n10222 & ~n10223 ;
  assign n10225 = ~n10218 & ~n10224 ;
  assign n10226 = ~n10217 & ~n10225 ;
  assign n10227 = ~n10208 & ~n10226 ;
  assign n10228 = ~n10207 & ~n10227 ;
  assign n10229 = ~n10196 & ~n10228 ;
  assign n10230 = n10196 & n10228 ;
  assign n10231 = ~n10146 & ~n10147 ;
  assign n10232 = ~n10153 & n10231 ;
  assign n10233 = n10153 & ~n10231 ;
  assign n10234 = ~n10232 & ~n10233 ;
  assign n10235 = ~n10185 & ~n10187 ;
  assign n10236 = ~n10186 & ~n10235 ;
  assign n10237 = ~n10142 & ~n10176 ;
  assign n10238 = n10142 & n10176 ;
  assign n10239 = ~n10148 & ~n10238 ;
  assign n10240 = ~n10237 & ~n10239 ;
  assign n10241 = n10236 & n10240 ;
  assign n10242 = ~n10236 & ~n10240 ;
  assign n10243 = ~n10136 & ~n10162 ;
  assign n10244 = ~n10163 & ~n10243 ;
  assign n10245 = ~n10242 & n10244 ;
  assign n10246 = ~n10241 & ~n10245 ;
  assign n10247 = ~n10234 & n10246 ;
  assign n10248 = n10234 & ~n10246 ;
  assign n10249 = ~n10183 & ~n10184 ;
  assign n10250 = ~n10191 & n10249 ;
  assign n10251 = n10191 & ~n10249 ;
  assign n10252 = ~n10250 & ~n10251 ;
  assign n10253 = ~n10248 & ~n10252 ;
  assign n10254 = ~n10247 & ~n10253 ;
  assign n10255 = ~n10230 & n10254 ;
  assign n10256 = ~n10229 & ~n10255 ;
  assign n10257 = \din[25]_pad  & ~sel_pad ;
  assign n10258 = ~n10185 & ~n10257 ;
  assign n10259 = n10185 & n10257 ;
  assign n10260 = ~n10258 & ~n10259 ;
  assign n10261 = ~n10136 & n10260 ;
  assign n10262 = n10136 & ~n10260 ;
  assign n10263 = ~n10261 & ~n10262 ;
  assign n10264 = n10221 & n10263 ;
  assign n10265 = ~n10221 & ~n10263 ;
  assign n10266 = ~n10197 & ~n10198 ;
  assign n10267 = ~n10140 & n10266 ;
  assign n10268 = n10140 & ~n10266 ;
  assign n10269 = ~n10267 & ~n10268 ;
  assign n10270 = ~n10265 & n10269 ;
  assign n10271 = ~n10264 & ~n10270 ;
  assign n10272 = \din[27]_pad  & ~sel_pad ;
  assign n10273 = n10166 & n10272 ;
  assign n10274 = ~n10166 & ~n10272 ;
  assign n10275 = ~n10273 & ~n10274 ;
  assign n10276 = ~n10257 & n10275 ;
  assign n10277 = n10257 & ~n10275 ;
  assign n10278 = ~n10276 & ~n10277 ;
  assign n10279 = ~n10175 & ~n10278 ;
  assign n10280 = n10175 & n10278 ;
  assign n10281 = ~n10279 & ~n10280 ;
  assign n10282 = n10191 & n10281 ;
  assign n10283 = ~n10191 & ~n10281 ;
  assign n10284 = ~n10282 & ~n10283 ;
  assign n10285 = n10271 & ~n10284 ;
  assign n10286 = ~n10271 & n10284 ;
  assign n10287 = ~n10285 & ~n10286 ;
  assign n10288 = ~n10140 & ~n10166 ;
  assign n10289 = \din[13]_pad  & n10140 ;
  assign n10290 = ~n10137 & ~n10289 ;
  assign n10291 = ~n10288 & ~n10290 ;
  assign n10292 = ~n10182 & n10291 ;
  assign n10293 = n10182 & ~n10291 ;
  assign n10294 = ~n10292 & ~n10293 ;
  assign n10295 = n10135 & n10157 ;
  assign n10296 = n10139 & ~n10272 ;
  assign n10297 = ~n10139 & n10272 ;
  assign n10298 = ~n10296 & ~n10297 ;
  assign n10299 = n10295 & ~n10298 ;
  assign n10300 = ~n10295 & n10298 ;
  assign n10301 = ~n10299 & ~n10300 ;
  assign n10302 = ~n10294 & n10301 ;
  assign n10303 = n10294 & ~n10301 ;
  assign n10304 = ~n10302 & ~n10303 ;
  assign n10305 = n10287 & n10304 ;
  assign n10306 = ~n10287 & ~n10304 ;
  assign n10307 = ~n10305 & ~n10306 ;
  assign n10308 = n10256 & n10307 ;
  assign n10309 = ~n10256 & ~n10307 ;
  assign n10310 = ~n10308 & ~n10309 ;
  assign n10311 = ~n10170 & ~n10193 ;
  assign n10312 = ~n10169 & ~n10311 ;
  assign n10313 = ~n10264 & ~n10265 ;
  assign n10314 = n10269 & n10313 ;
  assign n10315 = ~n10269 & ~n10313 ;
  assign n10316 = ~n10314 & ~n10315 ;
  assign n10317 = ~n10200 & ~n10240 ;
  assign n10318 = n10200 & n10240 ;
  assign n10319 = ~n10317 & ~n10318 ;
  assign n10320 = ~n10257 & n10319 ;
  assign n10321 = n10257 & ~n10319 ;
  assign n10322 = ~n10320 & ~n10321 ;
  assign n10323 = n10316 & n10322 ;
  assign n10324 = ~n10316 & ~n10322 ;
  assign n10325 = ~n10237 & ~n10238 ;
  assign n10326 = ~n10162 & n10325 ;
  assign n10327 = n10162 & ~n10325 ;
  assign n10328 = ~n10326 & ~n10327 ;
  assign n10329 = ~n10236 & n10328 ;
  assign n10330 = n10236 & ~n10328 ;
  assign n10331 = ~n10329 & ~n10330 ;
  assign n10332 = n10148 & n10150 ;
  assign n10333 = ~n10151 & ~n10332 ;
  assign n10334 = ~n10156 & n10333 ;
  assign n10335 = n10156 & ~n10333 ;
  assign n10336 = ~n10334 & ~n10335 ;
  assign n10337 = n10331 & n10336 ;
  assign n10338 = ~n10331 & ~n10336 ;
  assign n10339 = ~n10337 & ~n10338 ;
  assign n10340 = ~n10324 & n10339 ;
  assign n10341 = ~n10323 & ~n10340 ;
  assign n10342 = n10312 & ~n10341 ;
  assign n10343 = ~n10312 & n10341 ;
  assign n10344 = ~n10342 & ~n10343 ;
  assign n10345 = ~n10257 & ~n10318 ;
  assign n10346 = ~n10317 & ~n10345 ;
  assign n10347 = ~n10162 & ~n10238 ;
  assign n10348 = ~n10237 & ~n10347 ;
  assign n10349 = ~n10136 & ~n10259 ;
  assign n10350 = ~n10258 & ~n10349 ;
  assign n10351 = ~n10149 & ~n10156 ;
  assign n10352 = ~n10151 & ~n10351 ;
  assign n10353 = n10350 & n10352 ;
  assign n10354 = ~n10350 & ~n10352 ;
  assign n10355 = ~n10353 & ~n10354 ;
  assign n10356 = n10348 & ~n10355 ;
  assign n10357 = ~n10348 & n10355 ;
  assign n10358 = ~n10356 & ~n10357 ;
  assign n10359 = ~n10346 & n10358 ;
  assign n10360 = n10346 & ~n10358 ;
  assign n10361 = ~n10359 & ~n10360 ;
  assign n10362 = ~n10329 & ~n10336 ;
  assign n10363 = ~n10330 & ~n10362 ;
  assign n10364 = n10361 & ~n10363 ;
  assign n10365 = ~n10361 & n10363 ;
  assign n10366 = ~n10364 & ~n10365 ;
  assign n10367 = n10344 & ~n10366 ;
  assign n10368 = ~n10344 & n10366 ;
  assign n10369 = ~n10367 & ~n10368 ;
  assign n10370 = n10310 & ~n10369 ;
  assign n10371 = ~n10310 & n10369 ;
  assign n10372 = ~n10370 & ~n10371 ;
  assign n10373 = ~n10241 & ~n10242 ;
  assign n10374 = ~n10244 & n10373 ;
  assign n10375 = n10244 & ~n10373 ;
  assign n10376 = ~n10374 & ~n10375 ;
  assign n10377 = ~n10182 & n10352 ;
  assign n10378 = n10182 & ~n10352 ;
  assign n10379 = ~n10191 & ~n10378 ;
  assign n10380 = ~n10377 & ~n10379 ;
  assign n10381 = n10376 & n10380 ;
  assign n10382 = ~n10376 & ~n10380 ;
  assign n10383 = ~n10217 & ~n10218 ;
  assign n10384 = ~n10224 & n10383 ;
  assign n10385 = n10224 & ~n10383 ;
  assign n10386 = ~n10384 & ~n10385 ;
  assign n10387 = ~n10382 & ~n10386 ;
  assign n10388 = ~n10381 & ~n10387 ;
  assign n10389 = ~n10136 & ~n10238 ;
  assign n10390 = ~n10237 & ~n10389 ;
  assign n10391 = ~n10295 & ~n10390 ;
  assign n10392 = n10295 & n10390 ;
  assign n10393 = ~n10162 & ~n10166 ;
  assign n10394 = ~n10186 & ~n10288 ;
  assign n10395 = ~n10393 & n10394 ;
  assign n10396 = ~n10392 & ~n10395 ;
  assign n10397 = ~n10391 & ~n10396 ;
  assign n10398 = ~n10200 & n10266 ;
  assign n10399 = n10200 & ~n10266 ;
  assign n10400 = ~n10398 & ~n10399 ;
  assign n10401 = ~n10397 & n10400 ;
  assign n10402 = n10397 & ~n10400 ;
  assign n10403 = ~n10139 & ~n10166 ;
  assign n10404 = n10139 & n10166 ;
  assign n10405 = ~n10185 & ~n10404 ;
  assign n10406 = ~n10403 & ~n10405 ;
  assign n10407 = ~n10402 & ~n10406 ;
  assign n10408 = ~n10401 & ~n10407 ;
  assign n10409 = ~n10388 & ~n10408 ;
  assign n10410 = n10388 & n10408 ;
  assign n10411 = ~n10207 & ~n10208 ;
  assign n10412 = ~n10226 & n10411 ;
  assign n10413 = n10226 & ~n10411 ;
  assign n10414 = ~n10412 & ~n10413 ;
  assign n10415 = ~n10410 & ~n10414 ;
  assign n10416 = ~n10409 & ~n10415 ;
  assign n10417 = ~n10323 & ~n10324 ;
  assign n10418 = n10339 & n10417 ;
  assign n10419 = ~n10339 & ~n10417 ;
  assign n10420 = ~n10418 & ~n10419 ;
  assign n10421 = n10416 & ~n10420 ;
  assign n10422 = ~n10416 & n10420 ;
  assign n10423 = ~n10229 & ~n10230 ;
  assign n10424 = ~n10254 & n10423 ;
  assign n10425 = n10254 & ~n10423 ;
  assign n10426 = ~n10424 & ~n10425 ;
  assign n10427 = ~n10422 & ~n10426 ;
  assign n10428 = ~n10421 & ~n10427 ;
  assign n10429 = ~n10372 & n10428 ;
  assign n10430 = ~n10359 & ~n10363 ;
  assign n10431 = ~n10360 & ~n10430 ;
  assign n10432 = ~n10136 & n10325 ;
  assign n10433 = n10136 & ~n10325 ;
  assign n10434 = ~n10432 & ~n10433 ;
  assign n10435 = n10336 & n10434 ;
  assign n10436 = ~n10336 & ~n10434 ;
  assign n10437 = ~n10435 & ~n10436 ;
  assign n10438 = ~n10140 & n10275 ;
  assign n10439 = n10140 & ~n10275 ;
  assign n10440 = ~n10438 & ~n10439 ;
  assign n10441 = ~n10437 & n10440 ;
  assign n10442 = n10437 & ~n10440 ;
  assign n10443 = ~n10441 & ~n10442 ;
  assign n10444 = n10431 & ~n10443 ;
  assign n10445 = ~n10431 & n10443 ;
  assign n10446 = ~n10444 & ~n10445 ;
  assign n10447 = ~n10293 & n10301 ;
  assign n10448 = ~n10292 & ~n10447 ;
  assign n10449 = n10446 & n10448 ;
  assign n10450 = ~n10446 & ~n10448 ;
  assign n10451 = ~n10449 & ~n10450 ;
  assign n10452 = ~n10342 & n10366 ;
  assign n10453 = ~n10343 & ~n10452 ;
  assign n10454 = n10451 & n10453 ;
  assign n10455 = ~n10451 & ~n10453 ;
  assign n10456 = ~n10454 & ~n10455 ;
  assign n10457 = ~n10286 & ~n10304 ;
  assign n10458 = ~n10285 & ~n10457 ;
  assign n10459 = ~\din[13]_pad  & ~\din[27]_pad  ;
  assign n10460 = n10257 & ~n10459 ;
  assign n10461 = ~n10273 & ~n10460 ;
  assign n10462 = ~n10221 & ~n10461 ;
  assign n10463 = n10221 & n10461 ;
  assign n10464 = ~n10462 & ~n10463 ;
  assign n10465 = n10236 & n10464 ;
  assign n10466 = ~n10236 & ~n10464 ;
  assign n10467 = ~n10465 & ~n10466 ;
  assign n10468 = ~n10191 & ~n10280 ;
  assign n10469 = ~n10279 & ~n10468 ;
  assign n10470 = n10467 & ~n10469 ;
  assign n10471 = ~n10467 & n10469 ;
  assign n10472 = ~n10470 & ~n10471 ;
  assign n10473 = n10137 & ~n10319 ;
  assign n10474 = ~n10137 & n10319 ;
  assign n10475 = ~n10473 & ~n10474 ;
  assign n10476 = ~n10472 & n10475 ;
  assign n10477 = n10472 & ~n10475 ;
  assign n10478 = ~n10476 & ~n10477 ;
  assign n10479 = ~n10458 & n10478 ;
  assign n10480 = n10458 & ~n10478 ;
  assign n10481 = ~n10479 & ~n10480 ;
  assign n10482 = ~n10136 & n10157 ;
  assign n10483 = ~n10272 & ~n10482 ;
  assign n10484 = ~n10139 & ~n10295 ;
  assign n10485 = ~n10483 & ~n10484 ;
  assign n10486 = ~n10162 & n10260 ;
  assign n10487 = n10162 & ~n10260 ;
  assign n10488 = ~n10486 & ~n10487 ;
  assign n10489 = n10485 & ~n10488 ;
  assign n10490 = ~n10485 & n10488 ;
  assign n10491 = ~n10489 & ~n10490 ;
  assign n10492 = ~n10348 & ~n10353 ;
  assign n10493 = ~n10354 & ~n10492 ;
  assign n10494 = n10491 & ~n10493 ;
  assign n10495 = ~n10491 & n10493 ;
  assign n10496 = ~n10494 & ~n10495 ;
  assign n10497 = n10481 & ~n10496 ;
  assign n10498 = ~n10481 & n10496 ;
  assign n10499 = ~n10497 & ~n10498 ;
  assign n10500 = n10456 & ~n10499 ;
  assign n10501 = ~n10456 & n10499 ;
  assign n10502 = ~n10500 & ~n10501 ;
  assign n10503 = ~n10308 & ~n10369 ;
  assign n10504 = ~n10309 & ~n10503 ;
  assign n10505 = n10502 & n10504 ;
  assign n10506 = ~n10429 & ~n10505 ;
  assign n10507 = ~n10445 & n10448 ;
  assign n10508 = ~n10444 & ~n10507 ;
  assign n10509 = ~n10480 & ~n10496 ;
  assign n10510 = ~n10479 & ~n10509 ;
  assign n10511 = n10508 & ~n10510 ;
  assign n10512 = ~n10508 & n10510 ;
  assign n10513 = ~n10162 & ~n10259 ;
  assign n10514 = ~n10258 & ~n10513 ;
  assign n10515 = n10272 & ~n10288 ;
  assign n10516 = ~n10289 & ~n10515 ;
  assign n10517 = ~n10514 & n10516 ;
  assign n10518 = n10514 & ~n10516 ;
  assign n10519 = ~n10517 & ~n10518 ;
  assign n10520 = \din[29]_pad  & ~sel_pad ;
  assign n10521 = n10172 & ~n10520 ;
  assign n10522 = ~n10172 & n10520 ;
  assign n10523 = ~n10521 & ~n10522 ;
  assign n10524 = n10519 & n10523 ;
  assign n10525 = ~n10519 & ~n10523 ;
  assign n10526 = ~n10524 & ~n10525 ;
  assign n10527 = n10236 & ~n10463 ;
  assign n10528 = ~n10462 & ~n10527 ;
  assign n10529 = n10526 & n10528 ;
  assign n10530 = ~n10526 & ~n10528 ;
  assign n10531 = ~n10529 & ~n10530 ;
  assign n10532 = ~n10391 & ~n10392 ;
  assign n10533 = n10352 & ~n10532 ;
  assign n10534 = ~n10352 & n10532 ;
  assign n10535 = ~n10533 & ~n10534 ;
  assign n10536 = n10531 & ~n10535 ;
  assign n10537 = ~n10531 & n10535 ;
  assign n10538 = ~n10536 & ~n10537 ;
  assign n10539 = ~n10137 & ~n10240 ;
  assign n10540 = n10137 & n10240 ;
  assign n10541 = ~n10200 & ~n10540 ;
  assign n10542 = ~n10539 & ~n10541 ;
  assign n10543 = n10298 & n10520 ;
  assign n10544 = ~n10298 & ~n10520 ;
  assign n10545 = ~n10543 & ~n10544 ;
  assign n10546 = ~n10542 & n10545 ;
  assign n10547 = n10542 & ~n10545 ;
  assign n10548 = ~n10546 & ~n10547 ;
  assign n10549 = ~n10435 & ~n10440 ;
  assign n10550 = ~n10436 & ~n10549 ;
  assign n10551 = n10548 & ~n10550 ;
  assign n10552 = ~n10548 & n10550 ;
  assign n10553 = ~n10551 & ~n10552 ;
  assign n10554 = ~n10538 & ~n10553 ;
  assign n10555 = n10538 & n10553 ;
  assign n10556 = ~n10554 & ~n10555 ;
  assign n10557 = ~n10489 & ~n10493 ;
  assign n10558 = ~n10490 & ~n10557 ;
  assign n10559 = ~n10166 & n10260 ;
  assign n10560 = n10166 & ~n10260 ;
  assign n10561 = ~n10559 & ~n10560 ;
  assign n10562 = n10216 & n10561 ;
  assign n10563 = ~n10216 & ~n10561 ;
  assign n10564 = ~n10562 & ~n10563 ;
  assign n10565 = ~n10142 & n10188 ;
  assign n10566 = n10142 & ~n10188 ;
  assign n10567 = ~n10565 & ~n10566 ;
  assign n10568 = ~n10564 & n10567 ;
  assign n10569 = n10564 & ~n10567 ;
  assign n10570 = ~n10568 & ~n10569 ;
  assign n10571 = n10558 & n10570 ;
  assign n10572 = ~n10558 & ~n10570 ;
  assign n10573 = ~n10571 & ~n10572 ;
  assign n10574 = ~n10470 & n10475 ;
  assign n10575 = ~n10471 & ~n10574 ;
  assign n10576 = n10573 & ~n10575 ;
  assign n10577 = ~n10573 & n10575 ;
  assign n10578 = ~n10576 & ~n10577 ;
  assign n10579 = n10556 & ~n10578 ;
  assign n10580 = ~n10556 & n10578 ;
  assign n10581 = ~n10579 & ~n10580 ;
  assign n10582 = ~n10512 & n10581 ;
  assign n10583 = ~n10511 & ~n10582 ;
  assign n10584 = ~n10555 & n10578 ;
  assign n10585 = ~n10554 & ~n10584 ;
  assign n10586 = ~n10562 & ~n10567 ;
  assign n10587 = ~n10563 & ~n10586 ;
  assign n10588 = n10139 & ~n10191 ;
  assign n10589 = ~n10139 & n10191 ;
  assign n10590 = ~n10588 & ~n10589 ;
  assign n10591 = ~n10278 & n10590 ;
  assign n10592 = n10278 & ~n10590 ;
  assign n10593 = ~n10591 & ~n10592 ;
  assign n10594 = n10587 & ~n10593 ;
  assign n10595 = ~n10587 & n10593 ;
  assign n10596 = ~n10594 & ~n10595 ;
  assign n10597 = ~n10517 & ~n10523 ;
  assign n10598 = ~n10518 & ~n10597 ;
  assign n10599 = n10596 & ~n10598 ;
  assign n10600 = ~n10596 & n10598 ;
  assign n10601 = ~n10599 & ~n10600 ;
  assign n10602 = ~n10159 & ~n10520 ;
  assign n10603 = ~n10158 & ~n10602 ;
  assign n10604 = ~n10137 & ~n10520 ;
  assign n10605 = \din[29]_pad  & n10137 ;
  assign n10606 = ~n10604 & ~n10605 ;
  assign n10607 = n10603 & ~n10606 ;
  assign n10608 = ~n10603 & n10606 ;
  assign n10609 = ~n10607 & ~n10608 ;
  assign n10610 = ~n10352 & ~n10392 ;
  assign n10611 = ~n10391 & ~n10610 ;
  assign n10612 = n10609 & ~n10611 ;
  assign n10613 = ~n10609 & n10611 ;
  assign n10614 = ~n10612 & ~n10613 ;
  assign n10615 = ~n10166 & ~n10259 ;
  assign n10616 = ~n10258 & ~n10615 ;
  assign n10617 = ~n10153 & n10616 ;
  assign n10618 = n10153 & ~n10616 ;
  assign n10619 = ~n10617 & ~n10618 ;
  assign n10620 = ~n10141 & ~n10162 ;
  assign n10621 = ~n10143 & ~n10620 ;
  assign n10622 = n10619 & ~n10621 ;
  assign n10623 = ~n10619 & n10621 ;
  assign n10624 = ~n10622 & ~n10623 ;
  assign n10625 = n10614 & ~n10624 ;
  assign n10626 = ~n10614 & n10624 ;
  assign n10627 = ~n10625 & ~n10626 ;
  assign n10628 = n10601 & n10627 ;
  assign n10629 = ~n10601 & ~n10627 ;
  assign n10630 = ~n10628 & ~n10629 ;
  assign n10631 = ~n10571 & ~n10575 ;
  assign n10632 = ~n10572 & ~n10631 ;
  assign n10633 = n10630 & ~n10632 ;
  assign n10634 = ~n10630 & n10632 ;
  assign n10635 = ~n10633 & ~n10634 ;
  assign n10636 = n10585 & ~n10635 ;
  assign n10637 = ~n10585 & n10635 ;
  assign n10638 = ~n10636 & ~n10637 ;
  assign n10639 = ~n10546 & ~n10550 ;
  assign n10640 = ~n10547 & ~n10639 ;
  assign n10641 = ~n10272 & ~n10520 ;
  assign n10642 = n10139 & ~n10641 ;
  assign n10643 = \din[27]_pad  & n10520 ;
  assign n10644 = ~n10642 & ~n10643 ;
  assign n10645 = n10249 & ~n10644 ;
  assign n10646 = ~n10249 & n10644 ;
  assign n10647 = ~n10645 & ~n10646 ;
  assign n10648 = n10640 & ~n10647 ;
  assign n10649 = ~n10640 & n10647 ;
  assign n10650 = ~n10648 & ~n10649 ;
  assign n10651 = ~n10529 & ~n10535 ;
  assign n10652 = ~n10530 & ~n10651 ;
  assign n10653 = n10650 & ~n10652 ;
  assign n10654 = ~n10650 & n10652 ;
  assign n10655 = ~n10653 & ~n10654 ;
  assign n10656 = n10638 & ~n10655 ;
  assign n10657 = ~n10638 & n10655 ;
  assign n10658 = ~n10656 & ~n10657 ;
  assign n10659 = n10583 & n10658 ;
  assign n10660 = ~n10454 & n10499 ;
  assign n10661 = ~n10455 & ~n10660 ;
  assign n10662 = ~n10511 & ~n10512 ;
  assign n10663 = n10581 & n10662 ;
  assign n10664 = ~n10581 & ~n10662 ;
  assign n10665 = ~n10663 & ~n10664 ;
  assign n10666 = n10661 & ~n10665 ;
  assign n10667 = ~n10659 & ~n10666 ;
  assign n10668 = n10506 & n10667 ;
  assign n10669 = ~n10421 & ~n10422 ;
  assign n10670 = ~n10426 & n10669 ;
  assign n10671 = n10426 & ~n10669 ;
  assign n10672 = ~n10670 & ~n10671 ;
  assign n10673 = ~n10403 & ~n10404 ;
  assign n10674 = ~n10185 & n10673 ;
  assign n10675 = n10185 & ~n10673 ;
  assign n10676 = ~n10674 & ~n10675 ;
  assign n10677 = ~n10175 & ~n10676 ;
  assign n10678 = n10175 & n10676 ;
  assign n10679 = ~n10540 & ~n10621 ;
  assign n10680 = ~n10539 & ~n10679 ;
  assign n10681 = ~n10678 & n10680 ;
  assign n10682 = ~n10677 & ~n10681 ;
  assign n10683 = ~n10401 & ~n10402 ;
  assign n10684 = ~n10406 & n10683 ;
  assign n10685 = n10406 & ~n10683 ;
  assign n10686 = ~n10684 & ~n10685 ;
  assign n10687 = ~n10682 & ~n10686 ;
  assign n10688 = n10682 & n10686 ;
  assign n10689 = n10200 & ~n10435 ;
  assign n10690 = ~n10436 & ~n10689 ;
  assign n10691 = ~n10395 & n10532 ;
  assign n10692 = n10395 & ~n10532 ;
  assign n10693 = ~n10691 & ~n10692 ;
  assign n10694 = ~n10690 & ~n10693 ;
  assign n10695 = n10690 & n10693 ;
  assign n10696 = ~n10377 & ~n10378 ;
  assign n10697 = ~n10191 & n10696 ;
  assign n10698 = n10191 & ~n10696 ;
  assign n10699 = ~n10697 & ~n10698 ;
  assign n10700 = ~n10695 & n10699 ;
  assign n10701 = ~n10694 & ~n10700 ;
  assign n10702 = ~n10688 & ~n10701 ;
  assign n10703 = ~n10687 & ~n10702 ;
  assign n10704 = ~n10247 & ~n10248 ;
  assign n10705 = ~n10252 & n10704 ;
  assign n10706 = n10252 & ~n10704 ;
  assign n10707 = ~n10705 & ~n10706 ;
  assign n10708 = ~n10703 & ~n10707 ;
  assign n10709 = n10703 & n10707 ;
  assign n10710 = ~n10409 & ~n10410 ;
  assign n10711 = ~n10414 & n10710 ;
  assign n10712 = n10414 & ~n10710 ;
  assign n10713 = ~n10711 & ~n10712 ;
  assign n10714 = ~n10709 & ~n10713 ;
  assign n10715 = ~n10708 & ~n10714 ;
  assign n10716 = ~n10672 & n10715 ;
  assign n10717 = ~n10677 & ~n10678 ;
  assign n10718 = ~n10680 & n10717 ;
  assign n10719 = n10680 & ~n10717 ;
  assign n10720 = ~n10718 & ~n10719 ;
  assign n10721 = ~n10166 & n10188 ;
  assign n10722 = n10166 & ~n10188 ;
  assign n10723 = ~n10721 & ~n10722 ;
  assign n10724 = ~n10221 & ~n10723 ;
  assign n10725 = n10221 & n10723 ;
  assign n10726 = ~n10150 & ~n10156 ;
  assign n10727 = n10150 & n10156 ;
  assign n10728 = ~n10135 & ~n10727 ;
  assign n10729 = ~n10726 & ~n10728 ;
  assign n10730 = ~n10404 & ~n10729 ;
  assign n10731 = ~n10403 & ~n10730 ;
  assign n10732 = ~n10725 & n10731 ;
  assign n10733 = ~n10724 & ~n10732 ;
  assign n10734 = ~n10720 & ~n10733 ;
  assign n10735 = n10720 & n10733 ;
  assign n10736 = ~n10694 & ~n10695 ;
  assign n10737 = ~n10699 & n10736 ;
  assign n10738 = n10699 & ~n10736 ;
  assign n10739 = ~n10737 & ~n10738 ;
  assign n10740 = ~n10735 & ~n10739 ;
  assign n10741 = ~n10734 & ~n10740 ;
  assign n10742 = ~n10687 & ~n10688 ;
  assign n10743 = ~n10701 & n10742 ;
  assign n10744 = n10701 & ~n10742 ;
  assign n10745 = ~n10743 & ~n10744 ;
  assign n10746 = n10741 & ~n10745 ;
  assign n10747 = ~n10741 & n10745 ;
  assign n10748 = ~n10381 & ~n10382 ;
  assign n10749 = ~n10386 & n10748 ;
  assign n10750 = n10386 & ~n10748 ;
  assign n10751 = ~n10749 & ~n10750 ;
  assign n10752 = ~n10747 & n10751 ;
  assign n10753 = ~n10746 & ~n10752 ;
  assign n10754 = ~n10708 & ~n10709 ;
  assign n10755 = ~n10713 & n10754 ;
  assign n10756 = n10713 & ~n10754 ;
  assign n10757 = ~n10755 & ~n10756 ;
  assign n10758 = ~n10753 & ~n10757 ;
  assign n10759 = ~n10716 & ~n10758 ;
  assign n10760 = ~n10724 & ~n10725 ;
  assign n10761 = ~n10731 & n10760 ;
  assign n10762 = n10731 & ~n10760 ;
  assign n10763 = ~n10761 & ~n10762 ;
  assign n10764 = ~n10200 & n10437 ;
  assign n10765 = n10200 & ~n10437 ;
  assign n10766 = ~n10764 & ~n10765 ;
  assign n10767 = ~n10763 & ~n10766 ;
  assign n10768 = n10763 & n10766 ;
  assign n10769 = ~n10176 & ~n10200 ;
  assign n10770 = n10176 & n10200 ;
  assign n10771 = ~n10395 & ~n10770 ;
  assign n10772 = ~n10769 & ~n10771 ;
  assign n10773 = n10673 & ~n10729 ;
  assign n10774 = ~n10673 & n10729 ;
  assign n10775 = ~n10773 & ~n10774 ;
  assign n10776 = n10772 & ~n10775 ;
  assign n10777 = ~n10772 & n10775 ;
  assign n10778 = n10136 & n10157 ;
  assign n10779 = ~n10140 & ~n10148 ;
  assign n10780 = n10140 & n10148 ;
  assign n10781 = ~n10176 & ~n10780 ;
  assign n10782 = ~n10779 & ~n10781 ;
  assign n10783 = ~n10778 & ~n10782 ;
  assign n10784 = n10778 & n10782 ;
  assign n10785 = ~n10783 & ~n10784 ;
  assign n10786 = n10567 & n10785 ;
  assign n10787 = ~n10567 & ~n10785 ;
  assign n10788 = ~n10786 & ~n10787 ;
  assign n10789 = ~n10777 & ~n10788 ;
  assign n10790 = ~n10776 & ~n10789 ;
  assign n10791 = ~n10768 & ~n10790 ;
  assign n10792 = ~n10767 & ~n10791 ;
  assign n10793 = ~n10567 & ~n10783 ;
  assign n10794 = ~n10784 & ~n10793 ;
  assign n10795 = ~n10539 & ~n10540 ;
  assign n10796 = ~n10621 & n10795 ;
  assign n10797 = n10621 & ~n10795 ;
  assign n10798 = ~n10796 & ~n10797 ;
  assign n10799 = ~n10794 & ~n10798 ;
  assign n10800 = n10794 & n10798 ;
  assign n10801 = n10162 & n10166 ;
  assign n10802 = ~n10137 & ~n10801 ;
  assign n10803 = ~n10393 & ~n10802 ;
  assign n10804 = ~n10183 & ~n10803 ;
  assign n10805 = ~n10184 & ~n10804 ;
  assign n10806 = ~n10800 & n10805 ;
  assign n10807 = ~n10799 & ~n10806 ;
  assign n10808 = ~n10792 & ~n10807 ;
  assign n10809 = n10792 & n10807 ;
  assign n10810 = ~n10734 & ~n10735 ;
  assign n10811 = ~n10739 & n10810 ;
  assign n10812 = n10739 & ~n10810 ;
  assign n10813 = ~n10811 & ~n10812 ;
  assign n10814 = ~n10809 & n10813 ;
  assign n10815 = ~n10808 & ~n10814 ;
  assign n10816 = ~n10746 & ~n10747 ;
  assign n10817 = n10751 & n10816 ;
  assign n10818 = ~n10751 & ~n10816 ;
  assign n10819 = ~n10817 & ~n10818 ;
  assign n10820 = ~n10815 & ~n10819 ;
  assign n10821 = n10815 & n10819 ;
  assign n10822 = ~n10799 & ~n10800 ;
  assign n10823 = n10805 & n10822 ;
  assign n10824 = ~n10805 & ~n10822 ;
  assign n10825 = ~n10823 & ~n10824 ;
  assign n10826 = ~n10767 & ~n10768 ;
  assign n10827 = ~n10790 & n10826 ;
  assign n10828 = n10790 & ~n10826 ;
  assign n10829 = ~n10827 & ~n10828 ;
  assign n10830 = ~n10825 & ~n10829 ;
  assign n10831 = n10825 & n10829 ;
  assign n10832 = ~n10136 & ~n10157 ;
  assign n10833 = ~n10778 & ~n10832 ;
  assign n10834 = n10140 & n10179 ;
  assign n10835 = ~n10140 & ~n10179 ;
  assign n10836 = ~n10834 & ~n10835 ;
  assign n10837 = ~n10833 & n10836 ;
  assign n10838 = n10833 & ~n10836 ;
  assign n10839 = ~n10726 & ~n10727 ;
  assign n10840 = ~n10135 & n10839 ;
  assign n10841 = n10135 & ~n10839 ;
  assign n10842 = ~n10840 & ~n10841 ;
  assign n10843 = ~n10838 & n10842 ;
  assign n10844 = ~n10837 & ~n10843 ;
  assign n10845 = n10249 & ~n10803 ;
  assign n10846 = ~n10249 & n10803 ;
  assign n10847 = ~n10845 & ~n10846 ;
  assign n10848 = ~n10844 & n10847 ;
  assign n10849 = n10844 & ~n10847 ;
  assign n10850 = ~n10776 & ~n10777 ;
  assign n10851 = ~n10788 & n10850 ;
  assign n10852 = n10788 & ~n10850 ;
  assign n10853 = ~n10851 & ~n10852 ;
  assign n10854 = ~n10849 & ~n10853 ;
  assign n10855 = ~n10848 & ~n10854 ;
  assign n10856 = ~n10831 & ~n10855 ;
  assign n10857 = ~n10830 & ~n10856 ;
  assign n10858 = ~n10808 & ~n10809 ;
  assign n10859 = n10813 & n10858 ;
  assign n10860 = ~n10813 & ~n10858 ;
  assign n10861 = ~n10859 & ~n10860 ;
  assign n10862 = n10857 & n10861 ;
  assign n10863 = ~n10821 & n10862 ;
  assign n10864 = ~n10820 & ~n10863 ;
  assign n10865 = n10759 & ~n10864 ;
  assign n10866 = n10672 & ~n10715 ;
  assign n10867 = n10753 & n10757 ;
  assign n10868 = ~n10716 & n10867 ;
  assign n10869 = ~n10866 & ~n10868 ;
  assign n10870 = ~n10865 & n10869 ;
  assign n10871 = ~n10857 & ~n10861 ;
  assign n10872 = ~n10821 & ~n10871 ;
  assign n10873 = n10759 & n10872 ;
  assign n10918 = ~n10393 & ~n10801 ;
  assign n10919 = n10137 & ~n10918 ;
  assign n10920 = ~n10137 & n10918 ;
  assign n10921 = ~n10919 & ~n10920 ;
  assign n10943 = ~n10139 & ~n10200 ;
  assign n10881 = n10136 & n10148 ;
  assign n10944 = n10139 & n10200 ;
  assign n10945 = ~n10881 & ~n10944 ;
  assign n10946 = ~n10943 & ~n10945 ;
  assign n10947 = n10921 & ~n10946 ;
  assign n10948 = ~n10921 & n10946 ;
  assign n10949 = ~n10769 & ~n10770 ;
  assign n10950 = n10395 & ~n10949 ;
  assign n10951 = ~n10395 & n10949 ;
  assign n10952 = ~n10950 & ~n10951 ;
  assign n10953 = ~n10948 & n10952 ;
  assign n10954 = ~n10947 & ~n10953 ;
  assign n10955 = ~n10848 & ~n10849 ;
  assign n10956 = ~n10853 & n10955 ;
  assign n10957 = n10853 & ~n10955 ;
  assign n10958 = ~n10956 & ~n10957 ;
  assign n10959 = ~n10954 & n10958 ;
  assign n10960 = n10954 & ~n10958 ;
  assign n10961 = ~n10959 & ~n10960 ;
  assign n10962 = ~n10135 & ~n10187 ;
  assign n10963 = ~n10186 & ~n10962 ;
  assign n10964 = ~n10175 & n10963 ;
  assign n10965 = n10175 & ~n10963 ;
  assign n10966 = ~n10723 & ~n10965 ;
  assign n10967 = ~n10964 & ~n10966 ;
  assign n10968 = ~n10837 & ~n10838 ;
  assign n10969 = n10842 & n10968 ;
  assign n10970 = ~n10842 & ~n10968 ;
  assign n10971 = ~n10969 & ~n10970 ;
  assign n10972 = ~n10967 & ~n10971 ;
  assign n10973 = n10967 & n10971 ;
  assign n10974 = ~n10947 & ~n10948 ;
  assign n10975 = n10952 & n10974 ;
  assign n10976 = ~n10952 & ~n10974 ;
  assign n10977 = ~n10975 & ~n10976 ;
  assign n10978 = ~n10973 & ~n10977 ;
  assign n10979 = ~n10972 & ~n10978 ;
  assign n10980 = n10961 & ~n10979 ;
  assign n10981 = ~n10961 & n10979 ;
  assign n10982 = ~n10980 & ~n10981 ;
  assign n10882 = ~n10136 & ~n10148 ;
  assign n10883 = ~n10881 & ~n10882 ;
  assign n10983 = ~n10150 & n10158 ;
  assign n10984 = n10883 & ~n10983 ;
  assign n10985 = n10150 & n10159 ;
  assign n10986 = ~n10984 & ~n10985 ;
  assign n10987 = ~n10139 & ~n10801 ;
  assign n10988 = ~n10393 & ~n10987 ;
  assign n10989 = ~n10135 & n10188 ;
  assign n10990 = n10135 & ~n10188 ;
  assign n10991 = ~n10989 & ~n10990 ;
  assign n10992 = ~n10988 & n10991 ;
  assign n10993 = n10988 & ~n10991 ;
  assign n10994 = ~n10161 & ~n10881 ;
  assign n10995 = n10161 & n10881 ;
  assign n10996 = ~n10395 & ~n10995 ;
  assign n10997 = ~n10994 & ~n10996 ;
  assign n10998 = ~n10993 & ~n10997 ;
  assign n10999 = ~n10992 & ~n10998 ;
  assign n11000 = n10986 & ~n10999 ;
  assign n11001 = ~n10986 & n10999 ;
  assign n11002 = ~n10964 & ~n10965 ;
  assign n11003 = ~n10723 & n11002 ;
  assign n11004 = n10723 & ~n11002 ;
  assign n11005 = ~n11003 & ~n11004 ;
  assign n11006 = ~n11001 & ~n11005 ;
  assign n11007 = ~n11000 & ~n11006 ;
  assign n11008 = ~n10972 & ~n10973 ;
  assign n11009 = ~n10977 & n11008 ;
  assign n11010 = n10977 & ~n11008 ;
  assign n11011 = ~n11009 & ~n11010 ;
  assign n11012 = n11007 & n11011 ;
  assign n11013 = ~n11007 & ~n11011 ;
  assign n11014 = ~n10140 & ~n10149 ;
  assign n11015 = ~n10151 & ~n11014 ;
  assign n11016 = ~n10197 & ~n11015 ;
  assign n11017 = ~n10198 & ~n11016 ;
  assign n11018 = n10148 & n11017 ;
  assign n11019 = ~n10148 & ~n11017 ;
  assign n11020 = ~n10943 & ~n10944 ;
  assign n11021 = n10881 & ~n11020 ;
  assign n11022 = ~n10881 & n11020 ;
  assign n11023 = ~n11021 & ~n11022 ;
  assign n11024 = ~n11019 & ~n11023 ;
  assign n11025 = ~n11018 & ~n11024 ;
  assign n11026 = ~n11013 & ~n11025 ;
  assign n11027 = ~n11012 & ~n11026 ;
  assign n11028 = ~n10982 & n11027 ;
  assign n11029 = ~n10959 & ~n10979 ;
  assign n11030 = ~n10960 & ~n11029 ;
  assign n11031 = ~n10830 & ~n10831 ;
  assign n11032 = ~n10855 & n11031 ;
  assign n11033 = n10855 & ~n11031 ;
  assign n11034 = ~n11032 & ~n11033 ;
  assign n11035 = n11030 & n11034 ;
  assign n11036 = ~n11028 & ~n11035 ;
  assign n11037 = ~n10266 & n11015 ;
  assign n11038 = ~n10198 & n11016 ;
  assign n11039 = ~n11037 & ~n11038 ;
  assign n11040 = ~n10140 & n10333 ;
  assign n11041 = n10140 & ~n10333 ;
  assign n11042 = ~n11040 & ~n11041 ;
  assign n11043 = ~n10175 & ~n11042 ;
  assign n11044 = n10175 & n11042 ;
  assign n11045 = n10139 & ~n10918 ;
  assign n11046 = ~n10139 & n10918 ;
  assign n11047 = ~n11045 & ~n11046 ;
  assign n11048 = ~n11044 & ~n11047 ;
  assign n11049 = ~n11043 & ~n11048 ;
  assign n11050 = ~n11039 & ~n11049 ;
  assign n11051 = n11039 & n11049 ;
  assign n11052 = n10984 & ~n10985 ;
  assign n11053 = ~n10172 & ~n10839 ;
  assign n11054 = ~n10883 & n11053 ;
  assign n11055 = ~n11052 & ~n11054 ;
  assign n11056 = ~n11051 & n11055 ;
  assign n11057 = ~n11050 & ~n11056 ;
  assign n11058 = ~n11018 & ~n11019 ;
  assign n11059 = ~n11023 & n11058 ;
  assign n11060 = n11023 & ~n11058 ;
  assign n11061 = ~n11059 & ~n11060 ;
  assign n11062 = ~n11057 & n11061 ;
  assign n11063 = n11057 & ~n11061 ;
  assign n11064 = ~n11000 & ~n11001 ;
  assign n11065 = ~n11005 & n11064 ;
  assign n11066 = n11005 & ~n11064 ;
  assign n11067 = ~n11065 & ~n11066 ;
  assign n11068 = ~n11063 & ~n11067 ;
  assign n11069 = ~n11062 & ~n11068 ;
  assign n11070 = ~n11012 & ~n11013 ;
  assign n11071 = ~n11025 & n11070 ;
  assign n11072 = n11025 & ~n11070 ;
  assign n11073 = ~n11071 & ~n11072 ;
  assign n11074 = n11069 & ~n11073 ;
  assign n11103 = ~n11062 & ~n11063 ;
  assign n11105 = n11067 & n11103 ;
  assign n11104 = ~n11067 & ~n11103 ;
  assign n11075 = ~n10994 & ~n10995 ;
  assign n11076 = n10395 & ~n11075 ;
  assign n11077 = ~n10395 & n11075 ;
  assign n11078 = ~n11076 & ~n11077 ;
  assign n11079 = ~n10137 & ~n10156 ;
  assign n11080 = \din[15]_pad  & n10137 ;
  assign n11081 = ~n10148 & ~n10187 ;
  assign n11082 = ~n10186 & ~n11081 ;
  assign n11083 = ~n11080 & ~n11082 ;
  assign n11084 = ~n11079 & ~n11083 ;
  assign n11085 = n11078 & ~n11084 ;
  assign n11086 = ~n11078 & n11084 ;
  assign n11087 = ~n10224 & n10883 ;
  assign n11088 = n10224 & ~n10883 ;
  assign n11089 = ~n10723 & ~n11088 ;
  assign n11090 = ~n11087 & ~n11089 ;
  assign n11091 = ~n11086 & n11090 ;
  assign n11092 = ~n11085 & ~n11091 ;
  assign n11093 = ~n10992 & ~n10993 ;
  assign n11094 = ~n10997 & n11093 ;
  assign n11095 = n10997 & ~n11093 ;
  assign n11096 = ~n11094 & ~n11095 ;
  assign n11097 = ~n11092 & n11096 ;
  assign n11098 = ~n11050 & ~n11051 ;
  assign n11099 = ~n11055 & n11098 ;
  assign n11100 = n11055 & ~n11098 ;
  assign n11101 = ~n11099 & ~n11100 ;
  assign n11102 = ~n11097 & ~n11101 ;
  assign n11106 = n11092 & ~n11096 ;
  assign n11107 = ~n11102 & ~n11106 ;
  assign n11108 = ~n11104 & n11107 ;
  assign n11109 = ~n11105 & n11108 ;
  assign n11110 = ~n11074 & ~n11109 ;
  assign n11111 = n11036 & n11110 ;
  assign n10874 = ~n10148 & ~n10163 ;
  assign n10875 = ~n10243 & ~n10874 ;
  assign n10876 = n10139 & n10295 ;
  assign n10877 = ~n10484 & ~n10876 ;
  assign n10878 = n10875 & ~n10877 ;
  assign n10879 = ~n10875 & n10877 ;
  assign n10880 = ~n10878 & ~n10879 ;
  assign n10884 = ~n10162 & ~n10883 ;
  assign n10885 = n10221 & n10883 ;
  assign n10886 = ~n10884 & ~n10885 ;
  assign n10887 = ~n10880 & n10886 ;
  assign n10888 = n10880 & ~n10886 ;
  assign n10889 = ~n10148 & ~n10157 ;
  assign n10890 = n10148 & n10157 ;
  assign n10891 = ~n10889 & ~n10890 ;
  assign n10892 = ~n10166 & n10891 ;
  assign n10893 = n10166 & ~n10891 ;
  assign n10894 = ~n10892 & ~n10893 ;
  assign n10895 = ~n10723 & ~n10894 ;
  assign n10896 = n10723 & n10894 ;
  assign n10897 = ~n10895 & ~n10896 ;
  assign n10898 = \din[9]_pad  & n10157 ;
  assign n10899 = ~n10140 & ~n10898 ;
  assign n10900 = ~n10889 & ~n10899 ;
  assign n10901 = ~n10137 & ~n10900 ;
  assign n10902 = n10137 & n10900 ;
  assign n10903 = ~n10140 & ~n10902 ;
  assign n10904 = ~n10901 & ~n10903 ;
  assign n10905 = ~n10897 & n10904 ;
  assign n10906 = n10897 & ~n10904 ;
  assign n10907 = ~n10905 & ~n10906 ;
  assign n10908 = ~n10888 & ~n10907 ;
  assign n10909 = ~n10887 & ~n10908 ;
  assign n10910 = ~\din[13]_pad  & ~n10898 ;
  assign n10911 = ~n10889 & ~n10910 ;
  assign n10912 = n10395 & n10911 ;
  assign n10913 = ~n10395 & ~n10911 ;
  assign n10914 = ~n10912 & ~n10913 ;
  assign n10915 = ~n10833 & n10914 ;
  assign n10916 = n10833 & ~n10914 ;
  assign n10917 = ~n10915 & ~n10916 ;
  assign n10922 = ~n10779 & ~n10780 ;
  assign n10923 = ~n10135 & n10922 ;
  assign n10924 = n10135 & ~n10922 ;
  assign n10925 = ~n10923 & ~n10924 ;
  assign n10926 = n10921 & n10925 ;
  assign n10927 = ~n10921 & ~n10925 ;
  assign n10928 = ~n10926 & ~n10927 ;
  assign n10929 = ~n10482 & ~n10875 ;
  assign n10930 = ~n10484 & ~n10929 ;
  assign n10931 = n10928 & ~n10930 ;
  assign n10932 = ~n10928 & n10930 ;
  assign n10933 = ~n10931 & ~n10932 ;
  assign n10934 = n10917 & n10933 ;
  assign n10935 = ~n10917 & ~n10933 ;
  assign n10936 = ~n10934 & ~n10935 ;
  assign n10937 = ~n10895 & ~n10904 ;
  assign n10938 = ~n10896 & ~n10937 ;
  assign n10939 = n10936 & ~n10938 ;
  assign n10940 = ~n10936 & n10938 ;
  assign n10941 = ~n10939 & ~n10940 ;
  assign n10942 = n10909 & n10941 ;
  assign n11112 = ~n10934 & n10938 ;
  assign n11113 = ~n10935 & ~n11112 ;
  assign n11114 = ~n10162 & n10922 ;
  assign n11115 = n10162 & ~n10922 ;
  assign n11116 = ~n11114 & ~n11115 ;
  assign n11117 = ~n10135 & ~n10780 ;
  assign n11118 = ~n10779 & ~n11117 ;
  assign n11119 = n10157 & n11118 ;
  assign n11120 = ~n10157 & ~n11118 ;
  assign n11121 = ~n11119 & ~n11120 ;
  assign n11122 = ~n10926 & n10930 ;
  assign n11123 = ~n10927 & ~n11122 ;
  assign n11124 = n11121 & ~n11123 ;
  assign n11125 = ~n11121 & n11123 ;
  assign n11126 = ~n11124 & ~n11125 ;
  assign n11127 = ~n10673 & n10778 ;
  assign n11128 = n10673 & ~n10778 ;
  assign n11129 = ~n11127 & ~n11128 ;
  assign n11130 = n10803 & ~n11129 ;
  assign n11131 = ~n10803 & n11129 ;
  assign n11132 = ~n11130 & ~n11131 ;
  assign n11133 = n11126 & n11132 ;
  assign n11134 = ~n11126 & ~n11132 ;
  assign n11135 = ~n11133 & ~n11134 ;
  assign n11136 = ~n10833 & ~n10912 ;
  assign n11137 = ~n10913 & ~n11136 ;
  assign n11138 = n11135 & ~n11137 ;
  assign n11139 = ~n11135 & n11137 ;
  assign n11140 = ~n11138 & ~n11139 ;
  assign n11141 = n11116 & n11140 ;
  assign n11142 = ~n11116 & ~n11140 ;
  assign n11143 = ~n11141 & ~n11142 ;
  assign n11144 = n11113 & ~n11143 ;
  assign n11145 = ~n10942 & ~n11144 ;
  assign n11146 = n11111 & n11145 ;
  assign n11147 = n10873 & n11146 ;
  assign n11148 = n10870 & ~n11147 ;
  assign n11149 = n10668 & ~n11148 ;
  assign n11158 = ~n11069 & n11073 ;
  assign n11159 = n11036 & n11158 ;
  assign n11160 = ~n11030 & ~n11034 ;
  assign n11161 = n10982 & ~n11027 ;
  assign n11162 = ~n11035 & n11161 ;
  assign n11163 = ~n11160 & ~n11162 ;
  assign n11164 = ~n11159 & n11163 ;
  assign n11165 = ~n11113 & n11143 ;
  assign n11167 = ~n11043 & ~n11044 ;
  assign n11168 = ~n11047 & n11167 ;
  assign n11169 = n11047 & ~n11167 ;
  assign n11170 = ~n11168 & ~n11169 ;
  assign n11171 = ~n10166 & ~n10220 ;
  assign n11172 = ~n10484 & ~n11171 ;
  assign n11173 = ~n11116 & ~n11120 ;
  assign n11174 = ~n11119 & ~n11173 ;
  assign n11175 = ~n11172 & n11174 ;
  assign n11176 = n11172 & ~n11174 ;
  assign n11177 = ~n11175 & ~n11176 ;
  assign n11178 = ~n11079 & ~n11080 ;
  assign n11179 = n11082 & ~n11178 ;
  assign n11180 = ~n11079 & n11083 ;
  assign n11181 = ~n11179 & ~n11180 ;
  assign n11182 = n11177 & ~n11181 ;
  assign n11183 = ~n11177 & n11181 ;
  assign n11184 = ~n11182 & ~n11183 ;
  assign n11185 = ~n11170 & ~n11184 ;
  assign n11166 = ~n11130 & ~n11137 ;
  assign n11186 = ~n11131 & ~n11166 ;
  assign n11187 = ~n11185 & n11186 ;
  assign n11188 = ~n11087 & ~n11088 ;
  assign n11189 = ~n10723 & n11188 ;
  assign n11190 = n10723 & ~n11188 ;
  assign n11191 = ~n11189 & ~n11190 ;
  assign n11192 = n11184 & n11191 ;
  assign n11193 = ~n11187 & ~n11192 ;
  assign n11194 = ~n11176 & n11181 ;
  assign n11195 = ~n11175 & ~n11194 ;
  assign n11196 = ~n11170 & ~n11195 ;
  assign n11197 = n11170 & n11195 ;
  assign n11198 = ~n11196 & ~n11197 ;
  assign n11199 = ~n11085 & ~n11086 ;
  assign n11200 = n11090 & n11199 ;
  assign n11201 = ~n11090 & ~n11199 ;
  assign n11202 = ~n11200 & ~n11201 ;
  assign n11203 = ~n11198 & ~n11202 ;
  assign n11204 = n11198 & n11202 ;
  assign n11205 = ~n11203 & ~n11204 ;
  assign n11206 = ~n11193 & ~n11205 ;
  assign n11208 = ~n11097 & ~n11106 ;
  assign n11210 = n11101 & n11208 ;
  assign n11209 = ~n11101 & ~n11208 ;
  assign n11207 = ~n11196 & ~n11202 ;
  assign n11211 = ~n11197 & ~n11207 ;
  assign n11212 = ~n11209 & n11211 ;
  assign n11213 = ~n11210 & n11212 ;
  assign n11214 = n11206 & ~n11213 ;
  assign n11215 = ~n11165 & ~n11214 ;
  assign n11216 = n11111 & ~n11215 ;
  assign n11217 = n11164 & ~n11216 ;
  assign n11218 = n10873 & ~n11217 ;
  assign n11219 = n10668 & n11218 ;
  assign n11152 = ~n10502 & ~n10504 ;
  assign n11153 = n10372 & ~n10428 ;
  assign n11154 = ~n10505 & n11153 ;
  assign n11155 = ~n11152 & ~n11154 ;
  assign n11156 = n10667 & ~n11155 ;
  assign n11150 = ~n10661 & n10665 ;
  assign n11151 = ~n10659 & n11150 ;
  assign n11157 = ~n10583 & ~n10658 ;
  assign n11220 = ~n11151 & ~n11157 ;
  assign n11221 = ~n11156 & n11220 ;
  assign n11222 = ~n11219 & n11221 ;
  assign n11223 = ~n11149 & n11222 ;
  assign n11224 = ~n10637 & n10655 ;
  assign n11225 = ~n10636 & ~n11224 ;
  assign n11226 = n11223 & n11225 ;
  assign n11227 = ~n11223 & ~n11225 ;
  assign n11228 = ~n11226 & ~n11227 ;
  assign n11229 = ~n10184 & ~n10644 ;
  assign n11230 = ~n10183 & ~n11229 ;
  assign n11231 = ~n10648 & ~n10652 ;
  assign n11232 = ~n10649 & ~n11231 ;
  assign n11233 = ~n10274 & ~n10460 ;
  assign n11234 = ~n10275 & n10460 ;
  assign n11235 = ~n11233 & ~n11234 ;
  assign n11236 = n11232 & ~n11235 ;
  assign n11237 = ~n11232 & n11235 ;
  assign n11238 = ~n11236 & ~n11237 ;
  assign n11239 = n10949 & ~n11238 ;
  assign n11240 = ~n10949 & n11238 ;
  assign n11241 = ~n11239 & ~n11240 ;
  assign n11242 = n11230 & ~n11241 ;
  assign n11243 = ~n11230 & n11241 ;
  assign n11244 = ~n11242 & ~n11243 ;
  assign n11245 = ~n10603 & ~n10605 ;
  assign n11246 = ~n10604 & ~n11245 ;
  assign n11247 = n10142 & ~n10373 ;
  assign n11248 = ~n10142 & n10373 ;
  assign n11249 = ~n11247 & ~n11248 ;
  assign n11250 = n11246 & n11249 ;
  assign n11251 = ~n11246 & ~n11249 ;
  assign n11252 = ~n11250 & ~n11251 ;
  assign n11253 = ~n10278 & ~n10589 ;
  assign n11254 = ~n10138 & ~n10588 ;
  assign n11255 = ~n11253 & ~n11254 ;
  assign n11256 = ~n10138 & n11253 ;
  assign n11257 = ~n11255 & ~n11256 ;
  assign n11258 = n11252 & ~n11257 ;
  assign n11259 = ~n11252 & n11257 ;
  assign n11260 = ~n11258 & ~n11259 ;
  assign n11261 = n10523 & ~n11042 ;
  assign n11262 = ~n10523 & n11042 ;
  assign n11263 = ~n11261 & ~n11262 ;
  assign n11264 = n11260 & ~n11263 ;
  assign n11265 = ~n11260 & n11263 ;
  assign n11266 = ~n11264 & ~n11265 ;
  assign n11267 = n11244 & ~n11266 ;
  assign n11268 = ~n11244 & n11266 ;
  assign n11269 = ~n11267 & ~n11268 ;
  assign n11270 = ~n10594 & ~n10598 ;
  assign n11271 = ~n10595 & ~n11270 ;
  assign n11272 = ~n10617 & ~n10621 ;
  assign n11273 = ~n10618 & ~n11272 ;
  assign n11274 = ~n10628 & ~n10632 ;
  assign n11275 = ~n10629 & ~n11274 ;
  assign n11276 = ~n11273 & n11275 ;
  assign n11277 = n11273 & ~n11275 ;
  assign n11278 = ~n11276 & ~n11277 ;
  assign n11279 = ~n10488 & n11278 ;
  assign n11280 = n10488 & ~n11278 ;
  assign n11281 = ~n11279 & ~n11280 ;
  assign n11282 = n11271 & n11281 ;
  assign n11283 = ~n11271 & ~n11281 ;
  assign n11284 = ~n11282 & ~n11283 ;
  assign n11285 = ~n10612 & ~n10624 ;
  assign n11286 = ~n10613 & ~n11285 ;
  assign n11287 = n11284 & ~n11286 ;
  assign n11288 = ~n11284 & n11286 ;
  assign n11289 = ~n11287 & ~n11288 ;
  assign n11290 = n11269 & n11289 ;
  assign n11291 = ~n11269 & ~n11289 ;
  assign n11292 = ~n11290 & ~n11291 ;
  assign n11293 = ~n11228 & ~n11292 ;
  assign n11294 = n11228 & n11292 ;
  assign n11295 = ~n11293 & ~n11294 ;
  assign n11296 = ~n10134 & ~n11295 ;
  assign n11347 = \P2_buf1_reg[23]/NET0131  & n10134 ;
  assign n11348 = ~n10862 & ~n10871 ;
  assign n11349 = ~n11146 & n11217 ;
  assign n11351 = ~n11348 & n11349 ;
  assign n11350 = n11348 & ~n11349 ;
  assign n11352 = ~n10134 & ~n11350 ;
  assign n11353 = ~n11351 & n11352 ;
  assign n11354 = ~n11347 & ~n11353 ;
  assign n11355 = \P2_buf1_reg[21]/NET0131  & n10134 ;
  assign n11356 = ~n11028 & ~n11161 ;
  assign n11357 = n11110 & ~n11213 ;
  assign n11302 = ~n10909 & ~n10941 ;
  assign n11303 = ~n11165 & ~n11302 ;
  assign n11304 = ~n11206 & n11303 ;
  assign n11305 = ~n10148 & ~n10220 ;
  assign n11306 = ~n10484 & ~n11305 ;
  assign n11307 = ~n10221 & ~n10883 ;
  assign n11308 = ~n10885 & ~n11307 ;
  assign n11309 = ~n10901 & ~n10902 ;
  assign n11310 = n10140 & ~n11309 ;
  assign n11311 = ~n10140 & n11309 ;
  assign n11312 = ~n11310 & ~n11311 ;
  assign n11313 = n11308 & n11312 ;
  assign n11314 = ~n11308 & ~n11312 ;
  assign n11315 = ~n11313 & ~n11314 ;
  assign n11316 = n11306 & n11315 ;
  assign n11317 = ~n11306 & ~n11315 ;
  assign n11318 = ~n11316 & ~n11317 ;
  assign n11319 = n10139 & n10157 ;
  assign n11320 = ~n10219 & ~n11319 ;
  assign n11321 = ~n10883 & n11320 ;
  assign n11322 = n10883 & ~n11320 ;
  assign n11323 = ~n11321 & ~n11322 ;
  assign n11324 = ~\din[1]_pad  & ~\din[5]_pad  ;
  assign n11325 = n10135 & ~n11324 ;
  assign n11326 = ~n11323 & ~n11325 ;
  assign n11327 = n11323 & n11325 ;
  assign n11328 = ~n10140 & n10891 ;
  assign n11329 = n10140 & ~n10891 ;
  assign n11330 = ~n11328 & ~n11329 ;
  assign n11331 = ~n11327 & n11330 ;
  assign n11332 = ~n11326 & ~n11331 ;
  assign n11333 = ~n11318 & ~n11332 ;
  assign n11358 = n11304 & n11333 ;
  assign n11359 = n11357 & ~n11358 ;
  assign n11360 = ~n11158 & ~n11359 ;
  assign n11362 = ~n11356 & n11360 ;
  assign n11361 = n11356 & ~n11360 ;
  assign n11363 = ~n10134 & ~n11361 ;
  assign n11364 = ~n11362 & n11363 ;
  assign n11365 = ~n11355 & ~n11364 ;
  assign n11297 = \P2_buf1_reg[22]/NET0131  & n10134 ;
  assign n11298 = ~n11035 & ~n11160 ;
  assign n11299 = ~n11158 & ~n11161 ;
  assign n11300 = ~n11028 & ~n11074 ;
  assign n11301 = ~n11213 & n11300 ;
  assign n11334 = ~n10942 & ~n11333 ;
  assign n11335 = n11304 & ~n11334 ;
  assign n11336 = n11301 & ~n11335 ;
  assign n11337 = n11299 & ~n11336 ;
  assign n11339 = ~n11298 & n11337 ;
  assign n11338 = n11298 & ~n11337 ;
  assign n11340 = ~n10134 & ~n11338 ;
  assign n11341 = ~n11339 & n11340 ;
  assign n11342 = ~n11297 & ~n11341 ;
  assign n11366 = \P2_buf1_reg[20]/NET0131  & n10134 ;
  assign n11367 = ~n11074 & ~n11158 ;
  assign n11369 = n11213 & ~n11367 ;
  assign n11368 = ~n11213 & n11367 ;
  assign n11370 = ~n10134 & ~n11368 ;
  assign n11371 = ~n11369 & n11370 ;
  assign n11372 = ~n11366 & ~n11371 ;
  assign n11377 = \P2_buf1_reg[15]/NET0131  & n10134 ;
  assign n11378 = \P2_buf1_reg[5]/NET0131  & n10134 ;
  assign n11391 = ~n11377 & ~n11378 ;
  assign n11379 = \P2_buf1_reg[0]/NET0131  & n10134 ;
  assign n11380 = \P2_buf1_reg[1]/NET0131  & n10134 ;
  assign n11392 = ~n11379 & ~n11380 ;
  assign n11399 = n11391 & n11392 ;
  assign n11373 = \P2_buf1_reg[10]/NET0131  & n10134 ;
  assign n11374 = \P2_buf1_reg[3]/NET0131  & n10134 ;
  assign n11389 = ~n11373 & ~n11374 ;
  assign n11375 = \P2_buf1_reg[12]/NET0131  & n10134 ;
  assign n11376 = \P2_buf1_reg[4]/NET0131  & n10134 ;
  assign n11390 = ~n11375 & ~n11376 ;
  assign n11400 = n11389 & n11390 ;
  assign n11401 = n11399 & n11400 ;
  assign n11385 = \P2_buf1_reg[8]/NET0131  & n10134 ;
  assign n11386 = \P2_buf1_reg[9]/NET0131  & n10134 ;
  assign n11395 = ~n11385 & ~n11386 ;
  assign n11387 = \P2_buf1_reg[7]/NET0131  & n10134 ;
  assign n11388 = \P2_buf1_reg[11]/NET0131  & n10134 ;
  assign n11396 = ~n11387 & ~n11388 ;
  assign n11397 = n11395 & n11396 ;
  assign n11381 = \P2_buf1_reg[14]/NET0131  & n10134 ;
  assign n11382 = \P2_buf1_reg[2]/NET0131  & n10134 ;
  assign n11393 = ~n11381 & ~n11382 ;
  assign n11383 = \P2_buf1_reg[6]/NET0131  & n10134 ;
  assign n11384 = \P2_buf1_reg[13]/NET0131  & n10134 ;
  assign n11394 = ~n11383 & ~n11384 ;
  assign n11398 = n11393 & n11394 ;
  assign n11402 = n11397 & n11398 ;
  assign n11403 = n11401 & n11402 ;
  assign n11343 = \P2_buf1_reg[19]/NET0131  & n10134 ;
  assign n11344 = \P2_buf1_reg[17]/NET0131  & n10134 ;
  assign n11404 = ~n11343 & ~n11344 ;
  assign n11345 = \P2_buf1_reg[18]/NET0131  & n10134 ;
  assign n11346 = \P2_buf1_reg[16]/NET0131  & n10134 ;
  assign n11405 = ~n11345 & ~n11346 ;
  assign n11406 = n11404 & n11405 ;
  assign n11407 = n11403 & n11406 ;
  assign n11408 = n11372 & n11407 ;
  assign n11409 = n11342 & n11408 ;
  assign n11410 = n11365 & n11409 ;
  assign n11411 = n11354 & n11410 ;
  assign n11412 = n11296 & ~n11411 ;
  assign n11413 = ~\P2_buf1_reg[24]/NET0131  & n10134 ;
  assign n11414 = ~n10820 & ~n10821 ;
  assign n11415 = ~n10862 & ~n11160 ;
  assign n11416 = ~n10871 & ~n11035 ;
  assign n11417 = ~n11299 & n11416 ;
  assign n11418 = n11415 & ~n11417 ;
  assign n11419 = n11318 & n11332 ;
  assign n11420 = ~n11326 & ~n11327 ;
  assign n11421 = n11330 & n11420 ;
  assign n11422 = ~n11330 & ~n11420 ;
  assign n11423 = ~n11421 & ~n11422 ;
  assign n11424 = \din[5]_pad  & n10136 ;
  assign n11425 = ~n10482 & ~n11424 ;
  assign n11426 = ~n11423 & ~n11425 ;
  assign n11427 = ~n11333 & n11426 ;
  assign n11428 = ~n11419 & ~n11427 ;
  assign n11429 = n11303 & n11428 ;
  assign n11430 = n10138 & ~n10140 ;
  assign n11432 = ~\din[5]_pad  & ~n10881 ;
  assign n11433 = ~n10882 & ~n11432 ;
  assign n11434 = n10295 & n11433 ;
  assign n11435 = ~n10295 & ~n11433 ;
  assign n11444 = ~n11330 & ~n11435 ;
  assign n11445 = ~n11434 & ~n11444 ;
  assign n11447 = n11315 & n11445 ;
  assign n11446 = ~n11315 & ~n11445 ;
  assign n11431 = ~n10139 & ~n10902 ;
  assign n11436 = ~n11434 & ~n11435 ;
  assign n11437 = ~n11330 & n11436 ;
  assign n11438 = n11330 & ~n11436 ;
  assign n11439 = ~n11437 & ~n11438 ;
  assign n11440 = ~n11431 & n11439 ;
  assign n11441 = ~n10139 & ~n11439 ;
  assign n11442 = ~n10221 & ~n10901 ;
  assign n11443 = ~n11441 & n11442 ;
  assign n11448 = ~n11440 & ~n11443 ;
  assign n11449 = ~n11446 & n11448 ;
  assign n11450 = ~n11447 & n11449 ;
  assign n11451 = ~n11430 & ~n11450 ;
  assign n11452 = n11334 & n11451 ;
  assign n11453 = ~n11144 & n11452 ;
  assign n11454 = ~n11214 & ~n11453 ;
  assign n11455 = n11429 & n11454 ;
  assign n11456 = n11300 & n11416 ;
  assign n11457 = ~n11455 & n11456 ;
  assign n11458 = n11418 & ~n11457 ;
  assign n11460 = n11414 & n11458 ;
  assign n11459 = ~n11414 & ~n11458 ;
  assign n11461 = ~n10134 & ~n11459 ;
  assign n11462 = ~n11460 & n11461 ;
  assign n11463 = ~n11413 & ~n11462 ;
  assign n11464 = n11412 & n11463 ;
  assign n11465 = \P2_buf1_reg[25]/NET0131  & n10134 ;
  assign n11466 = ~n10758 & ~n10867 ;
  assign n11467 = n10872 & ~n11163 ;
  assign n11468 = n10864 & ~n11467 ;
  assign n11469 = n10872 & n11036 ;
  assign n11470 = n11423 & n11425 ;
  assign n11471 = ~n11430 & ~n11470 ;
  assign n11472 = ~n11333 & n11471 ;
  assign n11473 = ~n11206 & ~n11472 ;
  assign n11474 = n11429 & n11473 ;
  assign n11475 = n11357 & ~n11474 ;
  assign n11476 = ~n11158 & ~n11475 ;
  assign n11477 = n11469 & ~n11476 ;
  assign n11478 = n11468 & ~n11477 ;
  assign n11480 = ~n11466 & n11478 ;
  assign n11479 = n11466 & ~n11478 ;
  assign n11481 = ~n10134 & ~n11479 ;
  assign n11482 = ~n11480 & n11481 ;
  assign n11483 = ~n11465 & ~n11482 ;
  assign n11484 = n11464 & ~n11483 ;
  assign n11485 = \P2_buf1_reg[26]/NET0131  & n10134 ;
  assign n11486 = ~n10716 & ~n10866 ;
  assign n11487 = ~n10758 & ~n10821 ;
  assign n11488 = ~n11415 & n11487 ;
  assign n11489 = ~n10820 & ~n10867 ;
  assign n11490 = ~n10758 & ~n11489 ;
  assign n11491 = ~n11488 & ~n11490 ;
  assign n11492 = n11416 & n11487 ;
  assign n11493 = ~n10942 & n11419 ;
  assign n11494 = n11470 & ~n11493 ;
  assign n11495 = n11304 & n11494 ;
  assign n11496 = n11301 & ~n11495 ;
  assign n11497 = n11299 & ~n11496 ;
  assign n11498 = n11492 & ~n11497 ;
  assign n11499 = n11491 & ~n11498 ;
  assign n11501 = ~n11486 & n11499 ;
  assign n11500 = n11486 & ~n11499 ;
  assign n11502 = ~n10134 & ~n11500 ;
  assign n11503 = ~n11501 & n11502 ;
  assign n11504 = ~n11485 & ~n11503 ;
  assign n11505 = n11484 & ~n11504 ;
  assign n11506 = \P2_buf1_reg[27]/NET0131  & n10134 ;
  assign n11507 = ~n10429 & ~n11153 ;
  assign n11508 = n11428 & n11430 ;
  assign n11509 = ~n11333 & ~n11508 ;
  assign n11510 = ~n11144 & n11509 ;
  assign n11511 = n11304 & ~n11510 ;
  assign n11512 = n11111 & ~n11511 ;
  assign n11513 = n11164 & ~n11512 ;
  assign n11514 = n10873 & ~n11513 ;
  assign n11515 = n10870 & ~n11514 ;
  assign n11517 = ~n11507 & n11515 ;
  assign n11516 = n11507 & ~n11515 ;
  assign n11518 = ~n10134 & ~n11516 ;
  assign n11519 = ~n11517 & n11518 ;
  assign n11520 = ~n11506 & ~n11519 ;
  assign n11521 = n11505 & ~n11520 ;
  assign n11522 = \P2_buf1_reg[28]/NET0131  & n10134 ;
  assign n11523 = ~n10505 & ~n11152 ;
  assign n11524 = ~n10429 & n10866 ;
  assign n11525 = ~n11153 & ~n11524 ;
  assign n11526 = ~n10429 & ~n10716 ;
  assign n11527 = n11301 & n11492 ;
  assign n11528 = ~n11418 & n11487 ;
  assign n11529 = ~n11490 & ~n11528 ;
  assign n11530 = ~n11527 & n11529 ;
  assign n11531 = n11526 & ~n11530 ;
  assign n11532 = n11525 & ~n11531 ;
  assign n11534 = ~n11523 & n11532 ;
  assign n11533 = n11523 & ~n11532 ;
  assign n11535 = ~n10134 & ~n11533 ;
  assign n11536 = ~n11534 & n11535 ;
  assign n11537 = ~n11522 & ~n11536 ;
  assign n11538 = n11521 & ~n11537 ;
  assign n11539 = \P2_buf1_reg[29]/NET0131  & n10134 ;
  assign n11540 = ~n10666 & ~n11150 ;
  assign n11544 = n10759 & ~n11468 ;
  assign n11545 = n10869 & ~n11544 ;
  assign n11546 = n10506 & ~n11545 ;
  assign n11541 = n10506 & n10759 ;
  assign n11542 = ~n11360 & n11541 ;
  assign n11543 = n11469 & n11542 ;
  assign n11547 = n11155 & ~n11543 ;
  assign n11548 = ~n11546 & n11547 ;
  assign n11550 = ~n11540 & n11548 ;
  assign n11549 = n11540 & ~n11548 ;
  assign n11551 = ~n10134 & ~n11549 ;
  assign n11552 = ~n11550 & n11551 ;
  assign n11553 = ~n11539 & ~n11552 ;
  assign n11554 = n11538 & ~n11553 ;
  assign n11555 = \P2_buf1_reg[30]/NET0131  & n10134 ;
  assign n11556 = ~n10659 & ~n11157 ;
  assign n11557 = ~n11337 & n11492 ;
  assign n11558 = n11491 & ~n11557 ;
  assign n11559 = n11526 & ~n11558 ;
  assign n11560 = ~n11152 & n11525 ;
  assign n11561 = ~n11559 & n11560 ;
  assign n11562 = ~n10505 & ~n10666 ;
  assign n11563 = ~n11561 & n11562 ;
  assign n11564 = ~n11150 & ~n11563 ;
  assign n11566 = ~n11556 & n11564 ;
  assign n11565 = n11556 & ~n11564 ;
  assign n11567 = ~n10134 & ~n11565 ;
  assign n11568 = ~n11566 & n11567 ;
  assign n11569 = ~n11555 & ~n11568 ;
  assign n11570 = n11554 & ~n11569 ;
  assign n11571 = n11296 & ~n11570 ;
  assign n11572 = ~n11296 & n11570 ;
  assign n11573 = ~n11571 & ~n11572 ;
  assign n11574 = n10105 & ~n11573 ;
  assign n11575 = \P2_P1_InstQueueWr_Addr_reg[0]/NET0131  & ~\P2_P1_InstQueueWr_Addr_reg[1]/NET0131  ;
  assign n11576 = ~\P2_P1_InstQueueWr_Addr_reg[2]/NET0131  & n11575 ;
  assign n11577 = \P2_P1_InstQueueWr_Addr_reg[3]/NET0131  & n11576 ;
  assign n11578 = n11296 & ~n11403 ;
  assign n11579 = n11346 & n11578 ;
  assign n11580 = \P2_buf1_reg[17]/NET0131  & n11579 ;
  assign n11581 = n11345 & n11580 ;
  assign n11582 = \P2_buf1_reg[19]/NET0131  & n11581 ;
  assign n11583 = n11366 & n11582 ;
  assign n11584 = ~n11365 & n11583 ;
  assign n11585 = ~n11342 & n11584 ;
  assign n11586 = n11354 & ~n11585 ;
  assign n11587 = ~n11354 & n11585 ;
  assign n11588 = ~n11586 & ~n11587 ;
  assign n11589 = n11577 & n11588 ;
  assign n11590 = ~n11574 & ~n11589 ;
  assign n11591 = \P2_P1_DataWidth_reg[1]/NET0131  & ~n11590 ;
  assign n11592 = ~n10105 & ~n11577 ;
  assign n11593 = \P2_P1_DataWidth_reg[1]/NET0131  & ~n11592 ;
  assign n11594 = \P2_P1_InstQueueWr_Addr_reg[0]/NET0131  & \P2_P1_InstQueueWr_Addr_reg[1]/NET0131  ;
  assign n11595 = ~\P2_P1_InstQueueWr_Addr_reg[2]/NET0131  & n11594 ;
  assign n11596 = \P2_P1_InstQueueWr_Addr_reg[3]/NET0131  & n11595 ;
  assign n11597 = ~\P2_P1_InstQueueWr_Addr_reg[0]/NET0131  & \P2_P1_InstQueueWr_Addr_reg[1]/NET0131  ;
  assign n11598 = ~\P2_P1_InstQueueWr_Addr_reg[2]/NET0131  & n11597 ;
  assign n11599 = \P2_P1_InstQueueWr_Addr_reg[3]/NET0131  & n11598 ;
  assign n11600 = ~n11596 & ~n11599 ;
  assign n11601 = n11387 & ~n11600 ;
  assign n11602 = \P2_P1_InstQueue_reg[11][7]/NET0131  & ~n11596 ;
  assign n11603 = ~n11599 & n11602 ;
  assign n11604 = ~n11601 & ~n11603 ;
  assign n11605 = ~n11593 & ~n11604 ;
  assign n11606 = ~n11591 & ~n11605 ;
  assign n11607 = \P2_P1_State2_reg[1]/NET0131  & ~\P2_P1_State2_reg[2]/NET0131  ;
  assign n11608 = ~\P2_P1_State2_reg[3]/NET0131  & n11607 ;
  assign n11609 = ~\P2_P1_State2_reg[0]/NET0131  & n11608 ;
  assign n11610 = ~n11606 & n11609 ;
  assign n11649 = \P2_P1_InstQueueRd_Addr_reg[1]/NET0131  & \P2_P1_InstQueueRd_Addr_reg[2]/NET0131  ;
  assign n11650 = ~\P2_P1_InstQueueRd_Addr_reg[3]/NET0131  & n11649 ;
  assign n11651 = ~\P2_P1_InstQueueRd_Addr_reg[0]/NET0131  & n11650 ;
  assign n11652 = \P2_P1_InstQueue_reg[6][7]/NET0131  & n11651 ;
  assign n11645 = \P2_P1_InstQueueRd_Addr_reg[0]/NET0131  & \P2_P1_InstQueueRd_Addr_reg[1]/NET0131  ;
  assign n11646 = \P2_P1_InstQueueRd_Addr_reg[2]/NET0131  & n11645 ;
  assign n11647 = \P2_P1_InstQueueRd_Addr_reg[3]/NET0131  & n11646 ;
  assign n11648 = \P2_P1_InstQueue_reg[15][7]/NET0131  & n11647 ;
  assign n11632 = ~\P2_P1_InstQueueRd_Addr_reg[0]/NET0131  & \P2_P1_InstQueueRd_Addr_reg[1]/NET0131  ;
  assign n11633 = ~\P2_P1_InstQueueRd_Addr_reg[2]/NET0131  & \P2_P1_InstQueueRd_Addr_reg[3]/NET0131  ;
  assign n11634 = n11632 & n11633 ;
  assign n11635 = \P2_P1_InstQueue_reg[10][7]/NET0131  & n11634 ;
  assign n11636 = \P2_P1_InstQueueRd_Addr_reg[0]/NET0131  & ~\P2_P1_InstQueueRd_Addr_reg[1]/NET0131  ;
  assign n11637 = \P2_P1_InstQueueRd_Addr_reg[2]/NET0131  & ~\P2_P1_InstQueueRd_Addr_reg[3]/NET0131  ;
  assign n11638 = n11636 & n11637 ;
  assign n11639 = \P2_P1_InstQueue_reg[5][7]/NET0131  & n11638 ;
  assign n11675 = ~n11635 & ~n11639 ;
  assign n11685 = ~n11648 & n11675 ;
  assign n11686 = ~n11652 & n11685 ;
  assign n11658 = ~\P2_P1_InstQueueRd_Addr_reg[0]/NET0131  & ~\P2_P1_InstQueueRd_Addr_reg[1]/NET0131  ;
  assign n11667 = n11637 & n11658 ;
  assign n11668 = \P2_P1_InstQueue_reg[4][7]/NET0131  & n11667 ;
  assign n11653 = ~\P2_P1_InstQueueRd_Addr_reg[2]/NET0131  & ~\P2_P1_InstQueueRd_Addr_reg[3]/NET0131  ;
  assign n11669 = n11653 & n11658 ;
  assign n11670 = \P2_P1_InstQueue_reg[0][7]/NET0131  & n11669 ;
  assign n11680 = ~n11668 & ~n11670 ;
  assign n11671 = n11636 & n11653 ;
  assign n11672 = \P2_P1_InstQueue_reg[1][7]/NET0131  & n11671 ;
  assign n11640 = \P2_P1_InstQueueRd_Addr_reg[2]/NET0131  & \P2_P1_InstQueueRd_Addr_reg[3]/NET0131  ;
  assign n11673 = n11640 & n11658 ;
  assign n11674 = \P2_P1_InstQueue_reg[12][7]/NET0131  & n11673 ;
  assign n11681 = ~n11672 & ~n11674 ;
  assign n11682 = n11680 & n11681 ;
  assign n11659 = n11633 & n11658 ;
  assign n11660 = \P2_P1_InstQueue_reg[8][7]/NET0131  & n11659 ;
  assign n11661 = n11637 & n11645 ;
  assign n11662 = \P2_P1_InstQueue_reg[7][7]/NET0131  & n11661 ;
  assign n11678 = ~n11660 & ~n11662 ;
  assign n11663 = n11645 & n11653 ;
  assign n11664 = \P2_P1_InstQueue_reg[3][7]/NET0131  & n11663 ;
  assign n11665 = n11633 & n11645 ;
  assign n11666 = \P2_P1_InstQueue_reg[11][7]/NET0131  & n11665 ;
  assign n11679 = ~n11664 & ~n11666 ;
  assign n11683 = n11678 & n11679 ;
  assign n11641 = n11636 & n11640 ;
  assign n11642 = \P2_P1_InstQueue_reg[13][7]/NET0131  & n11641 ;
  assign n11643 = n11632 & n11640 ;
  assign n11644 = \P2_P1_InstQueue_reg[14][7]/NET0131  & n11643 ;
  assign n11676 = ~n11642 & ~n11644 ;
  assign n11654 = n11632 & n11653 ;
  assign n11655 = \P2_P1_InstQueue_reg[2][7]/NET0131  & n11654 ;
  assign n11656 = n11633 & n11636 ;
  assign n11657 = \P2_P1_InstQueue_reg[9][7]/NET0131  & n11656 ;
  assign n11677 = ~n11655 & ~n11657 ;
  assign n11684 = n11676 & n11677 ;
  assign n11687 = n11683 & n11684 ;
  assign n11688 = n11682 & n11687 ;
  assign n11689 = n11686 & n11688 ;
  assign n11690 = n11596 & ~n11689 ;
  assign n11691 = ~n11602 & ~n11690 ;
  assign n11615 = ~\P2_P1_State2_reg[1]/NET0131  & ~\P2_P1_State2_reg[2]/NET0131  ;
  assign n11624 = \P2_P1_State2_reg[3]/NET0131  & n11615 ;
  assign n11692 = ~\P2_P1_State2_reg[0]/NET0131  & n11624 ;
  assign n11693 = ~n11691 & n11692 ;
  assign n11611 = ~\P2_P1_State2_reg[0]/NET0131  & ~\P2_P1_State2_reg[3]/NET0131  ;
  assign n11612 = ~\P2_P1_State2_reg[1]/NET0131  & \P2_P1_State2_reg[2]/NET0131  ;
  assign n11613 = n11611 & n11612 ;
  assign n11614 = ~n11604 & n11613 ;
  assign n11622 = \P2_P1_State2_reg[0]/NET0131  & ~\P2_P1_State2_reg[3]/NET0131  ;
  assign n11623 = n11612 & n11622 ;
  assign n11625 = \P2_P1_State2_reg[0]/NET0131  & n11624 ;
  assign n11626 = ~n11623 & ~n11625 ;
  assign n11616 = n11611 & n11615 ;
  assign n11617 = \P2_P1_State2_reg[0]/NET0131  & n11615 ;
  assign n11618 = ~\P2_P1_State2_reg[3]/NET0131  & n11617 ;
  assign n11619 = ~n11616 & ~n11618 ;
  assign n11620 = \P2_P1_State2_reg[1]/NET0131  & \P2_P1_State2_reg[2]/NET0131  ;
  assign n11621 = ~\P2_P1_State2_reg[3]/NET0131  & n11620 ;
  assign n11627 = \P2_P1_State2_reg[0]/NET0131  & n11608 ;
  assign n11628 = ~n11621 & ~n11627 ;
  assign n11629 = n11619 & n11628 ;
  assign n11630 = n11626 & n11629 ;
  assign n11631 = \P2_P1_InstQueue_reg[11][7]/NET0131  & ~n11630 ;
  assign n11694 = ~n11614 & ~n11631 ;
  assign n11695 = ~n11693 & n11694 ;
  assign n11696 = ~n11610 & n11695 ;
  assign n11697 = n8736 & ~n8741 ;
  assign n11698 = \P1_P3_DataWidth_reg[1]/NET0131  & n9245 ;
  assign n11699 = ~n8734 & ~n9241 ;
  assign n11700 = ~n11698 & n11699 ;
  assign n11701 = ~n11697 & n11700 ;
  assign n11703 = n8375 & n10050 ;
  assign n11704 = n8372 & n10053 ;
  assign n11705 = ~n11703 & ~n11704 ;
  assign n11706 = \P1_P1_DataWidth_reg[1]/NET0131  & ~n11705 ;
  assign n11707 = \P1_P1_DataWidth_reg[1]/NET0131  & ~n8474 ;
  assign n11708 = ~n7913 & ~n8379 ;
  assign n11709 = \P1_P1_InstQueue_reg[0][3]/NET0131  & ~n8376 ;
  assign n11710 = ~n8378 & n11709 ;
  assign n11711 = ~n11708 & ~n11710 ;
  assign n11712 = ~n11707 & ~n11711 ;
  assign n11713 = ~n11706 & ~n11712 ;
  assign n11714 = n8282 & ~n11713 ;
  assign n11715 = n8287 & ~n11711 ;
  assign n11702 = \P1_P1_InstQueue_reg[0][3]/NET0131  & ~n8366 ;
  assign n11716 = n8376 & ~n10096 ;
  assign n11717 = ~n11709 & ~n11716 ;
  assign n11718 = n8350 & ~n11717 ;
  assign n11719 = ~n11702 & ~n11718 ;
  assign n11720 = ~n11715 & n11719 ;
  assign n11721 = ~n11714 & n11720 ;
  assign n11723 = n8139 & n10053 ;
  assign n11724 = n8407 & n10050 ;
  assign n11725 = ~n11723 & ~n11724 ;
  assign n11726 = \P1_P1_DataWidth_reg[1]/NET0131  & ~n11725 ;
  assign n11727 = ~n7913 & ~n8401 ;
  assign n11728 = \P1_P1_InstQueue_reg[10][3]/NET0131  & ~n8145 ;
  assign n11729 = ~n4327 & n11728 ;
  assign n11730 = ~n11727 & ~n11729 ;
  assign n11731 = ~n9418 & ~n11730 ;
  assign n11732 = ~n11726 & ~n11731 ;
  assign n11733 = n8282 & ~n11732 ;
  assign n11734 = n8287 & ~n11730 ;
  assign n11722 = \P1_P1_InstQueue_reg[10][3]/NET0131  & ~n8366 ;
  assign n11735 = n8145 & ~n10096 ;
  assign n11736 = ~n11728 & ~n11735 ;
  assign n11737 = n8350 & ~n11736 ;
  assign n11738 = ~n11722 & ~n11737 ;
  assign n11739 = ~n11734 & n11738 ;
  assign n11740 = ~n11733 & n11739 ;
  assign n11742 = n4327 & n10050 ;
  assign n11743 = n8145 & n10053 ;
  assign n11744 = ~n11742 & ~n11743 ;
  assign n11745 = \P1_P1_DataWidth_reg[1]/NET0131  & ~n11744 ;
  assign n11746 = \P1_P1_DataWidth_reg[1]/NET0131  & ~n8401 ;
  assign n11747 = ~n7913 & ~n8428 ;
  assign n11748 = \P1_P1_InstQueue_reg[12][3]/NET0131  & ~n8427 ;
  assign n11749 = ~n8142 & n11748 ;
  assign n11750 = ~n11747 & ~n11749 ;
  assign n11751 = ~n11746 & ~n11750 ;
  assign n11752 = ~n11745 & ~n11751 ;
  assign n11753 = n8282 & ~n11752 ;
  assign n11754 = n8287 & ~n11750 ;
  assign n11741 = \P1_P1_InstQueue_reg[12][3]/NET0131  & ~n8366 ;
  assign n11755 = n8427 & ~n10096 ;
  assign n11756 = ~n11748 & ~n11755 ;
  assign n11757 = n8350 & ~n11756 ;
  assign n11758 = ~n11741 & ~n11757 ;
  assign n11759 = ~n11754 & n11758 ;
  assign n11760 = ~n11753 & n11759 ;
  assign n11762 = n8145 & n10050 ;
  assign n11763 = n8142 & n10053 ;
  assign n11764 = ~n11762 & ~n11763 ;
  assign n11765 = \P1_P1_DataWidth_reg[1]/NET0131  & ~n11764 ;
  assign n11766 = \P1_P1_DataWidth_reg[1]/NET0131  & ~n8146 ;
  assign n11767 = ~n7913 & ~n8451 ;
  assign n11768 = \P1_P1_InstQueue_reg[13][3]/NET0131  & ~n8375 ;
  assign n11769 = ~n8427 & n11768 ;
  assign n11770 = ~n11767 & ~n11769 ;
  assign n11771 = ~n11766 & ~n11770 ;
  assign n11772 = ~n11765 & ~n11771 ;
  assign n11773 = n8282 & ~n11772 ;
  assign n11774 = n8287 & ~n11770 ;
  assign n11761 = \P1_P1_InstQueue_reg[13][3]/NET0131  & ~n8366 ;
  assign n11775 = n8375 & ~n10096 ;
  assign n11776 = ~n11768 & ~n11775 ;
  assign n11777 = n8350 & ~n11776 ;
  assign n11778 = ~n11761 & ~n11777 ;
  assign n11779 = ~n11774 & n11778 ;
  assign n11780 = ~n11773 & n11779 ;
  assign n11782 = n8142 & n10050 ;
  assign n11783 = n8427 & n10053 ;
  assign n11784 = ~n11782 & ~n11783 ;
  assign n11785 = \P1_P1_DataWidth_reg[1]/NET0131  & ~n11784 ;
  assign n11786 = \P1_P1_DataWidth_reg[1]/NET0131  & ~n8428 ;
  assign n11787 = ~n7913 & ~n8474 ;
  assign n11788 = \P1_P1_InstQueue_reg[14][3]/NET0131  & ~n8372 ;
  assign n11789 = ~n8375 & n11788 ;
  assign n11790 = ~n11787 & ~n11789 ;
  assign n11791 = ~n11786 & ~n11790 ;
  assign n11792 = ~n11785 & ~n11791 ;
  assign n11793 = n8282 & ~n11792 ;
  assign n11794 = n8287 & ~n11790 ;
  assign n11781 = \P1_P1_InstQueue_reg[14][3]/NET0131  & ~n8366 ;
  assign n11795 = n8372 & ~n10096 ;
  assign n11796 = ~n11788 & ~n11795 ;
  assign n11797 = n8350 & ~n11796 ;
  assign n11798 = ~n11781 & ~n11797 ;
  assign n11799 = ~n11794 & n11798 ;
  assign n11800 = ~n11793 & n11799 ;
  assign n11802 = n8427 & n10050 ;
  assign n11803 = n8375 & n10053 ;
  assign n11804 = ~n11802 & ~n11803 ;
  assign n11805 = \P1_P1_DataWidth_reg[1]/NET0131  & ~n11804 ;
  assign n11806 = \P1_P1_DataWidth_reg[1]/NET0131  & ~n8451 ;
  assign n11807 = ~n7913 & ~n8497 ;
  assign n11808 = \P1_P1_InstQueue_reg[15][3]/NET0131  & ~n8378 ;
  assign n11809 = ~n8372 & n11808 ;
  assign n11810 = ~n11807 & ~n11809 ;
  assign n11811 = ~n11806 & ~n11810 ;
  assign n11812 = ~n11805 & ~n11811 ;
  assign n11813 = n8282 & ~n11812 ;
  assign n11814 = n8287 & ~n11810 ;
  assign n11801 = \P1_P1_InstQueue_reg[15][3]/NET0131  & ~n8366 ;
  assign n11815 = n8378 & ~n10096 ;
  assign n11816 = ~n11808 & ~n11815 ;
  assign n11817 = n8350 & ~n11816 ;
  assign n11818 = ~n11801 & ~n11817 ;
  assign n11819 = ~n11814 & n11818 ;
  assign n11820 = ~n11813 & n11819 ;
  assign n11822 = n8372 & n10050 ;
  assign n11823 = n8378 & n10053 ;
  assign n11824 = ~n11822 & ~n11823 ;
  assign n11825 = \P1_P1_DataWidth_reg[1]/NET0131  & ~n11824 ;
  assign n11826 = \P1_P1_DataWidth_reg[1]/NET0131  & ~n8497 ;
  assign n11827 = ~n7913 & ~n8521 ;
  assign n11828 = \P1_P1_InstQueue_reg[1][3]/NET0131  & ~n8520 ;
  assign n11829 = ~n8376 & n11828 ;
  assign n11830 = ~n11827 & ~n11829 ;
  assign n11831 = ~n11826 & ~n11830 ;
  assign n11832 = ~n11825 & ~n11831 ;
  assign n11833 = n8282 & ~n11832 ;
  assign n11834 = n8287 & ~n11830 ;
  assign n11821 = \P1_P1_InstQueue_reg[1][3]/NET0131  & ~n8366 ;
  assign n11835 = n8520 & ~n10096 ;
  assign n11836 = ~n11828 & ~n11835 ;
  assign n11837 = n8350 & ~n11836 ;
  assign n11838 = ~n11821 & ~n11837 ;
  assign n11839 = ~n11834 & n11838 ;
  assign n11840 = ~n11833 & n11839 ;
  assign n11842 = n8376 & n10053 ;
  assign n11843 = n8378 & n10050 ;
  assign n11844 = ~n11842 & ~n11843 ;
  assign n11845 = \P1_P1_DataWidth_reg[1]/NET0131  & ~n11844 ;
  assign n11846 = \P1_P1_DataWidth_reg[1]/NET0131  & ~n8379 ;
  assign n11847 = ~n7913 & ~n8545 ;
  assign n11848 = \P1_P1_InstQueue_reg[2][3]/NET0131  & ~n8544 ;
  assign n11849 = ~n8520 & n11848 ;
  assign n11850 = ~n11847 & ~n11849 ;
  assign n11851 = ~n11846 & ~n11850 ;
  assign n11852 = ~n11845 & ~n11851 ;
  assign n11853 = n8282 & ~n11852 ;
  assign n11854 = n8287 & ~n11850 ;
  assign n11841 = \P1_P1_InstQueue_reg[2][3]/NET0131  & ~n8366 ;
  assign n11855 = n8544 & ~n10096 ;
  assign n11856 = ~n11848 & ~n11855 ;
  assign n11857 = n8350 & ~n11856 ;
  assign n11858 = ~n11841 & ~n11857 ;
  assign n11859 = ~n11854 & n11858 ;
  assign n11860 = ~n11853 & n11859 ;
  assign n11861 = \P2_P1_InstQueueWr_Addr_reg[2]/NET0131  & n11575 ;
  assign n11862 = \P2_P1_InstQueueWr_Addr_reg[3]/NET0131  & n11861 ;
  assign n11863 = ~n11573 & n11862 ;
  assign n11864 = \P2_P1_InstQueueWr_Addr_reg[2]/NET0131  & n11597 ;
  assign n11865 = \P2_P1_InstQueueWr_Addr_reg[3]/NET0131  & n11864 ;
  assign n11866 = n11588 & n11865 ;
  assign n11867 = ~n11863 & ~n11866 ;
  assign n11868 = \P2_P1_DataWidth_reg[1]/NET0131  & ~n11867 ;
  assign n11869 = ~n11862 & ~n11865 ;
  assign n11870 = \P2_P1_DataWidth_reg[1]/NET0131  & ~n11869 ;
  assign n11871 = ~\P2_P1_InstQueueWr_Addr_reg[3]/NET0131  & n10104 ;
  assign n11872 = \P2_P1_InstQueueWr_Addr_reg[2]/NET0131  & n11594 ;
  assign n11873 = \P2_P1_InstQueueWr_Addr_reg[3]/NET0131  & n11872 ;
  assign n11874 = ~n11871 & ~n11873 ;
  assign n11875 = n11387 & ~n11874 ;
  assign n11876 = \P2_P1_InstQueue_reg[0][7]/NET0131  & ~n11871 ;
  assign n11877 = ~n11873 & n11876 ;
  assign n11878 = ~n11875 & ~n11877 ;
  assign n11879 = ~n11870 & ~n11878 ;
  assign n11880 = ~n11868 & ~n11879 ;
  assign n11881 = n11609 & ~n11880 ;
  assign n11884 = ~n11689 & n11871 ;
  assign n11885 = ~n11876 & ~n11884 ;
  assign n11886 = n11692 & ~n11885 ;
  assign n11882 = n11613 & ~n11878 ;
  assign n11883 = \P2_P1_InstQueue_reg[0][7]/NET0131  & ~n11630 ;
  assign n11887 = ~n11882 & ~n11883 ;
  assign n11888 = ~n11886 & n11887 ;
  assign n11889 = ~n11881 & n11888 ;
  assign n11890 = n10105 & n11588 ;
  assign n11891 = ~\P2_P1_InstQueueWr_Addr_reg[3]/NET0131  & n11872 ;
  assign n11892 = ~n11573 & n11891 ;
  assign n11893 = ~n11890 & ~n11892 ;
  assign n11894 = \P2_P1_DataWidth_reg[1]/NET0131  & ~n11893 ;
  assign n11895 = ~n10105 & ~n11891 ;
  assign n11896 = \P2_P1_DataWidth_reg[1]/NET0131  & ~n11895 ;
  assign n11897 = ~n11577 & ~n11599 ;
  assign n11898 = n11387 & ~n11897 ;
  assign n11899 = \P2_P1_InstQueue_reg[10][7]/NET0131  & ~n11599 ;
  assign n11900 = ~n11577 & n11899 ;
  assign n11901 = ~n11898 & ~n11900 ;
  assign n11902 = ~n11896 & ~n11901 ;
  assign n11903 = ~n11894 & ~n11902 ;
  assign n11904 = n11609 & ~n11903 ;
  assign n11907 = n11599 & ~n11689 ;
  assign n11908 = ~n11899 & ~n11907 ;
  assign n11909 = n11692 & ~n11908 ;
  assign n11905 = n11613 & ~n11901 ;
  assign n11906 = \P2_P1_InstQueue_reg[10][7]/NET0131  & ~n11630 ;
  assign n11910 = ~n11905 & ~n11906 ;
  assign n11911 = ~n11909 & n11910 ;
  assign n11912 = ~n11904 & n11911 ;
  assign n11913 = ~n11573 & n11577 ;
  assign n11914 = n11588 & n11599 ;
  assign n11915 = ~n11913 & ~n11914 ;
  assign n11916 = \P2_P1_DataWidth_reg[1]/NET0131  & ~n11915 ;
  assign n11917 = \P2_P1_DataWidth_reg[1]/NET0131  & ~n11897 ;
  assign n11918 = \P2_P1_InstQueueWr_Addr_reg[2]/NET0131  & n10103 ;
  assign n11919 = \P2_P1_InstQueueWr_Addr_reg[3]/NET0131  & n11918 ;
  assign n11920 = ~n11596 & ~n11919 ;
  assign n11921 = n11387 & ~n11920 ;
  assign n11922 = \P2_P1_InstQueue_reg[12][7]/NET0131  & ~n11919 ;
  assign n11923 = ~n11596 & n11922 ;
  assign n11924 = ~n11921 & ~n11923 ;
  assign n11925 = ~n11917 & ~n11924 ;
  assign n11926 = ~n11916 & ~n11925 ;
  assign n11927 = n11609 & ~n11926 ;
  assign n11930 = ~n11689 & n11919 ;
  assign n11931 = ~n11922 & ~n11930 ;
  assign n11932 = n11692 & ~n11931 ;
  assign n11928 = n11613 & ~n11924 ;
  assign n11929 = \P2_P1_InstQueue_reg[12][7]/NET0131  & ~n11630 ;
  assign n11933 = ~n11928 & ~n11929 ;
  assign n11934 = ~n11932 & n11933 ;
  assign n11935 = ~n11927 & n11934 ;
  assign n11937 = n8376 & n10050 ;
  assign n11938 = n8520 & n10053 ;
  assign n11939 = ~n11937 & ~n11938 ;
  assign n11940 = \P1_P1_DataWidth_reg[1]/NET0131  & ~n11939 ;
  assign n11941 = \P1_P1_DataWidth_reg[1]/NET0131  & ~n8521 ;
  assign n11942 = ~n7913 & ~n8569 ;
  assign n11943 = \P1_P1_InstQueue_reg[3][3]/NET0131  & ~n8568 ;
  assign n11944 = ~n8544 & n11943 ;
  assign n11945 = ~n11942 & ~n11944 ;
  assign n11946 = ~n11941 & ~n11945 ;
  assign n11947 = ~n11940 & ~n11946 ;
  assign n11948 = n8282 & ~n11947 ;
  assign n11949 = n8287 & ~n11945 ;
  assign n11936 = \P1_P1_InstQueue_reg[3][3]/NET0131  & ~n8366 ;
  assign n11950 = n8568 & ~n10096 ;
  assign n11951 = ~n11943 & ~n11950 ;
  assign n11952 = n8350 & ~n11951 ;
  assign n11953 = ~n11936 & ~n11952 ;
  assign n11954 = ~n11949 & n11953 ;
  assign n11955 = ~n11948 & n11954 ;
  assign n11956 = ~n11573 & n11599 ;
  assign n11957 = n11588 & n11596 ;
  assign n11958 = ~n11956 & ~n11957 ;
  assign n11959 = \P2_P1_DataWidth_reg[1]/NET0131  & ~n11958 ;
  assign n11960 = \P2_P1_DataWidth_reg[1]/NET0131  & ~n11600 ;
  assign n11961 = ~n11862 & ~n11919 ;
  assign n11962 = n11387 & ~n11961 ;
  assign n11963 = \P2_P1_InstQueue_reg[13][7]/NET0131  & ~n11862 ;
  assign n11964 = ~n11919 & n11963 ;
  assign n11965 = ~n11962 & ~n11964 ;
  assign n11966 = ~n11960 & ~n11965 ;
  assign n11967 = ~n11959 & ~n11966 ;
  assign n11968 = n11609 & ~n11967 ;
  assign n11971 = ~n11689 & n11862 ;
  assign n11972 = ~n11963 & ~n11971 ;
  assign n11973 = n11692 & ~n11972 ;
  assign n11969 = n11613 & ~n11965 ;
  assign n11970 = \P2_P1_InstQueue_reg[13][7]/NET0131  & ~n11630 ;
  assign n11974 = ~n11969 & ~n11970 ;
  assign n11975 = ~n11973 & n11974 ;
  assign n11976 = ~n11968 & n11975 ;
  assign n11977 = ~n11573 & n11596 ;
  assign n11978 = n11588 & n11919 ;
  assign n11979 = ~n11977 & ~n11978 ;
  assign n11980 = \P2_P1_DataWidth_reg[1]/NET0131  & ~n11979 ;
  assign n11981 = \P2_P1_DataWidth_reg[1]/NET0131  & ~n11920 ;
  assign n11982 = n11387 & ~n11869 ;
  assign n11983 = \P2_P1_InstQueue_reg[14][7]/NET0131  & ~n11865 ;
  assign n11984 = ~n11862 & n11983 ;
  assign n11985 = ~n11982 & ~n11984 ;
  assign n11986 = ~n11981 & ~n11985 ;
  assign n11987 = ~n11980 & ~n11986 ;
  assign n11988 = n11609 & ~n11987 ;
  assign n11991 = ~n11689 & n11865 ;
  assign n11992 = ~n11983 & ~n11991 ;
  assign n11993 = n11692 & ~n11992 ;
  assign n11989 = n11613 & ~n11985 ;
  assign n11990 = \P2_P1_InstQueue_reg[14][7]/NET0131  & ~n11630 ;
  assign n11994 = ~n11989 & ~n11990 ;
  assign n11995 = ~n11993 & n11994 ;
  assign n11996 = ~n11988 & n11995 ;
  assign n11997 = ~n11573 & n11919 ;
  assign n11998 = n11588 & n11862 ;
  assign n11999 = ~n11997 & ~n11998 ;
  assign n12000 = \P2_P1_DataWidth_reg[1]/NET0131  & ~n11999 ;
  assign n12001 = \P2_P1_DataWidth_reg[1]/NET0131  & ~n11961 ;
  assign n12002 = ~n11865 & ~n11873 ;
  assign n12003 = n11387 & ~n12002 ;
  assign n12004 = \P2_P1_InstQueue_reg[15][7]/NET0131  & ~n11873 ;
  assign n12005 = ~n11865 & n12004 ;
  assign n12006 = ~n12003 & ~n12005 ;
  assign n12007 = ~n12001 & ~n12006 ;
  assign n12008 = ~n12000 & ~n12007 ;
  assign n12009 = n11609 & ~n12008 ;
  assign n12012 = ~n11689 & n11873 ;
  assign n12013 = ~n12004 & ~n12012 ;
  assign n12014 = n11692 & ~n12013 ;
  assign n12010 = n11613 & ~n12006 ;
  assign n12011 = \P2_P1_InstQueue_reg[15][7]/NET0131  & ~n11630 ;
  assign n12015 = ~n12010 & ~n12011 ;
  assign n12016 = ~n12014 & n12015 ;
  assign n12017 = ~n12009 & n12016 ;
  assign n12018 = ~n11573 & n11865 ;
  assign n12019 = n11588 & n11873 ;
  assign n12020 = ~n12018 & ~n12019 ;
  assign n12021 = \P2_P1_DataWidth_reg[1]/NET0131  & ~n12020 ;
  assign n12022 = \P2_P1_DataWidth_reg[1]/NET0131  & ~n12002 ;
  assign n12023 = ~\P2_P1_InstQueueWr_Addr_reg[3]/NET0131  & n11576 ;
  assign n12024 = ~n11871 & ~n12023 ;
  assign n12025 = n11387 & ~n12024 ;
  assign n12026 = \P2_P1_InstQueue_reg[1][7]/NET0131  & ~n12023 ;
  assign n12027 = ~n11871 & n12026 ;
  assign n12028 = ~n12025 & ~n12027 ;
  assign n12029 = ~n12022 & ~n12028 ;
  assign n12030 = ~n12021 & ~n12029 ;
  assign n12031 = n11609 & ~n12030 ;
  assign n12034 = ~n11689 & n12023 ;
  assign n12035 = ~n12026 & ~n12034 ;
  assign n12036 = n11692 & ~n12035 ;
  assign n12032 = n11613 & ~n12028 ;
  assign n12033 = \P2_P1_InstQueue_reg[1][7]/NET0131  & ~n11630 ;
  assign n12037 = ~n12032 & ~n12033 ;
  assign n12038 = ~n12036 & n12037 ;
  assign n12039 = ~n12031 & n12038 ;
  assign n12041 = n8520 & n10050 ;
  assign n12042 = n8544 & n10053 ;
  assign n12043 = ~n12041 & ~n12042 ;
  assign n12044 = \P1_P1_DataWidth_reg[1]/NET0131  & ~n12043 ;
  assign n12045 = \P1_P1_DataWidth_reg[1]/NET0131  & ~n8545 ;
  assign n12046 = ~n7913 & ~n8593 ;
  assign n12047 = \P1_P1_InstQueue_reg[4][3]/NET0131  & ~n8592 ;
  assign n12048 = ~n8568 & n12047 ;
  assign n12049 = ~n12046 & ~n12048 ;
  assign n12050 = ~n12045 & ~n12049 ;
  assign n12051 = ~n12044 & ~n12050 ;
  assign n12052 = n8282 & ~n12051 ;
  assign n12053 = n8287 & ~n12049 ;
  assign n12040 = \P1_P1_InstQueue_reg[4][3]/NET0131  & ~n8366 ;
  assign n12054 = n8592 & ~n10096 ;
  assign n12055 = ~n12047 & ~n12054 ;
  assign n12056 = n8350 & ~n12055 ;
  assign n12057 = ~n12040 & ~n12056 ;
  assign n12058 = ~n12053 & n12057 ;
  assign n12059 = ~n12052 & n12058 ;
  assign n12060 = n11588 & n11871 ;
  assign n12061 = ~n11573 & n11873 ;
  assign n12062 = ~n12060 & ~n12061 ;
  assign n12063 = \P2_P1_DataWidth_reg[1]/NET0131  & ~n12062 ;
  assign n12064 = \P2_P1_DataWidth_reg[1]/NET0131  & ~n11874 ;
  assign n12065 = ~\P2_P1_InstQueueWr_Addr_reg[3]/NET0131  & n11598 ;
  assign n12066 = ~n12023 & ~n12065 ;
  assign n12067 = n11387 & ~n12066 ;
  assign n12068 = \P2_P1_InstQueue_reg[2][7]/NET0131  & ~n12065 ;
  assign n12069 = ~n12023 & n12068 ;
  assign n12070 = ~n12067 & ~n12069 ;
  assign n12071 = ~n12064 & ~n12070 ;
  assign n12072 = ~n12063 & ~n12071 ;
  assign n12073 = n11609 & ~n12072 ;
  assign n12076 = ~n11689 & n12065 ;
  assign n12077 = ~n12068 & ~n12076 ;
  assign n12078 = n11692 & ~n12077 ;
  assign n12074 = n11613 & ~n12070 ;
  assign n12075 = \P2_P1_InstQueue_reg[2][7]/NET0131  & ~n11630 ;
  assign n12079 = ~n12074 & ~n12075 ;
  assign n12080 = ~n12078 & n12079 ;
  assign n12081 = ~n12073 & n12080 ;
  assign n12082 = ~n11573 & n11871 ;
  assign n12083 = n11588 & n12023 ;
  assign n12084 = ~n12082 & ~n12083 ;
  assign n12085 = \P2_P1_DataWidth_reg[1]/NET0131  & ~n12084 ;
  assign n12086 = \P2_P1_DataWidth_reg[1]/NET0131  & ~n12024 ;
  assign n12087 = ~\P2_P1_InstQueueWr_Addr_reg[3]/NET0131  & n11595 ;
  assign n12088 = ~n12065 & ~n12087 ;
  assign n12089 = n11387 & ~n12088 ;
  assign n12090 = \P2_P1_InstQueue_reg[3][7]/NET0131  & ~n12087 ;
  assign n12091 = ~n12065 & n12090 ;
  assign n12092 = ~n12089 & ~n12091 ;
  assign n12093 = ~n12086 & ~n12092 ;
  assign n12094 = ~n12085 & ~n12093 ;
  assign n12095 = n11609 & ~n12094 ;
  assign n12098 = ~n11689 & n12087 ;
  assign n12099 = ~n12090 & ~n12098 ;
  assign n12100 = n11692 & ~n12099 ;
  assign n12096 = n11613 & ~n12092 ;
  assign n12097 = \P2_P1_InstQueue_reg[3][7]/NET0131  & ~n11630 ;
  assign n12101 = ~n12096 & ~n12097 ;
  assign n12102 = ~n12100 & n12101 ;
  assign n12103 = ~n12095 & n12102 ;
  assign n12104 = ~n11573 & n12023 ;
  assign n12105 = n11588 & n12065 ;
  assign n12106 = ~n12104 & ~n12105 ;
  assign n12107 = \P2_P1_DataWidth_reg[1]/NET0131  & ~n12106 ;
  assign n12108 = \P2_P1_DataWidth_reg[1]/NET0131  & ~n12066 ;
  assign n12109 = ~\P2_P1_InstQueueWr_Addr_reg[3]/NET0131  & n11918 ;
  assign n12110 = ~n12087 & ~n12109 ;
  assign n12111 = n11387 & ~n12110 ;
  assign n12112 = \P2_P1_InstQueue_reg[4][7]/NET0131  & ~n12109 ;
  assign n12113 = ~n12087 & n12112 ;
  assign n12114 = ~n12111 & ~n12113 ;
  assign n12115 = ~n12108 & ~n12114 ;
  assign n12116 = ~n12107 & ~n12115 ;
  assign n12117 = n11609 & ~n12116 ;
  assign n12120 = ~n11689 & n12109 ;
  assign n12121 = ~n12112 & ~n12120 ;
  assign n12122 = n11692 & ~n12121 ;
  assign n12118 = n11613 & ~n12114 ;
  assign n12119 = \P2_P1_InstQueue_reg[4][7]/NET0131  & ~n11630 ;
  assign n12123 = ~n12118 & ~n12119 ;
  assign n12124 = ~n12122 & n12123 ;
  assign n12125 = ~n12117 & n12124 ;
  assign n12126 = ~n11573 & n12065 ;
  assign n12127 = n11588 & n12087 ;
  assign n12128 = ~n12126 & ~n12127 ;
  assign n12129 = \P2_P1_DataWidth_reg[1]/NET0131  & ~n12128 ;
  assign n12130 = \P2_P1_DataWidth_reg[1]/NET0131  & ~n12088 ;
  assign n12131 = ~\P2_P1_InstQueueWr_Addr_reg[3]/NET0131  & n11861 ;
  assign n12132 = ~n12109 & ~n12131 ;
  assign n12133 = n11387 & ~n12132 ;
  assign n12134 = \P2_P1_InstQueue_reg[5][7]/NET0131  & ~n12131 ;
  assign n12135 = ~n12109 & n12134 ;
  assign n12136 = ~n12133 & ~n12135 ;
  assign n12137 = ~n12130 & ~n12136 ;
  assign n12138 = ~n12129 & ~n12137 ;
  assign n12139 = n11609 & ~n12138 ;
  assign n12142 = ~n11689 & n12131 ;
  assign n12143 = ~n12134 & ~n12142 ;
  assign n12144 = n11692 & ~n12143 ;
  assign n12140 = n11613 & ~n12136 ;
  assign n12141 = \P2_P1_InstQueue_reg[5][7]/NET0131  & ~n11630 ;
  assign n12145 = ~n12140 & ~n12141 ;
  assign n12146 = ~n12144 & n12145 ;
  assign n12147 = ~n12139 & n12146 ;
  assign n12149 = n8544 & n10050 ;
  assign n12150 = n8568 & n10053 ;
  assign n12151 = ~n12149 & ~n12150 ;
  assign n12152 = \P1_P1_DataWidth_reg[1]/NET0131  & ~n12151 ;
  assign n12153 = \P1_P1_DataWidth_reg[1]/NET0131  & ~n8569 ;
  assign n12154 = ~n7913 & ~n8617 ;
  assign n12155 = \P1_P1_InstQueue_reg[5][3]/NET0131  & ~n8616 ;
  assign n12156 = ~n8592 & n12155 ;
  assign n12157 = ~n12154 & ~n12156 ;
  assign n12158 = ~n12153 & ~n12157 ;
  assign n12159 = ~n12152 & ~n12158 ;
  assign n12160 = n8282 & ~n12159 ;
  assign n12161 = n8287 & ~n12157 ;
  assign n12148 = \P1_P1_InstQueue_reg[5][3]/NET0131  & ~n8366 ;
  assign n12162 = n8616 & ~n10096 ;
  assign n12163 = ~n12155 & ~n12162 ;
  assign n12164 = n8350 & ~n12163 ;
  assign n12165 = ~n12148 & ~n12164 ;
  assign n12166 = ~n12161 & n12165 ;
  assign n12167 = ~n12160 & n12166 ;
  assign n12168 = ~n11573 & n12087 ;
  assign n12169 = n11588 & n12109 ;
  assign n12170 = ~n12168 & ~n12169 ;
  assign n12171 = \P2_P1_DataWidth_reg[1]/NET0131  & ~n12170 ;
  assign n12172 = \P2_P1_DataWidth_reg[1]/NET0131  & ~n12110 ;
  assign n12173 = ~\P2_P1_InstQueueWr_Addr_reg[3]/NET0131  & n11864 ;
  assign n12174 = ~n12131 & ~n12173 ;
  assign n12175 = n11387 & ~n12174 ;
  assign n12176 = \P2_P1_InstQueue_reg[6][7]/NET0131  & ~n12173 ;
  assign n12177 = ~n12131 & n12176 ;
  assign n12178 = ~n12175 & ~n12177 ;
  assign n12179 = ~n12172 & ~n12178 ;
  assign n12180 = ~n12171 & ~n12179 ;
  assign n12181 = n11609 & ~n12180 ;
  assign n12184 = ~n11689 & n12173 ;
  assign n12185 = ~n12176 & ~n12184 ;
  assign n12186 = n11692 & ~n12185 ;
  assign n12182 = n11613 & ~n12178 ;
  assign n12183 = \P2_P1_InstQueue_reg[6][7]/NET0131  & ~n11630 ;
  assign n12187 = ~n12182 & ~n12183 ;
  assign n12188 = ~n12186 & n12187 ;
  assign n12189 = ~n12181 & n12188 ;
  assign n12190 = ~n11573 & n12109 ;
  assign n12191 = n11588 & n12131 ;
  assign n12192 = ~n12190 & ~n12191 ;
  assign n12193 = \P2_P1_DataWidth_reg[1]/NET0131  & ~n12192 ;
  assign n12194 = \P2_P1_DataWidth_reg[1]/NET0131  & ~n12132 ;
  assign n12195 = ~n11891 & ~n12173 ;
  assign n12196 = n11387 & ~n12195 ;
  assign n12197 = \P2_P1_InstQueue_reg[7][7]/NET0131  & ~n11891 ;
  assign n12198 = ~n12173 & n12197 ;
  assign n12199 = ~n12196 & ~n12198 ;
  assign n12200 = ~n12194 & ~n12199 ;
  assign n12201 = ~n12193 & ~n12200 ;
  assign n12202 = n11609 & ~n12201 ;
  assign n12205 = ~n11689 & n11891 ;
  assign n12206 = ~n12197 & ~n12205 ;
  assign n12207 = n11692 & ~n12206 ;
  assign n12203 = n11613 & ~n12199 ;
  assign n12204 = \P2_P1_InstQueue_reg[7][7]/NET0131  & ~n11630 ;
  assign n12208 = ~n12203 & ~n12204 ;
  assign n12209 = ~n12207 & n12208 ;
  assign n12210 = ~n12202 & n12209 ;
  assign n12211 = ~n11573 & n12131 ;
  assign n12212 = n11588 & n12173 ;
  assign n12213 = ~n12211 & ~n12212 ;
  assign n12214 = \P2_P1_DataWidth_reg[1]/NET0131  & ~n12213 ;
  assign n12215 = \P2_P1_DataWidth_reg[1]/NET0131  & ~n12174 ;
  assign n12216 = n11387 & ~n11895 ;
  assign n12217 = \P2_P1_InstQueue_reg[8][7]/NET0131  & ~n10105 ;
  assign n12218 = ~n11891 & n12217 ;
  assign n12219 = ~n12216 & ~n12218 ;
  assign n12220 = ~n12215 & ~n12219 ;
  assign n12221 = ~n12214 & ~n12220 ;
  assign n12222 = n11609 & ~n12221 ;
  assign n12225 = n10105 & ~n11689 ;
  assign n12226 = ~n12217 & ~n12225 ;
  assign n12227 = n11692 & ~n12226 ;
  assign n12223 = n11613 & ~n12219 ;
  assign n12224 = \P2_P1_InstQueue_reg[8][7]/NET0131  & ~n11630 ;
  assign n12228 = ~n12223 & ~n12224 ;
  assign n12229 = ~n12227 & n12228 ;
  assign n12230 = ~n12222 & n12229 ;
  assign n12231 = ~n11573 & n12173 ;
  assign n12232 = n11588 & n11891 ;
  assign n12233 = ~n12231 & ~n12232 ;
  assign n12234 = \P2_P1_DataWidth_reg[1]/NET0131  & ~n12233 ;
  assign n12235 = \P2_P1_DataWidth_reg[1]/NET0131  & ~n12195 ;
  assign n12236 = n11387 & ~n11592 ;
  assign n12237 = \P2_P1_InstQueue_reg[9][7]/NET0131  & ~n11577 ;
  assign n12238 = ~n10105 & n12237 ;
  assign n12239 = ~n12236 & ~n12238 ;
  assign n12240 = ~n12235 & ~n12239 ;
  assign n12241 = ~n12234 & ~n12240 ;
  assign n12242 = n11609 & ~n12241 ;
  assign n12245 = n11577 & ~n11689 ;
  assign n12246 = ~n12237 & ~n12245 ;
  assign n12247 = n11692 & ~n12246 ;
  assign n12243 = n11613 & ~n12239 ;
  assign n12244 = \P2_P1_InstQueue_reg[9][7]/NET0131  & ~n11630 ;
  assign n12248 = ~n12243 & ~n12244 ;
  assign n12249 = ~n12247 & n12248 ;
  assign n12250 = ~n12242 & n12249 ;
  assign n12252 = n8568 & n10050 ;
  assign n12253 = n8592 & n10053 ;
  assign n12254 = ~n12252 & ~n12253 ;
  assign n12255 = \P1_P1_DataWidth_reg[1]/NET0131  & ~n12254 ;
  assign n12256 = \P1_P1_DataWidth_reg[1]/NET0131  & ~n8593 ;
  assign n12257 = ~n7913 & ~n8641 ;
  assign n12258 = \P1_P1_InstQueue_reg[6][3]/NET0131  & ~n8640 ;
  assign n12259 = ~n8616 & n12258 ;
  assign n12260 = ~n12257 & ~n12259 ;
  assign n12261 = ~n12256 & ~n12260 ;
  assign n12262 = ~n12255 & ~n12261 ;
  assign n12263 = n8282 & ~n12262 ;
  assign n12264 = n8287 & ~n12260 ;
  assign n12251 = \P1_P1_InstQueue_reg[6][3]/NET0131  & ~n8366 ;
  assign n12265 = n8640 & ~n10096 ;
  assign n12266 = ~n12258 & ~n12265 ;
  assign n12267 = n8350 & ~n12266 ;
  assign n12268 = ~n12251 & ~n12267 ;
  assign n12269 = ~n12264 & n12268 ;
  assign n12270 = ~n12263 & n12269 ;
  assign n12272 = n8592 & n10050 ;
  assign n12273 = n8616 & n10053 ;
  assign n12274 = ~n12272 & ~n12273 ;
  assign n12275 = \P1_P1_DataWidth_reg[1]/NET0131  & ~n12274 ;
  assign n12276 = \P1_P1_DataWidth_reg[1]/NET0131  & ~n8617 ;
  assign n12277 = ~n7913 & ~n8664 ;
  assign n12278 = \P1_P1_InstQueue_reg[7][3]/NET0131  & ~n8407 ;
  assign n12279 = ~n8640 & n12278 ;
  assign n12280 = ~n12277 & ~n12279 ;
  assign n12281 = ~n12276 & ~n12280 ;
  assign n12282 = ~n12275 & ~n12281 ;
  assign n12283 = n8282 & ~n12282 ;
  assign n12284 = n8287 & ~n12280 ;
  assign n12271 = \P1_P1_InstQueue_reg[7][3]/NET0131  & ~n8366 ;
  assign n12285 = n8407 & ~n10096 ;
  assign n12286 = ~n12278 & ~n12285 ;
  assign n12287 = n8350 & ~n12286 ;
  assign n12288 = ~n12271 & ~n12287 ;
  assign n12289 = ~n12284 & n12288 ;
  assign n12290 = ~n12283 & n12289 ;
  assign n12292 = n8616 & n10050 ;
  assign n12293 = n8640 & n10053 ;
  assign n12294 = ~n12292 & ~n12293 ;
  assign n12295 = \P1_P1_DataWidth_reg[1]/NET0131  & ~n12294 ;
  assign n12296 = \P1_P1_DataWidth_reg[1]/NET0131  & ~n8641 ;
  assign n12297 = ~n7913 & ~n8410 ;
  assign n12298 = \P1_P1_InstQueue_reg[8][3]/NET0131  & ~n8139 ;
  assign n12299 = ~n8407 & n12298 ;
  assign n12300 = ~n12297 & ~n12299 ;
  assign n12301 = ~n12296 & ~n12300 ;
  assign n12302 = ~n12295 & ~n12301 ;
  assign n12303 = n8282 & ~n12302 ;
  assign n12304 = n8287 & ~n12300 ;
  assign n12291 = \P1_P1_InstQueue_reg[8][3]/NET0131  & ~n8366 ;
  assign n12305 = n8139 & ~n10096 ;
  assign n12306 = ~n12298 & ~n12305 ;
  assign n12307 = n8350 & ~n12306 ;
  assign n12308 = ~n12291 & ~n12307 ;
  assign n12309 = ~n12304 & n12308 ;
  assign n12310 = ~n12303 & n12309 ;
  assign n12312 = n8640 & n10050 ;
  assign n12313 = n8407 & n10053 ;
  assign n12314 = ~n12312 & ~n12313 ;
  assign n12315 = \P1_P1_DataWidth_reg[1]/NET0131  & ~n12314 ;
  assign n12316 = \P1_P1_DataWidth_reg[1]/NET0131  & ~n8664 ;
  assign n12317 = ~n7913 & ~n8709 ;
  assign n12318 = \P1_P1_InstQueue_reg[9][3]/NET0131  & ~n4327 ;
  assign n12319 = ~n8139 & n12318 ;
  assign n12320 = ~n12317 & ~n12319 ;
  assign n12321 = ~n12316 & ~n12320 ;
  assign n12322 = ~n12315 & ~n12321 ;
  assign n12323 = n8282 & ~n12322 ;
  assign n12324 = n8287 & ~n12320 ;
  assign n12311 = \P1_P1_InstQueue_reg[9][3]/NET0131  & ~n8366 ;
  assign n12325 = n4327 & ~n10096 ;
  assign n12326 = ~n12318 & ~n12325 ;
  assign n12327 = n8350 & ~n12326 ;
  assign n12328 = ~n12311 & ~n12327 ;
  assign n12329 = ~n12324 & n12328 ;
  assign n12330 = ~n12323 & n12329 ;
  assign n12335 = ~n11372 & n11582 ;
  assign n12336 = n11372 & ~n11582 ;
  assign n12337 = ~n12335 & ~n12336 ;
  assign n12338 = ~n10105 & ~n12337 ;
  assign n12331 = ~n11521 & n11537 ;
  assign n12332 = ~n11538 & ~n12331 ;
  assign n12333 = n10105 & ~n12332 ;
  assign n12334 = n11593 & n11609 ;
  assign n12339 = ~n12333 & n12334 ;
  assign n12340 = ~n12338 & n12339 ;
  assign n12353 = \P2_P1_InstQueue_reg[6][4]/NET0131  & n11651 ;
  assign n12352 = \P2_P1_InstQueue_reg[15][4]/NET0131  & n11647 ;
  assign n12348 = \P2_P1_InstQueue_reg[5][4]/NET0131  & n11638 ;
  assign n12349 = \P2_P1_InstQueue_reg[0][4]/NET0131  & n11669 ;
  assign n12364 = ~n12348 & ~n12349 ;
  assign n12374 = ~n12352 & n12364 ;
  assign n12375 = ~n12353 & n12374 ;
  assign n12360 = \P2_P1_InstQueue_reg[8][4]/NET0131  & n11659 ;
  assign n12361 = \P2_P1_InstQueue_reg[11][4]/NET0131  & n11665 ;
  assign n12369 = ~n12360 & ~n12361 ;
  assign n12362 = \P2_P1_InstQueue_reg[3][4]/NET0131  & n11663 ;
  assign n12363 = \P2_P1_InstQueue_reg[9][4]/NET0131  & n11656 ;
  assign n12370 = ~n12362 & ~n12363 ;
  assign n12371 = n12369 & n12370 ;
  assign n12356 = \P2_P1_InstQueue_reg[4][4]/NET0131  & n11667 ;
  assign n12357 = \P2_P1_InstQueue_reg[7][4]/NET0131  & n11661 ;
  assign n12367 = ~n12356 & ~n12357 ;
  assign n12358 = \P2_P1_InstQueue_reg[12][4]/NET0131  & n11673 ;
  assign n12359 = \P2_P1_InstQueue_reg[13][4]/NET0131  & n11641 ;
  assign n12368 = ~n12358 & ~n12359 ;
  assign n12372 = n12367 & n12368 ;
  assign n12350 = \P2_P1_InstQueue_reg[10][4]/NET0131  & n11634 ;
  assign n12351 = \P2_P1_InstQueue_reg[14][4]/NET0131  & n11643 ;
  assign n12365 = ~n12350 & ~n12351 ;
  assign n12354 = \P2_P1_InstQueue_reg[1][4]/NET0131  & n11671 ;
  assign n12355 = \P2_P1_InstQueue_reg[2][4]/NET0131  & n11654 ;
  assign n12366 = ~n12354 & ~n12355 ;
  assign n12373 = n12365 & n12366 ;
  assign n12376 = n12372 & n12373 ;
  assign n12377 = n12371 & n12376 ;
  assign n12378 = n12375 & n12377 ;
  assign n12379 = n11596 & n12378 ;
  assign n12347 = ~\P2_P1_InstQueue_reg[11][4]/NET0131  & ~n11596 ;
  assign n12380 = n11692 & ~n12347 ;
  assign n12381 = ~n12379 & n12380 ;
  assign n12341 = ~n11609 & ~n11613 ;
  assign n12342 = n11593 & ~n11613 ;
  assign n12343 = ~n12341 & ~n12342 ;
  assign n12344 = n11600 & n12343 ;
  assign n12345 = n11630 & ~n12344 ;
  assign n12346 = \P2_P1_InstQueue_reg[11][4]/NET0131  & ~n12345 ;
  assign n12382 = n11376 & ~n11600 ;
  assign n12383 = n12343 & n12382 ;
  assign n12384 = ~n12346 & ~n12383 ;
  assign n12385 = ~n12381 & n12384 ;
  assign n12386 = ~n12340 & n12385 ;
  assign n12389 = ~n11862 & ~n12337 ;
  assign n12387 = n11862 & ~n12332 ;
  assign n12388 = n11609 & n11870 ;
  assign n12390 = ~n12387 & n12388 ;
  assign n12391 = ~n12389 & n12390 ;
  assign n12398 = n11871 & n12378 ;
  assign n12397 = ~\P2_P1_InstQueue_reg[0][4]/NET0131  & ~n11871 ;
  assign n12399 = n11692 & ~n12397 ;
  assign n12400 = ~n12398 & n12399 ;
  assign n12392 = ~n11613 & n11870 ;
  assign n12393 = ~n12341 & ~n12392 ;
  assign n12394 = n11874 & n12393 ;
  assign n12395 = n11630 & ~n12394 ;
  assign n12396 = \P2_P1_InstQueue_reg[0][4]/NET0131  & ~n12395 ;
  assign n12401 = n11376 & ~n11874 ;
  assign n12402 = n12393 & n12401 ;
  assign n12403 = ~n12396 & ~n12402 ;
  assign n12404 = ~n12400 & n12403 ;
  assign n12405 = ~n12391 & n12404 ;
  assign n12408 = ~n11891 & ~n12337 ;
  assign n12406 = n11891 & ~n12332 ;
  assign n12407 = n11609 & n11896 ;
  assign n12409 = ~n12406 & n12407 ;
  assign n12410 = ~n12408 & n12409 ;
  assign n12417 = n11599 & n12378 ;
  assign n12416 = ~\P2_P1_InstQueue_reg[10][4]/NET0131  & ~n11599 ;
  assign n12418 = n11692 & ~n12416 ;
  assign n12419 = ~n12417 & n12418 ;
  assign n12411 = ~n11613 & n11896 ;
  assign n12412 = ~n12341 & ~n12411 ;
  assign n12413 = n11897 & n12412 ;
  assign n12414 = n11630 & ~n12413 ;
  assign n12415 = \P2_P1_InstQueue_reg[10][4]/NET0131  & ~n12414 ;
  assign n12420 = n11376 & ~n11897 ;
  assign n12421 = n12412 & n12420 ;
  assign n12422 = ~n12415 & ~n12421 ;
  assign n12423 = ~n12419 & n12422 ;
  assign n12424 = ~n12410 & n12423 ;
  assign n12427 = ~n11577 & ~n12337 ;
  assign n12425 = n11577 & ~n12332 ;
  assign n12426 = n11609 & n11917 ;
  assign n12428 = ~n12425 & n12426 ;
  assign n12429 = ~n12427 & n12428 ;
  assign n12436 = n11919 & n12378 ;
  assign n12435 = ~\P2_P1_InstQueue_reg[12][4]/NET0131  & ~n11919 ;
  assign n12437 = n11692 & ~n12435 ;
  assign n12438 = ~n12436 & n12437 ;
  assign n12430 = ~n11613 & n11917 ;
  assign n12431 = ~n12341 & ~n12430 ;
  assign n12432 = n11920 & n12431 ;
  assign n12433 = n11630 & ~n12432 ;
  assign n12434 = \P2_P1_InstQueue_reg[12][4]/NET0131  & ~n12433 ;
  assign n12439 = n11376 & ~n11920 ;
  assign n12440 = n12431 & n12439 ;
  assign n12441 = ~n12434 & ~n12440 ;
  assign n12442 = ~n12438 & n12441 ;
  assign n12443 = ~n12429 & n12442 ;
  assign n12446 = ~n11599 & ~n12337 ;
  assign n12444 = n11599 & ~n12332 ;
  assign n12445 = n11609 & n11960 ;
  assign n12447 = ~n12444 & n12445 ;
  assign n12448 = ~n12446 & n12447 ;
  assign n12455 = n11862 & n12378 ;
  assign n12454 = ~\P2_P1_InstQueue_reg[13][4]/NET0131  & ~n11862 ;
  assign n12456 = n11692 & ~n12454 ;
  assign n12457 = ~n12455 & n12456 ;
  assign n12449 = ~n11613 & n11960 ;
  assign n12450 = ~n12341 & ~n12449 ;
  assign n12451 = n11961 & n12450 ;
  assign n12452 = n11630 & ~n12451 ;
  assign n12453 = \P2_P1_InstQueue_reg[13][4]/NET0131  & ~n12452 ;
  assign n12458 = n11376 & ~n11961 ;
  assign n12459 = n12450 & n12458 ;
  assign n12460 = ~n12453 & ~n12459 ;
  assign n12461 = ~n12457 & n12460 ;
  assign n12462 = ~n12448 & n12461 ;
  assign n12465 = ~n11596 & ~n12337 ;
  assign n12463 = n11596 & ~n12332 ;
  assign n12464 = n11609 & n11981 ;
  assign n12466 = ~n12463 & n12464 ;
  assign n12467 = ~n12465 & n12466 ;
  assign n12474 = n11865 & n12378 ;
  assign n12473 = ~\P2_P1_InstQueue_reg[14][4]/NET0131  & ~n11865 ;
  assign n12475 = n11692 & ~n12473 ;
  assign n12476 = ~n12474 & n12475 ;
  assign n12468 = ~n11613 & n11981 ;
  assign n12469 = ~n12341 & ~n12468 ;
  assign n12470 = n11869 & n12469 ;
  assign n12471 = n11630 & ~n12470 ;
  assign n12472 = \P2_P1_InstQueue_reg[14][4]/NET0131  & ~n12471 ;
  assign n12477 = n11376 & ~n11869 ;
  assign n12478 = n12469 & n12477 ;
  assign n12479 = ~n12472 & ~n12478 ;
  assign n12480 = ~n12476 & n12479 ;
  assign n12481 = ~n12467 & n12480 ;
  assign n12484 = ~n11919 & ~n12337 ;
  assign n12482 = n11919 & ~n12332 ;
  assign n12483 = n11609 & n12001 ;
  assign n12485 = ~n12482 & n12483 ;
  assign n12486 = ~n12484 & n12485 ;
  assign n12493 = n11873 & n12378 ;
  assign n12492 = ~\P2_P1_InstQueue_reg[15][4]/NET0131  & ~n11873 ;
  assign n12494 = n11692 & ~n12492 ;
  assign n12495 = ~n12493 & n12494 ;
  assign n12487 = ~n11613 & n12001 ;
  assign n12488 = ~n12341 & ~n12487 ;
  assign n12489 = n12002 & n12488 ;
  assign n12490 = n11630 & ~n12489 ;
  assign n12491 = \P2_P1_InstQueue_reg[15][4]/NET0131  & ~n12490 ;
  assign n12496 = n11376 & ~n12002 ;
  assign n12497 = n12488 & n12496 ;
  assign n12498 = ~n12491 & ~n12497 ;
  assign n12499 = ~n12495 & n12498 ;
  assign n12500 = ~n12486 & n12499 ;
  assign n12503 = ~n11865 & ~n12337 ;
  assign n12501 = n11865 & ~n12332 ;
  assign n12502 = n11609 & n12022 ;
  assign n12504 = ~n12501 & n12502 ;
  assign n12505 = ~n12503 & n12504 ;
  assign n12512 = n12023 & n12378 ;
  assign n12511 = ~\P2_P1_InstQueue_reg[1][4]/NET0131  & ~n12023 ;
  assign n12513 = n11692 & ~n12511 ;
  assign n12514 = ~n12512 & n12513 ;
  assign n12506 = ~n11613 & n12022 ;
  assign n12507 = ~n12341 & ~n12506 ;
  assign n12508 = n12024 & n12507 ;
  assign n12509 = n11630 & ~n12508 ;
  assign n12510 = \P2_P1_InstQueue_reg[1][4]/NET0131  & ~n12509 ;
  assign n12515 = n11376 & ~n12024 ;
  assign n12516 = n12507 & n12515 ;
  assign n12517 = ~n12510 & ~n12516 ;
  assign n12518 = ~n12514 & n12517 ;
  assign n12519 = ~n12505 & n12518 ;
  assign n12522 = ~n11873 & ~n12337 ;
  assign n12520 = n11873 & ~n12332 ;
  assign n12521 = n11609 & n12064 ;
  assign n12523 = ~n12520 & n12521 ;
  assign n12524 = ~n12522 & n12523 ;
  assign n12531 = n12065 & n12378 ;
  assign n12530 = ~\P2_P1_InstQueue_reg[2][4]/NET0131  & ~n12065 ;
  assign n12532 = n11692 & ~n12530 ;
  assign n12533 = ~n12531 & n12532 ;
  assign n12525 = ~n11613 & n12064 ;
  assign n12526 = ~n12341 & ~n12525 ;
  assign n12527 = n12066 & n12526 ;
  assign n12528 = n11630 & ~n12527 ;
  assign n12529 = \P2_P1_InstQueue_reg[2][4]/NET0131  & ~n12528 ;
  assign n12534 = n11376 & ~n12066 ;
  assign n12535 = n12526 & n12534 ;
  assign n12536 = ~n12529 & ~n12535 ;
  assign n12537 = ~n12533 & n12536 ;
  assign n12538 = ~n12524 & n12537 ;
  assign n12541 = ~n11871 & ~n12337 ;
  assign n12539 = n11871 & ~n12332 ;
  assign n12540 = n11609 & n12086 ;
  assign n12542 = ~n12539 & n12540 ;
  assign n12543 = ~n12541 & n12542 ;
  assign n12550 = n12087 & n12378 ;
  assign n12549 = ~\P2_P1_InstQueue_reg[3][4]/NET0131  & ~n12087 ;
  assign n12551 = n11692 & ~n12549 ;
  assign n12552 = ~n12550 & n12551 ;
  assign n12544 = ~n11613 & n12086 ;
  assign n12545 = ~n12341 & ~n12544 ;
  assign n12546 = n12088 & n12545 ;
  assign n12547 = n11630 & ~n12546 ;
  assign n12548 = \P2_P1_InstQueue_reg[3][4]/NET0131  & ~n12547 ;
  assign n12553 = n11376 & ~n12088 ;
  assign n12554 = n12545 & n12553 ;
  assign n12555 = ~n12548 & ~n12554 ;
  assign n12556 = ~n12552 & n12555 ;
  assign n12557 = ~n12543 & n12556 ;
  assign n12560 = ~n12023 & ~n12337 ;
  assign n12558 = n12023 & ~n12332 ;
  assign n12559 = n11609 & n12108 ;
  assign n12561 = ~n12558 & n12559 ;
  assign n12562 = ~n12560 & n12561 ;
  assign n12569 = n12109 & n12378 ;
  assign n12568 = ~\P2_P1_InstQueue_reg[4][4]/NET0131  & ~n12109 ;
  assign n12570 = n11692 & ~n12568 ;
  assign n12571 = ~n12569 & n12570 ;
  assign n12563 = ~n11613 & n12108 ;
  assign n12564 = ~n12341 & ~n12563 ;
  assign n12565 = n12110 & n12564 ;
  assign n12566 = n11630 & ~n12565 ;
  assign n12567 = \P2_P1_InstQueue_reg[4][4]/NET0131  & ~n12566 ;
  assign n12572 = n11376 & ~n12110 ;
  assign n12573 = n12564 & n12572 ;
  assign n12574 = ~n12567 & ~n12573 ;
  assign n12575 = ~n12571 & n12574 ;
  assign n12576 = ~n12562 & n12575 ;
  assign n12579 = ~n12065 & ~n12337 ;
  assign n12577 = n12065 & ~n12332 ;
  assign n12578 = n11609 & n12130 ;
  assign n12580 = ~n12577 & n12578 ;
  assign n12581 = ~n12579 & n12580 ;
  assign n12588 = n12131 & n12378 ;
  assign n12587 = ~\P2_P1_InstQueue_reg[5][4]/NET0131  & ~n12131 ;
  assign n12589 = n11692 & ~n12587 ;
  assign n12590 = ~n12588 & n12589 ;
  assign n12582 = ~n11613 & n12130 ;
  assign n12583 = ~n12341 & ~n12582 ;
  assign n12584 = n12132 & n12583 ;
  assign n12585 = n11630 & ~n12584 ;
  assign n12586 = \P2_P1_InstQueue_reg[5][4]/NET0131  & ~n12585 ;
  assign n12591 = n11376 & ~n12132 ;
  assign n12592 = n12583 & n12591 ;
  assign n12593 = ~n12586 & ~n12592 ;
  assign n12594 = ~n12590 & n12593 ;
  assign n12595 = ~n12581 & n12594 ;
  assign n12598 = ~n12087 & ~n12337 ;
  assign n12596 = n12087 & ~n12332 ;
  assign n12597 = n11609 & n12172 ;
  assign n12599 = ~n12596 & n12597 ;
  assign n12600 = ~n12598 & n12599 ;
  assign n12607 = n12173 & n12378 ;
  assign n12606 = ~\P2_P1_InstQueue_reg[6][4]/NET0131  & ~n12173 ;
  assign n12608 = n11692 & ~n12606 ;
  assign n12609 = ~n12607 & n12608 ;
  assign n12601 = ~n11613 & n12172 ;
  assign n12602 = ~n12341 & ~n12601 ;
  assign n12603 = n12174 & n12602 ;
  assign n12604 = n11630 & ~n12603 ;
  assign n12605 = \P2_P1_InstQueue_reg[6][4]/NET0131  & ~n12604 ;
  assign n12610 = n11376 & ~n12174 ;
  assign n12611 = n12602 & n12610 ;
  assign n12612 = ~n12605 & ~n12611 ;
  assign n12613 = ~n12609 & n12612 ;
  assign n12614 = ~n12600 & n12613 ;
  assign n12617 = ~n12109 & ~n12337 ;
  assign n12615 = n12109 & ~n12332 ;
  assign n12616 = n11609 & n12194 ;
  assign n12618 = ~n12615 & n12616 ;
  assign n12619 = ~n12617 & n12618 ;
  assign n12626 = n11891 & n12378 ;
  assign n12625 = ~\P2_P1_InstQueue_reg[7][4]/NET0131  & ~n11891 ;
  assign n12627 = n11692 & ~n12625 ;
  assign n12628 = ~n12626 & n12627 ;
  assign n12620 = ~n11613 & n12194 ;
  assign n12621 = ~n12341 & ~n12620 ;
  assign n12622 = n12195 & n12621 ;
  assign n12623 = n11630 & ~n12622 ;
  assign n12624 = \P2_P1_InstQueue_reg[7][4]/NET0131  & ~n12623 ;
  assign n12629 = n11376 & ~n12195 ;
  assign n12630 = n12621 & n12629 ;
  assign n12631 = ~n12624 & ~n12630 ;
  assign n12632 = ~n12628 & n12631 ;
  assign n12633 = ~n12619 & n12632 ;
  assign n12636 = ~n12131 & ~n12337 ;
  assign n12634 = n12131 & ~n12332 ;
  assign n12635 = n11609 & n12215 ;
  assign n12637 = ~n12634 & n12635 ;
  assign n12638 = ~n12636 & n12637 ;
  assign n12645 = n10105 & n12378 ;
  assign n12644 = ~\P2_P1_InstQueue_reg[8][4]/NET0131  & ~n10105 ;
  assign n12646 = n11692 & ~n12644 ;
  assign n12647 = ~n12645 & n12646 ;
  assign n12639 = ~n11613 & n12215 ;
  assign n12640 = ~n12341 & ~n12639 ;
  assign n12641 = n11895 & n12640 ;
  assign n12642 = n11630 & ~n12641 ;
  assign n12643 = \P2_P1_InstQueue_reg[8][4]/NET0131  & ~n12642 ;
  assign n12648 = n11376 & ~n11895 ;
  assign n12649 = n12640 & n12648 ;
  assign n12650 = ~n12643 & ~n12649 ;
  assign n12651 = ~n12647 & n12650 ;
  assign n12652 = ~n12638 & n12651 ;
  assign n12655 = ~n12173 & ~n12337 ;
  assign n12653 = n12173 & ~n12332 ;
  assign n12654 = n11609 & n12235 ;
  assign n12656 = ~n12653 & n12654 ;
  assign n12657 = ~n12655 & n12656 ;
  assign n12664 = n11577 & n12378 ;
  assign n12663 = ~\P2_P1_InstQueue_reg[9][4]/NET0131  & ~n11577 ;
  assign n12665 = n11692 & ~n12663 ;
  assign n12666 = ~n12664 & n12665 ;
  assign n12658 = ~n11613 & n12235 ;
  assign n12659 = ~n12341 & ~n12658 ;
  assign n12660 = n11592 & n12659 ;
  assign n12661 = n11630 & ~n12660 ;
  assign n12662 = \P2_P1_InstQueue_reg[9][4]/NET0131  & ~n12661 ;
  assign n12667 = n11376 & ~n11592 ;
  assign n12668 = n12659 & n12667 ;
  assign n12669 = ~n12662 & ~n12668 ;
  assign n12670 = ~n12666 & n12669 ;
  assign n12671 = ~n12657 & n12670 ;
  assign n12678 = ~n8191 & n8206 ;
  assign n12679 = ~n8207 & ~n12678 ;
  assign n12680 = n8139 & ~n12679 ;
  assign n12681 = ~n8053 & n8068 ;
  assign n12682 = ~n8069 & ~n12681 ;
  assign n12683 = ~n8139 & ~n12682 ;
  assign n12684 = ~n12680 & ~n12683 ;
  assign n12685 = n10057 & ~n12684 ;
  assign n12672 = n7947 & ~n8146 ;
  assign n12673 = \P1_P1_InstQueue_reg[11][2]/NET0131  & ~n8142 ;
  assign n12674 = ~n8145 & n12673 ;
  assign n12675 = ~n12672 & ~n12674 ;
  assign n12677 = ~n10057 & n12675 ;
  assign n12686 = n8282 & ~n12677 ;
  assign n12687 = ~n12685 & n12686 ;
  assign n12676 = n8287 & ~n12675 ;
  assign n12688 = \P1_P1_InstQueue_reg[14][2]/NET0131  & n8291 ;
  assign n12689 = \P1_P1_InstQueue_reg[2][2]/NET0131  & n8314 ;
  assign n12690 = \P1_P1_InstQueue_reg[13][2]/NET0131  & n8327 ;
  assign n12704 = ~n12689 & ~n12690 ;
  assign n12691 = \P1_P1_InstQueue_reg[11][2]/NET0131  & n8312 ;
  assign n12692 = \P1_P1_InstQueue_reg[3][2]/NET0131  & n8323 ;
  assign n12705 = ~n12691 & ~n12692 ;
  assign n12714 = n12704 & n12705 ;
  assign n12715 = ~n12688 & n12714 ;
  assign n12703 = \P1_P1_InstQueue_reg[9][2]/NET0131  & n8325 ;
  assign n12701 = \P1_P1_InstQueue_reg[1][2]/NET0131  & n8299 ;
  assign n12702 = \P1_P1_InstQueue_reg[4][2]/NET0131  & n8295 ;
  assign n12710 = ~n12701 & ~n12702 ;
  assign n12711 = ~n12703 & n12710 ;
  assign n12697 = \P1_P1_InstQueue_reg[6][2]/NET0131  & n8316 ;
  assign n12698 = \P1_P1_InstQueue_reg[15][2]/NET0131  & n8321 ;
  assign n12708 = ~n12697 & ~n12698 ;
  assign n12699 = \P1_P1_InstQueue_reg[7][2]/NET0131  & n8318 ;
  assign n12700 = \P1_P1_InstQueue_reg[10][2]/NET0131  & n8303 ;
  assign n12709 = ~n12699 & ~n12700 ;
  assign n12712 = n12708 & n12709 ;
  assign n12693 = \P1_P1_InstQueue_reg[8][2]/NET0131  & n8305 ;
  assign n12694 = \P1_P1_InstQueue_reg[0][2]/NET0131  & n8309 ;
  assign n12706 = ~n12693 & ~n12694 ;
  assign n12695 = \P1_P1_InstQueue_reg[12][2]/NET0131  & n8329 ;
  assign n12696 = \P1_P1_InstQueue_reg[5][2]/NET0131  & n8307 ;
  assign n12707 = ~n12695 & ~n12696 ;
  assign n12713 = n12706 & n12707 ;
  assign n12716 = n12712 & n12713 ;
  assign n12717 = n12711 & n12716 ;
  assign n12718 = n12715 & n12717 ;
  assign n12719 = n8142 & ~n12718 ;
  assign n12720 = ~n12673 & ~n12719 ;
  assign n12721 = n8350 & ~n12720 ;
  assign n12722 = \P1_P1_InstQueue_reg[11][2]/NET0131  & ~n8366 ;
  assign n12723 = ~n12721 & ~n12722 ;
  assign n12724 = ~n12676 & n12723 ;
  assign n12725 = ~n12687 & n12724 ;
  assign n12729 = ~n11505 & n11520 ;
  assign n12730 = ~n11521 & ~n12729 ;
  assign n12731 = n10105 & ~n12730 ;
  assign n12726 = ~n11343 & ~n11581 ;
  assign n12727 = ~n11582 & ~n12726 ;
  assign n12728 = ~n10105 & ~n12727 ;
  assign n12732 = n12334 & ~n12728 ;
  assign n12733 = ~n12731 & n12732 ;
  assign n12741 = \P2_P1_InstQueue_reg[6][3]/NET0131  & n11651 ;
  assign n12740 = \P2_P1_InstQueue_reg[15][3]/NET0131  & n11647 ;
  assign n12736 = \P2_P1_InstQueue_reg[4][3]/NET0131  & n11667 ;
  assign n12737 = \P2_P1_InstQueue_reg[2][3]/NET0131  & n11654 ;
  assign n12752 = ~n12736 & ~n12737 ;
  assign n12762 = ~n12740 & n12752 ;
  assign n12763 = ~n12741 & n12762 ;
  assign n12748 = \P2_P1_InstQueue_reg[11][3]/NET0131  & n11665 ;
  assign n12749 = \P2_P1_InstQueue_reg[12][3]/NET0131  & n11673 ;
  assign n12757 = ~n12748 & ~n12749 ;
  assign n12750 = \P2_P1_InstQueue_reg[1][3]/NET0131  & n11671 ;
  assign n12751 = \P2_P1_InstQueue_reg[10][3]/NET0131  & n11634 ;
  assign n12758 = ~n12750 & ~n12751 ;
  assign n12759 = n12757 & n12758 ;
  assign n12744 = \P2_P1_InstQueue_reg[3][3]/NET0131  & n11663 ;
  assign n12745 = \P2_P1_InstQueue_reg[7][3]/NET0131  & n11661 ;
  assign n12755 = ~n12744 & ~n12745 ;
  assign n12746 = \P2_P1_InstQueue_reg[13][3]/NET0131  & n11641 ;
  assign n12747 = \P2_P1_InstQueue_reg[5][3]/NET0131  & n11638 ;
  assign n12756 = ~n12746 & ~n12747 ;
  assign n12760 = n12755 & n12756 ;
  assign n12738 = \P2_P1_InstQueue_reg[0][3]/NET0131  & n11669 ;
  assign n12739 = \P2_P1_InstQueue_reg[14][3]/NET0131  & n11643 ;
  assign n12753 = ~n12738 & ~n12739 ;
  assign n12742 = \P2_P1_InstQueue_reg[8][3]/NET0131  & n11659 ;
  assign n12743 = \P2_P1_InstQueue_reg[9][3]/NET0131  & n11656 ;
  assign n12754 = ~n12742 & ~n12743 ;
  assign n12761 = n12753 & n12754 ;
  assign n12764 = n12760 & n12761 ;
  assign n12765 = n12759 & n12764 ;
  assign n12766 = n12763 & n12765 ;
  assign n12767 = n11596 & n12766 ;
  assign n12735 = ~\P2_P1_InstQueue_reg[11][3]/NET0131  & ~n11596 ;
  assign n12768 = n11692 & ~n12735 ;
  assign n12769 = ~n12767 & n12768 ;
  assign n12734 = \P2_P1_InstQueue_reg[11][3]/NET0131  & ~n12345 ;
  assign n12770 = n11374 & ~n11600 ;
  assign n12771 = n12343 & n12770 ;
  assign n12772 = ~n12734 & ~n12771 ;
  assign n12773 = ~n12769 & n12772 ;
  assign n12774 = ~n12733 & n12773 ;
  assign n12816 = ~n11554 & n11569 ;
  assign n12817 = ~n11570 & ~n12816 ;
  assign n12818 = n10105 & ~n12817 ;
  assign n12819 = n11342 & ~n11584 ;
  assign n12820 = ~n11585 & ~n12819 ;
  assign n12821 = ~n10105 & ~n12820 ;
  assign n12822 = ~n12818 & ~n12821 ;
  assign n12823 = n11593 & ~n12822 ;
  assign n12811 = n11383 & ~n11600 ;
  assign n12776 = \P2_P1_InstQueue_reg[11][6]/NET0131  & ~n11596 ;
  assign n12812 = ~n11599 & n12776 ;
  assign n12813 = ~n12811 & ~n12812 ;
  assign n12815 = ~n11593 & n12813 ;
  assign n12824 = n11609 & ~n12815 ;
  assign n12825 = ~n12823 & n12824 ;
  assign n12782 = \P2_P1_InstQueue_reg[6][6]/NET0131  & n11651 ;
  assign n12781 = \P2_P1_InstQueue_reg[15][6]/NET0131  & n11647 ;
  assign n12777 = \P2_P1_InstQueue_reg[10][6]/NET0131  & n11634 ;
  assign n12778 = \P2_P1_InstQueue_reg[5][6]/NET0131  & n11638 ;
  assign n12793 = ~n12777 & ~n12778 ;
  assign n12803 = ~n12781 & n12793 ;
  assign n12804 = ~n12782 & n12803 ;
  assign n12789 = \P2_P1_InstQueue_reg[13][6]/NET0131  & n11641 ;
  assign n12790 = \P2_P1_InstQueue_reg[11][6]/NET0131  & n11665 ;
  assign n12798 = ~n12789 & ~n12790 ;
  assign n12791 = \P2_P1_InstQueue_reg[1][6]/NET0131  & n11671 ;
  assign n12792 = \P2_P1_InstQueue_reg[12][6]/NET0131  & n11673 ;
  assign n12799 = ~n12791 & ~n12792 ;
  assign n12800 = n12798 & n12799 ;
  assign n12785 = \P2_P1_InstQueue_reg[8][6]/NET0131  & n11659 ;
  assign n12786 = \P2_P1_InstQueue_reg[7][6]/NET0131  & n11661 ;
  assign n12796 = ~n12785 & ~n12786 ;
  assign n12787 = \P2_P1_InstQueue_reg[0][6]/NET0131  & n11669 ;
  assign n12788 = \P2_P1_InstQueue_reg[2][6]/NET0131  & n11654 ;
  assign n12797 = ~n12787 & ~n12788 ;
  assign n12801 = n12796 & n12797 ;
  assign n12779 = \P2_P1_InstQueue_reg[4][6]/NET0131  & n11667 ;
  assign n12780 = \P2_P1_InstQueue_reg[14][6]/NET0131  & n11643 ;
  assign n12794 = ~n12779 & ~n12780 ;
  assign n12783 = \P2_P1_InstQueue_reg[3][6]/NET0131  & n11663 ;
  assign n12784 = \P2_P1_InstQueue_reg[9][6]/NET0131  & n11656 ;
  assign n12795 = ~n12783 & ~n12784 ;
  assign n12802 = n12794 & n12795 ;
  assign n12805 = n12801 & n12802 ;
  assign n12806 = n12800 & n12805 ;
  assign n12807 = n12804 & n12806 ;
  assign n12808 = n11596 & ~n12807 ;
  assign n12809 = ~n12776 & ~n12808 ;
  assign n12810 = n11692 & ~n12809 ;
  assign n12775 = \P2_P1_InstQueue_reg[11][6]/NET0131  & ~n11630 ;
  assign n12814 = n11613 & ~n12813 ;
  assign n12826 = ~n12775 & ~n12814 ;
  assign n12827 = ~n12810 & n12826 ;
  assign n12828 = ~n12825 & n12827 ;
  assign n12835 = n8375 & ~n12679 ;
  assign n12836 = ~n8375 & ~n12682 ;
  assign n12837 = ~n12835 & ~n12836 ;
  assign n12838 = n11707 & ~n12837 ;
  assign n12829 = n7947 & ~n8379 ;
  assign n12830 = \P1_P1_InstQueue_reg[0][2]/NET0131  & ~n8376 ;
  assign n12831 = ~n8378 & n12830 ;
  assign n12832 = ~n12829 & ~n12831 ;
  assign n12834 = ~n11707 & n12832 ;
  assign n12839 = n8282 & ~n12834 ;
  assign n12840 = ~n12838 & n12839 ;
  assign n12833 = n8287 & ~n12832 ;
  assign n12841 = n8376 & ~n12718 ;
  assign n12842 = ~n12830 & ~n12841 ;
  assign n12843 = n8350 & ~n12842 ;
  assign n12844 = \P1_P1_InstQueue_reg[0][2]/NET0131  & ~n8366 ;
  assign n12845 = ~n12843 & ~n12844 ;
  assign n12846 = ~n12833 & n12845 ;
  assign n12847 = ~n12840 & n12846 ;
  assign n12854 = n8407 & ~n12679 ;
  assign n12855 = ~n8407 & ~n12682 ;
  assign n12856 = ~n12854 & ~n12855 ;
  assign n12857 = n9418 & ~n12856 ;
  assign n12848 = n7947 & ~n8401 ;
  assign n12849 = \P1_P1_InstQueue_reg[10][2]/NET0131  & ~n8145 ;
  assign n12850 = ~n4327 & n12849 ;
  assign n12851 = ~n12848 & ~n12850 ;
  assign n12853 = ~n9418 & n12851 ;
  assign n12858 = n8282 & ~n12853 ;
  assign n12859 = ~n12857 & n12858 ;
  assign n12852 = n8287 & ~n12851 ;
  assign n12860 = n8145 & ~n12718 ;
  assign n12861 = ~n12849 & ~n12860 ;
  assign n12862 = n8350 & ~n12861 ;
  assign n12863 = \P1_P1_InstQueue_reg[10][2]/NET0131  & ~n8366 ;
  assign n12864 = ~n12862 & ~n12863 ;
  assign n12865 = ~n12852 & n12864 ;
  assign n12866 = ~n12859 & n12865 ;
  assign n12873 = n4327 & ~n12679 ;
  assign n12874 = ~n4327 & ~n12682 ;
  assign n12875 = ~n12873 & ~n12874 ;
  assign n12876 = n11746 & ~n12875 ;
  assign n12867 = n7947 & ~n8428 ;
  assign n12868 = \P1_P1_InstQueue_reg[12][2]/NET0131  & ~n8427 ;
  assign n12869 = ~n8142 & n12868 ;
  assign n12870 = ~n12867 & ~n12869 ;
  assign n12872 = ~n11746 & n12870 ;
  assign n12877 = n8282 & ~n12872 ;
  assign n12878 = ~n12876 & n12877 ;
  assign n12871 = n8287 & ~n12870 ;
  assign n12879 = n8427 & ~n12718 ;
  assign n12880 = ~n12868 & ~n12879 ;
  assign n12881 = n8350 & ~n12880 ;
  assign n12882 = \P1_P1_InstQueue_reg[12][2]/NET0131  & ~n8366 ;
  assign n12883 = ~n12881 & ~n12882 ;
  assign n12884 = ~n12871 & n12883 ;
  assign n12885 = ~n12878 & n12884 ;
  assign n12892 = n8145 & ~n12679 ;
  assign n12893 = ~n8145 & ~n12682 ;
  assign n12894 = ~n12892 & ~n12893 ;
  assign n12895 = n11766 & ~n12894 ;
  assign n12886 = n7947 & ~n8451 ;
  assign n12887 = \P1_P1_InstQueue_reg[13][2]/NET0131  & ~n8375 ;
  assign n12888 = ~n8427 & n12887 ;
  assign n12889 = ~n12886 & ~n12888 ;
  assign n12891 = ~n11766 & n12889 ;
  assign n12896 = n8282 & ~n12891 ;
  assign n12897 = ~n12895 & n12896 ;
  assign n12890 = n8287 & ~n12889 ;
  assign n12898 = n8375 & ~n12718 ;
  assign n12899 = ~n12887 & ~n12898 ;
  assign n12900 = n8350 & ~n12899 ;
  assign n12901 = \P1_P1_InstQueue_reg[13][2]/NET0131  & ~n8366 ;
  assign n12902 = ~n12900 & ~n12901 ;
  assign n12903 = ~n12890 & n12902 ;
  assign n12904 = ~n12897 & n12903 ;
  assign n12911 = n8142 & ~n12679 ;
  assign n12912 = ~n8142 & ~n12682 ;
  assign n12913 = ~n12911 & ~n12912 ;
  assign n12914 = n11786 & ~n12913 ;
  assign n12905 = n7947 & ~n8474 ;
  assign n12906 = \P1_P1_InstQueue_reg[14][2]/NET0131  & ~n8372 ;
  assign n12907 = ~n8375 & n12906 ;
  assign n12908 = ~n12905 & ~n12907 ;
  assign n12910 = ~n11786 & n12908 ;
  assign n12915 = n8282 & ~n12910 ;
  assign n12916 = ~n12914 & n12915 ;
  assign n12909 = n8287 & ~n12908 ;
  assign n12917 = n8372 & ~n12718 ;
  assign n12918 = ~n12906 & ~n12917 ;
  assign n12919 = n8350 & ~n12918 ;
  assign n12920 = \P1_P1_InstQueue_reg[14][2]/NET0131  & ~n8366 ;
  assign n12921 = ~n12919 & ~n12920 ;
  assign n12922 = ~n12909 & n12921 ;
  assign n12923 = ~n12916 & n12922 ;
  assign n12930 = n8427 & ~n12679 ;
  assign n12931 = ~n8427 & ~n12682 ;
  assign n12932 = ~n12930 & ~n12931 ;
  assign n12933 = n11806 & ~n12932 ;
  assign n12924 = n7947 & ~n8497 ;
  assign n12925 = \P1_P1_InstQueue_reg[15][2]/NET0131  & ~n8378 ;
  assign n12926 = ~n8372 & n12925 ;
  assign n12927 = ~n12924 & ~n12926 ;
  assign n12929 = ~n11806 & n12927 ;
  assign n12934 = n8282 & ~n12929 ;
  assign n12935 = ~n12933 & n12934 ;
  assign n12928 = n8287 & ~n12927 ;
  assign n12936 = n8378 & ~n12718 ;
  assign n12937 = ~n12925 & ~n12936 ;
  assign n12938 = n8350 & ~n12937 ;
  assign n12939 = \P1_P1_InstQueue_reg[15][2]/NET0131  & ~n8366 ;
  assign n12940 = ~n12938 & ~n12939 ;
  assign n12941 = ~n12928 & n12940 ;
  assign n12942 = ~n12935 & n12941 ;
  assign n12949 = n8372 & ~n12679 ;
  assign n12950 = ~n8372 & ~n12682 ;
  assign n12951 = ~n12949 & ~n12950 ;
  assign n12952 = n11826 & ~n12951 ;
  assign n12943 = n7947 & ~n8521 ;
  assign n12944 = \P1_P1_InstQueue_reg[1][2]/NET0131  & ~n8520 ;
  assign n12945 = ~n8376 & n12944 ;
  assign n12946 = ~n12943 & ~n12945 ;
  assign n12948 = ~n11826 & n12946 ;
  assign n12953 = n8282 & ~n12948 ;
  assign n12954 = ~n12952 & n12953 ;
  assign n12947 = n8287 & ~n12946 ;
  assign n12955 = n8520 & ~n12718 ;
  assign n12956 = ~n12944 & ~n12955 ;
  assign n12957 = n8350 & ~n12956 ;
  assign n12958 = \P1_P1_InstQueue_reg[1][2]/NET0131  & ~n8366 ;
  assign n12959 = ~n12957 & ~n12958 ;
  assign n12960 = ~n12947 & n12959 ;
  assign n12961 = ~n12954 & n12960 ;
  assign n12963 = n11862 & ~n12730 ;
  assign n12962 = ~n11862 & ~n12727 ;
  assign n12964 = n12388 & ~n12962 ;
  assign n12965 = ~n12963 & n12964 ;
  assign n12968 = n11871 & n12766 ;
  assign n12967 = ~\P2_P1_InstQueue_reg[0][3]/NET0131  & ~n11871 ;
  assign n12969 = n11692 & ~n12967 ;
  assign n12970 = ~n12968 & n12969 ;
  assign n12966 = \P2_P1_InstQueue_reg[0][3]/NET0131  & ~n12395 ;
  assign n12971 = n11374 & ~n11874 ;
  assign n12972 = n12393 & n12971 ;
  assign n12973 = ~n12966 & ~n12972 ;
  assign n12974 = ~n12970 & n12973 ;
  assign n12975 = ~n12965 & n12974 ;
  assign n12982 = n8378 & ~n12679 ;
  assign n12983 = ~n8378 & ~n12682 ;
  assign n12984 = ~n12982 & ~n12983 ;
  assign n12985 = n11846 & ~n12984 ;
  assign n12976 = n7947 & ~n8545 ;
  assign n12977 = \P1_P1_InstQueue_reg[2][2]/NET0131  & ~n8544 ;
  assign n12978 = ~n8520 & n12977 ;
  assign n12979 = ~n12976 & ~n12978 ;
  assign n12981 = ~n11846 & n12979 ;
  assign n12986 = n8282 & ~n12981 ;
  assign n12987 = ~n12985 & n12986 ;
  assign n12980 = n8287 & ~n12979 ;
  assign n12988 = n8544 & ~n12718 ;
  assign n12989 = ~n12977 & ~n12988 ;
  assign n12990 = n8350 & ~n12989 ;
  assign n12991 = \P1_P1_InstQueue_reg[2][2]/NET0131  & ~n8366 ;
  assign n12992 = ~n12990 & ~n12991 ;
  assign n12993 = ~n12980 & n12992 ;
  assign n12994 = ~n12987 & n12993 ;
  assign n13005 = n11862 & ~n12817 ;
  assign n13006 = ~n11862 & ~n12820 ;
  assign n13007 = ~n13005 & ~n13006 ;
  assign n13008 = n11870 & ~n13007 ;
  assign n13000 = n11383 & ~n11874 ;
  assign n12996 = \P2_P1_InstQueue_reg[0][6]/NET0131  & ~n11871 ;
  assign n13001 = ~n11873 & n12996 ;
  assign n13002 = ~n13000 & ~n13001 ;
  assign n13004 = ~n11870 & n13002 ;
  assign n13009 = n11609 & ~n13004 ;
  assign n13010 = ~n13008 & n13009 ;
  assign n12997 = n11871 & ~n12807 ;
  assign n12998 = ~n12996 & ~n12997 ;
  assign n12999 = n11692 & ~n12998 ;
  assign n12995 = \P2_P1_InstQueue_reg[0][6]/NET0131  & ~n11630 ;
  assign n13003 = n11613 & ~n13002 ;
  assign n13011 = ~n12995 & ~n13003 ;
  assign n13012 = ~n12999 & n13011 ;
  assign n13013 = ~n13010 & n13012 ;
  assign n13015 = n11891 & ~n12730 ;
  assign n13014 = ~n11891 & ~n12727 ;
  assign n13016 = n12407 & ~n13014 ;
  assign n13017 = ~n13015 & n13016 ;
  assign n13020 = n11599 & n12766 ;
  assign n13019 = ~\P2_P1_InstQueue_reg[10][3]/NET0131  & ~n11599 ;
  assign n13021 = n11692 & ~n13019 ;
  assign n13022 = ~n13020 & n13021 ;
  assign n13018 = \P2_P1_InstQueue_reg[10][3]/NET0131  & ~n12414 ;
  assign n13023 = n11374 & ~n11897 ;
  assign n13024 = n12412 & n13023 ;
  assign n13025 = ~n13018 & ~n13024 ;
  assign n13026 = ~n13022 & n13025 ;
  assign n13027 = ~n13017 & n13026 ;
  assign n13038 = n11891 & ~n12817 ;
  assign n13039 = ~n11891 & ~n12820 ;
  assign n13040 = ~n13038 & ~n13039 ;
  assign n13041 = n11896 & ~n13040 ;
  assign n13033 = n11383 & ~n11897 ;
  assign n13029 = \P2_P1_InstQueue_reg[10][6]/NET0131  & ~n11599 ;
  assign n13034 = ~n11577 & n13029 ;
  assign n13035 = ~n13033 & ~n13034 ;
  assign n13037 = ~n11896 & n13035 ;
  assign n13042 = n11609 & ~n13037 ;
  assign n13043 = ~n13041 & n13042 ;
  assign n13030 = n11599 & ~n12807 ;
  assign n13031 = ~n13029 & ~n13030 ;
  assign n13032 = n11692 & ~n13031 ;
  assign n13028 = \P2_P1_InstQueue_reg[10][6]/NET0131  & ~n11630 ;
  assign n13036 = n11613 & ~n13035 ;
  assign n13044 = ~n13028 & ~n13036 ;
  assign n13045 = ~n13032 & n13044 ;
  assign n13046 = ~n13043 & n13045 ;
  assign n13048 = n11577 & ~n12730 ;
  assign n13047 = ~n11577 & ~n12727 ;
  assign n13049 = n12426 & ~n13047 ;
  assign n13050 = ~n13048 & n13049 ;
  assign n13053 = n11919 & n12766 ;
  assign n13052 = ~\P2_P1_InstQueue_reg[12][3]/NET0131  & ~n11919 ;
  assign n13054 = n11692 & ~n13052 ;
  assign n13055 = ~n13053 & n13054 ;
  assign n13051 = \P2_P1_InstQueue_reg[12][3]/NET0131  & ~n12433 ;
  assign n13056 = n11374 & ~n11920 ;
  assign n13057 = n12431 & n13056 ;
  assign n13058 = ~n13051 & ~n13057 ;
  assign n13059 = ~n13055 & n13058 ;
  assign n13060 = ~n13050 & n13059 ;
  assign n13067 = n8376 & ~n12679 ;
  assign n13068 = ~n8376 & ~n12682 ;
  assign n13069 = ~n13067 & ~n13068 ;
  assign n13070 = n11941 & ~n13069 ;
  assign n13061 = n7947 & ~n8569 ;
  assign n13062 = \P1_P1_InstQueue_reg[3][2]/NET0131  & ~n8568 ;
  assign n13063 = ~n8544 & n13062 ;
  assign n13064 = ~n13061 & ~n13063 ;
  assign n13066 = ~n11941 & n13064 ;
  assign n13071 = n8282 & ~n13066 ;
  assign n13072 = ~n13070 & n13071 ;
  assign n13065 = n8287 & ~n13064 ;
  assign n13073 = n8568 & ~n12718 ;
  assign n13074 = ~n13062 & ~n13073 ;
  assign n13075 = n8350 & ~n13074 ;
  assign n13076 = \P1_P1_InstQueue_reg[3][2]/NET0131  & ~n8366 ;
  assign n13077 = ~n13075 & ~n13076 ;
  assign n13078 = ~n13065 & n13077 ;
  assign n13079 = ~n13072 & n13078 ;
  assign n13081 = n11599 & ~n12730 ;
  assign n13080 = ~n11599 & ~n12727 ;
  assign n13082 = n12445 & ~n13080 ;
  assign n13083 = ~n13081 & n13082 ;
  assign n13086 = n11862 & n12766 ;
  assign n13085 = ~\P2_P1_InstQueue_reg[13][3]/NET0131  & ~n11862 ;
  assign n13087 = n11692 & ~n13085 ;
  assign n13088 = ~n13086 & n13087 ;
  assign n13084 = \P2_P1_InstQueue_reg[13][3]/NET0131  & ~n12452 ;
  assign n13089 = n11374 & ~n11961 ;
  assign n13090 = n12450 & n13089 ;
  assign n13091 = ~n13084 & ~n13090 ;
  assign n13092 = ~n13088 & n13091 ;
  assign n13093 = ~n13083 & n13092 ;
  assign n13104 = n11599 & ~n12817 ;
  assign n13105 = ~n11599 & ~n12820 ;
  assign n13106 = ~n13104 & ~n13105 ;
  assign n13107 = n11960 & ~n13106 ;
  assign n13099 = n11383 & ~n11961 ;
  assign n13095 = \P2_P1_InstQueue_reg[13][6]/NET0131  & ~n11862 ;
  assign n13100 = ~n11919 & n13095 ;
  assign n13101 = ~n13099 & ~n13100 ;
  assign n13103 = ~n11960 & n13101 ;
  assign n13108 = n11609 & ~n13103 ;
  assign n13109 = ~n13107 & n13108 ;
  assign n13096 = n11862 & ~n12807 ;
  assign n13097 = ~n13095 & ~n13096 ;
  assign n13098 = n11692 & ~n13097 ;
  assign n13094 = \P2_P1_InstQueue_reg[13][6]/NET0131  & ~n11630 ;
  assign n13102 = n11613 & ~n13101 ;
  assign n13110 = ~n13094 & ~n13102 ;
  assign n13111 = ~n13098 & n13110 ;
  assign n13112 = ~n13109 & n13111 ;
  assign n13114 = n11596 & ~n12730 ;
  assign n13113 = ~n11596 & ~n12727 ;
  assign n13115 = n12464 & ~n13113 ;
  assign n13116 = ~n13114 & n13115 ;
  assign n13119 = n11865 & n12766 ;
  assign n13118 = ~\P2_P1_InstQueue_reg[14][3]/NET0131  & ~n11865 ;
  assign n13120 = n11692 & ~n13118 ;
  assign n13121 = ~n13119 & n13120 ;
  assign n13117 = \P2_P1_InstQueue_reg[14][3]/NET0131  & ~n12471 ;
  assign n13122 = n11374 & ~n11869 ;
  assign n13123 = n12469 & n13122 ;
  assign n13124 = ~n13117 & ~n13123 ;
  assign n13125 = ~n13121 & n13124 ;
  assign n13126 = ~n13116 & n13125 ;
  assign n13137 = n11596 & ~n12817 ;
  assign n13138 = ~n11596 & ~n12820 ;
  assign n13139 = ~n13137 & ~n13138 ;
  assign n13140 = n11981 & ~n13139 ;
  assign n13132 = n11383 & ~n11869 ;
  assign n13128 = \P2_P1_InstQueue_reg[14][6]/NET0131  & ~n11865 ;
  assign n13133 = ~n11862 & n13128 ;
  assign n13134 = ~n13132 & ~n13133 ;
  assign n13136 = ~n11981 & n13134 ;
  assign n13141 = n11609 & ~n13136 ;
  assign n13142 = ~n13140 & n13141 ;
  assign n13129 = n11865 & ~n12807 ;
  assign n13130 = ~n13128 & ~n13129 ;
  assign n13131 = n11692 & ~n13130 ;
  assign n13127 = \P2_P1_InstQueue_reg[14][6]/NET0131  & ~n11630 ;
  assign n13135 = n11613 & ~n13134 ;
  assign n13143 = ~n13127 & ~n13135 ;
  assign n13144 = ~n13131 & n13143 ;
  assign n13145 = ~n13142 & n13144 ;
  assign n13147 = n11919 & ~n12730 ;
  assign n13146 = ~n11919 & ~n12727 ;
  assign n13148 = n12483 & ~n13146 ;
  assign n13149 = ~n13147 & n13148 ;
  assign n13152 = n11873 & n12766 ;
  assign n13151 = ~\P2_P1_InstQueue_reg[15][3]/NET0131  & ~n11873 ;
  assign n13153 = n11692 & ~n13151 ;
  assign n13154 = ~n13152 & n13153 ;
  assign n13150 = \P2_P1_InstQueue_reg[15][3]/NET0131  & ~n12490 ;
  assign n13155 = n11374 & ~n12002 ;
  assign n13156 = n12488 & n13155 ;
  assign n13157 = ~n13150 & ~n13156 ;
  assign n13158 = ~n13154 & n13157 ;
  assign n13159 = ~n13149 & n13158 ;
  assign n13170 = n11919 & ~n12817 ;
  assign n13171 = ~n11919 & ~n12820 ;
  assign n13172 = ~n13170 & ~n13171 ;
  assign n13173 = n12001 & ~n13172 ;
  assign n13165 = n11383 & ~n12002 ;
  assign n13161 = \P2_P1_InstQueue_reg[15][6]/NET0131  & ~n11873 ;
  assign n13166 = ~n11865 & n13161 ;
  assign n13167 = ~n13165 & ~n13166 ;
  assign n13169 = ~n12001 & n13167 ;
  assign n13174 = n11609 & ~n13169 ;
  assign n13175 = ~n13173 & n13174 ;
  assign n13162 = n11873 & ~n12807 ;
  assign n13163 = ~n13161 & ~n13162 ;
  assign n13164 = n11692 & ~n13163 ;
  assign n13160 = \P2_P1_InstQueue_reg[15][6]/NET0131  & ~n11630 ;
  assign n13168 = n11613 & ~n13167 ;
  assign n13176 = ~n13160 & ~n13168 ;
  assign n13177 = ~n13164 & n13176 ;
  assign n13178 = ~n13175 & n13177 ;
  assign n13180 = n11865 & ~n12730 ;
  assign n13179 = ~n11865 & ~n12727 ;
  assign n13181 = n12502 & ~n13179 ;
  assign n13182 = ~n13180 & n13181 ;
  assign n13185 = n12023 & n12766 ;
  assign n13184 = ~\P2_P1_InstQueue_reg[1][3]/NET0131  & ~n12023 ;
  assign n13186 = n11692 & ~n13184 ;
  assign n13187 = ~n13185 & n13186 ;
  assign n13183 = \P2_P1_InstQueue_reg[1][3]/NET0131  & ~n12509 ;
  assign n13188 = n11374 & ~n12024 ;
  assign n13189 = n12507 & n13188 ;
  assign n13190 = ~n13183 & ~n13189 ;
  assign n13191 = ~n13187 & n13190 ;
  assign n13192 = ~n13182 & n13191 ;
  assign n13203 = n11865 & ~n12817 ;
  assign n13204 = ~n11865 & ~n12820 ;
  assign n13205 = ~n13203 & ~n13204 ;
  assign n13206 = n12022 & ~n13205 ;
  assign n13198 = n11383 & ~n12024 ;
  assign n13194 = \P2_P1_InstQueue_reg[1][6]/NET0131  & ~n12023 ;
  assign n13199 = ~n11871 & n13194 ;
  assign n13200 = ~n13198 & ~n13199 ;
  assign n13202 = ~n12022 & n13200 ;
  assign n13207 = n11609 & ~n13202 ;
  assign n13208 = ~n13206 & n13207 ;
  assign n13195 = n12023 & ~n12807 ;
  assign n13196 = ~n13194 & ~n13195 ;
  assign n13197 = n11692 & ~n13196 ;
  assign n13193 = \P2_P1_InstQueue_reg[1][6]/NET0131  & ~n11630 ;
  assign n13201 = n11613 & ~n13200 ;
  assign n13209 = ~n13193 & ~n13201 ;
  assign n13210 = ~n13197 & n13209 ;
  assign n13211 = ~n13208 & n13210 ;
  assign n13218 = n8520 & ~n12679 ;
  assign n13219 = ~n8520 & ~n12682 ;
  assign n13220 = ~n13218 & ~n13219 ;
  assign n13221 = n12045 & ~n13220 ;
  assign n13212 = n7947 & ~n8593 ;
  assign n13213 = \P1_P1_InstQueue_reg[4][2]/NET0131  & ~n8592 ;
  assign n13214 = ~n8568 & n13213 ;
  assign n13215 = ~n13212 & ~n13214 ;
  assign n13217 = ~n12045 & n13215 ;
  assign n13222 = n8282 & ~n13217 ;
  assign n13223 = ~n13221 & n13222 ;
  assign n13216 = n8287 & ~n13215 ;
  assign n13224 = n8592 & ~n12718 ;
  assign n13225 = ~n13213 & ~n13224 ;
  assign n13226 = n8350 & ~n13225 ;
  assign n13227 = \P1_P1_InstQueue_reg[4][2]/NET0131  & ~n8366 ;
  assign n13228 = ~n13226 & ~n13227 ;
  assign n13229 = ~n13216 & n13228 ;
  assign n13230 = ~n13223 & n13229 ;
  assign n13232 = n11873 & ~n12730 ;
  assign n13231 = ~n11873 & ~n12727 ;
  assign n13233 = n12521 & ~n13231 ;
  assign n13234 = ~n13232 & n13233 ;
  assign n13237 = n12065 & n12766 ;
  assign n13236 = ~\P2_P1_InstQueue_reg[2][3]/NET0131  & ~n12065 ;
  assign n13238 = n11692 & ~n13236 ;
  assign n13239 = ~n13237 & n13238 ;
  assign n13235 = \P2_P1_InstQueue_reg[2][3]/NET0131  & ~n12528 ;
  assign n13240 = n11374 & ~n12066 ;
  assign n13241 = n12526 & n13240 ;
  assign n13242 = ~n13235 & ~n13241 ;
  assign n13243 = ~n13239 & n13242 ;
  assign n13244 = ~n13234 & n13243 ;
  assign n13255 = n11873 & ~n12817 ;
  assign n13256 = ~n11873 & ~n12820 ;
  assign n13257 = ~n13255 & ~n13256 ;
  assign n13258 = n12064 & ~n13257 ;
  assign n13250 = n11383 & ~n12066 ;
  assign n13246 = \P2_P1_InstQueue_reg[2][6]/NET0131  & ~n12065 ;
  assign n13251 = ~n12023 & n13246 ;
  assign n13252 = ~n13250 & ~n13251 ;
  assign n13254 = ~n12064 & n13252 ;
  assign n13259 = n11609 & ~n13254 ;
  assign n13260 = ~n13258 & n13259 ;
  assign n13247 = n12065 & ~n12807 ;
  assign n13248 = ~n13246 & ~n13247 ;
  assign n13249 = n11692 & ~n13248 ;
  assign n13245 = \P2_P1_InstQueue_reg[2][6]/NET0131  & ~n11630 ;
  assign n13253 = n11613 & ~n13252 ;
  assign n13261 = ~n13245 & ~n13253 ;
  assign n13262 = ~n13249 & n13261 ;
  assign n13263 = ~n13260 & n13262 ;
  assign n13265 = n11871 & ~n12730 ;
  assign n13264 = ~n11871 & ~n12727 ;
  assign n13266 = n12540 & ~n13264 ;
  assign n13267 = ~n13265 & n13266 ;
  assign n13270 = n12087 & n12766 ;
  assign n13269 = ~\P2_P1_InstQueue_reg[3][3]/NET0131  & ~n12087 ;
  assign n13271 = n11692 & ~n13269 ;
  assign n13272 = ~n13270 & n13271 ;
  assign n13268 = \P2_P1_InstQueue_reg[3][3]/NET0131  & ~n12547 ;
  assign n13273 = n11374 & ~n12088 ;
  assign n13274 = n12545 & n13273 ;
  assign n13275 = ~n13268 & ~n13274 ;
  assign n13276 = ~n13272 & n13275 ;
  assign n13277 = ~n13267 & n13276 ;
  assign n13288 = n11871 & ~n12817 ;
  assign n13289 = ~n11871 & ~n12820 ;
  assign n13290 = ~n13288 & ~n13289 ;
  assign n13291 = n12086 & ~n13290 ;
  assign n13283 = n11383 & ~n12088 ;
  assign n13279 = \P2_P1_InstQueue_reg[3][6]/NET0131  & ~n12087 ;
  assign n13284 = ~n12065 & n13279 ;
  assign n13285 = ~n13283 & ~n13284 ;
  assign n13287 = ~n12086 & n13285 ;
  assign n13292 = n11609 & ~n13287 ;
  assign n13293 = ~n13291 & n13292 ;
  assign n13280 = n12087 & ~n12807 ;
  assign n13281 = ~n13279 & ~n13280 ;
  assign n13282 = n11692 & ~n13281 ;
  assign n13278 = \P2_P1_InstQueue_reg[3][6]/NET0131  & ~n11630 ;
  assign n13286 = n11613 & ~n13285 ;
  assign n13294 = ~n13278 & ~n13286 ;
  assign n13295 = ~n13282 & n13294 ;
  assign n13296 = ~n13293 & n13295 ;
  assign n13298 = n12023 & ~n12730 ;
  assign n13297 = ~n12023 & ~n12727 ;
  assign n13299 = n12559 & ~n13297 ;
  assign n13300 = ~n13298 & n13299 ;
  assign n13303 = n12109 & n12766 ;
  assign n13302 = ~\P2_P1_InstQueue_reg[4][3]/NET0131  & ~n12109 ;
  assign n13304 = n11692 & ~n13302 ;
  assign n13305 = ~n13303 & n13304 ;
  assign n13301 = \P2_P1_InstQueue_reg[4][3]/NET0131  & ~n12566 ;
  assign n13306 = n11374 & ~n12110 ;
  assign n13307 = n12564 & n13306 ;
  assign n13308 = ~n13301 & ~n13307 ;
  assign n13309 = ~n13305 & n13308 ;
  assign n13310 = ~n13300 & n13309 ;
  assign n13321 = n12023 & ~n12817 ;
  assign n13322 = ~n12023 & ~n12820 ;
  assign n13323 = ~n13321 & ~n13322 ;
  assign n13324 = n12108 & ~n13323 ;
  assign n13316 = n11383 & ~n12110 ;
  assign n13312 = \P2_P1_InstQueue_reg[4][6]/NET0131  & ~n12109 ;
  assign n13317 = ~n12087 & n13312 ;
  assign n13318 = ~n13316 & ~n13317 ;
  assign n13320 = ~n12108 & n13318 ;
  assign n13325 = n11609 & ~n13320 ;
  assign n13326 = ~n13324 & n13325 ;
  assign n13313 = n12109 & ~n12807 ;
  assign n13314 = ~n13312 & ~n13313 ;
  assign n13315 = n11692 & ~n13314 ;
  assign n13311 = \P2_P1_InstQueue_reg[4][6]/NET0131  & ~n11630 ;
  assign n13319 = n11613 & ~n13318 ;
  assign n13327 = ~n13311 & ~n13319 ;
  assign n13328 = ~n13315 & n13327 ;
  assign n13329 = ~n13326 & n13328 ;
  assign n13331 = n12065 & ~n12730 ;
  assign n13330 = ~n12065 & ~n12727 ;
  assign n13332 = n12578 & ~n13330 ;
  assign n13333 = ~n13331 & n13332 ;
  assign n13336 = n12131 & n12766 ;
  assign n13335 = ~\P2_P1_InstQueue_reg[5][3]/NET0131  & ~n12131 ;
  assign n13337 = n11692 & ~n13335 ;
  assign n13338 = ~n13336 & n13337 ;
  assign n13334 = \P2_P1_InstQueue_reg[5][3]/NET0131  & ~n12585 ;
  assign n13339 = n11374 & ~n12132 ;
  assign n13340 = n12583 & n13339 ;
  assign n13341 = ~n13334 & ~n13340 ;
  assign n13342 = ~n13338 & n13341 ;
  assign n13343 = ~n13333 & n13342 ;
  assign n13354 = n12065 & ~n12817 ;
  assign n13355 = ~n12065 & ~n12820 ;
  assign n13356 = ~n13354 & ~n13355 ;
  assign n13357 = n12130 & ~n13356 ;
  assign n13349 = n11383 & ~n12132 ;
  assign n13345 = \P2_P1_InstQueue_reg[5][6]/NET0131  & ~n12131 ;
  assign n13350 = ~n12109 & n13345 ;
  assign n13351 = ~n13349 & ~n13350 ;
  assign n13353 = ~n12130 & n13351 ;
  assign n13358 = n11609 & ~n13353 ;
  assign n13359 = ~n13357 & n13358 ;
  assign n13346 = n12131 & ~n12807 ;
  assign n13347 = ~n13345 & ~n13346 ;
  assign n13348 = n11692 & ~n13347 ;
  assign n13344 = \P2_P1_InstQueue_reg[5][6]/NET0131  & ~n11630 ;
  assign n13352 = n11613 & ~n13351 ;
  assign n13360 = ~n13344 & ~n13352 ;
  assign n13361 = ~n13348 & n13360 ;
  assign n13362 = ~n13359 & n13361 ;
  assign n13369 = n8544 & ~n12679 ;
  assign n13370 = ~n8544 & ~n12682 ;
  assign n13371 = ~n13369 & ~n13370 ;
  assign n13372 = n12153 & ~n13371 ;
  assign n13363 = n7947 & ~n8617 ;
  assign n13364 = \P1_P1_InstQueue_reg[5][2]/NET0131  & ~n8616 ;
  assign n13365 = ~n8592 & n13364 ;
  assign n13366 = ~n13363 & ~n13365 ;
  assign n13368 = ~n12153 & n13366 ;
  assign n13373 = n8282 & ~n13368 ;
  assign n13374 = ~n13372 & n13373 ;
  assign n13367 = n8287 & ~n13366 ;
  assign n13375 = n8616 & ~n12718 ;
  assign n13376 = ~n13364 & ~n13375 ;
  assign n13377 = n8350 & ~n13376 ;
  assign n13378 = \P1_P1_InstQueue_reg[5][2]/NET0131  & ~n8366 ;
  assign n13379 = ~n13377 & ~n13378 ;
  assign n13380 = ~n13367 & n13379 ;
  assign n13381 = ~n13374 & n13380 ;
  assign n13383 = n12087 & ~n12730 ;
  assign n13382 = ~n12087 & ~n12727 ;
  assign n13384 = n12597 & ~n13382 ;
  assign n13385 = ~n13383 & n13384 ;
  assign n13388 = n12173 & n12766 ;
  assign n13387 = ~\P2_P1_InstQueue_reg[6][3]/NET0131  & ~n12173 ;
  assign n13389 = n11692 & ~n13387 ;
  assign n13390 = ~n13388 & n13389 ;
  assign n13386 = \P2_P1_InstQueue_reg[6][3]/NET0131  & ~n12604 ;
  assign n13391 = n11374 & ~n12174 ;
  assign n13392 = n12602 & n13391 ;
  assign n13393 = ~n13386 & ~n13392 ;
  assign n13394 = ~n13390 & n13393 ;
  assign n13395 = ~n13385 & n13394 ;
  assign n13406 = n12087 & ~n12817 ;
  assign n13407 = ~n12087 & ~n12820 ;
  assign n13408 = ~n13406 & ~n13407 ;
  assign n13409 = n12172 & ~n13408 ;
  assign n13401 = n11383 & ~n12174 ;
  assign n13397 = \P2_P1_InstQueue_reg[6][6]/NET0131  & ~n12173 ;
  assign n13402 = ~n12131 & n13397 ;
  assign n13403 = ~n13401 & ~n13402 ;
  assign n13405 = ~n12172 & n13403 ;
  assign n13410 = n11609 & ~n13405 ;
  assign n13411 = ~n13409 & n13410 ;
  assign n13398 = n12173 & ~n12807 ;
  assign n13399 = ~n13397 & ~n13398 ;
  assign n13400 = n11692 & ~n13399 ;
  assign n13396 = \P2_P1_InstQueue_reg[6][6]/NET0131  & ~n11630 ;
  assign n13404 = n11613 & ~n13403 ;
  assign n13412 = ~n13396 & ~n13404 ;
  assign n13413 = ~n13400 & n13412 ;
  assign n13414 = ~n13411 & n13413 ;
  assign n13416 = n12109 & ~n12730 ;
  assign n13415 = ~n12109 & ~n12727 ;
  assign n13417 = n12616 & ~n13415 ;
  assign n13418 = ~n13416 & n13417 ;
  assign n13421 = n11891 & n12766 ;
  assign n13420 = ~\P2_P1_InstQueue_reg[7][3]/NET0131  & ~n11891 ;
  assign n13422 = n11692 & ~n13420 ;
  assign n13423 = ~n13421 & n13422 ;
  assign n13419 = \P2_P1_InstQueue_reg[7][3]/NET0131  & ~n12623 ;
  assign n13424 = n11374 & ~n12195 ;
  assign n13425 = n12621 & n13424 ;
  assign n13426 = ~n13419 & ~n13425 ;
  assign n13427 = ~n13423 & n13426 ;
  assign n13428 = ~n13418 & n13427 ;
  assign n13439 = n12109 & ~n12817 ;
  assign n13440 = ~n12109 & ~n12820 ;
  assign n13441 = ~n13439 & ~n13440 ;
  assign n13442 = n12194 & ~n13441 ;
  assign n13434 = n11383 & ~n12195 ;
  assign n13430 = \P2_P1_InstQueue_reg[7][6]/NET0131  & ~n11891 ;
  assign n13435 = ~n12173 & n13430 ;
  assign n13436 = ~n13434 & ~n13435 ;
  assign n13438 = ~n12194 & n13436 ;
  assign n13443 = n11609 & ~n13438 ;
  assign n13444 = ~n13442 & n13443 ;
  assign n13431 = n11891 & ~n12807 ;
  assign n13432 = ~n13430 & ~n13431 ;
  assign n13433 = n11692 & ~n13432 ;
  assign n13429 = \P2_P1_InstQueue_reg[7][6]/NET0131  & ~n11630 ;
  assign n13437 = n11613 & ~n13436 ;
  assign n13445 = ~n13429 & ~n13437 ;
  assign n13446 = ~n13433 & n13445 ;
  assign n13447 = ~n13444 & n13446 ;
  assign n13449 = n12131 & ~n12730 ;
  assign n13448 = ~n12131 & ~n12727 ;
  assign n13450 = n12635 & ~n13448 ;
  assign n13451 = ~n13449 & n13450 ;
  assign n13454 = n10105 & n12766 ;
  assign n13453 = ~\P2_P1_InstQueue_reg[8][3]/NET0131  & ~n10105 ;
  assign n13455 = n11692 & ~n13453 ;
  assign n13456 = ~n13454 & n13455 ;
  assign n13452 = \P2_P1_InstQueue_reg[8][3]/NET0131  & ~n12642 ;
  assign n13457 = n11374 & ~n11895 ;
  assign n13458 = n12640 & n13457 ;
  assign n13459 = ~n13452 & ~n13458 ;
  assign n13460 = ~n13456 & n13459 ;
  assign n13461 = ~n13451 & n13460 ;
  assign n13472 = n12131 & ~n12817 ;
  assign n13473 = ~n12131 & ~n12820 ;
  assign n13474 = ~n13472 & ~n13473 ;
  assign n13475 = n12215 & ~n13474 ;
  assign n13467 = n11383 & ~n11895 ;
  assign n13463 = \P2_P1_InstQueue_reg[8][6]/NET0131  & ~n10105 ;
  assign n13468 = ~n11891 & n13463 ;
  assign n13469 = ~n13467 & ~n13468 ;
  assign n13471 = ~n12215 & n13469 ;
  assign n13476 = n11609 & ~n13471 ;
  assign n13477 = ~n13475 & n13476 ;
  assign n13464 = n10105 & ~n12807 ;
  assign n13465 = ~n13463 & ~n13464 ;
  assign n13466 = n11692 & ~n13465 ;
  assign n13462 = \P2_P1_InstQueue_reg[8][6]/NET0131  & ~n11630 ;
  assign n13470 = n11613 & ~n13469 ;
  assign n13478 = ~n13462 & ~n13470 ;
  assign n13479 = ~n13466 & n13478 ;
  assign n13480 = ~n13477 & n13479 ;
  assign n13482 = n12173 & ~n12730 ;
  assign n13481 = ~n12173 & ~n12727 ;
  assign n13483 = n12654 & ~n13481 ;
  assign n13484 = ~n13482 & n13483 ;
  assign n13487 = n11577 & n12766 ;
  assign n13486 = ~\P2_P1_InstQueue_reg[9][3]/NET0131  & ~n11577 ;
  assign n13488 = n11692 & ~n13486 ;
  assign n13489 = ~n13487 & n13488 ;
  assign n13485 = \P2_P1_InstQueue_reg[9][3]/NET0131  & ~n12661 ;
  assign n13490 = n11374 & ~n11592 ;
  assign n13491 = n12659 & n13490 ;
  assign n13492 = ~n13485 & ~n13491 ;
  assign n13493 = ~n13489 & n13492 ;
  assign n13494 = ~n13484 & n13493 ;
  assign n13505 = n12173 & ~n12817 ;
  assign n13506 = ~n12173 & ~n12820 ;
  assign n13507 = ~n13505 & ~n13506 ;
  assign n13508 = n12235 & ~n13507 ;
  assign n13500 = n11383 & ~n11592 ;
  assign n13496 = \P2_P1_InstQueue_reg[9][6]/NET0131  & ~n11577 ;
  assign n13501 = ~n10105 & n13496 ;
  assign n13502 = ~n13500 & ~n13501 ;
  assign n13504 = ~n12235 & n13502 ;
  assign n13509 = n11609 & ~n13504 ;
  assign n13510 = ~n13508 & n13509 ;
  assign n13497 = n11577 & ~n12807 ;
  assign n13498 = ~n13496 & ~n13497 ;
  assign n13499 = n11692 & ~n13498 ;
  assign n13495 = \P2_P1_InstQueue_reg[9][6]/NET0131  & ~n11630 ;
  assign n13503 = n11613 & ~n13502 ;
  assign n13511 = ~n13495 & ~n13503 ;
  assign n13512 = ~n13499 & n13511 ;
  assign n13513 = ~n13510 & n13512 ;
  assign n13520 = n8568 & ~n12679 ;
  assign n13521 = ~n8568 & ~n12682 ;
  assign n13522 = ~n13520 & ~n13521 ;
  assign n13523 = n12256 & ~n13522 ;
  assign n13514 = n7947 & ~n8641 ;
  assign n13515 = \P1_P1_InstQueue_reg[6][2]/NET0131  & ~n8640 ;
  assign n13516 = ~n8616 & n13515 ;
  assign n13517 = ~n13514 & ~n13516 ;
  assign n13519 = ~n12256 & n13517 ;
  assign n13524 = n8282 & ~n13519 ;
  assign n13525 = ~n13523 & n13524 ;
  assign n13518 = n8287 & ~n13517 ;
  assign n13526 = n8640 & ~n12718 ;
  assign n13527 = ~n13515 & ~n13526 ;
  assign n13528 = n8350 & ~n13527 ;
  assign n13529 = \P1_P1_InstQueue_reg[6][2]/NET0131  & ~n8366 ;
  assign n13530 = ~n13528 & ~n13529 ;
  assign n13531 = ~n13518 & n13530 ;
  assign n13532 = ~n13525 & n13531 ;
  assign n13539 = n8592 & ~n12679 ;
  assign n13540 = ~n8592 & ~n12682 ;
  assign n13541 = ~n13539 & ~n13540 ;
  assign n13542 = n12276 & ~n13541 ;
  assign n13533 = n7947 & ~n8664 ;
  assign n13534 = \P1_P1_InstQueue_reg[7][2]/NET0131  & ~n8407 ;
  assign n13535 = ~n8640 & n13534 ;
  assign n13536 = ~n13533 & ~n13535 ;
  assign n13538 = ~n12276 & n13536 ;
  assign n13543 = n8282 & ~n13538 ;
  assign n13544 = ~n13542 & n13543 ;
  assign n13537 = n8287 & ~n13536 ;
  assign n13545 = n8407 & ~n12718 ;
  assign n13546 = ~n13534 & ~n13545 ;
  assign n13547 = n8350 & ~n13546 ;
  assign n13548 = \P1_P1_InstQueue_reg[7][2]/NET0131  & ~n8366 ;
  assign n13549 = ~n13547 & ~n13548 ;
  assign n13550 = ~n13537 & n13549 ;
  assign n13551 = ~n13544 & n13550 ;
  assign n13558 = n8616 & ~n12679 ;
  assign n13559 = ~n8616 & ~n12682 ;
  assign n13560 = ~n13558 & ~n13559 ;
  assign n13561 = n12296 & ~n13560 ;
  assign n13552 = n7947 & ~n8410 ;
  assign n13553 = \P1_P1_InstQueue_reg[8][2]/NET0131  & ~n8139 ;
  assign n13554 = ~n8407 & n13553 ;
  assign n13555 = ~n13552 & ~n13554 ;
  assign n13557 = ~n12296 & n13555 ;
  assign n13562 = n8282 & ~n13557 ;
  assign n13563 = ~n13561 & n13562 ;
  assign n13556 = n8287 & ~n13555 ;
  assign n13564 = n8139 & ~n12718 ;
  assign n13565 = ~n13553 & ~n13564 ;
  assign n13566 = n8350 & ~n13565 ;
  assign n13567 = \P1_P1_InstQueue_reg[8][2]/NET0131  & ~n8366 ;
  assign n13568 = ~n13566 & ~n13567 ;
  assign n13569 = ~n13556 & n13568 ;
  assign n13570 = ~n13563 & n13569 ;
  assign n13577 = n8640 & ~n12679 ;
  assign n13578 = ~n8640 & ~n12682 ;
  assign n13579 = ~n13577 & ~n13578 ;
  assign n13580 = n12316 & ~n13579 ;
  assign n13571 = n7947 & ~n8709 ;
  assign n13572 = \P1_P1_InstQueue_reg[9][2]/NET0131  & ~n4327 ;
  assign n13573 = ~n8139 & n13572 ;
  assign n13574 = ~n13571 & ~n13573 ;
  assign n13576 = ~n12316 & n13574 ;
  assign n13581 = n8282 & ~n13576 ;
  assign n13582 = ~n13580 & n13581 ;
  assign n13575 = n8287 & ~n13574 ;
  assign n13583 = n4327 & ~n12718 ;
  assign n13584 = ~n13572 & ~n13583 ;
  assign n13585 = n8350 & ~n13584 ;
  assign n13586 = \P1_P1_InstQueue_reg[9][2]/NET0131  & ~n8366 ;
  assign n13587 = ~n13585 & ~n13586 ;
  assign n13588 = ~n13575 & n13587 ;
  assign n13589 = ~n13582 & n13588 ;
  assign n13598 = ~n8094 & n8106 ;
  assign n13599 = ~n9311 & ~n13598 ;
  assign n13600 = n4327 & ~n13599 ;
  assign n13593 = ~n7933 & ~n8146 ;
  assign n13594 = \P1_P1_InstQueue_reg[11][5]/NET0131  & ~n8142 ;
  assign n13595 = ~n8145 & n13594 ;
  assign n13596 = ~n13593 & ~n13595 ;
  assign n13597 = ~n4327 & n13596 ;
  assign n13601 = ~n8139 & ~n13597 ;
  assign n13602 = ~n13600 & n13601 ;
  assign n13590 = ~n8234 & n8248 ;
  assign n13591 = ~n9322 & ~n13590 ;
  assign n13592 = n8139 & n13591 ;
  assign n13603 = \P1_P1_DataWidth_reg[1]/NET0131  & ~n13592 ;
  assign n13604 = ~n13602 & n13603 ;
  assign n13605 = ~\P1_P1_DataWidth_reg[1]/NET0131  & n13596 ;
  assign n13606 = n8282 & ~n13605 ;
  assign n13607 = ~n13604 & n13606 ;
  assign n13608 = n8287 & ~n13596 ;
  assign n13609 = \P1_P1_InstQueue_reg[14][5]/NET0131  & n8291 ;
  assign n13610 = \P1_P1_InstQueue_reg[3][5]/NET0131  & n8323 ;
  assign n13611 = \P1_P1_InstQueue_reg[1][5]/NET0131  & n8299 ;
  assign n13625 = ~n13610 & ~n13611 ;
  assign n13612 = \P1_P1_InstQueue_reg[11][5]/NET0131  & n8312 ;
  assign n13613 = \P1_P1_InstQueue_reg[8][5]/NET0131  & n8305 ;
  assign n13626 = ~n13612 & ~n13613 ;
  assign n13635 = n13625 & n13626 ;
  assign n13636 = ~n13609 & n13635 ;
  assign n13624 = \P1_P1_InstQueue_reg[10][5]/NET0131  & n8303 ;
  assign n13622 = \P1_P1_InstQueue_reg[13][5]/NET0131  & n8327 ;
  assign n13623 = \P1_P1_InstQueue_reg[0][5]/NET0131  & n8309 ;
  assign n13631 = ~n13622 & ~n13623 ;
  assign n13632 = ~n13624 & n13631 ;
  assign n13618 = \P1_P1_InstQueue_reg[6][5]/NET0131  & n8316 ;
  assign n13619 = \P1_P1_InstQueue_reg[7][5]/NET0131  & n8318 ;
  assign n13629 = ~n13618 & ~n13619 ;
  assign n13620 = \P1_P1_InstQueue_reg[15][5]/NET0131  & n8321 ;
  assign n13621 = \P1_P1_InstQueue_reg[5][5]/NET0131  & n8307 ;
  assign n13630 = ~n13620 & ~n13621 ;
  assign n13633 = n13629 & n13630 ;
  assign n13614 = \P1_P1_InstQueue_reg[4][5]/NET0131  & n8295 ;
  assign n13615 = \P1_P1_InstQueue_reg[12][5]/NET0131  & n8329 ;
  assign n13627 = ~n13614 & ~n13615 ;
  assign n13616 = \P1_P1_InstQueue_reg[9][5]/NET0131  & n8325 ;
  assign n13617 = \P1_P1_InstQueue_reg[2][5]/NET0131  & n8314 ;
  assign n13628 = ~n13616 & ~n13617 ;
  assign n13634 = n13627 & n13628 ;
  assign n13637 = n13633 & n13634 ;
  assign n13638 = n13632 & n13637 ;
  assign n13639 = n13636 & n13638 ;
  assign n13640 = n8142 & ~n13639 ;
  assign n13641 = ~n13594 & ~n13640 ;
  assign n13642 = n8350 & ~n13641 ;
  assign n13643 = \P1_P1_InstQueue_reg[11][5]/NET0131  & ~n8366 ;
  assign n13644 = ~n13642 & ~n13643 ;
  assign n13645 = ~n13608 & n13644 ;
  assign n13646 = ~n13607 & n13645 ;
  assign n13653 = n8372 & ~n13599 ;
  assign n13648 = ~n7933 & ~n8379 ;
  assign n13649 = \P1_P1_InstQueue_reg[0][5]/NET0131  & ~n8376 ;
  assign n13650 = ~n8378 & n13649 ;
  assign n13651 = ~n13648 & ~n13650 ;
  assign n13652 = ~n8372 & n13651 ;
  assign n13654 = ~n8375 & ~n13652 ;
  assign n13655 = ~n13653 & n13654 ;
  assign n13647 = n8375 & n13591 ;
  assign n13656 = \P1_P1_DataWidth_reg[1]/NET0131  & ~n13647 ;
  assign n13657 = ~n13655 & n13656 ;
  assign n13658 = ~\P1_P1_DataWidth_reg[1]/NET0131  & n13651 ;
  assign n13659 = n8282 & ~n13658 ;
  assign n13660 = ~n13657 & n13659 ;
  assign n13661 = n8287 & ~n13651 ;
  assign n13662 = n8376 & ~n13639 ;
  assign n13663 = ~n13649 & ~n13662 ;
  assign n13664 = n8350 & ~n13663 ;
  assign n13665 = \P1_P1_InstQueue_reg[0][5]/NET0131  & ~n8366 ;
  assign n13666 = ~n13664 & ~n13665 ;
  assign n13667 = ~n13661 & n13666 ;
  assign n13668 = ~n13660 & n13667 ;
  assign n13669 = n8407 & n13591 ;
  assign n13670 = n8139 & n13599 ;
  assign n13671 = ~n13669 & ~n13670 ;
  assign n13672 = \P1_P1_DataWidth_reg[1]/NET0131  & ~n13671 ;
  assign n13673 = ~n7933 & ~n8401 ;
  assign n13674 = \P1_P1_InstQueue_reg[10][5]/NET0131  & ~n8145 ;
  assign n13675 = ~n4327 & n13674 ;
  assign n13676 = ~n13673 & ~n13675 ;
  assign n13677 = ~n9418 & ~n13676 ;
  assign n13678 = ~n13672 & ~n13677 ;
  assign n13679 = n8282 & ~n13678 ;
  assign n13681 = n8287 & ~n13676 ;
  assign n13680 = \P1_P1_InstQueue_reg[10][5]/NET0131  & ~n8366 ;
  assign n13682 = n8145 & ~n13639 ;
  assign n13683 = ~n13674 & ~n13682 ;
  assign n13684 = n8350 & ~n13683 ;
  assign n13685 = ~n13680 & ~n13684 ;
  assign n13686 = ~n13681 & n13685 ;
  assign n13687 = ~n13679 & n13686 ;
  assign n13694 = n8145 & ~n13599 ;
  assign n13689 = ~n7933 & ~n8428 ;
  assign n13690 = \P1_P1_InstQueue_reg[12][5]/NET0131  & ~n8427 ;
  assign n13691 = ~n8142 & n13690 ;
  assign n13692 = ~n13689 & ~n13691 ;
  assign n13693 = ~n8145 & n13692 ;
  assign n13695 = ~n4327 & ~n13693 ;
  assign n13696 = ~n13694 & n13695 ;
  assign n13688 = n4327 & n13591 ;
  assign n13697 = \P1_P1_DataWidth_reg[1]/NET0131  & ~n13688 ;
  assign n13698 = ~n13696 & n13697 ;
  assign n13699 = ~\P1_P1_DataWidth_reg[1]/NET0131  & n13692 ;
  assign n13700 = n8282 & ~n13699 ;
  assign n13701 = ~n13698 & n13700 ;
  assign n13702 = n8287 & ~n13692 ;
  assign n13703 = n8427 & ~n13639 ;
  assign n13704 = ~n13690 & ~n13703 ;
  assign n13705 = n8350 & ~n13704 ;
  assign n13706 = \P1_P1_InstQueue_reg[12][5]/NET0131  & ~n8366 ;
  assign n13707 = ~n13705 & ~n13706 ;
  assign n13708 = ~n13702 & n13707 ;
  assign n13709 = ~n13701 & n13708 ;
  assign n13716 = n8142 & ~n13599 ;
  assign n13711 = ~n7933 & ~n8451 ;
  assign n13712 = \P1_P1_InstQueue_reg[13][5]/NET0131  & ~n8375 ;
  assign n13713 = ~n8427 & n13712 ;
  assign n13714 = ~n13711 & ~n13713 ;
  assign n13715 = ~n8142 & n13714 ;
  assign n13717 = ~n8145 & ~n13715 ;
  assign n13718 = ~n13716 & n13717 ;
  assign n13710 = n8145 & n13591 ;
  assign n13719 = \P1_P1_DataWidth_reg[1]/NET0131  & ~n13710 ;
  assign n13720 = ~n13718 & n13719 ;
  assign n13721 = ~\P1_P1_DataWidth_reg[1]/NET0131  & n13714 ;
  assign n13722 = n8282 & ~n13721 ;
  assign n13723 = ~n13720 & n13722 ;
  assign n13724 = n8287 & ~n13714 ;
  assign n13725 = n8375 & ~n13639 ;
  assign n13726 = ~n13712 & ~n13725 ;
  assign n13727 = n8350 & ~n13726 ;
  assign n13728 = \P1_P1_InstQueue_reg[13][5]/NET0131  & ~n8366 ;
  assign n13729 = ~n13727 & ~n13728 ;
  assign n13730 = ~n13724 & n13729 ;
  assign n13731 = ~n13723 & n13730 ;
  assign n13738 = n8427 & ~n13599 ;
  assign n13733 = ~n7933 & ~n8474 ;
  assign n13734 = \P1_P1_InstQueue_reg[14][5]/NET0131  & ~n8372 ;
  assign n13735 = ~n8375 & n13734 ;
  assign n13736 = ~n13733 & ~n13735 ;
  assign n13737 = ~n8427 & n13736 ;
  assign n13739 = ~n8142 & ~n13737 ;
  assign n13740 = ~n13738 & n13739 ;
  assign n13732 = n8142 & n13591 ;
  assign n13741 = \P1_P1_DataWidth_reg[1]/NET0131  & ~n13732 ;
  assign n13742 = ~n13740 & n13741 ;
  assign n13743 = ~\P1_P1_DataWidth_reg[1]/NET0131  & n13736 ;
  assign n13744 = n8282 & ~n13743 ;
  assign n13745 = ~n13742 & n13744 ;
  assign n13746 = n8287 & ~n13736 ;
  assign n13747 = n8372 & ~n13639 ;
  assign n13748 = ~n13734 & ~n13747 ;
  assign n13749 = n8350 & ~n13748 ;
  assign n13750 = \P1_P1_InstQueue_reg[14][5]/NET0131  & ~n8366 ;
  assign n13751 = ~n13749 & ~n13750 ;
  assign n13752 = ~n13746 & n13751 ;
  assign n13753 = ~n13745 & n13752 ;
  assign n13760 = n8375 & ~n13599 ;
  assign n13755 = ~n7933 & ~n8497 ;
  assign n13756 = \P1_P1_InstQueue_reg[15][5]/NET0131  & ~n8378 ;
  assign n13757 = ~n8372 & n13756 ;
  assign n13758 = ~n13755 & ~n13757 ;
  assign n13759 = ~n8375 & n13758 ;
  assign n13761 = ~n8427 & ~n13759 ;
  assign n13762 = ~n13760 & n13761 ;
  assign n13754 = n8427 & n13591 ;
  assign n13763 = \P1_P1_DataWidth_reg[1]/NET0131  & ~n13754 ;
  assign n13764 = ~n13762 & n13763 ;
  assign n13765 = ~\P1_P1_DataWidth_reg[1]/NET0131  & n13758 ;
  assign n13766 = n8282 & ~n13765 ;
  assign n13767 = ~n13764 & n13766 ;
  assign n13768 = n8287 & ~n13758 ;
  assign n13769 = n8378 & ~n13639 ;
  assign n13770 = ~n13756 & ~n13769 ;
  assign n13771 = n8350 & ~n13770 ;
  assign n13772 = \P1_P1_InstQueue_reg[15][5]/NET0131  & ~n8366 ;
  assign n13773 = ~n13771 & ~n13772 ;
  assign n13774 = ~n13768 & n13773 ;
  assign n13775 = ~n13767 & n13774 ;
  assign n13782 = n8378 & ~n13599 ;
  assign n13777 = ~n7933 & ~n8521 ;
  assign n13778 = \P1_P1_InstQueue_reg[1][5]/NET0131  & ~n8520 ;
  assign n13779 = ~n8376 & n13778 ;
  assign n13780 = ~n13777 & ~n13779 ;
  assign n13781 = ~n8378 & n13780 ;
  assign n13783 = ~n8372 & ~n13781 ;
  assign n13784 = ~n13782 & n13783 ;
  assign n13776 = n8372 & n13591 ;
  assign n13785 = \P1_P1_DataWidth_reg[1]/NET0131  & ~n13776 ;
  assign n13786 = ~n13784 & n13785 ;
  assign n13787 = ~\P1_P1_DataWidth_reg[1]/NET0131  & n13780 ;
  assign n13788 = n8282 & ~n13787 ;
  assign n13789 = ~n13786 & n13788 ;
  assign n13790 = n8287 & ~n13780 ;
  assign n13791 = n8520 & ~n13639 ;
  assign n13792 = ~n13778 & ~n13791 ;
  assign n13793 = n8350 & ~n13792 ;
  assign n13794 = \P1_P1_InstQueue_reg[1][5]/NET0131  & ~n8366 ;
  assign n13795 = ~n13793 & ~n13794 ;
  assign n13796 = ~n13790 & n13795 ;
  assign n13797 = ~n13789 & n13796 ;
  assign n13804 = n8376 & ~n13599 ;
  assign n13799 = ~n7933 & ~n8545 ;
  assign n13800 = \P1_P1_InstQueue_reg[2][5]/NET0131  & ~n8544 ;
  assign n13801 = ~n8520 & n13800 ;
  assign n13802 = ~n13799 & ~n13801 ;
  assign n13803 = ~n8376 & n13802 ;
  assign n13805 = ~n8378 & ~n13803 ;
  assign n13806 = ~n13804 & n13805 ;
  assign n13798 = n8378 & n13591 ;
  assign n13807 = \P1_P1_DataWidth_reg[1]/NET0131  & ~n13798 ;
  assign n13808 = ~n13806 & n13807 ;
  assign n13809 = ~\P1_P1_DataWidth_reg[1]/NET0131  & n13802 ;
  assign n13810 = n8282 & ~n13809 ;
  assign n13811 = ~n13808 & n13810 ;
  assign n13812 = n8287 & ~n13802 ;
  assign n13813 = n8544 & ~n13639 ;
  assign n13814 = ~n13800 & ~n13813 ;
  assign n13815 = n8350 & ~n13814 ;
  assign n13816 = \P1_P1_InstQueue_reg[2][5]/NET0131  & ~n8366 ;
  assign n13817 = ~n13815 & ~n13816 ;
  assign n13818 = ~n13812 & n13817 ;
  assign n13819 = ~n13811 & n13818 ;
  assign n13826 = n8520 & ~n13599 ;
  assign n13821 = ~n7933 & ~n8569 ;
  assign n13822 = \P1_P1_InstQueue_reg[3][5]/NET0131  & ~n8568 ;
  assign n13823 = ~n8544 & n13822 ;
  assign n13824 = ~n13821 & ~n13823 ;
  assign n13825 = ~n8520 & n13824 ;
  assign n13827 = ~n8376 & ~n13825 ;
  assign n13828 = ~n13826 & n13827 ;
  assign n13820 = n8376 & n13591 ;
  assign n13829 = \P1_P1_DataWidth_reg[1]/NET0131  & ~n13820 ;
  assign n13830 = ~n13828 & n13829 ;
  assign n13831 = ~\P1_P1_DataWidth_reg[1]/NET0131  & n13824 ;
  assign n13832 = n8282 & ~n13831 ;
  assign n13833 = ~n13830 & n13832 ;
  assign n13834 = n8287 & ~n13824 ;
  assign n13835 = n8568 & ~n13639 ;
  assign n13836 = ~n13822 & ~n13835 ;
  assign n13837 = n8350 & ~n13836 ;
  assign n13838 = \P1_P1_InstQueue_reg[3][5]/NET0131  & ~n8366 ;
  assign n13839 = ~n13837 & ~n13838 ;
  assign n13840 = ~n13834 & n13839 ;
  assign n13841 = ~n13833 & n13840 ;
  assign n13848 = n8544 & ~n13599 ;
  assign n13843 = ~n7933 & ~n8593 ;
  assign n13844 = \P1_P1_InstQueue_reg[4][5]/NET0131  & ~n8592 ;
  assign n13845 = ~n8568 & n13844 ;
  assign n13846 = ~n13843 & ~n13845 ;
  assign n13847 = ~n8544 & n13846 ;
  assign n13849 = ~n8520 & ~n13847 ;
  assign n13850 = ~n13848 & n13849 ;
  assign n13842 = n8520 & n13591 ;
  assign n13851 = \P1_P1_DataWidth_reg[1]/NET0131  & ~n13842 ;
  assign n13852 = ~n13850 & n13851 ;
  assign n13853 = ~\P1_P1_DataWidth_reg[1]/NET0131  & n13846 ;
  assign n13854 = n8282 & ~n13853 ;
  assign n13855 = ~n13852 & n13854 ;
  assign n13856 = n8287 & ~n13846 ;
  assign n13857 = n8592 & ~n13639 ;
  assign n13858 = ~n13844 & ~n13857 ;
  assign n13859 = n8350 & ~n13858 ;
  assign n13860 = \P1_P1_InstQueue_reg[4][5]/NET0131  & ~n8366 ;
  assign n13861 = ~n13859 & ~n13860 ;
  assign n13862 = ~n13856 & n13861 ;
  assign n13863 = ~n13855 & n13862 ;
  assign n13870 = n8568 & ~n13599 ;
  assign n13865 = ~n7933 & ~n8617 ;
  assign n13866 = \P1_P1_InstQueue_reg[5][5]/NET0131  & ~n8616 ;
  assign n13867 = ~n8592 & n13866 ;
  assign n13868 = ~n13865 & ~n13867 ;
  assign n13869 = ~n8568 & n13868 ;
  assign n13871 = ~n8544 & ~n13869 ;
  assign n13872 = ~n13870 & n13871 ;
  assign n13864 = n8544 & n13591 ;
  assign n13873 = \P1_P1_DataWidth_reg[1]/NET0131  & ~n13864 ;
  assign n13874 = ~n13872 & n13873 ;
  assign n13875 = ~\P1_P1_DataWidth_reg[1]/NET0131  & n13868 ;
  assign n13876 = n8282 & ~n13875 ;
  assign n13877 = ~n13874 & n13876 ;
  assign n13878 = n8287 & ~n13868 ;
  assign n13879 = n8616 & ~n13639 ;
  assign n13880 = ~n13866 & ~n13879 ;
  assign n13881 = n8350 & ~n13880 ;
  assign n13882 = \P1_P1_InstQueue_reg[5][5]/NET0131  & ~n8366 ;
  assign n13883 = ~n13881 & ~n13882 ;
  assign n13884 = ~n13878 & n13883 ;
  assign n13885 = ~n13877 & n13884 ;
  assign n13892 = n8592 & ~n13599 ;
  assign n13887 = ~n7933 & ~n8641 ;
  assign n13888 = \P1_P1_InstQueue_reg[6][5]/NET0131  & ~n8640 ;
  assign n13889 = ~n8616 & n13888 ;
  assign n13890 = ~n13887 & ~n13889 ;
  assign n13891 = ~n8592 & n13890 ;
  assign n13893 = ~n8568 & ~n13891 ;
  assign n13894 = ~n13892 & n13893 ;
  assign n13886 = n8568 & n13591 ;
  assign n13895 = \P1_P1_DataWidth_reg[1]/NET0131  & ~n13886 ;
  assign n13896 = ~n13894 & n13895 ;
  assign n13897 = ~\P1_P1_DataWidth_reg[1]/NET0131  & n13890 ;
  assign n13898 = n8282 & ~n13897 ;
  assign n13899 = ~n13896 & n13898 ;
  assign n13900 = n8287 & ~n13890 ;
  assign n13901 = n8640 & ~n13639 ;
  assign n13902 = ~n13888 & ~n13901 ;
  assign n13903 = n8350 & ~n13902 ;
  assign n13904 = \P1_P1_InstQueue_reg[6][5]/NET0131  & ~n8366 ;
  assign n13905 = ~n13903 & ~n13904 ;
  assign n13906 = ~n13900 & n13905 ;
  assign n13907 = ~n13899 & n13906 ;
  assign n13914 = n8616 & ~n13599 ;
  assign n13909 = ~n7933 & ~n8664 ;
  assign n13910 = \P1_P1_InstQueue_reg[7][5]/NET0131  & ~n8407 ;
  assign n13911 = ~n8640 & n13910 ;
  assign n13912 = ~n13909 & ~n13911 ;
  assign n13913 = ~n8616 & n13912 ;
  assign n13915 = ~n8592 & ~n13913 ;
  assign n13916 = ~n13914 & n13915 ;
  assign n13908 = n8592 & n13591 ;
  assign n13917 = \P1_P1_DataWidth_reg[1]/NET0131  & ~n13908 ;
  assign n13918 = ~n13916 & n13917 ;
  assign n13919 = ~\P1_P1_DataWidth_reg[1]/NET0131  & n13912 ;
  assign n13920 = n8282 & ~n13919 ;
  assign n13921 = ~n13918 & n13920 ;
  assign n13922 = n8287 & ~n13912 ;
  assign n13923 = n8407 & ~n13639 ;
  assign n13924 = ~n13910 & ~n13923 ;
  assign n13925 = n8350 & ~n13924 ;
  assign n13926 = \P1_P1_InstQueue_reg[7][5]/NET0131  & ~n8366 ;
  assign n13927 = ~n13925 & ~n13926 ;
  assign n13928 = ~n13922 & n13927 ;
  assign n13929 = ~n13921 & n13928 ;
  assign n13936 = n8640 & ~n13599 ;
  assign n13931 = ~n7933 & ~n8410 ;
  assign n13932 = \P1_P1_InstQueue_reg[8][5]/NET0131  & ~n8139 ;
  assign n13933 = ~n8407 & n13932 ;
  assign n13934 = ~n13931 & ~n13933 ;
  assign n13935 = ~n8640 & n13934 ;
  assign n13937 = ~n8616 & ~n13935 ;
  assign n13938 = ~n13936 & n13937 ;
  assign n13930 = n8616 & n13591 ;
  assign n13939 = \P1_P1_DataWidth_reg[1]/NET0131  & ~n13930 ;
  assign n13940 = ~n13938 & n13939 ;
  assign n13941 = ~\P1_P1_DataWidth_reg[1]/NET0131  & n13934 ;
  assign n13942 = n8282 & ~n13941 ;
  assign n13943 = ~n13940 & n13942 ;
  assign n13944 = n8287 & ~n13934 ;
  assign n13945 = n8139 & ~n13639 ;
  assign n13946 = ~n13932 & ~n13945 ;
  assign n13947 = n8350 & ~n13946 ;
  assign n13948 = \P1_P1_InstQueue_reg[8][5]/NET0131  & ~n8366 ;
  assign n13949 = ~n13947 & ~n13948 ;
  assign n13950 = ~n13944 & n13949 ;
  assign n13951 = ~n13943 & n13950 ;
  assign n13958 = n8407 & ~n13599 ;
  assign n13953 = ~n7933 & ~n8709 ;
  assign n13954 = \P1_P1_InstQueue_reg[9][5]/NET0131  & ~n4327 ;
  assign n13955 = ~n8139 & n13954 ;
  assign n13956 = ~n13953 & ~n13955 ;
  assign n13957 = ~n8407 & n13956 ;
  assign n13959 = ~n8640 & ~n13957 ;
  assign n13960 = ~n13958 & n13959 ;
  assign n13952 = n8640 & n13591 ;
  assign n13961 = \P1_P1_DataWidth_reg[1]/NET0131  & ~n13952 ;
  assign n13962 = ~n13960 & n13961 ;
  assign n13963 = ~\P1_P1_DataWidth_reg[1]/NET0131  & n13956 ;
  assign n13964 = n8282 & ~n13963 ;
  assign n13965 = ~n13962 & n13964 ;
  assign n13966 = n8287 & ~n13956 ;
  assign n13967 = n4327 & ~n13639 ;
  assign n13968 = ~n13954 & ~n13967 ;
  assign n13969 = n8350 & ~n13968 ;
  assign n13970 = \P1_P1_InstQueue_reg[9][5]/NET0131  & ~n8366 ;
  assign n13971 = ~n13969 & ~n13970 ;
  assign n13972 = ~n13966 & n13971 ;
  assign n13973 = ~n13965 & n13972 ;
  assign n13980 = ~n8178 & n8190 ;
  assign n13981 = ~n8191 & ~n13980 ;
  assign n13982 = n8139 & ~n13981 ;
  assign n13983 = ~n8040 & n8052 ;
  assign n13984 = ~n8053 & ~n13983 ;
  assign n13985 = ~n8139 & ~n13984 ;
  assign n13986 = ~n13982 & ~n13985 ;
  assign n13987 = n10057 & ~n13986 ;
  assign n13974 = n7920 & ~n8146 ;
  assign n13975 = \P1_P1_InstQueue_reg[11][1]/NET0131  & ~n8142 ;
  assign n13976 = ~n8145 & n13975 ;
  assign n13977 = ~n13974 & ~n13976 ;
  assign n13979 = ~n10057 & n13977 ;
  assign n13988 = n8282 & ~n13979 ;
  assign n13989 = ~n13987 & n13988 ;
  assign n13990 = \P1_P1_InstQueue_reg[14][1]/NET0131  & n8291 ;
  assign n13991 = \P1_P1_InstQueue_reg[3][1]/NET0131  & n8323 ;
  assign n13992 = \P1_P1_InstQueue_reg[8][1]/NET0131  & n8305 ;
  assign n14006 = ~n13991 & ~n13992 ;
  assign n13993 = \P1_P1_InstQueue_reg[12][1]/NET0131  & n8329 ;
  assign n13994 = \P1_P1_InstQueue_reg[13][1]/NET0131  & n8327 ;
  assign n14007 = ~n13993 & ~n13994 ;
  assign n14016 = n14006 & n14007 ;
  assign n14017 = ~n13990 & n14016 ;
  assign n14005 = \P1_P1_InstQueue_reg[2][1]/NET0131  & n8314 ;
  assign n14003 = \P1_P1_InstQueue_reg[4][1]/NET0131  & n8295 ;
  assign n14004 = \P1_P1_InstQueue_reg[0][1]/NET0131  & n8309 ;
  assign n14012 = ~n14003 & ~n14004 ;
  assign n14013 = ~n14005 & n14012 ;
  assign n13999 = \P1_P1_InstQueue_reg[6][1]/NET0131  & n8316 ;
  assign n14000 = \P1_P1_InstQueue_reg[7][1]/NET0131  & n8318 ;
  assign n14010 = ~n13999 & ~n14000 ;
  assign n14001 = \P1_P1_InstQueue_reg[15][1]/NET0131  & n8321 ;
  assign n14002 = \P1_P1_InstQueue_reg[11][1]/NET0131  & n8312 ;
  assign n14011 = ~n14001 & ~n14002 ;
  assign n14014 = n14010 & n14011 ;
  assign n13995 = \P1_P1_InstQueue_reg[9][1]/NET0131  & n8325 ;
  assign n13996 = \P1_P1_InstQueue_reg[5][1]/NET0131  & n8307 ;
  assign n14008 = ~n13995 & ~n13996 ;
  assign n13997 = \P1_P1_InstQueue_reg[1][1]/NET0131  & n8299 ;
  assign n13998 = \P1_P1_InstQueue_reg[10][1]/NET0131  & n8303 ;
  assign n14009 = ~n13997 & ~n13998 ;
  assign n14015 = n14008 & n14009 ;
  assign n14018 = n14014 & n14015 ;
  assign n14019 = n14013 & n14018 ;
  assign n14020 = n14017 & n14019 ;
  assign n14021 = n8142 & ~n14020 ;
  assign n14022 = ~n13975 & ~n14021 ;
  assign n14023 = n8350 & ~n14022 ;
  assign n13978 = n8287 & ~n13977 ;
  assign n14024 = \P1_P1_InstQueue_reg[11][1]/NET0131  & ~n8366 ;
  assign n14025 = ~n13978 & ~n14024 ;
  assign n14026 = ~n14023 & n14025 ;
  assign n14027 = ~n13989 & n14026 ;
  assign n14031 = ~n11345 & ~n11580 ;
  assign n14032 = ~n11581 & ~n14031 ;
  assign n14033 = ~n10105 & ~n14032 ;
  assign n14028 = ~n11484 & n11504 ;
  assign n14029 = ~n11505 & ~n14028 ;
  assign n14030 = n10105 & ~n14029 ;
  assign n14034 = n12334 & ~n14030 ;
  assign n14035 = ~n14033 & n14034 ;
  assign n14043 = \P2_P1_InstQueue_reg[6][2]/NET0131  & n11651 ;
  assign n14042 = \P2_P1_InstQueue_reg[15][2]/NET0131  & n11647 ;
  assign n14038 = \P2_P1_InstQueue_reg[11][2]/NET0131  & n11665 ;
  assign n14039 = \P2_P1_InstQueue_reg[13][2]/NET0131  & n11641 ;
  assign n14054 = ~n14038 & ~n14039 ;
  assign n14064 = ~n14042 & n14054 ;
  assign n14065 = ~n14043 & n14064 ;
  assign n14050 = \P2_P1_InstQueue_reg[0][2]/NET0131  & n11669 ;
  assign n14051 = \P2_P1_InstQueue_reg[9][2]/NET0131  & n11656 ;
  assign n14059 = ~n14050 & ~n14051 ;
  assign n14052 = \P2_P1_InstQueue_reg[2][2]/NET0131  & n11654 ;
  assign n14053 = \P2_P1_InstQueue_reg[4][2]/NET0131  & n11667 ;
  assign n14060 = ~n14052 & ~n14053 ;
  assign n14061 = n14059 & n14060 ;
  assign n14046 = \P2_P1_InstQueue_reg[5][2]/NET0131  & n11638 ;
  assign n14047 = \P2_P1_InstQueue_reg[7][2]/NET0131  & n11661 ;
  assign n14057 = ~n14046 & ~n14047 ;
  assign n14048 = \P2_P1_InstQueue_reg[12][2]/NET0131  & n11673 ;
  assign n14049 = \P2_P1_InstQueue_reg[8][2]/NET0131  & n11659 ;
  assign n14058 = ~n14048 & ~n14049 ;
  assign n14062 = n14057 & n14058 ;
  assign n14040 = \P2_P1_InstQueue_reg[10][2]/NET0131  & n11634 ;
  assign n14041 = \P2_P1_InstQueue_reg[14][2]/NET0131  & n11643 ;
  assign n14055 = ~n14040 & ~n14041 ;
  assign n14044 = \P2_P1_InstQueue_reg[1][2]/NET0131  & n11671 ;
  assign n14045 = \P2_P1_InstQueue_reg[3][2]/NET0131  & n11663 ;
  assign n14056 = ~n14044 & ~n14045 ;
  assign n14063 = n14055 & n14056 ;
  assign n14066 = n14062 & n14063 ;
  assign n14067 = n14061 & n14066 ;
  assign n14068 = n14065 & n14067 ;
  assign n14069 = n11596 & n14068 ;
  assign n14037 = ~\P2_P1_InstQueue_reg[11][2]/NET0131  & ~n11596 ;
  assign n14070 = n11692 & ~n14037 ;
  assign n14071 = ~n14069 & n14070 ;
  assign n14036 = \P2_P1_InstQueue_reg[11][2]/NET0131  & ~n12345 ;
  assign n14072 = n11382 & ~n11600 ;
  assign n14073 = n12343 & n14072 ;
  assign n14074 = ~n14036 & ~n14073 ;
  assign n14075 = ~n14071 & n14074 ;
  assign n14076 = ~n14035 & n14075 ;
  assign n14083 = n8375 & ~n13981 ;
  assign n14084 = ~n8375 & ~n13984 ;
  assign n14085 = ~n14083 & ~n14084 ;
  assign n14086 = n11707 & ~n14085 ;
  assign n14077 = n7920 & ~n8379 ;
  assign n14078 = \P1_P1_InstQueue_reg[0][1]/NET0131  & ~n8376 ;
  assign n14079 = ~n8378 & n14078 ;
  assign n14080 = ~n14077 & ~n14079 ;
  assign n14082 = ~n11707 & n14080 ;
  assign n14087 = n8282 & ~n14082 ;
  assign n14088 = ~n14086 & n14087 ;
  assign n14089 = n8376 & ~n14020 ;
  assign n14090 = ~n14078 & ~n14089 ;
  assign n14091 = n8350 & ~n14090 ;
  assign n14081 = n8287 & ~n14080 ;
  assign n14092 = \P1_P1_InstQueue_reg[0][1]/NET0131  & ~n8366 ;
  assign n14093 = ~n14081 & ~n14092 ;
  assign n14094 = ~n14091 & n14093 ;
  assign n14095 = ~n14088 & n14094 ;
  assign n14102 = n8407 & ~n13981 ;
  assign n14103 = ~n8407 & ~n13984 ;
  assign n14104 = ~n14102 & ~n14103 ;
  assign n14105 = n9418 & ~n14104 ;
  assign n14096 = n7920 & ~n8401 ;
  assign n14097 = \P1_P1_InstQueue_reg[10][1]/NET0131  & ~n8145 ;
  assign n14098 = ~n4327 & n14097 ;
  assign n14099 = ~n14096 & ~n14098 ;
  assign n14101 = ~n9418 & n14099 ;
  assign n14106 = n8282 & ~n14101 ;
  assign n14107 = ~n14105 & n14106 ;
  assign n14108 = n8145 & ~n14020 ;
  assign n14109 = ~n14097 & ~n14108 ;
  assign n14110 = n8350 & ~n14109 ;
  assign n14100 = n8287 & ~n14099 ;
  assign n14111 = \P1_P1_InstQueue_reg[10][1]/NET0131  & ~n8366 ;
  assign n14112 = ~n14100 & ~n14111 ;
  assign n14113 = ~n14110 & n14112 ;
  assign n14114 = ~n14107 & n14113 ;
  assign n14121 = n4327 & ~n13981 ;
  assign n14122 = ~n4327 & ~n13984 ;
  assign n14123 = ~n14121 & ~n14122 ;
  assign n14124 = n11746 & ~n14123 ;
  assign n14115 = n7920 & ~n8428 ;
  assign n14116 = \P1_P1_InstQueue_reg[12][1]/NET0131  & ~n8427 ;
  assign n14117 = ~n8142 & n14116 ;
  assign n14118 = ~n14115 & ~n14117 ;
  assign n14120 = ~n11746 & n14118 ;
  assign n14125 = n8282 & ~n14120 ;
  assign n14126 = ~n14124 & n14125 ;
  assign n14127 = n8427 & ~n14020 ;
  assign n14128 = ~n14116 & ~n14127 ;
  assign n14129 = n8350 & ~n14128 ;
  assign n14119 = n8287 & ~n14118 ;
  assign n14130 = \P1_P1_InstQueue_reg[12][1]/NET0131  & ~n8366 ;
  assign n14131 = ~n14119 & ~n14130 ;
  assign n14132 = ~n14129 & n14131 ;
  assign n14133 = ~n14126 & n14132 ;
  assign n14140 = n8145 & ~n13981 ;
  assign n14141 = ~n8145 & ~n13984 ;
  assign n14142 = ~n14140 & ~n14141 ;
  assign n14143 = n11766 & ~n14142 ;
  assign n14134 = n7920 & ~n8451 ;
  assign n14135 = \P1_P1_InstQueue_reg[13][1]/NET0131  & ~n8375 ;
  assign n14136 = ~n8427 & n14135 ;
  assign n14137 = ~n14134 & ~n14136 ;
  assign n14139 = ~n11766 & n14137 ;
  assign n14144 = n8282 & ~n14139 ;
  assign n14145 = ~n14143 & n14144 ;
  assign n14146 = n8375 & ~n14020 ;
  assign n14147 = ~n14135 & ~n14146 ;
  assign n14148 = n8350 & ~n14147 ;
  assign n14138 = n8287 & ~n14137 ;
  assign n14149 = \P1_P1_InstQueue_reg[13][1]/NET0131  & ~n8366 ;
  assign n14150 = ~n14138 & ~n14149 ;
  assign n14151 = ~n14148 & n14150 ;
  assign n14152 = ~n14145 & n14151 ;
  assign n14159 = n8142 & ~n13981 ;
  assign n14160 = ~n8142 & ~n13984 ;
  assign n14161 = ~n14159 & ~n14160 ;
  assign n14162 = n11786 & ~n14161 ;
  assign n14153 = n7920 & ~n8474 ;
  assign n14154 = \P1_P1_InstQueue_reg[14][1]/NET0131  & ~n8372 ;
  assign n14155 = ~n8375 & n14154 ;
  assign n14156 = ~n14153 & ~n14155 ;
  assign n14158 = ~n11786 & n14156 ;
  assign n14163 = n8282 & ~n14158 ;
  assign n14164 = ~n14162 & n14163 ;
  assign n14165 = n8372 & ~n14020 ;
  assign n14166 = ~n14154 & ~n14165 ;
  assign n14167 = n8350 & ~n14166 ;
  assign n14157 = n8287 & ~n14156 ;
  assign n14168 = \P1_P1_InstQueue_reg[14][1]/NET0131  & ~n8366 ;
  assign n14169 = ~n14157 & ~n14168 ;
  assign n14170 = ~n14167 & n14169 ;
  assign n14171 = ~n14164 & n14170 ;
  assign n14178 = n8427 & ~n13981 ;
  assign n14179 = ~n8427 & ~n13984 ;
  assign n14180 = ~n14178 & ~n14179 ;
  assign n14181 = n11806 & ~n14180 ;
  assign n14172 = n7920 & ~n8497 ;
  assign n14173 = \P1_P1_InstQueue_reg[15][1]/NET0131  & ~n8378 ;
  assign n14174 = ~n8372 & n14173 ;
  assign n14175 = ~n14172 & ~n14174 ;
  assign n14177 = ~n11806 & n14175 ;
  assign n14182 = n8282 & ~n14177 ;
  assign n14183 = ~n14181 & n14182 ;
  assign n14184 = n8378 & ~n14020 ;
  assign n14185 = ~n14173 & ~n14184 ;
  assign n14186 = n8350 & ~n14185 ;
  assign n14176 = n8287 & ~n14175 ;
  assign n14187 = \P1_P1_InstQueue_reg[15][1]/NET0131  & ~n8366 ;
  assign n14188 = ~n14176 & ~n14187 ;
  assign n14189 = ~n14186 & n14188 ;
  assign n14190 = ~n14183 & n14189 ;
  assign n14197 = n8372 & ~n13981 ;
  assign n14198 = ~n8372 & ~n13984 ;
  assign n14199 = ~n14197 & ~n14198 ;
  assign n14200 = n11826 & ~n14199 ;
  assign n14191 = n7920 & ~n8521 ;
  assign n14192 = \P1_P1_InstQueue_reg[1][1]/NET0131  & ~n8520 ;
  assign n14193 = ~n8376 & n14192 ;
  assign n14194 = ~n14191 & ~n14193 ;
  assign n14196 = ~n11826 & n14194 ;
  assign n14201 = n8282 & ~n14196 ;
  assign n14202 = ~n14200 & n14201 ;
  assign n14203 = n8520 & ~n14020 ;
  assign n14204 = ~n14192 & ~n14203 ;
  assign n14205 = n8350 & ~n14204 ;
  assign n14195 = n8287 & ~n14194 ;
  assign n14206 = \P1_P1_InstQueue_reg[1][1]/NET0131  & ~n8366 ;
  assign n14207 = ~n14195 & ~n14206 ;
  assign n14208 = ~n14205 & n14207 ;
  assign n14209 = ~n14202 & n14208 ;
  assign n14216 = n8378 & ~n13981 ;
  assign n14217 = ~n8378 & ~n13984 ;
  assign n14218 = ~n14216 & ~n14217 ;
  assign n14219 = n11846 & ~n14218 ;
  assign n14210 = n7920 & ~n8545 ;
  assign n14211 = \P1_P1_InstQueue_reg[2][1]/NET0131  & ~n8544 ;
  assign n14212 = ~n8520 & n14211 ;
  assign n14213 = ~n14210 & ~n14212 ;
  assign n14215 = ~n11846 & n14213 ;
  assign n14220 = n8282 & ~n14215 ;
  assign n14221 = ~n14219 & n14220 ;
  assign n14222 = n8544 & ~n14020 ;
  assign n14223 = ~n14211 & ~n14222 ;
  assign n14224 = n8350 & ~n14223 ;
  assign n14214 = n8287 & ~n14213 ;
  assign n14225 = \P1_P1_InstQueue_reg[2][1]/NET0131  & ~n8366 ;
  assign n14226 = ~n14214 & ~n14225 ;
  assign n14227 = ~n14224 & n14226 ;
  assign n14228 = ~n14221 & n14227 ;
  assign n14230 = ~n11862 & ~n14032 ;
  assign n14229 = n11862 & ~n14029 ;
  assign n14231 = n12388 & ~n14229 ;
  assign n14232 = ~n14230 & n14231 ;
  assign n14235 = n11871 & n14068 ;
  assign n14234 = ~\P2_P1_InstQueue_reg[0][2]/NET0131  & ~n11871 ;
  assign n14236 = n11692 & ~n14234 ;
  assign n14237 = ~n14235 & n14236 ;
  assign n14233 = \P2_P1_InstQueue_reg[0][2]/NET0131  & ~n12395 ;
  assign n14238 = n11382 & ~n11874 ;
  assign n14239 = n12393 & n14238 ;
  assign n14240 = ~n14233 & ~n14239 ;
  assign n14241 = ~n14237 & n14240 ;
  assign n14242 = ~n14232 & n14241 ;
  assign n14244 = ~n11891 & ~n14032 ;
  assign n14243 = n11891 & ~n14029 ;
  assign n14245 = n12407 & ~n14243 ;
  assign n14246 = ~n14244 & n14245 ;
  assign n14249 = n11599 & n14068 ;
  assign n14248 = ~\P2_P1_InstQueue_reg[10][2]/NET0131  & ~n11599 ;
  assign n14250 = n11692 & ~n14248 ;
  assign n14251 = ~n14249 & n14250 ;
  assign n14247 = \P2_P1_InstQueue_reg[10][2]/NET0131  & ~n12414 ;
  assign n14252 = n11382 & ~n11897 ;
  assign n14253 = n12412 & n14252 ;
  assign n14254 = ~n14247 & ~n14253 ;
  assign n14255 = ~n14251 & n14254 ;
  assign n14256 = ~n14246 & n14255 ;
  assign n14263 = n8376 & ~n13981 ;
  assign n14264 = ~n8376 & ~n13984 ;
  assign n14265 = ~n14263 & ~n14264 ;
  assign n14266 = n11941 & ~n14265 ;
  assign n14257 = n7920 & ~n8569 ;
  assign n14258 = \P1_P1_InstQueue_reg[3][1]/NET0131  & ~n8568 ;
  assign n14259 = ~n8544 & n14258 ;
  assign n14260 = ~n14257 & ~n14259 ;
  assign n14262 = ~n11941 & n14260 ;
  assign n14267 = n8282 & ~n14262 ;
  assign n14268 = ~n14266 & n14267 ;
  assign n14269 = n8568 & ~n14020 ;
  assign n14270 = ~n14258 & ~n14269 ;
  assign n14271 = n8350 & ~n14270 ;
  assign n14261 = n8287 & ~n14260 ;
  assign n14272 = \P1_P1_InstQueue_reg[3][1]/NET0131  & ~n8366 ;
  assign n14273 = ~n14261 & ~n14272 ;
  assign n14274 = ~n14271 & n14273 ;
  assign n14275 = ~n14268 & n14274 ;
  assign n14277 = ~n11577 & ~n14032 ;
  assign n14276 = n11577 & ~n14029 ;
  assign n14278 = n12426 & ~n14276 ;
  assign n14279 = ~n14277 & n14278 ;
  assign n14282 = n11919 & n14068 ;
  assign n14281 = ~\P2_P1_InstQueue_reg[12][2]/NET0131  & ~n11919 ;
  assign n14283 = n11692 & ~n14281 ;
  assign n14284 = ~n14282 & n14283 ;
  assign n14280 = \P2_P1_InstQueue_reg[12][2]/NET0131  & ~n12433 ;
  assign n14285 = n11382 & ~n11920 ;
  assign n14286 = n12431 & n14285 ;
  assign n14287 = ~n14280 & ~n14286 ;
  assign n14288 = ~n14284 & n14287 ;
  assign n14289 = ~n14279 & n14288 ;
  assign n14291 = ~n11599 & ~n14032 ;
  assign n14290 = n11599 & ~n14029 ;
  assign n14292 = n12445 & ~n14290 ;
  assign n14293 = ~n14291 & n14292 ;
  assign n14296 = n11862 & n14068 ;
  assign n14295 = ~\P2_P1_InstQueue_reg[13][2]/NET0131  & ~n11862 ;
  assign n14297 = n11692 & ~n14295 ;
  assign n14298 = ~n14296 & n14297 ;
  assign n14294 = \P2_P1_InstQueue_reg[13][2]/NET0131  & ~n12452 ;
  assign n14299 = n11382 & ~n11961 ;
  assign n14300 = n12450 & n14299 ;
  assign n14301 = ~n14294 & ~n14300 ;
  assign n14302 = ~n14298 & n14301 ;
  assign n14303 = ~n14293 & n14302 ;
  assign n14305 = ~n11596 & ~n14032 ;
  assign n14304 = n11596 & ~n14029 ;
  assign n14306 = n12464 & ~n14304 ;
  assign n14307 = ~n14305 & n14306 ;
  assign n14310 = n11865 & n14068 ;
  assign n14309 = ~\P2_P1_InstQueue_reg[14][2]/NET0131  & ~n11865 ;
  assign n14311 = n11692 & ~n14309 ;
  assign n14312 = ~n14310 & n14311 ;
  assign n14308 = \P2_P1_InstQueue_reg[14][2]/NET0131  & ~n12471 ;
  assign n14313 = n11382 & ~n11869 ;
  assign n14314 = n12469 & n14313 ;
  assign n14315 = ~n14308 & ~n14314 ;
  assign n14316 = ~n14312 & n14315 ;
  assign n14317 = ~n14307 & n14316 ;
  assign n14319 = ~n11919 & ~n14032 ;
  assign n14318 = n11919 & ~n14029 ;
  assign n14320 = n12483 & ~n14318 ;
  assign n14321 = ~n14319 & n14320 ;
  assign n14324 = n11873 & n14068 ;
  assign n14323 = ~\P2_P1_InstQueue_reg[15][2]/NET0131  & ~n11873 ;
  assign n14325 = n11692 & ~n14323 ;
  assign n14326 = ~n14324 & n14325 ;
  assign n14322 = \P2_P1_InstQueue_reg[15][2]/NET0131  & ~n12490 ;
  assign n14327 = n11382 & ~n12002 ;
  assign n14328 = n12488 & n14327 ;
  assign n14329 = ~n14322 & ~n14328 ;
  assign n14330 = ~n14326 & n14329 ;
  assign n14331 = ~n14321 & n14330 ;
  assign n14333 = ~n11865 & ~n14032 ;
  assign n14332 = n11865 & ~n14029 ;
  assign n14334 = n12502 & ~n14332 ;
  assign n14335 = ~n14333 & n14334 ;
  assign n14338 = n12023 & n14068 ;
  assign n14337 = ~\P2_P1_InstQueue_reg[1][2]/NET0131  & ~n12023 ;
  assign n14339 = n11692 & ~n14337 ;
  assign n14340 = ~n14338 & n14339 ;
  assign n14336 = \P2_P1_InstQueue_reg[1][2]/NET0131  & ~n12509 ;
  assign n14341 = n11382 & ~n12024 ;
  assign n14342 = n12507 & n14341 ;
  assign n14343 = ~n14336 & ~n14342 ;
  assign n14344 = ~n14340 & n14343 ;
  assign n14345 = ~n14335 & n14344 ;
  assign n14352 = n8520 & ~n13981 ;
  assign n14353 = ~n8520 & ~n13984 ;
  assign n14354 = ~n14352 & ~n14353 ;
  assign n14355 = n12045 & ~n14354 ;
  assign n14346 = n7920 & ~n8593 ;
  assign n14347 = \P1_P1_InstQueue_reg[4][1]/NET0131  & ~n8592 ;
  assign n14348 = ~n8568 & n14347 ;
  assign n14349 = ~n14346 & ~n14348 ;
  assign n14351 = ~n12045 & n14349 ;
  assign n14356 = n8282 & ~n14351 ;
  assign n14357 = ~n14355 & n14356 ;
  assign n14358 = n8592 & ~n14020 ;
  assign n14359 = ~n14347 & ~n14358 ;
  assign n14360 = n8350 & ~n14359 ;
  assign n14350 = n8287 & ~n14349 ;
  assign n14361 = \P1_P1_InstQueue_reg[4][1]/NET0131  & ~n8366 ;
  assign n14362 = ~n14350 & ~n14361 ;
  assign n14363 = ~n14360 & n14362 ;
  assign n14364 = ~n14357 & n14363 ;
  assign n14366 = ~n11873 & ~n14032 ;
  assign n14365 = n11873 & ~n14029 ;
  assign n14367 = n12521 & ~n14365 ;
  assign n14368 = ~n14366 & n14367 ;
  assign n14371 = n12065 & n14068 ;
  assign n14370 = ~\P2_P1_InstQueue_reg[2][2]/NET0131  & ~n12065 ;
  assign n14372 = n11692 & ~n14370 ;
  assign n14373 = ~n14371 & n14372 ;
  assign n14369 = \P2_P1_InstQueue_reg[2][2]/NET0131  & ~n12528 ;
  assign n14374 = n11382 & ~n12066 ;
  assign n14375 = n12526 & n14374 ;
  assign n14376 = ~n14369 & ~n14375 ;
  assign n14377 = ~n14373 & n14376 ;
  assign n14378 = ~n14368 & n14377 ;
  assign n14380 = ~n11871 & ~n14032 ;
  assign n14379 = n11871 & ~n14029 ;
  assign n14381 = n12540 & ~n14379 ;
  assign n14382 = ~n14380 & n14381 ;
  assign n14385 = n12087 & n14068 ;
  assign n14384 = ~\P2_P1_InstQueue_reg[3][2]/NET0131  & ~n12087 ;
  assign n14386 = n11692 & ~n14384 ;
  assign n14387 = ~n14385 & n14386 ;
  assign n14383 = \P2_P1_InstQueue_reg[3][2]/NET0131  & ~n12547 ;
  assign n14388 = n11382 & ~n12088 ;
  assign n14389 = n12545 & n14388 ;
  assign n14390 = ~n14383 & ~n14389 ;
  assign n14391 = ~n14387 & n14390 ;
  assign n14392 = ~n14382 & n14391 ;
  assign n14394 = ~n12023 & ~n14032 ;
  assign n14393 = n12023 & ~n14029 ;
  assign n14395 = n12559 & ~n14393 ;
  assign n14396 = ~n14394 & n14395 ;
  assign n14399 = n12109 & n14068 ;
  assign n14398 = ~\P2_P1_InstQueue_reg[4][2]/NET0131  & ~n12109 ;
  assign n14400 = n11692 & ~n14398 ;
  assign n14401 = ~n14399 & n14400 ;
  assign n14397 = \P2_P1_InstQueue_reg[4][2]/NET0131  & ~n12566 ;
  assign n14402 = n11382 & ~n12110 ;
  assign n14403 = n12564 & n14402 ;
  assign n14404 = ~n14397 & ~n14403 ;
  assign n14405 = ~n14401 & n14404 ;
  assign n14406 = ~n14396 & n14405 ;
  assign n14408 = ~n12065 & ~n14032 ;
  assign n14407 = n12065 & ~n14029 ;
  assign n14409 = n12578 & ~n14407 ;
  assign n14410 = ~n14408 & n14409 ;
  assign n14413 = n12131 & n14068 ;
  assign n14412 = ~\P2_P1_InstQueue_reg[5][2]/NET0131  & ~n12131 ;
  assign n14414 = n11692 & ~n14412 ;
  assign n14415 = ~n14413 & n14414 ;
  assign n14411 = \P2_P1_InstQueue_reg[5][2]/NET0131  & ~n12585 ;
  assign n14416 = n11382 & ~n12132 ;
  assign n14417 = n12583 & n14416 ;
  assign n14418 = ~n14411 & ~n14417 ;
  assign n14419 = ~n14415 & n14418 ;
  assign n14420 = ~n14410 & n14419 ;
  assign n14427 = n8544 & ~n13981 ;
  assign n14428 = ~n8544 & ~n13984 ;
  assign n14429 = ~n14427 & ~n14428 ;
  assign n14430 = n12153 & ~n14429 ;
  assign n14421 = n7920 & ~n8617 ;
  assign n14422 = \P1_P1_InstQueue_reg[5][1]/NET0131  & ~n8616 ;
  assign n14423 = ~n8592 & n14422 ;
  assign n14424 = ~n14421 & ~n14423 ;
  assign n14426 = ~n12153 & n14424 ;
  assign n14431 = n8282 & ~n14426 ;
  assign n14432 = ~n14430 & n14431 ;
  assign n14433 = n8616 & ~n14020 ;
  assign n14434 = ~n14422 & ~n14433 ;
  assign n14435 = n8350 & ~n14434 ;
  assign n14425 = n8287 & ~n14424 ;
  assign n14436 = \P1_P1_InstQueue_reg[5][1]/NET0131  & ~n8366 ;
  assign n14437 = ~n14425 & ~n14436 ;
  assign n14438 = ~n14435 & n14437 ;
  assign n14439 = ~n14432 & n14438 ;
  assign n14441 = ~n12087 & ~n14032 ;
  assign n14440 = n12087 & ~n14029 ;
  assign n14442 = n12597 & ~n14440 ;
  assign n14443 = ~n14441 & n14442 ;
  assign n14446 = n12173 & n14068 ;
  assign n14445 = ~\P2_P1_InstQueue_reg[6][2]/NET0131  & ~n12173 ;
  assign n14447 = n11692 & ~n14445 ;
  assign n14448 = ~n14446 & n14447 ;
  assign n14444 = \P2_P1_InstQueue_reg[6][2]/NET0131  & ~n12604 ;
  assign n14449 = n11382 & ~n12174 ;
  assign n14450 = n12602 & n14449 ;
  assign n14451 = ~n14444 & ~n14450 ;
  assign n14452 = ~n14448 & n14451 ;
  assign n14453 = ~n14443 & n14452 ;
  assign n14455 = ~n12109 & ~n14032 ;
  assign n14454 = n12109 & ~n14029 ;
  assign n14456 = n12616 & ~n14454 ;
  assign n14457 = ~n14455 & n14456 ;
  assign n14460 = n11891 & n14068 ;
  assign n14459 = ~\P2_P1_InstQueue_reg[7][2]/NET0131  & ~n11891 ;
  assign n14461 = n11692 & ~n14459 ;
  assign n14462 = ~n14460 & n14461 ;
  assign n14458 = \P2_P1_InstQueue_reg[7][2]/NET0131  & ~n12623 ;
  assign n14463 = n11382 & ~n12195 ;
  assign n14464 = n12621 & n14463 ;
  assign n14465 = ~n14458 & ~n14464 ;
  assign n14466 = ~n14462 & n14465 ;
  assign n14467 = ~n14457 & n14466 ;
  assign n14469 = ~n12131 & ~n14032 ;
  assign n14468 = n12131 & ~n14029 ;
  assign n14470 = n12635 & ~n14468 ;
  assign n14471 = ~n14469 & n14470 ;
  assign n14474 = n10105 & n14068 ;
  assign n14473 = ~\P2_P1_InstQueue_reg[8][2]/NET0131  & ~n10105 ;
  assign n14475 = n11692 & ~n14473 ;
  assign n14476 = ~n14474 & n14475 ;
  assign n14472 = \P2_P1_InstQueue_reg[8][2]/NET0131  & ~n12642 ;
  assign n14477 = n11382 & ~n11895 ;
  assign n14478 = n12640 & n14477 ;
  assign n14479 = ~n14472 & ~n14478 ;
  assign n14480 = ~n14476 & n14479 ;
  assign n14481 = ~n14471 & n14480 ;
  assign n14483 = ~n12173 & ~n14032 ;
  assign n14482 = n12173 & ~n14029 ;
  assign n14484 = n12654 & ~n14482 ;
  assign n14485 = ~n14483 & n14484 ;
  assign n14488 = n11577 & n14068 ;
  assign n14487 = ~\P2_P1_InstQueue_reg[9][2]/NET0131  & ~n11577 ;
  assign n14489 = n11692 & ~n14487 ;
  assign n14490 = ~n14488 & n14489 ;
  assign n14486 = \P2_P1_InstQueue_reg[9][2]/NET0131  & ~n12661 ;
  assign n14491 = n11382 & ~n11592 ;
  assign n14492 = n12659 & n14491 ;
  assign n14493 = ~n14486 & ~n14492 ;
  assign n14494 = ~n14490 & n14493 ;
  assign n14495 = ~n14485 & n14494 ;
  assign n14502 = n8568 & ~n13981 ;
  assign n14503 = ~n8568 & ~n13984 ;
  assign n14504 = ~n14502 & ~n14503 ;
  assign n14505 = n12256 & ~n14504 ;
  assign n14496 = n7920 & ~n8641 ;
  assign n14497 = \P1_P1_InstQueue_reg[6][1]/NET0131  & ~n8640 ;
  assign n14498 = ~n8616 & n14497 ;
  assign n14499 = ~n14496 & ~n14498 ;
  assign n14501 = ~n12256 & n14499 ;
  assign n14506 = n8282 & ~n14501 ;
  assign n14507 = ~n14505 & n14506 ;
  assign n14508 = n8640 & ~n14020 ;
  assign n14509 = ~n14497 & ~n14508 ;
  assign n14510 = n8350 & ~n14509 ;
  assign n14500 = n8287 & ~n14499 ;
  assign n14511 = \P1_P1_InstQueue_reg[6][1]/NET0131  & ~n8366 ;
  assign n14512 = ~n14500 & ~n14511 ;
  assign n14513 = ~n14510 & n14512 ;
  assign n14514 = ~n14507 & n14513 ;
  assign n14521 = n8592 & ~n13981 ;
  assign n14522 = ~n8592 & ~n13984 ;
  assign n14523 = ~n14521 & ~n14522 ;
  assign n14524 = n12276 & ~n14523 ;
  assign n14515 = n7920 & ~n8664 ;
  assign n14516 = \P1_P1_InstQueue_reg[7][1]/NET0131  & ~n8407 ;
  assign n14517 = ~n8640 & n14516 ;
  assign n14518 = ~n14515 & ~n14517 ;
  assign n14520 = ~n12276 & n14518 ;
  assign n14525 = n8282 & ~n14520 ;
  assign n14526 = ~n14524 & n14525 ;
  assign n14527 = n8407 & ~n14020 ;
  assign n14528 = ~n14516 & ~n14527 ;
  assign n14529 = n8350 & ~n14528 ;
  assign n14519 = n8287 & ~n14518 ;
  assign n14530 = \P1_P1_InstQueue_reg[7][1]/NET0131  & ~n8366 ;
  assign n14531 = ~n14519 & ~n14530 ;
  assign n14532 = ~n14529 & n14531 ;
  assign n14533 = ~n14526 & n14532 ;
  assign n14540 = n8616 & ~n13981 ;
  assign n14541 = ~n8616 & ~n13984 ;
  assign n14542 = ~n14540 & ~n14541 ;
  assign n14543 = n12296 & ~n14542 ;
  assign n14534 = n7920 & ~n8410 ;
  assign n14535 = \P1_P1_InstQueue_reg[8][1]/NET0131  & ~n8139 ;
  assign n14536 = ~n8407 & n14535 ;
  assign n14537 = ~n14534 & ~n14536 ;
  assign n14539 = ~n12296 & n14537 ;
  assign n14544 = n8282 & ~n14539 ;
  assign n14545 = ~n14543 & n14544 ;
  assign n14546 = n8139 & ~n14020 ;
  assign n14547 = ~n14535 & ~n14546 ;
  assign n14548 = n8350 & ~n14547 ;
  assign n14538 = n8287 & ~n14537 ;
  assign n14549 = \P1_P1_InstQueue_reg[8][1]/NET0131  & ~n8366 ;
  assign n14550 = ~n14538 & ~n14549 ;
  assign n14551 = ~n14548 & n14550 ;
  assign n14552 = ~n14545 & n14551 ;
  assign n14559 = n8640 & ~n13981 ;
  assign n14560 = ~n8640 & ~n13984 ;
  assign n14561 = ~n14559 & ~n14560 ;
  assign n14562 = n12316 & ~n14561 ;
  assign n14553 = n7920 & ~n8709 ;
  assign n14554 = \P1_P1_InstQueue_reg[9][1]/NET0131  & ~n4327 ;
  assign n14555 = ~n8139 & n14554 ;
  assign n14556 = ~n14553 & ~n14555 ;
  assign n14558 = ~n12316 & n14556 ;
  assign n14563 = n8282 & ~n14558 ;
  assign n14564 = ~n14562 & n14563 ;
  assign n14565 = n4327 & ~n14020 ;
  assign n14566 = ~n14554 & ~n14565 ;
  assign n14567 = n8350 & ~n14566 ;
  assign n14557 = n8287 & ~n14556 ;
  assign n14568 = \P1_P1_InstQueue_reg[9][1]/NET0131  & ~n8366 ;
  assign n14569 = ~n14557 & ~n14568 ;
  assign n14570 = ~n14567 & n14569 ;
  assign n14571 = ~n14564 & n14570 ;
  assign n14575 = n11365 & ~n11583 ;
  assign n14576 = ~n11584 & ~n14575 ;
  assign n14577 = ~n10105 & ~n14576 ;
  assign n14572 = ~n11538 & n11553 ;
  assign n14573 = ~n11554 & ~n14572 ;
  assign n14574 = n10105 & ~n14573 ;
  assign n14578 = n12334 & ~n14574 ;
  assign n14579 = ~n14577 & n14578 ;
  assign n14587 = \P2_P1_InstQueue_reg[6][5]/NET0131  & n11651 ;
  assign n14586 = \P2_P1_InstQueue_reg[15][5]/NET0131  & n11647 ;
  assign n14582 = \P2_P1_InstQueue_reg[11][5]/NET0131  & n11665 ;
  assign n14583 = \P2_P1_InstQueue_reg[10][5]/NET0131  & n11634 ;
  assign n14598 = ~n14582 & ~n14583 ;
  assign n14608 = ~n14586 & n14598 ;
  assign n14609 = ~n14587 & n14608 ;
  assign n14594 = \P2_P1_InstQueue_reg[0][5]/NET0131  & n11669 ;
  assign n14595 = \P2_P1_InstQueue_reg[9][5]/NET0131  & n11656 ;
  assign n14603 = ~n14594 & ~n14595 ;
  assign n14596 = \P2_P1_InstQueue_reg[2][5]/NET0131  & n11654 ;
  assign n14597 = \P2_P1_InstQueue_reg[4][5]/NET0131  & n11667 ;
  assign n14604 = ~n14596 & ~n14597 ;
  assign n14605 = n14603 & n14604 ;
  assign n14590 = \P2_P1_InstQueue_reg[12][5]/NET0131  & n11673 ;
  assign n14591 = \P2_P1_InstQueue_reg[7][5]/NET0131  & n11661 ;
  assign n14601 = ~n14590 & ~n14591 ;
  assign n14592 = \P2_P1_InstQueue_reg[5][5]/NET0131  & n11638 ;
  assign n14593 = \P2_P1_InstQueue_reg[8][5]/NET0131  & n11659 ;
  assign n14602 = ~n14592 & ~n14593 ;
  assign n14606 = n14601 & n14602 ;
  assign n14584 = \P2_P1_InstQueue_reg[1][5]/NET0131  & n11671 ;
  assign n14585 = \P2_P1_InstQueue_reg[14][5]/NET0131  & n11643 ;
  assign n14599 = ~n14584 & ~n14585 ;
  assign n14588 = \P2_P1_InstQueue_reg[13][5]/NET0131  & n11641 ;
  assign n14589 = \P2_P1_InstQueue_reg[3][5]/NET0131  & n11663 ;
  assign n14600 = ~n14588 & ~n14589 ;
  assign n14607 = n14599 & n14600 ;
  assign n14610 = n14606 & n14607 ;
  assign n14611 = n14605 & n14610 ;
  assign n14612 = n14609 & n14611 ;
  assign n14613 = n11596 & n14612 ;
  assign n14581 = ~\P2_P1_InstQueue_reg[11][5]/NET0131  & ~n11596 ;
  assign n14614 = n11692 & ~n14581 ;
  assign n14615 = ~n14613 & n14614 ;
  assign n14580 = \P2_P1_InstQueue_reg[11][5]/NET0131  & ~n12345 ;
  assign n14616 = n11378 & ~n11600 ;
  assign n14617 = n12343 & n14616 ;
  assign n14618 = ~n14580 & ~n14617 ;
  assign n14619 = ~n14615 & n14618 ;
  assign n14620 = ~n14579 & n14619 ;
  assign n14622 = ~n11891 & ~n14576 ;
  assign n14621 = n11891 & ~n14573 ;
  assign n14623 = n12407 & ~n14621 ;
  assign n14624 = ~n14622 & n14623 ;
  assign n14627 = n11599 & n14612 ;
  assign n14626 = ~\P2_P1_InstQueue_reg[10][5]/NET0131  & ~n11599 ;
  assign n14628 = n11692 & ~n14626 ;
  assign n14629 = ~n14627 & n14628 ;
  assign n14625 = \P2_P1_InstQueue_reg[10][5]/NET0131  & ~n12414 ;
  assign n14630 = n11378 & ~n11897 ;
  assign n14631 = n12412 & n14630 ;
  assign n14632 = ~n14625 & ~n14631 ;
  assign n14633 = ~n14629 & n14632 ;
  assign n14634 = ~n14624 & n14633 ;
  assign n14636 = ~n11596 & ~n14576 ;
  assign n14635 = n11596 & ~n14573 ;
  assign n14637 = n12464 & ~n14635 ;
  assign n14638 = ~n14636 & n14637 ;
  assign n14641 = n11865 & n14612 ;
  assign n14640 = ~\P2_P1_InstQueue_reg[14][5]/NET0131  & ~n11865 ;
  assign n14642 = n11692 & ~n14640 ;
  assign n14643 = ~n14641 & n14642 ;
  assign n14639 = \P2_P1_InstQueue_reg[14][5]/NET0131  & ~n12471 ;
  assign n14644 = n11378 & ~n11869 ;
  assign n14645 = n12469 & n14644 ;
  assign n14646 = ~n14639 & ~n14645 ;
  assign n14647 = ~n14643 & n14646 ;
  assign n14648 = ~n14638 & n14647 ;
  assign n14650 = ~n11871 & ~n14576 ;
  assign n14649 = n11871 & ~n14573 ;
  assign n14651 = n12540 & ~n14649 ;
  assign n14652 = ~n14650 & n14651 ;
  assign n14655 = n12087 & n14612 ;
  assign n14654 = ~\P2_P1_InstQueue_reg[3][5]/NET0131  & ~n12087 ;
  assign n14656 = n11692 & ~n14654 ;
  assign n14657 = ~n14655 & n14656 ;
  assign n14653 = \P2_P1_InstQueue_reg[3][5]/NET0131  & ~n12547 ;
  assign n14658 = n11378 & ~n12088 ;
  assign n14659 = n12545 & n14658 ;
  assign n14660 = ~n14653 & ~n14659 ;
  assign n14661 = ~n14657 & n14660 ;
  assign n14662 = ~n14652 & n14661 ;
  assign n14664 = ~n12023 & ~n14576 ;
  assign n14663 = n12023 & ~n14573 ;
  assign n14665 = n12559 & ~n14663 ;
  assign n14666 = ~n14664 & n14665 ;
  assign n14669 = n12109 & n14612 ;
  assign n14668 = ~\P2_P1_InstQueue_reg[4][5]/NET0131  & ~n12109 ;
  assign n14670 = n11692 & ~n14668 ;
  assign n14671 = ~n14669 & n14670 ;
  assign n14667 = \P2_P1_InstQueue_reg[4][5]/NET0131  & ~n12566 ;
  assign n14672 = n11378 & ~n12110 ;
  assign n14673 = n12564 & n14672 ;
  assign n14674 = ~n14667 & ~n14673 ;
  assign n14675 = ~n14671 & n14674 ;
  assign n14676 = ~n14666 & n14675 ;
  assign n14678 = ~n12065 & ~n14576 ;
  assign n14677 = n12065 & ~n14573 ;
  assign n14679 = n12578 & ~n14677 ;
  assign n14680 = ~n14678 & n14679 ;
  assign n14683 = n12131 & n14612 ;
  assign n14682 = ~\P2_P1_InstQueue_reg[5][5]/NET0131  & ~n12131 ;
  assign n14684 = n11692 & ~n14682 ;
  assign n14685 = ~n14683 & n14684 ;
  assign n14681 = \P2_P1_InstQueue_reg[5][5]/NET0131  & ~n12585 ;
  assign n14686 = n11378 & ~n12132 ;
  assign n14687 = n12583 & n14686 ;
  assign n14688 = ~n14681 & ~n14687 ;
  assign n14689 = ~n14685 & n14688 ;
  assign n14690 = ~n14680 & n14689 ;
  assign n14692 = ~n12173 & ~n14576 ;
  assign n14691 = n12173 & ~n14573 ;
  assign n14693 = n12654 & ~n14691 ;
  assign n14694 = ~n14692 & n14693 ;
  assign n14697 = n11577 & n14612 ;
  assign n14696 = ~\P2_P1_InstQueue_reg[9][5]/NET0131  & ~n11577 ;
  assign n14698 = n11692 & ~n14696 ;
  assign n14699 = ~n14697 & n14698 ;
  assign n14695 = \P2_P1_InstQueue_reg[9][5]/NET0131  & ~n12661 ;
  assign n14700 = n11378 & ~n11592 ;
  assign n14701 = n12659 & n14700 ;
  assign n14702 = ~n14695 & ~n14701 ;
  assign n14703 = ~n14699 & n14702 ;
  assign n14704 = ~n14694 & n14703 ;
  assign n14711 = ~n8162 & n8177 ;
  assign n14712 = ~n8178 & ~n14711 ;
  assign n14713 = n8139 & ~n14712 ;
  assign n14714 = ~n8025 & n8039 ;
  assign n14715 = ~n8040 & ~n14714 ;
  assign n14716 = ~n8139 & ~n14715 ;
  assign n14717 = ~n14713 & ~n14716 ;
  assign n14718 = n10057 & ~n14717 ;
  assign n14705 = ~n7924 & ~n8146 ;
  assign n14706 = \P1_P1_InstQueue_reg[11][0]/NET0131  & ~n8142 ;
  assign n14707 = ~n8145 & n14706 ;
  assign n14708 = ~n14705 & ~n14707 ;
  assign n14710 = ~n10057 & n14708 ;
  assign n14719 = n8282 & ~n14710 ;
  assign n14720 = ~n14718 & n14719 ;
  assign n14721 = \P1_P1_InstQueue_reg[14][0]/NET0131  & n8291 ;
  assign n14722 = \P1_P1_InstQueue_reg[1][0]/NET0131  & n8299 ;
  assign n14723 = \P1_P1_InstQueue_reg[8][0]/NET0131  & n8305 ;
  assign n14737 = ~n14722 & ~n14723 ;
  assign n14724 = \P1_P1_InstQueue_reg[4][0]/NET0131  & n8295 ;
  assign n14725 = \P1_P1_InstQueue_reg[3][0]/NET0131  & n8323 ;
  assign n14738 = ~n14724 & ~n14725 ;
  assign n14747 = n14737 & n14738 ;
  assign n14748 = ~n14721 & n14747 ;
  assign n14736 = \P1_P1_InstQueue_reg[9][0]/NET0131  & n8325 ;
  assign n14734 = \P1_P1_InstQueue_reg[13][0]/NET0131  & n8327 ;
  assign n14735 = \P1_P1_InstQueue_reg[10][0]/NET0131  & n8303 ;
  assign n14743 = ~n14734 & ~n14735 ;
  assign n14744 = ~n14736 & n14743 ;
  assign n14730 = \P1_P1_InstQueue_reg[6][0]/NET0131  & n8316 ;
  assign n14731 = \P1_P1_InstQueue_reg[15][0]/NET0131  & n8321 ;
  assign n14741 = ~n14730 & ~n14731 ;
  assign n14732 = \P1_P1_InstQueue_reg[7][0]/NET0131  & n8318 ;
  assign n14733 = \P1_P1_InstQueue_reg[2][0]/NET0131  & n8314 ;
  assign n14742 = ~n14732 & ~n14733 ;
  assign n14745 = n14741 & n14742 ;
  assign n14726 = \P1_P1_InstQueue_reg[11][0]/NET0131  & n8312 ;
  assign n14727 = \P1_P1_InstQueue_reg[0][0]/NET0131  & n8309 ;
  assign n14739 = ~n14726 & ~n14727 ;
  assign n14728 = \P1_P1_InstQueue_reg[12][0]/NET0131  & n8329 ;
  assign n14729 = \P1_P1_InstQueue_reg[5][0]/NET0131  & n8307 ;
  assign n14740 = ~n14728 & ~n14729 ;
  assign n14746 = n14739 & n14740 ;
  assign n14749 = n14745 & n14746 ;
  assign n14750 = n14744 & n14749 ;
  assign n14751 = n14748 & n14750 ;
  assign n14752 = n8142 & ~n14751 ;
  assign n14753 = ~n14706 & ~n14752 ;
  assign n14754 = n8350 & ~n14753 ;
  assign n14709 = n8287 & ~n14708 ;
  assign n14755 = \P1_P1_InstQueue_reg[11][0]/NET0131  & ~n8366 ;
  assign n14756 = ~n14709 & ~n14755 ;
  assign n14757 = ~n14754 & n14756 ;
  assign n14758 = ~n14720 & n14757 ;
  assign n14762 = ~n11464 & n11483 ;
  assign n14763 = ~n11484 & ~n14762 ;
  assign n14764 = n10105 & ~n14763 ;
  assign n14759 = ~n11344 & ~n11579 ;
  assign n14760 = ~n11580 & ~n14759 ;
  assign n14761 = ~n10105 & ~n14760 ;
  assign n14765 = n12334 & ~n14761 ;
  assign n14766 = ~n14764 & n14765 ;
  assign n14774 = \P2_P1_InstQueue_reg[6][1]/NET0131  & n11651 ;
  assign n14773 = \P2_P1_InstQueue_reg[15][1]/NET0131  & n11647 ;
  assign n14769 = \P2_P1_InstQueue_reg[10][1]/NET0131  & n11634 ;
  assign n14770 = \P2_P1_InstQueue_reg[3][1]/NET0131  & n11663 ;
  assign n14785 = ~n14769 & ~n14770 ;
  assign n14795 = ~n14773 & n14785 ;
  assign n14796 = ~n14774 & n14795 ;
  assign n14781 = \P2_P1_InstQueue_reg[1][1]/NET0131  & n11671 ;
  assign n14782 = \P2_P1_InstQueue_reg[9][1]/NET0131  & n11656 ;
  assign n14790 = ~n14781 & ~n14782 ;
  assign n14783 = \P2_P1_InstQueue_reg[12][1]/NET0131  & n11673 ;
  assign n14784 = \P2_P1_InstQueue_reg[5][1]/NET0131  & n11638 ;
  assign n14791 = ~n14783 & ~n14784 ;
  assign n14792 = n14790 & n14791 ;
  assign n14777 = \P2_P1_InstQueue_reg[8][1]/NET0131  & n11659 ;
  assign n14778 = \P2_P1_InstQueue_reg[7][1]/NET0131  & n11661 ;
  assign n14788 = ~n14777 & ~n14778 ;
  assign n14779 = \P2_P1_InstQueue_reg[0][1]/NET0131  & n11669 ;
  assign n14780 = \P2_P1_InstQueue_reg[11][1]/NET0131  & n11665 ;
  assign n14789 = ~n14779 & ~n14780 ;
  assign n14793 = n14788 & n14789 ;
  assign n14771 = \P2_P1_InstQueue_reg[13][1]/NET0131  & n11641 ;
  assign n14772 = \P2_P1_InstQueue_reg[14][1]/NET0131  & n11643 ;
  assign n14786 = ~n14771 & ~n14772 ;
  assign n14775 = \P2_P1_InstQueue_reg[4][1]/NET0131  & n11667 ;
  assign n14776 = \P2_P1_InstQueue_reg[2][1]/NET0131  & n11654 ;
  assign n14787 = ~n14775 & ~n14776 ;
  assign n14794 = n14786 & n14787 ;
  assign n14797 = n14793 & n14794 ;
  assign n14798 = n14792 & n14797 ;
  assign n14799 = n14796 & n14798 ;
  assign n14800 = n11596 & n14799 ;
  assign n14768 = ~\P2_P1_InstQueue_reg[11][1]/NET0131  & ~n11596 ;
  assign n14801 = n11692 & ~n14768 ;
  assign n14802 = ~n14800 & n14801 ;
  assign n14767 = \P2_P1_InstQueue_reg[11][1]/NET0131  & ~n12345 ;
  assign n14803 = n11380 & ~n11600 ;
  assign n14804 = n12343 & n14803 ;
  assign n14805 = ~n14767 & ~n14804 ;
  assign n14806 = ~n14802 & n14805 ;
  assign n14807 = ~n14766 & n14806 ;
  assign n14814 = n8375 & ~n14712 ;
  assign n14815 = ~n8375 & ~n14715 ;
  assign n14816 = ~n14814 & ~n14815 ;
  assign n14817 = n11707 & ~n14816 ;
  assign n14808 = ~n7924 & ~n8379 ;
  assign n14809 = \P1_P1_InstQueue_reg[0][0]/NET0131  & ~n8376 ;
  assign n14810 = ~n8378 & n14809 ;
  assign n14811 = ~n14808 & ~n14810 ;
  assign n14813 = ~n11707 & n14811 ;
  assign n14818 = n8282 & ~n14813 ;
  assign n14819 = ~n14817 & n14818 ;
  assign n14820 = n8376 & ~n14751 ;
  assign n14821 = ~n14809 & ~n14820 ;
  assign n14822 = n8350 & ~n14821 ;
  assign n14812 = n8287 & ~n14811 ;
  assign n14823 = \P1_P1_InstQueue_reg[0][0]/NET0131  & ~n8366 ;
  assign n14824 = ~n14812 & ~n14823 ;
  assign n14825 = ~n14822 & n14824 ;
  assign n14826 = ~n14819 & n14825 ;
  assign n14833 = n8407 & ~n14712 ;
  assign n14834 = ~n8407 & ~n14715 ;
  assign n14835 = ~n14833 & ~n14834 ;
  assign n14836 = n9418 & ~n14835 ;
  assign n14827 = ~n7924 & ~n8401 ;
  assign n14828 = \P1_P1_InstQueue_reg[10][0]/NET0131  & ~n8145 ;
  assign n14829 = ~n4327 & n14828 ;
  assign n14830 = ~n14827 & ~n14829 ;
  assign n14832 = ~n9418 & n14830 ;
  assign n14837 = n8282 & ~n14832 ;
  assign n14838 = ~n14836 & n14837 ;
  assign n14839 = n8145 & ~n14751 ;
  assign n14840 = ~n14828 & ~n14839 ;
  assign n14841 = n8350 & ~n14840 ;
  assign n14831 = n8287 & ~n14830 ;
  assign n14842 = \P1_P1_InstQueue_reg[10][0]/NET0131  & ~n8366 ;
  assign n14843 = ~n14831 & ~n14842 ;
  assign n14844 = ~n14841 & n14843 ;
  assign n14845 = ~n14838 & n14844 ;
  assign n14852 = n4327 & ~n14712 ;
  assign n14853 = ~n4327 & ~n14715 ;
  assign n14854 = ~n14852 & ~n14853 ;
  assign n14855 = n11746 & ~n14854 ;
  assign n14846 = ~n7924 & ~n8428 ;
  assign n14847 = \P1_P1_InstQueue_reg[12][0]/NET0131  & ~n8427 ;
  assign n14848 = ~n8142 & n14847 ;
  assign n14849 = ~n14846 & ~n14848 ;
  assign n14851 = ~n11746 & n14849 ;
  assign n14856 = n8282 & ~n14851 ;
  assign n14857 = ~n14855 & n14856 ;
  assign n14858 = n8427 & ~n14751 ;
  assign n14859 = ~n14847 & ~n14858 ;
  assign n14860 = n8350 & ~n14859 ;
  assign n14850 = n8287 & ~n14849 ;
  assign n14861 = \P1_P1_InstQueue_reg[12][0]/NET0131  & ~n8366 ;
  assign n14862 = ~n14850 & ~n14861 ;
  assign n14863 = ~n14860 & n14862 ;
  assign n14864 = ~n14857 & n14863 ;
  assign n14871 = n8145 & ~n14712 ;
  assign n14872 = ~n8145 & ~n14715 ;
  assign n14873 = ~n14871 & ~n14872 ;
  assign n14874 = n11766 & ~n14873 ;
  assign n14865 = ~n7924 & ~n8451 ;
  assign n14866 = \P1_P1_InstQueue_reg[13][0]/NET0131  & ~n8375 ;
  assign n14867 = ~n8427 & n14866 ;
  assign n14868 = ~n14865 & ~n14867 ;
  assign n14870 = ~n11766 & n14868 ;
  assign n14875 = n8282 & ~n14870 ;
  assign n14876 = ~n14874 & n14875 ;
  assign n14877 = n8375 & ~n14751 ;
  assign n14878 = ~n14866 & ~n14877 ;
  assign n14879 = n8350 & ~n14878 ;
  assign n14869 = n8287 & ~n14868 ;
  assign n14880 = \P1_P1_InstQueue_reg[13][0]/NET0131  & ~n8366 ;
  assign n14881 = ~n14869 & ~n14880 ;
  assign n14882 = ~n14879 & n14881 ;
  assign n14883 = ~n14876 & n14882 ;
  assign n14890 = n8142 & ~n14712 ;
  assign n14891 = ~n8142 & ~n14715 ;
  assign n14892 = ~n14890 & ~n14891 ;
  assign n14893 = n11786 & ~n14892 ;
  assign n14884 = ~n7924 & ~n8474 ;
  assign n14885 = \P1_P1_InstQueue_reg[14][0]/NET0131  & ~n8372 ;
  assign n14886 = ~n8375 & n14885 ;
  assign n14887 = ~n14884 & ~n14886 ;
  assign n14889 = ~n11786 & n14887 ;
  assign n14894 = n8282 & ~n14889 ;
  assign n14895 = ~n14893 & n14894 ;
  assign n14896 = n8372 & ~n14751 ;
  assign n14897 = ~n14885 & ~n14896 ;
  assign n14898 = n8350 & ~n14897 ;
  assign n14888 = n8287 & ~n14887 ;
  assign n14899 = \P1_P1_InstQueue_reg[14][0]/NET0131  & ~n8366 ;
  assign n14900 = ~n14888 & ~n14899 ;
  assign n14901 = ~n14898 & n14900 ;
  assign n14902 = ~n14895 & n14901 ;
  assign n14909 = n8427 & ~n14712 ;
  assign n14910 = ~n8427 & ~n14715 ;
  assign n14911 = ~n14909 & ~n14910 ;
  assign n14912 = n11806 & ~n14911 ;
  assign n14903 = ~n7924 & ~n8497 ;
  assign n14904 = \P1_P1_InstQueue_reg[15][0]/NET0131  & ~n8378 ;
  assign n14905 = ~n8372 & n14904 ;
  assign n14906 = ~n14903 & ~n14905 ;
  assign n14908 = ~n11806 & n14906 ;
  assign n14913 = n8282 & ~n14908 ;
  assign n14914 = ~n14912 & n14913 ;
  assign n14915 = n8378 & ~n14751 ;
  assign n14916 = ~n14904 & ~n14915 ;
  assign n14917 = n8350 & ~n14916 ;
  assign n14907 = n8287 & ~n14906 ;
  assign n14918 = \P1_P1_InstQueue_reg[15][0]/NET0131  & ~n8366 ;
  assign n14919 = ~n14907 & ~n14918 ;
  assign n14920 = ~n14917 & n14919 ;
  assign n14921 = ~n14914 & n14920 ;
  assign n14928 = n8372 & ~n14712 ;
  assign n14929 = ~n8372 & ~n14715 ;
  assign n14930 = ~n14928 & ~n14929 ;
  assign n14931 = n11826 & ~n14930 ;
  assign n14922 = ~n7924 & ~n8521 ;
  assign n14923 = \P1_P1_InstQueue_reg[1][0]/NET0131  & ~n8520 ;
  assign n14924 = ~n8376 & n14923 ;
  assign n14925 = ~n14922 & ~n14924 ;
  assign n14927 = ~n11826 & n14925 ;
  assign n14932 = n8282 & ~n14927 ;
  assign n14933 = ~n14931 & n14932 ;
  assign n14934 = n8520 & ~n14751 ;
  assign n14935 = ~n14923 & ~n14934 ;
  assign n14936 = n8350 & ~n14935 ;
  assign n14926 = n8287 & ~n14925 ;
  assign n14937 = \P1_P1_InstQueue_reg[1][0]/NET0131  & ~n8366 ;
  assign n14938 = ~n14926 & ~n14937 ;
  assign n14939 = ~n14936 & n14938 ;
  assign n14940 = ~n14933 & n14939 ;
  assign n14947 = n8378 & ~n14712 ;
  assign n14948 = ~n8378 & ~n14715 ;
  assign n14949 = ~n14947 & ~n14948 ;
  assign n14950 = n11846 & ~n14949 ;
  assign n14941 = ~n7924 & ~n8545 ;
  assign n14942 = \P1_P1_InstQueue_reg[2][0]/NET0131  & ~n8544 ;
  assign n14943 = ~n8520 & n14942 ;
  assign n14944 = ~n14941 & ~n14943 ;
  assign n14946 = ~n11846 & n14944 ;
  assign n14951 = n8282 & ~n14946 ;
  assign n14952 = ~n14950 & n14951 ;
  assign n14953 = n8544 & ~n14751 ;
  assign n14954 = ~n14942 & ~n14953 ;
  assign n14955 = n8350 & ~n14954 ;
  assign n14945 = n8287 & ~n14944 ;
  assign n14956 = \P1_P1_InstQueue_reg[2][0]/NET0131  & ~n8366 ;
  assign n14957 = ~n14945 & ~n14956 ;
  assign n14958 = ~n14955 & n14957 ;
  assign n14959 = ~n14952 & n14958 ;
  assign n14961 = n11862 & ~n14763 ;
  assign n14960 = ~n11862 & ~n14760 ;
  assign n14962 = n12388 & ~n14960 ;
  assign n14963 = ~n14961 & n14962 ;
  assign n14966 = n11871 & n14799 ;
  assign n14965 = ~\P2_P1_InstQueue_reg[0][1]/NET0131  & ~n11871 ;
  assign n14967 = n11692 & ~n14965 ;
  assign n14968 = ~n14966 & n14967 ;
  assign n14964 = \P2_P1_InstQueue_reg[0][1]/NET0131  & ~n12395 ;
  assign n14969 = n11380 & ~n11874 ;
  assign n14970 = n12393 & n14969 ;
  assign n14971 = ~n14964 & ~n14970 ;
  assign n14972 = ~n14968 & n14971 ;
  assign n14973 = ~n14963 & n14972 ;
  assign n14975 = n11891 & ~n14763 ;
  assign n14974 = ~n11891 & ~n14760 ;
  assign n14976 = n12407 & ~n14974 ;
  assign n14977 = ~n14975 & n14976 ;
  assign n14980 = n11599 & n14799 ;
  assign n14979 = ~\P2_P1_InstQueue_reg[10][1]/NET0131  & ~n11599 ;
  assign n14981 = n11692 & ~n14979 ;
  assign n14982 = ~n14980 & n14981 ;
  assign n14978 = \P2_P1_InstQueue_reg[10][1]/NET0131  & ~n12414 ;
  assign n14983 = n11380 & ~n11897 ;
  assign n14984 = n12412 & n14983 ;
  assign n14985 = ~n14978 & ~n14984 ;
  assign n14986 = ~n14982 & n14985 ;
  assign n14987 = ~n14977 & n14986 ;
  assign n14994 = n8376 & ~n14712 ;
  assign n14995 = ~n8376 & ~n14715 ;
  assign n14996 = ~n14994 & ~n14995 ;
  assign n14997 = n11941 & ~n14996 ;
  assign n14988 = ~n7924 & ~n8569 ;
  assign n14989 = \P1_P1_InstQueue_reg[3][0]/NET0131  & ~n8568 ;
  assign n14990 = ~n8544 & n14989 ;
  assign n14991 = ~n14988 & ~n14990 ;
  assign n14993 = ~n11941 & n14991 ;
  assign n14998 = n8282 & ~n14993 ;
  assign n14999 = ~n14997 & n14998 ;
  assign n15000 = n8568 & ~n14751 ;
  assign n15001 = ~n14989 & ~n15000 ;
  assign n15002 = n8350 & ~n15001 ;
  assign n14992 = n8287 & ~n14991 ;
  assign n15003 = \P1_P1_InstQueue_reg[3][0]/NET0131  & ~n8366 ;
  assign n15004 = ~n14992 & ~n15003 ;
  assign n15005 = ~n15002 & n15004 ;
  assign n15006 = ~n14999 & n15005 ;
  assign n15008 = n11577 & ~n14763 ;
  assign n15007 = ~n11577 & ~n14760 ;
  assign n15009 = n12426 & ~n15007 ;
  assign n15010 = ~n15008 & n15009 ;
  assign n15013 = n11919 & n14799 ;
  assign n15012 = ~\P2_P1_InstQueue_reg[12][1]/NET0131  & ~n11919 ;
  assign n15014 = n11692 & ~n15012 ;
  assign n15015 = ~n15013 & n15014 ;
  assign n15011 = \P2_P1_InstQueue_reg[12][1]/NET0131  & ~n12433 ;
  assign n15016 = n11380 & ~n11920 ;
  assign n15017 = n12431 & n15016 ;
  assign n15018 = ~n15011 & ~n15017 ;
  assign n15019 = ~n15015 & n15018 ;
  assign n15020 = ~n15010 & n15019 ;
  assign n15022 = n11599 & ~n14763 ;
  assign n15021 = ~n11599 & ~n14760 ;
  assign n15023 = n12445 & ~n15021 ;
  assign n15024 = ~n15022 & n15023 ;
  assign n15027 = n11862 & n14799 ;
  assign n15026 = ~\P2_P1_InstQueue_reg[13][1]/NET0131  & ~n11862 ;
  assign n15028 = n11692 & ~n15026 ;
  assign n15029 = ~n15027 & n15028 ;
  assign n15025 = \P2_P1_InstQueue_reg[13][1]/NET0131  & ~n12452 ;
  assign n15030 = n11380 & ~n11961 ;
  assign n15031 = n12450 & n15030 ;
  assign n15032 = ~n15025 & ~n15031 ;
  assign n15033 = ~n15029 & n15032 ;
  assign n15034 = ~n15024 & n15033 ;
  assign n15036 = n11596 & ~n14763 ;
  assign n15035 = ~n11596 & ~n14760 ;
  assign n15037 = n12464 & ~n15035 ;
  assign n15038 = ~n15036 & n15037 ;
  assign n15041 = n11865 & n14799 ;
  assign n15040 = ~\P2_P1_InstQueue_reg[14][1]/NET0131  & ~n11865 ;
  assign n15042 = n11692 & ~n15040 ;
  assign n15043 = ~n15041 & n15042 ;
  assign n15039 = \P2_P1_InstQueue_reg[14][1]/NET0131  & ~n12471 ;
  assign n15044 = n11380 & ~n11869 ;
  assign n15045 = n12469 & n15044 ;
  assign n15046 = ~n15039 & ~n15045 ;
  assign n15047 = ~n15043 & n15046 ;
  assign n15048 = ~n15038 & n15047 ;
  assign n15050 = n11919 & ~n14763 ;
  assign n15049 = ~n11919 & ~n14760 ;
  assign n15051 = n12483 & ~n15049 ;
  assign n15052 = ~n15050 & n15051 ;
  assign n15055 = n11873 & n14799 ;
  assign n15054 = ~\P2_P1_InstQueue_reg[15][1]/NET0131  & ~n11873 ;
  assign n15056 = n11692 & ~n15054 ;
  assign n15057 = ~n15055 & n15056 ;
  assign n15053 = \P2_P1_InstQueue_reg[15][1]/NET0131  & ~n12490 ;
  assign n15058 = n11380 & ~n12002 ;
  assign n15059 = n12488 & n15058 ;
  assign n15060 = ~n15053 & ~n15059 ;
  assign n15061 = ~n15057 & n15060 ;
  assign n15062 = ~n15052 & n15061 ;
  assign n15069 = n8520 & ~n14712 ;
  assign n15070 = ~n8520 & ~n14715 ;
  assign n15071 = ~n15069 & ~n15070 ;
  assign n15072 = n12045 & ~n15071 ;
  assign n15063 = ~n7924 & ~n8593 ;
  assign n15064 = \P1_P1_InstQueue_reg[4][0]/NET0131  & ~n8592 ;
  assign n15065 = ~n8568 & n15064 ;
  assign n15066 = ~n15063 & ~n15065 ;
  assign n15068 = ~n12045 & n15066 ;
  assign n15073 = n8282 & ~n15068 ;
  assign n15074 = ~n15072 & n15073 ;
  assign n15075 = n8592 & ~n14751 ;
  assign n15076 = ~n15064 & ~n15075 ;
  assign n15077 = n8350 & ~n15076 ;
  assign n15067 = n8287 & ~n15066 ;
  assign n15078 = \P1_P1_InstQueue_reg[4][0]/NET0131  & ~n8366 ;
  assign n15079 = ~n15067 & ~n15078 ;
  assign n15080 = ~n15077 & n15079 ;
  assign n15081 = ~n15074 & n15080 ;
  assign n15083 = n11865 & ~n14763 ;
  assign n15082 = ~n11865 & ~n14760 ;
  assign n15084 = n12502 & ~n15082 ;
  assign n15085 = ~n15083 & n15084 ;
  assign n15088 = n12023 & n14799 ;
  assign n15087 = ~\P2_P1_InstQueue_reg[1][1]/NET0131  & ~n12023 ;
  assign n15089 = n11692 & ~n15087 ;
  assign n15090 = ~n15088 & n15089 ;
  assign n15086 = \P2_P1_InstQueue_reg[1][1]/NET0131  & ~n12509 ;
  assign n15091 = n11380 & ~n12024 ;
  assign n15092 = n12507 & n15091 ;
  assign n15093 = ~n15086 & ~n15092 ;
  assign n15094 = ~n15090 & n15093 ;
  assign n15095 = ~n15085 & n15094 ;
  assign n15097 = n11873 & ~n14763 ;
  assign n15096 = ~n11873 & ~n14760 ;
  assign n15098 = n12521 & ~n15096 ;
  assign n15099 = ~n15097 & n15098 ;
  assign n15102 = n12065 & n14799 ;
  assign n15101 = ~\P2_P1_InstQueue_reg[2][1]/NET0131  & ~n12065 ;
  assign n15103 = n11692 & ~n15101 ;
  assign n15104 = ~n15102 & n15103 ;
  assign n15100 = \P2_P1_InstQueue_reg[2][1]/NET0131  & ~n12528 ;
  assign n15105 = n11380 & ~n12066 ;
  assign n15106 = n12526 & n15105 ;
  assign n15107 = ~n15100 & ~n15106 ;
  assign n15108 = ~n15104 & n15107 ;
  assign n15109 = ~n15099 & n15108 ;
  assign n15111 = n11871 & ~n14763 ;
  assign n15110 = ~n11871 & ~n14760 ;
  assign n15112 = n12540 & ~n15110 ;
  assign n15113 = ~n15111 & n15112 ;
  assign n15116 = n12087 & n14799 ;
  assign n15115 = ~\P2_P1_InstQueue_reg[3][1]/NET0131  & ~n12087 ;
  assign n15117 = n11692 & ~n15115 ;
  assign n15118 = ~n15116 & n15117 ;
  assign n15114 = \P2_P1_InstQueue_reg[3][1]/NET0131  & ~n12547 ;
  assign n15119 = n11380 & ~n12088 ;
  assign n15120 = n12545 & n15119 ;
  assign n15121 = ~n15114 & ~n15120 ;
  assign n15122 = ~n15118 & n15121 ;
  assign n15123 = ~n15113 & n15122 ;
  assign n15125 = n12023 & ~n14763 ;
  assign n15124 = ~n12023 & ~n14760 ;
  assign n15126 = n12559 & ~n15124 ;
  assign n15127 = ~n15125 & n15126 ;
  assign n15130 = n12109 & n14799 ;
  assign n15129 = ~\P2_P1_InstQueue_reg[4][1]/NET0131  & ~n12109 ;
  assign n15131 = n11692 & ~n15129 ;
  assign n15132 = ~n15130 & n15131 ;
  assign n15128 = \P2_P1_InstQueue_reg[4][1]/NET0131  & ~n12566 ;
  assign n15133 = n11380 & ~n12110 ;
  assign n15134 = n12564 & n15133 ;
  assign n15135 = ~n15128 & ~n15134 ;
  assign n15136 = ~n15132 & n15135 ;
  assign n15137 = ~n15127 & n15136 ;
  assign n15144 = n8544 & ~n14712 ;
  assign n15145 = ~n8544 & ~n14715 ;
  assign n15146 = ~n15144 & ~n15145 ;
  assign n15147 = n12153 & ~n15146 ;
  assign n15138 = ~n7924 & ~n8617 ;
  assign n15139 = \P1_P1_InstQueue_reg[5][0]/NET0131  & ~n8616 ;
  assign n15140 = ~n8592 & n15139 ;
  assign n15141 = ~n15138 & ~n15140 ;
  assign n15143 = ~n12153 & n15141 ;
  assign n15148 = n8282 & ~n15143 ;
  assign n15149 = ~n15147 & n15148 ;
  assign n15150 = n8616 & ~n14751 ;
  assign n15151 = ~n15139 & ~n15150 ;
  assign n15152 = n8350 & ~n15151 ;
  assign n15142 = n8287 & ~n15141 ;
  assign n15153 = \P1_P1_InstQueue_reg[5][0]/NET0131  & ~n8366 ;
  assign n15154 = ~n15142 & ~n15153 ;
  assign n15155 = ~n15152 & n15154 ;
  assign n15156 = ~n15149 & n15155 ;
  assign n15158 = n12065 & ~n14763 ;
  assign n15157 = ~n12065 & ~n14760 ;
  assign n15159 = n12578 & ~n15157 ;
  assign n15160 = ~n15158 & n15159 ;
  assign n15163 = n12131 & n14799 ;
  assign n15162 = ~\P2_P1_InstQueue_reg[5][1]/NET0131  & ~n12131 ;
  assign n15164 = n11692 & ~n15162 ;
  assign n15165 = ~n15163 & n15164 ;
  assign n15161 = \P2_P1_InstQueue_reg[5][1]/NET0131  & ~n12585 ;
  assign n15166 = n11380 & ~n12132 ;
  assign n15167 = n12583 & n15166 ;
  assign n15168 = ~n15161 & ~n15167 ;
  assign n15169 = ~n15165 & n15168 ;
  assign n15170 = ~n15160 & n15169 ;
  assign n15172 = n12087 & ~n14763 ;
  assign n15171 = ~n12087 & ~n14760 ;
  assign n15173 = n12597 & ~n15171 ;
  assign n15174 = ~n15172 & n15173 ;
  assign n15177 = n12173 & n14799 ;
  assign n15176 = ~\P2_P1_InstQueue_reg[6][1]/NET0131  & ~n12173 ;
  assign n15178 = n11692 & ~n15176 ;
  assign n15179 = ~n15177 & n15178 ;
  assign n15175 = \P2_P1_InstQueue_reg[6][1]/NET0131  & ~n12604 ;
  assign n15180 = n11380 & ~n12174 ;
  assign n15181 = n12602 & n15180 ;
  assign n15182 = ~n15175 & ~n15181 ;
  assign n15183 = ~n15179 & n15182 ;
  assign n15184 = ~n15174 & n15183 ;
  assign n15186 = n12109 & ~n14763 ;
  assign n15185 = ~n12109 & ~n14760 ;
  assign n15187 = n12616 & ~n15185 ;
  assign n15188 = ~n15186 & n15187 ;
  assign n15191 = n11891 & n14799 ;
  assign n15190 = ~\P2_P1_InstQueue_reg[7][1]/NET0131  & ~n11891 ;
  assign n15192 = n11692 & ~n15190 ;
  assign n15193 = ~n15191 & n15192 ;
  assign n15189 = \P2_P1_InstQueue_reg[7][1]/NET0131  & ~n12623 ;
  assign n15194 = n11380 & ~n12195 ;
  assign n15195 = n12621 & n15194 ;
  assign n15196 = ~n15189 & ~n15195 ;
  assign n15197 = ~n15193 & n15196 ;
  assign n15198 = ~n15188 & n15197 ;
  assign n15200 = n12131 & ~n14763 ;
  assign n15199 = ~n12131 & ~n14760 ;
  assign n15201 = n12635 & ~n15199 ;
  assign n15202 = ~n15200 & n15201 ;
  assign n15205 = n10105 & n14799 ;
  assign n15204 = ~\P2_P1_InstQueue_reg[8][1]/NET0131  & ~n10105 ;
  assign n15206 = n11692 & ~n15204 ;
  assign n15207 = ~n15205 & n15206 ;
  assign n15203 = \P2_P1_InstQueue_reg[8][1]/NET0131  & ~n12642 ;
  assign n15208 = n11380 & ~n11895 ;
  assign n15209 = n12640 & n15208 ;
  assign n15210 = ~n15203 & ~n15209 ;
  assign n15211 = ~n15207 & n15210 ;
  assign n15212 = ~n15202 & n15211 ;
  assign n15219 = n8568 & ~n14712 ;
  assign n15220 = ~n8568 & ~n14715 ;
  assign n15221 = ~n15219 & ~n15220 ;
  assign n15222 = n12256 & ~n15221 ;
  assign n15213 = ~n7924 & ~n8641 ;
  assign n15214 = \P1_P1_InstQueue_reg[6][0]/NET0131  & ~n8640 ;
  assign n15215 = ~n8616 & n15214 ;
  assign n15216 = ~n15213 & ~n15215 ;
  assign n15218 = ~n12256 & n15216 ;
  assign n15223 = n8282 & ~n15218 ;
  assign n15224 = ~n15222 & n15223 ;
  assign n15225 = n8640 & ~n14751 ;
  assign n15226 = ~n15214 & ~n15225 ;
  assign n15227 = n8350 & ~n15226 ;
  assign n15217 = n8287 & ~n15216 ;
  assign n15228 = \P1_P1_InstQueue_reg[6][0]/NET0131  & ~n8366 ;
  assign n15229 = ~n15217 & ~n15228 ;
  assign n15230 = ~n15227 & n15229 ;
  assign n15231 = ~n15224 & n15230 ;
  assign n15233 = n12173 & ~n14763 ;
  assign n15232 = ~n12173 & ~n14760 ;
  assign n15234 = n12654 & ~n15232 ;
  assign n15235 = ~n15233 & n15234 ;
  assign n15238 = n11577 & n14799 ;
  assign n15237 = ~\P2_P1_InstQueue_reg[9][1]/NET0131  & ~n11577 ;
  assign n15239 = n11692 & ~n15237 ;
  assign n15240 = ~n15238 & n15239 ;
  assign n15236 = \P2_P1_InstQueue_reg[9][1]/NET0131  & ~n12661 ;
  assign n15241 = n11380 & ~n11592 ;
  assign n15242 = n12659 & n15241 ;
  assign n15243 = ~n15236 & ~n15242 ;
  assign n15244 = ~n15240 & n15243 ;
  assign n15245 = ~n15235 & n15244 ;
  assign n15252 = n8592 & ~n14712 ;
  assign n15253 = ~n8592 & ~n14715 ;
  assign n15254 = ~n15252 & ~n15253 ;
  assign n15255 = n12276 & ~n15254 ;
  assign n15246 = ~n7924 & ~n8664 ;
  assign n15247 = \P1_P1_InstQueue_reg[7][0]/NET0131  & ~n8407 ;
  assign n15248 = ~n8640 & n15247 ;
  assign n15249 = ~n15246 & ~n15248 ;
  assign n15251 = ~n12276 & n15249 ;
  assign n15256 = n8282 & ~n15251 ;
  assign n15257 = ~n15255 & n15256 ;
  assign n15258 = n8407 & ~n14751 ;
  assign n15259 = ~n15247 & ~n15258 ;
  assign n15260 = n8350 & ~n15259 ;
  assign n15250 = n8287 & ~n15249 ;
  assign n15261 = \P1_P1_InstQueue_reg[7][0]/NET0131  & ~n8366 ;
  assign n15262 = ~n15250 & ~n15261 ;
  assign n15263 = ~n15260 & n15262 ;
  assign n15264 = ~n15257 & n15263 ;
  assign n15271 = n8616 & ~n14712 ;
  assign n15272 = ~n8616 & ~n14715 ;
  assign n15273 = ~n15271 & ~n15272 ;
  assign n15274 = n12296 & ~n15273 ;
  assign n15265 = ~n7924 & ~n8410 ;
  assign n15266 = \P1_P1_InstQueue_reg[8][0]/NET0131  & ~n8139 ;
  assign n15267 = ~n8407 & n15266 ;
  assign n15268 = ~n15265 & ~n15267 ;
  assign n15270 = ~n12296 & n15268 ;
  assign n15275 = n8282 & ~n15270 ;
  assign n15276 = ~n15274 & n15275 ;
  assign n15277 = n8139 & ~n14751 ;
  assign n15278 = ~n15266 & ~n15277 ;
  assign n15279 = n8350 & ~n15278 ;
  assign n15269 = n8287 & ~n15268 ;
  assign n15280 = \P1_P1_InstQueue_reg[8][0]/NET0131  & ~n8366 ;
  assign n15281 = ~n15269 & ~n15280 ;
  assign n15282 = ~n15279 & n15281 ;
  assign n15283 = ~n15276 & n15282 ;
  assign n15290 = n8640 & ~n14712 ;
  assign n15291 = ~n8640 & ~n14715 ;
  assign n15292 = ~n15290 & ~n15291 ;
  assign n15293 = n12316 & ~n15292 ;
  assign n15284 = ~n7924 & ~n8709 ;
  assign n15285 = \P1_P1_InstQueue_reg[9][0]/NET0131  & ~n4327 ;
  assign n15286 = ~n8139 & n15285 ;
  assign n15287 = ~n15284 & ~n15286 ;
  assign n15289 = ~n12316 & n15287 ;
  assign n15294 = n8282 & ~n15289 ;
  assign n15295 = ~n15293 & n15294 ;
  assign n15296 = n4327 & ~n14751 ;
  assign n15297 = ~n15285 & ~n15296 ;
  assign n15298 = n8350 & ~n15297 ;
  assign n15288 = n8287 & ~n15287 ;
  assign n15299 = \P1_P1_InstQueue_reg[9][0]/NET0131  & ~n8366 ;
  assign n15300 = ~n15288 & ~n15299 ;
  assign n15301 = ~n15298 & n15300 ;
  assign n15302 = ~n15295 & n15301 ;
  assign n15304 = ~n9218 & n9241 ;
  assign n15305 = ~\P1_P3_Flush_reg/NET0131  & \P1_P3_InstQueueRd_Addr_reg[1]/NET0131  ;
  assign n15306 = \P1_P3_Flush_reg/NET0131  & \P1_P3_InstAddrPointer_reg[0]/NET0131  ;
  assign n15307 = \P1_P3_InstAddrPointer_reg[0]/NET0131  & \P1_P3_InstAddrPointer_reg[1]/NET0131  ;
  assign n15308 = ~\P1_P3_InstAddrPointer_reg[0]/NET0131  & ~\P1_P3_InstAddrPointer_reg[1]/NET0131  ;
  assign n15309 = ~n15307 & ~n15308 ;
  assign n15310 = \P1_P3_InstAddrPointer_reg[31]/NET0131  & ~n15309 ;
  assign n15311 = ~\P1_P3_InstAddrPointer_reg[1]/NET0131  & ~\P1_P3_InstAddrPointer_reg[31]/NET0131  ;
  assign n15312 = ~n15310 & ~n15311 ;
  assign n15313 = n15306 & ~n15312 ;
  assign n15314 = ~n15305 & ~n15313 ;
  assign n15315 = n10037 & ~n15314 ;
  assign n15303 = ~n9207 & n10046 ;
  assign n15316 = ~n8734 & ~n9243 ;
  assign n15317 = ~n10031 & n15316 ;
  assign n15318 = \P1_P3_InstQueueRd_Addr_reg[1]/NET0131  & ~n15317 ;
  assign n15319 = ~n15303 & ~n15318 ;
  assign n15320 = ~n15315 & n15319 ;
  assign n15321 = ~n15304 & n15320 ;
  assign n15322 = \P1_P1_State2_reg[0]/NET0131  & n8353 ;
  assign n15323 = ~n8349 & ~n15322 ;
  assign n15324 = ~\P1_P1_State2_reg[2]/NET0131  & n8354 ;
  assign n15325 = ~n8356 & ~n15324 ;
  assign n15326 = n15323 & n15325 ;
  assign n15327 = \P1_P1_EAX_reg[31]/NET0131  & ~n15326 ;
  assign n15335 = \P1_ready11_reg/NET0131  & \P2_P1_ADS_n_reg/NET0131  ;
  assign n15723 = n7874 & ~n15335 ;
  assign n15336 = \P1_P1_InstQueueRd_Addr_reg[2]/NET0131  & ~\P1_P1_InstQueueWr_Addr_reg[2]/NET0131  ;
  assign n15337 = ~\P1_P1_InstQueueRd_Addr_reg[2]/NET0131  & \P1_P1_InstQueueWr_Addr_reg[2]/NET0131  ;
  assign n15338 = ~n15336 & ~n15337 ;
  assign n15339 = ~\P1_P1_InstQueueRd_Addr_reg[1]/NET0131  & \P1_P1_InstQueueWr_Addr_reg[1]/NET0131  ;
  assign n15340 = \P1_P1_InstQueueRd_Addr_reg[1]/NET0131  & ~\P1_P1_InstQueueWr_Addr_reg[1]/NET0131  ;
  assign n15341 = \P1_P1_InstQueueRd_Addr_reg[0]/NET0131  & ~\P1_P1_InstQueueWr_Addr_reg[0]/NET0131  ;
  assign n15342 = ~n15340 & ~n15341 ;
  assign n15343 = ~n15339 & ~n15342 ;
  assign n15344 = n15338 & n15343 ;
  assign n15345 = ~n15338 & ~n15343 ;
  assign n15346 = ~n15344 & ~n15345 ;
  assign n15347 = \P1_P1_InstQueueRd_Addr_reg[3]/NET0131  & ~\P1_P1_InstQueueWr_Addr_reg[3]/NET0131  ;
  assign n15348 = ~\P1_P1_InstQueueRd_Addr_reg[3]/NET0131  & \P1_P1_InstQueueWr_Addr_reg[3]/NET0131  ;
  assign n15349 = ~n15347 & ~n15348 ;
  assign n15350 = ~n15336 & ~n15343 ;
  assign n15351 = ~n15337 & ~n15350 ;
  assign n15352 = n15349 & n15351 ;
  assign n15353 = ~n15349 & ~n15351 ;
  assign n15354 = ~n15352 & ~n15353 ;
  assign n15355 = n15346 & n15354 ;
  assign n15356 = ~n15347 & ~n15351 ;
  assign n15357 = ~n15348 & ~n15356 ;
  assign n15358 = ~n15355 & ~n15357 ;
  assign n15359 = ~n15339 & ~n15340 ;
  assign n15360 = n15341 & ~n15359 ;
  assign n15361 = ~n15341 & n15359 ;
  assign n15362 = ~n15360 & ~n15361 ;
  assign n15363 = ~n15357 & n15362 ;
  assign n15364 = ~n15358 & ~n15363 ;
  assign n15378 = ~n8345 & ~n9362 ;
  assign n15379 = n9303 & ~n13639 ;
  assign n15380 = n15378 & n15379 ;
  assign n15375 = n10096 & n14751 ;
  assign n15381 = ~n12718 & n15375 ;
  assign n15382 = n15380 & n15381 ;
  assign n15724 = ~n15364 & n15382 ;
  assign n15722 = ~\P1_P1_EAX_reg[31]/NET0131  & n15335 ;
  assign n15725 = n14020 & ~n15722 ;
  assign n15726 = n15724 & n15725 ;
  assign n15727 = ~n15723 & n15726 ;
  assign n15331 = n9303 & n13639 ;
  assign n15373 = n8345 & ~n9362 ;
  assign n15374 = n15331 & n15373 ;
  assign n15368 = n12718 & n14020 ;
  assign n15376 = n15368 & n15375 ;
  assign n15377 = n15374 & n15376 ;
  assign n15388 = \P1_P1_EAX_reg[0]/NET0131  & \P1_P1_EAX_reg[1]/NET0131  ;
  assign n15389 = \P1_P1_EAX_reg[2]/NET0131  & n15388 ;
  assign n15390 = \P1_P1_EAX_reg[3]/NET0131  & n15389 ;
  assign n15391 = \P1_P1_EAX_reg[4]/NET0131  & n15390 ;
  assign n15392 = \P1_P1_EAX_reg[5]/NET0131  & n15391 ;
  assign n15393 = \P1_P1_EAX_reg[6]/NET0131  & n15392 ;
  assign n15394 = \P1_P1_EAX_reg[7]/NET0131  & n15393 ;
  assign n15395 = \P1_P1_EAX_reg[8]/NET0131  & n15394 ;
  assign n15396 = \P1_P1_EAX_reg[9]/NET0131  & n15395 ;
  assign n15397 = \P1_P1_EAX_reg[10]/NET0131  & n15396 ;
  assign n15398 = \P1_P1_EAX_reg[11]/NET0131  & n15397 ;
  assign n15399 = \P1_P1_EAX_reg[12]/NET0131  & n15398 ;
  assign n15400 = \P1_P1_EAX_reg[13]/NET0131  & n15399 ;
  assign n15401 = \P1_P1_EAX_reg[14]/NET0131  & n15400 ;
  assign n15402 = \P1_P1_EAX_reg[15]/NET0131  & n15401 ;
  assign n15403 = \P1_P1_EAX_reg[16]/NET0131  & n15402 ;
  assign n15406 = \P1_P1_EAX_reg[19]/NET0131  & \P1_P1_EAX_reg[20]/NET0131  ;
  assign n15407 = \P1_P1_EAX_reg[23]/NET0131  & \P1_P1_EAX_reg[24]/NET0131  ;
  assign n15408 = n15406 & n15407 ;
  assign n15404 = \P1_P1_EAX_reg[21]/NET0131  & \P1_P1_EAX_reg[22]/NET0131  ;
  assign n15405 = \P1_P1_EAX_reg[17]/NET0131  & \P1_P1_EAX_reg[18]/NET0131  ;
  assign n15409 = n15404 & n15405 ;
  assign n15410 = n15408 & n15409 ;
  assign n15411 = n15403 & n15410 ;
  assign n15412 = \P1_P1_EAX_reg[26]/NET0131  & \P1_P1_EAX_reg[27]/NET0131  ;
  assign n15413 = \P1_P1_EAX_reg[25]/NET0131  & \P1_P1_EAX_reg[28]/NET0131  ;
  assign n15414 = n15412 & n15413 ;
  assign n15415 = n15411 & n15414 ;
  assign n15416 = \P1_P1_EAX_reg[29]/NET0131  & \P1_P1_EAX_reg[30]/NET0131  ;
  assign n15417 = n15415 & n15416 ;
  assign n15418 = n15377 & ~n15417 ;
  assign n15328 = n12718 & ~n14020 ;
  assign n15329 = ~n10096 & ~n14751 ;
  assign n15330 = n15328 & n15329 ;
  assign n15332 = ~n8345 & n9362 ;
  assign n15333 = n15331 & n15332 ;
  assign n15334 = n15330 & n15333 ;
  assign n15365 = ~n15335 & ~n15364 ;
  assign n15366 = n15334 & ~n15365 ;
  assign n15383 = n14020 & n15382 ;
  assign n15384 = ~n15334 & ~n15383 ;
  assign n15369 = ~n9303 & n15332 ;
  assign n15370 = ~n13639 & n15369 ;
  assign n15367 = ~n10096 & n14751 ;
  assign n15371 = n15367 & n15368 ;
  assign n15372 = n15370 & n15371 ;
  assign n15385 = ~n15372 & ~n15377 ;
  assign n15386 = n15384 & n15385 ;
  assign n15387 = ~n15366 & ~n15386 ;
  assign n15419 = n15364 & n15383 ;
  assign n15420 = n15387 & ~n15419 ;
  assign n15421 = ~n15418 & n15420 ;
  assign n15422 = \P1_P1_EAX_reg[31]/NET0131  & ~n15421 ;
  assign n15423 = ~\P1_P1_InstQueueRd_Addr_reg[0]/NET0131  & \P1_P1_InstQueueWr_Addr_reg[0]/NET0131  ;
  assign n15424 = ~n15341 & ~n15423 ;
  assign n15425 = n15359 & n15424 ;
  assign n15426 = ~n15346 & ~n15425 ;
  assign n15427 = n15354 & ~n15426 ;
  assign n15428 = ~n15357 & ~n15427 ;
  assign n15430 = \P1_P1_InstQueue_reg[1][7]/NET0131  & n8291 ;
  assign n15431 = \P1_P1_InstQueue_reg[12][7]/NET0131  & n8325 ;
  assign n15432 = \P1_P1_InstQueue_reg[15][7]/NET0131  & n8329 ;
  assign n15446 = ~n15431 & ~n15432 ;
  assign n15433 = \P1_P1_InstQueue_reg[3][7]/NET0131  & n8309 ;
  assign n15434 = \P1_P1_InstQueue_reg[6][7]/NET0131  & n8323 ;
  assign n15447 = ~n15433 & ~n15434 ;
  assign n15456 = n15446 & n15447 ;
  assign n15457 = ~n15430 & n15456 ;
  assign n15445 = \P1_P1_InstQueue_reg[13][7]/NET0131  & n8303 ;
  assign n15443 = \P1_P1_InstQueue_reg[0][7]/NET0131  & n8327 ;
  assign n15444 = \P1_P1_InstQueue_reg[8][7]/NET0131  & n8307 ;
  assign n15452 = ~n15443 & ~n15444 ;
  assign n15453 = ~n15445 & n15452 ;
  assign n15439 = \P1_P1_InstQueue_reg[9][7]/NET0131  & n8316 ;
  assign n15440 = \P1_P1_InstQueue_reg[2][7]/NET0131  & n8321 ;
  assign n15450 = ~n15439 & ~n15440 ;
  assign n15441 = \P1_P1_InstQueue_reg[10][7]/NET0131  & n8318 ;
  assign n15442 = \P1_P1_InstQueue_reg[4][7]/NET0131  & n8299 ;
  assign n15451 = ~n15441 & ~n15442 ;
  assign n15454 = n15450 & n15451 ;
  assign n15435 = \P1_P1_InstQueue_reg[14][7]/NET0131  & n8312 ;
  assign n15436 = \P1_P1_InstQueue_reg[7][7]/NET0131  & n8295 ;
  assign n15448 = ~n15435 & ~n15436 ;
  assign n15437 = \P1_P1_InstQueue_reg[5][7]/NET0131  & n8314 ;
  assign n15438 = \P1_P1_InstQueue_reg[11][7]/NET0131  & n8305 ;
  assign n15449 = ~n15437 & ~n15438 ;
  assign n15455 = n15448 & n15449 ;
  assign n15458 = n15454 & n15455 ;
  assign n15459 = n15453 & n15458 ;
  assign n15460 = n15457 & n15459 ;
  assign n15461 = \P1_P1_InstQueue_reg[2][0]/NET0131  & n8291 ;
  assign n15462 = \P1_P1_InstQueue_reg[6][0]/NET0131  & n8314 ;
  assign n15463 = \P1_P1_InstQueue_reg[14][0]/NET0131  & n8303 ;
  assign n15477 = ~n15462 & ~n15463 ;
  assign n15464 = \P1_P1_InstQueue_reg[7][0]/NET0131  & n8323 ;
  assign n15465 = \P1_P1_InstQueue_reg[15][0]/NET0131  & n8312 ;
  assign n15478 = ~n15464 & ~n15465 ;
  assign n15487 = n15477 & n15478 ;
  assign n15488 = ~n15461 & n15487 ;
  assign n15476 = \P1_P1_InstQueue_reg[4][0]/NET0131  & n8309 ;
  assign n15474 = \P1_P1_InstQueue_reg[8][0]/NET0131  & n8295 ;
  assign n15475 = \P1_P1_InstQueue_reg[12][0]/NET0131  & n8305 ;
  assign n15483 = ~n15474 & ~n15475 ;
  assign n15484 = ~n15476 & n15483 ;
  assign n15470 = \P1_P1_InstQueue_reg[10][0]/NET0131  & n8316 ;
  assign n15471 = \P1_P1_InstQueue_reg[3][0]/NET0131  & n8321 ;
  assign n15481 = ~n15470 & ~n15471 ;
  assign n15472 = \P1_P1_InstQueue_reg[11][0]/NET0131  & n8318 ;
  assign n15473 = \P1_P1_InstQueue_reg[13][0]/NET0131  & n8325 ;
  assign n15482 = ~n15472 & ~n15473 ;
  assign n15485 = n15481 & n15482 ;
  assign n15466 = \P1_P1_InstQueue_reg[1][0]/NET0131  & n8327 ;
  assign n15467 = \P1_P1_InstQueue_reg[0][0]/NET0131  & n8329 ;
  assign n15479 = ~n15466 & ~n15467 ;
  assign n15468 = \P1_P1_InstQueue_reg[5][0]/NET0131  & n8299 ;
  assign n15469 = \P1_P1_InstQueue_reg[9][0]/NET0131  & n8307 ;
  assign n15480 = ~n15468 & ~n15469 ;
  assign n15486 = n15479 & n15480 ;
  assign n15489 = n15485 & n15486 ;
  assign n15490 = n15484 & n15489 ;
  assign n15491 = n15488 & n15490 ;
  assign n15492 = ~n15460 & ~n15491 ;
  assign n15493 = \P1_P1_InstQueue_reg[2][1]/NET0131  & n8291 ;
  assign n15494 = \P1_P1_InstQueue_reg[7][1]/NET0131  & n8323 ;
  assign n15495 = \P1_P1_InstQueue_reg[13][1]/NET0131  & n8325 ;
  assign n15509 = ~n15494 & ~n15495 ;
  assign n15496 = \P1_P1_InstQueue_reg[8][1]/NET0131  & n8295 ;
  assign n15497 = \P1_P1_InstQueue_reg[15][1]/NET0131  & n8312 ;
  assign n15510 = ~n15496 & ~n15497 ;
  assign n15519 = n15509 & n15510 ;
  assign n15520 = ~n15493 & n15519 ;
  assign n15508 = \P1_P1_InstQueue_reg[4][1]/NET0131  & n8309 ;
  assign n15506 = \P1_P1_InstQueue_reg[0][1]/NET0131  & n8329 ;
  assign n15507 = \P1_P1_InstQueue_reg[12][1]/NET0131  & n8305 ;
  assign n15515 = ~n15506 & ~n15507 ;
  assign n15516 = ~n15508 & n15515 ;
  assign n15502 = \P1_P1_InstQueue_reg[10][1]/NET0131  & n8316 ;
  assign n15503 = \P1_P1_InstQueue_reg[11][1]/NET0131  & n8318 ;
  assign n15513 = ~n15502 & ~n15503 ;
  assign n15504 = \P1_P1_InstQueue_reg[3][1]/NET0131  & n8321 ;
  assign n15505 = \P1_P1_InstQueue_reg[5][1]/NET0131  & n8299 ;
  assign n15514 = ~n15504 & ~n15505 ;
  assign n15517 = n15513 & n15514 ;
  assign n15498 = \P1_P1_InstQueue_reg[1][1]/NET0131  & n8327 ;
  assign n15499 = \P1_P1_InstQueue_reg[9][1]/NET0131  & n8307 ;
  assign n15511 = ~n15498 & ~n15499 ;
  assign n15500 = \P1_P1_InstQueue_reg[6][1]/NET0131  & n8314 ;
  assign n15501 = \P1_P1_InstQueue_reg[14][1]/NET0131  & n8303 ;
  assign n15512 = ~n15500 & ~n15501 ;
  assign n15518 = n15511 & n15512 ;
  assign n15521 = n15517 & n15518 ;
  assign n15522 = n15516 & n15521 ;
  assign n15523 = n15520 & n15522 ;
  assign n15524 = n15492 & ~n15523 ;
  assign n15525 = \P1_P1_InstQueue_reg[2][2]/NET0131  & n8291 ;
  assign n15526 = \P1_P1_InstQueue_reg[6][2]/NET0131  & n8314 ;
  assign n15527 = \P1_P1_InstQueue_reg[14][2]/NET0131  & n8303 ;
  assign n15541 = ~n15526 & ~n15527 ;
  assign n15528 = \P1_P1_InstQueue_reg[7][2]/NET0131  & n8323 ;
  assign n15529 = \P1_P1_InstQueue_reg[15][2]/NET0131  & n8312 ;
  assign n15542 = ~n15528 & ~n15529 ;
  assign n15551 = n15541 & n15542 ;
  assign n15552 = ~n15525 & n15551 ;
  assign n15540 = \P1_P1_InstQueue_reg[4][2]/NET0131  & n8309 ;
  assign n15538 = \P1_P1_InstQueue_reg[8][2]/NET0131  & n8295 ;
  assign n15539 = \P1_P1_InstQueue_reg[12][2]/NET0131  & n8305 ;
  assign n15547 = ~n15538 & ~n15539 ;
  assign n15548 = ~n15540 & n15547 ;
  assign n15534 = \P1_P1_InstQueue_reg[10][2]/NET0131  & n8316 ;
  assign n15535 = \P1_P1_InstQueue_reg[3][2]/NET0131  & n8321 ;
  assign n15545 = ~n15534 & ~n15535 ;
  assign n15536 = \P1_P1_InstQueue_reg[11][2]/NET0131  & n8318 ;
  assign n15537 = \P1_P1_InstQueue_reg[13][2]/NET0131  & n8325 ;
  assign n15546 = ~n15536 & ~n15537 ;
  assign n15549 = n15545 & n15546 ;
  assign n15530 = \P1_P1_InstQueue_reg[1][2]/NET0131  & n8327 ;
  assign n15531 = \P1_P1_InstQueue_reg[0][2]/NET0131  & n8329 ;
  assign n15543 = ~n15530 & ~n15531 ;
  assign n15532 = \P1_P1_InstQueue_reg[5][2]/NET0131  & n8299 ;
  assign n15533 = \P1_P1_InstQueue_reg[9][2]/NET0131  & n8307 ;
  assign n15544 = ~n15532 & ~n15533 ;
  assign n15550 = n15543 & n15544 ;
  assign n15553 = n15549 & n15550 ;
  assign n15554 = n15548 & n15553 ;
  assign n15555 = n15552 & n15554 ;
  assign n15556 = n15524 & ~n15555 ;
  assign n15557 = \P1_P1_InstQueue_reg[2][3]/NET0131  & n8291 ;
  assign n15558 = \P1_P1_InstQueue_reg[6][3]/NET0131  & n8314 ;
  assign n15559 = \P1_P1_InstQueue_reg[14][3]/NET0131  & n8303 ;
  assign n15573 = ~n15558 & ~n15559 ;
  assign n15560 = \P1_P1_InstQueue_reg[7][3]/NET0131  & n8323 ;
  assign n15561 = \P1_P1_InstQueue_reg[15][3]/NET0131  & n8312 ;
  assign n15574 = ~n15560 & ~n15561 ;
  assign n15583 = n15573 & n15574 ;
  assign n15584 = ~n15557 & n15583 ;
  assign n15572 = \P1_P1_InstQueue_reg[4][3]/NET0131  & n8309 ;
  assign n15570 = \P1_P1_InstQueue_reg[8][3]/NET0131  & n8295 ;
  assign n15571 = \P1_P1_InstQueue_reg[12][3]/NET0131  & n8305 ;
  assign n15579 = ~n15570 & ~n15571 ;
  assign n15580 = ~n15572 & n15579 ;
  assign n15566 = \P1_P1_InstQueue_reg[10][3]/NET0131  & n8316 ;
  assign n15567 = \P1_P1_InstQueue_reg[3][3]/NET0131  & n8321 ;
  assign n15577 = ~n15566 & ~n15567 ;
  assign n15568 = \P1_P1_InstQueue_reg[11][3]/NET0131  & n8318 ;
  assign n15569 = \P1_P1_InstQueue_reg[9][3]/NET0131  & n8307 ;
  assign n15578 = ~n15568 & ~n15569 ;
  assign n15581 = n15577 & n15578 ;
  assign n15562 = \P1_P1_InstQueue_reg[1][3]/NET0131  & n8327 ;
  assign n15563 = \P1_P1_InstQueue_reg[0][3]/NET0131  & n8329 ;
  assign n15575 = ~n15562 & ~n15563 ;
  assign n15564 = \P1_P1_InstQueue_reg[5][3]/NET0131  & n8299 ;
  assign n15565 = \P1_P1_InstQueue_reg[13][3]/NET0131  & n8325 ;
  assign n15576 = ~n15564 & ~n15565 ;
  assign n15582 = n15575 & n15576 ;
  assign n15585 = n15581 & n15582 ;
  assign n15586 = n15580 & n15585 ;
  assign n15587 = n15584 & n15586 ;
  assign n15588 = n15556 & ~n15587 ;
  assign n15589 = \P1_P1_InstQueue_reg[2][4]/NET0131  & n8291 ;
  assign n15590 = \P1_P1_InstQueue_reg[7][4]/NET0131  & n8323 ;
  assign n15591 = \P1_P1_InstQueue_reg[13][4]/NET0131  & n8325 ;
  assign n15605 = ~n15590 & ~n15591 ;
  assign n15592 = \P1_P1_InstQueue_reg[8][4]/NET0131  & n8295 ;
  assign n15593 = \P1_P1_InstQueue_reg[15][4]/NET0131  & n8312 ;
  assign n15606 = ~n15592 & ~n15593 ;
  assign n15615 = n15605 & n15606 ;
  assign n15616 = ~n15589 & n15615 ;
  assign n15604 = \P1_P1_InstQueue_reg[4][4]/NET0131  & n8309 ;
  assign n15602 = \P1_P1_InstQueue_reg[0][4]/NET0131  & n8329 ;
  assign n15603 = \P1_P1_InstQueue_reg[12][4]/NET0131  & n8305 ;
  assign n15611 = ~n15602 & ~n15603 ;
  assign n15612 = ~n15604 & n15611 ;
  assign n15598 = \P1_P1_InstQueue_reg[10][4]/NET0131  & n8316 ;
  assign n15599 = \P1_P1_InstQueue_reg[11][4]/NET0131  & n8318 ;
  assign n15609 = ~n15598 & ~n15599 ;
  assign n15600 = \P1_P1_InstQueue_reg[3][4]/NET0131  & n8321 ;
  assign n15601 = \P1_P1_InstQueue_reg[5][4]/NET0131  & n8299 ;
  assign n15610 = ~n15600 & ~n15601 ;
  assign n15613 = n15609 & n15610 ;
  assign n15594 = \P1_P1_InstQueue_reg[1][4]/NET0131  & n8327 ;
  assign n15595 = \P1_P1_InstQueue_reg[9][4]/NET0131  & n8307 ;
  assign n15607 = ~n15594 & ~n15595 ;
  assign n15596 = \P1_P1_InstQueue_reg[6][4]/NET0131  & n8314 ;
  assign n15597 = \P1_P1_InstQueue_reg[14][4]/NET0131  & n8303 ;
  assign n15608 = ~n15596 & ~n15597 ;
  assign n15614 = n15607 & n15608 ;
  assign n15617 = n15613 & n15614 ;
  assign n15618 = n15612 & n15617 ;
  assign n15619 = n15616 & n15618 ;
  assign n15620 = n15588 & ~n15619 ;
  assign n15621 = \P1_P1_InstQueue_reg[2][5]/NET0131  & n8291 ;
  assign n15622 = \P1_P1_InstQueue_reg[6][5]/NET0131  & n8314 ;
  assign n15623 = \P1_P1_InstQueue_reg[14][5]/NET0131  & n8303 ;
  assign n15637 = ~n15622 & ~n15623 ;
  assign n15624 = \P1_P1_InstQueue_reg[7][5]/NET0131  & n8323 ;
  assign n15625 = \P1_P1_InstQueue_reg[15][5]/NET0131  & n8312 ;
  assign n15638 = ~n15624 & ~n15625 ;
  assign n15647 = n15637 & n15638 ;
  assign n15648 = ~n15621 & n15647 ;
  assign n15636 = \P1_P1_InstQueue_reg[4][5]/NET0131  & n8309 ;
  assign n15634 = \P1_P1_InstQueue_reg[8][5]/NET0131  & n8295 ;
  assign n15635 = \P1_P1_InstQueue_reg[12][5]/NET0131  & n8305 ;
  assign n15643 = ~n15634 & ~n15635 ;
  assign n15644 = ~n15636 & n15643 ;
  assign n15630 = \P1_P1_InstQueue_reg[10][5]/NET0131  & n8316 ;
  assign n15631 = \P1_P1_InstQueue_reg[3][5]/NET0131  & n8321 ;
  assign n15641 = ~n15630 & ~n15631 ;
  assign n15632 = \P1_P1_InstQueue_reg[11][5]/NET0131  & n8318 ;
  assign n15633 = \P1_P1_InstQueue_reg[9][5]/NET0131  & n8307 ;
  assign n15642 = ~n15632 & ~n15633 ;
  assign n15645 = n15641 & n15642 ;
  assign n15626 = \P1_P1_InstQueue_reg[1][5]/NET0131  & n8327 ;
  assign n15627 = \P1_P1_InstQueue_reg[0][5]/NET0131  & n8329 ;
  assign n15639 = ~n15626 & ~n15627 ;
  assign n15628 = \P1_P1_InstQueue_reg[5][5]/NET0131  & n8299 ;
  assign n15629 = \P1_P1_InstQueue_reg[13][5]/NET0131  & n8325 ;
  assign n15640 = ~n15628 & ~n15629 ;
  assign n15646 = n15639 & n15640 ;
  assign n15649 = n15645 & n15646 ;
  assign n15650 = n15644 & n15649 ;
  assign n15651 = n15648 & n15650 ;
  assign n15652 = n15620 & ~n15651 ;
  assign n15653 = \P1_P1_InstQueue_reg[2][6]/NET0131  & n8291 ;
  assign n15654 = \P1_P1_InstQueue_reg[6][6]/NET0131  & n8314 ;
  assign n15655 = \P1_P1_InstQueue_reg[14][6]/NET0131  & n8303 ;
  assign n15669 = ~n15654 & ~n15655 ;
  assign n15656 = \P1_P1_InstQueue_reg[7][6]/NET0131  & n8323 ;
  assign n15657 = \P1_P1_InstQueue_reg[15][6]/NET0131  & n8312 ;
  assign n15670 = ~n15656 & ~n15657 ;
  assign n15679 = n15669 & n15670 ;
  assign n15680 = ~n15653 & n15679 ;
  assign n15668 = \P1_P1_InstQueue_reg[4][6]/NET0131  & n8309 ;
  assign n15666 = \P1_P1_InstQueue_reg[8][6]/NET0131  & n8295 ;
  assign n15667 = \P1_P1_InstQueue_reg[12][6]/NET0131  & n8305 ;
  assign n15675 = ~n15666 & ~n15667 ;
  assign n15676 = ~n15668 & n15675 ;
  assign n15662 = \P1_P1_InstQueue_reg[10][6]/NET0131  & n8316 ;
  assign n15663 = \P1_P1_InstQueue_reg[3][6]/NET0131  & n8321 ;
  assign n15673 = ~n15662 & ~n15663 ;
  assign n15664 = \P1_P1_InstQueue_reg[11][6]/NET0131  & n8318 ;
  assign n15665 = \P1_P1_InstQueue_reg[13][6]/NET0131  & n8325 ;
  assign n15674 = ~n15664 & ~n15665 ;
  assign n15677 = n15673 & n15674 ;
  assign n15658 = \P1_P1_InstQueue_reg[1][6]/NET0131  & n8327 ;
  assign n15659 = \P1_P1_InstQueue_reg[0][6]/NET0131  & n8329 ;
  assign n15671 = ~n15658 & ~n15659 ;
  assign n15660 = \P1_P1_InstQueue_reg[5][6]/NET0131  & n8299 ;
  assign n15661 = \P1_P1_InstQueue_reg[9][6]/NET0131  & n8307 ;
  assign n15672 = ~n15660 & ~n15661 ;
  assign n15678 = n15671 & n15672 ;
  assign n15681 = n15677 & n15678 ;
  assign n15682 = n15676 & n15681 ;
  assign n15683 = n15680 & n15682 ;
  assign n15684 = n15652 & ~n15683 ;
  assign n15685 = \P1_P1_InstQueue_reg[2][7]/NET0131  & n8291 ;
  assign n15686 = \P1_P1_InstQueue_reg[6][7]/NET0131  & n8314 ;
  assign n15687 = \P1_P1_InstQueue_reg[14][7]/NET0131  & n8303 ;
  assign n15701 = ~n15686 & ~n15687 ;
  assign n15688 = \P1_P1_InstQueue_reg[7][7]/NET0131  & n8323 ;
  assign n15689 = \P1_P1_InstQueue_reg[15][7]/NET0131  & n8312 ;
  assign n15702 = ~n15688 & ~n15689 ;
  assign n15711 = n15701 & n15702 ;
  assign n15712 = ~n15685 & n15711 ;
  assign n15700 = \P1_P1_InstQueue_reg[4][7]/NET0131  & n8309 ;
  assign n15698 = \P1_P1_InstQueue_reg[8][7]/NET0131  & n8295 ;
  assign n15699 = \P1_P1_InstQueue_reg[12][7]/NET0131  & n8305 ;
  assign n15707 = ~n15698 & ~n15699 ;
  assign n15708 = ~n15700 & n15707 ;
  assign n15694 = \P1_P1_InstQueue_reg[10][7]/NET0131  & n8316 ;
  assign n15695 = \P1_P1_InstQueue_reg[3][7]/NET0131  & n8321 ;
  assign n15705 = ~n15694 & ~n15695 ;
  assign n15696 = \P1_P1_InstQueue_reg[11][7]/NET0131  & n8318 ;
  assign n15697 = \P1_P1_InstQueue_reg[13][7]/NET0131  & n8325 ;
  assign n15706 = ~n15696 & ~n15697 ;
  assign n15709 = n15705 & n15706 ;
  assign n15690 = \P1_P1_InstQueue_reg[1][7]/NET0131  & n8327 ;
  assign n15691 = \P1_P1_InstQueue_reg[0][7]/NET0131  & n8329 ;
  assign n15703 = ~n15690 & ~n15691 ;
  assign n15692 = \P1_P1_InstQueue_reg[5][7]/NET0131  & n8299 ;
  assign n15693 = \P1_P1_InstQueue_reg[9][7]/NET0131  & n8307 ;
  assign n15704 = ~n15692 & ~n15693 ;
  assign n15710 = n15703 & n15704 ;
  assign n15713 = n15709 & n15710 ;
  assign n15714 = n15708 & n15713 ;
  assign n15715 = n15712 & n15714 ;
  assign n15716 = n15684 & ~n15715 ;
  assign n15717 = n15428 & ~n15716 ;
  assign n15429 = ~\P1_P1_EAX_reg[31]/NET0131  & ~n15428 ;
  assign n15718 = n15372 & ~n15429 ;
  assign n15719 = ~n15717 & n15718 ;
  assign n15720 = ~\P1_P1_EAX_reg[31]/NET0131  & n15377 ;
  assign n15721 = n15417 & n15720 ;
  assign n15728 = ~n15719 & ~n15721 ;
  assign n15729 = ~n15422 & n15728 ;
  assign n15730 = ~n15727 & n15729 ;
  assign n15731 = n8355 & ~n15730 ;
  assign n15732 = ~n15327 & ~n15731 ;
  assign n15734 = \P4_IR_reg[21]/NET0131  & \P4_IR_reg[22]/NET0131  ;
  assign n15735 = \P4_IR_reg[24]/NET0131  & \P4_IR_reg[25]/NET0131  ;
  assign n15736 = \P4_IR_reg[26]/NET0131  & n15735 ;
  assign n15737 = n15734 & ~n15736 ;
  assign n15733 = \P4_IR_reg[27]/NET0131  & \P4_IR_reg[28]/NET0131  ;
  assign n15738 = ~\P4_IR_reg[19]/NET0131  & ~\P4_IR_reg[20]/NET0131  ;
  assign n15739 = n15733 & n15738 ;
  assign n15740 = n15737 & n15739 ;
  assign n15741 = ~\P4_IR_reg[23]/NET0131  & ~n15740 ;
  assign n15742 = \P3_rd_reg/NET0131  & ~n15741 ;
  assign n15743 = \P4_B_reg/NET0131  & ~n15742 ;
  assign n15744 = \P3_rd_reg/NET0131  & \P4_IR_reg[23]/NET0131  ;
  assign n15745 = ~\P4_IR_reg[27]/NET0131  & ~\P4_IR_reg[28]/NET0131  ;
  assign n15746 = \P2_P3_Datao_reg[29]/NET0131  & ~n15745 ;
  assign n15753 = \P4_IR_reg[29]/NET0131  & \P4_IR_reg[30]/NET0131  ;
  assign n15754 = \P4_reg3_reg[3]/NET0131  & \P4_reg3_reg[4]/NET0131  ;
  assign n15755 = \P4_reg3_reg[5]/NET0131  & n15754 ;
  assign n15756 = \P4_reg3_reg[6]/NET0131  & n15755 ;
  assign n15757 = \P4_reg3_reg[7]/NET0131  & n15756 ;
  assign n15758 = \P4_reg3_reg[8]/NET0131  & n15757 ;
  assign n15759 = \P4_reg3_reg[9]/NET0131  & n15758 ;
  assign n15760 = \P4_reg3_reg[10]/NET0131  & n15759 ;
  assign n15761 = \P4_reg3_reg[11]/NET0131  & n15760 ;
  assign n15762 = \P4_reg3_reg[12]/NET0131  & n15761 ;
  assign n15763 = \P4_reg3_reg[13]/NET0131  & n15762 ;
  assign n15764 = \P4_reg3_reg[14]/NET0131  & \P4_reg3_reg[15]/NET0131  ;
  assign n15765 = n15763 & n15764 ;
  assign n15766 = \P4_reg3_reg[16]/NET0131  & n15765 ;
  assign n15767 = \P4_reg3_reg[17]/NET0131  & \P4_reg3_reg[18]/NET0131  ;
  assign n15768 = \P4_reg3_reg[19]/NET0131  & \P4_reg3_reg[20]/NET0131  ;
  assign n15769 = \P4_reg3_reg[21]/NET0131  & \P4_reg3_reg[22]/NET0131  ;
  assign n15770 = n15768 & n15769 ;
  assign n15771 = n15767 & n15770 ;
  assign n15772 = n15766 & n15771 ;
  assign n15773 = \P4_reg3_reg[23]/NET0131  & \P4_reg3_reg[24]/NET0131  ;
  assign n15774 = n15772 & n15773 ;
  assign n15775 = \P4_reg3_reg[25]/NET0131  & \P4_reg3_reg[26]/NET0131  ;
  assign n15776 = \P4_reg3_reg[27]/NET0131  & n15775 ;
  assign n15777 = n15774 & n15776 ;
  assign n15778 = \P4_reg3_reg[28]/NET0131  & n15777 ;
  assign n15779 = n15753 & n15778 ;
  assign n15751 = ~\P4_IR_reg[29]/NET0131  & \P4_IR_reg[30]/NET0131  ;
  assign n15752 = \P4_reg2_reg[29]/NET0131  & n15751 ;
  assign n15747 = \P4_IR_reg[29]/NET0131  & ~\P4_IR_reg[30]/NET0131  ;
  assign n15748 = \P4_reg1_reg[29]/NET0131  & n15747 ;
  assign n15749 = ~\P4_IR_reg[29]/NET0131  & ~\P4_IR_reg[30]/NET0131  ;
  assign n15750 = \P4_reg0_reg[29]/NET0131  & n15749 ;
  assign n15780 = ~n15748 & ~n15750 ;
  assign n15781 = ~n15752 & n15780 ;
  assign n15782 = ~n15779 & n15781 ;
  assign n15783 = ~n15746 & ~n15782 ;
  assign n15784 = n15746 & n15782 ;
  assign n15785 = \P2_P3_Datao_reg[28]/NET0131  & ~n15745 ;
  assign n15789 = ~\P4_reg3_reg[28]/NET0131  & ~n15777 ;
  assign n15790 = ~n15778 & ~n15789 ;
  assign n15791 = n15753 & n15790 ;
  assign n15788 = \P4_reg2_reg[28]/NET0131  & n15751 ;
  assign n15786 = \P4_reg1_reg[28]/NET0131  & n15747 ;
  assign n15787 = \P4_reg0_reg[28]/NET0131  & n15749 ;
  assign n15792 = ~n15786 & ~n15787 ;
  assign n15793 = ~n15788 & n15792 ;
  assign n15794 = ~n15791 & n15793 ;
  assign n15795 = n15785 & n15794 ;
  assign n15796 = ~n15784 & ~n15795 ;
  assign n15797 = ~n15785 & ~n15794 ;
  assign n15798 = \P2_P3_Datao_reg[27]/NET0131  & ~n15745 ;
  assign n15802 = \P4_reg3_reg[25]/NET0131  & n15774 ;
  assign n15803 = \P4_reg3_reg[26]/NET0131  & n15802 ;
  assign n15804 = ~\P4_reg3_reg[27]/NET0131  & ~n15803 ;
  assign n15805 = ~n15777 & ~n15804 ;
  assign n15806 = n15753 & n15805 ;
  assign n15801 = \P4_reg2_reg[27]/NET0131  & n15751 ;
  assign n15799 = \P4_reg0_reg[27]/NET0131  & n15749 ;
  assign n15800 = \P4_reg1_reg[27]/NET0131  & n15747 ;
  assign n15807 = ~n15799 & ~n15800 ;
  assign n15808 = ~n15801 & n15807 ;
  assign n15809 = ~n15806 & n15808 ;
  assign n15810 = n15798 & n15809 ;
  assign n15811 = \P2_P3_Datao_reg[26]/NET0131  & ~n15745 ;
  assign n15815 = ~\P4_reg3_reg[26]/NET0131  & ~n15802 ;
  assign n15816 = ~n15803 & ~n15815 ;
  assign n15817 = n15753 & n15816 ;
  assign n15814 = \P4_reg1_reg[26]/NET0131  & n15747 ;
  assign n15812 = \P4_reg0_reg[26]/NET0131  & n15749 ;
  assign n15813 = \P4_reg2_reg[26]/NET0131  & n15751 ;
  assign n15818 = ~n15812 & ~n15813 ;
  assign n15819 = ~n15814 & n15818 ;
  assign n15820 = ~n15817 & n15819 ;
  assign n15821 = n15811 & n15820 ;
  assign n15822 = ~n15810 & ~n15821 ;
  assign n15823 = \P2_P3_Datao_reg[25]/NET0131  & ~n15745 ;
  assign n15827 = ~\P4_reg3_reg[25]/NET0131  & ~n15774 ;
  assign n15828 = ~n15802 & ~n15827 ;
  assign n15829 = n15753 & n15828 ;
  assign n15826 = \P4_reg2_reg[25]/NET0131  & n15751 ;
  assign n15824 = \P4_reg1_reg[25]/NET0131  & n15747 ;
  assign n15825 = \P4_reg0_reg[25]/NET0131  & n15749 ;
  assign n15830 = ~n15824 & ~n15825 ;
  assign n15831 = ~n15826 & n15830 ;
  assign n15832 = ~n15829 & n15831 ;
  assign n15833 = n15823 & n15832 ;
  assign n15834 = \P2_P3_Datao_reg[24]/NET0131  & ~n15745 ;
  assign n15838 = \P4_reg3_reg[23]/NET0131  & n15772 ;
  assign n15839 = ~\P4_reg3_reg[24]/NET0131  & ~n15838 ;
  assign n15840 = ~n15774 & ~n15839 ;
  assign n15841 = n15753 & n15840 ;
  assign n15837 = \P4_reg1_reg[24]/NET0131  & n15747 ;
  assign n15835 = \P4_reg0_reg[24]/NET0131  & n15749 ;
  assign n15836 = \P4_reg2_reg[24]/NET0131  & n15751 ;
  assign n15842 = ~n15835 & ~n15836 ;
  assign n15843 = ~n15837 & n15842 ;
  assign n15844 = ~n15841 & n15843 ;
  assign n15845 = n15834 & n15844 ;
  assign n15846 = ~n15833 & ~n15845 ;
  assign n15847 = \P2_P3_Datao_reg[23]/NET0131  & ~n15745 ;
  assign n15851 = ~\P4_reg3_reg[23]/NET0131  & ~n15772 ;
  assign n15852 = ~n15838 & ~n15851 ;
  assign n15853 = n15753 & n15852 ;
  assign n15850 = \P4_reg0_reg[23]/NET0131  & n15749 ;
  assign n15848 = \P4_reg1_reg[23]/NET0131  & n15747 ;
  assign n15849 = \P4_reg2_reg[23]/NET0131  & n15751 ;
  assign n15854 = ~n15848 & ~n15849 ;
  assign n15855 = ~n15850 & n15854 ;
  assign n15856 = ~n15853 & n15855 ;
  assign n15857 = n15847 & n15856 ;
  assign n15858 = \P2_P3_Datao_reg[22]/NET0131  & ~n15745 ;
  assign n15862 = \P4_reg3_reg[17]/NET0131  & n15766 ;
  assign n15863 = \P4_reg3_reg[18]/NET0131  & n15862 ;
  assign n15864 = \P4_reg3_reg[19]/NET0131  & n15863 ;
  assign n15865 = \P4_reg3_reg[20]/NET0131  & n15864 ;
  assign n15866 = \P4_reg3_reg[21]/NET0131  & n15865 ;
  assign n15867 = ~\P4_reg3_reg[22]/NET0131  & ~n15866 ;
  assign n15868 = ~n15772 & ~n15867 ;
  assign n15869 = n15753 & n15868 ;
  assign n15861 = \P4_reg2_reg[22]/NET0131  & n15751 ;
  assign n15859 = \P4_reg0_reg[22]/NET0131  & n15749 ;
  assign n15860 = \P4_reg1_reg[22]/NET0131  & n15747 ;
  assign n15870 = ~n15859 & ~n15860 ;
  assign n15871 = ~n15861 & n15870 ;
  assign n15872 = ~n15869 & n15871 ;
  assign n15873 = n15858 & n15872 ;
  assign n15874 = ~n15857 & ~n15873 ;
  assign n15875 = \P2_P3_Datao_reg[21]/NET0131  & ~n15745 ;
  assign n15879 = ~\P4_reg3_reg[21]/NET0131  & ~n15865 ;
  assign n15880 = ~n15866 & ~n15879 ;
  assign n15881 = n15753 & n15880 ;
  assign n15878 = \P4_reg2_reg[21]/NET0131  & n15751 ;
  assign n15876 = \P4_reg1_reg[21]/NET0131  & n15747 ;
  assign n15877 = \P4_reg0_reg[21]/NET0131  & n15749 ;
  assign n15882 = ~n15876 & ~n15877 ;
  assign n15883 = ~n15878 & n15882 ;
  assign n15884 = ~n15881 & n15883 ;
  assign n15885 = n15875 & n15884 ;
  assign n15886 = \P2_P3_Datao_reg[20]/NET0131  & ~n15745 ;
  assign n15890 = ~\P4_reg3_reg[20]/NET0131  & ~n15864 ;
  assign n15891 = ~n15865 & ~n15890 ;
  assign n15892 = n15753 & n15891 ;
  assign n15889 = \P4_reg0_reg[20]/NET0131  & n15749 ;
  assign n15887 = \P4_reg2_reg[20]/NET0131  & n15751 ;
  assign n15888 = \P4_reg1_reg[20]/NET0131  & n15747 ;
  assign n15893 = ~n15887 & ~n15888 ;
  assign n15894 = ~n15889 & n15893 ;
  assign n15895 = ~n15892 & n15894 ;
  assign n15896 = n15886 & n15895 ;
  assign n15897 = ~n15885 & ~n15896 ;
  assign n15898 = \P2_P3_Datao_reg[19]/NET0131  & ~n15745 ;
  assign n15899 = \P4_IR_reg[19]/NET0131  & n15745 ;
  assign n15900 = ~n15898 & ~n15899 ;
  assign n15904 = ~\P4_reg3_reg[19]/NET0131  & ~n15863 ;
  assign n15905 = ~n15864 & ~n15904 ;
  assign n15906 = n15753 & n15905 ;
  assign n15903 = \P4_reg2_reg[19]/NET0131  & n15751 ;
  assign n15901 = \P4_reg0_reg[19]/NET0131  & n15749 ;
  assign n15902 = \P4_reg1_reg[19]/NET0131  & n15747 ;
  assign n15907 = ~n15901 & ~n15902 ;
  assign n15908 = ~n15903 & n15907 ;
  assign n15909 = ~n15906 & n15908 ;
  assign n15910 = ~n15900 & n15909 ;
  assign n15911 = \P2_P3_Datao_reg[18]/NET0131  & ~n15745 ;
  assign n15912 = \P4_IR_reg[18]/NET0131  & n15745 ;
  assign n15913 = ~n15911 & ~n15912 ;
  assign n15917 = ~\P4_reg3_reg[18]/NET0131  & ~n15862 ;
  assign n15918 = ~n15863 & ~n15917 ;
  assign n15919 = n15753 & n15918 ;
  assign n15916 = \P4_reg0_reg[18]/NET0131  & n15749 ;
  assign n15914 = \P4_reg1_reg[18]/NET0131  & n15747 ;
  assign n15915 = \P4_reg2_reg[18]/NET0131  & n15751 ;
  assign n15920 = ~n15914 & ~n15915 ;
  assign n15921 = ~n15916 & n15920 ;
  assign n15922 = ~n15919 & n15921 ;
  assign n15923 = ~n15913 & n15922 ;
  assign n15924 = ~n15910 & ~n15923 ;
  assign n15925 = \P2_P3_Datao_reg[17]/NET0131  & ~n15745 ;
  assign n15926 = \P4_IR_reg[17]/NET0131  & n15745 ;
  assign n15927 = ~n15925 & ~n15926 ;
  assign n15931 = ~\P4_reg3_reg[17]/NET0131  & ~n15766 ;
  assign n15932 = ~n15862 & ~n15931 ;
  assign n15933 = n15753 & n15932 ;
  assign n15930 = \P4_reg1_reg[17]/NET0131  & n15747 ;
  assign n15928 = \P4_reg0_reg[17]/NET0131  & n15749 ;
  assign n15929 = \P4_reg2_reg[17]/NET0131  & n15751 ;
  assign n15934 = ~n15928 & ~n15929 ;
  assign n15935 = ~n15930 & n15934 ;
  assign n15936 = ~n15933 & n15935 ;
  assign n15937 = ~n15927 & n15936 ;
  assign n15938 = \P2_P3_Datao_reg[16]/NET0131  & ~n15745 ;
  assign n15939 = \P4_IR_reg[16]/NET0131  & n15745 ;
  assign n15940 = ~n15938 & ~n15939 ;
  assign n15944 = ~\P4_reg3_reg[16]/NET0131  & ~n15765 ;
  assign n15945 = ~n15766 & ~n15944 ;
  assign n15946 = n15753 & n15945 ;
  assign n15943 = \P4_reg1_reg[16]/NET0131  & n15747 ;
  assign n15941 = \P4_reg0_reg[16]/NET0131  & n15749 ;
  assign n15942 = \P4_reg2_reg[16]/NET0131  & n15751 ;
  assign n15947 = ~n15941 & ~n15942 ;
  assign n15948 = ~n15943 & n15947 ;
  assign n15949 = ~n15946 & n15948 ;
  assign n15950 = ~n15940 & n15949 ;
  assign n15951 = ~n15937 & ~n15950 ;
  assign n15952 = \P2_P3_Datao_reg[13]/NET0131  & ~n15745 ;
  assign n15953 = \P4_IR_reg[13]/NET0131  & n15745 ;
  assign n15954 = ~n15952 & ~n15953 ;
  assign n15958 = ~\P4_reg3_reg[13]/NET0131  & ~n15762 ;
  assign n15959 = ~n15763 & ~n15958 ;
  assign n15960 = n15753 & n15959 ;
  assign n15957 = \P4_reg2_reg[13]/NET0131  & n15751 ;
  assign n15955 = \P4_reg1_reg[13]/NET0131  & n15747 ;
  assign n15956 = \P4_reg0_reg[13]/NET0131  & n15749 ;
  assign n15961 = ~n15955 & ~n15956 ;
  assign n15962 = ~n15957 & n15961 ;
  assign n15963 = ~n15960 & n15962 ;
  assign n15964 = n15954 & ~n15963 ;
  assign n15965 = \P2_P3_Datao_reg[12]/NET0131  & ~n15745 ;
  assign n15966 = \P4_IR_reg[12]/NET0131  & n15745 ;
  assign n15967 = ~n15965 & ~n15966 ;
  assign n15971 = ~\P4_reg3_reg[12]/NET0131  & ~n15761 ;
  assign n15972 = ~n15762 & ~n15971 ;
  assign n15973 = n15753 & n15972 ;
  assign n15970 = \P4_reg1_reg[12]/NET0131  & n15747 ;
  assign n15968 = \P4_reg2_reg[12]/NET0131  & n15751 ;
  assign n15969 = \P4_reg0_reg[12]/NET0131  & n15749 ;
  assign n15974 = ~n15968 & ~n15969 ;
  assign n15975 = ~n15970 & n15974 ;
  assign n15976 = ~n15973 & n15975 ;
  assign n15977 = n15967 & ~n15976 ;
  assign n15978 = ~n15964 & ~n15977 ;
  assign n15979 = ~n15967 & n15976 ;
  assign n15980 = \P2_P3_Datao_reg[11]/NET0131  & ~n15745 ;
  assign n15981 = \P4_IR_reg[11]/NET0131  & n15745 ;
  assign n15982 = ~n15980 & ~n15981 ;
  assign n15986 = ~\P4_reg3_reg[11]/NET0131  & ~n15760 ;
  assign n15987 = ~n15761 & ~n15986 ;
  assign n15988 = n15753 & n15987 ;
  assign n15985 = \P4_reg2_reg[11]/NET0131  & n15751 ;
  assign n15983 = \P4_reg0_reg[11]/NET0131  & n15749 ;
  assign n15984 = \P4_reg1_reg[11]/NET0131  & n15747 ;
  assign n15989 = ~n15983 & ~n15984 ;
  assign n15990 = ~n15985 & n15989 ;
  assign n15991 = ~n15988 & n15990 ;
  assign n15992 = ~n15982 & n15991 ;
  assign n15993 = ~n15979 & ~n15992 ;
  assign n15994 = n15982 & ~n15991 ;
  assign n15995 = \P2_P3_Datao_reg[10]/NET0131  & ~n15745 ;
  assign n15996 = \P4_IR_reg[10]/NET0131  & n15745 ;
  assign n15997 = ~n15995 & ~n15996 ;
  assign n16001 = ~\P4_reg3_reg[10]/NET0131  & ~n15759 ;
  assign n16002 = ~n15760 & ~n16001 ;
  assign n16003 = n15753 & n16002 ;
  assign n16000 = \P4_reg0_reg[10]/NET0131  & n15749 ;
  assign n15998 = \P4_reg1_reg[10]/NET0131  & n15747 ;
  assign n15999 = \P4_reg2_reg[10]/NET0131  & n15751 ;
  assign n16004 = ~n15998 & ~n15999 ;
  assign n16005 = ~n16000 & n16004 ;
  assign n16006 = ~n16003 & n16005 ;
  assign n16007 = n15997 & ~n16006 ;
  assign n16008 = ~n15994 & ~n16007 ;
  assign n16009 = ~n15997 & n16006 ;
  assign n16010 = \P2_P3_Datao_reg[9]/NET0131  & ~n15745 ;
  assign n16011 = \P4_IR_reg[9]/NET0131  & n15745 ;
  assign n16012 = ~n16010 & ~n16011 ;
  assign n16016 = ~\P4_reg3_reg[9]/NET0131  & ~n15758 ;
  assign n16017 = ~n15759 & ~n16016 ;
  assign n16018 = n15753 & n16017 ;
  assign n16015 = \P4_reg0_reg[9]/NET0131  & n15749 ;
  assign n16013 = \P4_reg1_reg[9]/NET0131  & n15747 ;
  assign n16014 = \P4_reg2_reg[9]/NET0131  & n15751 ;
  assign n16019 = ~n16013 & ~n16014 ;
  assign n16020 = ~n16015 & n16019 ;
  assign n16021 = ~n16018 & n16020 ;
  assign n16022 = ~n16012 & n16021 ;
  assign n16023 = n16012 & ~n16021 ;
  assign n16024 = \P2_P3_Datao_reg[8]/NET0131  & ~n15745 ;
  assign n16025 = \P4_IR_reg[8]/NET0131  & n15745 ;
  assign n16026 = ~n16024 & ~n16025 ;
  assign n16030 = ~\P4_reg3_reg[8]/NET0131  & ~n15757 ;
  assign n16031 = ~n15758 & ~n16030 ;
  assign n16032 = n15753 & n16031 ;
  assign n16029 = \P4_reg1_reg[8]/NET0131  & n15747 ;
  assign n16027 = \P4_reg2_reg[8]/NET0131  & n15751 ;
  assign n16028 = \P4_reg0_reg[8]/NET0131  & n15749 ;
  assign n16033 = ~n16027 & ~n16028 ;
  assign n16034 = ~n16029 & n16033 ;
  assign n16035 = ~n16032 & n16034 ;
  assign n16036 = ~n16026 & n16035 ;
  assign n16037 = \P2_P3_Datao_reg[5]/NET0131  & ~n15745 ;
  assign n16038 = \P4_IR_reg[5]/NET0131  & n15745 ;
  assign n16039 = ~n16037 & ~n16038 ;
  assign n16043 = ~\P4_reg3_reg[5]/NET0131  & ~n15754 ;
  assign n16044 = ~n15755 & ~n16043 ;
  assign n16045 = n15753 & n16044 ;
  assign n16042 = \P4_reg2_reg[5]/NET0131  & n15751 ;
  assign n16040 = \P4_reg1_reg[5]/NET0131  & n15747 ;
  assign n16041 = \P4_reg0_reg[5]/NET0131  & n15749 ;
  assign n16046 = ~n16040 & ~n16041 ;
  assign n16047 = ~n16042 & n16046 ;
  assign n16048 = ~n16045 & n16047 ;
  assign n16049 = ~n16039 & n16048 ;
  assign n16050 = \P2_P3_Datao_reg[4]/NET0131  & ~n15745 ;
  assign n16051 = \P4_IR_reg[4]/NET0131  & n15745 ;
  assign n16052 = ~n16050 & ~n16051 ;
  assign n16056 = ~\P4_reg3_reg[3]/NET0131  & ~\P4_reg3_reg[4]/NET0131  ;
  assign n16057 = ~n15754 & ~n16056 ;
  assign n16058 = n15753 & n16057 ;
  assign n16055 = \P4_reg0_reg[4]/NET0131  & n15749 ;
  assign n16053 = \P4_reg2_reg[4]/NET0131  & n15751 ;
  assign n16054 = \P4_reg1_reg[4]/NET0131  & n15747 ;
  assign n16059 = ~n16053 & ~n16054 ;
  assign n16060 = ~n16055 & n16059 ;
  assign n16061 = ~n16058 & n16060 ;
  assign n16062 = ~n16052 & n16061 ;
  assign n16063 = ~n16049 & ~n16062 ;
  assign n16064 = n16052 & ~n16061 ;
  assign n16065 = \P4_reg2_reg[3]/NET0131  & n15751 ;
  assign n16066 = ~\P4_reg3_reg[3]/NET0131  & n15753 ;
  assign n16069 = ~n16065 & ~n16066 ;
  assign n16067 = \P4_reg1_reg[3]/NET0131  & n15747 ;
  assign n16068 = \P4_reg0_reg[3]/NET0131  & n15749 ;
  assign n16070 = ~n16067 & ~n16068 ;
  assign n16071 = n16069 & n16070 ;
  assign n16072 = \P2_P3_Datao_reg[3]/NET0131  & ~n15745 ;
  assign n16073 = \P4_IR_reg[3]/NET0131  & n15745 ;
  assign n16074 = ~n16072 & ~n16073 ;
  assign n16075 = ~n16071 & n16074 ;
  assign n16076 = n16071 & ~n16074 ;
  assign n16077 = \P4_reg0_reg[2]/NET0131  & n15749 ;
  assign n16078 = \P4_reg3_reg[2]/NET0131  & n15753 ;
  assign n16081 = ~n16077 & ~n16078 ;
  assign n16079 = \P4_reg1_reg[2]/NET0131  & n15747 ;
  assign n16080 = \P4_reg2_reg[2]/NET0131  & n15751 ;
  assign n16082 = ~n16079 & ~n16080 ;
  assign n16083 = n16081 & n16082 ;
  assign n16084 = \P2_P3_Datao_reg[2]/NET0131  & ~n15745 ;
  assign n16085 = \P4_IR_reg[2]/NET0131  & n15745 ;
  assign n16086 = ~n16084 & ~n16085 ;
  assign n16087 = n16083 & ~n16086 ;
  assign n16088 = ~n16083 & n16086 ;
  assign n16089 = \P4_reg1_reg[1]/NET0131  & n15747 ;
  assign n16090 = \P4_reg0_reg[1]/NET0131  & n15749 ;
  assign n16093 = ~n16089 & ~n16090 ;
  assign n16091 = \P4_reg3_reg[1]/NET0131  & n15753 ;
  assign n16092 = \P4_reg2_reg[1]/NET0131  & n15751 ;
  assign n16094 = ~n16091 & ~n16092 ;
  assign n16095 = n16093 & n16094 ;
  assign n16096 = \P2_P3_Datao_reg[1]/NET0131  & ~n15745 ;
  assign n16097 = \P4_IR_reg[1]/NET0131  & n15745 ;
  assign n16098 = ~n16096 & ~n16097 ;
  assign n16099 = ~n16095 & n16098 ;
  assign n16100 = n16095 & ~n16098 ;
  assign n16101 = \P2_P3_Datao_reg[0]/NET0131  & ~n15745 ;
  assign n16102 = \P4_IR_reg[0]/NET0131  & n15745 ;
  assign n16103 = ~n16101 & ~n16102 ;
  assign n16104 = \P4_reg1_reg[0]/NET0131  & n15747 ;
  assign n16105 = \P4_reg0_reg[0]/NET0131  & n15749 ;
  assign n16108 = ~n16104 & ~n16105 ;
  assign n16106 = \P4_reg2_reg[0]/NET0131  & n15751 ;
  assign n16107 = \P4_reg3_reg[0]/NET0131  & n15753 ;
  assign n16109 = ~n16106 & ~n16107 ;
  assign n16110 = n16108 & n16109 ;
  assign n16111 = ~n16103 & n16110 ;
  assign n16112 = ~n16100 & ~n16111 ;
  assign n16113 = ~n16099 & ~n16112 ;
  assign n16114 = ~n16088 & n16113 ;
  assign n16115 = ~n16087 & ~n16114 ;
  assign n16116 = ~n16076 & n16115 ;
  assign n16117 = ~n16075 & ~n16116 ;
  assign n16118 = ~n16064 & n16117 ;
  assign n16119 = n16063 & ~n16118 ;
  assign n16120 = \P2_P3_Datao_reg[6]/NET0131  & ~n15745 ;
  assign n16121 = \P4_IR_reg[6]/NET0131  & n15745 ;
  assign n16122 = ~n16120 & ~n16121 ;
  assign n16126 = ~\P4_reg3_reg[6]/NET0131  & ~n15755 ;
  assign n16127 = ~n15756 & ~n16126 ;
  assign n16128 = n15753 & n16127 ;
  assign n16125 = \P4_reg0_reg[6]/NET0131  & n15749 ;
  assign n16123 = \P4_reg2_reg[6]/NET0131  & n15751 ;
  assign n16124 = \P4_reg1_reg[6]/NET0131  & n15747 ;
  assign n16129 = ~n16123 & ~n16124 ;
  assign n16130 = ~n16125 & n16129 ;
  assign n16131 = ~n16128 & n16130 ;
  assign n16132 = n16122 & ~n16131 ;
  assign n16133 = n16039 & ~n16048 ;
  assign n16134 = ~n16132 & ~n16133 ;
  assign n16135 = ~n16119 & n16134 ;
  assign n16136 = \P2_P3_Datao_reg[7]/NET0131  & ~n15745 ;
  assign n16137 = \P4_IR_reg[7]/NET0131  & n15745 ;
  assign n16138 = ~n16136 & ~n16137 ;
  assign n16142 = ~\P4_reg3_reg[7]/NET0131  & ~n15756 ;
  assign n16143 = ~n15757 & ~n16142 ;
  assign n16144 = n15753 & n16143 ;
  assign n16141 = \P4_reg2_reg[7]/NET0131  & n15751 ;
  assign n16139 = \P4_reg0_reg[7]/NET0131  & n15749 ;
  assign n16140 = \P4_reg1_reg[7]/NET0131  & n15747 ;
  assign n16145 = ~n16139 & ~n16140 ;
  assign n16146 = ~n16141 & n16145 ;
  assign n16147 = ~n16144 & n16146 ;
  assign n16148 = ~n16138 & n16147 ;
  assign n16149 = ~n16122 & n16131 ;
  assign n16150 = ~n16148 & ~n16149 ;
  assign n16151 = ~n16135 & n16150 ;
  assign n16152 = n16026 & ~n16035 ;
  assign n16153 = n16138 & ~n16147 ;
  assign n16154 = ~n16152 & ~n16153 ;
  assign n16155 = ~n16151 & n16154 ;
  assign n16156 = ~n16036 & ~n16155 ;
  assign n16157 = ~n16023 & ~n16156 ;
  assign n16158 = ~n16022 & ~n16157 ;
  assign n16159 = ~n16009 & n16158 ;
  assign n16160 = n16008 & ~n16159 ;
  assign n16161 = n15993 & ~n16160 ;
  assign n16162 = n15978 & ~n16161 ;
  assign n16163 = \P2_P3_Datao_reg[15]/NET0131  & ~n15745 ;
  assign n16164 = \P4_IR_reg[15]/NET0131  & n15745 ;
  assign n16165 = ~n16163 & ~n16164 ;
  assign n16169 = \P4_reg3_reg[14]/NET0131  & n15763 ;
  assign n16170 = ~\P4_reg3_reg[15]/NET0131  & ~n16169 ;
  assign n16171 = ~n15765 & ~n16170 ;
  assign n16172 = n15753 & n16171 ;
  assign n16168 = \P4_reg0_reg[15]/NET0131  & n15749 ;
  assign n16166 = \P4_reg2_reg[15]/NET0131  & n15751 ;
  assign n16167 = \P4_reg1_reg[15]/NET0131  & n15747 ;
  assign n16173 = ~n16166 & ~n16167 ;
  assign n16174 = ~n16168 & n16173 ;
  assign n16175 = ~n16172 & n16174 ;
  assign n16176 = ~n16165 & n16175 ;
  assign n16177 = \P2_P3_Datao_reg[14]/NET0131  & ~n15745 ;
  assign n16178 = \P4_IR_reg[14]/NET0131  & n15745 ;
  assign n16179 = ~n16177 & ~n16178 ;
  assign n16183 = ~\P4_reg3_reg[14]/NET0131  & ~n15763 ;
  assign n16184 = ~n16169 & ~n16183 ;
  assign n16185 = n15753 & n16184 ;
  assign n16182 = \P4_reg2_reg[14]/NET0131  & n15751 ;
  assign n16180 = \P4_reg1_reg[14]/NET0131  & n15747 ;
  assign n16181 = \P4_reg0_reg[14]/NET0131  & n15749 ;
  assign n16186 = ~n16180 & ~n16181 ;
  assign n16187 = ~n16182 & n16186 ;
  assign n16188 = ~n16185 & n16187 ;
  assign n16189 = ~n16179 & n16188 ;
  assign n16190 = ~n15954 & n15963 ;
  assign n16191 = ~n16189 & ~n16190 ;
  assign n16192 = ~n16176 & n16191 ;
  assign n16193 = ~n16162 & n16192 ;
  assign n16194 = n16165 & ~n16175 ;
  assign n16195 = n16179 & ~n16188 ;
  assign n16196 = ~n16194 & ~n16195 ;
  assign n16197 = ~n16176 & ~n16196 ;
  assign n16198 = ~n16193 & ~n16197 ;
  assign n16199 = n15951 & ~n16198 ;
  assign n16200 = n15927 & ~n15936 ;
  assign n16201 = n15940 & ~n15949 ;
  assign n16202 = ~n15937 & n16201 ;
  assign n16203 = ~n16200 & ~n16202 ;
  assign n16204 = ~n16199 & n16203 ;
  assign n16205 = n15924 & ~n16204 ;
  assign n16206 = n15900 & ~n15909 ;
  assign n16207 = n15913 & ~n15922 ;
  assign n16208 = ~n15910 & n16207 ;
  assign n16209 = ~n16206 & ~n16208 ;
  assign n16210 = ~n16205 & n16209 ;
  assign n16211 = n15897 & ~n16210 ;
  assign n16212 = ~n15875 & ~n15884 ;
  assign n16213 = ~n15886 & ~n15895 ;
  assign n16214 = ~n16212 & ~n16213 ;
  assign n16215 = ~n15885 & ~n16214 ;
  assign n16216 = ~n16211 & ~n16215 ;
  assign n16217 = n15874 & ~n16216 ;
  assign n16218 = ~n15847 & ~n15856 ;
  assign n16219 = ~n15858 & ~n15872 ;
  assign n16220 = ~n16218 & ~n16219 ;
  assign n16221 = ~n15857 & ~n16220 ;
  assign n16222 = ~n16217 & ~n16221 ;
  assign n16223 = n15846 & ~n16222 ;
  assign n16224 = n15822 & n16223 ;
  assign n16226 = ~n15823 & ~n15832 ;
  assign n16227 = ~n15834 & ~n15844 ;
  assign n16228 = ~n16226 & ~n16227 ;
  assign n16229 = ~n15833 & ~n16228 ;
  assign n16230 = ~n15821 & n16229 ;
  assign n16225 = ~n15798 & ~n15809 ;
  assign n16231 = ~n15811 & ~n15820 ;
  assign n16232 = ~n16225 & ~n16231 ;
  assign n16233 = ~n16230 & n16232 ;
  assign n16234 = ~n15810 & ~n16233 ;
  assign n16235 = ~n16224 & ~n16234 ;
  assign n16236 = ~n15797 & n16235 ;
  assign n16237 = n15796 & ~n16236 ;
  assign n16238 = ~n15783 & ~n16237 ;
  assign n16241 = \P4_reg1_reg[31]/NET0131  & n15747 ;
  assign n16239 = \P4_reg2_reg[31]/NET0131  & n15751 ;
  assign n16240 = \P4_reg0_reg[31]/NET0131  & n15749 ;
  assign n16242 = ~n16239 & ~n16240 ;
  assign n16243 = ~n16241 & n16242 ;
  assign n16244 = ~n15779 & n16243 ;
  assign n16245 = \P2_P3_Datao_reg[30]/NET0131  & ~n15745 ;
  assign n16246 = n16244 & ~n16245 ;
  assign n16247 = ~n16238 & n16246 ;
  assign n16248 = ~\P4_IR_reg[19]/NET0131  & ~n16247 ;
  assign n16249 = \P4_IR_reg[19]/NET0131  & n16247 ;
  assign n16250 = ~n16248 & ~n16249 ;
  assign n16435 = ~\P4_B_reg/NET0131  & n16250 ;
  assign n16436 = \P4_IR_reg[20]/NET0131  & n15734 ;
  assign n16437 = ~n16435 & n16436 ;
  assign n16299 = \P4_reg0_reg[30]/NET0131  & n15749 ;
  assign n16297 = \P4_reg2_reg[30]/NET0131  & n15751 ;
  assign n16298 = \P4_reg1_reg[30]/NET0131  & n15747 ;
  assign n16300 = ~n16297 & ~n16298 ;
  assign n16301 = ~n16299 & n16300 ;
  assign n16302 = ~n15779 & n16301 ;
  assign n16326 = n16245 & n16302 ;
  assign n16327 = n16244 & ~n16326 ;
  assign n16303 = ~n16245 & ~n16302 ;
  assign n16423 = n16238 & ~n16303 ;
  assign n16424 = n16327 & ~n16423 ;
  assign n16428 = ~\P4_IR_reg[20]/NET0131  & ~\P4_IR_reg[21]/NET0131  ;
  assign n16429 = ~\P4_IR_reg[19]/NET0131  & n16428 ;
  assign n16430 = ~n16424 & n16429 ;
  assign n16254 = \P4_IR_reg[19]/NET0131  & ~\P4_IR_reg[20]/NET0131  ;
  assign n16425 = ~\P4_IR_reg[21]/NET0131  & ~\P4_IR_reg[22]/NET0131  ;
  assign n16426 = n16254 & n16425 ;
  assign n16427 = n16424 & n16426 ;
  assign n16255 = \P4_B_reg/NET0131  & \P4_IR_reg[22]/NET0131  ;
  assign n16256 = ~n16254 & n16255 ;
  assign n16276 = n15834 & ~n15844 ;
  assign n16277 = ~n15834 & n15844 ;
  assign n16278 = ~n16276 & ~n16277 ;
  assign n16316 = ~n15910 & ~n16206 ;
  assign n16356 = ~n16278 & n16316 ;
  assign n16328 = ~n15783 & ~n15784 ;
  assign n16357 = n16327 & n16328 ;
  assign n16358 = n16356 & n16357 ;
  assign n16307 = n15847 & ~n15856 ;
  assign n16308 = ~n15847 & n15856 ;
  assign n16309 = ~n16307 & ~n16308 ;
  assign n16304 = ~n15913 & ~n15922 ;
  assign n16305 = n15913 & n15922 ;
  assign n16306 = ~n16304 & ~n16305 ;
  assign n16353 = ~n16303 & ~n16306 ;
  assign n16354 = ~n16309 & n16353 ;
  assign n16260 = n15823 & ~n15832 ;
  assign n16261 = ~n15823 & n15832 ;
  assign n16262 = ~n16260 & ~n16261 ;
  assign n16313 = ~n15927 & ~n15936 ;
  assign n16314 = n15927 & n15936 ;
  assign n16315 = ~n16313 & ~n16314 ;
  assign n16335 = ~n16189 & ~n16195 ;
  assign n16263 = ~n15954 & ~n15963 ;
  assign n16264 = n15954 & n15963 ;
  assign n16265 = ~n16263 & ~n16264 ;
  assign n16279 = n15967 & n15976 ;
  assign n16280 = ~n15967 & ~n15976 ;
  assign n16281 = ~n16279 & ~n16280 ;
  assign n16267 = ~n15982 & ~n15991 ;
  assign n16268 = n15982 & n15991 ;
  assign n16269 = ~n16267 & ~n16268 ;
  assign n16283 = ~n15997 & ~n16006 ;
  assign n16284 = n15997 & n16006 ;
  assign n16285 = ~n16283 & ~n16284 ;
  assign n16270 = n16012 & n16021 ;
  assign n16271 = ~n16012 & ~n16021 ;
  assign n16272 = ~n16270 & ~n16271 ;
  assign n16290 = ~n16026 & ~n16035 ;
  assign n16291 = n16026 & n16035 ;
  assign n16292 = ~n16290 & ~n16291 ;
  assign n16286 = ~n16148 & ~n16153 ;
  assign n16293 = ~n16132 & ~n16149 ;
  assign n16282 = ~n16087 & ~n16088 ;
  assign n16336 = n16112 & n16282 ;
  assign n16287 = ~n16075 & ~n16076 ;
  assign n16288 = n16103 & ~n16110 ;
  assign n16289 = ~n16099 & ~n16288 ;
  assign n16337 = n16287 & n16289 ;
  assign n16338 = n16336 & n16337 ;
  assign n16266 = ~n16062 & ~n16064 ;
  assign n16294 = n16039 & n16048 ;
  assign n16295 = ~n16039 & ~n16048 ;
  assign n16296 = ~n16294 & ~n16295 ;
  assign n16339 = n16266 & ~n16296 ;
  assign n16340 = n16338 & n16339 ;
  assign n16341 = n16293 & n16340 ;
  assign n16342 = n16286 & n16341 ;
  assign n16343 = ~n16292 & n16342 ;
  assign n16344 = ~n16272 & n16343 ;
  assign n16345 = ~n16285 & n16344 ;
  assign n16346 = ~n16269 & n16345 ;
  assign n16347 = ~n16281 & n16346 ;
  assign n16348 = ~n16265 & n16347 ;
  assign n16349 = n16335 & n16348 ;
  assign n16323 = ~n16165 & ~n16175 ;
  assign n16324 = n16165 & n16175 ;
  assign n16325 = ~n16323 & ~n16324 ;
  assign n16332 = ~n15940 & ~n15949 ;
  assign n16333 = n15940 & n15949 ;
  assign n16334 = ~n16332 & ~n16333 ;
  assign n16350 = ~n16325 & ~n16334 ;
  assign n16351 = n16349 & n16350 ;
  assign n16352 = ~n16315 & n16351 ;
  assign n16355 = ~n16262 & n16352 ;
  assign n16359 = n16354 & n16355 ;
  assign n16362 = n16358 & n16359 ;
  assign n16273 = n15875 & ~n15884 ;
  assign n16274 = ~n15875 & n15884 ;
  assign n16275 = ~n16273 & ~n16274 ;
  assign n16317 = n15798 & ~n15809 ;
  assign n16318 = ~n15798 & n15809 ;
  assign n16319 = ~n16317 & ~n16318 ;
  assign n16363 = ~n16275 & ~n16319 ;
  assign n16364 = n16362 & n16363 ;
  assign n16320 = n15858 & ~n15872 ;
  assign n16321 = ~n15858 & n15872 ;
  assign n16322 = ~n16320 & ~n16321 ;
  assign n16329 = ~n15811 & n15820 ;
  assign n16330 = n15811 & ~n15820 ;
  assign n16331 = ~n16329 & ~n16330 ;
  assign n16257 = n15886 & ~n15895 ;
  assign n16258 = ~n15886 & n15895 ;
  assign n16259 = ~n16257 & ~n16258 ;
  assign n16310 = ~n15785 & n15794 ;
  assign n16311 = n15785 & ~n15794 ;
  assign n16312 = ~n16310 & ~n16311 ;
  assign n16360 = ~n16259 & ~n16312 ;
  assign n16361 = ~n16331 & n16360 ;
  assign n16365 = ~n16322 & n16361 ;
  assign n16366 = n16364 & n16365 ;
  assign n16368 = \P4_IR_reg[19]/NET0131  & n16366 ;
  assign n16367 = ~\P4_IR_reg[19]/NET0131  & ~n16366 ;
  assign n16369 = \P4_IR_reg[20]/NET0131  & ~n16367 ;
  assign n16370 = ~n16368 & n16369 ;
  assign n16371 = ~n16256 & ~n16370 ;
  assign n16372 = ~\P4_IR_reg[21]/NET0131  & ~n16371 ;
  assign n16378 = ~n16212 & ~n16219 ;
  assign n16379 = ~n16206 & ~n16213 ;
  assign n16380 = ~n16200 & ~n16207 ;
  assign n16381 = ~n16009 & ~n16022 ;
  assign n16382 = ~n16087 & ~n16100 ;
  assign n16383 = ~n16289 & n16382 ;
  assign n16384 = ~n16075 & ~n16088 ;
  assign n16385 = ~n16383 & n16384 ;
  assign n16386 = ~n16076 & ~n16385 ;
  assign n16387 = ~n16064 & ~n16386 ;
  assign n16388 = n16063 & ~n16387 ;
  assign n16389 = n16134 & ~n16388 ;
  assign n16390 = n16150 & ~n16389 ;
  assign n16391 = n16154 & ~n16390 ;
  assign n16392 = ~n16036 & ~n16391 ;
  assign n16393 = ~n16023 & ~n16392 ;
  assign n16394 = n16381 & ~n16393 ;
  assign n16395 = n16008 & ~n16394 ;
  assign n16396 = n15993 & ~n16395 ;
  assign n16397 = n15978 & ~n16396 ;
  assign n16398 = n16192 & ~n16397 ;
  assign n16399 = ~n16197 & ~n16201 ;
  assign n16400 = ~n16398 & n16399 ;
  assign n16401 = n15951 & ~n16400 ;
  assign n16402 = n16380 & ~n16401 ;
  assign n16403 = n15924 & ~n16402 ;
  assign n16404 = n16379 & ~n16403 ;
  assign n16405 = n15897 & ~n16404 ;
  assign n16406 = n16378 & ~n16405 ;
  assign n16407 = n15874 & ~n16406 ;
  assign n16376 = ~n16226 & ~n16231 ;
  assign n16408 = ~n16218 & ~n16227 ;
  assign n16409 = n16376 & n16408 ;
  assign n16410 = ~n16407 & n16409 ;
  assign n16377 = ~n15846 & n16376 ;
  assign n16411 = n15822 & ~n16377 ;
  assign n16412 = ~n16410 & n16411 ;
  assign n16373 = ~n15783 & ~n16303 ;
  assign n16375 = ~n15797 & ~n16225 ;
  assign n16413 = n16373 & n16375 ;
  assign n16414 = ~n16412 & n16413 ;
  assign n16374 = ~n15796 & n16373 ;
  assign n16415 = n16327 & ~n16374 ;
  assign n16416 = ~n16414 & n16415 ;
  assign n16418 = \P4_IR_reg[19]/NET0131  & n16416 ;
  assign n16417 = ~\P4_IR_reg[19]/NET0131  & ~n16416 ;
  assign n16419 = ~n16255 & ~n16417 ;
  assign n16420 = ~n16418 & n16419 ;
  assign n16421 = ~\P4_IR_reg[20]/NET0131  & \P4_IR_reg[21]/NET0131  ;
  assign n16422 = ~n16420 & n16421 ;
  assign n16438 = ~n16372 & ~n16422 ;
  assign n16439 = ~n16427 & n16438 ;
  assign n16440 = ~n16430 & n16439 ;
  assign n16251 = \P4_IR_reg[20]/NET0131  & \P4_IR_reg[21]/NET0131  ;
  assign n16252 = ~\P4_IR_reg[22]/NET0131  & n16251 ;
  assign n16253 = ~n16250 & n16252 ;
  assign n16431 = ~\P4_B_reg/NET0131  & ~n16424 ;
  assign n16432 = \P4_IR_reg[19]/NET0131  & \P4_IR_reg[22]/NET0131  ;
  assign n16433 = n16428 & n16432 ;
  assign n16434 = ~n16431 & n16433 ;
  assign n16441 = ~n16253 & ~n16434 ;
  assign n16442 = n16440 & n16441 ;
  assign n16443 = ~n16437 & n16442 ;
  assign n16444 = n15744 & ~n16443 ;
  assign n16445 = ~n15743 & ~n16444 ;
  assign n16448 = \P1_P3_PhyAddrPointer_reg[1]/NET0131  & \P1_P3_PhyAddrPointer_reg[2]/NET0131  ;
  assign n16449 = ~\P1_P3_PhyAddrPointer_reg[3]/NET0131  & ~n16448 ;
  assign n16450 = \P1_P3_PhyAddrPointer_reg[3]/NET0131  & n16448 ;
  assign n16451 = ~n16449 & ~n16450 ;
  assign n16452 = ~\P1_P3_PhyAddrPointer_reg[0]/NET0131  & n16448 ;
  assign n16453 = \P1_P3_PhyAddrPointer_reg[2]/NET0131  & \P1_P3_PhyAddrPointer_reg[3]/NET0131  ;
  assign n16454 = \P1_P3_PhyAddrPointer_reg[4]/NET0131  & n16453 ;
  assign n16455 = \P1_P3_PhyAddrPointer_reg[5]/NET0131  & n16454 ;
  assign n16456 = \P1_P3_PhyAddrPointer_reg[6]/NET0131  & n16455 ;
  assign n16457 = \P1_P3_PhyAddrPointer_reg[7]/NET0131  & n16456 ;
  assign n16458 = \P1_P3_PhyAddrPointer_reg[8]/NET0131  & n16457 ;
  assign n16459 = \P1_P3_PhyAddrPointer_reg[9]/NET0131  & n16458 ;
  assign n16460 = \P1_P3_PhyAddrPointer_reg[10]/NET0131  & n16459 ;
  assign n16461 = \P1_P3_PhyAddrPointer_reg[11]/NET0131  & n16460 ;
  assign n16462 = \P1_P3_PhyAddrPointer_reg[12]/NET0131  & n16461 ;
  assign n16463 = \P1_P3_PhyAddrPointer_reg[13]/NET0131  & n16462 ;
  assign n16464 = \P1_P3_PhyAddrPointer_reg[14]/NET0131  & n16463 ;
  assign n16465 = \P1_P3_PhyAddrPointer_reg[15]/NET0131  & n16464 ;
  assign n16466 = \P1_P3_PhyAddrPointer_reg[16]/NET0131  & n16465 ;
  assign n16467 = \P1_P3_PhyAddrPointer_reg[17]/NET0131  & n16466 ;
  assign n16468 = \P1_P3_PhyAddrPointer_reg[18]/NET0131  & n16467 ;
  assign n16469 = \P1_P3_PhyAddrPointer_reg[19]/NET0131  & n16468 ;
  assign n16470 = \P1_P3_PhyAddrPointer_reg[20]/NET0131  & n16469 ;
  assign n16471 = \P1_P3_PhyAddrPointer_reg[21]/NET0131  & n16470 ;
  assign n16472 = \P1_P3_PhyAddrPointer_reg[22]/NET0131  & n16471 ;
  assign n16473 = \P1_P3_PhyAddrPointer_reg[23]/NET0131  & n16472 ;
  assign n16474 = \P1_P3_PhyAddrPointer_reg[24]/NET0131  & n16473 ;
  assign n16475 = \P1_P3_PhyAddrPointer_reg[25]/NET0131  & n16474 ;
  assign n16476 = \P1_P3_PhyAddrPointer_reg[26]/NET0131  & n16475 ;
  assign n16477 = \P1_P3_PhyAddrPointer_reg[27]/NET0131  & n16476 ;
  assign n16478 = \P1_P3_PhyAddrPointer_reg[28]/NET0131  & n16477 ;
  assign n16479 = \P1_P3_PhyAddrPointer_reg[29]/NET0131  & n16478 ;
  assign n16480 = \P1_P3_PhyAddrPointer_reg[30]/NET0131  & n16479 ;
  assign n16481 = \P1_P3_PhyAddrPointer_reg[1]/NET0131  & n16480 ;
  assign n16482 = ~\P1_P3_PhyAddrPointer_reg[31]/NET0131  & ~n16481 ;
  assign n16483 = \P1_P3_PhyAddrPointer_reg[31]/NET0131  & n16481 ;
  assign n16484 = ~n16482 & ~n16483 ;
  assign n16485 = ~n16452 & n16484 ;
  assign n16487 = ~n16451 & n16485 ;
  assign n16486 = n16451 & ~n16485 ;
  assign n16488 = ~\P1_P3_DataWidth_reg[1]/NET0131  & ~n16486 ;
  assign n16489 = ~n16487 & n16488 ;
  assign n16447 = \P1_P3_DataWidth_reg[1]/NET0131  & ~\P1_P3_rEIP_reg[3]/NET0131  ;
  assign n16490 = n9245 & ~n16447 ;
  assign n16491 = ~n16489 & n16490 ;
  assign n16497 = \P1_P3_rEIP_reg[3]/NET0131  & ~n9195 ;
  assign n16500 = ~n9075 & n9085 ;
  assign n16505 = ~\P1_P3_DataWidth_reg[1]/NET0131  & ~n8741 ;
  assign n16501 = ~\P1_P3_EBX_reg[0]/NET0131  & ~\P1_P3_EBX_reg[1]/NET0131  ;
  assign n16502 = ~\P1_P3_EBX_reg[2]/NET0131  & n16501 ;
  assign n16503 = \P1_P3_EBX_reg[31]/NET0131  & ~n16502 ;
  assign n16504 = \P1_P3_EBX_reg[3]/NET0131  & n16503 ;
  assign n16506 = ~\P1_P3_EBX_reg[3]/NET0131  & ~n16503 ;
  assign n16507 = ~n16504 & ~n16506 ;
  assign n16508 = ~n16505 & n16507 ;
  assign n16509 = \P1_P3_rEIP_reg[1]/NET0131  & \P1_P3_rEIP_reg[2]/NET0131  ;
  assign n16511 = ~\P1_P3_rEIP_reg[3]/NET0131  & ~n16509 ;
  assign n16510 = \P1_P3_rEIP_reg[3]/NET0131  & n16509 ;
  assign n16512 = ~\P1_P3_DataWidth_reg[1]/NET0131  & ~n16510 ;
  assign n16513 = ~n16511 & n16512 ;
  assign n16514 = ~n8741 & n16513 ;
  assign n16515 = ~n16508 & ~n16514 ;
  assign n16516 = n16500 & ~n16515 ;
  assign n16498 = ~n9075 & n9082 ;
  assign n16499 = ~n9180 & n16498 ;
  assign n16517 = ~\P1_P3_DataWidth_reg[1]/NET0131  & n9096 ;
  assign n16518 = \P1_P3_EBX_reg[3]/NET0131  & ~n16517 ;
  assign n16519 = n9096 & n16513 ;
  assign n16520 = ~n16518 & ~n16519 ;
  assign n16521 = n9236 & ~n16520 ;
  assign n16522 = ~n16499 & ~n16521 ;
  assign n16523 = ~n16516 & n16522 ;
  assign n16524 = ~n16497 & n16523 ;
  assign n16525 = n9241 & ~n16524 ;
  assign n16446 = \P1_P3_PhyAddrPointer_reg[3]/NET0131  & n10031 ;
  assign n16492 = ~\P1_P3_State2_reg[1]/NET0131  & n8734 ;
  assign n16493 = ~n8732 & ~n16492 ;
  assign n16494 = ~n10036 & ~n10046 ;
  assign n16495 = n16493 & n16494 ;
  assign n16496 = \P1_P3_rEIP_reg[3]/NET0131  & ~n16495 ;
  assign n16526 = ~n16446 & ~n16496 ;
  assign n16527 = ~n16525 & n16526 ;
  assign n16528 = ~n16491 & n16527 ;
  assign n16531 = \P1_P3_PhyAddrPointer_reg[1]/NET0131  & n16461 ;
  assign n16532 = \P1_P3_PhyAddrPointer_reg[12]/NET0131  & n16531 ;
  assign n16533 = \P1_P3_PhyAddrPointer_reg[13]/NET0131  & n16532 ;
  assign n16534 = \P1_P3_PhyAddrPointer_reg[14]/NET0131  & n16533 ;
  assign n16535 = \P1_P3_PhyAddrPointer_reg[15]/NET0131  & n16534 ;
  assign n16536 = \P1_P3_PhyAddrPointer_reg[16]/NET0131  & n16535 ;
  assign n16537 = \P1_P3_PhyAddrPointer_reg[17]/NET0131  & n16536 ;
  assign n16538 = \P1_P3_PhyAddrPointer_reg[18]/NET0131  & n16537 ;
  assign n16539 = \P1_P3_PhyAddrPointer_reg[19]/NET0131  & n16538 ;
  assign n16540 = ~\P1_P3_PhyAddrPointer_reg[20]/NET0131  & ~n16539 ;
  assign n16541 = \P1_P3_PhyAddrPointer_reg[1]/NET0131  & n16470 ;
  assign n16542 = ~n16540 & ~n16541 ;
  assign n16543 = ~\P1_P3_PhyAddrPointer_reg[19]/NET0131  & ~n16538 ;
  assign n16544 = ~n16539 & ~n16543 ;
  assign n16545 = ~\P1_P3_PhyAddrPointer_reg[17]/NET0131  & ~n16536 ;
  assign n16546 = ~n16537 & ~n16545 ;
  assign n16547 = ~\P1_P3_PhyAddrPointer_reg[0]/NET0131  & n16532 ;
  assign n16548 = \P1_P3_PhyAddrPointer_reg[13]/NET0131  & n16547 ;
  assign n16549 = n16465 & n16548 ;
  assign n16550 = \P1_P3_PhyAddrPointer_reg[16]/NET0131  & n16549 ;
  assign n16551 = ~n16546 & n16550 ;
  assign n16552 = ~\P1_P3_PhyAddrPointer_reg[18]/NET0131  & ~n16537 ;
  assign n16553 = ~n16538 & ~n16552 ;
  assign n16554 = n16551 & ~n16553 ;
  assign n16555 = ~n16544 & n16554 ;
  assign n16556 = n16484 & ~n16555 ;
  assign n16558 = n16542 & ~n16556 ;
  assign n16557 = ~n16542 & n16556 ;
  assign n16559 = ~\P1_P3_DataWidth_reg[1]/NET0131  & ~n16557 ;
  assign n16560 = ~n16558 & n16559 ;
  assign n16530 = \P1_P3_DataWidth_reg[1]/NET0131  & ~\P1_P3_rEIP_reg[20]/NET0131  ;
  assign n16561 = n9245 & ~n16530 ;
  assign n16562 = ~n16560 & n16561 ;
  assign n16596 = ~\P1_P3_EBX_reg[3]/NET0131  & n16502 ;
  assign n16597 = ~\P1_P3_EBX_reg[4]/NET0131  & n16596 ;
  assign n16598 = ~\P1_P3_EBX_reg[5]/NET0131  & n16597 ;
  assign n16599 = ~\P1_P3_EBX_reg[6]/NET0131  & n16598 ;
  assign n16600 = ~\P1_P3_EBX_reg[7]/NET0131  & n16599 ;
  assign n16601 = ~\P1_P3_EBX_reg[8]/NET0131  & n16600 ;
  assign n16602 = ~\P1_P3_EBX_reg[9]/NET0131  & n16601 ;
  assign n16603 = ~\P1_P3_EBX_reg[10]/NET0131  & n16602 ;
  assign n16604 = ~\P1_P3_EBX_reg[11]/NET0131  & n16603 ;
  assign n16605 = ~\P1_P3_EBX_reg[12]/NET0131  & n16604 ;
  assign n16606 = ~\P1_P3_EBX_reg[13]/NET0131  & n16605 ;
  assign n16607 = ~\P1_P3_EBX_reg[14]/NET0131  & n16606 ;
  assign n16608 = ~\P1_P3_EBX_reg[15]/NET0131  & n16607 ;
  assign n16609 = ~\P1_P3_EBX_reg[16]/NET0131  & n16608 ;
  assign n16610 = ~\P1_P3_EBX_reg[17]/NET0131  & n16609 ;
  assign n16611 = ~\P1_P3_EBX_reg[18]/NET0131  & n16610 ;
  assign n16612 = ~\P1_P3_EBX_reg[19]/NET0131  & n16611 ;
  assign n16613 = \P1_P3_EBX_reg[31]/NET0131  & ~n16612 ;
  assign n16615 = ~\P1_P3_EBX_reg[20]/NET0131  & n16613 ;
  assign n16614 = \P1_P3_EBX_reg[20]/NET0131  & ~n16613 ;
  assign n16616 = ~n16505 & ~n16614 ;
  assign n16617 = ~n16615 & n16616 ;
  assign n16570 = \P1_P3_rEIP_reg[4]/NET0131  & n16510 ;
  assign n16571 = \P1_P3_rEIP_reg[5]/NET0131  & n16570 ;
  assign n16572 = \P1_P3_rEIP_reg[6]/NET0131  & n16571 ;
  assign n16573 = \P1_P3_rEIP_reg[7]/NET0131  & n16572 ;
  assign n16574 = \P1_P3_rEIP_reg[8]/NET0131  & n16573 ;
  assign n16575 = \P1_P3_rEIP_reg[9]/NET0131  & n16574 ;
  assign n16576 = \P1_P3_rEIP_reg[10]/NET0131  & n16575 ;
  assign n16577 = \P1_P3_rEIP_reg[11]/NET0131  & n16576 ;
  assign n16578 = \P1_P3_rEIP_reg[12]/NET0131  & n16577 ;
  assign n16579 = \P1_P3_rEIP_reg[13]/NET0131  & n16578 ;
  assign n16580 = \P1_P3_rEIP_reg[14]/NET0131  & n16579 ;
  assign n16581 = \P1_P3_rEIP_reg[15]/NET0131  & n16580 ;
  assign n16582 = \P1_P3_rEIP_reg[16]/NET0131  & n16581 ;
  assign n16583 = \P1_P3_rEIP_reg[17]/NET0131  & n16582 ;
  assign n16584 = \P1_P3_rEIP_reg[18]/NET0131  & n16583 ;
  assign n16585 = \P1_P3_rEIP_reg[19]/NET0131  & n16584 ;
  assign n16586 = ~\P1_P3_rEIP_reg[20]/NET0131  & ~n16585 ;
  assign n16587 = \P1_P3_rEIP_reg[20]/NET0131  & n16585 ;
  assign n16588 = ~n16586 & ~n16587 ;
  assign n16589 = n16505 & ~n16588 ;
  assign n16618 = n16500 & ~n16589 ;
  assign n16619 = ~n16617 & n16618 ;
  assign n16564 = n9075 & ~n9115 ;
  assign n16565 = ~n9116 & ~n16564 ;
  assign n16566 = \P1_P3_rEIP_reg[20]/NET0131  & ~n16565 ;
  assign n16590 = ~\P1_P3_EBX_reg[20]/NET0131  & ~n16505 ;
  assign n16591 = n9162 & ~n16590 ;
  assign n16592 = ~n16589 & n16591 ;
  assign n16567 = ~n9075 & n9095 ;
  assign n16568 = \P1_P3_EBX_reg[20]/NET0131  & n16567 ;
  assign n16569 = \P1_P3_rEIP_reg[20]/NET0131  & n9075 ;
  assign n16593 = ~n16568 & ~n16569 ;
  assign n16594 = ~n16592 & n16593 ;
  assign n16595 = n9079 & ~n16594 ;
  assign n16620 = ~n16566 & ~n16595 ;
  assign n16621 = ~n16619 & n16620 ;
  assign n16622 = n9241 & ~n16621 ;
  assign n16529 = \P1_P3_PhyAddrPointer_reg[20]/NET0131  & n10031 ;
  assign n16563 = \P1_P3_rEIP_reg[20]/NET0131  & ~n16495 ;
  assign n16623 = ~n16529 & ~n16563 ;
  assign n16624 = ~n16622 & n16623 ;
  assign n16625 = ~n16562 & n16624 ;
  assign n16628 = ~\P1_P3_PhyAddrPointer_reg[21]/NET0131  & ~n16541 ;
  assign n16629 = \P1_P3_PhyAddrPointer_reg[1]/NET0131  & n16471 ;
  assign n16630 = ~n16628 & ~n16629 ;
  assign n16631 = ~n16542 & n16555 ;
  assign n16632 = n16484 & ~n16631 ;
  assign n16634 = n16630 & ~n16632 ;
  assign n16633 = ~n16630 & n16632 ;
  assign n16635 = ~\P1_P3_DataWidth_reg[1]/NET0131  & ~n16633 ;
  assign n16636 = ~n16634 & n16635 ;
  assign n16627 = \P1_P3_DataWidth_reg[1]/NET0131  & ~\P1_P3_rEIP_reg[21]/NET0131  ;
  assign n16637 = n9245 & ~n16627 ;
  assign n16638 = ~n16636 & n16637 ;
  assign n16640 = \P1_P3_rEIP_reg[21]/NET0131  & ~n9195 ;
  assign n16641 = ~\P1_P3_EBX_reg[21]/NET0131  & ~n16517 ;
  assign n16642 = n9079 & ~n16641 ;
  assign n16643 = ~\P1_P3_EBX_reg[20]/NET0131  & n16612 ;
  assign n16644 = \P1_P3_EBX_reg[31]/NET0131  & ~n16643 ;
  assign n16646 = ~\P1_P3_EBX_reg[21]/NET0131  & n16644 ;
  assign n16645 = \P1_P3_EBX_reg[21]/NET0131  & ~n16644 ;
  assign n16647 = ~n16505 & ~n16645 ;
  assign n16648 = ~n16646 & n16647 ;
  assign n16649 = n9085 & ~n16648 ;
  assign n16650 = ~n16642 & ~n16649 ;
  assign n16652 = ~\P1_P3_rEIP_reg[21]/NET0131  & ~n16587 ;
  assign n16653 = \P1_P3_rEIP_reg[21]/NET0131  & n16587 ;
  assign n16654 = ~n16652 & ~n16653 ;
  assign n16651 = n9095 & n16642 ;
  assign n16655 = n16505 & ~n16651 ;
  assign n16656 = ~n16654 & n16655 ;
  assign n16657 = ~n9075 & ~n16656 ;
  assign n16658 = ~n16650 & n16657 ;
  assign n16659 = ~n16640 & ~n16658 ;
  assign n16660 = n9241 & ~n16659 ;
  assign n16626 = \P1_P3_PhyAddrPointer_reg[21]/NET0131  & n10031 ;
  assign n16639 = \P1_P3_rEIP_reg[21]/NET0131  & ~n16495 ;
  assign n16661 = ~n16626 & ~n16639 ;
  assign n16662 = ~n16660 & n16661 ;
  assign n16663 = ~n16638 & n16662 ;
  assign n16666 = ~n16630 & n16631 ;
  assign n16667 = n16484 & ~n16666 ;
  assign n16668 = ~\P1_P3_PhyAddrPointer_reg[22]/NET0131  & ~n16629 ;
  assign n16669 = \P1_P3_PhyAddrPointer_reg[22]/NET0131  & n16629 ;
  assign n16670 = ~n16668 & ~n16669 ;
  assign n16672 = n16667 & ~n16670 ;
  assign n16671 = ~n16667 & n16670 ;
  assign n16673 = ~\P1_P3_DataWidth_reg[1]/NET0131  & ~n16671 ;
  assign n16674 = ~n16672 & n16673 ;
  assign n16665 = \P1_P3_DataWidth_reg[1]/NET0131  & ~\P1_P3_rEIP_reg[22]/NET0131  ;
  assign n16675 = n9245 & ~n16665 ;
  assign n16676 = ~n16674 & n16675 ;
  assign n16691 = ~\P1_P3_EBX_reg[21]/NET0131  & n16643 ;
  assign n16692 = \P1_P3_EBX_reg[31]/NET0131  & ~n16691 ;
  assign n16694 = ~\P1_P3_EBX_reg[22]/NET0131  & n16692 ;
  assign n16693 = \P1_P3_EBX_reg[22]/NET0131  & ~n16692 ;
  assign n16695 = ~n16505 & ~n16693 ;
  assign n16696 = ~n16694 & n16695 ;
  assign n16681 = ~\P1_P3_rEIP_reg[22]/NET0131  & ~n16653 ;
  assign n16682 = \P1_P3_rEIP_reg[22]/NET0131  & n16653 ;
  assign n16683 = ~n16681 & ~n16682 ;
  assign n16684 = n16505 & ~n16683 ;
  assign n16697 = n16500 & ~n16684 ;
  assign n16698 = ~n16696 & n16697 ;
  assign n16678 = \P1_P3_rEIP_reg[22]/NET0131  & ~n16565 ;
  assign n16685 = ~\P1_P3_EBX_reg[22]/NET0131  & ~n16505 ;
  assign n16686 = n9162 & ~n16685 ;
  assign n16687 = ~n16684 & n16686 ;
  assign n16679 = \P1_P3_EBX_reg[22]/NET0131  & n16567 ;
  assign n16680 = \P1_P3_rEIP_reg[22]/NET0131  & n9075 ;
  assign n16688 = ~n16679 & ~n16680 ;
  assign n16689 = ~n16687 & n16688 ;
  assign n16690 = n9079 & ~n16689 ;
  assign n16699 = ~n16678 & ~n16690 ;
  assign n16700 = ~n16698 & n16699 ;
  assign n16701 = n9241 & ~n16700 ;
  assign n16664 = \P1_P3_PhyAddrPointer_reg[22]/NET0131  & n10031 ;
  assign n16677 = \P1_P3_rEIP_reg[22]/NET0131  & ~n16495 ;
  assign n16702 = ~n16664 & ~n16677 ;
  assign n16703 = ~n16701 & n16702 ;
  assign n16704 = ~n16676 & n16703 ;
  assign n16707 = n16666 & ~n16670 ;
  assign n16708 = n16484 & ~n16707 ;
  assign n16709 = ~\P1_P3_PhyAddrPointer_reg[23]/NET0131  & ~n16669 ;
  assign n16710 = \P1_P3_PhyAddrPointer_reg[23]/NET0131  & n16669 ;
  assign n16711 = ~n16709 & ~n16710 ;
  assign n16713 = ~n16708 & n16711 ;
  assign n16712 = n16708 & ~n16711 ;
  assign n16714 = ~\P1_P3_DataWidth_reg[1]/NET0131  & ~n16712 ;
  assign n16715 = ~n16713 & n16714 ;
  assign n16706 = \P1_P3_DataWidth_reg[1]/NET0131  & ~\P1_P3_rEIP_reg[23]/NET0131  ;
  assign n16716 = n9245 & ~n16706 ;
  assign n16717 = ~n16715 & n16716 ;
  assign n16719 = \P1_P3_rEIP_reg[23]/NET0131  & ~n9195 ;
  assign n16720 = ~\P1_P3_EBX_reg[23]/NET0131  & ~n16517 ;
  assign n16721 = n9079 & ~n16720 ;
  assign n16722 = ~\P1_P3_EBX_reg[22]/NET0131  & n16691 ;
  assign n16723 = \P1_P3_EBX_reg[31]/NET0131  & ~n16722 ;
  assign n16725 = ~\P1_P3_EBX_reg[23]/NET0131  & n16723 ;
  assign n16724 = \P1_P3_EBX_reg[23]/NET0131  & ~n16723 ;
  assign n16726 = ~n16505 & ~n16724 ;
  assign n16727 = ~n16725 & n16726 ;
  assign n16728 = n9085 & ~n16727 ;
  assign n16729 = ~n16721 & ~n16728 ;
  assign n16731 = ~\P1_P3_rEIP_reg[23]/NET0131  & ~n16682 ;
  assign n16732 = \P1_P3_rEIP_reg[23]/NET0131  & n16682 ;
  assign n16733 = ~n16731 & ~n16732 ;
  assign n16730 = n9095 & n16721 ;
  assign n16734 = n16505 & ~n16730 ;
  assign n16735 = ~n16733 & n16734 ;
  assign n16736 = ~n9075 & ~n16735 ;
  assign n16737 = ~n16729 & n16736 ;
  assign n16738 = ~n16719 & ~n16737 ;
  assign n16739 = n9241 & ~n16738 ;
  assign n16705 = \P1_P3_PhyAddrPointer_reg[23]/NET0131  & n10031 ;
  assign n16718 = \P1_P3_rEIP_reg[23]/NET0131  & ~n16495 ;
  assign n16740 = ~n16705 & ~n16718 ;
  assign n16741 = ~n16739 & n16740 ;
  assign n16742 = ~n16717 & n16741 ;
  assign n16745 = n16707 & ~n16711 ;
  assign n16746 = n16484 & ~n16745 ;
  assign n16747 = ~\P1_P3_PhyAddrPointer_reg[24]/NET0131  & ~n16710 ;
  assign n16748 = \P1_P3_PhyAddrPointer_reg[24]/NET0131  & n16710 ;
  assign n16749 = ~n16747 & ~n16748 ;
  assign n16751 = n16746 & ~n16749 ;
  assign n16750 = ~n16746 & n16749 ;
  assign n16752 = ~\P1_P3_DataWidth_reg[1]/NET0131  & ~n16750 ;
  assign n16753 = ~n16751 & n16752 ;
  assign n16744 = \P1_P3_DataWidth_reg[1]/NET0131  & ~\P1_P3_rEIP_reg[24]/NET0131  ;
  assign n16754 = n9245 & ~n16744 ;
  assign n16755 = ~n16753 & n16754 ;
  assign n16758 = \P1_P3_DataWidth_reg[1]/NET0131  & \P1_P3_EBX_reg[24]/NET0131  ;
  assign n16760 = ~\P1_P3_rEIP_reg[24]/NET0131  & ~n16732 ;
  assign n16759 = \P1_P3_rEIP_reg[24]/NET0131  & n16732 ;
  assign n16761 = ~\P1_P3_DataWidth_reg[1]/NET0131  & ~n16759 ;
  assign n16762 = ~n16760 & n16761 ;
  assign n16763 = ~n16758 & ~n16762 ;
  assign n16764 = n9096 & ~n16763 ;
  assign n16765 = \P1_P3_EBX_reg[24]/NET0131  & ~n9095 ;
  assign n16766 = n8741 & n16765 ;
  assign n16767 = ~n16764 & ~n16766 ;
  assign n16768 = ~n9075 & ~n16767 ;
  assign n16757 = \P1_P3_EBX_reg[24]/NET0131  & n16567 ;
  assign n16769 = \P1_P3_rEIP_reg[24]/NET0131  & n9075 ;
  assign n16770 = ~n16757 & ~n16769 ;
  assign n16771 = ~n16768 & n16770 ;
  assign n16772 = n9079 & ~n16771 ;
  assign n16756 = \P1_P3_rEIP_reg[24]/NET0131  & ~n16565 ;
  assign n16773 = ~\P1_P3_EBX_reg[23]/NET0131  & n16722 ;
  assign n16774 = \P1_P3_EBX_reg[31]/NET0131  & ~n16773 ;
  assign n16776 = \P1_P3_EBX_reg[24]/NET0131  & n16774 ;
  assign n16775 = ~\P1_P3_EBX_reg[24]/NET0131  & ~n16774 ;
  assign n16777 = ~n16505 & ~n16775 ;
  assign n16778 = ~n16776 & n16777 ;
  assign n16779 = ~n8741 & n16762 ;
  assign n16780 = ~n16778 & ~n16779 ;
  assign n16781 = n16500 & ~n16780 ;
  assign n16782 = ~n16756 & ~n16781 ;
  assign n16783 = ~n16772 & n16782 ;
  assign n16784 = n9241 & ~n16783 ;
  assign n16743 = \P1_P3_PhyAddrPointer_reg[24]/NET0131  & n10031 ;
  assign n16785 = \P1_P3_rEIP_reg[24]/NET0131  & ~n16495 ;
  assign n16786 = ~n16743 & ~n16785 ;
  assign n16787 = ~n16784 & n16786 ;
  assign n16788 = ~n16755 & n16787 ;
  assign n16791 = n16745 & ~n16749 ;
  assign n16792 = ~\P1_P3_PhyAddrPointer_reg[25]/NET0131  & ~n16748 ;
  assign n16793 = \P1_P3_PhyAddrPointer_reg[1]/NET0131  & n16475 ;
  assign n16794 = ~n16792 & ~n16793 ;
  assign n16795 = n16791 & ~n16794 ;
  assign n16796 = n16484 & ~n16795 ;
  assign n16797 = ~\P1_P3_PhyAddrPointer_reg[26]/NET0131  & ~n16793 ;
  assign n16798 = \P1_P3_PhyAddrPointer_reg[26]/NET0131  & n16793 ;
  assign n16799 = ~n16797 & ~n16798 ;
  assign n16801 = n16796 & ~n16799 ;
  assign n16800 = ~n16796 & n16799 ;
  assign n16802 = ~\P1_P3_DataWidth_reg[1]/NET0131  & ~n16800 ;
  assign n16803 = ~n16801 & n16802 ;
  assign n16790 = \P1_P3_DataWidth_reg[1]/NET0131  & ~\P1_P3_rEIP_reg[26]/NET0131  ;
  assign n16804 = n9245 & ~n16790 ;
  assign n16805 = ~n16803 & n16804 ;
  assign n16812 = ~\P1_P3_EBX_reg[24]/NET0131  & n16773 ;
  assign n16813 = ~\P1_P3_EBX_reg[25]/NET0131  & n16812 ;
  assign n16814 = \P1_P3_EBX_reg[31]/NET0131  & ~n16813 ;
  assign n16816 = ~\P1_P3_EBX_reg[26]/NET0131  & n16814 ;
  assign n16815 = \P1_P3_EBX_reg[26]/NET0131  & ~n16814 ;
  assign n16817 = ~n16505 & ~n16815 ;
  assign n16818 = ~n16816 & n16817 ;
  assign n16807 = \P1_P3_rEIP_reg[25]/NET0131  & n16759 ;
  assign n16808 = ~\P1_P3_rEIP_reg[26]/NET0131  & ~n16807 ;
  assign n16809 = \P1_P3_rEIP_reg[26]/NET0131  & n16807 ;
  assign n16810 = ~n16808 & ~n16809 ;
  assign n16811 = n16505 & ~n16810 ;
  assign n16819 = n16500 & ~n16811 ;
  assign n16820 = ~n16818 & n16819 ;
  assign n16821 = \P1_P3_rEIP_reg[26]/NET0131  & ~n9195 ;
  assign n16823 = ~n9095 & n16811 ;
  assign n16822 = ~\P1_P3_EBX_reg[26]/NET0131  & ~n16517 ;
  assign n16824 = n9236 & ~n16822 ;
  assign n16825 = ~n16823 & n16824 ;
  assign n16826 = ~n16821 & ~n16825 ;
  assign n16827 = ~n16820 & n16826 ;
  assign n16828 = n9241 & ~n16827 ;
  assign n16789 = \P1_P3_PhyAddrPointer_reg[26]/NET0131  & n10031 ;
  assign n16806 = \P1_P3_rEIP_reg[26]/NET0131  & ~n16495 ;
  assign n16829 = ~n16789 & ~n16806 ;
  assign n16830 = ~n16828 & n16829 ;
  assign n16831 = ~n16805 & n16830 ;
  assign n16834 = ~\P1_P3_PhyAddrPointer_reg[27]/NET0131  & ~n16798 ;
  assign n16835 = \P1_P3_PhyAddrPointer_reg[27]/NET0131  & n16798 ;
  assign n16836 = ~n16834 & ~n16835 ;
  assign n16837 = n16795 & ~n16799 ;
  assign n16838 = n16484 & ~n16837 ;
  assign n16840 = n16836 & ~n16838 ;
  assign n16839 = ~n16836 & n16838 ;
  assign n16841 = ~\P1_P3_DataWidth_reg[1]/NET0131  & ~n16839 ;
  assign n16842 = ~n16840 & n16841 ;
  assign n16833 = \P1_P3_DataWidth_reg[1]/NET0131  & ~\P1_P3_rEIP_reg[27]/NET0131  ;
  assign n16843 = n9245 & ~n16833 ;
  assign n16844 = ~n16842 & n16843 ;
  assign n16859 = ~\P1_P3_EBX_reg[26]/NET0131  & n16813 ;
  assign n16860 = \P1_P3_EBX_reg[31]/NET0131  & ~n16859 ;
  assign n16862 = ~\P1_P3_EBX_reg[27]/NET0131  & n16860 ;
  assign n16861 = \P1_P3_EBX_reg[27]/NET0131  & ~n16860 ;
  assign n16863 = ~n16505 & ~n16861 ;
  assign n16864 = ~n16862 & n16863 ;
  assign n16849 = \P1_P3_rEIP_reg[27]/NET0131  & n16809 ;
  assign n16850 = ~\P1_P3_rEIP_reg[27]/NET0131  & ~n16809 ;
  assign n16851 = ~n16849 & ~n16850 ;
  assign n16852 = n16505 & ~n16851 ;
  assign n16865 = n16500 & ~n16852 ;
  assign n16866 = ~n16864 & n16865 ;
  assign n16846 = \P1_P3_rEIP_reg[27]/NET0131  & ~n16565 ;
  assign n16853 = ~\P1_P3_EBX_reg[27]/NET0131  & ~n16505 ;
  assign n16854 = n9162 & ~n16853 ;
  assign n16855 = ~n16852 & n16854 ;
  assign n16847 = \P1_P3_rEIP_reg[27]/NET0131  & n9075 ;
  assign n16848 = \P1_P3_EBX_reg[27]/NET0131  & n16567 ;
  assign n16856 = ~n16847 & ~n16848 ;
  assign n16857 = ~n16855 & n16856 ;
  assign n16858 = n9079 & ~n16857 ;
  assign n16867 = ~n16846 & ~n16858 ;
  assign n16868 = ~n16866 & n16867 ;
  assign n16869 = n9241 & ~n16868 ;
  assign n16832 = \P1_P3_PhyAddrPointer_reg[27]/NET0131  & n10031 ;
  assign n16845 = \P1_P3_rEIP_reg[27]/NET0131  & ~n16495 ;
  assign n16870 = ~n16832 & ~n16845 ;
  assign n16871 = ~n16869 & n16870 ;
  assign n16872 = ~n16844 & n16871 ;
  assign n16896 = ~n16836 & n16837 ;
  assign n16897 = n16484 & ~n16896 ;
  assign n16898 = ~\P1_P3_PhyAddrPointer_reg[28]/NET0131  & ~n16835 ;
  assign n16899 = \P1_P3_PhyAddrPointer_reg[28]/NET0131  & n16835 ;
  assign n16900 = ~n16898 & ~n16899 ;
  assign n16902 = ~n16897 & n16900 ;
  assign n16901 = n16897 & ~n16900 ;
  assign n16903 = ~\P1_P3_DataWidth_reg[1]/NET0131  & ~n16901 ;
  assign n16904 = ~n16902 & n16903 ;
  assign n16895 = \P1_P3_DataWidth_reg[1]/NET0131  & ~\P1_P3_rEIP_reg[28]/NET0131  ;
  assign n16905 = n9245 & ~n16895 ;
  assign n16906 = ~n16904 & n16905 ;
  assign n16878 = ~\P1_P3_EBX_reg[27]/NET0131  & n16859 ;
  assign n16879 = \P1_P3_EBX_reg[31]/NET0131  & ~n16878 ;
  assign n16881 = ~\P1_P3_EBX_reg[28]/NET0131  & n16879 ;
  assign n16880 = \P1_P3_EBX_reg[28]/NET0131  & ~n16879 ;
  assign n16882 = ~n16505 & ~n16880 ;
  assign n16883 = ~n16881 & n16882 ;
  assign n16874 = ~\P1_P3_rEIP_reg[28]/NET0131  & ~n16849 ;
  assign n16875 = \P1_P3_rEIP_reg[28]/NET0131  & n16849 ;
  assign n16876 = ~n16874 & ~n16875 ;
  assign n16877 = n16505 & ~n16876 ;
  assign n16884 = n16500 & ~n16877 ;
  assign n16885 = ~n16883 & n16884 ;
  assign n16886 = \P1_P3_rEIP_reg[28]/NET0131  & ~n9195 ;
  assign n16888 = ~n9095 & n16877 ;
  assign n16887 = ~\P1_P3_EBX_reg[28]/NET0131  & ~n16517 ;
  assign n16889 = n9236 & ~n16887 ;
  assign n16890 = ~n16888 & n16889 ;
  assign n16891 = ~n16886 & ~n16890 ;
  assign n16892 = ~n16885 & n16891 ;
  assign n16893 = n9241 & ~n16892 ;
  assign n16873 = \P1_P3_PhyAddrPointer_reg[28]/NET0131  & n10031 ;
  assign n16894 = \P1_P3_rEIP_reg[28]/NET0131  & ~n16495 ;
  assign n16907 = ~n16873 & ~n16894 ;
  assign n16908 = ~n16893 & n16907 ;
  assign n16909 = ~n16906 & n16908 ;
  assign n16912 = ~\P1_P3_PhyAddrPointer_reg[1]/NET0131  & ~\P1_P3_PhyAddrPointer_reg[2]/NET0131  ;
  assign n16913 = ~n16448 & ~n16912 ;
  assign n16914 = \P1_P3_PhyAddrPointer_reg[0]/NET0131  & n16484 ;
  assign n16915 = \P1_P3_PhyAddrPointer_reg[1]/NET0131  & ~n16914 ;
  assign n16916 = n16484 & ~n16915 ;
  assign n16918 = ~n16913 & n16916 ;
  assign n16917 = n16913 & ~n16916 ;
  assign n16919 = ~\P1_P3_DataWidth_reg[1]/NET0131  & ~n16917 ;
  assign n16920 = ~n16918 & n16919 ;
  assign n16911 = \P1_P3_DataWidth_reg[1]/NET0131  & ~\P1_P3_rEIP_reg[2]/NET0131  ;
  assign n16921 = n9245 & ~n16911 ;
  assign n16922 = ~n16920 & n16921 ;
  assign n16924 = \P1_P3_rEIP_reg[2]/NET0131  & ~n9195 ;
  assign n16926 = ~\P1_P3_rEIP_reg[1]/NET0131  & ~\P1_P3_rEIP_reg[2]/NET0131  ;
  assign n16927 = ~\P1_P3_DataWidth_reg[1]/NET0131  & ~n16509 ;
  assign n16928 = ~n16926 & n16927 ;
  assign n16929 = ~n8741 & n16928 ;
  assign n16930 = \P1_P3_EBX_reg[31]/NET0131  & ~n16501 ;
  assign n16931 = ~\P1_P3_EBX_reg[2]/NET0131  & ~n16930 ;
  assign n16932 = \P1_P3_EBX_reg[2]/NET0131  & n16930 ;
  assign n16933 = ~n16931 & ~n16932 ;
  assign n16934 = ~n16505 & n16933 ;
  assign n16935 = ~n16929 & ~n16934 ;
  assign n16936 = n16500 & ~n16935 ;
  assign n16925 = n9104 & n16498 ;
  assign n16937 = \P1_P3_EBX_reg[2]/NET0131  & ~n16517 ;
  assign n16938 = n9096 & n16928 ;
  assign n16939 = ~n16937 & ~n16938 ;
  assign n16940 = n9236 & ~n16939 ;
  assign n16941 = ~n16925 & ~n16940 ;
  assign n16942 = ~n16936 & n16941 ;
  assign n16943 = ~n16924 & n16942 ;
  assign n16944 = n9241 & ~n16943 ;
  assign n16910 = \P1_P3_PhyAddrPointer_reg[2]/NET0131  & n10031 ;
  assign n16923 = \P1_P3_rEIP_reg[2]/NET0131  & ~n16495 ;
  assign n16945 = ~n16910 & ~n16923 ;
  assign n16946 = ~n16944 & n16945 ;
  assign n16947 = ~n16922 & n16946 ;
  assign n16949 = ~n9160 & n9241 ;
  assign n16950 = n15306 & n15312 ;
  assign n16951 = ~n10038 & ~n16950 ;
  assign n16952 = n10037 & ~n16951 ;
  assign n16948 = n9104 & n10046 ;
  assign n16953 = \P1_P3_InstQueueRd_Addr_reg[2]/NET0131  & ~n15317 ;
  assign n16954 = ~n16948 & ~n16953 ;
  assign n16955 = ~n16952 & n16954 ;
  assign n16956 = ~n16949 & n16955 ;
  assign n16958 = ~n9189 & n9241 ;
  assign n16959 = ~\P1_P3_Flush_reg/NET0131  & \P1_P3_InstQueueRd_Addr_reg[3]/NET0131  ;
  assign n16960 = ~n16950 & ~n16959 ;
  assign n16961 = n10037 & ~n16960 ;
  assign n16957 = ~n9180 & n10046 ;
  assign n16962 = \P1_P3_InstQueueRd_Addr_reg[3]/NET0131  & ~n15317 ;
  assign n16963 = ~n16957 & ~n16962 ;
  assign n16964 = ~n16961 & n16963 ;
  assign n16965 = ~n16958 & n16964 ;
  assign n16966 = ~n8732 & ~n10030 ;
  assign n16967 = ~n8733 & ~n10037 ;
  assign n16968 = n16966 & n16967 ;
  assign n16969 = \P1_P3_EAX_reg[11]/NET0131  & ~n16968 ;
  assign n16972 = \P1_P3_EAX_reg[0]/NET0131  & \P1_P3_EAX_reg[1]/NET0131  ;
  assign n16973 = \P1_P3_EAX_reg[2]/NET0131  & n16972 ;
  assign n16974 = \P1_P3_EAX_reg[3]/NET0131  & n16973 ;
  assign n16975 = \P1_P3_EAX_reg[4]/NET0131  & n16974 ;
  assign n16976 = \P1_P3_EAX_reg[5]/NET0131  & n16975 ;
  assign n16977 = \P1_P3_EAX_reg[6]/NET0131  & n16976 ;
  assign n16978 = \P1_P3_EAX_reg[7]/NET0131  & n16977 ;
  assign n16979 = \P1_P3_EAX_reg[8]/NET0131  & n16978 ;
  assign n16980 = \P1_P3_EAX_reg[9]/NET0131  & n16979 ;
  assign n16981 = \P1_P3_EAX_reg[10]/NET0131  & n16980 ;
  assign n16982 = n9106 & n9111 ;
  assign n16983 = ~n16981 & n16982 ;
  assign n16984 = n9049 & n9060 ;
  assign n16985 = n9087 & ~n16982 ;
  assign n16986 = ~n9060 & ~n16985 ;
  assign n16987 = ~n16984 & ~n16986 ;
  assign n16988 = ~n9089 & ~n16987 ;
  assign n16989 = ~n16983 & n16988 ;
  assign n16990 = \P1_P3_EAX_reg[11]/NET0131  & ~n16989 ;
  assign n16995 = \P1_P3_InstQueue_reg[11][3]/NET0131  & n8763 ;
  assign n16996 = \P1_P3_InstQueue_reg[6][3]/NET0131  & n8745 ;
  assign n17009 = ~n16995 & ~n16996 ;
  assign n16997 = \P1_P3_InstQueue_reg[3][3]/NET0131  & n8777 ;
  assign n16998 = \P1_P3_InstQueue_reg[8][3]/NET0131  & n8754 ;
  assign n17010 = ~n16997 & ~n16998 ;
  assign n17017 = n17009 & n17010 ;
  assign n16991 = \P1_P3_InstQueue_reg[4][3]/NET0131  & n8752 ;
  assign n16992 = \P1_P3_InstQueue_reg[9][3]/NET0131  & n8748 ;
  assign n17007 = ~n16991 & ~n16992 ;
  assign n16993 = \P1_P3_InstQueue_reg[7][3]/NET0131  & n8779 ;
  assign n16994 = \P1_P3_InstQueue_reg[13][3]/NET0131  & n8765 ;
  assign n17008 = ~n16993 & ~n16994 ;
  assign n17018 = n17007 & n17008 ;
  assign n17019 = n17017 & n17018 ;
  assign n17003 = \P1_P3_InstQueue_reg[14][3]/NET0131  & n8760 ;
  assign n17004 = \P1_P3_InstQueue_reg[2][3]/NET0131  & n8767 ;
  assign n17013 = ~n17003 & ~n17004 ;
  assign n17005 = \P1_P3_InstQueue_reg[10][3]/NET0131  & n8769 ;
  assign n17006 = \P1_P3_InstQueue_reg[0][3]/NET0131  & n8781 ;
  assign n17014 = ~n17005 & ~n17006 ;
  assign n17015 = n17013 & n17014 ;
  assign n16999 = \P1_P3_InstQueue_reg[5][3]/NET0131  & n8771 ;
  assign n17000 = \P1_P3_InstQueue_reg[12][3]/NET0131  & n8757 ;
  assign n17011 = ~n16999 & ~n17000 ;
  assign n17001 = \P1_P3_InstQueue_reg[15][3]/NET0131  & n8775 ;
  assign n17002 = \P1_P3_InstQueue_reg[1][3]/NET0131  & n8773 ;
  assign n17012 = ~n17001 & ~n17002 ;
  assign n17016 = n17011 & n17012 ;
  assign n17020 = n17015 & n17016 ;
  assign n17021 = n17019 & n17020 ;
  assign n17022 = n16984 & ~n17021 ;
  assign n16970 = \P1_buf2_reg[11]/NET0131  & n9088 ;
  assign n16971 = ~n9087 & n16970 ;
  assign n17023 = ~\P1_P3_EAX_reg[11]/NET0131  & n16981 ;
  assign n17024 = n16982 & n17023 ;
  assign n17025 = ~n16971 & ~n17024 ;
  assign n17026 = ~n17022 & n17025 ;
  assign n17027 = ~n16990 & n17026 ;
  assign n17028 = n9241 & ~n17027 ;
  assign n17029 = ~n16969 & ~n17028 ;
  assign n17030 = n9241 & ~n16988 ;
  assign n17031 = n16968 & ~n17030 ;
  assign n17032 = \P1_P3_EAX_reg[12]/NET0131  & ~n17031 ;
  assign n17035 = \P1_P3_EAX_reg[11]/NET0131  & n16981 ;
  assign n17036 = ~\P1_P3_EAX_reg[12]/NET0131  & ~n17035 ;
  assign n17037 = \P1_P3_EAX_reg[12]/NET0131  & n17035 ;
  assign n17038 = n16982 & ~n17037 ;
  assign n17039 = ~n17036 & n17038 ;
  assign n17033 = \P1_buf2_reg[12]/NET0131  & n9088 ;
  assign n17034 = ~n9087 & n17033 ;
  assign n17044 = \P1_P3_InstQueue_reg[11][4]/NET0131  & n8763 ;
  assign n17045 = \P1_P3_InstQueue_reg[6][4]/NET0131  & n8745 ;
  assign n17058 = ~n17044 & ~n17045 ;
  assign n17046 = \P1_P3_InstQueue_reg[3][4]/NET0131  & n8777 ;
  assign n17047 = \P1_P3_InstQueue_reg[8][4]/NET0131  & n8754 ;
  assign n17059 = ~n17046 & ~n17047 ;
  assign n17066 = n17058 & n17059 ;
  assign n17040 = \P1_P3_InstQueue_reg[4][4]/NET0131  & n8752 ;
  assign n17041 = \P1_P3_InstQueue_reg[9][4]/NET0131  & n8748 ;
  assign n17056 = ~n17040 & ~n17041 ;
  assign n17042 = \P1_P3_InstQueue_reg[7][4]/NET0131  & n8779 ;
  assign n17043 = \P1_P3_InstQueue_reg[13][4]/NET0131  & n8765 ;
  assign n17057 = ~n17042 & ~n17043 ;
  assign n17067 = n17056 & n17057 ;
  assign n17068 = n17066 & n17067 ;
  assign n17052 = \P1_P3_InstQueue_reg[14][4]/NET0131  & n8760 ;
  assign n17053 = \P1_P3_InstQueue_reg[2][4]/NET0131  & n8767 ;
  assign n17062 = ~n17052 & ~n17053 ;
  assign n17054 = \P1_P3_InstQueue_reg[10][4]/NET0131  & n8769 ;
  assign n17055 = \P1_P3_InstQueue_reg[0][4]/NET0131  & n8781 ;
  assign n17063 = ~n17054 & ~n17055 ;
  assign n17064 = n17062 & n17063 ;
  assign n17048 = \P1_P3_InstQueue_reg[5][4]/NET0131  & n8771 ;
  assign n17049 = \P1_P3_InstQueue_reg[12][4]/NET0131  & n8757 ;
  assign n17060 = ~n17048 & ~n17049 ;
  assign n17050 = \P1_P3_InstQueue_reg[15][4]/NET0131  & n8775 ;
  assign n17051 = \P1_P3_InstQueue_reg[1][4]/NET0131  & n8773 ;
  assign n17061 = ~n17050 & ~n17051 ;
  assign n17065 = n17060 & n17061 ;
  assign n17069 = n17064 & n17065 ;
  assign n17070 = n17068 & n17069 ;
  assign n17071 = n16984 & ~n17070 ;
  assign n17072 = ~n17034 & ~n17071 ;
  assign n17073 = ~n17039 & n17072 ;
  assign n17074 = n9241 & ~n17073 ;
  assign n17075 = ~n17032 & ~n17074 ;
  assign n17076 = n9241 & n16987 ;
  assign n17077 = n16968 & ~n17076 ;
  assign n17078 = \P1_P3_EAX_reg[13]/NET0131  & ~n17077 ;
  assign n17081 = ~n9089 & ~n17038 ;
  assign n17082 = \P1_P3_EAX_reg[13]/NET0131  & ~n17081 ;
  assign n17115 = ~\P1_P3_EAX_reg[13]/NET0131  & n16982 ;
  assign n17116 = n17037 & n17115 ;
  assign n17079 = \P1_buf2_reg[13]/NET0131  & n9088 ;
  assign n17080 = ~n9087 & n17079 ;
  assign n17087 = \P1_P3_InstQueue_reg[11][5]/NET0131  & n8763 ;
  assign n17088 = \P1_P3_InstQueue_reg[6][5]/NET0131  & n8745 ;
  assign n17101 = ~n17087 & ~n17088 ;
  assign n17089 = \P1_P3_InstQueue_reg[3][5]/NET0131  & n8777 ;
  assign n17090 = \P1_P3_InstQueue_reg[8][5]/NET0131  & n8754 ;
  assign n17102 = ~n17089 & ~n17090 ;
  assign n17109 = n17101 & n17102 ;
  assign n17083 = \P1_P3_InstQueue_reg[4][5]/NET0131  & n8752 ;
  assign n17084 = \P1_P3_InstQueue_reg[9][5]/NET0131  & n8748 ;
  assign n17099 = ~n17083 & ~n17084 ;
  assign n17085 = \P1_P3_InstQueue_reg[7][5]/NET0131  & n8779 ;
  assign n17086 = \P1_P3_InstQueue_reg[13][5]/NET0131  & n8765 ;
  assign n17100 = ~n17085 & ~n17086 ;
  assign n17110 = n17099 & n17100 ;
  assign n17111 = n17109 & n17110 ;
  assign n17095 = \P1_P3_InstQueue_reg[14][5]/NET0131  & n8760 ;
  assign n17096 = \P1_P3_InstQueue_reg[2][5]/NET0131  & n8767 ;
  assign n17105 = ~n17095 & ~n17096 ;
  assign n17097 = \P1_P3_InstQueue_reg[10][5]/NET0131  & n8769 ;
  assign n17098 = \P1_P3_InstQueue_reg[0][5]/NET0131  & n8781 ;
  assign n17106 = ~n17097 & ~n17098 ;
  assign n17107 = n17105 & n17106 ;
  assign n17091 = \P1_P3_InstQueue_reg[5][5]/NET0131  & n8771 ;
  assign n17092 = \P1_P3_InstQueue_reg[12][5]/NET0131  & n8757 ;
  assign n17103 = ~n17091 & ~n17092 ;
  assign n17093 = \P1_P3_InstQueue_reg[15][5]/NET0131  & n8775 ;
  assign n17094 = \P1_P3_InstQueue_reg[1][5]/NET0131  & n8773 ;
  assign n17104 = ~n17093 & ~n17094 ;
  assign n17108 = n17103 & n17104 ;
  assign n17112 = n17107 & n17108 ;
  assign n17113 = n17111 & n17112 ;
  assign n17114 = n16984 & ~n17113 ;
  assign n17117 = ~n17080 & ~n17114 ;
  assign n17118 = ~n17116 & n17117 ;
  assign n17119 = ~n17082 & n17118 ;
  assign n17120 = n9241 & ~n17119 ;
  assign n17121 = ~n17078 & ~n17120 ;
  assign n17122 = \P1_P3_EAX_reg[10]/NET0131  & ~n16968 ;
  assign n17125 = \P1_P3_EAX_reg[10]/NET0131  & ~n16989 ;
  assign n17130 = \P1_P3_InstQueue_reg[3][2]/NET0131  & n8777 ;
  assign n17131 = \P1_P3_InstQueue_reg[10][2]/NET0131  & n8769 ;
  assign n17144 = ~n17130 & ~n17131 ;
  assign n17132 = \P1_P3_InstQueue_reg[11][2]/NET0131  & n8763 ;
  assign n17133 = \P1_P3_InstQueue_reg[5][2]/NET0131  & n8771 ;
  assign n17145 = ~n17132 & ~n17133 ;
  assign n17152 = n17144 & n17145 ;
  assign n17126 = \P1_P3_InstQueue_reg[6][2]/NET0131  & n8745 ;
  assign n17127 = \P1_P3_InstQueue_reg[9][2]/NET0131  & n8748 ;
  assign n17142 = ~n17126 & ~n17127 ;
  assign n17128 = \P1_P3_InstQueue_reg[14][2]/NET0131  & n8760 ;
  assign n17129 = \P1_P3_InstQueue_reg[13][2]/NET0131  & n8765 ;
  assign n17143 = ~n17128 & ~n17129 ;
  assign n17153 = n17142 & n17143 ;
  assign n17154 = n17152 & n17153 ;
  assign n17138 = \P1_P3_InstQueue_reg[4][2]/NET0131  & n8752 ;
  assign n17139 = \P1_P3_InstQueue_reg[7][2]/NET0131  & n8779 ;
  assign n17148 = ~n17138 & ~n17139 ;
  assign n17140 = \P1_P3_InstQueue_reg[2][2]/NET0131  & n8767 ;
  assign n17141 = \P1_P3_InstQueue_reg[0][2]/NET0131  & n8781 ;
  assign n17149 = ~n17140 & ~n17141 ;
  assign n17150 = n17148 & n17149 ;
  assign n17134 = \P1_P3_InstQueue_reg[8][2]/NET0131  & n8754 ;
  assign n17135 = \P1_P3_InstQueue_reg[12][2]/NET0131  & n8757 ;
  assign n17146 = ~n17134 & ~n17135 ;
  assign n17136 = \P1_P3_InstQueue_reg[15][2]/NET0131  & n8775 ;
  assign n17137 = \P1_P3_InstQueue_reg[1][2]/NET0131  & n8773 ;
  assign n17147 = ~n17136 & ~n17137 ;
  assign n17151 = n17146 & n17147 ;
  assign n17155 = n17150 & n17151 ;
  assign n17156 = n17154 & n17155 ;
  assign n17157 = n16984 & ~n17156 ;
  assign n17123 = \P1_buf2_reg[10]/NET0131  & n9088 ;
  assign n17124 = ~n9087 & n17123 ;
  assign n17158 = n16980 & n16983 ;
  assign n17159 = ~n17124 & ~n17158 ;
  assign n17160 = ~n17157 & n17159 ;
  assign n17161 = ~n17125 & n17160 ;
  assign n17162 = n9241 & ~n17161 ;
  assign n17163 = ~n17122 & ~n17162 ;
  assign n17164 = \P1_P3_EAX_reg[14]/NET0131  & ~n16968 ;
  assign n17165 = \P1_P3_EAX_reg[13]/NET0131  & n17037 ;
  assign n17166 = \P1_P3_EAX_reg[14]/NET0131  & n17165 ;
  assign n17167 = n16982 & ~n17166 ;
  assign n17169 = n16988 & ~n17167 ;
  assign n17170 = \P1_P3_EAX_reg[14]/NET0131  & ~n17169 ;
  assign n17168 = n17165 & n17167 ;
  assign n17175 = \P1_P3_InstQueue_reg[3][6]/NET0131  & n8777 ;
  assign n17176 = \P1_P3_InstQueue_reg[10][6]/NET0131  & n8769 ;
  assign n17189 = ~n17175 & ~n17176 ;
  assign n17177 = \P1_P3_InstQueue_reg[11][6]/NET0131  & n8763 ;
  assign n17178 = \P1_P3_InstQueue_reg[5][6]/NET0131  & n8771 ;
  assign n17190 = ~n17177 & ~n17178 ;
  assign n17197 = n17189 & n17190 ;
  assign n17171 = \P1_P3_InstQueue_reg[6][6]/NET0131  & n8745 ;
  assign n17172 = \P1_P3_InstQueue_reg[9][6]/NET0131  & n8748 ;
  assign n17187 = ~n17171 & ~n17172 ;
  assign n17173 = \P1_P3_InstQueue_reg[14][6]/NET0131  & n8760 ;
  assign n17174 = \P1_P3_InstQueue_reg[13][6]/NET0131  & n8765 ;
  assign n17188 = ~n17173 & ~n17174 ;
  assign n17198 = n17187 & n17188 ;
  assign n17199 = n17197 & n17198 ;
  assign n17183 = \P1_P3_InstQueue_reg[4][6]/NET0131  & n8752 ;
  assign n17184 = \P1_P3_InstQueue_reg[7][6]/NET0131  & n8779 ;
  assign n17193 = ~n17183 & ~n17184 ;
  assign n17185 = \P1_P3_InstQueue_reg[2][6]/NET0131  & n8767 ;
  assign n17186 = \P1_P3_InstQueue_reg[0][6]/NET0131  & n8781 ;
  assign n17194 = ~n17185 & ~n17186 ;
  assign n17195 = n17193 & n17194 ;
  assign n17179 = \P1_P3_InstQueue_reg[8][6]/NET0131  & n8754 ;
  assign n17180 = \P1_P3_InstQueue_reg[12][6]/NET0131  & n8757 ;
  assign n17191 = ~n17179 & ~n17180 ;
  assign n17181 = \P1_P3_InstQueue_reg[15][6]/NET0131  & n8775 ;
  assign n17182 = \P1_P3_InstQueue_reg[1][6]/NET0131  & n8773 ;
  assign n17192 = ~n17181 & ~n17182 ;
  assign n17196 = n17191 & n17192 ;
  assign n17200 = n17195 & n17196 ;
  assign n17201 = n17199 & n17200 ;
  assign n17202 = n16984 & ~n17201 ;
  assign n17203 = \P1_buf2_reg[14]/NET0131  & n9175 ;
  assign n17204 = ~n17202 & ~n17203 ;
  assign n17205 = ~n17168 & n17204 ;
  assign n17206 = ~n17170 & n17205 ;
  assign n17207 = n9241 & ~n17206 ;
  assign n17208 = ~n17164 & ~n17207 ;
  assign n17209 = \P1_P3_EAX_reg[15]/NET0131  & ~n16968 ;
  assign n17211 = \P1_P3_EAX_reg[15]/NET0131  & ~n17169 ;
  assign n17244 = ~\P1_P3_EAX_reg[15]/NET0131  & n16982 ;
  assign n17245 = n17166 & n17244 ;
  assign n17210 = \P1_buf2_reg[15]/NET0131  & n9175 ;
  assign n17216 = \P1_P3_InstQueue_reg[11][7]/NET0131  & n8763 ;
  assign n17217 = \P1_P3_InstQueue_reg[6][7]/NET0131  & n8745 ;
  assign n17230 = ~n17216 & ~n17217 ;
  assign n17218 = \P1_P3_InstQueue_reg[3][7]/NET0131  & n8777 ;
  assign n17219 = \P1_P3_InstQueue_reg[8][7]/NET0131  & n8754 ;
  assign n17231 = ~n17218 & ~n17219 ;
  assign n17238 = n17230 & n17231 ;
  assign n17212 = \P1_P3_InstQueue_reg[4][7]/NET0131  & n8752 ;
  assign n17213 = \P1_P3_InstQueue_reg[9][7]/NET0131  & n8748 ;
  assign n17228 = ~n17212 & ~n17213 ;
  assign n17214 = \P1_P3_InstQueue_reg[7][7]/NET0131  & n8779 ;
  assign n17215 = \P1_P3_InstQueue_reg[13][7]/NET0131  & n8765 ;
  assign n17229 = ~n17214 & ~n17215 ;
  assign n17239 = n17228 & n17229 ;
  assign n17240 = n17238 & n17239 ;
  assign n17224 = \P1_P3_InstQueue_reg[14][7]/NET0131  & n8760 ;
  assign n17225 = \P1_P3_InstQueue_reg[2][7]/NET0131  & n8767 ;
  assign n17234 = ~n17224 & ~n17225 ;
  assign n17226 = \P1_P3_InstQueue_reg[10][7]/NET0131  & n8769 ;
  assign n17227 = \P1_P3_InstQueue_reg[0][7]/NET0131  & n8781 ;
  assign n17235 = ~n17226 & ~n17227 ;
  assign n17236 = n17234 & n17235 ;
  assign n17220 = \P1_P3_InstQueue_reg[5][7]/NET0131  & n8771 ;
  assign n17221 = \P1_P3_InstQueue_reg[12][7]/NET0131  & n8757 ;
  assign n17232 = ~n17220 & ~n17221 ;
  assign n17222 = \P1_P3_InstQueue_reg[15][7]/NET0131  & n8775 ;
  assign n17223 = \P1_P3_InstQueue_reg[1][7]/NET0131  & n8773 ;
  assign n17233 = ~n17222 & ~n17223 ;
  assign n17237 = n17232 & n17233 ;
  assign n17241 = n17236 & n17237 ;
  assign n17242 = n17240 & n17241 ;
  assign n17243 = n16984 & ~n17242 ;
  assign n17246 = ~n17210 & ~n17243 ;
  assign n17247 = ~n17245 & n17246 ;
  assign n17248 = ~n17211 & n17247 ;
  assign n17249 = n9241 & ~n17248 ;
  assign n17250 = ~n17209 & ~n17249 ;
  assign n17251 = \P1_P3_EAX_reg[7]/NET0131  & ~n17031 ;
  assign n17284 = \P1_buf2_reg[7]/NET0131  & n9088 ;
  assign n17285 = ~n9087 & n17284 ;
  assign n17256 = \P1_P3_InstQueue_reg[6][7]/NET0131  & n8779 ;
  assign n17257 = \P1_P3_InstQueue_reg[13][7]/NET0131  & n8760 ;
  assign n17270 = ~n17256 & ~n17257 ;
  assign n17258 = \P1_P3_InstQueue_reg[5][7]/NET0131  & n8745 ;
  assign n17259 = \P1_P3_InstQueue_reg[4][7]/NET0131  & n8771 ;
  assign n17271 = ~n17258 & ~n17259 ;
  assign n17278 = n17270 & n17271 ;
  assign n17252 = \P1_P3_InstQueue_reg[11][7]/NET0131  & n8757 ;
  assign n17253 = \P1_P3_InstQueue_reg[8][7]/NET0131  & n8748 ;
  assign n17268 = ~n17252 & ~n17253 ;
  assign n17254 = \P1_P3_InstQueue_reg[2][7]/NET0131  & n8777 ;
  assign n17255 = \P1_P3_InstQueue_reg[12][7]/NET0131  & n8765 ;
  assign n17269 = ~n17254 & ~n17255 ;
  assign n17279 = n17268 & n17269 ;
  assign n17280 = n17278 & n17279 ;
  assign n17264 = \P1_P3_InstQueue_reg[9][7]/NET0131  & n8769 ;
  assign n17265 = \P1_P3_InstQueue_reg[14][7]/NET0131  & n8775 ;
  assign n17274 = ~n17264 & ~n17265 ;
  assign n17266 = \P1_P3_InstQueue_reg[1][7]/NET0131  & n8767 ;
  assign n17267 = \P1_P3_InstQueue_reg[15][7]/NET0131  & n8781 ;
  assign n17275 = ~n17266 & ~n17267 ;
  assign n17276 = n17274 & n17275 ;
  assign n17260 = \P1_P3_InstQueue_reg[7][7]/NET0131  & n8754 ;
  assign n17261 = \P1_P3_InstQueue_reg[3][7]/NET0131  & n8752 ;
  assign n17272 = ~n17260 & ~n17261 ;
  assign n17262 = \P1_P3_InstQueue_reg[10][7]/NET0131  & n8763 ;
  assign n17263 = \P1_P3_InstQueue_reg[0][7]/NET0131  & n8773 ;
  assign n17273 = ~n17262 & ~n17263 ;
  assign n17277 = n17272 & n17273 ;
  assign n17281 = n17276 & n17277 ;
  assign n17282 = n17280 & n17281 ;
  assign n17283 = n16984 & ~n17282 ;
  assign n17286 = ~\P1_P3_EAX_reg[7]/NET0131  & ~n16977 ;
  assign n17287 = ~n16978 & ~n17286 ;
  assign n17288 = n16982 & n17287 ;
  assign n17289 = ~n17283 & ~n17288 ;
  assign n17290 = ~n17285 & n17289 ;
  assign n17291 = n9241 & ~n17290 ;
  assign n17292 = ~n17251 & ~n17291 ;
  assign n17293 = \P1_P3_EAX_reg[8]/NET0131  & ~n17031 ;
  assign n17300 = \P1_P3_InstQueue_reg[3][0]/NET0131  & n8777 ;
  assign n17301 = \P1_P3_InstQueue_reg[10][0]/NET0131  & n8769 ;
  assign n17314 = ~n17300 & ~n17301 ;
  assign n17302 = \P1_P3_InstQueue_reg[11][0]/NET0131  & n8763 ;
  assign n17303 = \P1_P3_InstQueue_reg[5][0]/NET0131  & n8771 ;
  assign n17315 = ~n17302 & ~n17303 ;
  assign n17322 = n17314 & n17315 ;
  assign n17296 = \P1_P3_InstQueue_reg[6][0]/NET0131  & n8745 ;
  assign n17297 = \P1_P3_InstQueue_reg[9][0]/NET0131  & n8748 ;
  assign n17312 = ~n17296 & ~n17297 ;
  assign n17298 = \P1_P3_InstQueue_reg[14][0]/NET0131  & n8760 ;
  assign n17299 = \P1_P3_InstQueue_reg[13][0]/NET0131  & n8765 ;
  assign n17313 = ~n17298 & ~n17299 ;
  assign n17323 = n17312 & n17313 ;
  assign n17324 = n17322 & n17323 ;
  assign n17308 = \P1_P3_InstQueue_reg[4][0]/NET0131  & n8752 ;
  assign n17309 = \P1_P3_InstQueue_reg[7][0]/NET0131  & n8779 ;
  assign n17318 = ~n17308 & ~n17309 ;
  assign n17310 = \P1_P3_InstQueue_reg[2][0]/NET0131  & n8767 ;
  assign n17311 = \P1_P3_InstQueue_reg[0][0]/NET0131  & n8781 ;
  assign n17319 = ~n17310 & ~n17311 ;
  assign n17320 = n17318 & n17319 ;
  assign n17304 = \P1_P3_InstQueue_reg[8][0]/NET0131  & n8754 ;
  assign n17305 = \P1_P3_InstQueue_reg[12][0]/NET0131  & n8757 ;
  assign n17316 = ~n17304 & ~n17305 ;
  assign n17306 = \P1_P3_InstQueue_reg[15][0]/NET0131  & n8775 ;
  assign n17307 = \P1_P3_InstQueue_reg[1][0]/NET0131  & n8773 ;
  assign n17317 = ~n17306 & ~n17307 ;
  assign n17321 = n17316 & n17317 ;
  assign n17325 = n17320 & n17321 ;
  assign n17326 = n17324 & n17325 ;
  assign n17327 = n16984 & ~n17326 ;
  assign n17294 = \P1_buf2_reg[8]/NET0131  & n9088 ;
  assign n17295 = ~n9087 & n17294 ;
  assign n17328 = ~\P1_P3_EAX_reg[8]/NET0131  & ~n16978 ;
  assign n17329 = ~n16979 & ~n17328 ;
  assign n17330 = n16982 & n17329 ;
  assign n17331 = ~n17295 & ~n17330 ;
  assign n17332 = ~n17327 & n17331 ;
  assign n17333 = n9241 & ~n17332 ;
  assign n17334 = ~n17293 & ~n17333 ;
  assign n17335 = \P1_P3_EAX_reg[9]/NET0131  & ~n17031 ;
  assign n17342 = \P1_P3_InstQueue_reg[11][1]/NET0131  & n8763 ;
  assign n17343 = \P1_P3_InstQueue_reg[6][1]/NET0131  & n8745 ;
  assign n17356 = ~n17342 & ~n17343 ;
  assign n17344 = \P1_P3_InstQueue_reg[3][1]/NET0131  & n8777 ;
  assign n17345 = \P1_P3_InstQueue_reg[8][1]/NET0131  & n8754 ;
  assign n17357 = ~n17344 & ~n17345 ;
  assign n17364 = n17356 & n17357 ;
  assign n17338 = \P1_P3_InstQueue_reg[4][1]/NET0131  & n8752 ;
  assign n17339 = \P1_P3_InstQueue_reg[9][1]/NET0131  & n8748 ;
  assign n17354 = ~n17338 & ~n17339 ;
  assign n17340 = \P1_P3_InstQueue_reg[7][1]/NET0131  & n8779 ;
  assign n17341 = \P1_P3_InstQueue_reg[13][1]/NET0131  & n8765 ;
  assign n17355 = ~n17340 & ~n17341 ;
  assign n17365 = n17354 & n17355 ;
  assign n17366 = n17364 & n17365 ;
  assign n17350 = \P1_P3_InstQueue_reg[14][1]/NET0131  & n8760 ;
  assign n17351 = \P1_P3_InstQueue_reg[2][1]/NET0131  & n8767 ;
  assign n17360 = ~n17350 & ~n17351 ;
  assign n17352 = \P1_P3_InstQueue_reg[10][1]/NET0131  & n8769 ;
  assign n17353 = \P1_P3_InstQueue_reg[0][1]/NET0131  & n8781 ;
  assign n17361 = ~n17352 & ~n17353 ;
  assign n17362 = n17360 & n17361 ;
  assign n17346 = \P1_P3_InstQueue_reg[5][1]/NET0131  & n8771 ;
  assign n17347 = \P1_P3_InstQueue_reg[12][1]/NET0131  & n8757 ;
  assign n17358 = ~n17346 & ~n17347 ;
  assign n17348 = \P1_P3_InstQueue_reg[15][1]/NET0131  & n8775 ;
  assign n17349 = \P1_P3_InstQueue_reg[1][1]/NET0131  & n8773 ;
  assign n17359 = ~n17348 & ~n17349 ;
  assign n17363 = n17358 & n17359 ;
  assign n17367 = n17362 & n17363 ;
  assign n17368 = n17366 & n17367 ;
  assign n17369 = n16984 & ~n17368 ;
  assign n17336 = \P1_buf2_reg[9]/NET0131  & n9088 ;
  assign n17337 = ~n9087 & n17336 ;
  assign n17370 = ~\P1_P3_EAX_reg[9]/NET0131  & ~n16979 ;
  assign n17371 = ~n16980 & ~n17370 ;
  assign n17372 = n16982 & n17371 ;
  assign n17373 = ~n17337 & ~n17372 ;
  assign n17374 = ~n17369 & n17373 ;
  assign n17375 = n9241 & ~n17374 ;
  assign n17376 = ~n17335 & ~n17375 ;
  assign n17380 = ~n11346 & ~n11578 ;
  assign n17381 = ~n11579 & ~n17380 ;
  assign n17382 = ~n10105 & ~n17381 ;
  assign n17377 = ~n11412 & ~n11463 ;
  assign n17378 = ~n11464 & ~n17377 ;
  assign n17379 = n10105 & ~n17378 ;
  assign n17383 = n12334 & ~n17379 ;
  assign n17384 = ~n17382 & n17383 ;
  assign n17392 = \P2_P1_InstQueue_reg[6][0]/NET0131  & n11651 ;
  assign n17391 = \P2_P1_InstQueue_reg[15][0]/NET0131  & n11647 ;
  assign n17387 = \P2_P1_InstQueue_reg[11][0]/NET0131  & n11665 ;
  assign n17388 = \P2_P1_InstQueue_reg[10][0]/NET0131  & n11634 ;
  assign n17403 = ~n17387 & ~n17388 ;
  assign n17413 = ~n17391 & n17403 ;
  assign n17414 = ~n17392 & n17413 ;
  assign n17399 = \P2_P1_InstQueue_reg[0][0]/NET0131  & n11669 ;
  assign n17400 = \P2_P1_InstQueue_reg[9][0]/NET0131  & n11656 ;
  assign n17408 = ~n17399 & ~n17400 ;
  assign n17401 = \P2_P1_InstQueue_reg[2][0]/NET0131  & n11654 ;
  assign n17402 = \P2_P1_InstQueue_reg[4][0]/NET0131  & n11667 ;
  assign n17409 = ~n17401 & ~n17402 ;
  assign n17410 = n17408 & n17409 ;
  assign n17395 = \P2_P1_InstQueue_reg[12][0]/NET0131  & n11673 ;
  assign n17396 = \P2_P1_InstQueue_reg[7][0]/NET0131  & n11661 ;
  assign n17406 = ~n17395 & ~n17396 ;
  assign n17397 = \P2_P1_InstQueue_reg[1][0]/NET0131  & n11671 ;
  assign n17398 = \P2_P1_InstQueue_reg[5][0]/NET0131  & n11638 ;
  assign n17407 = ~n17397 & ~n17398 ;
  assign n17411 = n17406 & n17407 ;
  assign n17389 = \P2_P1_InstQueue_reg[8][0]/NET0131  & n11659 ;
  assign n17390 = \P2_P1_InstQueue_reg[14][0]/NET0131  & n11643 ;
  assign n17404 = ~n17389 & ~n17390 ;
  assign n17393 = \P2_P1_InstQueue_reg[13][0]/NET0131  & n11641 ;
  assign n17394 = \P2_P1_InstQueue_reg[3][0]/NET0131  & n11663 ;
  assign n17405 = ~n17393 & ~n17394 ;
  assign n17412 = n17404 & n17405 ;
  assign n17415 = n17411 & n17412 ;
  assign n17416 = n17410 & n17415 ;
  assign n17417 = n17414 & n17416 ;
  assign n17418 = n11596 & n17417 ;
  assign n17386 = ~\P2_P1_InstQueue_reg[11][0]/NET0131  & ~n11596 ;
  assign n17419 = n11692 & ~n17386 ;
  assign n17420 = ~n17418 & n17419 ;
  assign n17385 = \P2_P1_InstQueue_reg[11][0]/NET0131  & ~n12345 ;
  assign n17421 = n11379 & ~n11600 ;
  assign n17422 = n12343 & n17421 ;
  assign n17423 = ~n17385 & ~n17422 ;
  assign n17424 = ~n17420 & n17423 ;
  assign n17425 = ~n17384 & n17424 ;
  assign n17428 = ~\P1_P3_PhyAddrPointer_reg[15]/NET0131  & ~n16534 ;
  assign n17429 = ~n16535 & ~n17428 ;
  assign n17430 = ~\P1_P3_PhyAddrPointer_reg[0]/NET0131  & n16534 ;
  assign n17431 = n16484 & ~n17430 ;
  assign n17433 = n17429 & ~n17431 ;
  assign n17432 = ~n17429 & n17431 ;
  assign n17434 = ~\P1_P3_DataWidth_reg[1]/NET0131  & ~n17432 ;
  assign n17435 = ~n17433 & n17434 ;
  assign n17427 = \P1_P3_DataWidth_reg[1]/NET0131  & ~\P1_P3_rEIP_reg[15]/NET0131  ;
  assign n17436 = n9245 & ~n17427 ;
  assign n17437 = ~n17435 & n17436 ;
  assign n17438 = \P1_P3_rEIP_reg[15]/NET0131  & ~n9195 ;
  assign n17440 = ~\P1_P3_rEIP_reg[15]/NET0131  & ~n16580 ;
  assign n17441 = ~n16581 & ~n17440 ;
  assign n17442 = n16505 & ~n17441 ;
  assign n17443 = ~n9095 & n17442 ;
  assign n17439 = ~\P1_P3_EBX_reg[15]/NET0131  & ~n16517 ;
  assign n17444 = n9079 & ~n17439 ;
  assign n17445 = ~n17443 & n17444 ;
  assign n17446 = \P1_P3_EBX_reg[31]/NET0131  & ~n16607 ;
  assign n17448 = ~\P1_P3_EBX_reg[15]/NET0131  & n17446 ;
  assign n17447 = \P1_P3_EBX_reg[15]/NET0131  & ~n17446 ;
  assign n17449 = ~n16505 & ~n17447 ;
  assign n17450 = ~n17448 & n17449 ;
  assign n17451 = n9085 & ~n17442 ;
  assign n17452 = ~n17450 & n17451 ;
  assign n17453 = ~n17445 & ~n17452 ;
  assign n17454 = ~n9075 & ~n17453 ;
  assign n17455 = ~n17438 & ~n17454 ;
  assign n17456 = n9241 & ~n17455 ;
  assign n17458 = n8735 & n10047 ;
  assign n17459 = \P1_P3_rEIP_reg[15]/NET0131  & ~n17458 ;
  assign n17426 = n8733 & n10029 ;
  assign n17457 = \P1_P3_PhyAddrPointer_reg[15]/NET0131  & n10031 ;
  assign n17460 = ~n17426 & ~n17457 ;
  assign n17461 = ~n17459 & n17460 ;
  assign n17462 = ~n17456 & n17461 ;
  assign n17463 = ~n17437 & n17462 ;
  assign n17466 = n16484 & ~n16550 ;
  assign n17468 = ~n16546 & n17466 ;
  assign n17467 = n16546 & ~n17466 ;
  assign n17469 = ~\P1_P3_DataWidth_reg[1]/NET0131  & ~n17467 ;
  assign n17470 = ~n17468 & n17469 ;
  assign n17465 = \P1_P3_DataWidth_reg[1]/NET0131  & ~\P1_P3_rEIP_reg[17]/NET0131  ;
  assign n17471 = n9245 & ~n17465 ;
  assign n17472 = ~n17470 & n17471 ;
  assign n17473 = \P1_P3_rEIP_reg[17]/NET0131  & ~n9195 ;
  assign n17474 = ~\P1_P3_EBX_reg[17]/NET0131  & ~n16517 ;
  assign n17475 = n9079 & ~n17474 ;
  assign n17476 = \P1_P3_EBX_reg[31]/NET0131  & ~n16609 ;
  assign n17478 = ~\P1_P3_EBX_reg[17]/NET0131  & n17476 ;
  assign n17477 = \P1_P3_EBX_reg[17]/NET0131  & ~n17476 ;
  assign n17479 = ~n16505 & ~n17477 ;
  assign n17480 = ~n17478 & n17479 ;
  assign n17481 = n9085 & ~n17480 ;
  assign n17482 = ~n17475 & ~n17481 ;
  assign n17484 = ~\P1_P3_rEIP_reg[17]/NET0131  & ~n16582 ;
  assign n17485 = ~n16583 & ~n17484 ;
  assign n17483 = n9095 & n17475 ;
  assign n17486 = n16505 & ~n17483 ;
  assign n17487 = ~n17485 & n17486 ;
  assign n17488 = ~n9075 & ~n17487 ;
  assign n17489 = ~n17482 & n17488 ;
  assign n17490 = ~n17473 & ~n17489 ;
  assign n17491 = n9241 & ~n17490 ;
  assign n17464 = \P1_P3_rEIP_reg[17]/NET0131  & ~n17458 ;
  assign n17492 = \P1_P3_PhyAddrPointer_reg[17]/NET0131  & n10031 ;
  assign n17493 = ~n17426 & ~n17492 ;
  assign n17494 = ~n17464 & n17493 ;
  assign n17495 = ~n17491 & n17494 ;
  assign n17496 = ~n17472 & n17495 ;
  assign n17499 = n16484 & ~n16551 ;
  assign n17501 = ~n16553 & n17499 ;
  assign n17500 = n16553 & ~n17499 ;
  assign n17502 = ~\P1_P3_DataWidth_reg[1]/NET0131  & ~n17500 ;
  assign n17503 = ~n17501 & n17502 ;
  assign n17498 = \P1_P3_DataWidth_reg[1]/NET0131  & ~\P1_P3_rEIP_reg[18]/NET0131  ;
  assign n17504 = n9245 & ~n17498 ;
  assign n17505 = ~n17503 & n17504 ;
  assign n17506 = \P1_P3_rEIP_reg[18]/NET0131  & ~n9195 ;
  assign n17507 = ~\P1_P3_EBX_reg[18]/NET0131  & ~n16517 ;
  assign n17508 = n9079 & ~n17507 ;
  assign n17509 = \P1_P3_EBX_reg[31]/NET0131  & ~n16610 ;
  assign n17511 = ~\P1_P3_EBX_reg[18]/NET0131  & n17509 ;
  assign n17510 = \P1_P3_EBX_reg[18]/NET0131  & ~n17509 ;
  assign n17512 = ~n16505 & ~n17510 ;
  assign n17513 = ~n17511 & n17512 ;
  assign n17514 = n9085 & ~n17513 ;
  assign n17515 = ~n17508 & ~n17514 ;
  assign n17517 = ~\P1_P3_rEIP_reg[18]/NET0131  & ~n16583 ;
  assign n17518 = ~n16584 & ~n17517 ;
  assign n17516 = n9095 & n17508 ;
  assign n17519 = n16505 & ~n17516 ;
  assign n17520 = ~n17518 & n17519 ;
  assign n17521 = ~n9075 & ~n17520 ;
  assign n17522 = ~n17515 & n17521 ;
  assign n17523 = ~n17506 & ~n17522 ;
  assign n17524 = n9241 & ~n17523 ;
  assign n17497 = \P1_P3_rEIP_reg[18]/NET0131  & ~n17458 ;
  assign n17525 = \P1_P3_PhyAddrPointer_reg[18]/NET0131  & n10031 ;
  assign n17526 = ~n17426 & ~n17525 ;
  assign n17527 = ~n17497 & n17526 ;
  assign n17528 = ~n17524 & n17527 ;
  assign n17529 = ~n17505 & n17528 ;
  assign n17532 = ~\P1_P3_PhyAddrPointer_reg[4]/NET0131  & ~n16450 ;
  assign n17533 = \P1_P3_PhyAddrPointer_reg[1]/NET0131  & n16454 ;
  assign n17534 = ~n17532 & ~n17533 ;
  assign n17535 = \P1_P3_PhyAddrPointer_reg[3]/NET0131  & n16452 ;
  assign n17536 = n16484 & ~n17535 ;
  assign n17537 = ~n17534 & ~n17536 ;
  assign n17538 = n17534 & n17536 ;
  assign n17539 = ~n17537 & ~n17538 ;
  assign n17540 = ~\P1_P3_DataWidth_reg[1]/NET0131  & ~n17539 ;
  assign n17531 = \P1_P3_DataWidth_reg[1]/NET0131  & ~\P1_P3_rEIP_reg[4]/NET0131  ;
  assign n17541 = n9245 & ~n17531 ;
  assign n17542 = ~n17540 & n17541 ;
  assign n17549 = \P1_P3_rEIP_reg[4]/NET0131  & ~n9195 ;
  assign n17543 = ~\P1_P3_EBX_reg[4]/NET0131  & ~n16517 ;
  assign n17544 = ~\P1_P3_rEIP_reg[4]/NET0131  & ~n16510 ;
  assign n17545 = ~n16570 & ~n17544 ;
  assign n17546 = n16517 & ~n17545 ;
  assign n17547 = ~n17543 & ~n17546 ;
  assign n17548 = n9236 & n17547 ;
  assign n17550 = \P1_P3_EBX_reg[31]/NET0131  & ~n16596 ;
  assign n17552 = ~\P1_P3_EBX_reg[4]/NET0131  & n17550 ;
  assign n17551 = \P1_P3_EBX_reg[4]/NET0131  & ~n17550 ;
  assign n17553 = ~n16505 & ~n17551 ;
  assign n17554 = ~n17552 & n17553 ;
  assign n17555 = n16505 & ~n17545 ;
  assign n17556 = ~n17554 & ~n17555 ;
  assign n17557 = n16500 & n17556 ;
  assign n17558 = ~n17548 & ~n17557 ;
  assign n17559 = ~n17549 & n17558 ;
  assign n17560 = n9241 & ~n17559 ;
  assign n17530 = \P1_P3_rEIP_reg[4]/NET0131  & ~n17458 ;
  assign n17561 = \P1_P3_PhyAddrPointer_reg[4]/NET0131  & n10031 ;
  assign n17562 = ~n17426 & ~n17561 ;
  assign n17563 = ~n17530 & n17562 ;
  assign n17564 = ~n17560 & n17563 ;
  assign n17565 = ~n17542 & n17564 ;
  assign n17568 = \P1_P3_PhyAddrPointer_reg[5]/NET0131  & n17533 ;
  assign n17569 = ~\P1_P3_PhyAddrPointer_reg[6]/NET0131  & ~n17568 ;
  assign n17570 = \P1_P3_PhyAddrPointer_reg[6]/NET0131  & n17568 ;
  assign n17571 = ~n17569 & ~n17570 ;
  assign n17572 = ~\P1_P3_PhyAddrPointer_reg[0]/NET0131  & n17568 ;
  assign n17573 = n16484 & ~n17572 ;
  assign n17575 = ~n17571 & n17573 ;
  assign n17574 = n17571 & ~n17573 ;
  assign n17576 = ~\P1_P3_DataWidth_reg[1]/NET0131  & ~n17574 ;
  assign n17577 = ~n17575 & n17576 ;
  assign n17567 = \P1_P3_DataWidth_reg[1]/NET0131  & ~\P1_P3_rEIP_reg[6]/NET0131  ;
  assign n17578 = n9245 & ~n17567 ;
  assign n17579 = ~n17577 & n17578 ;
  assign n17580 = \P1_P3_rEIP_reg[6]/NET0131  & ~n9195 ;
  assign n17581 = ~\P1_P3_EBX_reg[6]/NET0131  & ~n16517 ;
  assign n17582 = ~\P1_P3_rEIP_reg[6]/NET0131  & ~n16571 ;
  assign n17583 = ~n16572 & ~n17582 ;
  assign n17584 = n16517 & ~n17583 ;
  assign n17585 = ~n17581 & ~n17584 ;
  assign n17586 = n9236 & n17585 ;
  assign n17587 = n16505 & ~n17583 ;
  assign n17588 = \P1_P3_EBX_reg[31]/NET0131  & ~n16598 ;
  assign n17590 = ~\P1_P3_EBX_reg[6]/NET0131  & n17588 ;
  assign n17589 = \P1_P3_EBX_reg[6]/NET0131  & ~n17588 ;
  assign n17591 = ~n16505 & ~n17589 ;
  assign n17592 = ~n17590 & n17591 ;
  assign n17593 = ~n17587 & ~n17592 ;
  assign n17594 = n16500 & n17593 ;
  assign n17595 = ~n17586 & ~n17594 ;
  assign n17596 = ~n17580 & n17595 ;
  assign n17597 = n9241 & ~n17596 ;
  assign n17566 = \P1_P3_rEIP_reg[6]/NET0131  & ~n17458 ;
  assign n17598 = \P1_P3_PhyAddrPointer_reg[6]/NET0131  & n10031 ;
  assign n17599 = ~n17426 & ~n17598 ;
  assign n17600 = ~n17566 & n17599 ;
  assign n17601 = ~n17597 & n17600 ;
  assign n17602 = ~n17579 & n17601 ;
  assign n17605 = ~\P1_P3_PhyAddrPointer_reg[7]/NET0131  & ~n17570 ;
  assign n17606 = \P1_P3_PhyAddrPointer_reg[7]/NET0131  & n17570 ;
  assign n17607 = ~n17605 & ~n17606 ;
  assign n17608 = ~\P1_P3_PhyAddrPointer_reg[0]/NET0131  & n17570 ;
  assign n17609 = n16484 & ~n17608 ;
  assign n17611 = ~n17607 & n17609 ;
  assign n17610 = n17607 & ~n17609 ;
  assign n17612 = ~\P1_P3_DataWidth_reg[1]/NET0131  & ~n17610 ;
  assign n17613 = ~n17611 & n17612 ;
  assign n17604 = \P1_P3_DataWidth_reg[1]/NET0131  & ~\P1_P3_rEIP_reg[7]/NET0131  ;
  assign n17614 = n9245 & ~n17604 ;
  assign n17615 = ~n17613 & n17614 ;
  assign n17616 = \P1_P3_rEIP_reg[7]/NET0131  & ~n9195 ;
  assign n17617 = ~\P1_P3_EBX_reg[7]/NET0131  & ~n16517 ;
  assign n17618 = ~\P1_P3_rEIP_reg[7]/NET0131  & ~n16572 ;
  assign n17619 = ~n16573 & ~n17618 ;
  assign n17620 = n16517 & ~n17619 ;
  assign n17621 = ~n17617 & ~n17620 ;
  assign n17622 = n9236 & n17621 ;
  assign n17623 = n16505 & ~n17619 ;
  assign n17624 = \P1_P3_EBX_reg[31]/NET0131  & ~n16599 ;
  assign n17626 = ~\P1_P3_EBX_reg[7]/NET0131  & n17624 ;
  assign n17625 = \P1_P3_EBX_reg[7]/NET0131  & ~n17624 ;
  assign n17627 = ~n16505 & ~n17625 ;
  assign n17628 = ~n17626 & n17627 ;
  assign n17629 = ~n17623 & ~n17628 ;
  assign n17630 = n16500 & n17629 ;
  assign n17631 = ~n17622 & ~n17630 ;
  assign n17632 = ~n17616 & n17631 ;
  assign n17633 = n9241 & ~n17632 ;
  assign n17603 = \P1_P3_rEIP_reg[7]/NET0131  & ~n17458 ;
  assign n17634 = \P1_P3_PhyAddrPointer_reg[7]/NET0131  & n10031 ;
  assign n17635 = ~n17426 & ~n17634 ;
  assign n17636 = ~n17603 & n17635 ;
  assign n17637 = ~n17633 & n17636 ;
  assign n17638 = ~n17615 & n17637 ;
  assign n17661 = \P1_P3_PhyAddrPointer_reg[1]/NET0131  & n16458 ;
  assign n17662 = \P1_P3_PhyAddrPointer_reg[9]/NET0131  & n17661 ;
  assign n17663 = ~\P1_P3_PhyAddrPointer_reg[10]/NET0131  & ~n17662 ;
  assign n17664 = \P1_P3_PhyAddrPointer_reg[10]/NET0131  & n17662 ;
  assign n17665 = ~n17663 & ~n17664 ;
  assign n17666 = \P1_P3_PhyAddrPointer_reg[7]/NET0131  & n17608 ;
  assign n17667 = n16459 & n17666 ;
  assign n17668 = n16484 & ~n17667 ;
  assign n17669 = ~n17665 & ~n17668 ;
  assign n17670 = n17665 & n17668 ;
  assign n17671 = ~n17669 & ~n17670 ;
  assign n17672 = ~\P1_P3_DataWidth_reg[1]/NET0131  & ~n17671 ;
  assign n17660 = \P1_P3_DataWidth_reg[1]/NET0131  & ~\P1_P3_rEIP_reg[10]/NET0131  ;
  assign n17673 = n9245 & ~n17660 ;
  assign n17674 = ~n17672 & n17673 ;
  assign n17640 = \P1_P3_rEIP_reg[10]/NET0131  & ~n9195 ;
  assign n17642 = ~\P1_P3_rEIP_reg[10]/NET0131  & ~n16575 ;
  assign n17643 = ~n16576 & ~n17642 ;
  assign n17644 = n16517 & ~n17643 ;
  assign n17641 = ~\P1_P3_EBX_reg[10]/NET0131  & ~n16517 ;
  assign n17645 = n9079 & ~n17641 ;
  assign n17646 = ~n17644 & n17645 ;
  assign n17648 = \P1_P3_EBX_reg[31]/NET0131  & ~n16602 ;
  assign n17650 = ~\P1_P3_EBX_reg[10]/NET0131  & n17648 ;
  assign n17649 = \P1_P3_EBX_reg[10]/NET0131  & ~n17648 ;
  assign n17651 = ~n16505 & ~n17649 ;
  assign n17652 = ~n17650 & n17651 ;
  assign n17647 = n16505 & ~n17643 ;
  assign n17653 = n9085 & ~n17647 ;
  assign n17654 = ~n17652 & n17653 ;
  assign n17655 = ~n17646 & ~n17654 ;
  assign n17656 = ~n9075 & ~n17655 ;
  assign n17657 = ~n17640 & ~n17656 ;
  assign n17658 = n9241 & ~n17657 ;
  assign n17639 = \P1_P3_rEIP_reg[10]/NET0131  & ~n17458 ;
  assign n17659 = \P1_P3_PhyAddrPointer_reg[10]/NET0131  & n10031 ;
  assign n17675 = ~n17426 & ~n17659 ;
  assign n17676 = ~n17639 & n17675 ;
  assign n17677 = ~n17658 & n17676 ;
  assign n17678 = ~n17674 & n17677 ;
  assign n17680 = ~\P1_P3_PhyAddrPointer_reg[11]/NET0131  & ~n17664 ;
  assign n17681 = ~n16531 & ~n17680 ;
  assign n17682 = ~n17665 & n17667 ;
  assign n17683 = n16484 & ~n17682 ;
  assign n17684 = ~n17681 & ~n17683 ;
  assign n17685 = n17681 & n17683 ;
  assign n17686 = ~n17684 & ~n17685 ;
  assign n17687 = ~\P1_P3_DataWidth_reg[1]/NET0131  & ~n17686 ;
  assign n17688 = \P1_P3_DataWidth_reg[1]/NET0131  & ~\P1_P3_rEIP_reg[11]/NET0131  ;
  assign n17689 = n9245 & ~n17688 ;
  assign n17690 = ~n17687 & n17689 ;
  assign n17691 = \P1_P3_rEIP_reg[11]/NET0131  & ~n9195 ;
  assign n17692 = \P1_P3_EBX_reg[31]/NET0131  & ~n16603 ;
  assign n17694 = \P1_P3_EBX_reg[11]/NET0131  & n17692 ;
  assign n17693 = ~\P1_P3_EBX_reg[11]/NET0131  & ~n17692 ;
  assign n17695 = ~n16505 & ~n17693 ;
  assign n17696 = ~n17694 & n17695 ;
  assign n17697 = ~\P1_P3_rEIP_reg[11]/NET0131  & ~n16576 ;
  assign n17698 = ~n16577 & ~n17697 ;
  assign n17699 = ~\P1_P3_DataWidth_reg[1]/NET0131  & n17698 ;
  assign n17700 = ~n8741 & n17699 ;
  assign n17701 = ~n17696 & ~n17700 ;
  assign n17702 = n9085 & ~n17701 ;
  assign n17703 = \P1_P3_EBX_reg[11]/NET0131  & ~n16517 ;
  assign n17704 = n9096 & n17699 ;
  assign n17705 = ~n17703 & ~n17704 ;
  assign n17706 = n9079 & ~n17705 ;
  assign n17707 = ~n17702 & ~n17706 ;
  assign n17708 = ~n9075 & ~n17707 ;
  assign n17709 = ~n17691 & ~n17708 ;
  assign n17710 = n9241 & ~n17709 ;
  assign n17679 = \P1_P3_rEIP_reg[11]/NET0131  & ~n17458 ;
  assign n17711 = \P1_P3_PhyAddrPointer_reg[11]/NET0131  & n10031 ;
  assign n17712 = ~n17426 & ~n17711 ;
  assign n17713 = ~n17679 & n17712 ;
  assign n17714 = ~n17710 & n17713 ;
  assign n17715 = ~n17690 & n17714 ;
  assign n17718 = ~\P1_P3_PhyAddrPointer_reg[12]/NET0131  & ~n16531 ;
  assign n17719 = ~n16532 & ~n17718 ;
  assign n17720 = n16484 & ~n17684 ;
  assign n17722 = n17719 & ~n17720 ;
  assign n17721 = ~n17719 & n17720 ;
  assign n17723 = ~\P1_P3_DataWidth_reg[1]/NET0131  & ~n17721 ;
  assign n17724 = ~n17722 & n17723 ;
  assign n17717 = \P1_P3_DataWidth_reg[1]/NET0131  & ~\P1_P3_rEIP_reg[12]/NET0131  ;
  assign n17725 = n9245 & ~n17717 ;
  assign n17726 = ~n17724 & n17725 ;
  assign n17727 = \P1_P3_rEIP_reg[12]/NET0131  & ~n9195 ;
  assign n17729 = ~\P1_P3_rEIP_reg[12]/NET0131  & ~n16577 ;
  assign n17730 = ~n16578 & ~n17729 ;
  assign n17731 = n16505 & ~n17730 ;
  assign n17732 = ~n9095 & n17731 ;
  assign n17728 = ~\P1_P3_EBX_reg[12]/NET0131  & ~n16517 ;
  assign n17733 = n9079 & ~n17728 ;
  assign n17734 = ~n17732 & n17733 ;
  assign n17735 = \P1_P3_EBX_reg[31]/NET0131  & ~n16604 ;
  assign n17737 = ~\P1_P3_EBX_reg[12]/NET0131  & n17735 ;
  assign n17736 = \P1_P3_EBX_reg[12]/NET0131  & ~n17735 ;
  assign n17738 = ~n16505 & ~n17736 ;
  assign n17739 = ~n17737 & n17738 ;
  assign n17740 = n9085 & ~n17731 ;
  assign n17741 = ~n17739 & n17740 ;
  assign n17742 = ~n17734 & ~n17741 ;
  assign n17743 = ~n9075 & ~n17742 ;
  assign n17744 = ~n17727 & ~n17743 ;
  assign n17745 = n9241 & ~n17744 ;
  assign n17716 = \P1_P3_rEIP_reg[12]/NET0131  & ~n17458 ;
  assign n17746 = \P1_P3_PhyAddrPointer_reg[12]/NET0131  & n10031 ;
  assign n17747 = ~n17426 & ~n17746 ;
  assign n17748 = ~n17716 & n17747 ;
  assign n17749 = ~n17745 & n17748 ;
  assign n17750 = ~n17726 & n17749 ;
  assign n17753 = ~\P1_P3_PhyAddrPointer_reg[13]/NET0131  & ~n16532 ;
  assign n17754 = ~n16533 & ~n17753 ;
  assign n17755 = n16484 & ~n16547 ;
  assign n17757 = n17754 & ~n17755 ;
  assign n17756 = ~n17754 & n17755 ;
  assign n17758 = ~\P1_P3_DataWidth_reg[1]/NET0131  & ~n17756 ;
  assign n17759 = ~n17757 & n17758 ;
  assign n17752 = \P1_P3_DataWidth_reg[1]/NET0131  & ~\P1_P3_rEIP_reg[13]/NET0131  ;
  assign n17760 = n9245 & ~n17752 ;
  assign n17761 = ~n17759 & n17760 ;
  assign n17774 = \P1_P3_EBX_reg[31]/NET0131  & ~n16605 ;
  assign n17776 = ~\P1_P3_EBX_reg[13]/NET0131  & n17774 ;
  assign n17775 = \P1_P3_EBX_reg[13]/NET0131  & ~n17774 ;
  assign n17777 = ~n16505 & ~n17775 ;
  assign n17778 = ~n17776 & n17777 ;
  assign n17765 = ~\P1_P3_rEIP_reg[13]/NET0131  & ~n16578 ;
  assign n17766 = ~n16579 & ~n17765 ;
  assign n17767 = n16505 & ~n17766 ;
  assign n17779 = n16500 & ~n17767 ;
  assign n17780 = ~n17778 & n17779 ;
  assign n17762 = \P1_P3_rEIP_reg[13]/NET0131  & ~n16565 ;
  assign n17768 = ~\P1_P3_EBX_reg[13]/NET0131  & ~n16505 ;
  assign n17769 = n9162 & ~n17768 ;
  assign n17770 = ~n17767 & n17769 ;
  assign n17763 = \P1_P3_rEIP_reg[13]/NET0131  & n9075 ;
  assign n17764 = \P1_P3_EBX_reg[13]/NET0131  & n16567 ;
  assign n17771 = ~n17763 & ~n17764 ;
  assign n17772 = ~n17770 & n17771 ;
  assign n17773 = n9079 & ~n17772 ;
  assign n17781 = ~n17762 & ~n17773 ;
  assign n17782 = ~n17780 & n17781 ;
  assign n17783 = n9241 & ~n17782 ;
  assign n17751 = \P1_P3_rEIP_reg[13]/NET0131  & ~n17458 ;
  assign n17784 = \P1_P3_PhyAddrPointer_reg[13]/NET0131  & n10031 ;
  assign n17785 = ~n17426 & ~n17784 ;
  assign n17786 = ~n17751 & n17785 ;
  assign n17787 = ~n17783 & n17786 ;
  assign n17788 = ~n17761 & n17787 ;
  assign n17791 = n16484 & ~n16548 ;
  assign n17792 = ~\P1_P3_PhyAddrPointer_reg[14]/NET0131  & ~n16533 ;
  assign n17793 = ~n16534 & ~n17792 ;
  assign n17795 = ~n17791 & n17793 ;
  assign n17794 = n17791 & ~n17793 ;
  assign n17796 = ~\P1_P3_DataWidth_reg[1]/NET0131  & ~n17794 ;
  assign n17797 = ~n17795 & n17796 ;
  assign n17790 = \P1_P3_DataWidth_reg[1]/NET0131  & ~\P1_P3_rEIP_reg[14]/NET0131  ;
  assign n17798 = n9245 & ~n17790 ;
  assign n17799 = ~n17797 & n17798 ;
  assign n17812 = \P1_P3_EBX_reg[31]/NET0131  & ~n16606 ;
  assign n17814 = ~\P1_P3_EBX_reg[14]/NET0131  & n17812 ;
  assign n17813 = \P1_P3_EBX_reg[14]/NET0131  & ~n17812 ;
  assign n17815 = ~n16505 & ~n17813 ;
  assign n17816 = ~n17814 & n17815 ;
  assign n17803 = ~\P1_P3_rEIP_reg[14]/NET0131  & ~n16579 ;
  assign n17804 = ~n16580 & ~n17803 ;
  assign n17805 = n16505 & ~n17804 ;
  assign n17817 = n16500 & ~n17805 ;
  assign n17818 = ~n17816 & n17817 ;
  assign n17800 = \P1_P3_rEIP_reg[14]/NET0131  & ~n16565 ;
  assign n17806 = ~\P1_P3_EBX_reg[14]/NET0131  & ~n16505 ;
  assign n17807 = n9162 & ~n17806 ;
  assign n17808 = ~n17805 & n17807 ;
  assign n17801 = \P1_P3_rEIP_reg[14]/NET0131  & n9075 ;
  assign n17802 = \P1_P3_EBX_reg[14]/NET0131  & n16567 ;
  assign n17809 = ~n17801 & ~n17802 ;
  assign n17810 = ~n17808 & n17809 ;
  assign n17811 = n9079 & ~n17810 ;
  assign n17819 = ~n17800 & ~n17811 ;
  assign n17820 = ~n17818 & n17819 ;
  assign n17821 = n9241 & ~n17820 ;
  assign n17789 = \P1_P3_rEIP_reg[14]/NET0131  & ~n17458 ;
  assign n17822 = \P1_P3_PhyAddrPointer_reg[14]/NET0131  & n10031 ;
  assign n17823 = ~n17426 & ~n17822 ;
  assign n17824 = ~n17789 & n17823 ;
  assign n17825 = ~n17821 & n17824 ;
  assign n17826 = ~n17799 & n17825 ;
  assign n17829 = ~\P1_P3_PhyAddrPointer_reg[16]/NET0131  & ~n16535 ;
  assign n17830 = ~n16536 & ~n17829 ;
  assign n17831 = n16484 & ~n16549 ;
  assign n17833 = n17830 & ~n17831 ;
  assign n17832 = ~n17830 & n17831 ;
  assign n17834 = ~\P1_P3_DataWidth_reg[1]/NET0131  & ~n17832 ;
  assign n17835 = ~n17833 & n17834 ;
  assign n17828 = \P1_P3_DataWidth_reg[1]/NET0131  & ~\P1_P3_rEIP_reg[16]/NET0131  ;
  assign n17836 = n9245 & ~n17828 ;
  assign n17837 = ~n17835 & n17836 ;
  assign n17841 = \P1_P3_EBX_reg[31]/NET0131  & ~n16608 ;
  assign n17843 = ~\P1_P3_EBX_reg[16]/NET0131  & n17841 ;
  assign n17842 = \P1_P3_EBX_reg[16]/NET0131  & ~n17841 ;
  assign n17844 = ~n16505 & ~n17842 ;
  assign n17845 = ~n17843 & n17844 ;
  assign n17838 = ~\P1_P3_rEIP_reg[16]/NET0131  & ~n16581 ;
  assign n17839 = ~n16582 & ~n17838 ;
  assign n17840 = n16505 & ~n17839 ;
  assign n17846 = n16500 & ~n17840 ;
  assign n17847 = ~n17845 & n17846 ;
  assign n17848 = \P1_P3_rEIP_reg[16]/NET0131  & ~n9195 ;
  assign n17850 = ~n9095 & n17840 ;
  assign n17849 = ~\P1_P3_EBX_reg[16]/NET0131  & ~n16517 ;
  assign n17851 = n9236 & ~n17849 ;
  assign n17852 = ~n17850 & n17851 ;
  assign n17853 = ~n17848 & ~n17852 ;
  assign n17854 = ~n17847 & n17853 ;
  assign n17855 = n9241 & ~n17854 ;
  assign n17827 = \P1_P3_rEIP_reg[16]/NET0131  & ~n17458 ;
  assign n17856 = \P1_P3_PhyAddrPointer_reg[16]/NET0131  & n10031 ;
  assign n17857 = ~n17426 & ~n17856 ;
  assign n17858 = ~n17827 & n17857 ;
  assign n17859 = ~n17855 & n17858 ;
  assign n17860 = ~n17837 & n17859 ;
  assign n17863 = n16484 & ~n16554 ;
  assign n17865 = ~n16544 & n17863 ;
  assign n17864 = n16544 & ~n17863 ;
  assign n17866 = ~\P1_P3_DataWidth_reg[1]/NET0131  & ~n17864 ;
  assign n17867 = ~n17865 & n17866 ;
  assign n17862 = \P1_P3_DataWidth_reg[1]/NET0131  & ~\P1_P3_rEIP_reg[19]/NET0131  ;
  assign n17868 = n9245 & ~n17862 ;
  assign n17869 = ~n17867 & n17868 ;
  assign n17882 = \P1_P3_EBX_reg[31]/NET0131  & ~n16611 ;
  assign n17884 = ~\P1_P3_EBX_reg[19]/NET0131  & n17882 ;
  assign n17883 = \P1_P3_EBX_reg[19]/NET0131  & ~n17882 ;
  assign n17885 = ~n16505 & ~n17883 ;
  assign n17886 = ~n17884 & n17885 ;
  assign n17873 = ~\P1_P3_rEIP_reg[19]/NET0131  & ~n16584 ;
  assign n17874 = ~n16585 & ~n17873 ;
  assign n17875 = n16505 & ~n17874 ;
  assign n17887 = n16500 & ~n17875 ;
  assign n17888 = ~n17886 & n17887 ;
  assign n17870 = \P1_P3_rEIP_reg[19]/NET0131  & ~n16565 ;
  assign n17876 = ~\P1_P3_EBX_reg[19]/NET0131  & ~n16505 ;
  assign n17877 = n9162 & ~n17876 ;
  assign n17878 = ~n17875 & n17877 ;
  assign n17871 = \P1_P3_EBX_reg[19]/NET0131  & n16567 ;
  assign n17872 = \P1_P3_rEIP_reg[19]/NET0131  & n9075 ;
  assign n17879 = ~n17871 & ~n17872 ;
  assign n17880 = ~n17878 & n17879 ;
  assign n17881 = n9079 & ~n17880 ;
  assign n17889 = ~n17870 & ~n17881 ;
  assign n17890 = ~n17888 & n17889 ;
  assign n17891 = n9241 & ~n17890 ;
  assign n17861 = \P1_P3_rEIP_reg[19]/NET0131  & ~n17458 ;
  assign n17892 = \P1_P3_PhyAddrPointer_reg[19]/NET0131  & n10031 ;
  assign n17893 = ~n17426 & ~n17892 ;
  assign n17894 = ~n17861 & n17893 ;
  assign n17895 = ~n17891 & n17894 ;
  assign n17896 = ~n17869 & n17895 ;
  assign n17899 = ~\P1_P3_PhyAddrPointer_reg[9]/NET0131  & ~n17661 ;
  assign n17900 = ~n17662 & ~n17899 ;
  assign n17901 = \P1_P3_PhyAddrPointer_reg[8]/NET0131  & n17666 ;
  assign n17902 = n16484 & ~n17901 ;
  assign n17904 = ~n17900 & n17902 ;
  assign n17903 = n17900 & ~n17902 ;
  assign n17905 = ~\P1_P3_DataWidth_reg[1]/NET0131  & ~n17903 ;
  assign n17906 = ~n17904 & n17905 ;
  assign n17898 = \P1_P3_DataWidth_reg[1]/NET0131  & ~\P1_P3_rEIP_reg[9]/NET0131  ;
  assign n17907 = n9245 & ~n17898 ;
  assign n17908 = ~n17906 & n17907 ;
  assign n17909 = \P1_P3_rEIP_reg[9]/NET0131  & ~n9195 ;
  assign n17910 = \P1_P3_EBX_reg[31]/NET0131  & ~n16601 ;
  assign n17912 = \P1_P3_EBX_reg[9]/NET0131  & n17910 ;
  assign n17911 = ~\P1_P3_EBX_reg[9]/NET0131  & ~n17910 ;
  assign n17913 = ~n16505 & ~n17911 ;
  assign n17914 = ~n17912 & n17913 ;
  assign n17915 = ~\P1_P3_rEIP_reg[9]/NET0131  & ~n16574 ;
  assign n17916 = ~n16575 & ~n17915 ;
  assign n17917 = ~\P1_P3_DataWidth_reg[1]/NET0131  & n17916 ;
  assign n17918 = ~n8741 & n17917 ;
  assign n17919 = ~n17914 & ~n17918 ;
  assign n17920 = n9085 & ~n17919 ;
  assign n17921 = \P1_P3_EBX_reg[9]/NET0131  & ~n16517 ;
  assign n17922 = n9096 & n17917 ;
  assign n17923 = ~n17921 & ~n17922 ;
  assign n17924 = n9079 & ~n17923 ;
  assign n17925 = ~n17920 & ~n17924 ;
  assign n17926 = ~n9075 & ~n17925 ;
  assign n17927 = ~n17909 & ~n17926 ;
  assign n17928 = n9241 & ~n17927 ;
  assign n17897 = \P1_P3_rEIP_reg[9]/NET0131  & ~n17458 ;
  assign n17929 = \P1_P3_PhyAddrPointer_reg[9]/NET0131  & n10031 ;
  assign n17930 = ~n17426 & ~n17929 ;
  assign n17931 = ~n17897 & n17930 ;
  assign n17932 = ~n17928 & n17931 ;
  assign n17933 = ~n17908 & n17932 ;
  assign n17936 = n16484 & ~n17666 ;
  assign n17937 = ~\P1_P3_PhyAddrPointer_reg[8]/NET0131  & ~n17606 ;
  assign n17938 = ~n17661 & ~n17937 ;
  assign n17940 = n17936 & ~n17938 ;
  assign n17939 = ~n17936 & n17938 ;
  assign n17941 = ~\P1_P3_DataWidth_reg[1]/NET0131  & ~n17939 ;
  assign n17942 = ~n17940 & n17941 ;
  assign n17935 = \P1_P3_DataWidth_reg[1]/NET0131  & ~\P1_P3_rEIP_reg[8]/NET0131  ;
  assign n17943 = n9245 & ~n17935 ;
  assign n17944 = ~n17942 & n17943 ;
  assign n17945 = \P1_P3_rEIP_reg[8]/NET0131  & ~n9195 ;
  assign n17946 = ~\P1_P3_EBX_reg[8]/NET0131  & ~n16517 ;
  assign n17947 = ~\P1_P3_rEIP_reg[8]/NET0131  & ~n16573 ;
  assign n17948 = ~n16574 & ~n17947 ;
  assign n17949 = n16517 & ~n17948 ;
  assign n17950 = ~n17946 & ~n17949 ;
  assign n17951 = n9079 & n17950 ;
  assign n17953 = \P1_P3_EBX_reg[31]/NET0131  & ~n16600 ;
  assign n17955 = \P1_P3_EBX_reg[8]/NET0131  & ~n17953 ;
  assign n17954 = ~\P1_P3_EBX_reg[8]/NET0131  & n17953 ;
  assign n17956 = ~n16505 & ~n17954 ;
  assign n17957 = ~n17955 & n17956 ;
  assign n17952 = n16505 & ~n17948 ;
  assign n17958 = n9085 & ~n17952 ;
  assign n17959 = ~n17957 & n17958 ;
  assign n17960 = ~n17951 & ~n17959 ;
  assign n17961 = ~n9075 & ~n17960 ;
  assign n17962 = ~n17945 & ~n17961 ;
  assign n17963 = n9241 & ~n17962 ;
  assign n17934 = \P1_P3_rEIP_reg[8]/NET0131  & ~n17458 ;
  assign n17964 = \P1_P3_PhyAddrPointer_reg[8]/NET0131  & n10031 ;
  assign n17965 = ~n17426 & ~n17964 ;
  assign n17966 = ~n17934 & n17965 ;
  assign n17967 = ~n17963 & n17966 ;
  assign n17968 = ~n17944 & n17967 ;
  assign n17970 = ~n11862 & ~n17381 ;
  assign n17969 = n11862 & ~n17378 ;
  assign n17971 = n12388 & ~n17969 ;
  assign n17972 = ~n17970 & n17971 ;
  assign n17975 = n11871 & n17417 ;
  assign n17974 = ~\P2_P1_InstQueue_reg[0][0]/NET0131  & ~n11871 ;
  assign n17976 = n11692 & ~n17974 ;
  assign n17977 = ~n17975 & n17976 ;
  assign n17973 = \P2_P1_InstQueue_reg[0][0]/NET0131  & ~n12395 ;
  assign n17978 = n11379 & ~n11874 ;
  assign n17979 = n12393 & n17978 ;
  assign n17980 = ~n17973 & ~n17979 ;
  assign n17981 = ~n17977 & n17980 ;
  assign n17982 = ~n17972 & n17981 ;
  assign n17984 = ~n11891 & ~n17381 ;
  assign n17983 = n11891 & ~n17378 ;
  assign n17985 = n12407 & ~n17983 ;
  assign n17986 = ~n17984 & n17985 ;
  assign n17989 = n11599 & n17417 ;
  assign n17988 = ~\P2_P1_InstQueue_reg[10][0]/NET0131  & ~n11599 ;
  assign n17990 = n11692 & ~n17988 ;
  assign n17991 = ~n17989 & n17990 ;
  assign n17987 = \P2_P1_InstQueue_reg[10][0]/NET0131  & ~n12414 ;
  assign n17992 = n11379 & ~n11897 ;
  assign n17993 = n12412 & n17992 ;
  assign n17994 = ~n17987 & ~n17993 ;
  assign n17995 = ~n17991 & n17994 ;
  assign n17996 = ~n17986 & n17995 ;
  assign n17998 = ~n11577 & ~n17381 ;
  assign n17997 = n11577 & ~n17378 ;
  assign n17999 = n12426 & ~n17997 ;
  assign n18000 = ~n17998 & n17999 ;
  assign n18003 = n11919 & n17417 ;
  assign n18002 = ~\P2_P1_InstQueue_reg[12][0]/NET0131  & ~n11919 ;
  assign n18004 = n11692 & ~n18002 ;
  assign n18005 = ~n18003 & n18004 ;
  assign n18001 = \P2_P1_InstQueue_reg[12][0]/NET0131  & ~n12433 ;
  assign n18006 = n11379 & ~n11920 ;
  assign n18007 = n12431 & n18006 ;
  assign n18008 = ~n18001 & ~n18007 ;
  assign n18009 = ~n18005 & n18008 ;
  assign n18010 = ~n18000 & n18009 ;
  assign n18012 = ~n11599 & ~n17381 ;
  assign n18011 = n11599 & ~n17378 ;
  assign n18013 = n12445 & ~n18011 ;
  assign n18014 = ~n18012 & n18013 ;
  assign n18017 = n11862 & n17417 ;
  assign n18016 = ~\P2_P1_InstQueue_reg[13][0]/NET0131  & ~n11862 ;
  assign n18018 = n11692 & ~n18016 ;
  assign n18019 = ~n18017 & n18018 ;
  assign n18015 = \P2_P1_InstQueue_reg[13][0]/NET0131  & ~n12452 ;
  assign n18020 = n11379 & ~n11961 ;
  assign n18021 = n12450 & n18020 ;
  assign n18022 = ~n18015 & ~n18021 ;
  assign n18023 = ~n18019 & n18022 ;
  assign n18024 = ~n18014 & n18023 ;
  assign n18026 = ~n11596 & ~n17381 ;
  assign n18025 = n11596 & ~n17378 ;
  assign n18027 = n12464 & ~n18025 ;
  assign n18028 = ~n18026 & n18027 ;
  assign n18031 = n11865 & n17417 ;
  assign n18030 = ~\P2_P1_InstQueue_reg[14][0]/NET0131  & ~n11865 ;
  assign n18032 = n11692 & ~n18030 ;
  assign n18033 = ~n18031 & n18032 ;
  assign n18029 = \P2_P1_InstQueue_reg[14][0]/NET0131  & ~n12471 ;
  assign n18034 = n11379 & ~n11869 ;
  assign n18035 = n12469 & n18034 ;
  assign n18036 = ~n18029 & ~n18035 ;
  assign n18037 = ~n18033 & n18036 ;
  assign n18038 = ~n18028 & n18037 ;
  assign n18040 = ~n11919 & ~n17381 ;
  assign n18039 = n11919 & ~n17378 ;
  assign n18041 = n12483 & ~n18039 ;
  assign n18042 = ~n18040 & n18041 ;
  assign n18045 = n11873 & n17417 ;
  assign n18044 = ~\P2_P1_InstQueue_reg[15][0]/NET0131  & ~n11873 ;
  assign n18046 = n11692 & ~n18044 ;
  assign n18047 = ~n18045 & n18046 ;
  assign n18043 = \P2_P1_InstQueue_reg[15][0]/NET0131  & ~n12490 ;
  assign n18048 = n11379 & ~n12002 ;
  assign n18049 = n12488 & n18048 ;
  assign n18050 = ~n18043 & ~n18049 ;
  assign n18051 = ~n18047 & n18050 ;
  assign n18052 = ~n18042 & n18051 ;
  assign n18054 = ~n11865 & ~n17381 ;
  assign n18053 = n11865 & ~n17378 ;
  assign n18055 = n12502 & ~n18053 ;
  assign n18056 = ~n18054 & n18055 ;
  assign n18059 = n12023 & n17417 ;
  assign n18058 = ~\P2_P1_InstQueue_reg[1][0]/NET0131  & ~n12023 ;
  assign n18060 = n11692 & ~n18058 ;
  assign n18061 = ~n18059 & n18060 ;
  assign n18057 = \P2_P1_InstQueue_reg[1][0]/NET0131  & ~n12509 ;
  assign n18062 = n11379 & ~n12024 ;
  assign n18063 = n12507 & n18062 ;
  assign n18064 = ~n18057 & ~n18063 ;
  assign n18065 = ~n18061 & n18064 ;
  assign n18066 = ~n18056 & n18065 ;
  assign n18068 = ~n11873 & ~n17381 ;
  assign n18067 = n11873 & ~n17378 ;
  assign n18069 = n12521 & ~n18067 ;
  assign n18070 = ~n18068 & n18069 ;
  assign n18073 = n12065 & n17417 ;
  assign n18072 = ~\P2_P1_InstQueue_reg[2][0]/NET0131  & ~n12065 ;
  assign n18074 = n11692 & ~n18072 ;
  assign n18075 = ~n18073 & n18074 ;
  assign n18071 = \P2_P1_InstQueue_reg[2][0]/NET0131  & ~n12528 ;
  assign n18076 = n11379 & ~n12066 ;
  assign n18077 = n12526 & n18076 ;
  assign n18078 = ~n18071 & ~n18077 ;
  assign n18079 = ~n18075 & n18078 ;
  assign n18080 = ~n18070 & n18079 ;
  assign n18082 = ~n11871 & ~n17381 ;
  assign n18081 = n11871 & ~n17378 ;
  assign n18083 = n12540 & ~n18081 ;
  assign n18084 = ~n18082 & n18083 ;
  assign n18087 = n12087 & n17417 ;
  assign n18086 = ~\P2_P1_InstQueue_reg[3][0]/NET0131  & ~n12087 ;
  assign n18088 = n11692 & ~n18086 ;
  assign n18089 = ~n18087 & n18088 ;
  assign n18085 = \P2_P1_InstQueue_reg[3][0]/NET0131  & ~n12547 ;
  assign n18090 = n11379 & ~n12088 ;
  assign n18091 = n12545 & n18090 ;
  assign n18092 = ~n18085 & ~n18091 ;
  assign n18093 = ~n18089 & n18092 ;
  assign n18094 = ~n18084 & n18093 ;
  assign n18096 = ~n12023 & ~n17381 ;
  assign n18095 = n12023 & ~n17378 ;
  assign n18097 = n12559 & ~n18095 ;
  assign n18098 = ~n18096 & n18097 ;
  assign n18101 = n12109 & n17417 ;
  assign n18100 = ~\P2_P1_InstQueue_reg[4][0]/NET0131  & ~n12109 ;
  assign n18102 = n11692 & ~n18100 ;
  assign n18103 = ~n18101 & n18102 ;
  assign n18099 = \P2_P1_InstQueue_reg[4][0]/NET0131  & ~n12566 ;
  assign n18104 = n11379 & ~n12110 ;
  assign n18105 = n12564 & n18104 ;
  assign n18106 = ~n18099 & ~n18105 ;
  assign n18107 = ~n18103 & n18106 ;
  assign n18108 = ~n18098 & n18107 ;
  assign n18110 = ~n12065 & ~n17381 ;
  assign n18109 = n12065 & ~n17378 ;
  assign n18111 = n12578 & ~n18109 ;
  assign n18112 = ~n18110 & n18111 ;
  assign n18115 = n12131 & n17417 ;
  assign n18114 = ~\P2_P1_InstQueue_reg[5][0]/NET0131  & ~n12131 ;
  assign n18116 = n11692 & ~n18114 ;
  assign n18117 = ~n18115 & n18116 ;
  assign n18113 = \P2_P1_InstQueue_reg[5][0]/NET0131  & ~n12585 ;
  assign n18118 = n11379 & ~n12132 ;
  assign n18119 = n12583 & n18118 ;
  assign n18120 = ~n18113 & ~n18119 ;
  assign n18121 = ~n18117 & n18120 ;
  assign n18122 = ~n18112 & n18121 ;
  assign n18124 = ~n12087 & ~n17381 ;
  assign n18123 = n12087 & ~n17378 ;
  assign n18125 = n12597 & ~n18123 ;
  assign n18126 = ~n18124 & n18125 ;
  assign n18129 = n12173 & n17417 ;
  assign n18128 = ~\P2_P1_InstQueue_reg[6][0]/NET0131  & ~n12173 ;
  assign n18130 = n11692 & ~n18128 ;
  assign n18131 = ~n18129 & n18130 ;
  assign n18127 = \P2_P1_InstQueue_reg[6][0]/NET0131  & ~n12604 ;
  assign n18132 = n11379 & ~n12174 ;
  assign n18133 = n12602 & n18132 ;
  assign n18134 = ~n18127 & ~n18133 ;
  assign n18135 = ~n18131 & n18134 ;
  assign n18136 = ~n18126 & n18135 ;
  assign n18138 = ~n12109 & ~n17381 ;
  assign n18137 = n12109 & ~n17378 ;
  assign n18139 = n12616 & ~n18137 ;
  assign n18140 = ~n18138 & n18139 ;
  assign n18143 = n11891 & n17417 ;
  assign n18142 = ~\P2_P1_InstQueue_reg[7][0]/NET0131  & ~n11891 ;
  assign n18144 = n11692 & ~n18142 ;
  assign n18145 = ~n18143 & n18144 ;
  assign n18141 = \P2_P1_InstQueue_reg[7][0]/NET0131  & ~n12623 ;
  assign n18146 = n11379 & ~n12195 ;
  assign n18147 = n12621 & n18146 ;
  assign n18148 = ~n18141 & ~n18147 ;
  assign n18149 = ~n18145 & n18148 ;
  assign n18150 = ~n18140 & n18149 ;
  assign n18152 = ~n12131 & ~n17381 ;
  assign n18151 = n12131 & ~n17378 ;
  assign n18153 = n12635 & ~n18151 ;
  assign n18154 = ~n18152 & n18153 ;
  assign n18157 = n10105 & n17417 ;
  assign n18156 = ~\P2_P1_InstQueue_reg[8][0]/NET0131  & ~n10105 ;
  assign n18158 = n11692 & ~n18156 ;
  assign n18159 = ~n18157 & n18158 ;
  assign n18155 = \P2_P1_InstQueue_reg[8][0]/NET0131  & ~n12642 ;
  assign n18160 = n11379 & ~n11895 ;
  assign n18161 = n12640 & n18160 ;
  assign n18162 = ~n18155 & ~n18161 ;
  assign n18163 = ~n18159 & n18162 ;
  assign n18164 = ~n18154 & n18163 ;
  assign n18166 = ~n12173 & ~n17381 ;
  assign n18165 = n12173 & ~n17378 ;
  assign n18167 = n12654 & ~n18165 ;
  assign n18168 = ~n18166 & n18167 ;
  assign n18171 = n11577 & n17417 ;
  assign n18170 = ~\P2_P1_InstQueue_reg[9][0]/NET0131  & ~n11577 ;
  assign n18172 = n11692 & ~n18170 ;
  assign n18173 = ~n18171 & n18172 ;
  assign n18169 = \P2_P1_InstQueue_reg[9][0]/NET0131  & ~n12661 ;
  assign n18174 = n11379 & ~n11592 ;
  assign n18175 = n12659 & n18174 ;
  assign n18176 = ~n18169 & ~n18175 ;
  assign n18177 = ~n18173 & n18176 ;
  assign n18178 = ~n18168 & n18177 ;
  assign n18180 = n9079 & n9162 ;
  assign n18181 = ~n16500 & ~n18180 ;
  assign n18185 = ~n16505 & ~n18181 ;
  assign n18186 = n9095 & n9236 ;
  assign n18187 = ~n18185 & ~n18186 ;
  assign n18188 = \P1_P3_EBX_reg[0]/NET0131  & ~n18187 ;
  assign n18179 = ~\P1_P3_InstQueueRd_Addr_reg[0]/NET0131  & n16498 ;
  assign n18182 = n16505 & ~n18181 ;
  assign n18183 = n9195 & ~n18182 ;
  assign n18184 = \P1_P3_rEIP_reg[0]/NET0131  & ~n18183 ;
  assign n18189 = ~n18179 & ~n18184 ;
  assign n18190 = ~n18188 & n18189 ;
  assign n18191 = n9241 & ~n18190 ;
  assign n18192 = ~n9246 & ~n10031 ;
  assign n18193 = \P1_P3_PhyAddrPointer_reg[0]/NET0131  & ~n18192 ;
  assign n18194 = ~n11698 & n16495 ;
  assign n18195 = \P1_P3_rEIP_reg[0]/NET0131  & ~n18194 ;
  assign n18196 = ~n18193 & ~n18195 ;
  assign n18197 = ~n18191 & n18196 ;
  assign n18200 = n16484 & ~n16791 ;
  assign n18202 = n16794 & ~n18200 ;
  assign n18201 = ~n16794 & n18200 ;
  assign n18203 = ~\P1_P3_DataWidth_reg[1]/NET0131  & ~n18201 ;
  assign n18204 = ~n18202 & n18203 ;
  assign n18199 = \P1_P3_DataWidth_reg[1]/NET0131  & ~\P1_P3_rEIP_reg[25]/NET0131  ;
  assign n18205 = n9245 & ~n18199 ;
  assign n18206 = ~n18204 & n18205 ;
  assign n18220 = \P1_P3_EBX_reg[31]/NET0131  & ~n16812 ;
  assign n18222 = ~\P1_P3_EBX_reg[25]/NET0131  & n18220 ;
  assign n18221 = \P1_P3_EBX_reg[25]/NET0131  & ~n18220 ;
  assign n18223 = ~n16505 & ~n18221 ;
  assign n18224 = ~n18222 & n18223 ;
  assign n18211 = ~\P1_P3_rEIP_reg[25]/NET0131  & ~n16759 ;
  assign n18212 = ~n16807 & ~n18211 ;
  assign n18213 = n16505 & ~n18212 ;
  assign n18225 = n16500 & ~n18213 ;
  assign n18226 = ~n18224 & n18225 ;
  assign n18208 = \P1_P3_rEIP_reg[25]/NET0131  & ~n16565 ;
  assign n18214 = ~\P1_P3_EBX_reg[25]/NET0131  & ~n16505 ;
  assign n18215 = n9162 & ~n18214 ;
  assign n18216 = ~n18213 & n18215 ;
  assign n18209 = \P1_P3_rEIP_reg[25]/NET0131  & n9075 ;
  assign n18210 = \P1_P3_EBX_reg[25]/NET0131  & n16567 ;
  assign n18217 = ~n18209 & ~n18210 ;
  assign n18218 = ~n18216 & n18217 ;
  assign n18219 = n9079 & ~n18218 ;
  assign n18227 = ~n18208 & ~n18219 ;
  assign n18228 = ~n18226 & n18227 ;
  assign n18229 = n9241 & ~n18228 ;
  assign n18198 = \P1_P3_PhyAddrPointer_reg[25]/NET0131  & n10031 ;
  assign n18207 = \P1_P3_rEIP_reg[25]/NET0131  & ~n16495 ;
  assign n18230 = ~n18198 & ~n18207 ;
  assign n18231 = ~n18229 & n18230 ;
  assign n18232 = ~n18206 & n18231 ;
  assign n18260 = n16896 & ~n16900 ;
  assign n18261 = n16484 & ~n18260 ;
  assign n18262 = ~\P1_P3_PhyAddrPointer_reg[29]/NET0131  & ~n16899 ;
  assign n18263 = \P1_P3_PhyAddrPointer_reg[1]/NET0131  & n16479 ;
  assign n18264 = ~n18262 & ~n18263 ;
  assign n18266 = ~n18261 & n18264 ;
  assign n18265 = n18261 & ~n18264 ;
  assign n18267 = ~\P1_P3_DataWidth_reg[1]/NET0131  & ~n18265 ;
  assign n18268 = ~n18266 & n18267 ;
  assign n18259 = \P1_P3_DataWidth_reg[1]/NET0131  & ~\P1_P3_rEIP_reg[29]/NET0131  ;
  assign n18269 = n9245 & ~n18259 ;
  assign n18270 = ~n18268 & n18269 ;
  assign n18248 = ~\P1_P3_EBX_reg[28]/NET0131  & n16878 ;
  assign n18249 = \P1_P3_EBX_reg[31]/NET0131  & ~n18248 ;
  assign n18251 = ~\P1_P3_EBX_reg[29]/NET0131  & n18249 ;
  assign n18250 = \P1_P3_EBX_reg[29]/NET0131  & ~n18249 ;
  assign n18252 = ~n16505 & ~n18250 ;
  assign n18253 = ~n18251 & n18252 ;
  assign n18238 = \P1_P3_rEIP_reg[29]/NET0131  & n16875 ;
  assign n18239 = ~\P1_P3_rEIP_reg[29]/NET0131  & ~n16875 ;
  assign n18240 = ~n18238 & ~n18239 ;
  assign n18241 = n16505 & ~n18240 ;
  assign n18254 = n16500 & ~n18241 ;
  assign n18255 = ~n18253 & n18254 ;
  assign n18235 = \P1_P3_rEIP_reg[29]/NET0131  & ~n16565 ;
  assign n18242 = ~\P1_P3_EBX_reg[29]/NET0131  & ~n16505 ;
  assign n18243 = n9162 & ~n18242 ;
  assign n18244 = ~n18241 & n18243 ;
  assign n18236 = \P1_P3_EBX_reg[29]/NET0131  & n16567 ;
  assign n18237 = \P1_P3_rEIP_reg[29]/NET0131  & n9075 ;
  assign n18245 = ~n18236 & ~n18237 ;
  assign n18246 = ~n18244 & n18245 ;
  assign n18247 = n9079 & ~n18246 ;
  assign n18256 = ~n18235 & ~n18247 ;
  assign n18257 = ~n18255 & n18256 ;
  assign n18258 = n9241 & ~n18257 ;
  assign n18233 = \P1_P3_PhyAddrPointer_reg[29]/NET0131  & n10031 ;
  assign n18234 = \P1_P3_rEIP_reg[29]/NET0131  & ~n16495 ;
  assign n18271 = ~n18233 & ~n18234 ;
  assign n18272 = ~n18258 & n18271 ;
  assign n18273 = ~n18270 & n18272 ;
  assign n18297 = n18260 & ~n18264 ;
  assign n18298 = n16484 & ~n18297 ;
  assign n18299 = ~\P1_P3_PhyAddrPointer_reg[30]/NET0131  & ~n18263 ;
  assign n18300 = ~n16481 & ~n18299 ;
  assign n18302 = ~n18298 & n18300 ;
  assign n18301 = n18298 & ~n18300 ;
  assign n18303 = ~\P1_P3_DataWidth_reg[1]/NET0131  & ~n18301 ;
  assign n18304 = ~n18302 & n18303 ;
  assign n18296 = \P1_P3_DataWidth_reg[1]/NET0131  & ~\P1_P3_rEIP_reg[30]/NET0131  ;
  assign n18305 = n9245 & ~n18296 ;
  assign n18306 = ~n18304 & n18305 ;
  assign n18280 = ~\P1_P3_EBX_reg[29]/NET0131  & n18248 ;
  assign n18281 = \P1_P3_EBX_reg[31]/NET0131  & ~n18280 ;
  assign n18283 = ~\P1_P3_EBX_reg[30]/NET0131  & n18281 ;
  assign n18282 = \P1_P3_EBX_reg[30]/NET0131  & ~n18281 ;
  assign n18284 = ~n16505 & ~n18282 ;
  assign n18285 = ~n18283 & n18284 ;
  assign n18276 = ~\P1_P3_rEIP_reg[30]/NET0131  & ~n18238 ;
  assign n18277 = \P1_P3_rEIP_reg[30]/NET0131  & n18238 ;
  assign n18278 = ~n18276 & ~n18277 ;
  assign n18279 = n16505 & ~n18278 ;
  assign n18286 = n16500 & ~n18279 ;
  assign n18287 = ~n18285 & n18286 ;
  assign n18288 = \P1_P3_rEIP_reg[30]/NET0131  & ~n9195 ;
  assign n18290 = ~n9095 & n18279 ;
  assign n18289 = ~\P1_P3_EBX_reg[30]/NET0131  & ~n16517 ;
  assign n18291 = n9236 & ~n18289 ;
  assign n18292 = ~n18290 & n18291 ;
  assign n18293 = ~n18288 & ~n18292 ;
  assign n18294 = ~n18287 & n18293 ;
  assign n18295 = n9241 & ~n18294 ;
  assign n18274 = \P1_P3_PhyAddrPointer_reg[30]/NET0131  & n10031 ;
  assign n18275 = \P1_P3_rEIP_reg[30]/NET0131  & ~n16495 ;
  assign n18307 = ~n18274 & ~n18275 ;
  assign n18308 = ~n18295 & n18307 ;
  assign n18309 = ~n18306 & n18308 ;
  assign n18322 = \P1_P3_EBX_reg[31]/NET0131  & ~n16517 ;
  assign n18316 = \P1_P3_rEIP_reg[31]/NET0131  & n18277 ;
  assign n18315 = ~\P1_P3_rEIP_reg[31]/NET0131  & ~n18277 ;
  assign n18317 = ~\P1_P3_DataWidth_reg[1]/NET0131  & ~n18315 ;
  assign n18318 = ~n18316 & n18317 ;
  assign n18323 = n9096 & n18318 ;
  assign n18324 = ~n18322 & ~n18323 ;
  assign n18325 = n9236 & ~n18324 ;
  assign n18311 = \P1_P3_rEIP_reg[31]/NET0131  & ~n9195 ;
  assign n18312 = ~\P1_P3_EBX_reg[30]/NET0131  & \P1_P3_EBX_reg[31]/NET0131  ;
  assign n18313 = ~n16505 & n18312 ;
  assign n18314 = n18280 & n18313 ;
  assign n18319 = ~n8741 & n18318 ;
  assign n18320 = ~n18314 & ~n18319 ;
  assign n18321 = n16500 & ~n18320 ;
  assign n18326 = ~n18311 & ~n18321 ;
  assign n18327 = ~n18325 & n18326 ;
  assign n18328 = n9241 & ~n18327 ;
  assign n18329 = \P1_P3_DataWidth_reg[1]/NET0131  & \P1_P3_rEIP_reg[31]/NET0131  ;
  assign n18330 = ~\P1_P3_DataWidth_reg[1]/NET0131  & ~n18300 ;
  assign n18331 = n16484 & n18297 ;
  assign n18332 = n18330 & n18331 ;
  assign n18333 = ~n18329 & ~n18332 ;
  assign n18334 = n9245 & ~n18333 ;
  assign n18310 = \P1_P3_PhyAddrPointer_reg[31]/NET0131  & n10031 ;
  assign n18335 = \P1_P3_rEIP_reg[31]/NET0131  & ~n16495 ;
  assign n18336 = ~n18310 & ~n18335 ;
  assign n18337 = ~n18334 & n18336 ;
  assign n18338 = ~n18328 & n18337 ;
  assign n18432 = ~\P1_P3_InstAddrPointer_reg[1]/NET0131  & n9176 ;
  assign n18433 = n9084 & ~n9147 ;
  assign n18434 = n8741 & ~n18433 ;
  assign n18435 = ~n9050 & ~n9135 ;
  assign n18436 = ~n9062 & n18435 ;
  assign n18437 = ~n9163 & n18436 ;
  assign n18438 = ~n18434 & n18437 ;
  assign n18439 = ~\P1_P3_InstAddrPointer_reg[0]/NET0131  & ~n9061 ;
  assign n18440 = \P1_P3_InstAddrPointer_reg[1]/NET0131  & ~n9073 ;
  assign n18441 = ~n18439 & n18440 ;
  assign n18442 = n18438 & n18441 ;
  assign n18443 = ~n18432 & ~n18442 ;
  assign n18349 = \P1_P3_InstQueue_reg[10][1]/NET0131  & n8763 ;
  assign n18350 = \P1_P3_InstQueue_reg[4][1]/NET0131  & n8771 ;
  assign n18363 = ~n18349 & ~n18350 ;
  assign n18351 = \P1_P3_InstQueue_reg[1][1]/NET0131  & n8767 ;
  assign n18352 = \P1_P3_InstQueue_reg[8][1]/NET0131  & n8748 ;
  assign n18364 = ~n18351 & ~n18352 ;
  assign n18371 = n18363 & n18364 ;
  assign n18345 = \P1_P3_InstQueue_reg[12][1]/NET0131  & n8765 ;
  assign n18346 = \P1_P3_InstQueue_reg[9][1]/NET0131  & n8769 ;
  assign n18361 = ~n18345 & ~n18346 ;
  assign n18347 = \P1_P3_InstQueue_reg[13][1]/NET0131  & n8760 ;
  assign n18348 = \P1_P3_InstQueue_reg[14][1]/NET0131  & n8775 ;
  assign n18362 = ~n18347 & ~n18348 ;
  assign n18372 = n18361 & n18362 ;
  assign n18373 = n18371 & n18372 ;
  assign n18357 = \P1_P3_InstQueue_reg[6][1]/NET0131  & n8779 ;
  assign n18358 = \P1_P3_InstQueue_reg[15][1]/NET0131  & n8781 ;
  assign n18367 = ~n18357 & ~n18358 ;
  assign n18359 = \P1_P3_InstQueue_reg[11][1]/NET0131  & n8757 ;
  assign n18360 = \P1_P3_InstQueue_reg[3][1]/NET0131  & n8752 ;
  assign n18368 = ~n18359 & ~n18360 ;
  assign n18369 = n18367 & n18368 ;
  assign n18353 = \P1_P3_InstQueue_reg[0][1]/NET0131  & n8773 ;
  assign n18354 = \P1_P3_InstQueue_reg[7][1]/NET0131  & n8754 ;
  assign n18365 = ~n18353 & ~n18354 ;
  assign n18355 = \P1_P3_InstQueue_reg[2][1]/NET0131  & n8777 ;
  assign n18356 = \P1_P3_InstQueue_reg[5][1]/NET0131  & n8745 ;
  assign n18366 = ~n18355 & ~n18356 ;
  assign n18370 = n18365 & n18366 ;
  assign n18374 = n18369 & n18370 ;
  assign n18375 = n18373 & n18374 ;
  assign n18376 = ~n15309 & n18375 ;
  assign n18377 = n15309 & ~n18375 ;
  assign n18378 = ~n18376 & ~n18377 ;
  assign n18383 = \P1_P3_InstQueue_reg[11][0]/NET0131  & n8757 ;
  assign n18384 = \P1_P3_InstQueue_reg[1][0]/NET0131  & n8767 ;
  assign n18397 = ~n18383 & ~n18384 ;
  assign n18385 = \P1_P3_InstQueue_reg[5][0]/NET0131  & n8745 ;
  assign n18386 = \P1_P3_InstQueue_reg[7][0]/NET0131  & n8754 ;
  assign n18398 = ~n18385 & ~n18386 ;
  assign n18405 = n18397 & n18398 ;
  assign n18379 = \P1_P3_InstQueue_reg[6][0]/NET0131  & n8779 ;
  assign n18380 = \P1_P3_InstQueue_reg[14][0]/NET0131  & n8775 ;
  assign n18395 = ~n18379 & ~n18380 ;
  assign n18381 = \P1_P3_InstQueue_reg[2][0]/NET0131  & n8777 ;
  assign n18382 = \P1_P3_InstQueue_reg[3][0]/NET0131  & n8752 ;
  assign n18396 = ~n18381 & ~n18382 ;
  assign n18406 = n18395 & n18396 ;
  assign n18407 = n18405 & n18406 ;
  assign n18391 = \P1_P3_InstQueue_reg[12][0]/NET0131  & n8765 ;
  assign n18392 = \P1_P3_InstQueue_reg[8][0]/NET0131  & n8748 ;
  assign n18401 = ~n18391 & ~n18392 ;
  assign n18393 = \P1_P3_InstQueue_reg[15][0]/NET0131  & n8781 ;
  assign n18394 = \P1_P3_InstQueue_reg[4][0]/NET0131  & n8771 ;
  assign n18402 = ~n18393 & ~n18394 ;
  assign n18403 = n18401 & n18402 ;
  assign n18387 = \P1_P3_InstQueue_reg[0][0]/NET0131  & n8773 ;
  assign n18388 = \P1_P3_InstQueue_reg[10][0]/NET0131  & n8763 ;
  assign n18399 = ~n18387 & ~n18388 ;
  assign n18389 = \P1_P3_InstQueue_reg[9][0]/NET0131  & n8769 ;
  assign n18390 = \P1_P3_InstQueue_reg[13][0]/NET0131  & n8760 ;
  assign n18400 = ~n18389 & ~n18390 ;
  assign n18404 = n18399 & n18400 ;
  assign n18408 = n18403 & n18404 ;
  assign n18409 = n18407 & n18408 ;
  assign n18410 = ~\P1_P3_InstAddrPointer_reg[0]/NET0131  & ~n18409 ;
  assign n18411 = ~n18378 & ~n18410 ;
  assign n18412 = ~\P1_P3_InstAddrPointer_reg[1]/NET0131  & ~n18375 ;
  assign n18413 = \P1_P3_InstAddrPointer_reg[1]/NET0131  & n18375 ;
  assign n18414 = ~n18412 & ~n18413 ;
  assign n18415 = n18410 & ~n18414 ;
  assign n18416 = ~n18411 & ~n18415 ;
  assign n18417 = n9191 & n18416 ;
  assign n18423 = \P1_P3_InstAddrPointer_reg[0]/NET0131  & n18409 ;
  assign n18425 = n18414 & n18423 ;
  assign n18424 = ~n18378 & ~n18423 ;
  assign n18426 = ~n17282 & ~n18424 ;
  assign n18427 = ~n18425 & n18426 ;
  assign n18418 = \P1_P3_InstAddrPointer_reg[0]/NET0131  & ~n18409 ;
  assign n18419 = ~n18414 & ~n18418 ;
  assign n18420 = n18414 & n18418 ;
  assign n18421 = ~n18419 & ~n18420 ;
  assign n18422 = n17282 & ~n18421 ;
  assign n18428 = n9192 & ~n18422 ;
  assign n18429 = ~n18427 & n18428 ;
  assign n18430 = ~n18417 & ~n18429 ;
  assign n18431 = ~n9221 & n15309 ;
  assign n18444 = n18430 & ~n18431 ;
  assign n18445 = ~n18443 & n18444 ;
  assign n18446 = n9241 & ~n18445 ;
  assign n18339 = \P1_P3_rEIP_reg[1]/NET0131  & n17426 ;
  assign n18340 = ~n9244 & ~n16492 ;
  assign n18341 = ~n10036 & n18340 ;
  assign n18342 = ~n8733 & n10029 ;
  assign n18343 = n18341 & ~n18342 ;
  assign n18344 = \P1_P3_InstAddrPointer_reg[1]/NET0131  & ~n18343 ;
  assign n18447 = ~n18339 & ~n18344 ;
  assign n18448 = ~n18446 & n18447 ;
  assign n18449 = ~n16110 & ~n16244 ;
  assign n18450 = ~n16095 & n18449 ;
  assign n18451 = ~n16083 & n18450 ;
  assign n18452 = ~n16071 & n18451 ;
  assign n18453 = ~n16061 & n18452 ;
  assign n18454 = ~n16048 & n18453 ;
  assign n18455 = ~n16131 & n18454 ;
  assign n18456 = ~n16147 & n18455 ;
  assign n18457 = ~n16035 & n18456 ;
  assign n18458 = ~n16021 & n18457 ;
  assign n18459 = ~n16006 & n18458 ;
  assign n18460 = ~n15991 & n18459 ;
  assign n18461 = ~n15976 & n18460 ;
  assign n18462 = ~n15963 & n18461 ;
  assign n18463 = ~n15949 & ~n16175 ;
  assign n18464 = ~n15936 & n18463 ;
  assign n18465 = ~n15922 & ~n16188 ;
  assign n18466 = n18464 & n18465 ;
  assign n18467 = n18462 & n18466 ;
  assign n18468 = ~n15895 & ~n15909 ;
  assign n18469 = ~n15884 & n18468 ;
  assign n18470 = n18467 & n18469 ;
  assign n18471 = ~n15856 & ~n15872 ;
  assign n18472 = n18470 & n18471 ;
  assign n18473 = ~n15832 & ~n15844 ;
  assign n18474 = n18472 & n18473 ;
  assign n18475 = ~n15809 & ~n15820 ;
  assign n18476 = n18474 & n18475 ;
  assign n18477 = n15794 & ~n18476 ;
  assign n18478 = ~n15794 & n18476 ;
  assign n18479 = ~n18477 & ~n18478 ;
  assign n18480 = ~\P4_IR_reg[28]/NET0131  & ~n18479 ;
  assign n18481 = \P4_IR_reg[28]/NET0131  & n15820 ;
  assign n18482 = ~n18480 & ~n18481 ;
  assign n18483 = n15734 & n15738 ;
  assign n18484 = n18482 & n18483 ;
  assign n18608 = ~n15896 & ~n16379 ;
  assign n18609 = ~n15923 & ~n16380 ;
  assign n18610 = ~n16036 & n16381 ;
  assign n18611 = ~n16155 & n18610 ;
  assign n18612 = ~n16007 & ~n16023 ;
  assign n18613 = ~n16009 & ~n18612 ;
  assign n18614 = ~n18611 & ~n18613 ;
  assign n18615 = n15993 & ~n18614 ;
  assign n18616 = ~n15977 & ~n15994 ;
  assign n18617 = ~n15979 & ~n18616 ;
  assign n18618 = ~n18615 & ~n18617 ;
  assign n18619 = n16191 & ~n18618 ;
  assign n18620 = ~n15964 & ~n16195 ;
  assign n18621 = ~n16189 & ~n18620 ;
  assign n18622 = ~n18619 & ~n18621 ;
  assign n18623 = ~n15950 & ~n16176 ;
  assign n18624 = ~n18622 & n18623 ;
  assign n18625 = ~n16194 & ~n16201 ;
  assign n18626 = ~n15950 & ~n18625 ;
  assign n18627 = ~n18624 & ~n18626 ;
  assign n18628 = ~n15923 & ~n15937 ;
  assign n18629 = ~n18627 & n18628 ;
  assign n18630 = ~n18609 & ~n18629 ;
  assign n18631 = ~n15896 & ~n15910 ;
  assign n18632 = ~n18630 & n18631 ;
  assign n18633 = ~n18608 & ~n18632 ;
  assign n18634 = ~n15885 & ~n18633 ;
  assign n18635 = n16378 & ~n18634 ;
  assign n18636 = n15874 & ~n18635 ;
  assign n18637 = n16408 & ~n18636 ;
  assign n18638 = n15846 & ~n18637 ;
  assign n18639 = n16376 & ~n18638 ;
  assign n18640 = ~n15821 & ~n18639 ;
  assign n18642 = ~n16319 & n18640 ;
  assign n18488 = ~n16251 & ~n16432 ;
  assign n18607 = ~n15734 & ~n18488 ;
  assign n18641 = n16319 & ~n18640 ;
  assign n18643 = n18607 & ~n18641 ;
  assign n18644 = ~n18642 & n18643 ;
  assign n18491 = ~n16261 & ~n16277 ;
  assign n18492 = ~n16329 & n18491 ;
  assign n18493 = ~n16276 & ~n16307 ;
  assign n18494 = ~n16274 & ~n16321 ;
  assign n18495 = n15900 & n15909 ;
  assign n18496 = ~n16258 & ~n18495 ;
  assign n18497 = n18494 & n18496 ;
  assign n18498 = ~n16305 & ~n16314 ;
  assign n18499 = n16323 & ~n16333 ;
  assign n18500 = ~n16332 & ~n18499 ;
  assign n18501 = n18498 & ~n18500 ;
  assign n18502 = ~n16305 & n16313 ;
  assign n18503 = ~n16304 & ~n18502 ;
  assign n18504 = ~n18501 & n18503 ;
  assign n18505 = ~n16324 & ~n16333 ;
  assign n18506 = n18498 & n18505 ;
  assign n18507 = n16179 & n16188 ;
  assign n18508 = ~n16264 & ~n18507 ;
  assign n18509 = n16267 & ~n16279 ;
  assign n18510 = ~n16280 & ~n18509 ;
  assign n18511 = n18508 & ~n18510 ;
  assign n18512 = ~n16179 & ~n16188 ;
  assign n18513 = n16263 & ~n18507 ;
  assign n18514 = ~n18512 & ~n18513 ;
  assign n18515 = ~n18511 & n18514 ;
  assign n18516 = ~n16268 & ~n16279 ;
  assign n18517 = n18508 & n18516 ;
  assign n18518 = ~n16138 & ~n16147 ;
  assign n18519 = ~n16290 & ~n18518 ;
  assign n18520 = ~n16270 & ~n16291 ;
  assign n18521 = ~n16284 & n18520 ;
  assign n18522 = ~n18519 & n18521 ;
  assign n18523 = n16271 & ~n16284 ;
  assign n18524 = ~n16283 & ~n18523 ;
  assign n18525 = ~n18522 & n18524 ;
  assign n18526 = n16138 & n16147 ;
  assign n18527 = n16122 & n16131 ;
  assign n18528 = ~n16122 & ~n16131 ;
  assign n18529 = n16052 & n16061 ;
  assign n18530 = ~n16052 & ~n16061 ;
  assign n18531 = n16071 & n16074 ;
  assign n18532 = ~n16071 & ~n16074 ;
  assign n18533 = n16083 & n16086 ;
  assign n18534 = ~n16083 & ~n16086 ;
  assign n18535 = n16095 & n16098 ;
  assign n18536 = ~n16095 & ~n16098 ;
  assign n18537 = ~n16103 & ~n16110 ;
  assign n18538 = ~n18536 & ~n18537 ;
  assign n18539 = ~n18535 & ~n18538 ;
  assign n18540 = ~n18534 & ~n18539 ;
  assign n18541 = ~n18533 & ~n18540 ;
  assign n18542 = ~n18532 & ~n18541 ;
  assign n18543 = ~n18531 & ~n18542 ;
  assign n18544 = ~n18530 & ~n18543 ;
  assign n18545 = ~n18529 & ~n18544 ;
  assign n18546 = ~n16295 & ~n18545 ;
  assign n18547 = ~n16294 & ~n18546 ;
  assign n18548 = ~n18528 & ~n18547 ;
  assign n18549 = ~n18527 & ~n18548 ;
  assign n18550 = ~n18526 & n18549 ;
  assign n18551 = n18521 & n18550 ;
  assign n18552 = n18525 & ~n18551 ;
  assign n18553 = n18517 & ~n18552 ;
  assign n18554 = n18515 & ~n18553 ;
  assign n18555 = n18506 & ~n18554 ;
  assign n18556 = n18504 & ~n18555 ;
  assign n18557 = n18497 & ~n18556 ;
  assign n18558 = ~n15900 & ~n15909 ;
  assign n18559 = ~n16258 & n18558 ;
  assign n18560 = ~n16257 & ~n18559 ;
  assign n18561 = n18494 & ~n18560 ;
  assign n18562 = n16273 & ~n16321 ;
  assign n18563 = ~n16320 & ~n18562 ;
  assign n18564 = ~n18561 & n18563 ;
  assign n18565 = ~n18557 & n18564 ;
  assign n18566 = ~n16308 & ~n18565 ;
  assign n18567 = n18493 & ~n18566 ;
  assign n18568 = n18492 & ~n18567 ;
  assign n18569 = n16260 & ~n16329 ;
  assign n18570 = ~n16330 & ~n18569 ;
  assign n18571 = ~n18568 & n18570 ;
  assign n18573 = ~n16319 & n18571 ;
  assign n18489 = ~n16425 & n18488 ;
  assign n18490 = ~n15734 & n18489 ;
  assign n18572 = n16319 & ~n18571 ;
  assign n18574 = n18490 & ~n18572 ;
  assign n18575 = ~n18573 & n18574 ;
  assign n18485 = \P4_IR_reg[20]/NET0131  & ~\P4_IR_reg[21]/NET0131  ;
  assign n18486 = ~\P4_IR_reg[22]/NET0131  & n18485 ;
  assign n18487 = n15798 & n18486 ;
  assign n18576 = n16098 & n16103 ;
  assign n18577 = n16086 & n18576 ;
  assign n18578 = n16074 & n18577 ;
  assign n18579 = n16052 & n18578 ;
  assign n18580 = n16039 & n18579 ;
  assign n18581 = n16122 & n18580 ;
  assign n18582 = n16138 & n18581 ;
  assign n18583 = n16026 & n18582 ;
  assign n18584 = n16012 & n18583 ;
  assign n18585 = n15997 & n18584 ;
  assign n18586 = n15982 & n18585 ;
  assign n18587 = n15967 & n18586 ;
  assign n18588 = n15954 & n18587 ;
  assign n18589 = n16179 & n18588 ;
  assign n18590 = n16165 & n18589 ;
  assign n18591 = n15940 & n18590 ;
  assign n18592 = n15927 & n18591 ;
  assign n18593 = n15913 & n18592 ;
  assign n18594 = n15900 & n18593 ;
  assign n18595 = ~n15886 & n18594 ;
  assign n18596 = ~n15875 & n18595 ;
  assign n18597 = ~n15858 & n18596 ;
  assign n18598 = ~n15847 & n18597 ;
  assign n18599 = ~n15834 & n18598 ;
  assign n18600 = ~n15823 & n18599 ;
  assign n18601 = ~n15811 & n18600 ;
  assign n18603 = ~n15798 & n18601 ;
  assign n18602 = n15798 & ~n18601 ;
  assign n18604 = n15738 & n16425 ;
  assign n18605 = ~n18602 & n18604 ;
  assign n18606 = ~n18603 & n18605 ;
  assign n18645 = ~n18487 & ~n18606 ;
  assign n18646 = ~n18575 & n18645 ;
  assign n18647 = ~n18644 & n18646 ;
  assign n18648 = ~n18484 & n18647 ;
  assign n18650 = ~\P4_IR_reg[25]/NET0131  & \P4_IR_reg[26]/NET0131  ;
  assign n18653 = ~\P4_B_reg/NET0131  & \P4_IR_reg[24]/NET0131  ;
  assign n18654 = n18650 & n18653 ;
  assign n18651 = \P4_B_reg/NET0131  & ~\P4_IR_reg[24]/NET0131  ;
  assign n18652 = n18650 & n18651 ;
  assign n18649 = \P4_IR_reg[26]/NET0131  & \P4_d_reg[0]/NET0131  ;
  assign n18655 = \P4_IR_reg[24]/NET0131  & ~\P4_IR_reg[26]/NET0131  ;
  assign n18656 = ~n18649 & ~n18655 ;
  assign n18657 = ~n18652 & n18656 ;
  assign n18658 = ~n18654 & n18657 ;
  assign n18659 = \P4_IR_reg[26]/NET0131  & \P4_d_reg[1]/NET0131  ;
  assign n18660 = \P4_IR_reg[25]/NET0131  & ~\P4_IR_reg[26]/NET0131  ;
  assign n18661 = ~n18659 & ~n18660 ;
  assign n18662 = ~n18652 & n18661 ;
  assign n18663 = ~n18654 & n18662 ;
  assign n18664 = ~n18658 & n18663 ;
  assign n18665 = \P3_rd_reg/NET0131  & ~\P4_IR_reg[23]/NET0131  ;
  assign n18666 = ~n15736 & n18665 ;
  assign n18667 = n18664 & n18666 ;
  assign n18668 = ~n18648 & n18667 ;
  assign n18669 = ~n16254 & n16425 ;
  assign n18670 = ~n18483 & ~n18669 ;
  assign n18671 = ~n18664 & ~n18670 ;
  assign n18672 = ~n18490 & ~n18607 ;
  assign n18673 = ~n18664 & ~n18672 ;
  assign n18674 = ~\P4_IR_reg[20]/NET0131  & n16425 ;
  assign n18675 = ~n15734 & ~n18674 ;
  assign n18676 = ~n15738 & ~n18675 ;
  assign n18677 = n18666 & ~n18676 ;
  assign n18678 = ~n18673 & n18677 ;
  assign n18679 = ~n18671 & n18678 ;
  assign n18680 = \P4_reg1_reg[27]/NET0131  & ~n18679 ;
  assign n18681 = ~n18668 & ~n18680 ;
  assign n18682 = \P4_reg1_reg[28]/NET0131  & ~n18679 ;
  assign n18683 = ~n16308 & ~n16321 ;
  assign n18684 = n18519 & ~n18550 ;
  assign n18685 = ~n16291 & ~n18684 ;
  assign n18686 = ~n16270 & n18685 ;
  assign n18687 = ~n16271 & ~n18686 ;
  assign n18688 = ~n16283 & n18687 ;
  assign n18689 = ~n16268 & ~n16284 ;
  assign n18690 = ~n18688 & n18689 ;
  assign n18691 = ~n16267 & ~n18690 ;
  assign n18692 = ~n16279 & ~n18691 ;
  assign n18693 = ~n16263 & ~n16280 ;
  assign n18694 = ~n18692 & n18693 ;
  assign n18695 = n18508 & ~n18694 ;
  assign n18696 = ~n16323 & ~n18512 ;
  assign n18697 = ~n18695 & n18696 ;
  assign n18698 = n18505 & ~n18697 ;
  assign n18699 = ~n16313 & ~n16332 ;
  assign n18700 = ~n18698 & n18699 ;
  assign n18701 = ~n18495 & n18498 ;
  assign n18702 = ~n18700 & n18701 ;
  assign n18703 = ~n16304 & ~n18558 ;
  assign n18704 = ~n18495 & ~n18703 ;
  assign n18705 = ~n18702 & ~n18704 ;
  assign n18706 = ~n16258 & ~n16274 ;
  assign n18707 = ~n18705 & n18706 ;
  assign n18708 = n18683 & n18707 ;
  assign n18709 = n16257 & ~n16274 ;
  assign n18710 = ~n16273 & ~n18709 ;
  assign n18711 = n18683 & ~n18710 ;
  assign n18712 = ~n16308 & n16320 ;
  assign n18713 = ~n16307 & ~n18712 ;
  assign n18714 = ~n18711 & n18713 ;
  assign n18715 = ~n18708 & n18714 ;
  assign n18716 = ~n16318 & n18492 ;
  assign n18717 = ~n18715 & n18716 ;
  assign n18718 = ~n16261 & n16276 ;
  assign n18719 = ~n16260 & ~n18718 ;
  assign n18720 = ~n16329 & ~n18719 ;
  assign n18721 = ~n16317 & ~n16330 ;
  assign n18722 = ~n18720 & n18721 ;
  assign n18723 = ~n16318 & ~n18722 ;
  assign n18724 = ~n18717 & ~n18723 ;
  assign n18726 = n16312 & ~n18724 ;
  assign n18725 = ~n16312 & n18724 ;
  assign n18727 = n18490 & ~n18725 ;
  assign n18728 = ~n18726 & n18727 ;
  assign n18735 = ~n16235 & ~n16312 ;
  assign n18734 = n16235 & n16312 ;
  assign n18736 = n18607 & ~n18734 ;
  assign n18737 = ~n18735 & n18736 ;
  assign n18729 = n15785 & n18486 ;
  assign n18731 = n15785 & ~n18603 ;
  assign n18730 = ~n15785 & n18603 ;
  assign n18732 = n18604 & ~n18730 ;
  assign n18733 = ~n18731 & n18732 ;
  assign n18738 = ~n18729 & ~n18733 ;
  assign n18739 = ~n18737 & n18738 ;
  assign n18740 = ~n18728 & n18739 ;
  assign n18741 = n15782 & ~n18478 ;
  assign n18742 = ~n15782 & ~n15794 ;
  assign n18743 = n18476 & n18742 ;
  assign n18744 = ~n18741 & ~n18743 ;
  assign n18745 = ~\P4_IR_reg[28]/NET0131  & ~n18744 ;
  assign n18746 = \P4_IR_reg[28]/NET0131  & n15809 ;
  assign n18747 = ~n18745 & ~n18746 ;
  assign n18748 = n18483 & n18747 ;
  assign n18749 = n18740 & ~n18748 ;
  assign n18750 = n18667 & ~n18749 ;
  assign n18751 = ~n18682 & ~n18750 ;
  assign n18752 = \P1_P3_EAX_reg[16]/NET0131  & ~n16968 ;
  assign n18753 = \P1_P3_EAX_reg[15]/NET0131  & n17166 ;
  assign n18754 = n16982 & ~n18753 ;
  assign n18755 = n16988 & ~n18754 ;
  assign n18756 = \P1_P3_EAX_reg[16]/NET0131  & ~n18755 ;
  assign n18757 = ~\P1_P3_EAX_reg[16]/NET0131  & n16982 ;
  assign n18758 = n18753 & n18757 ;
  assign n18763 = \P1_P3_InstQueue_reg[4][0]/NET0131  & n8777 ;
  assign n18764 = \P1_P3_InstQueue_reg[9][0]/NET0131  & n8754 ;
  assign n18777 = ~n18763 & ~n18764 ;
  assign n18765 = \P1_P3_InstQueue_reg[0][0]/NET0131  & n8775 ;
  assign n18766 = \P1_P3_InstQueue_reg[6][0]/NET0131  & n8771 ;
  assign n18778 = ~n18765 & ~n18766 ;
  assign n18785 = n18777 & n18778 ;
  assign n18759 = \P1_P3_InstQueue_reg[15][0]/NET0131  & n8760 ;
  assign n18760 = \P1_P3_InstQueue_reg[10][0]/NET0131  & n8748 ;
  assign n18775 = ~n18759 & ~n18760 ;
  assign n18761 = \P1_P3_InstQueue_reg[13][0]/NET0131  & n8757 ;
  assign n18762 = \P1_P3_InstQueue_reg[8][0]/NET0131  & n8779 ;
  assign n18776 = ~n18761 & ~n18762 ;
  assign n18786 = n18775 & n18776 ;
  assign n18787 = n18785 & n18786 ;
  assign n18771 = \P1_P3_InstQueue_reg[5][0]/NET0131  & n8752 ;
  assign n18772 = \P1_P3_InstQueue_reg[7][0]/NET0131  & n8745 ;
  assign n18781 = ~n18771 & ~n18772 ;
  assign n18773 = \P1_P3_InstQueue_reg[11][0]/NET0131  & n8769 ;
  assign n18774 = \P1_P3_InstQueue_reg[1][0]/NET0131  & n8781 ;
  assign n18782 = ~n18773 & ~n18774 ;
  assign n18783 = n18781 & n18782 ;
  assign n18767 = \P1_P3_InstQueue_reg[12][0]/NET0131  & n8763 ;
  assign n18768 = \P1_P3_InstQueue_reg[3][0]/NET0131  & n8767 ;
  assign n18779 = ~n18767 & ~n18768 ;
  assign n18769 = \P1_P3_InstQueue_reg[14][0]/NET0131  & n8765 ;
  assign n18770 = \P1_P3_InstQueue_reg[2][0]/NET0131  & n8773 ;
  assign n18780 = ~n18769 & ~n18770 ;
  assign n18784 = n18779 & n18780 ;
  assign n18788 = n18783 & n18784 ;
  assign n18789 = n18787 & n18788 ;
  assign n18790 = n16984 & ~n18789 ;
  assign n18791 = \P1_buf2_reg[0]/NET0131  & n9085 ;
  assign n18792 = \P1_buf2_reg[16]/NET0131  & n9086 ;
  assign n18793 = ~n18791 & ~n18792 ;
  assign n18794 = n9088 & ~n18793 ;
  assign n18795 = ~n18790 & ~n18794 ;
  assign n18796 = ~n18758 & n18795 ;
  assign n18797 = ~n18756 & n18796 ;
  assign n18798 = n9241 & ~n18797 ;
  assign n18799 = ~n18752 & ~n18798 ;
  assign n18800 = \P1_P3_EAX_reg[1]/NET0131  & ~n17031 ;
  assign n18802 = \P1_buf2_reg[1]/NET0131  & n9088 ;
  assign n18803 = ~n9087 & n18802 ;
  assign n18801 = n16984 & ~n18375 ;
  assign n18804 = ~\P1_P3_EAX_reg[0]/NET0131  & ~\P1_P3_EAX_reg[1]/NET0131  ;
  assign n18805 = ~n16972 & ~n18804 ;
  assign n18806 = n16982 & n18805 ;
  assign n18807 = ~n18801 & ~n18806 ;
  assign n18808 = ~n18803 & n18807 ;
  assign n18809 = n9241 & ~n18808 ;
  assign n18810 = ~n18800 & ~n18809 ;
  assign n18811 = \P1_P3_EAX_reg[18]/NET0131  & ~n16968 ;
  assign n18812 = \P1_P3_EAX_reg[16]/NET0131  & n18753 ;
  assign n18813 = \P1_P3_EAX_reg[17]/NET0131  & n18812 ;
  assign n18814 = n16982 & ~n18813 ;
  assign n18815 = n16988 & ~n18814 ;
  assign n18816 = \P1_P3_EAX_reg[18]/NET0131  & ~n18815 ;
  assign n18817 = ~\P1_P3_EAX_reg[18]/NET0131  & n16982 ;
  assign n18818 = n18813 & n18817 ;
  assign n18823 = \P1_P3_InstQueue_reg[6][2]/NET0131  & n8771 ;
  assign n18824 = \P1_P3_InstQueue_reg[14][2]/NET0131  & n8765 ;
  assign n18837 = ~n18823 & ~n18824 ;
  assign n18825 = \P1_P3_InstQueue_reg[11][2]/NET0131  & n8769 ;
  assign n18826 = \P1_P3_InstQueue_reg[5][2]/NET0131  & n8752 ;
  assign n18838 = ~n18825 & ~n18826 ;
  assign n18845 = n18837 & n18838 ;
  assign n18819 = \P1_P3_InstQueue_reg[4][2]/NET0131  & n8777 ;
  assign n18820 = \P1_P3_InstQueue_reg[10][2]/NET0131  & n8748 ;
  assign n18835 = ~n18819 & ~n18820 ;
  assign n18821 = \P1_P3_InstQueue_reg[0][2]/NET0131  & n8775 ;
  assign n18822 = \P1_P3_InstQueue_reg[8][2]/NET0131  & n8779 ;
  assign n18836 = ~n18821 & ~n18822 ;
  assign n18846 = n18835 & n18836 ;
  assign n18847 = n18845 & n18846 ;
  assign n18831 = \P1_P3_InstQueue_reg[13][2]/NET0131  & n8757 ;
  assign n18832 = \P1_P3_InstQueue_reg[12][2]/NET0131  & n8763 ;
  assign n18841 = ~n18831 & ~n18832 ;
  assign n18833 = \P1_P3_InstQueue_reg[7][2]/NET0131  & n8745 ;
  assign n18834 = \P1_P3_InstQueue_reg[1][2]/NET0131  & n8781 ;
  assign n18842 = ~n18833 & ~n18834 ;
  assign n18843 = n18841 & n18842 ;
  assign n18827 = \P1_P3_InstQueue_reg[15][2]/NET0131  & n8760 ;
  assign n18828 = \P1_P3_InstQueue_reg[3][2]/NET0131  & n8767 ;
  assign n18839 = ~n18827 & ~n18828 ;
  assign n18829 = \P1_P3_InstQueue_reg[9][2]/NET0131  & n8754 ;
  assign n18830 = \P1_P3_InstQueue_reg[2][2]/NET0131  & n8773 ;
  assign n18840 = ~n18829 & ~n18830 ;
  assign n18844 = n18839 & n18840 ;
  assign n18848 = n18843 & n18844 ;
  assign n18849 = n18847 & n18848 ;
  assign n18850 = n16984 & ~n18849 ;
  assign n18851 = \P1_buf2_reg[2]/NET0131  & n9085 ;
  assign n18852 = \P1_buf2_reg[18]/NET0131  & n9086 ;
  assign n18853 = ~n18851 & ~n18852 ;
  assign n18854 = n9088 & ~n18853 ;
  assign n18855 = ~n18850 & ~n18854 ;
  assign n18856 = ~n18818 & n18855 ;
  assign n18857 = ~n18816 & n18856 ;
  assign n18858 = n9241 & ~n18857 ;
  assign n18859 = ~n18811 & ~n18858 ;
  assign n18860 = \P1_P3_EAX_reg[2]/NET0131  & ~n17031 ;
  assign n18893 = \P1_buf2_reg[2]/NET0131  & n9175 ;
  assign n18865 = \P1_P3_InstQueue_reg[12][2]/NET0131  & n8765 ;
  assign n18866 = \P1_P3_InstQueue_reg[6][2]/NET0131  & n8779 ;
  assign n18879 = ~n18865 & ~n18866 ;
  assign n18867 = \P1_P3_InstQueue_reg[7][2]/NET0131  & n8754 ;
  assign n18868 = \P1_P3_InstQueue_reg[2][2]/NET0131  & n8777 ;
  assign n18880 = ~n18867 & ~n18868 ;
  assign n18887 = n18879 & n18880 ;
  assign n18861 = \P1_P3_InstQueue_reg[5][2]/NET0131  & n8745 ;
  assign n18862 = \P1_P3_InstQueue_reg[13][2]/NET0131  & n8760 ;
  assign n18877 = ~n18861 & ~n18862 ;
  assign n18863 = \P1_P3_InstQueue_reg[8][2]/NET0131  & n8748 ;
  assign n18864 = \P1_P3_InstQueue_reg[14][2]/NET0131  & n8775 ;
  assign n18878 = ~n18863 & ~n18864 ;
  assign n18888 = n18877 & n18878 ;
  assign n18889 = n18887 & n18888 ;
  assign n18873 = \P1_P3_InstQueue_reg[9][2]/NET0131  & n8769 ;
  assign n18874 = \P1_P3_InstQueue_reg[3][2]/NET0131  & n8752 ;
  assign n18883 = ~n18873 & ~n18874 ;
  assign n18875 = \P1_P3_InstQueue_reg[1][2]/NET0131  & n8767 ;
  assign n18876 = \P1_P3_InstQueue_reg[10][2]/NET0131  & n8763 ;
  assign n18884 = ~n18875 & ~n18876 ;
  assign n18885 = n18883 & n18884 ;
  assign n18869 = \P1_P3_InstQueue_reg[11][2]/NET0131  & n8757 ;
  assign n18870 = \P1_P3_InstQueue_reg[0][2]/NET0131  & n8773 ;
  assign n18881 = ~n18869 & ~n18870 ;
  assign n18871 = \P1_P3_InstQueue_reg[4][2]/NET0131  & n8771 ;
  assign n18872 = \P1_P3_InstQueue_reg[15][2]/NET0131  & n8781 ;
  assign n18882 = ~n18871 & ~n18872 ;
  assign n18886 = n18881 & n18882 ;
  assign n18890 = n18885 & n18886 ;
  assign n18891 = n18889 & n18890 ;
  assign n18892 = n16984 & ~n18891 ;
  assign n18894 = ~\P1_P3_EAX_reg[2]/NET0131  & ~n16972 ;
  assign n18895 = ~n16973 & ~n18894 ;
  assign n18896 = n16982 & n18895 ;
  assign n18897 = ~n18892 & ~n18896 ;
  assign n18898 = ~n18893 & n18897 ;
  assign n18899 = n9241 & ~n18898 ;
  assign n18900 = ~n18860 & ~n18899 ;
  assign n18901 = \P1_P3_EAX_reg[3]/NET0131  & ~n17031 ;
  assign n18934 = \P1_buf2_reg[3]/NET0131  & n9175 ;
  assign n18906 = \P1_P3_InstQueue_reg[14][3]/NET0131  & n8775 ;
  assign n18907 = \P1_P3_InstQueue_reg[7][3]/NET0131  & n8754 ;
  assign n18920 = ~n18906 & ~n18907 ;
  assign n18908 = \P1_P3_InstQueue_reg[13][3]/NET0131  & n8760 ;
  assign n18909 = \P1_P3_InstQueue_reg[12][3]/NET0131  & n8765 ;
  assign n18921 = ~n18908 & ~n18909 ;
  assign n18928 = n18920 & n18921 ;
  assign n18902 = \P1_P3_InstQueue_reg[11][3]/NET0131  & n8757 ;
  assign n18903 = \P1_P3_InstQueue_reg[8][3]/NET0131  & n8748 ;
  assign n18918 = ~n18902 & ~n18903 ;
  assign n18904 = \P1_P3_InstQueue_reg[2][3]/NET0131  & n8777 ;
  assign n18905 = \P1_P3_InstQueue_reg[5][3]/NET0131  & n8745 ;
  assign n18919 = ~n18904 & ~n18905 ;
  assign n18929 = n18918 & n18919 ;
  assign n18930 = n18928 & n18929 ;
  assign n18914 = \P1_P3_InstQueue_reg[3][3]/NET0131  & n8752 ;
  assign n18915 = \P1_P3_InstQueue_reg[1][3]/NET0131  & n8767 ;
  assign n18924 = ~n18914 & ~n18915 ;
  assign n18916 = \P1_P3_InstQueue_reg[10][3]/NET0131  & n8763 ;
  assign n18917 = \P1_P3_InstQueue_reg[15][3]/NET0131  & n8781 ;
  assign n18925 = ~n18916 & ~n18917 ;
  assign n18926 = n18924 & n18925 ;
  assign n18910 = \P1_P3_InstQueue_reg[6][3]/NET0131  & n8779 ;
  assign n18911 = \P1_P3_InstQueue_reg[9][3]/NET0131  & n8769 ;
  assign n18922 = ~n18910 & ~n18911 ;
  assign n18912 = \P1_P3_InstQueue_reg[4][3]/NET0131  & n8771 ;
  assign n18913 = \P1_P3_InstQueue_reg[0][3]/NET0131  & n8773 ;
  assign n18923 = ~n18912 & ~n18913 ;
  assign n18927 = n18922 & n18923 ;
  assign n18931 = n18926 & n18927 ;
  assign n18932 = n18930 & n18931 ;
  assign n18933 = n16984 & ~n18932 ;
  assign n18935 = ~\P1_P3_EAX_reg[3]/NET0131  & ~n16973 ;
  assign n18936 = ~n16974 & ~n18935 ;
  assign n18937 = n16982 & n18936 ;
  assign n18938 = ~n18933 & ~n18937 ;
  assign n18939 = ~n18934 & n18938 ;
  assign n18940 = n9241 & ~n18939 ;
  assign n18941 = ~n18901 & ~n18940 ;
  assign n18942 = \P1_P3_EAX_reg[4]/NET0131  & ~n17031 ;
  assign n18975 = \P1_buf2_reg[4]/NET0131  & n9175 ;
  assign n18947 = \P1_P3_InstQueue_reg[14][4]/NET0131  & n8775 ;
  assign n18948 = \P1_P3_InstQueue_reg[7][4]/NET0131  & n8754 ;
  assign n18961 = ~n18947 & ~n18948 ;
  assign n18949 = \P1_P3_InstQueue_reg[13][4]/NET0131  & n8760 ;
  assign n18950 = \P1_P3_InstQueue_reg[12][4]/NET0131  & n8765 ;
  assign n18962 = ~n18949 & ~n18950 ;
  assign n18969 = n18961 & n18962 ;
  assign n18943 = \P1_P3_InstQueue_reg[11][4]/NET0131  & n8757 ;
  assign n18944 = \P1_P3_InstQueue_reg[8][4]/NET0131  & n8748 ;
  assign n18959 = ~n18943 & ~n18944 ;
  assign n18945 = \P1_P3_InstQueue_reg[2][4]/NET0131  & n8777 ;
  assign n18946 = \P1_P3_InstQueue_reg[5][4]/NET0131  & n8745 ;
  assign n18960 = ~n18945 & ~n18946 ;
  assign n18970 = n18959 & n18960 ;
  assign n18971 = n18969 & n18970 ;
  assign n18955 = \P1_P3_InstQueue_reg[3][4]/NET0131  & n8752 ;
  assign n18956 = \P1_P3_InstQueue_reg[1][4]/NET0131  & n8767 ;
  assign n18965 = ~n18955 & ~n18956 ;
  assign n18957 = \P1_P3_InstQueue_reg[10][4]/NET0131  & n8763 ;
  assign n18958 = \P1_P3_InstQueue_reg[15][4]/NET0131  & n8781 ;
  assign n18966 = ~n18957 & ~n18958 ;
  assign n18967 = n18965 & n18966 ;
  assign n18951 = \P1_P3_InstQueue_reg[6][4]/NET0131  & n8779 ;
  assign n18952 = \P1_P3_InstQueue_reg[9][4]/NET0131  & n8769 ;
  assign n18963 = ~n18951 & ~n18952 ;
  assign n18953 = \P1_P3_InstQueue_reg[4][4]/NET0131  & n8771 ;
  assign n18954 = \P1_P3_InstQueue_reg[0][4]/NET0131  & n8773 ;
  assign n18964 = ~n18953 & ~n18954 ;
  assign n18968 = n18963 & n18964 ;
  assign n18972 = n18967 & n18968 ;
  assign n18973 = n18971 & n18972 ;
  assign n18974 = n16984 & ~n18973 ;
  assign n18976 = ~\P1_P3_EAX_reg[4]/NET0131  & ~n16974 ;
  assign n18977 = ~n16975 & ~n18976 ;
  assign n18978 = n16982 & n18977 ;
  assign n18979 = ~n18974 & ~n18978 ;
  assign n18980 = ~n18975 & n18979 ;
  assign n18981 = n9241 & ~n18980 ;
  assign n18982 = ~n18942 & ~n18981 ;
  assign n18983 = \P1_P3_EAX_reg[5]/NET0131  & ~n16968 ;
  assign n18985 = ~n16976 & n16982 ;
  assign n18986 = n16988 & ~n18985 ;
  assign n18987 = \P1_P3_EAX_reg[5]/NET0131  & ~n18986 ;
  assign n18984 = \P1_buf2_reg[5]/NET0131  & n9175 ;
  assign n18992 = \P1_P3_InstQueue_reg[6][5]/NET0131  & n8779 ;
  assign n18993 = \P1_P3_InstQueue_reg[13][5]/NET0131  & n8760 ;
  assign n19006 = ~n18992 & ~n18993 ;
  assign n18994 = \P1_P3_InstQueue_reg[5][5]/NET0131  & n8745 ;
  assign n18995 = \P1_P3_InstQueue_reg[4][5]/NET0131  & n8771 ;
  assign n19007 = ~n18994 & ~n18995 ;
  assign n19014 = n19006 & n19007 ;
  assign n18988 = \P1_P3_InstQueue_reg[11][5]/NET0131  & n8757 ;
  assign n18989 = \P1_P3_InstQueue_reg[8][5]/NET0131  & n8748 ;
  assign n19004 = ~n18988 & ~n18989 ;
  assign n18990 = \P1_P3_InstQueue_reg[2][5]/NET0131  & n8777 ;
  assign n18991 = \P1_P3_InstQueue_reg[12][5]/NET0131  & n8765 ;
  assign n19005 = ~n18990 & ~n18991 ;
  assign n19015 = n19004 & n19005 ;
  assign n19016 = n19014 & n19015 ;
  assign n19000 = \P1_P3_InstQueue_reg[9][5]/NET0131  & n8769 ;
  assign n19001 = \P1_P3_InstQueue_reg[14][5]/NET0131  & n8775 ;
  assign n19010 = ~n19000 & ~n19001 ;
  assign n19002 = \P1_P3_InstQueue_reg[1][5]/NET0131  & n8767 ;
  assign n19003 = \P1_P3_InstQueue_reg[15][5]/NET0131  & n8781 ;
  assign n19011 = ~n19002 & ~n19003 ;
  assign n19012 = n19010 & n19011 ;
  assign n18996 = \P1_P3_InstQueue_reg[7][5]/NET0131  & n8754 ;
  assign n18997 = \P1_P3_InstQueue_reg[3][5]/NET0131  & n8752 ;
  assign n19008 = ~n18996 & ~n18997 ;
  assign n18998 = \P1_P3_InstQueue_reg[10][5]/NET0131  & n8763 ;
  assign n18999 = \P1_P3_InstQueue_reg[0][5]/NET0131  & n8773 ;
  assign n19009 = ~n18998 & ~n18999 ;
  assign n19013 = n19008 & n19009 ;
  assign n19017 = n19012 & n19013 ;
  assign n19018 = n19016 & n19017 ;
  assign n19019 = n16984 & ~n19018 ;
  assign n19020 = n16975 & n18985 ;
  assign n19021 = ~n19019 & ~n19020 ;
  assign n19022 = ~n18984 & n19021 ;
  assign n19023 = ~n18987 & n19022 ;
  assign n19024 = n9241 & ~n19023 ;
  assign n19025 = ~n18983 & ~n19024 ;
  assign n19026 = \P1_P3_EAX_reg[6]/NET0131  & ~n16968 ;
  assign n19027 = ~n16987 & ~n18985 ;
  assign n19028 = \P1_P3_EAX_reg[6]/NET0131  & ~n19027 ;
  assign n19064 = ~\P1_buf2_reg[6]/NET0131  & n9088 ;
  assign n19063 = ~\P1_P3_EAX_reg[6]/NET0131  & ~n9088 ;
  assign n19065 = ~n9087 & ~n19063 ;
  assign n19066 = ~n19064 & n19065 ;
  assign n19029 = ~\P1_P3_EAX_reg[6]/NET0131  & n16976 ;
  assign n19030 = n16982 & n19029 ;
  assign n19035 = \P1_P3_InstQueue_reg[14][6]/NET0131  & n8775 ;
  assign n19036 = \P1_P3_InstQueue_reg[7][6]/NET0131  & n8754 ;
  assign n19049 = ~n19035 & ~n19036 ;
  assign n19037 = \P1_P3_InstQueue_reg[13][6]/NET0131  & n8760 ;
  assign n19038 = \P1_P3_InstQueue_reg[12][6]/NET0131  & n8765 ;
  assign n19050 = ~n19037 & ~n19038 ;
  assign n19057 = n19049 & n19050 ;
  assign n19031 = \P1_P3_InstQueue_reg[11][6]/NET0131  & n8757 ;
  assign n19032 = \P1_P3_InstQueue_reg[8][6]/NET0131  & n8748 ;
  assign n19047 = ~n19031 & ~n19032 ;
  assign n19033 = \P1_P3_InstQueue_reg[2][6]/NET0131  & n8777 ;
  assign n19034 = \P1_P3_InstQueue_reg[5][6]/NET0131  & n8745 ;
  assign n19048 = ~n19033 & ~n19034 ;
  assign n19058 = n19047 & n19048 ;
  assign n19059 = n19057 & n19058 ;
  assign n19043 = \P1_P3_InstQueue_reg[3][6]/NET0131  & n8752 ;
  assign n19044 = \P1_P3_InstQueue_reg[1][6]/NET0131  & n8767 ;
  assign n19053 = ~n19043 & ~n19044 ;
  assign n19045 = \P1_P3_InstQueue_reg[10][6]/NET0131  & n8763 ;
  assign n19046 = \P1_P3_InstQueue_reg[15][6]/NET0131  & n8781 ;
  assign n19054 = ~n19045 & ~n19046 ;
  assign n19055 = n19053 & n19054 ;
  assign n19039 = \P1_P3_InstQueue_reg[6][6]/NET0131  & n8779 ;
  assign n19040 = \P1_P3_InstQueue_reg[9][6]/NET0131  & n8769 ;
  assign n19051 = ~n19039 & ~n19040 ;
  assign n19041 = \P1_P3_InstQueue_reg[4][6]/NET0131  & n8771 ;
  assign n19042 = \P1_P3_InstQueue_reg[0][6]/NET0131  & n8773 ;
  assign n19052 = ~n19041 & ~n19042 ;
  assign n19056 = n19051 & n19052 ;
  assign n19060 = n19055 & n19056 ;
  assign n19061 = n19059 & n19060 ;
  assign n19062 = n16984 & ~n19061 ;
  assign n19067 = ~n19030 & ~n19062 ;
  assign n19068 = ~n19066 & n19067 ;
  assign n19069 = ~n19028 & n19068 ;
  assign n19070 = n9241 & ~n19069 ;
  assign n19071 = ~n19026 & ~n19070 ;
  assign n19073 = ~\P4_IR_reg[23]/NET0131  & n15736 ;
  assign n19074 = n16171 & n19073 ;
  assign n19075 = ~\P4_IR_reg[23]/NET0131  & ~n15736 ;
  assign n19077 = ~n16188 & n18462 ;
  assign n19078 = ~n16175 & n19077 ;
  assign n19079 = n15949 & ~n19078 ;
  assign n19080 = ~n15949 & n19078 ;
  assign n19081 = ~n19079 & ~n19080 ;
  assign n19082 = ~\P4_IR_reg[28]/NET0131  & ~n19081 ;
  assign n19083 = \P4_IR_reg[28]/NET0131  & n16188 ;
  assign n19084 = ~n19082 & ~n19083 ;
  assign n19085 = n18483 & n19084 ;
  assign n19104 = n15734 & ~n15738 ;
  assign n19076 = ~n18658 & ~n18663 ;
  assign n19105 = ~n15734 & ~n16425 ;
  assign n19106 = ~n15738 & ~n19105 ;
  assign n19107 = ~\P4_IR_reg[21]/NET0131  & ~n19105 ;
  assign n19108 = ~n19106 & ~n19107 ;
  assign n19109 = ~n18669 & ~n19108 ;
  assign n19110 = ~n19076 & ~n19109 ;
  assign n19111 = ~n19104 & ~n19110 ;
  assign n19112 = ~n19085 & n19111 ;
  assign n19113 = n16171 & ~n19112 ;
  assign n19095 = ~n16325 & n18554 ;
  assign n19094 = n16325 & ~n18554 ;
  assign n19096 = n18490 & ~n19094 ;
  assign n19097 = ~n19095 & n19096 ;
  assign n19091 = n16325 & n18622 ;
  assign n19090 = ~n16325 & ~n18622 ;
  assign n19092 = n18607 & ~n19090 ;
  assign n19093 = ~n19091 & n19092 ;
  assign n19086 = ~n16165 & n18486 ;
  assign n19087 = ~n16165 & ~n18589 ;
  assign n19088 = ~n18590 & n18604 ;
  assign n19089 = ~n19087 & n19088 ;
  assign n19098 = ~n19086 & ~n19089 ;
  assign n19099 = ~n19093 & n19098 ;
  assign n19100 = ~n19097 & n19099 ;
  assign n19101 = ~n19085 & n19100 ;
  assign n19102 = n19076 & ~n19101 ;
  assign n19103 = ~n16165 & n16426 ;
  assign n19114 = ~n19102 & ~n19103 ;
  assign n19115 = ~n19113 & n19114 ;
  assign n19116 = n19075 & ~n19115 ;
  assign n19117 = ~n19074 & ~n19116 ;
  assign n19118 = \P3_rd_reg/NET0131  & ~n19117 ;
  assign n19072 = ~\P3_rd_reg/NET0131  & \P4_reg3_reg[15]/NET0131  ;
  assign n19119 = n15744 & n16171 ;
  assign n19120 = ~n19072 & ~n19119 ;
  assign n19121 = ~n19118 & n19120 ;
  assign n19123 = ~\P1_P3_PhyAddrPointer_reg[1]/NET0131  & n16914 ;
  assign n19124 = ~n16915 & ~n19123 ;
  assign n19125 = ~\P1_P3_DataWidth_reg[1]/NET0131  & ~n19124 ;
  assign n19126 = \P1_P3_DataWidth_reg[1]/NET0131  & ~\P1_P3_rEIP_reg[1]/NET0131  ;
  assign n19127 = n9245 & ~n19126 ;
  assign n19128 = ~n19125 & n19127 ;
  assign n19130 = \P1_P3_rEIP_reg[1]/NET0131  & ~n9195 ;
  assign n19131 = \P1_P3_EBX_reg[1]/NET0131  & ~\P1_P3_EBX_reg[31]/NET0131  ;
  assign n19132 = \P1_P3_EBX_reg[0]/NET0131  & \P1_P3_EBX_reg[1]/NET0131  ;
  assign n19133 = n16930 & ~n19132 ;
  assign n19134 = ~n19131 & ~n19133 ;
  assign n19135 = ~n16505 & ~n19134 ;
  assign n19136 = ~\P1_P3_rEIP_reg[1]/NET0131  & n16505 ;
  assign n19137 = ~n19135 & ~n19136 ;
  assign n19138 = n9085 & ~n19137 ;
  assign n19139 = n9082 & ~n9207 ;
  assign n19140 = \P1_P3_EBX_reg[1]/NET0131  & ~n16517 ;
  assign n19141 = ~n9095 & n19136 ;
  assign n19142 = ~n19140 & ~n19141 ;
  assign n19143 = n9079 & ~n19142 ;
  assign n19144 = ~n19139 & ~n19143 ;
  assign n19145 = ~n19138 & n19144 ;
  assign n19146 = ~n9075 & ~n19145 ;
  assign n19147 = ~n19130 & ~n19146 ;
  assign n19148 = n9241 & ~n19147 ;
  assign n19122 = \P1_P3_PhyAddrPointer_reg[1]/NET0131  & n10031 ;
  assign n19129 = \P1_P3_rEIP_reg[1]/NET0131  & ~n16495 ;
  assign n19149 = ~n19122 & ~n19129 ;
  assign n19150 = ~n19148 & n19149 ;
  assign n19151 = ~n19128 & n19150 ;
  assign n19152 = ~n18648 & n19076 ;
  assign n19153 = n15798 & n16426 ;
  assign n19154 = ~n19152 & ~n19153 ;
  assign n19155 = n19075 & ~n19154 ;
  assign n19156 = n18489 & ~n19076 ;
  assign n19157 = n19076 & ~n19104 ;
  assign n19158 = n18488 & ~n18669 ;
  assign n19159 = ~n19157 & ~n19158 ;
  assign n19160 = ~n19156 & ~n19159 ;
  assign n19161 = ~n15736 & n19160 ;
  assign n19162 = ~\P4_IR_reg[23]/NET0131  & ~n19161 ;
  assign n19163 = n15805 & n19162 ;
  assign n19164 = ~n19155 & ~n19163 ;
  assign n19165 = \P3_rd_reg/NET0131  & ~n19164 ;
  assign n19166 = ~\P3_rd_reg/NET0131  & \P4_reg3_reg[27]/NET0131  ;
  assign n19167 = n15744 & n15805 ;
  assign n19168 = ~n19166 & ~n19167 ;
  assign n19169 = ~n19165 & n19168 ;
  assign n19170 = ~n18747 & n19076 ;
  assign n19171 = ~n15790 & ~n19076 ;
  assign n19172 = n18483 & ~n19171 ;
  assign n19173 = ~n19170 & n19172 ;
  assign n19174 = ~n18740 & n19076 ;
  assign n19175 = n15785 & n16426 ;
  assign n19176 = ~n15734 & n19156 ;
  assign n19177 = ~n19159 & ~n19176 ;
  assign n19178 = n15790 & ~n19177 ;
  assign n19179 = ~n19175 & ~n19178 ;
  assign n19180 = ~n19174 & n19179 ;
  assign n19181 = ~n19173 & n19180 ;
  assign n19182 = n19075 & ~n19181 ;
  assign n19183 = n15790 & n19073 ;
  assign n19184 = ~n19182 & ~n19183 ;
  assign n19185 = \P3_rd_reg/NET0131  & ~n19184 ;
  assign n19186 = ~\P3_rd_reg/NET0131  & \P4_reg3_reg[28]/NET0131  ;
  assign n19187 = n15744 & n15790 ;
  assign n19188 = ~n19186 & ~n19187 ;
  assign n19189 = ~n19185 & n19188 ;
  assign n19205 = \P1_P3_InstAddrPointer_reg[10]/NET0131  & n9072 ;
  assign n19191 = \P1_P3_InstAddrPointer_reg[1]/NET0131  & \P1_P3_InstAddrPointer_reg[2]/NET0131  ;
  assign n19192 = \P1_P3_InstAddrPointer_reg[3]/NET0131  & n19191 ;
  assign n19193 = \P1_P3_InstAddrPointer_reg[4]/NET0131  & n19192 ;
  assign n19194 = \P1_P3_InstAddrPointer_reg[5]/NET0131  & n19193 ;
  assign n19195 = \P1_P3_InstAddrPointer_reg[6]/NET0131  & n19194 ;
  assign n19258 = \P1_P3_InstAddrPointer_reg[7]/NET0131  & n19195 ;
  assign n19259 = \P1_P3_InstAddrPointer_reg[8]/NET0131  & n19258 ;
  assign n19260 = \P1_P3_InstAddrPointer_reg[9]/NET0131  & n19259 ;
  assign n19261 = ~\P1_P3_InstAddrPointer_reg[10]/NET0131  & ~n19260 ;
  assign n19201 = \P1_P3_InstAddrPointer_reg[10]/NET0131  & \P1_P3_InstAddrPointer_reg[9]/NET0131  ;
  assign n19262 = n19201 & n19259 ;
  assign n19263 = ~n19261 & ~n19262 ;
  assign n19264 = ~\P1_P3_InstAddrPointer_reg[8]/NET0131  & ~n19258 ;
  assign n19265 = ~n19259 & ~n19264 ;
  assign n19266 = ~\P1_P3_InstAddrPointer_reg[7]/NET0131  & ~n19195 ;
  assign n19267 = ~n19258 & ~n19266 ;
  assign n19268 = ~\P1_P3_InstAddrPointer_reg[6]/NET0131  & ~n19194 ;
  assign n19269 = ~n19195 & ~n19268 ;
  assign n19270 = ~n19061 & n19269 ;
  assign n19271 = n19061 & ~n19269 ;
  assign n19272 = ~\P1_P3_InstAddrPointer_reg[5]/NET0131  & ~n19193 ;
  assign n19273 = ~n19194 & ~n19272 ;
  assign n19274 = ~n19018 & n19273 ;
  assign n19275 = n19018 & ~n19273 ;
  assign n19276 = ~\P1_P3_InstAddrPointer_reg[4]/NET0131  & ~n19192 ;
  assign n19277 = ~n19193 & ~n19276 ;
  assign n19278 = n18973 & ~n19277 ;
  assign n19279 = ~\P1_P3_InstAddrPointer_reg[3]/NET0131  & ~n19191 ;
  assign n19280 = ~n19192 & ~n19279 ;
  assign n19281 = n18932 & ~n19280 ;
  assign n19282 = ~n18932 & n19280 ;
  assign n19283 = ~\P1_P3_InstAddrPointer_reg[1]/NET0131  & ~\P1_P3_InstAddrPointer_reg[2]/NET0131  ;
  assign n19284 = ~n19191 & ~n19283 ;
  assign n19285 = n18891 & ~n19284 ;
  assign n19286 = ~n18891 & n19284 ;
  assign n19287 = ~n18412 & ~n18418 ;
  assign n19288 = ~n18413 & ~n19287 ;
  assign n19289 = ~n19286 & ~n19288 ;
  assign n19290 = ~n19285 & ~n19289 ;
  assign n19291 = ~n19282 & ~n19290 ;
  assign n19292 = ~n19281 & ~n19291 ;
  assign n19293 = ~n19278 & n19292 ;
  assign n19294 = ~n18973 & n19277 ;
  assign n19295 = ~n19293 & ~n19294 ;
  assign n19296 = ~n19275 & ~n19295 ;
  assign n19297 = ~n19274 & ~n19296 ;
  assign n19298 = ~n19271 & ~n19297 ;
  assign n19299 = ~n19270 & ~n19298 ;
  assign n19300 = ~n19267 & n19299 ;
  assign n19301 = n19267 & ~n19299 ;
  assign n19302 = n17282 & ~n19301 ;
  assign n19303 = ~n19300 & ~n19302 ;
  assign n19304 = n19265 & n19303 ;
  assign n19305 = \P1_P3_InstAddrPointer_reg[9]/NET0131  & n19304 ;
  assign n19306 = ~n19263 & ~n19305 ;
  assign n19307 = \P1_P3_InstAddrPointer_reg[10]/NET0131  & n19305 ;
  assign n19308 = ~n19306 & ~n19307 ;
  assign n19309 = n17282 & ~n19308 ;
  assign n19196 = \P1_P3_InstAddrPointer_reg[0]/NET0131  & n19195 ;
  assign n19197 = \P1_P3_InstAddrPointer_reg[7]/NET0131  & n19196 ;
  assign n19198 = \P1_P3_InstAddrPointer_reg[8]/NET0131  & n19197 ;
  assign n19199 = \P1_P3_InstAddrPointer_reg[9]/NET0131  & n19198 ;
  assign n19200 = ~\P1_P3_InstAddrPointer_reg[10]/NET0131  & ~n19199 ;
  assign n19202 = n19198 & n19201 ;
  assign n19203 = ~n19200 & ~n19202 ;
  assign n19206 = ~\P1_P3_InstAddrPointer_reg[9]/NET0131  & ~n19198 ;
  assign n19207 = ~n19199 & ~n19206 ;
  assign n19208 = ~\P1_P3_InstAddrPointer_reg[8]/NET0131  & ~n19197 ;
  assign n19209 = ~n19198 & ~n19208 ;
  assign n19210 = ~\P1_P3_InstAddrPointer_reg[7]/NET0131  & ~n19196 ;
  assign n19211 = ~n19197 & ~n19210 ;
  assign n19212 = \P1_P3_InstAddrPointer_reg[0]/NET0131  & n19194 ;
  assign n19213 = ~\P1_P3_InstAddrPointer_reg[6]/NET0131  & ~n19212 ;
  assign n19214 = ~n19196 & ~n19213 ;
  assign n19215 = n19061 & ~n19214 ;
  assign n19216 = ~n19061 & n19214 ;
  assign n19217 = \P1_P3_InstAddrPointer_reg[0]/NET0131  & n19193 ;
  assign n19218 = ~\P1_P3_InstAddrPointer_reg[5]/NET0131  & ~n19217 ;
  assign n19219 = ~n19212 & ~n19218 ;
  assign n19220 = n19018 & ~n19219 ;
  assign n19221 = ~n19018 & n19219 ;
  assign n19222 = \P1_P3_InstAddrPointer_reg[0]/NET0131  & n19192 ;
  assign n19223 = ~\P1_P3_InstAddrPointer_reg[4]/NET0131  & ~n19222 ;
  assign n19224 = ~n19217 & ~n19223 ;
  assign n19225 = n18973 & ~n19224 ;
  assign n19226 = ~n18973 & n19224 ;
  assign n19227 = \P1_P3_InstAddrPointer_reg[2]/NET0131  & n15307 ;
  assign n19228 = ~\P1_P3_InstAddrPointer_reg[3]/NET0131  & ~n19227 ;
  assign n19229 = ~n19222 & ~n19228 ;
  assign n19230 = n18932 & ~n19229 ;
  assign n19231 = ~n18932 & n19229 ;
  assign n19232 = ~\P1_P3_InstAddrPointer_reg[2]/NET0131  & ~n15307 ;
  assign n19233 = ~n19227 & ~n19232 ;
  assign n19234 = n18891 & ~n19233 ;
  assign n19235 = ~n18376 & ~n18423 ;
  assign n19236 = ~n18377 & ~n19235 ;
  assign n19237 = ~n18891 & n19233 ;
  assign n19238 = n19236 & ~n19237 ;
  assign n19239 = ~n19234 & ~n19238 ;
  assign n19240 = ~n19231 & ~n19239 ;
  assign n19241 = ~n19230 & ~n19240 ;
  assign n19242 = ~n19226 & ~n19241 ;
  assign n19243 = ~n19225 & ~n19242 ;
  assign n19244 = ~n19221 & ~n19243 ;
  assign n19245 = ~n19220 & ~n19244 ;
  assign n19246 = ~n19216 & ~n19245 ;
  assign n19247 = ~n19215 & ~n19246 ;
  assign n19248 = n19211 & n19247 ;
  assign n19249 = ~n19211 & ~n19247 ;
  assign n19250 = ~n17282 & ~n19249 ;
  assign n19251 = ~n19248 & ~n19250 ;
  assign n19252 = ~n19209 & n19251 ;
  assign n19253 = ~n19207 & n19252 ;
  assign n19255 = ~n19203 & n19253 ;
  assign n19254 = n19203 & ~n19253 ;
  assign n19256 = ~n17282 & ~n19254 ;
  assign n19257 = ~n19255 & n19256 ;
  assign n19310 = ~n9072 & ~n19257 ;
  assign n19311 = ~n19309 & n19310 ;
  assign n19312 = ~n19205 & ~n19311 ;
  assign n19313 = n9064 & ~n19312 ;
  assign n19314 = \P1_P3_InstAddrPointer_reg[3]/NET0131  & ~n19232 ;
  assign n19315 = \P1_P3_InstAddrPointer_reg[4]/NET0131  & n19314 ;
  assign n19316 = \P1_P3_InstAddrPointer_reg[5]/NET0131  & n19315 ;
  assign n19317 = \P1_P3_InstAddrPointer_reg[6]/NET0131  & n19316 ;
  assign n19318 = \P1_P3_InstAddrPointer_reg[7]/NET0131  & n19317 ;
  assign n19320 = \P1_P3_InstAddrPointer_reg[8]/NET0131  & n19318 ;
  assign n19360 = \P1_P3_InstAddrPointer_reg[9]/NET0131  & n19320 ;
  assign n19361 = ~\P1_P3_InstAddrPointer_reg[10]/NET0131  & ~n19360 ;
  assign n19362 = n19201 & n19320 ;
  assign n19363 = ~n19361 & ~n19362 ;
  assign n19319 = ~\P1_P3_InstAddrPointer_reg[8]/NET0131  & ~n19318 ;
  assign n19321 = ~n19319 & ~n19320 ;
  assign n19322 = ~\P1_P3_InstAddrPointer_reg[7]/NET0131  & ~n19317 ;
  assign n19323 = ~n19318 & ~n19322 ;
  assign n19324 = ~n17282 & n19323 ;
  assign n19325 = n17282 & ~n19323 ;
  assign n19326 = ~\P1_P3_InstAddrPointer_reg[6]/NET0131  & ~n19316 ;
  assign n19327 = ~n19317 & ~n19326 ;
  assign n19328 = ~n19061 & n19327 ;
  assign n19329 = n19061 & ~n19327 ;
  assign n19330 = ~\P1_P3_InstAddrPointer_reg[5]/NET0131  & ~n19315 ;
  assign n19331 = ~n19316 & ~n19330 ;
  assign n19332 = ~n19018 & n19331 ;
  assign n19333 = n19018 & ~n19331 ;
  assign n19334 = ~\P1_P3_InstAddrPointer_reg[4]/NET0131  & ~n19314 ;
  assign n19335 = ~n19315 & ~n19334 ;
  assign n19336 = n18973 & ~n19335 ;
  assign n19337 = ~\P1_P3_InstAddrPointer_reg[3]/NET0131  & n19232 ;
  assign n19338 = ~n19314 & ~n19337 ;
  assign n19339 = ~n18932 & n19338 ;
  assign n19340 = n18932 & ~n19338 ;
  assign n19341 = ~n18891 & ~n19233 ;
  assign n19342 = n18891 & n19233 ;
  assign n19343 = ~n18377 & ~n18410 ;
  assign n19344 = ~n18376 & ~n19343 ;
  assign n19345 = ~n19342 & n19344 ;
  assign n19346 = ~n19341 & ~n19345 ;
  assign n19347 = ~n19340 & ~n19346 ;
  assign n19348 = ~n19339 & ~n19347 ;
  assign n19349 = ~n19336 & ~n19348 ;
  assign n19350 = ~n18973 & n19335 ;
  assign n19351 = ~n19349 & ~n19350 ;
  assign n19352 = ~n19333 & ~n19351 ;
  assign n19353 = ~n19332 & ~n19352 ;
  assign n19354 = ~n19329 & ~n19353 ;
  assign n19355 = ~n19328 & ~n19354 ;
  assign n19356 = ~n19325 & ~n19355 ;
  assign n19357 = ~n19324 & ~n19356 ;
  assign n19358 = n19321 & ~n19357 ;
  assign n19364 = \P1_P3_InstAddrPointer_reg[9]/NET0131  & n19358 ;
  assign n19365 = ~n19363 & ~n19364 ;
  assign n19359 = n19201 & n19358 ;
  assign n19366 = n9191 & ~n19359 ;
  assign n19367 = ~n19365 & n19366 ;
  assign n19368 = ~n8741 & ~n19263 ;
  assign n19369 = ~n9084 & ~n19368 ;
  assign n19370 = n18437 & ~n19369 ;
  assign n19371 = \P1_P3_InstAddrPointer_reg[10]/NET0131  & ~n19370 ;
  assign n19204 = ~n9133 & n19203 ;
  assign n19374 = ~\P1_P3_InstAddrPointer_reg[10]/NET0131  & n8741 ;
  assign n19375 = ~n19368 & ~n19374 ;
  assign n19376 = ~n9166 & n19375 ;
  assign n19372 = n9118 & n19263 ;
  assign n19373 = n9220 & n19363 ;
  assign n19377 = ~n19372 & ~n19373 ;
  assign n19378 = ~n19376 & n19377 ;
  assign n19379 = ~n19204 & n19378 ;
  assign n19380 = ~n19371 & n19379 ;
  assign n19381 = ~n19367 & n19380 ;
  assign n19382 = ~n19313 & n19381 ;
  assign n19383 = n9241 & ~n19382 ;
  assign n19190 = \P1_P3_rEIP_reg[10]/NET0131  & n17426 ;
  assign n19384 = \P1_P3_InstAddrPointer_reg[10]/NET0131  & ~n18343 ;
  assign n19385 = ~n19190 & ~n19384 ;
  assign n19386 = ~n19383 & n19385 ;
  assign n19392 = \P1_P3_InstAddrPointer_reg[11]/NET0131  & n9072 ;
  assign n19397 = ~\P1_P3_InstAddrPointer_reg[11]/NET0131  & ~n19202 ;
  assign n19398 = \P1_P3_InstAddrPointer_reg[11]/NET0131  & n19201 ;
  assign n19399 = n19198 & n19398 ;
  assign n19400 = ~n19397 & ~n19399 ;
  assign n19402 = n19255 & ~n19400 ;
  assign n19401 = ~n19255 & n19400 ;
  assign n19403 = ~n17282 & ~n19401 ;
  assign n19404 = ~n19402 & n19403 ;
  assign n19388 = ~\P1_P3_InstAddrPointer_reg[11]/NET0131  & ~n19262 ;
  assign n19389 = \P1_P3_InstAddrPointer_reg[11]/NET0131  & n19262 ;
  assign n19390 = ~n19388 & ~n19389 ;
  assign n19393 = ~n19307 & ~n19390 ;
  assign n19394 = n19307 & n19390 ;
  assign n19395 = ~n19393 & ~n19394 ;
  assign n19396 = n17282 & ~n19395 ;
  assign n19405 = ~n9072 & ~n19396 ;
  assign n19406 = ~n19404 & n19405 ;
  assign n19407 = ~n19392 & ~n19406 ;
  assign n19408 = n9064 & ~n19407 ;
  assign n19409 = ~\P1_P3_InstAddrPointer_reg[11]/NET0131  & ~n19362 ;
  assign n19410 = \P1_P3_InstAddrPointer_reg[11]/NET0131  & n19362 ;
  assign n19411 = ~n19409 & ~n19410 ;
  assign n19413 = ~n19359 & ~n19411 ;
  assign n19412 = n19359 & n19411 ;
  assign n19414 = n9191 & ~n19412 ;
  assign n19415 = ~n19413 & n19414 ;
  assign n19418 = ~n9167 & n18437 ;
  assign n19419 = \P1_P3_InstAddrPointer_reg[11]/NET0131  & ~n19418 ;
  assign n19417 = ~n9133 & n19400 ;
  assign n19391 = ~n9176 & n19390 ;
  assign n19416 = n9220 & n19411 ;
  assign n19420 = ~n19391 & ~n19416 ;
  assign n19421 = ~n19417 & n19420 ;
  assign n19422 = ~n19419 & n19421 ;
  assign n19423 = ~n19415 & n19422 ;
  assign n19424 = ~n19408 & n19423 ;
  assign n19425 = n9241 & ~n19424 ;
  assign n19387 = \P1_P3_rEIP_reg[11]/NET0131  & n17426 ;
  assign n19426 = \P1_P3_InstAddrPointer_reg[11]/NET0131  & ~n18343 ;
  assign n19427 = ~n19387 & ~n19426 ;
  assign n19428 = ~n19425 & n19427 ;
  assign n19435 = \P1_P3_InstAddrPointer_reg[12]/NET0131  & n19399 ;
  assign n19436 = ~\P1_P3_InstAddrPointer_reg[13]/NET0131  & ~n19435 ;
  assign n19437 = \P1_P3_InstAddrPointer_reg[12]/NET0131  & \P1_P3_InstAddrPointer_reg[13]/NET0131  ;
  assign n19438 = n19399 & n19437 ;
  assign n19439 = ~n19436 & ~n19438 ;
  assign n19440 = ~\P1_P3_InstAddrPointer_reg[12]/NET0131  & ~n19399 ;
  assign n19441 = ~n19435 & ~n19440 ;
  assign n19442 = n19402 & ~n19441 ;
  assign n19443 = ~n19439 & n19442 ;
  assign n19444 = n19439 & ~n19442 ;
  assign n19445 = ~n19443 & ~n19444 ;
  assign n19446 = ~n17282 & ~n19445 ;
  assign n19430 = \P1_P3_InstAddrPointer_reg[12]/NET0131  & n19389 ;
  assign n19431 = ~\P1_P3_InstAddrPointer_reg[13]/NET0131  & ~n19430 ;
  assign n19432 = \P1_P3_InstAddrPointer_reg[13]/NET0131  & n19430 ;
  assign n19433 = ~n19431 & ~n19432 ;
  assign n19447 = \P1_P3_InstAddrPointer_reg[12]/NET0131  & n19394 ;
  assign n19449 = ~n19433 & ~n19447 ;
  assign n19448 = n19433 & n19447 ;
  assign n19450 = n17282 & ~n19448 ;
  assign n19451 = ~n19449 & n19450 ;
  assign n19452 = ~n19446 & ~n19451 ;
  assign n19453 = ~n9072 & n19452 ;
  assign n19454 = ~\P1_P3_InstAddrPointer_reg[13]/NET0131  & n9072 ;
  assign n19455 = n9064 & ~n19454 ;
  assign n19456 = ~n19453 & n19455 ;
  assign n19457 = \P1_P3_InstAddrPointer_reg[12]/NET0131  & n19410 ;
  assign n19458 = ~\P1_P3_InstAddrPointer_reg[13]/NET0131  & ~n19457 ;
  assign n19459 = \P1_P3_InstAddrPointer_reg[13]/NET0131  & n19457 ;
  assign n19460 = ~n19458 & ~n19459 ;
  assign n19461 = \P1_P3_InstAddrPointer_reg[12]/NET0131  & n19412 ;
  assign n19463 = n19460 & n19461 ;
  assign n19462 = ~n19460 & ~n19461 ;
  assign n19464 = n9191 & ~n19462 ;
  assign n19465 = ~n19463 & n19464 ;
  assign n19468 = \P1_P3_InstAddrPointer_reg[13]/NET0131  & ~n19418 ;
  assign n19467 = ~n9133 & n19439 ;
  assign n19434 = ~n9176 & n19433 ;
  assign n19466 = n9220 & n19460 ;
  assign n19469 = ~n19434 & ~n19466 ;
  assign n19470 = ~n19467 & n19469 ;
  assign n19471 = ~n19468 & n19470 ;
  assign n19472 = ~n19465 & n19471 ;
  assign n19473 = ~n19456 & n19472 ;
  assign n19474 = n9241 & ~n19473 ;
  assign n19429 = \P1_P3_rEIP_reg[13]/NET0131  & n17426 ;
  assign n19475 = \P1_P3_InstAddrPointer_reg[13]/NET0131  & ~n18343 ;
  assign n19476 = ~n19429 & ~n19475 ;
  assign n19477 = ~n19474 & n19476 ;
  assign n19484 = \P1_P3_InstAddrPointer_reg[14]/NET0131  & n9072 ;
  assign n19489 = ~\P1_P3_InstAddrPointer_reg[14]/NET0131  & ~n19438 ;
  assign n19480 = \P1_P3_InstAddrPointer_reg[13]/NET0131  & \P1_P3_InstAddrPointer_reg[14]/NET0131  ;
  assign n19490 = n19435 & n19480 ;
  assign n19491 = ~n19489 & ~n19490 ;
  assign n19493 = ~n19443 & n19491 ;
  assign n19492 = n19443 & ~n19491 ;
  assign n19494 = ~n17282 & ~n19492 ;
  assign n19495 = ~n19493 & n19494 ;
  assign n19479 = ~\P1_P3_InstAddrPointer_reg[14]/NET0131  & ~n19432 ;
  assign n19481 = n19430 & n19480 ;
  assign n19482 = ~n19479 & ~n19481 ;
  assign n19485 = ~n19448 & ~n19482 ;
  assign n19486 = \P1_P3_InstAddrPointer_reg[14]/NET0131  & n19448 ;
  assign n19487 = ~n19485 & ~n19486 ;
  assign n19488 = n17282 & ~n19487 ;
  assign n19496 = ~n9072 & ~n19488 ;
  assign n19497 = ~n19495 & n19496 ;
  assign n19498 = ~n19484 & ~n19497 ;
  assign n19499 = n9064 & ~n19498 ;
  assign n19504 = \P1_P3_InstAddrPointer_reg[14]/NET0131  & n19463 ;
  assign n19500 = ~\P1_P3_InstAddrPointer_reg[14]/NET0131  & ~n19459 ;
  assign n19501 = \P1_P3_InstAddrPointer_reg[14]/NET0131  & n19459 ;
  assign n19502 = ~n19500 & ~n19501 ;
  assign n19503 = ~n19463 & ~n19502 ;
  assign n19505 = n9191 & ~n19503 ;
  assign n19506 = ~n19504 & n19505 ;
  assign n19512 = ~n9133 & n19491 ;
  assign n19507 = ~n9050 & ~n9193 ;
  assign n19508 = n9075 & ~n9116 ;
  assign n19509 = n19507 & ~n19508 ;
  assign n19510 = ~n9167 & n19509 ;
  assign n19511 = \P1_P3_InstAddrPointer_reg[14]/NET0131  & ~n19510 ;
  assign n19483 = ~n9176 & n19482 ;
  assign n19514 = n9049 & ~n19502 ;
  assign n19513 = ~\P1_P3_InstAddrPointer_reg[14]/NET0131  & ~n9049 ;
  assign n19515 = ~n9061 & ~n19513 ;
  assign n19516 = ~n19514 & n19515 ;
  assign n19517 = ~n19483 & ~n19516 ;
  assign n19518 = ~n19511 & n19517 ;
  assign n19519 = ~n19512 & n19518 ;
  assign n19520 = ~n19506 & n19519 ;
  assign n19521 = ~n19499 & n19520 ;
  assign n19522 = n9241 & ~n19521 ;
  assign n19478 = \P1_P3_rEIP_reg[14]/NET0131  & n17426 ;
  assign n19523 = \P1_P3_InstAddrPointer_reg[14]/NET0131  & ~n18343 ;
  assign n19524 = ~n19478 & ~n19523 ;
  assign n19525 = ~n19522 & n19524 ;
  assign n19528 = ~\P1_P3_InstAddrPointer_reg[15]/NET0131  & ~n19490 ;
  assign n19529 = \P1_P3_InstAddrPointer_reg[15]/NET0131  & n19490 ;
  assign n19530 = ~n19528 & ~n19529 ;
  assign n19531 = ~n19492 & n19530 ;
  assign n19532 = n19492 & ~n19530 ;
  assign n19533 = ~n19531 & ~n19532 ;
  assign n19534 = ~n17282 & ~n19533 ;
  assign n19535 = n19447 & n19480 ;
  assign n19540 = \P1_P3_InstAddrPointer_reg[15]/NET0131  & n19535 ;
  assign n19536 = ~\P1_P3_InstAddrPointer_reg[15]/NET0131  & ~n19481 ;
  assign n19537 = \P1_P3_InstAddrPointer_reg[15]/NET0131  & n19481 ;
  assign n19538 = ~n19536 & ~n19537 ;
  assign n19539 = ~n19535 & ~n19538 ;
  assign n19541 = n17282 & ~n19539 ;
  assign n19542 = ~n19540 & n19541 ;
  assign n19543 = ~n19534 & ~n19542 ;
  assign n19544 = ~n9072 & n19543 ;
  assign n19545 = ~\P1_P3_InstAddrPointer_reg[15]/NET0131  & n9072 ;
  assign n19546 = n9064 & ~n19545 ;
  assign n19547 = ~n19544 & n19546 ;
  assign n19548 = ~\P1_P3_InstAddrPointer_reg[15]/NET0131  & ~n19501 ;
  assign n19549 = \P1_P3_InstAddrPointer_reg[15]/NET0131  & n19501 ;
  assign n19550 = ~n19548 & ~n19549 ;
  assign n19556 = n19504 & n19550 ;
  assign n19555 = ~n19504 & ~n19550 ;
  assign n19557 = n9191 & ~n19555 ;
  assign n19558 = ~n19556 & n19557 ;
  assign n19553 = \P1_P3_InstAddrPointer_reg[15]/NET0131  & ~n19418 ;
  assign n19552 = ~n9133 & n19530 ;
  assign n19551 = n9220 & n19550 ;
  assign n19554 = ~n9176 & n19538 ;
  assign n19559 = ~n19551 & ~n19554 ;
  assign n19560 = ~n19552 & n19559 ;
  assign n19561 = ~n19553 & n19560 ;
  assign n19562 = ~n19558 & n19561 ;
  assign n19563 = ~n19547 & n19562 ;
  assign n19564 = n9241 & ~n19563 ;
  assign n19526 = \P1_P3_rEIP_reg[15]/NET0131  & n17426 ;
  assign n19527 = \P1_P3_InstAddrPointer_reg[15]/NET0131  & ~n18343 ;
  assign n19565 = ~n19526 & ~n19527 ;
  assign n19566 = ~n19564 & n19565 ;
  assign n19569 = \P1_P3_InstAddrPointer_reg[12]/NET0131  & n9072 ;
  assign n19575 = ~n19402 & n19441 ;
  assign n19576 = ~n17282 & ~n19442 ;
  assign n19577 = ~n19575 & n19576 ;
  assign n19570 = ~\P1_P3_InstAddrPointer_reg[12]/NET0131  & ~n19389 ;
  assign n19571 = ~n19430 & ~n19570 ;
  assign n19572 = ~n19394 & ~n19571 ;
  assign n19573 = ~n19447 & ~n19572 ;
  assign n19574 = n17282 & ~n19573 ;
  assign n19578 = ~n9072 & ~n19574 ;
  assign n19579 = ~n19577 & n19578 ;
  assign n19580 = ~n19569 & ~n19579 ;
  assign n19581 = n9064 & ~n19580 ;
  assign n19582 = ~\P1_P3_InstAddrPointer_reg[12]/NET0131  & ~n19410 ;
  assign n19583 = ~n19457 & ~n19582 ;
  assign n19584 = ~n19412 & ~n19583 ;
  assign n19585 = n9191 & ~n19461 ;
  assign n19586 = ~n19584 & n19585 ;
  assign n19568 = ~n9133 & n19441 ;
  assign n19587 = ~n9163 & n18435 ;
  assign n19588 = \P1_P3_InstAddrPointer_reg[12]/NET0131  & ~n19587 ;
  assign n19589 = ~\P1_P3_InstAddrPointer_reg[12]/NET0131  & n8741 ;
  assign n19590 = ~n8741 & ~n19571 ;
  assign n19591 = ~n19589 & ~n19590 ;
  assign n19592 = ~n9166 & n19591 ;
  assign n19594 = n9049 & ~n19583 ;
  assign n19593 = ~\P1_P3_InstAddrPointer_reg[12]/NET0131  & ~n9049 ;
  assign n19595 = ~n9061 & ~n19593 ;
  assign n19596 = ~n19594 & n19595 ;
  assign n19597 = n9118 & n19571 ;
  assign n19598 = ~n19596 & ~n19597 ;
  assign n19599 = ~n19592 & n19598 ;
  assign n19600 = ~n19588 & n19599 ;
  assign n19601 = ~n19568 & n19600 ;
  assign n19602 = ~n19586 & n19601 ;
  assign n19603 = ~n19581 & n19602 ;
  assign n19604 = n9241 & ~n19603 ;
  assign n19567 = \P1_P3_rEIP_reg[12]/NET0131  & n17426 ;
  assign n19605 = \P1_P3_InstAddrPointer_reg[12]/NET0131  & ~n18343 ;
  assign n19606 = ~n19567 & ~n19605 ;
  assign n19607 = ~n19604 & n19606 ;
  assign n19616 = \P1_P3_InstAddrPointer_reg[16]/NET0131  & n9072 ;
  assign n19609 = ~\P1_P3_InstAddrPointer_reg[16]/NET0131  & ~n19529 ;
  assign n19610 = \P1_P3_InstAddrPointer_reg[14]/NET0131  & \P1_P3_InstAddrPointer_reg[15]/NET0131  ;
  assign n19611 = \P1_P3_InstAddrPointer_reg[16]/NET0131  & n19610 ;
  assign n19612 = n19432 & n19611 ;
  assign n19613 = \P1_P3_InstAddrPointer_reg[0]/NET0131  & n19612 ;
  assign n19614 = ~n19609 & ~n19613 ;
  assign n19625 = ~n19532 & n19614 ;
  assign n19624 = n19532 & ~n19614 ;
  assign n19626 = ~n17282 & ~n19624 ;
  assign n19627 = ~n19625 & n19626 ;
  assign n19617 = ~\P1_P3_InstAddrPointer_reg[16]/NET0131  & ~n19537 ;
  assign n19618 = ~n19612 & ~n19617 ;
  assign n19619 = n19486 & n19538 ;
  assign n19620 = ~n19618 & ~n19619 ;
  assign n19621 = \P1_P3_InstAddrPointer_reg[16]/NET0131  & n19619 ;
  assign n19622 = ~n19620 & ~n19621 ;
  assign n19623 = n17282 & ~n19622 ;
  assign n19628 = ~n9072 & ~n19623 ;
  assign n19629 = ~n19627 & n19628 ;
  assign n19630 = ~n19616 & ~n19629 ;
  assign n19631 = n9064 & ~n19630 ;
  assign n19636 = \P1_P3_InstAddrPointer_reg[16]/NET0131  & n19556 ;
  assign n19632 = ~\P1_P3_InstAddrPointer_reg[16]/NET0131  & ~n19549 ;
  assign n19633 = n19459 & n19611 ;
  assign n19634 = ~n19632 & ~n19633 ;
  assign n19635 = ~n19556 & ~n19634 ;
  assign n19637 = n9191 & ~n19635 ;
  assign n19638 = ~n19636 & n19637 ;
  assign n19639 = ~n8741 & n19618 ;
  assign n19640 = \P1_P3_InstAddrPointer_reg[16]/NET0131  & n8741 ;
  assign n19641 = ~n19639 & ~n19640 ;
  assign n19642 = ~n9075 & n19641 ;
  assign n19643 = n9086 & ~n19642 ;
  assign n19644 = n9075 & n9085 ;
  assign n19645 = ~n9050 & ~n19644 ;
  assign n19646 = ~n9163 & n19645 ;
  assign n19647 = ~n19643 & n19646 ;
  assign n19648 = \P1_P3_InstAddrPointer_reg[16]/NET0131  & ~n19647 ;
  assign n19650 = n9049 & ~n19634 ;
  assign n19651 = ~\P1_P3_InstAddrPointer_reg[16]/NET0131  & ~n9049 ;
  assign n19652 = ~n9061 & ~n19651 ;
  assign n19653 = ~n19650 & n19652 ;
  assign n19615 = ~n9133 & n19614 ;
  assign n19649 = n9118 & n19618 ;
  assign n19654 = ~n9166 & ~n19641 ;
  assign n19655 = ~n19649 & ~n19654 ;
  assign n19656 = ~n19615 & n19655 ;
  assign n19657 = ~n19653 & n19656 ;
  assign n19658 = ~n19648 & n19657 ;
  assign n19659 = ~n19638 & n19658 ;
  assign n19660 = ~n19631 & n19659 ;
  assign n19661 = n9241 & ~n19660 ;
  assign n19608 = \P1_P3_rEIP_reg[16]/NET0131  & n17426 ;
  assign n19662 = \P1_P3_InstAddrPointer_reg[16]/NET0131  & ~n18343 ;
  assign n19663 = ~n19608 & ~n19662 ;
  assign n19664 = ~n19661 & n19663 ;
  assign n19671 = \P1_P3_InstAddrPointer_reg[17]/NET0131  & n9072 ;
  assign n19679 = ~\P1_P3_InstAddrPointer_reg[17]/NET0131  & ~n19613 ;
  assign n19667 = \P1_P3_InstAddrPointer_reg[16]/NET0131  & \P1_P3_InstAddrPointer_reg[17]/NET0131  ;
  assign n19672 = n19537 & n19667 ;
  assign n19680 = \P1_P3_InstAddrPointer_reg[0]/NET0131  & n19672 ;
  assign n19681 = ~n19679 & ~n19680 ;
  assign n19683 = ~n19624 & n19681 ;
  assign n19682 = n19624 & ~n19681 ;
  assign n19684 = ~n17282 & ~n19682 ;
  assign n19685 = ~n19683 & n19684 ;
  assign n19673 = ~\P1_P3_InstAddrPointer_reg[17]/NET0131  & ~n19612 ;
  assign n19674 = ~n19672 & ~n19673 ;
  assign n19675 = ~n19621 & ~n19674 ;
  assign n19676 = \P1_P3_InstAddrPointer_reg[17]/NET0131  & n19621 ;
  assign n19677 = ~n19675 & ~n19676 ;
  assign n19678 = n17282 & ~n19677 ;
  assign n19686 = ~n9072 & ~n19678 ;
  assign n19687 = ~n19685 & n19686 ;
  assign n19688 = ~n19671 & ~n19687 ;
  assign n19689 = n9064 & ~n19688 ;
  assign n19666 = ~\P1_P3_InstAddrPointer_reg[17]/NET0131  & ~n19633 ;
  assign n19668 = n19549 & n19667 ;
  assign n19669 = ~n19666 & ~n19668 ;
  assign n19691 = ~n19636 & ~n19669 ;
  assign n19690 = n19636 & n19669 ;
  assign n19692 = n9191 & ~n19690 ;
  assign n19693 = ~n19691 & n19692 ;
  assign n19696 = ~n9133 & n19681 ;
  assign n19694 = \P1_P3_InstAddrPointer_reg[17]/NET0131  & ~n19418 ;
  assign n19670 = n9220 & n19669 ;
  assign n19695 = ~n9176 & n19674 ;
  assign n19697 = ~n19670 & ~n19695 ;
  assign n19698 = ~n19694 & n19697 ;
  assign n19699 = ~n19696 & n19698 ;
  assign n19700 = ~n19693 & n19699 ;
  assign n19701 = ~n19689 & n19700 ;
  assign n19702 = n9241 & ~n19701 ;
  assign n19665 = \P1_P3_rEIP_reg[17]/NET0131  & n17426 ;
  assign n19703 = \P1_P3_InstAddrPointer_reg[17]/NET0131  & ~n18343 ;
  assign n19704 = ~n19665 & ~n19703 ;
  assign n19705 = ~n19702 & n19704 ;
  assign n19711 = \P1_P3_InstAddrPointer_reg[18]/NET0131  & n9072 ;
  assign n19707 = \P1_P3_InstAddrPointer_reg[18]/NET0131  & ~n19680 ;
  assign n19708 = ~\P1_P3_InstAddrPointer_reg[18]/NET0131  & n19680 ;
  assign n19709 = ~n19707 & ~n19708 ;
  assign n19722 = n19682 & n19709 ;
  assign n19721 = ~n19682 & ~n19709 ;
  assign n19723 = ~n17282 & ~n19721 ;
  assign n19724 = ~n19722 & n19723 ;
  assign n19712 = ~\P1_P3_InstAddrPointer_reg[18]/NET0131  & ~n19672 ;
  assign n19713 = \P1_P3_InstAddrPointer_reg[17]/NET0131  & \P1_P3_InstAddrPointer_reg[18]/NET0131  ;
  assign n19714 = n19612 & n19713 ;
  assign n19715 = ~n19712 & ~n19714 ;
  assign n19716 = ~n19676 & ~n19715 ;
  assign n19717 = \P1_P3_InstAddrPointer_reg[18]/NET0131  & n19667 ;
  assign n19718 = n19619 & n19717 ;
  assign n19719 = ~n19716 & ~n19718 ;
  assign n19720 = n17282 & ~n19719 ;
  assign n19725 = ~n9072 & ~n19720 ;
  assign n19726 = ~n19724 & n19725 ;
  assign n19727 = ~n19711 & ~n19726 ;
  assign n19728 = n9064 & ~n19727 ;
  assign n19733 = \P1_P3_InstAddrPointer_reg[18]/NET0131  & n19690 ;
  assign n19729 = ~\P1_P3_InstAddrPointer_reg[18]/NET0131  & ~n19668 ;
  assign n19730 = n19633 & n19713 ;
  assign n19731 = ~n19729 & ~n19730 ;
  assign n19732 = ~n19690 & ~n19731 ;
  assign n19734 = n9191 & ~n19732 ;
  assign n19735 = ~n19733 & n19734 ;
  assign n19742 = n9220 & n19731 ;
  assign n19710 = ~n9133 & ~n19709 ;
  assign n19739 = n9088 & ~n19715 ;
  assign n19736 = ~\P1_P3_InstAddrPointer_reg[18]/NET0131  & ~n9088 ;
  assign n19737 = ~n9165 & ~n16500 ;
  assign n19738 = ~n9086 & n19737 ;
  assign n19740 = ~n19736 & ~n19738 ;
  assign n19741 = ~n19739 & n19740 ;
  assign n19743 = n9118 & n19715 ;
  assign n19744 = ~n9062 & n19646 ;
  assign n19745 = \P1_P3_InstAddrPointer_reg[18]/NET0131  & ~n19744 ;
  assign n19746 = ~n19743 & ~n19745 ;
  assign n19747 = ~n19741 & n19746 ;
  assign n19748 = ~n19710 & n19747 ;
  assign n19749 = ~n19742 & n19748 ;
  assign n19750 = ~n19735 & n19749 ;
  assign n19751 = ~n19728 & n19750 ;
  assign n19752 = n9241 & ~n19751 ;
  assign n19706 = \P1_P3_rEIP_reg[18]/NET0131  & n17426 ;
  assign n19753 = \P1_P3_InstAddrPointer_reg[18]/NET0131  & ~n18343 ;
  assign n19754 = ~n19706 & ~n19753 ;
  assign n19755 = ~n19752 & n19754 ;
  assign n19761 = \P1_P3_InstAddrPointer_reg[19]/NET0131  & n9072 ;
  assign n19768 = n19529 & n19717 ;
  assign n19769 = ~\P1_P3_InstAddrPointer_reg[19]/NET0131  & ~n19768 ;
  assign n19770 = \P1_P3_InstAddrPointer_reg[19]/NET0131  & n19768 ;
  assign n19771 = ~n19769 & ~n19770 ;
  assign n19772 = ~n19722 & n19771 ;
  assign n19773 = n19709 & ~n19771 ;
  assign n19774 = n19682 & n19773 ;
  assign n19775 = ~n17282 & ~n19774 ;
  assign n19776 = ~n19772 & n19775 ;
  assign n19757 = ~\P1_P3_InstAddrPointer_reg[19]/NET0131  & ~n19714 ;
  assign n19758 = \P1_P3_InstAddrPointer_reg[19]/NET0131  & n19714 ;
  assign n19759 = ~n19757 & ~n19758 ;
  assign n19762 = n19618 & n19713 ;
  assign n19763 = n19540 & n19762 ;
  assign n19764 = n19759 & n19763 ;
  assign n19765 = ~n19759 & ~n19763 ;
  assign n19766 = ~n19764 & ~n19765 ;
  assign n19767 = n17282 & ~n19766 ;
  assign n19777 = ~n9072 & ~n19767 ;
  assign n19778 = ~n19776 & n19777 ;
  assign n19779 = ~n19761 & ~n19778 ;
  assign n19780 = n9064 & ~n19779 ;
  assign n19781 = ~\P1_P3_InstAddrPointer_reg[19]/NET0131  & ~n19730 ;
  assign n19782 = \P1_P3_InstAddrPointer_reg[19]/NET0131  & n19713 ;
  assign n19783 = n19611 & n19782 ;
  assign n19784 = n19459 & n19783 ;
  assign n19785 = ~n19781 & ~n19784 ;
  assign n19787 = ~n19733 & ~n19785 ;
  assign n19786 = n19733 & n19785 ;
  assign n19788 = n9191 & ~n19786 ;
  assign n19789 = ~n19787 & n19788 ;
  assign n19792 = \P1_P3_InstAddrPointer_reg[19]/NET0131  & ~n19418 ;
  assign n19791 = ~n9133 & n19771 ;
  assign n19760 = ~n9176 & n19759 ;
  assign n19790 = n9220 & n19785 ;
  assign n19793 = ~n19760 & ~n19790 ;
  assign n19794 = ~n19791 & n19793 ;
  assign n19795 = ~n19792 & n19794 ;
  assign n19796 = ~n19789 & n19795 ;
  assign n19797 = ~n19780 & n19796 ;
  assign n19798 = n9241 & ~n19797 ;
  assign n19756 = \P1_P3_rEIP_reg[19]/NET0131  & n17426 ;
  assign n19799 = \P1_P3_InstAddrPointer_reg[19]/NET0131  & ~n18343 ;
  assign n19800 = ~n19756 & ~n19799 ;
  assign n19801 = ~n19798 & n19800 ;
  assign n19807 = \P1_P3_InstAddrPointer_reg[20]/NET0131  & n9072 ;
  assign n19813 = ~\P1_P3_InstAddrPointer_reg[20]/NET0131  & ~n19770 ;
  assign n19814 = \P1_P3_InstAddrPointer_reg[20]/NET0131  & n19770 ;
  assign n19815 = ~n19813 & ~n19814 ;
  assign n19817 = ~n19774 & n19815 ;
  assign n19816 = n19774 & ~n19815 ;
  assign n19818 = ~n17282 & ~n19816 ;
  assign n19819 = ~n19817 & n19818 ;
  assign n19803 = \P1_P3_InstAddrPointer_reg[20]/NET0131  & ~n19758 ;
  assign n19804 = ~\P1_P3_InstAddrPointer_reg[20]/NET0131  & n19758 ;
  assign n19805 = ~n19803 & ~n19804 ;
  assign n19808 = n19718 & n19759 ;
  assign n19809 = n19805 & ~n19808 ;
  assign n19810 = \P1_P3_InstAddrPointer_reg[20]/NET0131  & n19808 ;
  assign n19811 = ~n19809 & ~n19810 ;
  assign n19812 = n17282 & ~n19811 ;
  assign n19820 = ~n9072 & ~n19812 ;
  assign n19821 = ~n19819 & n19820 ;
  assign n19822 = ~n19807 & ~n19821 ;
  assign n19823 = n9064 & ~n19822 ;
  assign n19828 = \P1_P3_InstAddrPointer_reg[20]/NET0131  & n19786 ;
  assign n19824 = \P1_P3_InstAddrPointer_reg[20]/NET0131  & ~n19784 ;
  assign n19825 = ~\P1_P3_InstAddrPointer_reg[20]/NET0131  & n19784 ;
  assign n19826 = ~n19824 & ~n19825 ;
  assign n19827 = ~n19786 & n19826 ;
  assign n19829 = n9191 & ~n19827 ;
  assign n19830 = ~n19828 & n19829 ;
  assign n19831 = ~n9061 & ~n19784 ;
  assign n19832 = n18438 & ~n19831 ;
  assign n19833 = \P1_P3_InstAddrPointer_reg[20]/NET0131  & ~n19832 ;
  assign n19835 = ~n9133 & n19815 ;
  assign n19806 = ~n9176 & ~n19805 ;
  assign n19834 = n9220 & ~n19826 ;
  assign n19836 = ~n19806 & ~n19834 ;
  assign n19837 = ~n19835 & n19836 ;
  assign n19838 = ~n19833 & n19837 ;
  assign n19839 = ~n19830 & n19838 ;
  assign n19840 = ~n19823 & n19839 ;
  assign n19841 = n9241 & ~n19840 ;
  assign n19802 = \P1_P3_rEIP_reg[20]/NET0131  & n17426 ;
  assign n19842 = \P1_P3_InstAddrPointer_reg[20]/NET0131  & ~n18343 ;
  assign n19843 = ~n19802 & ~n19842 ;
  assign n19844 = ~n19841 & n19843 ;
  assign n19860 = \P1_P3_InstAddrPointer_reg[21]/NET0131  & n9072 ;
  assign n19847 = \P1_P3_InstAddrPointer_reg[6]/NET0131  & \P1_P3_InstAddrPointer_reg[7]/NET0131  ;
  assign n19848 = \P1_P3_InstAddrPointer_reg[8]/NET0131  & n19847 ;
  assign n19849 = n19437 & n19848 ;
  assign n19850 = n19398 & n19849 ;
  assign n19846 = \P1_P3_InstAddrPointer_reg[20]/NET0131  & n19783 ;
  assign n19851 = \P1_P3_InstAddrPointer_reg[5]/NET0131  & n19846 ;
  assign n19852 = n19850 & n19851 ;
  assign n19865 = \P1_P3_InstAddrPointer_reg[0]/NET0131  & n19852 ;
  assign n19866 = \P1_P3_InstAddrPointer_reg[21]/NET0131  & ~n19865 ;
  assign n19854 = ~\P1_P3_InstAddrPointer_reg[21]/NET0131  & ~n19193 ;
  assign n19855 = \P1_P3_InstAddrPointer_reg[21]/NET0131  & n19193 ;
  assign n19856 = ~n19854 & ~n19855 ;
  assign n19857 = n19852 & n19856 ;
  assign n19867 = \P1_P3_InstAddrPointer_reg[0]/NET0131  & n19857 ;
  assign n19868 = ~n19866 & ~n19867 ;
  assign n19869 = ~n19816 & ~n19868 ;
  assign n19870 = ~n19815 & n19868 ;
  assign n19871 = n19774 & n19870 ;
  assign n19872 = ~n17282 & ~n19871 ;
  assign n19873 = ~n19869 & n19872 ;
  assign n19853 = \P1_P3_InstAddrPointer_reg[21]/NET0131  & ~n19852 ;
  assign n19858 = ~n19853 & ~n19857 ;
  assign n19861 = ~n19810 & n19858 ;
  assign n19862 = n19810 & ~n19858 ;
  assign n19863 = ~n19861 & ~n19862 ;
  assign n19864 = n17282 & ~n19863 ;
  assign n19874 = ~n9072 & ~n19864 ;
  assign n19875 = ~n19873 & n19874 ;
  assign n19876 = ~n19860 & ~n19875 ;
  assign n19877 = n9064 & ~n19876 ;
  assign n19878 = n19315 & n19852 ;
  assign n19879 = \P1_P3_InstAddrPointer_reg[21]/NET0131  & n19878 ;
  assign n19880 = ~\P1_P3_InstAddrPointer_reg[21]/NET0131  & ~n19878 ;
  assign n19881 = ~n19879 & ~n19880 ;
  assign n19883 = n19828 & n19881 ;
  assign n19882 = ~n19828 & ~n19881 ;
  assign n19884 = n9191 & ~n19882 ;
  assign n19885 = ~n19883 & n19884 ;
  assign n19888 = \P1_P3_InstAddrPointer_reg[21]/NET0131  & ~n19418 ;
  assign n19887 = ~n9133 & ~n19868 ;
  assign n19859 = ~n9176 & ~n19858 ;
  assign n19886 = n9220 & n19881 ;
  assign n19889 = ~n19859 & ~n19886 ;
  assign n19890 = ~n19887 & n19889 ;
  assign n19891 = ~n19888 & n19890 ;
  assign n19892 = ~n19885 & n19891 ;
  assign n19893 = ~n19877 & n19892 ;
  assign n19894 = n9241 & ~n19893 ;
  assign n19845 = \P1_P3_rEIP_reg[21]/NET0131  & n17426 ;
  assign n19895 = \P1_P3_InstAddrPointer_reg[21]/NET0131  & ~n18343 ;
  assign n19896 = ~n19845 & ~n19895 ;
  assign n19897 = ~n19894 & n19896 ;
  assign n19908 = \P1_P3_InstAddrPointer_reg[22]/NET0131  & n9072 ;
  assign n19900 = \P1_P3_InstAddrPointer_reg[21]/NET0131  & n19846 ;
  assign n19903 = ~\P1_P3_InstAddrPointer_reg[22]/NET0131  & n19900 ;
  assign n19915 = n19438 & n19903 ;
  assign n19916 = \P1_P3_InstAddrPointer_reg[0]/NET0131  & n19900 ;
  assign n19917 = n19432 & n19916 ;
  assign n19918 = \P1_P3_InstAddrPointer_reg[22]/NET0131  & ~n19917 ;
  assign n19919 = ~n19915 & ~n19918 ;
  assign n19921 = n19871 & n19919 ;
  assign n19920 = ~n19871 & ~n19919 ;
  assign n19922 = ~n17282 & ~n19920 ;
  assign n19923 = ~n19921 & n19922 ;
  assign n19899 = ~\P1_P3_InstAddrPointer_reg[22]/NET0131  & ~n19432 ;
  assign n19901 = n19850 & n19900 ;
  assign n19902 = \P1_P3_InstAddrPointer_reg[22]/NET0131  & ~n19901 ;
  assign n19904 = n19194 & ~n19903 ;
  assign n19905 = ~n19902 & n19904 ;
  assign n19906 = ~n19899 & ~n19905 ;
  assign n19909 = ~n19862 & ~n19906 ;
  assign n19910 = ~n19858 & n19906 ;
  assign n19911 = ~n19805 & n19910 ;
  assign n19912 = n19808 & n19911 ;
  assign n19913 = ~n19909 & ~n19912 ;
  assign n19914 = n17282 & ~n19913 ;
  assign n19924 = ~n9072 & ~n19914 ;
  assign n19925 = ~n19923 & n19924 ;
  assign n19926 = ~n19908 & ~n19925 ;
  assign n19927 = n9064 & ~n19926 ;
  assign n19928 = n19316 & n19901 ;
  assign n19929 = \P1_P3_InstAddrPointer_reg[22]/NET0131  & ~n19928 ;
  assign n19930 = n19459 & n19903 ;
  assign n19931 = ~n19929 & ~n19930 ;
  assign n19933 = ~n19883 & n19931 ;
  assign n19932 = n19883 & ~n19931 ;
  assign n19934 = n9191 & ~n19932 ;
  assign n19935 = ~n19933 & n19934 ;
  assign n19938 = \P1_P3_InstAddrPointer_reg[22]/NET0131  & ~n19418 ;
  assign n19937 = ~n9133 & ~n19919 ;
  assign n19907 = ~n9176 & n19906 ;
  assign n19936 = n9220 & ~n19931 ;
  assign n19939 = ~n19907 & ~n19936 ;
  assign n19940 = ~n19937 & n19939 ;
  assign n19941 = ~n19938 & n19940 ;
  assign n19942 = ~n19935 & n19941 ;
  assign n19943 = ~n19927 & n19942 ;
  assign n19944 = n9241 & ~n19943 ;
  assign n19898 = \P1_P3_rEIP_reg[22]/NET0131  & n17426 ;
  assign n19945 = \P1_P3_InstAddrPointer_reg[22]/NET0131  & ~n18343 ;
  assign n19946 = ~n19898 & ~n19945 ;
  assign n19947 = ~n19944 & n19946 ;
  assign n19956 = \P1_P3_InstAddrPointer_reg[23]/NET0131  & n9072 ;
  assign n19949 = \P1_P3_InstAddrPointer_reg[13]/NET0131  & \P1_P3_InstAddrPointer_reg[22]/NET0131  ;
  assign n19950 = n19900 & n19949 ;
  assign n19962 = n19435 & n19950 ;
  assign n19963 = ~\P1_P3_InstAddrPointer_reg[23]/NET0131  & ~n19962 ;
  assign n19964 = \P1_P3_InstAddrPointer_reg[23]/NET0131  & n19962 ;
  assign n19965 = ~n19963 & ~n19964 ;
  assign n19967 = ~n19921 & n19965 ;
  assign n19966 = n19921 & ~n19965 ;
  assign n19968 = ~n17282 & ~n19966 ;
  assign n19969 = ~n19967 & n19968 ;
  assign n19951 = n19430 & n19950 ;
  assign n19952 = ~\P1_P3_InstAddrPointer_reg[23]/NET0131  & ~n19951 ;
  assign n19953 = \P1_P3_InstAddrPointer_reg[23]/NET0131  & n19951 ;
  assign n19954 = ~n19952 & ~n19953 ;
  assign n19957 = n19912 & n19954 ;
  assign n19958 = n19764 & n19911 ;
  assign n19959 = ~n19954 & ~n19958 ;
  assign n19960 = ~n19957 & ~n19959 ;
  assign n19961 = n17282 & ~n19960 ;
  assign n19970 = ~n9072 & ~n19961 ;
  assign n19971 = ~n19969 & n19970 ;
  assign n19972 = ~n19956 & ~n19971 ;
  assign n19973 = n9064 & ~n19972 ;
  assign n19974 = n19457 & n19950 ;
  assign n19975 = ~\P1_P3_InstAddrPointer_reg[23]/NET0131  & ~n19974 ;
  assign n19976 = \P1_P3_InstAddrPointer_reg[23]/NET0131  & n19974 ;
  assign n19977 = ~n19975 & ~n19976 ;
  assign n19979 = ~n19932 & ~n19977 ;
  assign n19978 = n19932 & n19977 ;
  assign n19980 = n9191 & ~n19978 ;
  assign n19981 = ~n19979 & n19980 ;
  assign n19984 = \P1_P3_InstAddrPointer_reg[23]/NET0131  & ~n19418 ;
  assign n19983 = ~n9133 & n19965 ;
  assign n19955 = ~n9176 & n19954 ;
  assign n19982 = n9220 & n19977 ;
  assign n19985 = ~n19955 & ~n19982 ;
  assign n19986 = ~n19983 & n19985 ;
  assign n19987 = ~n19984 & n19986 ;
  assign n19988 = ~n19981 & n19987 ;
  assign n19989 = ~n19973 & n19988 ;
  assign n19990 = n9241 & ~n19989 ;
  assign n19948 = \P1_P3_rEIP_reg[23]/NET0131  & n17426 ;
  assign n19991 = \P1_P3_InstAddrPointer_reg[23]/NET0131  & ~n18343 ;
  assign n19992 = ~n19948 & ~n19991 ;
  assign n19993 = ~n19990 & n19992 ;
  assign n19999 = \P1_P3_InstAddrPointer_reg[24]/NET0131  & n9072 ;
  assign n19995 = \P1_P3_InstAddrPointer_reg[24]/NET0131  & ~n19964 ;
  assign n19996 = ~\P1_P3_InstAddrPointer_reg[24]/NET0131  & n19964 ;
  assign n19997 = ~n19995 & ~n19996 ;
  assign n20008 = ~n19966 & ~n19997 ;
  assign n20007 = n19966 & n19997 ;
  assign n20009 = ~n17282 & ~n20007 ;
  assign n20010 = ~n20008 & n20009 ;
  assign n20000 = ~\P1_P3_InstAddrPointer_reg[24]/NET0131  & ~n19953 ;
  assign n20001 = \P1_P3_InstAddrPointer_reg[24]/NET0131  & n19953 ;
  assign n20002 = ~n20000 & ~n20001 ;
  assign n20003 = ~n19957 & ~n20002 ;
  assign n20004 = \P1_P3_InstAddrPointer_reg[24]/NET0131  & n19957 ;
  assign n20005 = ~n20003 & ~n20004 ;
  assign n20006 = n17282 & ~n20005 ;
  assign n20011 = ~n9072 & ~n20006 ;
  assign n20012 = ~n20010 & n20011 ;
  assign n20013 = ~n19999 & ~n20012 ;
  assign n20014 = n9064 & ~n20013 ;
  assign n20019 = \P1_P3_InstAddrPointer_reg[24]/NET0131  & n19978 ;
  assign n20015 = ~\P1_P3_InstAddrPointer_reg[24]/NET0131  & ~n19976 ;
  assign n20016 = \P1_P3_InstAddrPointer_reg[24]/NET0131  & n19976 ;
  assign n20017 = ~n20015 & ~n20016 ;
  assign n20018 = ~n19978 & ~n20017 ;
  assign n20020 = n9191 & ~n20018 ;
  assign n20021 = ~n20019 & n20020 ;
  assign n20024 = ~n8741 & ~n20002 ;
  assign n20025 = ~n19737 & ~n20024 ;
  assign n20026 = n9086 & ~n9088 ;
  assign n20027 = n19744 & ~n20026 ;
  assign n20028 = ~n20025 & n20027 ;
  assign n20029 = \P1_P3_InstAddrPointer_reg[24]/NET0131  & ~n20028 ;
  assign n19998 = ~n9133 & ~n19997 ;
  assign n20022 = ~n9176 & n20002 ;
  assign n20023 = n9220 & n20017 ;
  assign n20030 = ~n20022 & ~n20023 ;
  assign n20031 = ~n19998 & n20030 ;
  assign n20032 = ~n20029 & n20031 ;
  assign n20033 = ~n20021 & n20032 ;
  assign n20034 = ~n20014 & n20033 ;
  assign n20035 = n9241 & ~n20034 ;
  assign n19994 = \P1_P3_rEIP_reg[24]/NET0131  & n17426 ;
  assign n20036 = \P1_P3_InstAddrPointer_reg[24]/NET0131  & ~n18343 ;
  assign n20037 = ~n19994 & ~n20036 ;
  assign n20038 = ~n20035 & n20037 ;
  assign n20044 = \P1_P3_InstAddrPointer_reg[25]/NET0131  & n9072 ;
  assign n20053 = \P1_P3_InstAddrPointer_reg[0]/NET0131  & n20001 ;
  assign n20054 = ~\P1_P3_InstAddrPointer_reg[25]/NET0131  & ~n20053 ;
  assign n20055 = \P1_P3_InstAddrPointer_reg[25]/NET0131  & n20053 ;
  assign n20056 = ~n20054 & ~n20055 ;
  assign n20057 = ~n20007 & n20056 ;
  assign n20058 = n19997 & ~n20056 ;
  assign n20059 = n19966 & n20058 ;
  assign n20060 = ~n17282 & ~n20059 ;
  assign n20061 = ~n20057 & n20060 ;
  assign n20045 = ~\P1_P3_InstAddrPointer_reg[25]/NET0131  & ~n20001 ;
  assign n20046 = \P1_P3_InstAddrPointer_reg[24]/NET0131  & \P1_P3_InstAddrPointer_reg[25]/NET0131  ;
  assign n20047 = n19953 & n20046 ;
  assign n20048 = ~n20045 & ~n20047 ;
  assign n20049 = ~n20004 & ~n20048 ;
  assign n20050 = n19957 & n20046 ;
  assign n20051 = ~n20049 & ~n20050 ;
  assign n20052 = n17282 & ~n20051 ;
  assign n20062 = ~n9072 & ~n20052 ;
  assign n20063 = ~n20061 & n20062 ;
  assign n20064 = ~n20044 & ~n20063 ;
  assign n20065 = n9064 & ~n20064 ;
  assign n20040 = ~\P1_P3_InstAddrPointer_reg[25]/NET0131  & ~n20016 ;
  assign n20041 = \P1_P3_InstAddrPointer_reg[25]/NET0131  & n20016 ;
  assign n20042 = ~n20040 & ~n20041 ;
  assign n20067 = n20019 & n20042 ;
  assign n20066 = ~n20019 & ~n20042 ;
  assign n20068 = n9191 & ~n20066 ;
  assign n20069 = ~n20067 & n20068 ;
  assign n20072 = ~n9133 & n20056 ;
  assign n20070 = \P1_P3_InstAddrPointer_reg[25]/NET0131  & ~n19418 ;
  assign n20043 = n9220 & n20042 ;
  assign n20071 = ~n9176 & n20048 ;
  assign n20073 = ~n20043 & ~n20071 ;
  assign n20074 = ~n20070 & n20073 ;
  assign n20075 = ~n20072 & n20074 ;
  assign n20076 = ~n20069 & n20075 ;
  assign n20077 = ~n20065 & n20076 ;
  assign n20078 = n9241 & ~n20077 ;
  assign n20039 = \P1_P3_rEIP_reg[25]/NET0131  & n17426 ;
  assign n20079 = \P1_P3_InstAddrPointer_reg[25]/NET0131  & ~n18343 ;
  assign n20080 = ~n20039 & ~n20079 ;
  assign n20081 = ~n20078 & n20080 ;
  assign n20084 = \P1_P3_InstAddrPointer_reg[26]/NET0131  & n9072 ;
  assign n20094 = n19964 & n20046 ;
  assign n20095 = ~\P1_P3_InstAddrPointer_reg[26]/NET0131  & ~n20094 ;
  assign n20096 = \P1_P3_InstAddrPointer_reg[26]/NET0131  & n20094 ;
  assign n20097 = ~n20095 & ~n20096 ;
  assign n20099 = ~n20059 & n20097 ;
  assign n20098 = n20059 & ~n20097 ;
  assign n20100 = ~n17282 & ~n20098 ;
  assign n20101 = ~n20099 & n20100 ;
  assign n20085 = ~\P1_P3_InstAddrPointer_reg[26]/NET0131  & ~n20047 ;
  assign n20086 = \P1_P3_InstAddrPointer_reg[26]/NET0131  & n20047 ;
  assign n20087 = ~n20085 & ~n20086 ;
  assign n20088 = ~n20050 & ~n20087 ;
  assign n20089 = n19954 & n20046 ;
  assign n20090 = n20087 & n20089 ;
  assign n20091 = n19912 & n20090 ;
  assign n20092 = ~n20088 & ~n20091 ;
  assign n20093 = n17282 & ~n20092 ;
  assign n20102 = ~n9072 & ~n20093 ;
  assign n20103 = ~n20101 & n20102 ;
  assign n20104 = ~n20084 & ~n20103 ;
  assign n20105 = n9064 & ~n20104 ;
  assign n20119 = \P1_P3_InstAddrPointer_reg[26]/NET0131  & n20067 ;
  assign n20114 = ~\P1_P3_InstAddrPointer_reg[26]/NET0131  & ~n20041 ;
  assign n20115 = \P1_P3_InstAddrPointer_reg[26]/NET0131  & n20041 ;
  assign n20116 = ~n20114 & ~n20115 ;
  assign n20118 = ~n20067 & ~n20116 ;
  assign n20120 = n9191 & ~n20118 ;
  assign n20121 = ~n20119 & n20120 ;
  assign n20106 = ~n9176 & n20087 ;
  assign n20107 = ~n9050 & ~n9089 ;
  assign n20108 = ~n9137 & n20107 ;
  assign n20109 = ~n9062 & n20108 ;
  assign n20110 = ~n9061 & ~n20041 ;
  assign n20111 = n20109 & ~n20110 ;
  assign n20112 = \P1_P3_InstAddrPointer_reg[26]/NET0131  & ~n20111 ;
  assign n20122 = ~n20106 & ~n20112 ;
  assign n20113 = ~n9133 & n20097 ;
  assign n20117 = n9220 & n20116 ;
  assign n20123 = ~n20113 & ~n20117 ;
  assign n20124 = n20122 & n20123 ;
  assign n20125 = ~n20121 & n20124 ;
  assign n20126 = ~n20105 & n20125 ;
  assign n20127 = n9241 & ~n20126 ;
  assign n20082 = \P1_P3_rEIP_reg[26]/NET0131  & n17426 ;
  assign n20083 = \P1_P3_InstAddrPointer_reg[26]/NET0131  & ~n18343 ;
  assign n20128 = ~n20082 & ~n20083 ;
  assign n20129 = ~n20127 & n20128 ;
  assign n20149 = \P1_P3_InstAddrPointer_reg[27]/NET0131  & n9072 ;
  assign n20140 = \P1_P3_InstAddrPointer_reg[26]/NET0131  & n20055 ;
  assign n20141 = ~\P1_P3_InstAddrPointer_reg[27]/NET0131  & ~n20140 ;
  assign n20142 = \P1_P3_InstAddrPointer_reg[27]/NET0131  & n20140 ;
  assign n20143 = ~n20141 & ~n20142 ;
  assign n20155 = ~n20098 & n20143 ;
  assign n20156 = ~n19965 & ~n20097 ;
  assign n20157 = n20058 & n20156 ;
  assign n20158 = ~n20143 & n20157 ;
  assign n20159 = n19921 & n20158 ;
  assign n20160 = ~n17282 & ~n20159 ;
  assign n20161 = ~n20155 & n20160 ;
  assign n20136 = \P1_P3_InstAddrPointer_reg[27]/NET0131  & n20086 ;
  assign n20137 = ~\P1_P3_InstAddrPointer_reg[27]/NET0131  & ~n20086 ;
  assign n20138 = ~n20136 & ~n20137 ;
  assign n20150 = n19958 & n20090 ;
  assign n20151 = ~n20138 & ~n20150 ;
  assign n20152 = n20138 & n20150 ;
  assign n20153 = ~n20151 & ~n20152 ;
  assign n20154 = n17282 & ~n20153 ;
  assign n20162 = ~n9072 & ~n20154 ;
  assign n20163 = ~n20161 & n20162 ;
  assign n20164 = ~n20149 & ~n20163 ;
  assign n20165 = n9064 & ~n20164 ;
  assign n20132 = ~\P1_P3_InstAddrPointer_reg[27]/NET0131  & ~n20115 ;
  assign n20133 = \P1_P3_InstAddrPointer_reg[27]/NET0131  & n20115 ;
  assign n20134 = ~n20132 & ~n20133 ;
  assign n20167 = ~n20119 & ~n20134 ;
  assign n20166 = n20119 & n20134 ;
  assign n20168 = n9191 & ~n20166 ;
  assign n20169 = ~n20167 & n20168 ;
  assign n20144 = ~n9133 & n20143 ;
  assign n20135 = n9220 & n20134 ;
  assign n20139 = ~n9176 & n20138 ;
  assign n20145 = ~n9088 & ~n9116 ;
  assign n20146 = ~n9062 & n19507 ;
  assign n20147 = ~n20145 & n20146 ;
  assign n20148 = \P1_P3_InstAddrPointer_reg[27]/NET0131  & ~n20147 ;
  assign n20170 = ~n20139 & ~n20148 ;
  assign n20171 = ~n20135 & n20170 ;
  assign n20172 = ~n20144 & n20171 ;
  assign n20173 = ~n20169 & n20172 ;
  assign n20174 = ~n20165 & n20173 ;
  assign n20175 = n9241 & ~n20174 ;
  assign n20130 = \P1_P3_rEIP_reg[27]/NET0131  & n17426 ;
  assign n20131 = \P1_P3_InstAddrPointer_reg[27]/NET0131  & ~n18343 ;
  assign n20176 = ~n20130 & ~n20131 ;
  assign n20177 = ~n20175 & n20176 ;
  assign n20201 = \P1_P3_InstAddrPointer_reg[28]/NET0131  & n20133 ;
  assign n20202 = ~\P1_P3_InstAddrPointer_reg[28]/NET0131  & ~n20133 ;
  assign n20203 = ~n20201 & ~n20202 ;
  assign n20209 = ~n20166 & ~n20203 ;
  assign n20208 = \P1_P3_InstAddrPointer_reg[28]/NET0131  & n20166 ;
  assign n20210 = n9191 & ~n20208 ;
  assign n20211 = ~n20209 & n20210 ;
  assign n20180 = \P1_P3_InstAddrPointer_reg[28]/NET0131  & n9072 ;
  assign n20189 = \P1_P3_InstAddrPointer_reg[27]/NET0131  & n20096 ;
  assign n20190 = \P1_P3_InstAddrPointer_reg[28]/NET0131  & n20189 ;
  assign n20191 = ~\P1_P3_InstAddrPointer_reg[28]/NET0131  & ~n20189 ;
  assign n20192 = ~n20190 & ~n20191 ;
  assign n20194 = n20159 & ~n20192 ;
  assign n20193 = ~n20159 & n20192 ;
  assign n20195 = ~n17282 & ~n20193 ;
  assign n20196 = ~n20194 & n20195 ;
  assign n20181 = ~\P1_P3_InstAddrPointer_reg[28]/NET0131  & ~n20136 ;
  assign n20182 = \P1_P3_InstAddrPointer_reg[28]/NET0131  & n20136 ;
  assign n20183 = ~n20181 & ~n20182 ;
  assign n20184 = \P1_P3_InstAddrPointer_reg[27]/NET0131  & n20091 ;
  assign n20185 = ~n20183 & ~n20184 ;
  assign n20186 = \P1_P3_InstAddrPointer_reg[28]/NET0131  & n20184 ;
  assign n20187 = ~n20185 & ~n20186 ;
  assign n20188 = n17282 & ~n20187 ;
  assign n20197 = ~n9072 & ~n20188 ;
  assign n20198 = ~n20196 & n20197 ;
  assign n20199 = ~n20180 & ~n20198 ;
  assign n20200 = n9064 & ~n20199 ;
  assign n20204 = n9220 & n20203 ;
  assign n20207 = ~n9176 & n20183 ;
  assign n20205 = ~n9133 & n20192 ;
  assign n20206 = \P1_P3_InstAddrPointer_reg[28]/NET0131  & ~n19418 ;
  assign n20212 = ~n20205 & ~n20206 ;
  assign n20213 = ~n20207 & n20212 ;
  assign n20214 = ~n20204 & n20213 ;
  assign n20215 = ~n20200 & n20214 ;
  assign n20216 = ~n20211 & n20215 ;
  assign n20217 = n9241 & ~n20216 ;
  assign n20178 = \P1_P3_rEIP_reg[28]/NET0131  & n17426 ;
  assign n20179 = \P1_P3_InstAddrPointer_reg[28]/NET0131  & ~n18343 ;
  assign n20218 = ~n20178 & ~n20179 ;
  assign n20219 = ~n20217 & n20218 ;
  assign n20247 = \P1_P3_InstAddrPointer_reg[29]/NET0131  & n20201 ;
  assign n20248 = ~\P1_P3_InstAddrPointer_reg[29]/NET0131  & ~n20201 ;
  assign n20249 = ~n20247 & ~n20248 ;
  assign n20253 = ~n20208 & ~n20249 ;
  assign n20251 = \P1_P3_InstAddrPointer_reg[29]/NET0131  & n20203 ;
  assign n20252 = n20166 & n20251 ;
  assign n20254 = n9191 & ~n20252 ;
  assign n20255 = ~n20253 & n20254 ;
  assign n20222 = \P1_P3_InstAddrPointer_reg[29]/NET0131  & n9072 ;
  assign n20231 = \P1_P3_InstAddrPointer_reg[29]/NET0131  & n20182 ;
  assign n20232 = ~\P1_P3_InstAddrPointer_reg[29]/NET0131  & ~n20182 ;
  assign n20233 = ~n20231 & ~n20232 ;
  assign n20234 = ~n20186 & ~n20233 ;
  assign n20235 = n20186 & n20233 ;
  assign n20236 = ~n20234 & ~n20235 ;
  assign n20237 = n17282 & ~n20236 ;
  assign n20223 = \P1_P3_InstAddrPointer_reg[29]/NET0131  & ~n20190 ;
  assign n20224 = ~\P1_P3_InstAddrPointer_reg[29]/NET0131  & n20190 ;
  assign n20225 = ~n20223 & ~n20224 ;
  assign n20226 = ~n20194 & ~n20225 ;
  assign n20227 = ~n20192 & n20225 ;
  assign n20228 = n20159 & n20227 ;
  assign n20229 = ~n17282 & ~n20228 ;
  assign n20230 = ~n20226 & n20229 ;
  assign n20238 = ~n9072 & ~n20230 ;
  assign n20239 = ~n20237 & n20238 ;
  assign n20240 = ~n20222 & ~n20239 ;
  assign n20241 = n9064 & ~n20240 ;
  assign n20250 = n9220 & n20249 ;
  assign n20243 = ~n9061 & ~n20201 ;
  assign n20244 = n20109 & ~n20243 ;
  assign n20245 = \P1_P3_InstAddrPointer_reg[29]/NET0131  & ~n20244 ;
  assign n20242 = ~n9133 & ~n20225 ;
  assign n20246 = ~n9176 & n20233 ;
  assign n20256 = ~n20242 & ~n20246 ;
  assign n20257 = ~n20245 & n20256 ;
  assign n20258 = ~n20250 & n20257 ;
  assign n20259 = ~n20241 & n20258 ;
  assign n20260 = ~n20255 & n20259 ;
  assign n20261 = n9241 & ~n20260 ;
  assign n20220 = \P1_P3_InstAddrPointer_reg[29]/NET0131  & ~n18343 ;
  assign n20221 = \P1_P3_rEIP_reg[29]/NET0131  & n17426 ;
  assign n20262 = ~n20220 & ~n20221 ;
  assign n20263 = ~n20261 & n20262 ;
  assign n20275 = ~n9073 & n19418 ;
  assign n20276 = \P1_P3_InstAddrPointer_reg[2]/NET0131  & ~n20275 ;
  assign n20274 = ~n9133 & n19233 ;
  assign n20277 = \P1_P3_InstAddrPointer_reg[2]/NET0131  & ~n9166 ;
  assign n20278 = n9176 & ~n20277 ;
  assign n20279 = n19284 & ~n20278 ;
  assign n20266 = ~n19234 & ~n19237 ;
  assign n20267 = ~n19344 & n20266 ;
  assign n20268 = n19344 & ~n20266 ;
  assign n20269 = ~n20267 & ~n20268 ;
  assign n20270 = n9021 & n20269 ;
  assign n20271 = ~n9061 & ~n19233 ;
  assign n20272 = ~n20270 & ~n20271 ;
  assign n20273 = n9049 & ~n20272 ;
  assign n20284 = ~n19285 & ~n19286 ;
  assign n20285 = ~n19288 & ~n20284 ;
  assign n20286 = n19288 & n20284 ;
  assign n20287 = ~n20285 & ~n20286 ;
  assign n20288 = n17282 & ~n20287 ;
  assign n20281 = ~n19234 & n19238 ;
  assign n20280 = ~n19236 & ~n20266 ;
  assign n20282 = ~n17282 & ~n20280 ;
  assign n20283 = ~n20281 & n20282 ;
  assign n20289 = n9192 & ~n20283 ;
  assign n20290 = ~n20288 & n20289 ;
  assign n20291 = ~n20273 & ~n20290 ;
  assign n20292 = ~n20279 & n20291 ;
  assign n20293 = ~n20274 & n20292 ;
  assign n20294 = ~n20276 & n20293 ;
  assign n20295 = n9241 & ~n20294 ;
  assign n20264 = \P1_P3_rEIP_reg[2]/NET0131  & n17426 ;
  assign n20265 = \P1_P3_InstAddrPointer_reg[2]/NET0131  & ~n18343 ;
  assign n20296 = ~n20264 & ~n20265 ;
  assign n20297 = ~n20295 & n20296 ;
  assign n20311 = ~\P1_P3_InstAddrPointer_reg[30]/NET0131  & ~n20247 ;
  assign n20312 = \P1_P3_InstAddrPointer_reg[30]/NET0131  & n20247 ;
  assign n20313 = ~n20311 & ~n20312 ;
  assign n20315 = n20252 & n20313 ;
  assign n20314 = ~n20252 & ~n20313 ;
  assign n20316 = n9191 & ~n20314 ;
  assign n20317 = ~n20315 & n20316 ;
  assign n20304 = \P1_P3_InstAddrPointer_reg[0]/NET0131  & n20231 ;
  assign n20305 = ~\P1_P3_InstAddrPointer_reg[30]/NET0131  & ~n20304 ;
  assign n20306 = \P1_P3_InstAddrPointer_reg[30]/NET0131  & n20304 ;
  assign n20307 = ~n20305 & ~n20306 ;
  assign n20318 = ~n20228 & n20307 ;
  assign n20319 = n20228 & ~n20307 ;
  assign n20320 = ~n20318 & ~n20319 ;
  assign n20321 = ~n17282 & ~n20320 ;
  assign n20300 = \P1_P3_InstAddrPointer_reg[30]/NET0131  & n20231 ;
  assign n20301 = ~\P1_P3_InstAddrPointer_reg[30]/NET0131  & ~n20231 ;
  assign n20302 = ~n20300 & ~n20301 ;
  assign n20323 = ~n20235 & ~n20302 ;
  assign n20322 = \P1_P3_InstAddrPointer_reg[30]/NET0131  & n20235 ;
  assign n20324 = n17282 & ~n20322 ;
  assign n20325 = ~n20323 & n20324 ;
  assign n20326 = ~n20321 & ~n20325 ;
  assign n20327 = n9192 & ~n20326 ;
  assign n20328 = n9220 & n20313 ;
  assign n20308 = ~n9133 & n20307 ;
  assign n20303 = ~n9176 & n20302 ;
  assign n20309 = n9074 & n20108 ;
  assign n20310 = \P1_P3_InstAddrPointer_reg[30]/NET0131  & ~n20309 ;
  assign n20329 = ~n20303 & ~n20310 ;
  assign n20330 = ~n20308 & n20329 ;
  assign n20331 = ~n20328 & n20330 ;
  assign n20332 = ~n20327 & n20331 ;
  assign n20333 = ~n20317 & n20332 ;
  assign n20334 = n9241 & ~n20333 ;
  assign n20298 = \P1_P3_InstAddrPointer_reg[30]/NET0131  & ~n18343 ;
  assign n20299 = \P1_P3_rEIP_reg[30]/NET0131  & n17426 ;
  assign n20335 = ~n20298 & ~n20299 ;
  assign n20336 = ~n20334 & n20335 ;
  assign n20371 = \P1_P3_InstAddrPointer_reg[31]/NET0131  & n20315 ;
  assign n20364 = ~\P1_P3_InstAddrPointer_reg[31]/NET0131  & ~n20312 ;
  assign n20365 = \P1_P3_InstAddrPointer_reg[31]/NET0131  & n20312 ;
  assign n20366 = ~n20364 & ~n20365 ;
  assign n20370 = ~n20315 & ~n20366 ;
  assign n20372 = n9191 & ~n20370 ;
  assign n20373 = ~n20371 & n20372 ;
  assign n20337 = \P1_P3_InstAddrPointer_reg[31]/NET0131  & n9072 ;
  assign n20348 = \P1_P3_InstAddrPointer_reg[31]/NET0131  & ~n20306 ;
  assign n20349 = ~\P1_P3_InstAddrPointer_reg[31]/NET0131  & n20306 ;
  assign n20350 = ~n20348 & ~n20349 ;
  assign n20352 = n20319 & n20350 ;
  assign n20351 = ~n20319 & ~n20350 ;
  assign n20353 = ~n17282 & ~n20351 ;
  assign n20354 = ~n20352 & n20353 ;
  assign n20338 = ~\P1_P3_InstAddrPointer_reg[31]/NET0131  & ~n20300 ;
  assign n20339 = \P1_P3_InstAddrPointer_reg[31]/NET0131  & n20300 ;
  assign n20340 = ~n20338 & ~n20339 ;
  assign n20341 = \P1_P3_InstAddrPointer_reg[29]/NET0131  & n20183 ;
  assign n20342 = n20302 & n20341 ;
  assign n20343 = n20152 & n20342 ;
  assign n20345 = ~n20340 & n20343 ;
  assign n20344 = n20340 & ~n20343 ;
  assign n20346 = n17282 & ~n20344 ;
  assign n20347 = ~n20345 & n20346 ;
  assign n20355 = ~n9072 & ~n20347 ;
  assign n20356 = ~n20354 & n20355 ;
  assign n20357 = ~n20337 & ~n20356 ;
  assign n20358 = n9064 & ~n20357 ;
  assign n20367 = ~\P1_P3_InstAddrPointer_reg[31]/NET0131  & ~n9049 ;
  assign n20368 = ~n9061 & ~n20367 ;
  assign n20369 = n20366 & n20368 ;
  assign n20360 = ~n9133 & ~n20350 ;
  assign n20359 = ~n9176 & n20340 ;
  assign n20361 = n9086 & ~n20300 ;
  assign n20362 = n20147 & ~n20361 ;
  assign n20363 = \P1_P3_InstAddrPointer_reg[31]/NET0131  & ~n20362 ;
  assign n20374 = ~n20359 & ~n20363 ;
  assign n20375 = ~n20360 & n20374 ;
  assign n20376 = ~n20369 & n20375 ;
  assign n20377 = ~n20358 & n20376 ;
  assign n20378 = ~n20373 & n20377 ;
  assign n20379 = n9241 & ~n20378 ;
  assign n20380 = \P1_P3_InstAddrPointer_reg[31]/NET0131  & ~n18343 ;
  assign n20381 = \P1_P3_rEIP_reg[31]/NET0131  & n17426 ;
  assign n20382 = ~n20380 & ~n20381 ;
  assign n20383 = ~n20379 & n20382 ;
  assign n20411 = ~n9133 & n19229 ;
  assign n20389 = ~n19230 & ~n19231 ;
  assign n20391 = ~n19239 & n20389 ;
  assign n20390 = n19239 & ~n20389 ;
  assign n20392 = ~n17282 & ~n20390 ;
  assign n20393 = ~n20391 & n20392 ;
  assign n20394 = ~n19281 & ~n19282 ;
  assign n20396 = ~n19290 & n20394 ;
  assign n20395 = n19290 & ~n20394 ;
  assign n20397 = n17282 & ~n20395 ;
  assign n20398 = ~n20396 & n20397 ;
  assign n20399 = ~n20393 & ~n20398 ;
  assign n20400 = ~n9072 & ~n20399 ;
  assign n20401 = ~\P1_P3_InstAddrPointer_reg[3]/NET0131  & n9072 ;
  assign n20402 = n9064 & ~n20401 ;
  assign n20403 = ~n20400 & n20402 ;
  assign n20412 = ~n9061 & n19232 ;
  assign n20413 = n18436 & ~n20412 ;
  assign n20414 = \P1_P3_InstAddrPointer_reg[3]/NET0131  & ~n20413 ;
  assign n20407 = ~n8741 & ~n19280 ;
  assign n20408 = ~\P1_P3_InstAddrPointer_reg[3]/NET0131  & n8741 ;
  assign n20409 = ~n20407 & ~n20408 ;
  assign n20410 = n9147 & n20409 ;
  assign n20386 = ~\P1_P3_InstAddrPointer_reg[3]/NET0131  & ~n9097 ;
  assign n20387 = ~n9084 & ~n20386 ;
  assign n20388 = ~n9097 & n20387 ;
  assign n20404 = n9220 & n19338 ;
  assign n20420 = ~n20388 & ~n20404 ;
  assign n20421 = ~n20410 & n20420 ;
  assign n20405 = ~n9118 & ~n20387 ;
  assign n20406 = n19280 & ~n20405 ;
  assign n20415 = ~n19339 & ~n19340 ;
  assign n20417 = ~n19346 & n20415 ;
  assign n20416 = n19346 & ~n20415 ;
  assign n20418 = n9191 & ~n20416 ;
  assign n20419 = ~n20417 & n20418 ;
  assign n20422 = ~n20406 & ~n20419 ;
  assign n20423 = n20421 & n20422 ;
  assign n20424 = ~n20414 & n20423 ;
  assign n20425 = ~n20403 & n20424 ;
  assign n20426 = ~n20411 & n20425 ;
  assign n20427 = n9241 & ~n20426 ;
  assign n20384 = \P1_P3_rEIP_reg[3]/NET0131  & n17426 ;
  assign n20385 = \P1_P3_InstAddrPointer_reg[3]/NET0131  & ~n18343 ;
  assign n20428 = ~n20384 & ~n20385 ;
  assign n20429 = ~n20427 & n20428 ;
  assign n20433 = \P1_P3_InstAddrPointer_reg[4]/NET0131  & n9072 ;
  assign n20436 = n19293 & ~n19294 ;
  assign n20434 = ~n19278 & ~n19294 ;
  assign n20435 = ~n19292 & ~n20434 ;
  assign n20437 = ~n9072 & ~n20435 ;
  assign n20438 = ~n20436 & n20437 ;
  assign n20439 = ~n20433 & ~n20438 ;
  assign n20440 = n9064 & ~n20439 ;
  assign n20447 = ~n9133 & n19224 ;
  assign n20450 = n19349 & ~n19350 ;
  assign n20448 = ~n19336 & ~n19350 ;
  assign n20449 = n19348 & ~n20448 ;
  assign n20451 = n9191 & ~n20449 ;
  assign n20452 = ~n20450 & n20451 ;
  assign n20441 = ~n9137 & n18435 ;
  assign n20442 = \P1_P3_InstAddrPointer_reg[4]/NET0131  & ~n20441 ;
  assign n20432 = ~n9174 & n19277 ;
  assign n20443 = ~\P1_P3_InstAddrPointer_reg[4]/NET0131  & n8741 ;
  assign n20444 = ~n8741 & ~n19277 ;
  assign n20445 = ~n20443 & ~n20444 ;
  assign n20446 = n9147 & n20445 ;
  assign n20453 = n9049 & ~n19335 ;
  assign n20454 = ~\P1_P3_InstAddrPointer_reg[4]/NET0131  & ~n9049 ;
  assign n20455 = ~n20453 & ~n20454 ;
  assign n20456 = ~n9061 & n20455 ;
  assign n20457 = ~n20446 & ~n20456 ;
  assign n20458 = ~n20432 & n20457 ;
  assign n20459 = ~n20442 & n20458 ;
  assign n20460 = ~n20452 & n20459 ;
  assign n20461 = ~n20447 & n20460 ;
  assign n20462 = ~n20440 & n20461 ;
  assign n20463 = n9241 & ~n20462 ;
  assign n20430 = \P1_P3_rEIP_reg[4]/NET0131  & n17426 ;
  assign n20431 = \P1_P3_InstAddrPointer_reg[4]/NET0131  & ~n18343 ;
  assign n20464 = ~n20430 & ~n20431 ;
  assign n20465 = ~n20463 & n20464 ;
  assign n20476 = \P1_P3_InstAddrPointer_reg[5]/NET0131  & n9072 ;
  assign n20482 = ~n19220 & ~n19221 ;
  assign n20484 = ~n19243 & n20482 ;
  assign n20483 = n19243 & ~n20482 ;
  assign n20485 = ~n17282 & ~n20483 ;
  assign n20486 = ~n20484 & n20485 ;
  assign n20477 = ~n19274 & ~n19275 ;
  assign n20479 = n19295 & n20477 ;
  assign n20478 = ~n19295 & ~n20477 ;
  assign n20480 = n17282 & ~n20478 ;
  assign n20481 = ~n20479 & n20480 ;
  assign n20487 = ~n9072 & ~n20481 ;
  assign n20488 = ~n20486 & n20487 ;
  assign n20489 = ~n20476 & ~n20488 ;
  assign n20490 = n9064 & ~n20489 ;
  assign n20470 = ~n19332 & ~n19333 ;
  assign n20472 = ~n19351 & n20470 ;
  assign n20471 = n19351 & ~n20470 ;
  assign n20473 = n9191 & ~n20471 ;
  assign n20474 = ~n20472 & n20473 ;
  assign n20475 = ~n9133 & n19219 ;
  assign n20469 = \P1_P3_InstAddrPointer_reg[5]/NET0131  & ~n19418 ;
  assign n20467 = ~n9176 & n19273 ;
  assign n20468 = n9220 & n19331 ;
  assign n20491 = ~n20467 & ~n20468 ;
  assign n20492 = ~n20469 & n20491 ;
  assign n20493 = ~n20475 & n20492 ;
  assign n20494 = ~n20474 & n20493 ;
  assign n20495 = ~n20490 & n20494 ;
  assign n20496 = n9241 & ~n20495 ;
  assign n20466 = \P1_P3_rEIP_reg[5]/NET0131  & n17426 ;
  assign n20497 = \P1_P3_InstAddrPointer_reg[5]/NET0131  & ~n18343 ;
  assign n20498 = ~n20466 & ~n20497 ;
  assign n20499 = ~n20496 & n20498 ;
  assign n20502 = \P1_P3_InstAddrPointer_reg[6]/NET0131  & n9072 ;
  assign n20508 = ~n19215 & ~n19216 ;
  assign n20510 = ~n19245 & n20508 ;
  assign n20509 = n19245 & ~n20508 ;
  assign n20511 = ~n17282 & ~n20509 ;
  assign n20512 = ~n20510 & n20511 ;
  assign n20503 = ~n19270 & ~n19271 ;
  assign n20505 = n19297 & n20503 ;
  assign n20504 = ~n19297 & ~n20503 ;
  assign n20506 = n17282 & ~n20504 ;
  assign n20507 = ~n20505 & n20506 ;
  assign n20513 = ~n9072 & ~n20507 ;
  assign n20514 = ~n20512 & n20513 ;
  assign n20515 = ~n20502 & ~n20514 ;
  assign n20516 = n9064 & ~n20515 ;
  assign n20520 = ~n19328 & n19354 ;
  assign n20518 = ~n19328 & ~n19329 ;
  assign n20519 = n19353 & ~n20518 ;
  assign n20521 = n9191 & ~n20519 ;
  assign n20522 = ~n20520 & n20521 ;
  assign n20517 = ~n9133 & n19214 ;
  assign n20501 = \P1_P3_InstAddrPointer_reg[6]/NET0131  & ~n18435 ;
  assign n20528 = ~n8741 & ~n19269 ;
  assign n20529 = ~\P1_P3_InstAddrPointer_reg[6]/NET0131  & n8741 ;
  assign n20530 = ~n20528 & ~n20529 ;
  assign n20531 = n9147 & n20530 ;
  assign n20524 = n9097 & ~n19269 ;
  assign n20523 = ~\P1_P3_InstAddrPointer_reg[6]/NET0131  & ~n9097 ;
  assign n20525 = ~n9084 & ~n20523 ;
  assign n20526 = ~n20524 & n20525 ;
  assign n20527 = n9118 & n19269 ;
  assign n20532 = ~\P1_P3_InstAddrPointer_reg[6]/NET0131  & ~n9049 ;
  assign n20533 = n9049 & ~n19327 ;
  assign n20534 = ~n20532 & ~n20533 ;
  assign n20535 = ~n9061 & n20534 ;
  assign n20536 = ~n20527 & ~n20535 ;
  assign n20537 = ~n20526 & n20536 ;
  assign n20538 = ~n20531 & n20537 ;
  assign n20539 = ~n20501 & n20538 ;
  assign n20540 = ~n20517 & n20539 ;
  assign n20541 = ~n20522 & n20540 ;
  assign n20542 = ~n20516 & n20541 ;
  assign n20543 = n9241 & ~n20542 ;
  assign n20500 = \P1_P3_rEIP_reg[6]/NET0131  & n17426 ;
  assign n20544 = \P1_P3_InstAddrPointer_reg[6]/NET0131  & ~n18343 ;
  assign n20545 = ~n20500 & ~n20544 ;
  assign n20546 = ~n20543 & n20545 ;
  assign n20549 = \P1_P3_InstAddrPointer_reg[7]/NET0131  & n9072 ;
  assign n20552 = ~n19248 & n19250 ;
  assign n20550 = ~n19300 & ~n19301 ;
  assign n20551 = n17282 & ~n20550 ;
  assign n20553 = ~n9072 & ~n20551 ;
  assign n20554 = ~n20552 & n20553 ;
  assign n20555 = ~n20549 & ~n20554 ;
  assign n20556 = n9064 & ~n20555 ;
  assign n20557 = ~n19324 & ~n19325 ;
  assign n20559 = ~n19355 & n20557 ;
  assign n20558 = n19355 & ~n20557 ;
  assign n20560 = n9191 & ~n20558 ;
  assign n20561 = ~n20559 & n20560 ;
  assign n20575 = ~n9133 & n19211 ;
  assign n20548 = \P1_P3_InstAddrPointer_reg[7]/NET0131  & ~n18435 ;
  assign n20571 = n9097 & ~n19267 ;
  assign n20570 = ~\P1_P3_InstAddrPointer_reg[7]/NET0131  & ~n9097 ;
  assign n20572 = ~n9084 & ~n20570 ;
  assign n20573 = ~n20571 & n20572 ;
  assign n20562 = ~n8741 & ~n19267 ;
  assign n20563 = ~\P1_P3_InstAddrPointer_reg[7]/NET0131  & n8741 ;
  assign n20564 = ~n20562 & ~n20563 ;
  assign n20565 = n9147 & n20564 ;
  assign n20566 = ~\P1_P3_InstAddrPointer_reg[7]/NET0131  & ~n9049 ;
  assign n20567 = n9049 & ~n19323 ;
  assign n20568 = ~n20566 & ~n20567 ;
  assign n20569 = ~n9061 & n20568 ;
  assign n20574 = n9118 & n19267 ;
  assign n20576 = ~n20569 & ~n20574 ;
  assign n20577 = ~n20565 & n20576 ;
  assign n20578 = ~n20573 & n20577 ;
  assign n20579 = ~n20548 & n20578 ;
  assign n20580 = ~n20575 & n20579 ;
  assign n20581 = ~n20561 & n20580 ;
  assign n20582 = ~n20556 & n20581 ;
  assign n20583 = n9241 & ~n20582 ;
  assign n20547 = \P1_P3_rEIP_reg[7]/NET0131  & n17426 ;
  assign n20584 = \P1_P3_InstAddrPointer_reg[7]/NET0131  & ~n18343 ;
  assign n20585 = ~n20547 & ~n20584 ;
  assign n20586 = ~n20583 & n20585 ;
  assign n20589 = \P1_P3_InstAddrPointer_reg[8]/NET0131  & n9072 ;
  assign n20593 = ~n19265 & ~n19303 ;
  assign n20594 = ~n19304 & ~n20593 ;
  assign n20595 = n17282 & ~n20594 ;
  assign n20590 = n19209 & ~n19251 ;
  assign n20591 = ~n17282 & ~n19252 ;
  assign n20592 = ~n20590 & n20591 ;
  assign n20596 = ~n9072 & ~n20592 ;
  assign n20597 = ~n20595 & n20596 ;
  assign n20598 = ~n20589 & ~n20597 ;
  assign n20599 = n9064 & ~n20598 ;
  assign n20600 = ~n19321 & n19357 ;
  assign n20601 = n9191 & ~n19358 ;
  assign n20602 = ~n20600 & n20601 ;
  assign n20607 = \P1_P3_InstAddrPointer_reg[8]/NET0131  & ~n18438 ;
  assign n20588 = ~n9133 & n19209 ;
  assign n20603 = ~n9084 & ~n19258 ;
  assign n20604 = n9176 & ~n20603 ;
  assign n20605 = n19265 & ~n20604 ;
  assign n20606 = n9220 & n19321 ;
  assign n20608 = ~n20605 & ~n20606 ;
  assign n20609 = ~n20588 & n20608 ;
  assign n20610 = ~n20607 & n20609 ;
  assign n20611 = ~n20602 & n20610 ;
  assign n20612 = ~n20599 & n20611 ;
  assign n20613 = n9241 & ~n20612 ;
  assign n20587 = \P1_P3_rEIP_reg[8]/NET0131  & n17426 ;
  assign n20614 = \P1_P3_InstAddrPointer_reg[8]/NET0131  & ~n18343 ;
  assign n20615 = ~n20587 & ~n20614 ;
  assign n20616 = ~n20613 & n20615 ;
  assign n20621 = \P1_P3_InstAddrPointer_reg[9]/NET0131  & n9072 ;
  assign n20625 = ~\P1_P3_InstAddrPointer_reg[9]/NET0131  & ~n19259 ;
  assign n20626 = ~n19260 & ~n20625 ;
  assign n20627 = ~n19304 & ~n20626 ;
  assign n20628 = ~n19305 & ~n20627 ;
  assign n20629 = n17282 & ~n20628 ;
  assign n20622 = n19207 & ~n19252 ;
  assign n20623 = ~n17282 & ~n19253 ;
  assign n20624 = ~n20622 & n20623 ;
  assign n20630 = ~n9072 & ~n20624 ;
  assign n20631 = ~n20629 & n20630 ;
  assign n20632 = ~n20621 & ~n20631 ;
  assign n20633 = n9064 & ~n20632 ;
  assign n20618 = ~\P1_P3_InstAddrPointer_reg[9]/NET0131  & ~n19320 ;
  assign n20619 = ~n19360 & ~n20618 ;
  assign n20634 = ~n19358 & ~n20619 ;
  assign n20635 = n9191 & ~n19364 ;
  assign n20636 = ~n20634 & n20635 ;
  assign n20645 = ~n9133 & n19207 ;
  assign n20637 = ~n9061 & ~n19320 ;
  assign n20638 = n18436 & ~n20637 ;
  assign n20639 = \P1_P3_InstAddrPointer_reg[9]/NET0131  & ~n20638 ;
  assign n20640 = ~\P1_P3_InstAddrPointer_reg[9]/NET0131  & ~n9097 ;
  assign n20641 = ~n9084 & ~n20640 ;
  assign n20643 = ~n9118 & ~n20641 ;
  assign n20644 = n20626 & ~n20643 ;
  assign n20646 = ~\P1_P3_InstAddrPointer_reg[9]/NET0131  & n8741 ;
  assign n20647 = ~n8741 & ~n20626 ;
  assign n20648 = ~n20646 & ~n20647 ;
  assign n20649 = n9147 & n20648 ;
  assign n20620 = n9220 & n20619 ;
  assign n20642 = ~n9097 & n20641 ;
  assign n20650 = ~n20620 & ~n20642 ;
  assign n20651 = ~n20649 & n20650 ;
  assign n20652 = ~n20644 & n20651 ;
  assign n20653 = ~n20639 & n20652 ;
  assign n20654 = ~n20645 & n20653 ;
  assign n20655 = ~n20636 & n20654 ;
  assign n20656 = ~n20633 & n20655 ;
  assign n20657 = n9241 & ~n20656 ;
  assign n20617 = \P1_P3_rEIP_reg[9]/NET0131  & n17426 ;
  assign n20658 = \P1_P3_InstAddrPointer_reg[9]/NET0131  & ~n18343 ;
  assign n20659 = ~n20617 & ~n20658 ;
  assign n20660 = ~n20657 & n20659 ;
  assign n20661 = n18658 & n18663 ;
  assign n20662 = ~n18676 & n20661 ;
  assign n20663 = n18666 & n20662 ;
  assign n20664 = \P4_reg0_reg[27]/NET0131  & ~n20663 ;
  assign n20665 = n18666 & n20661 ;
  assign n20666 = ~n18648 & n20665 ;
  assign n20667 = ~n20664 & ~n20666 ;
  assign n20668 = ~n18749 & n20665 ;
  assign n20669 = \P4_reg0_reg[28]/NET0131  & ~n20663 ;
  assign n20670 = ~n20668 & ~n20669 ;
  assign n20671 = \P4_reg2_reg[27]/NET0131  & ~n18665 ;
  assign n20672 = \P4_reg2_reg[27]/NET0131  & n19073 ;
  assign n20673 = n18658 & ~n18663 ;
  assign n20674 = ~n18482 & n20673 ;
  assign n20675 = ~\P4_reg2_reg[27]/NET0131  & ~n20673 ;
  assign n20676 = n18483 & ~n20675 ;
  assign n20677 = ~n20674 & n20676 ;
  assign n20684 = ~n18647 & n20673 ;
  assign n20678 = ~n19104 & n20673 ;
  assign n20679 = ~n19158 & ~n20678 ;
  assign n20680 = n18489 & ~n20673 ;
  assign n20681 = ~n15734 & n20680 ;
  assign n20682 = ~n20679 & ~n20681 ;
  assign n20683 = \P4_reg2_reg[27]/NET0131  & ~n20682 ;
  assign n20685 = n15805 & n16426 ;
  assign n20686 = ~n20683 & ~n20685 ;
  assign n20687 = ~n20684 & n20686 ;
  assign n20688 = ~n20677 & n20687 ;
  assign n20689 = n19075 & ~n20688 ;
  assign n20690 = ~n20672 & ~n20689 ;
  assign n20691 = \P3_rd_reg/NET0131  & ~n20690 ;
  assign n20692 = ~n20671 & ~n20691 ;
  assign n21073 = \P1_P1_ADS_n_reg/NET0131  & \P2_ready11_reg/NET0131  ;
  assign n21086 = ~n11296 & ~n21073 ;
  assign n21063 = n12378 & ~n14612 ;
  assign n21064 = ~n11689 & ~n12807 ;
  assign n21065 = n21063 & n21064 ;
  assign n21017 = n12766 & n17417 ;
  assign n21066 = ~n14068 & n21017 ;
  assign n21067 = n21065 & n21066 ;
  assign n20709 = ~\P2_P1_InstQueueRd_Addr_reg[3]/NET0131  & \P2_P1_InstQueueWr_Addr_reg[3]/NET0131  ;
  assign n20710 = \P2_P1_InstQueueRd_Addr_reg[3]/NET0131  & ~\P2_P1_InstQueueWr_Addr_reg[3]/NET0131  ;
  assign n20700 = ~\P2_P1_InstQueueRd_Addr_reg[2]/NET0131  & \P2_P1_InstQueueWr_Addr_reg[2]/NET0131  ;
  assign n20701 = \P2_P1_InstQueueRd_Addr_reg[2]/NET0131  & ~\P2_P1_InstQueueWr_Addr_reg[2]/NET0131  ;
  assign n20693 = ~\P2_P1_InstQueueRd_Addr_reg[1]/NET0131  & \P2_P1_InstQueueWr_Addr_reg[1]/NET0131  ;
  assign n20694 = \P2_P1_InstQueueRd_Addr_reg[1]/NET0131  & ~\P2_P1_InstQueueWr_Addr_reg[1]/NET0131  ;
  assign n20696 = \P2_P1_InstQueueRd_Addr_reg[0]/NET0131  & ~\P2_P1_InstQueueWr_Addr_reg[0]/NET0131  ;
  assign n20703 = ~n20694 & ~n20696 ;
  assign n20704 = ~n20693 & ~n20703 ;
  assign n20712 = ~n20701 & ~n20704 ;
  assign n20713 = ~n20700 & ~n20712 ;
  assign n20718 = ~n20710 & ~n20713 ;
  assign n20719 = ~n20709 & ~n20718 ;
  assign n20702 = ~n20700 & ~n20701 ;
  assign n20705 = n20702 & n20704 ;
  assign n20706 = ~n20702 & ~n20704 ;
  assign n20707 = ~n20705 & ~n20706 ;
  assign n20711 = ~n20709 & ~n20710 ;
  assign n20714 = n20711 & n20713 ;
  assign n20715 = ~n20711 & ~n20713 ;
  assign n20716 = ~n20714 & ~n20715 ;
  assign n21075 = n20707 & n20716 ;
  assign n21076 = ~n20719 & ~n21075 ;
  assign n20695 = ~n20693 & ~n20694 ;
  assign n21077 = n20695 & ~n20696 ;
  assign n21078 = ~n20695 & n20696 ;
  assign n21079 = ~n21077 & ~n21078 ;
  assign n21080 = ~n20719 & n21079 ;
  assign n21081 = ~n21076 & ~n21080 ;
  assign n21087 = n21067 & ~n21081 ;
  assign n21088 = ~\P2_P1_EAX_reg[31]/NET0131  & n21073 ;
  assign n21089 = n14799 & ~n21088 ;
  assign n21090 = n21087 & n21089 ;
  assign n21091 = ~n21086 & n21090 ;
  assign n21023 = \P2_P1_EAX_reg[0]/NET0131  & \P2_P1_EAX_reg[1]/NET0131  ;
  assign n21024 = \P2_P1_EAX_reg[2]/NET0131  & n21023 ;
  assign n21025 = \P2_P1_EAX_reg[3]/NET0131  & n21024 ;
  assign n21026 = \P2_P1_EAX_reg[4]/NET0131  & n21025 ;
  assign n21027 = \P2_P1_EAX_reg[5]/NET0131  & n21026 ;
  assign n21028 = \P2_P1_EAX_reg[6]/NET0131  & n21027 ;
  assign n21029 = \P2_P1_EAX_reg[7]/NET0131  & n21028 ;
  assign n21030 = \P2_P1_EAX_reg[8]/NET0131  & n21029 ;
  assign n21031 = \P2_P1_EAX_reg[9]/NET0131  & n21030 ;
  assign n21032 = \P2_P1_EAX_reg[10]/NET0131  & n21031 ;
  assign n21033 = \P2_P1_EAX_reg[11]/NET0131  & n21032 ;
  assign n21034 = \P2_P1_EAX_reg[12]/NET0131  & n21033 ;
  assign n21035 = \P2_P1_EAX_reg[13]/NET0131  & n21034 ;
  assign n21036 = \P2_P1_EAX_reg[14]/NET0131  & n21035 ;
  assign n21037 = \P2_P1_EAX_reg[15]/NET0131  & n21036 ;
  assign n21038 = \P2_P1_EAX_reg[16]/NET0131  & n21037 ;
  assign n21039 = \P2_P1_EAX_reg[17]/NET0131  & n21038 ;
  assign n21040 = \P2_P1_EAX_reg[18]/NET0131  & n21039 ;
  assign n21041 = \P2_P1_EAX_reg[19]/NET0131  & n21040 ;
  assign n21042 = \P2_P1_EAX_reg[20]/NET0131  & n21041 ;
  assign n21043 = \P2_P1_EAX_reg[21]/NET0131  & n21042 ;
  assign n21044 = \P2_P1_EAX_reg[22]/NET0131  & n21043 ;
  assign n21045 = \P2_P1_EAX_reg[23]/NET0131  & n21044 ;
  assign n21046 = \P2_P1_EAX_reg[24]/NET0131  & n21045 ;
  assign n21047 = \P2_P1_EAX_reg[25]/NET0131  & n21046 ;
  assign n21048 = \P2_P1_EAX_reg[26]/NET0131  & n21047 ;
  assign n21049 = \P2_P1_EAX_reg[27]/NET0131  & n21048 ;
  assign n21050 = \P2_P1_EAX_reg[28]/NET0131  & n21049 ;
  assign n21051 = \P2_P1_EAX_reg[29]/NET0131  & n21050 ;
  assign n21052 = \P2_P1_EAX_reg[30]/NET0131  & n21051 ;
  assign n21054 = \P2_P1_EAX_reg[31]/NET0131  & n21052 ;
  assign n20722 = n14068 & n14799 ;
  assign n21018 = n20722 & n21017 ;
  assign n21019 = n12378 & n14612 ;
  assign n21020 = n11689 & ~n12807 ;
  assign n21021 = n21019 & n21020 ;
  assign n21022 = n21018 & n21021 ;
  assign n21053 = ~\P2_P1_EAX_reg[31]/NET0131  & ~n21052 ;
  assign n21055 = n21022 & ~n21053 ;
  assign n21056 = ~n21054 & n21055 ;
  assign n20697 = ~\P2_P1_InstQueueRd_Addr_reg[0]/NET0131  & \P2_P1_InstQueueWr_Addr_reg[0]/NET0131  ;
  assign n20698 = ~n20696 & ~n20697 ;
  assign n20699 = n20695 & n20698 ;
  assign n20708 = ~n20699 & ~n20707 ;
  assign n20717 = ~n20708 & n20716 ;
  assign n20720 = ~n20717 & ~n20719 ;
  assign n20723 = ~n11689 & ~n12378 ;
  assign n20724 = n12807 & n20723 ;
  assign n20725 = ~n14612 & n20724 ;
  assign n20721 = ~n12766 & n17417 ;
  assign n20726 = n20721 & n20722 ;
  assign n20727 = n20725 & n20726 ;
  assign n20728 = n20720 & n20727 ;
  assign n20734 = \P2_P1_InstQueue_reg[9][7]/NET0131  & n11651 ;
  assign n20733 = \P2_P1_InstQueue_reg[2][7]/NET0131  & n11647 ;
  assign n20729 = \P2_P1_InstQueue_reg[14][7]/NET0131  & n11665 ;
  assign n20730 = \P2_P1_InstQueue_reg[3][7]/NET0131  & n11669 ;
  assign n20745 = ~n20729 & ~n20730 ;
  assign n20755 = ~n20733 & n20745 ;
  assign n20756 = ~n20734 & n20755 ;
  assign n20741 = \P2_P1_InstQueue_reg[0][7]/NET0131  & n11641 ;
  assign n20742 = \P2_P1_InstQueue_reg[8][7]/NET0131  & n11638 ;
  assign n20750 = ~n20741 & ~n20742 ;
  assign n20743 = \P2_P1_InstQueue_reg[15][7]/NET0131  & n11673 ;
  assign n20744 = \P2_P1_InstQueue_reg[13][7]/NET0131  & n11634 ;
  assign n20751 = ~n20743 & ~n20744 ;
  assign n20752 = n20750 & n20751 ;
  assign n20737 = \P2_P1_InstQueue_reg[4][7]/NET0131  & n11671 ;
  assign n20738 = \P2_P1_InstQueue_reg[10][7]/NET0131  & n11661 ;
  assign n20748 = ~n20737 & ~n20738 ;
  assign n20739 = \P2_P1_InstQueue_reg[12][7]/NET0131  & n11656 ;
  assign n20740 = \P2_P1_InstQueue_reg[7][7]/NET0131  & n11667 ;
  assign n20749 = ~n20739 & ~n20740 ;
  assign n20753 = n20748 & n20749 ;
  assign n20731 = \P2_P1_InstQueue_reg[6][7]/NET0131  & n11663 ;
  assign n20732 = \P2_P1_InstQueue_reg[1][7]/NET0131  & n11643 ;
  assign n20746 = ~n20731 & ~n20732 ;
  assign n20735 = \P2_P1_InstQueue_reg[11][7]/NET0131  & n11659 ;
  assign n20736 = \P2_P1_InstQueue_reg[5][7]/NET0131  & n11654 ;
  assign n20747 = ~n20735 & ~n20736 ;
  assign n20754 = n20746 & n20747 ;
  assign n20757 = n20753 & n20754 ;
  assign n20758 = n20752 & n20757 ;
  assign n20759 = n20756 & n20758 ;
  assign n20765 = \P2_P1_InstQueue_reg[10][0]/NET0131  & n11651 ;
  assign n20764 = \P2_P1_InstQueue_reg[3][0]/NET0131  & n11647 ;
  assign n20760 = \P2_P1_InstQueue_reg[5][0]/NET0131  & n11671 ;
  assign n20761 = \P2_P1_InstQueue_reg[1][0]/NET0131  & n11641 ;
  assign n20776 = ~n20760 & ~n20761 ;
  assign n20786 = ~n20764 & n20776 ;
  assign n20787 = ~n20765 & n20786 ;
  assign n20772 = \P2_P1_InstQueue_reg[9][0]/NET0131  & n11638 ;
  assign n20773 = \P2_P1_InstQueue_reg[7][0]/NET0131  & n11663 ;
  assign n20781 = ~n20772 & ~n20773 ;
  assign n20774 = \P2_P1_InstQueue_reg[4][0]/NET0131  & n11669 ;
  assign n20775 = \P2_P1_InstQueue_reg[12][0]/NET0131  & n11659 ;
  assign n20782 = ~n20774 & ~n20775 ;
  assign n20783 = n20781 & n20782 ;
  assign n20768 = \P2_P1_InstQueue_reg[8][0]/NET0131  & n11667 ;
  assign n20769 = \P2_P1_InstQueue_reg[11][0]/NET0131  & n11661 ;
  assign n20779 = ~n20768 & ~n20769 ;
  assign n20770 = \P2_P1_InstQueue_reg[0][0]/NET0131  & n11673 ;
  assign n20771 = \P2_P1_InstQueue_reg[15][0]/NET0131  & n11665 ;
  assign n20780 = ~n20770 & ~n20771 ;
  assign n20784 = n20779 & n20780 ;
  assign n20762 = \P2_P1_InstQueue_reg[6][0]/NET0131  & n11654 ;
  assign n20763 = \P2_P1_InstQueue_reg[2][0]/NET0131  & n11643 ;
  assign n20777 = ~n20762 & ~n20763 ;
  assign n20766 = \P2_P1_InstQueue_reg[13][0]/NET0131  & n11656 ;
  assign n20767 = \P2_P1_InstQueue_reg[14][0]/NET0131  & n11634 ;
  assign n20778 = ~n20766 & ~n20767 ;
  assign n20785 = n20777 & n20778 ;
  assign n20788 = n20784 & n20785 ;
  assign n20789 = n20783 & n20788 ;
  assign n20790 = n20787 & n20789 ;
  assign n20791 = ~n20759 & ~n20790 ;
  assign n20797 = \P2_P1_InstQueue_reg[10][1]/NET0131  & n11651 ;
  assign n20796 = \P2_P1_InstQueue_reg[3][1]/NET0131  & n11647 ;
  assign n20792 = \P2_P1_InstQueue_reg[5][1]/NET0131  & n11671 ;
  assign n20793 = \P2_P1_InstQueue_reg[1][1]/NET0131  & n11641 ;
  assign n20808 = ~n20792 & ~n20793 ;
  assign n20818 = ~n20796 & n20808 ;
  assign n20819 = ~n20797 & n20818 ;
  assign n20804 = \P2_P1_InstQueue_reg[9][1]/NET0131  & n11638 ;
  assign n20805 = \P2_P1_InstQueue_reg[7][1]/NET0131  & n11663 ;
  assign n20813 = ~n20804 & ~n20805 ;
  assign n20806 = \P2_P1_InstQueue_reg[4][1]/NET0131  & n11669 ;
  assign n20807 = \P2_P1_InstQueue_reg[12][1]/NET0131  & n11659 ;
  assign n20814 = ~n20806 & ~n20807 ;
  assign n20815 = n20813 & n20814 ;
  assign n20800 = \P2_P1_InstQueue_reg[8][1]/NET0131  & n11667 ;
  assign n20801 = \P2_P1_InstQueue_reg[11][1]/NET0131  & n11661 ;
  assign n20811 = ~n20800 & ~n20801 ;
  assign n20802 = \P2_P1_InstQueue_reg[0][1]/NET0131  & n11673 ;
  assign n20803 = \P2_P1_InstQueue_reg[15][1]/NET0131  & n11665 ;
  assign n20812 = ~n20802 & ~n20803 ;
  assign n20816 = n20811 & n20812 ;
  assign n20794 = \P2_P1_InstQueue_reg[6][1]/NET0131  & n11654 ;
  assign n20795 = \P2_P1_InstQueue_reg[2][1]/NET0131  & n11643 ;
  assign n20809 = ~n20794 & ~n20795 ;
  assign n20798 = \P2_P1_InstQueue_reg[13][1]/NET0131  & n11656 ;
  assign n20799 = \P2_P1_InstQueue_reg[14][1]/NET0131  & n11634 ;
  assign n20810 = ~n20798 & ~n20799 ;
  assign n20817 = n20809 & n20810 ;
  assign n20820 = n20816 & n20817 ;
  assign n20821 = n20815 & n20820 ;
  assign n20822 = n20819 & n20821 ;
  assign n20823 = n20791 & ~n20822 ;
  assign n20829 = \P2_P1_InstQueue_reg[10][2]/NET0131  & n11651 ;
  assign n20828 = \P2_P1_InstQueue_reg[3][2]/NET0131  & n11647 ;
  assign n20824 = \P2_P1_InstQueue_reg[5][2]/NET0131  & n11671 ;
  assign n20825 = \P2_P1_InstQueue_reg[1][2]/NET0131  & n11641 ;
  assign n20840 = ~n20824 & ~n20825 ;
  assign n20850 = ~n20828 & n20840 ;
  assign n20851 = ~n20829 & n20850 ;
  assign n20836 = \P2_P1_InstQueue_reg[9][2]/NET0131  & n11638 ;
  assign n20837 = \P2_P1_InstQueue_reg[7][2]/NET0131  & n11663 ;
  assign n20845 = ~n20836 & ~n20837 ;
  assign n20838 = \P2_P1_InstQueue_reg[4][2]/NET0131  & n11669 ;
  assign n20839 = \P2_P1_InstQueue_reg[12][2]/NET0131  & n11659 ;
  assign n20846 = ~n20838 & ~n20839 ;
  assign n20847 = n20845 & n20846 ;
  assign n20832 = \P2_P1_InstQueue_reg[8][2]/NET0131  & n11667 ;
  assign n20833 = \P2_P1_InstQueue_reg[11][2]/NET0131  & n11661 ;
  assign n20843 = ~n20832 & ~n20833 ;
  assign n20834 = \P2_P1_InstQueue_reg[0][2]/NET0131  & n11673 ;
  assign n20835 = \P2_P1_InstQueue_reg[15][2]/NET0131  & n11665 ;
  assign n20844 = ~n20834 & ~n20835 ;
  assign n20848 = n20843 & n20844 ;
  assign n20826 = \P2_P1_InstQueue_reg[6][2]/NET0131  & n11654 ;
  assign n20827 = \P2_P1_InstQueue_reg[2][2]/NET0131  & n11643 ;
  assign n20841 = ~n20826 & ~n20827 ;
  assign n20830 = \P2_P1_InstQueue_reg[13][2]/NET0131  & n11656 ;
  assign n20831 = \P2_P1_InstQueue_reg[14][2]/NET0131  & n11634 ;
  assign n20842 = ~n20830 & ~n20831 ;
  assign n20849 = n20841 & n20842 ;
  assign n20852 = n20848 & n20849 ;
  assign n20853 = n20847 & n20852 ;
  assign n20854 = n20851 & n20853 ;
  assign n20855 = n20823 & ~n20854 ;
  assign n20861 = \P2_P1_InstQueue_reg[10][3]/NET0131  & n11651 ;
  assign n20860 = \P2_P1_InstQueue_reg[3][3]/NET0131  & n11647 ;
  assign n20856 = \P2_P1_InstQueue_reg[5][3]/NET0131  & n11671 ;
  assign n20857 = \P2_P1_InstQueue_reg[1][3]/NET0131  & n11641 ;
  assign n20872 = ~n20856 & ~n20857 ;
  assign n20882 = ~n20860 & n20872 ;
  assign n20883 = ~n20861 & n20882 ;
  assign n20868 = \P2_P1_InstQueue_reg[9][3]/NET0131  & n11638 ;
  assign n20869 = \P2_P1_InstQueue_reg[7][3]/NET0131  & n11663 ;
  assign n20877 = ~n20868 & ~n20869 ;
  assign n20870 = \P2_P1_InstQueue_reg[4][3]/NET0131  & n11669 ;
  assign n20871 = \P2_P1_InstQueue_reg[12][3]/NET0131  & n11659 ;
  assign n20878 = ~n20870 & ~n20871 ;
  assign n20879 = n20877 & n20878 ;
  assign n20864 = \P2_P1_InstQueue_reg[8][3]/NET0131  & n11667 ;
  assign n20865 = \P2_P1_InstQueue_reg[11][3]/NET0131  & n11661 ;
  assign n20875 = ~n20864 & ~n20865 ;
  assign n20866 = \P2_P1_InstQueue_reg[0][3]/NET0131  & n11673 ;
  assign n20867 = \P2_P1_InstQueue_reg[15][3]/NET0131  & n11665 ;
  assign n20876 = ~n20866 & ~n20867 ;
  assign n20880 = n20875 & n20876 ;
  assign n20858 = \P2_P1_InstQueue_reg[6][3]/NET0131  & n11654 ;
  assign n20859 = \P2_P1_InstQueue_reg[2][3]/NET0131  & n11643 ;
  assign n20873 = ~n20858 & ~n20859 ;
  assign n20862 = \P2_P1_InstQueue_reg[13][3]/NET0131  & n11656 ;
  assign n20863 = \P2_P1_InstQueue_reg[14][3]/NET0131  & n11634 ;
  assign n20874 = ~n20862 & ~n20863 ;
  assign n20881 = n20873 & n20874 ;
  assign n20884 = n20880 & n20881 ;
  assign n20885 = n20879 & n20884 ;
  assign n20886 = n20883 & n20885 ;
  assign n20887 = n20855 & ~n20886 ;
  assign n20893 = \P2_P1_InstQueue_reg[10][4]/NET0131  & n11651 ;
  assign n20892 = \P2_P1_InstQueue_reg[3][4]/NET0131  & n11647 ;
  assign n20888 = \P2_P1_InstQueue_reg[5][4]/NET0131  & n11671 ;
  assign n20889 = \P2_P1_InstQueue_reg[1][4]/NET0131  & n11641 ;
  assign n20904 = ~n20888 & ~n20889 ;
  assign n20914 = ~n20892 & n20904 ;
  assign n20915 = ~n20893 & n20914 ;
  assign n20900 = \P2_P1_InstQueue_reg[9][4]/NET0131  & n11638 ;
  assign n20901 = \P2_P1_InstQueue_reg[7][4]/NET0131  & n11663 ;
  assign n20909 = ~n20900 & ~n20901 ;
  assign n20902 = \P2_P1_InstQueue_reg[4][4]/NET0131  & n11669 ;
  assign n20903 = \P2_P1_InstQueue_reg[12][4]/NET0131  & n11659 ;
  assign n20910 = ~n20902 & ~n20903 ;
  assign n20911 = n20909 & n20910 ;
  assign n20896 = \P2_P1_InstQueue_reg[8][4]/NET0131  & n11667 ;
  assign n20897 = \P2_P1_InstQueue_reg[11][4]/NET0131  & n11661 ;
  assign n20907 = ~n20896 & ~n20897 ;
  assign n20898 = \P2_P1_InstQueue_reg[0][4]/NET0131  & n11673 ;
  assign n20899 = \P2_P1_InstQueue_reg[15][4]/NET0131  & n11665 ;
  assign n20908 = ~n20898 & ~n20899 ;
  assign n20912 = n20907 & n20908 ;
  assign n20890 = \P2_P1_InstQueue_reg[6][4]/NET0131  & n11654 ;
  assign n20891 = \P2_P1_InstQueue_reg[2][4]/NET0131  & n11643 ;
  assign n20905 = ~n20890 & ~n20891 ;
  assign n20894 = \P2_P1_InstQueue_reg[13][4]/NET0131  & n11656 ;
  assign n20895 = \P2_P1_InstQueue_reg[14][4]/NET0131  & n11634 ;
  assign n20906 = ~n20894 & ~n20895 ;
  assign n20913 = n20905 & n20906 ;
  assign n20916 = n20912 & n20913 ;
  assign n20917 = n20911 & n20916 ;
  assign n20918 = n20915 & n20917 ;
  assign n20919 = n20887 & ~n20918 ;
  assign n20925 = \P2_P1_InstQueue_reg[10][5]/NET0131  & n11651 ;
  assign n20924 = \P2_P1_InstQueue_reg[3][5]/NET0131  & n11647 ;
  assign n20920 = \P2_P1_InstQueue_reg[1][5]/NET0131  & n11641 ;
  assign n20921 = \P2_P1_InstQueue_reg[8][5]/NET0131  & n11667 ;
  assign n20936 = ~n20920 & ~n20921 ;
  assign n20946 = ~n20924 & n20936 ;
  assign n20947 = ~n20925 & n20946 ;
  assign n20932 = \P2_P1_InstQueue_reg[14][5]/NET0131  & n11634 ;
  assign n20933 = \P2_P1_InstQueue_reg[4][5]/NET0131  & n11669 ;
  assign n20941 = ~n20932 & ~n20933 ;
  assign n20934 = \P2_P1_InstQueue_reg[5][5]/NET0131  & n11671 ;
  assign n20935 = \P2_P1_InstQueue_reg[12][5]/NET0131  & n11659 ;
  assign n20942 = ~n20934 & ~n20935 ;
  assign n20943 = n20941 & n20942 ;
  assign n20928 = \P2_P1_InstQueue_reg[9][5]/NET0131  & n11638 ;
  assign n20929 = \P2_P1_InstQueue_reg[11][5]/NET0131  & n11661 ;
  assign n20939 = ~n20928 & ~n20929 ;
  assign n20930 = \P2_P1_InstQueue_reg[6][5]/NET0131  & n11654 ;
  assign n20931 = \P2_P1_InstQueue_reg[15][5]/NET0131  & n11665 ;
  assign n20940 = ~n20930 & ~n20931 ;
  assign n20944 = n20939 & n20940 ;
  assign n20922 = \P2_P1_InstQueue_reg[7][5]/NET0131  & n11663 ;
  assign n20923 = \P2_P1_InstQueue_reg[2][5]/NET0131  & n11643 ;
  assign n20937 = ~n20922 & ~n20923 ;
  assign n20926 = \P2_P1_InstQueue_reg[13][5]/NET0131  & n11656 ;
  assign n20927 = \P2_P1_InstQueue_reg[0][5]/NET0131  & n11673 ;
  assign n20938 = ~n20926 & ~n20927 ;
  assign n20945 = n20937 & n20938 ;
  assign n20948 = n20944 & n20945 ;
  assign n20949 = n20943 & n20948 ;
  assign n20950 = n20947 & n20949 ;
  assign n20951 = n20919 & ~n20950 ;
  assign n20957 = \P2_P1_InstQueue_reg[10][6]/NET0131  & n11651 ;
  assign n20956 = \P2_P1_InstQueue_reg[3][6]/NET0131  & n11647 ;
  assign n20952 = \P2_P1_InstQueue_reg[1][6]/NET0131  & n11641 ;
  assign n20953 = \P2_P1_InstQueue_reg[8][6]/NET0131  & n11667 ;
  assign n20968 = ~n20952 & ~n20953 ;
  assign n20978 = ~n20956 & n20968 ;
  assign n20979 = ~n20957 & n20978 ;
  assign n20964 = \P2_P1_InstQueue_reg[14][6]/NET0131  & n11634 ;
  assign n20965 = \P2_P1_InstQueue_reg[4][6]/NET0131  & n11669 ;
  assign n20973 = ~n20964 & ~n20965 ;
  assign n20966 = \P2_P1_InstQueue_reg[5][6]/NET0131  & n11671 ;
  assign n20967 = \P2_P1_InstQueue_reg[12][6]/NET0131  & n11659 ;
  assign n20974 = ~n20966 & ~n20967 ;
  assign n20975 = n20973 & n20974 ;
  assign n20960 = \P2_P1_InstQueue_reg[9][6]/NET0131  & n11638 ;
  assign n20961 = \P2_P1_InstQueue_reg[11][6]/NET0131  & n11661 ;
  assign n20971 = ~n20960 & ~n20961 ;
  assign n20962 = \P2_P1_InstQueue_reg[6][6]/NET0131  & n11654 ;
  assign n20963 = \P2_P1_InstQueue_reg[15][6]/NET0131  & n11665 ;
  assign n20972 = ~n20962 & ~n20963 ;
  assign n20976 = n20971 & n20972 ;
  assign n20954 = \P2_P1_InstQueue_reg[7][6]/NET0131  & n11663 ;
  assign n20955 = \P2_P1_InstQueue_reg[2][6]/NET0131  & n11643 ;
  assign n20969 = ~n20954 & ~n20955 ;
  assign n20958 = \P2_P1_InstQueue_reg[13][6]/NET0131  & n11656 ;
  assign n20959 = \P2_P1_InstQueue_reg[0][6]/NET0131  & n11673 ;
  assign n20970 = ~n20958 & ~n20959 ;
  assign n20977 = n20969 & n20970 ;
  assign n20980 = n20976 & n20977 ;
  assign n20981 = n20975 & n20980 ;
  assign n20982 = n20979 & n20981 ;
  assign n20983 = n20951 & ~n20982 ;
  assign n20989 = \P2_P1_InstQueue_reg[10][7]/NET0131  & n11651 ;
  assign n20988 = \P2_P1_InstQueue_reg[3][7]/NET0131  & n11647 ;
  assign n20984 = \P2_P1_InstQueue_reg[15][7]/NET0131  & n11665 ;
  assign n20985 = \P2_P1_InstQueue_reg[7][7]/NET0131  & n11663 ;
  assign n21000 = ~n20984 & ~n20985 ;
  assign n21010 = ~n20988 & n21000 ;
  assign n21011 = ~n20989 & n21010 ;
  assign n20996 = \P2_P1_InstQueue_reg[12][7]/NET0131  & n11659 ;
  assign n20997 = \P2_P1_InstQueue_reg[5][7]/NET0131  & n11671 ;
  assign n21005 = ~n20996 & ~n20997 ;
  assign n20998 = \P2_P1_InstQueue_reg[1][7]/NET0131  & n11641 ;
  assign n20999 = \P2_P1_InstQueue_reg[8][7]/NET0131  & n11667 ;
  assign n21006 = ~n20998 & ~n20999 ;
  assign n21007 = n21005 & n21006 ;
  assign n20992 = \P2_P1_InstQueue_reg[6][7]/NET0131  & n11654 ;
  assign n20993 = \P2_P1_InstQueue_reg[11][7]/NET0131  & n11661 ;
  assign n21003 = ~n20992 & ~n20993 ;
  assign n20994 = \P2_P1_InstQueue_reg[9][7]/NET0131  & n11638 ;
  assign n20995 = \P2_P1_InstQueue_reg[4][7]/NET0131  & n11669 ;
  assign n21004 = ~n20994 & ~n20995 ;
  assign n21008 = n21003 & n21004 ;
  assign n20986 = \P2_P1_InstQueue_reg[0][7]/NET0131  & n11673 ;
  assign n20987 = \P2_P1_InstQueue_reg[2][7]/NET0131  & n11643 ;
  assign n21001 = ~n20986 & ~n20987 ;
  assign n20990 = \P2_P1_InstQueue_reg[14][7]/NET0131  & n11634 ;
  assign n20991 = \P2_P1_InstQueue_reg[13][7]/NET0131  & n11656 ;
  assign n21002 = ~n20990 & ~n20991 ;
  assign n21009 = n21001 & n21002 ;
  assign n21012 = n21008 & n21009 ;
  assign n21013 = n21007 & n21012 ;
  assign n21014 = n21011 & n21013 ;
  assign n21015 = n20983 & ~n21014 ;
  assign n21016 = n20728 & n21015 ;
  assign n21057 = ~n12766 & ~n17417 ;
  assign n21058 = n14068 & ~n14799 ;
  assign n21059 = n21057 & n21058 ;
  assign n21060 = n12807 & n21019 ;
  assign n21061 = ~n11689 & n21060 ;
  assign n21062 = n21059 & n21061 ;
  assign n21068 = n14799 & n21067 ;
  assign n21069 = ~n21062 & ~n21068 ;
  assign n21070 = ~n21022 & n21069 ;
  assign n21071 = ~n20727 & ~n21070 ;
  assign n21072 = ~n20728 & ~n21071 ;
  assign n21074 = n21062 & n21073 ;
  assign n21082 = ~n21069 & n21081 ;
  assign n21083 = ~n21074 & ~n21082 ;
  assign n21084 = ~n21072 & n21083 ;
  assign n21085 = \P2_P1_EAX_reg[31]/NET0131  & ~n21084 ;
  assign n21092 = ~n21016 & ~n21085 ;
  assign n21093 = ~n21056 & n21092 ;
  assign n21094 = ~n21091 & n21093 ;
  assign n21095 = n11623 & ~n21094 ;
  assign n21096 = \P2_P1_State2_reg[0]/NET0131  & n11621 ;
  assign n21097 = ~n11624 & ~n21096 ;
  assign n21098 = ~\P2_P1_State2_reg[2]/NET0131  & n11622 ;
  assign n21099 = ~n11611 & ~n21098 ;
  assign n21100 = n21097 & n21099 ;
  assign n21101 = \P2_P1_EAX_reg[31]/NET0131  & ~n21100 ;
  assign n21102 = ~n21095 & ~n21101 ;
  assign n21103 = \P1_P3_EAX_reg[0]/NET0131  & ~n17031 ;
  assign n21104 = \P1_buf2_reg[0]/NET0131  & n9175 ;
  assign n21105 = n16984 & ~n18409 ;
  assign n21106 = ~\P1_P3_EAX_reg[0]/NET0131  & n16982 ;
  assign n21107 = ~n21105 & ~n21106 ;
  assign n21108 = ~n21104 & n21107 ;
  assign n21109 = n9241 & ~n21108 ;
  assign n21110 = ~n21103 & ~n21109 ;
  assign n21111 = \P1_P3_EAX_reg[17]/NET0131  & ~n16968 ;
  assign n21113 = n16982 & ~n18812 ;
  assign n21114 = ~n16987 & ~n21113 ;
  assign n21115 = \P1_P3_EAX_reg[17]/NET0131  & ~n21114 ;
  assign n21112 = n18812 & n18814 ;
  assign n21148 = \P1_P3_EAX_reg[17]/NET0131  & ~n9088 ;
  assign n21151 = \P1_buf2_reg[17]/NET0131  & n9088 ;
  assign n21152 = ~n21148 & ~n21151 ;
  assign n21153 = n9086 & ~n21152 ;
  assign n21120 = \P1_P3_InstQueue_reg[6][1]/NET0131  & n8771 ;
  assign n21121 = \P1_P3_InstQueue_reg[14][1]/NET0131  & n8765 ;
  assign n21134 = ~n21120 & ~n21121 ;
  assign n21122 = \P1_P3_InstQueue_reg[11][1]/NET0131  & n8769 ;
  assign n21123 = \P1_P3_InstQueue_reg[5][1]/NET0131  & n8752 ;
  assign n21135 = ~n21122 & ~n21123 ;
  assign n21142 = n21134 & n21135 ;
  assign n21116 = \P1_P3_InstQueue_reg[4][1]/NET0131  & n8777 ;
  assign n21117 = \P1_P3_InstQueue_reg[10][1]/NET0131  & n8748 ;
  assign n21132 = ~n21116 & ~n21117 ;
  assign n21118 = \P1_P3_InstQueue_reg[0][1]/NET0131  & n8775 ;
  assign n21119 = \P1_P3_InstQueue_reg[8][1]/NET0131  & n8779 ;
  assign n21133 = ~n21118 & ~n21119 ;
  assign n21143 = n21132 & n21133 ;
  assign n21144 = n21142 & n21143 ;
  assign n21128 = \P1_P3_InstQueue_reg[13][1]/NET0131  & n8757 ;
  assign n21129 = \P1_P3_InstQueue_reg[12][1]/NET0131  & n8763 ;
  assign n21138 = ~n21128 & ~n21129 ;
  assign n21130 = \P1_P3_InstQueue_reg[7][1]/NET0131  & n8745 ;
  assign n21131 = \P1_P3_InstQueue_reg[1][1]/NET0131  & n8781 ;
  assign n21139 = ~n21130 & ~n21131 ;
  assign n21140 = n21138 & n21139 ;
  assign n21124 = \P1_P3_InstQueue_reg[15][1]/NET0131  & n8760 ;
  assign n21125 = \P1_P3_InstQueue_reg[3][1]/NET0131  & n8767 ;
  assign n21136 = ~n21124 & ~n21125 ;
  assign n21126 = \P1_P3_InstQueue_reg[9][1]/NET0131  & n8754 ;
  assign n21127 = \P1_P3_InstQueue_reg[2][1]/NET0131  & n8773 ;
  assign n21137 = ~n21126 & ~n21127 ;
  assign n21141 = n21136 & n21137 ;
  assign n21145 = n21140 & n21141 ;
  assign n21146 = n21144 & n21145 ;
  assign n21147 = n16984 & ~n21146 ;
  assign n21149 = ~n18802 & ~n21148 ;
  assign n21150 = n9085 & ~n21149 ;
  assign n21154 = ~n21147 & ~n21150 ;
  assign n21155 = ~n21153 & n21154 ;
  assign n21156 = ~n21112 & n21155 ;
  assign n21157 = ~n21115 & n21156 ;
  assign n21158 = n9241 & ~n21157 ;
  assign n21159 = ~n21111 & ~n21158 ;
  assign n21161 = \P1_P3_EAX_reg[18]/NET0131  & n18813 ;
  assign n21162 = \P1_P3_EAX_reg[19]/NET0131  & n21161 ;
  assign n21163 = n16982 & ~n21162 ;
  assign n21164 = ~\P1_P3_EAX_reg[19]/NET0131  & ~n21161 ;
  assign n21165 = n21163 & ~n21164 ;
  assign n21160 = \P1_P3_EAX_reg[19]/NET0131  & ~n16988 ;
  assign n21166 = \P1_buf2_reg[19]/NET0131  & n9086 ;
  assign n21167 = \P1_buf2_reg[3]/NET0131  & n9085 ;
  assign n21168 = ~n21166 & ~n21167 ;
  assign n21169 = n9088 & ~n21168 ;
  assign n21174 = \P1_P3_InstQueue_reg[8][3]/NET0131  & n8779 ;
  assign n21175 = \P1_P3_InstQueue_reg[9][3]/NET0131  & n8754 ;
  assign n21188 = ~n21174 & ~n21175 ;
  assign n21176 = \P1_P3_InstQueue_reg[15][3]/NET0131  & n8760 ;
  assign n21177 = \P1_P3_InstQueue_reg[14][3]/NET0131  & n8765 ;
  assign n21189 = ~n21176 & ~n21177 ;
  assign n21196 = n21188 & n21189 ;
  assign n21170 = \P1_P3_InstQueue_reg[7][3]/NET0131  & n8745 ;
  assign n21171 = \P1_P3_InstQueue_reg[10][3]/NET0131  & n8748 ;
  assign n21186 = ~n21170 & ~n21171 ;
  assign n21172 = \P1_P3_InstQueue_reg[5][3]/NET0131  & n8752 ;
  assign n21173 = \P1_P3_InstQueue_reg[6][3]/NET0131  & n8771 ;
  assign n21187 = ~n21172 & ~n21173 ;
  assign n21197 = n21186 & n21187 ;
  assign n21198 = n21196 & n21197 ;
  assign n21182 = \P1_P3_InstQueue_reg[4][3]/NET0131  & n8777 ;
  assign n21183 = \P1_P3_InstQueue_reg[0][3]/NET0131  & n8775 ;
  assign n21192 = ~n21182 & ~n21183 ;
  assign n21184 = \P1_P3_InstQueue_reg[3][3]/NET0131  & n8767 ;
  assign n21185 = \P1_P3_InstQueue_reg[1][3]/NET0131  & n8781 ;
  assign n21193 = ~n21184 & ~n21185 ;
  assign n21194 = n21192 & n21193 ;
  assign n21178 = \P1_P3_InstQueue_reg[12][3]/NET0131  & n8763 ;
  assign n21179 = \P1_P3_InstQueue_reg[11][3]/NET0131  & n8769 ;
  assign n21190 = ~n21178 & ~n21179 ;
  assign n21180 = \P1_P3_InstQueue_reg[13][3]/NET0131  & n8757 ;
  assign n21181 = \P1_P3_InstQueue_reg[2][3]/NET0131  & n8773 ;
  assign n21191 = ~n21180 & ~n21181 ;
  assign n21195 = n21190 & n21191 ;
  assign n21199 = n21194 & n21195 ;
  assign n21200 = n21198 & n21199 ;
  assign n21201 = n16984 & ~n21200 ;
  assign n21202 = ~n21169 & ~n21201 ;
  assign n21203 = ~n21160 & n21202 ;
  assign n21204 = ~n21165 & n21203 ;
  assign n21205 = n9241 & ~n21204 ;
  assign n21206 = \P1_P3_EAX_reg[19]/NET0131  & ~n16968 ;
  assign n21207 = ~n21205 & ~n21206 ;
  assign n21208 = \P1_P3_EAX_reg[20]/NET0131  & ~n17077 ;
  assign n21209 = ~n9089 & ~n21163 ;
  assign n21210 = \P1_P3_EAX_reg[20]/NET0131  & ~n21209 ;
  assign n21211 = ~\P1_P3_EAX_reg[20]/NET0131  & n16982 ;
  assign n21212 = n21162 & n21211 ;
  assign n21217 = \P1_P3_InstQueue_reg[12][4]/NET0131  & n8763 ;
  assign n21218 = \P1_P3_InstQueue_reg[11][4]/NET0131  & n8769 ;
  assign n21231 = ~n21217 & ~n21218 ;
  assign n21219 = \P1_P3_InstQueue_reg[7][4]/NET0131  & n8745 ;
  assign n21220 = \P1_P3_InstQueue_reg[6][4]/NET0131  & n8771 ;
  assign n21232 = ~n21219 & ~n21220 ;
  assign n21239 = n21231 & n21232 ;
  assign n21213 = \P1_P3_InstQueue_reg[3][4]/NET0131  & n8767 ;
  assign n21214 = \P1_P3_InstQueue_reg[10][4]/NET0131  & n8748 ;
  assign n21229 = ~n21213 & ~n21214 ;
  assign n21215 = \P1_P3_InstQueue_reg[8][4]/NET0131  & n8779 ;
  assign n21216 = \P1_P3_InstQueue_reg[13][4]/NET0131  & n8757 ;
  assign n21230 = ~n21215 & ~n21216 ;
  assign n21240 = n21229 & n21230 ;
  assign n21241 = n21239 & n21240 ;
  assign n21225 = \P1_P3_InstQueue_reg[0][4]/NET0131  & n8775 ;
  assign n21226 = \P1_P3_InstQueue_reg[4][4]/NET0131  & n8777 ;
  assign n21235 = ~n21225 & ~n21226 ;
  assign n21227 = \P1_P3_InstQueue_reg[5][4]/NET0131  & n8752 ;
  assign n21228 = \P1_P3_InstQueue_reg[1][4]/NET0131  & n8781 ;
  assign n21236 = ~n21227 & ~n21228 ;
  assign n21237 = n21235 & n21236 ;
  assign n21221 = \P1_P3_InstQueue_reg[14][4]/NET0131  & n8765 ;
  assign n21222 = \P1_P3_InstQueue_reg[9][4]/NET0131  & n8754 ;
  assign n21233 = ~n21221 & ~n21222 ;
  assign n21223 = \P1_P3_InstQueue_reg[15][4]/NET0131  & n8760 ;
  assign n21224 = \P1_P3_InstQueue_reg[2][4]/NET0131  & n8773 ;
  assign n21234 = ~n21223 & ~n21224 ;
  assign n21238 = n21233 & n21234 ;
  assign n21242 = n21237 & n21238 ;
  assign n21243 = n21241 & n21242 ;
  assign n21244 = n16984 & ~n21243 ;
  assign n21245 = \P1_buf2_reg[4]/NET0131  & n9085 ;
  assign n21246 = \P1_buf2_reg[20]/NET0131  & n9086 ;
  assign n21247 = ~n21245 & ~n21246 ;
  assign n21248 = n9088 & ~n21247 ;
  assign n21249 = ~n21244 & ~n21248 ;
  assign n21250 = ~n21212 & n21249 ;
  assign n21251 = ~n21210 & n21250 ;
  assign n21252 = n9241 & ~n21251 ;
  assign n21253 = ~n21208 & ~n21252 ;
  assign n21254 = \P1_P3_EAX_reg[21]/NET0131  & ~n16968 ;
  assign n21256 = \P1_P3_EAX_reg[20]/NET0131  & n21162 ;
  assign n21258 = ~\P1_P3_EAX_reg[21]/NET0131  & ~n21256 ;
  assign n21257 = \P1_P3_EAX_reg[21]/NET0131  & n21256 ;
  assign n21259 = n16982 & ~n21257 ;
  assign n21260 = ~n21258 & n21259 ;
  assign n21255 = \P1_P3_EAX_reg[21]/NET0131  & ~n16988 ;
  assign n21261 = \P1_buf2_reg[5]/NET0131  & n9085 ;
  assign n21262 = \P1_buf2_reg[21]/NET0131  & n9086 ;
  assign n21263 = ~n21261 & ~n21262 ;
  assign n21264 = n9088 & ~n21263 ;
  assign n21269 = \P1_P3_InstQueue_reg[6][5]/NET0131  & n8771 ;
  assign n21270 = \P1_P3_InstQueue_reg[14][5]/NET0131  & n8765 ;
  assign n21283 = ~n21269 & ~n21270 ;
  assign n21271 = \P1_P3_InstQueue_reg[11][5]/NET0131  & n8769 ;
  assign n21272 = \P1_P3_InstQueue_reg[5][5]/NET0131  & n8752 ;
  assign n21284 = ~n21271 & ~n21272 ;
  assign n21291 = n21283 & n21284 ;
  assign n21265 = \P1_P3_InstQueue_reg[4][5]/NET0131  & n8777 ;
  assign n21266 = \P1_P3_InstQueue_reg[10][5]/NET0131  & n8748 ;
  assign n21281 = ~n21265 & ~n21266 ;
  assign n21267 = \P1_P3_InstQueue_reg[0][5]/NET0131  & n8775 ;
  assign n21268 = \P1_P3_InstQueue_reg[8][5]/NET0131  & n8779 ;
  assign n21282 = ~n21267 & ~n21268 ;
  assign n21292 = n21281 & n21282 ;
  assign n21293 = n21291 & n21292 ;
  assign n21277 = \P1_P3_InstQueue_reg[13][5]/NET0131  & n8757 ;
  assign n21278 = \P1_P3_InstQueue_reg[12][5]/NET0131  & n8763 ;
  assign n21287 = ~n21277 & ~n21278 ;
  assign n21279 = \P1_P3_InstQueue_reg[7][5]/NET0131  & n8745 ;
  assign n21280 = \P1_P3_InstQueue_reg[1][5]/NET0131  & n8781 ;
  assign n21288 = ~n21279 & ~n21280 ;
  assign n21289 = n21287 & n21288 ;
  assign n21273 = \P1_P3_InstQueue_reg[15][5]/NET0131  & n8760 ;
  assign n21274 = \P1_P3_InstQueue_reg[3][5]/NET0131  & n8767 ;
  assign n21285 = ~n21273 & ~n21274 ;
  assign n21275 = \P1_P3_InstQueue_reg[9][5]/NET0131  & n8754 ;
  assign n21276 = \P1_P3_InstQueue_reg[2][5]/NET0131  & n8773 ;
  assign n21286 = ~n21275 & ~n21276 ;
  assign n21290 = n21285 & n21286 ;
  assign n21294 = n21289 & n21290 ;
  assign n21295 = n21293 & n21294 ;
  assign n21296 = n16984 & ~n21295 ;
  assign n21297 = ~n21264 & ~n21296 ;
  assign n21298 = ~n21255 & n21297 ;
  assign n21299 = ~n21260 & n21298 ;
  assign n21300 = n9241 & ~n21299 ;
  assign n21301 = ~n21254 & ~n21300 ;
  assign n21302 = \P1_P3_EAX_reg[22]/NET0131  & ~n16968 ;
  assign n21304 = \P1_P3_EAX_reg[21]/NET0131  & \P1_P3_EAX_reg[22]/NET0131  ;
  assign n21305 = n21256 & n21304 ;
  assign n21306 = n16982 & ~n21305 ;
  assign n21307 = ~\P1_P3_EAX_reg[22]/NET0131  & ~n21257 ;
  assign n21308 = n21306 & ~n21307 ;
  assign n21303 = \P1_P3_EAX_reg[22]/NET0131  & ~n16988 ;
  assign n21309 = \P1_buf2_reg[6]/NET0131  & n9085 ;
  assign n21310 = \P1_buf2_reg[22]/NET0131  & n9086 ;
  assign n21311 = ~n21309 & ~n21310 ;
  assign n21312 = n9088 & ~n21311 ;
  assign n21317 = \P1_P3_InstQueue_reg[6][6]/NET0131  & n8771 ;
  assign n21318 = \P1_P3_InstQueue_reg[14][6]/NET0131  & n8765 ;
  assign n21331 = ~n21317 & ~n21318 ;
  assign n21319 = \P1_P3_InstQueue_reg[11][6]/NET0131  & n8769 ;
  assign n21320 = \P1_P3_InstQueue_reg[5][6]/NET0131  & n8752 ;
  assign n21332 = ~n21319 & ~n21320 ;
  assign n21339 = n21331 & n21332 ;
  assign n21313 = \P1_P3_InstQueue_reg[4][6]/NET0131  & n8777 ;
  assign n21314 = \P1_P3_InstQueue_reg[10][6]/NET0131  & n8748 ;
  assign n21329 = ~n21313 & ~n21314 ;
  assign n21315 = \P1_P3_InstQueue_reg[0][6]/NET0131  & n8775 ;
  assign n21316 = \P1_P3_InstQueue_reg[8][6]/NET0131  & n8779 ;
  assign n21330 = ~n21315 & ~n21316 ;
  assign n21340 = n21329 & n21330 ;
  assign n21341 = n21339 & n21340 ;
  assign n21325 = \P1_P3_InstQueue_reg[13][6]/NET0131  & n8757 ;
  assign n21326 = \P1_P3_InstQueue_reg[12][6]/NET0131  & n8763 ;
  assign n21335 = ~n21325 & ~n21326 ;
  assign n21327 = \P1_P3_InstQueue_reg[7][6]/NET0131  & n8745 ;
  assign n21328 = \P1_P3_InstQueue_reg[1][6]/NET0131  & n8781 ;
  assign n21336 = ~n21327 & ~n21328 ;
  assign n21337 = n21335 & n21336 ;
  assign n21321 = \P1_P3_InstQueue_reg[15][6]/NET0131  & n8760 ;
  assign n21322 = \P1_P3_InstQueue_reg[3][6]/NET0131  & n8767 ;
  assign n21333 = ~n21321 & ~n21322 ;
  assign n21323 = \P1_P3_InstQueue_reg[9][6]/NET0131  & n8754 ;
  assign n21324 = \P1_P3_InstQueue_reg[2][6]/NET0131  & n8773 ;
  assign n21334 = ~n21323 & ~n21324 ;
  assign n21338 = n21333 & n21334 ;
  assign n21342 = n21337 & n21338 ;
  assign n21343 = n21341 & n21342 ;
  assign n21344 = n16984 & ~n21343 ;
  assign n21345 = ~n21312 & ~n21344 ;
  assign n21346 = ~n21303 & n21345 ;
  assign n21347 = ~n21308 & n21346 ;
  assign n21348 = n9241 & ~n21347 ;
  assign n21349 = ~n21302 & ~n21348 ;
  assign n21350 = \P1_P3_EAX_reg[23]/NET0131  & ~n16968 ;
  assign n21417 = ~n16987 & ~n21306 ;
  assign n21418 = \P1_P3_EAX_reg[23]/NET0131  & ~n21417 ;
  assign n21425 = ~\P1_P3_EAX_reg[23]/NET0131  & n16982 ;
  assign n21426 = n21305 & n21425 ;
  assign n21419 = \P1_P3_EAX_reg[23]/NET0131  & ~n9088 ;
  assign n21423 = ~n17284 & ~n21419 ;
  assign n21424 = n9085 & ~n21423 ;
  assign n21355 = \P1_P3_InstQueue_reg[15][7]/NET0131  & n8760 ;
  assign n21356 = \P1_P3_InstQueue_reg[13][7]/NET0131  & n8757 ;
  assign n21369 = ~n21355 & ~n21356 ;
  assign n21357 = \P1_P3_InstQueue_reg[8][7]/NET0131  & n8779 ;
  assign n21358 = \P1_P3_InstQueue_reg[14][7]/NET0131  & n8765 ;
  assign n21370 = ~n21357 & ~n21358 ;
  assign n21377 = n21369 & n21370 ;
  assign n21351 = \P1_P3_InstQueue_reg[0][7]/NET0131  & n8775 ;
  assign n21352 = \P1_P3_InstQueue_reg[10][7]/NET0131  & n8748 ;
  assign n21367 = ~n21351 & ~n21352 ;
  assign n21353 = \P1_P3_InstQueue_reg[7][7]/NET0131  & n8745 ;
  assign n21354 = \P1_P3_InstQueue_reg[3][7]/NET0131  & n8767 ;
  assign n21368 = ~n21353 & ~n21354 ;
  assign n21378 = n21367 & n21368 ;
  assign n21379 = n21377 & n21378 ;
  assign n21363 = \P1_P3_InstQueue_reg[4][7]/NET0131  & n8777 ;
  assign n21364 = \P1_P3_InstQueue_reg[12][7]/NET0131  & n8763 ;
  assign n21373 = ~n21363 & ~n21364 ;
  assign n21365 = \P1_P3_InstQueue_reg[5][7]/NET0131  & n8752 ;
  assign n21366 = \P1_P3_InstQueue_reg[1][7]/NET0131  & n8781 ;
  assign n21374 = ~n21365 & ~n21366 ;
  assign n21375 = n21373 & n21374 ;
  assign n21359 = \P1_P3_InstQueue_reg[11][7]/NET0131  & n8769 ;
  assign n21360 = \P1_P3_InstQueue_reg[6][7]/NET0131  & n8771 ;
  assign n21371 = ~n21359 & ~n21360 ;
  assign n21361 = \P1_P3_InstQueue_reg[9][7]/NET0131  & n8754 ;
  assign n21362 = \P1_P3_InstQueue_reg[2][7]/NET0131  & n8773 ;
  assign n21372 = ~n21361 & ~n21362 ;
  assign n21376 = n21371 & n21372 ;
  assign n21380 = n21375 & n21376 ;
  assign n21381 = n21379 & n21380 ;
  assign n21386 = \P1_P3_InstQueue_reg[0][0]/NET0131  & n8760 ;
  assign n21387 = \P1_P3_InstQueue_reg[6][0]/NET0131  & n8752 ;
  assign n21400 = ~n21386 & ~n21387 ;
  assign n21388 = \P1_P3_InstQueue_reg[12][0]/NET0131  & n8769 ;
  assign n21389 = \P1_P3_InstQueue_reg[10][0]/NET0131  & n8754 ;
  assign n21401 = ~n21388 & ~n21389 ;
  assign n21408 = n21400 & n21401 ;
  assign n21382 = \P1_P3_InstQueue_reg[13][0]/NET0131  & n8763 ;
  assign n21383 = \P1_P3_InstQueue_reg[11][0]/NET0131  & n8748 ;
  assign n21398 = ~n21382 & ~n21383 ;
  assign n21384 = \P1_P3_InstQueue_reg[9][0]/NET0131  & n8779 ;
  assign n21385 = \P1_P3_InstQueue_reg[14][0]/NET0131  & n8757 ;
  assign n21399 = ~n21384 & ~n21385 ;
  assign n21409 = n21398 & n21399 ;
  assign n21410 = n21408 & n21409 ;
  assign n21394 = \P1_P3_InstQueue_reg[4][0]/NET0131  & n8767 ;
  assign n21395 = \P1_P3_InstQueue_reg[5][0]/NET0131  & n8777 ;
  assign n21404 = ~n21394 & ~n21395 ;
  assign n21396 = \P1_P3_InstQueue_reg[1][0]/NET0131  & n8775 ;
  assign n21397 = \P1_P3_InstQueue_reg[2][0]/NET0131  & n8781 ;
  assign n21405 = ~n21396 & ~n21397 ;
  assign n21406 = n21404 & n21405 ;
  assign n21390 = \P1_P3_InstQueue_reg[7][0]/NET0131  & n8771 ;
  assign n21391 = \P1_P3_InstQueue_reg[15][0]/NET0131  & n8765 ;
  assign n21402 = ~n21390 & ~n21391 ;
  assign n21392 = \P1_P3_InstQueue_reg[8][0]/NET0131  & n8745 ;
  assign n21393 = \P1_P3_InstQueue_reg[3][0]/NET0131  & n8773 ;
  assign n21403 = ~n21392 & ~n21393 ;
  assign n21407 = n21402 & n21403 ;
  assign n21411 = n21406 & n21407 ;
  assign n21412 = n21410 & n21411 ;
  assign n21413 = n21381 & n21412 ;
  assign n21414 = ~n21381 & ~n21412 ;
  assign n21415 = ~n21413 & ~n21414 ;
  assign n21416 = n16984 & n21415 ;
  assign n21420 = \P1_buf2_reg[23]/NET0131  & n9088 ;
  assign n21421 = ~n21419 & ~n21420 ;
  assign n21422 = n9086 & ~n21421 ;
  assign n21427 = ~n21416 & ~n21422 ;
  assign n21428 = ~n21424 & n21427 ;
  assign n21429 = ~n21426 & n21428 ;
  assign n21430 = ~n21418 & n21429 ;
  assign n21431 = n9241 & ~n21430 ;
  assign n21432 = ~n21350 & ~n21431 ;
  assign n21433 = \P1_P3_EAX_reg[24]/NET0131  & ~n17077 ;
  assign n21470 = \P1_P3_EAX_reg[18]/NET0131  & \P1_P3_EAX_reg[19]/NET0131  ;
  assign n21471 = \P1_P3_EAX_reg[20]/NET0131  & \P1_P3_EAX_reg[23]/NET0131  ;
  assign n21472 = n21470 & n21471 ;
  assign n21469 = \P1_P3_EAX_reg[16]/NET0131  & \P1_P3_EAX_reg[17]/NET0131  ;
  assign n21473 = n21304 & n21469 ;
  assign n21474 = n21472 & n21473 ;
  assign n21475 = n18753 & n21474 ;
  assign n21477 = ~\P1_P3_EAX_reg[24]/NET0131  & ~n21475 ;
  assign n21476 = \P1_P3_EAX_reg[24]/NET0131  & n21475 ;
  assign n21478 = n16982 & ~n21476 ;
  assign n21479 = ~n21477 & n21478 ;
  assign n21480 = \P1_P3_EAX_reg[24]/NET0131  & ~n9088 ;
  assign n21484 = ~n17294 & ~n21480 ;
  assign n21485 = n9085 & ~n21484 ;
  assign n21438 = \P1_P3_InstQueue_reg[9][1]/NET0131  & n8779 ;
  assign n21439 = \P1_P3_InstQueue_reg[14][1]/NET0131  & n8757 ;
  assign n21452 = ~n21438 & ~n21439 ;
  assign n21440 = \P1_P3_InstQueue_reg[1][1]/NET0131  & n8775 ;
  assign n21441 = \P1_P3_InstQueue_reg[10][1]/NET0131  & n8754 ;
  assign n21453 = ~n21440 & ~n21441 ;
  assign n21460 = n21452 & n21453 ;
  assign n21434 = \P1_P3_InstQueue_reg[6][1]/NET0131  & n8752 ;
  assign n21435 = \P1_P3_InstQueue_reg[11][1]/NET0131  & n8748 ;
  assign n21450 = ~n21434 & ~n21435 ;
  assign n21436 = \P1_P3_InstQueue_reg[12][1]/NET0131  & n8769 ;
  assign n21437 = \P1_P3_InstQueue_reg[13][1]/NET0131  & n8763 ;
  assign n21451 = ~n21436 & ~n21437 ;
  assign n21461 = n21450 & n21451 ;
  assign n21462 = n21460 & n21461 ;
  assign n21446 = \P1_P3_InstQueue_reg[8][1]/NET0131  & n8745 ;
  assign n21447 = \P1_P3_InstQueue_reg[7][1]/NET0131  & n8771 ;
  assign n21456 = ~n21446 & ~n21447 ;
  assign n21448 = \P1_P3_InstQueue_reg[0][1]/NET0131  & n8760 ;
  assign n21449 = \P1_P3_InstQueue_reg[2][1]/NET0131  & n8781 ;
  assign n21457 = ~n21448 & ~n21449 ;
  assign n21458 = n21456 & n21457 ;
  assign n21442 = \P1_P3_InstQueue_reg[5][1]/NET0131  & n8777 ;
  assign n21443 = \P1_P3_InstQueue_reg[4][1]/NET0131  & n8767 ;
  assign n21454 = ~n21442 & ~n21443 ;
  assign n21444 = \P1_P3_InstQueue_reg[15][1]/NET0131  & n8765 ;
  assign n21445 = \P1_P3_InstQueue_reg[3][1]/NET0131  & n8773 ;
  assign n21455 = ~n21444 & ~n21445 ;
  assign n21459 = n21454 & n21455 ;
  assign n21463 = n21458 & n21459 ;
  assign n21464 = n21462 & n21463 ;
  assign n21465 = ~n21414 & n21464 ;
  assign n21466 = n21414 & ~n21464 ;
  assign n21467 = ~n21465 & ~n21466 ;
  assign n21468 = n16984 & n21467 ;
  assign n21481 = \P1_buf2_reg[24]/NET0131  & n9088 ;
  assign n21482 = ~n21480 & ~n21481 ;
  assign n21483 = n9086 & ~n21482 ;
  assign n21486 = ~n21468 & ~n21483 ;
  assign n21487 = ~n21485 & n21486 ;
  assign n21488 = ~n21479 & n21487 ;
  assign n21489 = n9241 & ~n21488 ;
  assign n21490 = ~n21433 & ~n21489 ;
  assign n21491 = \P1_P3_EAX_reg[29]/NET0131  & ~n16968 ;
  assign n21492 = \P1_P3_EAX_reg[24]/NET0131  & \P1_P3_EAX_reg[25]/NET0131  ;
  assign n21493 = \P1_P3_EAX_reg[26]/NET0131  & \P1_P3_EAX_reg[27]/NET0131  ;
  assign n21494 = n21492 & n21493 ;
  assign n21495 = n21474 & n21494 ;
  assign n21496 = n18753 & n21495 ;
  assign n21497 = \P1_P3_EAX_reg[28]/NET0131  & n21496 ;
  assign n21498 = n16982 & ~n21497 ;
  assign n21499 = ~n16987 & ~n21498 ;
  assign n21500 = \P1_P3_EAX_reg[29]/NET0131  & ~n21499 ;
  assign n21501 = n16982 & n21496 ;
  assign n21502 = \P1_P3_EAX_reg[28]/NET0131  & ~\P1_P3_EAX_reg[29]/NET0131  ;
  assign n21503 = n21501 & n21502 ;
  assign n21508 = \P1_P3_InstQueue_reg[0][2]/NET0131  & n8760 ;
  assign n21509 = \P1_P3_InstQueue_reg[6][2]/NET0131  & n8752 ;
  assign n21522 = ~n21508 & ~n21509 ;
  assign n21510 = \P1_P3_InstQueue_reg[12][2]/NET0131  & n8769 ;
  assign n21511 = \P1_P3_InstQueue_reg[10][2]/NET0131  & n8754 ;
  assign n21523 = ~n21510 & ~n21511 ;
  assign n21530 = n21522 & n21523 ;
  assign n21504 = \P1_P3_InstQueue_reg[13][2]/NET0131  & n8763 ;
  assign n21505 = \P1_P3_InstQueue_reg[11][2]/NET0131  & n8748 ;
  assign n21520 = ~n21504 & ~n21505 ;
  assign n21506 = \P1_P3_InstQueue_reg[9][2]/NET0131  & n8779 ;
  assign n21507 = \P1_P3_InstQueue_reg[14][2]/NET0131  & n8757 ;
  assign n21521 = ~n21506 & ~n21507 ;
  assign n21531 = n21520 & n21521 ;
  assign n21532 = n21530 & n21531 ;
  assign n21516 = \P1_P3_InstQueue_reg[4][2]/NET0131  & n8767 ;
  assign n21517 = \P1_P3_InstQueue_reg[5][2]/NET0131  & n8777 ;
  assign n21526 = ~n21516 & ~n21517 ;
  assign n21518 = \P1_P3_InstQueue_reg[1][2]/NET0131  & n8775 ;
  assign n21519 = \P1_P3_InstQueue_reg[2][2]/NET0131  & n8781 ;
  assign n21527 = ~n21518 & ~n21519 ;
  assign n21528 = n21526 & n21527 ;
  assign n21512 = \P1_P3_InstQueue_reg[7][2]/NET0131  & n8771 ;
  assign n21513 = \P1_P3_InstQueue_reg[15][2]/NET0131  & n8765 ;
  assign n21524 = ~n21512 & ~n21513 ;
  assign n21514 = \P1_P3_InstQueue_reg[8][2]/NET0131  & n8745 ;
  assign n21515 = \P1_P3_InstQueue_reg[3][2]/NET0131  & n8773 ;
  assign n21525 = ~n21514 & ~n21515 ;
  assign n21529 = n21524 & n21525 ;
  assign n21533 = n21528 & n21529 ;
  assign n21534 = n21532 & n21533 ;
  assign n21535 = n21466 & ~n21534 ;
  assign n21540 = \P1_P3_InstQueue_reg[0][3]/NET0131  & n8760 ;
  assign n21541 = \P1_P3_InstQueue_reg[6][3]/NET0131  & n8752 ;
  assign n21554 = ~n21540 & ~n21541 ;
  assign n21542 = \P1_P3_InstQueue_reg[12][3]/NET0131  & n8769 ;
  assign n21543 = \P1_P3_InstQueue_reg[10][3]/NET0131  & n8754 ;
  assign n21555 = ~n21542 & ~n21543 ;
  assign n21562 = n21554 & n21555 ;
  assign n21536 = \P1_P3_InstQueue_reg[13][3]/NET0131  & n8763 ;
  assign n21537 = \P1_P3_InstQueue_reg[11][3]/NET0131  & n8748 ;
  assign n21552 = ~n21536 & ~n21537 ;
  assign n21538 = \P1_P3_InstQueue_reg[9][3]/NET0131  & n8779 ;
  assign n21539 = \P1_P3_InstQueue_reg[14][3]/NET0131  & n8757 ;
  assign n21553 = ~n21538 & ~n21539 ;
  assign n21563 = n21552 & n21553 ;
  assign n21564 = n21562 & n21563 ;
  assign n21548 = \P1_P3_InstQueue_reg[4][3]/NET0131  & n8767 ;
  assign n21549 = \P1_P3_InstQueue_reg[5][3]/NET0131  & n8777 ;
  assign n21558 = ~n21548 & ~n21549 ;
  assign n21550 = \P1_P3_InstQueue_reg[1][3]/NET0131  & n8775 ;
  assign n21551 = \P1_P3_InstQueue_reg[2][3]/NET0131  & n8781 ;
  assign n21559 = ~n21550 & ~n21551 ;
  assign n21560 = n21558 & n21559 ;
  assign n21544 = \P1_P3_InstQueue_reg[7][3]/NET0131  & n8771 ;
  assign n21545 = \P1_P3_InstQueue_reg[15][3]/NET0131  & n8765 ;
  assign n21556 = ~n21544 & ~n21545 ;
  assign n21546 = \P1_P3_InstQueue_reg[8][3]/NET0131  & n8745 ;
  assign n21547 = \P1_P3_InstQueue_reg[3][3]/NET0131  & n8773 ;
  assign n21557 = ~n21546 & ~n21547 ;
  assign n21561 = n21556 & n21557 ;
  assign n21565 = n21560 & n21561 ;
  assign n21566 = n21564 & n21565 ;
  assign n21567 = n21535 & ~n21566 ;
  assign n21572 = \P1_P3_InstQueue_reg[0][4]/NET0131  & n8760 ;
  assign n21573 = \P1_P3_InstQueue_reg[6][4]/NET0131  & n8752 ;
  assign n21586 = ~n21572 & ~n21573 ;
  assign n21574 = \P1_P3_InstQueue_reg[12][4]/NET0131  & n8769 ;
  assign n21575 = \P1_P3_InstQueue_reg[10][4]/NET0131  & n8754 ;
  assign n21587 = ~n21574 & ~n21575 ;
  assign n21594 = n21586 & n21587 ;
  assign n21568 = \P1_P3_InstQueue_reg[13][4]/NET0131  & n8763 ;
  assign n21569 = \P1_P3_InstQueue_reg[11][4]/NET0131  & n8748 ;
  assign n21584 = ~n21568 & ~n21569 ;
  assign n21570 = \P1_P3_InstQueue_reg[9][4]/NET0131  & n8779 ;
  assign n21571 = \P1_P3_InstQueue_reg[14][4]/NET0131  & n8757 ;
  assign n21585 = ~n21570 & ~n21571 ;
  assign n21595 = n21584 & n21585 ;
  assign n21596 = n21594 & n21595 ;
  assign n21580 = \P1_P3_InstQueue_reg[4][4]/NET0131  & n8767 ;
  assign n21581 = \P1_P3_InstQueue_reg[5][4]/NET0131  & n8777 ;
  assign n21590 = ~n21580 & ~n21581 ;
  assign n21582 = \P1_P3_InstQueue_reg[1][4]/NET0131  & n8775 ;
  assign n21583 = \P1_P3_InstQueue_reg[2][4]/NET0131  & n8781 ;
  assign n21591 = ~n21582 & ~n21583 ;
  assign n21592 = n21590 & n21591 ;
  assign n21576 = \P1_P3_InstQueue_reg[7][4]/NET0131  & n8771 ;
  assign n21577 = \P1_P3_InstQueue_reg[15][4]/NET0131  & n8765 ;
  assign n21588 = ~n21576 & ~n21577 ;
  assign n21578 = \P1_P3_InstQueue_reg[8][4]/NET0131  & n8745 ;
  assign n21579 = \P1_P3_InstQueue_reg[3][4]/NET0131  & n8773 ;
  assign n21589 = ~n21578 & ~n21579 ;
  assign n21593 = n21588 & n21589 ;
  assign n21597 = n21592 & n21593 ;
  assign n21598 = n21596 & n21597 ;
  assign n21599 = n21567 & ~n21598 ;
  assign n21604 = \P1_P3_InstQueue_reg[4][5]/NET0131  & n8767 ;
  assign n21605 = \P1_P3_InstQueue_reg[14][5]/NET0131  & n8757 ;
  assign n21618 = ~n21604 & ~n21605 ;
  assign n21606 = \P1_P3_InstQueue_reg[5][5]/NET0131  & n8777 ;
  assign n21607 = \P1_P3_InstQueue_reg[10][5]/NET0131  & n8754 ;
  assign n21619 = ~n21606 & ~n21607 ;
  assign n21626 = n21618 & n21619 ;
  assign n21600 = \P1_P3_InstQueue_reg[1][5]/NET0131  & n8775 ;
  assign n21601 = \P1_P3_InstQueue_reg[11][5]/NET0131  & n8748 ;
  assign n21616 = ~n21600 & ~n21601 ;
  assign n21602 = \P1_P3_InstQueue_reg[8][5]/NET0131  & n8745 ;
  assign n21603 = \P1_P3_InstQueue_reg[15][5]/NET0131  & n8765 ;
  assign n21617 = ~n21602 & ~n21603 ;
  assign n21627 = n21616 & n21617 ;
  assign n21628 = n21626 & n21627 ;
  assign n21612 = \P1_P3_InstQueue_reg[0][5]/NET0131  & n8760 ;
  assign n21613 = \P1_P3_InstQueue_reg[6][5]/NET0131  & n8752 ;
  assign n21622 = ~n21612 & ~n21613 ;
  assign n21614 = \P1_P3_InstQueue_reg[12][5]/NET0131  & n8769 ;
  assign n21615 = \P1_P3_InstQueue_reg[2][5]/NET0131  & n8781 ;
  assign n21623 = ~n21614 & ~n21615 ;
  assign n21624 = n21622 & n21623 ;
  assign n21608 = \P1_P3_InstQueue_reg[13][5]/NET0131  & n8763 ;
  assign n21609 = \P1_P3_InstQueue_reg[7][5]/NET0131  & n8771 ;
  assign n21620 = ~n21608 & ~n21609 ;
  assign n21610 = \P1_P3_InstQueue_reg[9][5]/NET0131  & n8779 ;
  assign n21611 = \P1_P3_InstQueue_reg[3][5]/NET0131  & n8773 ;
  assign n21621 = ~n21610 & ~n21611 ;
  assign n21625 = n21620 & n21621 ;
  assign n21629 = n21624 & n21625 ;
  assign n21630 = n21628 & n21629 ;
  assign n21631 = n21599 & ~n21630 ;
  assign n21636 = \P1_P3_InstQueue_reg[4][6]/NET0131  & n8767 ;
  assign n21637 = \P1_P3_InstQueue_reg[14][6]/NET0131  & n8757 ;
  assign n21650 = ~n21636 & ~n21637 ;
  assign n21638 = \P1_P3_InstQueue_reg[5][6]/NET0131  & n8777 ;
  assign n21639 = \P1_P3_InstQueue_reg[10][6]/NET0131  & n8754 ;
  assign n21651 = ~n21638 & ~n21639 ;
  assign n21658 = n21650 & n21651 ;
  assign n21632 = \P1_P3_InstQueue_reg[1][6]/NET0131  & n8775 ;
  assign n21633 = \P1_P3_InstQueue_reg[11][6]/NET0131  & n8748 ;
  assign n21648 = ~n21632 & ~n21633 ;
  assign n21634 = \P1_P3_InstQueue_reg[8][6]/NET0131  & n8745 ;
  assign n21635 = \P1_P3_InstQueue_reg[15][6]/NET0131  & n8765 ;
  assign n21649 = ~n21634 & ~n21635 ;
  assign n21659 = n21648 & n21649 ;
  assign n21660 = n21658 & n21659 ;
  assign n21644 = \P1_P3_InstQueue_reg[0][6]/NET0131  & n8760 ;
  assign n21645 = \P1_P3_InstQueue_reg[6][6]/NET0131  & n8752 ;
  assign n21654 = ~n21644 & ~n21645 ;
  assign n21646 = \P1_P3_InstQueue_reg[12][6]/NET0131  & n8769 ;
  assign n21647 = \P1_P3_InstQueue_reg[2][6]/NET0131  & n8781 ;
  assign n21655 = ~n21646 & ~n21647 ;
  assign n21656 = n21654 & n21655 ;
  assign n21640 = \P1_P3_InstQueue_reg[13][6]/NET0131  & n8763 ;
  assign n21641 = \P1_P3_InstQueue_reg[7][6]/NET0131  & n8771 ;
  assign n21652 = ~n21640 & ~n21641 ;
  assign n21642 = \P1_P3_InstQueue_reg[9][6]/NET0131  & n8779 ;
  assign n21643 = \P1_P3_InstQueue_reg[3][6]/NET0131  & n8773 ;
  assign n21653 = ~n21642 & ~n21643 ;
  assign n21657 = n21652 & n21653 ;
  assign n21661 = n21656 & n21657 ;
  assign n21662 = n21660 & n21661 ;
  assign n21663 = ~n21631 & n21662 ;
  assign n21664 = n21631 & ~n21662 ;
  assign n21665 = ~n21663 & ~n21664 ;
  assign n21666 = n16984 & n21665 ;
  assign n21667 = \P1_P3_EAX_reg[29]/NET0131  & ~n9088 ;
  assign n21668 = ~n17079 & ~n21667 ;
  assign n21669 = n9085 & ~n21668 ;
  assign n21670 = \P1_buf2_reg[29]/NET0131  & n9088 ;
  assign n21671 = ~n21667 & ~n21670 ;
  assign n21672 = n9086 & ~n21671 ;
  assign n21673 = ~n21669 & ~n21672 ;
  assign n21674 = ~n21666 & n21673 ;
  assign n21675 = ~n21503 & n21674 ;
  assign n21676 = ~n21500 & n21675 ;
  assign n21677 = n9241 & ~n21676 ;
  assign n21678 = ~n21491 & ~n21677 ;
  assign n21680 = \P1_P3_EAX_reg[28]/NET0131  & \P1_P3_EAX_reg[29]/NET0131  ;
  assign n21681 = n21496 & n21680 ;
  assign n21682 = ~\P1_P3_EAX_reg[30]/NET0131  & ~n21681 ;
  assign n21683 = \P1_P3_EAX_reg[30]/NET0131  & n21681 ;
  assign n21684 = n16982 & ~n21683 ;
  assign n21685 = ~n21682 & n21684 ;
  assign n21690 = \P1_P3_InstQueue_reg[0][7]/NET0131  & n8760 ;
  assign n21691 = \P1_P3_InstQueue_reg[6][7]/NET0131  & n8752 ;
  assign n21704 = ~n21690 & ~n21691 ;
  assign n21692 = \P1_P3_InstQueue_reg[12][7]/NET0131  & n8769 ;
  assign n21693 = \P1_P3_InstQueue_reg[10][7]/NET0131  & n8754 ;
  assign n21705 = ~n21692 & ~n21693 ;
  assign n21712 = n21704 & n21705 ;
  assign n21686 = \P1_P3_InstQueue_reg[13][7]/NET0131  & n8763 ;
  assign n21687 = \P1_P3_InstQueue_reg[11][7]/NET0131  & n8748 ;
  assign n21702 = ~n21686 & ~n21687 ;
  assign n21688 = \P1_P3_InstQueue_reg[9][7]/NET0131  & n8779 ;
  assign n21689 = \P1_P3_InstQueue_reg[14][7]/NET0131  & n8757 ;
  assign n21703 = ~n21688 & ~n21689 ;
  assign n21713 = n21702 & n21703 ;
  assign n21714 = n21712 & n21713 ;
  assign n21698 = \P1_P3_InstQueue_reg[4][7]/NET0131  & n8767 ;
  assign n21699 = \P1_P3_InstQueue_reg[5][7]/NET0131  & n8777 ;
  assign n21708 = ~n21698 & ~n21699 ;
  assign n21700 = \P1_P3_InstQueue_reg[1][7]/NET0131  & n8775 ;
  assign n21701 = \P1_P3_InstQueue_reg[2][7]/NET0131  & n8781 ;
  assign n21709 = ~n21700 & ~n21701 ;
  assign n21710 = n21708 & n21709 ;
  assign n21694 = \P1_P3_InstQueue_reg[7][7]/NET0131  & n8771 ;
  assign n21695 = \P1_P3_InstQueue_reg[15][7]/NET0131  & n8765 ;
  assign n21706 = ~n21694 & ~n21695 ;
  assign n21696 = \P1_P3_InstQueue_reg[8][7]/NET0131  & n8745 ;
  assign n21697 = \P1_P3_InstQueue_reg[3][7]/NET0131  & n8773 ;
  assign n21707 = ~n21696 & ~n21697 ;
  assign n21711 = n21706 & n21707 ;
  assign n21715 = n21710 & n21711 ;
  assign n21716 = n21714 & n21715 ;
  assign n21717 = n21664 & ~n21716 ;
  assign n21718 = ~n21664 & n21716 ;
  assign n21719 = ~n21717 & ~n21718 ;
  assign n21720 = n16984 & n21719 ;
  assign n21679 = \P1_P3_EAX_reg[30]/NET0131  & ~n16988 ;
  assign n21721 = \P1_buf2_reg[14]/NET0131  & n9085 ;
  assign n21722 = \P1_buf2_reg[30]/NET0131  & n9086 ;
  assign n21723 = ~n21721 & ~n21722 ;
  assign n21724 = n9088 & ~n21723 ;
  assign n21725 = ~n21679 & ~n21724 ;
  assign n21726 = ~n21720 & n21725 ;
  assign n21727 = ~n21685 & n21726 ;
  assign n21728 = n9241 & ~n21727 ;
  assign n21729 = \P1_P3_EAX_reg[30]/NET0131  & ~n16968 ;
  assign n21730 = ~n21728 & ~n21729 ;
  assign n21733 = ~\P1_P3_PhyAddrPointer_reg[5]/NET0131  & ~n17533 ;
  assign n21734 = ~n17568 & ~n21733 ;
  assign n21735 = \P1_P3_PhyAddrPointer_reg[4]/NET0131  & n17535 ;
  assign n21736 = n16484 & ~n21735 ;
  assign n21738 = ~n21734 & n21736 ;
  assign n21737 = n21734 & ~n21736 ;
  assign n21739 = ~\P1_P3_DataWidth_reg[1]/NET0131  & ~n21737 ;
  assign n21740 = ~n21738 & n21739 ;
  assign n21732 = \P1_P3_DataWidth_reg[1]/NET0131  & ~\P1_P3_rEIP_reg[5]/NET0131  ;
  assign n21741 = n9245 & ~n21732 ;
  assign n21742 = ~n21740 & n21741 ;
  assign n21743 = \P1_P3_rEIP_reg[5]/NET0131  & ~n9195 ;
  assign n21744 = ~\P1_P3_rEIP_reg[5]/NET0131  & ~n16570 ;
  assign n21745 = ~n16571 & ~n21744 ;
  assign n21746 = n16505 & ~n21745 ;
  assign n21747 = ~n9095 & n21746 ;
  assign n21748 = ~\P1_P3_EBX_reg[5]/NET0131  & ~n16517 ;
  assign n21749 = ~n21747 & ~n21748 ;
  assign n21750 = n9236 & n21749 ;
  assign n21751 = \P1_P3_EBX_reg[31]/NET0131  & ~n16597 ;
  assign n21753 = ~\P1_P3_EBX_reg[5]/NET0131  & n21751 ;
  assign n21752 = \P1_P3_EBX_reg[5]/NET0131  & ~n21751 ;
  assign n21754 = ~n16505 & ~n21752 ;
  assign n21755 = ~n21753 & n21754 ;
  assign n21756 = ~n21746 & ~n21755 ;
  assign n21757 = n16500 & n21756 ;
  assign n21758 = ~n21750 & ~n21757 ;
  assign n21759 = ~n21743 & n21758 ;
  assign n21760 = n9241 & ~n21759 ;
  assign n21731 = \P1_P3_rEIP_reg[5]/NET0131  & ~n17458 ;
  assign n21761 = \P1_P3_PhyAddrPointer_reg[5]/NET0131  & n10031 ;
  assign n21762 = ~n17426 & ~n21761 ;
  assign n21763 = ~n21731 & n21762 ;
  assign n21764 = ~n21760 & n21763 ;
  assign n21765 = ~n21742 & n21764 ;
  assign n21772 = ~\P1_P3_RequestPending_reg/NET0131  & ~n9195 ;
  assign n21773 = n9088 & ~n9116 ;
  assign n21774 = ~n21772 & ~n21773 ;
  assign n21775 = ~n9075 & ~n9084 ;
  assign n21776 = n9095 & n21775 ;
  assign n21777 = ~n9237 & ~n21776 ;
  assign n21778 = ~n21774 & n21777 ;
  assign n21779 = n9241 & ~n21778 ;
  assign n21766 = ~\P1_P3_State2_reg[0]/NET0131  & ~n8741 ;
  assign n21767 = n10036 & ~n21766 ;
  assign n21768 = ~n10030 & ~n21767 ;
  assign n21769 = \P1_P3_RequestPending_reg/NET0131  & ~n21768 ;
  assign n21770 = ~\P1_P3_State2_reg[0]/NET0131  & \P1_P3_State2_reg[1]/NET0131  ;
  assign n21771 = n9243 & ~n21770 ;
  assign n21780 = ~n21769 & ~n21771 ;
  assign n21781 = ~n21779 & n21780 ;
  assign n21782 = \P4_reg2_reg[29]/NET0131  & ~n18665 ;
  assign n21783 = \P4_reg2_reg[29]/NET0131  & n19073 ;
  assign n21784 = \P4_IR_reg[28]/NET0131  & ~n15794 ;
  assign n21789 = ~n16302 & n18743 ;
  assign n21785 = n16302 & ~n18743 ;
  assign n21786 = \P4_IR_reg[27]/NET0131  & ~\P4_IR_reg[28]/NET0131  ;
  assign n21787 = ~\P4_B_reg/NET0131  & n21786 ;
  assign n21788 = ~n15745 & ~n21787 ;
  assign n21790 = ~n21785 & ~n21788 ;
  assign n21791 = ~n21789 & n21790 ;
  assign n21792 = ~n21784 & ~n21791 ;
  assign n21793 = n20673 & n21792 ;
  assign n21794 = ~\P4_reg2_reg[29]/NET0131  & ~n20673 ;
  assign n21795 = n18483 & ~n21794 ;
  assign n21796 = ~n21793 & n21795 ;
  assign n21830 = ~n15810 & n18640 ;
  assign n21831 = n16375 & ~n21830 ;
  assign n21832 = ~n15795 & ~n21831 ;
  assign n21834 = ~n16328 & ~n21832 ;
  assign n21833 = n16328 & n21832 ;
  assign n21835 = n18607 & ~n21833 ;
  assign n21836 = ~n21834 & n21835 ;
  assign n21798 = n18516 & n18521 ;
  assign n21799 = ~n18684 & n21798 ;
  assign n21797 = n18516 & ~n18524 ;
  assign n21800 = n18510 & ~n21797 ;
  assign n21801 = ~n21799 & n21800 ;
  assign n21802 = n18505 & n18508 ;
  assign n21803 = ~n21801 & n21802 ;
  assign n21804 = n18505 & ~n18514 ;
  assign n21805 = n18500 & ~n21804 ;
  assign n21806 = ~n21803 & n21805 ;
  assign n21807 = n18498 & ~n21806 ;
  assign n21808 = n18503 & ~n21807 ;
  assign n21809 = n18496 & ~n21808 ;
  assign n21810 = n18560 & ~n21809 ;
  assign n21811 = n18494 & ~n21810 ;
  assign n21812 = n18563 & ~n21811 ;
  assign n21813 = ~n16308 & ~n21812 ;
  assign n21814 = n18493 & ~n21813 ;
  assign n21815 = n18492 & ~n21814 ;
  assign n21816 = n18570 & ~n21815 ;
  assign n21817 = ~n16318 & ~n21816 ;
  assign n21818 = ~n16311 & ~n16317 ;
  assign n21819 = ~n21817 & n21818 ;
  assign n21820 = ~n16310 & ~n21819 ;
  assign n21822 = ~n16328 & n21820 ;
  assign n21821 = n16328 & ~n21820 ;
  assign n21823 = n18490 & ~n21821 ;
  assign n21824 = ~n21822 & n21823 ;
  assign n21825 = n15746 & n18486 ;
  assign n21827 = n15746 & ~n18730 ;
  assign n21826 = ~n15746 & n18730 ;
  assign n21828 = n18604 & ~n21826 ;
  assign n21829 = ~n21827 & n21828 ;
  assign n21837 = ~n21825 & ~n21829 ;
  assign n21838 = ~n21824 & n21837 ;
  assign n21839 = ~n21836 & n21838 ;
  assign n21840 = n20673 & ~n21839 ;
  assign n21841 = n15778 & n16426 ;
  assign n21842 = \P4_reg2_reg[29]/NET0131  & ~n20682 ;
  assign n21843 = ~n21841 & ~n21842 ;
  assign n21844 = ~n21840 & n21843 ;
  assign n21845 = ~n21796 & n21844 ;
  assign n21846 = n19075 & ~n21845 ;
  assign n21847 = ~n21783 & ~n21846 ;
  assign n21848 = \P3_rd_reg/NET0131  & ~n21847 ;
  assign n21849 = ~n21782 & ~n21848 ;
  assign n21850 = n18483 & ~n20661 ;
  assign n21851 = ~n19108 & ~n20662 ;
  assign n21852 = ~n18672 & ~n20661 ;
  assign n21853 = n18666 & ~n21852 ;
  assign n21854 = ~n21851 & n21853 ;
  assign n21855 = ~n21850 & n21854 ;
  assign n21856 = \P4_reg0_reg[15]/NET0131  & ~n21855 ;
  assign n21857 = ~n19101 & n20665 ;
  assign n21858 = ~n21856 & ~n21857 ;
  assign n21859 = \P4_reg1_reg[15]/NET0131  & ~n18679 ;
  assign n21860 = n18667 & ~n19101 ;
  assign n21861 = ~n21859 & ~n21860 ;
  assign n21865 = \P4_reg1_reg[23]/NET0131  & ~n18664 ;
  assign n21866 = ~n15844 & n18472 ;
  assign n21867 = n15844 & ~n18472 ;
  assign n21868 = ~n21866 & ~n21867 ;
  assign n21869 = ~\P4_IR_reg[28]/NET0131  & ~n21868 ;
  assign n21870 = \P4_IR_reg[28]/NET0131  & n15872 ;
  assign n21871 = ~n21869 & ~n21870 ;
  assign n21872 = n18667 & n21871 ;
  assign n21873 = ~n21865 & ~n21872 ;
  assign n21874 = n18483 & ~n21873 ;
  assign n21862 = ~n18664 & n18669 ;
  assign n21863 = n18678 & ~n21862 ;
  assign n21864 = \P4_reg1_reg[23]/NET0131  & ~n21863 ;
  assign n21879 = ~n16190 & ~n18618 ;
  assign n21880 = n18620 & ~n21879 ;
  assign n21881 = ~n16176 & ~n16189 ;
  assign n21882 = ~n21880 & n21881 ;
  assign n21883 = n18625 & ~n21882 ;
  assign n21884 = n15951 & ~n21883 ;
  assign n21885 = n16380 & ~n21884 ;
  assign n21886 = n15924 & ~n21885 ;
  assign n21887 = n16379 & ~n21886 ;
  assign n21888 = n15897 & ~n21887 ;
  assign n21889 = n16378 & ~n21888 ;
  assign n21890 = ~n15873 & ~n21889 ;
  assign n21891 = n16309 & n21890 ;
  assign n21892 = ~n16309 & ~n21890 ;
  assign n21893 = ~n21891 & ~n21892 ;
  assign n21894 = n18607 & ~n21893 ;
  assign n21895 = n18497 & n18506 ;
  assign n21900 = n18517 & n18551 ;
  assign n21901 = n21895 & n21900 ;
  assign n21896 = n18517 & ~n18525 ;
  assign n21897 = n18515 & ~n21896 ;
  assign n21898 = n21895 & ~n21897 ;
  assign n21899 = n18497 & ~n18504 ;
  assign n21902 = n18564 & ~n21899 ;
  assign n21903 = ~n21898 & n21902 ;
  assign n21904 = ~n21901 & n21903 ;
  assign n21906 = n16309 & ~n21904 ;
  assign n21905 = ~n16309 & n21904 ;
  assign n21907 = n18490 & ~n21905 ;
  assign n21908 = ~n21906 & n21907 ;
  assign n21875 = n15847 & n18486 ;
  assign n21876 = n15847 & ~n18597 ;
  assign n21877 = ~n18598 & ~n21876 ;
  assign n21878 = n18604 & n21877 ;
  assign n21909 = ~n21875 & ~n21878 ;
  assign n21910 = ~n21908 & n21909 ;
  assign n21911 = ~n21894 & n21910 ;
  assign n21912 = n18667 & ~n21911 ;
  assign n21913 = ~n21864 & ~n21912 ;
  assign n21914 = ~n21874 & n21913 ;
  assign n21915 = \P4_reg2_reg[15]/NET0131  & ~n18665 ;
  assign n21916 = \P4_reg2_reg[15]/NET0131  & n19073 ;
  assign n21918 = ~n19084 & n20673 ;
  assign n21919 = ~\P4_reg2_reg[15]/NET0131  & ~n20673 ;
  assign n21920 = n18483 & ~n21919 ;
  assign n21921 = ~n21918 & n21920 ;
  assign n21922 = ~n19100 & n20673 ;
  assign n21917 = \P4_reg2_reg[15]/NET0131  & ~n20682 ;
  assign n21923 = n16171 & n16426 ;
  assign n21924 = ~n21917 & ~n21923 ;
  assign n21925 = ~n21922 & n21924 ;
  assign n21926 = ~n21921 & n21925 ;
  assign n21927 = n19075 & ~n21926 ;
  assign n21928 = ~n21916 & ~n21927 ;
  assign n21929 = \P3_rd_reg/NET0131  & ~n21928 ;
  assign n21930 = ~n21915 & ~n21929 ;
  assign n21931 = \P1_P3_EAX_reg[28]/NET0131  & ~n16968 ;
  assign n21936 = n16982 & ~n21496 ;
  assign n21937 = ~n16987 & ~n21936 ;
  assign n21938 = \P1_P3_EAX_reg[28]/NET0131  & ~n21937 ;
  assign n21944 = ~\P1_P3_EAX_reg[28]/NET0131  & n21501 ;
  assign n21939 = ~n21599 & n21630 ;
  assign n21940 = ~n21631 & ~n21939 ;
  assign n21941 = n16984 & n21940 ;
  assign n21932 = \P1_P3_EAX_reg[28]/NET0131  & ~n9088 ;
  assign n21933 = \P1_buf2_reg[28]/NET0131  & n9088 ;
  assign n21934 = ~n21932 & ~n21933 ;
  assign n21935 = n9086 & ~n21934 ;
  assign n21942 = ~n17033 & ~n21932 ;
  assign n21943 = n9085 & ~n21942 ;
  assign n21945 = ~n21935 & ~n21943 ;
  assign n21946 = ~n21941 & n21945 ;
  assign n21947 = ~n21944 & n21946 ;
  assign n21948 = ~n21938 & n21947 ;
  assign n21949 = n9241 & ~n21948 ;
  assign n21950 = ~n21931 & ~n21949 ;
  assign n21951 = \P1_P3_EAX_reg[31]/NET0131  & ~n16968 ;
  assign n21956 = ~n9060 & n16985 ;
  assign n21957 = ~n9089 & ~n21956 ;
  assign n21958 = ~n21684 & n21957 ;
  assign n21959 = \P1_P3_EAX_reg[31]/NET0131  & ~n21958 ;
  assign n21953 = n9049 & ~n21717 ;
  assign n21952 = ~\P1_P3_EAX_reg[31]/NET0131  & ~n9049 ;
  assign n21954 = n9060 & ~n21952 ;
  assign n21955 = ~n21953 & n21954 ;
  assign n21960 = ~\P1_P3_EAX_reg[31]/NET0131  & n16982 ;
  assign n21961 = n21683 & n21960 ;
  assign n21962 = ~n21955 & ~n21961 ;
  assign n21963 = ~n21959 & n21962 ;
  assign n21964 = n9241 & ~n21963 ;
  assign n21965 = ~n21951 & ~n21964 ;
  assign n21966 = ~n9199 & n9241 ;
  assign n21967 = \P1_P3_Flush_reg/NET0131  & ~n16968 ;
  assign n21968 = ~n21966 & ~n21967 ;
  assign n21969 = ~n9101 & n9241 ;
  assign n21970 = \P1_P3_More_reg/NET0131  & ~n16968 ;
  assign n21971 = ~n21969 & ~n21970 ;
  assign n21972 = ~\P3_rd_reg/NET0131  & \P4_reg3_reg[11]/NET0131  ;
  assign n21973 = ~n15982 & n16426 ;
  assign n21974 = n15976 & ~n18460 ;
  assign n21975 = ~n18461 & ~n21974 ;
  assign n21976 = ~\P4_IR_reg[28]/NET0131  & ~n21975 ;
  assign n21977 = \P4_IR_reg[28]/NET0131  & n16006 ;
  assign n21978 = ~n21976 & ~n21977 ;
  assign n21979 = n18483 & n21978 ;
  assign n21989 = ~n16269 & n18552 ;
  assign n21988 = n16269 & ~n18552 ;
  assign n21990 = n18490 & ~n21988 ;
  assign n21991 = ~n21989 & n21990 ;
  assign n21985 = n16269 & n18614 ;
  assign n21984 = ~n16269 & ~n18614 ;
  assign n21986 = n18607 & ~n21984 ;
  assign n21987 = ~n21985 & n21986 ;
  assign n21980 = ~n15982 & n18486 ;
  assign n21981 = ~n15982 & ~n18585 ;
  assign n21982 = ~n18586 & n18604 ;
  assign n21983 = ~n21981 & n21982 ;
  assign n21992 = ~n21980 & ~n21983 ;
  assign n21993 = ~n21987 & n21992 ;
  assign n21994 = ~n21991 & n21993 ;
  assign n21995 = ~n21979 & n21994 ;
  assign n21996 = n19076 & ~n21995 ;
  assign n21997 = ~n21973 & ~n21996 ;
  assign n21998 = n19075 & ~n21997 ;
  assign n21999 = n19075 & ~n19104 ;
  assign n22000 = ~n18607 & ~n18669 ;
  assign n22001 = ~n19076 & ~n22000 ;
  assign n22002 = ~n19156 & ~n22001 ;
  assign n22003 = n21999 & n22002 ;
  assign n22004 = n15987 & ~n22003 ;
  assign n22005 = ~n21998 & ~n22004 ;
  assign n22006 = \P3_rd_reg/NET0131  & ~n22005 ;
  assign n22007 = ~n21972 & ~n22006 ;
  assign n22008 = ~\P3_rd_reg/NET0131  & \P4_reg3_reg[12]/NET0131  ;
  assign n22009 = ~n15967 & n16426 ;
  assign n22020 = ~n16281 & n18691 ;
  assign n22019 = n16281 & ~n18691 ;
  assign n22021 = n18490 & ~n22019 ;
  assign n22022 = ~n22020 & n22021 ;
  assign n22011 = ~n15992 & ~n16160 ;
  assign n22013 = n16281 & ~n22011 ;
  assign n22012 = ~n16281 & n22011 ;
  assign n22014 = n18607 & ~n22012 ;
  assign n22015 = ~n22013 & n22014 ;
  assign n22010 = ~n15967 & n18486 ;
  assign n22016 = ~n15967 & ~n18586 ;
  assign n22017 = ~n18587 & n18604 ;
  assign n22018 = ~n22016 & n22017 ;
  assign n22023 = ~n22010 & ~n22018 ;
  assign n22024 = ~n22015 & n22023 ;
  assign n22025 = ~n22022 & n22024 ;
  assign n22026 = n15963 & ~n18461 ;
  assign n22027 = ~n18462 & ~n22026 ;
  assign n22028 = ~\P4_IR_reg[28]/NET0131  & ~n22027 ;
  assign n22029 = \P4_IR_reg[28]/NET0131  & n15991 ;
  assign n22030 = n18483 & ~n22029 ;
  assign n22031 = ~n22028 & n22030 ;
  assign n22032 = n22025 & ~n22031 ;
  assign n22033 = n19076 & ~n22032 ;
  assign n22034 = ~n22009 & ~n22033 ;
  assign n22035 = n19075 & ~n22034 ;
  assign n22036 = n15972 & ~n22003 ;
  assign n22037 = ~n22035 & ~n22036 ;
  assign n22038 = \P3_rd_reg/NET0131  & ~n22037 ;
  assign n22039 = ~n22008 & ~n22038 ;
  assign n22040 = ~\P3_rd_reg/NET0131  & \P4_reg3_reg[16]/NET0131  ;
  assign n22041 = ~n15940 & n16426 ;
  assign n22042 = n15936 & ~n19080 ;
  assign n22043 = n18464 & n19077 ;
  assign n22044 = ~n22042 & ~n22043 ;
  assign n22045 = ~\P4_IR_reg[28]/NET0131  & ~n22044 ;
  assign n22046 = \P4_IR_reg[28]/NET0131  & n16175 ;
  assign n22047 = ~n22045 & ~n22046 ;
  assign n22048 = n18483 & n22047 ;
  assign n22052 = ~n16332 & n18698 ;
  assign n22050 = ~n16324 & ~n18697 ;
  assign n22051 = ~n16334 & ~n22050 ;
  assign n22053 = n18490 & ~n22051 ;
  assign n22054 = ~n22052 & n22053 ;
  assign n22059 = n16198 & n16334 ;
  assign n22058 = ~n16198 & ~n16334 ;
  assign n22060 = n18607 & ~n22058 ;
  assign n22061 = ~n22059 & n22060 ;
  assign n22049 = ~n15940 & n18486 ;
  assign n22055 = ~n15940 & ~n18590 ;
  assign n22056 = ~n18591 & n18604 ;
  assign n22057 = ~n22055 & n22056 ;
  assign n22062 = ~n22049 & ~n22057 ;
  assign n22063 = ~n22061 & n22062 ;
  assign n22064 = ~n22054 & n22063 ;
  assign n22065 = ~n22048 & n22064 ;
  assign n22066 = n19076 & ~n22065 ;
  assign n22067 = ~n22041 & ~n22066 ;
  assign n22068 = n19075 & ~n22067 ;
  assign n22069 = n15945 & ~n22003 ;
  assign n22070 = ~n22068 & ~n22069 ;
  assign n22071 = \P3_rd_reg/NET0131  & ~n22070 ;
  assign n22072 = ~n22040 & ~n22071 ;
  assign n22073 = ~\P3_rd_reg/NET0131  & \P4_reg3_reg[7]/NET0131  ;
  assign n22074 = ~n16138 & n16426 ;
  assign n22075 = n16035 & ~n18456 ;
  assign n22076 = ~n18457 & ~n22075 ;
  assign n22077 = ~\P4_IR_reg[28]/NET0131  & ~n22076 ;
  assign n22078 = \P4_IR_reg[28]/NET0131  & n16131 ;
  assign n22079 = ~n22077 & ~n22078 ;
  assign n22080 = n18483 & n22079 ;
  assign n22091 = ~n16286 & n18549 ;
  assign n22090 = n16286 & ~n18549 ;
  assign n22092 = n18490 & ~n22090 ;
  assign n22093 = ~n22091 & n22092 ;
  assign n22084 = n16151 & ~n16153 ;
  assign n22082 = ~n16135 & ~n16149 ;
  assign n22083 = ~n16286 & ~n22082 ;
  assign n22085 = n18607 & ~n22083 ;
  assign n22086 = ~n22084 & n22085 ;
  assign n22081 = ~n16138 & n18486 ;
  assign n22087 = ~n16138 & ~n18581 ;
  assign n22088 = ~n18582 & n18604 ;
  assign n22089 = ~n22087 & n22088 ;
  assign n22094 = ~n22081 & ~n22089 ;
  assign n22095 = ~n22086 & n22094 ;
  assign n22096 = ~n22093 & n22095 ;
  assign n22097 = ~n22080 & n22096 ;
  assign n22098 = n19076 & ~n22097 ;
  assign n22099 = ~n22074 & ~n22098 ;
  assign n22100 = n19075 & ~n22099 ;
  assign n22101 = n16143 & ~n22003 ;
  assign n22102 = ~n22100 & ~n22101 ;
  assign n22103 = \P3_rd_reg/NET0131  & ~n22102 ;
  assign n22104 = ~n22073 & ~n22103 ;
  assign n22108 = ~\P1_P3_State_reg[2]/NET0131  & hold_pad ;
  assign n22109 = ~n8741 & ~n22108 ;
  assign n22110 = ~\P1_P3_State_reg[0]/NET0131  & ~\P1_P3_State_reg[2]/NET0131  ;
  assign n22111 = \P1_P3_State_reg[1]/NET0131  & ~n22110 ;
  assign n22112 = ~n22109 & n22111 ;
  assign n22105 = \P1_P3_State_reg[2]/NET0131  & hold_pad ;
  assign n22106 = \P1_P3_RequestPending_reg/NET0131  & \P1_P3_State_reg[0]/NET0131  ;
  assign n22107 = ~n22105 & n22106 ;
  assign n22113 = n9095 & ~n22107 ;
  assign n22114 = ~n22112 & n22113 ;
  assign n22115 = \P1_P3_State_reg[2]/NET0131  & n9091 ;
  assign n22116 = ~\P1_P3_State_reg[0]/NET0131  & na_pad ;
  assign n22117 = \P1_P3_State_reg[2]/NET0131  & ~n22116 ;
  assign n22118 = \P1_P3_State_reg[0]/NET0131  & ~n8741 ;
  assign n22119 = ~n22117 & ~n22118 ;
  assign n22120 = ~hold_pad & ~n22119 ;
  assign n22121 = \P1_P3_State_reg[0]/NET0131  & ~\P1_P3_State_reg[1]/NET0131  ;
  assign n22122 = ~\P1_P3_State_reg[2]/NET0131  & n22121 ;
  assign n22123 = ~n22120 & ~n22122 ;
  assign n22124 = \P1_P3_RequestPending_reg/NET0131  & ~n22123 ;
  assign n22125 = ~n22115 & ~n22124 ;
  assign n22126 = n15816 & n19073 ;
  assign n22127 = n15811 & n18486 ;
  assign n22128 = ~n18707 & n18710 ;
  assign n22129 = n18491 & n18683 ;
  assign n22130 = ~n22128 & n22129 ;
  assign n22131 = n18491 & ~n18713 ;
  assign n22132 = n18719 & ~n22131 ;
  assign n22133 = ~n22130 & n22132 ;
  assign n22135 = n16331 & ~n22133 ;
  assign n22134 = ~n16331 & n22133 ;
  assign n22136 = n18490 & ~n22134 ;
  assign n22137 = ~n22135 & n22136 ;
  assign n22138 = ~n16223 & ~n16229 ;
  assign n22140 = n16331 & n22138 ;
  assign n22139 = ~n16331 & ~n22138 ;
  assign n22141 = n18607 & ~n22139 ;
  assign n22142 = ~n22140 & n22141 ;
  assign n22143 = n15811 & ~n18600 ;
  assign n22144 = ~n18601 & n18604 ;
  assign n22145 = ~n22143 & n22144 ;
  assign n22146 = ~n22142 & ~n22145 ;
  assign n22147 = ~n22137 & n22146 ;
  assign n22148 = ~n22127 & n22147 ;
  assign n22149 = ~n15820 & n18474 ;
  assign n22150 = n15809 & ~n22149 ;
  assign n22151 = ~n18476 & ~n22150 ;
  assign n22152 = ~\P4_IR_reg[28]/NET0131  & ~n22151 ;
  assign n22153 = \P4_IR_reg[28]/NET0131  & n15832 ;
  assign n22154 = ~n22152 & ~n22153 ;
  assign n22155 = n18483 & n22154 ;
  assign n22156 = n22148 & ~n22155 ;
  assign n22157 = n19076 & ~n22156 ;
  assign n22158 = n15811 & n16426 ;
  assign n22159 = n18483 & ~n19076 ;
  assign n22160 = n19177 & ~n22159 ;
  assign n22161 = n15816 & ~n22160 ;
  assign n22162 = ~n22158 & ~n22161 ;
  assign n22163 = ~n22157 & n22162 ;
  assign n22164 = n19075 & ~n22163 ;
  assign n22165 = ~n22126 & ~n22164 ;
  assign n22166 = \P3_rd_reg/NET0131  & ~n22165 ;
  assign n22167 = n15744 & n15816 ;
  assign n22168 = ~\P3_rd_reg/NET0131  & \P4_reg3_reg[26]/NET0131  ;
  assign n22169 = ~n22167 & ~n22168 ;
  assign n22170 = ~n22166 & n22169 ;
  assign n22171 = ~n16426 & ~n20673 ;
  assign n22172 = n18666 & ~n19104 ;
  assign n22173 = ~n22171 & n22172 ;
  assign n22174 = \P4_reg2_reg[31]/NET0131  & ~n22173 ;
  assign n22175 = ~n16245 & n21826 ;
  assign n22176 = n18604 & ~n22175 ;
  assign n22178 = ~n16244 & n21789 ;
  assign n22177 = n16244 & ~n21789 ;
  assign n22179 = n18483 & ~n21788 ;
  assign n22180 = ~n22177 & n22179 ;
  assign n22181 = ~n22178 & n22180 ;
  assign n22182 = ~n22176 & ~n22181 ;
  assign n22183 = n20673 & ~n22182 ;
  assign n22184 = ~n21841 & ~n22183 ;
  assign n22185 = n18666 & ~n22184 ;
  assign n22186 = ~n22174 & ~n22185 ;
  assign n22188 = n15852 & n19073 ;
  assign n22192 = n15852 & ~n19076 ;
  assign n22193 = n19076 & n21871 ;
  assign n22194 = ~n22192 & ~n22193 ;
  assign n22195 = n18483 & ~n22194 ;
  assign n22196 = n21893 & ~n21908 ;
  assign n22197 = n19076 & ~n22196 ;
  assign n22198 = ~n22192 & ~n22197 ;
  assign n22199 = ~n18607 & ~n19176 ;
  assign n22200 = ~n21908 & n22199 ;
  assign n22201 = ~n22198 & ~n22200 ;
  assign n22202 = n19076 & n21877 ;
  assign n22203 = ~n22192 & ~n22202 ;
  assign n22204 = n18604 & ~n22203 ;
  assign n22189 = n18486 & n19076 ;
  assign n22190 = ~n16426 & ~n22189 ;
  assign n22191 = n15847 & ~n22190 ;
  assign n22205 = ~n18486 & ~n19104 ;
  assign n22206 = ~n19157 & ~n22205 ;
  assign n22207 = n15852 & n22206 ;
  assign n22208 = ~n22191 & ~n22207 ;
  assign n22209 = ~n22204 & n22208 ;
  assign n22210 = ~n22201 & n22209 ;
  assign n22211 = ~n22195 & n22210 ;
  assign n22212 = n19075 & ~n22211 ;
  assign n22213 = ~n22188 & ~n22212 ;
  assign n22214 = \P3_rd_reg/NET0131  & ~n22213 ;
  assign n22187 = ~\P3_rd_reg/NET0131  & \P4_reg3_reg[23]/NET0131  ;
  assign n22215 = n15744 & n15852 ;
  assign n22216 = ~n22187 & ~n22215 ;
  assign n22217 = ~n22214 & n22216 ;
  assign n22218 = \P4_reg2_reg[24]/NET0131  & ~n18665 ;
  assign n22237 = \P4_IR_reg[28]/NET0131  & ~n15856 ;
  assign n22238 = n15832 & ~n21866 ;
  assign n22239 = ~\P4_IR_reg[28]/NET0131  & ~n18474 ;
  assign n22240 = ~n22238 & n22239 ;
  assign n22241 = ~n22237 & ~n22240 ;
  assign n22242 = n20673 & n22241 ;
  assign n22243 = ~\P4_reg2_reg[24]/NET0131  & ~n20673 ;
  assign n22244 = n18483 & ~n22243 ;
  assign n22245 = ~n22242 & n22244 ;
  assign n22229 = ~n16278 & n18715 ;
  assign n22228 = n16278 & ~n18715 ;
  assign n22230 = n18490 & ~n22228 ;
  assign n22231 = ~n22229 & n22230 ;
  assign n22225 = ~n16222 & ~n16278 ;
  assign n22224 = n16222 & n16278 ;
  assign n22226 = n18607 & ~n22224 ;
  assign n22227 = ~n22225 & n22226 ;
  assign n22220 = n15834 & n18486 ;
  assign n22221 = n15834 & ~n18598 ;
  assign n22222 = ~n18599 & n18604 ;
  assign n22223 = ~n22221 & n22222 ;
  assign n22232 = ~n22220 & ~n22223 ;
  assign n22233 = ~n22227 & n22232 ;
  assign n22234 = ~n22231 & n22233 ;
  assign n22235 = n20673 & ~n22234 ;
  assign n22219 = \P4_reg2_reg[24]/NET0131  & ~n20682 ;
  assign n22236 = n15840 & n16426 ;
  assign n22246 = ~n22219 & ~n22236 ;
  assign n22247 = ~n22235 & n22246 ;
  assign n22248 = ~n22245 & n22247 ;
  assign n22249 = n19075 & ~n22248 ;
  assign n22250 = \P4_reg2_reg[24]/NET0131  & n19073 ;
  assign n22251 = ~n22249 & ~n22250 ;
  assign n22252 = \P3_rd_reg/NET0131  & ~n22251 ;
  assign n22253 = ~n22218 & ~n22252 ;
  assign n22254 = \P4_reg2_reg[26]/NET0131  & n19073 ;
  assign n22255 = \P4_reg2_reg[26]/NET0131  & ~n20673 ;
  assign n22256 = n20673 & n22154 ;
  assign n22257 = ~n22255 & ~n22256 ;
  assign n22258 = n18483 & ~n22257 ;
  assign n22263 = n20673 & ~n22147 ;
  assign n22264 = n15816 & n16426 ;
  assign n22259 = n18488 & ~n18604 ;
  assign n22260 = ~n20681 & n22259 ;
  assign n22261 = ~n20678 & ~n22260 ;
  assign n22262 = \P4_reg2_reg[26]/NET0131  & n22261 ;
  assign n22265 = n15811 & n20673 ;
  assign n22266 = ~n22255 & ~n22265 ;
  assign n22267 = n18486 & ~n22266 ;
  assign n22268 = ~n22262 & ~n22267 ;
  assign n22269 = ~n22264 & n22268 ;
  assign n22270 = ~n22263 & n22269 ;
  assign n22271 = ~n22258 & n22270 ;
  assign n22272 = n19075 & ~n22271 ;
  assign n22273 = ~n22254 & ~n22272 ;
  assign n22274 = \P3_rd_reg/NET0131  & ~n22273 ;
  assign n22275 = \P4_reg2_reg[26]/NET0131  & ~n18665 ;
  assign n22276 = ~n22274 & ~n22275 ;
  assign n22277 = \P4_reg0_reg[11]/NET0131  & ~n21855 ;
  assign n22278 = n20665 & ~n21995 ;
  assign n22279 = ~n22277 & ~n22278 ;
  assign n22281 = \P4_reg0_reg[23]/NET0131  & ~n20661 ;
  assign n22282 = n20665 & n21871 ;
  assign n22283 = ~n22281 & ~n22282 ;
  assign n22284 = n18483 & ~n22283 ;
  assign n22280 = \P4_reg0_reg[23]/NET0131  & ~n21854 ;
  assign n22285 = n20665 & ~n21911 ;
  assign n22286 = ~n22280 & ~n22285 ;
  assign n22287 = ~n22284 & n22286 ;
  assign n22289 = \P4_reg0_reg[26]/NET0131  & ~n20661 ;
  assign n22290 = n20665 & n22154 ;
  assign n22291 = ~n22289 & ~n22290 ;
  assign n22292 = n18483 & ~n22291 ;
  assign n22288 = n20665 & ~n22148 ;
  assign n22293 = \P4_reg0_reg[26]/NET0131  & ~n21854 ;
  assign n22294 = ~n22288 & ~n22293 ;
  assign n22295 = ~n22292 & n22294 ;
  assign n22296 = \P4_reg1_reg[24]/NET0131  & ~n18679 ;
  assign n22297 = n18483 & ~n22241 ;
  assign n22298 = n22234 & ~n22297 ;
  assign n22299 = n18667 & ~n22298 ;
  assign n22300 = ~n22296 & ~n22299 ;
  assign n22301 = n18667 & ~n22156 ;
  assign n22302 = ~n18670 & n22127 ;
  assign n22303 = n18679 & ~n22302 ;
  assign n22304 = \P4_reg1_reg[26]/NET0131  & ~n22303 ;
  assign n22305 = ~n22301 & ~n22304 ;
  assign n22306 = \P4_reg2_reg[23]/NET0131  & ~n18665 ;
  assign n22308 = \P4_reg2_reg[23]/NET0131  & ~n20673 ;
  assign n22309 = n20673 & n21871 ;
  assign n22310 = ~n22308 & ~n22309 ;
  assign n22311 = n18483 & ~n22310 ;
  assign n22312 = n20673 & ~n22196 ;
  assign n22313 = ~n22308 & ~n22312 ;
  assign n22314 = ~n18607 & ~n20681 ;
  assign n22315 = ~n21908 & n22314 ;
  assign n22316 = ~n22313 & ~n22315 ;
  assign n22317 = n20673 & n21877 ;
  assign n22318 = ~n22308 & ~n22317 ;
  assign n22319 = n18604 & ~n22318 ;
  assign n22307 = n15852 & n16426 ;
  assign n22320 = n20673 & n21875 ;
  assign n22321 = ~n20678 & ~n22205 ;
  assign n22322 = \P4_reg2_reg[23]/NET0131  & n22321 ;
  assign n22323 = ~n22320 & ~n22322 ;
  assign n22324 = ~n22307 & n22323 ;
  assign n22325 = ~n22319 & n22324 ;
  assign n22326 = ~n22316 & n22325 ;
  assign n22327 = ~n22311 & n22326 ;
  assign n22328 = n19075 & ~n22327 ;
  assign n22329 = \P4_reg2_reg[23]/NET0131  & n19073 ;
  assign n22330 = ~n22328 & ~n22329 ;
  assign n22331 = \P3_rd_reg/NET0131  & ~n22330 ;
  assign n22332 = ~n22306 & ~n22331 ;
  assign n22333 = \P2_P1_EAX_reg[30]/NET0131  & ~n21100 ;
  assign n22337 = ~n21073 & ~n21081 ;
  assign n22338 = ~n11569 & n22337 ;
  assign n22339 = \P2_P1_EAX_reg[30]/NET0131  & ~n22337 ;
  assign n22340 = ~n22338 & ~n22339 ;
  assign n22341 = n21068 & ~n22340 ;
  assign n22342 = n21022 & ~n21051 ;
  assign n22343 = ~n21072 & ~n22342 ;
  assign n22344 = \P2_P1_EAX_reg[30]/NET0131  & ~n22343 ;
  assign n22348 = ~\P2_P1_EAX_reg[30]/NET0131  & n21022 ;
  assign n22349 = n21051 & n22348 ;
  assign n22334 = ~n20983 & n21014 ;
  assign n22335 = ~n21015 & ~n22334 ;
  assign n22336 = n20728 & n22335 ;
  assign n22345 = n11381 & n22337 ;
  assign n22346 = ~n22339 & ~n22345 ;
  assign n22347 = n21062 & ~n22346 ;
  assign n22350 = ~n22336 & ~n22347 ;
  assign n22351 = ~n22349 & n22350 ;
  assign n22352 = ~n22344 & n22351 ;
  assign n22353 = ~n22341 & n22352 ;
  assign n22354 = n11623 & ~n22353 ;
  assign n22355 = ~n22333 & ~n22354 ;
  assign n22356 = \P1_P3_EAX_reg[25]/NET0131  & ~n16968 ;
  assign n22360 = \P1_P3_EAX_reg[25]/NET0131  & n21476 ;
  assign n22361 = n16982 & ~n22360 ;
  assign n22362 = ~n16987 & ~n22361 ;
  assign n22363 = \P1_P3_EAX_reg[25]/NET0131  & ~n22362 ;
  assign n22364 = n21476 & n22361 ;
  assign n22365 = \P1_P3_EAX_reg[25]/NET0131  & ~n9088 ;
  assign n22368 = \P1_buf2_reg[25]/NET0131  & n9088 ;
  assign n22369 = ~n22365 & ~n22368 ;
  assign n22370 = n9086 & ~n22369 ;
  assign n22357 = ~n21466 & n21534 ;
  assign n22358 = ~n21535 & ~n22357 ;
  assign n22359 = n16984 & n22358 ;
  assign n22366 = ~n17336 & ~n22365 ;
  assign n22367 = n9085 & ~n22366 ;
  assign n22371 = ~n22359 & ~n22367 ;
  assign n22372 = ~n22370 & n22371 ;
  assign n22373 = ~n22364 & n22372 ;
  assign n22374 = ~n22363 & n22373 ;
  assign n22375 = n9241 & ~n22374 ;
  assign n22376 = ~n22356 & ~n22375 ;
  assign n22377 = \P1_P3_EAX_reg[26]/NET0131  & ~n16968 ;
  assign n22381 = \P1_P3_EAX_reg[26]/NET0131  & ~n22362 ;
  assign n22388 = ~\P1_P3_EAX_reg[26]/NET0131  & n16982 ;
  assign n22389 = n22360 & n22388 ;
  assign n22382 = \P1_P3_EAX_reg[26]/NET0131  & ~n9088 ;
  assign n22386 = ~n17123 & ~n22382 ;
  assign n22387 = n9085 & ~n22386 ;
  assign n22378 = ~n21535 & n21566 ;
  assign n22379 = ~n21567 & ~n22378 ;
  assign n22380 = n16984 & n22379 ;
  assign n22383 = \P1_buf2_reg[26]/NET0131  & n9088 ;
  assign n22384 = ~n22382 & ~n22383 ;
  assign n22385 = n9086 & ~n22384 ;
  assign n22390 = ~n22380 & ~n22385 ;
  assign n22391 = ~n22387 & n22390 ;
  assign n22392 = ~n22389 & n22391 ;
  assign n22393 = ~n22381 & n22392 ;
  assign n22394 = n9241 & ~n22393 ;
  assign n22395 = ~n22377 & ~n22394 ;
  assign n22396 = \P1_P3_EAX_reg[27]/NET0131  & ~n16968 ;
  assign n22399 = \P1_P3_EAX_reg[27]/NET0131  & ~n21937 ;
  assign n22397 = \P1_P3_EAX_reg[26]/NET0131  & n21936 ;
  assign n22398 = n22360 & n22397 ;
  assign n22400 = \P1_P3_EAX_reg[27]/NET0131  & ~n9088 ;
  assign n22406 = \P1_buf2_reg[27]/NET0131  & n9088 ;
  assign n22407 = ~n22400 & ~n22406 ;
  assign n22408 = n9086 & ~n22407 ;
  assign n22401 = ~n16970 & ~n22400 ;
  assign n22402 = n9085 & ~n22401 ;
  assign n22403 = ~n21567 & n21598 ;
  assign n22404 = ~n21599 & ~n22403 ;
  assign n22405 = n16984 & n22404 ;
  assign n22409 = ~n22402 & ~n22405 ;
  assign n22410 = ~n22408 & n22409 ;
  assign n22411 = ~n22398 & n22410 ;
  assign n22412 = ~n22399 & n22411 ;
  assign n22413 = n9241 & ~n22412 ;
  assign n22414 = ~n22396 & ~n22413 ;
  assign n22417 = n16002 & n19073 ;
  assign n22420 = ~n15997 & n18486 ;
  assign n22429 = ~n16285 & n18687 ;
  assign n22428 = n16285 & ~n18687 ;
  assign n22430 = n18490 & ~n22428 ;
  assign n22431 = ~n22429 & n22430 ;
  assign n22421 = ~n15997 & ~n18584 ;
  assign n22422 = ~n18585 & n18604 ;
  assign n22423 = ~n22421 & n22422 ;
  assign n22425 = n16158 & ~n16285 ;
  assign n22424 = ~n16158 & n16285 ;
  assign n22426 = n18607 & ~n22424 ;
  assign n22427 = ~n22425 & n22426 ;
  assign n22432 = ~n22423 & ~n22427 ;
  assign n22433 = ~n22431 & n22432 ;
  assign n22434 = ~n22420 & n22433 ;
  assign n22435 = n15991 & ~n18459 ;
  assign n22436 = ~n18460 & ~n22435 ;
  assign n22437 = ~\P4_IR_reg[28]/NET0131  & ~n22436 ;
  assign n22438 = \P4_IR_reg[28]/NET0131  & n16021 ;
  assign n22439 = ~n22437 & ~n22438 ;
  assign n22440 = n18483 & n22439 ;
  assign n22441 = n22434 & ~n22440 ;
  assign n22442 = n19076 & ~n22441 ;
  assign n22418 = ~n15997 & n16426 ;
  assign n22419 = n16002 & ~n22160 ;
  assign n22443 = ~n22418 & ~n22419 ;
  assign n22444 = ~n22442 & n22443 ;
  assign n22445 = n19075 & ~n22444 ;
  assign n22446 = ~n22417 & ~n22445 ;
  assign n22447 = \P3_rd_reg/NET0131  & ~n22446 ;
  assign n22415 = ~\P3_rd_reg/NET0131  & \P4_reg3_reg[10]/NET0131  ;
  assign n22416 = n15744 & n16002 ;
  assign n22448 = ~n22415 & ~n22416 ;
  assign n22449 = ~n22447 & n22448 ;
  assign n22450 = ~\P3_rd_reg/NET0131  & \P4_reg3_reg[14]/NET0131  ;
  assign n22451 = ~n16179 & n16426 ;
  assign n22452 = n16175 & ~n19077 ;
  assign n22453 = ~n19078 & ~n22452 ;
  assign n22454 = ~\P4_IR_reg[28]/NET0131  & ~n22453 ;
  assign n22455 = \P4_IR_reg[28]/NET0131  & n15963 ;
  assign n22456 = ~n22454 & ~n22455 ;
  assign n22457 = n18483 & n22456 ;
  assign n22459 = ~n16264 & ~n18694 ;
  assign n22461 = n16335 & ~n22459 ;
  assign n22460 = ~n16335 & n22459 ;
  assign n22462 = n18490 & ~n22460 ;
  assign n22463 = ~n22461 & n22462 ;
  assign n22464 = ~n16162 & ~n16190 ;
  assign n22466 = ~n16335 & ~n22464 ;
  assign n22465 = n16335 & n22464 ;
  assign n22467 = n18607 & ~n22465 ;
  assign n22468 = ~n22466 & n22467 ;
  assign n22458 = ~n16179 & n18486 ;
  assign n22469 = ~n16179 & ~n18588 ;
  assign n22470 = ~n18589 & n18604 ;
  assign n22471 = ~n22469 & n22470 ;
  assign n22472 = ~n22458 & ~n22471 ;
  assign n22473 = ~n22468 & n22472 ;
  assign n22474 = ~n22463 & n22473 ;
  assign n22475 = ~n22457 & n22474 ;
  assign n22476 = n19076 & ~n22475 ;
  assign n22477 = ~n22451 & ~n22476 ;
  assign n22478 = n19075 & ~n22477 ;
  assign n22479 = n16184 & ~n22003 ;
  assign n22480 = ~n22478 & ~n22479 ;
  assign n22481 = \P3_rd_reg/NET0131  & ~n22480 ;
  assign n22482 = ~n22450 & ~n22481 ;
  assign n22484 = n15891 & n19073 ;
  assign n22486 = \P4_IR_reg[28]/NET0131  & ~n15909 ;
  assign n22487 = ~n15909 & n18467 ;
  assign n22488 = ~n15895 & n22487 ;
  assign n22489 = n15884 & ~n22488 ;
  assign n22490 = ~\P4_IR_reg[28]/NET0131  & ~n18470 ;
  assign n22491 = ~n22489 & n22490 ;
  assign n22492 = ~n22486 & ~n22491 ;
  assign n22493 = n18483 & ~n22492 ;
  assign n22504 = n16259 & ~n18705 ;
  assign n22503 = ~n16259 & n18705 ;
  assign n22505 = n18490 & ~n22503 ;
  assign n22506 = ~n22504 & n22505 ;
  assign n22495 = n16210 & n16259 ;
  assign n22494 = ~n16210 & ~n16259 ;
  assign n22496 = n18607 & ~n22494 ;
  assign n22497 = ~n22495 & n22496 ;
  assign n22498 = n15886 & n18486 ;
  assign n22499 = n15886 & ~n18594 ;
  assign n22500 = ~n18595 & n18604 ;
  assign n22501 = ~n22499 & n22500 ;
  assign n22502 = ~n22498 & ~n22501 ;
  assign n22507 = ~n22497 & n22502 ;
  assign n22508 = ~n22506 & n22507 ;
  assign n22509 = ~n22493 & n22508 ;
  assign n22510 = n19076 & ~n22509 ;
  assign n22485 = n15886 & n16426 ;
  assign n22511 = n15891 & ~n22160 ;
  assign n22512 = ~n22485 & ~n22511 ;
  assign n22513 = ~n22510 & n22512 ;
  assign n22514 = n19075 & ~n22513 ;
  assign n22515 = ~n22484 & ~n22514 ;
  assign n22516 = \P3_rd_reg/NET0131  & ~n22515 ;
  assign n22483 = ~\P3_rd_reg/NET0131  & \P4_reg3_reg[20]/NET0131  ;
  assign n22517 = n15744 & n15891 ;
  assign n22518 = ~n22483 & ~n22517 ;
  assign n22519 = ~n22516 & n22518 ;
  assign n22520 = ~\P3_rd_reg/NET0131  & \P4_reg3_reg[19]/NET0131  ;
  assign n22521 = ~n15900 & n16426 ;
  assign n22522 = n15895 & ~n22487 ;
  assign n22523 = ~n22488 & ~n22522 ;
  assign n22524 = ~\P4_IR_reg[28]/NET0131  & ~n22523 ;
  assign n22525 = \P4_IR_reg[28]/NET0131  & n15922 ;
  assign n22526 = ~n22524 & ~n22525 ;
  assign n22527 = n18483 & n22526 ;
  assign n22537 = ~n16316 & n18630 ;
  assign n22536 = n16316 & ~n18630 ;
  assign n22538 = n18607 & ~n22536 ;
  assign n22539 = ~n22537 & n22538 ;
  assign n22533 = ~n16316 & ~n18556 ;
  assign n22532 = n16316 & n18556 ;
  assign n22534 = n18490 & ~n22532 ;
  assign n22535 = ~n22533 & n22534 ;
  assign n22528 = ~n15900 & n18486 ;
  assign n22529 = ~n15900 & ~n18593 ;
  assign n22530 = ~n18594 & n18604 ;
  assign n22531 = ~n22529 & n22530 ;
  assign n22540 = ~n22528 & ~n22531 ;
  assign n22541 = ~n22535 & n22540 ;
  assign n22542 = ~n22539 & n22541 ;
  assign n22543 = ~n22527 & n22542 ;
  assign n22544 = n19076 & ~n22543 ;
  assign n22545 = ~n22521 & ~n22544 ;
  assign n22546 = n19075 & ~n22545 ;
  assign n22547 = n15905 & ~n22003 ;
  assign n22548 = ~n22546 & ~n22547 ;
  assign n22549 = \P3_rd_reg/NET0131  & ~n22548 ;
  assign n22550 = ~n22520 & ~n22549 ;
  assign n22551 = ~\P3_rd_reg/NET0131  & \P4_reg3_reg[24]/NET0131  ;
  assign n22552 = n15834 & n16426 ;
  assign n22553 = n19076 & ~n22298 ;
  assign n22554 = ~n22552 & ~n22553 ;
  assign n22555 = n19075 & ~n22554 ;
  assign n22556 = n15840 & ~n22003 ;
  assign n22557 = ~n22555 & ~n22556 ;
  assign n22558 = \P3_rd_reg/NET0131  & ~n22557 ;
  assign n22559 = ~n22551 & ~n22558 ;
  assign n22560 = \P4_reg2_reg[20]/NET0131  & ~n18665 ;
  assign n22561 = \P4_reg2_reg[20]/NET0131  & n19073 ;
  assign n22563 = n20673 & ~n22509 ;
  assign n22562 = n15891 & n16426 ;
  assign n22564 = ~n19106 & ~n20673 ;
  assign n22565 = ~n22321 & ~n22564 ;
  assign n22566 = \P4_reg2_reg[20]/NET0131  & ~n22565 ;
  assign n22567 = ~n22562 & ~n22566 ;
  assign n22568 = ~n22563 & n22567 ;
  assign n22569 = n19075 & ~n22568 ;
  assign n22570 = ~n22561 & ~n22569 ;
  assign n22571 = \P3_rd_reg/NET0131  & ~n22570 ;
  assign n22572 = ~n22560 & ~n22571 ;
  assign n22573 = n18666 & ~n20680 ;
  assign n22574 = ~n20679 & n22573 ;
  assign n22575 = \P4_reg2_reg[22]/NET0131  & ~n22574 ;
  assign n22576 = n15868 & n16426 ;
  assign n22577 = ~n15872 & n18470 ;
  assign n22578 = n15856 & ~n22577 ;
  assign n22579 = ~n18472 & ~n22578 ;
  assign n22580 = ~\P4_IR_reg[28]/NET0131  & ~n22579 ;
  assign n22581 = \P4_IR_reg[28]/NET0131  & n15884 ;
  assign n22582 = ~n22580 & ~n22581 ;
  assign n22583 = n18483 & n22582 ;
  assign n22593 = ~n16322 & n22128 ;
  assign n22592 = n16322 & ~n22128 ;
  assign n22594 = n18490 & ~n22592 ;
  assign n22595 = ~n22593 & n22594 ;
  assign n22589 = ~n16216 & ~n16322 ;
  assign n22588 = n16216 & n16322 ;
  assign n22590 = n18607 & ~n22588 ;
  assign n22591 = ~n22589 & n22590 ;
  assign n22584 = n15858 & n18486 ;
  assign n22585 = n15858 & ~n18596 ;
  assign n22586 = ~n18597 & n18604 ;
  assign n22587 = ~n22585 & n22586 ;
  assign n22596 = ~n22584 & ~n22587 ;
  assign n22597 = ~n22591 & n22596 ;
  assign n22598 = ~n22595 & n22597 ;
  assign n22599 = ~n22583 & n22598 ;
  assign n22600 = n20673 & ~n22599 ;
  assign n22601 = ~n22576 & ~n22600 ;
  assign n22602 = n18666 & ~n22601 ;
  assign n22603 = ~n22575 & ~n22602 ;
  assign n22604 = \P4_reg0_reg[12]/NET0131  & ~n21855 ;
  assign n22605 = n20665 & ~n22032 ;
  assign n22606 = ~n22604 & ~n22605 ;
  assign n22607 = \P4_reg0_reg[16]/NET0131  & ~n21855 ;
  assign n22608 = n20665 & ~n22065 ;
  assign n22609 = ~n22607 & ~n22608 ;
  assign n22610 = \P4_reg0_reg[19]/NET0131  & ~n21855 ;
  assign n22611 = n20665 & ~n22543 ;
  assign n22612 = ~n22610 & ~n22611 ;
  assign n22613 = \P4_reg0_reg[20]/NET0131  & ~n18665 ;
  assign n22614 = \P4_reg0_reg[20]/NET0131  & n19073 ;
  assign n22622 = n20661 & n22492 ;
  assign n22617 = ~\P4_reg0_reg[20]/NET0131  & ~n20661 ;
  assign n22623 = n18483 & ~n22617 ;
  assign n22624 = ~n22622 & n22623 ;
  assign n22618 = n20661 & ~n22497 ;
  assign n22619 = ~n22506 & n22618 ;
  assign n22620 = ~n18672 & ~n22617 ;
  assign n22621 = ~n22619 & n22620 ;
  assign n22615 = \P4_reg0_reg[20]/NET0131  & n21851 ;
  assign n22616 = n20661 & ~n22502 ;
  assign n22625 = ~n22615 & ~n22616 ;
  assign n22626 = ~n22621 & n22625 ;
  assign n22627 = ~n22624 & n22626 ;
  assign n22628 = n19075 & ~n22627 ;
  assign n22629 = ~n22614 & ~n22628 ;
  assign n22630 = \P3_rd_reg/NET0131  & ~n22629 ;
  assign n22631 = ~n22613 & ~n22630 ;
  assign n22632 = \P4_reg0_reg[24]/NET0131  & ~n21855 ;
  assign n22633 = n20665 & ~n22298 ;
  assign n22634 = ~n22632 & ~n22633 ;
  assign n22635 = \P4_reg0_reg[29]/NET0131  & ~n21855 ;
  assign n22636 = n18483 & ~n21792 ;
  assign n22637 = n21839 & ~n22636 ;
  assign n22638 = n20665 & ~n22637 ;
  assign n22639 = ~n22635 & ~n22638 ;
  assign n22640 = \P4_reg0_reg[30]/NET0131  & ~n18665 ;
  assign n22641 = \P4_reg0_reg[30]/NET0131  & n19073 ;
  assign n22642 = \P4_reg0_reg[30]/NET0131  & ~n20662 ;
  assign n22643 = n16245 & n18486 ;
  assign n22644 = n16245 & ~n21826 ;
  assign n22645 = n22176 & ~n22644 ;
  assign n22646 = ~n22643 & ~n22645 ;
  assign n22647 = ~n22181 & n22646 ;
  assign n22648 = n20661 & ~n22647 ;
  assign n22649 = ~n22642 & ~n22648 ;
  assign n22650 = n19075 & ~n22649 ;
  assign n22651 = ~n22641 & ~n22650 ;
  assign n22652 = \P3_rd_reg/NET0131  & ~n22651 ;
  assign n22653 = ~n22640 & ~n22652 ;
  assign n22654 = n20665 & ~n22182 ;
  assign n22655 = \P4_reg0_reg[31]/NET0131  & ~n20663 ;
  assign n22656 = ~n22654 & ~n22655 ;
  assign n22657 = \P4_reg0_reg[7]/NET0131  & ~n21855 ;
  assign n22658 = n20665 & ~n22097 ;
  assign n22659 = ~n22657 & ~n22658 ;
  assign n22660 = \P4_reg1_reg[11]/NET0131  & ~n18679 ;
  assign n22661 = n18667 & ~n21995 ;
  assign n22662 = ~n22660 & ~n22661 ;
  assign n22663 = \P4_reg1_reg[12]/NET0131  & ~n18679 ;
  assign n22664 = n18667 & ~n22032 ;
  assign n22665 = ~n22663 & ~n22664 ;
  assign n22666 = \P4_reg1_reg[16]/NET0131  & ~n18679 ;
  assign n22667 = n18667 & ~n22065 ;
  assign n22668 = ~n22666 & ~n22667 ;
  assign n22669 = \P4_reg1_reg[19]/NET0131  & ~n18679 ;
  assign n22670 = n18667 & ~n22543 ;
  assign n22671 = ~n22669 & ~n22670 ;
  assign n22673 = \P4_reg1_reg[22]/NET0131  & ~n18664 ;
  assign n22674 = n18667 & n22582 ;
  assign n22675 = ~n22673 & ~n22674 ;
  assign n22676 = n18483 & ~n22675 ;
  assign n22672 = n18667 & ~n22598 ;
  assign n22677 = \P4_reg1_reg[22]/NET0131  & ~n21863 ;
  assign n22678 = ~n22672 & ~n22677 ;
  assign n22679 = ~n22676 & n22678 ;
  assign n22680 = \P4_reg1_reg[29]/NET0131  & ~n18679 ;
  assign n22681 = n18667 & ~n22637 ;
  assign n22682 = ~n22680 & ~n22681 ;
  assign n22683 = \P4_reg1_reg[30]/NET0131  & ~n18665 ;
  assign n22684 = \P4_reg1_reg[30]/NET0131  & n19073 ;
  assign n22685 = n18664 & ~n18676 ;
  assign n22686 = \P4_reg1_reg[30]/NET0131  & ~n22685 ;
  assign n22687 = n18664 & ~n22647 ;
  assign n22688 = ~n22686 & ~n22687 ;
  assign n22689 = n19075 & ~n22688 ;
  assign n22690 = ~n22684 & ~n22689 ;
  assign n22691 = \P3_rd_reg/NET0131  & ~n22690 ;
  assign n22692 = ~n22683 & ~n22691 ;
  assign n22693 = n18667 & ~n22182 ;
  assign n22694 = n18664 & n18677 ;
  assign n22695 = \P4_reg1_reg[31]/NET0131  & ~n22694 ;
  assign n22696 = ~n22693 & ~n22695 ;
  assign n22697 = n18667 & ~n22097 ;
  assign n22698 = ~n18664 & ~n19109 ;
  assign n22699 = n18677 & ~n22698 ;
  assign n22700 = \P4_reg1_reg[7]/NET0131  & ~n22699 ;
  assign n22701 = ~n22697 & ~n22700 ;
  assign n22702 = \P4_reg2_reg[11]/NET0131  & ~n18665 ;
  assign n22703 = \P4_reg2_reg[11]/NET0131  & n19073 ;
  assign n22705 = n20673 & ~n21978 ;
  assign n22706 = ~\P4_reg2_reg[11]/NET0131  & ~n20673 ;
  assign n22707 = n18483 & ~n22706 ;
  assign n22708 = ~n22705 & n22707 ;
  assign n22709 = n20673 & ~n21994 ;
  assign n22704 = n15987 & n16426 ;
  assign n22710 = \P4_reg2_reg[11]/NET0131  & ~n20682 ;
  assign n22711 = ~n22704 & ~n22710 ;
  assign n22712 = ~n22709 & n22711 ;
  assign n22713 = ~n22708 & n22712 ;
  assign n22714 = n19075 & ~n22713 ;
  assign n22715 = ~n22703 & ~n22714 ;
  assign n22716 = \P3_rd_reg/NET0131  & ~n22715 ;
  assign n22717 = ~n22702 & ~n22716 ;
  assign n22718 = n15972 & n16426 ;
  assign n22719 = ~\P4_reg2_reg[12]/NET0131  & ~n20673 ;
  assign n22720 = n20673 & ~n22025 ;
  assign n22721 = n22573 & ~n22720 ;
  assign n22722 = ~n22031 & n22721 ;
  assign n22723 = ~n22719 & ~n22722 ;
  assign n22724 = ~n22718 & ~n22723 ;
  assign n22725 = ~\P4_reg2_reg[12]/NET0131  & ~n18666 ;
  assign n22726 = ~n22724 & ~n22725 ;
  assign n22727 = \P4_reg2_reg[12]/NET0131  & n20679 ;
  assign n22728 = ~n22726 & ~n22727 ;
  assign n22729 = \P4_reg2_reg[16]/NET0131  & ~n18665 ;
  assign n22730 = \P4_reg2_reg[16]/NET0131  & n19073 ;
  assign n22732 = n20673 & ~n22047 ;
  assign n22733 = ~\P4_reg2_reg[16]/NET0131  & ~n20673 ;
  assign n22734 = n18483 & ~n22733 ;
  assign n22735 = ~n22732 & n22734 ;
  assign n22736 = n20673 & ~n22064 ;
  assign n22731 = n15945 & n16426 ;
  assign n22737 = \P4_reg2_reg[16]/NET0131  & ~n20682 ;
  assign n22738 = ~n22731 & ~n22737 ;
  assign n22739 = ~n22736 & n22738 ;
  assign n22740 = ~n22735 & n22739 ;
  assign n22741 = n19075 & ~n22740 ;
  assign n22742 = ~n22730 & ~n22741 ;
  assign n22743 = \P3_rd_reg/NET0131  & ~n22742 ;
  assign n22744 = ~n22729 & ~n22743 ;
  assign n22745 = \P4_reg2_reg[19]/NET0131  & ~n18665 ;
  assign n22746 = \P4_reg2_reg[19]/NET0131  & n19073 ;
  assign n22748 = n20673 & ~n22526 ;
  assign n22749 = ~\P4_reg2_reg[19]/NET0131  & ~n20673 ;
  assign n22750 = n18483 & ~n22749 ;
  assign n22751 = ~n22748 & n22750 ;
  assign n22752 = n20673 & ~n22542 ;
  assign n22747 = n15905 & n16426 ;
  assign n22753 = \P4_reg2_reg[19]/NET0131  & ~n20682 ;
  assign n22754 = ~n22747 & ~n22753 ;
  assign n22755 = ~n22752 & n22754 ;
  assign n22756 = ~n22751 & n22755 ;
  assign n22757 = n19075 & ~n22756 ;
  assign n22758 = ~n22746 & ~n22757 ;
  assign n22759 = \P3_rd_reg/NET0131  & ~n22758 ;
  assign n22760 = ~n22745 & ~n22759 ;
  assign n22761 = n18604 & ~n20673 ;
  assign n22762 = n18666 & ~n22761 ;
  assign n22763 = \P4_reg2_reg[30]/NET0131  & ~n22762 ;
  assign n22770 = ~n22181 & ~n22645 ;
  assign n22771 = n20673 & ~n22770 ;
  assign n22765 = ~n16245 & n20673 ;
  assign n22764 = ~\P4_reg2_reg[30]/NET0131  & ~n20673 ;
  assign n22766 = n18486 & ~n22764 ;
  assign n22767 = ~n22765 & n22766 ;
  assign n22768 = \P4_reg2_reg[30]/NET0131  & ~n16425 ;
  assign n22769 = ~n20678 & n22768 ;
  assign n22772 = ~n22767 & ~n22769 ;
  assign n22773 = ~n21841 & n22772 ;
  assign n22774 = ~n22771 & n22773 ;
  assign n22775 = n18666 & ~n22774 ;
  assign n22776 = ~n22763 & ~n22775 ;
  assign n22777 = \P4_reg2_reg[7]/NET0131  & ~n18665 ;
  assign n22778 = \P4_reg2_reg[7]/NET0131  & n19073 ;
  assign n22780 = n20673 & ~n22079 ;
  assign n22781 = ~\P4_reg2_reg[7]/NET0131  & ~n20673 ;
  assign n22782 = n18483 & ~n22781 ;
  assign n22783 = ~n22780 & n22782 ;
  assign n22784 = n20673 & ~n22096 ;
  assign n22779 = \P4_reg2_reg[7]/NET0131  & ~n20682 ;
  assign n22785 = n16143 & n16426 ;
  assign n22786 = ~n22779 & ~n22785 ;
  assign n22787 = ~n22784 & n22786 ;
  assign n22788 = ~n22783 & n22787 ;
  assign n22789 = n19075 & ~n22788 ;
  assign n22790 = ~n22778 & ~n22789 ;
  assign n22791 = \P3_rd_reg/NET0131  & ~n22790 ;
  assign n22792 = ~n22777 & ~n22791 ;
  assign n22793 = \P2_P1_EAX_reg[28]/NET0131  & ~n21100 ;
  assign n22797 = ~n11537 & n22337 ;
  assign n22798 = \P2_P1_EAX_reg[28]/NET0131  & ~n22337 ;
  assign n22799 = ~n22797 & ~n22798 ;
  assign n22800 = n21068 & ~n22799 ;
  assign n22801 = n21022 & ~n21049 ;
  assign n22802 = ~n21072 & ~n22801 ;
  assign n22803 = \P2_P1_EAX_reg[28]/NET0131  & ~n22802 ;
  assign n22807 = ~\P2_P1_EAX_reg[28]/NET0131  & n21022 ;
  assign n22808 = n21049 & n22807 ;
  assign n22794 = ~n20919 & n20950 ;
  assign n22795 = ~n20951 & ~n22794 ;
  assign n22796 = n20728 & n22795 ;
  assign n22804 = n11375 & n22337 ;
  assign n22805 = ~n22798 & ~n22804 ;
  assign n22806 = n21062 & ~n22805 ;
  assign n22809 = ~n22796 & ~n22806 ;
  assign n22810 = ~n22808 & n22809 ;
  assign n22811 = ~n22803 & n22810 ;
  assign n22812 = ~n22800 & n22811 ;
  assign n22813 = n11623 & ~n22812 ;
  assign n22814 = ~n22793 & ~n22813 ;
  assign n22815 = \P1_P1_EAX_reg[28]/NET0131  & ~n15326 ;
  assign n22839 = n8223 & n15365 ;
  assign n22838 = ~\P1_P1_EAX_reg[28]/NET0131  & ~n15365 ;
  assign n22840 = n15383 & ~n22838 ;
  assign n22841 = ~n22839 & n22840 ;
  assign n22834 = n7985 & n15365 ;
  assign n22835 = n15334 & n22834 ;
  assign n22820 = \P1_P1_EAX_reg[24]/NET0131  & \P1_P1_EAX_reg[25]/NET0131  ;
  assign n22821 = \P1_P1_EAX_reg[17]/NET0131  & n15403 ;
  assign n22822 = \P1_P1_EAX_reg[18]/NET0131  & n22821 ;
  assign n22823 = \P1_P1_EAX_reg[19]/NET0131  & n22822 ;
  assign n22824 = \P1_P1_EAX_reg[20]/NET0131  & n22823 ;
  assign n22825 = n15404 & n22824 ;
  assign n22826 = \P1_P1_EAX_reg[23]/NET0131  & n22825 ;
  assign n22827 = n22820 & n22826 ;
  assign n22828 = n15412 & n22827 ;
  assign n22829 = n15377 & ~n22828 ;
  assign n22830 = n15372 & ~n15428 ;
  assign n22831 = n15387 & ~n22830 ;
  assign n22832 = ~n22829 & n22831 ;
  assign n22833 = \P1_P1_EAX_reg[28]/NET0131  & ~n22832 ;
  assign n22816 = ~n15620 & n15651 ;
  assign n22817 = ~n15652 & ~n22816 ;
  assign n22818 = n15372 & n15428 ;
  assign n22819 = n22817 & n22818 ;
  assign n22836 = ~\P1_P1_EAX_reg[28]/NET0131  & n15377 ;
  assign n22837 = n22828 & n22836 ;
  assign n22842 = ~n22819 & ~n22837 ;
  assign n22843 = ~n22833 & n22842 ;
  assign n22844 = ~n22835 & n22843 ;
  assign n22845 = ~n22841 & n22844 ;
  assign n22846 = n8355 & ~n22845 ;
  assign n22847 = ~n22815 & ~n22846 ;
  assign n22862 = n8270 & n15365 ;
  assign n22861 = ~\P1_P1_EAX_reg[30]/NET0131  & ~n15365 ;
  assign n22863 = n15383 & ~n22861 ;
  assign n22864 = ~n22862 & n22863 ;
  assign n22858 = ~n7925 & ~n7995 ;
  assign n22859 = n15365 & ~n22858 ;
  assign n22860 = n15334 & n22859 ;
  assign n22848 = \P1_P1_EAX_reg[28]/NET0131  & \P1_P1_EAX_reg[29]/NET0131  ;
  assign n22849 = n22828 & n22848 ;
  assign n22850 = n15377 & ~n22849 ;
  assign n22851 = n22831 & ~n22850 ;
  assign n22852 = \P1_P1_EAX_reg[30]/NET0131  & ~n22851 ;
  assign n22853 = ~\P1_P1_EAX_reg[30]/NET0131  & n15377 ;
  assign n22854 = n22849 & n22853 ;
  assign n22855 = ~n15684 & n15715 ;
  assign n22856 = ~n15716 & ~n22855 ;
  assign n22857 = n22818 & n22856 ;
  assign n22865 = ~n22854 & ~n22857 ;
  assign n22866 = ~n22852 & n22865 ;
  assign n22867 = ~n22860 & n22866 ;
  assign n22868 = ~n22864 & n22867 ;
  assign n22869 = n8355 & ~n22868 ;
  assign n22870 = \P1_P1_EAX_reg[30]/NET0131  & ~n15326 ;
  assign n22871 = ~n22869 & ~n22870 ;
  assign n22872 = ~n10029 & n18341 ;
  assign n22873 = \P1_P3_uWord_reg[14]/NET0131  & ~n22872 ;
  assign n22874 = ~n8741 & n21721 ;
  assign n22876 = ~\P1_P3_EAX_reg[12]/NET0131  & ~\P1_P3_EAX_reg[13]/NET0131  ;
  assign n22877 = ~\P1_P3_EAX_reg[14]/NET0131  & ~\P1_P3_EAX_reg[15]/NET0131  ;
  assign n22884 = n22876 & n22877 ;
  assign n22875 = ~\P1_P3_EAX_reg[10]/NET0131  & ~\P1_P3_EAX_reg[11]/NET0131  ;
  assign n22885 = n18804 & n22875 ;
  assign n22886 = n22884 & n22885 ;
  assign n22880 = ~\P1_P3_EAX_reg[6]/NET0131  & ~\P1_P3_EAX_reg[7]/NET0131  ;
  assign n22881 = ~\P1_P3_EAX_reg[8]/NET0131  & ~\P1_P3_EAX_reg[9]/NET0131  ;
  assign n22882 = n22880 & n22881 ;
  assign n22878 = ~\P1_P3_EAX_reg[2]/NET0131  & ~\P1_P3_EAX_reg[3]/NET0131  ;
  assign n22879 = ~\P1_P3_EAX_reg[4]/NET0131  & ~\P1_P3_EAX_reg[5]/NET0131  ;
  assign n22883 = n22878 & n22879 ;
  assign n22887 = n22882 & n22883 ;
  assign n22888 = n22886 & n22887 ;
  assign n22889 = \P1_P3_EAX_reg[31]/NET0131  & n21680 ;
  assign n22890 = n21495 & n22889 ;
  assign n22891 = ~n22888 & n22890 ;
  assign n22892 = ~\P1_P3_EAX_reg[30]/NET0131  & ~n22891 ;
  assign n22893 = \P1_P3_EAX_reg[30]/NET0131  & n22891 ;
  assign n22894 = ~n22892 & ~n22893 ;
  assign n22895 = n9079 & n22894 ;
  assign n22896 = ~n22874 & ~n22895 ;
  assign n22897 = ~n9075 & ~n22896 ;
  assign n22898 = n8741 & n9085 ;
  assign n22899 = ~n9236 & ~n16500 ;
  assign n22900 = ~n22898 & ~n22899 ;
  assign n22901 = \P1_P3_uWord_reg[14]/NET0131  & ~n22900 ;
  assign n22902 = ~n22897 & ~n22901 ;
  assign n22903 = n9241 & ~n22902 ;
  assign n22904 = ~n22873 & ~n22903 ;
  assign n22907 = ~\P4_reg3_reg[3]/NET0131  & n19073 ;
  assign n22914 = n16061 & ~n18452 ;
  assign n22915 = ~n18453 & ~n22914 ;
  assign n22916 = ~\P4_IR_reg[28]/NET0131  & ~n22915 ;
  assign n22917 = \P4_IR_reg[28]/NET0131  & n16083 ;
  assign n22918 = ~n22916 & ~n22917 ;
  assign n22919 = n19076 & ~n22918 ;
  assign n22910 = \P4_reg3_reg[3]/NET0131  & ~n19076 ;
  assign n22920 = n18483 & ~n22910 ;
  assign n22921 = ~n22919 & n22920 ;
  assign n22923 = n16287 & ~n18541 ;
  assign n22922 = ~n16287 & n18541 ;
  assign n22924 = n18490 & ~n22922 ;
  assign n22925 = ~n22923 & n22924 ;
  assign n22927 = ~n16115 & ~n16287 ;
  assign n22926 = n16115 & n16287 ;
  assign n22928 = n18607 & ~n22926 ;
  assign n22929 = ~n22927 & n22928 ;
  assign n22930 = ~n22925 & ~n22929 ;
  assign n22931 = n19076 & n22930 ;
  assign n22932 = ~n18672 & ~n22910 ;
  assign n22933 = ~n22931 & n22932 ;
  assign n22934 = ~n16074 & ~n18577 ;
  assign n22935 = ~n18578 & ~n22934 ;
  assign n22936 = n19076 & ~n22935 ;
  assign n22937 = n18604 & ~n22910 ;
  assign n22938 = ~n22936 & n22937 ;
  assign n22911 = n16074 & n19076 ;
  assign n22912 = n18486 & ~n22910 ;
  assign n22913 = ~n22911 & n22912 ;
  assign n22908 = ~n16074 & n16426 ;
  assign n22909 = ~\P4_reg3_reg[3]/NET0131  & n19104 ;
  assign n22939 = ~n22908 & ~n22909 ;
  assign n22940 = ~n22913 & n22939 ;
  assign n22941 = ~n22938 & n22940 ;
  assign n22942 = ~n22933 & n22941 ;
  assign n22943 = ~n22921 & n22942 ;
  assign n22944 = n19075 & ~n22943 ;
  assign n22945 = ~n22907 & ~n22944 ;
  assign n22946 = \P3_rd_reg/NET0131  & ~n22945 ;
  assign n22905 = ~\P4_reg3_reg[3]/NET0131  & n15744 ;
  assign n22906 = ~\P3_rd_reg/NET0131  & \P4_reg3_reg[3]/NET0131  ;
  assign n22947 = ~n22905 & ~n22906 ;
  assign n22948 = ~n22946 & n22947 ;
  assign n22949 = ~\P3_rd_reg/NET0131  & \P4_reg3_reg[6]/NET0131  ;
  assign n22950 = ~n16122 & n16426 ;
  assign n22951 = n16147 & ~n18455 ;
  assign n22952 = ~n18456 & ~n22951 ;
  assign n22953 = ~\P4_IR_reg[28]/NET0131  & ~n22952 ;
  assign n22954 = \P4_IR_reg[28]/NET0131  & n16048 ;
  assign n22955 = ~n22953 & ~n22954 ;
  assign n22956 = n18483 & n22955 ;
  assign n22967 = ~n16293 & n18547 ;
  assign n22966 = n16293 & ~n18547 ;
  assign n22968 = n18490 & ~n22966 ;
  assign n22969 = ~n22967 & n22968 ;
  assign n22958 = ~n16119 & ~n16133 ;
  assign n22960 = n16293 & ~n22958 ;
  assign n22959 = ~n16293 & n22958 ;
  assign n22961 = n18607 & ~n22959 ;
  assign n22962 = ~n22960 & n22961 ;
  assign n22957 = ~n16122 & n18486 ;
  assign n22963 = ~n16122 & ~n18580 ;
  assign n22964 = ~n18581 & n18604 ;
  assign n22965 = ~n22963 & n22964 ;
  assign n22970 = ~n22957 & ~n22965 ;
  assign n22971 = ~n22962 & n22970 ;
  assign n22972 = ~n22969 & n22971 ;
  assign n22973 = ~n22956 & n22972 ;
  assign n22974 = n19076 & ~n22973 ;
  assign n22975 = ~n22950 & ~n22974 ;
  assign n22976 = n19075 & ~n22975 ;
  assign n22977 = n16127 & ~n22003 ;
  assign n22978 = ~n22976 & ~n22977 ;
  assign n22979 = \P3_rd_reg/NET0131  & ~n22978 ;
  assign n22980 = ~n22949 & ~n22979 ;
  assign n22981 = ~\P3_rd_reg/NET0131  & \P4_reg3_reg[8]/NET0131  ;
  assign n22982 = ~n16026 & n16426 ;
  assign n22984 = n16021 & ~n18457 ;
  assign n22985 = ~n18458 & ~n22984 ;
  assign n22986 = ~\P4_IR_reg[28]/NET0131  & ~n22985 ;
  assign n22987 = \P4_IR_reg[28]/NET0131  & n16147 ;
  assign n22988 = n18483 & ~n22987 ;
  assign n22989 = ~n22986 & n22988 ;
  assign n22990 = ~n18518 & ~n18550 ;
  assign n22992 = ~n16292 & n22990 ;
  assign n22991 = n16292 & ~n22990 ;
  assign n22993 = n18490 & ~n22991 ;
  assign n22994 = ~n22992 & n22993 ;
  assign n22995 = ~n16151 & ~n16153 ;
  assign n22997 = ~n16292 & ~n22995 ;
  assign n22996 = n16292 & n22995 ;
  assign n22998 = n18607 & ~n22996 ;
  assign n22999 = ~n22997 & n22998 ;
  assign n22983 = ~n16026 & n18486 ;
  assign n23000 = ~n16026 & ~n18582 ;
  assign n23001 = ~n18583 & n18604 ;
  assign n23002 = ~n23000 & n23001 ;
  assign n23003 = ~n22983 & ~n23002 ;
  assign n23004 = ~n22999 & n23003 ;
  assign n23005 = ~n22994 & n23004 ;
  assign n23006 = ~n22989 & n23005 ;
  assign n23007 = n19076 & ~n23006 ;
  assign n23008 = ~n22982 & ~n23007 ;
  assign n23009 = n19075 & ~n23008 ;
  assign n23010 = n16031 & ~n22003 ;
  assign n23011 = ~n23009 & ~n23010 ;
  assign n23012 = \P3_rd_reg/NET0131  & ~n23011 ;
  assign n23013 = ~n22981 & ~n23012 ;
  assign n23014 = \P1_P3_State_reg[0]/NET0131  & hold_pad ;
  assign n23015 = \P1_P3_State_reg[1]/NET0131  & ~n22118 ;
  assign n23016 = ~n23014 & ~n23015 ;
  assign n23017 = \P1_P3_State_reg[2]/NET0131  & ~n23016 ;
  assign n23018 = \P1_P3_State_reg[0]/NET0131  & \P1_P3_State_reg[1]/NET0131  ;
  assign n23019 = ~\P1_P3_State_reg[2]/NET0131  & n23018 ;
  assign n23020 = ~\P1_P3_RequestPending_reg/NET0131  & ~hold_pad ;
  assign n23021 = n23019 & ~n23020 ;
  assign n23022 = n8741 & n23021 ;
  assign n23023 = ~n9094 & ~n23022 ;
  assign n23024 = ~na_pad & ~n23023 ;
  assign n23025 = ~\P1_P3_RequestPending_reg/NET0131  & ~\P1_P3_State_reg[1]/NET0131  ;
  assign n23026 = n23014 & n23025 ;
  assign n23027 = ~n23024 & ~n23026 ;
  assign n23028 = ~n23017 & n23027 ;
  assign n23029 = n15918 & ~n21999 ;
  assign n23031 = ~n16314 & ~n18700 ;
  assign n23032 = n16306 & ~n23031 ;
  assign n23033 = ~n16306 & n23031 ;
  assign n23034 = ~n23032 & ~n23033 ;
  assign n23035 = n18490 & ~n23034 ;
  assign n23037 = n16204 & n16306 ;
  assign n23036 = ~n16204 & ~n16306 ;
  assign n23038 = n18607 & ~n23036 ;
  assign n23039 = ~n23037 & n23038 ;
  assign n23040 = ~n23035 & ~n23039 ;
  assign n23041 = n15909 & ~n18467 ;
  assign n23042 = ~n22487 & ~n23041 ;
  assign n23043 = ~\P4_IR_reg[28]/NET0131  & ~n23042 ;
  assign n23044 = \P4_IR_reg[28]/NET0131  & n15936 ;
  assign n23045 = ~n23043 & ~n23044 ;
  assign n23046 = n18483 & n23045 ;
  assign n23047 = ~n15913 & ~n18592 ;
  assign n23048 = ~n18593 & ~n23047 ;
  assign n23049 = n18604 & n23048 ;
  assign n23050 = ~n23046 & ~n23049 ;
  assign n23051 = n23040 & n23050 ;
  assign n23052 = n19076 & ~n23051 ;
  assign n23030 = ~n15913 & ~n22190 ;
  assign n23053 = n15918 & ~n22002 ;
  assign n23054 = ~n23030 & ~n23053 ;
  assign n23055 = ~n23052 & n23054 ;
  assign n23056 = n19075 & ~n23055 ;
  assign n23057 = ~n23029 & ~n23056 ;
  assign n23058 = \P3_rd_reg/NET0131  & ~n23057 ;
  assign n23059 = ~\P3_rd_reg/NET0131  & \P4_reg3_reg[18]/NET0131  ;
  assign n23060 = ~n23058 & ~n23059 ;
  assign n23061 = n15828 & n19073 ;
  assign n23083 = n15820 & ~n18474 ;
  assign n23084 = ~n22149 & ~n23083 ;
  assign n23085 = ~\P4_IR_reg[28]/NET0131  & ~n23084 ;
  assign n23086 = \P4_IR_reg[28]/NET0131  & n15844 ;
  assign n23087 = ~n23085 & ~n23086 ;
  assign n23088 = n19076 & ~n23087 ;
  assign n23082 = ~n15828 & ~n19076 ;
  assign n23089 = n18483 & ~n23082 ;
  assign n23090 = ~n23088 & n23089 ;
  assign n23063 = n15823 & ~n18599 ;
  assign n23064 = ~n18600 & ~n23063 ;
  assign n23065 = n18604 & n23064 ;
  assign n23067 = ~n15845 & ~n18637 ;
  assign n23069 = ~n16262 & n23067 ;
  assign n23068 = n16262 & ~n23067 ;
  assign n23070 = n18607 & ~n23068 ;
  assign n23071 = ~n23069 & n23070 ;
  assign n23066 = n15823 & n18486 ;
  assign n23072 = ~n16277 & ~n21814 ;
  assign n23074 = ~n16262 & ~n23072 ;
  assign n23073 = n16262 & n23072 ;
  assign n23075 = n18490 & ~n23073 ;
  assign n23076 = ~n23074 & n23075 ;
  assign n23077 = ~n23066 & ~n23076 ;
  assign n23078 = ~n23071 & n23077 ;
  assign n23079 = ~n23065 & n23078 ;
  assign n23080 = n19076 & ~n23079 ;
  assign n23062 = n15823 & n16426 ;
  assign n23081 = n15828 & ~n19177 ;
  assign n23091 = ~n23062 & ~n23081 ;
  assign n23092 = ~n23080 & n23091 ;
  assign n23093 = ~n23090 & n23092 ;
  assign n23094 = n19075 & ~n23093 ;
  assign n23095 = ~n23061 & ~n23094 ;
  assign n23096 = \P3_rd_reg/NET0131  & ~n23095 ;
  assign n23097 = n15744 & n15828 ;
  assign n23098 = ~\P3_rd_reg/NET0131  & \P4_reg3_reg[25]/NET0131  ;
  assign n23099 = ~n23097 & ~n23098 ;
  assign n23100 = ~n23096 & n23099 ;
  assign n23101 = ~\P3_rd_reg/NET0131  & \P4_reg3_reg[22]/NET0131  ;
  assign n23102 = n15858 & n16426 ;
  assign n23103 = n19076 & ~n22599 ;
  assign n23104 = ~n23102 & ~n23103 ;
  assign n23105 = n19075 & ~n23104 ;
  assign n23106 = n15868 & ~n22003 ;
  assign n23107 = ~n23105 & ~n23106 ;
  assign n23108 = \P3_rd_reg/NET0131  & ~n23107 ;
  assign n23109 = ~n23101 & ~n23108 ;
  assign n23110 = \P4_reg2_reg[10]/NET0131  & ~n18665 ;
  assign n23111 = \P4_reg2_reg[10]/NET0131  & n19073 ;
  assign n23113 = \P4_reg2_reg[10]/NET0131  & ~n20673 ;
  assign n23114 = n20673 & n22439 ;
  assign n23115 = ~n23113 & ~n23114 ;
  assign n23116 = n18483 & ~n23115 ;
  assign n23117 = n20673 & ~n22433 ;
  assign n23118 = \P4_reg2_reg[10]/NET0131  & n22261 ;
  assign n23112 = n16002 & n16426 ;
  assign n23119 = ~n15997 & n20673 ;
  assign n23120 = ~n23113 & ~n23119 ;
  assign n23121 = n18486 & ~n23120 ;
  assign n23122 = ~n23112 & ~n23121 ;
  assign n23123 = ~n23118 & n23122 ;
  assign n23124 = ~n23117 & n23123 ;
  assign n23125 = ~n23116 & n23124 ;
  assign n23126 = n19075 & ~n23125 ;
  assign n23127 = ~n23111 & ~n23126 ;
  assign n23128 = \P3_rd_reg/NET0131  & ~n23127 ;
  assign n23129 = ~n23110 & ~n23128 ;
  assign n23131 = \P4_reg0_reg[14]/NET0131  & ~n20661 ;
  assign n23132 = n20665 & n22456 ;
  assign n23133 = ~n23131 & ~n23132 ;
  assign n23134 = n18483 & ~n23133 ;
  assign n23130 = n20665 & ~n22474 ;
  assign n23135 = \P4_reg0_reg[14]/NET0131  & ~n21854 ;
  assign n23136 = ~n23130 & ~n23135 ;
  assign n23137 = ~n23134 & n23136 ;
  assign n23138 = \P4_reg0_reg[22]/NET0131  & ~n21855 ;
  assign n23139 = n20665 & ~n22599 ;
  assign n23140 = ~n23138 & ~n23139 ;
  assign n23141 = \P4_reg1_reg[14]/NET0131  & ~n18679 ;
  assign n23142 = n18667 & ~n22475 ;
  assign n23143 = ~n23141 & ~n23142 ;
  assign n23145 = \P4_reg1_reg[20]/NET0131  & ~n18664 ;
  assign n23146 = n18667 & ~n22492 ;
  assign n23147 = ~n23145 & ~n23146 ;
  assign n23148 = n18483 & ~n23147 ;
  assign n23144 = \P4_reg1_reg[20]/NET0131  & ~n21863 ;
  assign n23149 = n18667 & ~n22508 ;
  assign n23150 = ~n23144 & ~n23149 ;
  assign n23151 = ~n23148 & n23150 ;
  assign n23152 = n16184 & n16426 ;
  assign n23153 = n20673 & ~n22475 ;
  assign n23154 = ~n23152 & ~n23153 ;
  assign n23155 = n18666 & ~n23154 ;
  assign n23156 = \P4_reg2_reg[14]/NET0131  & ~n22574 ;
  assign n23157 = ~n23155 & ~n23156 ;
  assign n23158 = \P2_P1_EAX_reg[29]/NET0131  & ~n21100 ;
  assign n23171 = n11553 & n22337 ;
  assign n23170 = ~\P2_P1_EAX_reg[29]/NET0131  & ~n22337 ;
  assign n23172 = n21068 & ~n23170 ;
  assign n23173 = ~n23171 & n23172 ;
  assign n23159 = ~\P2_P1_EAX_reg[29]/NET0131  & ~n21050 ;
  assign n23160 = n22342 & ~n23159 ;
  assign n23161 = n21062 & ~n22337 ;
  assign n23162 = ~n21072 & ~n23161 ;
  assign n23163 = \P2_P1_EAX_reg[29]/NET0131  & ~n23162 ;
  assign n23164 = ~n20951 & n20982 ;
  assign n23165 = ~n20983 & ~n23164 ;
  assign n23166 = n20728 & n23165 ;
  assign n23167 = n21062 & ~n21073 ;
  assign n23168 = n11384 & n23167 ;
  assign n23169 = ~n21081 & n23168 ;
  assign n23174 = ~n23166 & ~n23169 ;
  assign n23175 = ~n23163 & n23174 ;
  assign n23176 = ~n23160 & n23175 ;
  assign n23177 = ~n23173 & n23176 ;
  assign n23178 = n11623 & ~n23177 ;
  assign n23179 = ~n23158 & ~n23178 ;
  assign n23183 = ~n8248 & n15365 ;
  assign n23184 = \P1_P1_EAX_reg[29]/NET0131  & ~n15365 ;
  assign n23185 = ~n23183 & ~n23184 ;
  assign n23186 = n15383 & ~n23185 ;
  assign n23187 = ~n8007 & n15365 ;
  assign n23188 = ~n23184 & ~n23187 ;
  assign n23189 = n15334 & ~n23188 ;
  assign n23190 = ~n15386 & ~n22830 ;
  assign n23191 = n15377 & ~n15415 ;
  assign n23192 = n23190 & ~n23191 ;
  assign n23193 = \P1_P1_EAX_reg[29]/NET0131  & ~n23192 ;
  assign n23180 = ~n15652 & n15683 ;
  assign n23181 = ~n15684 & ~n23180 ;
  assign n23182 = n22818 & n23181 ;
  assign n23194 = n15377 & n15411 ;
  assign n23195 = ~\P1_P1_EAX_reg[29]/NET0131  & n15414 ;
  assign n23196 = n23194 & n23195 ;
  assign n23197 = ~n23182 & ~n23196 ;
  assign n23198 = ~n23193 & n23197 ;
  assign n23199 = ~n23189 & n23198 ;
  assign n23200 = ~n23186 & n23199 ;
  assign n23201 = n8355 & ~n23200 ;
  assign n23202 = \P1_P1_EAX_reg[29]/NET0131  & ~n15326 ;
  assign n23203 = ~n23201 & ~n23202 ;
  assign n23204 = ~\P3_rd_reg/NET0131  & \P4_reg3_reg[13]/NET0131  ;
  assign n23205 = ~n15954 & n16426 ;
  assign n23206 = n16188 & ~n18462 ;
  assign n23207 = ~n19077 & ~n23206 ;
  assign n23208 = ~\P4_IR_reg[28]/NET0131  & ~n23207 ;
  assign n23209 = \P4_IR_reg[28]/NET0131  & n15976 ;
  assign n23210 = ~n23208 & ~n23209 ;
  assign n23211 = n18483 & n23210 ;
  assign n23221 = ~n16265 & n21801 ;
  assign n23220 = n16265 & ~n21801 ;
  assign n23222 = n18490 & ~n23220 ;
  assign n23223 = ~n23221 & n23222 ;
  assign n23217 = n16265 & n18618 ;
  assign n23216 = ~n16265 & ~n18618 ;
  assign n23218 = n18607 & ~n23216 ;
  assign n23219 = ~n23217 & n23218 ;
  assign n23212 = ~n15954 & n18486 ;
  assign n23213 = ~n15954 & ~n18587 ;
  assign n23214 = ~n18588 & n18604 ;
  assign n23215 = ~n23213 & n23214 ;
  assign n23224 = ~n23212 & ~n23215 ;
  assign n23225 = ~n23219 & n23224 ;
  assign n23226 = ~n23223 & n23225 ;
  assign n23227 = ~n23211 & n23226 ;
  assign n23228 = n19076 & ~n23227 ;
  assign n23229 = ~n23205 & ~n23228 ;
  assign n23230 = n19075 & ~n23229 ;
  assign n23231 = n15959 & ~n22003 ;
  assign n23232 = ~n23230 & ~n23231 ;
  assign n23233 = \P3_rd_reg/NET0131  & ~n23232 ;
  assign n23234 = ~n23204 & ~n23233 ;
  assign n23236 = n15932 & n19073 ;
  assign n23238 = n16315 & ~n21806 ;
  assign n23239 = ~n16315 & n21806 ;
  assign n23240 = ~n23238 & ~n23239 ;
  assign n23241 = n18490 & n23240 ;
  assign n23247 = n16315 & n18627 ;
  assign n23246 = ~n16315 & ~n18627 ;
  assign n23248 = n18607 & ~n23246 ;
  assign n23249 = ~n23247 & n23248 ;
  assign n23242 = ~n15927 & n18486 ;
  assign n23243 = ~n15927 & ~n18591 ;
  assign n23244 = ~n18592 & n18604 ;
  assign n23245 = ~n23243 & n23244 ;
  assign n23250 = ~n23242 & ~n23245 ;
  assign n23251 = ~n23249 & n23250 ;
  assign n23252 = ~n23241 & n23251 ;
  assign n23253 = \P4_IR_reg[28]/NET0131  & ~n15949 ;
  assign n23254 = n15922 & ~n22043 ;
  assign n23255 = ~\P4_IR_reg[28]/NET0131  & ~n18467 ;
  assign n23256 = ~n23254 & n23255 ;
  assign n23257 = ~n23253 & ~n23256 ;
  assign n23258 = n18483 & ~n23257 ;
  assign n23259 = n23252 & ~n23258 ;
  assign n23260 = n19076 & ~n23259 ;
  assign n23237 = ~n15927 & n16426 ;
  assign n23261 = n15932 & ~n22160 ;
  assign n23262 = ~n23237 & ~n23261 ;
  assign n23263 = ~n23260 & n23262 ;
  assign n23264 = n19075 & ~n23263 ;
  assign n23265 = ~n23236 & ~n23264 ;
  assign n23266 = \P3_rd_reg/NET0131  & ~n23265 ;
  assign n23235 = n15744 & n15932 ;
  assign n23267 = ~\P3_rd_reg/NET0131  & \P4_reg3_reg[17]/NET0131  ;
  assign n23268 = ~n23235 & ~n23267 ;
  assign n23269 = ~n23266 & n23268 ;
  assign n23270 = ~\P4_reg3_reg[1]/NET0131  & ~n19076 ;
  assign n23271 = n16083 & ~n18450 ;
  assign n23272 = ~n18451 & ~n23271 ;
  assign n23273 = ~\P4_IR_reg[28]/NET0131  & ~n23272 ;
  assign n23274 = \P4_IR_reg[28]/NET0131  & n16110 ;
  assign n23275 = ~n23273 & ~n23274 ;
  assign n23276 = n19076 & ~n23275 ;
  assign n23277 = n18483 & ~n23276 ;
  assign n23278 = ~n16098 & n18486 ;
  assign n23279 = ~n16098 & ~n16103 ;
  assign n23280 = ~n18576 & ~n23279 ;
  assign n23281 = n18604 & n23280 ;
  assign n23282 = ~n16099 & ~n16100 ;
  assign n23284 = ~n16111 & n23282 ;
  assign n23283 = n16111 & ~n23282 ;
  assign n23285 = n18607 & ~n23283 ;
  assign n23286 = ~n23284 & n23285 ;
  assign n23288 = n18537 & ~n23282 ;
  assign n23287 = ~n18537 & n23282 ;
  assign n23289 = n18490 & ~n23287 ;
  assign n23290 = ~n23288 & n23289 ;
  assign n23291 = ~n23286 & ~n23290 ;
  assign n23292 = ~n23281 & n23291 ;
  assign n23293 = ~n23278 & n23292 ;
  assign n23294 = n19076 & ~n23293 ;
  assign n23295 = n18666 & ~n23294 ;
  assign n23296 = ~n23277 & n23295 ;
  assign n23297 = ~n23270 & ~n23296 ;
  assign n23298 = ~n16098 & n16426 ;
  assign n23299 = \P4_reg3_reg[1]/NET0131  & ~n19177 ;
  assign n23300 = ~n23298 & ~n23299 ;
  assign n23301 = ~n23297 & n23300 ;
  assign n23302 = ~\P4_reg3_reg[1]/NET0131  & ~n18666 ;
  assign n23303 = ~n23301 & ~n23302 ;
  assign n23304 = ~n16086 & n16426 ;
  assign n23305 = n16071 & ~n18451 ;
  assign n23306 = ~n18452 & ~n23305 ;
  assign n23307 = ~\P4_IR_reg[28]/NET0131  & ~n23306 ;
  assign n23308 = \P4_IR_reg[28]/NET0131  & n16095 ;
  assign n23309 = ~n23307 & ~n23308 ;
  assign n23310 = n18483 & n23309 ;
  assign n23320 = n16113 & ~n16282 ;
  assign n23319 = ~n16113 & n16282 ;
  assign n23321 = n18607 & ~n23319 ;
  assign n23322 = ~n23320 & n23321 ;
  assign n23316 = ~n16282 & n18539 ;
  assign n23315 = n16282 & ~n18539 ;
  assign n23317 = n18490 & ~n23315 ;
  assign n23318 = ~n23316 & n23317 ;
  assign n23311 = ~n16086 & n18486 ;
  assign n23312 = ~n16086 & ~n18576 ;
  assign n23313 = ~n18577 & n18604 ;
  assign n23314 = ~n23312 & n23313 ;
  assign n23323 = ~n23311 & ~n23314 ;
  assign n23324 = ~n23318 & n23323 ;
  assign n23325 = ~n23322 & n23324 ;
  assign n23326 = ~n23310 & n23325 ;
  assign n23327 = n19076 & ~n23326 ;
  assign n23328 = ~n23304 & ~n23327 ;
  assign n23329 = n18666 & ~n23328 ;
  assign n23330 = \P3_rd_reg/NET0131  & n22003 ;
  assign n23331 = \P4_reg3_reg[2]/NET0131  & ~n23330 ;
  assign n23332 = ~n23329 & ~n23331 ;
  assign n23333 = ~\P3_rd_reg/NET0131  & \P4_reg3_reg[5]/NET0131  ;
  assign n23334 = ~n16039 & n16426 ;
  assign n23335 = n16131 & ~n18454 ;
  assign n23336 = ~n18455 & ~n23335 ;
  assign n23337 = ~\P4_IR_reg[28]/NET0131  & ~n23336 ;
  assign n23338 = \P4_IR_reg[28]/NET0131  & n16061 ;
  assign n23339 = ~n23337 & ~n23338 ;
  assign n23340 = n18483 & n23339 ;
  assign n23351 = n16296 & n18545 ;
  assign n23350 = ~n16296 & ~n18545 ;
  assign n23352 = n18490 & ~n23350 ;
  assign n23353 = ~n23351 & n23352 ;
  assign n23342 = ~n16062 & ~n16118 ;
  assign n23344 = n16296 & ~n23342 ;
  assign n23343 = ~n16296 & n23342 ;
  assign n23345 = n18607 & ~n23343 ;
  assign n23346 = ~n23344 & n23345 ;
  assign n23341 = ~n16039 & n18486 ;
  assign n23347 = ~n16039 & ~n18579 ;
  assign n23348 = ~n18580 & n18604 ;
  assign n23349 = ~n23347 & n23348 ;
  assign n23354 = ~n23341 & ~n23349 ;
  assign n23355 = ~n23346 & n23354 ;
  assign n23356 = ~n23353 & n23355 ;
  assign n23357 = ~n23340 & n23356 ;
  assign n23358 = n19076 & ~n23357 ;
  assign n23359 = ~n23334 & ~n23358 ;
  assign n23360 = n19075 & ~n23359 ;
  assign n23361 = n16044 & ~n22003 ;
  assign n23362 = ~n23360 & ~n23361 ;
  assign n23363 = \P3_rd_reg/NET0131  & ~n23362 ;
  assign n23364 = ~n23333 & ~n23363 ;
  assign n23366 = n16017 & n19073 ;
  assign n23368 = ~n16012 & ~n18583 ;
  assign n23369 = ~n18584 & ~n23368 ;
  assign n23370 = n18604 & n23369 ;
  assign n23377 = n16272 & n18685 ;
  assign n23376 = ~n16272 & ~n18685 ;
  assign n23378 = n18490 & ~n23376 ;
  assign n23379 = ~n23377 & n23378 ;
  assign n23371 = ~n16012 & n18486 ;
  assign n23373 = ~n16156 & n16272 ;
  assign n23372 = n16156 & ~n16272 ;
  assign n23374 = n18607 & ~n23372 ;
  assign n23375 = ~n23373 & n23374 ;
  assign n23380 = ~n23371 & ~n23375 ;
  assign n23381 = ~n23379 & n23380 ;
  assign n23382 = ~n23370 & n23381 ;
  assign n23383 = n16006 & ~n18458 ;
  assign n23384 = ~n18459 & ~n23383 ;
  assign n23385 = ~\P4_IR_reg[28]/NET0131  & ~n23384 ;
  assign n23386 = \P4_IR_reg[28]/NET0131  & n16035 ;
  assign n23387 = ~n23385 & ~n23386 ;
  assign n23388 = n18483 & n23387 ;
  assign n23389 = n23382 & ~n23388 ;
  assign n23390 = n19076 & ~n23389 ;
  assign n23367 = ~n16012 & n16426 ;
  assign n23391 = n16017 & ~n22160 ;
  assign n23392 = ~n23367 & ~n23391 ;
  assign n23393 = ~n23390 & n23392 ;
  assign n23394 = n19075 & ~n23393 ;
  assign n23395 = ~n23366 & ~n23394 ;
  assign n23396 = \P3_rd_reg/NET0131  & ~n23395 ;
  assign n23365 = n15744 & n16017 ;
  assign n23397 = ~\P3_rd_reg/NET0131  & \P4_reg3_reg[9]/NET0131  ;
  assign n23398 = ~n23365 & ~n23397 ;
  assign n23399 = ~n23396 & n23398 ;
  assign n23401 = \P4_reg0_reg[10]/NET0131  & ~n20661 ;
  assign n23402 = n20665 & n22439 ;
  assign n23403 = ~n23401 & ~n23402 ;
  assign n23404 = n18483 & ~n23403 ;
  assign n23400 = n20665 & ~n22434 ;
  assign n23405 = \P4_reg0_reg[10]/NET0131  & ~n21854 ;
  assign n23406 = ~n23400 & ~n23405 ;
  assign n23407 = ~n23404 & n23406 ;
  assign n23408 = \P4_reg0_reg[18]/NET0131  & ~n18665 ;
  assign n23409 = \P4_reg0_reg[18]/NET0131  & n19073 ;
  assign n23410 = \P4_reg0_reg[18]/NET0131  & ~n20661 ;
  assign n23411 = n20661 & n23045 ;
  assign n23412 = ~n23410 & ~n23411 ;
  assign n23413 = n18483 & ~n23412 ;
  assign n23418 = ~n15913 & n18486 ;
  assign n23419 = n23040 & ~n23418 ;
  assign n23420 = n20661 & ~n23419 ;
  assign n23414 = ~n18676 & ~n21852 ;
  assign n23415 = n18486 & ~n20661 ;
  assign n23416 = n23414 & ~n23415 ;
  assign n23417 = \P4_reg0_reg[18]/NET0131  & ~n23416 ;
  assign n23421 = n20661 & n23048 ;
  assign n23422 = ~n23410 & ~n23421 ;
  assign n23423 = n18604 & ~n23422 ;
  assign n23424 = ~n23417 & ~n23423 ;
  assign n23425 = ~n23420 & n23424 ;
  assign n23426 = ~n23413 & n23425 ;
  assign n23427 = n19075 & ~n23426 ;
  assign n23428 = ~n23409 & ~n23427 ;
  assign n23429 = \P3_rd_reg/NET0131  & ~n23428 ;
  assign n23430 = ~n23408 & ~n23429 ;
  assign n23431 = \P4_reg0_reg[25]/NET0131  & ~n21855 ;
  assign n23432 = n18483 & n23087 ;
  assign n23433 = n23079 & ~n23432 ;
  assign n23434 = n20665 & ~n23433 ;
  assign n23435 = ~n23431 & ~n23434 ;
  assign n23436 = n18483 & n22918 ;
  assign n23437 = ~n16074 & n18486 ;
  assign n23438 = n18604 & n22935 ;
  assign n23439 = ~n23437 & ~n23438 ;
  assign n23440 = n22930 & n23439 ;
  assign n23441 = ~n23436 & n23440 ;
  assign n23442 = n20665 & ~n23441 ;
  assign n23443 = \P4_reg0_reg[3]/NET0131  & ~n21855 ;
  assign n23444 = ~n23442 & ~n23443 ;
  assign n23445 = n20665 & ~n22973 ;
  assign n23446 = \P4_reg0_reg[6]/NET0131  & ~n21855 ;
  assign n23447 = ~n23445 & ~n23446 ;
  assign n23448 = n20665 & ~n23006 ;
  assign n23449 = \P4_reg0_reg[8]/NET0131  & ~n21855 ;
  assign n23450 = ~n23448 & ~n23449 ;
  assign n23452 = \P4_reg1_reg[10]/NET0131  & ~n18664 ;
  assign n23453 = n18667 & n22439 ;
  assign n23454 = ~n23452 & ~n23453 ;
  assign n23455 = n18483 & ~n23454 ;
  assign n23451 = n18667 & ~n22434 ;
  assign n23456 = \P4_reg1_reg[10]/NET0131  & ~n21863 ;
  assign n23457 = ~n23451 & ~n23456 ;
  assign n23458 = ~n23455 & n23457 ;
  assign n23459 = ~\P4_reg1_reg[18]/NET0131  & ~n18667 ;
  assign n23461 = ~n18490 & n18664 ;
  assign n23462 = ~n18672 & ~n23461 ;
  assign n23463 = ~n23034 & n23462 ;
  assign n23460 = \P4_reg1_reg[18]/NET0131  & ~n22685 ;
  assign n23464 = ~n23418 & ~n23460 ;
  assign n23465 = ~n23463 & n23464 ;
  assign n23466 = n23050 & n23465 ;
  assign n23467 = ~n18486 & n18675 ;
  assign n23468 = ~n18664 & n23467 ;
  assign n23469 = ~n23462 & n23468 ;
  assign n23470 = ~n23466 & ~n23469 ;
  assign n23471 = n18666 & ~n23039 ;
  assign n23472 = ~n23470 & n23471 ;
  assign n23473 = ~n23459 & ~n23472 ;
  assign n23474 = n18667 & ~n23433 ;
  assign n23475 = \P4_reg1_reg[25]/NET0131  & ~n18679 ;
  assign n23476 = ~n23474 & ~n23475 ;
  assign n23477 = \P4_reg1_reg[3]/NET0131  & ~n18679 ;
  assign n23478 = n18667 & ~n23441 ;
  assign n23479 = ~n23477 & ~n23478 ;
  assign n23480 = \P4_reg1_reg[6]/NET0131  & ~n18679 ;
  assign n23481 = n18667 & ~n22973 ;
  assign n23482 = ~n23480 & ~n23481 ;
  assign n23483 = \P4_reg1_reg[8]/NET0131  & ~n18679 ;
  assign n23484 = n18667 & ~n23006 ;
  assign n23485 = ~n23483 & ~n23484 ;
  assign n23486 = \P4_reg2_reg[18]/NET0131  & ~n18665 ;
  assign n23487 = \P4_reg2_reg[18]/NET0131  & n19073 ;
  assign n23491 = \P4_reg2_reg[18]/NET0131  & ~n20673 ;
  assign n23492 = n20673 & n23045 ;
  assign n23493 = ~n23491 & ~n23492 ;
  assign n23494 = n18483 & ~n23493 ;
  assign n23495 = n20673 & ~n23419 ;
  assign n23496 = n20673 & n23048 ;
  assign n23497 = ~n23491 & ~n23496 ;
  assign n23498 = n18604 & ~n23497 ;
  assign n23488 = ~n18672 & ~n20673 ;
  assign n23489 = ~n22321 & ~n23488 ;
  assign n23490 = \P4_reg2_reg[18]/NET0131  & ~n23489 ;
  assign n23499 = n15918 & n16426 ;
  assign n23500 = ~n23490 & ~n23499 ;
  assign n23501 = ~n23498 & n23500 ;
  assign n23502 = ~n23495 & n23501 ;
  assign n23503 = ~n23494 & n23502 ;
  assign n23504 = n19075 & ~n23503 ;
  assign n23505 = ~n23487 & ~n23504 ;
  assign n23506 = \P3_rd_reg/NET0131  & ~n23505 ;
  assign n23507 = ~n23486 & ~n23506 ;
  assign n23508 = \P4_reg2_reg[25]/NET0131  & ~n18665 ;
  assign n23510 = \P4_reg2_reg[25]/NET0131  & ~n20673 ;
  assign n23511 = n20673 & n23087 ;
  assign n23512 = ~n23510 & ~n23511 ;
  assign n23513 = n18483 & ~n23512 ;
  assign n23514 = n20673 & ~n23078 ;
  assign n23515 = n20673 & n23064 ;
  assign n23516 = ~n23510 & ~n23515 ;
  assign n23517 = n18604 & ~n23516 ;
  assign n23509 = \P4_reg2_reg[25]/NET0131  & ~n23489 ;
  assign n23518 = n15828 & n16426 ;
  assign n23519 = ~n23509 & ~n23518 ;
  assign n23520 = ~n23517 & n23519 ;
  assign n23521 = ~n23514 & n23520 ;
  assign n23522 = ~n23513 & n23521 ;
  assign n23523 = n19075 & ~n23522 ;
  assign n23524 = \P4_reg2_reg[25]/NET0131  & n19073 ;
  assign n23525 = ~n23523 & ~n23524 ;
  assign n23526 = \P3_rd_reg/NET0131  & ~n23525 ;
  assign n23527 = ~n23508 & ~n23526 ;
  assign n23528 = ~\P4_reg2_reg[3]/NET0131  & ~n20673 ;
  assign n23529 = n20673 & ~n22918 ;
  assign n23530 = n18483 & ~n23529 ;
  assign n23531 = n20673 & ~n23440 ;
  assign n23532 = n18666 & ~n23531 ;
  assign n23533 = ~n23530 & n23532 ;
  assign n23534 = ~n23528 & ~n23533 ;
  assign n23535 = ~\P4_reg3_reg[3]/NET0131  & n16426 ;
  assign n23536 = ~n23534 & ~n23535 ;
  assign n23537 = n18666 & ~n23536 ;
  assign n23538 = ~\P4_reg2_reg[3]/NET0131  & ~n23537 ;
  assign n23539 = n20682 & n23536 ;
  assign n23540 = ~n23538 & ~n23539 ;
  assign n23541 = \P4_reg2_reg[6]/NET0131  & ~n18665 ;
  assign n23542 = \P4_reg2_reg[6]/NET0131  & n19073 ;
  assign n23544 = n20673 & ~n22955 ;
  assign n23545 = ~\P4_reg2_reg[6]/NET0131  & ~n20673 ;
  assign n23546 = n18483 & ~n23545 ;
  assign n23547 = ~n23544 & n23546 ;
  assign n23548 = n20673 & ~n22972 ;
  assign n23543 = \P4_reg2_reg[6]/NET0131  & ~n20682 ;
  assign n23549 = n16127 & n16426 ;
  assign n23550 = ~n23543 & ~n23549 ;
  assign n23551 = ~n23548 & n23550 ;
  assign n23552 = ~n23547 & n23551 ;
  assign n23553 = n19075 & ~n23552 ;
  assign n23554 = ~n23542 & ~n23553 ;
  assign n23555 = \P3_rd_reg/NET0131  & ~n23554 ;
  assign n23556 = ~n23541 & ~n23555 ;
  assign n23557 = \P4_reg2_reg[8]/NET0131  & ~n22574 ;
  assign n23558 = n16031 & n16426 ;
  assign n23559 = n20673 & ~n23006 ;
  assign n23560 = ~n23558 & ~n23559 ;
  assign n23561 = n18666 & ~n23560 ;
  assign n23562 = ~n23557 & ~n23561 ;
  assign n23563 = \P1_P1_EAX_reg[26]/NET0131  & ~n15326 ;
  assign n23565 = n8206 & n15365 ;
  assign n23564 = ~\P1_P1_EAX_reg[26]/NET0131  & ~n15365 ;
  assign n23566 = n15383 & ~n23564 ;
  assign n23567 = ~n23565 & n23566 ;
  assign n23580 = ~n7966 & n15365 ;
  assign n23581 = n15334 & n23580 ;
  assign n23571 = n15377 & ~n22827 ;
  assign n23572 = n15387 & ~n23571 ;
  assign n23573 = \P1_P1_EAX_reg[26]/NET0131  & ~n23572 ;
  assign n23568 = n15377 & n22826 ;
  assign n23569 = ~\P1_P1_EAX_reg[26]/NET0131  & n22820 ;
  assign n23570 = n23568 & n23569 ;
  assign n23574 = \P1_P1_EAX_reg[26]/NET0131  & ~n15428 ;
  assign n23575 = ~n15556 & n15587 ;
  assign n23576 = n15428 & ~n15588 ;
  assign n23577 = ~n23575 & n23576 ;
  assign n23578 = ~n23574 & ~n23577 ;
  assign n23579 = n15372 & ~n23578 ;
  assign n23582 = ~n23570 & ~n23579 ;
  assign n23583 = ~n23573 & n23582 ;
  assign n23584 = ~n23581 & n23583 ;
  assign n23585 = ~n23567 & n23584 ;
  assign n23586 = n8355 & ~n23585 ;
  assign n23587 = ~n23563 & ~n23586 ;
  assign n23588 = ~\P3_rd_reg/NET0131  & \P4_reg3_reg[4]/NET0131  ;
  assign n23589 = ~n16052 & n16426 ;
  assign n23590 = n16048 & ~n18453 ;
  assign n23591 = ~n18454 & ~n23590 ;
  assign n23592 = ~\P4_IR_reg[28]/NET0131  & ~n23591 ;
  assign n23593 = \P4_IR_reg[28]/NET0131  & n16071 ;
  assign n23594 = ~n23592 & ~n23593 ;
  assign n23595 = n18483 & n23594 ;
  assign n23605 = n16117 & ~n16266 ;
  assign n23604 = ~n16117 & n16266 ;
  assign n23606 = n18607 & ~n23604 ;
  assign n23607 = ~n23605 & n23606 ;
  assign n23601 = ~n16266 & n18543 ;
  assign n23600 = n16266 & ~n18543 ;
  assign n23602 = n18490 & ~n23600 ;
  assign n23603 = ~n23601 & n23602 ;
  assign n23596 = ~n16052 & n18486 ;
  assign n23597 = ~n16052 & ~n18578 ;
  assign n23598 = ~n18579 & n18604 ;
  assign n23599 = ~n23597 & n23598 ;
  assign n23608 = ~n23596 & ~n23599 ;
  assign n23609 = ~n23603 & n23608 ;
  assign n23610 = ~n23607 & n23609 ;
  assign n23611 = ~n23595 & n23610 ;
  assign n23612 = n19076 & ~n23611 ;
  assign n23613 = ~n23589 & ~n23612 ;
  assign n23614 = n19075 & ~n23613 ;
  assign n23615 = n16057 & ~n22003 ;
  assign n23616 = ~n23614 & ~n23615 ;
  assign n23617 = \P3_rd_reg/NET0131  & ~n23616 ;
  assign n23618 = ~n23588 & ~n23617 ;
  assign n23620 = n15880 & n19073 ;
  assign n23640 = n15872 & ~n18470 ;
  assign n23641 = ~n22577 & ~n23640 ;
  assign n23642 = ~\P4_IR_reg[28]/NET0131  & ~n23641 ;
  assign n23643 = \P4_IR_reg[28]/NET0131  & n15895 ;
  assign n23644 = ~n23642 & ~n23643 ;
  assign n23645 = n19076 & ~n23644 ;
  assign n23639 = ~n15880 & ~n19076 ;
  assign n23646 = n18483 & ~n23639 ;
  assign n23647 = ~n23645 & n23646 ;
  assign n23622 = n15875 & ~n18595 ;
  assign n23623 = ~n18596 & ~n23622 ;
  assign n23624 = n18604 & n23623 ;
  assign n23625 = n15875 & n18486 ;
  assign n23627 = n16275 & n18633 ;
  assign n23626 = ~n16275 & ~n18633 ;
  assign n23628 = n18607 & ~n23626 ;
  assign n23629 = ~n23627 & n23628 ;
  assign n23631 = ~n16275 & n21810 ;
  assign n23630 = n16275 & ~n21810 ;
  assign n23632 = n18490 & ~n23630 ;
  assign n23633 = ~n23631 & n23632 ;
  assign n23634 = ~n23629 & ~n23633 ;
  assign n23635 = ~n23625 & n23634 ;
  assign n23636 = ~n23624 & n23635 ;
  assign n23637 = n19076 & ~n23636 ;
  assign n23621 = n15880 & ~n19177 ;
  assign n23638 = n15875 & n16426 ;
  assign n23648 = ~n23621 & ~n23638 ;
  assign n23649 = ~n23637 & n23648 ;
  assign n23650 = ~n23647 & n23649 ;
  assign n23651 = n19075 & ~n23650 ;
  assign n23652 = ~n23620 & ~n23651 ;
  assign n23653 = \P3_rd_reg/NET0131  & ~n23652 ;
  assign n23619 = ~\P3_rd_reg/NET0131  & \P4_reg3_reg[21]/NET0131  ;
  assign n23654 = n15744 & n15880 ;
  assign n23655 = ~n23619 & ~n23654 ;
  assign n23656 = ~n23653 & n23655 ;
  assign n23657 = \P4_reg2_reg[21]/NET0131  & ~n18665 ;
  assign n23658 = \P4_reg2_reg[21]/NET0131  & n19073 ;
  assign n23660 = \P4_reg2_reg[21]/NET0131  & ~n20673 ;
  assign n23661 = n20673 & n23644 ;
  assign n23662 = ~n23660 & ~n23661 ;
  assign n23663 = n18483 & ~n23662 ;
  assign n23664 = n20673 & ~n23635 ;
  assign n23665 = n20673 & n23623 ;
  assign n23666 = ~n23660 & ~n23665 ;
  assign n23667 = n18604 & ~n23666 ;
  assign n23659 = \P4_reg2_reg[21]/NET0131  & ~n23489 ;
  assign n23668 = n15880 & n16426 ;
  assign n23669 = ~n23659 & ~n23668 ;
  assign n23670 = ~n23667 & n23669 ;
  assign n23671 = ~n23664 & n23670 ;
  assign n23672 = ~n23663 & n23671 ;
  assign n23673 = n19075 & ~n23672 ;
  assign n23674 = ~n23658 & ~n23673 ;
  assign n23675 = \P3_rd_reg/NET0131  & ~n23674 ;
  assign n23676 = ~n23657 & ~n23675 ;
  assign n23677 = n20665 & ~n23259 ;
  assign n23678 = ~n18670 & ~n20661 ;
  assign n23679 = n18666 & ~n23678 ;
  assign n23680 = n23414 & n23679 ;
  assign n23681 = ~n23249 & n23680 ;
  assign n23682 = \P4_reg0_reg[17]/NET0131  & ~n23681 ;
  assign n23683 = ~n23677 & ~n23682 ;
  assign n23684 = \P4_reg0_reg[1]/NET0131  & ~n18665 ;
  assign n23685 = \P4_reg0_reg[1]/NET0131  & n19073 ;
  assign n23686 = \P4_reg0_reg[1]/NET0131  & ~n20661 ;
  assign n23687 = n20661 & n23275 ;
  assign n23688 = ~n23686 & ~n23687 ;
  assign n23689 = n18483 & ~n23688 ;
  assign n23693 = n20661 & ~n23292 ;
  assign n23690 = n18604 & ~n20661 ;
  assign n23691 = n23414 & ~n23690 ;
  assign n23692 = \P4_reg0_reg[1]/NET0131  & ~n23691 ;
  assign n23694 = ~n16098 & n20661 ;
  assign n23695 = ~n23686 & ~n23694 ;
  assign n23696 = n18486 & ~n23695 ;
  assign n23697 = ~n23692 & ~n23696 ;
  assign n23698 = ~n23693 & n23697 ;
  assign n23699 = ~n23689 & n23698 ;
  assign n23700 = n19075 & ~n23699 ;
  assign n23701 = ~n23685 & ~n23700 ;
  assign n23702 = \P3_rd_reg/NET0131  & ~n23701 ;
  assign n23703 = ~n23684 & ~n23702 ;
  assign n23705 = \P4_reg0_reg[21]/NET0131  & ~n20661 ;
  assign n23706 = n20665 & n23644 ;
  assign n23707 = ~n23705 & ~n23706 ;
  assign n23708 = n18483 & ~n23707 ;
  assign n23704 = n20665 & ~n23636 ;
  assign n23709 = \P4_reg0_reg[21]/NET0131  & ~n21854 ;
  assign n23710 = ~n23704 & ~n23709 ;
  assign n23711 = ~n23708 & n23710 ;
  assign n23712 = n20665 & ~n23326 ;
  assign n23713 = \P4_reg0_reg[2]/NET0131  & ~n21855 ;
  assign n23714 = ~n23712 & ~n23713 ;
  assign n23715 = n20665 & ~n23357 ;
  assign n23716 = \P4_reg0_reg[5]/NET0131  & ~n21855 ;
  assign n23717 = ~n23715 & ~n23716 ;
  assign n23719 = \P4_reg0_reg[9]/NET0131  & ~n20661 ;
  assign n23720 = n20665 & n23387 ;
  assign n23721 = ~n23719 & ~n23720 ;
  assign n23722 = n18483 & ~n23721 ;
  assign n23718 = n20665 & ~n23382 ;
  assign n23723 = \P4_reg0_reg[9]/NET0131  & ~n21854 ;
  assign n23724 = ~n23718 & ~n23723 ;
  assign n23725 = ~n23722 & n23724 ;
  assign n23726 = \P2_P1_EAX_reg[24]/NET0131  & ~n21100 ;
  assign n23730 = n11463 & n22337 ;
  assign n23731 = \P2_P1_EAX_reg[24]/NET0131  & ~n22337 ;
  assign n23732 = ~n23730 & ~n23731 ;
  assign n23733 = n21068 & ~n23732 ;
  assign n23734 = n21022 & ~n21045 ;
  assign n23735 = ~n21072 & ~n23734 ;
  assign n23736 = \P2_P1_EAX_reg[24]/NET0131  & ~n23735 ;
  assign n23740 = n21022 & n21044 ;
  assign n23741 = \P2_P1_EAX_reg[23]/NET0131  & ~\P2_P1_EAX_reg[24]/NET0131  ;
  assign n23742 = n23740 & n23741 ;
  assign n23727 = ~n20791 & n20822 ;
  assign n23728 = ~n20823 & ~n23727 ;
  assign n23729 = n20728 & n23728 ;
  assign n23737 = n11385 & n22337 ;
  assign n23738 = ~n23731 & ~n23737 ;
  assign n23739 = n21062 & ~n23738 ;
  assign n23743 = ~n23729 & ~n23739 ;
  assign n23744 = ~n23742 & n23743 ;
  assign n23745 = ~n23736 & n23744 ;
  assign n23746 = ~n23733 & n23745 ;
  assign n23747 = n11623 & ~n23746 ;
  assign n23748 = ~n23726 & ~n23747 ;
  assign n23749 = \P4_reg1_reg[17]/NET0131  & ~n18664 ;
  assign n23750 = n18667 & ~n23257 ;
  assign n23751 = ~n23749 & ~n23750 ;
  assign n23752 = n18483 & ~n23751 ;
  assign n23753 = n23240 & n23462 ;
  assign n23754 = n23251 & ~n23753 ;
  assign n23755 = n18667 & ~n23754 ;
  assign n23756 = n21863 & ~n23249 ;
  assign n23757 = \P4_reg1_reg[17]/NET0131  & ~n23756 ;
  assign n23758 = ~n23755 & ~n23757 ;
  assign n23759 = ~n23752 & n23758 ;
  assign n23761 = \P4_reg1_reg[1]/NET0131  & ~n18664 ;
  assign n23762 = n18667 & n23275 ;
  assign n23763 = ~n23761 & ~n23762 ;
  assign n23764 = n18483 & ~n23763 ;
  assign n23760 = \P4_reg1_reg[1]/NET0131  & ~n18678 ;
  assign n23768 = n18664 & ~n23291 ;
  assign n23765 = ~n16098 & n18664 ;
  assign n23766 = ~n23761 & ~n23765 ;
  assign n23767 = n18486 & ~n23766 ;
  assign n23769 = n18664 & n23280 ;
  assign n23770 = ~n23761 & ~n23769 ;
  assign n23771 = n18604 & ~n23770 ;
  assign n23772 = ~n23767 & ~n23771 ;
  assign n23773 = ~n23768 & n23772 ;
  assign n23774 = n18666 & ~n23773 ;
  assign n23775 = ~n23760 & ~n23774 ;
  assign n23776 = ~n23764 & n23775 ;
  assign n23777 = \P4_reg1_reg[2]/NET0131  & ~n18679 ;
  assign n23778 = n18667 & ~n23326 ;
  assign n23779 = ~n23777 & ~n23778 ;
  assign n23780 = \P2_P1_EAX_reg[25]/NET0131  & ~n21100 ;
  assign n23784 = ~n11483 & n22337 ;
  assign n23785 = \P2_P1_EAX_reg[25]/NET0131  & ~n22337 ;
  assign n23786 = ~n23784 & ~n23785 ;
  assign n23787 = n21068 & ~n23786 ;
  assign n23788 = ~\P2_P1_EAX_reg[25]/NET0131  & ~n21046 ;
  assign n23789 = n21022 & ~n21047 ;
  assign n23790 = ~n23788 & n23789 ;
  assign n23791 = \P2_P1_EAX_reg[25]/NET0131  & n21072 ;
  assign n23781 = ~n20823 & n20854 ;
  assign n23782 = ~n20855 & ~n23781 ;
  assign n23783 = n20728 & n23782 ;
  assign n23792 = n11386 & n22337 ;
  assign n23793 = ~n23785 & ~n23792 ;
  assign n23794 = n21062 & ~n23793 ;
  assign n23795 = ~n23783 & ~n23794 ;
  assign n23796 = ~n23791 & n23795 ;
  assign n23797 = ~n23790 & n23796 ;
  assign n23798 = ~n23787 & n23797 ;
  assign n23799 = n11623 & ~n23798 ;
  assign n23800 = ~n23780 & ~n23799 ;
  assign n23801 = \P4_reg1_reg[5]/NET0131  & ~n18679 ;
  assign n23802 = n18667 & ~n23357 ;
  assign n23803 = ~n23801 & ~n23802 ;
  assign n23804 = \P4_reg2_reg[13]/NET0131  & ~n18665 ;
  assign n23805 = \P4_reg2_reg[13]/NET0131  & n19073 ;
  assign n23807 = n20673 & ~n23210 ;
  assign n23808 = ~\P4_reg2_reg[13]/NET0131  & ~n20673 ;
  assign n23809 = n18483 & ~n23808 ;
  assign n23810 = ~n23807 & n23809 ;
  assign n23811 = n20673 & ~n23226 ;
  assign n23806 = \P4_reg2_reg[13]/NET0131  & ~n20682 ;
  assign n23812 = n15959 & n16426 ;
  assign n23813 = ~n23806 & ~n23812 ;
  assign n23814 = ~n23811 & n23813 ;
  assign n23815 = ~n23810 & n23814 ;
  assign n23816 = n19075 & ~n23815 ;
  assign n23817 = ~n23805 & ~n23816 ;
  assign n23818 = \P3_rd_reg/NET0131  & ~n23817 ;
  assign n23819 = ~n23804 & ~n23818 ;
  assign n23820 = \P2_P1_EAX_reg[26]/NET0131  & ~n21100 ;
  assign n23832 = n11504 & n22337 ;
  assign n23831 = ~\P2_P1_EAX_reg[26]/NET0131  & ~n22337 ;
  assign n23833 = n21068 & ~n23831 ;
  assign n23834 = ~n23832 & n23833 ;
  assign n23825 = n23162 & ~n23789 ;
  assign n23826 = \P2_P1_EAX_reg[26]/NET0131  & ~n23825 ;
  assign n23827 = ~\P2_P1_EAX_reg[26]/NET0131  & n21022 ;
  assign n23828 = n21047 & n23827 ;
  assign n23821 = ~n20855 & n20886 ;
  assign n23822 = n20720 & ~n20887 ;
  assign n23823 = ~n23821 & n23822 ;
  assign n23824 = n20727 & n23823 ;
  assign n23829 = n11373 & ~n21081 ;
  assign n23830 = n23167 & n23829 ;
  assign n23835 = ~n23824 & ~n23830 ;
  assign n23836 = ~n23828 & n23835 ;
  assign n23837 = ~n23826 & n23836 ;
  assign n23838 = ~n23834 & n23837 ;
  assign n23839 = n11623 & ~n23838 ;
  assign n23840 = ~n23820 & ~n23839 ;
  assign n23843 = n18666 & n20673 ;
  assign n23844 = ~n23257 & n23843 ;
  assign n23845 = \P4_reg2_reg[17]/NET0131  & ~n20673 ;
  assign n23846 = ~n23844 & ~n23845 ;
  assign n23847 = n18483 & ~n23846 ;
  assign n23841 = n18666 & n20682 ;
  assign n23842 = \P4_reg2_reg[17]/NET0131  & ~n23841 ;
  assign n23848 = n20673 & ~n23252 ;
  assign n23849 = n15932 & n16426 ;
  assign n23850 = ~n23848 & ~n23849 ;
  assign n23851 = n18666 & ~n23850 ;
  assign n23852 = ~n23842 & ~n23851 ;
  assign n23853 = ~n23847 & n23852 ;
  assign n23857 = ~n11520 & n22337 ;
  assign n23858 = \P2_P1_EAX_reg[27]/NET0131  & ~n22337 ;
  assign n23859 = ~n23857 & ~n23858 ;
  assign n23860 = n21068 & ~n23859 ;
  assign n23861 = \P2_P1_EAX_reg[27]/NET0131  & ~n22802 ;
  assign n23862 = n21048 & n22801 ;
  assign n23854 = ~n20887 & n20918 ;
  assign n23855 = ~n20919 & ~n23854 ;
  assign n23856 = n20728 & n23855 ;
  assign n23863 = n11388 & n22337 ;
  assign n23864 = ~n23858 & ~n23863 ;
  assign n23865 = n21062 & ~n23864 ;
  assign n23866 = ~n23856 & ~n23865 ;
  assign n23867 = ~n23862 & n23866 ;
  assign n23868 = ~n23861 & n23867 ;
  assign n23869 = ~n23860 & n23868 ;
  assign n23870 = n11623 & ~n23869 ;
  assign n23871 = \P2_P1_EAX_reg[27]/NET0131  & ~n21100 ;
  assign n23872 = ~n23870 & ~n23871 ;
  assign n23873 = \P4_reg2_reg[2]/NET0131  & ~n18665 ;
  assign n23874 = \P4_reg2_reg[2]/NET0131  & n19073 ;
  assign n23876 = n20673 & ~n23309 ;
  assign n23877 = ~\P4_reg2_reg[2]/NET0131  & ~n20673 ;
  assign n23878 = n18483 & ~n23877 ;
  assign n23879 = ~n23876 & n23878 ;
  assign n23880 = n20673 & ~n23325 ;
  assign n23875 = \P4_reg2_reg[2]/NET0131  & ~n20682 ;
  assign n23881 = \P4_reg3_reg[2]/NET0131  & n16426 ;
  assign n23882 = ~n23875 & ~n23881 ;
  assign n23883 = ~n23880 & n23882 ;
  assign n23884 = ~n23879 & n23883 ;
  assign n23885 = n19075 & ~n23884 ;
  assign n23886 = ~n23874 & ~n23885 ;
  assign n23887 = \P3_rd_reg/NET0131  & ~n23886 ;
  assign n23888 = ~n23873 & ~n23887 ;
  assign n23889 = \P4_reg2_reg[5]/NET0131  & ~n18665 ;
  assign n23890 = \P4_reg2_reg[5]/NET0131  & n19073 ;
  assign n23892 = n20673 & ~n23339 ;
  assign n23893 = ~\P4_reg2_reg[5]/NET0131  & ~n20673 ;
  assign n23894 = n18483 & ~n23893 ;
  assign n23895 = ~n23892 & n23894 ;
  assign n23896 = n20673 & ~n23356 ;
  assign n23891 = \P4_reg2_reg[5]/NET0131  & ~n20682 ;
  assign n23897 = n16044 & n16426 ;
  assign n23898 = ~n23891 & ~n23897 ;
  assign n23899 = ~n23896 & n23898 ;
  assign n23900 = ~n23895 & n23899 ;
  assign n23901 = n19075 & ~n23900 ;
  assign n23902 = ~n23890 & ~n23901 ;
  assign n23903 = \P3_rd_reg/NET0131  & ~n23902 ;
  assign n23904 = ~n23889 & ~n23903 ;
  assign n23905 = \P4_reg2_reg[9]/NET0131  & ~n18665 ;
  assign n23906 = \P4_reg2_reg[9]/NET0131  & n19073 ;
  assign n23908 = n20673 & ~n23389 ;
  assign n23907 = n16017 & n16426 ;
  assign n23909 = n18483 & ~n20673 ;
  assign n23910 = n20682 & ~n23909 ;
  assign n23911 = \P4_reg2_reg[9]/NET0131  & ~n23910 ;
  assign n23912 = ~n23907 & ~n23911 ;
  assign n23913 = ~n23908 & n23912 ;
  assign n23914 = n19075 & ~n23913 ;
  assign n23915 = ~n23906 & ~n23914 ;
  assign n23916 = \P3_rd_reg/NET0131  & ~n23915 ;
  assign n23917 = ~n23905 & ~n23916 ;
  assign n23922 = ~n8177 & n15365 ;
  assign n23923 = \P1_P1_EAX_reg[24]/NET0131  & ~n15365 ;
  assign n23924 = ~n23922 & ~n23923 ;
  assign n23925 = n15383 & ~n23924 ;
  assign n23926 = ~n7891 & n15365 ;
  assign n23927 = ~n23923 & ~n23926 ;
  assign n23928 = n15334 & ~n23927 ;
  assign n23929 = n15377 & ~n22826 ;
  assign n23930 = ~n22830 & ~n23929 ;
  assign n23931 = \P1_P1_EAX_reg[24]/NET0131  & ~n23930 ;
  assign n23932 = ~\P1_P1_EAX_reg[24]/NET0131  & n23568 ;
  assign n23918 = ~n15492 & n15523 ;
  assign n23919 = n15428 & ~n15524 ;
  assign n23920 = ~n23918 & n23919 ;
  assign n23921 = n15372 & n23920 ;
  assign n23933 = \P1_P1_EAX_reg[24]/NET0131  & n15386 ;
  assign n23934 = ~n23921 & ~n23933 ;
  assign n23935 = ~n23932 & n23934 ;
  assign n23936 = ~n23931 & n23935 ;
  assign n23937 = ~n23928 & n23936 ;
  assign n23938 = ~n23925 & n23937 ;
  assign n23939 = n8355 & ~n23938 ;
  assign n23940 = \P1_P1_EAX_reg[24]/NET0131  & ~n15326 ;
  assign n23941 = ~n23939 & ~n23940 ;
  assign n23942 = \P1_P1_EAX_reg[25]/NET0131  & ~n15326 ;
  assign n23954 = n8190 & n15365 ;
  assign n23953 = ~\P1_P1_EAX_reg[25]/NET0131  & ~n15365 ;
  assign n23955 = n15383 & ~n23953 ;
  assign n23956 = ~n23954 & n23955 ;
  assign n23946 = n15334 & ~n15335 ;
  assign n23947 = ~n15364 & n23946 ;
  assign n23948 = n7955 & n23947 ;
  assign n23949 = n15377 & ~n15411 ;
  assign n23950 = n22831 & ~n23949 ;
  assign n23951 = \P1_P1_EAX_reg[25]/NET0131  & ~n23950 ;
  assign n23943 = ~n15524 & n15555 ;
  assign n23944 = ~n15556 & ~n23943 ;
  assign n23945 = n22818 & n23944 ;
  assign n23952 = ~\P1_P1_EAX_reg[25]/NET0131  & n23194 ;
  assign n23957 = ~n23945 & ~n23952 ;
  assign n23958 = ~n23951 & n23957 ;
  assign n23959 = ~n23948 & n23958 ;
  assign n23960 = ~n23956 & n23959 ;
  assign n23961 = n8355 & ~n23960 ;
  assign n23962 = ~n23942 & ~n23961 ;
  assign n23966 = ~n8232 & n15365 ;
  assign n23967 = \P1_P1_EAX_reg[27]/NET0131  & ~n15365 ;
  assign n23968 = ~n23966 & ~n23967 ;
  assign n23969 = n15383 & ~n23968 ;
  assign n23970 = n7974 & n15365 ;
  assign n23971 = ~n23967 & ~n23970 ;
  assign n23972 = n15334 & ~n23971 ;
  assign n23973 = \P1_P1_EAX_reg[25]/NET0131  & \P1_P1_EAX_reg[26]/NET0131  ;
  assign n23974 = n15411 & n23973 ;
  assign n23975 = n15377 & ~n23974 ;
  assign n23976 = n23190 & ~n23975 ;
  assign n23977 = \P1_P1_EAX_reg[27]/NET0131  & ~n23976 ;
  assign n23963 = ~n15588 & n15619 ;
  assign n23964 = ~n15620 & ~n23963 ;
  assign n23965 = n22818 & n23964 ;
  assign n23978 = ~\P1_P1_EAX_reg[27]/NET0131  & n23973 ;
  assign n23979 = n23194 & n23978 ;
  assign n23980 = ~n23965 & ~n23979 ;
  assign n23981 = ~n23977 & n23980 ;
  assign n23982 = ~n23972 & n23981 ;
  assign n23983 = ~n23969 & n23982 ;
  assign n23984 = n8355 & ~n23983 ;
  assign n23985 = \P1_P1_EAX_reg[27]/NET0131  & ~n15326 ;
  assign n23986 = ~n23984 & ~n23985 ;
  assign n23987 = \P4_reg3_reg[0]/NET0131  & ~n18665 ;
  assign n23988 = \P4_reg3_reg[0]/NET0131  & n19073 ;
  assign n23991 = ~n16103 & n18669 ;
  assign n23992 = ~n16111 & ~n16288 ;
  assign n23993 = ~n18672 & ~n23992 ;
  assign n23994 = ~n23991 & ~n23993 ;
  assign n23995 = n16095 & ~n18449 ;
  assign n23996 = ~\P4_IR_reg[28]/NET0131  & ~n18450 ;
  assign n23997 = ~n23995 & n23996 ;
  assign n23998 = n18483 & n23997 ;
  assign n23999 = n23994 & ~n23998 ;
  assign n24000 = n19076 & ~n23999 ;
  assign n23989 = ~n16103 & n16426 ;
  assign n23990 = \P4_reg3_reg[0]/NET0131  & ~n19160 ;
  assign n24001 = ~n23989 & ~n23990 ;
  assign n24002 = ~n24000 & n24001 ;
  assign n24003 = n19075 & ~n24002 ;
  assign n24004 = ~n23988 & ~n24003 ;
  assign n24005 = \P3_rd_reg/NET0131  & ~n24004 ;
  assign n24006 = ~n23987 & ~n24005 ;
  assign n24007 = n20665 & ~n23227 ;
  assign n24008 = \P4_reg0_reg[13]/NET0131  & ~n21855 ;
  assign n24009 = ~n24007 & ~n24008 ;
  assign n24010 = n20665 & ~n23611 ;
  assign n24011 = \P4_reg0_reg[4]/NET0131  & ~n21855 ;
  assign n24012 = ~n24010 & ~n24011 ;
  assign n24013 = \P4_reg1_reg[13]/NET0131  & ~n18679 ;
  assign n24014 = n18667 & ~n23227 ;
  assign n24015 = ~n24013 & ~n24014 ;
  assign n24016 = \P4_reg1_reg[21]/NET0131  & ~n18665 ;
  assign n24017 = \P4_reg1_reg[21]/NET0131  & n19073 ;
  assign n24018 = \P4_reg1_reg[21]/NET0131  & ~n18664 ;
  assign n24019 = n18664 & n23644 ;
  assign n24020 = ~n24018 & ~n24019 ;
  assign n24021 = n18483 & ~n24020 ;
  assign n24022 = ~n23624 & n23634 ;
  assign n24023 = n18664 & ~n24022 ;
  assign n24024 = n15875 & n18664 ;
  assign n24025 = ~n24018 & ~n24024 ;
  assign n24026 = n18486 & ~n24025 ;
  assign n24027 = ~n16429 & ~n19105 ;
  assign n24028 = ~n18676 & n24027 ;
  assign n24029 = \P4_reg1_reg[21]/NET0131  & ~n24028 ;
  assign n24030 = ~n22685 & n24029 ;
  assign n24031 = ~n24026 & ~n24030 ;
  assign n24032 = ~n24023 & n24031 ;
  assign n24033 = ~n24021 & n24032 ;
  assign n24034 = n19075 & ~n24033 ;
  assign n24035 = ~n24017 & ~n24034 ;
  assign n24036 = \P3_rd_reg/NET0131  & ~n24035 ;
  assign n24037 = ~n24016 & ~n24036 ;
  assign n24038 = \P4_reg1_reg[4]/NET0131  & ~n18679 ;
  assign n24039 = n18667 & ~n23611 ;
  assign n24040 = ~n24038 & ~n24039 ;
  assign n24041 = \P4_reg1_reg[9]/NET0131  & ~n18665 ;
  assign n24042 = \P4_reg1_reg[9]/NET0131  & ~n18664 ;
  assign n24043 = n18664 & n23387 ;
  assign n24044 = ~n24042 & ~n24043 ;
  assign n24045 = n18483 & ~n24044 ;
  assign n24050 = n18664 & ~n23381 ;
  assign n24046 = n18486 & ~n18664 ;
  assign n24047 = ~n18673 & ~n18676 ;
  assign n24048 = ~n24046 & n24047 ;
  assign n24049 = \P4_reg1_reg[9]/NET0131  & ~n24048 ;
  assign n24051 = n18664 & n23369 ;
  assign n24052 = ~n24042 & ~n24051 ;
  assign n24053 = n18604 & ~n24052 ;
  assign n24054 = ~n24049 & ~n24053 ;
  assign n24055 = ~n24050 & n24054 ;
  assign n24056 = ~n24045 & n24055 ;
  assign n24057 = n19075 & ~n24056 ;
  assign n24058 = \P4_reg1_reg[9]/NET0131  & n19073 ;
  assign n24059 = ~n24057 & ~n24058 ;
  assign n24060 = \P3_rd_reg/NET0131  & ~n24059 ;
  assign n24061 = ~n24041 & ~n24060 ;
  assign n24062 = \P4_reg2_reg[1]/NET0131  & ~n18665 ;
  assign n24063 = \P4_reg2_reg[1]/NET0131  & n19073 ;
  assign n24068 = n20673 & ~n23275 ;
  assign n24067 = ~\P4_reg2_reg[1]/NET0131  & ~n20673 ;
  assign n24069 = n18483 & ~n24067 ;
  assign n24070 = ~n24068 & n24069 ;
  assign n24065 = n20673 & ~n23293 ;
  assign n24064 = \P4_reg2_reg[1]/NET0131  & ~n20682 ;
  assign n24066 = \P4_reg3_reg[1]/NET0131  & n16426 ;
  assign n24071 = ~n24064 & ~n24066 ;
  assign n24072 = ~n24065 & n24071 ;
  assign n24073 = ~n24070 & n24072 ;
  assign n24074 = n19075 & ~n24073 ;
  assign n24075 = ~n24063 & ~n24074 ;
  assign n24076 = \P3_rd_reg/NET0131  & ~n24075 ;
  assign n24077 = ~n24062 & ~n24076 ;
  assign n24078 = \P4_reg2_reg[4]/NET0131  & ~n18665 ;
  assign n24079 = \P4_reg2_reg[4]/NET0131  & n19073 ;
  assign n24081 = n20673 & ~n23594 ;
  assign n24082 = ~\P4_reg2_reg[4]/NET0131  & ~n20673 ;
  assign n24083 = n18483 & ~n24082 ;
  assign n24084 = ~n24081 & n24083 ;
  assign n24085 = n20673 & ~n23610 ;
  assign n24080 = n16057 & n16426 ;
  assign n24086 = \P4_reg2_reg[4]/NET0131  & ~n20682 ;
  assign n24087 = ~n24080 & ~n24086 ;
  assign n24088 = ~n24085 & n24087 ;
  assign n24089 = ~n24084 & n24088 ;
  assign n24090 = n19075 & ~n24089 ;
  assign n24091 = ~n24079 & ~n24090 ;
  assign n24092 = \P3_rd_reg/NET0131  & ~n24091 ;
  assign n24093 = ~n24078 & ~n24092 ;
  assign n24095 = \P4_reg0_reg[0]/NET0131  & ~n20661 ;
  assign n24096 = n20665 & n23997 ;
  assign n24097 = ~n24095 & ~n24096 ;
  assign n24098 = n18483 & ~n24097 ;
  assign n24094 = n20665 & ~n23994 ;
  assign n24099 = \P4_reg0_reg[0]/NET0131  & ~n21854 ;
  assign n24100 = ~n24094 & ~n24099 ;
  assign n24101 = ~n24098 & n24100 ;
  assign n24102 = \P2_P1_EAX_reg[23]/NET0131  & ~n21100 ;
  assign n24106 = ~n11354 & n22337 ;
  assign n24107 = \P2_P1_EAX_reg[23]/NET0131  & ~n22337 ;
  assign n24108 = ~n24106 & ~n24107 ;
  assign n24109 = n21068 & ~n24108 ;
  assign n24114 = n21022 & ~n21044 ;
  assign n24115 = ~n21072 & ~n24114 ;
  assign n24116 = \P2_P1_EAX_reg[23]/NET0131  & ~n24115 ;
  assign n24113 = ~\P2_P1_EAX_reg[23]/NET0131  & n23740 ;
  assign n24103 = n20759 & n20790 ;
  assign n24104 = ~n20791 & ~n24103 ;
  assign n24105 = n20728 & n24104 ;
  assign n24110 = n11387 & n22337 ;
  assign n24111 = ~n24107 & ~n24110 ;
  assign n24112 = n21062 & ~n24111 ;
  assign n24117 = ~n24105 & ~n24112 ;
  assign n24118 = ~n24113 & n24117 ;
  assign n24119 = ~n24116 & n24118 ;
  assign n24120 = ~n24109 & n24119 ;
  assign n24121 = n11623 & ~n24120 ;
  assign n24122 = ~n24102 & ~n24121 ;
  assign n24123 = \P4_reg1_reg[0]/NET0131  & ~n18679 ;
  assign n24124 = n18667 & ~n23999 ;
  assign n24125 = ~n24123 & ~n24124 ;
  assign n24127 = ~n8132 & n15365 ;
  assign n24128 = \P1_P1_EAX_reg[23]/NET0131  & ~n15365 ;
  assign n24129 = ~n24127 & ~n24128 ;
  assign n24130 = n15383 & ~n24129 ;
  assign n24133 = n7899 & n15365 ;
  assign n24134 = ~n24128 & ~n24133 ;
  assign n24135 = n15334 & ~n24134 ;
  assign n24131 = ~\P1_P1_EAX_reg[23]/NET0131  & ~n22825 ;
  assign n24132 = n23929 & ~n24131 ;
  assign n24126 = \P1_P1_EAX_reg[23]/NET0131  & ~n23190 ;
  assign n24136 = n15460 & n15491 ;
  assign n24137 = n15428 & ~n15492 ;
  assign n24138 = ~n24136 & n24137 ;
  assign n24139 = n15372 & n24138 ;
  assign n24140 = ~n24126 & ~n24139 ;
  assign n24141 = ~n24132 & n24140 ;
  assign n24142 = ~n24135 & n24141 ;
  assign n24143 = ~n24130 & n24142 ;
  assign n24144 = n8355 & ~n24143 ;
  assign n24145 = \P1_P1_EAX_reg[23]/NET0131  & ~n15326 ;
  assign n24146 = ~n24144 & ~n24145 ;
  assign n24148 = \P4_reg2_reg[0]/NET0131  & ~n20673 ;
  assign n24149 = n23843 & n23997 ;
  assign n24150 = ~n24148 & ~n24149 ;
  assign n24151 = n18483 & ~n24150 ;
  assign n24147 = \P4_reg2_reg[0]/NET0131  & ~n23841 ;
  assign n24152 = \P4_reg3_reg[0]/NET0131  & n16426 ;
  assign n24153 = n20673 & ~n23994 ;
  assign n24154 = ~n24152 & ~n24153 ;
  assign n24155 = n18666 & ~n24154 ;
  assign n24156 = ~n24147 & ~n24155 ;
  assign n24157 = ~n24151 & n24156 ;
  assign n24159 = ~n8121 & n15365 ;
  assign n24160 = \P1_P1_EAX_reg[22]/NET0131  & ~n15365 ;
  assign n24161 = ~n24159 & ~n24160 ;
  assign n24162 = n15383 & ~n24161 ;
  assign n24167 = n7906 & n15365 ;
  assign n24168 = ~n24160 & ~n24167 ;
  assign n24169 = n15334 & ~n24168 ;
  assign n24163 = \P1_P1_EAX_reg[21]/NET0131  & n22824 ;
  assign n24164 = ~\P1_P1_EAX_reg[22]/NET0131  & ~n24163 ;
  assign n24165 = n15377 & ~n22825 ;
  assign n24166 = ~n24164 & n24165 ;
  assign n24158 = \P1_P1_EAX_reg[22]/NET0131  & ~n23190 ;
  assign n24170 = \P1_P1_InstQueue_reg[1][6]/NET0131  & n8291 ;
  assign n24171 = \P1_P1_InstQueue_reg[6][6]/NET0131  & n8323 ;
  assign n24172 = \P1_P1_InstQueue_reg[8][6]/NET0131  & n8307 ;
  assign n24186 = ~n24171 & ~n24172 ;
  assign n24173 = \P1_P1_InstQueue_reg[15][6]/NET0131  & n8329 ;
  assign n24174 = \P1_P1_InstQueue_reg[14][6]/NET0131  & n8312 ;
  assign n24187 = ~n24173 & ~n24174 ;
  assign n24196 = n24186 & n24187 ;
  assign n24197 = ~n24170 & n24196 ;
  assign n24185 = \P1_P1_InstQueue_reg[13][6]/NET0131  & n8303 ;
  assign n24183 = \P1_P1_InstQueue_reg[5][6]/NET0131  & n8314 ;
  assign n24184 = \P1_P1_InstQueue_reg[3][6]/NET0131  & n8309 ;
  assign n24192 = ~n24183 & ~n24184 ;
  assign n24193 = ~n24185 & n24192 ;
  assign n24179 = \P1_P1_InstQueue_reg[9][6]/NET0131  & n8316 ;
  assign n24180 = \P1_P1_InstQueue_reg[10][6]/NET0131  & n8318 ;
  assign n24190 = ~n24179 & ~n24180 ;
  assign n24181 = \P1_P1_InstQueue_reg[2][6]/NET0131  & n8321 ;
  assign n24182 = \P1_P1_InstQueue_reg[0][6]/NET0131  & n8327 ;
  assign n24191 = ~n24181 & ~n24182 ;
  assign n24194 = n24190 & n24191 ;
  assign n24175 = \P1_P1_InstQueue_reg[7][6]/NET0131  & n8295 ;
  assign n24176 = \P1_P1_InstQueue_reg[12][6]/NET0131  & n8325 ;
  assign n24188 = ~n24175 & ~n24176 ;
  assign n24177 = \P1_P1_InstQueue_reg[4][6]/NET0131  & n8299 ;
  assign n24178 = \P1_P1_InstQueue_reg[11][6]/NET0131  & n8305 ;
  assign n24189 = ~n24177 & ~n24178 ;
  assign n24195 = n24188 & n24189 ;
  assign n24198 = n24194 & n24195 ;
  assign n24199 = n24193 & n24198 ;
  assign n24200 = n24197 & n24199 ;
  assign n24201 = n22818 & ~n24200 ;
  assign n24202 = ~n24158 & ~n24201 ;
  assign n24203 = ~n24166 & n24202 ;
  assign n24204 = ~n24169 & n24203 ;
  assign n24205 = ~n24162 & n24204 ;
  assign n24206 = n8355 & ~n24205 ;
  assign n24207 = \P1_P1_EAX_reg[22]/NET0131  & ~n15326 ;
  assign n24208 = ~n24206 & ~n24207 ;
  assign n24209 = \P2_P1_EAX_reg[21]/NET0131  & ~n21100 ;
  assign n24242 = ~n11365 & n22337 ;
  assign n24243 = \P2_P1_EAX_reg[21]/NET0131  & ~n22337 ;
  assign n24244 = ~n24242 & ~n24243 ;
  assign n24245 = n21068 & ~n24244 ;
  assign n24246 = n21022 & ~n21042 ;
  assign n24247 = ~n21072 & ~n24246 ;
  assign n24248 = \P2_P1_EAX_reg[21]/NET0131  & ~n24247 ;
  assign n24252 = ~\P2_P1_EAX_reg[21]/NET0131  & n21022 ;
  assign n24253 = n21042 & n24252 ;
  assign n24221 = \P2_P1_InstQueue_reg[9][5]/NET0131  & n11651 ;
  assign n24214 = \P2_P1_InstQueue_reg[2][5]/NET0131  & n11647 ;
  assign n24210 = \P2_P1_InstQueue_reg[5][5]/NET0131  & n11654 ;
  assign n24211 = \P2_P1_InstQueue_reg[13][5]/NET0131  & n11634 ;
  assign n24226 = ~n24210 & ~n24211 ;
  assign n24236 = ~n24214 & n24226 ;
  assign n24237 = ~n24221 & n24236 ;
  assign n24222 = \P2_P1_InstQueue_reg[11][5]/NET0131  & n11659 ;
  assign n24223 = \P2_P1_InstQueue_reg[12][5]/NET0131  & n11656 ;
  assign n24231 = ~n24222 & ~n24223 ;
  assign n24224 = \P2_P1_InstQueue_reg[7][5]/NET0131  & n11667 ;
  assign n24225 = \P2_P1_InstQueue_reg[8][5]/NET0131  & n11638 ;
  assign n24232 = ~n24224 & ~n24225 ;
  assign n24233 = n24231 & n24232 ;
  assign n24217 = \P2_P1_InstQueue_reg[14][5]/NET0131  & n11665 ;
  assign n24218 = \P2_P1_InstQueue_reg[6][5]/NET0131  & n11663 ;
  assign n24229 = ~n24217 & ~n24218 ;
  assign n24219 = \P2_P1_InstQueue_reg[10][5]/NET0131  & n11661 ;
  assign n24220 = \P2_P1_InstQueue_reg[3][5]/NET0131  & n11669 ;
  assign n24230 = ~n24219 & ~n24220 ;
  assign n24234 = n24229 & n24230 ;
  assign n24212 = \P2_P1_InstQueue_reg[15][5]/NET0131  & n11673 ;
  assign n24213 = \P2_P1_InstQueue_reg[1][5]/NET0131  & n11643 ;
  assign n24227 = ~n24212 & ~n24213 ;
  assign n24215 = \P2_P1_InstQueue_reg[0][5]/NET0131  & n11641 ;
  assign n24216 = \P2_P1_InstQueue_reg[4][5]/NET0131  & n11671 ;
  assign n24228 = ~n24215 & ~n24216 ;
  assign n24235 = n24227 & n24228 ;
  assign n24238 = n24234 & n24235 ;
  assign n24239 = n24233 & n24238 ;
  assign n24240 = n24237 & n24239 ;
  assign n24241 = n20728 & ~n24240 ;
  assign n24249 = n11378 & n22337 ;
  assign n24250 = ~n24243 & ~n24249 ;
  assign n24251 = n21062 & ~n24250 ;
  assign n24254 = ~n24241 & ~n24251 ;
  assign n24255 = ~n24253 & n24254 ;
  assign n24256 = ~n24248 & n24255 ;
  assign n24257 = ~n24245 & n24256 ;
  assign n24258 = n11623 & ~n24257 ;
  assign n24259 = ~n24209 & ~n24258 ;
  assign n24292 = ~n11342 & n22337 ;
  assign n24293 = \P2_P1_EAX_reg[22]/NET0131  & ~n22337 ;
  assign n24294 = ~n24292 & ~n24293 ;
  assign n24295 = n21068 & ~n24294 ;
  assign n24296 = \P2_P1_EAX_reg[22]/NET0131  & ~n24115 ;
  assign n24297 = n21043 & n24114 ;
  assign n24271 = \P2_P1_InstQueue_reg[9][6]/NET0131  & n11651 ;
  assign n24264 = \P2_P1_InstQueue_reg[2][6]/NET0131  & n11647 ;
  assign n24260 = \P2_P1_InstQueue_reg[5][6]/NET0131  & n11654 ;
  assign n24261 = \P2_P1_InstQueue_reg[13][6]/NET0131  & n11634 ;
  assign n24276 = ~n24260 & ~n24261 ;
  assign n24286 = ~n24264 & n24276 ;
  assign n24287 = ~n24271 & n24286 ;
  assign n24272 = \P2_P1_InstQueue_reg[11][6]/NET0131  & n11659 ;
  assign n24273 = \P2_P1_InstQueue_reg[12][6]/NET0131  & n11656 ;
  assign n24281 = ~n24272 & ~n24273 ;
  assign n24274 = \P2_P1_InstQueue_reg[7][6]/NET0131  & n11667 ;
  assign n24275 = \P2_P1_InstQueue_reg[8][6]/NET0131  & n11638 ;
  assign n24282 = ~n24274 & ~n24275 ;
  assign n24283 = n24281 & n24282 ;
  assign n24267 = \P2_P1_InstQueue_reg[14][6]/NET0131  & n11665 ;
  assign n24268 = \P2_P1_InstQueue_reg[6][6]/NET0131  & n11663 ;
  assign n24279 = ~n24267 & ~n24268 ;
  assign n24269 = \P2_P1_InstQueue_reg[10][6]/NET0131  & n11661 ;
  assign n24270 = \P2_P1_InstQueue_reg[3][6]/NET0131  & n11669 ;
  assign n24280 = ~n24269 & ~n24270 ;
  assign n24284 = n24279 & n24280 ;
  assign n24262 = \P2_P1_InstQueue_reg[15][6]/NET0131  & n11673 ;
  assign n24263 = \P2_P1_InstQueue_reg[1][6]/NET0131  & n11643 ;
  assign n24277 = ~n24262 & ~n24263 ;
  assign n24265 = \P2_P1_InstQueue_reg[0][6]/NET0131  & n11641 ;
  assign n24266 = \P2_P1_InstQueue_reg[4][6]/NET0131  & n11671 ;
  assign n24278 = ~n24265 & ~n24266 ;
  assign n24285 = n24277 & n24278 ;
  assign n24288 = n24284 & n24285 ;
  assign n24289 = n24283 & n24288 ;
  assign n24290 = n24287 & n24289 ;
  assign n24291 = n20728 & ~n24290 ;
  assign n24298 = n11383 & n22337 ;
  assign n24299 = ~n24293 & ~n24298 ;
  assign n24300 = n21062 & ~n24299 ;
  assign n24301 = ~n24291 & ~n24300 ;
  assign n24302 = ~n24297 & n24301 ;
  assign n24303 = ~n24296 & n24302 ;
  assign n24304 = ~n24295 & n24303 ;
  assign n24305 = n11623 & ~n24304 ;
  assign n24306 = \P2_P1_EAX_reg[22]/NET0131  & ~n21100 ;
  assign n24307 = ~n24305 & ~n24306 ;
  assign n24308 = \P1_P1_EAX_reg[14]/NET0131  & ~n15326 ;
  assign n24341 = ~n15364 & ~n15384 ;
  assign n24342 = ~n15335 & n24341 ;
  assign n24343 = ~n22858 & n24342 ;
  assign n24344 = n15377 & ~n15400 ;
  assign n24345 = ~n15365 & ~n15384 ;
  assign n24346 = n23190 & ~n24345 ;
  assign n24347 = ~n24344 & n24346 ;
  assign n24348 = \P1_P1_EAX_reg[14]/NET0131  & ~n24347 ;
  assign n24309 = \P1_P1_InstQueue_reg[0][6]/NET0131  & n8291 ;
  assign n24310 = \P1_P1_InstQueue_reg[13][6]/NET0131  & n8312 ;
  assign n24311 = \P1_P1_InstQueue_reg[2][6]/NET0131  & n8309 ;
  assign n24325 = ~n24310 & ~n24311 ;
  assign n24312 = \P1_P1_InstQueue_reg[15][6]/NET0131  & n8327 ;
  assign n24313 = \P1_P1_InstQueue_reg[4][6]/NET0131  & n8314 ;
  assign n24326 = ~n24312 & ~n24313 ;
  assign n24335 = n24325 & n24326 ;
  assign n24336 = ~n24309 & n24335 ;
  assign n24324 = \P1_P1_InstQueue_reg[7][6]/NET0131  & n8307 ;
  assign n24322 = \P1_P1_InstQueue_reg[11][6]/NET0131  & n8325 ;
  assign n24323 = \P1_P1_InstQueue_reg[6][6]/NET0131  & n8295 ;
  assign n24331 = ~n24322 & ~n24323 ;
  assign n24332 = ~n24324 & n24331 ;
  assign n24318 = \P1_P1_InstQueue_reg[8][6]/NET0131  & n8316 ;
  assign n24319 = \P1_P1_InstQueue_reg[1][6]/NET0131  & n8321 ;
  assign n24329 = ~n24318 & ~n24319 ;
  assign n24320 = \P1_P1_InstQueue_reg[9][6]/NET0131  & n8318 ;
  assign n24321 = \P1_P1_InstQueue_reg[12][6]/NET0131  & n8303 ;
  assign n24330 = ~n24320 & ~n24321 ;
  assign n24333 = n24329 & n24330 ;
  assign n24314 = \P1_P1_InstQueue_reg[10][6]/NET0131  & n8305 ;
  assign n24315 = \P1_P1_InstQueue_reg[14][6]/NET0131  & n8329 ;
  assign n24327 = ~n24314 & ~n24315 ;
  assign n24316 = \P1_P1_InstQueue_reg[5][6]/NET0131  & n8323 ;
  assign n24317 = \P1_P1_InstQueue_reg[3][6]/NET0131  & n8299 ;
  assign n24328 = ~n24316 & ~n24317 ;
  assign n24334 = n24327 & n24328 ;
  assign n24337 = n24333 & n24334 ;
  assign n24338 = n24332 & n24337 ;
  assign n24339 = n24336 & n24338 ;
  assign n24340 = n22818 & ~n24339 ;
  assign n24349 = ~\P1_P1_EAX_reg[14]/NET0131  & n15377 ;
  assign n24350 = n15400 & n24349 ;
  assign n24351 = ~n24340 & ~n24350 ;
  assign n24352 = ~n24348 & n24351 ;
  assign n24353 = ~n24343 & n24352 ;
  assign n24354 = n8355 & ~n24353 ;
  assign n24355 = ~n24308 & ~n24354 ;
  assign n24358 = ~n7926 & ~n8000 ;
  assign n24359 = n24342 & ~n24358 ;
  assign n24356 = n15377 & ~n15402 ;
  assign n24360 = n24346 & ~n24356 ;
  assign n24361 = \P1_P1_EAX_reg[15]/NET0131  & ~n24360 ;
  assign n24357 = n15401 & n24356 ;
  assign n24362 = \P1_P1_InstQueue_reg[0][7]/NET0131  & n8291 ;
  assign n24363 = \P1_P1_InstQueue_reg[5][7]/NET0131  & n8323 ;
  assign n24364 = \P1_P1_InstQueue_reg[4][7]/NET0131  & n8314 ;
  assign n24378 = ~n24363 & ~n24364 ;
  assign n24365 = \P1_P1_InstQueue_reg[6][7]/NET0131  & n8295 ;
  assign n24366 = \P1_P1_InstQueue_reg[12][7]/NET0131  & n8303 ;
  assign n24379 = ~n24365 & ~n24366 ;
  assign n24388 = n24378 & n24379 ;
  assign n24389 = ~n24362 & n24388 ;
  assign n24377 = \P1_P1_InstQueue_reg[7][7]/NET0131  & n8307 ;
  assign n24375 = \P1_P1_InstQueue_reg[10][7]/NET0131  & n8305 ;
  assign n24376 = \P1_P1_InstQueue_reg[2][7]/NET0131  & n8309 ;
  assign n24384 = ~n24375 & ~n24376 ;
  assign n24385 = ~n24377 & n24384 ;
  assign n24371 = \P1_P1_InstQueue_reg[8][7]/NET0131  & n8316 ;
  assign n24372 = \P1_P1_InstQueue_reg[9][7]/NET0131  & n8318 ;
  assign n24382 = ~n24371 & ~n24372 ;
  assign n24373 = \P1_P1_InstQueue_reg[1][7]/NET0131  & n8321 ;
  assign n24374 = \P1_P1_InstQueue_reg[15][7]/NET0131  & n8327 ;
  assign n24383 = ~n24373 & ~n24374 ;
  assign n24386 = n24382 & n24383 ;
  assign n24367 = \P1_P1_InstQueue_reg[13][7]/NET0131  & n8312 ;
  assign n24368 = \P1_P1_InstQueue_reg[14][7]/NET0131  & n8329 ;
  assign n24380 = ~n24367 & ~n24368 ;
  assign n24369 = \P1_P1_InstQueue_reg[11][7]/NET0131  & n8325 ;
  assign n24370 = \P1_P1_InstQueue_reg[3][7]/NET0131  & n8299 ;
  assign n24381 = ~n24369 & ~n24370 ;
  assign n24387 = n24380 & n24381 ;
  assign n24390 = n24386 & n24387 ;
  assign n24391 = n24385 & n24390 ;
  assign n24392 = n24389 & n24391 ;
  assign n24393 = n22818 & ~n24392 ;
  assign n24394 = ~n24357 & ~n24393 ;
  assign n24395 = ~n24361 & n24394 ;
  assign n24396 = ~n24359 & n24395 ;
  assign n24397 = n8355 & ~n24396 ;
  assign n24398 = \P1_P1_EAX_reg[15]/NET0131  & ~n15326 ;
  assign n24399 = ~n24397 & ~n24398 ;
  assign n24432 = ~n8106 & n15365 ;
  assign n24433 = \P1_P1_EAX_reg[21]/NET0131  & ~n15365 ;
  assign n24434 = ~n24432 & ~n24433 ;
  assign n24435 = n15383 & ~n24434 ;
  assign n24436 = ~\P1_P1_EAX_reg[21]/NET0131  & ~n22824 ;
  assign n24437 = n15377 & ~n24163 ;
  assign n24438 = ~n24436 & n24437 ;
  assign n24439 = ~n7933 & n15365 ;
  assign n24440 = ~n24433 & ~n24439 ;
  assign n24441 = n15334 & ~n24440 ;
  assign n24400 = \P1_P1_InstQueue_reg[1][5]/NET0131  & n8291 ;
  assign n24401 = \P1_P1_InstQueue_reg[14][5]/NET0131  & n8312 ;
  assign n24402 = \P1_P1_InstQueue_reg[0][5]/NET0131  & n8327 ;
  assign n24416 = ~n24401 & ~n24402 ;
  assign n24403 = \P1_P1_InstQueue_reg[13][5]/NET0131  & n8303 ;
  assign n24404 = \P1_P1_InstQueue_reg[6][5]/NET0131  & n8323 ;
  assign n24417 = ~n24403 & ~n24404 ;
  assign n24426 = n24416 & n24417 ;
  assign n24427 = ~n24400 & n24426 ;
  assign n24415 = \P1_P1_InstQueue_reg[11][5]/NET0131  & n8305 ;
  assign n24413 = \P1_P1_InstQueue_reg[5][5]/NET0131  & n8314 ;
  assign n24414 = \P1_P1_InstQueue_reg[12][5]/NET0131  & n8325 ;
  assign n24422 = ~n24413 & ~n24414 ;
  assign n24423 = ~n24415 & n24422 ;
  assign n24409 = \P1_P1_InstQueue_reg[9][5]/NET0131  & n8316 ;
  assign n24410 = \P1_P1_InstQueue_reg[2][5]/NET0131  & n8321 ;
  assign n24420 = ~n24409 & ~n24410 ;
  assign n24411 = \P1_P1_InstQueue_reg[10][5]/NET0131  & n8318 ;
  assign n24412 = \P1_P1_InstQueue_reg[7][5]/NET0131  & n8295 ;
  assign n24421 = ~n24411 & ~n24412 ;
  assign n24424 = n24420 & n24421 ;
  assign n24405 = \P1_P1_InstQueue_reg[15][5]/NET0131  & n8329 ;
  assign n24406 = \P1_P1_InstQueue_reg[8][5]/NET0131  & n8307 ;
  assign n24418 = ~n24405 & ~n24406 ;
  assign n24407 = \P1_P1_InstQueue_reg[4][5]/NET0131  & n8299 ;
  assign n24408 = \P1_P1_InstQueue_reg[3][5]/NET0131  & n8309 ;
  assign n24419 = ~n24407 & ~n24408 ;
  assign n24425 = n24418 & n24419 ;
  assign n24428 = n24424 & n24425 ;
  assign n24429 = n24423 & n24428 ;
  assign n24430 = n24427 & n24429 ;
  assign n24431 = n22818 & ~n24430 ;
  assign n24442 = \P1_P1_EAX_reg[21]/NET0131  & ~n23190 ;
  assign n24443 = ~n24431 & ~n24442 ;
  assign n24444 = ~n24441 & n24443 ;
  assign n24445 = ~n24438 & n24444 ;
  assign n24446 = ~n24435 & n24445 ;
  assign n24447 = n8355 & ~n24446 ;
  assign n24448 = \P1_P1_EAX_reg[21]/NET0131  & ~n15326 ;
  assign n24449 = ~n24447 & ~n24448 ;
  assign n24482 = ~\P2_P1_EAX_reg[19]/NET0131  & ~n21040 ;
  assign n24483 = n21022 & ~n21041 ;
  assign n24484 = ~n24482 & n24483 ;
  assign n24485 = \P2_P1_EAX_reg[19]/NET0131  & n21072 ;
  assign n24486 = \P2_P1_EAX_reg[19]/NET0131  & ~n22337 ;
  assign n24490 = n11343 & n22337 ;
  assign n24491 = ~n24486 & ~n24490 ;
  assign n24492 = n21068 & ~n24491 ;
  assign n24461 = \P2_P1_InstQueue_reg[9][3]/NET0131  & n11651 ;
  assign n24454 = \P2_P1_InstQueue_reg[2][3]/NET0131  & n11647 ;
  assign n24450 = \P2_P1_InstQueue_reg[5][3]/NET0131  & n11654 ;
  assign n24451 = \P2_P1_InstQueue_reg[13][3]/NET0131  & n11634 ;
  assign n24466 = ~n24450 & ~n24451 ;
  assign n24476 = ~n24454 & n24466 ;
  assign n24477 = ~n24461 & n24476 ;
  assign n24462 = \P2_P1_InstQueue_reg[11][3]/NET0131  & n11659 ;
  assign n24463 = \P2_P1_InstQueue_reg[12][3]/NET0131  & n11656 ;
  assign n24471 = ~n24462 & ~n24463 ;
  assign n24464 = \P2_P1_InstQueue_reg[7][3]/NET0131  & n11667 ;
  assign n24465 = \P2_P1_InstQueue_reg[8][3]/NET0131  & n11638 ;
  assign n24472 = ~n24464 & ~n24465 ;
  assign n24473 = n24471 & n24472 ;
  assign n24457 = \P2_P1_InstQueue_reg[14][3]/NET0131  & n11665 ;
  assign n24458 = \P2_P1_InstQueue_reg[6][3]/NET0131  & n11663 ;
  assign n24469 = ~n24457 & ~n24458 ;
  assign n24459 = \P2_P1_InstQueue_reg[10][3]/NET0131  & n11661 ;
  assign n24460 = \P2_P1_InstQueue_reg[3][3]/NET0131  & n11669 ;
  assign n24470 = ~n24459 & ~n24460 ;
  assign n24474 = n24469 & n24470 ;
  assign n24452 = \P2_P1_InstQueue_reg[15][3]/NET0131  & n11673 ;
  assign n24453 = \P2_P1_InstQueue_reg[1][3]/NET0131  & n11643 ;
  assign n24467 = ~n24452 & ~n24453 ;
  assign n24455 = \P2_P1_InstQueue_reg[0][3]/NET0131  & n11641 ;
  assign n24456 = \P2_P1_InstQueue_reg[4][3]/NET0131  & n11671 ;
  assign n24468 = ~n24455 & ~n24456 ;
  assign n24475 = n24467 & n24468 ;
  assign n24478 = n24474 & n24475 ;
  assign n24479 = n24473 & n24478 ;
  assign n24480 = n24477 & n24479 ;
  assign n24481 = n20728 & ~n24480 ;
  assign n24487 = n11374 & n22337 ;
  assign n24488 = ~n24486 & ~n24487 ;
  assign n24489 = n21062 & ~n24488 ;
  assign n24493 = ~n24481 & ~n24489 ;
  assign n24494 = ~n24492 & n24493 ;
  assign n24495 = ~n24485 & n24494 ;
  assign n24496 = ~n24484 & n24495 ;
  assign n24497 = n11623 & ~n24496 ;
  assign n24498 = \P2_P1_EAX_reg[19]/NET0131  & ~n21100 ;
  assign n24499 = ~n24497 & ~n24498 ;
  assign n24508 = n23947 & ~n24358 ;
  assign n24500 = n15334 & n15335 ;
  assign n24501 = n15329 & n15368 ;
  assign n24502 = n15333 & n24501 ;
  assign n24503 = ~n15364 & n24502 ;
  assign n24504 = n15334 & ~n15364 ;
  assign n24505 = ~n24503 & ~n24504 ;
  assign n24506 = ~n24500 & ~n24505 ;
  assign n24507 = \P1_P1_lWord_reg[15]/NET0131  & ~n24506 ;
  assign n24509 = \P1_P1_EAX_reg[15]/NET0131  & n24503 ;
  assign n24510 = ~n24507 & ~n24509 ;
  assign n24511 = ~n24508 & n24510 ;
  assign n24512 = n8355 & ~n24511 ;
  assign n24513 = ~n8348 & ~n15325 ;
  assign n24514 = n15323 & ~n24513 ;
  assign n24515 = n8360 & n24514 ;
  assign n24516 = \P1_P1_lWord_reg[15]/NET0131  & ~n24515 ;
  assign n24517 = ~n24512 & ~n24516 ;
  assign n24518 = \P1_P1_EAX_reg[13]/NET0131  & ~n15326 ;
  assign n24519 = ~n8007 & n24342 ;
  assign n24520 = \P1_P1_EAX_reg[13]/NET0131  & ~n24347 ;
  assign n24521 = \P1_P1_InstQueue_reg[0][5]/NET0131  & n8291 ;
  assign n24522 = \P1_P1_InstQueue_reg[10][5]/NET0131  & n8305 ;
  assign n24523 = \P1_P1_InstQueue_reg[6][5]/NET0131  & n8295 ;
  assign n24537 = ~n24522 & ~n24523 ;
  assign n24524 = \P1_P1_InstQueue_reg[5][5]/NET0131  & n8323 ;
  assign n24525 = \P1_P1_InstQueue_reg[13][5]/NET0131  & n8312 ;
  assign n24538 = ~n24524 & ~n24525 ;
  assign n24547 = n24537 & n24538 ;
  assign n24548 = ~n24521 & n24547 ;
  assign n24536 = \P1_P1_InstQueue_reg[15][5]/NET0131  & n8327 ;
  assign n24534 = \P1_P1_InstQueue_reg[14][5]/NET0131  & n8329 ;
  assign n24535 = \P1_P1_InstQueue_reg[12][5]/NET0131  & n8303 ;
  assign n24543 = ~n24534 & ~n24535 ;
  assign n24544 = ~n24536 & n24543 ;
  assign n24530 = \P1_P1_InstQueue_reg[8][5]/NET0131  & n8316 ;
  assign n24531 = \P1_P1_InstQueue_reg[1][5]/NET0131  & n8321 ;
  assign n24541 = ~n24530 & ~n24531 ;
  assign n24532 = \P1_P1_InstQueue_reg[9][5]/NET0131  & n8318 ;
  assign n24533 = \P1_P1_InstQueue_reg[4][5]/NET0131  & n8314 ;
  assign n24542 = ~n24532 & ~n24533 ;
  assign n24545 = n24541 & n24542 ;
  assign n24526 = \P1_P1_InstQueue_reg[2][5]/NET0131  & n8309 ;
  assign n24527 = \P1_P1_InstQueue_reg[11][5]/NET0131  & n8325 ;
  assign n24539 = ~n24526 & ~n24527 ;
  assign n24528 = \P1_P1_InstQueue_reg[7][5]/NET0131  & n8307 ;
  assign n24529 = \P1_P1_InstQueue_reg[3][5]/NET0131  & n8299 ;
  assign n24540 = ~n24528 & ~n24529 ;
  assign n24546 = n24539 & n24540 ;
  assign n24549 = n24545 & n24546 ;
  assign n24550 = n24544 & n24549 ;
  assign n24551 = n24548 & n24550 ;
  assign n24552 = n22818 & ~n24551 ;
  assign n24553 = n15399 & n24344 ;
  assign n24554 = ~n24552 & ~n24553 ;
  assign n24555 = ~n24520 & n24554 ;
  assign n24556 = ~n24519 & n24555 ;
  assign n24557 = n8355 & ~n24556 ;
  assign n24558 = ~n24518 & ~n24557 ;
  assign n24559 = \P1_P1_EAX_reg[18]/NET0131  & ~n15326 ;
  assign n24561 = n8068 & n15365 ;
  assign n24560 = ~\P1_P1_EAX_reg[18]/NET0131  & ~n15365 ;
  assign n24562 = n15383 & ~n24560 ;
  assign n24563 = ~n24561 & n24562 ;
  assign n24566 = n15377 & ~n22821 ;
  assign n24567 = n22831 & ~n24566 ;
  assign n24568 = \P1_P1_EAX_reg[18]/NET0131  & ~n24567 ;
  assign n24564 = ~\P1_P1_EAX_reg[18]/NET0131  & n15377 ;
  assign n24565 = n22821 & n24564 ;
  assign n24569 = \P1_P1_InstQueue_reg[1][2]/NET0131  & n8291 ;
  assign n24570 = \P1_P1_InstQueue_reg[4][2]/NET0131  & n8299 ;
  assign n24571 = \P1_P1_InstQueue_reg[5][2]/NET0131  & n8314 ;
  assign n24585 = ~n24570 & ~n24571 ;
  assign n24572 = \P1_P1_InstQueue_reg[11][2]/NET0131  & n8305 ;
  assign n24573 = \P1_P1_InstQueue_reg[14][2]/NET0131  & n8312 ;
  assign n24586 = ~n24572 & ~n24573 ;
  assign n24595 = n24585 & n24586 ;
  assign n24596 = ~n24569 & n24595 ;
  assign n24584 = \P1_P1_InstQueue_reg[13][2]/NET0131  & n8303 ;
  assign n24582 = \P1_P1_InstQueue_reg[12][2]/NET0131  & n8325 ;
  assign n24583 = \P1_P1_InstQueue_reg[3][2]/NET0131  & n8309 ;
  assign n24591 = ~n24582 & ~n24583 ;
  assign n24592 = ~n24584 & n24591 ;
  assign n24578 = \P1_P1_InstQueue_reg[9][2]/NET0131  & n8316 ;
  assign n24579 = \P1_P1_InstQueue_reg[2][2]/NET0131  & n8321 ;
  assign n24589 = ~n24578 & ~n24579 ;
  assign n24580 = \P1_P1_InstQueue_reg[10][2]/NET0131  & n8318 ;
  assign n24581 = \P1_P1_InstQueue_reg[6][2]/NET0131  & n8323 ;
  assign n24590 = ~n24580 & ~n24581 ;
  assign n24593 = n24589 & n24590 ;
  assign n24574 = \P1_P1_InstQueue_reg[15][2]/NET0131  & n8329 ;
  assign n24575 = \P1_P1_InstQueue_reg[8][2]/NET0131  & n8307 ;
  assign n24587 = ~n24574 & ~n24575 ;
  assign n24576 = \P1_P1_InstQueue_reg[7][2]/NET0131  & n8295 ;
  assign n24577 = \P1_P1_InstQueue_reg[0][2]/NET0131  & n8327 ;
  assign n24588 = ~n24576 & ~n24577 ;
  assign n24594 = n24587 & n24588 ;
  assign n24597 = n24593 & n24594 ;
  assign n24598 = n24592 & n24597 ;
  assign n24599 = n24596 & n24598 ;
  assign n24600 = n22818 & ~n24599 ;
  assign n24601 = n7947 & n23947 ;
  assign n24602 = ~n24600 & ~n24601 ;
  assign n24603 = ~n24565 & n24602 ;
  assign n24604 = ~n24568 & n24603 ;
  assign n24605 = ~n24563 & n24604 ;
  assign n24606 = n8355 & ~n24605 ;
  assign n24607 = ~n24559 & ~n24606 ;
  assign n24640 = ~n8077 & n15365 ;
  assign n24641 = \P1_P1_EAX_reg[19]/NET0131  & ~n15365 ;
  assign n24642 = ~n24640 & ~n24641 ;
  assign n24643 = n15383 & ~n24642 ;
  assign n24644 = n15377 & ~n22823 ;
  assign n24645 = n23190 & ~n24644 ;
  assign n24646 = \P1_P1_EAX_reg[19]/NET0131  & ~n24645 ;
  assign n24647 = n22822 & n24644 ;
  assign n24608 = \P1_P1_InstQueue_reg[1][3]/NET0131  & n8291 ;
  assign n24609 = \P1_P1_InstQueue_reg[3][3]/NET0131  & n8309 ;
  assign n24610 = \P1_P1_InstQueue_reg[6][3]/NET0131  & n8323 ;
  assign n24624 = ~n24609 & ~n24610 ;
  assign n24611 = \P1_P1_InstQueue_reg[13][3]/NET0131  & n8303 ;
  assign n24612 = \P1_P1_InstQueue_reg[12][3]/NET0131  & n8325 ;
  assign n24625 = ~n24611 & ~n24612 ;
  assign n24634 = n24624 & n24625 ;
  assign n24635 = ~n24608 & n24634 ;
  assign n24623 = \P1_P1_InstQueue_reg[4][3]/NET0131  & n8299 ;
  assign n24621 = \P1_P1_InstQueue_reg[11][3]/NET0131  & n8305 ;
  assign n24622 = \P1_P1_InstQueue_reg[8][3]/NET0131  & n8307 ;
  assign n24630 = ~n24621 & ~n24622 ;
  assign n24631 = ~n24623 & n24630 ;
  assign n24617 = \P1_P1_InstQueue_reg[9][3]/NET0131  & n8316 ;
  assign n24618 = \P1_P1_InstQueue_reg[2][3]/NET0131  & n8321 ;
  assign n24628 = ~n24617 & ~n24618 ;
  assign n24619 = \P1_P1_InstQueue_reg[10][3]/NET0131  & n8318 ;
  assign n24620 = \P1_P1_InstQueue_reg[14][3]/NET0131  & n8312 ;
  assign n24629 = ~n24619 & ~n24620 ;
  assign n24632 = n24628 & n24629 ;
  assign n24613 = \P1_P1_InstQueue_reg[15][3]/NET0131  & n8329 ;
  assign n24614 = \P1_P1_InstQueue_reg[5][3]/NET0131  & n8314 ;
  assign n24626 = ~n24613 & ~n24614 ;
  assign n24615 = \P1_P1_InstQueue_reg[7][3]/NET0131  & n8295 ;
  assign n24616 = \P1_P1_InstQueue_reg[0][3]/NET0131  & n8327 ;
  assign n24627 = ~n24615 & ~n24616 ;
  assign n24633 = n24626 & n24627 ;
  assign n24636 = n24632 & n24633 ;
  assign n24637 = n24631 & n24636 ;
  assign n24638 = n24635 & n24637 ;
  assign n24639 = n22818 & ~n24638 ;
  assign n24648 = ~n7913 & n15365 ;
  assign n24649 = ~n24641 & ~n24648 ;
  assign n24650 = n15334 & ~n24649 ;
  assign n24651 = ~n24639 & ~n24650 ;
  assign n24652 = ~n24647 & n24651 ;
  assign n24653 = ~n24646 & n24652 ;
  assign n24654 = ~n24643 & n24653 ;
  assign n24655 = n8355 & ~n24654 ;
  assign n24656 = \P1_P1_EAX_reg[19]/NET0131  & ~n15326 ;
  assign n24657 = ~n24655 & ~n24656 ;
  assign n24658 = \P1_P1_EAX_reg[20]/NET0131  & ~n15326 ;
  assign n24691 = ~n8092 & n15365 ;
  assign n24692 = \P1_P1_EAX_reg[20]/NET0131  & ~n15365 ;
  assign n24693 = ~n24691 & ~n24692 ;
  assign n24694 = n15383 & ~n24693 ;
  assign n24695 = \P1_P1_EAX_reg[20]/NET0131  & ~n24645 ;
  assign n24696 = ~n7940 & n15365 ;
  assign n24697 = ~n24692 & ~n24696 ;
  assign n24698 = n15334 & ~n24697 ;
  assign n24659 = \P1_P1_InstQueue_reg[1][4]/NET0131  & n8291 ;
  assign n24660 = \P1_P1_InstQueue_reg[11][4]/NET0131  & n8305 ;
  assign n24661 = \P1_P1_InstQueue_reg[3][4]/NET0131  & n8309 ;
  assign n24675 = ~n24660 & ~n24661 ;
  assign n24662 = \P1_P1_InstQueue_reg[15][4]/NET0131  & n8329 ;
  assign n24663 = \P1_P1_InstQueue_reg[6][4]/NET0131  & n8323 ;
  assign n24676 = ~n24662 & ~n24663 ;
  assign n24685 = n24675 & n24676 ;
  assign n24686 = ~n24659 & n24685 ;
  assign n24674 = \P1_P1_InstQueue_reg[8][4]/NET0131  & n8307 ;
  assign n24672 = \P1_P1_InstQueue_reg[4][4]/NET0131  & n8299 ;
  assign n24673 = \P1_P1_InstQueue_reg[13][4]/NET0131  & n8303 ;
  assign n24681 = ~n24672 & ~n24673 ;
  assign n24682 = ~n24674 & n24681 ;
  assign n24668 = \P1_P1_InstQueue_reg[9][4]/NET0131  & n8316 ;
  assign n24669 = \P1_P1_InstQueue_reg[2][4]/NET0131  & n8321 ;
  assign n24679 = ~n24668 & ~n24669 ;
  assign n24670 = \P1_P1_InstQueue_reg[10][4]/NET0131  & n8318 ;
  assign n24671 = \P1_P1_InstQueue_reg[5][4]/NET0131  & n8314 ;
  assign n24680 = ~n24670 & ~n24671 ;
  assign n24683 = n24679 & n24680 ;
  assign n24664 = \P1_P1_InstQueue_reg[7][4]/NET0131  & n8295 ;
  assign n24665 = \P1_P1_InstQueue_reg[12][4]/NET0131  & n8325 ;
  assign n24677 = ~n24664 & ~n24665 ;
  assign n24666 = \P1_P1_InstQueue_reg[14][4]/NET0131  & n8312 ;
  assign n24667 = \P1_P1_InstQueue_reg[0][4]/NET0131  & n8327 ;
  assign n24678 = ~n24666 & ~n24667 ;
  assign n24684 = n24677 & n24678 ;
  assign n24687 = n24683 & n24684 ;
  assign n24688 = n24682 & n24687 ;
  assign n24689 = n24686 & n24688 ;
  assign n24690 = n22818 & ~n24689 ;
  assign n24699 = ~\P1_P1_EAX_reg[20]/NET0131  & n15377 ;
  assign n24700 = n22823 & n24699 ;
  assign n24701 = ~n24690 & ~n24700 ;
  assign n24702 = ~n24698 & n24701 ;
  assign n24703 = ~n24695 & n24702 ;
  assign n24704 = ~n24694 & n24703 ;
  assign n24705 = n8355 & ~n24704 ;
  assign n24706 = ~n24658 & ~n24705 ;
  assign n24707 = \P2_P1_EAX_reg[14]/NET0131  & ~n21100 ;
  assign n24710 = n21022 & ~n21035 ;
  assign n24711 = ~n21069 & ~n22337 ;
  assign n24712 = ~n21072 & ~n24711 ;
  assign n24713 = ~n24710 & n24712 ;
  assign n24714 = \P2_P1_EAX_reg[14]/NET0131  & ~n24713 ;
  assign n24708 = ~n21069 & n22337 ;
  assign n24709 = n11381 & n24708 ;
  assign n24720 = \P2_P1_InstQueue_reg[8][6]/NET0131  & n11651 ;
  assign n24719 = \P2_P1_InstQueue_reg[1][6]/NET0131  & n11647 ;
  assign n24715 = \P2_P1_InstQueue_reg[4][6]/NET0131  & n11654 ;
  assign n24716 = \P2_P1_InstQueue_reg[7][6]/NET0131  & n11638 ;
  assign n24731 = ~n24715 & ~n24716 ;
  assign n24741 = ~n24719 & n24731 ;
  assign n24742 = ~n24720 & n24741 ;
  assign n24727 = \P2_P1_InstQueue_reg[13][6]/NET0131  & n11665 ;
  assign n24728 = \P2_P1_InstQueue_reg[5][6]/NET0131  & n11663 ;
  assign n24736 = ~n24727 & ~n24728 ;
  assign n24729 = \P2_P1_InstQueue_reg[3][6]/NET0131  & n11671 ;
  assign n24730 = \P2_P1_InstQueue_reg[11][6]/NET0131  & n11656 ;
  assign n24737 = ~n24729 & ~n24730 ;
  assign n24738 = n24736 & n24737 ;
  assign n24723 = \P2_P1_InstQueue_reg[12][6]/NET0131  & n11634 ;
  assign n24724 = \P2_P1_InstQueue_reg[9][6]/NET0131  & n11661 ;
  assign n24734 = ~n24723 & ~n24724 ;
  assign n24725 = \P2_P1_InstQueue_reg[10][6]/NET0131  & n11659 ;
  assign n24726 = \P2_P1_InstQueue_reg[6][6]/NET0131  & n11667 ;
  assign n24735 = ~n24725 & ~n24726 ;
  assign n24739 = n24734 & n24735 ;
  assign n24717 = \P2_P1_InstQueue_reg[14][6]/NET0131  & n11673 ;
  assign n24718 = \P2_P1_InstQueue_reg[0][6]/NET0131  & n11643 ;
  assign n24732 = ~n24717 & ~n24718 ;
  assign n24721 = \P2_P1_InstQueue_reg[2][6]/NET0131  & n11669 ;
  assign n24722 = \P2_P1_InstQueue_reg[15][6]/NET0131  & n11641 ;
  assign n24733 = ~n24721 & ~n24722 ;
  assign n24740 = n24732 & n24733 ;
  assign n24743 = n24739 & n24740 ;
  assign n24744 = n24738 & n24743 ;
  assign n24745 = n24742 & n24744 ;
  assign n24746 = n20728 & ~n24745 ;
  assign n24747 = ~\P2_P1_EAX_reg[14]/NET0131  & n21022 ;
  assign n24748 = n21035 & n24747 ;
  assign n24749 = ~n24746 & ~n24748 ;
  assign n24750 = ~n24709 & n24749 ;
  assign n24751 = ~n24714 & n24750 ;
  assign n24752 = n11623 & ~n24751 ;
  assign n24753 = ~n24707 & ~n24752 ;
  assign n24754 = \P2_P1_EAX_reg[15]/NET0131  & ~n21100 ;
  assign n24756 = n21022 & ~n21036 ;
  assign n24757 = n24712 & ~n24756 ;
  assign n24758 = \P2_P1_EAX_reg[15]/NET0131  & ~n24757 ;
  assign n24791 = ~\P2_P1_EAX_reg[15]/NET0131  & n21022 ;
  assign n24792 = n21036 & n24791 ;
  assign n24755 = n11377 & n24708 ;
  assign n24764 = \P2_P1_InstQueue_reg[8][7]/NET0131  & n11651 ;
  assign n24763 = \P2_P1_InstQueue_reg[1][7]/NET0131  & n11647 ;
  assign n24759 = \P2_P1_InstQueue_reg[4][7]/NET0131  & n11654 ;
  assign n24760 = \P2_P1_InstQueue_reg[7][7]/NET0131  & n11638 ;
  assign n24775 = ~n24759 & ~n24760 ;
  assign n24785 = ~n24763 & n24775 ;
  assign n24786 = ~n24764 & n24785 ;
  assign n24771 = \P2_P1_InstQueue_reg[13][7]/NET0131  & n11665 ;
  assign n24772 = \P2_P1_InstQueue_reg[5][7]/NET0131  & n11663 ;
  assign n24780 = ~n24771 & ~n24772 ;
  assign n24773 = \P2_P1_InstQueue_reg[3][7]/NET0131  & n11671 ;
  assign n24774 = \P2_P1_InstQueue_reg[11][7]/NET0131  & n11656 ;
  assign n24781 = ~n24773 & ~n24774 ;
  assign n24782 = n24780 & n24781 ;
  assign n24767 = \P2_P1_InstQueue_reg[12][7]/NET0131  & n11634 ;
  assign n24768 = \P2_P1_InstQueue_reg[9][7]/NET0131  & n11661 ;
  assign n24778 = ~n24767 & ~n24768 ;
  assign n24769 = \P2_P1_InstQueue_reg[10][7]/NET0131  & n11659 ;
  assign n24770 = \P2_P1_InstQueue_reg[6][7]/NET0131  & n11667 ;
  assign n24779 = ~n24769 & ~n24770 ;
  assign n24783 = n24778 & n24779 ;
  assign n24761 = \P2_P1_InstQueue_reg[14][7]/NET0131  & n11673 ;
  assign n24762 = \P2_P1_InstQueue_reg[0][7]/NET0131  & n11643 ;
  assign n24776 = ~n24761 & ~n24762 ;
  assign n24765 = \P2_P1_InstQueue_reg[2][7]/NET0131  & n11669 ;
  assign n24766 = \P2_P1_InstQueue_reg[15][7]/NET0131  & n11641 ;
  assign n24777 = ~n24765 & ~n24766 ;
  assign n24784 = n24776 & n24777 ;
  assign n24787 = n24783 & n24784 ;
  assign n24788 = n24782 & n24787 ;
  assign n24789 = n24786 & n24788 ;
  assign n24790 = n20728 & ~n24789 ;
  assign n24793 = ~n24755 & ~n24790 ;
  assign n24794 = ~n24792 & n24793 ;
  assign n24795 = ~n24758 & n24794 ;
  assign n24796 = n11623 & ~n24795 ;
  assign n24797 = ~n24754 & ~n24796 ;
  assign n24830 = ~\P2_P1_EAX_reg[18]/NET0131  & ~n21039 ;
  assign n24831 = n21022 & ~n21040 ;
  assign n24832 = ~n24830 & n24831 ;
  assign n24833 = \P2_P1_EAX_reg[18]/NET0131  & n21072 ;
  assign n24834 = \P2_P1_EAX_reg[18]/NET0131  & ~n22337 ;
  assign n24838 = n11382 & n22337 ;
  assign n24839 = ~n24834 & ~n24838 ;
  assign n24840 = n21062 & ~n24839 ;
  assign n24809 = \P2_P1_InstQueue_reg[9][2]/NET0131  & n11651 ;
  assign n24802 = \P2_P1_InstQueue_reg[2][2]/NET0131  & n11647 ;
  assign n24798 = \P2_P1_InstQueue_reg[5][2]/NET0131  & n11654 ;
  assign n24799 = \P2_P1_InstQueue_reg[13][2]/NET0131  & n11634 ;
  assign n24814 = ~n24798 & ~n24799 ;
  assign n24824 = ~n24802 & n24814 ;
  assign n24825 = ~n24809 & n24824 ;
  assign n24810 = \P2_P1_InstQueue_reg[11][2]/NET0131  & n11659 ;
  assign n24811 = \P2_P1_InstQueue_reg[12][2]/NET0131  & n11656 ;
  assign n24819 = ~n24810 & ~n24811 ;
  assign n24812 = \P2_P1_InstQueue_reg[7][2]/NET0131  & n11667 ;
  assign n24813 = \P2_P1_InstQueue_reg[8][2]/NET0131  & n11638 ;
  assign n24820 = ~n24812 & ~n24813 ;
  assign n24821 = n24819 & n24820 ;
  assign n24805 = \P2_P1_InstQueue_reg[14][2]/NET0131  & n11665 ;
  assign n24806 = \P2_P1_InstQueue_reg[6][2]/NET0131  & n11663 ;
  assign n24817 = ~n24805 & ~n24806 ;
  assign n24807 = \P2_P1_InstQueue_reg[10][2]/NET0131  & n11661 ;
  assign n24808 = \P2_P1_InstQueue_reg[3][2]/NET0131  & n11669 ;
  assign n24818 = ~n24807 & ~n24808 ;
  assign n24822 = n24817 & n24818 ;
  assign n24800 = \P2_P1_InstQueue_reg[15][2]/NET0131  & n11673 ;
  assign n24801 = \P2_P1_InstQueue_reg[1][2]/NET0131  & n11643 ;
  assign n24815 = ~n24800 & ~n24801 ;
  assign n24803 = \P2_P1_InstQueue_reg[0][2]/NET0131  & n11641 ;
  assign n24804 = \P2_P1_InstQueue_reg[4][2]/NET0131  & n11671 ;
  assign n24816 = ~n24803 & ~n24804 ;
  assign n24823 = n24815 & n24816 ;
  assign n24826 = n24822 & n24823 ;
  assign n24827 = n24821 & n24826 ;
  assign n24828 = n24825 & n24827 ;
  assign n24829 = n20728 & ~n24828 ;
  assign n24835 = n11345 & n22337 ;
  assign n24836 = ~n24834 & ~n24835 ;
  assign n24837 = n21068 & ~n24836 ;
  assign n24841 = ~n24829 & ~n24837 ;
  assign n24842 = ~n24840 & n24841 ;
  assign n24843 = ~n24833 & n24842 ;
  assign n24844 = ~n24832 & n24843 ;
  assign n24845 = n11623 & ~n24844 ;
  assign n24846 = \P2_P1_EAX_reg[18]/NET0131  & ~n21100 ;
  assign n24847 = ~n24845 & ~n24846 ;
  assign n24880 = ~n11372 & n22337 ;
  assign n24881 = \P2_P1_EAX_reg[20]/NET0131  & ~n22337 ;
  assign n24882 = ~n24880 & ~n24881 ;
  assign n24883 = n21068 & ~n24882 ;
  assign n24884 = ~\P2_P1_EAX_reg[20]/NET0131  & ~n21041 ;
  assign n24885 = n24246 & ~n24884 ;
  assign n24886 = \P2_P1_EAX_reg[20]/NET0131  & n21072 ;
  assign n24859 = \P2_P1_InstQueue_reg[9][4]/NET0131  & n11651 ;
  assign n24852 = \P2_P1_InstQueue_reg[2][4]/NET0131  & n11647 ;
  assign n24848 = \P2_P1_InstQueue_reg[5][4]/NET0131  & n11654 ;
  assign n24849 = \P2_P1_InstQueue_reg[13][4]/NET0131  & n11634 ;
  assign n24864 = ~n24848 & ~n24849 ;
  assign n24874 = ~n24852 & n24864 ;
  assign n24875 = ~n24859 & n24874 ;
  assign n24860 = \P2_P1_InstQueue_reg[11][4]/NET0131  & n11659 ;
  assign n24861 = \P2_P1_InstQueue_reg[12][4]/NET0131  & n11656 ;
  assign n24869 = ~n24860 & ~n24861 ;
  assign n24862 = \P2_P1_InstQueue_reg[7][4]/NET0131  & n11667 ;
  assign n24863 = \P2_P1_InstQueue_reg[8][4]/NET0131  & n11638 ;
  assign n24870 = ~n24862 & ~n24863 ;
  assign n24871 = n24869 & n24870 ;
  assign n24855 = \P2_P1_InstQueue_reg[14][4]/NET0131  & n11665 ;
  assign n24856 = \P2_P1_InstQueue_reg[6][4]/NET0131  & n11663 ;
  assign n24867 = ~n24855 & ~n24856 ;
  assign n24857 = \P2_P1_InstQueue_reg[10][4]/NET0131  & n11661 ;
  assign n24858 = \P2_P1_InstQueue_reg[3][4]/NET0131  & n11669 ;
  assign n24868 = ~n24857 & ~n24858 ;
  assign n24872 = n24867 & n24868 ;
  assign n24850 = \P2_P1_InstQueue_reg[15][4]/NET0131  & n11673 ;
  assign n24851 = \P2_P1_InstQueue_reg[1][4]/NET0131  & n11643 ;
  assign n24865 = ~n24850 & ~n24851 ;
  assign n24853 = \P2_P1_InstQueue_reg[0][4]/NET0131  & n11641 ;
  assign n24854 = \P2_P1_InstQueue_reg[4][4]/NET0131  & n11671 ;
  assign n24866 = ~n24853 & ~n24854 ;
  assign n24873 = n24865 & n24866 ;
  assign n24876 = n24872 & n24873 ;
  assign n24877 = n24871 & n24876 ;
  assign n24878 = n24875 & n24877 ;
  assign n24879 = n20728 & ~n24878 ;
  assign n24887 = n11376 & n22337 ;
  assign n24888 = ~n24881 & ~n24887 ;
  assign n24889 = n21062 & ~n24888 ;
  assign n24890 = ~n24879 & ~n24889 ;
  assign n24891 = ~n24886 & n24890 ;
  assign n24892 = ~n24885 & n24891 ;
  assign n24893 = ~n24883 & n24892 ;
  assign n24894 = n11623 & ~n24893 ;
  assign n24895 = \P2_P1_EAX_reg[20]/NET0131  & ~n21100 ;
  assign n24896 = ~n24894 & ~n24895 ;
  assign n24897 = n20722 & n21057 ;
  assign n24898 = n21061 & n24897 ;
  assign n24899 = ~n21081 & n24898 ;
  assign n24901 = n21062 & ~n21081 ;
  assign n24902 = ~n24899 & ~n24901 ;
  assign n24903 = \P2_P1_lWord_reg[15]/NET0131  & n24902 ;
  assign n24900 = \P2_P1_EAX_reg[15]/NET0131  & n24899 ;
  assign n24904 = n11377 & n22337 ;
  assign n24905 = \P2_P1_lWord_reg[15]/NET0131  & n21073 ;
  assign n24906 = ~n24904 & ~n24905 ;
  assign n24907 = n21062 & ~n24906 ;
  assign n24908 = ~n24900 & ~n24907 ;
  assign n24909 = ~n24903 & n24908 ;
  assign n24910 = n11623 & ~n24909 ;
  assign n24911 = ~n11615 & ~n21099 ;
  assign n24912 = n21097 & ~n24911 ;
  assign n24913 = n11619 & n24912 ;
  assign n24914 = \P2_P1_lWord_reg[15]/NET0131  & ~n24913 ;
  assign n24915 = ~n24910 & ~n24914 ;
  assign n24916 = \P1_P1_lWord_reg[14]/NET0131  & ~n24515 ;
  assign n24917 = \P1_P1_lWord_reg[14]/NET0131  & ~n24506 ;
  assign n24918 = \P1_P1_EAX_reg[14]/NET0131  & n24503 ;
  assign n24919 = ~n24917 & ~n24918 ;
  assign n24920 = ~n22860 & n24919 ;
  assign n24921 = n8355 & ~n24920 ;
  assign n24922 = ~n24916 & ~n24921 ;
  assign n24923 = \P1_P1_EAX_reg[12]/NET0131  & ~n15326 ;
  assign n24924 = n7985 & n24342 ;
  assign n24925 = n15377 & ~n15398 ;
  assign n24926 = n24346 & ~n24925 ;
  assign n24927 = \P1_P1_EAX_reg[12]/NET0131  & ~n24926 ;
  assign n24928 = \P1_P1_InstQueue_reg[0][4]/NET0131  & n8291 ;
  assign n24929 = \P1_P1_InstQueue_reg[13][4]/NET0131  & n8312 ;
  assign n24930 = \P1_P1_InstQueue_reg[10][4]/NET0131  & n8305 ;
  assign n24944 = ~n24929 & ~n24930 ;
  assign n24931 = \P1_P1_InstQueue_reg[14][4]/NET0131  & n8329 ;
  assign n24932 = \P1_P1_InstQueue_reg[15][4]/NET0131  & n8327 ;
  assign n24945 = ~n24931 & ~n24932 ;
  assign n24954 = n24944 & n24945 ;
  assign n24955 = ~n24928 & n24954 ;
  assign n24943 = \P1_P1_InstQueue_reg[12][4]/NET0131  & n8303 ;
  assign n24941 = \P1_P1_InstQueue_reg[2][4]/NET0131  & n8309 ;
  assign n24942 = \P1_P1_InstQueue_reg[4][4]/NET0131  & n8314 ;
  assign n24950 = ~n24941 & ~n24942 ;
  assign n24951 = ~n24943 & n24950 ;
  assign n24937 = \P1_P1_InstQueue_reg[8][4]/NET0131  & n8316 ;
  assign n24938 = \P1_P1_InstQueue_reg[9][4]/NET0131  & n8318 ;
  assign n24948 = ~n24937 & ~n24938 ;
  assign n24939 = \P1_P1_InstQueue_reg[1][4]/NET0131  & n8321 ;
  assign n24940 = \P1_P1_InstQueue_reg[5][4]/NET0131  & n8323 ;
  assign n24949 = ~n24939 & ~n24940 ;
  assign n24952 = n24948 & n24949 ;
  assign n24933 = \P1_P1_InstQueue_reg[7][4]/NET0131  & n8307 ;
  assign n24934 = \P1_P1_InstQueue_reg[6][4]/NET0131  & n8295 ;
  assign n24946 = ~n24933 & ~n24934 ;
  assign n24935 = \P1_P1_InstQueue_reg[11][4]/NET0131  & n8325 ;
  assign n24936 = \P1_P1_InstQueue_reg[3][4]/NET0131  & n8299 ;
  assign n24947 = ~n24935 & ~n24936 ;
  assign n24953 = n24946 & n24947 ;
  assign n24956 = n24952 & n24953 ;
  assign n24957 = n24951 & n24956 ;
  assign n24958 = n24955 & n24957 ;
  assign n24959 = n22818 & ~n24958 ;
  assign n24960 = ~\P1_P1_EAX_reg[12]/NET0131  & n15377 ;
  assign n24961 = n15398 & n24960 ;
  assign n24962 = ~n24959 & ~n24961 ;
  assign n24963 = ~n24927 & n24962 ;
  assign n24964 = ~n24924 & n24963 ;
  assign n24965 = n8355 & ~n24964 ;
  assign n24966 = ~n24923 & ~n24965 ;
  assign n24967 = \P1_P1_EAX_reg[16]/NET0131  & ~n15326 ;
  assign n24970 = n8039 & n15365 ;
  assign n24969 = ~\P1_P1_EAX_reg[16]/NET0131  & ~n15365 ;
  assign n24971 = n15383 & ~n24969 ;
  assign n24972 = ~n24970 & n24971 ;
  assign n24973 = n22831 & ~n24356 ;
  assign n24974 = \P1_P1_EAX_reg[16]/NET0131  & ~n24973 ;
  assign n25007 = ~\P1_P1_EAX_reg[16]/NET0131  & n15377 ;
  assign n25008 = n15402 & n25007 ;
  assign n24968 = ~n7924 & n23947 ;
  assign n24975 = \P1_P1_InstQueue_reg[1][0]/NET0131  & n8291 ;
  assign n24976 = \P1_P1_InstQueue_reg[14][0]/NET0131  & n8312 ;
  assign n24977 = \P1_P1_InstQueue_reg[4][0]/NET0131  & n8299 ;
  assign n24991 = ~n24976 & ~n24977 ;
  assign n24978 = \P1_P1_InstQueue_reg[6][0]/NET0131  & n8323 ;
  assign n24979 = \P1_P1_InstQueue_reg[3][0]/NET0131  & n8309 ;
  assign n24992 = ~n24978 & ~n24979 ;
  assign n25001 = n24991 & n24992 ;
  assign n25002 = ~n24975 & n25001 ;
  assign n24990 = \P1_P1_InstQueue_reg[8][0]/NET0131  & n8307 ;
  assign n24988 = \P1_P1_InstQueue_reg[11][0]/NET0131  & n8305 ;
  assign n24989 = \P1_P1_InstQueue_reg[12][0]/NET0131  & n8325 ;
  assign n24997 = ~n24988 & ~n24989 ;
  assign n24998 = ~n24990 & n24997 ;
  assign n24984 = \P1_P1_InstQueue_reg[9][0]/NET0131  & n8316 ;
  assign n24985 = \P1_P1_InstQueue_reg[2][0]/NET0131  & n8321 ;
  assign n24995 = ~n24984 & ~n24985 ;
  assign n24986 = \P1_P1_InstQueue_reg[10][0]/NET0131  & n8318 ;
  assign n24987 = \P1_P1_InstQueue_reg[15][0]/NET0131  & n8329 ;
  assign n24996 = ~n24986 & ~n24987 ;
  assign n24999 = n24995 & n24996 ;
  assign n24980 = \P1_P1_InstQueue_reg[7][0]/NET0131  & n8295 ;
  assign n24981 = \P1_P1_InstQueue_reg[13][0]/NET0131  & n8303 ;
  assign n24993 = ~n24980 & ~n24981 ;
  assign n24982 = \P1_P1_InstQueue_reg[0][0]/NET0131  & n8327 ;
  assign n24983 = \P1_P1_InstQueue_reg[5][0]/NET0131  & n8314 ;
  assign n24994 = ~n24982 & ~n24983 ;
  assign n25000 = n24993 & n24994 ;
  assign n25003 = n24999 & n25000 ;
  assign n25004 = n24998 & n25003 ;
  assign n25005 = n25002 & n25004 ;
  assign n25006 = n22818 & ~n25005 ;
  assign n25009 = ~n24968 & ~n25006 ;
  assign n25010 = ~n25008 & n25009 ;
  assign n25011 = ~n24974 & n25010 ;
  assign n25012 = ~n24972 & n25011 ;
  assign n25013 = n8355 & ~n25012 ;
  assign n25014 = ~n24967 & ~n25013 ;
  assign n25015 = \P1_P1_EAX_reg[17]/NET0131  & ~n15326 ;
  assign n25053 = n8052 & n15365 ;
  assign n25052 = ~\P1_P1_EAX_reg[17]/NET0131  & ~n15365 ;
  assign n25054 = n15383 & ~n25052 ;
  assign n25055 = ~n25053 & n25054 ;
  assign n25016 = \P1_P1_EAX_reg[17]/NET0131  & ~n24567 ;
  assign n25017 = n15403 & n24566 ;
  assign n25018 = \P1_P1_InstQueue_reg[1][1]/NET0131  & n8291 ;
  assign n25019 = \P1_P1_InstQueue_reg[13][1]/NET0131  & n8303 ;
  assign n25020 = \P1_P1_InstQueue_reg[3][1]/NET0131  & n8309 ;
  assign n25034 = ~n25019 & ~n25020 ;
  assign n25021 = \P1_P1_InstQueue_reg[5][1]/NET0131  & n8314 ;
  assign n25022 = \P1_P1_InstQueue_reg[14][1]/NET0131  & n8312 ;
  assign n25035 = ~n25021 & ~n25022 ;
  assign n25044 = n25034 & n25035 ;
  assign n25045 = ~n25018 & n25044 ;
  assign n25033 = \P1_P1_InstQueue_reg[4][1]/NET0131  & n8299 ;
  assign n25031 = \P1_P1_InstQueue_reg[11][1]/NET0131  & n8305 ;
  assign n25032 = \P1_P1_InstQueue_reg[6][1]/NET0131  & n8323 ;
  assign n25040 = ~n25031 & ~n25032 ;
  assign n25041 = ~n25033 & n25040 ;
  assign n25027 = \P1_P1_InstQueue_reg[9][1]/NET0131  & n8316 ;
  assign n25028 = \P1_P1_InstQueue_reg[10][1]/NET0131  & n8318 ;
  assign n25038 = ~n25027 & ~n25028 ;
  assign n25029 = \P1_P1_InstQueue_reg[2][1]/NET0131  & n8321 ;
  assign n25030 = \P1_P1_InstQueue_reg[0][1]/NET0131  & n8327 ;
  assign n25039 = ~n25029 & ~n25030 ;
  assign n25042 = n25038 & n25039 ;
  assign n25023 = \P1_P1_InstQueue_reg[7][1]/NET0131  & n8295 ;
  assign n25024 = \P1_P1_InstQueue_reg[12][1]/NET0131  & n8325 ;
  assign n25036 = ~n25023 & ~n25024 ;
  assign n25025 = \P1_P1_InstQueue_reg[8][1]/NET0131  & n8307 ;
  assign n25026 = \P1_P1_InstQueue_reg[15][1]/NET0131  & n8329 ;
  assign n25037 = ~n25025 & ~n25026 ;
  assign n25043 = n25036 & n25037 ;
  assign n25046 = n25042 & n25043 ;
  assign n25047 = n25041 & n25046 ;
  assign n25048 = n25045 & n25047 ;
  assign n25049 = n22818 & ~n25048 ;
  assign n25050 = n7920 & n23946 ;
  assign n25051 = ~n15364 & n25050 ;
  assign n25056 = ~n25049 & ~n25051 ;
  assign n25057 = ~n25017 & n25056 ;
  assign n25058 = ~n25016 & n25057 ;
  assign n25059 = ~n25055 & n25058 ;
  assign n25060 = n8355 & ~n25059 ;
  assign n25061 = ~n25015 & ~n25060 ;
  assign n25062 = \P2_P1_EAX_reg[13]/NET0131  & ~n21100 ;
  assign n25064 = \P2_P1_EAX_reg[13]/NET0131  & ~n24713 ;
  assign n25065 = n11384 & n24708 ;
  assign n25063 = n21034 & n24710 ;
  assign n25071 = \P2_P1_InstQueue_reg[8][5]/NET0131  & n11651 ;
  assign n25070 = \P2_P1_InstQueue_reg[1][5]/NET0131  & n11647 ;
  assign n25066 = \P2_P1_InstQueue_reg[4][5]/NET0131  & n11654 ;
  assign n25067 = \P2_P1_InstQueue_reg[7][5]/NET0131  & n11638 ;
  assign n25082 = ~n25066 & ~n25067 ;
  assign n25092 = ~n25070 & n25082 ;
  assign n25093 = ~n25071 & n25092 ;
  assign n25078 = \P2_P1_InstQueue_reg[13][5]/NET0131  & n11665 ;
  assign n25079 = \P2_P1_InstQueue_reg[5][5]/NET0131  & n11663 ;
  assign n25087 = ~n25078 & ~n25079 ;
  assign n25080 = \P2_P1_InstQueue_reg[3][5]/NET0131  & n11671 ;
  assign n25081 = \P2_P1_InstQueue_reg[11][5]/NET0131  & n11656 ;
  assign n25088 = ~n25080 & ~n25081 ;
  assign n25089 = n25087 & n25088 ;
  assign n25074 = \P2_P1_InstQueue_reg[12][5]/NET0131  & n11634 ;
  assign n25075 = \P2_P1_InstQueue_reg[9][5]/NET0131  & n11661 ;
  assign n25085 = ~n25074 & ~n25075 ;
  assign n25076 = \P2_P1_InstQueue_reg[10][5]/NET0131  & n11659 ;
  assign n25077 = \P2_P1_InstQueue_reg[6][5]/NET0131  & n11667 ;
  assign n25086 = ~n25076 & ~n25077 ;
  assign n25090 = n25085 & n25086 ;
  assign n25068 = \P2_P1_InstQueue_reg[14][5]/NET0131  & n11673 ;
  assign n25069 = \P2_P1_InstQueue_reg[0][5]/NET0131  & n11643 ;
  assign n25083 = ~n25068 & ~n25069 ;
  assign n25072 = \P2_P1_InstQueue_reg[2][5]/NET0131  & n11669 ;
  assign n25073 = \P2_P1_InstQueue_reg[15][5]/NET0131  & n11641 ;
  assign n25084 = ~n25072 & ~n25073 ;
  assign n25091 = n25083 & n25084 ;
  assign n25094 = n25090 & n25091 ;
  assign n25095 = n25089 & n25094 ;
  assign n25096 = n25093 & n25095 ;
  assign n25097 = n20728 & ~n25096 ;
  assign n25098 = ~n25063 & ~n25097 ;
  assign n25099 = ~n25065 & n25098 ;
  assign n25100 = ~n25064 & n25099 ;
  assign n25101 = n11623 & ~n25100 ;
  assign n25102 = ~n25062 & ~n25101 ;
  assign n25103 = \P2_P1_EAX_reg[17]/NET0131  & ~n21100 ;
  assign n25136 = n21022 & ~n21038 ;
  assign n25137 = ~n21072 & ~n25136 ;
  assign n25138 = \P2_P1_EAX_reg[17]/NET0131  & ~n25137 ;
  assign n25146 = ~\P2_P1_EAX_reg[17]/NET0131  & n21022 ;
  assign n25147 = n21038 & n25146 ;
  assign n25139 = \P2_P1_EAX_reg[17]/NET0131  & ~n22337 ;
  assign n25143 = n11344 & n22337 ;
  assign n25144 = ~n25139 & ~n25143 ;
  assign n25145 = n21068 & ~n25144 ;
  assign n25115 = \P2_P1_InstQueue_reg[9][1]/NET0131  & n11651 ;
  assign n25108 = \P2_P1_InstQueue_reg[2][1]/NET0131  & n11647 ;
  assign n25104 = \P2_P1_InstQueue_reg[5][1]/NET0131  & n11654 ;
  assign n25105 = \P2_P1_InstQueue_reg[13][1]/NET0131  & n11634 ;
  assign n25120 = ~n25104 & ~n25105 ;
  assign n25130 = ~n25108 & n25120 ;
  assign n25131 = ~n25115 & n25130 ;
  assign n25116 = \P2_P1_InstQueue_reg[11][1]/NET0131  & n11659 ;
  assign n25117 = \P2_P1_InstQueue_reg[12][1]/NET0131  & n11656 ;
  assign n25125 = ~n25116 & ~n25117 ;
  assign n25118 = \P2_P1_InstQueue_reg[7][1]/NET0131  & n11667 ;
  assign n25119 = \P2_P1_InstQueue_reg[8][1]/NET0131  & n11638 ;
  assign n25126 = ~n25118 & ~n25119 ;
  assign n25127 = n25125 & n25126 ;
  assign n25111 = \P2_P1_InstQueue_reg[14][1]/NET0131  & n11665 ;
  assign n25112 = \P2_P1_InstQueue_reg[6][1]/NET0131  & n11663 ;
  assign n25123 = ~n25111 & ~n25112 ;
  assign n25113 = \P2_P1_InstQueue_reg[10][1]/NET0131  & n11661 ;
  assign n25114 = \P2_P1_InstQueue_reg[3][1]/NET0131  & n11669 ;
  assign n25124 = ~n25113 & ~n25114 ;
  assign n25128 = n25123 & n25124 ;
  assign n25106 = \P2_P1_InstQueue_reg[15][1]/NET0131  & n11673 ;
  assign n25107 = \P2_P1_InstQueue_reg[1][1]/NET0131  & n11643 ;
  assign n25121 = ~n25106 & ~n25107 ;
  assign n25109 = \P2_P1_InstQueue_reg[0][1]/NET0131  & n11641 ;
  assign n25110 = \P2_P1_InstQueue_reg[4][1]/NET0131  & n11671 ;
  assign n25122 = ~n25109 & ~n25110 ;
  assign n25129 = n25121 & n25122 ;
  assign n25132 = n25128 & n25129 ;
  assign n25133 = n25127 & n25132 ;
  assign n25134 = n25131 & n25133 ;
  assign n25135 = n20728 & ~n25134 ;
  assign n25140 = n11380 & n22337 ;
  assign n25141 = ~n25139 & ~n25140 ;
  assign n25142 = n21062 & ~n25141 ;
  assign n25148 = ~n25135 & ~n25142 ;
  assign n25149 = ~n25145 & n25148 ;
  assign n25150 = ~n25147 & n25149 ;
  assign n25151 = ~n25138 & n25150 ;
  assign n25152 = n11623 & ~n25151 ;
  assign n25153 = ~n25103 & ~n25152 ;
  assign n25154 = ~n21074 & ~n24902 ;
  assign n25155 = n11623 & ~n25154 ;
  assign n25156 = n24913 & ~n25155 ;
  assign n25157 = \P2_P1_lWord_reg[14]/NET0131  & ~n25156 ;
  assign n25158 = n11381 & n23167 ;
  assign n25159 = \P2_P1_EAX_reg[14]/NET0131  & n24898 ;
  assign n25160 = ~n25158 & ~n25159 ;
  assign n25161 = n11623 & ~n21081 ;
  assign n25162 = ~n25160 & n25161 ;
  assign n25163 = ~n25157 & ~n25162 ;
  assign n25164 = n8355 & ~n24506 ;
  assign n25165 = n24515 & ~n25164 ;
  assign n25166 = \P1_P1_lWord_reg[13]/NET0131  & ~n25165 ;
  assign n25167 = \P1_P1_EAX_reg[13]/NET0131  & n24503 ;
  assign n25168 = ~n8007 & n23947 ;
  assign n25169 = ~n25167 & ~n25168 ;
  assign n25170 = n8355 & ~n25169 ;
  assign n25171 = ~n25166 & ~n25170 ;
  assign n25172 = \P2_P1_EAX_reg[12]/NET0131  & ~n21100 ;
  assign n25175 = n21022 & ~n21033 ;
  assign n25176 = ~n21072 & ~n25175 ;
  assign n25177 = \P2_P1_EAX_reg[12]/NET0131  & ~n25176 ;
  assign n25210 = \P2_P1_EAX_reg[12]/NET0131  & ~n22337 ;
  assign n25211 = ~n22804 & ~n25210 ;
  assign n25212 = ~n21069 & ~n25211 ;
  assign n25173 = ~\P2_P1_EAX_reg[12]/NET0131  & n21022 ;
  assign n25174 = n21033 & n25173 ;
  assign n25183 = \P2_P1_InstQueue_reg[8][4]/NET0131  & n11651 ;
  assign n25182 = \P2_P1_InstQueue_reg[1][4]/NET0131  & n11647 ;
  assign n25178 = \P2_P1_InstQueue_reg[4][4]/NET0131  & n11654 ;
  assign n25179 = \P2_P1_InstQueue_reg[7][4]/NET0131  & n11638 ;
  assign n25194 = ~n25178 & ~n25179 ;
  assign n25204 = ~n25182 & n25194 ;
  assign n25205 = ~n25183 & n25204 ;
  assign n25190 = \P2_P1_InstQueue_reg[13][4]/NET0131  & n11665 ;
  assign n25191 = \P2_P1_InstQueue_reg[5][4]/NET0131  & n11663 ;
  assign n25199 = ~n25190 & ~n25191 ;
  assign n25192 = \P2_P1_InstQueue_reg[3][4]/NET0131  & n11671 ;
  assign n25193 = \P2_P1_InstQueue_reg[11][4]/NET0131  & n11656 ;
  assign n25200 = ~n25192 & ~n25193 ;
  assign n25201 = n25199 & n25200 ;
  assign n25186 = \P2_P1_InstQueue_reg[12][4]/NET0131  & n11634 ;
  assign n25187 = \P2_P1_InstQueue_reg[9][4]/NET0131  & n11661 ;
  assign n25197 = ~n25186 & ~n25187 ;
  assign n25188 = \P2_P1_InstQueue_reg[10][4]/NET0131  & n11659 ;
  assign n25189 = \P2_P1_InstQueue_reg[6][4]/NET0131  & n11667 ;
  assign n25198 = ~n25188 & ~n25189 ;
  assign n25202 = n25197 & n25198 ;
  assign n25180 = \P2_P1_InstQueue_reg[14][4]/NET0131  & n11673 ;
  assign n25181 = \P2_P1_InstQueue_reg[0][4]/NET0131  & n11643 ;
  assign n25195 = ~n25180 & ~n25181 ;
  assign n25184 = \P2_P1_InstQueue_reg[2][4]/NET0131  & n11669 ;
  assign n25185 = \P2_P1_InstQueue_reg[15][4]/NET0131  & n11641 ;
  assign n25196 = ~n25184 & ~n25185 ;
  assign n25203 = n25195 & n25196 ;
  assign n25206 = n25202 & n25203 ;
  assign n25207 = n25201 & n25206 ;
  assign n25208 = n25205 & n25207 ;
  assign n25209 = n20728 & ~n25208 ;
  assign n25213 = ~n25174 & ~n25209 ;
  assign n25214 = ~n25212 & n25213 ;
  assign n25215 = ~n25177 & n25214 ;
  assign n25216 = n11623 & ~n25215 ;
  assign n25217 = ~n25172 & ~n25216 ;
  assign n25250 = ~\P2_P1_EAX_reg[16]/NET0131  & ~n21037 ;
  assign n25251 = n25136 & ~n25250 ;
  assign n25252 = \P2_P1_EAX_reg[16]/NET0131  & n21072 ;
  assign n25253 = \P2_P1_EAX_reg[16]/NET0131  & ~n22337 ;
  assign n25257 = n11346 & n22337 ;
  assign n25258 = ~n25253 & ~n25257 ;
  assign n25259 = n21068 & ~n25258 ;
  assign n25223 = \P2_P1_InstQueue_reg[9][0]/NET0131  & n11651 ;
  assign n25222 = \P2_P1_InstQueue_reg[2][0]/NET0131  & n11647 ;
  assign n25218 = \P2_P1_InstQueue_reg[0][0]/NET0131  & n11641 ;
  assign n25219 = \P2_P1_InstQueue_reg[12][0]/NET0131  & n11656 ;
  assign n25234 = ~n25218 & ~n25219 ;
  assign n25244 = ~n25222 & n25234 ;
  assign n25245 = ~n25223 & n25244 ;
  assign n25230 = \P2_P1_InstQueue_reg[6][0]/NET0131  & n11663 ;
  assign n25231 = \P2_P1_InstQueue_reg[13][0]/NET0131  & n11634 ;
  assign n25239 = ~n25230 & ~n25231 ;
  assign n25232 = \P2_P1_InstQueue_reg[11][0]/NET0131  & n11659 ;
  assign n25233 = \P2_P1_InstQueue_reg[4][0]/NET0131  & n11671 ;
  assign n25240 = ~n25232 & ~n25233 ;
  assign n25241 = n25239 & n25240 ;
  assign n25226 = \P2_P1_InstQueue_reg[5][0]/NET0131  & n11654 ;
  assign n25227 = \P2_P1_InstQueue_reg[10][0]/NET0131  & n11661 ;
  assign n25237 = ~n25226 & ~n25227 ;
  assign n25228 = \P2_P1_InstQueue_reg[14][0]/NET0131  & n11665 ;
  assign n25229 = \P2_P1_InstQueue_reg[8][0]/NET0131  & n11638 ;
  assign n25238 = ~n25228 & ~n25229 ;
  assign n25242 = n25237 & n25238 ;
  assign n25220 = \P2_P1_InstQueue_reg[3][0]/NET0131  & n11669 ;
  assign n25221 = \P2_P1_InstQueue_reg[1][0]/NET0131  & n11643 ;
  assign n25235 = ~n25220 & ~n25221 ;
  assign n25224 = \P2_P1_InstQueue_reg[15][0]/NET0131  & n11673 ;
  assign n25225 = \P2_P1_InstQueue_reg[7][0]/NET0131  & n11667 ;
  assign n25236 = ~n25224 & ~n25225 ;
  assign n25243 = n25235 & n25236 ;
  assign n25246 = n25242 & n25243 ;
  assign n25247 = n25241 & n25246 ;
  assign n25248 = n25245 & n25247 ;
  assign n25249 = n20728 & ~n25248 ;
  assign n25254 = n11379 & n22337 ;
  assign n25255 = ~n25253 & ~n25254 ;
  assign n25256 = n21062 & ~n25255 ;
  assign n25260 = ~n25249 & ~n25256 ;
  assign n25261 = ~n25259 & n25260 ;
  assign n25262 = ~n25252 & n25261 ;
  assign n25263 = ~n25251 & n25262 ;
  assign n25264 = n11623 & ~n25263 ;
  assign n25265 = \P2_P1_EAX_reg[16]/NET0131  & ~n21100 ;
  assign n25266 = ~n25264 & ~n25265 ;
  assign n25267 = \P2_P1_lWord_reg[13]/NET0131  & ~n25156 ;
  assign n25268 = \P2_P1_EAX_reg[13]/NET0131  & n24898 ;
  assign n25269 = ~n23168 & ~n25268 ;
  assign n25270 = n25161 & ~n25269 ;
  assign n25271 = ~n25267 & ~n25270 ;
  assign n25272 = \P1_P1_lWord_reg[12]/NET0131  & ~n24515 ;
  assign n25274 = \P1_P1_lWord_reg[12]/NET0131  & n15335 ;
  assign n25275 = ~n22834 & ~n25274 ;
  assign n25276 = n15334 & ~n25275 ;
  assign n25273 = \P1_P1_EAX_reg[12]/NET0131  & n24503 ;
  assign n25277 = \P1_P1_lWord_reg[12]/NET0131  & n24505 ;
  assign n25278 = ~n25273 & ~n25277 ;
  assign n25279 = ~n25276 & n25278 ;
  assign n25280 = n8355 & ~n25279 ;
  assign n25281 = ~n25272 & ~n25280 ;
  assign n25282 = \P2_P1_lWord_reg[12]/NET0131  & ~n25156 ;
  assign n25283 = n11375 & n23167 ;
  assign n25284 = \P2_P1_EAX_reg[12]/NET0131  & n24898 ;
  assign n25285 = ~n25283 & ~n25284 ;
  assign n25286 = n25161 & ~n25285 ;
  assign n25287 = ~n25282 & ~n25286 ;
  assign n25288 = \P1_P1_EAX_reg[11]/NET0131  & ~n15326 ;
  assign n25289 = ~n15384 & n23970 ;
  assign n25290 = n15377 & ~n15397 ;
  assign n25291 = n24346 & ~n25290 ;
  assign n25292 = \P1_P1_EAX_reg[11]/NET0131  & ~n25291 ;
  assign n25293 = \P1_P1_InstQueue_reg[0][3]/NET0131  & n8291 ;
  assign n25294 = \P1_P1_InstQueue_reg[5][3]/NET0131  & n8323 ;
  assign n25295 = \P1_P1_InstQueue_reg[15][3]/NET0131  & n8327 ;
  assign n25309 = ~n25294 & ~n25295 ;
  assign n25296 = \P1_P1_InstQueue_reg[14][3]/NET0131  & n8329 ;
  assign n25297 = \P1_P1_InstQueue_reg[13][3]/NET0131  & n8312 ;
  assign n25310 = ~n25296 & ~n25297 ;
  assign n25319 = n25309 & n25310 ;
  assign n25320 = ~n25293 & n25319 ;
  assign n25308 = \P1_P1_InstQueue_reg[11][3]/NET0131  & n8325 ;
  assign n25306 = \P1_P1_InstQueue_reg[3][3]/NET0131  & n8299 ;
  assign n25307 = \P1_P1_InstQueue_reg[10][3]/NET0131  & n8305 ;
  assign n25315 = ~n25306 & ~n25307 ;
  assign n25316 = ~n25308 & n25315 ;
  assign n25302 = \P1_P1_InstQueue_reg[8][3]/NET0131  & n8316 ;
  assign n25303 = \P1_P1_InstQueue_reg[9][3]/NET0131  & n8318 ;
  assign n25313 = ~n25302 & ~n25303 ;
  assign n25304 = \P1_P1_InstQueue_reg[1][3]/NET0131  & n8321 ;
  assign n25305 = \P1_P1_InstQueue_reg[2][3]/NET0131  & n8309 ;
  assign n25314 = ~n25304 & ~n25305 ;
  assign n25317 = n25313 & n25314 ;
  assign n25298 = \P1_P1_InstQueue_reg[12][3]/NET0131  & n8303 ;
  assign n25299 = \P1_P1_InstQueue_reg[7][3]/NET0131  & n8307 ;
  assign n25311 = ~n25298 & ~n25299 ;
  assign n25300 = \P1_P1_InstQueue_reg[4][3]/NET0131  & n8314 ;
  assign n25301 = \P1_P1_InstQueue_reg[6][3]/NET0131  & n8295 ;
  assign n25312 = ~n25300 & ~n25301 ;
  assign n25318 = n25311 & n25312 ;
  assign n25321 = n25317 & n25318 ;
  assign n25322 = n25316 & n25321 ;
  assign n25323 = n25320 & n25322 ;
  assign n25324 = n22818 & ~n25323 ;
  assign n25325 = n15397 & n24925 ;
  assign n25326 = ~n25324 & ~n25325 ;
  assign n25327 = ~n25292 & n25326 ;
  assign n25328 = ~n25289 & n25327 ;
  assign n25329 = n8355 & ~n25328 ;
  assign n25330 = ~n25288 & ~n25329 ;
  assign n25331 = \P1_P1_uWord_reg[14]/NET0131  & ~n24515 ;
  assign n25363 = n15335 & ~n15364 ;
  assign n25364 = \P1_P1_uWord_reg[14]/NET0131  & n25363 ;
  assign n25365 = ~n22859 & ~n25364 ;
  assign n25366 = n15334 & ~n25365 ;
  assign n25334 = ~\P1_P1_EAX_reg[13]/NET0131  & ~\P1_P1_EAX_reg[14]/NET0131  ;
  assign n25335 = ~\P1_P1_EAX_reg[15]/NET0131  & ~\P1_P1_EAX_reg[1]/NET0131  ;
  assign n25342 = n25334 & n25335 ;
  assign n25332 = ~\P1_P1_EAX_reg[0]/NET0131  & ~\P1_P1_EAX_reg[10]/NET0131  ;
  assign n25333 = ~\P1_P1_EAX_reg[11]/NET0131  & ~\P1_P1_EAX_reg[12]/NET0131  ;
  assign n25343 = n25332 & n25333 ;
  assign n25344 = n25342 & n25343 ;
  assign n25338 = ~\P1_P1_EAX_reg[6]/NET0131  & ~\P1_P1_EAX_reg[7]/NET0131  ;
  assign n25339 = ~\P1_P1_EAX_reg[8]/NET0131  & ~\P1_P1_EAX_reg[9]/NET0131  ;
  assign n25340 = n25338 & n25339 ;
  assign n25336 = ~\P1_P1_EAX_reg[2]/NET0131  & ~\P1_P1_EAX_reg[3]/NET0131  ;
  assign n25337 = ~\P1_P1_EAX_reg[4]/NET0131  & ~\P1_P1_EAX_reg[5]/NET0131  ;
  assign n25341 = n25336 & n25337 ;
  assign n25345 = n25340 & n25341 ;
  assign n25346 = n25344 & n25345 ;
  assign n25347 = \P1_P1_EAX_reg[31]/NET0131  & ~n25346 ;
  assign n25348 = \P1_P1_EAX_reg[16]/NET0131  & n25347 ;
  assign n25349 = \P1_P1_EAX_reg[17]/NET0131  & n25348 ;
  assign n25350 = \P1_P1_EAX_reg[18]/NET0131  & n25349 ;
  assign n25351 = \P1_P1_EAX_reg[19]/NET0131  & n25350 ;
  assign n25352 = \P1_P1_EAX_reg[20]/NET0131  & n25351 ;
  assign n25353 = \P1_P1_EAX_reg[21]/NET0131  & n25352 ;
  assign n25354 = \P1_P1_EAX_reg[22]/NET0131  & n25353 ;
  assign n25355 = \P1_P1_EAX_reg[23]/NET0131  & n25354 ;
  assign n25356 = n22820 & n25355 ;
  assign n25357 = n15412 & n25356 ;
  assign n25358 = n22848 & n25357 ;
  assign n25360 = \P1_P1_EAX_reg[30]/NET0131  & n25358 ;
  assign n25359 = ~\P1_P1_EAX_reg[30]/NET0131  & ~n25358 ;
  assign n25361 = n24503 & ~n25359 ;
  assign n25362 = ~n25360 & n25361 ;
  assign n25367 = \P1_P1_uWord_reg[14]/NET0131  & n24505 ;
  assign n25368 = ~n25362 & ~n25367 ;
  assign n25369 = ~n25366 & n25368 ;
  assign n25370 = n8355 & ~n25369 ;
  assign n25371 = ~n25331 & ~n25370 ;
  assign n25372 = \P2_P1_EAX_reg[11]/NET0131  & ~n21100 ;
  assign n25374 = \P2_P1_EAX_reg[11]/NET0131  & ~n25176 ;
  assign n25407 = \P2_P1_EAX_reg[11]/NET0131  & ~n22337 ;
  assign n25408 = ~n23863 & ~n25407 ;
  assign n25409 = ~n21069 & ~n25408 ;
  assign n25373 = n21032 & n25175 ;
  assign n25380 = \P2_P1_InstQueue_reg[8][3]/NET0131  & n11651 ;
  assign n25379 = \P2_P1_InstQueue_reg[1][3]/NET0131  & n11647 ;
  assign n25375 = \P2_P1_InstQueue_reg[7][3]/NET0131  & n11638 ;
  assign n25376 = \P2_P1_InstQueue_reg[4][3]/NET0131  & n11654 ;
  assign n25391 = ~n25375 & ~n25376 ;
  assign n25401 = ~n25379 & n25391 ;
  assign n25402 = ~n25380 & n25401 ;
  assign n25387 = \P2_P1_InstQueue_reg[3][3]/NET0131  & n11671 ;
  assign n25388 = \P2_P1_InstQueue_reg[6][3]/NET0131  & n11667 ;
  assign n25396 = ~n25387 & ~n25388 ;
  assign n25389 = \P2_P1_InstQueue_reg[12][3]/NET0131  & n11634 ;
  assign n25390 = \P2_P1_InstQueue_reg[15][3]/NET0131  & n11641 ;
  assign n25397 = ~n25389 & ~n25390 ;
  assign n25398 = n25396 & n25397 ;
  assign n25383 = \P2_P1_InstQueue_reg[2][3]/NET0131  & n11669 ;
  assign n25384 = \P2_P1_InstQueue_reg[9][3]/NET0131  & n11661 ;
  assign n25394 = ~n25383 & ~n25384 ;
  assign n25385 = \P2_P1_InstQueue_reg[10][3]/NET0131  & n11659 ;
  assign n25386 = \P2_P1_InstQueue_reg[13][3]/NET0131  & n11665 ;
  assign n25395 = ~n25385 & ~n25386 ;
  assign n25399 = n25394 & n25395 ;
  assign n25377 = \P2_P1_InstQueue_reg[11][3]/NET0131  & n11656 ;
  assign n25378 = \P2_P1_InstQueue_reg[0][3]/NET0131  & n11643 ;
  assign n25392 = ~n25377 & ~n25378 ;
  assign n25381 = \P2_P1_InstQueue_reg[5][3]/NET0131  & n11663 ;
  assign n25382 = \P2_P1_InstQueue_reg[14][3]/NET0131  & n11673 ;
  assign n25393 = ~n25381 & ~n25382 ;
  assign n25400 = n25392 & n25393 ;
  assign n25403 = n25399 & n25400 ;
  assign n25404 = n25398 & n25403 ;
  assign n25405 = n25402 & n25404 ;
  assign n25406 = n20728 & ~n25405 ;
  assign n25410 = ~n25373 & ~n25406 ;
  assign n25411 = ~n25409 & n25410 ;
  assign n25412 = ~n25374 & n25411 ;
  assign n25413 = n11623 & ~n25412 ;
  assign n25414 = ~n25372 & ~n25413 ;
  assign n25451 = \P1_P2_InstQueueRd_Addr_reg[1]/NET0131  & \P1_P2_InstQueueRd_Addr_reg[2]/NET0131  ;
  assign n25452 = ~\P1_P2_InstQueueRd_Addr_reg[3]/NET0131  & n25451 ;
  assign n25453 = ~\P1_P2_InstQueueRd_Addr_reg[0]/NET0131  & n25452 ;
  assign n25454 = \P1_P2_InstQueue_reg[6][5]/NET0131  & n25453 ;
  assign n25433 = \P1_P2_InstQueueRd_Addr_reg[0]/NET0131  & \P1_P2_InstQueueRd_Addr_reg[1]/NET0131  ;
  assign n25434 = \P1_P2_InstQueueRd_Addr_reg[2]/NET0131  & n25433 ;
  assign n25435 = ~\P1_P2_InstQueueRd_Addr_reg[3]/NET0131  & n25434 ;
  assign n25436 = \P1_P2_InstQueue_reg[7][5]/NET0131  & n25435 ;
  assign n25420 = \P1_P2_InstQueueRd_Addr_reg[2]/NET0131  & \P1_P2_InstQueueRd_Addr_reg[3]/NET0131  ;
  assign n25421 = ~\P1_P2_InstQueueRd_Addr_reg[0]/NET0131  & ~\P1_P2_InstQueueRd_Addr_reg[1]/NET0131  ;
  assign n25422 = n25420 & n25421 ;
  assign n25423 = \P1_P2_InstQueue_reg[12][5]/NET0131  & n25422 ;
  assign n25424 = ~\P1_P2_InstQueueRd_Addr_reg[2]/NET0131  & ~\P1_P2_InstQueueRd_Addr_reg[3]/NET0131  ;
  assign n25425 = n25421 & n25424 ;
  assign n25426 = \P1_P2_InstQueue_reg[0][5]/NET0131  & n25425 ;
  assign n25463 = ~n25423 & ~n25426 ;
  assign n25473 = ~n25436 & n25463 ;
  assign n25474 = ~n25454 & n25473 ;
  assign n25439 = ~\P1_P2_InstQueueRd_Addr_reg[2]/NET0131  & \P1_P2_InstQueueRd_Addr_reg[3]/NET0131  ;
  assign n25455 = n25421 & n25439 ;
  assign n25456 = \P1_P2_InstQueue_reg[8][5]/NET0131  & n25455 ;
  assign n25427 = \P1_P2_InstQueueRd_Addr_reg[0]/NET0131  & ~\P1_P2_InstQueueRd_Addr_reg[1]/NET0131  ;
  assign n25457 = n25427 & n25439 ;
  assign n25458 = \P1_P2_InstQueue_reg[9][5]/NET0131  & n25457 ;
  assign n25468 = ~n25456 & ~n25458 ;
  assign n25459 = n25433 & n25439 ;
  assign n25460 = \P1_P2_InstQueue_reg[11][5]/NET0131  & n25459 ;
  assign n25448 = \P1_P2_InstQueueRd_Addr_reg[2]/NET0131  & ~\P1_P2_InstQueueRd_Addr_reg[3]/NET0131  ;
  assign n25461 = n25421 & n25448 ;
  assign n25462 = \P1_P2_InstQueue_reg[4][5]/NET0131  & n25461 ;
  assign n25469 = ~n25460 & ~n25462 ;
  assign n25470 = n25468 & n25469 ;
  assign n25442 = n25420 & n25427 ;
  assign n25443 = \P1_P2_InstQueue_reg[13][5]/NET0131  & n25442 ;
  assign n25430 = ~\P1_P2_InstQueueRd_Addr_reg[0]/NET0131  & \P1_P2_InstQueueRd_Addr_reg[1]/NET0131  ;
  assign n25444 = n25424 & n25430 ;
  assign n25445 = \P1_P2_InstQueue_reg[2][5]/NET0131  & n25444 ;
  assign n25466 = ~n25443 & ~n25445 ;
  assign n25446 = n25420 & n25433 ;
  assign n25447 = \P1_P2_InstQueue_reg[15][5]/NET0131  & n25446 ;
  assign n25449 = n25427 & n25448 ;
  assign n25450 = \P1_P2_InstQueue_reg[5][5]/NET0131  & n25449 ;
  assign n25467 = ~n25447 & ~n25450 ;
  assign n25471 = n25466 & n25467 ;
  assign n25428 = n25424 & n25427 ;
  assign n25429 = \P1_P2_InstQueue_reg[1][5]/NET0131  & n25428 ;
  assign n25431 = n25420 & n25430 ;
  assign n25432 = \P1_P2_InstQueue_reg[14][5]/NET0131  & n25431 ;
  assign n25464 = ~n25429 & ~n25432 ;
  assign n25437 = n25424 & n25433 ;
  assign n25438 = \P1_P2_InstQueue_reg[3][5]/NET0131  & n25437 ;
  assign n25440 = n25430 & n25439 ;
  assign n25441 = \P1_P2_InstQueue_reg[10][5]/NET0131  & n25440 ;
  assign n25465 = ~n25438 & ~n25441 ;
  assign n25472 = n25464 & n25465 ;
  assign n25475 = n25471 & n25472 ;
  assign n25476 = n25470 & n25475 ;
  assign n25477 = n25474 & n25476 ;
  assign n25489 = \P1_P2_InstQueue_reg[6][4]/NET0131  & n25453 ;
  assign n25482 = \P1_P2_InstQueue_reg[7][4]/NET0131  & n25435 ;
  assign n25478 = \P1_P2_InstQueue_reg[0][4]/NET0131  & n25425 ;
  assign n25479 = \P1_P2_InstQueue_reg[8][4]/NET0131  & n25455 ;
  assign n25494 = ~n25478 & ~n25479 ;
  assign n25504 = ~n25482 & n25494 ;
  assign n25505 = ~n25489 & n25504 ;
  assign n25490 = \P1_P2_InstQueue_reg[1][4]/NET0131  & n25428 ;
  assign n25491 = \P1_P2_InstQueue_reg[2][4]/NET0131  & n25444 ;
  assign n25499 = ~n25490 & ~n25491 ;
  assign n25492 = \P1_P2_InstQueue_reg[10][4]/NET0131  & n25440 ;
  assign n25493 = \P1_P2_InstQueue_reg[13][4]/NET0131  & n25442 ;
  assign n25500 = ~n25492 & ~n25493 ;
  assign n25501 = n25499 & n25500 ;
  assign n25485 = \P1_P2_InstQueue_reg[12][4]/NET0131  & n25422 ;
  assign n25486 = \P1_P2_InstQueue_reg[3][4]/NET0131  & n25437 ;
  assign n25497 = ~n25485 & ~n25486 ;
  assign n25487 = \P1_P2_InstQueue_reg[15][4]/NET0131  & n25446 ;
  assign n25488 = \P1_P2_InstQueue_reg[5][4]/NET0131  & n25449 ;
  assign n25498 = ~n25487 & ~n25488 ;
  assign n25502 = n25497 & n25498 ;
  assign n25480 = \P1_P2_InstQueue_reg[4][4]/NET0131  & n25461 ;
  assign n25481 = \P1_P2_InstQueue_reg[14][4]/NET0131  & n25431 ;
  assign n25495 = ~n25480 & ~n25481 ;
  assign n25483 = \P1_P2_InstQueue_reg[9][4]/NET0131  & n25457 ;
  assign n25484 = \P1_P2_InstQueue_reg[11][4]/NET0131  & n25459 ;
  assign n25496 = ~n25483 & ~n25484 ;
  assign n25503 = n25495 & n25496 ;
  assign n25506 = n25502 & n25503 ;
  assign n25507 = n25501 & n25506 ;
  assign n25508 = n25505 & n25507 ;
  assign n25509 = ~n25477 & n25508 ;
  assign n25521 = \P1_P2_InstQueue_reg[6][7]/NET0131  & n25453 ;
  assign n25514 = \P1_P2_InstQueue_reg[7][7]/NET0131  & n25435 ;
  assign n25510 = \P1_P2_InstQueue_reg[0][7]/NET0131  & n25425 ;
  assign n25511 = \P1_P2_InstQueue_reg[10][7]/NET0131  & n25440 ;
  assign n25526 = ~n25510 & ~n25511 ;
  assign n25536 = ~n25514 & n25526 ;
  assign n25537 = ~n25521 & n25536 ;
  assign n25522 = \P1_P2_InstQueue_reg[9][7]/NET0131  & n25457 ;
  assign n25523 = \P1_P2_InstQueue_reg[12][7]/NET0131  & n25422 ;
  assign n25531 = ~n25522 & ~n25523 ;
  assign n25524 = \P1_P2_InstQueue_reg[13][7]/NET0131  & n25442 ;
  assign n25525 = \P1_P2_InstQueue_reg[5][7]/NET0131  & n25449 ;
  assign n25532 = ~n25524 & ~n25525 ;
  assign n25533 = n25531 & n25532 ;
  assign n25517 = \P1_P2_InstQueue_reg[8][7]/NET0131  & n25455 ;
  assign n25518 = \P1_P2_InstQueue_reg[4][7]/NET0131  & n25461 ;
  assign n25529 = ~n25517 & ~n25518 ;
  assign n25519 = \P1_P2_InstQueue_reg[15][7]/NET0131  & n25446 ;
  assign n25520 = \P1_P2_InstQueue_reg[2][7]/NET0131  & n25444 ;
  assign n25530 = ~n25519 & ~n25520 ;
  assign n25534 = n25529 & n25530 ;
  assign n25512 = \P1_P2_InstQueue_reg[1][7]/NET0131  & n25428 ;
  assign n25513 = \P1_P2_InstQueue_reg[14][7]/NET0131  & n25431 ;
  assign n25527 = ~n25512 & ~n25513 ;
  assign n25515 = \P1_P2_InstQueue_reg[3][7]/NET0131  & n25437 ;
  assign n25516 = \P1_P2_InstQueue_reg[11][7]/NET0131  & n25459 ;
  assign n25528 = ~n25515 & ~n25516 ;
  assign n25535 = n25527 & n25528 ;
  assign n25538 = n25534 & n25535 ;
  assign n25539 = n25533 & n25538 ;
  assign n25540 = n25537 & n25539 ;
  assign n25552 = \P1_P2_InstQueue_reg[6][6]/NET0131  & n25453 ;
  assign n25545 = \P1_P2_InstQueue_reg[7][6]/NET0131  & n25435 ;
  assign n25541 = \P1_P2_InstQueue_reg[13][6]/NET0131  & n25442 ;
  assign n25542 = \P1_P2_InstQueue_reg[8][6]/NET0131  & n25455 ;
  assign n25557 = ~n25541 & ~n25542 ;
  assign n25567 = ~n25545 & n25557 ;
  assign n25568 = ~n25552 & n25567 ;
  assign n25553 = \P1_P2_InstQueue_reg[9][6]/NET0131  & n25457 ;
  assign n25554 = \P1_P2_InstQueue_reg[5][6]/NET0131  & n25449 ;
  assign n25562 = ~n25553 & ~n25554 ;
  assign n25555 = \P1_P2_InstQueue_reg[10][6]/NET0131  & n25440 ;
  assign n25556 = \P1_P2_InstQueue_reg[1][6]/NET0131  & n25428 ;
  assign n25563 = ~n25555 & ~n25556 ;
  assign n25564 = n25562 & n25563 ;
  assign n25548 = \P1_P2_InstQueue_reg[2][6]/NET0131  & n25444 ;
  assign n25549 = \P1_P2_InstQueue_reg[11][6]/NET0131  & n25459 ;
  assign n25560 = ~n25548 & ~n25549 ;
  assign n25550 = \P1_P2_InstQueue_reg[15][6]/NET0131  & n25446 ;
  assign n25551 = \P1_P2_InstQueue_reg[12][6]/NET0131  & n25422 ;
  assign n25561 = ~n25550 & ~n25551 ;
  assign n25565 = n25560 & n25561 ;
  assign n25543 = \P1_P2_InstQueue_reg[0][6]/NET0131  & n25425 ;
  assign n25544 = \P1_P2_InstQueue_reg[14][6]/NET0131  & n25431 ;
  assign n25558 = ~n25543 & ~n25544 ;
  assign n25546 = \P1_P2_InstQueue_reg[4][6]/NET0131  & n25461 ;
  assign n25547 = \P1_P2_InstQueue_reg[3][6]/NET0131  & n25437 ;
  assign n25559 = ~n25546 & ~n25547 ;
  assign n25566 = n25558 & n25559 ;
  assign n25569 = n25565 & n25566 ;
  assign n25570 = n25564 & n25569 ;
  assign n25571 = n25568 & n25570 ;
  assign n25572 = ~n25540 & ~n25571 ;
  assign n25573 = n25509 & n25572 ;
  assign n25585 = \P1_P2_InstQueue_reg[6][2]/NET0131  & n25453 ;
  assign n25578 = \P1_P2_InstQueue_reg[7][2]/NET0131  & n25435 ;
  assign n25574 = \P1_P2_InstQueue_reg[0][2]/NET0131  & n25425 ;
  assign n25575 = \P1_P2_InstQueue_reg[2][2]/NET0131  & n25444 ;
  assign n25590 = ~n25574 & ~n25575 ;
  assign n25600 = ~n25578 & n25590 ;
  assign n25601 = ~n25585 & n25600 ;
  assign n25586 = \P1_P2_InstQueue_reg[12][2]/NET0131  & n25422 ;
  assign n25587 = \P1_P2_InstQueue_reg[1][2]/NET0131  & n25428 ;
  assign n25595 = ~n25586 & ~n25587 ;
  assign n25588 = \P1_P2_InstQueue_reg[10][2]/NET0131  & n25440 ;
  assign n25589 = \P1_P2_InstQueue_reg[13][2]/NET0131  & n25442 ;
  assign n25596 = ~n25588 & ~n25589 ;
  assign n25597 = n25595 & n25596 ;
  assign n25581 = \P1_P2_InstQueue_reg[5][2]/NET0131  & n25449 ;
  assign n25582 = \P1_P2_InstQueue_reg[3][2]/NET0131  & n25437 ;
  assign n25593 = ~n25581 & ~n25582 ;
  assign n25583 = \P1_P2_InstQueue_reg[15][2]/NET0131  & n25446 ;
  assign n25584 = \P1_P2_InstQueue_reg[8][2]/NET0131  & n25455 ;
  assign n25594 = ~n25583 & ~n25584 ;
  assign n25598 = n25593 & n25594 ;
  assign n25576 = \P1_P2_InstQueue_reg[4][2]/NET0131  & n25461 ;
  assign n25577 = \P1_P2_InstQueue_reg[14][2]/NET0131  & n25431 ;
  assign n25591 = ~n25576 & ~n25577 ;
  assign n25579 = \P1_P2_InstQueue_reg[9][2]/NET0131  & n25457 ;
  assign n25580 = \P1_P2_InstQueue_reg[11][2]/NET0131  & n25459 ;
  assign n25592 = ~n25579 & ~n25580 ;
  assign n25599 = n25591 & n25592 ;
  assign n25602 = n25598 & n25599 ;
  assign n25603 = n25597 & n25602 ;
  assign n25604 = n25601 & n25603 ;
  assign n25616 = \P1_P2_InstQueue_reg[6][1]/NET0131  & n25453 ;
  assign n25609 = \P1_P2_InstQueue_reg[7][1]/NET0131  & n25435 ;
  assign n25605 = \P1_P2_InstQueue_reg[0][1]/NET0131  & n25425 ;
  assign n25606 = \P1_P2_InstQueue_reg[2][1]/NET0131  & n25444 ;
  assign n25621 = ~n25605 & ~n25606 ;
  assign n25631 = ~n25609 & n25621 ;
  assign n25632 = ~n25616 & n25631 ;
  assign n25617 = \P1_P2_InstQueue_reg[12][1]/NET0131  & n25422 ;
  assign n25618 = \P1_P2_InstQueue_reg[1][1]/NET0131  & n25428 ;
  assign n25626 = ~n25617 & ~n25618 ;
  assign n25619 = \P1_P2_InstQueue_reg[10][1]/NET0131  & n25440 ;
  assign n25620 = \P1_P2_InstQueue_reg[13][1]/NET0131  & n25442 ;
  assign n25627 = ~n25619 & ~n25620 ;
  assign n25628 = n25626 & n25627 ;
  assign n25612 = \P1_P2_InstQueue_reg[5][1]/NET0131  & n25449 ;
  assign n25613 = \P1_P2_InstQueue_reg[3][1]/NET0131  & n25437 ;
  assign n25624 = ~n25612 & ~n25613 ;
  assign n25614 = \P1_P2_InstQueue_reg[15][1]/NET0131  & n25446 ;
  assign n25615 = \P1_P2_InstQueue_reg[8][1]/NET0131  & n25455 ;
  assign n25625 = ~n25614 & ~n25615 ;
  assign n25629 = n25624 & n25625 ;
  assign n25607 = \P1_P2_InstQueue_reg[4][1]/NET0131  & n25461 ;
  assign n25608 = \P1_P2_InstQueue_reg[14][1]/NET0131  & n25431 ;
  assign n25622 = ~n25607 & ~n25608 ;
  assign n25610 = \P1_P2_InstQueue_reg[9][1]/NET0131  & n25457 ;
  assign n25611 = \P1_P2_InstQueue_reg[11][1]/NET0131  & n25459 ;
  assign n25623 = ~n25610 & ~n25611 ;
  assign n25630 = n25622 & n25623 ;
  assign n25633 = n25629 & n25630 ;
  assign n25634 = n25628 & n25633 ;
  assign n25635 = n25632 & n25634 ;
  assign n25636 = n25604 & ~n25635 ;
  assign n25648 = \P1_P2_InstQueue_reg[6][0]/NET0131  & n25453 ;
  assign n25641 = \P1_P2_InstQueue_reg[7][0]/NET0131  & n25435 ;
  assign n25637 = \P1_P2_InstQueue_reg[2][0]/NET0131  & n25444 ;
  assign n25638 = \P1_P2_InstQueue_reg[10][0]/NET0131  & n25440 ;
  assign n25653 = ~n25637 & ~n25638 ;
  assign n25663 = ~n25641 & n25653 ;
  assign n25664 = ~n25648 & n25663 ;
  assign n25649 = \P1_P2_InstQueue_reg[5][0]/NET0131  & n25449 ;
  assign n25650 = \P1_P2_InstQueue_reg[9][0]/NET0131  & n25457 ;
  assign n25658 = ~n25649 & ~n25650 ;
  assign n25651 = \P1_P2_InstQueue_reg[11][0]/NET0131  & n25459 ;
  assign n25652 = \P1_P2_InstQueue_reg[4][0]/NET0131  & n25461 ;
  assign n25659 = ~n25651 & ~n25652 ;
  assign n25660 = n25658 & n25659 ;
  assign n25644 = \P1_P2_InstQueue_reg[0][0]/NET0131  & n25425 ;
  assign n25645 = \P1_P2_InstQueue_reg[12][0]/NET0131  & n25422 ;
  assign n25656 = ~n25644 & ~n25645 ;
  assign n25646 = \P1_P2_InstQueue_reg[15][0]/NET0131  & n25446 ;
  assign n25647 = \P1_P2_InstQueue_reg[8][0]/NET0131  & n25455 ;
  assign n25657 = ~n25646 & ~n25647 ;
  assign n25661 = n25656 & n25657 ;
  assign n25639 = \P1_P2_InstQueue_reg[1][0]/NET0131  & n25428 ;
  assign n25640 = \P1_P2_InstQueue_reg[14][0]/NET0131  & n25431 ;
  assign n25654 = ~n25639 & ~n25640 ;
  assign n25642 = \P1_P2_InstQueue_reg[3][0]/NET0131  & n25437 ;
  assign n25643 = \P1_P2_InstQueue_reg[13][0]/NET0131  & n25442 ;
  assign n25655 = ~n25642 & ~n25643 ;
  assign n25662 = n25654 & n25655 ;
  assign n25665 = n25661 & n25662 ;
  assign n25666 = n25660 & n25665 ;
  assign n25667 = n25664 & n25666 ;
  assign n25668 = n25636 & ~n25667 ;
  assign n25680 = \P1_P2_InstQueue_reg[6][3]/NET0131  & n25453 ;
  assign n25673 = \P1_P2_InstQueue_reg[7][3]/NET0131  & n25435 ;
  assign n25669 = \P1_P2_InstQueue_reg[0][3]/NET0131  & n25425 ;
  assign n25670 = \P1_P2_InstQueue_reg[2][3]/NET0131  & n25444 ;
  assign n25685 = ~n25669 & ~n25670 ;
  assign n25695 = ~n25673 & n25685 ;
  assign n25696 = ~n25680 & n25695 ;
  assign n25681 = \P1_P2_InstQueue_reg[1][3]/NET0131  & n25428 ;
  assign n25682 = \P1_P2_InstQueue_reg[12][3]/NET0131  & n25422 ;
  assign n25690 = ~n25681 & ~n25682 ;
  assign n25683 = \P1_P2_InstQueue_reg[10][3]/NET0131  & n25440 ;
  assign n25684 = \P1_P2_InstQueue_reg[13][3]/NET0131  & n25442 ;
  assign n25691 = ~n25683 & ~n25684 ;
  assign n25692 = n25690 & n25691 ;
  assign n25676 = \P1_P2_InstQueue_reg[5][3]/NET0131  & n25449 ;
  assign n25677 = \P1_P2_InstQueue_reg[11][3]/NET0131  & n25459 ;
  assign n25688 = ~n25676 & ~n25677 ;
  assign n25678 = \P1_P2_InstQueue_reg[15][3]/NET0131  & n25446 ;
  assign n25679 = \P1_P2_InstQueue_reg[8][3]/NET0131  & n25455 ;
  assign n25689 = ~n25678 & ~n25679 ;
  assign n25693 = n25688 & n25689 ;
  assign n25671 = \P1_P2_InstQueue_reg[4][3]/NET0131  & n25461 ;
  assign n25672 = \P1_P2_InstQueue_reg[14][3]/NET0131  & n25431 ;
  assign n25686 = ~n25671 & ~n25672 ;
  assign n25674 = \P1_P2_InstQueue_reg[9][3]/NET0131  & n25457 ;
  assign n25675 = \P1_P2_InstQueue_reg[3][3]/NET0131  & n25437 ;
  assign n25687 = ~n25674 & ~n25675 ;
  assign n25694 = n25686 & n25687 ;
  assign n25697 = n25693 & n25694 ;
  assign n25698 = n25692 & n25697 ;
  assign n25699 = n25696 & n25698 ;
  assign n25700 = n25668 & ~n25699 ;
  assign n25701 = n25573 & n25700 ;
  assign n25740 = n25604 & n25635 ;
  assign n25749 = ~n25667 & ~n25699 ;
  assign n25750 = n25740 & n25749 ;
  assign n25751 = n25573 & n25750 ;
  assign n25784 = ~n25701 & ~n25751 ;
  assign n25754 = n25477 & n25508 ;
  assign n25755 = n25571 & n25754 ;
  assign n25756 = ~n25540 & n25755 ;
  assign n25776 = n25700 & n25756 ;
  assign n25757 = n25750 & n25756 ;
  assign n25758 = ~n25604 & n25699 ;
  assign n25759 = n25509 & n25667 ;
  assign n25760 = n25758 & n25759 ;
  assign n25761 = n25572 & n25760 ;
  assign n25785 = ~n25757 & ~n25761 ;
  assign n25786 = ~n25776 & n25785 ;
  assign n25795 = n25667 & n25699 ;
  assign n25796 = n25740 & n25795 ;
  assign n25807 = n25477 & n25572 ;
  assign n25808 = n25796 & n25807 ;
  assign n25809 = n25786 & ~n25808 ;
  assign n25810 = n25784 & n25809 ;
  assign n25735 = ~n25508 & ~n25540 ;
  assign n25736 = n25571 & n25735 ;
  assign n25737 = ~n25477 & n25736 ;
  assign n25738 = n25700 & n25737 ;
  assign n25739 = n25667 & ~n25699 ;
  assign n25741 = n25739 & n25740 ;
  assign n25742 = n25737 & n25741 ;
  assign n25743 = ~n25738 & ~n25742 ;
  assign n25713 = ~\P1_P2_InstQueueRd_Addr_reg[3]/NET0131  & \P1_P2_InstQueueWr_Addr_reg[3]/NET0131  ;
  assign n25714 = \P1_P2_InstQueueRd_Addr_reg[3]/NET0131  & ~\P1_P2_InstQueueWr_Addr_reg[3]/NET0131  ;
  assign n25702 = ~\P1_P2_InstQueueRd_Addr_reg[2]/NET0131  & \P1_P2_InstQueueWr_Addr_reg[2]/NET0131  ;
  assign n25703 = \P1_P2_InstQueueRd_Addr_reg[2]/NET0131  & ~\P1_P2_InstQueueWr_Addr_reg[2]/NET0131  ;
  assign n25705 = ~\P1_P2_InstQueueRd_Addr_reg[1]/NET0131  & \P1_P2_InstQueueWr_Addr_reg[1]/NET0131  ;
  assign n25706 = \P1_P2_InstQueueRd_Addr_reg[1]/NET0131  & ~\P1_P2_InstQueueWr_Addr_reg[1]/NET0131  ;
  assign n25707 = \P1_P2_InstQueueRd_Addr_reg[0]/NET0131  & ~\P1_P2_InstQueueWr_Addr_reg[0]/NET0131  ;
  assign n25708 = ~n25706 & ~n25707 ;
  assign n25709 = ~n25705 & ~n25708 ;
  assign n25716 = ~n25703 & ~n25709 ;
  assign n25717 = ~n25702 & ~n25716 ;
  assign n25722 = ~n25714 & ~n25717 ;
  assign n25723 = ~n25713 & ~n25722 ;
  assign n25715 = ~n25713 & ~n25714 ;
  assign n25718 = n25715 & n25717 ;
  assign n25719 = ~n25715 & ~n25717 ;
  assign n25720 = ~n25718 & ~n25719 ;
  assign n25704 = ~n25702 & ~n25703 ;
  assign n25710 = n25704 & n25709 ;
  assign n25711 = ~n25704 & ~n25709 ;
  assign n25712 = ~n25710 & ~n25711 ;
  assign n25725 = ~\P1_P2_InstQueueRd_Addr_reg[0]/NET0131  & \P1_P2_InstQueueWr_Addr_reg[0]/NET0131  ;
  assign n25726 = ~n25707 & ~n25725 ;
  assign n25727 = ~n25705 & ~n25706 ;
  assign n25744 = n25726 & n25727 ;
  assign n25745 = ~n25712 & ~n25744 ;
  assign n25746 = n25720 & ~n25745 ;
  assign n25747 = ~n25723 & ~n25746 ;
  assign n25748 = ~n25743 & ~n25747 ;
  assign n25892 = \P1_P2_InstQueueRd_Addr_reg[0]/NET0131  & ~n25748 ;
  assign n25900 = n25810 & n25892 ;
  assign n25792 = n25540 & ~n25571 ;
  assign n25793 = n25754 & n25792 ;
  assign n25794 = ~n25736 & ~n25793 ;
  assign n25797 = ~n25794 & n25796 ;
  assign n25798 = n25636 & n25739 ;
  assign n25799 = n25573 & n25798 ;
  assign n25804 = ~n25797 & ~n25799 ;
  assign n25800 = ~n25635 & n25792 ;
  assign n25801 = n25760 & n25800 ;
  assign n25802 = n25668 & n25699 ;
  assign n25803 = n25793 & n25802 ;
  assign n25805 = ~n25801 & ~n25803 ;
  assign n25806 = n25804 & n25805 ;
  assign n25811 = n25743 & n25806 ;
  assign n25812 = n25810 & n25811 ;
  assign n25813 = n25540 & n25635 ;
  assign n25814 = n25758 & n25813 ;
  assign n25815 = n25755 & n25814 ;
  assign n25816 = ~n25812 & ~n25815 ;
  assign n25817 = n25806 & n25816 ;
  assign n25887 = ~n25743 & n25747 ;
  assign n25901 = n25817 & ~n25887 ;
  assign n25902 = ~\P1_P2_InstQueueRd_Addr_reg[0]/NET0131  & n25901 ;
  assign n25903 = ~n25900 & ~n25902 ;
  assign n25415 = \P1_ready12_reg/NET0131  & \P1_ready21_reg/NET0131  ;
  assign n25721 = n25712 & n25720 ;
  assign n25724 = ~n25721 & ~n25723 ;
  assign n25728 = n25707 & ~n25727 ;
  assign n25729 = ~n25707 & n25727 ;
  assign n25730 = ~n25728 & ~n25729 ;
  assign n25731 = ~n25723 & n25730 ;
  assign n25770 = ~n25724 & ~n25731 ;
  assign n25773 = ~n25415 & ~n25770 ;
  assign n25774 = n25635 & n25761 ;
  assign n25826 = ~n25774 & ~n25776 ;
  assign n25762 = ~n25635 & n25761 ;
  assign n25763 = ~n25757 & ~n25762 ;
  assign n25764 = ~\P1_P2_State_reg[0]/NET0131  & \P1_P2_State_reg[1]/NET0131  ;
  assign n25765 = ~\P1_P2_State_reg[2]/NET0131  & n25764 ;
  assign n25766 = ~\P1_P2_State_reg[0]/NET0131  & ~\P1_P2_State_reg[1]/NET0131  ;
  assign n25767 = \P1_P2_State_reg[2]/NET0131  & n25766 ;
  assign n25768 = ~n25765 & ~n25767 ;
  assign n25827 = ~n25763 & ~n25768 ;
  assign n25828 = n25826 & ~n25827 ;
  assign n25829 = n25773 & ~n25828 ;
  assign n25830 = ~n25808 & ~n25829 ;
  assign n25888 = n25806 & ~n25887 ;
  assign n25889 = \P1_P2_InstQueueRd_Addr_reg[0]/NET0131  & ~n25888 ;
  assign n25890 = n25830 & ~n25889 ;
  assign n25891 = ~\P1_P2_InstQueueRd_Addr_reg[1]/NET0131  & ~n25890 ;
  assign n25885 = ~n25427 & ~n25430 ;
  assign n25886 = ~n25816 & ~n25885 ;
  assign n25893 = ~n25811 & ~n25892 ;
  assign n25769 = ~n25415 & ~n25768 ;
  assign n25771 = n25769 & ~n25770 ;
  assign n25772 = ~n25763 & ~n25771 ;
  assign n25775 = ~n25773 & n25774 ;
  assign n25777 = ~n25773 & n25776 ;
  assign n25778 = ~n25775 & ~n25777 ;
  assign n25779 = ~n25772 & n25778 ;
  assign n25894 = n25779 & n25784 ;
  assign n25895 = ~n25893 & n25894 ;
  assign n25896 = \P1_P2_InstQueueRd_Addr_reg[1]/NET0131  & ~n25895 ;
  assign n25897 = ~n25886 & ~n25896 ;
  assign n25898 = ~n25891 & n25897 ;
  assign n25899 = ~\P1_P2_InstQueueWr_Addr_reg[1]/NET0131  & ~n25898 ;
  assign n25904 = \P1_P2_InstQueueWr_Addr_reg[0]/NET0131  & ~n25899 ;
  assign n25905 = ~n25903 & n25904 ;
  assign n25818 = ~\P1_P2_InstQueueRd_Addr_reg[2]/NET0131  & ~n25433 ;
  assign n25819 = ~n25434 & ~n25818 ;
  assign n25820 = ~n25817 & n25819 ;
  assign n25831 = ~\P1_P2_InstQueueRd_Addr_reg[1]/NET0131  & ~\P1_P2_InstQueueRd_Addr_reg[2]/NET0131  ;
  assign n25832 = ~n25451 & ~n25831 ;
  assign n25833 = ~n25830 & n25832 ;
  assign n25787 = ~n25763 & n25768 ;
  assign n25788 = n25773 & ~n25787 ;
  assign n25789 = ~n25786 & ~n25788 ;
  assign n25790 = n25784 & ~n25789 ;
  assign n25791 = \P1_P2_InstQueueRd_Addr_reg[2]/NET0131  & ~n25790 ;
  assign n25821 = n25747 & ~n25818 ;
  assign n25822 = ~n25434 & n25821 ;
  assign n25823 = ~\P1_P2_InstQueueRd_Addr_reg[2]/NET0131  & ~n25747 ;
  assign n25824 = ~n25822 & ~n25823 ;
  assign n25825 = ~n25743 & n25824 ;
  assign n25834 = ~n25791 & ~n25825 ;
  assign n25835 = ~n25833 & n25834 ;
  assign n25836 = ~n25820 & n25835 ;
  assign n25884 = \P1_P2_InstQueueWr_Addr_reg[2]/NET0131  & n25836 ;
  assign n25857 = \P1_P2_InstQueueRd_Addr_reg[3]/NET0131  & ~n25434 ;
  assign n25858 = ~n25435 & ~n25857 ;
  assign n25859 = ~n25817 & ~n25858 ;
  assign n25846 = ~n25770 & n25776 ;
  assign n25847 = ~n25770 & n25827 ;
  assign n25848 = ~n25846 & ~n25847 ;
  assign n25837 = \P1_P2_InstQueueRd_Addr_reg[3]/NET0131  & ~n25451 ;
  assign n25838 = ~n25452 & ~n25837 ;
  assign n25849 = ~n25415 & ~n25838 ;
  assign n25850 = \P1_P2_InstQueueRd_Addr_reg[3]/NET0131  & n25415 ;
  assign n25851 = ~n25849 & ~n25850 ;
  assign n25852 = ~n25848 & ~n25851 ;
  assign n25841 = ~n25768 & ~n25770 ;
  assign n25842 = ~n25763 & ~n25841 ;
  assign n25840 = n25770 & n25776 ;
  assign n25843 = n25784 & ~n25840 ;
  assign n25844 = ~n25842 & n25843 ;
  assign n25845 = \P1_P2_InstQueueRd_Addr_reg[3]/NET0131  & ~n25844 ;
  assign n25860 = ~\P1_P2_InstQueueRd_Addr_reg[3]/NET0131  & n25770 ;
  assign n25861 = ~n25770 & n25851 ;
  assign n25862 = ~n25860 & ~n25861 ;
  assign n25863 = n25774 & n25862 ;
  assign n25839 = n25808 & ~n25838 ;
  assign n25853 = ~\P1_P2_InstQueueRd_Addr_reg[3]/NET0131  & ~n25821 ;
  assign n25854 = \P1_P2_InstQueueRd_Addr_reg[3]/NET0131  & n25821 ;
  assign n25855 = ~n25853 & ~n25854 ;
  assign n25856 = ~n25743 & n25855 ;
  assign n25864 = ~n25839 & ~n25856 ;
  assign n25865 = ~n25863 & n25864 ;
  assign n25866 = ~n25845 & n25865 ;
  assign n25867 = ~n25852 & n25866 ;
  assign n25868 = ~n25859 & n25867 ;
  assign n25869 = \P1_P2_InstQueueWr_Addr_reg[3]/NET0131  & n25868 ;
  assign n25906 = \P1_P2_InstQueueWr_Addr_reg[1]/NET0131  & n25898 ;
  assign n25907 = ~n25869 & ~n25906 ;
  assign n25908 = ~n25884 & n25907 ;
  assign n25909 = ~n25905 & n25908 ;
  assign n25872 = \P1_P2_InstQueueWr_Addr_reg[3]/NET0131  & n25836 ;
  assign n25873 = ~n25868 & ~n25872 ;
  assign n25870 = ~\P1_P2_InstQueueWr_Addr_reg[2]/NET0131  & ~n25836 ;
  assign n25871 = ~n25869 & n25870 ;
  assign n25780 = ~\P1_P2_More_reg/NET0131  & ~n25770 ;
  assign n25781 = ~n25779 & ~n25780 ;
  assign n25732 = ~n25726 & n25731 ;
  assign n25733 = ~n25724 & ~n25732 ;
  assign n25734 = n25701 & n25733 ;
  assign n25752 = ~n25747 & n25751 ;
  assign n25753 = ~n25748 & ~n25752 ;
  assign n25782 = ~n25734 & n25753 ;
  assign n25783 = ~n25781 & n25782 ;
  assign n25875 = ~n25770 & ~n25826 ;
  assign n25876 = n25415 & n25875 ;
  assign n25877 = ~n25763 & ~n25770 ;
  assign n25878 = ~n25769 & n25877 ;
  assign n25879 = ~n25876 & ~n25878 ;
  assign n25880 = \P1_P2_Flush_reg/NET0131  & ~n25879 ;
  assign n25874 = n25701 & ~n25733 ;
  assign n25881 = n25747 & n25751 ;
  assign n25882 = ~n25874 & ~n25881 ;
  assign n25883 = ~n25880 & n25882 ;
  assign n25910 = n25783 & n25883 ;
  assign n25911 = ~n25871 & n25910 ;
  assign n25912 = ~n25873 & n25911 ;
  assign n25913 = ~n25909 & n25912 ;
  assign n25914 = ~\P1_P2_DataWidth_reg[1]/NET0131  & n25757 ;
  assign n25915 = n25771 & n25914 ;
  assign n25916 = n25913 & ~n25915 ;
  assign n25416 = \P1_P2_State2_reg[0]/NET0131  & ~\P1_P2_State2_reg[3]/NET0131  ;
  assign n25917 = ~\P1_P2_State2_reg[1]/NET0131  & \P1_P2_State2_reg[2]/NET0131  ;
  assign n25918 = n25416 & n25917 ;
  assign n25919 = ~n25916 & n25918 ;
  assign n25920 = \P1_P2_State2_reg[1]/NET0131  & \P1_P2_State2_reg[2]/NET0131  ;
  assign n25921 = ~\P1_P2_State2_reg[3]/NET0131  & n25920 ;
  assign n25922 = ~\P1_P2_State2_reg[0]/NET0131  & n25921 ;
  assign n25923 = \P1_P2_State2_reg[1]/NET0131  & ~\P1_P2_State2_reg[2]/NET0131  ;
  assign n25924 = ~\P1_P2_State2_reg[3]/NET0131  & n25923 ;
  assign n25925 = \P1_P2_State2_reg[0]/NET0131  & n25924 ;
  assign n25926 = ~n25922 & ~n25925 ;
  assign n25927 = n25415 & ~n25926 ;
  assign n25417 = ~\P1_P2_State2_reg[2]/NET0131  & n25416 ;
  assign n25418 = ~\P1_P2_State2_reg[1]/NET0131  & n25417 ;
  assign n25419 = ~n25415 & n25418 ;
  assign n25928 = ~\P1_P2_State2_reg[0]/NET0131  & n25924 ;
  assign n25929 = ~\P1_P2_DataWidth_reg[1]/NET0131  & n25928 ;
  assign n25930 = ~n25419 & ~n25929 ;
  assign n25931 = ~n25927 & n25930 ;
  assign n25932 = ~n25919 & n25931 ;
  assign n25936 = ~n25415 & ~n25926 ;
  assign n25933 = \P1_P2_DataWidth_reg[1]/NET0131  & n25928 ;
  assign n25934 = ~\P1_P2_State2_reg[0]/NET0131  & ~\P1_P2_State2_reg[3]/NET0131  ;
  assign n25935 = \P1_P2_State2_reg[2]/NET0131  & n25934 ;
  assign n25937 = ~n25918 & ~n25935 ;
  assign n25938 = ~n25933 & n25937 ;
  assign n25939 = ~n25936 & n25938 ;
  assign n25944 = n21058 & n21065 ;
  assign n25945 = n21057 & n25944 ;
  assign n25963 = n21065 & n24897 ;
  assign n25982 = ~n25945 & ~n25963 ;
  assign n25983 = n14612 & n21064 ;
  assign n25984 = n21018 & n25983 ;
  assign n25985 = n25982 & ~n25984 ;
  assign n25951 = ~n14799 & n21067 ;
  assign n25952 = ~n24898 & ~n25951 ;
  assign n25986 = n20725 & n21059 ;
  assign n25987 = ~n20727 & ~n25986 ;
  assign n25988 = n25952 & n25987 ;
  assign n25989 = n21070 & n25988 ;
  assign n25990 = n25985 & n25989 ;
  assign n25969 = ~n20724 & ~n21021 ;
  assign n25970 = n21018 & ~n25969 ;
  assign n25975 = n11689 & n12766 ;
  assign n25976 = ~n14068 & n14799 ;
  assign n25977 = n25975 & n25976 ;
  assign n25978 = n21060 & n25977 ;
  assign n25979 = n12766 & ~n17417 ;
  assign n25980 = n21058 & n25979 ;
  assign n25981 = n21021 & n25980 ;
  assign n25991 = ~n25978 & ~n25981 ;
  assign n25992 = ~n25970 & n25991 ;
  assign n25971 = ~n14799 & n21020 ;
  assign n25972 = n21063 & n25971 ;
  assign n25973 = n21066 & n25972 ;
  assign n25974 = n20721 & n25944 ;
  assign n25993 = ~n25973 & ~n25974 ;
  assign n25994 = n25992 & n25993 ;
  assign n25995 = ~n25990 & n25994 ;
  assign n26068 = n20720 & ~n25987 ;
  assign n26069 = n25995 & ~n26068 ;
  assign n26070 = ~n11645 & ~n11658 ;
  assign n26071 = ~n26069 & n26070 ;
  assign n26036 = ~n21082 & n25982 ;
  assign n26053 = ~n20720 & ~n25987 ;
  assign n26072 = ~n25987 & n26070 ;
  assign n26073 = ~n26053 & ~n26072 ;
  assign n26074 = n26036 & n26073 ;
  assign n26075 = \P2_P1_InstQueueRd_Addr_reg[1]/NET0131  & ~n26074 ;
  assign n25949 = ~n21069 & ~n21081 ;
  assign n26064 = ~\P2_P1_InstQueueRd_Addr_reg[1]/NET0131  & ~n21073 ;
  assign n26065 = \P2_P1_InstQueueRd_Addr_reg[1]/NET0131  & n21073 ;
  assign n26066 = ~n26064 & ~n26065 ;
  assign n26067 = n25949 & ~n26066 ;
  assign n26076 = ~\P2_P1_InstQueueRd_Addr_reg[1]/NET0131  & n25984 ;
  assign n25954 = ~\P2_P1_State_reg[0]/NET0131  & \P2_P1_State_reg[1]/NET0131  ;
  assign n25955 = ~\P2_P1_State_reg[2]/NET0131  & n25954 ;
  assign n25956 = ~\P2_P1_State_reg[0]/NET0131  & ~\P2_P1_State_reg[1]/NET0131  ;
  assign n25957 = \P2_P1_State_reg[2]/NET0131  & n25956 ;
  assign n25958 = ~n25955 & ~n25957 ;
  assign n26006 = ~n21081 & ~n25958 ;
  assign n26077 = ~\P2_P1_InstQueueRd_Addr_reg[1]/NET0131  & ~n26006 ;
  assign n26078 = n26006 & n26066 ;
  assign n26079 = ~n26077 & ~n26078 ;
  assign n26080 = ~n25952 & n26079 ;
  assign n26081 = ~n26076 & ~n26080 ;
  assign n26082 = ~n26067 & n26081 ;
  assign n26083 = ~n26075 & n26082 ;
  assign n26084 = ~n26071 & n26083 ;
  assign n26085 = ~\P2_P1_InstQueueWr_Addr_reg[1]/NET0131  & ~n26084 ;
  assign n26086 = ~\P2_P1_InstQueueRd_Addr_reg[0]/NET0131  & n26069 ;
  assign n26089 = \P2_P1_InstQueueRd_Addr_reg[0]/NET0131  & n25985 ;
  assign n26087 = ~n21062 & ~n21067 ;
  assign n26088 = ~n24898 & n26087 ;
  assign n26090 = ~n26053 & n26088 ;
  assign n26091 = n26089 & n26090 ;
  assign n26092 = ~n26086 & ~n26091 ;
  assign n26093 = \P2_P1_InstQueueWr_Addr_reg[0]/NET0131  & ~n26092 ;
  assign n26094 = ~n26085 & n26093 ;
  assign n26095 = \P2_P1_InstQueueWr_Addr_reg[1]/NET0131  & n26084 ;
  assign n25967 = \P2_P1_InstQueueRd_Addr_reg[3]/NET0131  & ~n11646 ;
  assign n25968 = ~n11661 & ~n25967 ;
  assign n25996 = ~n25968 & ~n25995 ;
  assign n25997 = ~\P2_P1_InstQueueRd_Addr_reg[3]/NET0131  & n21081 ;
  assign n25998 = \P2_P1_InstQueueRd_Addr_reg[3]/NET0131  & ~n11649 ;
  assign n25999 = ~n11650 & ~n25998 ;
  assign n26000 = ~n21073 & ~n25999 ;
  assign n26001 = \P2_P1_InstQueueRd_Addr_reg[3]/NET0131  & n21073 ;
  assign n26002 = ~n26000 & ~n26001 ;
  assign n26003 = ~n21081 & n26002 ;
  assign n26004 = ~n25997 & ~n26003 ;
  assign n26005 = ~n21069 & n26004 ;
  assign n26018 = n25984 & ~n25999 ;
  assign n26019 = ~n26005 & ~n26018 ;
  assign n26017 = \P2_P1_InstQueueRd_Addr_reg[3]/NET0131  & ~n25982 ;
  assign n26007 = n26002 & n26006 ;
  assign n26008 = ~\P2_P1_InstQueueRd_Addr_reg[3]/NET0131  & ~n26006 ;
  assign n26009 = ~n26007 & ~n26008 ;
  assign n26010 = ~n25952 & n26009 ;
  assign n26011 = ~\P2_P1_InstQueueRd_Addr_reg[2]/NET0131  & ~n11645 ;
  assign n26012 = n20720 & ~n26011 ;
  assign n26013 = ~\P2_P1_InstQueueRd_Addr_reg[3]/NET0131  & ~n26012 ;
  assign n26014 = \P2_P1_InstQueueRd_Addr_reg[3]/NET0131  & n26012 ;
  assign n26015 = ~n26013 & ~n26014 ;
  assign n26016 = ~n25987 & n26015 ;
  assign n26020 = ~n26010 & ~n26016 ;
  assign n26021 = ~n26017 & n26020 ;
  assign n26022 = n26019 & n26021 ;
  assign n26023 = ~n25996 & n26022 ;
  assign n26024 = \P2_P1_InstQueueWr_Addr_reg[3]/NET0131  & n26023 ;
  assign n26028 = ~n11646 & ~n26011 ;
  assign n26029 = ~n25995 & n26028 ;
  assign n26037 = ~n25952 & ~n26006 ;
  assign n26038 = n26036 & ~n26037 ;
  assign n26039 = \P2_P1_InstQueueRd_Addr_reg[2]/NET0131  & ~n26038 ;
  assign n26030 = ~n25952 & n26006 ;
  assign n26031 = ~n25949 & ~n26030 ;
  assign n26025 = ~\P2_P1_InstQueueRd_Addr_reg[1]/NET0131  & ~\P2_P1_InstQueueRd_Addr_reg[2]/NET0131  ;
  assign n26026 = ~n11649 & ~n26025 ;
  assign n26032 = ~n21073 & ~n26026 ;
  assign n26033 = ~\P2_P1_InstQueueRd_Addr_reg[2]/NET0131  & n21073 ;
  assign n26034 = ~n26032 & ~n26033 ;
  assign n26035 = ~n26031 & n26034 ;
  assign n26027 = n25984 & n26026 ;
  assign n26040 = ~\P2_P1_InstQueueRd_Addr_reg[2]/NET0131  & ~n20720 ;
  assign n26041 = n20720 & n26028 ;
  assign n26042 = ~n26040 & ~n26041 ;
  assign n26043 = ~n25987 & n26042 ;
  assign n26044 = ~n26027 & ~n26043 ;
  assign n26045 = ~n26035 & n26044 ;
  assign n26046 = ~n26039 & n26045 ;
  assign n26047 = ~n26029 & n26046 ;
  assign n26063 = \P2_P1_InstQueueWr_Addr_reg[2]/NET0131  & n26047 ;
  assign n26096 = ~n26024 & ~n26063 ;
  assign n26097 = ~n26095 & n26096 ;
  assign n26098 = ~n26094 & n26097 ;
  assign n26050 = \P2_P1_InstQueueWr_Addr_reg[3]/NET0131  & n26047 ;
  assign n26051 = ~n26023 & ~n26050 ;
  assign n26048 = ~\P2_P1_InstQueueWr_Addr_reg[2]/NET0131  & ~n26047 ;
  assign n26049 = ~n26024 & n26048 ;
  assign n25950 = n21073 & n25949 ;
  assign n25953 = ~n21081 & ~n25952 ;
  assign n25959 = ~n21073 & ~n25958 ;
  assign n25960 = n25953 & ~n25959 ;
  assign n25961 = ~n25950 & ~n25960 ;
  assign n25962 = \P2_P1_Flush_reg/NET0131  & ~n25961 ;
  assign n25946 = ~n20698 & n21080 ;
  assign n25947 = ~n21076 & ~n25946 ;
  assign n25948 = n25945 & ~n25947 ;
  assign n25964 = n20720 & n25963 ;
  assign n25965 = ~n25948 & ~n25964 ;
  assign n25966 = ~n25962 & n25965 ;
  assign n26052 = n25945 & n25947 ;
  assign n26054 = ~n20720 & n25963 ;
  assign n26055 = ~n26053 & ~n26054 ;
  assign n26056 = ~n26052 & n26055 ;
  assign n26059 = ~n24711 & n25952 ;
  assign n26057 = ~n21081 & n25959 ;
  assign n26058 = ~\P2_P1_More_reg/NET0131  & ~n21081 ;
  assign n26060 = ~n26057 & ~n26058 ;
  assign n26061 = ~n26059 & n26060 ;
  assign n26062 = n26056 & ~n26061 ;
  assign n26099 = n25966 & n26062 ;
  assign n26100 = ~n26049 & n26099 ;
  assign n26101 = ~n26051 & n26100 ;
  assign n26102 = ~n26098 & n26101 ;
  assign n26103 = ~\P2_P1_DataWidth_reg[1]/NET0131  & n25959 ;
  assign n26104 = n24898 & n26103 ;
  assign n26105 = ~n21081 & n26104 ;
  assign n26106 = n26102 & ~n26105 ;
  assign n26107 = n11623 & ~n26106 ;
  assign n25940 = \P2_P1_State2_reg[2]/NET0131  & n11611 ;
  assign n25941 = ~n21098 & ~n25940 ;
  assign n25942 = \P2_P1_State2_reg[1]/NET0131  & ~n25941 ;
  assign n25943 = n21073 & n25942 ;
  assign n26108 = ~\P2_P1_DataWidth_reg[1]/NET0131  & n11609 ;
  assign n26109 = n11618 & ~n21073 ;
  assign n26110 = ~n26108 & ~n26109 ;
  assign n26111 = ~n25943 & n26110 ;
  assign n26112 = ~n26107 & n26111 ;
  assign n26154 = ~\P1_P1_State_reg[0]/NET0131  & \P1_P1_State_reg[1]/NET0131  ;
  assign n26155 = ~\P1_P1_State_reg[2]/NET0131  & n26154 ;
  assign n26156 = ~\P1_P1_State_reg[0]/NET0131  & ~\P1_P1_State_reg[1]/NET0131  ;
  assign n26157 = \P1_P1_State_reg[2]/NET0131  & n26156 ;
  assign n26158 = ~n26155 & ~n26157 ;
  assign n26159 = ~n14020 & n15382 ;
  assign n26160 = ~n24502 & ~n26159 ;
  assign n26161 = ~n15364 & ~n26160 ;
  assign n26162 = ~n26158 & n26161 ;
  assign n26163 = ~n24341 & ~n26162 ;
  assign n26164 = \P1_P1_InstQueueRd_Addr_reg[2]/NET0131  & ~n26160 ;
  assign n26165 = n26163 & ~n26164 ;
  assign n26179 = n15335 & ~n26165 ;
  assign n26124 = n15380 & n24501 ;
  assign n26125 = n15328 & n15380 ;
  assign n26126 = n15329 & n26125 ;
  assign n26127 = ~n26124 & ~n26126 ;
  assign n26174 = n15334 & n15364 ;
  assign n26175 = ~n15364 & ~n26158 ;
  assign n26176 = ~n26160 & ~n26175 ;
  assign n26177 = ~n26174 & ~n26176 ;
  assign n26178 = n26127 & n26177 ;
  assign n26180 = ~n15419 & n26178 ;
  assign n26181 = ~n26179 & n26180 ;
  assign n26182 = \P1_P1_InstQueueRd_Addr_reg[2]/NET0131  & ~n26181 ;
  assign n26128 = n13639 & n15378 ;
  assign n26129 = n15376 & n26128 ;
  assign n26166 = ~n15335 & ~n26165 ;
  assign n26167 = ~n26129 & ~n26166 ;
  assign n26153 = ~\P1_P1_InstQueueRd_Addr_reg[1]/NET0131  & ~\P1_P1_InstQueueRd_Addr_reg[2]/NET0131  ;
  assign n26168 = ~n8289 & ~n26153 ;
  assign n26169 = ~n26167 & n26168 ;
  assign n26117 = ~\P1_P1_InstQueueRd_Addr_reg[2]/NET0131  & ~n8311 ;
  assign n26118 = \P1_P1_InstQueueRd_Addr_reg[2]/NET0131  & n8311 ;
  assign n26119 = ~n26117 & ~n26118 ;
  assign n26122 = n15330 & n15370 ;
  assign n26123 = ~n15372 & ~n26122 ;
  assign n26130 = ~n15334 & ~n15382 ;
  assign n26131 = ~n24502 & n26130 ;
  assign n26132 = ~n26129 & n26131 ;
  assign n26133 = n26127 & n26132 ;
  assign n26134 = n26123 & n26133 ;
  assign n26120 = ~n15369 & ~n15374 ;
  assign n26121 = n15376 & ~n26120 ;
  assign n26140 = n10096 & ~n12718 ;
  assign n26141 = n14020 & n26140 ;
  assign n26139 = n8345 & n9362 ;
  assign n26142 = n15331 & n26139 ;
  assign n26143 = n26141 & n26142 ;
  assign n26144 = n10096 & ~n14751 ;
  assign n26145 = n15328 & n26144 ;
  assign n26146 = n15374 & n26145 ;
  assign n26147 = ~n26143 & ~n26146 ;
  assign n26148 = ~n26121 & n26147 ;
  assign n26135 = ~n14020 & n15373 ;
  assign n26136 = n15379 & n26135 ;
  assign n26137 = n15381 & n26136 ;
  assign n26138 = n15367 & n26125 ;
  assign n26149 = ~n26137 & ~n26138 ;
  assign n26150 = n26148 & n26149 ;
  assign n26151 = ~n26134 & n26150 ;
  assign n26152 = n26119 & ~n26151 ;
  assign n26170 = ~\P1_P1_InstQueueRd_Addr_reg[2]/NET0131  & ~n15428 ;
  assign n26171 = n15428 & n26119 ;
  assign n26172 = ~n26170 & ~n26171 ;
  assign n26173 = ~n26123 & n26172 ;
  assign n26183 = ~n26152 & ~n26173 ;
  assign n26184 = ~n26169 & n26183 ;
  assign n26185 = ~n26182 & n26184 ;
  assign n26187 = ~\P1_P1_InstQueueWr_Addr_reg[2]/NET0131  & ~n26185 ;
  assign n26191 = ~n8293 & ~n8311 ;
  assign n26192 = n15428 & ~n26123 ;
  assign n26193 = n26151 & ~n26192 ;
  assign n26194 = \P1_P1_InstQueueRd_Addr_reg[1]/NET0131  & ~n26123 ;
  assign n26195 = n26193 & ~n26194 ;
  assign n26196 = n26191 & ~n26195 ;
  assign n26188 = ~n15335 & ~n26163 ;
  assign n26189 = ~n26129 & ~n26188 ;
  assign n26190 = ~\P1_P1_InstQueueRd_Addr_reg[1]/NET0131  & ~n26189 ;
  assign n26200 = n15335 & ~n26163 ;
  assign n26197 = ~n15428 & ~n26123 ;
  assign n26198 = \P1_P1_InstQueueRd_Addr_reg[0]/NET0131  & n26197 ;
  assign n26199 = ~n15365 & n15383 ;
  assign n26201 = ~n26198 & ~n26199 ;
  assign n26202 = n26178 & n26201 ;
  assign n26203 = ~n26200 & n26202 ;
  assign n26204 = \P1_P1_InstQueueRd_Addr_reg[1]/NET0131  & ~n26203 ;
  assign n26205 = ~n26190 & ~n26204 ;
  assign n26206 = ~n26196 & n26205 ;
  assign n26207 = \P1_P1_InstQueueWr_Addr_reg[1]/NET0131  & n26206 ;
  assign n26208 = ~\P1_P1_InstQueueWr_Addr_reg[1]/NET0131  & ~n26206 ;
  assign n26209 = ~\P1_P1_InstQueueRd_Addr_reg[0]/NET0131  & n26193 ;
  assign n26210 = \P1_P1_InstQueueRd_Addr_reg[0]/NET0131  & ~n26197 ;
  assign n26211 = n26133 & n26210 ;
  assign n26212 = ~n26209 & ~n26211 ;
  assign n26213 = \P1_P1_InstQueueWr_Addr_reg[0]/NET0131  & ~n26212 ;
  assign n26214 = ~n26208 & n26213 ;
  assign n26215 = ~n26207 & ~n26214 ;
  assign n26216 = ~n26187 & ~n26215 ;
  assign n26186 = \P1_P1_InstQueueWr_Addr_reg[2]/NET0131  & n26185 ;
  assign n26237 = \P1_P1_InstQueueRd_Addr_reg[3]/NET0131  & ~n26118 ;
  assign n26238 = ~n8318 & ~n26237 ;
  assign n26239 = ~n26151 & ~n26238 ;
  assign n26217 = ~\P1_P1_InstQueueRd_Addr_reg[3]/NET0131  & ~n8289 ;
  assign n26218 = ~n8290 & ~n26217 ;
  assign n26220 = ~n15335 & n26218 ;
  assign n26221 = \P1_P1_InstQueueRd_Addr_reg[3]/NET0131  & n15335 ;
  assign n26222 = ~n26220 & ~n26221 ;
  assign n26223 = ~n26160 & ~n26222 ;
  assign n26224 = n26178 & ~n26223 ;
  assign n26225 = \P1_P1_InstQueueRd_Addr_reg[3]/NET0131  & ~n26224 ;
  assign n26235 = ~n24504 & ~n26162 ;
  assign n26236 = ~n26222 & ~n26235 ;
  assign n26230 = n15428 & ~n26117 ;
  assign n26231 = ~\P1_P1_InstQueueRd_Addr_reg[3]/NET0131  & ~n26230 ;
  assign n26232 = \P1_P1_InstQueueRd_Addr_reg[3]/NET0131  & n26230 ;
  assign n26233 = ~n26231 & ~n26232 ;
  assign n26234 = ~n26123 & n26233 ;
  assign n26219 = n26129 & n26218 ;
  assign n26226 = ~\P1_P1_InstQueueRd_Addr_reg[3]/NET0131  & n15364 ;
  assign n26227 = ~n15364 & n26222 ;
  assign n26228 = ~n26226 & ~n26227 ;
  assign n26229 = n15383 & n26228 ;
  assign n26240 = ~n26219 & ~n26229 ;
  assign n26241 = ~n26234 & n26240 ;
  assign n26242 = ~n26236 & n26241 ;
  assign n26243 = ~n26225 & n26242 ;
  assign n26244 = ~n26239 & n26243 ;
  assign n26245 = \P1_P1_InstQueueWr_Addr_reg[3]/NET0131  & n26244 ;
  assign n26246 = ~n26186 & ~n26245 ;
  assign n26247 = ~n26216 & n26246 ;
  assign n26260 = \P1_P1_InstQueueWr_Addr_reg[3]/NET0131  & n26185 ;
  assign n26261 = ~n26244 & ~n26260 ;
  assign n26253 = ~\P1_P1_More_reg/NET0131  & ~n15364 ;
  assign n26254 = n15365 & ~n26158 ;
  assign n26255 = ~n26160 & ~n26254 ;
  assign n26256 = ~n24345 & ~n26255 ;
  assign n26257 = ~n26253 & ~n26256 ;
  assign n26248 = n15363 & ~n15424 ;
  assign n26249 = ~n15358 & ~n26248 ;
  assign n26250 = n26126 & n26249 ;
  assign n26251 = ~n15428 & n26124 ;
  assign n26252 = ~n26197 & ~n26251 ;
  assign n26258 = ~n26250 & n26252 ;
  assign n26259 = ~n26257 & n26258 ;
  assign n26264 = ~n15335 & ~n26158 ;
  assign n26265 = n26161 & ~n26264 ;
  assign n26266 = ~n15384 & n25363 ;
  assign n26267 = ~n26265 & ~n26266 ;
  assign n26268 = \P1_P1_Flush_reg/NET0131  & ~n26267 ;
  assign n26262 = n26126 & ~n26249 ;
  assign n26263 = n15428 & n26124 ;
  assign n26269 = ~n26262 & ~n26263 ;
  assign n26270 = ~n26268 & n26269 ;
  assign n26271 = n26259 & n26270 ;
  assign n26272 = ~n26261 & n26271 ;
  assign n26273 = ~n26247 & n26272 ;
  assign n26274 = ~\P1_P1_DataWidth_reg[1]/NET0131  & ~n15335 ;
  assign n26275 = ~n26158 & n26274 ;
  assign n26276 = n24503 & n26275 ;
  assign n26277 = ~\P1_P1_State2_reg[1]/NET0131  & ~n26276 ;
  assign n26278 = n26273 & n26277 ;
  assign n26279 = n8355 & ~n26278 ;
  assign n26113 = \P1_P1_State2_reg[2]/NET0131  & n8356 ;
  assign n26114 = ~n15324 & ~n26113 ;
  assign n26115 = \P1_P1_State2_reg[1]/NET0131  & ~n26114 ;
  assign n26116 = n15335 & n26115 ;
  assign n26280 = ~\P1_P1_DataWidth_reg[1]/NET0131  & n8282 ;
  assign n26281 = n8359 & ~n15335 ;
  assign n26282 = ~n26280 & ~n26281 ;
  assign n26283 = ~n26116 & n26282 ;
  assign n26284 = ~n26279 & n26283 ;
  assign n26701 = \P2_P2_InstQueueRd_Addr_reg[1]/NET0131  & \P2_P2_InstQueueRd_Addr_reg[2]/NET0131  ;
  assign n26312 = \P2_P2_InstQueueRd_Addr_reg[2]/NET0131  & \P2_P2_InstQueueRd_Addr_reg[3]/NET0131  ;
  assign n26329 = \P2_P2_InstQueueRd_Addr_reg[1]/NET0131  & n26312 ;
  assign n26330 = ~\P2_P2_InstQueueRd_Addr_reg[0]/NET0131  & n26329 ;
  assign n26462 = \P2_P2_InstQueue_reg[14][2]/NET0131  & n26330 ;
  assign n26309 = \P2_P2_InstQueueRd_Addr_reg[0]/NET0131  & \P2_P2_InstQueueRd_Addr_reg[1]/NET0131  ;
  assign n26324 = \P2_P2_InstQueueRd_Addr_reg[2]/NET0131  & n26309 ;
  assign n26325 = \P2_P2_InstQueueRd_Addr_reg[3]/NET0131  & n26324 ;
  assign n26460 = \P2_P2_InstQueue_reg[15][2]/NET0131  & n26325 ;
  assign n26298 = \P2_P2_InstQueueRd_Addr_reg[2]/NET0131  & ~\P2_P2_InstQueueRd_Addr_reg[3]/NET0131  ;
  assign n26299 = ~\P2_P2_InstQueueRd_Addr_reg[0]/NET0131  & \P2_P2_InstQueueRd_Addr_reg[1]/NET0131  ;
  assign n26300 = n26298 & n26299 ;
  assign n26451 = \P2_P2_InstQueue_reg[6][2]/NET0131  & n26300 ;
  assign n26306 = ~\P2_P2_InstQueueRd_Addr_reg[0]/NET0131  & ~\P2_P2_InstQueueRd_Addr_reg[1]/NET0131  ;
  assign n26307 = n26298 & n26306 ;
  assign n26452 = \P2_P2_InstQueue_reg[4][2]/NET0131  & n26307 ;
  assign n26467 = ~n26451 & ~n26452 ;
  assign n26477 = ~n26460 & n26467 ;
  assign n26478 = ~n26462 & n26477 ;
  assign n26315 = ~\P2_P2_InstQueueRd_Addr_reg[2]/NET0131  & ~\P2_P2_InstQueueRd_Addr_reg[3]/NET0131  ;
  assign n26322 = n26306 & n26315 ;
  assign n26463 = \P2_P2_InstQueue_reg[0][2]/NET0131  & n26322 ;
  assign n26302 = ~\P2_P2_InstQueueRd_Addr_reg[2]/NET0131  & \P2_P2_InstQueueRd_Addr_reg[3]/NET0131  ;
  assign n26334 = n26302 & n26306 ;
  assign n26464 = \P2_P2_InstQueue_reg[8][2]/NET0131  & n26334 ;
  assign n26472 = ~n26463 & ~n26464 ;
  assign n26320 = n26299 & n26302 ;
  assign n26465 = \P2_P2_InstQueue_reg[10][2]/NET0131  & n26320 ;
  assign n26332 = n26309 & n26315 ;
  assign n26466 = \P2_P2_InstQueue_reg[3][2]/NET0131  & n26332 ;
  assign n26473 = ~n26465 & ~n26466 ;
  assign n26474 = n26472 & n26473 ;
  assign n26303 = \P2_P2_InstQueueRd_Addr_reg[0]/NET0131  & ~\P2_P2_InstQueueRd_Addr_reg[1]/NET0131  ;
  assign n26336 = n26303 & n26312 ;
  assign n26457 = \P2_P2_InstQueue_reg[13][2]/NET0131  & n26336 ;
  assign n26338 = n26303 & n26315 ;
  assign n26458 = \P2_P2_InstQueue_reg[1][2]/NET0131  & n26338 ;
  assign n26470 = ~n26457 & ~n26458 ;
  assign n26316 = n26299 & n26315 ;
  assign n26459 = \P2_P2_InstQueue_reg[2][2]/NET0131  & n26316 ;
  assign n26327 = n26298 & n26309 ;
  assign n26461 = \P2_P2_InstQueue_reg[7][2]/NET0131  & n26327 ;
  assign n26471 = ~n26459 & ~n26461 ;
  assign n26475 = n26470 & n26471 ;
  assign n26313 = n26306 & n26312 ;
  assign n26453 = \P2_P2_InstQueue_reg[12][2]/NET0131  & n26313 ;
  assign n26310 = n26302 & n26309 ;
  assign n26454 = \P2_P2_InstQueue_reg[11][2]/NET0131  & n26310 ;
  assign n26468 = ~n26453 & ~n26454 ;
  assign n26304 = n26302 & n26303 ;
  assign n26455 = \P2_P2_InstQueue_reg[9][2]/NET0131  & n26304 ;
  assign n26318 = n26298 & n26303 ;
  assign n26456 = \P2_P2_InstQueue_reg[5][2]/NET0131  & n26318 ;
  assign n26469 = ~n26455 & ~n26456 ;
  assign n26476 = n26468 & n26469 ;
  assign n26479 = n26475 & n26476 ;
  assign n26480 = n26474 & n26479 ;
  assign n26481 = n26478 & n26480 ;
  assign n26493 = \P2_P2_InstQueue_reg[14][1]/NET0131  & n26330 ;
  assign n26491 = \P2_P2_InstQueue_reg[15][1]/NET0131  & n26325 ;
  assign n26482 = \P2_P2_InstQueue_reg[6][1]/NET0131  & n26300 ;
  assign n26483 = \P2_P2_InstQueue_reg[4][1]/NET0131  & n26307 ;
  assign n26498 = ~n26482 & ~n26483 ;
  assign n26508 = ~n26491 & n26498 ;
  assign n26509 = ~n26493 & n26508 ;
  assign n26494 = \P2_P2_InstQueue_reg[0][1]/NET0131  & n26322 ;
  assign n26495 = \P2_P2_InstQueue_reg[12][1]/NET0131  & n26313 ;
  assign n26503 = ~n26494 & ~n26495 ;
  assign n26496 = \P2_P2_InstQueue_reg[10][1]/NET0131  & n26320 ;
  assign n26497 = \P2_P2_InstQueue_reg[3][1]/NET0131  & n26332 ;
  assign n26504 = ~n26496 & ~n26497 ;
  assign n26505 = n26503 & n26504 ;
  assign n26488 = \P2_P2_InstQueue_reg[13][1]/NET0131  & n26336 ;
  assign n26489 = \P2_P2_InstQueue_reg[1][1]/NET0131  & n26338 ;
  assign n26501 = ~n26488 & ~n26489 ;
  assign n26490 = \P2_P2_InstQueue_reg[5][1]/NET0131  & n26318 ;
  assign n26492 = \P2_P2_InstQueue_reg[7][1]/NET0131  & n26327 ;
  assign n26502 = ~n26490 & ~n26492 ;
  assign n26506 = n26501 & n26502 ;
  assign n26484 = \P2_P2_InstQueue_reg[2][1]/NET0131  & n26316 ;
  assign n26485 = \P2_P2_InstQueue_reg[11][1]/NET0131  & n26310 ;
  assign n26499 = ~n26484 & ~n26485 ;
  assign n26486 = \P2_P2_InstQueue_reg[9][1]/NET0131  & n26304 ;
  assign n26487 = \P2_P2_InstQueue_reg[8][1]/NET0131  & n26334 ;
  assign n26500 = ~n26486 & ~n26487 ;
  assign n26507 = n26499 & n26500 ;
  assign n26510 = n26506 & n26507 ;
  assign n26511 = n26505 & n26510 ;
  assign n26512 = n26509 & n26511 ;
  assign n26580 = n26481 & n26512 ;
  assign n26525 = \P2_P2_InstQueue_reg[14][0]/NET0131  & n26330 ;
  assign n26523 = \P2_P2_InstQueue_reg[15][0]/NET0131  & n26325 ;
  assign n26514 = \P2_P2_InstQueue_reg[6][0]/NET0131  & n26300 ;
  assign n26515 = \P2_P2_InstQueue_reg[9][0]/NET0131  & n26304 ;
  assign n26530 = ~n26514 & ~n26515 ;
  assign n26540 = ~n26523 & n26530 ;
  assign n26541 = ~n26525 & n26540 ;
  assign n26526 = \P2_P2_InstQueue_reg[11][0]/NET0131  & n26310 ;
  assign n26527 = \P2_P2_InstQueue_reg[8][0]/NET0131  & n26334 ;
  assign n26535 = ~n26526 & ~n26527 ;
  assign n26528 = \P2_P2_InstQueue_reg[13][0]/NET0131  & n26336 ;
  assign n26529 = \P2_P2_InstQueue_reg[1][0]/NET0131  & n26338 ;
  assign n26536 = ~n26528 & ~n26529 ;
  assign n26537 = n26535 & n26536 ;
  assign n26520 = \P2_P2_InstQueue_reg[5][0]/NET0131  & n26318 ;
  assign n26521 = \P2_P2_InstQueue_reg[10][0]/NET0131  & n26320 ;
  assign n26533 = ~n26520 & ~n26521 ;
  assign n26522 = \P2_P2_InstQueue_reg[0][0]/NET0131  & n26322 ;
  assign n26524 = \P2_P2_InstQueue_reg[7][0]/NET0131  & n26327 ;
  assign n26534 = ~n26522 & ~n26524 ;
  assign n26538 = n26533 & n26534 ;
  assign n26516 = \P2_P2_InstQueue_reg[4][0]/NET0131  & n26307 ;
  assign n26517 = \P2_P2_InstQueue_reg[3][0]/NET0131  & n26332 ;
  assign n26531 = ~n26516 & ~n26517 ;
  assign n26518 = \P2_P2_InstQueue_reg[2][0]/NET0131  & n26316 ;
  assign n26519 = \P2_P2_InstQueue_reg[12][0]/NET0131  & n26313 ;
  assign n26532 = ~n26518 & ~n26519 ;
  assign n26539 = n26531 & n26532 ;
  assign n26542 = n26538 & n26539 ;
  assign n26543 = n26537 & n26542 ;
  assign n26544 = n26541 & n26543 ;
  assign n26557 = \P2_P2_InstQueue_reg[14][3]/NET0131  & n26330 ;
  assign n26555 = \P2_P2_InstQueue_reg[15][3]/NET0131  & n26325 ;
  assign n26546 = \P2_P2_InstQueue_reg[6][3]/NET0131  & n26300 ;
  assign n26547 = \P2_P2_InstQueue_reg[9][3]/NET0131  & n26304 ;
  assign n26562 = ~n26546 & ~n26547 ;
  assign n26572 = ~n26555 & n26562 ;
  assign n26573 = ~n26557 & n26572 ;
  assign n26558 = \P2_P2_InstQueue_reg[11][3]/NET0131  & n26310 ;
  assign n26559 = \P2_P2_InstQueue_reg[8][3]/NET0131  & n26334 ;
  assign n26567 = ~n26558 & ~n26559 ;
  assign n26560 = \P2_P2_InstQueue_reg[13][3]/NET0131  & n26336 ;
  assign n26561 = \P2_P2_InstQueue_reg[1][3]/NET0131  & n26338 ;
  assign n26568 = ~n26560 & ~n26561 ;
  assign n26569 = n26567 & n26568 ;
  assign n26552 = \P2_P2_InstQueue_reg[5][3]/NET0131  & n26318 ;
  assign n26553 = \P2_P2_InstQueue_reg[10][3]/NET0131  & n26320 ;
  assign n26565 = ~n26552 & ~n26553 ;
  assign n26554 = \P2_P2_InstQueue_reg[0][3]/NET0131  & n26322 ;
  assign n26556 = \P2_P2_InstQueue_reg[7][3]/NET0131  & n26327 ;
  assign n26566 = ~n26554 & ~n26556 ;
  assign n26570 = n26565 & n26566 ;
  assign n26548 = \P2_P2_InstQueue_reg[4][3]/NET0131  & n26307 ;
  assign n26549 = \P2_P2_InstQueue_reg[3][3]/NET0131  & n26332 ;
  assign n26563 = ~n26548 & ~n26549 ;
  assign n26550 = \P2_P2_InstQueue_reg[12][3]/NET0131  & n26313 ;
  assign n26551 = \P2_P2_InstQueue_reg[2][3]/NET0131  & n26316 ;
  assign n26564 = ~n26550 & ~n26551 ;
  assign n26571 = n26563 & n26564 ;
  assign n26574 = n26570 & n26571 ;
  assign n26575 = n26569 & n26574 ;
  assign n26576 = n26573 & n26575 ;
  assign n26668 = n26544 & n26576 ;
  assign n26669 = n26580 & n26668 ;
  assign n26430 = \P2_P2_InstQueue_reg[14][5]/NET0131  & n26330 ;
  assign n26428 = \P2_P2_InstQueue_reg[15][5]/NET0131  & n26325 ;
  assign n26419 = \P2_P2_InstQueue_reg[6][5]/NET0131  & n26300 ;
  assign n26420 = \P2_P2_InstQueue_reg[4][5]/NET0131  & n26307 ;
  assign n26435 = ~n26419 & ~n26420 ;
  assign n26445 = ~n26428 & n26435 ;
  assign n26446 = ~n26430 & n26445 ;
  assign n26431 = \P2_P2_InstQueue_reg[0][5]/NET0131  & n26322 ;
  assign n26432 = \P2_P2_InstQueue_reg[12][5]/NET0131  & n26313 ;
  assign n26440 = ~n26431 & ~n26432 ;
  assign n26433 = \P2_P2_InstQueue_reg[10][5]/NET0131  & n26320 ;
  assign n26434 = \P2_P2_InstQueue_reg[3][5]/NET0131  & n26332 ;
  assign n26441 = ~n26433 & ~n26434 ;
  assign n26442 = n26440 & n26441 ;
  assign n26425 = \P2_P2_InstQueue_reg[13][5]/NET0131  & n26336 ;
  assign n26426 = \P2_P2_InstQueue_reg[1][5]/NET0131  & n26338 ;
  assign n26438 = ~n26425 & ~n26426 ;
  assign n26427 = \P2_P2_InstQueue_reg[5][5]/NET0131  & n26318 ;
  assign n26429 = \P2_P2_InstQueue_reg[7][5]/NET0131  & n26327 ;
  assign n26439 = ~n26427 & ~n26429 ;
  assign n26443 = n26438 & n26439 ;
  assign n26421 = \P2_P2_InstQueue_reg[2][5]/NET0131  & n26316 ;
  assign n26422 = \P2_P2_InstQueue_reg[11][5]/NET0131  & n26310 ;
  assign n26436 = ~n26421 & ~n26422 ;
  assign n26423 = \P2_P2_InstQueue_reg[9][5]/NET0131  & n26304 ;
  assign n26424 = \P2_P2_InstQueue_reg[8][5]/NET0131  & n26334 ;
  assign n26437 = ~n26423 & ~n26424 ;
  assign n26444 = n26436 & n26437 ;
  assign n26447 = n26443 & n26444 ;
  assign n26448 = n26442 & n26447 ;
  assign n26449 = n26446 & n26448 ;
  assign n26331 = \P2_P2_InstQueue_reg[14][7]/NET0131  & n26330 ;
  assign n26326 = \P2_P2_InstQueue_reg[15][7]/NET0131  & n26325 ;
  assign n26301 = \P2_P2_InstQueue_reg[6][7]/NET0131  & n26300 ;
  assign n26305 = \P2_P2_InstQueue_reg[9][7]/NET0131  & n26304 ;
  assign n26340 = ~n26301 & ~n26305 ;
  assign n26350 = ~n26326 & n26340 ;
  assign n26351 = ~n26331 & n26350 ;
  assign n26333 = \P2_P2_InstQueue_reg[3][7]/NET0131  & n26332 ;
  assign n26335 = \P2_P2_InstQueue_reg[8][7]/NET0131  & n26334 ;
  assign n26345 = ~n26333 & ~n26335 ;
  assign n26337 = \P2_P2_InstQueue_reg[13][7]/NET0131  & n26336 ;
  assign n26339 = \P2_P2_InstQueue_reg[1][7]/NET0131  & n26338 ;
  assign n26346 = ~n26337 & ~n26339 ;
  assign n26347 = n26345 & n26346 ;
  assign n26319 = \P2_P2_InstQueue_reg[5][7]/NET0131  & n26318 ;
  assign n26321 = \P2_P2_InstQueue_reg[10][7]/NET0131  & n26320 ;
  assign n26343 = ~n26319 & ~n26321 ;
  assign n26323 = \P2_P2_InstQueue_reg[0][7]/NET0131  & n26322 ;
  assign n26328 = \P2_P2_InstQueue_reg[7][7]/NET0131  & n26327 ;
  assign n26344 = ~n26323 & ~n26328 ;
  assign n26348 = n26343 & n26344 ;
  assign n26308 = \P2_P2_InstQueue_reg[4][7]/NET0131  & n26307 ;
  assign n26311 = \P2_P2_InstQueue_reg[11][7]/NET0131  & n26310 ;
  assign n26341 = ~n26308 & ~n26311 ;
  assign n26314 = \P2_P2_InstQueue_reg[12][7]/NET0131  & n26313 ;
  assign n26317 = \P2_P2_InstQueue_reg[2][7]/NET0131  & n26316 ;
  assign n26342 = ~n26314 & ~n26317 ;
  assign n26349 = n26341 & n26342 ;
  assign n26352 = n26348 & n26349 ;
  assign n26353 = n26347 & n26352 ;
  assign n26354 = n26351 & n26353 ;
  assign n26366 = \P2_P2_InstQueue_reg[14][6]/NET0131  & n26330 ;
  assign n26364 = \P2_P2_InstQueue_reg[15][6]/NET0131  & n26325 ;
  assign n26355 = \P2_P2_InstQueue_reg[6][6]/NET0131  & n26300 ;
  assign n26356 = \P2_P2_InstQueue_reg[5][6]/NET0131  & n26318 ;
  assign n26371 = ~n26355 & ~n26356 ;
  assign n26381 = ~n26364 & n26371 ;
  assign n26382 = ~n26366 & n26381 ;
  assign n26367 = \P2_P2_InstQueue_reg[3][6]/NET0131  & n26332 ;
  assign n26368 = \P2_P2_InstQueue_reg[4][6]/NET0131  & n26307 ;
  assign n26376 = ~n26367 & ~n26368 ;
  assign n26369 = \P2_P2_InstQueue_reg[13][6]/NET0131  & n26336 ;
  assign n26370 = \P2_P2_InstQueue_reg[9][6]/NET0131  & n26304 ;
  assign n26377 = ~n26369 & ~n26370 ;
  assign n26378 = n26376 & n26377 ;
  assign n26361 = \P2_P2_InstQueue_reg[2][6]/NET0131  & n26316 ;
  assign n26362 = \P2_P2_InstQueue_reg[8][6]/NET0131  & n26334 ;
  assign n26374 = ~n26361 & ~n26362 ;
  assign n26363 = \P2_P2_InstQueue_reg[10][6]/NET0131  & n26320 ;
  assign n26365 = \P2_P2_InstQueue_reg[7][6]/NET0131  & n26327 ;
  assign n26375 = ~n26363 & ~n26365 ;
  assign n26379 = n26374 & n26375 ;
  assign n26357 = \P2_P2_InstQueue_reg[1][6]/NET0131  & n26338 ;
  assign n26358 = \P2_P2_InstQueue_reg[11][6]/NET0131  & n26310 ;
  assign n26372 = ~n26357 & ~n26358 ;
  assign n26359 = \P2_P2_InstQueue_reg[12][6]/NET0131  & n26313 ;
  assign n26360 = \P2_P2_InstQueue_reg[0][6]/NET0131  & n26322 ;
  assign n26373 = ~n26359 & ~n26360 ;
  assign n26380 = n26372 & n26373 ;
  assign n26383 = n26379 & n26380 ;
  assign n26384 = n26378 & n26383 ;
  assign n26385 = n26382 & n26384 ;
  assign n26613 = ~n26354 & ~n26385 ;
  assign n26677 = n26449 & n26613 ;
  assign n26678 = n26669 & n26677 ;
  assign n26513 = n26481 & ~n26512 ;
  assign n26545 = n26513 & ~n26544 ;
  assign n26577 = n26545 & ~n26576 ;
  assign n26386 = ~n26354 & n26385 ;
  assign n26398 = \P2_P2_InstQueue_reg[14][4]/NET0131  & n26330 ;
  assign n26396 = \P2_P2_InstQueue_reg[15][4]/NET0131  & n26325 ;
  assign n26387 = \P2_P2_InstQueue_reg[6][4]/NET0131  & n26300 ;
  assign n26388 = \P2_P2_InstQueue_reg[9][4]/NET0131  & n26304 ;
  assign n26403 = ~n26387 & ~n26388 ;
  assign n26413 = ~n26396 & n26403 ;
  assign n26414 = ~n26398 & n26413 ;
  assign n26399 = \P2_P2_InstQueue_reg[2][4]/NET0131  & n26316 ;
  assign n26400 = \P2_P2_InstQueue_reg[4][4]/NET0131  & n26307 ;
  assign n26408 = ~n26399 & ~n26400 ;
  assign n26401 = \P2_P2_InstQueue_reg[1][4]/NET0131  & n26338 ;
  assign n26402 = \P2_P2_InstQueue_reg[12][4]/NET0131  & n26313 ;
  assign n26409 = ~n26401 & ~n26402 ;
  assign n26410 = n26408 & n26409 ;
  assign n26393 = \P2_P2_InstQueue_reg[11][4]/NET0131  & n26310 ;
  assign n26394 = \P2_P2_InstQueue_reg[3][4]/NET0131  & n26332 ;
  assign n26406 = ~n26393 & ~n26394 ;
  assign n26395 = \P2_P2_InstQueue_reg[10][4]/NET0131  & n26320 ;
  assign n26397 = \P2_P2_InstQueue_reg[7][4]/NET0131  & n26327 ;
  assign n26407 = ~n26395 & ~n26397 ;
  assign n26411 = n26406 & n26407 ;
  assign n26389 = \P2_P2_InstQueue_reg[0][4]/NET0131  & n26322 ;
  assign n26390 = \P2_P2_InstQueue_reg[8][4]/NET0131  & n26334 ;
  assign n26404 = ~n26389 & ~n26390 ;
  assign n26391 = \P2_P2_InstQueue_reg[13][4]/NET0131  & n26336 ;
  assign n26392 = \P2_P2_InstQueue_reg[5][4]/NET0131  & n26318 ;
  assign n26405 = ~n26391 & ~n26392 ;
  assign n26412 = n26404 & n26405 ;
  assign n26415 = n26411 & n26412 ;
  assign n26416 = n26410 & n26415 ;
  assign n26417 = n26414 & n26416 ;
  assign n26631 = n26417 & n26449 ;
  assign n26632 = n26386 & n26631 ;
  assign n26633 = n26577 & n26632 ;
  assign n26634 = ~n26481 & n26576 ;
  assign n26614 = n26417 & ~n26449 ;
  assign n26635 = n26544 & n26614 ;
  assign n26636 = n26634 & n26635 ;
  assign n26637 = n26613 & n26636 ;
  assign n26638 = n26512 & n26637 ;
  assign n26639 = ~n26633 & ~n26638 ;
  assign n26584 = ~\P2_P2_InstQueueRd_Addr_reg[3]/NET0131  & \P2_P2_InstQueueWr_Addr_reg[3]/NET0131  ;
  assign n26585 = \P2_P2_InstQueueRd_Addr_reg[3]/NET0131  & ~\P2_P2_InstQueueWr_Addr_reg[3]/NET0131  ;
  assign n26587 = ~\P2_P2_InstQueueRd_Addr_reg[2]/NET0131  & \P2_P2_InstQueueWr_Addr_reg[2]/NET0131  ;
  assign n26588 = \P2_P2_InstQueueRd_Addr_reg[2]/NET0131  & ~\P2_P2_InstQueueWr_Addr_reg[2]/NET0131  ;
  assign n26589 = ~\P2_P2_InstQueueRd_Addr_reg[1]/NET0131  & \P2_P2_InstQueueWr_Addr_reg[1]/NET0131  ;
  assign n26590 = \P2_P2_InstQueueRd_Addr_reg[1]/NET0131  & ~\P2_P2_InstQueueWr_Addr_reg[1]/NET0131  ;
  assign n26591 = \P2_P2_InstQueueRd_Addr_reg[0]/NET0131  & ~\P2_P2_InstQueueWr_Addr_reg[0]/NET0131  ;
  assign n26592 = ~n26590 & ~n26591 ;
  assign n26593 = ~n26589 & ~n26592 ;
  assign n26594 = ~n26588 & ~n26593 ;
  assign n26595 = ~n26587 & ~n26594 ;
  assign n26609 = ~n26585 & ~n26595 ;
  assign n26610 = ~n26584 & ~n26609 ;
  assign n26586 = ~n26584 & ~n26585 ;
  assign n26596 = n26586 & n26595 ;
  assign n26597 = ~n26586 & ~n26595 ;
  assign n26598 = ~n26596 & ~n26597 ;
  assign n26599 = ~n26587 & ~n26588 ;
  assign n26600 = n26593 & n26599 ;
  assign n26601 = ~n26593 & ~n26599 ;
  assign n26602 = ~n26600 & ~n26601 ;
  assign n26622 = n26598 & n26602 ;
  assign n26623 = ~n26610 & ~n26622 ;
  assign n26603 = ~n26589 & ~n26590 ;
  assign n26624 = n26591 & ~n26603 ;
  assign n26625 = ~n26591 & n26603 ;
  assign n26626 = ~n26624 & ~n26625 ;
  assign n26627 = ~n26610 & n26626 ;
  assign n26640 = ~n26623 & ~n26627 ;
  assign n26697 = ~n26639 & ~n26640 ;
  assign n26646 = ~\P2_P2_State_reg[0]/NET0131  & \P2_P2_State_reg[1]/NET0131  ;
  assign n26647 = ~\P2_P2_State_reg[2]/NET0131  & n26646 ;
  assign n26648 = ~\P2_P2_State_reg[0]/NET0131  & ~\P2_P2_State_reg[1]/NET0131  ;
  assign n26649 = \P2_P2_State_reg[2]/NET0131  & n26648 ;
  assign n26650 = ~n26647 & ~n26649 ;
  assign n26616 = ~n26544 & ~n26576 ;
  assign n26617 = n26580 & n26616 ;
  assign n26643 = n26617 & n26632 ;
  assign n26644 = ~n26512 & n26637 ;
  assign n26645 = ~n26643 & ~n26644 ;
  assign n26698 = ~n26640 & ~n26645 ;
  assign n26699 = ~n26650 & n26698 ;
  assign n26700 = ~n26697 & ~n26699 ;
  assign n26723 = ~n26678 & n26700 ;
  assign n26286 = \P2_ready12_reg/NET0131  & \P2_ready21_reg/NET0131  ;
  assign n26724 = n26286 & ~n26678 ;
  assign n26725 = ~n26723 & ~n26724 ;
  assign n26726 = n26701 & n26725 ;
  assign n26727 = ~\P2_P2_InstQueueRd_Addr_reg[3]/NET0131  & ~n26726 ;
  assign n26729 = n26286 & ~n26700 ;
  assign n26730 = n26329 & ~n26729 ;
  assign n26731 = ~n26723 & ~n26730 ;
  assign n26728 = ~n26639 & n26640 ;
  assign n26615 = n26613 & n26614 ;
  assign n26618 = n26615 & n26617 ;
  assign n26621 = n26577 & n26615 ;
  assign n26676 = ~n26618 & ~n26621 ;
  assign n26692 = ~n26640 & ~n26650 ;
  assign n26693 = ~n26645 & ~n26692 ;
  assign n26732 = n26676 & ~n26693 ;
  assign n26733 = ~n26728 & n26732 ;
  assign n26734 = ~n26731 & n26733 ;
  assign n26735 = ~n26727 & ~n26734 ;
  assign n26659 = n26354 & n26631 ;
  assign n26660 = ~n26385 & n26659 ;
  assign n26661 = n26545 & n26576 ;
  assign n26662 = n26660 & n26661 ;
  assign n26663 = n26354 & ~n26385 ;
  assign n26664 = ~n26512 & n26663 ;
  assign n26665 = n26636 & n26664 ;
  assign n26666 = ~n26662 & ~n26665 ;
  assign n26679 = ~n26637 & ~n26643 ;
  assign n26680 = ~n26633 & n26679 ;
  assign n26681 = ~n26678 & n26680 ;
  assign n26682 = n26676 & n26681 ;
  assign n26418 = n26386 & ~n26417 ;
  assign n26450 = n26418 & ~n26449 ;
  assign n26578 = n26450 & n26577 ;
  assign n26579 = n26544 & ~n26576 ;
  assign n26581 = n26579 & n26580 ;
  assign n26582 = n26450 & n26581 ;
  assign n26583 = ~n26578 & ~n26582 ;
  assign n26683 = n26583 & n26666 ;
  assign n26684 = n26682 & n26683 ;
  assign n26667 = ~n26418 & ~n26660 ;
  assign n26670 = ~n26667 & n26669 ;
  assign n26671 = n26513 & n26579 ;
  assign n26672 = n26615 & n26671 ;
  assign n26673 = n26385 & n26512 ;
  assign n26674 = n26634 & n26673 ;
  assign n26675 = n26659 & n26674 ;
  assign n26685 = ~n26672 & ~n26675 ;
  assign n26686 = ~n26670 & n26685 ;
  assign n26687 = ~n26684 & n26686 ;
  assign n26688 = n26666 & n26687 ;
  assign n26720 = \P2_P2_InstQueueRd_Addr_reg[3]/NET0131  & ~n26324 ;
  assign n26721 = ~n26327 & ~n26720 ;
  assign n26722 = ~n26688 & ~n26721 ;
  assign n26604 = ~\P2_P2_InstQueueRd_Addr_reg[0]/NET0131  & \P2_P2_InstQueueWr_Addr_reg[0]/NET0131  ;
  assign n26605 = ~n26591 & ~n26604 ;
  assign n26606 = n26603 & n26605 ;
  assign n26607 = ~n26602 & ~n26606 ;
  assign n26608 = n26598 & ~n26607 ;
  assign n26611 = ~n26608 & ~n26610 ;
  assign n26689 = ~\P2_P2_InstQueueRd_Addr_reg[2]/NET0131  & ~n26309 ;
  assign n26736 = n26611 & ~n26689 ;
  assign n26737 = ~\P2_P2_InstQueueRd_Addr_reg[3]/NET0131  & ~n26736 ;
  assign n26738 = \P2_P2_InstQueueRd_Addr_reg[3]/NET0131  & n26736 ;
  assign n26739 = ~n26737 & ~n26738 ;
  assign n26740 = ~n26583 & n26739 ;
  assign n26741 = ~n26722 & ~n26740 ;
  assign n26742 = ~n26735 & n26741 ;
  assign n26752 = \P2_P2_InstQueueWr_Addr_reg[3]/NET0131  & n26742 ;
  assign n26756 = ~n26306 & ~n26309 ;
  assign n26757 = ~n26583 & n26611 ;
  assign n26758 = n26666 & ~n26757 ;
  assign n26759 = n26687 & n26758 ;
  assign n26760 = n26756 & ~n26759 ;
  assign n26641 = ~n26286 & ~n26640 ;
  assign n26761 = ~n26639 & n26641 ;
  assign n26762 = ~n26678 & ~n26761 ;
  assign n26651 = ~n26286 & ~n26650 ;
  assign n26763 = n26651 & n26698 ;
  assign n26764 = n26762 & ~n26763 ;
  assign n26765 = ~\P2_P2_InstQueueRd_Addr_reg[1]/NET0131  & n26764 ;
  assign n26612 = ~n26583 & ~n26611 ;
  assign n26652 = ~n26640 & n26651 ;
  assign n26653 = ~n26645 & ~n26652 ;
  assign n26766 = ~n26612 & ~n26653 ;
  assign n26642 = ~n26639 & ~n26641 ;
  assign n26694 = ~n26642 & n26676 ;
  assign n26767 = \P2_P2_InstQueueRd_Addr_reg[1]/NET0131  & n26694 ;
  assign n26768 = n26766 & n26767 ;
  assign n26769 = ~n26765 & ~n26768 ;
  assign n26770 = ~n26760 & ~n26769 ;
  assign n26771 = ~\P2_P2_InstQueueWr_Addr_reg[1]/NET0131  & ~n26770 ;
  assign n26772 = ~\P2_P2_InstQueueRd_Addr_reg[0]/NET0131  & n26759 ;
  assign n26773 = \P2_P2_InstQueueRd_Addr_reg[0]/NET0131  & ~n26612 ;
  assign n26774 = n26682 & n26773 ;
  assign n26775 = ~n26772 & ~n26774 ;
  assign n26776 = \P2_P2_InstQueueWr_Addr_reg[0]/NET0131  & ~n26775 ;
  assign n26777 = ~n26771 & n26776 ;
  assign n26690 = ~n26324 & ~n26689 ;
  assign n26691 = ~n26688 & n26690 ;
  assign n26702 = ~\P2_P2_InstQueueRd_Addr_reg[1]/NET0131  & ~\P2_P2_InstQueueRd_Addr_reg[2]/NET0131  ;
  assign n26703 = ~n26701 & ~n26702 ;
  assign n26704 = ~n26286 & ~n26703 ;
  assign n26705 = ~\P2_P2_InstQueueRd_Addr_reg[2]/NET0131  & n26286 ;
  assign n26706 = ~n26704 & ~n26705 ;
  assign n26707 = ~n26700 & n26706 ;
  assign n26695 = ~n26693 & n26694 ;
  assign n26696 = \P2_P2_InstQueueRd_Addr_reg[2]/NET0131  & ~n26695 ;
  assign n26708 = ~\P2_P2_InstQueueRd_Addr_reg[1]/NET0131  & ~n26639 ;
  assign n26709 = ~n26678 & ~n26708 ;
  assign n26710 = n26703 & ~n26709 ;
  assign n26711 = ~\P2_P2_InstQueueRd_Addr_reg[2]/NET0131  & ~n26611 ;
  assign n26712 = n26611 & n26690 ;
  assign n26713 = ~n26711 & ~n26712 ;
  assign n26714 = ~n26583 & n26713 ;
  assign n26715 = ~n26710 & ~n26714 ;
  assign n26716 = ~n26696 & n26715 ;
  assign n26717 = ~n26707 & n26716 ;
  assign n26718 = ~n26691 & n26717 ;
  assign n26755 = \P2_P2_InstQueueWr_Addr_reg[2]/NET0131  & n26718 ;
  assign n26778 = \P2_P2_InstQueueWr_Addr_reg[1]/NET0131  & n26770 ;
  assign n26779 = ~n26755 & ~n26778 ;
  assign n26780 = ~n26777 & n26779 ;
  assign n26781 = ~n26752 & n26780 ;
  assign n26753 = ~\P2_P2_InstQueueWr_Addr_reg[2]/NET0131  & ~n26718 ;
  assign n26754 = ~n26752 & n26753 ;
  assign n26719 = \P2_P2_InstQueueWr_Addr_reg[3]/NET0131  & n26718 ;
  assign n26743 = ~n26719 & ~n26742 ;
  assign n26654 = ~n26642 & ~n26653 ;
  assign n26655 = ~\P2_P2_More_reg/NET0131  & ~n26640 ;
  assign n26656 = ~n26654 & ~n26655 ;
  assign n26619 = ~n26611 & n26618 ;
  assign n26620 = ~n26612 & ~n26619 ;
  assign n26628 = ~n26605 & n26627 ;
  assign n26629 = ~n26623 & ~n26628 ;
  assign n26630 = n26621 & n26629 ;
  assign n26657 = n26620 & ~n26630 ;
  assign n26658 = ~n26656 & n26657 ;
  assign n26745 = n26286 & n26697 ;
  assign n26746 = ~n26651 & n26698 ;
  assign n26747 = ~n26745 & ~n26746 ;
  assign n26748 = \P2_P2_Flush_reg/NET0131  & ~n26747 ;
  assign n26744 = n26611 & n26618 ;
  assign n26749 = n26621 & ~n26629 ;
  assign n26750 = ~n26744 & ~n26749 ;
  assign n26751 = ~n26748 & n26750 ;
  assign n26782 = n26658 & n26751 ;
  assign n26783 = ~n26743 & n26782 ;
  assign n26784 = ~n26754 & n26783 ;
  assign n26785 = ~n26781 & n26784 ;
  assign n26786 = ~n26640 & n26643 ;
  assign n26787 = ~\P2_P2_DataWidth_reg[1]/NET0131  & n26786 ;
  assign n26788 = n26651 & n26787 ;
  assign n26789 = n26785 & ~n26788 ;
  assign n26790 = \P2_P2_State2_reg[0]/NET0131  & ~\P2_P2_State2_reg[3]/NET0131  ;
  assign n26791 = ~\P2_P2_State2_reg[1]/NET0131  & \P2_P2_State2_reg[2]/NET0131  ;
  assign n26792 = n26790 & n26791 ;
  assign n26793 = ~n26789 & n26792 ;
  assign n26285 = ~\P2_P2_State2_reg[0]/NET0131  & ~\P2_P2_State2_reg[3]/NET0131  ;
  assign n26287 = \P2_P2_State2_reg[1]/NET0131  & \P2_P2_State2_reg[2]/NET0131  ;
  assign n26288 = n26286 & n26287 ;
  assign n26289 = n26285 & n26288 ;
  assign n26290 = ~\P2_P2_State2_reg[1]/NET0131  & ~\P2_P2_State2_reg[2]/NET0131  ;
  assign n26291 = \P2_P2_State2_reg[0]/NET0131  & n26290 ;
  assign n26292 = ~\P2_P2_State2_reg[3]/NET0131  & n26291 ;
  assign n26293 = ~n26286 & n26292 ;
  assign n26796 = ~n26289 & ~n26293 ;
  assign n26294 = \P2_P2_State2_reg[1]/NET0131  & ~\P2_P2_State2_reg[2]/NET0131  ;
  assign n26295 = ~\P2_P2_State2_reg[3]/NET0131  & n26294 ;
  assign n26296 = \P2_P2_State2_reg[0]/NET0131  & n26295 ;
  assign n26297 = n26286 & n26296 ;
  assign n26794 = ~\P2_P2_State2_reg[0]/NET0131  & n26295 ;
  assign n26795 = ~\P2_P2_DataWidth_reg[1]/NET0131  & n26794 ;
  assign n26797 = ~n26297 & ~n26795 ;
  assign n26798 = n26796 & n26797 ;
  assign n26799 = ~n26793 & n26798 ;
  assign n26801 = ~n26286 & n26296 ;
  assign n26800 = \P2_P2_DataWidth_reg[1]/NET0131  & n26794 ;
  assign n26802 = \P2_P2_State2_reg[2]/NET0131  & n26285 ;
  assign n26803 = ~n26792 & ~n26802 ;
  assign n26804 = ~n26800 & n26803 ;
  assign n26805 = ~n26801 & n26804 ;
  assign n26835 = \P2_P3_InstQueueRd_Addr_reg[0]/NET0131  & \P2_P3_InstQueueRd_Addr_reg[1]/NET0131  ;
  assign n26836 = \P2_P3_InstQueueRd_Addr_reg[2]/NET0131  & n26835 ;
  assign n26837 = \P2_P3_InstQueueRd_Addr_reg[3]/NET0131  & n26836 ;
  assign n26838 = \P2_P3_InstQueue_reg[15][5]/NET0131  & n26837 ;
  assign n26810 = ~\P2_P3_InstQueueRd_Addr_reg[2]/NET0131  & ~\P2_P3_InstQueueRd_Addr_reg[3]/NET0131  ;
  assign n26811 = ~\P2_P3_InstQueueRd_Addr_reg[0]/NET0131  & ~\P2_P3_InstQueueRd_Addr_reg[1]/NET0131  ;
  assign n26812 = n26810 & n26811 ;
  assign n26813 = \P2_P3_InstQueue_reg[0][5]/NET0131  & n26812 ;
  assign n26814 = \P2_P3_InstQueueRd_Addr_reg[2]/NET0131  & ~\P2_P3_InstQueueRd_Addr_reg[3]/NET0131  ;
  assign n26815 = n26811 & n26814 ;
  assign n26816 = \P2_P3_InstQueue_reg[4][5]/NET0131  & n26815 ;
  assign n26851 = ~n26813 & ~n26816 ;
  assign n26860 = ~n26838 & n26851 ;
  assign n26839 = ~\P2_P3_InstQueueRd_Addr_reg[3]/NET0131  & n26836 ;
  assign n26840 = \P2_P3_InstQueue_reg[7][5]/NET0131  & n26839 ;
  assign n26806 = \P2_P3_InstQueueRd_Addr_reg[1]/NET0131  & \P2_P3_InstQueueRd_Addr_reg[2]/NET0131  ;
  assign n26808 = \P2_P3_InstQueueRd_Addr_reg[3]/NET0131  & n26806 ;
  assign n26845 = ~\P2_P3_InstQueueRd_Addr_reg[0]/NET0131  & n26808 ;
  assign n26846 = \P2_P3_InstQueue_reg[14][5]/NET0131  & n26845 ;
  assign n26861 = ~n26840 & ~n26846 ;
  assign n26862 = n26860 & n26861 ;
  assign n26817 = ~\P2_P3_InstQueueRd_Addr_reg[2]/NET0131  & \P2_P3_InstQueueRd_Addr_reg[3]/NET0131  ;
  assign n26849 = n26817 & n26835 ;
  assign n26850 = \P2_P3_InstQueue_reg[11][5]/NET0131  & n26849 ;
  assign n26818 = ~\P2_P3_InstQueueRd_Addr_reg[0]/NET0131  & \P2_P3_InstQueueRd_Addr_reg[1]/NET0131  ;
  assign n26843 = n26810 & n26818 ;
  assign n26844 = \P2_P3_InstQueue_reg[2][5]/NET0131  & n26843 ;
  assign n26847 = n26810 & n26835 ;
  assign n26848 = \P2_P3_InstQueue_reg[3][5]/NET0131  & n26847 ;
  assign n26856 = ~n26844 & ~n26848 ;
  assign n26857 = ~n26850 & n26856 ;
  assign n26824 = \P2_P3_InstQueueRd_Addr_reg[2]/NET0131  & \P2_P3_InstQueueRd_Addr_reg[3]/NET0131  ;
  assign n26829 = n26811 & n26824 ;
  assign n26830 = \P2_P3_InstQueue_reg[12][5]/NET0131  & n26829 ;
  assign n26821 = \P2_P3_InstQueueRd_Addr_reg[0]/NET0131  & ~\P2_P3_InstQueueRd_Addr_reg[1]/NET0131  ;
  assign n26831 = n26810 & n26821 ;
  assign n26832 = \P2_P3_InstQueue_reg[1][5]/NET0131  & n26831 ;
  assign n26854 = ~n26830 & ~n26832 ;
  assign n26833 = n26817 & n26821 ;
  assign n26834 = \P2_P3_InstQueue_reg[9][5]/NET0131  & n26833 ;
  assign n26841 = n26814 & n26818 ;
  assign n26842 = \P2_P3_InstQueue_reg[6][5]/NET0131  & n26841 ;
  assign n26855 = ~n26834 & ~n26842 ;
  assign n26858 = n26854 & n26855 ;
  assign n26819 = n26817 & n26818 ;
  assign n26820 = \P2_P3_InstQueue_reg[10][5]/NET0131  & n26819 ;
  assign n26822 = n26814 & n26821 ;
  assign n26823 = \P2_P3_InstQueue_reg[5][5]/NET0131  & n26822 ;
  assign n26852 = ~n26820 & ~n26823 ;
  assign n26825 = n26821 & n26824 ;
  assign n26826 = \P2_P3_InstQueue_reg[13][5]/NET0131  & n26825 ;
  assign n26827 = n26811 & n26817 ;
  assign n26828 = \P2_P3_InstQueue_reg[8][5]/NET0131  & n26827 ;
  assign n26853 = ~n26826 & ~n26828 ;
  assign n26859 = n26852 & n26853 ;
  assign n26863 = n26858 & n26859 ;
  assign n26864 = n26857 & n26863 ;
  assign n26865 = n26862 & n26864 ;
  assign n27070 = \P2_P3_InstQueue_reg[15][4]/NET0131  & n26837 ;
  assign n27061 = \P2_P3_InstQueue_reg[11][4]/NET0131  & n26849 ;
  assign n27062 = \P2_P3_InstQueue_reg[0][4]/NET0131  & n26812 ;
  assign n27077 = ~n27061 & ~n27062 ;
  assign n27086 = ~n27070 & n27077 ;
  assign n27071 = \P2_P3_InstQueue_reg[7][4]/NET0131  & n26839 ;
  assign n27074 = \P2_P3_InstQueue_reg[14][4]/NET0131  & n26845 ;
  assign n27087 = ~n27071 & ~n27074 ;
  assign n27088 = n27086 & n27087 ;
  assign n27076 = \P2_P3_InstQueue_reg[10][4]/NET0131  & n26819 ;
  assign n27073 = \P2_P3_InstQueue_reg[2][4]/NET0131  & n26843 ;
  assign n27075 = \P2_P3_InstQueue_reg[5][4]/NET0131  & n26822 ;
  assign n27082 = ~n27073 & ~n27075 ;
  assign n27083 = ~n27076 & n27082 ;
  assign n27067 = \P2_P3_InstQueue_reg[8][4]/NET0131  & n26827 ;
  assign n27068 = \P2_P3_InstQueue_reg[4][4]/NET0131  & n26815 ;
  assign n27080 = ~n27067 & ~n27068 ;
  assign n27069 = \P2_P3_InstQueue_reg[3][4]/NET0131  & n26847 ;
  assign n27072 = \P2_P3_InstQueue_reg[6][4]/NET0131  & n26841 ;
  assign n27081 = ~n27069 & ~n27072 ;
  assign n27084 = n27080 & n27081 ;
  assign n27063 = \P2_P3_InstQueue_reg[9][4]/NET0131  & n26833 ;
  assign n27064 = \P2_P3_InstQueue_reg[1][4]/NET0131  & n26831 ;
  assign n27078 = ~n27063 & ~n27064 ;
  assign n27065 = \P2_P3_InstQueue_reg[13][4]/NET0131  & n26825 ;
  assign n27066 = \P2_P3_InstQueue_reg[12][4]/NET0131  & n26829 ;
  assign n27079 = ~n27065 & ~n27066 ;
  assign n27085 = n27078 & n27079 ;
  assign n27089 = n27084 & n27085 ;
  assign n27090 = n27083 & n27089 ;
  assign n27091 = n27088 & n27090 ;
  assign n26875 = \P2_P3_InstQueue_reg[15][7]/NET0131  & n26837 ;
  assign n26866 = \P2_P3_InstQueue_reg[11][7]/NET0131  & n26849 ;
  assign n26867 = \P2_P3_InstQueue_reg[0][7]/NET0131  & n26812 ;
  assign n26882 = ~n26866 & ~n26867 ;
  assign n26891 = ~n26875 & n26882 ;
  assign n26876 = \P2_P3_InstQueue_reg[7][7]/NET0131  & n26839 ;
  assign n26879 = \P2_P3_InstQueue_reg[14][7]/NET0131  & n26845 ;
  assign n26892 = ~n26876 & ~n26879 ;
  assign n26893 = n26891 & n26892 ;
  assign n26881 = \P2_P3_InstQueue_reg[10][7]/NET0131  & n26819 ;
  assign n26878 = \P2_P3_InstQueue_reg[2][7]/NET0131  & n26843 ;
  assign n26880 = \P2_P3_InstQueue_reg[5][7]/NET0131  & n26822 ;
  assign n26887 = ~n26878 & ~n26880 ;
  assign n26888 = ~n26881 & n26887 ;
  assign n26872 = \P2_P3_InstQueue_reg[8][7]/NET0131  & n26827 ;
  assign n26873 = \P2_P3_InstQueue_reg[4][7]/NET0131  & n26815 ;
  assign n26885 = ~n26872 & ~n26873 ;
  assign n26874 = \P2_P3_InstQueue_reg[12][7]/NET0131  & n26829 ;
  assign n26877 = \P2_P3_InstQueue_reg[6][7]/NET0131  & n26841 ;
  assign n26886 = ~n26874 & ~n26877 ;
  assign n26889 = n26885 & n26886 ;
  assign n26868 = \P2_P3_InstQueue_reg[9][7]/NET0131  & n26833 ;
  assign n26869 = \P2_P3_InstQueue_reg[1][7]/NET0131  & n26831 ;
  assign n26883 = ~n26868 & ~n26869 ;
  assign n26870 = \P2_P3_InstQueue_reg[13][7]/NET0131  & n26825 ;
  assign n26871 = \P2_P3_InstQueue_reg[3][7]/NET0131  & n26847 ;
  assign n26884 = ~n26870 & ~n26871 ;
  assign n26890 = n26883 & n26884 ;
  assign n26894 = n26889 & n26890 ;
  assign n26895 = n26888 & n26894 ;
  assign n26896 = n26893 & n26895 ;
  assign n26906 = \P2_P3_InstQueue_reg[15][6]/NET0131  & n26837 ;
  assign n26897 = \P2_P3_InstQueue_reg[11][6]/NET0131  & n26849 ;
  assign n26898 = \P2_P3_InstQueue_reg[4][6]/NET0131  & n26815 ;
  assign n26913 = ~n26897 & ~n26898 ;
  assign n26922 = ~n26906 & n26913 ;
  assign n26907 = \P2_P3_InstQueue_reg[7][6]/NET0131  & n26839 ;
  assign n26910 = \P2_P3_InstQueue_reg[14][6]/NET0131  & n26845 ;
  assign n26923 = ~n26907 & ~n26910 ;
  assign n26924 = n26922 & n26923 ;
  assign n26912 = \P2_P3_InstQueue_reg[13][6]/NET0131  & n26825 ;
  assign n26909 = \P2_P3_InstQueue_reg[2][6]/NET0131  & n26843 ;
  assign n26911 = \P2_P3_InstQueue_reg[5][6]/NET0131  & n26822 ;
  assign n26918 = ~n26909 & ~n26911 ;
  assign n26919 = ~n26912 & n26918 ;
  assign n26903 = \P2_P3_InstQueue_reg[8][6]/NET0131  & n26827 ;
  assign n26904 = \P2_P3_InstQueue_reg[10][6]/NET0131  & n26819 ;
  assign n26916 = ~n26903 & ~n26904 ;
  assign n26905 = \P2_P3_InstQueue_reg[3][6]/NET0131  & n26847 ;
  assign n26908 = \P2_P3_InstQueue_reg[6][6]/NET0131  & n26841 ;
  assign n26917 = ~n26905 & ~n26908 ;
  assign n26920 = n26916 & n26917 ;
  assign n26899 = \P2_P3_InstQueue_reg[0][6]/NET0131  & n26812 ;
  assign n26900 = \P2_P3_InstQueue_reg[1][6]/NET0131  & n26831 ;
  assign n26914 = ~n26899 & ~n26900 ;
  assign n26901 = \P2_P3_InstQueue_reg[9][6]/NET0131  & n26833 ;
  assign n26902 = \P2_P3_InstQueue_reg[12][6]/NET0131  & n26829 ;
  assign n26915 = ~n26901 & ~n26902 ;
  assign n26921 = n26914 & n26915 ;
  assign n26925 = n26920 & n26921 ;
  assign n26926 = n26919 & n26925 ;
  assign n26927 = n26924 & n26926 ;
  assign n27102 = ~n26896 & n26927 ;
  assign n27103 = ~n27091 & n27102 ;
  assign n27104 = ~n26865 & n27103 ;
  assign n27032 = \P2_P3_InstQueue_reg[14][3]/NET0131  & n26845 ;
  assign n27024 = \P2_P3_InstQueue_reg[13][3]/NET0131  & n26825 ;
  assign n27025 = \P2_P3_InstQueue_reg[3][3]/NET0131  & n26847 ;
  assign n27040 = ~n27024 & ~n27025 ;
  assign n27049 = ~n27032 & n27040 ;
  assign n27034 = \P2_P3_InstQueue_reg[15][3]/NET0131  & n26837 ;
  assign n27035 = \P2_P3_InstQueue_reg[7][3]/NET0131  & n26839 ;
  assign n27050 = ~n27034 & ~n27035 ;
  assign n27051 = n27049 & n27050 ;
  assign n27039 = \P2_P3_InstQueue_reg[8][3]/NET0131  & n26827 ;
  assign n27037 = \P2_P3_InstQueue_reg[5][3]/NET0131  & n26822 ;
  assign n27038 = \P2_P3_InstQueue_reg[11][3]/NET0131  & n26849 ;
  assign n27045 = ~n27037 & ~n27038 ;
  assign n27046 = ~n27039 & n27045 ;
  assign n27030 = \P2_P3_InstQueue_reg[4][3]/NET0131  & n26815 ;
  assign n27031 = \P2_P3_InstQueue_reg[10][3]/NET0131  & n26819 ;
  assign n27043 = ~n27030 & ~n27031 ;
  assign n27033 = \P2_P3_InstQueue_reg[6][3]/NET0131  & n26841 ;
  assign n27036 = \P2_P3_InstQueue_reg[9][3]/NET0131  & n26833 ;
  assign n27044 = ~n27033 & ~n27036 ;
  assign n27047 = n27043 & n27044 ;
  assign n27026 = \P2_P3_InstQueue_reg[2][3]/NET0131  & n26843 ;
  assign n27027 = \P2_P3_InstQueue_reg[1][3]/NET0131  & n26831 ;
  assign n27041 = ~n27026 & ~n27027 ;
  assign n27028 = \P2_P3_InstQueue_reg[12][3]/NET0131  & n26829 ;
  assign n27029 = \P2_P3_InstQueue_reg[0][3]/NET0131  & n26812 ;
  assign n27042 = ~n27028 & ~n27029 ;
  assign n27048 = n27041 & n27042 ;
  assign n27052 = n27047 & n27048 ;
  assign n27053 = n27046 & n27052 ;
  assign n27054 = n27051 & n27053 ;
  assign n27000 = \P2_P3_InstQueue_reg[14][0]/NET0131  & n26845 ;
  assign n26992 = \P2_P3_InstQueue_reg[13][0]/NET0131  & n26825 ;
  assign n26993 = \P2_P3_InstQueue_reg[3][0]/NET0131  & n26847 ;
  assign n27008 = ~n26992 & ~n26993 ;
  assign n27017 = ~n27000 & n27008 ;
  assign n27002 = \P2_P3_InstQueue_reg[15][0]/NET0131  & n26837 ;
  assign n27003 = \P2_P3_InstQueue_reg[7][0]/NET0131  & n26839 ;
  assign n27018 = ~n27002 & ~n27003 ;
  assign n27019 = n27017 & n27018 ;
  assign n27007 = \P2_P3_InstQueue_reg[8][0]/NET0131  & n26827 ;
  assign n27005 = \P2_P3_InstQueue_reg[1][0]/NET0131  & n26831 ;
  assign n27006 = \P2_P3_InstQueue_reg[11][0]/NET0131  & n26849 ;
  assign n27013 = ~n27005 & ~n27006 ;
  assign n27014 = ~n27007 & n27013 ;
  assign n26998 = \P2_P3_InstQueue_reg[4][0]/NET0131  & n26815 ;
  assign n26999 = \P2_P3_InstQueue_reg[10][0]/NET0131  & n26819 ;
  assign n27011 = ~n26998 & ~n26999 ;
  assign n27001 = \P2_P3_InstQueue_reg[6][0]/NET0131  & n26841 ;
  assign n27004 = \P2_P3_InstQueue_reg[9][0]/NET0131  & n26833 ;
  assign n27012 = ~n27001 & ~n27004 ;
  assign n27015 = n27011 & n27012 ;
  assign n26994 = \P2_P3_InstQueue_reg[2][0]/NET0131  & n26843 ;
  assign n26995 = \P2_P3_InstQueue_reg[5][0]/NET0131  & n26822 ;
  assign n27009 = ~n26994 & ~n26995 ;
  assign n26996 = \P2_P3_InstQueue_reg[12][0]/NET0131  & n26829 ;
  assign n26997 = \P2_P3_InstQueue_reg[0][0]/NET0131  & n26812 ;
  assign n27010 = ~n26996 & ~n26997 ;
  assign n27016 = n27009 & n27010 ;
  assign n27020 = n27015 & n27016 ;
  assign n27021 = n27014 & n27020 ;
  assign n27022 = n27019 & n27021 ;
  assign n26938 = \P2_P3_InstQueue_reg[15][2]/NET0131  & n26837 ;
  assign n26929 = \P2_P3_InstQueue_reg[11][2]/NET0131  & n26849 ;
  assign n26930 = \P2_P3_InstQueue_reg[0][2]/NET0131  & n26812 ;
  assign n26945 = ~n26929 & ~n26930 ;
  assign n26954 = ~n26938 & n26945 ;
  assign n26939 = \P2_P3_InstQueue_reg[7][2]/NET0131  & n26839 ;
  assign n26942 = \P2_P3_InstQueue_reg[14][2]/NET0131  & n26845 ;
  assign n26955 = ~n26939 & ~n26942 ;
  assign n26956 = n26954 & n26955 ;
  assign n26944 = \P2_P3_InstQueue_reg[10][2]/NET0131  & n26819 ;
  assign n26941 = \P2_P3_InstQueue_reg[2][2]/NET0131  & n26843 ;
  assign n26943 = \P2_P3_InstQueue_reg[5][2]/NET0131  & n26822 ;
  assign n26950 = ~n26941 & ~n26943 ;
  assign n26951 = ~n26944 & n26950 ;
  assign n26935 = \P2_P3_InstQueue_reg[8][2]/NET0131  & n26827 ;
  assign n26936 = \P2_P3_InstQueue_reg[4][2]/NET0131  & n26815 ;
  assign n26948 = ~n26935 & ~n26936 ;
  assign n26937 = \P2_P3_InstQueue_reg[3][2]/NET0131  & n26847 ;
  assign n26940 = \P2_P3_InstQueue_reg[6][2]/NET0131  & n26841 ;
  assign n26949 = ~n26937 & ~n26940 ;
  assign n26952 = n26948 & n26949 ;
  assign n26931 = \P2_P3_InstQueue_reg[9][2]/NET0131  & n26833 ;
  assign n26932 = \P2_P3_InstQueue_reg[1][2]/NET0131  & n26831 ;
  assign n26946 = ~n26931 & ~n26932 ;
  assign n26933 = \P2_P3_InstQueue_reg[13][2]/NET0131  & n26825 ;
  assign n26934 = \P2_P3_InstQueue_reg[12][2]/NET0131  & n26829 ;
  assign n26947 = ~n26933 & ~n26934 ;
  assign n26953 = n26946 & n26947 ;
  assign n26957 = n26952 & n26953 ;
  assign n26958 = n26951 & n26957 ;
  assign n26959 = n26956 & n26958 ;
  assign n26969 = \P2_P3_InstQueue_reg[15][1]/NET0131  & n26837 ;
  assign n26960 = \P2_P3_InstQueue_reg[11][1]/NET0131  & n26849 ;
  assign n26961 = \P2_P3_InstQueue_reg[0][1]/NET0131  & n26812 ;
  assign n26976 = ~n26960 & ~n26961 ;
  assign n26985 = ~n26969 & n26976 ;
  assign n26970 = \P2_P3_InstQueue_reg[7][1]/NET0131  & n26839 ;
  assign n26973 = \P2_P3_InstQueue_reg[14][1]/NET0131  & n26845 ;
  assign n26986 = ~n26970 & ~n26973 ;
  assign n26987 = n26985 & n26986 ;
  assign n26975 = \P2_P3_InstQueue_reg[10][1]/NET0131  & n26819 ;
  assign n26972 = \P2_P3_InstQueue_reg[2][1]/NET0131  & n26843 ;
  assign n26974 = \P2_P3_InstQueue_reg[5][1]/NET0131  & n26822 ;
  assign n26981 = ~n26972 & ~n26974 ;
  assign n26982 = ~n26975 & n26981 ;
  assign n26966 = \P2_P3_InstQueue_reg[8][1]/NET0131  & n26827 ;
  assign n26967 = \P2_P3_InstQueue_reg[4][1]/NET0131  & n26815 ;
  assign n26979 = ~n26966 & ~n26967 ;
  assign n26968 = \P2_P3_InstQueue_reg[3][1]/NET0131  & n26847 ;
  assign n26971 = \P2_P3_InstQueue_reg[6][1]/NET0131  & n26841 ;
  assign n26980 = ~n26968 & ~n26971 ;
  assign n26983 = n26979 & n26980 ;
  assign n26962 = \P2_P3_InstQueue_reg[9][1]/NET0131  & n26833 ;
  assign n26963 = \P2_P3_InstQueue_reg[1][1]/NET0131  & n26831 ;
  assign n26977 = ~n26962 & ~n26963 ;
  assign n26964 = \P2_P3_InstQueue_reg[13][1]/NET0131  & n26825 ;
  assign n26965 = \P2_P3_InstQueue_reg[12][1]/NET0131  & n26829 ;
  assign n26978 = ~n26964 & ~n26965 ;
  assign n26984 = n26977 & n26978 ;
  assign n26988 = n26983 & n26984 ;
  assign n26989 = n26982 & n26988 ;
  assign n26990 = n26987 & n26989 ;
  assign n27105 = n26959 & ~n26990 ;
  assign n27106 = ~n27022 & n27105 ;
  assign n27107 = ~n27054 & n27106 ;
  assign n27108 = n27104 & n27107 ;
  assign n26991 = n26959 & n26990 ;
  assign n27023 = n26991 & n27022 ;
  assign n27109 = n27023 & ~n27054 ;
  assign n27110 = n27104 & n27109 ;
  assign n27111 = ~n27108 & ~n27110 ;
  assign n27112 = ~n27022 & ~n27054 ;
  assign n27113 = n26991 & n27112 ;
  assign n26928 = ~n26896 & ~n26927 ;
  assign n27114 = ~n26865 & n27091 ;
  assign n27115 = n26928 & n27114 ;
  assign n27116 = n27113 & n27115 ;
  assign n27117 = n27107 & n27115 ;
  assign n27118 = ~n27116 & ~n27117 ;
  assign n27055 = n27023 & n27054 ;
  assign n27056 = n26865 & n26928 ;
  assign n27057 = n27055 & n27056 ;
  assign n27119 = n26865 & n27091 ;
  assign n27120 = n27102 & n27119 ;
  assign n27122 = n27107 & n27120 ;
  assign n27121 = n27113 & n27120 ;
  assign n27092 = ~n26959 & n27054 ;
  assign n27123 = n27022 & n27092 ;
  assign n27124 = n27115 & n27123 ;
  assign n27125 = ~n27121 & ~n27124 ;
  assign n27126 = ~n27122 & n27125 ;
  assign n27127 = ~n27057 & n27126 ;
  assign n27128 = n27118 & n27127 ;
  assign n27129 = n27111 & n27128 ;
  assign n27093 = ~n26865 & ~n26927 ;
  assign n27094 = ~n26990 & n27022 ;
  assign n27095 = n27093 & n27094 ;
  assign n27096 = n26865 & n26927 ;
  assign n27097 = n26990 & n27096 ;
  assign n27098 = ~n27095 & ~n27097 ;
  assign n27099 = n26896 & n27091 ;
  assign n27100 = n27092 & n27099 ;
  assign n27101 = ~n27098 & n27100 ;
  assign n27136 = n27022 & ~n27054 ;
  assign n27137 = n27105 & n27136 ;
  assign n27138 = n27115 & n27137 ;
  assign n27139 = ~n27101 & ~n27138 ;
  assign n27130 = n26896 & ~n26927 ;
  assign n27131 = n27119 & n27130 ;
  assign n27132 = n27054 & n27106 ;
  assign n27133 = n27131 & n27132 ;
  assign n27134 = ~n27103 & ~n27131 ;
  assign n27135 = n27055 & ~n27134 ;
  assign n27140 = ~n27133 & ~n27135 ;
  assign n27141 = n27139 & n27140 ;
  assign n27142 = ~n27129 & n27141 ;
  assign n27149 = ~\P2_P3_InstQueueRd_Addr_reg[3]/NET0131  & \P2_P3_InstQueueWr_Addr_reg[3]/NET0131  ;
  assign n27150 = \P2_P3_InstQueueRd_Addr_reg[3]/NET0131  & ~\P2_P3_InstQueueWr_Addr_reg[3]/NET0131  ;
  assign n27152 = ~\P2_P3_InstQueueRd_Addr_reg[2]/NET0131  & \P2_P3_InstQueueWr_Addr_reg[2]/NET0131  ;
  assign n27153 = \P2_P3_InstQueueRd_Addr_reg[2]/NET0131  & ~\P2_P3_InstQueueWr_Addr_reg[2]/NET0131  ;
  assign n27154 = ~\P2_P3_InstQueueRd_Addr_reg[1]/NET0131  & \P2_P3_InstQueueWr_Addr_reg[1]/NET0131  ;
  assign n27155 = \P2_P3_InstQueueRd_Addr_reg[0]/NET0131  & ~\P2_P3_InstQueueWr_Addr_reg[0]/NET0131  ;
  assign n27156 = \P2_P3_InstQueueRd_Addr_reg[1]/NET0131  & ~\P2_P3_InstQueueWr_Addr_reg[1]/NET0131  ;
  assign n27157 = ~n27155 & ~n27156 ;
  assign n27158 = ~n27154 & ~n27157 ;
  assign n27159 = ~n27153 & ~n27158 ;
  assign n27160 = ~n27152 & ~n27159 ;
  assign n27169 = ~n27150 & ~n27160 ;
  assign n27170 = ~n27149 & ~n27169 ;
  assign n27151 = ~n27149 & ~n27150 ;
  assign n27161 = n27151 & n27160 ;
  assign n27162 = ~n27151 & ~n27160 ;
  assign n27163 = ~n27161 & ~n27162 ;
  assign n27164 = ~n27152 & ~n27153 ;
  assign n27165 = n27158 & ~n27164 ;
  assign n27166 = ~n27158 & n27164 ;
  assign n27167 = ~n27165 & ~n27166 ;
  assign n27172 = ~n27154 & ~n27156 ;
  assign n27174 = ~n27155 & n27172 ;
  assign n27202 = ~\P2_P3_InstQueueRd_Addr_reg[0]/NET0131  & \P2_P3_InstQueueWr_Addr_reg[0]/NET0131  ;
  assign n27203 = n27174 & ~n27202 ;
  assign n27204 = n27167 & ~n27203 ;
  assign n27205 = n27163 & ~n27204 ;
  assign n27206 = ~n27170 & ~n27205 ;
  assign n27219 = ~n27111 & n27206 ;
  assign n27220 = n27142 & ~n27219 ;
  assign n27221 = ~n26811 & ~n26835 ;
  assign n27222 = ~n27220 & n27221 ;
  assign n27188 = ~\P2_P3_ADS_n_reg/NET0131  & \P2_P3_D_C_n_reg/NET0131  ;
  assign n27189 = \P2_P3_M_IO_n_reg/NET0131  & \P2_P3_W_R_n_reg/NET0131  ;
  assign n27190 = \P4_rd_reg/NET0131  & n27189 ;
  assign n27191 = n27188 & n27190 ;
  assign n27192 = \P2_ready22_reg/NET0131  & ~n27191 ;
  assign n27168 = n27163 & ~n27167 ;
  assign n27171 = ~n27168 & ~n27170 ;
  assign n27173 = n27155 & ~n27172 ;
  assign n27175 = ~n27173 & ~n27174 ;
  assign n27176 = ~n27170 & n27175 ;
  assign n27177 = ~n27171 & ~n27176 ;
  assign n27144 = ~\P2_P3_State_reg[0]/NET0131  & \P2_P3_State_reg[1]/NET0131  ;
  assign n27145 = ~\P2_P3_State_reg[2]/NET0131  & n27144 ;
  assign n27146 = ~\P2_P3_State_reg[0]/NET0131  & ~\P2_P3_State_reg[1]/NET0131  ;
  assign n27147 = \P2_P3_State_reg[2]/NET0131  & n27146 ;
  assign n27148 = ~n27145 & ~n27147 ;
  assign n27179 = ~n26990 & n27124 ;
  assign n27180 = ~n27121 & ~n27179 ;
  assign n27199 = ~n27148 & ~n27180 ;
  assign n27223 = ~n27177 & n27199 ;
  assign n27224 = ~n27192 & n27223 ;
  assign n27225 = ~n27057 & ~n27224 ;
  assign n27186 = n26990 & n27124 ;
  assign n27226 = ~n27122 & ~n27186 ;
  assign n27227 = ~n27177 & ~n27192 ;
  assign n27228 = ~n27226 & n27227 ;
  assign n27229 = n27225 & ~n27228 ;
  assign n27230 = ~\P2_P3_InstQueueRd_Addr_reg[1]/NET0131  & n27229 ;
  assign n27231 = ~n27111 & ~n27206 ;
  assign n27178 = ~n27148 & ~n27177 ;
  assign n27232 = n27178 & ~n27192 ;
  assign n27233 = ~n27180 & ~n27232 ;
  assign n27234 = ~n27226 & ~n27227 ;
  assign n27235 = ~n27233 & ~n27234 ;
  assign n27236 = ~n27231 & n27235 ;
  assign n27237 = \P2_P3_InstQueueRd_Addr_reg[1]/NET0131  & n27118 ;
  assign n27238 = n27236 & n27237 ;
  assign n27239 = ~n27230 & ~n27238 ;
  assign n27240 = ~n27222 & ~n27239 ;
  assign n27241 = ~\P2_P3_InstQueueWr_Addr_reg[1]/NET0131  & ~n27240 ;
  assign n27242 = ~\P2_P3_InstQueueRd_Addr_reg[0]/NET0131  & n27220 ;
  assign n27243 = \P2_P3_InstQueueRd_Addr_reg[0]/NET0131  & ~n27231 ;
  assign n27244 = n27128 & n27243 ;
  assign n27245 = ~n27242 & ~n27244 ;
  assign n27246 = \P2_P3_InstQueueWr_Addr_reg[0]/NET0131  & ~n27245 ;
  assign n27247 = ~n27241 & n27246 ;
  assign n27271 = \P2_P3_InstQueueWr_Addr_reg[1]/NET0131  & n27240 ;
  assign n27059 = \P2_P3_InstQueueRd_Addr_reg[3]/NET0131  & ~n26836 ;
  assign n27060 = ~n26839 & ~n27059 ;
  assign n27143 = ~n27060 & ~n27142 ;
  assign n27181 = ~n27178 & ~n27180 ;
  assign n27182 = n27118 & ~n27181 ;
  assign n27183 = n27122 & n27177 ;
  assign n27184 = n27182 & ~n27183 ;
  assign n27185 = \P2_P3_InstQueueRd_Addr_reg[3]/NET0131  & ~n27184 ;
  assign n26807 = ~\P2_P3_InstQueueRd_Addr_reg[3]/NET0131  & ~n26806 ;
  assign n26809 = ~n26807 & ~n26808 ;
  assign n27193 = ~n26809 & ~n27192 ;
  assign n27194 = ~\P2_P3_InstQueueRd_Addr_reg[3]/NET0131  & n27192 ;
  assign n27195 = ~n27193 & ~n27194 ;
  assign n27196 = ~n27177 & n27195 ;
  assign n27200 = ~n27122 & ~n27199 ;
  assign n27201 = n27196 & ~n27200 ;
  assign n27207 = ~\P2_P3_InstQueueRd_Addr_reg[2]/NET0131  & ~n26835 ;
  assign n27208 = n27206 & ~n27207 ;
  assign n27209 = ~\P2_P3_InstQueueRd_Addr_reg[3]/NET0131  & ~n27208 ;
  assign n27210 = \P2_P3_InstQueueRd_Addr_reg[3]/NET0131  & n27208 ;
  assign n27211 = ~n27209 & ~n27210 ;
  assign n27212 = ~n27111 & n27211 ;
  assign n27058 = n26809 & n27057 ;
  assign n27187 = \P2_P3_InstQueueRd_Addr_reg[3]/NET0131  & n27177 ;
  assign n27197 = ~n27187 & ~n27196 ;
  assign n27198 = n27186 & ~n27197 ;
  assign n27213 = ~n27058 & ~n27198 ;
  assign n27214 = ~n27212 & n27213 ;
  assign n27215 = ~n27201 & n27214 ;
  assign n27216 = ~n27185 & n27215 ;
  assign n27217 = ~n27143 & n27216 ;
  assign n27218 = \P2_P3_InstQueueWr_Addr_reg[3]/NET0131  & n27217 ;
  assign n27251 = ~n26836 & ~n27207 ;
  assign n27252 = ~n27142 & n27251 ;
  assign n27256 = ~n27177 & ~n27226 ;
  assign n27257 = ~n27223 & ~n27256 ;
  assign n27248 = ~\P2_P3_InstQueueRd_Addr_reg[1]/NET0131  & ~\P2_P3_InstQueueRd_Addr_reg[2]/NET0131  ;
  assign n27249 = ~n26806 & ~n27248 ;
  assign n27258 = ~n27192 & ~n27249 ;
  assign n27259 = ~\P2_P3_InstQueueRd_Addr_reg[2]/NET0131  & n27192 ;
  assign n27260 = ~n27258 & ~n27259 ;
  assign n27261 = ~n27257 & n27260 ;
  assign n27253 = n27177 & ~n27226 ;
  assign n27254 = n27182 & ~n27253 ;
  assign n27255 = \P2_P3_InstQueueRd_Addr_reg[2]/NET0131  & ~n27254 ;
  assign n27250 = n27057 & n27249 ;
  assign n27262 = ~\P2_P3_InstQueueRd_Addr_reg[2]/NET0131  & ~n27206 ;
  assign n27263 = n27206 & n27251 ;
  assign n27264 = ~n27262 & ~n27263 ;
  assign n27265 = ~n27111 & n27264 ;
  assign n27266 = ~n27250 & ~n27265 ;
  assign n27267 = ~n27255 & n27266 ;
  assign n27268 = ~n27261 & n27267 ;
  assign n27269 = ~n27252 & n27268 ;
  assign n27270 = \P2_P3_InstQueueWr_Addr_reg[2]/NET0131  & n27269 ;
  assign n27272 = ~n27218 & ~n27270 ;
  assign n27273 = ~n27271 & n27272 ;
  assign n27274 = ~n27247 & n27273 ;
  assign n27289 = \P2_P3_InstQueueWr_Addr_reg[3]/NET0131  & n27269 ;
  assign n27290 = ~n27217 & ~n27289 ;
  assign n27287 = ~\P2_P3_InstQueueWr_Addr_reg[2]/NET0131  & ~n27218 ;
  assign n27288 = ~n27269 & n27287 ;
  assign n27275 = n27148 & ~n27180 ;
  assign n27276 = ~n27192 & ~n27275 ;
  assign n27277 = ~n27126 & ~n27177 ;
  assign n27278 = \P2_P3_Flush_reg/NET0131  & n27277 ;
  assign n27279 = ~n27276 & n27278 ;
  assign n27280 = n27116 & n27206 ;
  assign n27281 = ~n27172 & ~n27202 ;
  assign n27282 = ~n27171 & n27281 ;
  assign n27283 = ~n27177 & ~n27282 ;
  assign n27284 = n27117 & n27283 ;
  assign n27285 = ~n27280 & ~n27284 ;
  assign n27286 = ~n27279 & n27285 ;
  assign n27291 = ~\P2_P3_More_reg/NET0131  & ~n27177 ;
  assign n27292 = ~n27235 & ~n27291 ;
  assign n27293 = n27117 & ~n27283 ;
  assign n27294 = n27116 & ~n27206 ;
  assign n27295 = ~n27231 & ~n27294 ;
  assign n27296 = ~n27293 & n27295 ;
  assign n27297 = ~n27292 & n27296 ;
  assign n27298 = n27286 & n27297 ;
  assign n27299 = ~n27288 & n27298 ;
  assign n27300 = ~n27290 & n27299 ;
  assign n27301 = ~n27274 & n27300 ;
  assign n27302 = ~\P2_P3_DataWidth_reg[1]/NET0131  & ~n27192 ;
  assign n27303 = n27121 & n27178 ;
  assign n27304 = n27302 & n27303 ;
  assign n27305 = n27301 & ~n27304 ;
  assign n27306 = \P2_P3_State2_reg[0]/NET0131  & ~\P2_P3_State2_reg[3]/NET0131  ;
  assign n27307 = ~\P2_P3_State2_reg[1]/NET0131  & \P2_P3_State2_reg[2]/NET0131  ;
  assign n27308 = n27306 & n27307 ;
  assign n27309 = ~n27305 & n27308 ;
  assign n27310 = ~\P2_P3_State2_reg[2]/NET0131  & n27306 ;
  assign n27317 = ~\P2_P3_State2_reg[0]/NET0131  & ~\P2_P3_State2_reg[3]/NET0131  ;
  assign n27318 = \P2_P3_State2_reg[2]/NET0131  & n27317 ;
  assign n27319 = ~n27310 & ~n27318 ;
  assign n27320 = \P2_P3_State2_reg[1]/NET0131  & ~n27319 ;
  assign n27321 = n27192 & n27320 ;
  assign n27311 = ~\P2_P3_State2_reg[1]/NET0131  & n27310 ;
  assign n27312 = ~n27192 & n27311 ;
  assign n27313 = \P2_P3_State2_reg[1]/NET0131  & ~\P2_P3_State2_reg[2]/NET0131  ;
  assign n27314 = ~\P2_P3_State2_reg[3]/NET0131  & n27313 ;
  assign n27315 = ~\P2_P3_State2_reg[0]/NET0131  & n27314 ;
  assign n27316 = ~\P2_P3_DataWidth_reg[1]/NET0131  & n27315 ;
  assign n27322 = ~n27312 & ~n27316 ;
  assign n27323 = ~n27321 & n27322 ;
  assign n27324 = ~n27309 & n27323 ;
  assign n27326 = \P2_P3_State2_reg[0]/NET0131  & n27314 ;
  assign n27327 = ~n27192 & n27326 ;
  assign n27325 = \P2_P3_DataWidth_reg[1]/NET0131  & n27315 ;
  assign n27328 = ~n27308 & ~n27318 ;
  assign n27329 = ~n27325 & n27328 ;
  assign n27330 = ~n27327 & n27329 ;
  assign n27331 = \P1_P1_EAX_reg[10]/NET0131  & ~n15326 ;
  assign n27332 = ~n15384 & n23580 ;
  assign n27333 = \P1_P1_EAX_reg[10]/NET0131  & ~n25291 ;
  assign n27334 = \P1_P1_InstQueue_reg[0][2]/NET0131  & n8291 ;
  assign n27335 = \P1_P1_InstQueue_reg[5][2]/NET0131  & n8323 ;
  assign n27336 = \P1_P1_InstQueue_reg[4][2]/NET0131  & n8314 ;
  assign n27350 = ~n27335 & ~n27336 ;
  assign n27337 = \P1_P1_InstQueue_reg[6][2]/NET0131  & n8295 ;
  assign n27338 = \P1_P1_InstQueue_reg[12][2]/NET0131  & n8303 ;
  assign n27351 = ~n27337 & ~n27338 ;
  assign n27360 = n27350 & n27351 ;
  assign n27361 = ~n27334 & n27360 ;
  assign n27349 = \P1_P1_InstQueue_reg[7][2]/NET0131  & n8307 ;
  assign n27347 = \P1_P1_InstQueue_reg[10][2]/NET0131  & n8305 ;
  assign n27348 = \P1_P1_InstQueue_reg[2][2]/NET0131  & n8309 ;
  assign n27356 = ~n27347 & ~n27348 ;
  assign n27357 = ~n27349 & n27356 ;
  assign n27343 = \P1_P1_InstQueue_reg[8][2]/NET0131  & n8316 ;
  assign n27344 = \P1_P1_InstQueue_reg[9][2]/NET0131  & n8318 ;
  assign n27354 = ~n27343 & ~n27344 ;
  assign n27345 = \P1_P1_InstQueue_reg[1][2]/NET0131  & n8321 ;
  assign n27346 = \P1_P1_InstQueue_reg[15][2]/NET0131  & n8327 ;
  assign n27355 = ~n27345 & ~n27346 ;
  assign n27358 = n27354 & n27355 ;
  assign n27339 = \P1_P1_InstQueue_reg[13][2]/NET0131  & n8312 ;
  assign n27340 = \P1_P1_InstQueue_reg[14][2]/NET0131  & n8329 ;
  assign n27352 = ~n27339 & ~n27340 ;
  assign n27341 = \P1_P1_InstQueue_reg[11][2]/NET0131  & n8325 ;
  assign n27342 = \P1_P1_InstQueue_reg[3][2]/NET0131  & n8299 ;
  assign n27353 = ~n27341 & ~n27342 ;
  assign n27359 = n27352 & n27353 ;
  assign n27362 = n27358 & n27359 ;
  assign n27363 = n27357 & n27362 ;
  assign n27364 = n27361 & n27363 ;
  assign n27365 = n22818 & ~n27364 ;
  assign n27366 = n15396 & n25290 ;
  assign n27367 = ~n27365 & ~n27366 ;
  assign n27368 = ~n27333 & n27367 ;
  assign n27369 = ~n27332 & n27368 ;
  assign n27370 = n8355 & ~n27369 ;
  assign n27371 = ~n27331 & ~n27370 ;
  assign n27374 = ~\P2_P1_EAX_reg[13]/NET0131  & ~\P2_P1_EAX_reg[14]/NET0131  ;
  assign n27375 = ~\P2_P1_EAX_reg[15]/NET0131  & ~\P2_P1_EAX_reg[1]/NET0131  ;
  assign n27382 = n27374 & n27375 ;
  assign n27372 = ~\P2_P1_EAX_reg[0]/NET0131  & ~\P2_P1_EAX_reg[10]/NET0131  ;
  assign n27373 = ~\P2_P1_EAX_reg[11]/NET0131  & ~\P2_P1_EAX_reg[12]/NET0131  ;
  assign n27383 = n27372 & n27373 ;
  assign n27384 = n27382 & n27383 ;
  assign n27378 = ~\P2_P1_EAX_reg[6]/NET0131  & ~\P2_P1_EAX_reg[7]/NET0131  ;
  assign n27379 = ~\P2_P1_EAX_reg[8]/NET0131  & ~\P2_P1_EAX_reg[9]/NET0131  ;
  assign n27380 = n27378 & n27379 ;
  assign n27376 = ~\P2_P1_EAX_reg[2]/NET0131  & ~\P2_P1_EAX_reg[3]/NET0131  ;
  assign n27377 = ~\P2_P1_EAX_reg[4]/NET0131  & ~\P2_P1_EAX_reg[5]/NET0131  ;
  assign n27381 = n27376 & n27377 ;
  assign n27385 = n27380 & n27381 ;
  assign n27386 = n27384 & n27385 ;
  assign n27387 = \P2_P1_EAX_reg[31]/NET0131  & ~n27386 ;
  assign n27388 = \P2_P1_EAX_reg[16]/NET0131  & n27387 ;
  assign n27389 = \P2_P1_EAX_reg[17]/NET0131  & n27388 ;
  assign n27390 = \P2_P1_EAX_reg[18]/NET0131  & n27389 ;
  assign n27391 = \P2_P1_EAX_reg[19]/NET0131  & n27390 ;
  assign n27392 = \P2_P1_EAX_reg[20]/NET0131  & n27391 ;
  assign n27393 = \P2_P1_EAX_reg[21]/NET0131  & n27392 ;
  assign n27394 = \P2_P1_EAX_reg[22]/NET0131  & n27393 ;
  assign n27395 = \P2_P1_EAX_reg[23]/NET0131  & n27394 ;
  assign n27396 = \P2_P1_EAX_reg[24]/NET0131  & n27395 ;
  assign n27397 = \P2_P1_EAX_reg[25]/NET0131  & n27396 ;
  assign n27398 = \P2_P1_EAX_reg[26]/NET0131  & n27397 ;
  assign n27399 = \P2_P1_EAX_reg[27]/NET0131  & n27398 ;
  assign n27400 = \P2_P1_EAX_reg[28]/NET0131  & n27399 ;
  assign n27401 = \P2_P1_EAX_reg[29]/NET0131  & n27400 ;
  assign n27403 = \P2_P1_EAX_reg[30]/NET0131  & n27401 ;
  assign n27402 = ~\P2_P1_EAX_reg[30]/NET0131  & ~n27401 ;
  assign n27404 = n24898 & ~n27402 ;
  assign n27405 = ~n27403 & n27404 ;
  assign n27406 = ~n25158 & ~n27405 ;
  assign n27407 = ~n21081 & ~n27406 ;
  assign n27408 = \P2_P1_uWord_reg[14]/NET0131  & ~n25154 ;
  assign n27409 = ~n27407 & ~n27408 ;
  assign n27410 = n11623 & ~n27409 ;
  assign n27411 = \P2_P1_uWord_reg[14]/NET0131  & ~n24913 ;
  assign n27412 = ~n27410 & ~n27411 ;
  assign n27413 = \P1_P1_lWord_reg[11]/NET0131  & ~n25165 ;
  assign n27414 = \P1_P1_EAX_reg[11]/NET0131  & n24503 ;
  assign n27415 = n7974 & n23947 ;
  assign n27416 = ~n27414 & ~n27415 ;
  assign n27417 = n8355 & ~n27416 ;
  assign n27418 = ~n27413 & ~n27417 ;
  assign n27419 = \P1_P1_uWord_reg[13]/NET0131  & ~n24515 ;
  assign n27421 = \P1_P1_uWord_reg[13]/NET0131  & n25363 ;
  assign n27422 = ~n23187 & ~n27421 ;
  assign n27423 = n15334 & ~n27422 ;
  assign n27420 = \P1_P1_uWord_reg[13]/NET0131  & n24505 ;
  assign n27424 = n15410 & n25348 ;
  assign n27425 = \P1_P1_EAX_reg[25]/NET0131  & n27424 ;
  assign n27426 = \P1_P1_EAX_reg[26]/NET0131  & n27425 ;
  assign n27427 = \P1_P1_EAX_reg[27]/NET0131  & n27426 ;
  assign n27428 = \P1_P1_EAX_reg[28]/NET0131  & n27427 ;
  assign n27429 = ~\P1_P1_EAX_reg[29]/NET0131  & ~n27428 ;
  assign n27430 = \P1_P1_EAX_reg[29]/NET0131  & n27428 ;
  assign n27431 = ~n27429 & ~n27430 ;
  assign n27432 = n24503 & n27431 ;
  assign n27433 = ~n27420 & ~n27432 ;
  assign n27434 = ~n27423 & n27433 ;
  assign n27435 = n8355 & ~n27434 ;
  assign n27436 = ~n27419 & ~n27435 ;
  assign n27437 = n11623 & ~n24712 ;
  assign n27438 = n21100 & ~n27437 ;
  assign n27439 = \P2_P1_EAX_reg[10]/NET0131  & ~n27438 ;
  assign n27472 = n11373 & n24708 ;
  assign n27445 = \P2_P1_InstQueue_reg[8][2]/NET0131  & n11651 ;
  assign n27444 = \P2_P1_InstQueue_reg[1][2]/NET0131  & n11647 ;
  assign n27440 = \P2_P1_InstQueue_reg[4][2]/NET0131  & n11654 ;
  assign n27441 = \P2_P1_InstQueue_reg[7][2]/NET0131  & n11638 ;
  assign n27456 = ~n27440 & ~n27441 ;
  assign n27466 = ~n27444 & n27456 ;
  assign n27467 = ~n27445 & n27466 ;
  assign n27452 = \P2_P1_InstQueue_reg[13][2]/NET0131  & n11665 ;
  assign n27453 = \P2_P1_InstQueue_reg[5][2]/NET0131  & n11663 ;
  assign n27461 = ~n27452 & ~n27453 ;
  assign n27454 = \P2_P1_InstQueue_reg[3][2]/NET0131  & n11671 ;
  assign n27455 = \P2_P1_InstQueue_reg[11][2]/NET0131  & n11656 ;
  assign n27462 = ~n27454 & ~n27455 ;
  assign n27463 = n27461 & n27462 ;
  assign n27448 = \P2_P1_InstQueue_reg[12][2]/NET0131  & n11634 ;
  assign n27449 = \P2_P1_InstQueue_reg[9][2]/NET0131  & n11661 ;
  assign n27459 = ~n27448 & ~n27449 ;
  assign n27450 = \P2_P1_InstQueue_reg[10][2]/NET0131  & n11659 ;
  assign n27451 = \P2_P1_InstQueue_reg[6][2]/NET0131  & n11667 ;
  assign n27460 = ~n27450 & ~n27451 ;
  assign n27464 = n27459 & n27460 ;
  assign n27442 = \P2_P1_InstQueue_reg[14][2]/NET0131  & n11673 ;
  assign n27443 = \P2_P1_InstQueue_reg[0][2]/NET0131  & n11643 ;
  assign n27457 = ~n27442 & ~n27443 ;
  assign n27446 = \P2_P1_InstQueue_reg[2][2]/NET0131  & n11669 ;
  assign n27447 = \P2_P1_InstQueue_reg[15][2]/NET0131  & n11641 ;
  assign n27458 = ~n27446 & ~n27447 ;
  assign n27465 = n27457 & n27458 ;
  assign n27468 = n27464 & n27465 ;
  assign n27469 = n27463 & n27468 ;
  assign n27470 = n27467 & n27469 ;
  assign n27471 = n20728 & ~n27470 ;
  assign n27473 = ~\P2_P1_EAX_reg[10]/NET0131  & ~n21031 ;
  assign n27474 = ~n21032 & ~n27473 ;
  assign n27475 = n21022 & n27474 ;
  assign n27476 = ~n27471 & ~n27475 ;
  assign n27477 = ~n27472 & n27476 ;
  assign n27478 = n11623 & ~n27477 ;
  assign n27479 = ~n27439 & ~n27478 ;
  assign n27480 = n26102 & n26105 ;
  assign n27481 = n11623 & ~n27480 ;
  assign n27483 = ~\P2_P1_Flush_reg/NET0131  & \P2_P1_InstQueueRd_Addr_reg[2]/NET0131  ;
  assign n27484 = \P2_P1_InstQueueRd_Addr_reg[3]/NET0131  & ~n11658 ;
  assign n27485 = n27483 & n27484 ;
  assign n27486 = n21096 & ~n27485 ;
  assign n27487 = n11620 & n21073 ;
  assign n27488 = n11611 & ~n27487 ;
  assign n27482 = n21073 & n21098 ;
  assign n27489 = ~n11625 & ~n27482 ;
  assign n27490 = ~n27488 & n27489 ;
  assign n27491 = ~n27486 & n27490 ;
  assign n27492 = ~n27481 & n27491 ;
  assign n27493 = \P2_P1_EAX_reg[9]/NET0131  & ~n27438 ;
  assign n27526 = n11386 & n24708 ;
  assign n27499 = \P2_P1_InstQueue_reg[8][1]/NET0131  & n11651 ;
  assign n27498 = \P2_P1_InstQueue_reg[1][1]/NET0131  & n11647 ;
  assign n27494 = \P2_P1_InstQueue_reg[7][1]/NET0131  & n11638 ;
  assign n27495 = \P2_P1_InstQueue_reg[4][1]/NET0131  & n11654 ;
  assign n27510 = ~n27494 & ~n27495 ;
  assign n27520 = ~n27498 & n27510 ;
  assign n27521 = ~n27499 & n27520 ;
  assign n27506 = \P2_P1_InstQueue_reg[3][1]/NET0131  & n11671 ;
  assign n27507 = \P2_P1_InstQueue_reg[6][1]/NET0131  & n11667 ;
  assign n27515 = ~n27506 & ~n27507 ;
  assign n27508 = \P2_P1_InstQueue_reg[12][1]/NET0131  & n11634 ;
  assign n27509 = \P2_P1_InstQueue_reg[15][1]/NET0131  & n11641 ;
  assign n27516 = ~n27508 & ~n27509 ;
  assign n27517 = n27515 & n27516 ;
  assign n27502 = \P2_P1_InstQueue_reg[2][1]/NET0131  & n11669 ;
  assign n27503 = \P2_P1_InstQueue_reg[9][1]/NET0131  & n11661 ;
  assign n27513 = ~n27502 & ~n27503 ;
  assign n27504 = \P2_P1_InstQueue_reg[10][1]/NET0131  & n11659 ;
  assign n27505 = \P2_P1_InstQueue_reg[13][1]/NET0131  & n11665 ;
  assign n27514 = ~n27504 & ~n27505 ;
  assign n27518 = n27513 & n27514 ;
  assign n27496 = \P2_P1_InstQueue_reg[11][1]/NET0131  & n11656 ;
  assign n27497 = \P2_P1_InstQueue_reg[0][1]/NET0131  & n11643 ;
  assign n27511 = ~n27496 & ~n27497 ;
  assign n27500 = \P2_P1_InstQueue_reg[5][1]/NET0131  & n11663 ;
  assign n27501 = \P2_P1_InstQueue_reg[14][1]/NET0131  & n11673 ;
  assign n27512 = ~n27500 & ~n27501 ;
  assign n27519 = n27511 & n27512 ;
  assign n27522 = n27518 & n27519 ;
  assign n27523 = n27517 & n27522 ;
  assign n27524 = n27521 & n27523 ;
  assign n27525 = n20728 & ~n27524 ;
  assign n27527 = ~\P2_P1_EAX_reg[9]/NET0131  & ~n21030 ;
  assign n27528 = ~n21031 & ~n27527 ;
  assign n27529 = n21022 & n27528 ;
  assign n27530 = ~n27525 & ~n27529 ;
  assign n27531 = ~n27526 & n27530 ;
  assign n27532 = n11623 & ~n27531 ;
  assign n27533 = ~n27493 & ~n27532 ;
  assign n27534 = \P2_P1_lWord_reg[11]/NET0131  & ~n25156 ;
  assign n27535 = n11388 & n23167 ;
  assign n27536 = \P2_P1_EAX_reg[11]/NET0131  & n24898 ;
  assign n27537 = ~n27535 & ~n27536 ;
  assign n27538 = n25161 & ~n27537 ;
  assign n27539 = ~n27534 & ~n27538 ;
  assign n27540 = \P2_P1_uWord_reg[13]/NET0131  & ~n24913 ;
  assign n27542 = ~\P2_P1_EAX_reg[29]/NET0131  & ~n27400 ;
  assign n27543 = n24898 & ~n27401 ;
  assign n27544 = ~n27542 & n27543 ;
  assign n27545 = ~n21081 & n27544 ;
  assign n27541 = \P2_P1_uWord_reg[13]/NET0131  & ~n25154 ;
  assign n27546 = ~n23169 & ~n27541 ;
  assign n27547 = ~n27545 & n27546 ;
  assign n27548 = n11623 & ~n27547 ;
  assign n27549 = ~n27540 & ~n27548 ;
  assign n27550 = n8355 & ~n24346 ;
  assign n27551 = n15326 & ~n27550 ;
  assign n27552 = \P1_P1_EAX_reg[9]/NET0131  & ~n27551 ;
  assign n27553 = n7955 & n24342 ;
  assign n27554 = \P1_P1_InstQueue_reg[0][1]/NET0131  & n8291 ;
  assign n27555 = \P1_P1_InstQueue_reg[10][1]/NET0131  & n8305 ;
  assign n27556 = \P1_P1_InstQueue_reg[6][1]/NET0131  & n8295 ;
  assign n27570 = ~n27555 & ~n27556 ;
  assign n27557 = \P1_P1_InstQueue_reg[13][1]/NET0131  & n8312 ;
  assign n27558 = \P1_P1_InstQueue_reg[5][1]/NET0131  & n8323 ;
  assign n27571 = ~n27557 & ~n27558 ;
  assign n27580 = n27570 & n27571 ;
  assign n27581 = ~n27554 & n27580 ;
  assign n27569 = \P1_P1_InstQueue_reg[12][1]/NET0131  & n8303 ;
  assign n27567 = \P1_P1_InstQueue_reg[3][1]/NET0131  & n8299 ;
  assign n27568 = \P1_P1_InstQueue_reg[14][1]/NET0131  & n8329 ;
  assign n27576 = ~n27567 & ~n27568 ;
  assign n27577 = ~n27569 & n27576 ;
  assign n27563 = \P1_P1_InstQueue_reg[8][1]/NET0131  & n8316 ;
  assign n27564 = \P1_P1_InstQueue_reg[1][1]/NET0131  & n8321 ;
  assign n27574 = ~n27563 & ~n27564 ;
  assign n27565 = \P1_P1_InstQueue_reg[9][1]/NET0131  & n8318 ;
  assign n27566 = \P1_P1_InstQueue_reg[4][1]/NET0131  & n8314 ;
  assign n27575 = ~n27565 & ~n27566 ;
  assign n27578 = n27574 & n27575 ;
  assign n27559 = \P1_P1_InstQueue_reg[7][1]/NET0131  & n8307 ;
  assign n27560 = \P1_P1_InstQueue_reg[11][1]/NET0131  & n8325 ;
  assign n27572 = ~n27559 & ~n27560 ;
  assign n27561 = \P1_P1_InstQueue_reg[2][1]/NET0131  & n8309 ;
  assign n27562 = \P1_P1_InstQueue_reg[15][1]/NET0131  & n8327 ;
  assign n27573 = ~n27561 & ~n27562 ;
  assign n27579 = n27572 & n27573 ;
  assign n27582 = n27578 & n27579 ;
  assign n27583 = n27577 & n27582 ;
  assign n27584 = n27581 & n27583 ;
  assign n27585 = n22818 & ~n27584 ;
  assign n27586 = ~\P1_P1_EAX_reg[9]/NET0131  & ~n15395 ;
  assign n27587 = ~n15396 & ~n27586 ;
  assign n27588 = n15377 & n27587 ;
  assign n27589 = ~n27585 & ~n27588 ;
  assign n27590 = ~n27553 & n27589 ;
  assign n27591 = n8355 & ~n27590 ;
  assign n27592 = ~n27552 & ~n27591 ;
  assign n27593 = \P1_P1_uWord_reg[12]/NET0131  & ~n24515 ;
  assign n27598 = \P1_P1_uWord_reg[12]/NET0131  & n25363 ;
  assign n27599 = ~n22834 & ~n27598 ;
  assign n27600 = n15334 & ~n27599 ;
  assign n27595 = \P1_P1_EAX_reg[28]/NET0131  & n25357 ;
  assign n27594 = ~\P1_P1_EAX_reg[28]/NET0131  & ~n25357 ;
  assign n27596 = n24503 & ~n27594 ;
  assign n27597 = ~n27595 & n27596 ;
  assign n27601 = \P1_P1_uWord_reg[12]/NET0131  & n24505 ;
  assign n27602 = ~n27597 & ~n27601 ;
  assign n27603 = ~n27600 & n27602 ;
  assign n27604 = n8355 & ~n27603 ;
  assign n27605 = ~n27593 & ~n27604 ;
  assign n27606 = ~\P1_P2_State2_reg[1]/NET0131  & ~\P1_P2_State2_reg[2]/NET0131  ;
  assign n27607 = \P1_P2_State2_reg[3]/NET0131  & n27606 ;
  assign n27608 = ~\P1_P2_State2_reg[0]/NET0131  & n27607 ;
  assign n27609 = \P1_P2_State2_reg[0]/NET0131  & n25921 ;
  assign n27610 = ~n27608 & ~n27609 ;
  assign n27611 = ~n8350 & ~n15322 ;
  assign n27612 = \P2_P2_State2_reg[3]/NET0131  & n26290 ;
  assign n27613 = ~\P2_P2_State2_reg[0]/NET0131  & n27612 ;
  assign n27614 = ~\P2_P2_State2_reg[3]/NET0131  & n26287 ;
  assign n27615 = \P2_P2_State2_reg[0]/NET0131  & n27614 ;
  assign n27616 = ~n27613 & ~n27615 ;
  assign n27617 = n26273 & n26276 ;
  assign n27618 = n8355 & ~n27617 ;
  assign n27620 = ~\P1_P1_Flush_reg/NET0131  & \P1_P1_InstQueueRd_Addr_reg[2]/NET0131  ;
  assign n27621 = \P1_P1_InstQueueRd_Addr_reg[3]/NET0131  & ~n8293 ;
  assign n27622 = n27620 & n27621 ;
  assign n27623 = n15322 & ~n27622 ;
  assign n27624 = n8352 & n15335 ;
  assign n27625 = n8356 & ~n27624 ;
  assign n27619 = n15324 & n15335 ;
  assign n27626 = ~n8361 & ~n27619 ;
  assign n27627 = ~n27625 & n27626 ;
  assign n27628 = ~n27623 & n27627 ;
  assign n27629 = ~n27618 & n27628 ;
  assign n27630 = ~\P2_P2_DataWidth_reg[1]/NET0131  & n26652 ;
  assign n27631 = \P2_P2_State2_reg[0]/NET0131  & ~n27630 ;
  assign n27632 = n26643 & ~n27631 ;
  assign n27633 = n26785 & n27632 ;
  assign n27634 = n26792 & ~n27633 ;
  assign n27639 = ~\P2_P2_Flush_reg/NET0131  & \P2_P2_InstQueueRd_Addr_reg[2]/NET0131  ;
  assign n27640 = \P2_P2_InstQueueRd_Addr_reg[3]/NET0131  & ~n26306 ;
  assign n27641 = n27639 & n27640 ;
  assign n27642 = n27615 & ~n27641 ;
  assign n27638 = n26285 & ~n26288 ;
  assign n27635 = ~\P2_P2_State2_reg[2]/NET0131  & n26790 ;
  assign n27636 = n26286 & n27635 ;
  assign n27637 = \P2_P2_State2_reg[0]/NET0131  & n27612 ;
  assign n27643 = ~n27636 & ~n27637 ;
  assign n27644 = ~n27638 & n27643 ;
  assign n27645 = ~n27642 & n27644 ;
  assign n27646 = ~n27634 & n27645 ;
  assign n27647 = n27301 & n27304 ;
  assign n27648 = n27308 & ~n27647 ;
  assign n27653 = \P2_P3_State2_reg[1]/NET0131  & \P2_P3_State2_reg[2]/NET0131  ;
  assign n27654 = n27192 & n27653 ;
  assign n27655 = n27317 & ~n27654 ;
  assign n27652 = n27192 & n27310 ;
  assign n27649 = ~\P2_P3_State2_reg[1]/NET0131  & ~\P2_P3_State2_reg[2]/NET0131  ;
  assign n27650 = \P2_P3_State2_reg[3]/NET0131  & n27649 ;
  assign n27651 = \P2_P3_State2_reg[0]/NET0131  & n27650 ;
  assign n27656 = ~\P2_P3_State2_reg[3]/NET0131  & n27653 ;
  assign n27657 = \P2_P3_State2_reg[0]/NET0131  & n27656 ;
  assign n27658 = ~\P2_P3_Flush_reg/NET0131  & \P2_P3_InstQueueRd_Addr_reg[2]/NET0131  ;
  assign n27659 = \P2_P3_InstQueueRd_Addr_reg[3]/NET0131  & ~n26811 ;
  assign n27660 = n27658 & n27659 ;
  assign n27661 = n27657 & ~n27660 ;
  assign n27662 = ~n27651 & ~n27661 ;
  assign n27663 = ~n27652 & n27662 ;
  assign n27664 = ~n27655 & n27663 ;
  assign n27665 = ~n27648 & n27664 ;
  assign n27666 = n25913 & n25915 ;
  assign n27667 = n25918 & ~n27666 ;
  assign n27670 = ~\P1_P2_Flush_reg/NET0131  & \P1_P2_InstQueueRd_Addr_reg[2]/NET0131  ;
  assign n27671 = \P1_P2_InstQueueRd_Addr_reg[3]/NET0131  & ~n25421 ;
  assign n27672 = n27670 & n27671 ;
  assign n27673 = n27609 & ~n27672 ;
  assign n27675 = \P1_P2_State2_reg[0]/NET0131  & n27607 ;
  assign n27668 = n25415 & n25920 ;
  assign n27669 = n25934 & ~n27668 ;
  assign n27674 = n25415 & n25417 ;
  assign n27676 = ~n27669 & ~n27674 ;
  assign n27677 = ~n27675 & n27676 ;
  assign n27678 = ~n27673 & n27677 ;
  assign n27679 = ~n27667 & n27678 ;
  assign n27681 = \P2_P1_DataWidth_reg[1]/NET0131  & n11609 ;
  assign n27680 = n11627 & ~n21073 ;
  assign n27682 = ~n11623 & ~n25940 ;
  assign n27683 = ~n27680 & n27682 ;
  assign n27684 = ~n27681 & n27683 ;
  assign n27685 = \P2_P1_EAX_reg[8]/NET0131  & ~n27438 ;
  assign n27718 = ~n21069 & n23737 ;
  assign n27691 = \P2_P1_InstQueue_reg[8][0]/NET0131  & n11651 ;
  assign n27690 = \P2_P1_InstQueue_reg[1][0]/NET0131  & n11647 ;
  assign n27686 = \P2_P1_InstQueue_reg[4][0]/NET0131  & n11654 ;
  assign n27687 = \P2_P1_InstQueue_reg[7][0]/NET0131  & n11638 ;
  assign n27702 = ~n27686 & ~n27687 ;
  assign n27712 = ~n27690 & n27702 ;
  assign n27713 = ~n27691 & n27712 ;
  assign n27698 = \P2_P1_InstQueue_reg[13][0]/NET0131  & n11665 ;
  assign n27699 = \P2_P1_InstQueue_reg[5][0]/NET0131  & n11663 ;
  assign n27707 = ~n27698 & ~n27699 ;
  assign n27700 = \P2_P1_InstQueue_reg[3][0]/NET0131  & n11671 ;
  assign n27701 = \P2_P1_InstQueue_reg[11][0]/NET0131  & n11656 ;
  assign n27708 = ~n27700 & ~n27701 ;
  assign n27709 = n27707 & n27708 ;
  assign n27694 = \P2_P1_InstQueue_reg[12][0]/NET0131  & n11634 ;
  assign n27695 = \P2_P1_InstQueue_reg[9][0]/NET0131  & n11661 ;
  assign n27705 = ~n27694 & ~n27695 ;
  assign n27696 = \P2_P1_InstQueue_reg[10][0]/NET0131  & n11659 ;
  assign n27697 = \P2_P1_InstQueue_reg[6][0]/NET0131  & n11667 ;
  assign n27706 = ~n27696 & ~n27697 ;
  assign n27710 = n27705 & n27706 ;
  assign n27688 = \P2_P1_InstQueue_reg[14][0]/NET0131  & n11673 ;
  assign n27689 = \P2_P1_InstQueue_reg[0][0]/NET0131  & n11643 ;
  assign n27703 = ~n27688 & ~n27689 ;
  assign n27692 = \P2_P1_InstQueue_reg[2][0]/NET0131  & n11669 ;
  assign n27693 = \P2_P1_InstQueue_reg[15][0]/NET0131  & n11641 ;
  assign n27704 = ~n27692 & ~n27693 ;
  assign n27711 = n27703 & n27704 ;
  assign n27714 = n27710 & n27711 ;
  assign n27715 = n27709 & n27714 ;
  assign n27716 = n27713 & n27715 ;
  assign n27717 = n20728 & ~n27716 ;
  assign n27719 = ~\P2_P1_EAX_reg[8]/NET0131  & ~n21029 ;
  assign n27720 = ~n21030 & ~n27719 ;
  assign n27721 = n21022 & n27720 ;
  assign n27722 = ~n27717 & ~n27721 ;
  assign n27723 = ~n27718 & n27722 ;
  assign n27724 = n11623 & ~n27723 ;
  assign n27725 = ~n27685 & ~n27724 ;
  assign n27726 = \P2_P1_lWord_reg[10]/NET0131  & ~n25156 ;
  assign n27727 = \P2_P1_EAX_reg[10]/NET0131  & n24899 ;
  assign n27728 = ~n23830 & ~n27727 ;
  assign n27729 = n11623 & ~n27728 ;
  assign n27730 = ~n27726 & ~n27729 ;
  assign n27731 = ~\P2_P1_EAX_reg[28]/NET0131  & ~n27399 ;
  assign n27732 = ~n27400 & ~n27731 ;
  assign n27733 = n24898 & n27732 ;
  assign n27734 = ~n25283 & ~n27733 ;
  assign n27735 = ~n21081 & ~n27734 ;
  assign n27736 = \P2_P1_uWord_reg[12]/NET0131  & ~n25154 ;
  assign n27737 = ~n27735 & ~n27736 ;
  assign n27738 = n11623 & ~n27737 ;
  assign n27739 = \P2_P1_uWord_reg[12]/NET0131  & ~n24913 ;
  assign n27740 = ~n27738 & ~n27739 ;
  assign n27741 = \P1_P1_lWord_reg[10]/NET0131  & ~n25165 ;
  assign n27742 = \P1_P1_EAX_reg[10]/NET0131  & n24503 ;
  assign n27743 = ~n23581 & ~n27742 ;
  assign n27744 = n8355 & ~n27743 ;
  assign n27745 = ~n27741 & ~n27744 ;
  assign n27746 = \P1_P1_EAX_reg[8]/NET0131  & ~n27551 ;
  assign n27747 = ~n7891 & n24342 ;
  assign n27748 = \P1_P1_InstQueue_reg[0][0]/NET0131  & n8291 ;
  assign n27749 = \P1_P1_InstQueue_reg[5][0]/NET0131  & n8323 ;
  assign n27750 = \P1_P1_InstQueue_reg[2][0]/NET0131  & n8309 ;
  assign n27764 = ~n27749 & ~n27750 ;
  assign n27751 = \P1_P1_InstQueue_reg[7][0]/NET0131  & n8307 ;
  assign n27752 = \P1_P1_InstQueue_reg[15][0]/NET0131  & n8327 ;
  assign n27765 = ~n27751 & ~n27752 ;
  assign n27774 = n27764 & n27765 ;
  assign n27775 = ~n27748 & n27774 ;
  assign n27763 = \P1_P1_InstQueue_reg[14][0]/NET0131  & n8329 ;
  assign n27761 = \P1_P1_InstQueue_reg[12][0]/NET0131  & n8303 ;
  assign n27762 = \P1_P1_InstQueue_reg[10][0]/NET0131  & n8305 ;
  assign n27770 = ~n27761 & ~n27762 ;
  assign n27771 = ~n27763 & n27770 ;
  assign n27757 = \P1_P1_InstQueue_reg[8][0]/NET0131  & n8316 ;
  assign n27758 = \P1_P1_InstQueue_reg[9][0]/NET0131  & n8318 ;
  assign n27768 = ~n27757 & ~n27758 ;
  assign n27759 = \P1_P1_InstQueue_reg[1][0]/NET0131  & n8321 ;
  assign n27760 = \P1_P1_InstQueue_reg[11][0]/NET0131  & n8325 ;
  assign n27769 = ~n27759 & ~n27760 ;
  assign n27772 = n27768 & n27769 ;
  assign n27753 = \P1_P1_InstQueue_reg[4][0]/NET0131  & n8314 ;
  assign n27754 = \P1_P1_InstQueue_reg[6][0]/NET0131  & n8295 ;
  assign n27766 = ~n27753 & ~n27754 ;
  assign n27755 = \P1_P1_InstQueue_reg[13][0]/NET0131  & n8312 ;
  assign n27756 = \P1_P1_InstQueue_reg[3][0]/NET0131  & n8299 ;
  assign n27767 = ~n27755 & ~n27756 ;
  assign n27773 = n27766 & n27767 ;
  assign n27776 = n27772 & n27773 ;
  assign n27777 = n27771 & n27776 ;
  assign n27778 = n27775 & n27777 ;
  assign n27779 = n22818 & ~n27778 ;
  assign n27780 = ~\P1_P1_EAX_reg[8]/NET0131  & ~n15394 ;
  assign n27781 = ~n15395 & ~n27780 ;
  assign n27782 = n15377 & n27781 ;
  assign n27783 = ~n27779 & ~n27782 ;
  assign n27784 = ~n27747 & n27783 ;
  assign n27785 = n8355 & ~n27784 ;
  assign n27786 = ~n27746 & ~n27785 ;
  assign n27787 = ~n11692 & ~n21096 ;
  assign n27788 = ~\P2_P3_State2_reg[0]/NET0131  & n27650 ;
  assign n27789 = ~n27657 & ~n27788 ;
  assign n27792 = ~n15335 & n26115 ;
  assign n27791 = \P1_P1_DataWidth_reg[1]/NET0131  & n8282 ;
  assign n27790 = ~\P1_P1_State2_reg[0]/NET0131  & n8353 ;
  assign n27793 = ~n8286 & ~n27790 ;
  assign n27794 = ~n27791 & n27793 ;
  assign n27795 = ~n27792 & n27794 ;
  assign n27796 = ~\P3_rd_reg/NET0131  & \P4_reg3_reg[2]/NET0131  ;
  assign n27797 = \P4_addr_reg[2]/NET0131  & n15737 ;
  assign n27799 = \P4_IR_reg[0]/NET0131  & \P4_reg2_reg[0]/NET0131  ;
  assign n27798 = ~\P4_IR_reg[0]/NET0131  & ~\P4_reg2_reg[0]/NET0131  ;
  assign n27800 = n15733 & ~n27798 ;
  assign n27801 = ~n27799 & n27800 ;
  assign n27804 = ~\P4_IR_reg[27]/NET0131  & \P4_IR_reg[28]/NET0131  ;
  assign n27802 = \P4_IR_reg[0]/NET0131  & \P4_reg1_reg[0]/NET0131  ;
  assign n27803 = ~\P4_IR_reg[0]/NET0131  & ~\P4_reg1_reg[0]/NET0131  ;
  assign n27805 = ~n27802 & ~n27803 ;
  assign n27806 = n27804 & n27805 ;
  assign n27807 = ~n27801 & ~n27806 ;
  assign n27808 = \P4_IR_reg[0]/NET0131  & n21786 ;
  assign n27809 = ~n16102 & ~n27808 ;
  assign n27810 = n27807 & n27809 ;
  assign n27811 = n15736 & ~n27810 ;
  assign n27812 = ~n27797 & ~n27811 ;
  assign n27813 = ~\P4_IR_reg[23]/NET0131  & ~n27812 ;
  assign n27814 = ~n15734 & ~n15736 ;
  assign n27815 = ~\P4_IR_reg[23]/NET0131  & ~n27814 ;
  assign n27829 = \P4_IR_reg[2]/NET0131  & \P4_reg2_reg[2]/NET0131  ;
  assign n27830 = ~\P4_IR_reg[2]/NET0131  & ~\P4_reg2_reg[2]/NET0131  ;
  assign n27831 = ~n27829 & ~n27830 ;
  assign n27832 = ~\P4_IR_reg[1]/NET0131  & ~\P4_reg2_reg[1]/NET0131  ;
  assign n27833 = \P4_IR_reg[1]/NET0131  & \P4_reg2_reg[1]/NET0131  ;
  assign n27834 = ~n27799 & ~n27833 ;
  assign n27835 = ~n27832 & ~n27834 ;
  assign n27837 = n27831 & n27835 ;
  assign n27836 = ~n27831 & ~n27835 ;
  assign n27838 = n15733 & ~n27836 ;
  assign n27839 = ~n27837 & n27838 ;
  assign n27817 = \P4_IR_reg[2]/NET0131  & \P4_reg1_reg[2]/NET0131  ;
  assign n27818 = ~\P4_IR_reg[2]/NET0131  & ~\P4_reg1_reg[2]/NET0131  ;
  assign n27819 = ~n27817 & ~n27818 ;
  assign n27820 = ~\P4_IR_reg[1]/NET0131  & ~\P4_reg1_reg[1]/NET0131  ;
  assign n27821 = \P4_IR_reg[1]/NET0131  & \P4_reg1_reg[1]/NET0131  ;
  assign n27822 = ~n27802 & ~n27821 ;
  assign n27823 = ~n27820 & ~n27822 ;
  assign n27825 = n27819 & n27823 ;
  assign n27824 = ~n27819 & ~n27823 ;
  assign n27826 = n27804 & ~n27824 ;
  assign n27827 = ~n27825 & n27826 ;
  assign n27816 = \P4_addr_reg[2]/NET0131  & n15745 ;
  assign n27828 = \P4_IR_reg[2]/NET0131  & n21786 ;
  assign n27840 = ~n27816 & ~n27828 ;
  assign n27841 = ~n27827 & n27840 ;
  assign n27842 = ~n27839 & n27841 ;
  assign n27843 = ~n27815 & ~n27842 ;
  assign n27844 = ~n27813 & ~n27843 ;
  assign n27845 = \P3_rd_reg/NET0131  & ~n27844 ;
  assign n27846 = ~n27796 & ~n27845 ;
  assign n27847 = \P4_addr_reg[4]/NET0131  & ~n15736 ;
  assign n27848 = n15734 & n27847 ;
  assign n27849 = ~n27811 & ~n27848 ;
  assign n27850 = ~\P4_IR_reg[23]/NET0131  & ~n27849 ;
  assign n27851 = n27815 & ~n27847 ;
  assign n27867 = \P4_IR_reg[4]/NET0131  & \P4_reg1_reg[4]/NET0131  ;
  assign n27868 = ~\P4_IR_reg[4]/NET0131  & ~\P4_reg1_reg[4]/NET0131  ;
  assign n27869 = ~n27867 & ~n27868 ;
  assign n27870 = ~\P4_IR_reg[3]/NET0131  & ~\P4_reg1_reg[3]/NET0131  ;
  assign n27871 = \P4_IR_reg[3]/NET0131  & \P4_reg1_reg[3]/NET0131  ;
  assign n27872 = ~n27817 & ~n27823 ;
  assign n27873 = ~n27818 & ~n27872 ;
  assign n27874 = ~n27871 & ~n27873 ;
  assign n27875 = ~n27870 & ~n27874 ;
  assign n27877 = n27869 & n27875 ;
  assign n27876 = ~n27869 & ~n27875 ;
  assign n27878 = n27804 & ~n27876 ;
  assign n27879 = ~n27877 & n27878 ;
  assign n27854 = \P4_IR_reg[4]/NET0131  & \P4_reg2_reg[4]/NET0131  ;
  assign n27855 = ~\P4_IR_reg[4]/NET0131  & ~\P4_reg2_reg[4]/NET0131  ;
  assign n27856 = ~n27854 & ~n27855 ;
  assign n27857 = ~\P4_IR_reg[3]/NET0131  & ~\P4_reg2_reg[3]/NET0131  ;
  assign n27858 = \P4_IR_reg[3]/NET0131  & \P4_reg2_reg[3]/NET0131  ;
  assign n27859 = ~n27829 & ~n27835 ;
  assign n27860 = ~n27830 & ~n27859 ;
  assign n27861 = ~n27858 & ~n27860 ;
  assign n27862 = ~n27857 & ~n27861 ;
  assign n27864 = n27856 & n27862 ;
  assign n27863 = ~n27856 & ~n27862 ;
  assign n27865 = n15733 & ~n27863 ;
  assign n27866 = ~n27864 & n27865 ;
  assign n27852 = \P4_addr_reg[4]/NET0131  & n15745 ;
  assign n27853 = \P4_IR_reg[4]/NET0131  & n21786 ;
  assign n27880 = ~n27852 & ~n27853 ;
  assign n27881 = ~n27866 & n27880 ;
  assign n27882 = ~n27879 & n27881 ;
  assign n27883 = ~n27851 & ~n27882 ;
  assign n27884 = ~n27850 & ~n27883 ;
  assign n27885 = \P3_rd_reg/NET0131  & ~n27884 ;
  assign n27886 = ~n23588 & ~n27885 ;
  assign n27887 = \P2_P1_lWord_reg[9]/NET0131  & ~n25156 ;
  assign n27888 = \P2_P1_EAX_reg[9]/NET0131  & n24899 ;
  assign n27889 = n21062 & n23792 ;
  assign n27890 = ~n27888 & ~n27889 ;
  assign n27891 = n11623 & ~n27890 ;
  assign n27892 = ~n27887 & ~n27891 ;
  assign n27893 = \P1_P1_lWord_reg[9]/NET0131  & ~n25165 ;
  assign n27894 = \P1_P1_EAX_reg[9]/NET0131  & n24503 ;
  assign n27895 = ~n23948 & ~n27894 ;
  assign n27896 = n8355 & ~n27895 ;
  assign n27897 = ~n27893 & ~n27896 ;
  assign n27943 = ~\P1_P2_InstQueueWr_Addr_reg[0]/NET0131  & ~\P1_P2_InstQueueWr_Addr_reg[1]/NET0131  ;
  assign n27944 = ~\P1_P2_InstQueueWr_Addr_reg[2]/NET0131  & n27943 ;
  assign n27945 = \P1_P2_InstQueueWr_Addr_reg[3]/NET0131  & n27944 ;
  assign n27915 = ~\P1_P2_Address_reg[26]/NET0131  & ~\P1_P2_Address_reg[27]/NET0131  ;
  assign n27916 = ~\P1_P2_Address_reg[28]/NET0131  & ~\P1_P2_Address_reg[2]/NET0131  ;
  assign n27922 = n27915 & n27916 ;
  assign n27913 = ~\P1_P2_Address_reg[22]/NET0131  & ~\P1_P2_Address_reg[23]/NET0131  ;
  assign n27914 = ~\P1_P2_Address_reg[24]/NET0131  & ~\P1_P2_Address_reg[25]/NET0131  ;
  assign n27923 = n27913 & n27914 ;
  assign n27929 = n27922 & n27923 ;
  assign n27919 = ~\P1_P2_Address_reg[7]/NET0131  & ~\P1_P2_Address_reg[8]/NET0131  ;
  assign n27920 = ~\P1_P2_Address_reg[9]/NET0131  & n27919 ;
  assign n27917 = ~\P1_P2_Address_reg[3]/NET0131  & ~\P1_P2_Address_reg[4]/NET0131  ;
  assign n27918 = ~\P1_P2_Address_reg[5]/NET0131  & ~\P1_P2_Address_reg[6]/NET0131  ;
  assign n27921 = n27917 & n27918 ;
  assign n27930 = n27920 & n27921 ;
  assign n27931 = n27929 & n27930 ;
  assign n27906 = ~\P1_P2_Address_reg[0]/NET0131  & ~\P1_P2_Address_reg[10]/NET0131  ;
  assign n27907 = ~\P1_P2_Address_reg[11]/NET0131  & ~\P1_P2_Address_reg[12]/NET0131  ;
  assign n27908 = ~\P1_P2_Address_reg[13]/NET0131  & ~\P1_P2_Address_reg[14]/NET0131  ;
  assign n27926 = n27907 & n27908 ;
  assign n27927 = n27906 & n27926 ;
  assign n27911 = ~\P1_P2_Address_reg[19]/NET0131  & ~\P1_P2_Address_reg[1]/NET0131  ;
  assign n27912 = ~\P1_P2_Address_reg[20]/NET0131  & ~\P1_P2_Address_reg[21]/NET0131  ;
  assign n27924 = n27911 & n27912 ;
  assign n27909 = ~\P1_P2_Address_reg[15]/NET0131  & ~\P1_P2_Address_reg[16]/NET0131  ;
  assign n27910 = ~\P1_P2_Address_reg[17]/NET0131  & ~\P1_P2_Address_reg[18]/NET0131  ;
  assign n27925 = n27909 & n27910 ;
  assign n27928 = n27924 & n27925 ;
  assign n27932 = n27927 & n27928 ;
  assign n27933 = n27931 & n27932 ;
  assign n27934 = \P1_P2_Address_reg[29]/NET0131  & ~n27933 ;
  assign n27946 = \P1_buf2_reg[28]/NET0131  & ~n27934 ;
  assign n27947 = \P1_buf1_reg[28]/NET0131  & n27934 ;
  assign n27948 = ~n27946 & ~n27947 ;
  assign n27949 = n27945 & ~n27948 ;
  assign n27950 = \P1_P2_InstQueueWr_Addr_reg[0]/NET0131  & ~\P1_P2_InstQueueWr_Addr_reg[1]/NET0131  ;
  assign n27951 = ~\P1_P2_InstQueueWr_Addr_reg[2]/NET0131  & n27950 ;
  assign n27952 = \P1_P2_InstQueueWr_Addr_reg[3]/NET0131  & n27951 ;
  assign n27953 = \P1_buf2_reg[20]/NET0131  & ~n27934 ;
  assign n27954 = \P1_buf1_reg[20]/NET0131  & n27934 ;
  assign n27955 = ~n27953 & ~n27954 ;
  assign n27956 = n27952 & ~n27955 ;
  assign n27957 = ~n27949 & ~n27956 ;
  assign n27958 = \P1_P2_DataWidth_reg[1]/NET0131  & ~n27957 ;
  assign n27899 = \P1_P2_InstQueueWr_Addr_reg[0]/NET0131  & \P1_P2_InstQueueWr_Addr_reg[1]/NET0131  ;
  assign n27900 = ~\P1_P2_InstQueueWr_Addr_reg[2]/NET0131  & n27899 ;
  assign n27901 = \P1_P2_InstQueueWr_Addr_reg[3]/NET0131  & n27900 ;
  assign n27902 = ~\P1_P2_InstQueueWr_Addr_reg[0]/NET0131  & \P1_P2_InstQueueWr_Addr_reg[1]/NET0131  ;
  assign n27903 = ~\P1_P2_InstQueueWr_Addr_reg[2]/NET0131  & n27902 ;
  assign n27904 = \P1_P2_InstQueueWr_Addr_reg[3]/NET0131  & n27903 ;
  assign n27905 = ~n27901 & ~n27904 ;
  assign n27935 = \P1_buf2_reg[4]/NET0131  & ~n27934 ;
  assign n27936 = \P1_buf1_reg[4]/NET0131  & n27934 ;
  assign n27937 = ~n27935 & ~n27936 ;
  assign n27938 = ~n27905 & ~n27937 ;
  assign n27939 = \P1_P2_InstQueue_reg[11][4]/NET0131  & ~n27901 ;
  assign n27940 = ~n27904 & n27939 ;
  assign n27941 = ~n27938 & ~n27940 ;
  assign n27959 = ~n27945 & ~n27952 ;
  assign n27960 = \P1_P2_DataWidth_reg[1]/NET0131  & ~n27959 ;
  assign n27961 = ~n27941 & ~n27960 ;
  assign n27962 = ~n27958 & ~n27961 ;
  assign n27963 = n25928 & ~n27962 ;
  assign n27964 = ~n25508 & n27901 ;
  assign n27965 = ~n27939 & ~n27964 ;
  assign n27966 = n27608 & ~n27965 ;
  assign n27898 = ~\P1_P2_State2_reg[1]/NET0131  & n25935 ;
  assign n27942 = n27898 & ~n27941 ;
  assign n27967 = n25934 & n27606 ;
  assign n27968 = ~n25418 & ~n27967 ;
  assign n27969 = ~n27675 & n27968 ;
  assign n27970 = ~n25921 & ~n25925 ;
  assign n27971 = ~n25918 & n27970 ;
  assign n27972 = n27969 & n27971 ;
  assign n27973 = \P1_P2_InstQueue_reg[11][4]/NET0131  & ~n27972 ;
  assign n27974 = ~n27942 & ~n27973 ;
  assign n27975 = ~n27966 & n27974 ;
  assign n27976 = ~n27963 & n27975 ;
  assign n28025 = ~\P2_P2_InstQueueWr_Addr_reg[0]/NET0131  & ~\P2_P2_InstQueueWr_Addr_reg[1]/NET0131  ;
  assign n28026 = ~\P2_P2_InstQueueWr_Addr_reg[2]/NET0131  & n28025 ;
  assign n28027 = \P2_P2_InstQueueWr_Addr_reg[3]/NET0131  & n28026 ;
  assign n27994 = ~\P2_P2_Address_reg[26]/NET0131  & ~\P2_P2_Address_reg[27]/NET0131  ;
  assign n27995 = ~\P2_P2_Address_reg[28]/NET0131  & ~\P2_P2_Address_reg[2]/NET0131  ;
  assign n28001 = n27994 & n27995 ;
  assign n27992 = ~\P2_P2_Address_reg[22]/NET0131  & ~\P2_P2_Address_reg[23]/NET0131  ;
  assign n27993 = ~\P2_P2_Address_reg[24]/NET0131  & ~\P2_P2_Address_reg[25]/NET0131  ;
  assign n28002 = n27992 & n27993 ;
  assign n28008 = n28001 & n28002 ;
  assign n27998 = ~\P2_P2_Address_reg[7]/NET0131  & ~\P2_P2_Address_reg[8]/NET0131  ;
  assign n27999 = ~\P2_P2_Address_reg[9]/NET0131  & n27998 ;
  assign n27996 = ~\P2_P2_Address_reg[3]/NET0131  & ~\P2_P2_Address_reg[4]/NET0131  ;
  assign n27997 = ~\P2_P2_Address_reg[5]/NET0131  & ~\P2_P2_Address_reg[6]/NET0131  ;
  assign n28000 = n27996 & n27997 ;
  assign n28009 = n27999 & n28000 ;
  assign n28010 = n28008 & n28009 ;
  assign n27985 = ~\P2_P2_Address_reg[0]/NET0131  & ~\P2_P2_Address_reg[10]/NET0131  ;
  assign n27986 = ~\P2_P2_Address_reg[11]/NET0131  & ~\P2_P2_Address_reg[12]/NET0131  ;
  assign n27987 = ~\P2_P2_Address_reg[13]/NET0131  & ~\P2_P2_Address_reg[14]/NET0131  ;
  assign n28005 = n27986 & n27987 ;
  assign n28006 = n27985 & n28005 ;
  assign n27990 = ~\P2_P2_Address_reg[19]/NET0131  & ~\P2_P2_Address_reg[1]/NET0131  ;
  assign n27991 = ~\P2_P2_Address_reg[20]/NET0131  & ~\P2_P2_Address_reg[21]/NET0131  ;
  assign n28003 = n27990 & n27991 ;
  assign n27988 = ~\P2_P2_Address_reg[15]/NET0131  & ~\P2_P2_Address_reg[16]/NET0131  ;
  assign n27989 = ~\P2_P2_Address_reg[17]/NET0131  & ~\P2_P2_Address_reg[18]/NET0131  ;
  assign n28004 = n27988 & n27989 ;
  assign n28007 = n28003 & n28004 ;
  assign n28011 = n28006 & n28007 ;
  assign n28012 = n28010 & n28011 ;
  assign n28013 = \P2_P2_Address_reg[29]/NET0131  & ~n28012 ;
  assign n28028 = \P2_buf2_reg[28]/NET0131  & ~n28013 ;
  assign n28029 = \P2_buf1_reg[28]/NET0131  & n28013 ;
  assign n28030 = ~n28028 & ~n28029 ;
  assign n28031 = n28027 & ~n28030 ;
  assign n28032 = \P2_P2_InstQueueWr_Addr_reg[0]/NET0131  & ~\P2_P2_InstQueueWr_Addr_reg[1]/NET0131  ;
  assign n28033 = ~\P2_P2_InstQueueWr_Addr_reg[2]/NET0131  & n28032 ;
  assign n28034 = \P2_P2_InstQueueWr_Addr_reg[3]/NET0131  & n28033 ;
  assign n28035 = \P2_buf2_reg[20]/NET0131  & ~n28013 ;
  assign n28036 = \P2_buf1_reg[20]/NET0131  & n28013 ;
  assign n28037 = ~n28035 & ~n28036 ;
  assign n28038 = n28034 & ~n28037 ;
  assign n28039 = ~n28031 & ~n28038 ;
  assign n28040 = \P2_P2_DataWidth_reg[1]/NET0131  & ~n28039 ;
  assign n27978 = \P2_P2_InstQueueWr_Addr_reg[0]/NET0131  & \P2_P2_InstQueueWr_Addr_reg[1]/NET0131  ;
  assign n27979 = ~\P2_P2_InstQueueWr_Addr_reg[2]/NET0131  & n27978 ;
  assign n27980 = \P2_P2_InstQueueWr_Addr_reg[3]/NET0131  & n27979 ;
  assign n27981 = ~\P2_P2_InstQueueWr_Addr_reg[0]/NET0131  & \P2_P2_InstQueueWr_Addr_reg[1]/NET0131  ;
  assign n27982 = ~\P2_P2_InstQueueWr_Addr_reg[2]/NET0131  & n27981 ;
  assign n27983 = \P2_P2_InstQueueWr_Addr_reg[3]/NET0131  & n27982 ;
  assign n27984 = ~n27980 & ~n27983 ;
  assign n28014 = \P2_buf2_reg[4]/NET0131  & ~n28013 ;
  assign n28015 = \P2_buf1_reg[4]/NET0131  & n28013 ;
  assign n28016 = ~n28014 & ~n28015 ;
  assign n28017 = ~n27984 & ~n28016 ;
  assign n28018 = \P2_P2_InstQueue_reg[11][4]/NET0131  & ~n27980 ;
  assign n28019 = ~n27983 & n28018 ;
  assign n28020 = ~n28017 & ~n28019 ;
  assign n28041 = ~n28027 & ~n28034 ;
  assign n28042 = \P2_P2_DataWidth_reg[1]/NET0131  & ~n28041 ;
  assign n28043 = ~n28020 & ~n28042 ;
  assign n28044 = ~n28040 & ~n28043 ;
  assign n28045 = n26794 & ~n28044 ;
  assign n28022 = ~n26417 & n27980 ;
  assign n28023 = ~n28018 & ~n28022 ;
  assign n28024 = n27613 & ~n28023 ;
  assign n27977 = ~\P2_P2_State2_reg[1]/NET0131  & n26802 ;
  assign n28021 = n27977 & ~n28020 ;
  assign n28046 = n26285 & n26290 ;
  assign n28047 = ~n26291 & ~n28046 ;
  assign n28048 = ~n26792 & ~n27614 ;
  assign n28049 = ~n26296 & n28048 ;
  assign n28050 = n28047 & n28049 ;
  assign n28051 = \P2_P2_InstQueue_reg[11][4]/NET0131  & ~n28050 ;
  assign n28052 = ~n28021 & ~n28051 ;
  assign n28053 = ~n28024 & n28052 ;
  assign n28054 = ~n28045 & n28053 ;
  assign n28064 = \P1_P2_InstQueueWr_Addr_reg[2]/NET0131  & n27950 ;
  assign n28065 = \P1_P2_InstQueueWr_Addr_reg[3]/NET0131  & n28064 ;
  assign n28066 = ~n27948 & n28065 ;
  assign n28067 = \P1_P2_InstQueueWr_Addr_reg[2]/NET0131  & n27902 ;
  assign n28068 = \P1_P2_InstQueueWr_Addr_reg[3]/NET0131  & n28067 ;
  assign n28069 = ~n27955 & n28068 ;
  assign n28070 = ~n28066 & ~n28069 ;
  assign n28071 = \P1_P2_DataWidth_reg[1]/NET0131  & ~n28070 ;
  assign n28055 = ~\P1_P2_InstQueueWr_Addr_reg[3]/NET0131  & n27944 ;
  assign n28056 = \P1_P2_InstQueueWr_Addr_reg[2]/NET0131  & n27899 ;
  assign n28057 = \P1_P2_InstQueueWr_Addr_reg[3]/NET0131  & n28056 ;
  assign n28058 = ~n28055 & ~n28057 ;
  assign n28059 = ~n27937 & ~n28058 ;
  assign n28060 = \P1_P2_InstQueue_reg[0][4]/NET0131  & ~n28055 ;
  assign n28061 = ~n28057 & n28060 ;
  assign n28062 = ~n28059 & ~n28061 ;
  assign n28072 = ~n28065 & ~n28068 ;
  assign n28073 = \P1_P2_DataWidth_reg[1]/NET0131  & ~n28072 ;
  assign n28074 = ~n28062 & ~n28073 ;
  assign n28075 = ~n28071 & ~n28074 ;
  assign n28076 = n25928 & ~n28075 ;
  assign n28077 = ~n25508 & n28055 ;
  assign n28078 = ~n28060 & ~n28077 ;
  assign n28079 = n27608 & ~n28078 ;
  assign n28063 = n27898 & ~n28062 ;
  assign n28080 = \P1_P2_InstQueue_reg[0][4]/NET0131  & ~n27972 ;
  assign n28081 = ~n28063 & ~n28080 ;
  assign n28082 = ~n28079 & n28081 ;
  assign n28083 = ~n28076 & n28082 ;
  assign n28090 = ~\P1_P2_InstQueueWr_Addr_reg[3]/NET0131  & n28056 ;
  assign n28091 = ~n27948 & n28090 ;
  assign n28092 = n27945 & ~n27955 ;
  assign n28093 = ~n28091 & ~n28092 ;
  assign n28094 = \P1_P2_DataWidth_reg[1]/NET0131  & ~n28093 ;
  assign n28084 = ~n27904 & ~n27952 ;
  assign n28085 = ~n27937 & ~n28084 ;
  assign n28086 = \P1_P2_InstQueue_reg[10][4]/NET0131  & ~n27904 ;
  assign n28087 = ~n27952 & n28086 ;
  assign n28088 = ~n28085 & ~n28087 ;
  assign n28095 = ~n27945 & ~n28090 ;
  assign n28096 = \P1_P2_DataWidth_reg[1]/NET0131  & ~n28095 ;
  assign n28097 = ~n28088 & ~n28096 ;
  assign n28098 = ~n28094 & ~n28097 ;
  assign n28099 = n25928 & ~n28098 ;
  assign n28100 = ~n25508 & n27904 ;
  assign n28101 = ~n28086 & ~n28100 ;
  assign n28102 = n27608 & ~n28101 ;
  assign n28089 = n27898 & ~n28088 ;
  assign n28103 = \P1_P2_InstQueue_reg[10][4]/NET0131  & ~n27972 ;
  assign n28104 = ~n28089 & ~n28103 ;
  assign n28105 = ~n28102 & n28104 ;
  assign n28106 = ~n28099 & n28105 ;
  assign n28115 = ~n27948 & n27952 ;
  assign n28116 = n27904 & ~n27955 ;
  assign n28117 = ~n28115 & ~n28116 ;
  assign n28118 = \P1_P2_DataWidth_reg[1]/NET0131  & ~n28117 ;
  assign n28107 = \P1_P2_InstQueueWr_Addr_reg[2]/NET0131  & n27943 ;
  assign n28108 = \P1_P2_InstQueueWr_Addr_reg[3]/NET0131  & n28107 ;
  assign n28109 = ~n27901 & ~n28108 ;
  assign n28110 = ~n27937 & ~n28109 ;
  assign n28111 = \P1_P2_InstQueue_reg[12][4]/NET0131  & ~n28108 ;
  assign n28112 = ~n27901 & n28111 ;
  assign n28113 = ~n28110 & ~n28112 ;
  assign n28119 = \P1_P2_DataWidth_reg[1]/NET0131  & ~n28084 ;
  assign n28120 = ~n28113 & ~n28119 ;
  assign n28121 = ~n28118 & ~n28120 ;
  assign n28122 = n25928 & ~n28121 ;
  assign n28123 = ~n25508 & n28108 ;
  assign n28124 = ~n28111 & ~n28123 ;
  assign n28125 = n27608 & ~n28124 ;
  assign n28114 = n27898 & ~n28113 ;
  assign n28126 = \P1_P2_InstQueue_reg[12][4]/NET0131  & ~n27972 ;
  assign n28127 = ~n28114 & ~n28126 ;
  assign n28128 = ~n28125 & n28127 ;
  assign n28129 = ~n28122 & n28128 ;
  assign n28136 = n27904 & ~n27948 ;
  assign n28137 = n27901 & ~n27955 ;
  assign n28138 = ~n28136 & ~n28137 ;
  assign n28139 = \P1_P2_DataWidth_reg[1]/NET0131  & ~n28138 ;
  assign n28130 = ~n28065 & ~n28108 ;
  assign n28131 = ~n27937 & ~n28130 ;
  assign n28132 = \P1_P2_InstQueue_reg[13][4]/NET0131  & ~n28065 ;
  assign n28133 = ~n28108 & n28132 ;
  assign n28134 = ~n28131 & ~n28133 ;
  assign n28140 = \P1_P2_DataWidth_reg[1]/NET0131  & ~n27905 ;
  assign n28141 = ~n28134 & ~n28140 ;
  assign n28142 = ~n28139 & ~n28141 ;
  assign n28143 = n25928 & ~n28142 ;
  assign n28144 = ~n25508 & n28065 ;
  assign n28145 = ~n28132 & ~n28144 ;
  assign n28146 = n27608 & ~n28145 ;
  assign n28135 = n27898 & ~n28134 ;
  assign n28147 = \P1_P2_InstQueue_reg[13][4]/NET0131  & ~n27972 ;
  assign n28148 = ~n28135 & ~n28147 ;
  assign n28149 = ~n28146 & n28148 ;
  assign n28150 = ~n28143 & n28149 ;
  assign n28156 = n27901 & ~n27948 ;
  assign n28157 = ~n27955 & n28108 ;
  assign n28158 = ~n28156 & ~n28157 ;
  assign n28159 = \P1_P2_DataWidth_reg[1]/NET0131  & ~n28158 ;
  assign n28151 = ~n27937 & ~n28072 ;
  assign n28152 = \P1_P2_InstQueue_reg[14][4]/NET0131  & ~n28068 ;
  assign n28153 = ~n28065 & n28152 ;
  assign n28154 = ~n28151 & ~n28153 ;
  assign n28160 = \P1_P2_DataWidth_reg[1]/NET0131  & ~n28109 ;
  assign n28161 = ~n28154 & ~n28160 ;
  assign n28162 = ~n28159 & ~n28161 ;
  assign n28163 = n25928 & ~n28162 ;
  assign n28164 = ~n25508 & n28068 ;
  assign n28165 = ~n28152 & ~n28164 ;
  assign n28166 = n27608 & ~n28165 ;
  assign n28155 = n27898 & ~n28154 ;
  assign n28167 = \P1_P2_InstQueue_reg[14][4]/NET0131  & ~n27972 ;
  assign n28168 = ~n28155 & ~n28167 ;
  assign n28169 = ~n28166 & n28168 ;
  assign n28170 = ~n28163 & n28169 ;
  assign n28177 = ~n27948 & n28108 ;
  assign n28178 = ~n27955 & n28065 ;
  assign n28179 = ~n28177 & ~n28178 ;
  assign n28180 = \P1_P2_DataWidth_reg[1]/NET0131  & ~n28179 ;
  assign n28171 = ~n28057 & ~n28068 ;
  assign n28172 = ~n27937 & ~n28171 ;
  assign n28173 = \P1_P2_InstQueue_reg[15][4]/NET0131  & ~n28057 ;
  assign n28174 = ~n28068 & n28173 ;
  assign n28175 = ~n28172 & ~n28174 ;
  assign n28181 = \P1_P2_DataWidth_reg[1]/NET0131  & ~n28130 ;
  assign n28182 = ~n28175 & ~n28181 ;
  assign n28183 = ~n28180 & ~n28182 ;
  assign n28184 = n25928 & ~n28183 ;
  assign n28185 = ~n25508 & n28057 ;
  assign n28186 = ~n28173 & ~n28185 ;
  assign n28187 = n27608 & ~n28186 ;
  assign n28176 = n27898 & ~n28175 ;
  assign n28188 = \P1_P2_InstQueue_reg[15][4]/NET0131  & ~n27972 ;
  assign n28189 = ~n28176 & ~n28188 ;
  assign n28190 = ~n28187 & n28189 ;
  assign n28191 = ~n28184 & n28190 ;
  assign n28199 = ~n27948 & n28068 ;
  assign n28200 = ~n27955 & n28057 ;
  assign n28201 = ~n28199 & ~n28200 ;
  assign n28202 = \P1_P2_DataWidth_reg[1]/NET0131  & ~n28201 ;
  assign n28192 = ~\P1_P2_InstQueueWr_Addr_reg[3]/NET0131  & n27951 ;
  assign n28193 = ~n28055 & ~n28192 ;
  assign n28194 = ~n27937 & ~n28193 ;
  assign n28195 = \P1_P2_InstQueue_reg[1][4]/NET0131  & ~n28192 ;
  assign n28196 = ~n28055 & n28195 ;
  assign n28197 = ~n28194 & ~n28196 ;
  assign n28203 = \P1_P2_DataWidth_reg[1]/NET0131  & ~n28171 ;
  assign n28204 = ~n28197 & ~n28203 ;
  assign n28205 = ~n28202 & ~n28204 ;
  assign n28206 = n25928 & ~n28205 ;
  assign n28207 = ~n25508 & n28192 ;
  assign n28208 = ~n28195 & ~n28207 ;
  assign n28209 = n27608 & ~n28208 ;
  assign n28198 = n27898 & ~n28197 ;
  assign n28210 = \P1_P2_InstQueue_reg[1][4]/NET0131  & ~n27972 ;
  assign n28211 = ~n28198 & ~n28210 ;
  assign n28212 = ~n28209 & n28211 ;
  assign n28213 = ~n28206 & n28212 ;
  assign n28221 = ~n27948 & n28057 ;
  assign n28222 = ~n27955 & n28055 ;
  assign n28223 = ~n28221 & ~n28222 ;
  assign n28224 = \P1_P2_DataWidth_reg[1]/NET0131  & ~n28223 ;
  assign n28214 = ~\P1_P2_InstQueueWr_Addr_reg[3]/NET0131  & n27903 ;
  assign n28215 = ~n28192 & ~n28214 ;
  assign n28216 = ~n27937 & ~n28215 ;
  assign n28217 = \P1_P2_InstQueue_reg[2][4]/NET0131  & ~n28214 ;
  assign n28218 = ~n28192 & n28217 ;
  assign n28219 = ~n28216 & ~n28218 ;
  assign n28225 = \P1_P2_DataWidth_reg[1]/NET0131  & ~n28058 ;
  assign n28226 = ~n28219 & ~n28225 ;
  assign n28227 = ~n28224 & ~n28226 ;
  assign n28228 = n25928 & ~n28227 ;
  assign n28229 = ~n25508 & n28214 ;
  assign n28230 = ~n28217 & ~n28229 ;
  assign n28231 = n27608 & ~n28230 ;
  assign n28220 = n27898 & ~n28219 ;
  assign n28232 = \P1_P2_InstQueue_reg[2][4]/NET0131  & ~n27972 ;
  assign n28233 = ~n28220 & ~n28232 ;
  assign n28234 = ~n28231 & n28233 ;
  assign n28235 = ~n28228 & n28234 ;
  assign n28243 = ~n27948 & n28055 ;
  assign n28244 = ~n27955 & n28192 ;
  assign n28245 = ~n28243 & ~n28244 ;
  assign n28246 = \P1_P2_DataWidth_reg[1]/NET0131  & ~n28245 ;
  assign n28236 = ~\P1_P2_InstQueueWr_Addr_reg[3]/NET0131  & n27900 ;
  assign n28237 = ~n28214 & ~n28236 ;
  assign n28238 = ~n27937 & ~n28237 ;
  assign n28239 = \P1_P2_InstQueue_reg[3][4]/NET0131  & ~n28236 ;
  assign n28240 = ~n28214 & n28239 ;
  assign n28241 = ~n28238 & ~n28240 ;
  assign n28247 = \P1_P2_DataWidth_reg[1]/NET0131  & ~n28193 ;
  assign n28248 = ~n28241 & ~n28247 ;
  assign n28249 = ~n28246 & ~n28248 ;
  assign n28250 = n25928 & ~n28249 ;
  assign n28251 = ~n25508 & n28236 ;
  assign n28252 = ~n28239 & ~n28251 ;
  assign n28253 = n27608 & ~n28252 ;
  assign n28242 = n27898 & ~n28241 ;
  assign n28254 = \P1_P2_InstQueue_reg[3][4]/NET0131  & ~n27972 ;
  assign n28255 = ~n28242 & ~n28254 ;
  assign n28256 = ~n28253 & n28255 ;
  assign n28257 = ~n28250 & n28256 ;
  assign n28265 = ~n27948 & n28192 ;
  assign n28266 = ~n27955 & n28214 ;
  assign n28267 = ~n28265 & ~n28266 ;
  assign n28268 = \P1_P2_DataWidth_reg[1]/NET0131  & ~n28267 ;
  assign n28258 = ~\P1_P2_InstQueueWr_Addr_reg[3]/NET0131  & n28107 ;
  assign n28259 = ~n28236 & ~n28258 ;
  assign n28260 = ~n27937 & ~n28259 ;
  assign n28261 = \P1_P2_InstQueue_reg[4][4]/NET0131  & ~n28258 ;
  assign n28262 = ~n28236 & n28261 ;
  assign n28263 = ~n28260 & ~n28262 ;
  assign n28269 = \P1_P2_DataWidth_reg[1]/NET0131  & ~n28215 ;
  assign n28270 = ~n28263 & ~n28269 ;
  assign n28271 = ~n28268 & ~n28270 ;
  assign n28272 = n25928 & ~n28271 ;
  assign n28273 = ~n25508 & n28258 ;
  assign n28274 = ~n28261 & ~n28273 ;
  assign n28275 = n27608 & ~n28274 ;
  assign n28264 = n27898 & ~n28263 ;
  assign n28276 = \P1_P2_InstQueue_reg[4][4]/NET0131  & ~n27972 ;
  assign n28277 = ~n28264 & ~n28276 ;
  assign n28278 = ~n28275 & n28277 ;
  assign n28279 = ~n28272 & n28278 ;
  assign n28287 = ~n27948 & n28214 ;
  assign n28288 = ~n27955 & n28236 ;
  assign n28289 = ~n28287 & ~n28288 ;
  assign n28290 = \P1_P2_DataWidth_reg[1]/NET0131  & ~n28289 ;
  assign n28280 = ~\P1_P2_InstQueueWr_Addr_reg[3]/NET0131  & n28064 ;
  assign n28281 = ~n28258 & ~n28280 ;
  assign n28282 = ~n27937 & ~n28281 ;
  assign n28283 = \P1_P2_InstQueue_reg[5][4]/NET0131  & ~n28280 ;
  assign n28284 = ~n28258 & n28283 ;
  assign n28285 = ~n28282 & ~n28284 ;
  assign n28291 = \P1_P2_DataWidth_reg[1]/NET0131  & ~n28237 ;
  assign n28292 = ~n28285 & ~n28291 ;
  assign n28293 = ~n28290 & ~n28292 ;
  assign n28294 = n25928 & ~n28293 ;
  assign n28295 = ~n25508 & n28280 ;
  assign n28296 = ~n28283 & ~n28295 ;
  assign n28297 = n27608 & ~n28296 ;
  assign n28286 = n27898 & ~n28285 ;
  assign n28298 = \P1_P2_InstQueue_reg[5][4]/NET0131  & ~n27972 ;
  assign n28299 = ~n28286 & ~n28298 ;
  assign n28300 = ~n28297 & n28299 ;
  assign n28301 = ~n28294 & n28300 ;
  assign n28309 = ~n27948 & n28236 ;
  assign n28310 = ~n27955 & n28258 ;
  assign n28311 = ~n28309 & ~n28310 ;
  assign n28312 = \P1_P2_DataWidth_reg[1]/NET0131  & ~n28311 ;
  assign n28302 = ~\P1_P2_InstQueueWr_Addr_reg[3]/NET0131  & n28067 ;
  assign n28303 = ~n28280 & ~n28302 ;
  assign n28304 = ~n27937 & ~n28303 ;
  assign n28305 = \P1_P2_InstQueue_reg[6][4]/NET0131  & ~n28302 ;
  assign n28306 = ~n28280 & n28305 ;
  assign n28307 = ~n28304 & ~n28306 ;
  assign n28313 = \P1_P2_DataWidth_reg[1]/NET0131  & ~n28259 ;
  assign n28314 = ~n28307 & ~n28313 ;
  assign n28315 = ~n28312 & ~n28314 ;
  assign n28316 = n25928 & ~n28315 ;
  assign n28317 = ~n25508 & n28302 ;
  assign n28318 = ~n28305 & ~n28317 ;
  assign n28319 = n27608 & ~n28318 ;
  assign n28308 = n27898 & ~n28307 ;
  assign n28320 = \P1_P2_InstQueue_reg[6][4]/NET0131  & ~n27972 ;
  assign n28321 = ~n28308 & ~n28320 ;
  assign n28322 = ~n28319 & n28321 ;
  assign n28323 = ~n28316 & n28322 ;
  assign n28330 = ~n27948 & n28258 ;
  assign n28331 = ~n27955 & n28280 ;
  assign n28332 = ~n28330 & ~n28331 ;
  assign n28333 = \P1_P2_DataWidth_reg[1]/NET0131  & ~n28332 ;
  assign n28324 = ~n28090 & ~n28302 ;
  assign n28325 = ~n27937 & ~n28324 ;
  assign n28326 = \P1_P2_InstQueue_reg[7][4]/NET0131  & ~n28090 ;
  assign n28327 = ~n28302 & n28326 ;
  assign n28328 = ~n28325 & ~n28327 ;
  assign n28334 = \P1_P2_DataWidth_reg[1]/NET0131  & ~n28281 ;
  assign n28335 = ~n28328 & ~n28334 ;
  assign n28336 = ~n28333 & ~n28335 ;
  assign n28337 = n25928 & ~n28336 ;
  assign n28338 = ~n25508 & n28090 ;
  assign n28339 = ~n28326 & ~n28338 ;
  assign n28340 = n27608 & ~n28339 ;
  assign n28329 = n27898 & ~n28328 ;
  assign n28341 = \P1_P2_InstQueue_reg[7][4]/NET0131  & ~n27972 ;
  assign n28342 = ~n28329 & ~n28341 ;
  assign n28343 = ~n28340 & n28342 ;
  assign n28344 = ~n28337 & n28343 ;
  assign n28350 = ~n27948 & n28280 ;
  assign n28351 = ~n27955 & n28302 ;
  assign n28352 = ~n28350 & ~n28351 ;
  assign n28353 = \P1_P2_DataWidth_reg[1]/NET0131  & ~n28352 ;
  assign n28345 = ~n27937 & ~n28095 ;
  assign n28346 = \P1_P2_InstQueue_reg[8][4]/NET0131  & ~n27945 ;
  assign n28347 = ~n28090 & n28346 ;
  assign n28348 = ~n28345 & ~n28347 ;
  assign n28354 = \P1_P2_DataWidth_reg[1]/NET0131  & ~n28303 ;
  assign n28355 = ~n28348 & ~n28354 ;
  assign n28356 = ~n28353 & ~n28355 ;
  assign n28357 = n25928 & ~n28356 ;
  assign n28358 = ~n25508 & n27945 ;
  assign n28359 = ~n28346 & ~n28358 ;
  assign n28360 = n27608 & ~n28359 ;
  assign n28349 = n27898 & ~n28348 ;
  assign n28361 = \P1_P2_InstQueue_reg[8][4]/NET0131  & ~n27972 ;
  assign n28362 = ~n28349 & ~n28361 ;
  assign n28363 = ~n28360 & n28362 ;
  assign n28364 = ~n28357 & n28363 ;
  assign n28370 = ~n27948 & n28302 ;
  assign n28371 = ~n27955 & n28090 ;
  assign n28372 = ~n28370 & ~n28371 ;
  assign n28373 = \P1_P2_DataWidth_reg[1]/NET0131  & ~n28372 ;
  assign n28365 = ~n27937 & ~n27959 ;
  assign n28366 = \P1_P2_InstQueue_reg[9][4]/NET0131  & ~n27952 ;
  assign n28367 = ~n27945 & n28366 ;
  assign n28368 = ~n28365 & ~n28367 ;
  assign n28374 = \P1_P2_DataWidth_reg[1]/NET0131  & ~n28324 ;
  assign n28375 = ~n28368 & ~n28374 ;
  assign n28376 = ~n28373 & ~n28375 ;
  assign n28377 = n25928 & ~n28376 ;
  assign n28378 = ~n25508 & n27952 ;
  assign n28379 = ~n28366 & ~n28378 ;
  assign n28380 = n27608 & ~n28379 ;
  assign n28369 = n27898 & ~n28368 ;
  assign n28381 = \P1_P2_InstQueue_reg[9][4]/NET0131  & ~n27972 ;
  assign n28382 = ~n28369 & ~n28381 ;
  assign n28383 = ~n28380 & n28382 ;
  assign n28384 = ~n28377 & n28383 ;
  assign n28397 = \P2_P2_InstQueueWr_Addr_reg[2]/NET0131  & n28032 ;
  assign n28398 = \P2_P2_InstQueueWr_Addr_reg[3]/NET0131  & n28397 ;
  assign n28399 = ~n28030 & n28398 ;
  assign n28400 = \P2_P2_InstQueueWr_Addr_reg[2]/NET0131  & n27981 ;
  assign n28401 = \P2_P2_InstQueueWr_Addr_reg[3]/NET0131  & n28400 ;
  assign n28402 = ~n28037 & n28401 ;
  assign n28403 = ~n28399 & ~n28402 ;
  assign n28404 = \P2_P2_DataWidth_reg[1]/NET0131  & ~n28403 ;
  assign n28385 = ~\P2_P2_InstQueueWr_Addr_reg[3]/NET0131  & n28026 ;
  assign n28386 = \P2_P2_InstQueueWr_Addr_reg[2]/NET0131  & n27978 ;
  assign n28387 = \P2_P2_InstQueueWr_Addr_reg[3]/NET0131  & n28386 ;
  assign n28388 = ~n28385 & ~n28387 ;
  assign n28389 = ~n28016 & ~n28388 ;
  assign n28390 = \P2_P2_InstQueue_reg[0][4]/NET0131  & ~n28385 ;
  assign n28391 = ~n28387 & n28390 ;
  assign n28392 = ~n28389 & ~n28391 ;
  assign n28405 = ~n28398 & ~n28401 ;
  assign n28406 = \P2_P2_DataWidth_reg[1]/NET0131  & ~n28405 ;
  assign n28407 = ~n28392 & ~n28406 ;
  assign n28408 = ~n28404 & ~n28407 ;
  assign n28409 = n26794 & ~n28408 ;
  assign n28394 = ~n26417 & n28385 ;
  assign n28395 = ~n28390 & ~n28394 ;
  assign n28396 = n27613 & ~n28395 ;
  assign n28393 = n27977 & ~n28392 ;
  assign n28410 = \P2_P2_InstQueue_reg[0][4]/NET0131  & ~n28050 ;
  assign n28411 = ~n28393 & ~n28410 ;
  assign n28412 = ~n28396 & n28411 ;
  assign n28413 = ~n28409 & n28412 ;
  assign n28423 = ~\P2_P2_InstQueueWr_Addr_reg[3]/NET0131  & n28386 ;
  assign n28424 = ~n28030 & n28423 ;
  assign n28425 = n28027 & ~n28037 ;
  assign n28426 = ~n28424 & ~n28425 ;
  assign n28427 = \P2_P2_DataWidth_reg[1]/NET0131  & ~n28426 ;
  assign n28414 = ~n27983 & ~n28034 ;
  assign n28415 = ~n28016 & ~n28414 ;
  assign n28416 = \P2_P2_InstQueue_reg[10][4]/NET0131  & ~n27983 ;
  assign n28417 = ~n28034 & n28416 ;
  assign n28418 = ~n28415 & ~n28417 ;
  assign n28428 = ~n28027 & ~n28423 ;
  assign n28429 = \P2_P2_DataWidth_reg[1]/NET0131  & ~n28428 ;
  assign n28430 = ~n28418 & ~n28429 ;
  assign n28431 = ~n28427 & ~n28430 ;
  assign n28432 = n26794 & ~n28431 ;
  assign n28420 = ~n26417 & n27983 ;
  assign n28421 = ~n28416 & ~n28420 ;
  assign n28422 = n27613 & ~n28421 ;
  assign n28419 = n27977 & ~n28418 ;
  assign n28433 = \P2_P2_InstQueue_reg[10][4]/NET0131  & ~n28050 ;
  assign n28434 = ~n28419 & ~n28433 ;
  assign n28435 = ~n28422 & n28434 ;
  assign n28436 = ~n28432 & n28435 ;
  assign n28448 = ~n28030 & n28034 ;
  assign n28449 = n27983 & ~n28037 ;
  assign n28450 = ~n28448 & ~n28449 ;
  assign n28451 = \P2_P2_DataWidth_reg[1]/NET0131  & ~n28450 ;
  assign n28437 = \P2_P2_InstQueueWr_Addr_reg[2]/NET0131  & n28025 ;
  assign n28438 = \P2_P2_InstQueueWr_Addr_reg[3]/NET0131  & n28437 ;
  assign n28439 = ~n27980 & ~n28438 ;
  assign n28440 = ~n28016 & ~n28439 ;
  assign n28441 = \P2_P2_InstQueue_reg[12][4]/NET0131  & ~n28438 ;
  assign n28442 = ~n27980 & n28441 ;
  assign n28443 = ~n28440 & ~n28442 ;
  assign n28452 = \P2_P2_DataWidth_reg[1]/NET0131  & ~n28414 ;
  assign n28453 = ~n28443 & ~n28452 ;
  assign n28454 = ~n28451 & ~n28453 ;
  assign n28455 = n26794 & ~n28454 ;
  assign n28445 = ~n26417 & n28438 ;
  assign n28446 = ~n28441 & ~n28445 ;
  assign n28447 = n27613 & ~n28446 ;
  assign n28444 = n27977 & ~n28443 ;
  assign n28456 = \P2_P2_InstQueue_reg[12][4]/NET0131  & ~n28050 ;
  assign n28457 = ~n28444 & ~n28456 ;
  assign n28458 = ~n28447 & n28457 ;
  assign n28459 = ~n28455 & n28458 ;
  assign n28469 = n27983 & ~n28030 ;
  assign n28470 = n27980 & ~n28037 ;
  assign n28471 = ~n28469 & ~n28470 ;
  assign n28472 = \P2_P2_DataWidth_reg[1]/NET0131  & ~n28471 ;
  assign n28460 = ~n28398 & ~n28438 ;
  assign n28461 = ~n28016 & ~n28460 ;
  assign n28462 = \P2_P2_InstQueue_reg[13][4]/NET0131  & ~n28398 ;
  assign n28463 = ~n28438 & n28462 ;
  assign n28464 = ~n28461 & ~n28463 ;
  assign n28473 = \P2_P2_DataWidth_reg[1]/NET0131  & ~n27984 ;
  assign n28474 = ~n28464 & ~n28473 ;
  assign n28475 = ~n28472 & ~n28474 ;
  assign n28476 = n26794 & ~n28475 ;
  assign n28466 = ~n26417 & n28398 ;
  assign n28467 = ~n28462 & ~n28466 ;
  assign n28468 = n27613 & ~n28467 ;
  assign n28465 = n27977 & ~n28464 ;
  assign n28477 = \P2_P2_InstQueue_reg[13][4]/NET0131  & ~n28050 ;
  assign n28478 = ~n28465 & ~n28477 ;
  assign n28479 = ~n28468 & n28478 ;
  assign n28480 = ~n28476 & n28479 ;
  assign n28489 = n27980 & ~n28030 ;
  assign n28490 = ~n28037 & n28438 ;
  assign n28491 = ~n28489 & ~n28490 ;
  assign n28492 = \P2_P2_DataWidth_reg[1]/NET0131  & ~n28491 ;
  assign n28481 = ~n28016 & ~n28405 ;
  assign n28482 = \P2_P2_InstQueue_reg[14][4]/NET0131  & ~n28401 ;
  assign n28483 = ~n28398 & n28482 ;
  assign n28484 = ~n28481 & ~n28483 ;
  assign n28493 = \P2_P2_DataWidth_reg[1]/NET0131  & ~n28439 ;
  assign n28494 = ~n28484 & ~n28493 ;
  assign n28495 = ~n28492 & ~n28494 ;
  assign n28496 = n26794 & ~n28495 ;
  assign n28486 = ~n26417 & n28401 ;
  assign n28487 = ~n28482 & ~n28486 ;
  assign n28488 = n27613 & ~n28487 ;
  assign n28485 = n27977 & ~n28484 ;
  assign n28497 = \P2_P2_InstQueue_reg[14][4]/NET0131  & ~n28050 ;
  assign n28498 = ~n28485 & ~n28497 ;
  assign n28499 = ~n28488 & n28498 ;
  assign n28500 = ~n28496 & n28499 ;
  assign n28510 = ~n28030 & n28438 ;
  assign n28511 = ~n28037 & n28398 ;
  assign n28512 = ~n28510 & ~n28511 ;
  assign n28513 = \P2_P2_DataWidth_reg[1]/NET0131  & ~n28512 ;
  assign n28501 = ~n28387 & ~n28401 ;
  assign n28502 = ~n28016 & ~n28501 ;
  assign n28503 = \P2_P2_InstQueue_reg[15][4]/NET0131  & ~n28387 ;
  assign n28504 = ~n28401 & n28503 ;
  assign n28505 = ~n28502 & ~n28504 ;
  assign n28514 = \P2_P2_DataWidth_reg[1]/NET0131  & ~n28460 ;
  assign n28515 = ~n28505 & ~n28514 ;
  assign n28516 = ~n28513 & ~n28515 ;
  assign n28517 = n26794 & ~n28516 ;
  assign n28507 = ~n26417 & n28387 ;
  assign n28508 = ~n28503 & ~n28507 ;
  assign n28509 = n27613 & ~n28508 ;
  assign n28506 = n27977 & ~n28505 ;
  assign n28518 = \P2_P2_InstQueue_reg[15][4]/NET0131  & ~n28050 ;
  assign n28519 = ~n28506 & ~n28518 ;
  assign n28520 = ~n28509 & n28519 ;
  assign n28521 = ~n28517 & n28520 ;
  assign n28532 = ~n28030 & n28401 ;
  assign n28533 = ~n28037 & n28387 ;
  assign n28534 = ~n28532 & ~n28533 ;
  assign n28535 = \P2_P2_DataWidth_reg[1]/NET0131  & ~n28534 ;
  assign n28522 = ~\P2_P2_InstQueueWr_Addr_reg[3]/NET0131  & n28033 ;
  assign n28523 = ~n28385 & ~n28522 ;
  assign n28524 = ~n28016 & ~n28523 ;
  assign n28525 = \P2_P2_InstQueue_reg[1][4]/NET0131  & ~n28522 ;
  assign n28526 = ~n28385 & n28525 ;
  assign n28527 = ~n28524 & ~n28526 ;
  assign n28536 = \P2_P2_DataWidth_reg[1]/NET0131  & ~n28501 ;
  assign n28537 = ~n28527 & ~n28536 ;
  assign n28538 = ~n28535 & ~n28537 ;
  assign n28539 = n26794 & ~n28538 ;
  assign n28529 = ~n26417 & n28522 ;
  assign n28530 = ~n28525 & ~n28529 ;
  assign n28531 = n27613 & ~n28530 ;
  assign n28528 = n27977 & ~n28527 ;
  assign n28540 = \P2_P2_InstQueue_reg[1][4]/NET0131  & ~n28050 ;
  assign n28541 = ~n28528 & ~n28540 ;
  assign n28542 = ~n28531 & n28541 ;
  assign n28543 = ~n28539 & n28542 ;
  assign n28554 = ~n28030 & n28387 ;
  assign n28555 = ~n28037 & n28385 ;
  assign n28556 = ~n28554 & ~n28555 ;
  assign n28557 = \P2_P2_DataWidth_reg[1]/NET0131  & ~n28556 ;
  assign n28544 = ~\P2_P2_InstQueueWr_Addr_reg[3]/NET0131  & n27982 ;
  assign n28545 = ~n28522 & ~n28544 ;
  assign n28546 = ~n28016 & ~n28545 ;
  assign n28547 = \P2_P2_InstQueue_reg[2][4]/NET0131  & ~n28544 ;
  assign n28548 = ~n28522 & n28547 ;
  assign n28549 = ~n28546 & ~n28548 ;
  assign n28558 = \P2_P2_DataWidth_reg[1]/NET0131  & ~n28388 ;
  assign n28559 = ~n28549 & ~n28558 ;
  assign n28560 = ~n28557 & ~n28559 ;
  assign n28561 = n26794 & ~n28560 ;
  assign n28551 = ~n26417 & n28544 ;
  assign n28552 = ~n28547 & ~n28551 ;
  assign n28553 = n27613 & ~n28552 ;
  assign n28550 = n27977 & ~n28549 ;
  assign n28562 = \P2_P2_InstQueue_reg[2][4]/NET0131  & ~n28050 ;
  assign n28563 = ~n28550 & ~n28562 ;
  assign n28564 = ~n28553 & n28563 ;
  assign n28565 = ~n28561 & n28564 ;
  assign n28576 = ~n28030 & n28385 ;
  assign n28577 = ~n28037 & n28522 ;
  assign n28578 = ~n28576 & ~n28577 ;
  assign n28579 = \P2_P2_DataWidth_reg[1]/NET0131  & ~n28578 ;
  assign n28566 = ~\P2_P2_InstQueueWr_Addr_reg[3]/NET0131  & n27979 ;
  assign n28567 = ~n28544 & ~n28566 ;
  assign n28568 = ~n28016 & ~n28567 ;
  assign n28569 = \P2_P2_InstQueue_reg[3][4]/NET0131  & ~n28566 ;
  assign n28570 = ~n28544 & n28569 ;
  assign n28571 = ~n28568 & ~n28570 ;
  assign n28580 = \P2_P2_DataWidth_reg[1]/NET0131  & ~n28523 ;
  assign n28581 = ~n28571 & ~n28580 ;
  assign n28582 = ~n28579 & ~n28581 ;
  assign n28583 = n26794 & ~n28582 ;
  assign n28573 = ~n26417 & n28566 ;
  assign n28574 = ~n28569 & ~n28573 ;
  assign n28575 = n27613 & ~n28574 ;
  assign n28572 = n27977 & ~n28571 ;
  assign n28584 = \P2_P2_InstQueue_reg[3][4]/NET0131  & ~n28050 ;
  assign n28585 = ~n28572 & ~n28584 ;
  assign n28586 = ~n28575 & n28585 ;
  assign n28587 = ~n28583 & n28586 ;
  assign n28598 = ~n28030 & n28522 ;
  assign n28599 = ~n28037 & n28544 ;
  assign n28600 = ~n28598 & ~n28599 ;
  assign n28601 = \P2_P2_DataWidth_reg[1]/NET0131  & ~n28600 ;
  assign n28588 = ~\P2_P2_InstQueueWr_Addr_reg[3]/NET0131  & n28437 ;
  assign n28589 = ~n28566 & ~n28588 ;
  assign n28590 = ~n28016 & ~n28589 ;
  assign n28591 = \P2_P2_InstQueue_reg[4][4]/NET0131  & ~n28588 ;
  assign n28592 = ~n28566 & n28591 ;
  assign n28593 = ~n28590 & ~n28592 ;
  assign n28602 = \P2_P2_DataWidth_reg[1]/NET0131  & ~n28545 ;
  assign n28603 = ~n28593 & ~n28602 ;
  assign n28604 = ~n28601 & ~n28603 ;
  assign n28605 = n26794 & ~n28604 ;
  assign n28595 = ~n26417 & n28588 ;
  assign n28596 = ~n28591 & ~n28595 ;
  assign n28597 = n27613 & ~n28596 ;
  assign n28594 = n27977 & ~n28593 ;
  assign n28606 = \P2_P2_InstQueue_reg[4][4]/NET0131  & ~n28050 ;
  assign n28607 = ~n28594 & ~n28606 ;
  assign n28608 = ~n28597 & n28607 ;
  assign n28609 = ~n28605 & n28608 ;
  assign n28620 = ~n28030 & n28544 ;
  assign n28621 = ~n28037 & n28566 ;
  assign n28622 = ~n28620 & ~n28621 ;
  assign n28623 = \P2_P2_DataWidth_reg[1]/NET0131  & ~n28622 ;
  assign n28610 = ~\P2_P2_InstQueueWr_Addr_reg[3]/NET0131  & n28397 ;
  assign n28611 = ~n28588 & ~n28610 ;
  assign n28612 = ~n28016 & ~n28611 ;
  assign n28613 = \P2_P2_InstQueue_reg[5][4]/NET0131  & ~n28610 ;
  assign n28614 = ~n28588 & n28613 ;
  assign n28615 = ~n28612 & ~n28614 ;
  assign n28624 = \P2_P2_DataWidth_reg[1]/NET0131  & ~n28567 ;
  assign n28625 = ~n28615 & ~n28624 ;
  assign n28626 = ~n28623 & ~n28625 ;
  assign n28627 = n26794 & ~n28626 ;
  assign n28617 = ~n26417 & n28610 ;
  assign n28618 = ~n28613 & ~n28617 ;
  assign n28619 = n27613 & ~n28618 ;
  assign n28616 = n27977 & ~n28615 ;
  assign n28628 = \P2_P2_InstQueue_reg[5][4]/NET0131  & ~n28050 ;
  assign n28629 = ~n28616 & ~n28628 ;
  assign n28630 = ~n28619 & n28629 ;
  assign n28631 = ~n28627 & n28630 ;
  assign n28642 = ~n28030 & n28566 ;
  assign n28643 = ~n28037 & n28588 ;
  assign n28644 = ~n28642 & ~n28643 ;
  assign n28645 = \P2_P2_DataWidth_reg[1]/NET0131  & ~n28644 ;
  assign n28632 = ~\P2_P2_InstQueueWr_Addr_reg[3]/NET0131  & n28400 ;
  assign n28633 = ~n28610 & ~n28632 ;
  assign n28634 = ~n28016 & ~n28633 ;
  assign n28635 = \P2_P2_InstQueue_reg[6][4]/NET0131  & ~n28632 ;
  assign n28636 = ~n28610 & n28635 ;
  assign n28637 = ~n28634 & ~n28636 ;
  assign n28646 = \P2_P2_DataWidth_reg[1]/NET0131  & ~n28589 ;
  assign n28647 = ~n28637 & ~n28646 ;
  assign n28648 = ~n28645 & ~n28647 ;
  assign n28649 = n26794 & ~n28648 ;
  assign n28639 = ~n26417 & n28632 ;
  assign n28640 = ~n28635 & ~n28639 ;
  assign n28641 = n27613 & ~n28640 ;
  assign n28638 = n27977 & ~n28637 ;
  assign n28650 = \P2_P2_InstQueue_reg[6][4]/NET0131  & ~n28050 ;
  assign n28651 = ~n28638 & ~n28650 ;
  assign n28652 = ~n28641 & n28651 ;
  assign n28653 = ~n28649 & n28652 ;
  assign n28663 = ~n28030 & n28588 ;
  assign n28664 = ~n28037 & n28610 ;
  assign n28665 = ~n28663 & ~n28664 ;
  assign n28666 = \P2_P2_DataWidth_reg[1]/NET0131  & ~n28665 ;
  assign n28654 = ~n28423 & ~n28632 ;
  assign n28655 = ~n28016 & ~n28654 ;
  assign n28656 = \P2_P2_InstQueue_reg[7][4]/NET0131  & ~n28423 ;
  assign n28657 = ~n28632 & n28656 ;
  assign n28658 = ~n28655 & ~n28657 ;
  assign n28667 = \P2_P2_DataWidth_reg[1]/NET0131  & ~n28611 ;
  assign n28668 = ~n28658 & ~n28667 ;
  assign n28669 = ~n28666 & ~n28668 ;
  assign n28670 = n26794 & ~n28669 ;
  assign n28660 = ~n26417 & n28423 ;
  assign n28661 = ~n28656 & ~n28660 ;
  assign n28662 = n27613 & ~n28661 ;
  assign n28659 = n27977 & ~n28658 ;
  assign n28671 = \P2_P2_InstQueue_reg[7][4]/NET0131  & ~n28050 ;
  assign n28672 = ~n28659 & ~n28671 ;
  assign n28673 = ~n28662 & n28672 ;
  assign n28674 = ~n28670 & n28673 ;
  assign n28683 = ~n28030 & n28610 ;
  assign n28684 = ~n28037 & n28632 ;
  assign n28685 = ~n28683 & ~n28684 ;
  assign n28686 = \P2_P2_DataWidth_reg[1]/NET0131  & ~n28685 ;
  assign n28675 = ~n28016 & ~n28428 ;
  assign n28676 = \P2_P2_InstQueue_reg[8][4]/NET0131  & ~n28027 ;
  assign n28677 = ~n28423 & n28676 ;
  assign n28678 = ~n28675 & ~n28677 ;
  assign n28687 = \P2_P2_DataWidth_reg[1]/NET0131  & ~n28633 ;
  assign n28688 = ~n28678 & ~n28687 ;
  assign n28689 = ~n28686 & ~n28688 ;
  assign n28690 = n26794 & ~n28689 ;
  assign n28680 = ~n26417 & n28027 ;
  assign n28681 = ~n28676 & ~n28680 ;
  assign n28682 = n27613 & ~n28681 ;
  assign n28679 = n27977 & ~n28678 ;
  assign n28691 = \P2_P2_InstQueue_reg[8][4]/NET0131  & ~n28050 ;
  assign n28692 = ~n28679 & ~n28691 ;
  assign n28693 = ~n28682 & n28692 ;
  assign n28694 = ~n28690 & n28693 ;
  assign n28703 = ~n28030 & n28632 ;
  assign n28704 = ~n28037 & n28423 ;
  assign n28705 = ~n28703 & ~n28704 ;
  assign n28706 = \P2_P2_DataWidth_reg[1]/NET0131  & ~n28705 ;
  assign n28695 = ~n28016 & ~n28041 ;
  assign n28696 = \P2_P2_InstQueue_reg[9][4]/NET0131  & ~n28034 ;
  assign n28697 = ~n28027 & n28696 ;
  assign n28698 = ~n28695 & ~n28697 ;
  assign n28707 = \P2_P2_DataWidth_reg[1]/NET0131  & ~n28654 ;
  assign n28708 = ~n28698 & ~n28707 ;
  assign n28709 = ~n28706 & ~n28708 ;
  assign n28710 = n26794 & ~n28709 ;
  assign n28700 = ~n26417 & n28034 ;
  assign n28701 = ~n28696 & ~n28700 ;
  assign n28702 = n27613 & ~n28701 ;
  assign n28699 = n27977 & ~n28698 ;
  assign n28711 = \P2_P2_InstQueue_reg[9][4]/NET0131  & ~n28050 ;
  assign n28712 = ~n28699 & ~n28711 ;
  assign n28713 = ~n28702 & n28712 ;
  assign n28714 = ~n28710 & n28713 ;
  assign n28715 = \P2_P1_lWord_reg[8]/NET0131  & ~n25156 ;
  assign n28716 = \P2_P1_EAX_reg[8]/NET0131  & n24899 ;
  assign n28717 = n11385 & ~n21073 ;
  assign n28718 = n24901 & n28717 ;
  assign n28719 = ~n28716 & ~n28718 ;
  assign n28720 = n11623 & ~n28719 ;
  assign n28721 = ~n28715 & ~n28720 ;
  assign n28722 = \P1_P1_lWord_reg[8]/NET0131  & ~n25165 ;
  assign n28723 = \P1_P1_EAX_reg[8]/NET0131  & n24503 ;
  assign n28724 = ~n7891 & n23947 ;
  assign n28725 = ~n28723 & ~n28724 ;
  assign n28726 = n8355 & ~n28725 ;
  assign n28727 = ~n28722 & ~n28726 ;
  assign n28728 = \P1_P1_uWord_reg[11]/NET0131  & ~n24515 ;
  assign n28732 = \P1_P1_uWord_reg[11]/NET0131  & n25363 ;
  assign n28733 = ~n23970 & ~n28732 ;
  assign n28734 = n15334 & ~n28733 ;
  assign n28729 = ~\P1_P1_EAX_reg[27]/NET0131  & ~n27426 ;
  assign n28730 = ~n27427 & ~n28729 ;
  assign n28731 = n24503 & n28730 ;
  assign n28735 = \P1_P1_uWord_reg[11]/NET0131  & n24505 ;
  assign n28736 = ~n28731 & ~n28735 ;
  assign n28737 = ~n28734 & n28736 ;
  assign n28738 = n8355 & ~n28737 ;
  assign n28739 = ~n28728 & ~n28738 ;
  assign n28740 = ~\P4_addr_reg[11]/NET0131  & n15734 ;
  assign n28741 = n18666 & ~n28740 ;
  assign n28743 = ~n15744 & ~n28741 ;
  assign n28779 = \P4_IR_reg[11]/NET0131  & \P4_reg1_reg[11]/NET0131  ;
  assign n28780 = ~\P4_IR_reg[11]/NET0131  & ~\P4_reg1_reg[11]/NET0131  ;
  assign n28781 = ~n28779 & ~n28780 ;
  assign n28782 = ~\P4_IR_reg[10]/NET0131  & ~\P4_reg1_reg[10]/NET0131  ;
  assign n28783 = \P4_IR_reg[10]/NET0131  & \P4_reg1_reg[10]/NET0131  ;
  assign n28784 = ~\P4_IR_reg[9]/NET0131  & ~\P4_reg1_reg[9]/NET0131  ;
  assign n28785 = \P4_IR_reg[9]/NET0131  & \P4_reg1_reg[9]/NET0131  ;
  assign n28786 = ~\P4_IR_reg[8]/NET0131  & ~\P4_reg1_reg[8]/NET0131  ;
  assign n28787 = \P4_IR_reg[8]/NET0131  & \P4_reg1_reg[8]/NET0131  ;
  assign n28788 = ~\P4_IR_reg[7]/NET0131  & ~\P4_reg1_reg[7]/NET0131  ;
  assign n28789 = \P4_IR_reg[7]/NET0131  & \P4_reg1_reg[7]/NET0131  ;
  assign n28790 = ~\P4_IR_reg[6]/NET0131  & ~\P4_reg1_reg[6]/NET0131  ;
  assign n28791 = \P4_IR_reg[6]/NET0131  & \P4_reg1_reg[6]/NET0131  ;
  assign n28792 = ~\P4_IR_reg[5]/NET0131  & ~\P4_reg1_reg[5]/NET0131  ;
  assign n28793 = \P4_IR_reg[5]/NET0131  & \P4_reg1_reg[5]/NET0131  ;
  assign n28794 = ~n27867 & ~n27875 ;
  assign n28795 = ~n27868 & ~n28794 ;
  assign n28796 = ~n28793 & ~n28795 ;
  assign n28797 = ~n28792 & ~n28796 ;
  assign n28798 = ~n28791 & ~n28797 ;
  assign n28799 = ~n28790 & ~n28798 ;
  assign n28800 = ~n28789 & ~n28799 ;
  assign n28801 = ~n28788 & ~n28800 ;
  assign n28802 = ~n28787 & ~n28801 ;
  assign n28803 = ~n28786 & ~n28802 ;
  assign n28804 = ~n28785 & ~n28803 ;
  assign n28805 = ~n28784 & ~n28804 ;
  assign n28806 = ~n28783 & ~n28805 ;
  assign n28807 = ~n28782 & ~n28806 ;
  assign n28809 = n28781 & n28807 ;
  assign n28808 = ~n28781 & ~n28807 ;
  assign n28810 = n27804 & ~n28808 ;
  assign n28811 = ~n28809 & n28810 ;
  assign n28745 = \P4_IR_reg[11]/NET0131  & \P4_reg2_reg[11]/NET0131  ;
  assign n28746 = ~\P4_IR_reg[11]/NET0131  & ~\P4_reg2_reg[11]/NET0131  ;
  assign n28747 = ~n28745 & ~n28746 ;
  assign n28748 = ~\P4_IR_reg[10]/NET0131  & ~\P4_reg2_reg[10]/NET0131  ;
  assign n28749 = \P4_IR_reg[10]/NET0131  & \P4_reg2_reg[10]/NET0131  ;
  assign n28750 = ~\P4_IR_reg[9]/NET0131  & ~\P4_reg2_reg[9]/NET0131  ;
  assign n28751 = \P4_IR_reg[9]/NET0131  & \P4_reg2_reg[9]/NET0131  ;
  assign n28752 = ~\P4_IR_reg[8]/NET0131  & ~\P4_reg2_reg[8]/NET0131  ;
  assign n28753 = \P4_IR_reg[8]/NET0131  & \P4_reg2_reg[8]/NET0131  ;
  assign n28754 = ~\P4_IR_reg[7]/NET0131  & ~\P4_reg2_reg[7]/NET0131  ;
  assign n28755 = \P4_IR_reg[7]/NET0131  & \P4_reg2_reg[7]/NET0131  ;
  assign n28756 = ~\P4_IR_reg[6]/NET0131  & ~\P4_reg2_reg[6]/NET0131  ;
  assign n28757 = \P4_IR_reg[6]/NET0131  & \P4_reg2_reg[6]/NET0131  ;
  assign n28758 = ~\P4_IR_reg[5]/NET0131  & ~\P4_reg2_reg[5]/NET0131  ;
  assign n28759 = \P4_IR_reg[5]/NET0131  & \P4_reg2_reg[5]/NET0131  ;
  assign n28760 = ~n27854 & ~n27862 ;
  assign n28761 = ~n27855 & ~n28760 ;
  assign n28762 = ~n28759 & ~n28761 ;
  assign n28763 = ~n28758 & ~n28762 ;
  assign n28764 = ~n28757 & ~n28763 ;
  assign n28765 = ~n28756 & ~n28764 ;
  assign n28766 = ~n28755 & ~n28765 ;
  assign n28767 = ~n28754 & ~n28766 ;
  assign n28768 = ~n28753 & ~n28767 ;
  assign n28769 = ~n28752 & ~n28768 ;
  assign n28770 = ~n28751 & ~n28769 ;
  assign n28771 = ~n28750 & ~n28770 ;
  assign n28772 = ~n28749 & ~n28771 ;
  assign n28773 = ~n28748 & ~n28772 ;
  assign n28775 = n28747 & n28773 ;
  assign n28774 = ~n28747 & ~n28773 ;
  assign n28776 = n15733 & ~n28774 ;
  assign n28777 = ~n28775 & n28776 ;
  assign n28744 = \P4_addr_reg[11]/NET0131  & n15745 ;
  assign n28778 = \P4_IR_reg[11]/NET0131  & n21786 ;
  assign n28812 = ~n28744 & ~n28778 ;
  assign n28813 = ~n28777 & n28812 ;
  assign n28814 = ~n28811 & n28813 ;
  assign n28815 = ~n28743 & ~n28814 ;
  assign n28742 = n15734 & n28741 ;
  assign n28816 = ~n21972 & ~n28742 ;
  assign n28817 = ~n28815 & n28816 ;
  assign n28818 = ~\P4_addr_reg[13]/NET0131  & n15734 ;
  assign n28819 = n18666 & ~n28818 ;
  assign n28821 = ~n15744 & ~n28819 ;
  assign n28837 = \P4_IR_reg[13]/NET0131  & \P4_reg2_reg[13]/NET0131  ;
  assign n28838 = ~\P4_IR_reg[13]/NET0131  & ~\P4_reg2_reg[13]/NET0131  ;
  assign n28839 = ~n28837 & ~n28838 ;
  assign n28840 = ~\P4_IR_reg[12]/NET0131  & ~\P4_reg2_reg[12]/NET0131  ;
  assign n28841 = \P4_IR_reg[12]/NET0131  & \P4_reg2_reg[12]/NET0131  ;
  assign n28842 = ~n28745 & ~n28773 ;
  assign n28843 = ~n28746 & ~n28842 ;
  assign n28844 = ~n28841 & ~n28843 ;
  assign n28845 = ~n28840 & ~n28844 ;
  assign n28847 = n28839 & n28845 ;
  assign n28846 = ~n28839 & ~n28845 ;
  assign n28848 = n15733 & ~n28846 ;
  assign n28849 = ~n28847 & n28848 ;
  assign n28823 = \P4_IR_reg[13]/NET0131  & \P4_reg1_reg[13]/NET0131  ;
  assign n28824 = ~\P4_IR_reg[13]/NET0131  & ~\P4_reg1_reg[13]/NET0131  ;
  assign n28825 = ~n28823 & ~n28824 ;
  assign n28826 = ~\P4_IR_reg[12]/NET0131  & ~\P4_reg1_reg[12]/NET0131  ;
  assign n28827 = \P4_IR_reg[12]/NET0131  & \P4_reg1_reg[12]/NET0131  ;
  assign n28828 = ~n28779 & ~n28807 ;
  assign n28829 = ~n28780 & ~n28828 ;
  assign n28830 = ~n28827 & ~n28829 ;
  assign n28831 = ~n28826 & ~n28830 ;
  assign n28833 = n28825 & n28831 ;
  assign n28832 = ~n28825 & ~n28831 ;
  assign n28834 = n27804 & ~n28832 ;
  assign n28835 = ~n28833 & n28834 ;
  assign n28822 = \P4_IR_reg[13]/NET0131  & n21786 ;
  assign n28836 = \P4_addr_reg[13]/NET0131  & n15745 ;
  assign n28850 = ~n28822 & ~n28836 ;
  assign n28851 = ~n28835 & n28850 ;
  assign n28852 = ~n28849 & n28851 ;
  assign n28853 = ~n28821 & ~n28852 ;
  assign n28820 = n15734 & n28819 ;
  assign n28854 = ~n23204 & ~n28820 ;
  assign n28855 = ~n28853 & n28854 ;
  assign n28856 = ~\P4_addr_reg[5]/NET0131  & n15734 ;
  assign n28857 = n18666 & ~n28856 ;
  assign n28859 = ~n15744 & ~n28857 ;
  assign n28867 = ~n28758 & ~n28759 ;
  assign n28869 = n28761 & n28867 ;
  assign n28868 = ~n28761 & ~n28867 ;
  assign n28870 = n15733 & ~n28868 ;
  assign n28871 = ~n28869 & n28870 ;
  assign n28861 = ~n28792 & ~n28793 ;
  assign n28863 = n28795 & n28861 ;
  assign n28862 = ~n28795 & ~n28861 ;
  assign n28864 = n27804 & ~n28862 ;
  assign n28865 = ~n28863 & n28864 ;
  assign n28860 = \P4_IR_reg[5]/NET0131  & n21786 ;
  assign n28866 = \P4_addr_reg[5]/NET0131  & n15745 ;
  assign n28872 = ~n28860 & ~n28866 ;
  assign n28873 = ~n28865 & n28872 ;
  assign n28874 = ~n28871 & n28873 ;
  assign n28875 = ~n28859 & ~n28874 ;
  assign n28858 = n15734 & n28857 ;
  assign n28876 = ~n23333 & ~n28858 ;
  assign n28877 = ~n28875 & n28876 ;
  assign n28878 = ~\P4_addr_reg[8]/NET0131  & n15734 ;
  assign n28879 = n18666 & ~n28878 ;
  assign n28881 = ~n15744 & ~n28879 ;
  assign n28889 = ~n28786 & ~n28787 ;
  assign n28891 = n28801 & n28889 ;
  assign n28890 = ~n28801 & ~n28889 ;
  assign n28892 = n27804 & ~n28890 ;
  assign n28893 = ~n28891 & n28892 ;
  assign n28883 = ~n28752 & ~n28753 ;
  assign n28885 = n28767 & n28883 ;
  assign n28884 = ~n28767 & ~n28883 ;
  assign n28886 = n15733 & ~n28884 ;
  assign n28887 = ~n28885 & n28886 ;
  assign n28882 = \P4_IR_reg[8]/NET0131  & n21786 ;
  assign n28888 = \P4_addr_reg[8]/NET0131  & n15745 ;
  assign n28894 = ~n28882 & ~n28888 ;
  assign n28895 = ~n28887 & n28894 ;
  assign n28896 = ~n28893 & n28895 ;
  assign n28897 = ~n28881 & ~n28896 ;
  assign n28880 = n15734 & n28879 ;
  assign n28898 = ~n22981 & ~n28880 ;
  assign n28899 = ~n28897 & n28898 ;
  assign n28900 = ~\P4_addr_reg[9]/NET0131  & n15734 ;
  assign n28901 = n18666 & ~n28900 ;
  assign n28903 = ~n15744 & ~n28901 ;
  assign n28911 = ~n28784 & ~n28785 ;
  assign n28913 = n28803 & n28911 ;
  assign n28912 = ~n28803 & ~n28911 ;
  assign n28914 = n27804 & ~n28912 ;
  assign n28915 = ~n28913 & n28914 ;
  assign n28905 = ~n28750 & ~n28751 ;
  assign n28907 = n28769 & n28905 ;
  assign n28906 = ~n28769 & ~n28905 ;
  assign n28908 = n15733 & ~n28906 ;
  assign n28909 = ~n28907 & n28908 ;
  assign n28904 = \P4_addr_reg[9]/NET0131  & n15745 ;
  assign n28910 = \P4_IR_reg[9]/NET0131  & n21786 ;
  assign n28916 = ~n28904 & ~n28910 ;
  assign n28917 = ~n28909 & n28916 ;
  assign n28918 = ~n28915 & n28917 ;
  assign n28919 = ~n28903 & ~n28918 ;
  assign n28902 = n15734 & n28901 ;
  assign n28920 = ~n23397 & ~n28902 ;
  assign n28921 = ~n28919 & n28920 ;
  assign n28929 = \P1_buf2_reg[7]/NET0131  & ~n27934 ;
  assign n28930 = \P1_buf1_reg[7]/NET0131  & n27934 ;
  assign n28931 = ~n28929 & ~n28930 ;
  assign n28932 = ~n27905 & ~n28931 ;
  assign n28923 = \P1_P2_InstQueue_reg[11][7]/NET0131  & ~n27901 ;
  assign n28933 = ~n27904 & n28923 ;
  assign n28934 = ~n28932 & ~n28933 ;
  assign n28927 = ~n27898 & n27960 ;
  assign n28928 = ~n25928 & ~n27898 ;
  assign n28935 = ~n28927 & ~n28928 ;
  assign n28936 = ~n28934 & n28935 ;
  assign n28924 = ~n25540 & n27901 ;
  assign n28925 = ~n28923 & ~n28924 ;
  assign n28926 = n27608 & ~n28925 ;
  assign n28922 = \P1_P2_InstQueue_reg[11][7]/NET0131  & ~n27972 ;
  assign n28937 = \P1_buf2_reg[23]/NET0131  & ~n27934 ;
  assign n28938 = \P1_buf1_reg[23]/NET0131  & n27934 ;
  assign n28939 = ~n28937 & ~n28938 ;
  assign n28940 = \P1_P2_DataWidth_reg[1]/NET0131  & ~n28939 ;
  assign n28941 = n25928 & n27952 ;
  assign n28942 = n28940 & n28941 ;
  assign n28943 = ~n28922 & ~n28942 ;
  assign n28944 = ~n28926 & n28943 ;
  assign n28945 = ~n28936 & n28944 ;
  assign n28953 = \P2_P2_InstQueue_reg[11][7]/NET0131  & ~n27980 ;
  assign n28958 = ~n26354 & n27980 ;
  assign n28959 = ~n28953 & ~n28958 ;
  assign n28960 = n27613 & ~n28959 ;
  assign n28949 = \P2_buf2_reg[7]/NET0131  & ~n28013 ;
  assign n28950 = \P2_buf1_reg[7]/NET0131  & n28013 ;
  assign n28951 = ~n28949 & ~n28950 ;
  assign n28952 = ~n27984 & ~n28951 ;
  assign n28954 = ~n27983 & n28953 ;
  assign n28955 = ~n28952 & ~n28954 ;
  assign n28947 = ~n27977 & n28042 ;
  assign n28948 = ~n26794 & ~n27977 ;
  assign n28956 = ~n28947 & ~n28948 ;
  assign n28957 = ~n28955 & n28956 ;
  assign n28946 = \P2_P2_InstQueue_reg[11][7]/NET0131  & ~n28050 ;
  assign n28961 = \P2_buf2_reg[23]/NET0131  & ~n28013 ;
  assign n28962 = \P2_buf1_reg[23]/NET0131  & n28013 ;
  assign n28963 = ~n28961 & ~n28962 ;
  assign n28964 = \P2_P2_DataWidth_reg[1]/NET0131  & ~n28963 ;
  assign n28965 = n26794 & n28034 ;
  assign n28966 = n28964 & n28965 ;
  assign n28967 = ~n28946 & ~n28966 ;
  assign n28968 = ~n28957 & n28967 ;
  assign n28969 = ~n28960 & n28968 ;
  assign n28970 = ~\P4_addr_reg[10]/NET0131  & n15734 ;
  assign n28971 = n18666 & ~n28970 ;
  assign n28973 = ~n15744 & ~n28971 ;
  assign n28981 = ~n28748 & ~n28749 ;
  assign n28983 = n28771 & n28981 ;
  assign n28982 = ~n28771 & ~n28981 ;
  assign n28984 = n15733 & ~n28982 ;
  assign n28985 = ~n28983 & n28984 ;
  assign n28975 = ~n28782 & ~n28783 ;
  assign n28977 = n28805 & n28975 ;
  assign n28976 = ~n28805 & ~n28975 ;
  assign n28978 = n27804 & ~n28976 ;
  assign n28979 = ~n28977 & n28978 ;
  assign n28974 = \P4_IR_reg[10]/NET0131  & n21786 ;
  assign n28980 = \P4_addr_reg[10]/NET0131  & n15745 ;
  assign n28986 = ~n28974 & ~n28980 ;
  assign n28987 = ~n28979 & n28986 ;
  assign n28988 = ~n28985 & n28987 ;
  assign n28989 = ~n28973 & ~n28988 ;
  assign n28972 = n15734 & n28971 ;
  assign n28990 = ~n22415 & ~n28972 ;
  assign n28991 = ~n28989 & n28990 ;
  assign n28998 = ~n28058 & ~n28931 ;
  assign n28993 = \P1_P2_InstQueue_reg[0][7]/NET0131  & ~n28055 ;
  assign n28999 = ~n28057 & n28993 ;
  assign n29000 = ~n28998 & ~n28999 ;
  assign n28997 = ~n27898 & n28073 ;
  assign n29001 = ~n28928 & ~n28997 ;
  assign n29002 = ~n29000 & n29001 ;
  assign n28994 = ~n25540 & n28055 ;
  assign n28995 = ~n28993 & ~n28994 ;
  assign n28996 = n27608 & ~n28995 ;
  assign n28992 = \P1_P2_InstQueue_reg[0][7]/NET0131  & ~n27972 ;
  assign n29003 = n25928 & n28068 ;
  assign n29004 = n28940 & n29003 ;
  assign n29005 = ~n28992 & ~n29004 ;
  assign n29006 = ~n28996 & n29005 ;
  assign n29007 = ~n29002 & n29006 ;
  assign n29014 = ~n28084 & ~n28931 ;
  assign n29009 = \P1_P2_InstQueue_reg[10][7]/NET0131  & ~n27904 ;
  assign n29015 = ~n27952 & n29009 ;
  assign n29016 = ~n29014 & ~n29015 ;
  assign n29013 = ~n27898 & n28096 ;
  assign n29017 = ~n28928 & ~n29013 ;
  assign n29018 = ~n29016 & n29017 ;
  assign n29010 = ~n25540 & n27904 ;
  assign n29011 = ~n29009 & ~n29010 ;
  assign n29012 = n27608 & ~n29011 ;
  assign n29008 = \P1_P2_InstQueue_reg[10][7]/NET0131  & ~n27972 ;
  assign n29019 = n25928 & n27945 ;
  assign n29020 = n28940 & n29019 ;
  assign n29021 = ~n29008 & ~n29020 ;
  assign n29022 = ~n29012 & n29021 ;
  assign n29023 = ~n29018 & n29022 ;
  assign n29030 = ~n28109 & ~n28931 ;
  assign n29025 = \P1_P2_InstQueue_reg[12][7]/NET0131  & ~n28108 ;
  assign n29031 = ~n27901 & n29025 ;
  assign n29032 = ~n29030 & ~n29031 ;
  assign n29029 = ~n27898 & n28119 ;
  assign n29033 = ~n28928 & ~n29029 ;
  assign n29034 = ~n29032 & n29033 ;
  assign n29026 = ~n25540 & n28108 ;
  assign n29027 = ~n29025 & ~n29026 ;
  assign n29028 = n27608 & ~n29027 ;
  assign n29024 = \P1_P2_InstQueue_reg[12][7]/NET0131  & ~n27972 ;
  assign n29035 = n25928 & n27904 ;
  assign n29036 = n28940 & n29035 ;
  assign n29037 = ~n29024 & ~n29036 ;
  assign n29038 = ~n29028 & n29037 ;
  assign n29039 = ~n29034 & n29038 ;
  assign n29046 = ~n28130 & ~n28931 ;
  assign n29041 = \P1_P2_InstQueue_reg[13][7]/NET0131  & ~n28065 ;
  assign n29047 = ~n28108 & n29041 ;
  assign n29048 = ~n29046 & ~n29047 ;
  assign n29045 = ~n27898 & n28140 ;
  assign n29049 = ~n28928 & ~n29045 ;
  assign n29050 = ~n29048 & n29049 ;
  assign n29042 = ~n25540 & n28065 ;
  assign n29043 = ~n29041 & ~n29042 ;
  assign n29044 = n27608 & ~n29043 ;
  assign n29040 = \P1_P2_InstQueue_reg[13][7]/NET0131  & ~n27972 ;
  assign n29051 = n25928 & n27901 ;
  assign n29052 = n28940 & n29051 ;
  assign n29053 = ~n29040 & ~n29052 ;
  assign n29054 = ~n29044 & n29053 ;
  assign n29055 = ~n29050 & n29054 ;
  assign n29062 = ~n28072 & ~n28931 ;
  assign n29057 = \P1_P2_InstQueue_reg[14][7]/NET0131  & ~n28068 ;
  assign n29063 = ~n28065 & n29057 ;
  assign n29064 = ~n29062 & ~n29063 ;
  assign n29061 = ~n27898 & n28160 ;
  assign n29065 = ~n28928 & ~n29061 ;
  assign n29066 = ~n29064 & n29065 ;
  assign n29058 = ~n25540 & n28068 ;
  assign n29059 = ~n29057 & ~n29058 ;
  assign n29060 = n27608 & ~n29059 ;
  assign n29056 = \P1_P2_InstQueue_reg[14][7]/NET0131  & ~n27972 ;
  assign n29067 = n25928 & n28108 ;
  assign n29068 = n28940 & n29067 ;
  assign n29069 = ~n29056 & ~n29068 ;
  assign n29070 = ~n29060 & n29069 ;
  assign n29071 = ~n29066 & n29070 ;
  assign n29078 = ~n28171 & ~n28931 ;
  assign n29073 = \P1_P2_InstQueue_reg[15][7]/NET0131  & ~n28057 ;
  assign n29079 = ~n28068 & n29073 ;
  assign n29080 = ~n29078 & ~n29079 ;
  assign n29077 = ~n27898 & n28181 ;
  assign n29081 = ~n28928 & ~n29077 ;
  assign n29082 = ~n29080 & n29081 ;
  assign n29074 = ~n25540 & n28057 ;
  assign n29075 = ~n29073 & ~n29074 ;
  assign n29076 = n27608 & ~n29075 ;
  assign n29072 = \P1_P2_InstQueue_reg[15][7]/NET0131  & ~n27972 ;
  assign n29083 = n25928 & n28065 ;
  assign n29084 = n28940 & n29083 ;
  assign n29085 = ~n29072 & ~n29084 ;
  assign n29086 = ~n29076 & n29085 ;
  assign n29087 = ~n29082 & n29086 ;
  assign n29094 = ~n28193 & ~n28931 ;
  assign n29089 = \P1_P2_InstQueue_reg[1][7]/NET0131  & ~n28192 ;
  assign n29095 = ~n28055 & n29089 ;
  assign n29096 = ~n29094 & ~n29095 ;
  assign n29093 = ~n27898 & n28203 ;
  assign n29097 = ~n28928 & ~n29093 ;
  assign n29098 = ~n29096 & n29097 ;
  assign n29090 = ~n25540 & n28192 ;
  assign n29091 = ~n29089 & ~n29090 ;
  assign n29092 = n27608 & ~n29091 ;
  assign n29088 = \P1_P2_InstQueue_reg[1][7]/NET0131  & ~n27972 ;
  assign n29099 = n25928 & n28057 ;
  assign n29100 = n28940 & n29099 ;
  assign n29101 = ~n29088 & ~n29100 ;
  assign n29102 = ~n29092 & n29101 ;
  assign n29103 = ~n29098 & n29102 ;
  assign n29110 = ~n28215 & ~n28931 ;
  assign n29105 = \P1_P2_InstQueue_reg[2][7]/NET0131  & ~n28214 ;
  assign n29111 = ~n28192 & n29105 ;
  assign n29112 = ~n29110 & ~n29111 ;
  assign n29109 = ~n27898 & n28225 ;
  assign n29113 = ~n28928 & ~n29109 ;
  assign n29114 = ~n29112 & n29113 ;
  assign n29106 = ~n25540 & n28214 ;
  assign n29107 = ~n29105 & ~n29106 ;
  assign n29108 = n27608 & ~n29107 ;
  assign n29104 = \P1_P2_InstQueue_reg[2][7]/NET0131  & ~n27972 ;
  assign n29115 = n25928 & n28055 ;
  assign n29116 = n28940 & n29115 ;
  assign n29117 = ~n29104 & ~n29116 ;
  assign n29118 = ~n29108 & n29117 ;
  assign n29119 = ~n29114 & n29118 ;
  assign n29126 = ~n28237 & ~n28931 ;
  assign n29121 = \P1_P2_InstQueue_reg[3][7]/NET0131  & ~n28236 ;
  assign n29127 = ~n28214 & n29121 ;
  assign n29128 = ~n29126 & ~n29127 ;
  assign n29125 = ~n27898 & n28247 ;
  assign n29129 = ~n28928 & ~n29125 ;
  assign n29130 = ~n29128 & n29129 ;
  assign n29122 = ~n25540 & n28236 ;
  assign n29123 = ~n29121 & ~n29122 ;
  assign n29124 = n27608 & ~n29123 ;
  assign n29120 = \P1_P2_InstQueue_reg[3][7]/NET0131  & ~n27972 ;
  assign n29131 = n25928 & n28192 ;
  assign n29132 = n28940 & n29131 ;
  assign n29133 = ~n29120 & ~n29132 ;
  assign n29134 = ~n29124 & n29133 ;
  assign n29135 = ~n29130 & n29134 ;
  assign n29142 = ~n28259 & ~n28931 ;
  assign n29137 = \P1_P2_InstQueue_reg[4][7]/NET0131  & ~n28258 ;
  assign n29143 = ~n28236 & n29137 ;
  assign n29144 = ~n29142 & ~n29143 ;
  assign n29141 = ~n27898 & n28269 ;
  assign n29145 = ~n28928 & ~n29141 ;
  assign n29146 = ~n29144 & n29145 ;
  assign n29138 = ~n25540 & n28258 ;
  assign n29139 = ~n29137 & ~n29138 ;
  assign n29140 = n27608 & ~n29139 ;
  assign n29136 = \P1_P2_InstQueue_reg[4][7]/NET0131  & ~n27972 ;
  assign n29147 = n25928 & n28214 ;
  assign n29148 = n28940 & n29147 ;
  assign n29149 = ~n29136 & ~n29148 ;
  assign n29150 = ~n29140 & n29149 ;
  assign n29151 = ~n29146 & n29150 ;
  assign n29158 = ~n28281 & ~n28931 ;
  assign n29153 = \P1_P2_InstQueue_reg[5][7]/NET0131  & ~n28280 ;
  assign n29159 = ~n28258 & n29153 ;
  assign n29160 = ~n29158 & ~n29159 ;
  assign n29157 = ~n27898 & n28291 ;
  assign n29161 = ~n28928 & ~n29157 ;
  assign n29162 = ~n29160 & n29161 ;
  assign n29154 = ~n25540 & n28280 ;
  assign n29155 = ~n29153 & ~n29154 ;
  assign n29156 = n27608 & ~n29155 ;
  assign n29152 = \P1_P2_InstQueue_reg[5][7]/NET0131  & ~n27972 ;
  assign n29163 = n25928 & n28236 ;
  assign n29164 = n28940 & n29163 ;
  assign n29165 = ~n29152 & ~n29164 ;
  assign n29166 = ~n29156 & n29165 ;
  assign n29167 = ~n29162 & n29166 ;
  assign n29174 = ~n28303 & ~n28931 ;
  assign n29169 = \P1_P2_InstQueue_reg[6][7]/NET0131  & ~n28302 ;
  assign n29175 = ~n28280 & n29169 ;
  assign n29176 = ~n29174 & ~n29175 ;
  assign n29173 = ~n27898 & n28313 ;
  assign n29177 = ~n28928 & ~n29173 ;
  assign n29178 = ~n29176 & n29177 ;
  assign n29170 = ~n25540 & n28302 ;
  assign n29171 = ~n29169 & ~n29170 ;
  assign n29172 = n27608 & ~n29171 ;
  assign n29168 = \P1_P2_InstQueue_reg[6][7]/NET0131  & ~n27972 ;
  assign n29179 = n25928 & n28258 ;
  assign n29180 = n28940 & n29179 ;
  assign n29181 = ~n29168 & ~n29180 ;
  assign n29182 = ~n29172 & n29181 ;
  assign n29183 = ~n29178 & n29182 ;
  assign n29190 = ~n28324 & ~n28931 ;
  assign n29185 = \P1_P2_InstQueue_reg[7][7]/NET0131  & ~n28090 ;
  assign n29191 = ~n28302 & n29185 ;
  assign n29192 = ~n29190 & ~n29191 ;
  assign n29189 = ~n27898 & n28334 ;
  assign n29193 = ~n28928 & ~n29189 ;
  assign n29194 = ~n29192 & n29193 ;
  assign n29186 = ~n25540 & n28090 ;
  assign n29187 = ~n29185 & ~n29186 ;
  assign n29188 = n27608 & ~n29187 ;
  assign n29184 = \P1_P2_InstQueue_reg[7][7]/NET0131  & ~n27972 ;
  assign n29195 = n25928 & n28280 ;
  assign n29196 = n28940 & n29195 ;
  assign n29197 = ~n29184 & ~n29196 ;
  assign n29198 = ~n29188 & n29197 ;
  assign n29199 = ~n29194 & n29198 ;
  assign n29206 = ~n28095 & ~n28931 ;
  assign n29201 = \P1_P2_InstQueue_reg[8][7]/NET0131  & ~n27945 ;
  assign n29207 = ~n28090 & n29201 ;
  assign n29208 = ~n29206 & ~n29207 ;
  assign n29205 = ~n27898 & n28354 ;
  assign n29209 = ~n28928 & ~n29205 ;
  assign n29210 = ~n29208 & n29209 ;
  assign n29202 = ~n25540 & n27945 ;
  assign n29203 = ~n29201 & ~n29202 ;
  assign n29204 = n27608 & ~n29203 ;
  assign n29200 = \P1_P2_InstQueue_reg[8][7]/NET0131  & ~n27972 ;
  assign n29211 = n25928 & n28302 ;
  assign n29212 = n28940 & n29211 ;
  assign n29213 = ~n29200 & ~n29212 ;
  assign n29214 = ~n29204 & n29213 ;
  assign n29215 = ~n29210 & n29214 ;
  assign n29222 = ~n27959 & ~n28931 ;
  assign n29217 = \P1_P2_InstQueue_reg[9][7]/NET0131  & ~n27952 ;
  assign n29223 = ~n27945 & n29217 ;
  assign n29224 = ~n29222 & ~n29223 ;
  assign n29221 = ~n27898 & n28374 ;
  assign n29225 = ~n28928 & ~n29221 ;
  assign n29226 = ~n29224 & n29225 ;
  assign n29218 = ~n25540 & n27952 ;
  assign n29219 = ~n29217 & ~n29218 ;
  assign n29220 = n27608 & ~n29219 ;
  assign n29216 = \P1_P2_InstQueue_reg[9][7]/NET0131  & ~n27972 ;
  assign n29227 = n25928 & n28090 ;
  assign n29228 = n28940 & n29227 ;
  assign n29229 = ~n29216 & ~n29228 ;
  assign n29230 = ~n29220 & n29229 ;
  assign n29231 = ~n29226 & n29230 ;
  assign n29235 = \P2_P2_InstQueue_reg[0][7]/NET0131  & ~n28385 ;
  assign n29240 = ~n26354 & n28385 ;
  assign n29241 = ~n29235 & ~n29240 ;
  assign n29242 = n27613 & ~n29241 ;
  assign n29234 = ~n28388 & ~n28951 ;
  assign n29236 = ~n28387 & n29235 ;
  assign n29237 = ~n29234 & ~n29236 ;
  assign n29233 = ~n27977 & n28406 ;
  assign n29238 = ~n28948 & ~n29233 ;
  assign n29239 = ~n29237 & n29238 ;
  assign n29232 = \P2_P2_InstQueue_reg[0][7]/NET0131  & ~n28050 ;
  assign n29243 = n26794 & n28401 ;
  assign n29244 = n28964 & n29243 ;
  assign n29245 = ~n29232 & ~n29244 ;
  assign n29246 = ~n29239 & n29245 ;
  assign n29247 = ~n29242 & n29246 ;
  assign n29251 = \P2_P2_InstQueue_reg[10][7]/NET0131  & ~n27983 ;
  assign n29256 = ~n26354 & n27983 ;
  assign n29257 = ~n29251 & ~n29256 ;
  assign n29258 = n27613 & ~n29257 ;
  assign n29250 = ~n28414 & ~n28951 ;
  assign n29252 = ~n28034 & n29251 ;
  assign n29253 = ~n29250 & ~n29252 ;
  assign n29249 = ~n27977 & n28429 ;
  assign n29254 = ~n28948 & ~n29249 ;
  assign n29255 = ~n29253 & n29254 ;
  assign n29248 = \P2_P2_InstQueue_reg[10][7]/NET0131  & ~n28050 ;
  assign n29259 = n26794 & n28027 ;
  assign n29260 = n28964 & n29259 ;
  assign n29261 = ~n29248 & ~n29260 ;
  assign n29262 = ~n29255 & n29261 ;
  assign n29263 = ~n29258 & n29262 ;
  assign n29267 = \P2_P2_InstQueue_reg[12][7]/NET0131  & ~n28438 ;
  assign n29272 = ~n26354 & n28438 ;
  assign n29273 = ~n29267 & ~n29272 ;
  assign n29274 = n27613 & ~n29273 ;
  assign n29266 = ~n28439 & ~n28951 ;
  assign n29268 = ~n27980 & n29267 ;
  assign n29269 = ~n29266 & ~n29268 ;
  assign n29265 = ~n27977 & n28452 ;
  assign n29270 = ~n28948 & ~n29265 ;
  assign n29271 = ~n29269 & n29270 ;
  assign n29264 = \P2_P2_InstQueue_reg[12][7]/NET0131  & ~n28050 ;
  assign n29275 = n26794 & n27983 ;
  assign n29276 = n28964 & n29275 ;
  assign n29277 = ~n29264 & ~n29276 ;
  assign n29278 = ~n29271 & n29277 ;
  assign n29279 = ~n29274 & n29278 ;
  assign n29283 = \P2_P2_InstQueue_reg[13][7]/NET0131  & ~n28398 ;
  assign n29288 = ~n26354 & n28398 ;
  assign n29289 = ~n29283 & ~n29288 ;
  assign n29290 = n27613 & ~n29289 ;
  assign n29282 = ~n28460 & ~n28951 ;
  assign n29284 = ~n28438 & n29283 ;
  assign n29285 = ~n29282 & ~n29284 ;
  assign n29281 = ~n27977 & n28473 ;
  assign n29286 = ~n28948 & ~n29281 ;
  assign n29287 = ~n29285 & n29286 ;
  assign n29280 = \P2_P2_InstQueue_reg[13][7]/NET0131  & ~n28050 ;
  assign n29291 = n26794 & n27980 ;
  assign n29292 = n28964 & n29291 ;
  assign n29293 = ~n29280 & ~n29292 ;
  assign n29294 = ~n29287 & n29293 ;
  assign n29295 = ~n29290 & n29294 ;
  assign n29299 = \P2_P2_InstQueue_reg[14][7]/NET0131  & ~n28401 ;
  assign n29304 = ~n26354 & n28401 ;
  assign n29305 = ~n29299 & ~n29304 ;
  assign n29306 = n27613 & ~n29305 ;
  assign n29298 = ~n28405 & ~n28951 ;
  assign n29300 = ~n28398 & n29299 ;
  assign n29301 = ~n29298 & ~n29300 ;
  assign n29297 = ~n27977 & n28493 ;
  assign n29302 = ~n28948 & ~n29297 ;
  assign n29303 = ~n29301 & n29302 ;
  assign n29296 = \P2_P2_InstQueue_reg[14][7]/NET0131  & ~n28050 ;
  assign n29307 = n26794 & n28438 ;
  assign n29308 = n28964 & n29307 ;
  assign n29309 = ~n29296 & ~n29308 ;
  assign n29310 = ~n29303 & n29309 ;
  assign n29311 = ~n29306 & n29310 ;
  assign n29315 = \P2_P2_InstQueue_reg[15][7]/NET0131  & ~n28387 ;
  assign n29320 = ~n26354 & n28387 ;
  assign n29321 = ~n29315 & ~n29320 ;
  assign n29322 = n27613 & ~n29321 ;
  assign n29314 = ~n28501 & ~n28951 ;
  assign n29316 = ~n28401 & n29315 ;
  assign n29317 = ~n29314 & ~n29316 ;
  assign n29313 = ~n27977 & n28514 ;
  assign n29318 = ~n28948 & ~n29313 ;
  assign n29319 = ~n29317 & n29318 ;
  assign n29312 = \P2_P2_InstQueue_reg[15][7]/NET0131  & ~n28050 ;
  assign n29323 = n26794 & n28398 ;
  assign n29324 = n28964 & n29323 ;
  assign n29325 = ~n29312 & ~n29324 ;
  assign n29326 = ~n29319 & n29325 ;
  assign n29327 = ~n29322 & n29326 ;
  assign n29331 = \P2_P2_InstQueue_reg[1][7]/NET0131  & ~n28522 ;
  assign n29336 = ~n26354 & n28522 ;
  assign n29337 = ~n29331 & ~n29336 ;
  assign n29338 = n27613 & ~n29337 ;
  assign n29330 = ~n28523 & ~n28951 ;
  assign n29332 = ~n28385 & n29331 ;
  assign n29333 = ~n29330 & ~n29332 ;
  assign n29329 = ~n27977 & n28536 ;
  assign n29334 = ~n28948 & ~n29329 ;
  assign n29335 = ~n29333 & n29334 ;
  assign n29328 = \P2_P2_InstQueue_reg[1][7]/NET0131  & ~n28050 ;
  assign n29339 = n26794 & n28387 ;
  assign n29340 = n28964 & n29339 ;
  assign n29341 = ~n29328 & ~n29340 ;
  assign n29342 = ~n29335 & n29341 ;
  assign n29343 = ~n29338 & n29342 ;
  assign n29347 = \P2_P2_InstQueue_reg[2][7]/NET0131  & ~n28544 ;
  assign n29352 = ~n26354 & n28544 ;
  assign n29353 = ~n29347 & ~n29352 ;
  assign n29354 = n27613 & ~n29353 ;
  assign n29346 = ~n28545 & ~n28951 ;
  assign n29348 = ~n28522 & n29347 ;
  assign n29349 = ~n29346 & ~n29348 ;
  assign n29345 = ~n27977 & n28558 ;
  assign n29350 = ~n28948 & ~n29345 ;
  assign n29351 = ~n29349 & n29350 ;
  assign n29344 = \P2_P2_InstQueue_reg[2][7]/NET0131  & ~n28050 ;
  assign n29355 = n26794 & n28385 ;
  assign n29356 = n28964 & n29355 ;
  assign n29357 = ~n29344 & ~n29356 ;
  assign n29358 = ~n29351 & n29357 ;
  assign n29359 = ~n29354 & n29358 ;
  assign n29363 = \P2_P2_InstQueue_reg[3][7]/NET0131  & ~n28566 ;
  assign n29368 = ~n26354 & n28566 ;
  assign n29369 = ~n29363 & ~n29368 ;
  assign n29370 = n27613 & ~n29369 ;
  assign n29362 = ~n28567 & ~n28951 ;
  assign n29364 = ~n28544 & n29363 ;
  assign n29365 = ~n29362 & ~n29364 ;
  assign n29361 = ~n27977 & n28580 ;
  assign n29366 = ~n28948 & ~n29361 ;
  assign n29367 = ~n29365 & n29366 ;
  assign n29360 = \P2_P2_InstQueue_reg[3][7]/NET0131  & ~n28050 ;
  assign n29371 = n26794 & n28522 ;
  assign n29372 = n28964 & n29371 ;
  assign n29373 = ~n29360 & ~n29372 ;
  assign n29374 = ~n29367 & n29373 ;
  assign n29375 = ~n29370 & n29374 ;
  assign n29379 = \P2_P2_InstQueue_reg[4][7]/NET0131  & ~n28588 ;
  assign n29384 = ~n26354 & n28588 ;
  assign n29385 = ~n29379 & ~n29384 ;
  assign n29386 = n27613 & ~n29385 ;
  assign n29378 = ~n28589 & ~n28951 ;
  assign n29380 = ~n28566 & n29379 ;
  assign n29381 = ~n29378 & ~n29380 ;
  assign n29377 = ~n27977 & n28602 ;
  assign n29382 = ~n28948 & ~n29377 ;
  assign n29383 = ~n29381 & n29382 ;
  assign n29376 = \P2_P2_InstQueue_reg[4][7]/NET0131  & ~n28050 ;
  assign n29387 = n26794 & n28544 ;
  assign n29388 = n28964 & n29387 ;
  assign n29389 = ~n29376 & ~n29388 ;
  assign n29390 = ~n29383 & n29389 ;
  assign n29391 = ~n29386 & n29390 ;
  assign n29395 = \P2_P2_InstQueue_reg[5][7]/NET0131  & ~n28610 ;
  assign n29400 = ~n26354 & n28610 ;
  assign n29401 = ~n29395 & ~n29400 ;
  assign n29402 = n27613 & ~n29401 ;
  assign n29394 = ~n28611 & ~n28951 ;
  assign n29396 = ~n28588 & n29395 ;
  assign n29397 = ~n29394 & ~n29396 ;
  assign n29393 = ~n27977 & n28624 ;
  assign n29398 = ~n28948 & ~n29393 ;
  assign n29399 = ~n29397 & n29398 ;
  assign n29392 = \P2_P2_InstQueue_reg[5][7]/NET0131  & ~n28050 ;
  assign n29403 = n26794 & n28566 ;
  assign n29404 = n28964 & n29403 ;
  assign n29405 = ~n29392 & ~n29404 ;
  assign n29406 = ~n29399 & n29405 ;
  assign n29407 = ~n29402 & n29406 ;
  assign n29411 = \P2_P2_InstQueue_reg[6][7]/NET0131  & ~n28632 ;
  assign n29416 = ~n26354 & n28632 ;
  assign n29417 = ~n29411 & ~n29416 ;
  assign n29418 = n27613 & ~n29417 ;
  assign n29410 = ~n28633 & ~n28951 ;
  assign n29412 = ~n28610 & n29411 ;
  assign n29413 = ~n29410 & ~n29412 ;
  assign n29409 = ~n27977 & n28646 ;
  assign n29414 = ~n28948 & ~n29409 ;
  assign n29415 = ~n29413 & n29414 ;
  assign n29408 = \P2_P2_InstQueue_reg[6][7]/NET0131  & ~n28050 ;
  assign n29419 = n26794 & n28588 ;
  assign n29420 = n28964 & n29419 ;
  assign n29421 = ~n29408 & ~n29420 ;
  assign n29422 = ~n29415 & n29421 ;
  assign n29423 = ~n29418 & n29422 ;
  assign n29427 = \P2_P2_InstQueue_reg[7][7]/NET0131  & ~n28423 ;
  assign n29432 = ~n26354 & n28423 ;
  assign n29433 = ~n29427 & ~n29432 ;
  assign n29434 = n27613 & ~n29433 ;
  assign n29426 = ~n28654 & ~n28951 ;
  assign n29428 = ~n28632 & n29427 ;
  assign n29429 = ~n29426 & ~n29428 ;
  assign n29425 = ~n27977 & n28667 ;
  assign n29430 = ~n28948 & ~n29425 ;
  assign n29431 = ~n29429 & n29430 ;
  assign n29424 = \P2_P2_InstQueue_reg[7][7]/NET0131  & ~n28050 ;
  assign n29435 = n26794 & n28610 ;
  assign n29436 = n28964 & n29435 ;
  assign n29437 = ~n29424 & ~n29436 ;
  assign n29438 = ~n29431 & n29437 ;
  assign n29439 = ~n29434 & n29438 ;
  assign n29443 = \P2_P2_InstQueue_reg[8][7]/NET0131  & ~n28027 ;
  assign n29448 = ~n26354 & n28027 ;
  assign n29449 = ~n29443 & ~n29448 ;
  assign n29450 = n27613 & ~n29449 ;
  assign n29442 = ~n28428 & ~n28951 ;
  assign n29444 = ~n28423 & n29443 ;
  assign n29445 = ~n29442 & ~n29444 ;
  assign n29441 = ~n27977 & n28687 ;
  assign n29446 = ~n28948 & ~n29441 ;
  assign n29447 = ~n29445 & n29446 ;
  assign n29440 = \P2_P2_InstQueue_reg[8][7]/NET0131  & ~n28050 ;
  assign n29451 = n26794 & n28632 ;
  assign n29452 = n28964 & n29451 ;
  assign n29453 = ~n29440 & ~n29452 ;
  assign n29454 = ~n29447 & n29453 ;
  assign n29455 = ~n29450 & n29454 ;
  assign n29459 = \P2_P2_InstQueue_reg[9][7]/NET0131  & ~n28034 ;
  assign n29464 = ~n26354 & n28034 ;
  assign n29465 = ~n29459 & ~n29464 ;
  assign n29466 = n27613 & ~n29465 ;
  assign n29458 = ~n28041 & ~n28951 ;
  assign n29460 = ~n28027 & n29459 ;
  assign n29461 = ~n29458 & ~n29460 ;
  assign n29457 = ~n27977 & n28707 ;
  assign n29462 = ~n28948 & ~n29457 ;
  assign n29463 = ~n29461 & n29462 ;
  assign n29456 = \P2_P2_InstQueue_reg[9][7]/NET0131  & ~n28050 ;
  assign n29467 = n26794 & n28423 ;
  assign n29468 = n28964 & n29467 ;
  assign n29469 = ~n29456 & ~n29468 ;
  assign n29470 = ~n29463 & n29469 ;
  assign n29471 = ~n29466 & n29470 ;
  assign n29472 = \P2_P1_EAX_reg[7]/NET0131  & ~n27438 ;
  assign n29505 = n11387 & n24708 ;
  assign n29478 = \P2_P1_InstQueue_reg[7][7]/NET0131  & n11651 ;
  assign n29477 = \P2_P1_InstQueue_reg[0][7]/NET0131  & n11647 ;
  assign n29473 = \P2_P1_InstQueue_reg[12][7]/NET0131  & n11665 ;
  assign n29474 = \P2_P1_InstQueue_reg[2][7]/NET0131  & n11671 ;
  assign n29489 = ~n29473 & ~n29474 ;
  assign n29499 = ~n29477 & n29489 ;
  assign n29500 = ~n29478 & n29499 ;
  assign n29485 = \P2_P1_InstQueue_reg[11][7]/NET0131  & n11634 ;
  assign n29486 = \P2_P1_InstQueue_reg[5][7]/NET0131  & n11667 ;
  assign n29494 = ~n29485 & ~n29486 ;
  assign n29487 = \P2_P1_InstQueue_reg[1][7]/NET0131  & n11669 ;
  assign n29488 = \P2_P1_InstQueue_reg[14][7]/NET0131  & n11641 ;
  assign n29495 = ~n29487 & ~n29488 ;
  assign n29496 = n29494 & n29495 ;
  assign n29481 = \P2_P1_InstQueue_reg[9][7]/NET0131  & n11659 ;
  assign n29482 = \P2_P1_InstQueue_reg[8][7]/NET0131  & n11661 ;
  assign n29492 = ~n29481 & ~n29482 ;
  assign n29483 = \P2_P1_InstQueue_reg[10][7]/NET0131  & n11656 ;
  assign n29484 = \P2_P1_InstQueue_reg[13][7]/NET0131  & n11673 ;
  assign n29493 = ~n29483 & ~n29484 ;
  assign n29497 = n29492 & n29493 ;
  assign n29475 = \P2_P1_InstQueue_reg[6][7]/NET0131  & n11638 ;
  assign n29476 = \P2_P1_InstQueue_reg[15][7]/NET0131  & n11643 ;
  assign n29490 = ~n29475 & ~n29476 ;
  assign n29479 = \P2_P1_InstQueue_reg[3][7]/NET0131  & n11654 ;
  assign n29480 = \P2_P1_InstQueue_reg[4][7]/NET0131  & n11663 ;
  assign n29491 = ~n29479 & ~n29480 ;
  assign n29498 = n29490 & n29491 ;
  assign n29501 = n29497 & n29498 ;
  assign n29502 = n29496 & n29501 ;
  assign n29503 = n29500 & n29502 ;
  assign n29504 = n20728 & ~n29503 ;
  assign n29506 = ~\P2_P1_EAX_reg[7]/NET0131  & ~n21028 ;
  assign n29507 = ~n21029 & ~n29506 ;
  assign n29508 = n21022 & n29507 ;
  assign n29509 = ~n29504 & ~n29508 ;
  assign n29510 = ~n29505 & n29509 ;
  assign n29511 = n11623 & ~n29510 ;
  assign n29512 = ~n29472 & ~n29511 ;
  assign n29513 = ~\P2_P1_EAX_reg[27]/NET0131  & ~n27398 ;
  assign n29514 = ~n27399 & ~n29513 ;
  assign n29515 = n24898 & n29514 ;
  assign n29516 = ~n27535 & ~n29515 ;
  assign n29517 = ~n21081 & ~n29516 ;
  assign n29518 = \P2_P1_uWord_reg[11]/NET0131  & ~n25154 ;
  assign n29519 = ~n29517 & ~n29518 ;
  assign n29520 = n11623 & ~n29519 ;
  assign n29521 = \P2_P1_uWord_reg[11]/NET0131  & ~n24913 ;
  assign n29522 = ~n29520 & ~n29521 ;
  assign n29523 = \P1_P1_EAX_reg[7]/NET0131  & ~n15326 ;
  assign n29525 = \P1_P1_EAX_reg[7]/NET0131  & ~n15365 ;
  assign n29526 = ~n24133 & ~n29525 ;
  assign n29527 = ~n15384 & ~n29526 ;
  assign n29524 = \P1_P1_EAX_reg[7]/NET0131  & ~n23190 ;
  assign n29528 = \P1_P1_InstQueue_reg[15][7]/NET0131  & n8291 ;
  assign n29529 = \P1_P1_InstQueue_reg[12][7]/NET0131  & n8312 ;
  assign n29530 = \P1_P1_InstQueue_reg[2][7]/NET0131  & n8299 ;
  assign n29544 = ~n29529 & ~n29530 ;
  assign n29531 = \P1_P1_InstQueue_reg[11][7]/NET0131  & n8303 ;
  assign n29532 = \P1_P1_InstQueue_reg[1][7]/NET0131  & n8309 ;
  assign n29545 = ~n29531 & ~n29532 ;
  assign n29554 = n29544 & n29545 ;
  assign n29555 = ~n29528 & n29554 ;
  assign n29543 = \P1_P1_InstQueue_reg[6][7]/NET0131  & n8307 ;
  assign n29541 = \P1_P1_InstQueue_reg[10][7]/NET0131  & n8325 ;
  assign n29542 = \P1_P1_InstQueue_reg[5][7]/NET0131  & n8295 ;
  assign n29550 = ~n29541 & ~n29542 ;
  assign n29551 = ~n29543 & n29550 ;
  assign n29537 = \P1_P1_InstQueue_reg[7][7]/NET0131  & n8316 ;
  assign n29538 = \P1_P1_InstQueue_reg[0][7]/NET0131  & n8321 ;
  assign n29548 = ~n29537 & ~n29538 ;
  assign n29539 = \P1_P1_InstQueue_reg[8][7]/NET0131  & n8318 ;
  assign n29540 = \P1_P1_InstQueue_reg[3][7]/NET0131  & n8314 ;
  assign n29549 = ~n29539 & ~n29540 ;
  assign n29552 = n29548 & n29549 ;
  assign n29533 = \P1_P1_InstQueue_reg[13][7]/NET0131  & n8329 ;
  assign n29534 = \P1_P1_InstQueue_reg[14][7]/NET0131  & n8327 ;
  assign n29546 = ~n29533 & ~n29534 ;
  assign n29535 = \P1_P1_InstQueue_reg[4][7]/NET0131  & n8323 ;
  assign n29536 = \P1_P1_InstQueue_reg[9][7]/NET0131  & n8305 ;
  assign n29547 = ~n29535 & ~n29536 ;
  assign n29553 = n29546 & n29547 ;
  assign n29556 = n29552 & n29553 ;
  assign n29557 = n29551 & n29556 ;
  assign n29558 = n29555 & n29557 ;
  assign n29559 = n22818 & ~n29558 ;
  assign n29560 = ~\P1_P1_EAX_reg[7]/NET0131  & ~n15393 ;
  assign n29561 = ~n15394 & ~n29560 ;
  assign n29562 = n15377 & n29561 ;
  assign n29563 = ~n29559 & ~n29562 ;
  assign n29564 = ~n29524 & n29563 ;
  assign n29565 = ~n29527 & n29564 ;
  assign n29566 = n8355 & ~n29565 ;
  assign n29567 = ~n29523 & ~n29566 ;
  assign n29568 = ~\P4_addr_reg[12]/NET0131  & n15734 ;
  assign n29569 = n18666 & ~n29568 ;
  assign n29571 = ~n15744 & ~n29569 ;
  assign n29579 = ~n28840 & ~n28841 ;
  assign n29581 = n28843 & n29579 ;
  assign n29580 = ~n28843 & ~n29579 ;
  assign n29582 = n15733 & ~n29580 ;
  assign n29583 = ~n29581 & n29582 ;
  assign n29573 = ~n28826 & ~n28827 ;
  assign n29575 = n28829 & n29573 ;
  assign n29574 = ~n28829 & ~n29573 ;
  assign n29576 = n27804 & ~n29574 ;
  assign n29577 = ~n29575 & n29576 ;
  assign n29572 = \P4_IR_reg[12]/NET0131  & n21786 ;
  assign n29578 = \P4_addr_reg[12]/NET0131  & n15745 ;
  assign n29584 = ~n29572 & ~n29578 ;
  assign n29585 = ~n29577 & n29584 ;
  assign n29586 = ~n29583 & n29585 ;
  assign n29587 = ~n29571 & ~n29586 ;
  assign n29570 = n15734 & n29569 ;
  assign n29588 = ~n22008 & ~n29570 ;
  assign n29589 = ~n29587 & n29588 ;
  assign n29590 = ~\P4_addr_reg[14]/NET0131  & n15734 ;
  assign n29591 = n18666 & ~n29590 ;
  assign n29593 = ~n15744 & ~n29591 ;
  assign n29605 = \P4_IR_reg[14]/NET0131  & \P4_reg2_reg[14]/NET0131  ;
  assign n29606 = ~\P4_IR_reg[14]/NET0131  & ~\P4_reg2_reg[14]/NET0131  ;
  assign n29607 = ~n29605 & ~n29606 ;
  assign n29608 = ~n28837 & ~n28845 ;
  assign n29609 = ~n28838 & ~n29608 ;
  assign n29611 = n29607 & n29609 ;
  assign n29610 = ~n29607 & ~n29609 ;
  assign n29612 = n15733 & ~n29610 ;
  assign n29613 = ~n29611 & n29612 ;
  assign n29595 = \P4_IR_reg[14]/NET0131  & \P4_reg1_reg[14]/NET0131  ;
  assign n29596 = ~\P4_IR_reg[14]/NET0131  & ~\P4_reg1_reg[14]/NET0131  ;
  assign n29597 = ~n29595 & ~n29596 ;
  assign n29598 = ~n28823 & ~n28831 ;
  assign n29599 = ~n28824 & ~n29598 ;
  assign n29601 = n29597 & n29599 ;
  assign n29600 = ~n29597 & ~n29599 ;
  assign n29602 = n27804 & ~n29600 ;
  assign n29603 = ~n29601 & n29602 ;
  assign n29594 = \P4_addr_reg[14]/NET0131  & n15745 ;
  assign n29604 = \P4_IR_reg[14]/NET0131  & n21786 ;
  assign n29614 = ~n29594 & ~n29604 ;
  assign n29615 = ~n29603 & n29614 ;
  assign n29616 = ~n29613 & n29615 ;
  assign n29617 = ~n29593 & ~n29616 ;
  assign n29592 = n15734 & n29591 ;
  assign n29618 = ~n22450 & ~n29592 ;
  assign n29619 = ~n29617 & n29618 ;
  assign n29620 = ~\P4_addr_reg[15]/NET0131  & n15734 ;
  assign n29621 = n18666 & ~n29620 ;
  assign n29623 = ~n15744 & ~n29621 ;
  assign n29635 = \P4_IR_reg[15]/NET0131  & \P4_reg2_reg[15]/NET0131  ;
  assign n29636 = ~\P4_IR_reg[15]/NET0131  & ~\P4_reg2_reg[15]/NET0131  ;
  assign n29637 = ~n29635 & ~n29636 ;
  assign n29638 = ~n29605 & ~n29609 ;
  assign n29639 = ~n29606 & ~n29638 ;
  assign n29641 = n29637 & n29639 ;
  assign n29640 = ~n29637 & ~n29639 ;
  assign n29642 = n15733 & ~n29640 ;
  assign n29643 = ~n29641 & n29642 ;
  assign n29625 = \P4_IR_reg[15]/NET0131  & \P4_reg1_reg[15]/NET0131  ;
  assign n29626 = ~\P4_IR_reg[15]/NET0131  & ~\P4_reg1_reg[15]/NET0131  ;
  assign n29627 = ~n29625 & ~n29626 ;
  assign n29628 = ~n29595 & ~n29599 ;
  assign n29629 = ~n29596 & ~n29628 ;
  assign n29631 = n29627 & n29629 ;
  assign n29630 = ~n29627 & ~n29629 ;
  assign n29632 = n27804 & ~n29630 ;
  assign n29633 = ~n29631 & n29632 ;
  assign n29624 = \P4_IR_reg[15]/NET0131  & n21786 ;
  assign n29634 = \P4_addr_reg[15]/NET0131  & n15745 ;
  assign n29644 = ~n29624 & ~n29634 ;
  assign n29645 = ~n29633 & n29644 ;
  assign n29646 = ~n29643 & n29645 ;
  assign n29647 = ~n29623 & ~n29646 ;
  assign n29622 = n15734 & n29621 ;
  assign n29648 = ~n19072 & ~n29622 ;
  assign n29649 = ~n29647 & n29648 ;
  assign n29650 = ~\P4_addr_reg[16]/NET0131  & n15734 ;
  assign n29651 = n18666 & ~n29650 ;
  assign n29653 = ~n15744 & ~n29651 ;
  assign n29665 = \P4_IR_reg[16]/NET0131  & \P4_reg1_reg[16]/NET0131  ;
  assign n29666 = ~\P4_IR_reg[16]/NET0131  & ~\P4_reg1_reg[16]/NET0131  ;
  assign n29667 = ~n29665 & ~n29666 ;
  assign n29668 = ~n29625 & ~n29629 ;
  assign n29669 = ~n29626 & ~n29668 ;
  assign n29671 = n29667 & n29669 ;
  assign n29670 = ~n29667 & ~n29669 ;
  assign n29672 = n27804 & ~n29670 ;
  assign n29673 = ~n29671 & n29672 ;
  assign n29655 = \P4_IR_reg[16]/NET0131  & \P4_reg2_reg[16]/NET0131  ;
  assign n29656 = ~\P4_IR_reg[16]/NET0131  & ~\P4_reg2_reg[16]/NET0131  ;
  assign n29657 = ~n29655 & ~n29656 ;
  assign n29658 = ~n29635 & ~n29639 ;
  assign n29659 = ~n29636 & ~n29658 ;
  assign n29661 = n29657 & n29659 ;
  assign n29660 = ~n29657 & ~n29659 ;
  assign n29662 = n15733 & ~n29660 ;
  assign n29663 = ~n29661 & n29662 ;
  assign n29654 = \P4_addr_reg[16]/NET0131  & n15745 ;
  assign n29664 = \P4_IR_reg[16]/NET0131  & n21786 ;
  assign n29674 = ~n29654 & ~n29664 ;
  assign n29675 = ~n29663 & n29674 ;
  assign n29676 = ~n29673 & n29675 ;
  assign n29677 = ~n29653 & ~n29676 ;
  assign n29652 = n15734 & n29651 ;
  assign n29678 = ~n22040 & ~n29652 ;
  assign n29679 = ~n29677 & n29678 ;
  assign n29680 = ~\P4_addr_reg[17]/NET0131  & n15734 ;
  assign n29681 = n18666 & ~n29680 ;
  assign n29683 = ~n15744 & ~n29681 ;
  assign n29695 = \P4_IR_reg[17]/NET0131  & \P4_reg2_reg[17]/NET0131  ;
  assign n29696 = ~\P4_IR_reg[17]/NET0131  & ~\P4_reg2_reg[17]/NET0131  ;
  assign n29697 = ~n29695 & ~n29696 ;
  assign n29698 = ~n29655 & ~n29659 ;
  assign n29699 = ~n29656 & ~n29698 ;
  assign n29701 = n29697 & n29699 ;
  assign n29700 = ~n29697 & ~n29699 ;
  assign n29702 = n15733 & ~n29700 ;
  assign n29703 = ~n29701 & n29702 ;
  assign n29685 = \P4_IR_reg[17]/NET0131  & \P4_reg1_reg[17]/NET0131  ;
  assign n29686 = ~\P4_IR_reg[17]/NET0131  & ~\P4_reg1_reg[17]/NET0131  ;
  assign n29687 = ~n29685 & ~n29686 ;
  assign n29688 = ~n29665 & ~n29669 ;
  assign n29689 = ~n29666 & ~n29688 ;
  assign n29691 = n29687 & n29689 ;
  assign n29690 = ~n29687 & ~n29689 ;
  assign n29692 = n27804 & ~n29690 ;
  assign n29693 = ~n29691 & n29692 ;
  assign n29684 = \P4_IR_reg[17]/NET0131  & n21786 ;
  assign n29694 = \P4_addr_reg[17]/NET0131  & n15745 ;
  assign n29704 = ~n29684 & ~n29694 ;
  assign n29705 = ~n29693 & n29704 ;
  assign n29706 = ~n29703 & n29705 ;
  assign n29707 = ~n29683 & ~n29706 ;
  assign n29682 = n15734 & n29681 ;
  assign n29708 = ~n23267 & ~n29682 ;
  assign n29709 = ~n29707 & n29708 ;
  assign n29710 = ~\P4_addr_reg[18]/NET0131  & n15734 ;
  assign n29711 = n18666 & ~n29710 ;
  assign n29713 = ~n15744 & ~n29711 ;
  assign n29715 = ~n29695 & ~n29699 ;
  assign n29716 = ~n29696 & ~n29715 ;
  assign n29717 = \P4_IR_reg[18]/NET0131  & n29716 ;
  assign n29718 = ~\P4_IR_reg[18]/NET0131  & ~n29716 ;
  assign n29719 = ~n29717 & ~n29718 ;
  assign n29721 = ~\P4_reg2_reg[18]/NET0131  & ~n29719 ;
  assign n29720 = \P4_reg2_reg[18]/NET0131  & n29719 ;
  assign n29722 = n15733 & ~n29720 ;
  assign n29723 = ~n29721 & n29722 ;
  assign n29725 = ~\P4_IR_reg[18]/NET0131  & ~\P4_reg1_reg[18]/NET0131  ;
  assign n29726 = \P4_IR_reg[18]/NET0131  & \P4_reg1_reg[18]/NET0131  ;
  assign n29727 = ~n29725 & ~n29726 ;
  assign n29728 = ~n29685 & ~n29689 ;
  assign n29729 = ~n29686 & ~n29728 ;
  assign n29731 = n29727 & n29729 ;
  assign n29730 = ~n29727 & ~n29729 ;
  assign n29732 = n27804 & ~n29730 ;
  assign n29733 = ~n29731 & n29732 ;
  assign n29714 = \P4_addr_reg[18]/NET0131  & n15745 ;
  assign n29724 = \P4_IR_reg[18]/NET0131  & n21786 ;
  assign n29734 = ~n29714 & ~n29724 ;
  assign n29735 = ~n29733 & n29734 ;
  assign n29736 = ~n29723 & n29735 ;
  assign n29737 = ~n29713 & ~n29736 ;
  assign n29712 = n15734 & n29711 ;
  assign n29738 = ~n23059 & ~n29712 ;
  assign n29739 = ~n29737 & n29738 ;
  assign n29741 = \P3_rd_reg/NET0131  & ~n27815 ;
  assign n29749 = ~n27820 & ~n27821 ;
  assign n29751 = n27802 & n29749 ;
  assign n29750 = ~n27802 & ~n29749 ;
  assign n29752 = n27804 & ~n29750 ;
  assign n29753 = ~n29751 & n29752 ;
  assign n29743 = ~n27832 & ~n27833 ;
  assign n29745 = n27799 & n29743 ;
  assign n29744 = ~n27799 & ~n29743 ;
  assign n29746 = n15733 & ~n29744 ;
  assign n29747 = ~n29745 & n29746 ;
  assign n29742 = \P4_addr_reg[1]/NET0131  & n15745 ;
  assign n29748 = \P4_IR_reg[1]/NET0131  & n21786 ;
  assign n29754 = ~n29742 & ~n29748 ;
  assign n29755 = ~n29747 & n29754 ;
  assign n29756 = ~n29753 & n29755 ;
  assign n29757 = n29741 & ~n29756 ;
  assign n29740 = ~\P3_rd_reg/NET0131  & \P4_reg3_reg[1]/NET0131  ;
  assign n29758 = \P4_addr_reg[1]/NET0131  & n18665 ;
  assign n29759 = n15737 & n29758 ;
  assign n29760 = ~n29740 & ~n29759 ;
  assign n29761 = ~n29757 & n29760 ;
  assign n29769 = ~n27870 & ~n27871 ;
  assign n29771 = n27873 & n29769 ;
  assign n29770 = ~n27873 & ~n29769 ;
  assign n29772 = n27804 & ~n29770 ;
  assign n29773 = ~n29771 & n29772 ;
  assign n29764 = ~n27857 & ~n27858 ;
  assign n29766 = n27860 & n29764 ;
  assign n29765 = ~n27860 & ~n29764 ;
  assign n29767 = n15733 & ~n29765 ;
  assign n29768 = ~n29766 & n29767 ;
  assign n29762 = \P4_addr_reg[3]/NET0131  & n15745 ;
  assign n29763 = \P4_IR_reg[3]/NET0131  & n21786 ;
  assign n29774 = ~n29762 & ~n29763 ;
  assign n29775 = ~n29768 & n29774 ;
  assign n29776 = ~n29773 & n29775 ;
  assign n29779 = ~n15734 & n29776 ;
  assign n29778 = ~\P4_addr_reg[3]/NET0131  & n15734 ;
  assign n29780 = n18666 & ~n29778 ;
  assign n29781 = ~n29779 & n29780 ;
  assign n29777 = n15744 & ~n29776 ;
  assign n29782 = ~n22906 & ~n29777 ;
  assign n29783 = ~n29781 & n29782 ;
  assign n29784 = ~\P4_addr_reg[6]/NET0131  & n15734 ;
  assign n29785 = n18666 & ~n29784 ;
  assign n29787 = ~n15744 & ~n29785 ;
  assign n29795 = ~n28790 & ~n28791 ;
  assign n29797 = n28797 & n29795 ;
  assign n29796 = ~n28797 & ~n29795 ;
  assign n29798 = n27804 & ~n29796 ;
  assign n29799 = ~n29797 & n29798 ;
  assign n29789 = ~n28756 & ~n28757 ;
  assign n29791 = n28763 & n29789 ;
  assign n29790 = ~n28763 & ~n29789 ;
  assign n29792 = n15733 & ~n29790 ;
  assign n29793 = ~n29791 & n29792 ;
  assign n29788 = \P4_addr_reg[6]/NET0131  & n15745 ;
  assign n29794 = \P4_IR_reg[6]/NET0131  & n21786 ;
  assign n29800 = ~n29788 & ~n29794 ;
  assign n29801 = ~n29793 & n29800 ;
  assign n29802 = ~n29799 & n29801 ;
  assign n29803 = ~n29787 & ~n29802 ;
  assign n29786 = n15734 & n29785 ;
  assign n29804 = ~n22949 & ~n29786 ;
  assign n29805 = ~n29803 & n29804 ;
  assign n29806 = ~\P4_addr_reg[7]/NET0131  & n15734 ;
  assign n29807 = n18666 & ~n29806 ;
  assign n29809 = ~n15744 & ~n29807 ;
  assign n29817 = ~n28788 & ~n28789 ;
  assign n29819 = n28799 & n29817 ;
  assign n29818 = ~n28799 & ~n29817 ;
  assign n29820 = n27804 & ~n29818 ;
  assign n29821 = ~n29819 & n29820 ;
  assign n29811 = ~n28754 & ~n28755 ;
  assign n29813 = n28765 & n29811 ;
  assign n29812 = ~n28765 & ~n29811 ;
  assign n29814 = n15733 & ~n29812 ;
  assign n29815 = ~n29813 & n29814 ;
  assign n29810 = \P4_addr_reg[7]/NET0131  & n15745 ;
  assign n29816 = \P4_IR_reg[7]/NET0131  & n21786 ;
  assign n29822 = ~n29810 & ~n29816 ;
  assign n29823 = ~n29815 & n29822 ;
  assign n29824 = ~n29821 & n29823 ;
  assign n29825 = ~n29809 & ~n29824 ;
  assign n29808 = n15734 & n29807 ;
  assign n29826 = ~n22073 & ~n29808 ;
  assign n29827 = ~n29825 & n29826 ;
  assign n29828 = ~n15745 & ~n27815 ;
  assign n29829 = \P3_rd_reg/NET0131  & ~n29828 ;
  assign n29838 = \P1_buf2_reg[27]/NET0131  & ~n27934 ;
  assign n29839 = \P1_buf1_reg[27]/NET0131  & n27934 ;
  assign n29840 = ~n29838 & ~n29839 ;
  assign n29841 = n27945 & ~n29840 ;
  assign n29842 = \P1_buf2_reg[19]/NET0131  & ~n27934 ;
  assign n29843 = \P1_buf1_reg[19]/NET0131  & n27934 ;
  assign n29844 = ~n29842 & ~n29843 ;
  assign n29845 = n27952 & ~n29844 ;
  assign n29846 = ~n29841 & ~n29845 ;
  assign n29847 = \P1_P2_DataWidth_reg[1]/NET0131  & ~n29846 ;
  assign n29830 = \P1_buf2_reg[3]/NET0131  & ~n27934 ;
  assign n29831 = \P1_buf1_reg[3]/NET0131  & n27934 ;
  assign n29832 = ~n29830 & ~n29831 ;
  assign n29833 = ~n27905 & ~n29832 ;
  assign n29834 = \P1_P2_InstQueue_reg[11][3]/NET0131  & ~n27901 ;
  assign n29835 = ~n27904 & n29834 ;
  assign n29836 = ~n29833 & ~n29835 ;
  assign n29848 = ~n27960 & ~n29836 ;
  assign n29849 = ~n29847 & ~n29848 ;
  assign n29850 = n25928 & ~n29849 ;
  assign n29851 = ~n25699 & n27901 ;
  assign n29852 = ~n29834 & ~n29851 ;
  assign n29853 = n27608 & ~n29852 ;
  assign n29837 = n27898 & ~n29836 ;
  assign n29854 = \P1_P2_InstQueue_reg[11][3]/NET0131  & ~n27972 ;
  assign n29855 = ~n29837 & ~n29854 ;
  assign n29856 = ~n29853 & n29855 ;
  assign n29857 = ~n29850 & n29856 ;
  assign n29866 = \P1_buf2_reg[29]/NET0131  & ~n27934 ;
  assign n29867 = \P1_buf1_reg[29]/NET0131  & n27934 ;
  assign n29868 = ~n29866 & ~n29867 ;
  assign n29869 = n27945 & ~n29868 ;
  assign n29870 = \P1_buf2_reg[21]/NET0131  & ~n27934 ;
  assign n29871 = \P1_buf1_reg[21]/NET0131  & n27934 ;
  assign n29872 = ~n29870 & ~n29871 ;
  assign n29873 = n27952 & ~n29872 ;
  assign n29874 = ~n29869 & ~n29873 ;
  assign n29875 = \P1_P2_DataWidth_reg[1]/NET0131  & ~n29874 ;
  assign n29858 = \P1_buf2_reg[5]/NET0131  & ~n27934 ;
  assign n29859 = \P1_buf1_reg[5]/NET0131  & n27934 ;
  assign n29860 = ~n29858 & ~n29859 ;
  assign n29861 = ~n27905 & ~n29860 ;
  assign n29862 = \P1_P2_InstQueue_reg[11][5]/NET0131  & ~n27901 ;
  assign n29863 = ~n27904 & n29862 ;
  assign n29864 = ~n29861 & ~n29863 ;
  assign n29876 = ~n27960 & ~n29864 ;
  assign n29877 = ~n29875 & ~n29876 ;
  assign n29878 = n25928 & ~n29877 ;
  assign n29879 = ~n25477 & n27901 ;
  assign n29880 = ~n29862 & ~n29879 ;
  assign n29881 = n27608 & ~n29880 ;
  assign n29865 = n27898 & ~n29864 ;
  assign n29882 = \P1_P2_InstQueue_reg[11][5]/NET0131  & ~n27972 ;
  assign n29883 = ~n29865 & ~n29882 ;
  assign n29884 = ~n29881 & n29883 ;
  assign n29885 = ~n29878 & n29884 ;
  assign n29897 = \P2_buf2_reg[27]/NET0131  & ~n28013 ;
  assign n29898 = \P2_buf1_reg[27]/NET0131  & n28013 ;
  assign n29899 = ~n29897 & ~n29898 ;
  assign n29900 = n28027 & ~n29899 ;
  assign n29901 = \P2_buf2_reg[19]/NET0131  & ~n28013 ;
  assign n29902 = \P2_buf1_reg[19]/NET0131  & n28013 ;
  assign n29903 = ~n29901 & ~n29902 ;
  assign n29904 = n28034 & ~n29903 ;
  assign n29905 = ~n29900 & ~n29904 ;
  assign n29906 = \P2_P2_DataWidth_reg[1]/NET0131  & ~n29905 ;
  assign n29886 = \P2_buf2_reg[3]/NET0131  & ~n28013 ;
  assign n29887 = \P2_buf1_reg[3]/NET0131  & n28013 ;
  assign n29888 = ~n29886 & ~n29887 ;
  assign n29889 = ~n27984 & ~n29888 ;
  assign n29890 = \P2_P2_InstQueue_reg[11][3]/NET0131  & ~n27980 ;
  assign n29891 = ~n27983 & n29890 ;
  assign n29892 = ~n29889 & ~n29891 ;
  assign n29907 = ~n28042 & ~n29892 ;
  assign n29908 = ~n29906 & ~n29907 ;
  assign n29909 = n26794 & ~n29908 ;
  assign n29894 = ~n26576 & n27980 ;
  assign n29895 = ~n29890 & ~n29894 ;
  assign n29896 = n27613 & ~n29895 ;
  assign n29893 = n27977 & ~n29892 ;
  assign n29910 = \P2_P2_InstQueue_reg[11][3]/NET0131  & ~n28050 ;
  assign n29911 = ~n29893 & ~n29910 ;
  assign n29912 = ~n29896 & n29911 ;
  assign n29913 = ~n29909 & n29912 ;
  assign n29915 = \P4_addr_reg[0]/NET0131  & n15745 ;
  assign n29916 = ~n27808 & ~n29915 ;
  assign n29917 = n27807 & n29916 ;
  assign n29918 = n29741 & ~n29917 ;
  assign n29914 = ~\P3_rd_reg/NET0131  & \P4_reg3_reg[0]/NET0131  ;
  assign n29919 = \P4_addr_reg[0]/NET0131  & n18665 ;
  assign n29920 = n15737 & n29919 ;
  assign n29921 = ~n29914 & ~n29920 ;
  assign n29922 = ~n29918 & n29921 ;
  assign n29928 = n28065 & ~n29840 ;
  assign n29929 = n28068 & ~n29844 ;
  assign n29930 = ~n29928 & ~n29929 ;
  assign n29931 = \P1_P2_DataWidth_reg[1]/NET0131  & ~n29930 ;
  assign n29923 = ~n28058 & ~n29832 ;
  assign n29924 = \P1_P2_InstQueue_reg[0][3]/NET0131  & ~n28055 ;
  assign n29925 = ~n28057 & n29924 ;
  assign n29926 = ~n29923 & ~n29925 ;
  assign n29932 = ~n28073 & ~n29926 ;
  assign n29933 = ~n29931 & ~n29932 ;
  assign n29934 = n25928 & ~n29933 ;
  assign n29935 = ~n25699 & n28055 ;
  assign n29936 = ~n29924 & ~n29935 ;
  assign n29937 = n27608 & ~n29936 ;
  assign n29927 = n27898 & ~n29926 ;
  assign n29938 = \P1_P2_InstQueue_reg[0][3]/NET0131  & ~n27972 ;
  assign n29939 = ~n29927 & ~n29938 ;
  assign n29940 = ~n29937 & n29939 ;
  assign n29941 = ~n29934 & n29940 ;
  assign n29947 = n28065 & ~n29868 ;
  assign n29948 = n28068 & ~n29872 ;
  assign n29949 = ~n29947 & ~n29948 ;
  assign n29950 = \P1_P2_DataWidth_reg[1]/NET0131  & ~n29949 ;
  assign n29942 = ~n28058 & ~n29860 ;
  assign n29943 = \P1_P2_InstQueue_reg[0][5]/NET0131  & ~n28055 ;
  assign n29944 = ~n28057 & n29943 ;
  assign n29945 = ~n29942 & ~n29944 ;
  assign n29951 = ~n28073 & ~n29945 ;
  assign n29952 = ~n29950 & ~n29951 ;
  assign n29953 = n25928 & ~n29952 ;
  assign n29954 = ~n25477 & n28055 ;
  assign n29955 = ~n29943 & ~n29954 ;
  assign n29956 = n27608 & ~n29955 ;
  assign n29946 = n27898 & ~n29945 ;
  assign n29957 = \P1_P2_InstQueue_reg[0][5]/NET0131  & ~n27972 ;
  assign n29958 = ~n29946 & ~n29957 ;
  assign n29959 = ~n29956 & n29958 ;
  assign n29960 = ~n29953 & n29959 ;
  assign n29966 = n28090 & ~n29840 ;
  assign n29967 = n27945 & ~n29844 ;
  assign n29968 = ~n29966 & ~n29967 ;
  assign n29969 = \P1_P2_DataWidth_reg[1]/NET0131  & ~n29968 ;
  assign n29961 = ~n28084 & ~n29832 ;
  assign n29962 = \P1_P2_InstQueue_reg[10][3]/NET0131  & ~n27904 ;
  assign n29963 = ~n27952 & n29962 ;
  assign n29964 = ~n29961 & ~n29963 ;
  assign n29970 = ~n28096 & ~n29964 ;
  assign n29971 = ~n29969 & ~n29970 ;
  assign n29972 = n25928 & ~n29971 ;
  assign n29973 = ~n25699 & n27904 ;
  assign n29974 = ~n29962 & ~n29973 ;
  assign n29975 = n27608 & ~n29974 ;
  assign n29965 = n27898 & ~n29964 ;
  assign n29976 = \P1_P2_InstQueue_reg[10][3]/NET0131  & ~n27972 ;
  assign n29977 = ~n29965 & ~n29976 ;
  assign n29978 = ~n29975 & n29977 ;
  assign n29979 = ~n29972 & n29978 ;
  assign n29985 = n28090 & ~n29868 ;
  assign n29986 = n27945 & ~n29872 ;
  assign n29987 = ~n29985 & ~n29986 ;
  assign n29988 = \P1_P2_DataWidth_reg[1]/NET0131  & ~n29987 ;
  assign n29980 = ~n28084 & ~n29860 ;
  assign n29981 = \P1_P2_InstQueue_reg[10][5]/NET0131  & ~n27904 ;
  assign n29982 = ~n27952 & n29981 ;
  assign n29983 = ~n29980 & ~n29982 ;
  assign n29989 = ~n28096 & ~n29983 ;
  assign n29990 = ~n29988 & ~n29989 ;
  assign n29991 = n25928 & ~n29990 ;
  assign n29992 = ~n25477 & n27904 ;
  assign n29993 = ~n29981 & ~n29992 ;
  assign n29994 = n27608 & ~n29993 ;
  assign n29984 = n27898 & ~n29983 ;
  assign n29995 = \P1_P2_InstQueue_reg[10][5]/NET0131  & ~n27972 ;
  assign n29996 = ~n29984 & ~n29995 ;
  assign n29997 = ~n29994 & n29996 ;
  assign n29998 = ~n29991 & n29997 ;
  assign n30004 = n27952 & ~n29840 ;
  assign n30005 = n27904 & ~n29844 ;
  assign n30006 = ~n30004 & ~n30005 ;
  assign n30007 = \P1_P2_DataWidth_reg[1]/NET0131  & ~n30006 ;
  assign n29999 = ~n28109 & ~n29832 ;
  assign n30000 = \P1_P2_InstQueue_reg[12][3]/NET0131  & ~n28108 ;
  assign n30001 = ~n27901 & n30000 ;
  assign n30002 = ~n29999 & ~n30001 ;
  assign n30008 = ~n28119 & ~n30002 ;
  assign n30009 = ~n30007 & ~n30008 ;
  assign n30010 = n25928 & ~n30009 ;
  assign n30011 = ~n25699 & n28108 ;
  assign n30012 = ~n30000 & ~n30011 ;
  assign n30013 = n27608 & ~n30012 ;
  assign n30003 = n27898 & ~n30002 ;
  assign n30014 = \P1_P2_InstQueue_reg[12][3]/NET0131  & ~n27972 ;
  assign n30015 = ~n30003 & ~n30014 ;
  assign n30016 = ~n30013 & n30015 ;
  assign n30017 = ~n30010 & n30016 ;
  assign n30023 = n27952 & ~n29868 ;
  assign n30024 = n27904 & ~n29872 ;
  assign n30025 = ~n30023 & ~n30024 ;
  assign n30026 = \P1_P2_DataWidth_reg[1]/NET0131  & ~n30025 ;
  assign n30018 = ~n28109 & ~n29860 ;
  assign n30019 = \P1_P2_InstQueue_reg[12][5]/NET0131  & ~n28108 ;
  assign n30020 = ~n27901 & n30019 ;
  assign n30021 = ~n30018 & ~n30020 ;
  assign n30027 = ~n28119 & ~n30021 ;
  assign n30028 = ~n30026 & ~n30027 ;
  assign n30029 = n25928 & ~n30028 ;
  assign n30030 = ~n25477 & n28108 ;
  assign n30031 = ~n30019 & ~n30030 ;
  assign n30032 = n27608 & ~n30031 ;
  assign n30022 = n27898 & ~n30021 ;
  assign n30033 = \P1_P2_InstQueue_reg[12][5]/NET0131  & ~n27972 ;
  assign n30034 = ~n30022 & ~n30033 ;
  assign n30035 = ~n30032 & n30034 ;
  assign n30036 = ~n30029 & n30035 ;
  assign n30042 = n27904 & ~n29840 ;
  assign n30043 = n27901 & ~n29844 ;
  assign n30044 = ~n30042 & ~n30043 ;
  assign n30045 = \P1_P2_DataWidth_reg[1]/NET0131  & ~n30044 ;
  assign n30037 = ~n28130 & ~n29832 ;
  assign n30038 = \P1_P2_InstQueue_reg[13][3]/NET0131  & ~n28065 ;
  assign n30039 = ~n28108 & n30038 ;
  assign n30040 = ~n30037 & ~n30039 ;
  assign n30046 = ~n28140 & ~n30040 ;
  assign n30047 = ~n30045 & ~n30046 ;
  assign n30048 = n25928 & ~n30047 ;
  assign n30049 = ~n25699 & n28065 ;
  assign n30050 = ~n30038 & ~n30049 ;
  assign n30051 = n27608 & ~n30050 ;
  assign n30041 = n27898 & ~n30040 ;
  assign n30052 = \P1_P2_InstQueue_reg[13][3]/NET0131  & ~n27972 ;
  assign n30053 = ~n30041 & ~n30052 ;
  assign n30054 = ~n30051 & n30053 ;
  assign n30055 = ~n30048 & n30054 ;
  assign n30061 = n27904 & ~n29868 ;
  assign n30062 = n27901 & ~n29872 ;
  assign n30063 = ~n30061 & ~n30062 ;
  assign n30064 = \P1_P2_DataWidth_reg[1]/NET0131  & ~n30063 ;
  assign n30056 = ~n28130 & ~n29860 ;
  assign n30057 = \P1_P2_InstQueue_reg[13][5]/NET0131  & ~n28065 ;
  assign n30058 = ~n28108 & n30057 ;
  assign n30059 = ~n30056 & ~n30058 ;
  assign n30065 = ~n28140 & ~n30059 ;
  assign n30066 = ~n30064 & ~n30065 ;
  assign n30067 = n25928 & ~n30066 ;
  assign n30068 = ~n25477 & n28065 ;
  assign n30069 = ~n30057 & ~n30068 ;
  assign n30070 = n27608 & ~n30069 ;
  assign n30060 = n27898 & ~n30059 ;
  assign n30071 = \P1_P2_InstQueue_reg[13][5]/NET0131  & ~n27972 ;
  assign n30072 = ~n30060 & ~n30071 ;
  assign n30073 = ~n30070 & n30072 ;
  assign n30074 = ~n30067 & n30073 ;
  assign n30080 = n27901 & ~n29840 ;
  assign n30081 = n28108 & ~n29844 ;
  assign n30082 = ~n30080 & ~n30081 ;
  assign n30083 = \P1_P2_DataWidth_reg[1]/NET0131  & ~n30082 ;
  assign n30075 = ~n28072 & ~n29832 ;
  assign n30076 = \P1_P2_InstQueue_reg[14][3]/NET0131  & ~n28068 ;
  assign n30077 = ~n28065 & n30076 ;
  assign n30078 = ~n30075 & ~n30077 ;
  assign n30084 = ~n28160 & ~n30078 ;
  assign n30085 = ~n30083 & ~n30084 ;
  assign n30086 = n25928 & ~n30085 ;
  assign n30087 = ~n25699 & n28068 ;
  assign n30088 = ~n30076 & ~n30087 ;
  assign n30089 = n27608 & ~n30088 ;
  assign n30079 = n27898 & ~n30078 ;
  assign n30090 = \P1_P2_InstQueue_reg[14][3]/NET0131  & ~n27972 ;
  assign n30091 = ~n30079 & ~n30090 ;
  assign n30092 = ~n30089 & n30091 ;
  assign n30093 = ~n30086 & n30092 ;
  assign n30099 = n27901 & ~n29868 ;
  assign n30100 = n28108 & ~n29872 ;
  assign n30101 = ~n30099 & ~n30100 ;
  assign n30102 = \P1_P2_DataWidth_reg[1]/NET0131  & ~n30101 ;
  assign n30094 = ~n28072 & ~n29860 ;
  assign n30095 = \P1_P2_InstQueue_reg[14][5]/NET0131  & ~n28068 ;
  assign n30096 = ~n28065 & n30095 ;
  assign n30097 = ~n30094 & ~n30096 ;
  assign n30103 = ~n28160 & ~n30097 ;
  assign n30104 = ~n30102 & ~n30103 ;
  assign n30105 = n25928 & ~n30104 ;
  assign n30106 = ~n25477 & n28068 ;
  assign n30107 = ~n30095 & ~n30106 ;
  assign n30108 = n27608 & ~n30107 ;
  assign n30098 = n27898 & ~n30097 ;
  assign n30109 = \P1_P2_InstQueue_reg[14][5]/NET0131  & ~n27972 ;
  assign n30110 = ~n30098 & ~n30109 ;
  assign n30111 = ~n30108 & n30110 ;
  assign n30112 = ~n30105 & n30111 ;
  assign n30118 = n28108 & ~n29840 ;
  assign n30119 = n28065 & ~n29844 ;
  assign n30120 = ~n30118 & ~n30119 ;
  assign n30121 = \P1_P2_DataWidth_reg[1]/NET0131  & ~n30120 ;
  assign n30113 = ~n28171 & ~n29832 ;
  assign n30114 = \P1_P2_InstQueue_reg[15][3]/NET0131  & ~n28057 ;
  assign n30115 = ~n28068 & n30114 ;
  assign n30116 = ~n30113 & ~n30115 ;
  assign n30122 = ~n28181 & ~n30116 ;
  assign n30123 = ~n30121 & ~n30122 ;
  assign n30124 = n25928 & ~n30123 ;
  assign n30125 = ~n25699 & n28057 ;
  assign n30126 = ~n30114 & ~n30125 ;
  assign n30127 = n27608 & ~n30126 ;
  assign n30117 = n27898 & ~n30116 ;
  assign n30128 = \P1_P2_InstQueue_reg[15][3]/NET0131  & ~n27972 ;
  assign n30129 = ~n30117 & ~n30128 ;
  assign n30130 = ~n30127 & n30129 ;
  assign n30131 = ~n30124 & n30130 ;
  assign n30137 = n28108 & ~n29868 ;
  assign n30138 = n28065 & ~n29872 ;
  assign n30139 = ~n30137 & ~n30138 ;
  assign n30140 = \P1_P2_DataWidth_reg[1]/NET0131  & ~n30139 ;
  assign n30132 = ~n28171 & ~n29860 ;
  assign n30133 = \P1_P2_InstQueue_reg[15][5]/NET0131  & ~n28057 ;
  assign n30134 = ~n28068 & n30133 ;
  assign n30135 = ~n30132 & ~n30134 ;
  assign n30141 = ~n28181 & ~n30135 ;
  assign n30142 = ~n30140 & ~n30141 ;
  assign n30143 = n25928 & ~n30142 ;
  assign n30144 = ~n25477 & n28057 ;
  assign n30145 = ~n30133 & ~n30144 ;
  assign n30146 = n27608 & ~n30145 ;
  assign n30136 = n27898 & ~n30135 ;
  assign n30147 = \P1_P2_InstQueue_reg[15][5]/NET0131  & ~n27972 ;
  assign n30148 = ~n30136 & ~n30147 ;
  assign n30149 = ~n30146 & n30148 ;
  assign n30150 = ~n30143 & n30149 ;
  assign n30156 = n28068 & ~n29840 ;
  assign n30157 = n28057 & ~n29844 ;
  assign n30158 = ~n30156 & ~n30157 ;
  assign n30159 = \P1_P2_DataWidth_reg[1]/NET0131  & ~n30158 ;
  assign n30151 = ~n28193 & ~n29832 ;
  assign n30152 = \P1_P2_InstQueue_reg[1][3]/NET0131  & ~n28192 ;
  assign n30153 = ~n28055 & n30152 ;
  assign n30154 = ~n30151 & ~n30153 ;
  assign n30160 = ~n28203 & ~n30154 ;
  assign n30161 = ~n30159 & ~n30160 ;
  assign n30162 = n25928 & ~n30161 ;
  assign n30163 = ~n25699 & n28192 ;
  assign n30164 = ~n30152 & ~n30163 ;
  assign n30165 = n27608 & ~n30164 ;
  assign n30155 = n27898 & ~n30154 ;
  assign n30166 = \P1_P2_InstQueue_reg[1][3]/NET0131  & ~n27972 ;
  assign n30167 = ~n30155 & ~n30166 ;
  assign n30168 = ~n30165 & n30167 ;
  assign n30169 = ~n30162 & n30168 ;
  assign n30175 = n28068 & ~n29868 ;
  assign n30176 = n28057 & ~n29872 ;
  assign n30177 = ~n30175 & ~n30176 ;
  assign n30178 = \P1_P2_DataWidth_reg[1]/NET0131  & ~n30177 ;
  assign n30170 = ~n28193 & ~n29860 ;
  assign n30171 = \P1_P2_InstQueue_reg[1][5]/NET0131  & ~n28192 ;
  assign n30172 = ~n28055 & n30171 ;
  assign n30173 = ~n30170 & ~n30172 ;
  assign n30179 = ~n28203 & ~n30173 ;
  assign n30180 = ~n30178 & ~n30179 ;
  assign n30181 = n25928 & ~n30180 ;
  assign n30182 = ~n25477 & n28192 ;
  assign n30183 = ~n30171 & ~n30182 ;
  assign n30184 = n27608 & ~n30183 ;
  assign n30174 = n27898 & ~n30173 ;
  assign n30185 = \P1_P2_InstQueue_reg[1][5]/NET0131  & ~n27972 ;
  assign n30186 = ~n30174 & ~n30185 ;
  assign n30187 = ~n30184 & n30186 ;
  assign n30188 = ~n30181 & n30187 ;
  assign n30194 = n28057 & ~n29840 ;
  assign n30195 = n28055 & ~n29844 ;
  assign n30196 = ~n30194 & ~n30195 ;
  assign n30197 = \P1_P2_DataWidth_reg[1]/NET0131  & ~n30196 ;
  assign n30189 = ~n28215 & ~n29832 ;
  assign n30190 = \P1_P2_InstQueue_reg[2][3]/NET0131  & ~n28214 ;
  assign n30191 = ~n28192 & n30190 ;
  assign n30192 = ~n30189 & ~n30191 ;
  assign n30198 = ~n28225 & ~n30192 ;
  assign n30199 = ~n30197 & ~n30198 ;
  assign n30200 = n25928 & ~n30199 ;
  assign n30201 = ~n25699 & n28214 ;
  assign n30202 = ~n30190 & ~n30201 ;
  assign n30203 = n27608 & ~n30202 ;
  assign n30193 = n27898 & ~n30192 ;
  assign n30204 = \P1_P2_InstQueue_reg[2][3]/NET0131  & ~n27972 ;
  assign n30205 = ~n30193 & ~n30204 ;
  assign n30206 = ~n30203 & n30205 ;
  assign n30207 = ~n30200 & n30206 ;
  assign n30213 = n28057 & ~n29868 ;
  assign n30214 = n28055 & ~n29872 ;
  assign n30215 = ~n30213 & ~n30214 ;
  assign n30216 = \P1_P2_DataWidth_reg[1]/NET0131  & ~n30215 ;
  assign n30208 = ~n28215 & ~n29860 ;
  assign n30209 = \P1_P2_InstQueue_reg[2][5]/NET0131  & ~n28214 ;
  assign n30210 = ~n28192 & n30209 ;
  assign n30211 = ~n30208 & ~n30210 ;
  assign n30217 = ~n28225 & ~n30211 ;
  assign n30218 = ~n30216 & ~n30217 ;
  assign n30219 = n25928 & ~n30218 ;
  assign n30220 = ~n25477 & n28214 ;
  assign n30221 = ~n30209 & ~n30220 ;
  assign n30222 = n27608 & ~n30221 ;
  assign n30212 = n27898 & ~n30211 ;
  assign n30223 = \P1_P2_InstQueue_reg[2][5]/NET0131  & ~n27972 ;
  assign n30224 = ~n30212 & ~n30223 ;
  assign n30225 = ~n30222 & n30224 ;
  assign n30226 = ~n30219 & n30225 ;
  assign n30232 = n28055 & ~n29840 ;
  assign n30233 = n28192 & ~n29844 ;
  assign n30234 = ~n30232 & ~n30233 ;
  assign n30235 = \P1_P2_DataWidth_reg[1]/NET0131  & ~n30234 ;
  assign n30227 = ~n28237 & ~n29832 ;
  assign n30228 = \P1_P2_InstQueue_reg[3][3]/NET0131  & ~n28236 ;
  assign n30229 = ~n28214 & n30228 ;
  assign n30230 = ~n30227 & ~n30229 ;
  assign n30236 = ~n28247 & ~n30230 ;
  assign n30237 = ~n30235 & ~n30236 ;
  assign n30238 = n25928 & ~n30237 ;
  assign n30239 = ~n25699 & n28236 ;
  assign n30240 = ~n30228 & ~n30239 ;
  assign n30241 = n27608 & ~n30240 ;
  assign n30231 = n27898 & ~n30230 ;
  assign n30242 = \P1_P2_InstQueue_reg[3][3]/NET0131  & ~n27972 ;
  assign n30243 = ~n30231 & ~n30242 ;
  assign n30244 = ~n30241 & n30243 ;
  assign n30245 = ~n30238 & n30244 ;
  assign n30251 = n28055 & ~n29868 ;
  assign n30252 = n28192 & ~n29872 ;
  assign n30253 = ~n30251 & ~n30252 ;
  assign n30254 = \P1_P2_DataWidth_reg[1]/NET0131  & ~n30253 ;
  assign n30246 = ~n28237 & ~n29860 ;
  assign n30247 = \P1_P2_InstQueue_reg[3][5]/NET0131  & ~n28236 ;
  assign n30248 = ~n28214 & n30247 ;
  assign n30249 = ~n30246 & ~n30248 ;
  assign n30255 = ~n28247 & ~n30249 ;
  assign n30256 = ~n30254 & ~n30255 ;
  assign n30257 = n25928 & ~n30256 ;
  assign n30258 = ~n25477 & n28236 ;
  assign n30259 = ~n30247 & ~n30258 ;
  assign n30260 = n27608 & ~n30259 ;
  assign n30250 = n27898 & ~n30249 ;
  assign n30261 = \P1_P2_InstQueue_reg[3][5]/NET0131  & ~n27972 ;
  assign n30262 = ~n30250 & ~n30261 ;
  assign n30263 = ~n30260 & n30262 ;
  assign n30264 = ~n30257 & n30263 ;
  assign n30270 = n28192 & ~n29840 ;
  assign n30271 = n28214 & ~n29844 ;
  assign n30272 = ~n30270 & ~n30271 ;
  assign n30273 = \P1_P2_DataWidth_reg[1]/NET0131  & ~n30272 ;
  assign n30265 = ~n28259 & ~n29832 ;
  assign n30266 = \P1_P2_InstQueue_reg[4][3]/NET0131  & ~n28258 ;
  assign n30267 = ~n28236 & n30266 ;
  assign n30268 = ~n30265 & ~n30267 ;
  assign n30274 = ~n28269 & ~n30268 ;
  assign n30275 = ~n30273 & ~n30274 ;
  assign n30276 = n25928 & ~n30275 ;
  assign n30277 = ~n25699 & n28258 ;
  assign n30278 = ~n30266 & ~n30277 ;
  assign n30279 = n27608 & ~n30278 ;
  assign n30269 = n27898 & ~n30268 ;
  assign n30280 = \P1_P2_InstQueue_reg[4][3]/NET0131  & ~n27972 ;
  assign n30281 = ~n30269 & ~n30280 ;
  assign n30282 = ~n30279 & n30281 ;
  assign n30283 = ~n30276 & n30282 ;
  assign n30289 = n28192 & ~n29868 ;
  assign n30290 = n28214 & ~n29872 ;
  assign n30291 = ~n30289 & ~n30290 ;
  assign n30292 = \P1_P2_DataWidth_reg[1]/NET0131  & ~n30291 ;
  assign n30284 = ~n28259 & ~n29860 ;
  assign n30285 = \P1_P2_InstQueue_reg[4][5]/NET0131  & ~n28258 ;
  assign n30286 = ~n28236 & n30285 ;
  assign n30287 = ~n30284 & ~n30286 ;
  assign n30293 = ~n28269 & ~n30287 ;
  assign n30294 = ~n30292 & ~n30293 ;
  assign n30295 = n25928 & ~n30294 ;
  assign n30296 = ~n25477 & n28258 ;
  assign n30297 = ~n30285 & ~n30296 ;
  assign n30298 = n27608 & ~n30297 ;
  assign n30288 = n27898 & ~n30287 ;
  assign n30299 = \P1_P2_InstQueue_reg[4][5]/NET0131  & ~n27972 ;
  assign n30300 = ~n30288 & ~n30299 ;
  assign n30301 = ~n30298 & n30300 ;
  assign n30302 = ~n30295 & n30301 ;
  assign n30308 = n28214 & ~n29840 ;
  assign n30309 = n28236 & ~n29844 ;
  assign n30310 = ~n30308 & ~n30309 ;
  assign n30311 = \P1_P2_DataWidth_reg[1]/NET0131  & ~n30310 ;
  assign n30303 = ~n28281 & ~n29832 ;
  assign n30304 = \P1_P2_InstQueue_reg[5][3]/NET0131  & ~n28280 ;
  assign n30305 = ~n28258 & n30304 ;
  assign n30306 = ~n30303 & ~n30305 ;
  assign n30312 = ~n28291 & ~n30306 ;
  assign n30313 = ~n30311 & ~n30312 ;
  assign n30314 = n25928 & ~n30313 ;
  assign n30315 = ~n25699 & n28280 ;
  assign n30316 = ~n30304 & ~n30315 ;
  assign n30317 = n27608 & ~n30316 ;
  assign n30307 = n27898 & ~n30306 ;
  assign n30318 = \P1_P2_InstQueue_reg[5][3]/NET0131  & ~n27972 ;
  assign n30319 = ~n30307 & ~n30318 ;
  assign n30320 = ~n30317 & n30319 ;
  assign n30321 = ~n30314 & n30320 ;
  assign n30327 = n28214 & ~n29868 ;
  assign n30328 = n28236 & ~n29872 ;
  assign n30329 = ~n30327 & ~n30328 ;
  assign n30330 = \P1_P2_DataWidth_reg[1]/NET0131  & ~n30329 ;
  assign n30322 = ~n28281 & ~n29860 ;
  assign n30323 = \P1_P2_InstQueue_reg[5][5]/NET0131  & ~n28280 ;
  assign n30324 = ~n28258 & n30323 ;
  assign n30325 = ~n30322 & ~n30324 ;
  assign n30331 = ~n28291 & ~n30325 ;
  assign n30332 = ~n30330 & ~n30331 ;
  assign n30333 = n25928 & ~n30332 ;
  assign n30334 = ~n25477 & n28280 ;
  assign n30335 = ~n30323 & ~n30334 ;
  assign n30336 = n27608 & ~n30335 ;
  assign n30326 = n27898 & ~n30325 ;
  assign n30337 = \P1_P2_InstQueue_reg[5][5]/NET0131  & ~n27972 ;
  assign n30338 = ~n30326 & ~n30337 ;
  assign n30339 = ~n30336 & n30338 ;
  assign n30340 = ~n30333 & n30339 ;
  assign n30346 = n28236 & ~n29840 ;
  assign n30347 = n28258 & ~n29844 ;
  assign n30348 = ~n30346 & ~n30347 ;
  assign n30349 = \P1_P2_DataWidth_reg[1]/NET0131  & ~n30348 ;
  assign n30341 = ~n28303 & ~n29832 ;
  assign n30342 = \P1_P2_InstQueue_reg[6][3]/NET0131  & ~n28302 ;
  assign n30343 = ~n28280 & n30342 ;
  assign n30344 = ~n30341 & ~n30343 ;
  assign n30350 = ~n28313 & ~n30344 ;
  assign n30351 = ~n30349 & ~n30350 ;
  assign n30352 = n25928 & ~n30351 ;
  assign n30353 = ~n25699 & n28302 ;
  assign n30354 = ~n30342 & ~n30353 ;
  assign n30355 = n27608 & ~n30354 ;
  assign n30345 = n27898 & ~n30344 ;
  assign n30356 = \P1_P2_InstQueue_reg[6][3]/NET0131  & ~n27972 ;
  assign n30357 = ~n30345 & ~n30356 ;
  assign n30358 = ~n30355 & n30357 ;
  assign n30359 = ~n30352 & n30358 ;
  assign n30365 = n28236 & ~n29868 ;
  assign n30366 = n28258 & ~n29872 ;
  assign n30367 = ~n30365 & ~n30366 ;
  assign n30368 = \P1_P2_DataWidth_reg[1]/NET0131  & ~n30367 ;
  assign n30360 = ~n28303 & ~n29860 ;
  assign n30361 = \P1_P2_InstQueue_reg[6][5]/NET0131  & ~n28302 ;
  assign n30362 = ~n28280 & n30361 ;
  assign n30363 = ~n30360 & ~n30362 ;
  assign n30369 = ~n28313 & ~n30363 ;
  assign n30370 = ~n30368 & ~n30369 ;
  assign n30371 = n25928 & ~n30370 ;
  assign n30372 = ~n25477 & n28302 ;
  assign n30373 = ~n30361 & ~n30372 ;
  assign n30374 = n27608 & ~n30373 ;
  assign n30364 = n27898 & ~n30363 ;
  assign n30375 = \P1_P2_InstQueue_reg[6][5]/NET0131  & ~n27972 ;
  assign n30376 = ~n30364 & ~n30375 ;
  assign n30377 = ~n30374 & n30376 ;
  assign n30378 = ~n30371 & n30377 ;
  assign n30384 = n28258 & ~n29840 ;
  assign n30385 = n28280 & ~n29844 ;
  assign n30386 = ~n30384 & ~n30385 ;
  assign n30387 = \P1_P2_DataWidth_reg[1]/NET0131  & ~n30386 ;
  assign n30379 = ~n28324 & ~n29832 ;
  assign n30380 = \P1_P2_InstQueue_reg[7][3]/NET0131  & ~n28090 ;
  assign n30381 = ~n28302 & n30380 ;
  assign n30382 = ~n30379 & ~n30381 ;
  assign n30388 = ~n28334 & ~n30382 ;
  assign n30389 = ~n30387 & ~n30388 ;
  assign n30390 = n25928 & ~n30389 ;
  assign n30391 = ~n25699 & n28090 ;
  assign n30392 = ~n30380 & ~n30391 ;
  assign n30393 = n27608 & ~n30392 ;
  assign n30383 = n27898 & ~n30382 ;
  assign n30394 = \P1_P2_InstQueue_reg[7][3]/NET0131  & ~n27972 ;
  assign n30395 = ~n30383 & ~n30394 ;
  assign n30396 = ~n30393 & n30395 ;
  assign n30397 = ~n30390 & n30396 ;
  assign n30403 = n28258 & ~n29868 ;
  assign n30404 = n28280 & ~n29872 ;
  assign n30405 = ~n30403 & ~n30404 ;
  assign n30406 = \P1_P2_DataWidth_reg[1]/NET0131  & ~n30405 ;
  assign n30398 = ~n28324 & ~n29860 ;
  assign n30399 = \P1_P2_InstQueue_reg[7][5]/NET0131  & ~n28090 ;
  assign n30400 = ~n28302 & n30399 ;
  assign n30401 = ~n30398 & ~n30400 ;
  assign n30407 = ~n28334 & ~n30401 ;
  assign n30408 = ~n30406 & ~n30407 ;
  assign n30409 = n25928 & ~n30408 ;
  assign n30410 = ~n25477 & n28090 ;
  assign n30411 = ~n30399 & ~n30410 ;
  assign n30412 = n27608 & ~n30411 ;
  assign n30402 = n27898 & ~n30401 ;
  assign n30413 = \P1_P2_InstQueue_reg[7][5]/NET0131  & ~n27972 ;
  assign n30414 = ~n30402 & ~n30413 ;
  assign n30415 = ~n30412 & n30414 ;
  assign n30416 = ~n30409 & n30415 ;
  assign n30422 = n28280 & ~n29840 ;
  assign n30423 = n28302 & ~n29844 ;
  assign n30424 = ~n30422 & ~n30423 ;
  assign n30425 = \P1_P2_DataWidth_reg[1]/NET0131  & ~n30424 ;
  assign n30417 = ~n28095 & ~n29832 ;
  assign n30418 = \P1_P2_InstQueue_reg[8][3]/NET0131  & ~n27945 ;
  assign n30419 = ~n28090 & n30418 ;
  assign n30420 = ~n30417 & ~n30419 ;
  assign n30426 = ~n28354 & ~n30420 ;
  assign n30427 = ~n30425 & ~n30426 ;
  assign n30428 = n25928 & ~n30427 ;
  assign n30429 = ~n25699 & n27945 ;
  assign n30430 = ~n30418 & ~n30429 ;
  assign n30431 = n27608 & ~n30430 ;
  assign n30421 = n27898 & ~n30420 ;
  assign n30432 = \P1_P2_InstQueue_reg[8][3]/NET0131  & ~n27972 ;
  assign n30433 = ~n30421 & ~n30432 ;
  assign n30434 = ~n30431 & n30433 ;
  assign n30435 = ~n30428 & n30434 ;
  assign n30441 = n28280 & ~n29868 ;
  assign n30442 = n28302 & ~n29872 ;
  assign n30443 = ~n30441 & ~n30442 ;
  assign n30444 = \P1_P2_DataWidth_reg[1]/NET0131  & ~n30443 ;
  assign n30436 = ~n28095 & ~n29860 ;
  assign n30437 = \P1_P2_InstQueue_reg[8][5]/NET0131  & ~n27945 ;
  assign n30438 = ~n28090 & n30437 ;
  assign n30439 = ~n30436 & ~n30438 ;
  assign n30445 = ~n28354 & ~n30439 ;
  assign n30446 = ~n30444 & ~n30445 ;
  assign n30447 = n25928 & ~n30446 ;
  assign n30448 = ~n25477 & n27945 ;
  assign n30449 = ~n30437 & ~n30448 ;
  assign n30450 = n27608 & ~n30449 ;
  assign n30440 = n27898 & ~n30439 ;
  assign n30451 = \P1_P2_InstQueue_reg[8][5]/NET0131  & ~n27972 ;
  assign n30452 = ~n30440 & ~n30451 ;
  assign n30453 = ~n30450 & n30452 ;
  assign n30454 = ~n30447 & n30453 ;
  assign n30460 = n28302 & ~n29840 ;
  assign n30461 = n28090 & ~n29844 ;
  assign n30462 = ~n30460 & ~n30461 ;
  assign n30463 = \P1_P2_DataWidth_reg[1]/NET0131  & ~n30462 ;
  assign n30455 = ~n27959 & ~n29832 ;
  assign n30456 = \P1_P2_InstQueue_reg[9][3]/NET0131  & ~n27952 ;
  assign n30457 = ~n27945 & n30456 ;
  assign n30458 = ~n30455 & ~n30457 ;
  assign n30464 = ~n28374 & ~n30458 ;
  assign n30465 = ~n30463 & ~n30464 ;
  assign n30466 = n25928 & ~n30465 ;
  assign n30467 = ~n25699 & n27952 ;
  assign n30468 = ~n30456 & ~n30467 ;
  assign n30469 = n27608 & ~n30468 ;
  assign n30459 = n27898 & ~n30458 ;
  assign n30470 = \P1_P2_InstQueue_reg[9][3]/NET0131  & ~n27972 ;
  assign n30471 = ~n30459 & ~n30470 ;
  assign n30472 = ~n30469 & n30471 ;
  assign n30473 = ~n30466 & n30472 ;
  assign n30479 = n28302 & ~n29868 ;
  assign n30480 = n28090 & ~n29872 ;
  assign n30481 = ~n30479 & ~n30480 ;
  assign n30482 = \P1_P2_DataWidth_reg[1]/NET0131  & ~n30481 ;
  assign n30474 = ~n27959 & ~n29860 ;
  assign n30475 = \P1_P2_InstQueue_reg[9][5]/NET0131  & ~n27952 ;
  assign n30476 = ~n27945 & n30475 ;
  assign n30477 = ~n30474 & ~n30476 ;
  assign n30483 = ~n28374 & ~n30477 ;
  assign n30484 = ~n30482 & ~n30483 ;
  assign n30485 = n25928 & ~n30484 ;
  assign n30486 = ~n25477 & n27952 ;
  assign n30487 = ~n30475 & ~n30486 ;
  assign n30488 = n27608 & ~n30487 ;
  assign n30478 = n27898 & ~n30477 ;
  assign n30489 = \P1_P2_InstQueue_reg[9][5]/NET0131  & ~n27972 ;
  assign n30490 = ~n30478 & ~n30489 ;
  assign n30491 = ~n30488 & n30490 ;
  assign n30492 = ~n30485 & n30491 ;
  assign n30501 = n28398 & ~n29899 ;
  assign n30502 = n28401 & ~n29903 ;
  assign n30503 = ~n30501 & ~n30502 ;
  assign n30504 = \P2_P2_DataWidth_reg[1]/NET0131  & ~n30503 ;
  assign n30493 = ~n28388 & ~n29888 ;
  assign n30494 = \P2_P2_InstQueue_reg[0][3]/NET0131  & ~n28385 ;
  assign n30495 = ~n28387 & n30494 ;
  assign n30496 = ~n30493 & ~n30495 ;
  assign n30505 = ~n28406 & ~n30496 ;
  assign n30506 = ~n30504 & ~n30505 ;
  assign n30507 = n26794 & ~n30506 ;
  assign n30498 = ~n26576 & n28385 ;
  assign n30499 = ~n30494 & ~n30498 ;
  assign n30500 = n27613 & ~n30499 ;
  assign n30497 = n27977 & ~n30496 ;
  assign n30508 = \P2_P2_InstQueue_reg[0][3]/NET0131  & ~n28050 ;
  assign n30509 = ~n30497 & ~n30508 ;
  assign n30510 = ~n30500 & n30509 ;
  assign n30511 = ~n30507 & n30510 ;
  assign n30520 = n28423 & ~n29899 ;
  assign n30521 = n28027 & ~n29903 ;
  assign n30522 = ~n30520 & ~n30521 ;
  assign n30523 = \P2_P2_DataWidth_reg[1]/NET0131  & ~n30522 ;
  assign n30512 = ~n28414 & ~n29888 ;
  assign n30513 = \P2_P2_InstQueue_reg[10][3]/NET0131  & ~n27983 ;
  assign n30514 = ~n28034 & n30513 ;
  assign n30515 = ~n30512 & ~n30514 ;
  assign n30524 = ~n28429 & ~n30515 ;
  assign n30525 = ~n30523 & ~n30524 ;
  assign n30526 = n26794 & ~n30525 ;
  assign n30517 = ~n26576 & n27983 ;
  assign n30518 = ~n30513 & ~n30517 ;
  assign n30519 = n27613 & ~n30518 ;
  assign n30516 = n27977 & ~n30515 ;
  assign n30527 = \P2_P2_InstQueue_reg[10][3]/NET0131  & ~n28050 ;
  assign n30528 = ~n30516 & ~n30527 ;
  assign n30529 = ~n30519 & n30528 ;
  assign n30530 = ~n30526 & n30529 ;
  assign n30539 = n28034 & ~n29899 ;
  assign n30540 = n27983 & ~n29903 ;
  assign n30541 = ~n30539 & ~n30540 ;
  assign n30542 = \P2_P2_DataWidth_reg[1]/NET0131  & ~n30541 ;
  assign n30531 = ~n28439 & ~n29888 ;
  assign n30532 = \P2_P2_InstQueue_reg[12][3]/NET0131  & ~n28438 ;
  assign n30533 = ~n27980 & n30532 ;
  assign n30534 = ~n30531 & ~n30533 ;
  assign n30543 = ~n28452 & ~n30534 ;
  assign n30544 = ~n30542 & ~n30543 ;
  assign n30545 = n26794 & ~n30544 ;
  assign n30536 = ~n26576 & n28438 ;
  assign n30537 = ~n30532 & ~n30536 ;
  assign n30538 = n27613 & ~n30537 ;
  assign n30535 = n27977 & ~n30534 ;
  assign n30546 = \P2_P2_InstQueue_reg[12][3]/NET0131  & ~n28050 ;
  assign n30547 = ~n30535 & ~n30546 ;
  assign n30548 = ~n30538 & n30547 ;
  assign n30549 = ~n30545 & n30548 ;
  assign n30558 = n27983 & ~n29899 ;
  assign n30559 = n27980 & ~n29903 ;
  assign n30560 = ~n30558 & ~n30559 ;
  assign n30561 = \P2_P2_DataWidth_reg[1]/NET0131  & ~n30560 ;
  assign n30550 = ~n28460 & ~n29888 ;
  assign n30551 = \P2_P2_InstQueue_reg[13][3]/NET0131  & ~n28398 ;
  assign n30552 = ~n28438 & n30551 ;
  assign n30553 = ~n30550 & ~n30552 ;
  assign n30562 = ~n28473 & ~n30553 ;
  assign n30563 = ~n30561 & ~n30562 ;
  assign n30564 = n26794 & ~n30563 ;
  assign n30555 = ~n26576 & n28398 ;
  assign n30556 = ~n30551 & ~n30555 ;
  assign n30557 = n27613 & ~n30556 ;
  assign n30554 = n27977 & ~n30553 ;
  assign n30565 = \P2_P2_InstQueue_reg[13][3]/NET0131  & ~n28050 ;
  assign n30566 = ~n30554 & ~n30565 ;
  assign n30567 = ~n30557 & n30566 ;
  assign n30568 = ~n30564 & n30567 ;
  assign n30577 = n27980 & ~n29899 ;
  assign n30578 = n28438 & ~n29903 ;
  assign n30579 = ~n30577 & ~n30578 ;
  assign n30580 = \P2_P2_DataWidth_reg[1]/NET0131  & ~n30579 ;
  assign n30569 = ~n28405 & ~n29888 ;
  assign n30570 = \P2_P2_InstQueue_reg[14][3]/NET0131  & ~n28401 ;
  assign n30571 = ~n28398 & n30570 ;
  assign n30572 = ~n30569 & ~n30571 ;
  assign n30581 = ~n28493 & ~n30572 ;
  assign n30582 = ~n30580 & ~n30581 ;
  assign n30583 = n26794 & ~n30582 ;
  assign n30574 = ~n26576 & n28401 ;
  assign n30575 = ~n30570 & ~n30574 ;
  assign n30576 = n27613 & ~n30575 ;
  assign n30573 = n27977 & ~n30572 ;
  assign n30584 = \P2_P2_InstQueue_reg[14][3]/NET0131  & ~n28050 ;
  assign n30585 = ~n30573 & ~n30584 ;
  assign n30586 = ~n30576 & n30585 ;
  assign n30587 = ~n30583 & n30586 ;
  assign n30596 = n28438 & ~n29899 ;
  assign n30597 = n28398 & ~n29903 ;
  assign n30598 = ~n30596 & ~n30597 ;
  assign n30599 = \P2_P2_DataWidth_reg[1]/NET0131  & ~n30598 ;
  assign n30588 = ~n28501 & ~n29888 ;
  assign n30589 = \P2_P2_InstQueue_reg[15][3]/NET0131  & ~n28387 ;
  assign n30590 = ~n28401 & n30589 ;
  assign n30591 = ~n30588 & ~n30590 ;
  assign n30600 = ~n28514 & ~n30591 ;
  assign n30601 = ~n30599 & ~n30600 ;
  assign n30602 = n26794 & ~n30601 ;
  assign n30593 = ~n26576 & n28387 ;
  assign n30594 = ~n30589 & ~n30593 ;
  assign n30595 = n27613 & ~n30594 ;
  assign n30592 = n27977 & ~n30591 ;
  assign n30603 = \P2_P2_InstQueue_reg[15][3]/NET0131  & ~n28050 ;
  assign n30604 = ~n30592 & ~n30603 ;
  assign n30605 = ~n30595 & n30604 ;
  assign n30606 = ~n30602 & n30605 ;
  assign n30615 = n28401 & ~n29899 ;
  assign n30616 = n28387 & ~n29903 ;
  assign n30617 = ~n30615 & ~n30616 ;
  assign n30618 = \P2_P2_DataWidth_reg[1]/NET0131  & ~n30617 ;
  assign n30607 = ~n28523 & ~n29888 ;
  assign n30608 = \P2_P2_InstQueue_reg[1][3]/NET0131  & ~n28522 ;
  assign n30609 = ~n28385 & n30608 ;
  assign n30610 = ~n30607 & ~n30609 ;
  assign n30619 = ~n28536 & ~n30610 ;
  assign n30620 = ~n30618 & ~n30619 ;
  assign n30621 = n26794 & ~n30620 ;
  assign n30612 = ~n26576 & n28522 ;
  assign n30613 = ~n30608 & ~n30612 ;
  assign n30614 = n27613 & ~n30613 ;
  assign n30611 = n27977 & ~n30610 ;
  assign n30622 = \P2_P2_InstQueue_reg[1][3]/NET0131  & ~n28050 ;
  assign n30623 = ~n30611 & ~n30622 ;
  assign n30624 = ~n30614 & n30623 ;
  assign n30625 = ~n30621 & n30624 ;
  assign n30634 = n28387 & ~n29899 ;
  assign n30635 = n28385 & ~n29903 ;
  assign n30636 = ~n30634 & ~n30635 ;
  assign n30637 = \P2_P2_DataWidth_reg[1]/NET0131  & ~n30636 ;
  assign n30626 = ~n28545 & ~n29888 ;
  assign n30627 = \P2_P2_InstQueue_reg[2][3]/NET0131  & ~n28544 ;
  assign n30628 = ~n28522 & n30627 ;
  assign n30629 = ~n30626 & ~n30628 ;
  assign n30638 = ~n28558 & ~n30629 ;
  assign n30639 = ~n30637 & ~n30638 ;
  assign n30640 = n26794 & ~n30639 ;
  assign n30631 = ~n26576 & n28544 ;
  assign n30632 = ~n30627 & ~n30631 ;
  assign n30633 = n27613 & ~n30632 ;
  assign n30630 = n27977 & ~n30629 ;
  assign n30641 = \P2_P2_InstQueue_reg[2][3]/NET0131  & ~n28050 ;
  assign n30642 = ~n30630 & ~n30641 ;
  assign n30643 = ~n30633 & n30642 ;
  assign n30644 = ~n30640 & n30643 ;
  assign n30653 = n28385 & ~n29899 ;
  assign n30654 = n28522 & ~n29903 ;
  assign n30655 = ~n30653 & ~n30654 ;
  assign n30656 = \P2_P2_DataWidth_reg[1]/NET0131  & ~n30655 ;
  assign n30645 = ~n28567 & ~n29888 ;
  assign n30646 = \P2_P2_InstQueue_reg[3][3]/NET0131  & ~n28566 ;
  assign n30647 = ~n28544 & n30646 ;
  assign n30648 = ~n30645 & ~n30647 ;
  assign n30657 = ~n28580 & ~n30648 ;
  assign n30658 = ~n30656 & ~n30657 ;
  assign n30659 = n26794 & ~n30658 ;
  assign n30650 = ~n26576 & n28566 ;
  assign n30651 = ~n30646 & ~n30650 ;
  assign n30652 = n27613 & ~n30651 ;
  assign n30649 = n27977 & ~n30648 ;
  assign n30660 = \P2_P2_InstQueue_reg[3][3]/NET0131  & ~n28050 ;
  assign n30661 = ~n30649 & ~n30660 ;
  assign n30662 = ~n30652 & n30661 ;
  assign n30663 = ~n30659 & n30662 ;
  assign n30672 = n28522 & ~n29899 ;
  assign n30673 = n28544 & ~n29903 ;
  assign n30674 = ~n30672 & ~n30673 ;
  assign n30675 = \P2_P2_DataWidth_reg[1]/NET0131  & ~n30674 ;
  assign n30664 = ~n28589 & ~n29888 ;
  assign n30665 = \P2_P2_InstQueue_reg[4][3]/NET0131  & ~n28588 ;
  assign n30666 = ~n28566 & n30665 ;
  assign n30667 = ~n30664 & ~n30666 ;
  assign n30676 = ~n28602 & ~n30667 ;
  assign n30677 = ~n30675 & ~n30676 ;
  assign n30678 = n26794 & ~n30677 ;
  assign n30669 = ~n26576 & n28588 ;
  assign n30670 = ~n30665 & ~n30669 ;
  assign n30671 = n27613 & ~n30670 ;
  assign n30668 = n27977 & ~n30667 ;
  assign n30679 = \P2_P2_InstQueue_reg[4][3]/NET0131  & ~n28050 ;
  assign n30680 = ~n30668 & ~n30679 ;
  assign n30681 = ~n30671 & n30680 ;
  assign n30682 = ~n30678 & n30681 ;
  assign n30691 = n28544 & ~n29899 ;
  assign n30692 = n28566 & ~n29903 ;
  assign n30693 = ~n30691 & ~n30692 ;
  assign n30694 = \P2_P2_DataWidth_reg[1]/NET0131  & ~n30693 ;
  assign n30683 = ~n28611 & ~n29888 ;
  assign n30684 = \P2_P2_InstQueue_reg[5][3]/NET0131  & ~n28610 ;
  assign n30685 = ~n28588 & n30684 ;
  assign n30686 = ~n30683 & ~n30685 ;
  assign n30695 = ~n28624 & ~n30686 ;
  assign n30696 = ~n30694 & ~n30695 ;
  assign n30697 = n26794 & ~n30696 ;
  assign n30688 = ~n26576 & n28610 ;
  assign n30689 = ~n30684 & ~n30688 ;
  assign n30690 = n27613 & ~n30689 ;
  assign n30687 = n27977 & ~n30686 ;
  assign n30698 = \P2_P2_InstQueue_reg[5][3]/NET0131  & ~n28050 ;
  assign n30699 = ~n30687 & ~n30698 ;
  assign n30700 = ~n30690 & n30699 ;
  assign n30701 = ~n30697 & n30700 ;
  assign n30710 = n28566 & ~n29899 ;
  assign n30711 = n28588 & ~n29903 ;
  assign n30712 = ~n30710 & ~n30711 ;
  assign n30713 = \P2_P2_DataWidth_reg[1]/NET0131  & ~n30712 ;
  assign n30702 = ~n28633 & ~n29888 ;
  assign n30703 = \P2_P2_InstQueue_reg[6][3]/NET0131  & ~n28632 ;
  assign n30704 = ~n28610 & n30703 ;
  assign n30705 = ~n30702 & ~n30704 ;
  assign n30714 = ~n28646 & ~n30705 ;
  assign n30715 = ~n30713 & ~n30714 ;
  assign n30716 = n26794 & ~n30715 ;
  assign n30707 = ~n26576 & n28632 ;
  assign n30708 = ~n30703 & ~n30707 ;
  assign n30709 = n27613 & ~n30708 ;
  assign n30706 = n27977 & ~n30705 ;
  assign n30717 = \P2_P2_InstQueue_reg[6][3]/NET0131  & ~n28050 ;
  assign n30718 = ~n30706 & ~n30717 ;
  assign n30719 = ~n30709 & n30718 ;
  assign n30720 = ~n30716 & n30719 ;
  assign n30729 = n28588 & ~n29899 ;
  assign n30730 = n28610 & ~n29903 ;
  assign n30731 = ~n30729 & ~n30730 ;
  assign n30732 = \P2_P2_DataWidth_reg[1]/NET0131  & ~n30731 ;
  assign n30721 = ~n28654 & ~n29888 ;
  assign n30722 = \P2_P2_InstQueue_reg[7][3]/NET0131  & ~n28423 ;
  assign n30723 = ~n28632 & n30722 ;
  assign n30724 = ~n30721 & ~n30723 ;
  assign n30733 = ~n28667 & ~n30724 ;
  assign n30734 = ~n30732 & ~n30733 ;
  assign n30735 = n26794 & ~n30734 ;
  assign n30726 = ~n26576 & n28423 ;
  assign n30727 = ~n30722 & ~n30726 ;
  assign n30728 = n27613 & ~n30727 ;
  assign n30725 = n27977 & ~n30724 ;
  assign n30736 = \P2_P2_InstQueue_reg[7][3]/NET0131  & ~n28050 ;
  assign n30737 = ~n30725 & ~n30736 ;
  assign n30738 = ~n30728 & n30737 ;
  assign n30739 = ~n30735 & n30738 ;
  assign n30748 = n28610 & ~n29899 ;
  assign n30749 = n28632 & ~n29903 ;
  assign n30750 = ~n30748 & ~n30749 ;
  assign n30751 = \P2_P2_DataWidth_reg[1]/NET0131  & ~n30750 ;
  assign n30740 = ~n28428 & ~n29888 ;
  assign n30741 = \P2_P2_InstQueue_reg[8][3]/NET0131  & ~n28027 ;
  assign n30742 = ~n28423 & n30741 ;
  assign n30743 = ~n30740 & ~n30742 ;
  assign n30752 = ~n28687 & ~n30743 ;
  assign n30753 = ~n30751 & ~n30752 ;
  assign n30754 = n26794 & ~n30753 ;
  assign n30745 = ~n26576 & n28027 ;
  assign n30746 = ~n30741 & ~n30745 ;
  assign n30747 = n27613 & ~n30746 ;
  assign n30744 = n27977 & ~n30743 ;
  assign n30755 = \P2_P2_InstQueue_reg[8][3]/NET0131  & ~n28050 ;
  assign n30756 = ~n30744 & ~n30755 ;
  assign n30757 = ~n30747 & n30756 ;
  assign n30758 = ~n30754 & n30757 ;
  assign n30767 = n28632 & ~n29899 ;
  assign n30768 = n28423 & ~n29903 ;
  assign n30769 = ~n30767 & ~n30768 ;
  assign n30770 = \P2_P2_DataWidth_reg[1]/NET0131  & ~n30769 ;
  assign n30759 = ~n28041 & ~n29888 ;
  assign n30760 = \P2_P2_InstQueue_reg[9][3]/NET0131  & ~n28034 ;
  assign n30761 = ~n28027 & n30760 ;
  assign n30762 = ~n30759 & ~n30761 ;
  assign n30771 = ~n28707 & ~n30762 ;
  assign n30772 = ~n30770 & ~n30771 ;
  assign n30773 = n26794 & ~n30772 ;
  assign n30764 = ~n26576 & n28034 ;
  assign n30765 = ~n30760 & ~n30764 ;
  assign n30766 = n27613 & ~n30765 ;
  assign n30763 = n27977 & ~n30762 ;
  assign n30774 = \P2_P2_InstQueue_reg[9][3]/NET0131  & ~n28050 ;
  assign n30775 = ~n30763 & ~n30774 ;
  assign n30776 = ~n30766 & n30775 ;
  assign n30777 = ~n30773 & n30776 ;
  assign n30778 = \P1_P2_InstAddrPointer_reg[31]/NET0131  & n25733 ;
  assign n30810 = \P1_P2_InstAddrPointer_reg[27]/NET0131  & \P1_P2_InstAddrPointer_reg[28]/NET0131  ;
  assign n31170 = \P1_P2_InstAddrPointer_reg[29]/NET0131  & n30810 ;
  assign n30811 = \P1_P2_InstAddrPointer_reg[1]/NET0131  & \P1_P2_InstAddrPointer_reg[2]/NET0131  ;
  assign n30812 = \P1_P2_InstAddrPointer_reg[3]/NET0131  & n30811 ;
  assign n30813 = \P1_P2_InstAddrPointer_reg[4]/NET0131  & n30812 ;
  assign n30814 = \P1_P2_InstAddrPointer_reg[5]/NET0131  & n30813 ;
  assign n30815 = \P1_P2_InstAddrPointer_reg[6]/NET0131  & n30814 ;
  assign n30816 = \P1_P2_InstAddrPointer_reg[7]/NET0131  & n30815 ;
  assign n30817 = \P1_P2_InstAddrPointer_reg[22]/NET0131  & \P1_P2_InstAddrPointer_reg[23]/NET0131  ;
  assign n30818 = \P1_P2_InstAddrPointer_reg[18]/NET0131  & \P1_P2_InstAddrPointer_reg[19]/NET0131  ;
  assign n30819 = \P1_P2_InstAddrPointer_reg[17]/NET0131  & n30818 ;
  assign n30820 = \P1_P2_InstAddrPointer_reg[20]/NET0131  & n30819 ;
  assign n30821 = \P1_P2_InstAddrPointer_reg[15]/NET0131  & \P1_P2_InstAddrPointer_reg[16]/NET0131  ;
  assign n30822 = \P1_P2_InstAddrPointer_reg[21]/NET0131  & n30821 ;
  assign n30823 = n30820 & n30822 ;
  assign n30824 = n30817 & n30823 ;
  assign n30825 = \P1_P2_InstAddrPointer_reg[12]/NET0131  & \P1_P2_InstAddrPointer_reg[13]/NET0131  ;
  assign n30826 = \P1_P2_InstAddrPointer_reg[14]/NET0131  & n30825 ;
  assign n30827 = \P1_P2_InstAddrPointer_reg[10]/NET0131  & \P1_P2_InstAddrPointer_reg[9]/NET0131  ;
  assign n30828 = \P1_P2_InstAddrPointer_reg[11]/NET0131  & \P1_P2_InstAddrPointer_reg[8]/NET0131  ;
  assign n30829 = n30827 & n30828 ;
  assign n30830 = n30826 & n30829 ;
  assign n30831 = n30824 & n30830 ;
  assign n30832 = \P1_P2_InstAddrPointer_reg[24]/NET0131  & n30831 ;
  assign n30833 = n30816 & n30832 ;
  assign n30834 = \P1_P2_InstAddrPointer_reg[25]/NET0131  & n30833 ;
  assign n30835 = \P1_P2_InstAddrPointer_reg[26]/NET0131  & n30834 ;
  assign n31180 = \P1_P2_InstAddrPointer_reg[0]/NET0131  & n30835 ;
  assign n31181 = n31170 & n31180 ;
  assign n31182 = \P1_P2_InstAddrPointer_reg[30]/NET0131  & n31181 ;
  assign n31183 = \P1_P2_InstAddrPointer_reg[31]/NET0131  & ~n31182 ;
  assign n31184 = ~\P1_P2_InstAddrPointer_reg[31]/NET0131  & n31182 ;
  assign n31185 = ~n31183 & ~n31184 ;
  assign n30848 = n30816 & n30829 ;
  assign n31123 = n30825 & n30848 ;
  assign n31159 = \P1_P2_InstAddrPointer_reg[24]/NET0131  & \P1_P2_InstAddrPointer_reg[25]/NET0131  ;
  assign n31160 = \P1_P2_InstAddrPointer_reg[14]/NET0131  & n31159 ;
  assign n31161 = n30824 & n31160 ;
  assign n31162 = n31123 & n31161 ;
  assign n31163 = \P1_P2_InstAddrPointer_reg[26]/NET0131  & n31162 ;
  assign n31171 = n31163 & n31170 ;
  assign n31186 = \P1_P2_InstAddrPointer_reg[0]/NET0131  & n31171 ;
  assign n31187 = \P1_P2_InstAddrPointer_reg[30]/NET0131  & ~n31186 ;
  assign n31188 = ~\P1_P2_InstAddrPointer_reg[30]/NET0131  & n31186 ;
  assign n31189 = ~n31187 & ~n31188 ;
  assign n30846 = \P1_P2_InstAddrPointer_reg[15]/NET0131  & n30826 ;
  assign n30847 = \P1_P2_InstAddrPointer_reg[16]/NET0131  & n30846 ;
  assign n31190 = \P1_P2_InstAddrPointer_reg[0]/NET0131  & n30848 ;
  assign n31191 = n30847 & n31190 ;
  assign n31192 = n30820 & n31191 ;
  assign n31193 = ~\P1_P2_InstAddrPointer_reg[21]/NET0131  & ~n31192 ;
  assign n30844 = n30816 & n30830 ;
  assign n30845 = n30823 & n30844 ;
  assign n31194 = \P1_P2_InstAddrPointer_reg[0]/NET0131  & n30845 ;
  assign n31195 = ~n31193 & ~n31194 ;
  assign n31196 = \P1_P2_InstAddrPointer_reg[0]/NET0131  & \P1_P2_InstAddrPointer_reg[1]/NET0131  ;
  assign n31197 = \P1_P2_InstAddrPointer_reg[2]/NET0131  & n31196 ;
  assign n31198 = \P1_P2_InstAddrPointer_reg[3]/NET0131  & n31197 ;
  assign n31199 = \P1_P2_InstAddrPointer_reg[4]/NET0131  & n31198 ;
  assign n31200 = \P1_P2_InstAddrPointer_reg[5]/NET0131  & n31199 ;
  assign n31201 = \P1_P2_InstAddrPointer_reg[6]/NET0131  & n31200 ;
  assign n31202 = \P1_P2_InstAddrPointer_reg[7]/NET0131  & n31201 ;
  assign n31203 = \P1_P2_InstAddrPointer_reg[8]/NET0131  & n31202 ;
  assign n31204 = \P1_P2_InstAddrPointer_reg[9]/NET0131  & n31203 ;
  assign n31205 = ~\P1_P2_InstAddrPointer_reg[10]/NET0131  & ~n31204 ;
  assign n31206 = n30827 & n31203 ;
  assign n31207 = ~n31205 & ~n31206 ;
  assign n31208 = ~\P1_P2_InstAddrPointer_reg[9]/NET0131  & ~n31203 ;
  assign n31209 = ~n31204 & ~n31208 ;
  assign n31210 = ~\P1_P2_InstAddrPointer_reg[8]/NET0131  & ~n31202 ;
  assign n31211 = ~n31203 & ~n31210 ;
  assign n31212 = ~\P1_P2_InstAddrPointer_reg[7]/NET0131  & ~n31201 ;
  assign n31213 = ~n31202 & ~n31212 ;
  assign n30869 = \P1_P2_InstQueue_reg[7][6]/NET0131  & n25453 ;
  assign n30862 = \P1_P2_InstQueue_reg[8][6]/NET0131  & n25435 ;
  assign n30858 = \P1_P2_InstQueue_reg[6][6]/NET0131  & n25449 ;
  assign n30859 = \P1_P2_InstQueue_reg[14][6]/NET0131  & n25442 ;
  assign n30874 = ~n30858 & ~n30859 ;
  assign n30884 = ~n30862 & n30874 ;
  assign n30885 = ~n30869 & n30884 ;
  assign n30870 = \P1_P2_InstQueue_reg[3][6]/NET0131  & n25444 ;
  assign n30871 = \P1_P2_InstQueue_reg[13][6]/NET0131  & n25422 ;
  assign n30879 = ~n30870 & ~n30871 ;
  assign n30872 = \P1_P2_InstQueue_reg[4][6]/NET0131  & n25437 ;
  assign n30873 = \P1_P2_InstQueue_reg[11][6]/NET0131  & n25440 ;
  assign n30880 = ~n30872 & ~n30873 ;
  assign n30881 = n30879 & n30880 ;
  assign n30865 = \P1_P2_InstQueue_reg[2][6]/NET0131  & n25428 ;
  assign n30866 = \P1_P2_InstQueue_reg[9][6]/NET0131  & n25455 ;
  assign n30877 = ~n30865 & ~n30866 ;
  assign n30867 = \P1_P2_InstQueue_reg[0][6]/NET0131  & n25446 ;
  assign n30868 = \P1_P2_InstQueue_reg[10][6]/NET0131  & n25457 ;
  assign n30878 = ~n30867 & ~n30868 ;
  assign n30882 = n30877 & n30878 ;
  assign n30860 = \P1_P2_InstQueue_reg[12][6]/NET0131  & n25459 ;
  assign n30861 = \P1_P2_InstQueue_reg[15][6]/NET0131  & n25431 ;
  assign n30875 = ~n30860 & ~n30861 ;
  assign n30863 = \P1_P2_InstQueue_reg[1][6]/NET0131  & n25425 ;
  assign n30864 = \P1_P2_InstQueue_reg[5][6]/NET0131  & n25461 ;
  assign n30876 = ~n30863 & ~n30864 ;
  assign n30883 = n30875 & n30876 ;
  assign n30886 = n30882 & n30883 ;
  assign n30887 = n30881 & n30886 ;
  assign n30888 = n30885 & n30887 ;
  assign n31214 = ~\P1_P2_InstAddrPointer_reg[6]/NET0131  & ~n31200 ;
  assign n31215 = ~n31201 & ~n31214 ;
  assign n31216 = ~n30888 & n31215 ;
  assign n31217 = n30888 & ~n31215 ;
  assign n30904 = \P1_P2_InstQueue_reg[7][5]/NET0131  & n25453 ;
  assign n30897 = \P1_P2_InstQueue_reg[8][5]/NET0131  & n25435 ;
  assign n30893 = \P1_P2_InstQueue_reg[11][5]/NET0131  & n25440 ;
  assign n30894 = \P1_P2_InstQueue_reg[9][5]/NET0131  & n25455 ;
  assign n30909 = ~n30893 & ~n30894 ;
  assign n30919 = ~n30897 & n30909 ;
  assign n30920 = ~n30904 & n30919 ;
  assign n30905 = \P1_P2_InstQueue_reg[14][5]/NET0131  & n25442 ;
  assign n30906 = \P1_P2_InstQueue_reg[13][5]/NET0131  & n25422 ;
  assign n30914 = ~n30905 & ~n30906 ;
  assign n30907 = \P1_P2_InstQueue_reg[4][5]/NET0131  & n25437 ;
  assign n30908 = \P1_P2_InstQueue_reg[3][5]/NET0131  & n25444 ;
  assign n30915 = ~n30907 & ~n30908 ;
  assign n30916 = n30914 & n30915 ;
  assign n30900 = \P1_P2_InstQueue_reg[2][5]/NET0131  & n25428 ;
  assign n30901 = \P1_P2_InstQueue_reg[1][5]/NET0131  & n25425 ;
  assign n30912 = ~n30900 & ~n30901 ;
  assign n30902 = \P1_P2_InstQueue_reg[0][5]/NET0131  & n25446 ;
  assign n30903 = \P1_P2_InstQueue_reg[5][5]/NET0131  & n25461 ;
  assign n30913 = ~n30902 & ~n30903 ;
  assign n30917 = n30912 & n30913 ;
  assign n30895 = \P1_P2_InstQueue_reg[10][5]/NET0131  & n25457 ;
  assign n30896 = \P1_P2_InstQueue_reg[15][5]/NET0131  & n25431 ;
  assign n30910 = ~n30895 & ~n30896 ;
  assign n30898 = \P1_P2_InstQueue_reg[6][5]/NET0131  & n25449 ;
  assign n30899 = \P1_P2_InstQueue_reg[12][5]/NET0131  & n25459 ;
  assign n30911 = ~n30898 & ~n30899 ;
  assign n30918 = n30910 & n30911 ;
  assign n30921 = n30917 & n30918 ;
  assign n30922 = n30916 & n30921 ;
  assign n30923 = n30920 & n30922 ;
  assign n31218 = ~\P1_P2_InstAddrPointer_reg[5]/NET0131  & ~n31199 ;
  assign n31219 = ~n31200 & ~n31218 ;
  assign n31220 = ~n30923 & n31219 ;
  assign n31221 = n30923 & ~n31219 ;
  assign n30939 = \P1_P2_InstQueue_reg[7][4]/NET0131  & n25453 ;
  assign n30932 = \P1_P2_InstQueue_reg[8][4]/NET0131  & n25435 ;
  assign n30928 = \P1_P2_InstQueue_reg[6][4]/NET0131  & n25449 ;
  assign n30929 = \P1_P2_InstQueue_reg[2][4]/NET0131  & n25428 ;
  assign n30944 = ~n30928 & ~n30929 ;
  assign n30954 = ~n30932 & n30944 ;
  assign n30955 = ~n30939 & n30954 ;
  assign n30940 = \P1_P2_InstQueue_reg[11][4]/NET0131  & n25440 ;
  assign n30941 = \P1_P2_InstQueue_reg[1][4]/NET0131  & n25425 ;
  assign n30949 = ~n30940 & ~n30941 ;
  assign n30942 = \P1_P2_InstQueue_reg[4][4]/NET0131  & n25437 ;
  assign n30943 = \P1_P2_InstQueue_reg[9][4]/NET0131  & n25455 ;
  assign n30950 = ~n30942 & ~n30943 ;
  assign n30951 = n30949 & n30950 ;
  assign n30935 = \P1_P2_InstQueue_reg[13][4]/NET0131  & n25422 ;
  assign n30936 = \P1_P2_InstQueue_reg[3][4]/NET0131  & n25444 ;
  assign n30947 = ~n30935 & ~n30936 ;
  assign n30937 = \P1_P2_InstQueue_reg[0][4]/NET0131  & n25446 ;
  assign n30938 = \P1_P2_InstQueue_reg[10][4]/NET0131  & n25457 ;
  assign n30948 = ~n30937 & ~n30938 ;
  assign n30952 = n30947 & n30948 ;
  assign n30930 = \P1_P2_InstQueue_reg[14][4]/NET0131  & n25442 ;
  assign n30931 = \P1_P2_InstQueue_reg[15][4]/NET0131  & n25431 ;
  assign n30945 = ~n30930 & ~n30931 ;
  assign n30933 = \P1_P2_InstQueue_reg[12][4]/NET0131  & n25459 ;
  assign n30934 = \P1_P2_InstQueue_reg[5][4]/NET0131  & n25461 ;
  assign n30946 = ~n30933 & ~n30934 ;
  assign n30953 = n30945 & n30946 ;
  assign n30956 = n30952 & n30953 ;
  assign n30957 = n30951 & n30956 ;
  assign n30958 = n30955 & n30957 ;
  assign n31222 = ~\P1_P2_InstAddrPointer_reg[4]/NET0131  & ~n31198 ;
  assign n31223 = ~n31199 & ~n31222 ;
  assign n31224 = ~n30958 & n31223 ;
  assign n31225 = n30958 & ~n31223 ;
  assign n30974 = \P1_P2_InstQueue_reg[7][3]/NET0131  & n25453 ;
  assign n30967 = \P1_P2_InstQueue_reg[8][3]/NET0131  & n25435 ;
  assign n30963 = \P1_P2_InstQueue_reg[11][3]/NET0131  & n25440 ;
  assign n30964 = \P1_P2_InstQueue_reg[1][3]/NET0131  & n25425 ;
  assign n30979 = ~n30963 & ~n30964 ;
  assign n30989 = ~n30967 & n30979 ;
  assign n30990 = ~n30974 & n30989 ;
  assign n30975 = \P1_P2_InstQueue_reg[9][3]/NET0131  & n25455 ;
  assign n30976 = \P1_P2_InstQueue_reg[14][3]/NET0131  & n25442 ;
  assign n30984 = ~n30975 & ~n30976 ;
  assign n30977 = \P1_P2_InstQueue_reg[4][3]/NET0131  & n25437 ;
  assign n30978 = \P1_P2_InstQueue_reg[6][3]/NET0131  & n25449 ;
  assign n30985 = ~n30977 & ~n30978 ;
  assign n30986 = n30984 & n30985 ;
  assign n30970 = \P1_P2_InstQueue_reg[2][3]/NET0131  & n25428 ;
  assign n30971 = \P1_P2_InstQueue_reg[10][3]/NET0131  & n25457 ;
  assign n30982 = ~n30970 & ~n30971 ;
  assign n30972 = \P1_P2_InstQueue_reg[0][3]/NET0131  & n25446 ;
  assign n30973 = \P1_P2_InstQueue_reg[13][3]/NET0131  & n25422 ;
  assign n30983 = ~n30972 & ~n30973 ;
  assign n30987 = n30982 & n30983 ;
  assign n30965 = \P1_P2_InstQueue_reg[12][3]/NET0131  & n25459 ;
  assign n30966 = \P1_P2_InstQueue_reg[15][3]/NET0131  & n25431 ;
  assign n30980 = ~n30965 & ~n30966 ;
  assign n30968 = \P1_P2_InstQueue_reg[3][3]/NET0131  & n25444 ;
  assign n30969 = \P1_P2_InstQueue_reg[5][3]/NET0131  & n25461 ;
  assign n30981 = ~n30968 & ~n30969 ;
  assign n30988 = n30980 & n30981 ;
  assign n30991 = n30987 & n30988 ;
  assign n30992 = n30986 & n30991 ;
  assign n30993 = n30990 & n30992 ;
  assign n31226 = ~\P1_P2_InstAddrPointer_reg[3]/NET0131  & ~n31197 ;
  assign n31227 = ~n31198 & ~n31226 ;
  assign n31228 = ~n30993 & n31227 ;
  assign n31229 = n30993 & ~n31227 ;
  assign n31002 = \P1_P2_InstQueue_reg[8][2]/NET0131  & n25435 ;
  assign n30999 = \P1_P2_InstQueue_reg[7][2]/NET0131  & n25453 ;
  assign n30998 = \P1_P2_InstQueue_reg[1][2]/NET0131  & n25425 ;
  assign n31000 = \P1_P2_InstQueue_reg[4][2]/NET0131  & n25437 ;
  assign n31014 = ~n30998 & ~n31000 ;
  assign n31024 = ~n30999 & n31014 ;
  assign n31025 = ~n31002 & n31024 ;
  assign n31010 = \P1_P2_InstQueue_reg[13][2]/NET0131  & n25422 ;
  assign n31011 = \P1_P2_InstQueue_reg[14][2]/NET0131  & n25442 ;
  assign n31019 = ~n31010 & ~n31011 ;
  assign n31012 = \P1_P2_InstQueue_reg[11][2]/NET0131  & n25440 ;
  assign n31013 = \P1_P2_InstQueue_reg[2][2]/NET0131  & n25428 ;
  assign n31020 = ~n31012 & ~n31013 ;
  assign n31021 = n31019 & n31020 ;
  assign n31006 = \P1_P2_InstQueue_reg[10][2]/NET0131  & n25457 ;
  assign n31007 = \P1_P2_InstQueue_reg[6][2]/NET0131  & n25449 ;
  assign n31017 = ~n31006 & ~n31007 ;
  assign n31008 = \P1_P2_InstQueue_reg[0][2]/NET0131  & n25446 ;
  assign n31009 = \P1_P2_InstQueue_reg[9][2]/NET0131  & n25455 ;
  assign n31018 = ~n31008 & ~n31009 ;
  assign n31022 = n31017 & n31018 ;
  assign n31001 = \P1_P2_InstQueue_reg[15][2]/NET0131  & n25431 ;
  assign n31003 = \P1_P2_InstQueue_reg[12][2]/NET0131  & n25459 ;
  assign n31015 = ~n31001 & ~n31003 ;
  assign n31004 = \P1_P2_InstQueue_reg[5][2]/NET0131  & n25461 ;
  assign n31005 = \P1_P2_InstQueue_reg[3][2]/NET0131  & n25444 ;
  assign n31016 = ~n31004 & ~n31005 ;
  assign n31023 = n31015 & n31016 ;
  assign n31026 = n31022 & n31023 ;
  assign n31027 = n31021 & n31026 ;
  assign n31028 = n31025 & n31027 ;
  assign n31230 = ~\P1_P2_InstAddrPointer_reg[2]/NET0131  & ~n31196 ;
  assign n31231 = ~n31197 & ~n31230 ;
  assign n31232 = ~n31028 & n31231 ;
  assign n31233 = n31028 & ~n31231 ;
  assign n31043 = \P1_P2_InstQueue_reg[7][1]/NET0131  & n25453 ;
  assign n31031 = \P1_P2_InstQueue_reg[8][1]/NET0131  & n25435 ;
  assign n31032 = \P1_P2_InstQueue_reg[9][1]/NET0131  & n25455 ;
  assign n31033 = \P1_P2_InstQueue_reg[6][1]/NET0131  & n25449 ;
  assign n31047 = ~n31032 & ~n31033 ;
  assign n31057 = ~n31031 & n31047 ;
  assign n31058 = ~n31043 & n31057 ;
  assign n31042 = \P1_P2_InstQueue_reg[0][1]/NET0131  & n25446 ;
  assign n31044 = \P1_P2_InstQueue_reg[2][1]/NET0131  & n25428 ;
  assign n31052 = ~n31042 & ~n31044 ;
  assign n31045 = \P1_P2_InstQueue_reg[11][1]/NET0131  & n25440 ;
  assign n31046 = \P1_P2_InstQueue_reg[5][1]/NET0131  & n25461 ;
  assign n31053 = ~n31045 & ~n31046 ;
  assign n31054 = n31052 & n31053 ;
  assign n31038 = \P1_P2_InstQueue_reg[1][1]/NET0131  & n25425 ;
  assign n31039 = \P1_P2_InstQueue_reg[13][1]/NET0131  & n25422 ;
  assign n31050 = ~n31038 & ~n31039 ;
  assign n31040 = \P1_P2_InstQueue_reg[10][1]/NET0131  & n25457 ;
  assign n31041 = \P1_P2_InstQueue_reg[14][1]/NET0131  & n25442 ;
  assign n31051 = ~n31040 & ~n31041 ;
  assign n31055 = n31050 & n31051 ;
  assign n31034 = \P1_P2_InstQueue_reg[12][1]/NET0131  & n25459 ;
  assign n31035 = \P1_P2_InstQueue_reg[15][1]/NET0131  & n25431 ;
  assign n31048 = ~n31034 & ~n31035 ;
  assign n31036 = \P1_P2_InstQueue_reg[4][1]/NET0131  & n25437 ;
  assign n31037 = \P1_P2_InstQueue_reg[3][1]/NET0131  & n25444 ;
  assign n31049 = ~n31036 & ~n31037 ;
  assign n31056 = n31048 & n31049 ;
  assign n31059 = n31055 & n31056 ;
  assign n31060 = n31054 & n31059 ;
  assign n31061 = n31058 & n31060 ;
  assign n31062 = ~\P1_P2_InstAddrPointer_reg[1]/NET0131  & ~n31061 ;
  assign n31063 = \P1_P2_InstAddrPointer_reg[1]/NET0131  & n31061 ;
  assign n31076 = \P1_P2_InstQueue_reg[7][0]/NET0131  & n25453 ;
  assign n31064 = \P1_P2_InstQueue_reg[8][0]/NET0131  & n25435 ;
  assign n31065 = \P1_P2_InstQueue_reg[2][0]/NET0131  & n25428 ;
  assign n31066 = \P1_P2_InstQueue_reg[12][0]/NET0131  & n25459 ;
  assign n31080 = ~n31065 & ~n31066 ;
  assign n31090 = ~n31064 & n31080 ;
  assign n31091 = ~n31076 & n31090 ;
  assign n31075 = \P1_P2_InstQueue_reg[0][0]/NET0131  & n25446 ;
  assign n31077 = \P1_P2_InstQueue_reg[4][0]/NET0131  & n25437 ;
  assign n31085 = ~n31075 & ~n31077 ;
  assign n31078 = \P1_P2_InstQueue_reg[11][0]/NET0131  & n25440 ;
  assign n31079 = \P1_P2_InstQueue_reg[10][0]/NET0131  & n25457 ;
  assign n31086 = ~n31078 & ~n31079 ;
  assign n31087 = n31085 & n31086 ;
  assign n31071 = \P1_P2_InstQueue_reg[13][0]/NET0131  & n25422 ;
  assign n31072 = \P1_P2_InstQueue_reg[5][0]/NET0131  & n25461 ;
  assign n31083 = ~n31071 & ~n31072 ;
  assign n31073 = \P1_P2_InstQueue_reg[6][0]/NET0131  & n25449 ;
  assign n31074 = \P1_P2_InstQueue_reg[3][0]/NET0131  & n25444 ;
  assign n31084 = ~n31073 & ~n31074 ;
  assign n31088 = n31083 & n31084 ;
  assign n31067 = \P1_P2_InstQueue_reg[9][0]/NET0131  & n25455 ;
  assign n31068 = \P1_P2_InstQueue_reg[15][0]/NET0131  & n25431 ;
  assign n31081 = ~n31067 & ~n31068 ;
  assign n31069 = \P1_P2_InstQueue_reg[1][0]/NET0131  & n25425 ;
  assign n31070 = \P1_P2_InstQueue_reg[14][0]/NET0131  & n25442 ;
  assign n31082 = ~n31069 & ~n31070 ;
  assign n31089 = n31081 & n31082 ;
  assign n31092 = n31088 & n31089 ;
  assign n31093 = n31087 & n31092 ;
  assign n31094 = n31091 & n31093 ;
  assign n31095 = \P1_P2_InstAddrPointer_reg[0]/NET0131  & ~n31094 ;
  assign n31096 = ~n31063 & n31095 ;
  assign n31097 = ~n31062 & ~n31096 ;
  assign n31234 = ~\P1_P2_InstAddrPointer_reg[0]/NET0131  & \P1_P2_InstAddrPointer_reg[1]/NET0131  ;
  assign n31235 = n31097 & ~n31234 ;
  assign n31236 = ~n31233 & ~n31235 ;
  assign n31237 = ~n31232 & ~n31236 ;
  assign n31238 = ~n31229 & ~n31237 ;
  assign n31239 = ~n31228 & ~n31238 ;
  assign n31240 = ~n31225 & ~n31239 ;
  assign n31241 = ~n31224 & ~n31240 ;
  assign n31242 = ~n31221 & ~n31241 ;
  assign n31243 = ~n31220 & ~n31242 ;
  assign n31244 = ~n31217 & ~n31243 ;
  assign n31245 = ~n31216 & ~n31244 ;
  assign n31246 = n31213 & ~n31245 ;
  assign n30790 = \P1_P2_InstQueue_reg[7][7]/NET0131  & n25453 ;
  assign n30783 = \P1_P2_InstQueue_reg[8][7]/NET0131  & n25435 ;
  assign n30779 = \P1_P2_InstQueue_reg[10][7]/NET0131  & n25457 ;
  assign n30780 = \P1_P2_InstQueue_reg[2][7]/NET0131  & n25428 ;
  assign n30795 = ~n30779 & ~n30780 ;
  assign n30805 = ~n30783 & n30795 ;
  assign n30806 = ~n30790 & n30805 ;
  assign n30791 = \P1_P2_InstQueue_reg[11][7]/NET0131  & n25440 ;
  assign n30792 = \P1_P2_InstQueue_reg[14][7]/NET0131  & n25442 ;
  assign n30800 = ~n30791 & ~n30792 ;
  assign n30793 = \P1_P2_InstQueue_reg[6][7]/NET0131  & n25449 ;
  assign n30794 = \P1_P2_InstQueue_reg[1][7]/NET0131  & n25425 ;
  assign n30801 = ~n30793 & ~n30794 ;
  assign n30802 = n30800 & n30801 ;
  assign n30786 = \P1_P2_InstQueue_reg[13][7]/NET0131  & n25422 ;
  assign n30787 = \P1_P2_InstQueue_reg[9][7]/NET0131  & n25455 ;
  assign n30798 = ~n30786 & ~n30787 ;
  assign n30788 = \P1_P2_InstQueue_reg[0][7]/NET0131  & n25446 ;
  assign n30789 = \P1_P2_InstQueue_reg[5][7]/NET0131  & n25461 ;
  assign n30799 = ~n30788 & ~n30789 ;
  assign n30803 = n30798 & n30799 ;
  assign n30781 = \P1_P2_InstQueue_reg[3][7]/NET0131  & n25444 ;
  assign n30782 = \P1_P2_InstQueue_reg[15][7]/NET0131  & n25431 ;
  assign n30796 = ~n30781 & ~n30782 ;
  assign n30784 = \P1_P2_InstQueue_reg[4][7]/NET0131  & n25437 ;
  assign n30785 = \P1_P2_InstQueue_reg[12][7]/NET0131  & n25459 ;
  assign n30797 = ~n30784 & ~n30785 ;
  assign n30804 = n30796 & n30797 ;
  assign n30807 = n30803 & n30804 ;
  assign n30808 = n30802 & n30807 ;
  assign n30809 = n30806 & n30808 ;
  assign n31247 = ~n31213 & n31245 ;
  assign n31248 = ~n30809 & ~n31247 ;
  assign n31249 = ~n31246 & ~n31248 ;
  assign n31250 = ~n31211 & n31249 ;
  assign n31251 = ~n31209 & n31250 ;
  assign n31252 = ~n31207 & n31251 ;
  assign n31253 = ~\P1_P2_InstAddrPointer_reg[11]/NET0131  & ~n31206 ;
  assign n31254 = ~n31190 & ~n31253 ;
  assign n31255 = n31252 & ~n31254 ;
  assign n31256 = ~\P1_P2_InstAddrPointer_reg[12]/NET0131  & ~n31190 ;
  assign n31257 = \P1_P2_InstAddrPointer_reg[11]/NET0131  & \P1_P2_InstAddrPointer_reg[12]/NET0131  ;
  assign n31258 = n31206 & n31257 ;
  assign n31259 = ~n31256 & ~n31258 ;
  assign n31260 = n31255 & ~n31259 ;
  assign n31261 = ~\P1_P2_InstAddrPointer_reg[13]/NET0131  & ~n31258 ;
  assign n31262 = n30825 & n31190 ;
  assign n31263 = ~n31261 & ~n31262 ;
  assign n31264 = n31260 & ~n31263 ;
  assign n31265 = ~\P1_P2_InstAddrPointer_reg[14]/NET0131  & ~n31262 ;
  assign n31266 = \P1_P2_InstAddrPointer_reg[0]/NET0131  & n30844 ;
  assign n31267 = ~n31265 & ~n31266 ;
  assign n31268 = n31264 & ~n31267 ;
  assign n31269 = ~\P1_P2_InstAddrPointer_reg[15]/NET0131  & ~n31266 ;
  assign n31270 = n30846 & n31190 ;
  assign n31271 = ~n31269 & ~n31270 ;
  assign n31272 = n31268 & ~n31271 ;
  assign n31273 = ~\P1_P2_InstAddrPointer_reg[16]/NET0131  & ~n31270 ;
  assign n31274 = ~n31191 & ~n31273 ;
  assign n31275 = n31272 & ~n31274 ;
  assign n30849 = n30847 & n30848 ;
  assign n31128 = n30819 & n30849 ;
  assign n31276 = \P1_P2_InstAddrPointer_reg[0]/NET0131  & n31128 ;
  assign n31280 = \P1_P2_InstAddrPointer_reg[17]/NET0131  & n31191 ;
  assign n31282 = \P1_P2_InstAddrPointer_reg[18]/NET0131  & n31280 ;
  assign n31283 = ~\P1_P2_InstAddrPointer_reg[19]/NET0131  & ~n31282 ;
  assign n31284 = ~n31276 & ~n31283 ;
  assign n31285 = ~\P1_P2_InstAddrPointer_reg[18]/NET0131  & ~n31280 ;
  assign n31286 = ~n31282 & ~n31285 ;
  assign n31287 = ~n31284 & ~n31286 ;
  assign n31277 = ~\P1_P2_InstAddrPointer_reg[20]/NET0131  & ~n31276 ;
  assign n31278 = ~n31192 & ~n31277 ;
  assign n31279 = ~\P1_P2_InstAddrPointer_reg[17]/NET0131  & ~n31191 ;
  assign n31281 = ~n31279 & ~n31280 ;
  assign n31288 = ~n31278 & ~n31281 ;
  assign n31289 = n31287 & n31288 ;
  assign n31290 = n31275 & n31289 ;
  assign n31291 = ~n31195 & n31290 ;
  assign n31292 = ~\P1_P2_InstAddrPointer_reg[22]/NET0131  & ~n31194 ;
  assign n31293 = \P1_P2_InstAddrPointer_reg[22]/NET0131  & n31194 ;
  assign n31294 = ~n31292 & ~n31293 ;
  assign n31295 = n31291 & ~n31294 ;
  assign n31296 = n30817 & n31194 ;
  assign n31297 = \P1_P2_InstAddrPointer_reg[24]/NET0131  & n31296 ;
  assign n31298 = ~\P1_P2_InstAddrPointer_reg[25]/NET0131  & ~n31297 ;
  assign n31299 = \P1_P2_InstAddrPointer_reg[25]/NET0131  & n31297 ;
  assign n31300 = ~n31298 & ~n31299 ;
  assign n31301 = ~\P1_P2_InstAddrPointer_reg[23]/NET0131  & ~n31293 ;
  assign n31302 = ~n31296 & ~n31301 ;
  assign n31303 = \P1_P2_InstAddrPointer_reg[24]/NET0131  & ~n31202 ;
  assign n31304 = ~\P1_P2_InstAddrPointer_reg[24]/NET0131  & ~n30831 ;
  assign n31305 = ~n30832 & ~n31304 ;
  assign n31306 = n31202 & n31305 ;
  assign n31307 = ~n31303 & ~n31306 ;
  assign n31308 = ~n31302 & n31307 ;
  assign n31309 = ~n31300 & n31308 ;
  assign n31310 = n31295 & n31309 ;
  assign n31311 = n30810 & n31180 ;
  assign n31318 = \P1_P2_InstAddrPointer_reg[27]/NET0131  & n31180 ;
  assign n31319 = ~\P1_P2_InstAddrPointer_reg[28]/NET0131  & ~n31318 ;
  assign n31320 = ~n31311 & ~n31319 ;
  assign n31321 = ~\P1_P2_InstAddrPointer_reg[27]/NET0131  & ~n31180 ;
  assign n31322 = ~n31318 & ~n31321 ;
  assign n31323 = ~n31320 & ~n31322 ;
  assign n31312 = ~\P1_P2_InstAddrPointer_reg[29]/NET0131  & ~n31311 ;
  assign n31313 = ~n31181 & ~n31312 ;
  assign n31314 = n31161 & n31262 ;
  assign n31315 = \P1_P2_InstAddrPointer_reg[26]/NET0131  & ~n31314 ;
  assign n31316 = ~\P1_P2_InstAddrPointer_reg[26]/NET0131  & n31314 ;
  assign n31317 = ~n31315 & ~n31316 ;
  assign n31324 = ~n31313 & n31317 ;
  assign n31325 = n31323 & n31324 ;
  assign n31326 = n31310 & n31325 ;
  assign n31327 = n31189 & n31326 ;
  assign n31329 = n31185 & n31327 ;
  assign n31328 = ~n31185 & ~n31327 ;
  assign n31330 = ~n30809 & ~n31328 ;
  assign n31331 = ~n31329 & n31330 ;
  assign n30836 = n30810 & n30835 ;
  assign n30837 = \P1_P2_InstAddrPointer_reg[29]/NET0131  & n30836 ;
  assign n30838 = \P1_P2_InstAddrPointer_reg[30]/NET0131  & n30837 ;
  assign n30839 = \P1_P2_InstAddrPointer_reg[31]/NET0131  & ~n30838 ;
  assign n30840 = ~\P1_P2_InstAddrPointer_reg[31]/NET0131  & n30838 ;
  assign n30841 = ~n30839 & ~n30840 ;
  assign n30842 = ~\P1_P2_InstAddrPointer_reg[29]/NET0131  & ~n30836 ;
  assign n30843 = ~n30837 & ~n30842 ;
  assign n30850 = n30820 & n30849 ;
  assign n30851 = ~\P1_P2_InstAddrPointer_reg[21]/NET0131  & ~n30850 ;
  assign n30852 = ~n30845 & ~n30851 ;
  assign n30853 = \P1_P2_InstAddrPointer_reg[8]/NET0131  & n30816 ;
  assign n30854 = ~\P1_P2_InstAddrPointer_reg[8]/NET0131  & ~n30816 ;
  assign n30855 = ~n30853 & ~n30854 ;
  assign n30856 = ~\P1_P2_InstAddrPointer_reg[6]/NET0131  & ~n30814 ;
  assign n30857 = ~n30815 & ~n30856 ;
  assign n30889 = n30857 & ~n30888 ;
  assign n30890 = ~n30857 & n30888 ;
  assign n30891 = ~\P1_P2_InstAddrPointer_reg[5]/NET0131  & ~n30813 ;
  assign n30892 = ~n30814 & ~n30891 ;
  assign n30924 = n30892 & ~n30923 ;
  assign n30925 = ~n30892 & n30923 ;
  assign n30926 = ~\P1_P2_InstAddrPointer_reg[4]/NET0131  & ~n30812 ;
  assign n30927 = ~n30813 & ~n30926 ;
  assign n30959 = n30927 & ~n30958 ;
  assign n30960 = ~n30927 & n30958 ;
  assign n30961 = ~\P1_P2_InstAddrPointer_reg[3]/NET0131  & ~n30811 ;
  assign n30962 = ~n30812 & ~n30961 ;
  assign n30994 = n30962 & ~n30993 ;
  assign n30995 = ~n30962 & n30993 ;
  assign n30996 = ~\P1_P2_InstAddrPointer_reg[1]/NET0131  & ~\P1_P2_InstAddrPointer_reg[2]/NET0131  ;
  assign n30997 = ~n30811 & ~n30996 ;
  assign n31029 = n30997 & ~n31028 ;
  assign n31030 = ~n30997 & n31028 ;
  assign n31098 = ~n31030 & ~n31097 ;
  assign n31099 = ~n31029 & ~n31098 ;
  assign n31100 = ~n30995 & ~n31099 ;
  assign n31101 = ~n30994 & ~n31100 ;
  assign n31102 = ~n30960 & ~n31101 ;
  assign n31103 = ~n30959 & ~n31102 ;
  assign n31104 = ~n30925 & ~n31103 ;
  assign n31105 = ~n30924 & ~n31104 ;
  assign n31106 = ~n30890 & ~n31105 ;
  assign n31107 = ~n30889 & ~n31106 ;
  assign n31108 = ~\P1_P2_InstAddrPointer_reg[7]/NET0131  & ~n30815 ;
  assign n31109 = ~n30816 & ~n31108 ;
  assign n31110 = ~n31107 & n31109 ;
  assign n31111 = n31107 & ~n31109 ;
  assign n31112 = ~n30809 & ~n31111 ;
  assign n31113 = ~n31110 & ~n31112 ;
  assign n31114 = n30855 & ~n31113 ;
  assign n31115 = \P1_P2_InstAddrPointer_reg[9]/NET0131  & n31114 ;
  assign n31116 = \P1_P2_InstAddrPointer_reg[9]/NET0131  & n30853 ;
  assign n31117 = ~\P1_P2_InstAddrPointer_reg[10]/NET0131  & ~n31116 ;
  assign n31118 = \P1_P2_InstAddrPointer_reg[10]/NET0131  & n31116 ;
  assign n31119 = ~n31117 & ~n31118 ;
  assign n31120 = n31115 & n31119 ;
  assign n31121 = \P1_P2_InstAddrPointer_reg[11]/NET0131  & n31120 ;
  assign n31122 = n30825 & n31121 ;
  assign n31124 = ~\P1_P2_InstAddrPointer_reg[14]/NET0131  & ~n31123 ;
  assign n31125 = ~n30844 & ~n31124 ;
  assign n31126 = n31122 & n31125 ;
  assign n31127 = \P1_P2_InstAddrPointer_reg[15]/NET0131  & n31126 ;
  assign n31131 = \P1_P2_InstAddrPointer_reg[17]/NET0131  & n30849 ;
  assign n31132 = \P1_P2_InstAddrPointer_reg[18]/NET0131  & n31131 ;
  assign n31133 = ~\P1_P2_InstAddrPointer_reg[19]/NET0131  & ~n31132 ;
  assign n31134 = ~n31128 & ~n31133 ;
  assign n31135 = n30846 & n30848 ;
  assign n31136 = ~\P1_P2_InstAddrPointer_reg[16]/NET0131  & ~n31135 ;
  assign n31137 = ~n30849 & ~n31136 ;
  assign n31138 = \P1_P2_InstAddrPointer_reg[17]/NET0131  & n31137 ;
  assign n31129 = ~\P1_P2_InstAddrPointer_reg[20]/NET0131  & ~n31128 ;
  assign n31130 = ~n30850 & ~n31129 ;
  assign n31139 = \P1_P2_InstAddrPointer_reg[18]/NET0131  & n31130 ;
  assign n31140 = n31138 & n31139 ;
  assign n31141 = n31134 & n31140 ;
  assign n31142 = n31127 & n31141 ;
  assign n31143 = n30852 & n31142 ;
  assign n31144 = \P1_P2_InstAddrPointer_reg[22]/NET0131  & n30845 ;
  assign n31147 = ~\P1_P2_InstAddrPointer_reg[23]/NET0131  & ~n31144 ;
  assign n31148 = n30824 & n30844 ;
  assign n31149 = ~n31147 & ~n31148 ;
  assign n31145 = ~\P1_P2_InstAddrPointer_reg[22]/NET0131  & ~n30845 ;
  assign n31146 = ~n31144 & ~n31145 ;
  assign n31150 = \P1_P2_InstAddrPointer_reg[24]/NET0131  & n31146 ;
  assign n31151 = n31149 & n31150 ;
  assign n31152 = n31143 & n31151 ;
  assign n31153 = ~\P1_P2_InstAddrPointer_reg[25]/NET0131  & ~n30833 ;
  assign n31154 = ~n30834 & ~n31153 ;
  assign n31155 = n31152 & n31154 ;
  assign n31156 = \P1_P2_InstAddrPointer_reg[27]/NET0131  & n30835 ;
  assign n31157 = ~\P1_P2_InstAddrPointer_reg[27]/NET0131  & ~n30835 ;
  assign n31158 = ~n31156 & ~n31157 ;
  assign n31164 = ~\P1_P2_InstAddrPointer_reg[26]/NET0131  & ~n31162 ;
  assign n31165 = ~n31163 & ~n31164 ;
  assign n31166 = \P1_P2_InstAddrPointer_reg[28]/NET0131  & n31165 ;
  assign n31167 = n31158 & n31166 ;
  assign n31168 = n31155 & n31167 ;
  assign n31169 = n30843 & n31168 ;
  assign n31172 = ~\P1_P2_InstAddrPointer_reg[30]/NET0131  & ~n31171 ;
  assign n31173 = \P1_P2_InstAddrPointer_reg[30]/NET0131  & n31171 ;
  assign n31174 = ~n31172 & ~n31173 ;
  assign n31175 = n31169 & n31174 ;
  assign n31177 = n30841 & n31175 ;
  assign n31176 = ~n30841 & ~n31175 ;
  assign n31178 = n30809 & ~n31176 ;
  assign n31179 = ~n31177 & n31178 ;
  assign n31332 = ~n25733 & ~n31179 ;
  assign n31333 = ~n31331 & n31332 ;
  assign n31334 = ~n30778 & ~n31333 ;
  assign n31335 = n25701 & ~n31334 ;
  assign n31336 = \P1_P2_InstAddrPointer_reg[3]/NET0131  & ~n31230 ;
  assign n31337 = \P1_P2_InstAddrPointer_reg[4]/NET0131  & n31336 ;
  assign n31338 = \P1_P2_InstAddrPointer_reg[5]/NET0131  & n31337 ;
  assign n31339 = \P1_P2_InstAddrPointer_reg[6]/NET0131  & n31338 ;
  assign n31340 = \P1_P2_InstAddrPointer_reg[7]/NET0131  & n31339 ;
  assign n31341 = n30830 & n31340 ;
  assign n31342 = n30824 & n31341 ;
  assign n31343 = n31159 & n31342 ;
  assign n31344 = \P1_P2_InstAddrPointer_reg[26]/NET0131  & n31343 ;
  assign n31345 = n31170 & n31344 ;
  assign n31346 = \P1_P2_InstAddrPointer_reg[30]/NET0131  & n31345 ;
  assign n31347 = \P1_P2_InstAddrPointer_reg[31]/NET0131  & ~n31346 ;
  assign n31348 = ~\P1_P2_InstAddrPointer_reg[31]/NET0131  & n31346 ;
  assign n31349 = ~n31347 & ~n31348 ;
  assign n31350 = n30829 & n31340 ;
  assign n31351 = n30825 & n31350 ;
  assign n31352 = n31161 & n31351 ;
  assign n31353 = \P1_P2_InstAddrPointer_reg[26]/NET0131  & n31352 ;
  assign n31354 = n31170 & n31353 ;
  assign n31355 = \P1_P2_InstAddrPointer_reg[30]/NET0131  & ~n31354 ;
  assign n31356 = ~\P1_P2_InstAddrPointer_reg[30]/NET0131  & n31354 ;
  assign n31357 = ~n31355 & ~n31356 ;
  assign n31358 = n30846 & n31350 ;
  assign n31359 = \P1_P2_InstAddrPointer_reg[16]/NET0131  & n31358 ;
  assign n31360 = n30819 & n31359 ;
  assign n31361 = ~\P1_P2_InstAddrPointer_reg[20]/NET0131  & ~n31360 ;
  assign n31362 = n30820 & n31359 ;
  assign n31363 = ~n31361 & ~n31362 ;
  assign n31364 = \P1_P2_InstAddrPointer_reg[8]/NET0131  & n31340 ;
  assign n31365 = n30827 & n31364 ;
  assign n31366 = n31257 & n31365 ;
  assign n31367 = ~\P1_P2_InstAddrPointer_reg[13]/NET0131  & ~n31366 ;
  assign n31368 = ~n31351 & ~n31367 ;
  assign n31369 = ~\P1_P2_InstAddrPointer_reg[8]/NET0131  & ~n31340 ;
  assign n31370 = ~n31364 & ~n31369 ;
  assign n31371 = ~\P1_P2_InstAddrPointer_reg[7]/NET0131  & ~n31339 ;
  assign n31372 = ~n31340 & ~n31371 ;
  assign n31373 = ~n30809 & n31372 ;
  assign n31374 = n30809 & ~n31372 ;
  assign n31375 = ~\P1_P2_InstAddrPointer_reg[6]/NET0131  & ~n31338 ;
  assign n31376 = ~n31339 & ~n31375 ;
  assign n31377 = ~n30888 & n31376 ;
  assign n31378 = n30888 & ~n31376 ;
  assign n31379 = ~\P1_P2_InstAddrPointer_reg[5]/NET0131  & ~n31337 ;
  assign n31380 = ~n31338 & ~n31379 ;
  assign n31381 = ~n30923 & n31380 ;
  assign n31382 = n30923 & ~n31380 ;
  assign n31383 = ~\P1_P2_InstAddrPointer_reg[4]/NET0131  & ~n31336 ;
  assign n31384 = ~n31337 & ~n31383 ;
  assign n31385 = ~n30958 & n31384 ;
  assign n31386 = n30958 & ~n31384 ;
  assign n31387 = ~\P1_P2_InstAddrPointer_reg[3]/NET0131  & n31230 ;
  assign n31388 = ~n31336 & ~n31387 ;
  assign n31389 = ~n30993 & n31388 ;
  assign n31390 = n30993 & ~n31388 ;
  assign n31391 = ~n31028 & ~n31231 ;
  assign n31392 = n31028 & n31231 ;
  assign n31393 = \P1_P2_InstAddrPointer_reg[0]/NET0131  & ~\P1_P2_InstAddrPointer_reg[1]/NET0131  ;
  assign n31394 = ~n31234 & ~n31393 ;
  assign n31395 = ~n31061 & ~n31394 ;
  assign n31396 = n31061 & n31394 ;
  assign n31397 = ~\P1_P2_InstAddrPointer_reg[0]/NET0131  & ~n31094 ;
  assign n31398 = ~n31396 & n31397 ;
  assign n31399 = ~n31395 & ~n31398 ;
  assign n31400 = ~n31392 & ~n31399 ;
  assign n31401 = ~n31391 & ~n31400 ;
  assign n31402 = ~n31390 & ~n31401 ;
  assign n31403 = ~n31389 & ~n31402 ;
  assign n31404 = ~n31386 & ~n31403 ;
  assign n31405 = ~n31385 & ~n31404 ;
  assign n31406 = ~n31382 & ~n31405 ;
  assign n31407 = ~n31381 & ~n31406 ;
  assign n31408 = ~n31378 & ~n31407 ;
  assign n31409 = ~n31377 & ~n31408 ;
  assign n31410 = ~n31374 & ~n31409 ;
  assign n31411 = ~n31373 & ~n31410 ;
  assign n31412 = n31370 & ~n31411 ;
  assign n31413 = \P1_P2_InstAddrPointer_reg[9]/NET0131  & n31412 ;
  assign n31414 = \P1_P2_InstAddrPointer_reg[9]/NET0131  & n31364 ;
  assign n31415 = ~\P1_P2_InstAddrPointer_reg[10]/NET0131  & ~n31414 ;
  assign n31416 = ~n31365 & ~n31415 ;
  assign n31417 = n31413 & n31416 ;
  assign n31418 = n31257 & n31417 ;
  assign n31419 = n31368 & n31418 ;
  assign n31420 = \P1_P2_InstAddrPointer_reg[14]/NET0131  & n31419 ;
  assign n31421 = ~\P1_P2_InstAddrPointer_reg[15]/NET0131  & ~n31341 ;
  assign n31422 = ~n31358 & ~n31421 ;
  assign n31423 = n31420 & n31422 ;
  assign n31424 = \P1_P2_InstAddrPointer_reg[16]/NET0131  & n31423 ;
  assign n31425 = \P1_P2_InstAddrPointer_reg[17]/NET0131  & n31359 ;
  assign n31426 = ~\P1_P2_InstAddrPointer_reg[17]/NET0131  & ~n31359 ;
  assign n31427 = ~n31425 & ~n31426 ;
  assign n31428 = \P1_P2_InstAddrPointer_reg[18]/NET0131  & n31427 ;
  assign n31429 = n31424 & n31428 ;
  assign n31430 = \P1_P2_InstAddrPointer_reg[19]/NET0131  & n31429 ;
  assign n31431 = n31363 & n31430 ;
  assign n31432 = \P1_P2_InstAddrPointer_reg[21]/NET0131  & n31431 ;
  assign n31433 = n30823 & n31341 ;
  assign n31434 = \P1_P2_InstAddrPointer_reg[22]/NET0131  & n31433 ;
  assign n31435 = ~\P1_P2_InstAddrPointer_reg[22]/NET0131  & ~n31433 ;
  assign n31436 = ~n31434 & ~n31435 ;
  assign n31437 = n31432 & n31436 ;
  assign n31438 = \P1_P2_InstAddrPointer_reg[23]/NET0131  & n31437 ;
  assign n31439 = ~n31305 & n31340 ;
  assign n31440 = ~\P1_P2_InstAddrPointer_reg[24]/NET0131  & ~n31340 ;
  assign n31441 = ~n31439 & ~n31440 ;
  assign n31442 = n31438 & n31441 ;
  assign n31446 = ~\P1_P2_InstAddrPointer_reg[26]/NET0131  & ~n31352 ;
  assign n31447 = ~n31353 & ~n31446 ;
  assign n31443 = n30832 & n31340 ;
  assign n31444 = ~\P1_P2_InstAddrPointer_reg[25]/NET0131  & ~n31443 ;
  assign n31445 = ~n31343 & ~n31444 ;
  assign n31448 = \P1_P2_InstAddrPointer_reg[27]/NET0131  & n31445 ;
  assign n31449 = n31447 & n31448 ;
  assign n31450 = n31442 & n31449 ;
  assign n31451 = \P1_P2_InstAddrPointer_reg[28]/NET0131  & n31450 ;
  assign n31452 = \P1_P2_InstAddrPointer_reg[27]/NET0131  & n31344 ;
  assign n31453 = \P1_P2_InstAddrPointer_reg[28]/NET0131  & n31452 ;
  assign n31454 = ~\P1_P2_InstAddrPointer_reg[29]/NET0131  & ~n31453 ;
  assign n31455 = ~n31345 & ~n31454 ;
  assign n31456 = n31451 & n31455 ;
  assign n31457 = ~n31357 & n31456 ;
  assign n31459 = n31349 & ~n31457 ;
  assign n31458 = ~n31349 & n31457 ;
  assign n31460 = n25881 & ~n31458 ;
  assign n31461 = ~n31459 & n31460 ;
  assign n31462 = ~n25817 & ~n31185 ;
  assign n31470 = n25415 & n25776 ;
  assign n31471 = \P1_P2_InstAddrPointer_reg[31]/NET0131  & n31470 ;
  assign n31472 = ~n25415 & ~n30841 ;
  assign n31473 = ~n25828 & n31472 ;
  assign n31474 = ~n31471 & ~n31473 ;
  assign n31475 = ~n25770 & ~n31474 ;
  assign n31466 = ~n25775 & ~n25840 ;
  assign n31467 = n25753 & ~n25772 ;
  assign n31468 = n31466 & n31467 ;
  assign n31469 = \P1_P2_InstAddrPointer_reg[31]/NET0131  & ~n31468 ;
  assign n31463 = \P1_P2_InstAddrPointer_reg[31]/NET0131  & ~n25763 ;
  assign n31464 = ~n25808 & ~n31463 ;
  assign n31465 = ~n30841 & ~n31464 ;
  assign n31476 = n25887 & ~n31349 ;
  assign n31477 = ~n31465 & ~n31476 ;
  assign n31478 = ~n31469 & n31477 ;
  assign n31479 = ~n31475 & n31478 ;
  assign n31480 = ~n31462 & n31479 ;
  assign n31481 = ~n31461 & n31480 ;
  assign n31482 = ~n31335 & n31481 ;
  assign n31483 = n25918 & ~n31482 ;
  assign n31484 = ~n25934 & n27606 ;
  assign n31485 = ~n25921 & ~n25924 ;
  assign n31486 = ~n27898 & n31485 ;
  assign n31487 = ~n31484 & n31486 ;
  assign n31488 = \P1_P2_InstAddrPointer_reg[31]/NET0131  & ~n31487 ;
  assign n31489 = \P1_P2_rEIP_reg[31]/NET0131  & n27967 ;
  assign n31490 = ~n31488 & ~n31489 ;
  assign n31491 = ~n31483 & n31490 ;
  assign n31492 = \P2_P1_InstAddrPointer_reg[31]/NET0131  & n25947 ;
  assign n31493 = \P2_P1_InstAddrPointer_reg[7]/NET0131  & \P2_P1_InstAddrPointer_reg[8]/NET0131  ;
  assign n31494 = \P2_P1_InstAddrPointer_reg[10]/NET0131  & \P2_P1_InstAddrPointer_reg[9]/NET0131  ;
  assign n31495 = n31493 & n31494 ;
  assign n31496 = \P2_P1_InstAddrPointer_reg[6]/NET0131  & n31495 ;
  assign n31497 = \P2_P1_InstAddrPointer_reg[5]/NET0131  & n31496 ;
  assign n31498 = \P2_P1_InstAddrPointer_reg[1]/NET0131  & \P2_P1_InstAddrPointer_reg[2]/NET0131  ;
  assign n31499 = \P2_P1_InstAddrPointer_reg[3]/NET0131  & n31498 ;
  assign n31500 = \P2_P1_InstAddrPointer_reg[4]/NET0131  & n31499 ;
  assign n31501 = n31497 & n31500 ;
  assign n31502 = \P2_P1_InstAddrPointer_reg[11]/NET0131  & n31501 ;
  assign n31505 = \P2_P1_InstAddrPointer_reg[13]/NET0131  & \P2_P1_InstAddrPointer_reg[14]/NET0131  ;
  assign n31506 = \P2_P1_InstAddrPointer_reg[12]/NET0131  & n31505 ;
  assign n31507 = \P2_P1_InstAddrPointer_reg[15]/NET0131  & n31506 ;
  assign n31508 = \P2_P1_InstAddrPointer_reg[16]/NET0131  & n31507 ;
  assign n31509 = \P2_P1_InstAddrPointer_reg[17]/NET0131  & n31508 ;
  assign n31503 = \P2_P1_InstAddrPointer_reg[18]/NET0131  & \P2_P1_InstAddrPointer_reg[19]/NET0131  ;
  assign n31504 = \P2_P1_InstAddrPointer_reg[20]/NET0131  & n31503 ;
  assign n31510 = \P2_P1_InstAddrPointer_reg[21]/NET0131  & \P2_P1_InstAddrPointer_reg[22]/NET0131  ;
  assign n31511 = n31504 & n31510 ;
  assign n31512 = n31509 & n31511 ;
  assign n31513 = n31502 & n31512 ;
  assign n31514 = \P2_P1_InstAddrPointer_reg[23]/NET0131  & n31513 ;
  assign n31515 = \P2_P1_InstAddrPointer_reg[24]/NET0131  & n31514 ;
  assign n31516 = \P2_P1_InstAddrPointer_reg[25]/NET0131  & n31515 ;
  assign n31517 = \P2_P1_InstAddrPointer_reg[26]/NET0131  & n31516 ;
  assign n31518 = \P2_P1_InstAddrPointer_reg[27]/NET0131  & n31517 ;
  assign n31519 = \P2_P1_InstAddrPointer_reg[28]/NET0131  & n31518 ;
  assign n31520 = \P2_P1_InstAddrPointer_reg[29]/NET0131  & n31519 ;
  assign n31521 = \P2_P1_InstAddrPointer_reg[30]/NET0131  & n31520 ;
  assign n31522 = ~\P2_P1_InstAddrPointer_reg[30]/NET0131  & ~n31520 ;
  assign n31523 = ~n31521 & ~n31522 ;
  assign n31524 = \P2_P1_InstAddrPointer_reg[11]/NET0131  & n31509 ;
  assign n31525 = n31504 & n31524 ;
  assign n31526 = n31497 & n31525 ;
  assign n31527 = \P2_P1_InstAddrPointer_reg[21]/NET0131  & ~n31526 ;
  assign n31528 = ~\P2_P1_InstAddrPointer_reg[21]/NET0131  & ~n31500 ;
  assign n31529 = \P2_P1_InstAddrPointer_reg[21]/NET0131  & n31500 ;
  assign n31530 = ~n31528 & ~n31529 ;
  assign n31531 = n31526 & n31530 ;
  assign n31532 = ~n31527 & ~n31531 ;
  assign n31533 = n31502 & n31508 ;
  assign n31534 = ~\P2_P1_InstAddrPointer_reg[17]/NET0131  & ~n31533 ;
  assign n31535 = n31502 & n31509 ;
  assign n31536 = ~n31534 & ~n31535 ;
  assign n31537 = \P2_P1_InstAddrPointer_reg[11]/NET0131  & \P2_P1_InstAddrPointer_reg[12]/NET0131  ;
  assign n31538 = n31501 & n31537 ;
  assign n31539 = \P2_P1_InstAddrPointer_reg[13]/NET0131  & n31538 ;
  assign n31540 = ~\P2_P1_InstAddrPointer_reg[13]/NET0131  & ~n31538 ;
  assign n31541 = ~n31539 & ~n31540 ;
  assign n31542 = \P2_P1_InstAddrPointer_reg[5]/NET0131  & n31500 ;
  assign n31543 = \P2_P1_InstAddrPointer_reg[6]/NET0131  & n31542 ;
  assign n31544 = \P2_P1_InstAddrPointer_reg[7]/NET0131  & n31543 ;
  assign n31545 = ~\P2_P1_InstAddrPointer_reg[7]/NET0131  & ~n31543 ;
  assign n31546 = ~n31544 & ~n31545 ;
  assign n31547 = ~\P2_P1_InstAddrPointer_reg[6]/NET0131  & ~n31542 ;
  assign n31548 = ~n31543 & ~n31547 ;
  assign n31554 = \P2_P1_InstQueue_reg[7][6]/NET0131  & n11651 ;
  assign n31553 = \P2_P1_InstQueue_reg[0][6]/NET0131  & n11647 ;
  assign n31549 = \P2_P1_InstQueue_reg[2][6]/NET0131  & n11671 ;
  assign n31550 = \P2_P1_InstQueue_reg[4][6]/NET0131  & n11663 ;
  assign n31565 = ~n31549 & ~n31550 ;
  assign n31575 = ~n31553 & n31565 ;
  assign n31576 = ~n31554 & n31575 ;
  assign n31561 = \P2_P1_InstQueue_reg[1][6]/NET0131  & n11669 ;
  assign n31562 = \P2_P1_InstQueue_reg[6][6]/NET0131  & n11638 ;
  assign n31570 = ~n31561 & ~n31562 ;
  assign n31563 = \P2_P1_InstQueue_reg[10][6]/NET0131  & n11656 ;
  assign n31564 = \P2_P1_InstQueue_reg[3][6]/NET0131  & n11654 ;
  assign n31571 = ~n31563 & ~n31564 ;
  assign n31572 = n31570 & n31571 ;
  assign n31557 = \P2_P1_InstQueue_reg[11][6]/NET0131  & n11634 ;
  assign n31558 = \P2_P1_InstQueue_reg[8][6]/NET0131  & n11661 ;
  assign n31568 = ~n31557 & ~n31558 ;
  assign n31559 = \P2_P1_InstQueue_reg[5][6]/NET0131  & n11667 ;
  assign n31560 = \P2_P1_InstQueue_reg[12][6]/NET0131  & n11665 ;
  assign n31569 = ~n31559 & ~n31560 ;
  assign n31573 = n31568 & n31569 ;
  assign n31551 = \P2_P1_InstQueue_reg[14][6]/NET0131  & n11641 ;
  assign n31552 = \P2_P1_InstQueue_reg[15][6]/NET0131  & n11643 ;
  assign n31566 = ~n31551 & ~n31552 ;
  assign n31555 = \P2_P1_InstQueue_reg[9][6]/NET0131  & n11659 ;
  assign n31556 = \P2_P1_InstQueue_reg[13][6]/NET0131  & n11673 ;
  assign n31567 = ~n31555 & ~n31556 ;
  assign n31574 = n31566 & n31567 ;
  assign n31577 = n31573 & n31574 ;
  assign n31578 = n31572 & n31577 ;
  assign n31579 = n31576 & n31578 ;
  assign n31580 = n31548 & ~n31579 ;
  assign n31581 = ~n31548 & n31579 ;
  assign n31582 = ~\P2_P1_InstAddrPointer_reg[5]/NET0131  & ~n31500 ;
  assign n31583 = ~n31542 & ~n31582 ;
  assign n31589 = \P2_P1_InstQueue_reg[7][5]/NET0131  & n11651 ;
  assign n31588 = \P2_P1_InstQueue_reg[0][5]/NET0131  & n11647 ;
  assign n31584 = \P2_P1_InstQueue_reg[10][5]/NET0131  & n11656 ;
  assign n31585 = \P2_P1_InstQueue_reg[3][5]/NET0131  & n11654 ;
  assign n31600 = ~n31584 & ~n31585 ;
  assign n31610 = ~n31588 & n31600 ;
  assign n31611 = ~n31589 & n31610 ;
  assign n31596 = \P2_P1_InstQueue_reg[6][5]/NET0131  & n11638 ;
  assign n31597 = \P2_P1_InstQueue_reg[13][5]/NET0131  & n11673 ;
  assign n31605 = ~n31596 & ~n31597 ;
  assign n31598 = \P2_P1_InstQueue_reg[14][5]/NET0131  & n11641 ;
  assign n31599 = \P2_P1_InstQueue_reg[4][5]/NET0131  & n11663 ;
  assign n31606 = ~n31598 & ~n31599 ;
  assign n31607 = n31605 & n31606 ;
  assign n31592 = \P2_P1_InstQueue_reg[11][5]/NET0131  & n11634 ;
  assign n31593 = \P2_P1_InstQueue_reg[8][5]/NET0131  & n11661 ;
  assign n31603 = ~n31592 & ~n31593 ;
  assign n31594 = \P2_P1_InstQueue_reg[5][5]/NET0131  & n11667 ;
  assign n31595 = \P2_P1_InstQueue_reg[12][5]/NET0131  & n11665 ;
  assign n31604 = ~n31594 & ~n31595 ;
  assign n31608 = n31603 & n31604 ;
  assign n31586 = \P2_P1_InstQueue_reg[9][5]/NET0131  & n11659 ;
  assign n31587 = \P2_P1_InstQueue_reg[15][5]/NET0131  & n11643 ;
  assign n31601 = ~n31586 & ~n31587 ;
  assign n31590 = \P2_P1_InstQueue_reg[1][5]/NET0131  & n11669 ;
  assign n31591 = \P2_P1_InstQueue_reg[2][5]/NET0131  & n11671 ;
  assign n31602 = ~n31590 & ~n31591 ;
  assign n31609 = n31601 & n31602 ;
  assign n31612 = n31608 & n31609 ;
  assign n31613 = n31607 & n31612 ;
  assign n31614 = n31611 & n31613 ;
  assign n31615 = ~n31583 & n31614 ;
  assign n31616 = n31583 & ~n31614 ;
  assign n31617 = ~\P2_P1_InstAddrPointer_reg[4]/NET0131  & ~n31499 ;
  assign n31618 = ~n31500 & ~n31617 ;
  assign n31624 = \P2_P1_InstQueue_reg[7][4]/NET0131  & n11651 ;
  assign n31623 = \P2_P1_InstQueue_reg[0][4]/NET0131  & n11647 ;
  assign n31619 = \P2_P1_InstQueue_reg[12][4]/NET0131  & n11665 ;
  assign n31620 = \P2_P1_InstQueue_reg[2][4]/NET0131  & n11671 ;
  assign n31635 = ~n31619 & ~n31620 ;
  assign n31645 = ~n31623 & n31635 ;
  assign n31646 = ~n31624 & n31645 ;
  assign n31631 = \P2_P1_InstQueue_reg[5][4]/NET0131  & n11667 ;
  assign n31632 = \P2_P1_InstQueue_reg[14][4]/NET0131  & n11641 ;
  assign n31640 = ~n31631 & ~n31632 ;
  assign n31633 = \P2_P1_InstQueue_reg[1][4]/NET0131  & n11669 ;
  assign n31634 = \P2_P1_InstQueue_reg[9][4]/NET0131  & n11659 ;
  assign n31641 = ~n31633 & ~n31634 ;
  assign n31642 = n31640 & n31641 ;
  assign n31627 = \P2_P1_InstQueue_reg[10][4]/NET0131  & n11656 ;
  assign n31628 = \P2_P1_InstQueue_reg[8][4]/NET0131  & n11661 ;
  assign n31638 = ~n31627 & ~n31628 ;
  assign n31629 = \P2_P1_InstQueue_reg[11][4]/NET0131  & n11634 ;
  assign n31630 = \P2_P1_InstQueue_reg[3][4]/NET0131  & n11654 ;
  assign n31639 = ~n31629 & ~n31630 ;
  assign n31643 = n31638 & n31639 ;
  assign n31621 = \P2_P1_InstQueue_reg[4][4]/NET0131  & n11663 ;
  assign n31622 = \P2_P1_InstQueue_reg[15][4]/NET0131  & n11643 ;
  assign n31636 = ~n31621 & ~n31622 ;
  assign n31625 = \P2_P1_InstQueue_reg[13][4]/NET0131  & n11673 ;
  assign n31626 = \P2_P1_InstQueue_reg[6][4]/NET0131  & n11638 ;
  assign n31637 = ~n31625 & ~n31626 ;
  assign n31644 = n31636 & n31637 ;
  assign n31647 = n31643 & n31644 ;
  assign n31648 = n31642 & n31647 ;
  assign n31649 = n31646 & n31648 ;
  assign n31650 = n31618 & ~n31649 ;
  assign n31651 = ~n31618 & n31649 ;
  assign n31652 = ~\P2_P1_InstAddrPointer_reg[3]/NET0131  & ~n31498 ;
  assign n31653 = ~n31499 & ~n31652 ;
  assign n31659 = \P2_P1_InstQueue_reg[7][3]/NET0131  & n11651 ;
  assign n31658 = \P2_P1_InstQueue_reg[0][3]/NET0131  & n11647 ;
  assign n31654 = \P2_P1_InstQueue_reg[4][3]/NET0131  & n11663 ;
  assign n31655 = \P2_P1_InstQueue_reg[2][3]/NET0131  & n11671 ;
  assign n31670 = ~n31654 & ~n31655 ;
  assign n31680 = ~n31658 & n31670 ;
  assign n31681 = ~n31659 & n31680 ;
  assign n31666 = \P2_P1_InstQueue_reg[12][3]/NET0131  & n11665 ;
  assign n31667 = \P2_P1_InstQueue_reg[13][3]/NET0131  & n11673 ;
  assign n31675 = ~n31666 & ~n31667 ;
  assign n31668 = \P2_P1_InstQueue_reg[5][3]/NET0131  & n11667 ;
  assign n31669 = \P2_P1_InstQueue_reg[11][3]/NET0131  & n11634 ;
  assign n31676 = ~n31668 & ~n31669 ;
  assign n31677 = n31675 & n31676 ;
  assign n31662 = \P2_P1_InstQueue_reg[14][3]/NET0131  & n11641 ;
  assign n31663 = \P2_P1_InstQueue_reg[8][3]/NET0131  & n11661 ;
  assign n31673 = ~n31662 & ~n31663 ;
  assign n31664 = \P2_P1_InstQueue_reg[6][3]/NET0131  & n11638 ;
  assign n31665 = \P2_P1_InstQueue_reg[1][3]/NET0131  & n11669 ;
  assign n31674 = ~n31664 & ~n31665 ;
  assign n31678 = n31673 & n31674 ;
  assign n31656 = \P2_P1_InstQueue_reg[3][3]/NET0131  & n11654 ;
  assign n31657 = \P2_P1_InstQueue_reg[15][3]/NET0131  & n11643 ;
  assign n31671 = ~n31656 & ~n31657 ;
  assign n31660 = \P2_P1_InstQueue_reg[10][3]/NET0131  & n11656 ;
  assign n31661 = \P2_P1_InstQueue_reg[9][3]/NET0131  & n11659 ;
  assign n31672 = ~n31660 & ~n31661 ;
  assign n31679 = n31671 & n31672 ;
  assign n31682 = n31678 & n31679 ;
  assign n31683 = n31677 & n31682 ;
  assign n31684 = n31681 & n31683 ;
  assign n31685 = n31653 & ~n31684 ;
  assign n31686 = ~n31653 & n31684 ;
  assign n31687 = ~\P2_P1_InstAddrPointer_reg[1]/NET0131  & ~\P2_P1_InstAddrPointer_reg[2]/NET0131  ;
  assign n31688 = ~n31498 & ~n31687 ;
  assign n31696 = \P2_P1_InstQueue_reg[7][2]/NET0131  & n11651 ;
  assign n31691 = \P2_P1_InstQueue_reg[0][2]/NET0131  & n11647 ;
  assign n31689 = \P2_P1_InstQueue_reg[2][2]/NET0131  & n11671 ;
  assign n31690 = \P2_P1_InstQueue_reg[12][2]/NET0131  & n11665 ;
  assign n31705 = ~n31689 & ~n31690 ;
  assign n31715 = ~n31691 & n31705 ;
  assign n31716 = ~n31696 & n31715 ;
  assign n31701 = \P2_P1_InstQueue_reg[3][2]/NET0131  & n11654 ;
  assign n31702 = \P2_P1_InstQueue_reg[4][2]/NET0131  & n11663 ;
  assign n31710 = ~n31701 & ~n31702 ;
  assign n31703 = \P2_P1_InstQueue_reg[14][2]/NET0131  & n11641 ;
  assign n31704 = \P2_P1_InstQueue_reg[5][2]/NET0131  & n11667 ;
  assign n31711 = ~n31703 & ~n31704 ;
  assign n31712 = n31710 & n31711 ;
  assign n31697 = \P2_P1_InstQueue_reg[10][2]/NET0131  & n11656 ;
  assign n31698 = \P2_P1_InstQueue_reg[9][2]/NET0131  & n11659 ;
  assign n31708 = ~n31697 & ~n31698 ;
  assign n31699 = \P2_P1_InstQueue_reg[8][2]/NET0131  & n11661 ;
  assign n31700 = \P2_P1_InstQueue_reg[11][2]/NET0131  & n11634 ;
  assign n31709 = ~n31699 & ~n31700 ;
  assign n31713 = n31708 & n31709 ;
  assign n31692 = \P2_P1_InstQueue_reg[6][2]/NET0131  & n11638 ;
  assign n31693 = \P2_P1_InstQueue_reg[15][2]/NET0131  & n11643 ;
  assign n31706 = ~n31692 & ~n31693 ;
  assign n31694 = \P2_P1_InstQueue_reg[13][2]/NET0131  & n11673 ;
  assign n31695 = \P2_P1_InstQueue_reg[1][2]/NET0131  & n11669 ;
  assign n31707 = ~n31694 & ~n31695 ;
  assign n31714 = n31706 & n31707 ;
  assign n31717 = n31713 & n31714 ;
  assign n31718 = n31712 & n31717 ;
  assign n31719 = n31716 & n31718 ;
  assign n31720 = n31688 & ~n31719 ;
  assign n31721 = ~n31688 & n31719 ;
  assign n31734 = \P2_P1_InstQueue_reg[7][1]/NET0131  & n11651 ;
  assign n31722 = \P2_P1_InstQueue_reg[0][1]/NET0131  & n11647 ;
  assign n31723 = \P2_P1_InstQueue_reg[14][1]/NET0131  & n11641 ;
  assign n31724 = \P2_P1_InstQueue_reg[9][1]/NET0131  & n11659 ;
  assign n31738 = ~n31723 & ~n31724 ;
  assign n31748 = ~n31722 & n31738 ;
  assign n31749 = ~n31734 & n31748 ;
  assign n31733 = \P2_P1_InstQueue_reg[8][1]/NET0131  & n11661 ;
  assign n31735 = \P2_P1_InstQueue_reg[6][1]/NET0131  & n11638 ;
  assign n31743 = ~n31733 & ~n31735 ;
  assign n31736 = \P2_P1_InstQueue_reg[4][1]/NET0131  & n11663 ;
  assign n31737 = \P2_P1_InstQueue_reg[3][1]/NET0131  & n11654 ;
  assign n31744 = ~n31736 & ~n31737 ;
  assign n31745 = n31743 & n31744 ;
  assign n31729 = \P2_P1_InstQueue_reg[5][1]/NET0131  & n11667 ;
  assign n31730 = \P2_P1_InstQueue_reg[11][1]/NET0131  & n11634 ;
  assign n31741 = ~n31729 & ~n31730 ;
  assign n31731 = \P2_P1_InstQueue_reg[1][1]/NET0131  & n11669 ;
  assign n31732 = \P2_P1_InstQueue_reg[10][1]/NET0131  & n11656 ;
  assign n31742 = ~n31731 & ~n31732 ;
  assign n31746 = n31741 & n31742 ;
  assign n31725 = \P2_P1_InstQueue_reg[2][1]/NET0131  & n11671 ;
  assign n31726 = \P2_P1_InstQueue_reg[15][1]/NET0131  & n11643 ;
  assign n31739 = ~n31725 & ~n31726 ;
  assign n31727 = \P2_P1_InstQueue_reg[13][1]/NET0131  & n11673 ;
  assign n31728 = \P2_P1_InstQueue_reg[12][1]/NET0131  & n11665 ;
  assign n31740 = ~n31727 & ~n31728 ;
  assign n31747 = n31739 & n31740 ;
  assign n31750 = n31746 & n31747 ;
  assign n31751 = n31745 & n31750 ;
  assign n31752 = n31749 & n31751 ;
  assign n31753 = ~\P2_P1_InstAddrPointer_reg[1]/NET0131  & ~n31752 ;
  assign n31754 = \P2_P1_InstAddrPointer_reg[1]/NET0131  & n31752 ;
  assign n31767 = \P2_P1_InstQueue_reg[7][0]/NET0131  & n11651 ;
  assign n31755 = \P2_P1_InstQueue_reg[0][0]/NET0131  & n11647 ;
  assign n31756 = \P2_P1_InstQueue_reg[14][0]/NET0131  & n11641 ;
  assign n31757 = \P2_P1_InstQueue_reg[9][0]/NET0131  & n11659 ;
  assign n31771 = ~n31756 & ~n31757 ;
  assign n31781 = ~n31755 & n31771 ;
  assign n31782 = ~n31767 & n31781 ;
  assign n31766 = \P2_P1_InstQueue_reg[8][0]/NET0131  & n11661 ;
  assign n31768 = \P2_P1_InstQueue_reg[6][0]/NET0131  & n11638 ;
  assign n31776 = ~n31766 & ~n31768 ;
  assign n31769 = \P2_P1_InstQueue_reg[4][0]/NET0131  & n11663 ;
  assign n31770 = \P2_P1_InstQueue_reg[3][0]/NET0131  & n11654 ;
  assign n31777 = ~n31769 & ~n31770 ;
  assign n31778 = n31776 & n31777 ;
  assign n31762 = \P2_P1_InstQueue_reg[2][0]/NET0131  & n11671 ;
  assign n31763 = \P2_P1_InstQueue_reg[11][0]/NET0131  & n11634 ;
  assign n31774 = ~n31762 & ~n31763 ;
  assign n31764 = \P2_P1_InstQueue_reg[5][0]/NET0131  & n11667 ;
  assign n31765 = \P2_P1_InstQueue_reg[10][0]/NET0131  & n11656 ;
  assign n31775 = ~n31764 & ~n31765 ;
  assign n31779 = n31774 & n31775 ;
  assign n31758 = \P2_P1_InstQueue_reg[1][0]/NET0131  & n11669 ;
  assign n31759 = \P2_P1_InstQueue_reg[15][0]/NET0131  & n11643 ;
  assign n31772 = ~n31758 & ~n31759 ;
  assign n31760 = \P2_P1_InstQueue_reg[13][0]/NET0131  & n11673 ;
  assign n31761 = \P2_P1_InstQueue_reg[12][0]/NET0131  & n11665 ;
  assign n31773 = ~n31760 & ~n31761 ;
  assign n31780 = n31772 & n31773 ;
  assign n31783 = n31779 & n31780 ;
  assign n31784 = n31778 & n31783 ;
  assign n31785 = n31782 & n31784 ;
  assign n31786 = \P2_P1_InstAddrPointer_reg[0]/NET0131  & ~n31785 ;
  assign n31787 = ~n31754 & n31786 ;
  assign n31788 = ~n31753 & ~n31787 ;
  assign n31789 = ~n31721 & ~n31788 ;
  assign n31790 = ~n31720 & ~n31789 ;
  assign n31791 = ~n31686 & ~n31790 ;
  assign n31792 = ~n31685 & ~n31791 ;
  assign n31793 = ~n31651 & ~n31792 ;
  assign n31794 = ~n31650 & ~n31793 ;
  assign n31795 = ~n31616 & n31794 ;
  assign n31796 = ~n31615 & ~n31795 ;
  assign n31797 = ~n31581 & n31796 ;
  assign n31798 = ~n31580 & ~n31797 ;
  assign n31799 = n31546 & ~n31798 ;
  assign n31800 = n29503 & ~n31799 ;
  assign n31801 = ~\P2_P1_InstAddrPointer_reg[8]/NET0131  & ~n31544 ;
  assign n31802 = n31493 & n31543 ;
  assign n31803 = ~n31801 & ~n31802 ;
  assign n31804 = ~n31546 & n31798 ;
  assign n31805 = n31803 & ~n31804 ;
  assign n31806 = ~n31800 & n31805 ;
  assign n31807 = \P2_P1_InstAddrPointer_reg[9]/NET0131  & n31806 ;
  assign n31808 = \P2_P1_InstAddrPointer_reg[9]/NET0131  & n31802 ;
  assign n31809 = ~\P2_P1_InstAddrPointer_reg[10]/NET0131  & ~n31808 ;
  assign n31810 = ~n31501 & ~n31809 ;
  assign n31811 = n31807 & n31810 ;
  assign n31812 = n31537 & n31811 ;
  assign n31813 = n31541 & n31812 ;
  assign n31814 = \P2_P1_InstAddrPointer_reg[14]/NET0131  & n31813 ;
  assign n31815 = n31502 & n31506 ;
  assign n31816 = \P2_P1_InstAddrPointer_reg[15]/NET0131  & ~n31815 ;
  assign n31817 = ~\P2_P1_InstAddrPointer_reg[15]/NET0131  & n31815 ;
  assign n31818 = ~n31816 & ~n31817 ;
  assign n31819 = n31814 & ~n31818 ;
  assign n31820 = \P2_P1_InstAddrPointer_reg[16]/NET0131  & ~n31502 ;
  assign n31821 = ~\P2_P1_InstAddrPointer_reg[16]/NET0131  & ~n31507 ;
  assign n31822 = ~n31508 & ~n31821 ;
  assign n31823 = n31502 & n31822 ;
  assign n31824 = ~n31820 & ~n31823 ;
  assign n31825 = n31819 & ~n31824 ;
  assign n31826 = n31536 & n31825 ;
  assign n31827 = \P2_P1_InstAddrPointer_reg[18]/NET0131  & n31524 ;
  assign n31828 = \P2_P1_InstAddrPointer_reg[19]/NET0131  & n31495 ;
  assign n31829 = n31543 & n31828 ;
  assign n31830 = n31827 & n31829 ;
  assign n31831 = ~\P2_P1_InstAddrPointer_reg[20]/NET0131  & ~n31830 ;
  assign n31832 = \P2_P1_InstAddrPointer_reg[20]/NET0131  & n31830 ;
  assign n31833 = ~n31831 & ~n31832 ;
  assign n31834 = n31501 & n31827 ;
  assign n31835 = \P2_P1_InstAddrPointer_reg[19]/NET0131  & ~n31834 ;
  assign n31836 = ~\P2_P1_InstAddrPointer_reg[18]/NET0131  & ~n31535 ;
  assign n31837 = n31835 & ~n31836 ;
  assign n31838 = n31833 & n31837 ;
  assign n31839 = n31826 & n31838 ;
  assign n31840 = ~n31532 & n31839 ;
  assign n31841 = \P2_P1_InstAddrPointer_reg[21]/NET0131  & n31496 ;
  assign n31842 = n31525 & n31841 ;
  assign n31843 = ~\P2_P1_InstAddrPointer_reg[22]/NET0131  & n31842 ;
  assign n31844 = \P2_P1_InstAddrPointer_reg[22]/NET0131  & ~n31842 ;
  assign n31845 = ~n31843 & ~n31844 ;
  assign n31846 = n31542 & ~n31845 ;
  assign n31847 = \P2_P1_InstAddrPointer_reg[22]/NET0131  & ~n31542 ;
  assign n31848 = ~n31846 & ~n31847 ;
  assign n31849 = n31840 & ~n31848 ;
  assign n31850 = ~\P2_P1_InstAddrPointer_reg[23]/NET0131  & ~n31513 ;
  assign n31851 = ~n31514 & ~n31850 ;
  assign n31852 = n31849 & n31851 ;
  assign n31853 = \P2_P1_InstAddrPointer_reg[24]/NET0131  & n31852 ;
  assign n31854 = ~\P2_P1_InstAddrPointer_reg[25]/NET0131  & ~n31515 ;
  assign n31855 = ~n31516 & ~n31854 ;
  assign n31856 = \P2_P1_InstAddrPointer_reg[26]/NET0131  & n31855 ;
  assign n31857 = n31853 & n31856 ;
  assign n31858 = ~\P2_P1_InstAddrPointer_reg[27]/NET0131  & ~n31517 ;
  assign n31859 = ~n31518 & ~n31858 ;
  assign n31860 = \P2_P1_InstAddrPointer_reg[28]/NET0131  & \P2_P1_InstAddrPointer_reg[29]/NET0131  ;
  assign n31861 = n31859 & n31860 ;
  assign n31862 = n31857 & n31861 ;
  assign n31863 = n31523 & n31862 ;
  assign n31868 = ~\P2_P1_InstAddrPointer_reg[31]/NET0131  & n31863 ;
  assign n31864 = ~\P2_P1_InstAddrPointer_reg[31]/NET0131  & ~n31521 ;
  assign n31865 = \P2_P1_InstAddrPointer_reg[31]/NET0131  & n31521 ;
  assign n31866 = ~n31864 & ~n31865 ;
  assign n31867 = ~n31863 & n31866 ;
  assign n31869 = n29503 & ~n31867 ;
  assign n31870 = ~n31868 & n31869 ;
  assign n31872 = \P2_P1_InstAddrPointer_reg[0]/NET0131  & \P2_P1_InstAddrPointer_reg[1]/NET0131  ;
  assign n31873 = \P2_P1_InstAddrPointer_reg[2]/NET0131  & n31872 ;
  assign n31874 = \P2_P1_InstAddrPointer_reg[3]/NET0131  & n31873 ;
  assign n31875 = \P2_P1_InstAddrPointer_reg[4]/NET0131  & \P2_P1_InstAddrPointer_reg[5]/NET0131  ;
  assign n31876 = n31874 & n31875 ;
  assign n31886 = \P2_P1_InstAddrPointer_reg[6]/NET0131  & n31876 ;
  assign n31887 = \P2_P1_InstAddrPointer_reg[7]/NET0131  & n31886 ;
  assign n31888 = ~\P2_P1_InstAddrPointer_reg[8]/NET0131  & ~n31887 ;
  assign n31889 = n31493 & n31886 ;
  assign n31890 = ~n31888 & ~n31889 ;
  assign n31891 = ~\P2_P1_InstAddrPointer_reg[7]/NET0131  & ~n31886 ;
  assign n31892 = ~n31887 & ~n31891 ;
  assign n31893 = n29503 & ~n31892 ;
  assign n31894 = ~n29503 & n31892 ;
  assign n31895 = ~\P2_P1_InstAddrPointer_reg[6]/NET0131  & ~n31876 ;
  assign n31896 = ~n31886 & ~n31895 ;
  assign n31897 = n31579 & ~n31896 ;
  assign n31898 = ~n31579 & n31896 ;
  assign n31899 = \P2_P1_InstAddrPointer_reg[4]/NET0131  & n31874 ;
  assign n31900 = ~\P2_P1_InstAddrPointer_reg[5]/NET0131  & ~n31899 ;
  assign n31901 = ~n31876 & ~n31900 ;
  assign n31902 = n31614 & ~n31901 ;
  assign n31903 = ~n31614 & n31901 ;
  assign n31904 = ~\P2_P1_InstAddrPointer_reg[4]/NET0131  & ~n31874 ;
  assign n31905 = ~n31899 & ~n31904 ;
  assign n31906 = ~n31649 & n31905 ;
  assign n31907 = n31649 & ~n31905 ;
  assign n31908 = ~\P2_P1_InstAddrPointer_reg[3]/NET0131  & ~n31873 ;
  assign n31909 = ~n31874 & ~n31908 ;
  assign n31910 = ~n31684 & n31909 ;
  assign n31911 = n31684 & ~n31909 ;
  assign n31912 = ~\P2_P1_InstAddrPointer_reg[2]/NET0131  & ~n31872 ;
  assign n31913 = ~n31873 & ~n31912 ;
  assign n31914 = ~n31719 & n31913 ;
  assign n31915 = n31719 & ~n31913 ;
  assign n31916 = ~\P2_P1_InstAddrPointer_reg[0]/NET0131  & \P2_P1_InstAddrPointer_reg[1]/NET0131  ;
  assign n31917 = n31788 & ~n31916 ;
  assign n31918 = ~n31915 & ~n31917 ;
  assign n31919 = ~n31914 & ~n31918 ;
  assign n31920 = ~n31911 & ~n31919 ;
  assign n31921 = ~n31910 & ~n31920 ;
  assign n31922 = ~n31907 & ~n31921 ;
  assign n31923 = ~n31906 & ~n31922 ;
  assign n31924 = ~n31903 & n31923 ;
  assign n31925 = ~n31902 & ~n31924 ;
  assign n31926 = ~n31898 & ~n31925 ;
  assign n31927 = ~n31897 & ~n31926 ;
  assign n31928 = ~n31894 & ~n31927 ;
  assign n31929 = ~n31893 & ~n31928 ;
  assign n31930 = ~n31890 & ~n31929 ;
  assign n31931 = ~\P2_P1_InstAddrPointer_reg[9]/NET0131  & ~n31889 ;
  assign n31932 = \P2_P1_InstAddrPointer_reg[0]/NET0131  & n31808 ;
  assign n31933 = ~n31931 & ~n31932 ;
  assign n31934 = n31930 & ~n31933 ;
  assign n31877 = n31496 & n31876 ;
  assign n31935 = ~\P2_P1_InstAddrPointer_reg[10]/NET0131  & ~n31932 ;
  assign n31936 = ~n31877 & ~n31935 ;
  assign n31937 = n31934 & ~n31936 ;
  assign n31878 = \P2_P1_InstAddrPointer_reg[11]/NET0131  & n31877 ;
  assign n31938 = ~\P2_P1_InstAddrPointer_reg[11]/NET0131  & ~n31877 ;
  assign n31939 = ~n31878 & ~n31938 ;
  assign n31940 = n31937 & ~n31939 ;
  assign n31941 = ~\P2_P1_InstAddrPointer_reg[12]/NET0131  & ~n31878 ;
  assign n31942 = \P2_P1_InstAddrPointer_reg[0]/NET0131  & n31538 ;
  assign n31943 = ~n31941 & ~n31942 ;
  assign n31944 = n31940 & ~n31943 ;
  assign n31945 = \P2_P1_InstAddrPointer_reg[0]/NET0131  & n31539 ;
  assign n31947 = \P2_P1_InstAddrPointer_reg[14]/NET0131  & n31945 ;
  assign n31954 = ~\P2_P1_InstAddrPointer_reg[15]/NET0131  & ~n31947 ;
  assign n31955 = \P2_P1_InstAddrPointer_reg[15]/NET0131  & n31947 ;
  assign n31956 = ~n31954 & ~n31955 ;
  assign n31946 = ~\P2_P1_InstAddrPointer_reg[14]/NET0131  & ~n31945 ;
  assign n31948 = ~n31946 & ~n31947 ;
  assign n31949 = ~\P2_P1_InstAddrPointer_reg[13]/NET0131  & ~n31942 ;
  assign n31950 = ~n31945 & ~n31949 ;
  assign n31951 = \P2_P1_InstAddrPointer_reg[16]/NET0131  & ~n31878 ;
  assign n31952 = n31822 & n31878 ;
  assign n31953 = ~n31951 & ~n31952 ;
  assign n31957 = ~n31950 & n31953 ;
  assign n31958 = ~n31948 & n31957 ;
  assign n31959 = ~n31956 & n31958 ;
  assign n31960 = n31944 & n31959 ;
  assign n31965 = \P2_P1_InstAddrPointer_reg[16]/NET0131  & n31955 ;
  assign n31966 = \P2_P1_InstAddrPointer_reg[17]/NET0131  & ~n31965 ;
  assign n31967 = ~\P2_P1_InstAddrPointer_reg[17]/NET0131  & n31965 ;
  assign n31968 = ~n31966 & ~n31967 ;
  assign n31961 = \P2_P1_InstAddrPointer_reg[0]/NET0131  & n31526 ;
  assign n31962 = \P2_P1_InstAddrPointer_reg[21]/NET0131  & ~n31961 ;
  assign n31963 = \P2_P1_InstAddrPointer_reg[0]/NET0131  & n31531 ;
  assign n31964 = ~n31962 & ~n31963 ;
  assign n31969 = n31827 & n31877 ;
  assign n31970 = \P2_P1_InstAddrPointer_reg[19]/NET0131  & n31969 ;
  assign n31976 = ~\P2_P1_InstAddrPointer_reg[20]/NET0131  & ~n31970 ;
  assign n31977 = \P2_P1_InstAddrPointer_reg[20]/NET0131  & n31970 ;
  assign n31978 = ~n31976 & ~n31977 ;
  assign n31971 = ~\P2_P1_InstAddrPointer_reg[19]/NET0131  & ~n31969 ;
  assign n31972 = ~n31970 & ~n31971 ;
  assign n31973 = \P2_P1_InstAddrPointer_reg[0]/NET0131  & n31535 ;
  assign n31974 = ~\P2_P1_InstAddrPointer_reg[18]/NET0131  & ~n31973 ;
  assign n31975 = ~n31969 & ~n31974 ;
  assign n31979 = ~n31972 & ~n31975 ;
  assign n31980 = ~n31978 & n31979 ;
  assign n31981 = n31964 & n31980 ;
  assign n31982 = n31968 & n31981 ;
  assign n31983 = n31960 & n31982 ;
  assign n31871 = \P2_P1_InstAddrPointer_reg[23]/NET0131  & n31512 ;
  assign n31879 = n31871 & n31878 ;
  assign n31880 = \P2_P1_InstAddrPointer_reg[0]/NET0131  & n31513 ;
  assign n31881 = ~\P2_P1_InstAddrPointer_reg[23]/NET0131  & ~n31880 ;
  assign n31882 = ~n31879 & ~n31881 ;
  assign n31883 = \P2_P1_InstAddrPointer_reg[22]/NET0131  & ~n31876 ;
  assign n31884 = \P2_P1_InstAddrPointer_reg[0]/NET0131  & n31846 ;
  assign n31885 = ~n31883 & ~n31884 ;
  assign n31984 = ~n31882 & n31885 ;
  assign n31985 = n31983 & n31984 ;
  assign n31986 = ~\P2_P1_InstAddrPointer_reg[24]/NET0131  & ~n31879 ;
  assign n31987 = \P2_P1_InstAddrPointer_reg[0]/NET0131  & n31515 ;
  assign n31988 = ~n31986 & ~n31987 ;
  assign n31989 = n31985 & ~n31988 ;
  assign n31990 = ~\P2_P1_InstAddrPointer_reg[25]/NET0131  & ~n31987 ;
  assign n31991 = \P2_P1_InstAddrPointer_reg[25]/NET0131  & n31987 ;
  assign n31992 = ~n31990 & ~n31991 ;
  assign n31993 = n31989 & ~n31992 ;
  assign n31994 = ~\P2_P1_InstAddrPointer_reg[26]/NET0131  & ~n31991 ;
  assign n31995 = \P2_P1_InstAddrPointer_reg[26]/NET0131  & n31991 ;
  assign n31996 = ~n31994 & ~n31995 ;
  assign n31997 = n31993 & ~n31996 ;
  assign n31998 = ~\P2_P1_InstAddrPointer_reg[27]/NET0131  & ~n31995 ;
  assign n31999 = \P2_P1_InstAddrPointer_reg[0]/NET0131  & n31518 ;
  assign n32000 = ~n31998 & ~n31999 ;
  assign n32001 = n31997 & ~n32000 ;
  assign n32002 = ~\P2_P1_InstAddrPointer_reg[28]/NET0131  & ~n31999 ;
  assign n32003 = \P2_P1_InstAddrPointer_reg[0]/NET0131  & n31519 ;
  assign n32004 = ~n32002 & ~n32003 ;
  assign n32005 = n32001 & ~n32004 ;
  assign n32006 = ~\P2_P1_InstAddrPointer_reg[29]/NET0131  & ~n32003 ;
  assign n32007 = \P2_P1_InstAddrPointer_reg[29]/NET0131  & n32003 ;
  assign n32008 = ~n32006 & ~n32007 ;
  assign n32009 = n32005 & ~n32008 ;
  assign n32010 = ~\P2_P1_InstAddrPointer_reg[30]/NET0131  & ~n32007 ;
  assign n32011 = \P2_P1_InstAddrPointer_reg[30]/NET0131  & n32007 ;
  assign n32012 = ~n32010 & ~n32011 ;
  assign n32013 = n32009 & ~n32012 ;
  assign n32014 = \P2_P1_InstAddrPointer_reg[31]/NET0131  & ~n32011 ;
  assign n32015 = ~\P2_P1_InstAddrPointer_reg[31]/NET0131  & n32011 ;
  assign n32016 = ~n32014 & ~n32015 ;
  assign n32018 = n32013 & n32016 ;
  assign n32017 = ~n32013 & ~n32016 ;
  assign n32019 = ~n29503 & ~n32017 ;
  assign n32020 = ~n32018 & n32019 ;
  assign n32021 = ~n25947 & ~n32020 ;
  assign n32022 = ~n31870 & n32021 ;
  assign n32023 = ~n31492 & ~n32022 ;
  assign n32024 = n25945 & ~n32023 ;
  assign n32030 = \P2_P1_InstAddrPointer_reg[3]/NET0131  & ~n31912 ;
  assign n32031 = \P2_P1_InstAddrPointer_reg[4]/NET0131  & n32030 ;
  assign n32032 = n31526 & n32031 ;
  assign n32033 = \P2_P1_InstAddrPointer_reg[21]/NET0131  & n32032 ;
  assign n32034 = \P2_P1_InstAddrPointer_reg[22]/NET0131  & n32033 ;
  assign n32035 = \P2_P1_InstAddrPointer_reg[23]/NET0131  & n32034 ;
  assign n32036 = \P2_P1_InstAddrPointer_reg[24]/NET0131  & n32035 ;
  assign n32037 = \P2_P1_InstAddrPointer_reg[25]/NET0131  & n32036 ;
  assign n32038 = \P2_P1_InstAddrPointer_reg[26]/NET0131  & n32037 ;
  assign n32039 = \P2_P1_InstAddrPointer_reg[27]/NET0131  & n32038 ;
  assign n32040 = \P2_P1_InstAddrPointer_reg[28]/NET0131  & n32039 ;
  assign n32041 = ~\P2_P1_InstAddrPointer_reg[28]/NET0131  & ~n32039 ;
  assign n32042 = ~n32040 & ~n32041 ;
  assign n32043 = ~\P2_P1_InstAddrPointer_reg[25]/NET0131  & ~n32036 ;
  assign n32044 = ~n32037 & ~n32043 ;
  assign n32045 = \P2_P1_InstAddrPointer_reg[5]/NET0131  & n32031 ;
  assign n32046 = \P2_P1_InstAddrPointer_reg[6]/NET0131  & n32045 ;
  assign n32047 = \P2_P1_InstAddrPointer_reg[7]/NET0131  & n32046 ;
  assign n32048 = \P2_P1_InstAddrPointer_reg[8]/NET0131  & n32047 ;
  assign n32049 = \P2_P1_InstAddrPointer_reg[9]/NET0131  & n32048 ;
  assign n32050 = \P2_P1_InstAddrPointer_reg[10]/NET0131  & n32049 ;
  assign n32051 = n31537 & n32050 ;
  assign n32052 = \P2_P1_InstAddrPointer_reg[13]/NET0131  & n32051 ;
  assign n32053 = ~\P2_P1_InstAddrPointer_reg[13]/NET0131  & ~n32051 ;
  assign n32054 = ~n32052 & ~n32053 ;
  assign n32055 = \P2_P1_InstAddrPointer_reg[11]/NET0131  & n32050 ;
  assign n32056 = ~\P2_P1_InstAddrPointer_reg[11]/NET0131  & ~n32050 ;
  assign n32057 = ~n32055 & ~n32056 ;
  assign n32058 = ~\P2_P1_InstAddrPointer_reg[8]/NET0131  & ~n32047 ;
  assign n32059 = ~n32048 & ~n32058 ;
  assign n32060 = ~\P2_P1_InstAddrPointer_reg[7]/NET0131  & ~n32046 ;
  assign n32061 = ~n32047 & ~n32060 ;
  assign n32062 = ~n29503 & n32061 ;
  assign n32063 = n29503 & ~n32061 ;
  assign n32064 = ~\P2_P1_InstAddrPointer_reg[6]/NET0131  & ~n32045 ;
  assign n32065 = ~n32046 & ~n32064 ;
  assign n32066 = ~n31579 & n32065 ;
  assign n32067 = n31579 & ~n32065 ;
  assign n32068 = ~\P2_P1_InstAddrPointer_reg[5]/NET0131  & ~n32031 ;
  assign n32069 = ~n32045 & ~n32068 ;
  assign n32070 = ~n31614 & n32069 ;
  assign n32071 = n31614 & ~n32069 ;
  assign n32072 = ~\P2_P1_InstAddrPointer_reg[4]/NET0131  & ~n32030 ;
  assign n32073 = ~n32031 & ~n32072 ;
  assign n32074 = ~n31649 & n32073 ;
  assign n32075 = n31649 & ~n32073 ;
  assign n32076 = ~\P2_P1_InstAddrPointer_reg[3]/NET0131  & n31912 ;
  assign n32077 = ~n32030 & ~n32076 ;
  assign n32078 = ~n31684 & n32077 ;
  assign n32079 = n31684 & ~n32077 ;
  assign n32080 = ~n31719 & ~n31913 ;
  assign n32081 = n31719 & n31913 ;
  assign n32082 = \P2_P1_InstAddrPointer_reg[0]/NET0131  & ~\P2_P1_InstAddrPointer_reg[1]/NET0131  ;
  assign n32083 = ~n31916 & ~n32082 ;
  assign n32084 = ~n31752 & ~n32083 ;
  assign n32085 = n31752 & n32083 ;
  assign n32086 = ~\P2_P1_InstAddrPointer_reg[0]/NET0131  & ~n31785 ;
  assign n32087 = ~n32085 & n32086 ;
  assign n32088 = ~n32084 & ~n32087 ;
  assign n32089 = ~n32081 & ~n32088 ;
  assign n32090 = ~n32080 & ~n32089 ;
  assign n32091 = ~n32079 & ~n32090 ;
  assign n32092 = ~n32078 & ~n32091 ;
  assign n32093 = ~n32075 & ~n32092 ;
  assign n32094 = ~n32074 & ~n32093 ;
  assign n32095 = ~n32071 & ~n32094 ;
  assign n32096 = ~n32070 & ~n32095 ;
  assign n32097 = ~n32067 & ~n32096 ;
  assign n32098 = ~n32066 & ~n32097 ;
  assign n32099 = ~n32063 & ~n32098 ;
  assign n32100 = ~n32062 & ~n32099 ;
  assign n32101 = n32059 & ~n32100 ;
  assign n32102 = \P2_P1_InstAddrPointer_reg[9]/NET0131  & n32101 ;
  assign n32103 = \P2_P1_InstAddrPointer_reg[10]/NET0131  & n32102 ;
  assign n32104 = n32057 & n32103 ;
  assign n32105 = \P2_P1_InstAddrPointer_reg[12]/NET0131  & n32104 ;
  assign n32106 = n32054 & n32105 ;
  assign n32107 = \P2_P1_InstAddrPointer_reg[15]/NET0131  & \P2_P1_InstAddrPointer_reg[16]/NET0131  ;
  assign n32108 = ~\P2_P1_InstAddrPointer_reg[14]/NET0131  & ~n32052 ;
  assign n32109 = n31505 & n32051 ;
  assign n32110 = ~n32108 & ~n32109 ;
  assign n32111 = n32107 & n32110 ;
  assign n32112 = n32106 & n32111 ;
  assign n32113 = n32107 & n32109 ;
  assign n32114 = ~\P2_P1_InstAddrPointer_reg[17]/NET0131  & ~n32113 ;
  assign n32115 = n31524 & n32050 ;
  assign n32116 = ~n32114 & ~n32115 ;
  assign n32117 = n32112 & n32116 ;
  assign n32121 = n31503 & n32115 ;
  assign n32122 = ~\P2_P1_InstAddrPointer_reg[20]/NET0131  & ~n32121 ;
  assign n32123 = n31504 & n32115 ;
  assign n32124 = ~n32122 & ~n32123 ;
  assign n32118 = ~\P2_P1_InstAddrPointer_reg[18]/NET0131  & ~n32115 ;
  assign n32119 = \P2_P1_InstAddrPointer_reg[18]/NET0131  & n32115 ;
  assign n32120 = ~n32118 & ~n32119 ;
  assign n32125 = \P2_P1_InstAddrPointer_reg[19]/NET0131  & n32120 ;
  assign n32126 = n32124 & n32125 ;
  assign n32127 = n32117 & n32126 ;
  assign n32128 = ~\P2_P1_InstAddrPointer_reg[21]/NET0131  & ~n32032 ;
  assign n32129 = ~n32033 & ~n32128 ;
  assign n32130 = n32127 & n32129 ;
  assign n32134 = n31871 & n32055 ;
  assign n32135 = \P2_P1_InstAddrPointer_reg[24]/NET0131  & ~n32134 ;
  assign n32136 = ~\P2_P1_InstAddrPointer_reg[24]/NET0131  & n32134 ;
  assign n32137 = ~n32135 & ~n32136 ;
  assign n32131 = ~n31845 & n32045 ;
  assign n32132 = \P2_P1_InstAddrPointer_reg[22]/NET0131  & ~n32045 ;
  assign n32133 = ~n32131 & ~n32132 ;
  assign n32138 = ~\P2_P1_InstAddrPointer_reg[23]/NET0131  & ~n32034 ;
  assign n32139 = ~n32035 & ~n32138 ;
  assign n32140 = ~n32133 & n32139 ;
  assign n32141 = ~n32137 & n32140 ;
  assign n32142 = n32130 & n32141 ;
  assign n32143 = n32044 & n32142 ;
  assign n32144 = \P2_P1_InstAddrPointer_reg[26]/NET0131  & n32143 ;
  assign n32145 = \P2_P1_InstAddrPointer_reg[27]/NET0131  & n32144 ;
  assign n32146 = n32042 & n32145 ;
  assign n32147 = \P2_P1_InstAddrPointer_reg[29]/NET0131  & n32146 ;
  assign n32148 = \P2_P1_InstAddrPointer_reg[30]/NET0131  & n32147 ;
  assign n32150 = \P2_P1_InstAddrPointer_reg[29]/NET0131  & n32040 ;
  assign n32151 = \P2_P1_InstAddrPointer_reg[30]/NET0131  & n32150 ;
  assign n32152 = ~\P2_P1_InstAddrPointer_reg[31]/NET0131  & ~n32151 ;
  assign n32153 = \P2_P1_InstAddrPointer_reg[31]/NET0131  & n32151 ;
  assign n32154 = ~n32152 & ~n32153 ;
  assign n32155 = ~n32148 & ~n32154 ;
  assign n32149 = \P2_P1_InstAddrPointer_reg[31]/NET0131  & n32148 ;
  assign n32156 = n25964 & ~n32149 ;
  assign n32157 = ~n32155 & n32156 ;
  assign n32162 = n26068 & n32154 ;
  assign n32161 = ~n25995 & ~n32016 ;
  assign n32026 = n21073 & ~n26031 ;
  assign n32025 = ~n21082 & n26055 ;
  assign n32027 = ~n26037 & n32025 ;
  assign n32028 = ~n32026 & n32027 ;
  assign n32029 = \P2_P1_InstAddrPointer_reg[31]/NET0131  & ~n32028 ;
  assign n32158 = ~n21073 & ~n26031 ;
  assign n32159 = ~n25984 & ~n32158 ;
  assign n32160 = n31866 & ~n32159 ;
  assign n32163 = ~n32029 & ~n32160 ;
  assign n32164 = ~n32161 & n32163 ;
  assign n32165 = ~n32162 & n32164 ;
  assign n32166 = ~n32157 & n32165 ;
  assign n32167 = ~n32024 & n32166 ;
  assign n32168 = n11623 & ~n32167 ;
  assign n32169 = ~n11611 & n11615 ;
  assign n32170 = ~n11608 & ~n11613 ;
  assign n32171 = ~n11621 & n32170 ;
  assign n32172 = ~n32169 & n32171 ;
  assign n32173 = \P2_P1_InstAddrPointer_reg[31]/NET0131  & ~n32172 ;
  assign n32174 = \P2_P1_rEIP_reg[31]/NET0131  & n11616 ;
  assign n32175 = ~n32173 & ~n32174 ;
  assign n32176 = ~n32168 & n32175 ;
  assign n32564 = \P2_P2_InstAddrPointer_reg[27]/NET0131  & \P2_P2_InstAddrPointer_reg[28]/NET0131  ;
  assign n32178 = \P2_P2_InstAddrPointer_reg[21]/NET0131  & \P2_P2_InstAddrPointer_reg[22]/NET0131  ;
  assign n32179 = \P2_P2_InstAddrPointer_reg[17]/NET0131  & \P2_P2_InstAddrPointer_reg[18]/NET0131  ;
  assign n32180 = \P2_P2_InstAddrPointer_reg[15]/NET0131  & \P2_P2_InstAddrPointer_reg[16]/NET0131  ;
  assign n32181 = n32179 & n32180 ;
  assign n32182 = \P2_P2_InstAddrPointer_reg[19]/NET0131  & n32181 ;
  assign n32183 = \P2_P2_InstAddrPointer_reg[20]/NET0131  & n32182 ;
  assign n32188 = \P2_P2_InstAddrPointer_reg[11]/NET0131  & \P2_P2_InstAddrPointer_reg[12]/NET0131  ;
  assign n32189 = \P2_P2_InstAddrPointer_reg[10]/NET0131  & n32188 ;
  assign n32190 = \P2_P2_InstAddrPointer_reg[9]/NET0131  & n32189 ;
  assign n32191 = \P2_P2_InstAddrPointer_reg[13]/NET0131  & \P2_P2_InstAddrPointer_reg[6]/NET0131  ;
  assign n32192 = \P2_P2_InstAddrPointer_reg[7]/NET0131  & \P2_P2_InstAddrPointer_reg[8]/NET0131  ;
  assign n32193 = n32191 & n32192 ;
  assign n32194 = n32190 & n32193 ;
  assign n32584 = \P2_P2_InstAddrPointer_reg[0]/NET0131  & \P2_P2_InstAddrPointer_reg[1]/NET0131  ;
  assign n32603 = ~\P2_P2_InstAddrPointer_reg[2]/NET0131  & ~n32584 ;
  assign n32720 = \P2_P2_InstAddrPointer_reg[3]/NET0131  & ~n32603 ;
  assign n32721 = \P2_P2_InstAddrPointer_reg[4]/NET0131  & n32720 ;
  assign n32722 = \P2_P2_InstAddrPointer_reg[5]/NET0131  & n32721 ;
  assign n32723 = n32194 & n32722 ;
  assign n32724 = \P2_P2_InstAddrPointer_reg[14]/NET0131  & n32723 ;
  assign n32725 = n32183 & n32724 ;
  assign n32726 = n32178 & n32725 ;
  assign n32727 = \P2_P2_InstAddrPointer_reg[23]/NET0131  & n32726 ;
  assign n32728 = \P2_P2_InstAddrPointer_reg[24]/NET0131  & \P2_P2_InstAddrPointer_reg[25]/NET0131  ;
  assign n32729 = n32727 & n32728 ;
  assign n32730 = \P2_P2_InstAddrPointer_reg[26]/NET0131  & n32729 ;
  assign n32731 = n32564 & n32730 ;
  assign n32732 = \P2_P2_InstAddrPointer_reg[29]/NET0131  & n32731 ;
  assign n32733 = \P2_P2_InstAddrPointer_reg[30]/NET0131  & n32732 ;
  assign n32734 = ~\P2_P2_InstAddrPointer_reg[31]/NET0131  & ~n32733 ;
  assign n32735 = \P2_P2_InstAddrPointer_reg[31]/NET0131  & n32733 ;
  assign n32736 = ~n32734 & ~n32735 ;
  assign n32748 = ~\P2_P2_InstAddrPointer_reg[30]/NET0131  & ~n32732 ;
  assign n32749 = ~n32733 & ~n32748 ;
  assign n32750 = ~\P2_P2_InstAddrPointer_reg[23]/NET0131  & ~n32726 ;
  assign n32751 = ~n32727 & ~n32750 ;
  assign n32752 = \P2_P2_InstAddrPointer_reg[15]/NET0131  & n32724 ;
  assign n32753 = \P2_P2_InstAddrPointer_reg[16]/NET0131  & n32752 ;
  assign n32754 = \P2_P2_InstAddrPointer_reg[17]/NET0131  & n32753 ;
  assign n32755 = ~\P2_P2_InstAddrPointer_reg[17]/NET0131  & ~n32753 ;
  assign n32756 = ~n32754 & ~n32755 ;
  assign n32757 = \P2_P2_InstAddrPointer_reg[6]/NET0131  & n32722 ;
  assign n32758 = \P2_P2_InstAddrPointer_reg[7]/NET0131  & n32757 ;
  assign n32759 = \P2_P2_InstAddrPointer_reg[8]/NET0131  & n32758 ;
  assign n32760 = \P2_P2_InstAddrPointer_reg[9]/NET0131  & n32759 ;
  assign n32761 = ~\P2_P2_InstAddrPointer_reg[10]/NET0131  & ~n32760 ;
  assign n32762 = \P2_P2_InstAddrPointer_reg[10]/NET0131  & n32760 ;
  assign n32763 = ~n32761 & ~n32762 ;
  assign n32764 = ~\P2_P2_InstAddrPointer_reg[8]/NET0131  & ~n32758 ;
  assign n32765 = ~n32759 & ~n32764 ;
  assign n32491 = \P2_P2_InstQueue_reg[15][7]/NET0131  & n26330 ;
  assign n32489 = \P2_P2_InstQueue_reg[0][7]/NET0131  & n26325 ;
  assign n32480 = \P2_P2_InstQueue_reg[7][7]/NET0131  & n26300 ;
  assign n32481 = \P2_P2_InstQueue_reg[10][7]/NET0131  & n26304 ;
  assign n32496 = ~n32480 & ~n32481 ;
  assign n32506 = ~n32489 & n32496 ;
  assign n32507 = ~n32491 & n32506 ;
  assign n32492 = \P2_P2_InstQueue_reg[3][7]/NET0131  & n26316 ;
  assign n32493 = \P2_P2_InstQueue_reg[11][7]/NET0131  & n26320 ;
  assign n32501 = ~n32492 & ~n32493 ;
  assign n32494 = \P2_P2_InstQueue_reg[14][7]/NET0131  & n26336 ;
  assign n32495 = \P2_P2_InstQueue_reg[1][7]/NET0131  & n26322 ;
  assign n32502 = ~n32494 & ~n32495 ;
  assign n32503 = n32501 & n32502 ;
  assign n32486 = \P2_P2_InstQueue_reg[9][7]/NET0131  & n26334 ;
  assign n32487 = \P2_P2_InstQueue_reg[13][7]/NET0131  & n26313 ;
  assign n32499 = ~n32486 & ~n32487 ;
  assign n32488 = \P2_P2_InstQueue_reg[5][7]/NET0131  & n26307 ;
  assign n32490 = \P2_P2_InstQueue_reg[8][7]/NET0131  & n26327 ;
  assign n32500 = ~n32488 & ~n32490 ;
  assign n32504 = n32499 & n32500 ;
  assign n32482 = \P2_P2_InstQueue_reg[4][7]/NET0131  & n26332 ;
  assign n32483 = \P2_P2_InstQueue_reg[2][7]/NET0131  & n26338 ;
  assign n32497 = ~n32482 & ~n32483 ;
  assign n32484 = \P2_P2_InstQueue_reg[6][7]/NET0131  & n26318 ;
  assign n32485 = \P2_P2_InstQueue_reg[12][7]/NET0131  & n26310 ;
  assign n32498 = ~n32484 & ~n32485 ;
  assign n32505 = n32497 & n32498 ;
  assign n32508 = n32504 & n32505 ;
  assign n32509 = n32503 & n32508 ;
  assign n32510 = n32507 & n32509 ;
  assign n32766 = ~\P2_P2_InstAddrPointer_reg[7]/NET0131  & ~n32757 ;
  assign n32767 = ~n32758 & ~n32766 ;
  assign n32768 = ~n32510 & n32767 ;
  assign n32769 = n32510 & ~n32767 ;
  assign n32240 = \P2_P2_InstQueue_reg[15][6]/NET0131  & n26330 ;
  assign n32238 = \P2_P2_InstQueue_reg[0][6]/NET0131  & n26325 ;
  assign n32229 = \P2_P2_InstQueue_reg[7][6]/NET0131  & n26300 ;
  assign n32230 = \P2_P2_InstQueue_reg[10][6]/NET0131  & n26304 ;
  assign n32245 = ~n32229 & ~n32230 ;
  assign n32255 = ~n32238 & n32245 ;
  assign n32256 = ~n32240 & n32255 ;
  assign n32241 = \P2_P2_InstQueue_reg[11][6]/NET0131  & n26320 ;
  assign n32242 = \P2_P2_InstQueue_reg[13][6]/NET0131  & n26313 ;
  assign n32250 = ~n32241 & ~n32242 ;
  assign n32243 = \P2_P2_InstQueue_reg[6][6]/NET0131  & n26318 ;
  assign n32244 = \P2_P2_InstQueue_reg[14][6]/NET0131  & n26336 ;
  assign n32251 = ~n32243 & ~n32244 ;
  assign n32252 = n32250 & n32251 ;
  assign n32235 = \P2_P2_InstQueue_reg[12][6]/NET0131  & n26310 ;
  assign n32236 = \P2_P2_InstQueue_reg[1][6]/NET0131  & n26322 ;
  assign n32248 = ~n32235 & ~n32236 ;
  assign n32237 = \P2_P2_InstQueue_reg[3][6]/NET0131  & n26316 ;
  assign n32239 = \P2_P2_InstQueue_reg[8][6]/NET0131  & n26327 ;
  assign n32249 = ~n32237 & ~n32239 ;
  assign n32253 = n32248 & n32249 ;
  assign n32231 = \P2_P2_InstQueue_reg[9][6]/NET0131  & n26334 ;
  assign n32232 = \P2_P2_InstQueue_reg[4][6]/NET0131  & n26332 ;
  assign n32246 = ~n32231 & ~n32232 ;
  assign n32233 = \P2_P2_InstQueue_reg[2][6]/NET0131  & n26338 ;
  assign n32234 = \P2_P2_InstQueue_reg[5][6]/NET0131  & n26307 ;
  assign n32247 = ~n32233 & ~n32234 ;
  assign n32254 = n32246 & n32247 ;
  assign n32257 = n32253 & n32254 ;
  assign n32258 = n32252 & n32257 ;
  assign n32259 = n32256 & n32258 ;
  assign n32770 = ~\P2_P2_InstAddrPointer_reg[6]/NET0131  & ~n32722 ;
  assign n32771 = ~n32757 & ~n32770 ;
  assign n32772 = ~n32259 & n32771 ;
  assign n32773 = n32259 & ~n32771 ;
  assign n32275 = \P2_P2_InstQueue_reg[15][5]/NET0131  & n26330 ;
  assign n32273 = \P2_P2_InstQueue_reg[0][5]/NET0131  & n26325 ;
  assign n32264 = \P2_P2_InstQueue_reg[7][5]/NET0131  & n26300 ;
  assign n32265 = \P2_P2_InstQueue_reg[6][5]/NET0131  & n26318 ;
  assign n32280 = ~n32264 & ~n32265 ;
  assign n32290 = ~n32273 & n32280 ;
  assign n32291 = ~n32275 & n32290 ;
  assign n32276 = \P2_P2_InstQueue_reg[3][5]/NET0131  & n26316 ;
  assign n32277 = \P2_P2_InstQueue_reg[11][5]/NET0131  & n26320 ;
  assign n32285 = ~n32276 & ~n32277 ;
  assign n32278 = \P2_P2_InstQueue_reg[1][5]/NET0131  & n26322 ;
  assign n32279 = \P2_P2_InstQueue_reg[12][5]/NET0131  & n26310 ;
  assign n32286 = ~n32278 & ~n32279 ;
  assign n32287 = n32285 & n32286 ;
  assign n32270 = \P2_P2_InstQueue_reg[10][5]/NET0131  & n26304 ;
  assign n32271 = \P2_P2_InstQueue_reg[5][5]/NET0131  & n26307 ;
  assign n32283 = ~n32270 & ~n32271 ;
  assign n32272 = \P2_P2_InstQueue_reg[4][5]/NET0131  & n26332 ;
  assign n32274 = \P2_P2_InstQueue_reg[8][5]/NET0131  & n26327 ;
  assign n32284 = ~n32272 & ~n32274 ;
  assign n32288 = n32283 & n32284 ;
  assign n32266 = \P2_P2_InstQueue_reg[9][5]/NET0131  & n26334 ;
  assign n32267 = \P2_P2_InstQueue_reg[2][5]/NET0131  & n26338 ;
  assign n32281 = ~n32266 & ~n32267 ;
  assign n32268 = \P2_P2_InstQueue_reg[14][5]/NET0131  & n26336 ;
  assign n32269 = \P2_P2_InstQueue_reg[13][5]/NET0131  & n26313 ;
  assign n32282 = ~n32268 & ~n32269 ;
  assign n32289 = n32281 & n32282 ;
  assign n32292 = n32288 & n32289 ;
  assign n32293 = n32287 & n32292 ;
  assign n32294 = n32291 & n32293 ;
  assign n32774 = ~\P2_P2_InstAddrPointer_reg[5]/NET0131  & ~n32721 ;
  assign n32775 = ~n32722 & ~n32774 ;
  assign n32776 = ~n32294 & n32775 ;
  assign n32777 = n32294 & ~n32775 ;
  assign n32310 = \P2_P2_InstQueue_reg[15][4]/NET0131  & n26330 ;
  assign n32308 = \P2_P2_InstQueue_reg[0][4]/NET0131  & n26325 ;
  assign n32299 = \P2_P2_InstQueue_reg[7][4]/NET0131  & n26300 ;
  assign n32300 = \P2_P2_InstQueue_reg[11][4]/NET0131  & n26320 ;
  assign n32315 = ~n32299 & ~n32300 ;
  assign n32325 = ~n32308 & n32315 ;
  assign n32326 = ~n32310 & n32325 ;
  assign n32311 = \P2_P2_InstQueue_reg[1][4]/NET0131  & n26322 ;
  assign n32312 = \P2_P2_InstQueue_reg[5][4]/NET0131  & n26307 ;
  assign n32320 = ~n32311 & ~n32312 ;
  assign n32313 = \P2_P2_InstQueue_reg[14][4]/NET0131  & n26336 ;
  assign n32314 = \P2_P2_InstQueue_reg[3][4]/NET0131  & n26316 ;
  assign n32321 = ~n32313 & ~n32314 ;
  assign n32322 = n32320 & n32321 ;
  assign n32305 = \P2_P2_InstQueue_reg[2][4]/NET0131  & n26338 ;
  assign n32306 = \P2_P2_InstQueue_reg[6][4]/NET0131  & n26318 ;
  assign n32318 = ~n32305 & ~n32306 ;
  assign n32307 = \P2_P2_InstQueue_reg[4][4]/NET0131  & n26332 ;
  assign n32309 = \P2_P2_InstQueue_reg[8][4]/NET0131  & n26327 ;
  assign n32319 = ~n32307 & ~n32309 ;
  assign n32323 = n32318 & n32319 ;
  assign n32301 = \P2_P2_InstQueue_reg[10][4]/NET0131  & n26304 ;
  assign n32302 = \P2_P2_InstQueue_reg[9][4]/NET0131  & n26334 ;
  assign n32316 = ~n32301 & ~n32302 ;
  assign n32303 = \P2_P2_InstQueue_reg[12][4]/NET0131  & n26310 ;
  assign n32304 = \P2_P2_InstQueue_reg[13][4]/NET0131  & n26313 ;
  assign n32317 = ~n32303 & ~n32304 ;
  assign n32324 = n32316 & n32317 ;
  assign n32327 = n32323 & n32324 ;
  assign n32328 = n32322 & n32327 ;
  assign n32329 = n32326 & n32328 ;
  assign n32778 = ~\P2_P2_InstAddrPointer_reg[4]/NET0131  & ~n32720 ;
  assign n32779 = ~n32721 & ~n32778 ;
  assign n32780 = ~n32329 & n32779 ;
  assign n32781 = n32329 & ~n32779 ;
  assign n32345 = \P2_P2_InstQueue_reg[15][3]/NET0131  & n26330 ;
  assign n32343 = \P2_P2_InstQueue_reg[0][3]/NET0131  & n26325 ;
  assign n32334 = \P2_P2_InstQueue_reg[7][3]/NET0131  & n26300 ;
  assign n32335 = \P2_P2_InstQueue_reg[11][3]/NET0131  & n26320 ;
  assign n32350 = ~n32334 & ~n32335 ;
  assign n32360 = ~n32343 & n32350 ;
  assign n32361 = ~n32345 & n32360 ;
  assign n32346 = \P2_P2_InstQueue_reg[1][3]/NET0131  & n26322 ;
  assign n32347 = \P2_P2_InstQueue_reg[5][3]/NET0131  & n26307 ;
  assign n32355 = ~n32346 & ~n32347 ;
  assign n32348 = \P2_P2_InstQueue_reg[14][3]/NET0131  & n26336 ;
  assign n32349 = \P2_P2_InstQueue_reg[3][3]/NET0131  & n26316 ;
  assign n32356 = ~n32348 & ~n32349 ;
  assign n32357 = n32355 & n32356 ;
  assign n32340 = \P2_P2_InstQueue_reg[2][3]/NET0131  & n26338 ;
  assign n32341 = \P2_P2_InstQueue_reg[6][3]/NET0131  & n26318 ;
  assign n32353 = ~n32340 & ~n32341 ;
  assign n32342 = \P2_P2_InstQueue_reg[4][3]/NET0131  & n26332 ;
  assign n32344 = \P2_P2_InstQueue_reg[8][3]/NET0131  & n26327 ;
  assign n32354 = ~n32342 & ~n32344 ;
  assign n32358 = n32353 & n32354 ;
  assign n32336 = \P2_P2_InstQueue_reg[10][3]/NET0131  & n26304 ;
  assign n32337 = \P2_P2_InstQueue_reg[9][3]/NET0131  & n26334 ;
  assign n32351 = ~n32336 & ~n32337 ;
  assign n32338 = \P2_P2_InstQueue_reg[12][3]/NET0131  & n26310 ;
  assign n32339 = \P2_P2_InstQueue_reg[13][3]/NET0131  & n26313 ;
  assign n32352 = ~n32338 & ~n32339 ;
  assign n32359 = n32351 & n32352 ;
  assign n32362 = n32358 & n32359 ;
  assign n32363 = n32357 & n32362 ;
  assign n32364 = n32361 & n32363 ;
  assign n32782 = ~\P2_P2_InstAddrPointer_reg[3]/NET0131  & n32603 ;
  assign n32783 = ~n32720 & ~n32782 ;
  assign n32784 = n32364 & ~n32783 ;
  assign n32785 = ~n32364 & n32783 ;
  assign n32381 = \P2_P2_InstQueue_reg[15][2]/NET0131  & n26330 ;
  assign n32374 = \P2_P2_InstQueue_reg[0][2]/NET0131  & n26325 ;
  assign n32369 = \P2_P2_InstQueue_reg[7][2]/NET0131  & n26300 ;
  assign n32370 = \P2_P2_InstQueue_reg[14][2]/NET0131  & n26336 ;
  assign n32385 = ~n32369 & ~n32370 ;
  assign n32395 = ~n32374 & n32385 ;
  assign n32396 = ~n32381 & n32395 ;
  assign n32380 = \P2_P2_InstQueue_reg[4][2]/NET0131  & n26332 ;
  assign n32382 = \P2_P2_InstQueue_reg[6][2]/NET0131  & n26318 ;
  assign n32390 = ~n32380 & ~n32382 ;
  assign n32383 = \P2_P2_InstQueue_reg[1][2]/NET0131  & n26322 ;
  assign n32384 = \P2_P2_InstQueue_reg[9][2]/NET0131  & n26334 ;
  assign n32391 = ~n32383 & ~n32384 ;
  assign n32392 = n32390 & n32391 ;
  assign n32376 = \P2_P2_InstQueue_reg[3][2]/NET0131  & n26316 ;
  assign n32377 = \P2_P2_InstQueue_reg[12][2]/NET0131  & n26310 ;
  assign n32388 = ~n32376 & ~n32377 ;
  assign n32378 = \P2_P2_InstQueue_reg[13][2]/NET0131  & n26313 ;
  assign n32379 = \P2_P2_InstQueue_reg[2][2]/NET0131  & n26338 ;
  assign n32389 = ~n32378 & ~n32379 ;
  assign n32393 = n32388 & n32389 ;
  assign n32371 = \P2_P2_InstQueue_reg[8][2]/NET0131  & n26327 ;
  assign n32372 = \P2_P2_InstQueue_reg[11][2]/NET0131  & n26320 ;
  assign n32386 = ~n32371 & ~n32372 ;
  assign n32373 = \P2_P2_InstQueue_reg[5][2]/NET0131  & n26307 ;
  assign n32375 = \P2_P2_InstQueue_reg[10][2]/NET0131  & n26304 ;
  assign n32387 = ~n32373 & ~n32375 ;
  assign n32394 = n32386 & n32387 ;
  assign n32397 = n32393 & n32394 ;
  assign n32398 = n32392 & n32397 ;
  assign n32399 = n32396 & n32398 ;
  assign n32585 = \P2_P2_InstAddrPointer_reg[2]/NET0131  & n32584 ;
  assign n32604 = ~n32585 & ~n32603 ;
  assign n32786 = n32399 & n32604 ;
  assign n32787 = ~n32399 & ~n32604 ;
  assign n32403 = \P2_P2_InstQueue_reg[0][1]/NET0131  & n26325 ;
  assign n32402 = \P2_P2_InstQueue_reg[15][1]/NET0131  & n26330 ;
  assign n32404 = \P2_P2_InstQueue_reg[9][1]/NET0131  & n26334 ;
  assign n32405 = \P2_P2_InstQueue_reg[2][1]/NET0131  & n26338 ;
  assign n32418 = ~n32404 & ~n32405 ;
  assign n32428 = ~n32402 & n32418 ;
  assign n32429 = ~n32403 & n32428 ;
  assign n32414 = \P2_P2_InstQueue_reg[12][1]/NET0131  & n26310 ;
  assign n32415 = \P2_P2_InstQueue_reg[11][1]/NET0131  & n26320 ;
  assign n32423 = ~n32414 & ~n32415 ;
  assign n32416 = \P2_P2_InstQueue_reg[1][1]/NET0131  & n26322 ;
  assign n32417 = \P2_P2_InstQueue_reg[14][1]/NET0131  & n26336 ;
  assign n32424 = ~n32416 & ~n32417 ;
  assign n32425 = n32423 & n32424 ;
  assign n32410 = \P2_P2_InstQueue_reg[7][1]/NET0131  & n26300 ;
  assign n32411 = \P2_P2_InstQueue_reg[3][1]/NET0131  & n26316 ;
  assign n32421 = ~n32410 & ~n32411 ;
  assign n32412 = \P2_P2_InstQueue_reg[6][1]/NET0131  & n26318 ;
  assign n32413 = \P2_P2_InstQueue_reg[5][1]/NET0131  & n26307 ;
  assign n32422 = ~n32412 & ~n32413 ;
  assign n32426 = n32421 & n32422 ;
  assign n32406 = \P2_P2_InstQueue_reg[8][1]/NET0131  & n26327 ;
  assign n32407 = \P2_P2_InstQueue_reg[10][1]/NET0131  & n26304 ;
  assign n32419 = ~n32406 & ~n32407 ;
  assign n32408 = \P2_P2_InstQueue_reg[13][1]/NET0131  & n26313 ;
  assign n32409 = \P2_P2_InstQueue_reg[4][1]/NET0131  & n26332 ;
  assign n32420 = ~n32408 & ~n32409 ;
  assign n32427 = n32419 & n32420 ;
  assign n32430 = n32426 & n32427 ;
  assign n32431 = n32425 & n32430 ;
  assign n32432 = n32429 & n32431 ;
  assign n32607 = ~\P2_P2_InstAddrPointer_reg[0]/NET0131  & ~\P2_P2_InstAddrPointer_reg[1]/NET0131  ;
  assign n32608 = ~n32584 & ~n32607 ;
  assign n32609 = n32432 & ~n32608 ;
  assign n32788 = ~n32432 & n32608 ;
  assign n32436 = \P2_P2_InstQueue_reg[0][0]/NET0131  & n26325 ;
  assign n32435 = \P2_P2_InstQueue_reg[15][0]/NET0131  & n26330 ;
  assign n32437 = \P2_P2_InstQueue_reg[1][0]/NET0131  & n26322 ;
  assign n32438 = \P2_P2_InstQueue_reg[4][0]/NET0131  & n26332 ;
  assign n32451 = ~n32437 & ~n32438 ;
  assign n32461 = ~n32435 & n32451 ;
  assign n32462 = ~n32436 & n32461 ;
  assign n32447 = \P2_P2_InstQueue_reg[6][0]/NET0131  & n26318 ;
  assign n32448 = \P2_P2_InstQueue_reg[11][0]/NET0131  & n26320 ;
  assign n32456 = ~n32447 & ~n32448 ;
  assign n32449 = \P2_P2_InstQueue_reg[13][0]/NET0131  & n26313 ;
  assign n32450 = \P2_P2_InstQueue_reg[5][0]/NET0131  & n26307 ;
  assign n32457 = ~n32449 & ~n32450 ;
  assign n32458 = n32456 & n32457 ;
  assign n32443 = \P2_P2_InstQueue_reg[7][0]/NET0131  & n26300 ;
  assign n32444 = \P2_P2_InstQueue_reg[10][0]/NET0131  & n26304 ;
  assign n32454 = ~n32443 & ~n32444 ;
  assign n32445 = \P2_P2_InstQueue_reg[2][0]/NET0131  & n26338 ;
  assign n32446 = \P2_P2_InstQueue_reg[9][0]/NET0131  & n26334 ;
  assign n32455 = ~n32445 & ~n32446 ;
  assign n32459 = n32454 & n32455 ;
  assign n32439 = \P2_P2_InstQueue_reg[8][0]/NET0131  & n26327 ;
  assign n32440 = \P2_P2_InstQueue_reg[3][0]/NET0131  & n26316 ;
  assign n32452 = ~n32439 & ~n32440 ;
  assign n32441 = \P2_P2_InstQueue_reg[14][0]/NET0131  & n26336 ;
  assign n32442 = \P2_P2_InstQueue_reg[12][0]/NET0131  & n26310 ;
  assign n32453 = ~n32441 & ~n32442 ;
  assign n32460 = n32452 & n32453 ;
  assign n32463 = n32459 & n32460 ;
  assign n32464 = n32458 & n32463 ;
  assign n32465 = n32462 & n32464 ;
  assign n32789 = ~\P2_P2_InstAddrPointer_reg[0]/NET0131  & ~n32465 ;
  assign n32790 = ~n32788 & ~n32789 ;
  assign n32791 = ~n32609 & ~n32790 ;
  assign n32792 = ~n32787 & ~n32791 ;
  assign n32793 = ~n32786 & ~n32792 ;
  assign n32794 = ~n32785 & ~n32793 ;
  assign n32795 = ~n32784 & ~n32794 ;
  assign n32796 = ~n32781 & n32795 ;
  assign n32797 = ~n32780 & ~n32796 ;
  assign n32798 = ~n32777 & ~n32797 ;
  assign n32799 = ~n32776 & ~n32798 ;
  assign n32800 = ~n32773 & ~n32799 ;
  assign n32801 = ~n32772 & ~n32800 ;
  assign n32802 = ~n32769 & ~n32801 ;
  assign n32803 = ~n32768 & ~n32802 ;
  assign n32804 = n32765 & ~n32803 ;
  assign n32805 = \P2_P2_InstAddrPointer_reg[9]/NET0131  & n32804 ;
  assign n32806 = n32763 & n32805 ;
  assign n32807 = n32188 & n32806 ;
  assign n32808 = n32189 & n32760 ;
  assign n32809 = ~\P2_P2_InstAddrPointer_reg[13]/NET0131  & ~n32808 ;
  assign n32810 = ~n32723 & ~n32809 ;
  assign n32811 = n32807 & n32810 ;
  assign n32812 = \P2_P2_InstAddrPointer_reg[14]/NET0131  & n32811 ;
  assign n32813 = ~\P2_P2_InstAddrPointer_reg[15]/NET0131  & ~n32724 ;
  assign n32814 = ~n32752 & ~n32813 ;
  assign n32815 = n32812 & n32814 ;
  assign n32816 = \P2_P2_InstAddrPointer_reg[16]/NET0131  & n32815 ;
  assign n32817 = n32756 & n32816 ;
  assign n32818 = \P2_P2_InstAddrPointer_reg[18]/NET0131  & n32817 ;
  assign n32819 = n32179 & n32753 ;
  assign n32820 = ~\P2_P2_InstAddrPointer_reg[19]/NET0131  & ~n32819 ;
  assign n32821 = \P2_P2_InstAddrPointer_reg[19]/NET0131  & n32819 ;
  assign n32822 = ~n32820 & ~n32821 ;
  assign n32823 = n32818 & n32822 ;
  assign n32824 = \P2_P2_InstAddrPointer_reg[20]/NET0131  & n32823 ;
  assign n32825 = ~\P2_P2_InstAddrPointer_reg[21]/NET0131  & ~n32725 ;
  assign n32534 = \P2_P2_InstAddrPointer_reg[21]/NET0131  & n32183 ;
  assign n32826 = n32534 & n32724 ;
  assign n32827 = ~n32825 & ~n32826 ;
  assign n32828 = n32824 & n32827 ;
  assign n32829 = \P2_P2_InstAddrPointer_reg[22]/NET0131  & n32828 ;
  assign n32830 = n32751 & n32829 ;
  assign n32831 = ~\P2_P2_InstAddrPointer_reg[24]/NET0131  & ~n32727 ;
  assign n32832 = \P2_P2_InstAddrPointer_reg[24]/NET0131  & n32727 ;
  assign n32833 = ~n32831 & ~n32832 ;
  assign n32834 = \P2_P2_InstAddrPointer_reg[25]/NET0131  & n32833 ;
  assign n32835 = n32830 & n32834 ;
  assign n32836 = ~\P2_P2_InstAddrPointer_reg[26]/NET0131  & ~n32729 ;
  assign n32837 = ~n32730 & ~n32836 ;
  assign n32838 = n32835 & n32837 ;
  assign n32839 = \P2_P2_InstAddrPointer_reg[27]/NET0131  & n32838 ;
  assign n32840 = \P2_P2_InstAddrPointer_reg[27]/NET0131  & n32730 ;
  assign n32841 = ~\P2_P2_InstAddrPointer_reg[28]/NET0131  & ~n32840 ;
  assign n32842 = ~n32731 & ~n32841 ;
  assign n32843 = \P2_P2_InstAddrPointer_reg[29]/NET0131  & n32842 ;
  assign n32844 = n32839 & n32843 ;
  assign n32845 = n32749 & n32844 ;
  assign n32847 = ~n32736 & ~n32845 ;
  assign n32846 = \P2_P2_InstAddrPointer_reg[31]/NET0131  & n32845 ;
  assign n32848 = n26744 & ~n32846 ;
  assign n32849 = ~n32847 & n32848 ;
  assign n32177 = \P2_P2_InstAddrPointer_reg[31]/NET0131  & n26629 ;
  assign n32184 = \P2_P2_InstAddrPointer_reg[1]/NET0131  & \P2_P2_InstAddrPointer_reg[2]/NET0131  ;
  assign n32185 = \P2_P2_InstAddrPointer_reg[3]/NET0131  & n32184 ;
  assign n32186 = \P2_P2_InstAddrPointer_reg[4]/NET0131  & n32185 ;
  assign n32187 = \P2_P2_InstAddrPointer_reg[5]/NET0131  & n32186 ;
  assign n32195 = \P2_P2_InstAddrPointer_reg[14]/NET0131  & n32194 ;
  assign n32196 = n32187 & n32195 ;
  assign n32197 = n32183 & n32196 ;
  assign n32198 = n32178 & n32197 ;
  assign n32199 = \P2_P2_InstAddrPointer_reg[23]/NET0131  & n32198 ;
  assign n32200 = \P2_P2_InstAddrPointer_reg[24]/NET0131  & n32199 ;
  assign n32201 = \P2_P2_InstAddrPointer_reg[25]/NET0131  & n32200 ;
  assign n32202 = \P2_P2_InstAddrPointer_reg[26]/NET0131  & n32201 ;
  assign n32203 = \P2_P2_InstAddrPointer_reg[27]/NET0131  & n32202 ;
  assign n32204 = \P2_P2_InstAddrPointer_reg[28]/NET0131  & n32203 ;
  assign n32205 = \P2_P2_InstAddrPointer_reg[29]/NET0131  & n32204 ;
  assign n32206 = ~\P2_P2_InstAddrPointer_reg[29]/NET0131  & ~n32204 ;
  assign n32207 = ~n32205 & ~n32206 ;
  assign n32208 = \P2_P2_InstAddrPointer_reg[28]/NET0131  & n32207 ;
  assign n32209 = ~\P2_P2_InstAddrPointer_reg[27]/NET0131  & ~n32202 ;
  assign n32210 = ~n32203 & ~n32209 ;
  assign n32211 = \P2_P2_InstAddrPointer_reg[15]/NET0131  & n32196 ;
  assign n32212 = ~\P2_P2_InstAddrPointer_reg[15]/NET0131  & ~n32196 ;
  assign n32213 = ~n32211 & ~n32212 ;
  assign n32214 = n32187 & n32194 ;
  assign n32215 = \P2_P2_InstAddrPointer_reg[6]/NET0131  & n32187 ;
  assign n32216 = \P2_P2_InstAddrPointer_reg[7]/NET0131  & n32215 ;
  assign n32217 = \P2_P2_InstAddrPointer_reg[8]/NET0131  & n32216 ;
  assign n32218 = n32190 & n32217 ;
  assign n32219 = ~\P2_P2_InstAddrPointer_reg[13]/NET0131  & ~n32218 ;
  assign n32220 = ~n32214 & ~n32219 ;
  assign n32221 = \P2_P2_InstAddrPointer_reg[9]/NET0131  & n32217 ;
  assign n32222 = \P2_P2_InstAddrPointer_reg[10]/NET0131  & n32221 ;
  assign n32223 = ~\P2_P2_InstAddrPointer_reg[10]/NET0131  & ~n32221 ;
  assign n32224 = ~n32222 & ~n32223 ;
  assign n32225 = ~\P2_P2_InstAddrPointer_reg[7]/NET0131  & ~n32215 ;
  assign n32226 = ~n32216 & ~n32225 ;
  assign n32227 = ~\P2_P2_InstAddrPointer_reg[6]/NET0131  & ~n32187 ;
  assign n32228 = ~n32215 & ~n32227 ;
  assign n32260 = n32228 & ~n32259 ;
  assign n32261 = ~n32228 & n32259 ;
  assign n32262 = ~\P2_P2_InstAddrPointer_reg[5]/NET0131  & ~n32186 ;
  assign n32263 = ~n32187 & ~n32262 ;
  assign n32295 = n32263 & ~n32294 ;
  assign n32296 = ~n32263 & n32294 ;
  assign n32297 = ~\P2_P2_InstAddrPointer_reg[4]/NET0131  & ~n32185 ;
  assign n32298 = ~n32186 & ~n32297 ;
  assign n32330 = n32298 & ~n32329 ;
  assign n32331 = ~n32298 & n32329 ;
  assign n32332 = ~\P2_P2_InstAddrPointer_reg[3]/NET0131  & ~n32184 ;
  assign n32333 = ~n32185 & ~n32332 ;
  assign n32365 = n32333 & ~n32364 ;
  assign n32366 = ~n32333 & n32364 ;
  assign n32367 = ~\P2_P2_InstAddrPointer_reg[1]/NET0131  & ~\P2_P2_InstAddrPointer_reg[2]/NET0131  ;
  assign n32368 = ~n32184 & ~n32367 ;
  assign n32400 = n32368 & ~n32399 ;
  assign n32401 = ~n32368 & n32399 ;
  assign n32433 = ~\P2_P2_InstAddrPointer_reg[1]/NET0131  & ~n32432 ;
  assign n32434 = \P2_P2_InstAddrPointer_reg[1]/NET0131  & n32432 ;
  assign n32466 = \P2_P2_InstAddrPointer_reg[0]/NET0131  & ~n32465 ;
  assign n32467 = ~n32434 & n32466 ;
  assign n32468 = ~n32433 & ~n32467 ;
  assign n32469 = ~n32401 & ~n32468 ;
  assign n32470 = ~n32400 & ~n32469 ;
  assign n32471 = ~n32366 & ~n32470 ;
  assign n32472 = ~n32365 & ~n32471 ;
  assign n32473 = ~n32331 & ~n32472 ;
  assign n32474 = ~n32330 & ~n32473 ;
  assign n32475 = ~n32296 & ~n32474 ;
  assign n32476 = ~n32295 & ~n32475 ;
  assign n32477 = ~n32261 & ~n32476 ;
  assign n32478 = ~n32260 & ~n32477 ;
  assign n32479 = n32226 & ~n32478 ;
  assign n32511 = ~n32479 & n32510 ;
  assign n32512 = ~\P2_P2_InstAddrPointer_reg[8]/NET0131  & ~n32216 ;
  assign n32513 = ~n32217 & ~n32512 ;
  assign n32514 = ~n32226 & n32478 ;
  assign n32515 = n32513 & ~n32514 ;
  assign n32516 = ~n32511 & n32515 ;
  assign n32517 = \P2_P2_InstAddrPointer_reg[9]/NET0131  & n32516 ;
  assign n32518 = n32224 & n32517 ;
  assign n32519 = n32188 & n32518 ;
  assign n32520 = n32220 & n32519 ;
  assign n32521 = \P2_P2_InstAddrPointer_reg[14]/NET0131  & n32520 ;
  assign n32522 = n32213 & n32521 ;
  assign n32523 = \P2_P2_InstAddrPointer_reg[16]/NET0131  & n32211 ;
  assign n32524 = ~\P2_P2_InstAddrPointer_reg[16]/NET0131  & ~n32211 ;
  assign n32525 = ~n32523 & ~n32524 ;
  assign n32526 = n32179 & n32525 ;
  assign n32527 = \P2_P2_InstAddrPointer_reg[19]/NET0131  & n32526 ;
  assign n32528 = n32522 & n32527 ;
  assign n32529 = n32182 & n32196 ;
  assign n32530 = ~\P2_P2_InstAddrPointer_reg[20]/NET0131  & ~n32529 ;
  assign n32531 = ~n32197 & ~n32530 ;
  assign n32532 = n32528 & n32531 ;
  assign n32533 = \P2_P2_InstAddrPointer_reg[21]/NET0131  & n32532 ;
  assign n32542 = ~\P2_P2_InstAddrPointer_reg[23]/NET0131  & ~n32198 ;
  assign n32543 = ~n32199 & ~n32542 ;
  assign n32535 = n32195 & n32534 ;
  assign n32536 = \P2_P2_InstAddrPointer_reg[22]/NET0131  & ~n32535 ;
  assign n32537 = ~\P2_P2_InstAddrPointer_reg[22]/NET0131  & n32535 ;
  assign n32538 = ~n32536 & ~n32537 ;
  assign n32539 = n32187 & ~n32538 ;
  assign n32540 = \P2_P2_InstAddrPointer_reg[22]/NET0131  & ~n32187 ;
  assign n32541 = ~n32539 & ~n32540 ;
  assign n32544 = \P2_P2_InstAddrPointer_reg[24]/NET0131  & ~n32541 ;
  assign n32545 = n32543 & n32544 ;
  assign n32546 = n32533 & n32545 ;
  assign n32547 = ~\P2_P2_InstAddrPointer_reg[25]/NET0131  & ~n32200 ;
  assign n32548 = ~n32201 & ~n32547 ;
  assign n32549 = n32546 & n32548 ;
  assign n32550 = \P2_P2_InstAddrPointer_reg[26]/NET0131  & n32549 ;
  assign n32551 = n32210 & n32550 ;
  assign n32552 = n32208 & n32551 ;
  assign n32553 = \P2_P2_InstAddrPointer_reg[30]/NET0131  & n32205 ;
  assign n32554 = ~\P2_P2_InstAddrPointer_reg[30]/NET0131  & ~n32205 ;
  assign n32555 = ~n32553 & ~n32554 ;
  assign n32556 = n32552 & n32555 ;
  assign n32561 = ~\P2_P2_InstAddrPointer_reg[31]/NET0131  & n32556 ;
  assign n32557 = ~\P2_P2_InstAddrPointer_reg[31]/NET0131  & n32553 ;
  assign n32558 = \P2_P2_InstAddrPointer_reg[31]/NET0131  & ~n32553 ;
  assign n32559 = ~n32557 & ~n32558 ;
  assign n32560 = ~n32556 & ~n32559 ;
  assign n32562 = n32510 & ~n32560 ;
  assign n32563 = ~n32561 & n32562 ;
  assign n32565 = \P2_P2_InstAddrPointer_reg[0]/NET0131  & n32200 ;
  assign n32566 = \P2_P2_InstAddrPointer_reg[25]/NET0131  & n32565 ;
  assign n32567 = \P2_P2_InstAddrPointer_reg[26]/NET0131  & n32566 ;
  assign n32568 = n32564 & n32567 ;
  assign n32569 = \P2_P2_InstAddrPointer_reg[29]/NET0131  & n32568 ;
  assign n32570 = \P2_P2_InstAddrPointer_reg[30]/NET0131  & n32569 ;
  assign n32571 = \P2_P2_InstAddrPointer_reg[31]/NET0131  & ~n32570 ;
  assign n32572 = \P2_P2_InstAddrPointer_reg[0]/NET0131  & n32557 ;
  assign n32573 = ~n32571 & ~n32572 ;
  assign n32574 = ~\P2_P2_InstAddrPointer_reg[25]/NET0131  & ~n32565 ;
  assign n32575 = ~n32566 & ~n32574 ;
  assign n32576 = \P2_P2_InstAddrPointer_reg[0]/NET0131  & n32199 ;
  assign n32577 = ~\P2_P2_InstAddrPointer_reg[24]/NET0131  & ~n32576 ;
  assign n32578 = ~n32565 & ~n32577 ;
  assign n32579 = \P2_P2_InstAddrPointer_reg[11]/NET0131  & n32222 ;
  assign n32580 = \P2_P2_InstAddrPointer_reg[0]/NET0131  & n32579 ;
  assign n32581 = ~\P2_P2_InstAddrPointer_reg[12]/NET0131  & ~n32580 ;
  assign n32582 = \P2_P2_InstAddrPointer_reg[0]/NET0131  & n32218 ;
  assign n32583 = ~n32581 & ~n32582 ;
  assign n32586 = \P2_P2_InstAddrPointer_reg[3]/NET0131  & n32585 ;
  assign n32587 = \P2_P2_InstAddrPointer_reg[4]/NET0131  & n32586 ;
  assign n32588 = \P2_P2_InstAddrPointer_reg[5]/NET0131  & n32587 ;
  assign n32589 = \P2_P2_InstAddrPointer_reg[6]/NET0131  & n32588 ;
  assign n32590 = ~\P2_P2_InstAddrPointer_reg[7]/NET0131  & ~n32589 ;
  assign n32591 = \P2_P2_InstAddrPointer_reg[7]/NET0131  & n32589 ;
  assign n32592 = ~n32590 & ~n32591 ;
  assign n32593 = ~\P2_P2_InstAddrPointer_reg[6]/NET0131  & ~n32588 ;
  assign n32594 = ~n32589 & ~n32593 ;
  assign n32595 = ~n32259 & n32594 ;
  assign n32596 = n32259 & ~n32594 ;
  assign n32597 = ~\P2_P2_InstAddrPointer_reg[5]/NET0131  & ~n32587 ;
  assign n32598 = ~n32588 & ~n32597 ;
  assign n32599 = n32294 & ~n32598 ;
  assign n32600 = ~\P2_P2_InstAddrPointer_reg[3]/NET0131  & ~n32585 ;
  assign n32601 = ~n32586 & ~n32600 ;
  assign n32602 = ~n32364 & n32601 ;
  assign n32605 = ~n32399 & n32604 ;
  assign n32606 = n32399 & ~n32604 ;
  assign n32610 = \P2_P2_InstAddrPointer_reg[0]/NET0131  & n32465 ;
  assign n32611 = ~n32433 & n32610 ;
  assign n32612 = ~n32609 & ~n32611 ;
  assign n32613 = ~n32606 & n32612 ;
  assign n32614 = ~n32605 & ~n32613 ;
  assign n32615 = ~n32602 & n32614 ;
  assign n32616 = n32364 & ~n32601 ;
  assign n32617 = ~\P2_P2_InstAddrPointer_reg[4]/NET0131  & ~n32586 ;
  assign n32618 = ~n32587 & ~n32617 ;
  assign n32619 = n32329 & ~n32618 ;
  assign n32620 = ~n32616 & ~n32619 ;
  assign n32621 = ~n32615 & n32620 ;
  assign n32622 = ~n32294 & n32598 ;
  assign n32623 = ~n32329 & n32618 ;
  assign n32624 = ~n32622 & ~n32623 ;
  assign n32625 = ~n32621 & n32624 ;
  assign n32626 = ~n32599 & ~n32625 ;
  assign n32627 = ~n32596 & n32626 ;
  assign n32628 = ~n32595 & ~n32627 ;
  assign n32629 = n32592 & ~n32628 ;
  assign n32630 = ~n32592 & n32628 ;
  assign n32631 = ~n32510 & ~n32630 ;
  assign n32632 = ~n32629 & ~n32631 ;
  assign n32633 = ~\P2_P2_InstAddrPointer_reg[8]/NET0131  & ~n32591 ;
  assign n32634 = \P2_P2_InstAddrPointer_reg[8]/NET0131  & n32591 ;
  assign n32635 = ~n32633 & ~n32634 ;
  assign n32636 = n32632 & ~n32635 ;
  assign n32637 = ~\P2_P2_InstAddrPointer_reg[9]/NET0131  & ~n32634 ;
  assign n32638 = \P2_P2_InstAddrPointer_reg[0]/NET0131  & n32221 ;
  assign n32639 = ~n32637 & ~n32638 ;
  assign n32640 = n32636 & ~n32639 ;
  assign n32641 = ~\P2_P2_InstAddrPointer_reg[10]/NET0131  & ~n32638 ;
  assign n32642 = \P2_P2_InstAddrPointer_reg[0]/NET0131  & n32222 ;
  assign n32643 = ~n32641 & ~n32642 ;
  assign n32644 = ~\P2_P2_InstAddrPointer_reg[11]/NET0131  & ~n32642 ;
  assign n32645 = ~n32580 & ~n32644 ;
  assign n32646 = ~n32643 & ~n32645 ;
  assign n32647 = n32640 & n32646 ;
  assign n32648 = ~n32583 & n32647 ;
  assign n32649 = n32194 & n32588 ;
  assign n32650 = ~\P2_P2_InstAddrPointer_reg[14]/NET0131  & ~n32649 ;
  assign n32651 = n32195 & n32588 ;
  assign n32652 = ~n32650 & ~n32651 ;
  assign n32653 = ~\P2_P2_InstAddrPointer_reg[13]/NET0131  & ~n32582 ;
  assign n32654 = ~n32649 & ~n32653 ;
  assign n32655 = ~n32652 & ~n32654 ;
  assign n32656 = n32648 & n32655 ;
  assign n32657 = ~\P2_P2_InstAddrPointer_reg[15]/NET0131  & ~n32651 ;
  assign n32658 = \P2_P2_InstAddrPointer_reg[15]/NET0131  & n32651 ;
  assign n32659 = ~n32657 & ~n32658 ;
  assign n32660 = ~\P2_P2_InstAddrPointer_reg[16]/NET0131  & ~n32658 ;
  assign n32661 = \P2_P2_InstAddrPointer_reg[16]/NET0131  & n32658 ;
  assign n32662 = ~n32660 & ~n32661 ;
  assign n32663 = ~n32659 & ~n32662 ;
  assign n32664 = n32656 & n32663 ;
  assign n32665 = ~\P2_P2_InstAddrPointer_reg[17]/NET0131  & ~n32661 ;
  assign n32666 = \P2_P2_InstAddrPointer_reg[17]/NET0131  & n32661 ;
  assign n32667 = ~n32665 & ~n32666 ;
  assign n32668 = n32664 & ~n32667 ;
  assign n32669 = n32181 & n32196 ;
  assign n32670 = \P2_P2_InstAddrPointer_reg[0]/NET0131  & n32669 ;
  assign n32671 = ~\P2_P2_InstAddrPointer_reg[19]/NET0131  & ~n32670 ;
  assign n32672 = n32182 & n32651 ;
  assign n32673 = ~n32671 & ~n32672 ;
  assign n32674 = ~\P2_P2_InstAddrPointer_reg[18]/NET0131  & ~n32666 ;
  assign n32675 = ~n32670 & ~n32674 ;
  assign n32676 = ~n32673 & ~n32675 ;
  assign n32677 = n32668 & n32676 ;
  assign n32681 = \P2_P2_InstAddrPointer_reg[0]/NET0131  & n32197 ;
  assign n32682 = n32178 & n32681 ;
  assign n32683 = ~\P2_P2_InstAddrPointer_reg[23]/NET0131  & ~n32682 ;
  assign n32684 = ~n32576 & ~n32683 ;
  assign n32678 = \P2_P2_InstAddrPointer_reg[22]/NET0131  & ~n32588 ;
  assign n32679 = \P2_P2_InstAddrPointer_reg[0]/NET0131  & n32539 ;
  assign n32680 = ~n32678 & ~n32679 ;
  assign n32685 = \P2_P2_InstAddrPointer_reg[21]/NET0131  & ~n32681 ;
  assign n32686 = ~\P2_P2_InstAddrPointer_reg[21]/NET0131  & n32681 ;
  assign n32687 = ~n32685 & ~n32686 ;
  assign n32688 = ~\P2_P2_InstAddrPointer_reg[20]/NET0131  & ~n32672 ;
  assign n32689 = ~n32681 & ~n32688 ;
  assign n32690 = n32687 & ~n32689 ;
  assign n32691 = n32680 & n32690 ;
  assign n32692 = ~n32684 & n32691 ;
  assign n32693 = n32677 & n32692 ;
  assign n32694 = ~n32578 & n32693 ;
  assign n32695 = ~n32575 & n32694 ;
  assign n32696 = ~\P2_P2_InstAddrPointer_reg[26]/NET0131  & ~n32566 ;
  assign n32697 = ~n32567 & ~n32696 ;
  assign n32698 = n32695 & ~n32697 ;
  assign n32699 = ~\P2_P2_InstAddrPointer_reg[27]/NET0131  & ~n32567 ;
  assign n32700 = \P2_P2_InstAddrPointer_reg[0]/NET0131  & n32203 ;
  assign n32701 = ~n32699 & ~n32700 ;
  assign n32702 = n32698 & ~n32701 ;
  assign n32703 = ~\P2_P2_InstAddrPointer_reg[28]/NET0131  & ~n32700 ;
  assign n32704 = ~n32568 & ~n32703 ;
  assign n32705 = n32702 & ~n32704 ;
  assign n32706 = ~\P2_P2_InstAddrPointer_reg[29]/NET0131  & ~n32568 ;
  assign n32707 = ~n32569 & ~n32706 ;
  assign n32708 = n32705 & ~n32707 ;
  assign n32709 = ~\P2_P2_InstAddrPointer_reg[30]/NET0131  & ~n32569 ;
  assign n32710 = ~n32570 & ~n32709 ;
  assign n32711 = n32708 & ~n32710 ;
  assign n32713 = n32573 & n32711 ;
  assign n32712 = ~n32573 & ~n32711 ;
  assign n32714 = ~n32510 & ~n32712 ;
  assign n32715 = ~n32713 & n32714 ;
  assign n32716 = ~n26629 & ~n32715 ;
  assign n32717 = ~n32563 & n32716 ;
  assign n32718 = ~n32177 & ~n32717 ;
  assign n32719 = n26621 & ~n32718 ;
  assign n32737 = n26757 & n32736 ;
  assign n32738 = n26725 & ~n32559 ;
  assign n32850 = ~n32737 & ~n32738 ;
  assign n32739 = ~n26688 & ~n32573 ;
  assign n32740 = n26640 & ~n26679 ;
  assign n32741 = n26633 & n26640 ;
  assign n32742 = n26620 & ~n32741 ;
  assign n32743 = ~n26645 & n26650 ;
  assign n32744 = n32742 & ~n32743 ;
  assign n32745 = ~n32740 & n32744 ;
  assign n32746 = ~n26729 & n32745 ;
  assign n32747 = \P2_P2_InstAddrPointer_reg[31]/NET0131  & ~n32746 ;
  assign n32851 = ~n32739 & ~n32747 ;
  assign n32852 = n32850 & n32851 ;
  assign n32853 = ~n32719 & n32852 ;
  assign n32854 = ~n32849 & n32853 ;
  assign n32855 = n26792 & ~n32854 ;
  assign n32856 = \P2_P2_rEIP_reg[31]/NET0131  & n28046 ;
  assign n32857 = ~n26285 & n26290 ;
  assign n32858 = ~n26295 & ~n27614 ;
  assign n32859 = ~n32857 & n32858 ;
  assign n32860 = ~n27977 & n32859 ;
  assign n32861 = \P2_P2_InstAddrPointer_reg[31]/NET0131  & ~n32860 ;
  assign n32862 = ~n32856 & ~n32861 ;
  assign n32863 = ~n32855 & n32862 ;
  assign n32872 = \P2_P3_InstAddrPointer_reg[0]/NET0131  & \P2_P3_InstAddrPointer_reg[1]/NET0131  ;
  assign n32873 = ~\P2_P3_InstAddrPointer_reg[2]/NET0131  & ~n32872 ;
  assign n32874 = \P2_P3_InstAddrPointer_reg[3]/NET0131  & ~n32873 ;
  assign n32875 = \P2_P3_InstAddrPointer_reg[4]/NET0131  & n32874 ;
  assign n32876 = \P2_P3_InstAddrPointer_reg[5]/NET0131  & n32875 ;
  assign n32877 = \P2_P3_InstAddrPointer_reg[6]/NET0131  & n32876 ;
  assign n32878 = \P2_P3_InstAddrPointer_reg[7]/NET0131  & n32877 ;
  assign n32879 = \P2_P3_InstAddrPointer_reg[8]/NET0131  & n32878 ;
  assign n32880 = \P2_P3_InstAddrPointer_reg[9]/NET0131  & n32879 ;
  assign n32881 = \P2_P3_InstAddrPointer_reg[10]/NET0131  & n32880 ;
  assign n32882 = \P2_P3_InstAddrPointer_reg[11]/NET0131  & n32881 ;
  assign n32883 = \P2_P3_InstAddrPointer_reg[12]/NET0131  & n32882 ;
  assign n32884 = \P2_P3_InstAddrPointer_reg[13]/NET0131  & \P2_P3_InstAddrPointer_reg[14]/NET0131  ;
  assign n32885 = n32883 & n32884 ;
  assign n32886 = \P2_P3_InstAddrPointer_reg[15]/NET0131  & n32885 ;
  assign n32887 = \P2_P3_InstAddrPointer_reg[16]/NET0131  & n32886 ;
  assign n32888 = \P2_P3_InstAddrPointer_reg[18]/NET0131  & \P2_P3_InstAddrPointer_reg[19]/NET0131  ;
  assign n32889 = \P2_P3_InstAddrPointer_reg[17]/NET0131  & n32888 ;
  assign n32890 = n32887 & n32889 ;
  assign n32891 = \P2_P3_InstAddrPointer_reg[20]/NET0131  & n32890 ;
  assign n32892 = \P2_P3_InstAddrPointer_reg[21]/NET0131  & \P2_P3_InstAddrPointer_reg[22]/NET0131  ;
  assign n32893 = \P2_P3_InstAddrPointer_reg[23]/NET0131  & n32892 ;
  assign n32894 = n32891 & n32893 ;
  assign n32895 = \P2_P3_InstAddrPointer_reg[24]/NET0131  & n32894 ;
  assign n32896 = \P2_P3_InstAddrPointer_reg[25]/NET0131  & n32895 ;
  assign n32897 = \P2_P3_InstAddrPointer_reg[26]/NET0131  & n32896 ;
  assign n32898 = \P2_P3_InstAddrPointer_reg[27]/NET0131  & n32897 ;
  assign n32899 = \P2_P3_InstAddrPointer_reg[28]/NET0131  & n32898 ;
  assign n32900 = \P2_P3_InstAddrPointer_reg[29]/NET0131  & n32899 ;
  assign n32901 = \P2_P3_InstAddrPointer_reg[30]/NET0131  & n32900 ;
  assign n32902 = ~\P2_P3_InstAddrPointer_reg[31]/NET0131  & ~n32901 ;
  assign n32903 = \P2_P3_InstAddrPointer_reg[31]/NET0131  & n32901 ;
  assign n32904 = ~n32902 & ~n32903 ;
  assign n33418 = \P2_P3_InstAddrPointer_reg[21]/NET0131  & n32891 ;
  assign n33419 = \P2_P3_InstAddrPointer_reg[22]/NET0131  & n33418 ;
  assign n33420 = ~\P2_P3_InstAddrPointer_reg[23]/NET0131  & ~n33419 ;
  assign n33421 = ~n32894 & ~n33420 ;
  assign n33422 = \P2_P3_InstAddrPointer_reg[22]/NET0131  & n33421 ;
  assign n33423 = ~\P2_P3_InstAddrPointer_reg[20]/NET0131  & ~n32890 ;
  assign n33424 = ~n32891 & ~n33423 ;
  assign n33425 = ~\P2_P3_InstAddrPointer_reg[15]/NET0131  & ~n32885 ;
  assign n33426 = ~n32886 & ~n33425 ;
  assign n33427 = \P2_P3_InstAddrPointer_reg[13]/NET0131  & n32883 ;
  assign n33428 = ~\P2_P3_InstAddrPointer_reg[13]/NET0131  & ~n32883 ;
  assign n33429 = ~n33427 & ~n33428 ;
  assign n33430 = ~\P2_P3_InstAddrPointer_reg[8]/NET0131  & ~n32878 ;
  assign n33431 = ~n32879 & ~n33430 ;
  assign n33221 = \P2_P3_InstQueue_reg[0][7]/NET0131  & n26837 ;
  assign n33212 = \P2_P3_InstQueue_reg[10][7]/NET0131  & n26833 ;
  assign n33213 = \P2_P3_InstQueue_reg[11][7]/NET0131  & n26819 ;
  assign n33228 = ~n33212 & ~n33213 ;
  assign n33237 = ~n33221 & n33228 ;
  assign n33222 = \P2_P3_InstQueue_reg[8][7]/NET0131  & n26839 ;
  assign n33225 = \P2_P3_InstQueue_reg[15][7]/NET0131  & n26845 ;
  assign n33238 = ~n33222 & ~n33225 ;
  assign n33239 = n33237 & n33238 ;
  assign n33227 = \P2_P3_InstQueue_reg[4][7]/NET0131  & n26847 ;
  assign n33224 = \P2_P3_InstQueue_reg[3][7]/NET0131  & n26843 ;
  assign n33226 = \P2_P3_InstQueue_reg[13][7]/NET0131  & n26829 ;
  assign n33233 = ~n33224 & ~n33226 ;
  assign n33234 = ~n33227 & n33233 ;
  assign n33218 = \P2_P3_InstQueue_reg[5][7]/NET0131  & n26815 ;
  assign n33219 = \P2_P3_InstQueue_reg[12][7]/NET0131  & n26849 ;
  assign n33231 = ~n33218 & ~n33219 ;
  assign n33220 = \P2_P3_InstQueue_reg[9][7]/NET0131  & n26827 ;
  assign n33223 = \P2_P3_InstQueue_reg[7][7]/NET0131  & n26841 ;
  assign n33232 = ~n33220 & ~n33223 ;
  assign n33235 = n33231 & n33232 ;
  assign n33214 = \P2_P3_InstQueue_reg[1][7]/NET0131  & n26812 ;
  assign n33215 = \P2_P3_InstQueue_reg[6][7]/NET0131  & n26822 ;
  assign n33229 = ~n33214 & ~n33215 ;
  assign n33216 = \P2_P3_InstQueue_reg[14][7]/NET0131  & n26825 ;
  assign n33217 = \P2_P3_InstQueue_reg[2][7]/NET0131  & n26831 ;
  assign n33230 = ~n33216 & ~n33217 ;
  assign n33236 = n33229 & n33230 ;
  assign n33240 = n33235 & n33236 ;
  assign n33241 = n33234 & n33240 ;
  assign n33242 = n33239 & n33241 ;
  assign n33432 = ~\P2_P3_InstAddrPointer_reg[7]/NET0131  & ~n32877 ;
  assign n33433 = ~n32878 & ~n33432 ;
  assign n33434 = ~n33242 & n33433 ;
  assign n33435 = n33242 & ~n33433 ;
  assign n32969 = \P2_P3_InstQueue_reg[0][6]/NET0131  & n26837 ;
  assign n32960 = \P2_P3_InstQueue_reg[2][6]/NET0131  & n26831 ;
  assign n32961 = \P2_P3_InstQueue_reg[11][6]/NET0131  & n26819 ;
  assign n32976 = ~n32960 & ~n32961 ;
  assign n32985 = ~n32969 & n32976 ;
  assign n32970 = \P2_P3_InstQueue_reg[8][6]/NET0131  & n26839 ;
  assign n32973 = \P2_P3_InstQueue_reg[15][6]/NET0131  & n26845 ;
  assign n32986 = ~n32970 & ~n32973 ;
  assign n32987 = n32985 & n32986 ;
  assign n32975 = \P2_P3_InstQueue_reg[4][6]/NET0131  & n26847 ;
  assign n32972 = \P2_P3_InstQueue_reg[5][6]/NET0131  & n26815 ;
  assign n32974 = \P2_P3_InstQueue_reg[10][6]/NET0131  & n26833 ;
  assign n32981 = ~n32972 & ~n32974 ;
  assign n32982 = ~n32975 & n32981 ;
  assign n32966 = \P2_P3_InstQueue_reg[1][6]/NET0131  & n26812 ;
  assign n32967 = \P2_P3_InstQueue_reg[13][6]/NET0131  & n26829 ;
  assign n32979 = ~n32966 & ~n32967 ;
  assign n32968 = \P2_P3_InstQueue_reg[12][6]/NET0131  & n26849 ;
  assign n32971 = \P2_P3_InstQueue_reg[7][6]/NET0131  & n26841 ;
  assign n32980 = ~n32968 & ~n32971 ;
  assign n32983 = n32979 & n32980 ;
  assign n32962 = \P2_P3_InstQueue_reg[9][6]/NET0131  & n26827 ;
  assign n32963 = \P2_P3_InstQueue_reg[6][6]/NET0131  & n26822 ;
  assign n32977 = ~n32962 & ~n32963 ;
  assign n32964 = \P2_P3_InstQueue_reg[14][6]/NET0131  & n26825 ;
  assign n32965 = \P2_P3_InstQueue_reg[3][6]/NET0131  & n26843 ;
  assign n32978 = ~n32964 & ~n32965 ;
  assign n32984 = n32977 & n32978 ;
  assign n32988 = n32983 & n32984 ;
  assign n32989 = n32982 & n32988 ;
  assign n32990 = n32987 & n32989 ;
  assign n33436 = ~\P2_P3_InstAddrPointer_reg[6]/NET0131  & ~n32876 ;
  assign n33437 = ~n32877 & ~n33436 ;
  assign n33438 = ~n32990 & n33437 ;
  assign n33439 = n32990 & ~n33437 ;
  assign n33003 = \P2_P3_InstQueue_reg[15][5]/NET0131  & n26845 ;
  assign n32995 = \P2_P3_InstQueue_reg[9][5]/NET0131  & n26827 ;
  assign n32996 = \P2_P3_InstQueue_reg[10][5]/NET0131  & n26833 ;
  assign n33011 = ~n32995 & ~n32996 ;
  assign n33020 = ~n33003 & n33011 ;
  assign n33005 = \P2_P3_InstQueue_reg[0][5]/NET0131  & n26837 ;
  assign n33006 = \P2_P3_InstQueue_reg[8][5]/NET0131  & n26839 ;
  assign n33021 = ~n33005 & ~n33006 ;
  assign n33022 = n33020 & n33021 ;
  assign n33010 = \P2_P3_InstQueue_reg[5][5]/NET0131  & n26815 ;
  assign n33008 = \P2_P3_InstQueue_reg[6][5]/NET0131  & n26822 ;
  assign n33009 = \P2_P3_InstQueue_reg[4][5]/NET0131  & n26847 ;
  assign n33016 = ~n33008 & ~n33009 ;
  assign n33017 = ~n33010 & n33016 ;
  assign n33001 = \P2_P3_InstQueue_reg[2][5]/NET0131  & n26831 ;
  assign n33002 = \P2_P3_InstQueue_reg[11][5]/NET0131  & n26819 ;
  assign n33014 = ~n33001 & ~n33002 ;
  assign n33004 = \P2_P3_InstQueue_reg[7][5]/NET0131  & n26841 ;
  assign n33007 = \P2_P3_InstQueue_reg[12][5]/NET0131  & n26849 ;
  assign n33015 = ~n33004 & ~n33007 ;
  assign n33018 = n33014 & n33015 ;
  assign n32997 = \P2_P3_InstQueue_reg[3][5]/NET0131  & n26843 ;
  assign n32998 = \P2_P3_InstQueue_reg[1][5]/NET0131  & n26812 ;
  assign n33012 = ~n32997 & ~n32998 ;
  assign n32999 = \P2_P3_InstQueue_reg[13][5]/NET0131  & n26829 ;
  assign n33000 = \P2_P3_InstQueue_reg[14][5]/NET0131  & n26825 ;
  assign n33013 = ~n32999 & ~n33000 ;
  assign n33019 = n33012 & n33013 ;
  assign n33023 = n33018 & n33019 ;
  assign n33024 = n33017 & n33023 ;
  assign n33025 = n33022 & n33024 ;
  assign n33440 = ~\P2_P3_InstAddrPointer_reg[5]/NET0131  & ~n32875 ;
  assign n33441 = ~n32876 & ~n33440 ;
  assign n33442 = ~n33025 & n33441 ;
  assign n33443 = n33025 & ~n33441 ;
  assign n33039 = \P2_P3_InstQueue_reg[0][4]/NET0131  & n26837 ;
  assign n33030 = \P2_P3_InstQueue_reg[2][4]/NET0131  & n26831 ;
  assign n33031 = \P2_P3_InstQueue_reg[11][4]/NET0131  & n26819 ;
  assign n33046 = ~n33030 & ~n33031 ;
  assign n33055 = ~n33039 & n33046 ;
  assign n33040 = \P2_P3_InstQueue_reg[8][4]/NET0131  & n26839 ;
  assign n33043 = \P2_P3_InstQueue_reg[15][4]/NET0131  & n26845 ;
  assign n33056 = ~n33040 & ~n33043 ;
  assign n33057 = n33055 & n33056 ;
  assign n33045 = \P2_P3_InstQueue_reg[4][4]/NET0131  & n26847 ;
  assign n33042 = \P2_P3_InstQueue_reg[5][4]/NET0131  & n26815 ;
  assign n33044 = \P2_P3_InstQueue_reg[10][4]/NET0131  & n26833 ;
  assign n33051 = ~n33042 & ~n33044 ;
  assign n33052 = ~n33045 & n33051 ;
  assign n33036 = \P2_P3_InstQueue_reg[1][4]/NET0131  & n26812 ;
  assign n33037 = \P2_P3_InstQueue_reg[13][4]/NET0131  & n26829 ;
  assign n33049 = ~n33036 & ~n33037 ;
  assign n33038 = \P2_P3_InstQueue_reg[12][4]/NET0131  & n26849 ;
  assign n33041 = \P2_P3_InstQueue_reg[7][4]/NET0131  & n26841 ;
  assign n33050 = ~n33038 & ~n33041 ;
  assign n33053 = n33049 & n33050 ;
  assign n33032 = \P2_P3_InstQueue_reg[9][4]/NET0131  & n26827 ;
  assign n33033 = \P2_P3_InstQueue_reg[6][4]/NET0131  & n26822 ;
  assign n33047 = ~n33032 & ~n33033 ;
  assign n33034 = \P2_P3_InstQueue_reg[14][4]/NET0131  & n26825 ;
  assign n33035 = \P2_P3_InstQueue_reg[3][4]/NET0131  & n26843 ;
  assign n33048 = ~n33034 & ~n33035 ;
  assign n33054 = n33047 & n33048 ;
  assign n33058 = n33053 & n33054 ;
  assign n33059 = n33052 & n33058 ;
  assign n33060 = n33057 & n33059 ;
  assign n33444 = ~\P2_P3_InstAddrPointer_reg[4]/NET0131  & ~n32874 ;
  assign n33445 = ~n32875 & ~n33444 ;
  assign n33446 = ~n33060 & n33445 ;
  assign n33447 = n33060 & ~n33445 ;
  assign n33073 = \P2_P3_InstQueue_reg[15][3]/NET0131  & n26845 ;
  assign n33065 = \P2_P3_InstQueue_reg[14][3]/NET0131  & n26825 ;
  assign n33066 = \P2_P3_InstQueue_reg[6][3]/NET0131  & n26822 ;
  assign n33081 = ~n33065 & ~n33066 ;
  assign n33090 = ~n33073 & n33081 ;
  assign n33075 = \P2_P3_InstQueue_reg[0][3]/NET0131  & n26837 ;
  assign n33076 = \P2_P3_InstQueue_reg[8][3]/NET0131  & n26839 ;
  assign n33091 = ~n33075 & ~n33076 ;
  assign n33092 = n33090 & n33091 ;
  assign n33080 = \P2_P3_InstQueue_reg[2][3]/NET0131  & n26831 ;
  assign n33078 = \P2_P3_InstQueue_reg[10][3]/NET0131  & n26833 ;
  assign n33079 = \P2_P3_InstQueue_reg[13][3]/NET0131  & n26829 ;
  assign n33086 = ~n33078 & ~n33079 ;
  assign n33087 = ~n33080 & n33086 ;
  assign n33071 = \P2_P3_InstQueue_reg[1][3]/NET0131  & n26812 ;
  assign n33072 = \P2_P3_InstQueue_reg[11][3]/NET0131  & n26819 ;
  assign n33084 = ~n33071 & ~n33072 ;
  assign n33074 = \P2_P3_InstQueue_reg[7][3]/NET0131  & n26841 ;
  assign n33077 = \P2_P3_InstQueue_reg[12][3]/NET0131  & n26849 ;
  assign n33085 = ~n33074 & ~n33077 ;
  assign n33088 = n33084 & n33085 ;
  assign n33067 = \P2_P3_InstQueue_reg[3][3]/NET0131  & n26843 ;
  assign n33068 = \P2_P3_InstQueue_reg[5][3]/NET0131  & n26815 ;
  assign n33082 = ~n33067 & ~n33068 ;
  assign n33069 = \P2_P3_InstQueue_reg[4][3]/NET0131  & n26847 ;
  assign n33070 = \P2_P3_InstQueue_reg[9][3]/NET0131  & n26827 ;
  assign n33083 = ~n33069 & ~n33070 ;
  assign n33089 = n33082 & n33083 ;
  assign n33093 = n33088 & n33089 ;
  assign n33094 = n33087 & n33093 ;
  assign n33095 = n33092 & n33094 ;
  assign n33448 = ~\P2_P3_InstAddrPointer_reg[3]/NET0131  & n32873 ;
  assign n33449 = ~n32874 & ~n33448 ;
  assign n33450 = ~n33095 & n33449 ;
  assign n33451 = n33095 & ~n33449 ;
  assign n33109 = \P2_P3_InstQueue_reg[0][2]/NET0131  & n26837 ;
  assign n33100 = \P2_P3_InstQueue_reg[2][2]/NET0131  & n26831 ;
  assign n33101 = \P2_P3_InstQueue_reg[3][2]/NET0131  & n26843 ;
  assign n33116 = ~n33100 & ~n33101 ;
  assign n33125 = ~n33109 & n33116 ;
  assign n33110 = \P2_P3_InstQueue_reg[8][2]/NET0131  & n26839 ;
  assign n33113 = \P2_P3_InstQueue_reg[15][2]/NET0131  & n26845 ;
  assign n33126 = ~n33110 & ~n33113 ;
  assign n33127 = n33125 & n33126 ;
  assign n33115 = \P2_P3_InstQueue_reg[13][2]/NET0131  & n26829 ;
  assign n33112 = \P2_P3_InstQueue_reg[4][2]/NET0131  & n26847 ;
  assign n33114 = \P2_P3_InstQueue_reg[14][2]/NET0131  & n26825 ;
  assign n33121 = ~n33112 & ~n33114 ;
  assign n33122 = ~n33115 & n33121 ;
  assign n33106 = \P2_P3_InstQueue_reg[12][2]/NET0131  & n26849 ;
  assign n33107 = \P2_P3_InstQueue_reg[11][2]/NET0131  & n26819 ;
  assign n33119 = ~n33106 & ~n33107 ;
  assign n33108 = \P2_P3_InstQueue_reg[9][2]/NET0131  & n26827 ;
  assign n33111 = \P2_P3_InstQueue_reg[7][2]/NET0131  & n26841 ;
  assign n33120 = ~n33108 & ~n33111 ;
  assign n33123 = n33119 & n33120 ;
  assign n33102 = \P2_P3_InstQueue_reg[10][2]/NET0131  & n26833 ;
  assign n33103 = \P2_P3_InstQueue_reg[5][2]/NET0131  & n26815 ;
  assign n33117 = ~n33102 & ~n33103 ;
  assign n33104 = \P2_P3_InstQueue_reg[1][2]/NET0131  & n26812 ;
  assign n33105 = \P2_P3_InstQueue_reg[6][2]/NET0131  & n26822 ;
  assign n33118 = ~n33104 & ~n33105 ;
  assign n33124 = n33117 & n33118 ;
  assign n33128 = n33123 & n33124 ;
  assign n33129 = n33122 & n33128 ;
  assign n33130 = n33127 & n33129 ;
  assign n33306 = \P2_P3_InstAddrPointer_reg[2]/NET0131  & n32872 ;
  assign n33311 = ~n32873 & ~n33306 ;
  assign n33452 = ~n33130 & ~n33311 ;
  assign n33453 = n33130 & n33311 ;
  assign n33134 = \P2_P3_InstQueue_reg[15][1]/NET0131  & n26845 ;
  assign n33133 = \P2_P3_InstQueue_reg[10][1]/NET0131  & n26833 ;
  assign n33135 = \P2_P3_InstQueue_reg[9][1]/NET0131  & n26827 ;
  assign n33149 = ~n33133 & ~n33135 ;
  assign n33158 = ~n33134 & n33149 ;
  assign n33138 = \P2_P3_InstQueue_reg[0][1]/NET0131  & n26837 ;
  assign n33142 = \P2_P3_InstQueue_reg[8][1]/NET0131  & n26839 ;
  assign n33159 = ~n33138 & ~n33142 ;
  assign n33160 = n33158 & n33159 ;
  assign n33148 = \P2_P3_InstQueue_reg[6][1]/NET0131  & n26822 ;
  assign n33146 = \P2_P3_InstQueue_reg[1][1]/NET0131  & n26812 ;
  assign n33147 = \P2_P3_InstQueue_reg[3][1]/NET0131  & n26843 ;
  assign n33154 = ~n33146 & ~n33147 ;
  assign n33155 = ~n33148 & n33154 ;
  assign n33141 = \P2_P3_InstQueue_reg[4][1]/NET0131  & n26847 ;
  assign n33143 = \P2_P3_InstQueue_reg[11][1]/NET0131  & n26819 ;
  assign n33152 = ~n33141 & ~n33143 ;
  assign n33144 = \P2_P3_InstQueue_reg[14][1]/NET0131  & n26825 ;
  assign n33145 = \P2_P3_InstQueue_reg[13][1]/NET0131  & n26829 ;
  assign n33153 = ~n33144 & ~n33145 ;
  assign n33156 = n33152 & n33153 ;
  assign n33136 = \P2_P3_InstQueue_reg[12][1]/NET0131  & n26849 ;
  assign n33137 = \P2_P3_InstQueue_reg[5][1]/NET0131  & n26815 ;
  assign n33150 = ~n33136 & ~n33137 ;
  assign n33139 = \P2_P3_InstQueue_reg[7][1]/NET0131  & n26841 ;
  assign n33140 = \P2_P3_InstQueue_reg[2][1]/NET0131  & n26831 ;
  assign n33151 = ~n33139 & ~n33140 ;
  assign n33157 = n33150 & n33151 ;
  assign n33161 = n33156 & n33157 ;
  assign n33162 = n33155 & n33161 ;
  assign n33163 = n33160 & n33162 ;
  assign n33314 = ~\P2_P3_InstAddrPointer_reg[0]/NET0131  & \P2_P3_InstAddrPointer_reg[1]/NET0131  ;
  assign n33454 = \P2_P3_InstAddrPointer_reg[0]/NET0131  & ~\P2_P3_InstAddrPointer_reg[1]/NET0131  ;
  assign n33455 = ~n33314 & ~n33454 ;
  assign n33456 = ~n33163 & ~n33455 ;
  assign n33457 = n33163 & n33455 ;
  assign n33167 = \P2_P3_InstQueue_reg[15][0]/NET0131  & n26845 ;
  assign n33166 = \P2_P3_InstQueue_reg[6][0]/NET0131  & n26822 ;
  assign n33168 = \P2_P3_InstQueue_reg[11][0]/NET0131  & n26819 ;
  assign n33182 = ~n33166 & ~n33168 ;
  assign n33191 = ~n33167 & n33182 ;
  assign n33171 = \P2_P3_InstQueue_reg[0][0]/NET0131  & n26837 ;
  assign n33175 = \P2_P3_InstQueue_reg[8][0]/NET0131  & n26839 ;
  assign n33192 = ~n33171 & ~n33175 ;
  assign n33193 = n33191 & n33192 ;
  assign n33181 = \P2_P3_InstQueue_reg[5][0]/NET0131  & n26815 ;
  assign n33179 = \P2_P3_InstQueue_reg[4][0]/NET0131  & n26847 ;
  assign n33180 = \P2_P3_InstQueue_reg[12][0]/NET0131  & n26849 ;
  assign n33187 = ~n33179 & ~n33180 ;
  assign n33188 = ~n33181 & n33187 ;
  assign n33174 = \P2_P3_InstQueue_reg[3][0]/NET0131  & n26843 ;
  assign n33176 = \P2_P3_InstQueue_reg[14][0]/NET0131  & n26825 ;
  assign n33185 = ~n33174 & ~n33176 ;
  assign n33177 = \P2_P3_InstQueue_reg[9][0]/NET0131  & n26827 ;
  assign n33178 = \P2_P3_InstQueue_reg[1][0]/NET0131  & n26812 ;
  assign n33186 = ~n33177 & ~n33178 ;
  assign n33189 = n33185 & n33186 ;
  assign n33169 = \P2_P3_InstQueue_reg[13][0]/NET0131  & n26829 ;
  assign n33170 = \P2_P3_InstQueue_reg[10][0]/NET0131  & n26833 ;
  assign n33183 = ~n33169 & ~n33170 ;
  assign n33172 = \P2_P3_InstQueue_reg[7][0]/NET0131  & n26841 ;
  assign n33173 = \P2_P3_InstQueue_reg[2][0]/NET0131  & n26831 ;
  assign n33184 = ~n33172 & ~n33173 ;
  assign n33190 = n33183 & n33184 ;
  assign n33194 = n33189 & n33190 ;
  assign n33195 = n33188 & n33194 ;
  assign n33196 = n33193 & n33195 ;
  assign n33458 = ~\P2_P3_InstAddrPointer_reg[0]/NET0131  & ~n33196 ;
  assign n33459 = ~n33457 & n33458 ;
  assign n33460 = ~n33456 & ~n33459 ;
  assign n33461 = ~n33453 & ~n33460 ;
  assign n33462 = ~n33452 & ~n33461 ;
  assign n33463 = ~n33451 & ~n33462 ;
  assign n33464 = ~n33450 & ~n33463 ;
  assign n33465 = ~n33447 & ~n33464 ;
  assign n33466 = ~n33446 & ~n33465 ;
  assign n33467 = ~n33443 & ~n33466 ;
  assign n33468 = ~n33442 & ~n33467 ;
  assign n33469 = ~n33439 & ~n33468 ;
  assign n33470 = ~n33438 & ~n33469 ;
  assign n33471 = ~n33435 & ~n33470 ;
  assign n33472 = ~n33434 & ~n33471 ;
  assign n33473 = n33431 & ~n33472 ;
  assign n33474 = \P2_P3_InstAddrPointer_reg[9]/NET0131  & n33473 ;
  assign n33475 = ~\P2_P3_InstAddrPointer_reg[10]/NET0131  & ~n32880 ;
  assign n33476 = ~n32881 & ~n33475 ;
  assign n33477 = n33474 & n33476 ;
  assign n33478 = \P2_P3_InstAddrPointer_reg[11]/NET0131  & n33477 ;
  assign n33479 = \P2_P3_InstAddrPointer_reg[12]/NET0131  & n33478 ;
  assign n33480 = n33429 & n33479 ;
  assign n33481 = \P2_P3_InstAddrPointer_reg[14]/NET0131  & n33480 ;
  assign n33482 = n33426 & n33481 ;
  assign n33483 = \P2_P3_InstAddrPointer_reg[16]/NET0131  & n33482 ;
  assign n33484 = \P2_P3_InstAddrPointer_reg[17]/NET0131  & n32887 ;
  assign n33485 = ~\P2_P3_InstAddrPointer_reg[17]/NET0131  & ~n32887 ;
  assign n33486 = ~n33484 & ~n33485 ;
  assign n33487 = n32888 & n33486 ;
  assign n33488 = n33483 & n33487 ;
  assign n33489 = n33424 & n33488 ;
  assign n33490 = \P2_P3_InstAddrPointer_reg[21]/NET0131  & n33489 ;
  assign n33491 = n33422 & n33490 ;
  assign n33492 = \P2_P3_InstAddrPointer_reg[24]/NET0131  & n33491 ;
  assign n32906 = \P2_P3_InstAddrPointer_reg[26]/NET0131  & \P2_P3_InstAddrPointer_reg[27]/NET0131  ;
  assign n33493 = ~\P2_P3_InstAddrPointer_reg[25]/NET0131  & ~n32895 ;
  assign n33494 = ~n32896 & ~n33493 ;
  assign n33495 = n32906 & n33494 ;
  assign n33496 = n33492 & n33495 ;
  assign n33497 = ~\P2_P3_InstAddrPointer_reg[28]/NET0131  & ~n32898 ;
  assign n33498 = ~n32899 & ~n33497 ;
  assign n33499 = n33496 & n33498 ;
  assign n33500 = \P2_P3_InstAddrPointer_reg[29]/NET0131  & n33499 ;
  assign n33501 = \P2_P3_InstAddrPointer_reg[30]/NET0131  & n33500 ;
  assign n33503 = ~n32904 & ~n33501 ;
  assign n33502 = \P2_P3_InstAddrPointer_reg[31]/NET0131  & n33501 ;
  assign n33504 = n27280 & ~n33502 ;
  assign n33505 = ~n33503 & n33504 ;
  assign n32907 = \P2_P3_InstAddrPointer_reg[24]/NET0131  & n32893 ;
  assign n32908 = \P2_P3_InstAddrPointer_reg[1]/NET0131  & \P2_P3_InstAddrPointer_reg[2]/NET0131  ;
  assign n32909 = \P2_P3_InstAddrPointer_reg[3]/NET0131  & n32908 ;
  assign n32910 = \P2_P3_InstAddrPointer_reg[4]/NET0131  & n32909 ;
  assign n32911 = \P2_P3_InstAddrPointer_reg[5]/NET0131  & n32910 ;
  assign n32912 = \P2_P3_InstAddrPointer_reg[6]/NET0131  & n32911 ;
  assign n32913 = \P2_P3_InstAddrPointer_reg[7]/NET0131  & n32912 ;
  assign n32914 = \P2_P3_InstAddrPointer_reg[8]/NET0131  & n32913 ;
  assign n32915 = \P2_P3_InstAddrPointer_reg[9]/NET0131  & n32914 ;
  assign n32916 = \P2_P3_InstAddrPointer_reg[10]/NET0131  & n32915 ;
  assign n32917 = \P2_P3_InstAddrPointer_reg[11]/NET0131  & n32916 ;
  assign n32918 = \P2_P3_InstAddrPointer_reg[12]/NET0131  & n32917 ;
  assign n32919 = n32884 & n32918 ;
  assign n32920 = \P2_P3_InstAddrPointer_reg[15]/NET0131  & n32919 ;
  assign n32921 = \P2_P3_InstAddrPointer_reg[16]/NET0131  & n32920 ;
  assign n32922 = n32889 & n32921 ;
  assign n32923 = \P2_P3_InstAddrPointer_reg[20]/NET0131  & n32922 ;
  assign n32924 = n32907 & n32923 ;
  assign n32925 = \P2_P3_InstAddrPointer_reg[25]/NET0131  & n32924 ;
  assign n32948 = ~\P2_P3_InstAddrPointer_reg[25]/NET0131  & ~n32924 ;
  assign n32949 = ~n32925 & ~n32948 ;
  assign n32950 = n32906 & n32949 ;
  assign n32951 = ~\P2_P3_InstAddrPointer_reg[15]/NET0131  & ~n32919 ;
  assign n32952 = ~n32920 & ~n32951 ;
  assign n32953 = \P2_P3_InstAddrPointer_reg[13]/NET0131  & n32918 ;
  assign n32954 = ~\P2_P3_InstAddrPointer_reg[13]/NET0131  & ~n32918 ;
  assign n32955 = ~n32953 & ~n32954 ;
  assign n32956 = ~\P2_P3_InstAddrPointer_reg[7]/NET0131  & ~n32912 ;
  assign n32957 = ~n32913 & ~n32956 ;
  assign n32958 = ~\P2_P3_InstAddrPointer_reg[6]/NET0131  & ~n32911 ;
  assign n32959 = ~n32912 & ~n32958 ;
  assign n32991 = n32959 & ~n32990 ;
  assign n32992 = ~n32959 & n32990 ;
  assign n32993 = ~\P2_P3_InstAddrPointer_reg[5]/NET0131  & ~n32910 ;
  assign n32994 = ~n32911 & ~n32993 ;
  assign n33026 = n32994 & ~n33025 ;
  assign n33027 = ~n32994 & n33025 ;
  assign n33028 = ~\P2_P3_InstAddrPointer_reg[4]/NET0131  & ~n32909 ;
  assign n33029 = ~n32910 & ~n33028 ;
  assign n33061 = n33029 & ~n33060 ;
  assign n33062 = ~n33029 & n33060 ;
  assign n33063 = ~\P2_P3_InstAddrPointer_reg[3]/NET0131  & ~n32908 ;
  assign n33064 = ~n32909 & ~n33063 ;
  assign n33096 = n33064 & ~n33095 ;
  assign n33097 = ~n33064 & n33095 ;
  assign n33098 = ~\P2_P3_InstAddrPointer_reg[1]/NET0131  & ~\P2_P3_InstAddrPointer_reg[2]/NET0131  ;
  assign n33099 = ~n32908 & ~n33098 ;
  assign n33131 = n33099 & ~n33130 ;
  assign n33132 = ~n33099 & n33130 ;
  assign n33164 = ~\P2_P3_InstAddrPointer_reg[1]/NET0131  & ~n33163 ;
  assign n33165 = \P2_P3_InstAddrPointer_reg[1]/NET0131  & n33163 ;
  assign n33197 = \P2_P3_InstAddrPointer_reg[0]/NET0131  & ~n33196 ;
  assign n33198 = ~n33165 & n33197 ;
  assign n33199 = ~n33164 & ~n33198 ;
  assign n33200 = ~n33132 & ~n33199 ;
  assign n33201 = ~n33131 & ~n33200 ;
  assign n33202 = ~n33097 & ~n33201 ;
  assign n33203 = ~n33096 & ~n33202 ;
  assign n33204 = ~n33062 & ~n33203 ;
  assign n33205 = ~n33061 & ~n33204 ;
  assign n33206 = ~n33027 & ~n33205 ;
  assign n33207 = ~n33026 & ~n33206 ;
  assign n33208 = ~n32992 & ~n33207 ;
  assign n33209 = ~n32991 & ~n33208 ;
  assign n33210 = n32957 & ~n33209 ;
  assign n33211 = ~n32957 & n33209 ;
  assign n33243 = ~n33211 & ~n33242 ;
  assign n33244 = ~n33210 & ~n33243 ;
  assign n33245 = ~\P2_P3_InstAddrPointer_reg[8]/NET0131  & ~n32913 ;
  assign n33246 = ~n32914 & ~n33245 ;
  assign n33247 = ~n33244 & n33246 ;
  assign n33248 = \P2_P3_InstAddrPointer_reg[9]/NET0131  & n33247 ;
  assign n33249 = ~\P2_P3_InstAddrPointer_reg[10]/NET0131  & ~n32915 ;
  assign n33250 = ~n32916 & ~n33249 ;
  assign n33251 = n33248 & n33250 ;
  assign n33252 = \P2_P3_InstAddrPointer_reg[11]/NET0131  & n33251 ;
  assign n33253 = \P2_P3_InstAddrPointer_reg[12]/NET0131  & n33252 ;
  assign n33254 = n32955 & n33253 ;
  assign n33255 = \P2_P3_InstAddrPointer_reg[14]/NET0131  & n33254 ;
  assign n33256 = n32952 & n33255 ;
  assign n33257 = ~\P2_P3_InstAddrPointer_reg[16]/NET0131  & ~n32920 ;
  assign n33258 = ~n32921 & ~n33257 ;
  assign n33259 = n32889 & n33258 ;
  assign n33260 = n33256 & n33259 ;
  assign n33261 = ~\P2_P3_InstAddrPointer_reg[20]/NET0131  & ~n32922 ;
  assign n33262 = ~n32923 & ~n33261 ;
  assign n33263 = n33260 & n33262 ;
  assign n33264 = n32907 & n33263 ;
  assign n33265 = n32950 & n33264 ;
  assign n32926 = n32906 & n32925 ;
  assign n32927 = \P2_P3_InstAddrPointer_reg[28]/NET0131  & n32926 ;
  assign n33266 = ~\P2_P3_InstAddrPointer_reg[28]/NET0131  & ~n32926 ;
  assign n33267 = ~n32927 & ~n33266 ;
  assign n33268 = n33265 & n33267 ;
  assign n33269 = \P2_P3_InstAddrPointer_reg[29]/NET0131  & n33268 ;
  assign n33270 = \P2_P3_InstAddrPointer_reg[30]/NET0131  & n33269 ;
  assign n33272 = \P2_P3_InstAddrPointer_reg[31]/NET0131  & n33270 ;
  assign n32928 = \P2_P3_InstAddrPointer_reg[29]/NET0131  & n32927 ;
  assign n32935 = \P2_P3_InstAddrPointer_reg[30]/NET0131  & n32928 ;
  assign n32936 = ~\P2_P3_InstAddrPointer_reg[31]/NET0131  & ~n32935 ;
  assign n32937 = \P2_P3_InstAddrPointer_reg[31]/NET0131  & n32935 ;
  assign n32938 = ~n32936 & ~n32937 ;
  assign n33271 = ~n32938 & ~n33270 ;
  assign n33273 = n33242 & ~n33271 ;
  assign n33274 = ~n33272 & n33273 ;
  assign n32929 = \P2_P3_InstAddrPointer_reg[0]/NET0131  & n32928 ;
  assign n32930 = \P2_P3_InstAddrPointer_reg[30]/NET0131  & n32929 ;
  assign n32931 = \P2_P3_InstAddrPointer_reg[31]/NET0131  & ~n32930 ;
  assign n32932 = ~\P2_P3_InstAddrPointer_reg[31]/NET0131  & n32930 ;
  assign n32933 = ~n32931 & ~n32932 ;
  assign n33275 = \P2_P3_InstAddrPointer_reg[0]/NET0131  & n32923 ;
  assign n33276 = n32892 & n33275 ;
  assign n33277 = ~\P2_P3_InstAddrPointer_reg[23]/NET0131  & ~n33276 ;
  assign n33278 = n32893 & n33275 ;
  assign n33279 = ~n33277 & ~n33278 ;
  assign n33280 = \P2_P3_InstAddrPointer_reg[0]/NET0131  & n32913 ;
  assign n33281 = \P2_P3_InstAddrPointer_reg[8]/NET0131  & n33280 ;
  assign n33282 = \P2_P3_InstAddrPointer_reg[9]/NET0131  & n33281 ;
  assign n33283 = \P2_P3_InstAddrPointer_reg[10]/NET0131  & n33282 ;
  assign n33284 = ~\P2_P3_InstAddrPointer_reg[11]/NET0131  & ~n33283 ;
  assign n33285 = \P2_P3_InstAddrPointer_reg[11]/NET0131  & n33283 ;
  assign n33286 = ~n33284 & ~n33285 ;
  assign n33287 = \P2_P3_InstAddrPointer_reg[0]/NET0131  & n32912 ;
  assign n33288 = ~\P2_P3_InstAddrPointer_reg[7]/NET0131  & ~n33287 ;
  assign n33289 = ~n33280 & ~n33288 ;
  assign n33290 = \P2_P3_InstAddrPointer_reg[0]/NET0131  & n32911 ;
  assign n33291 = ~\P2_P3_InstAddrPointer_reg[6]/NET0131  & ~n33290 ;
  assign n33292 = ~n33287 & ~n33291 ;
  assign n33293 = n32990 & ~n33292 ;
  assign n33294 = \P2_P3_InstAddrPointer_reg[0]/NET0131  & n32910 ;
  assign n33295 = ~\P2_P3_InstAddrPointer_reg[5]/NET0131  & ~n33294 ;
  assign n33296 = ~n33290 & ~n33295 ;
  assign n33299 = n33025 & ~n33296 ;
  assign n33300 = ~n33293 & ~n33299 ;
  assign n33301 = \P2_P3_InstAddrPointer_reg[0]/NET0131  & n32909 ;
  assign n33302 = ~\P2_P3_InstAddrPointer_reg[4]/NET0131  & ~n33301 ;
  assign n33303 = ~n33294 & ~n33302 ;
  assign n33304 = n33060 & ~n33303 ;
  assign n33305 = ~n33060 & n33303 ;
  assign n33307 = ~\P2_P3_InstAddrPointer_reg[3]/NET0131  & ~n33306 ;
  assign n33308 = ~n33301 & ~n33307 ;
  assign n33309 = n33095 & ~n33308 ;
  assign n33310 = ~n33095 & n33308 ;
  assign n33312 = ~n33130 & n33311 ;
  assign n33313 = n33130 & ~n33311 ;
  assign n33315 = n33199 & ~n33314 ;
  assign n33316 = ~n33313 & ~n33315 ;
  assign n33317 = ~n33312 & ~n33316 ;
  assign n33318 = ~n33310 & n33317 ;
  assign n33319 = ~n33309 & ~n33318 ;
  assign n33320 = ~n33305 & ~n33319 ;
  assign n33321 = ~n33304 & ~n33320 ;
  assign n33322 = n33300 & n33321 ;
  assign n33297 = ~n33025 & n33296 ;
  assign n33298 = ~n33293 & n33297 ;
  assign n33323 = ~n32990 & n33292 ;
  assign n33324 = ~n33298 & ~n33323 ;
  assign n33325 = ~n33322 & n33324 ;
  assign n33326 = ~n33289 & n33325 ;
  assign n33327 = ~n33242 & ~n33326 ;
  assign n33328 = n33289 & ~n33325 ;
  assign n33329 = ~\P2_P3_InstAddrPointer_reg[8]/NET0131  & ~n33280 ;
  assign n33330 = ~n33281 & ~n33329 ;
  assign n33331 = ~n33328 & ~n33330 ;
  assign n33332 = ~n33327 & n33331 ;
  assign n33333 = ~\P2_P3_InstAddrPointer_reg[9]/NET0131  & ~n33281 ;
  assign n33334 = ~n33282 & ~n33333 ;
  assign n33335 = ~\P2_P3_InstAddrPointer_reg[10]/NET0131  & ~n33282 ;
  assign n33336 = ~n33283 & ~n33335 ;
  assign n33337 = ~n33334 & ~n33336 ;
  assign n33338 = n33332 & n33337 ;
  assign n33339 = ~n33286 & n33338 ;
  assign n33340 = ~\P2_P3_InstAddrPointer_reg[12]/NET0131  & ~n33285 ;
  assign n33341 = \P2_P3_InstAddrPointer_reg[12]/NET0131  & n33285 ;
  assign n33342 = ~n33340 & ~n33341 ;
  assign n33343 = n33339 & ~n33342 ;
  assign n33344 = ~\P2_P3_InstAddrPointer_reg[13]/NET0131  & ~n33341 ;
  assign n33345 = \P2_P3_InstAddrPointer_reg[13]/NET0131  & n33341 ;
  assign n33346 = ~n33344 & ~n33345 ;
  assign n33347 = ~\P2_P3_InstAddrPointer_reg[14]/NET0131  & ~n33345 ;
  assign n33348 = \P2_P3_InstAddrPointer_reg[0]/NET0131  & n32919 ;
  assign n33349 = ~n33347 & ~n33348 ;
  assign n33350 = ~n33346 & ~n33349 ;
  assign n33351 = n33343 & n33350 ;
  assign n33352 = \P2_P3_InstAddrPointer_reg[15]/NET0131  & n33348 ;
  assign n33353 = ~\P2_P3_InstAddrPointer_reg[16]/NET0131  & ~n33352 ;
  assign n33354 = \P2_P3_InstAddrPointer_reg[0]/NET0131  & n32921 ;
  assign n33355 = ~n33353 & ~n33354 ;
  assign n33356 = ~\P2_P3_InstAddrPointer_reg[15]/NET0131  & ~n33348 ;
  assign n33357 = ~n33352 & ~n33356 ;
  assign n33358 = ~n33355 & ~n33357 ;
  assign n33359 = n33351 & n33358 ;
  assign n33360 = \P2_P3_InstAddrPointer_reg[17]/NET0131  & n32921 ;
  assign n33361 = \P2_P3_InstAddrPointer_reg[18]/NET0131  & n33360 ;
  assign n33362 = \P2_P3_InstAddrPointer_reg[0]/NET0131  & n33361 ;
  assign n33363 = ~\P2_P3_InstAddrPointer_reg[19]/NET0131  & ~n33362 ;
  assign n33364 = n32889 & n33354 ;
  assign n33365 = ~n33363 & ~n33364 ;
  assign n33366 = ~\P2_P3_InstAddrPointer_reg[20]/NET0131  & ~n33364 ;
  assign n33367 = ~n33275 & ~n33366 ;
  assign n33378 = ~n33365 & ~n33367 ;
  assign n33368 = ~\P2_P3_InstAddrPointer_reg[21]/NET0131  & ~n33275 ;
  assign n33369 = \P2_P3_InstAddrPointer_reg[21]/NET0131  & n32923 ;
  assign n33370 = \P2_P3_InstAddrPointer_reg[0]/NET0131  & n33369 ;
  assign n33371 = ~n33368 & ~n33370 ;
  assign n33372 = \P2_P3_InstAddrPointer_reg[0]/NET0131  & n33360 ;
  assign n33373 = ~\P2_P3_InstAddrPointer_reg[18]/NET0131  & ~n33372 ;
  assign n33374 = ~n33362 & ~n33373 ;
  assign n33375 = ~\P2_P3_InstAddrPointer_reg[17]/NET0131  & ~n33354 ;
  assign n33376 = ~n33372 & ~n33375 ;
  assign n33377 = ~n33374 & ~n33376 ;
  assign n33379 = ~n33371 & n33377 ;
  assign n33380 = n33378 & n33379 ;
  assign n33381 = n33359 & n33380 ;
  assign n33382 = ~\P2_P3_InstAddrPointer_reg[22]/NET0131  & ~n33370 ;
  assign n33383 = ~n33276 & ~n33382 ;
  assign n33384 = n33381 & ~n33383 ;
  assign n33385 = ~n33279 & n33384 ;
  assign n33386 = ~\P2_P3_InstAddrPointer_reg[24]/NET0131  & ~n33278 ;
  assign n33387 = \P2_P3_InstAddrPointer_reg[0]/NET0131  & n32924 ;
  assign n33388 = ~n33386 & ~n33387 ;
  assign n33389 = n33385 & ~n33388 ;
  assign n33390 = ~\P2_P3_InstAddrPointer_reg[25]/NET0131  & ~n33387 ;
  assign n33391 = \P2_P3_InstAddrPointer_reg[0]/NET0131  & n32925 ;
  assign n33392 = ~n33390 & ~n33391 ;
  assign n33393 = n33389 & ~n33392 ;
  assign n33394 = ~\P2_P3_InstAddrPointer_reg[26]/NET0131  & ~n33391 ;
  assign n33395 = \P2_P3_InstAddrPointer_reg[26]/NET0131  & n33391 ;
  assign n33396 = ~n33394 & ~n33395 ;
  assign n33397 = n33393 & ~n33396 ;
  assign n33398 = ~\P2_P3_InstAddrPointer_reg[27]/NET0131  & ~n33395 ;
  assign n33399 = n32906 & n33391 ;
  assign n33400 = ~n33398 & ~n33399 ;
  assign n33401 = n33397 & ~n33400 ;
  assign n33402 = ~\P2_P3_InstAddrPointer_reg[28]/NET0131  & ~n33399 ;
  assign n33403 = \P2_P3_InstAddrPointer_reg[28]/NET0131  & n33399 ;
  assign n33404 = ~n33402 & ~n33403 ;
  assign n33405 = n33401 & ~n33404 ;
  assign n33406 = ~\P2_P3_InstAddrPointer_reg[29]/NET0131  & ~n33403 ;
  assign n33407 = ~n32929 & ~n33406 ;
  assign n33408 = n33405 & ~n33407 ;
  assign n33409 = ~\P2_P3_InstAddrPointer_reg[30]/NET0131  & ~n32929 ;
  assign n33410 = ~n32930 & ~n33409 ;
  assign n33411 = n33408 & ~n33410 ;
  assign n33413 = n32933 & ~n33411 ;
  assign n33412 = ~n32933 & n33411 ;
  assign n33414 = ~n33242 & ~n33412 ;
  assign n33415 = ~n33413 & n33414 ;
  assign n33416 = ~n33274 & ~n33415 ;
  assign n33417 = n27284 & ~n33416 ;
  assign n32905 = n27219 & n32904 ;
  assign n32934 = ~n27142 & ~n32933 ;
  assign n32939 = ~n27229 & n32938 ;
  assign n32940 = ~n27257 & ~n32935 ;
  assign n32941 = n27192 & ~n27257 ;
  assign n32942 = ~n27126 & n27177 ;
  assign n32943 = ~n27275 & ~n32942 ;
  assign n32944 = n27296 & n32943 ;
  assign n32945 = ~n32941 & n32944 ;
  assign n32946 = ~n32940 & n32945 ;
  assign n32947 = \P2_P3_InstAddrPointer_reg[31]/NET0131  & ~n32946 ;
  assign n33506 = ~n32939 & ~n32947 ;
  assign n33507 = ~n32934 & n33506 ;
  assign n33508 = ~n32905 & n33507 ;
  assign n33509 = ~n33417 & n33508 ;
  assign n33510 = ~n33505 & n33509 ;
  assign n33511 = n27308 & ~n33510 ;
  assign n32864 = n27317 & n27649 ;
  assign n32865 = \P2_P3_rEIP_reg[31]/NET0131  & n32864 ;
  assign n32866 = ~n27317 & n27649 ;
  assign n32867 = n27307 & n27317 ;
  assign n32868 = ~n27314 & ~n27656 ;
  assign n32869 = ~n32867 & n32868 ;
  assign n32870 = ~n32866 & n32869 ;
  assign n32871 = \P2_P3_InstAddrPointer_reg[31]/NET0131  & ~n32870 ;
  assign n33512 = ~n32865 & ~n32871 ;
  assign n33513 = ~n33511 & n33512 ;
  assign n33514 = \P1_P1_InstAddrPointer_reg[31]/NET0131  & n26249 ;
  assign n33833 = \P1_P1_InstAddrPointer_reg[15]/NET0131  & \P1_P1_InstAddrPointer_reg[16]/NET0131  ;
  assign n33520 = \P1_P1_InstAddrPointer_reg[11]/NET0131  & \P1_P1_InstAddrPointer_reg[12]/NET0131  ;
  assign n33521 = \P1_P1_InstAddrPointer_reg[10]/NET0131  & n33520 ;
  assign n33522 = \P1_P1_InstAddrPointer_reg[1]/NET0131  & \P1_P1_InstAddrPointer_reg[2]/NET0131  ;
  assign n33523 = \P1_P1_InstAddrPointer_reg[3]/NET0131  & n33522 ;
  assign n33524 = \P1_P1_InstAddrPointer_reg[4]/NET0131  & n33523 ;
  assign n33525 = \P1_P1_InstAddrPointer_reg[5]/NET0131  & n33524 ;
  assign n33526 = \P1_P1_InstAddrPointer_reg[6]/NET0131  & n33525 ;
  assign n33527 = \P1_P1_InstAddrPointer_reg[7]/NET0131  & n33526 ;
  assign n33528 = \P1_P1_InstAddrPointer_reg[8]/NET0131  & n33527 ;
  assign n33529 = \P1_P1_InstAddrPointer_reg[9]/NET0131  & n33528 ;
  assign n33530 = n33521 & n33529 ;
  assign n33877 = \P1_P1_InstAddrPointer_reg[0]/NET0131  & n33530 ;
  assign n33878 = \P1_P1_InstAddrPointer_reg[13]/NET0131  & n33877 ;
  assign n33879 = \P1_P1_InstAddrPointer_reg[14]/NET0131  & n33878 ;
  assign n33880 = n33833 & n33879 ;
  assign n33881 = ~\P1_P1_InstAddrPointer_reg[17]/NET0131  & ~n33880 ;
  assign n33519 = \P1_P1_InstAddrPointer_reg[13]/NET0131  & \P1_P1_InstAddrPointer_reg[14]/NET0131  ;
  assign n33531 = n33519 & n33530 ;
  assign n33532 = \P1_P1_InstAddrPointer_reg[15]/NET0131  & n33531 ;
  assign n33533 = \P1_P1_InstAddrPointer_reg[16]/NET0131  & n33532 ;
  assign n33823 = \P1_P1_InstAddrPointer_reg[17]/NET0131  & n33533 ;
  assign n33882 = \P1_P1_InstAddrPointer_reg[0]/NET0131  & n33823 ;
  assign n33883 = ~n33881 & ~n33882 ;
  assign n33884 = \P1_P1_InstAddrPointer_reg[15]/NET0131  & n33879 ;
  assign n33885 = ~\P1_P1_InstAddrPointer_reg[15]/NET0131  & ~n33879 ;
  assign n33886 = ~n33884 & ~n33885 ;
  assign n33832 = \P1_P1_InstAddrPointer_reg[8]/NET0131  & \P1_P1_InstAddrPointer_reg[9]/NET0131  ;
  assign n33887 = \P1_P1_InstAddrPointer_reg[0]/NET0131  & \P1_P1_InstAddrPointer_reg[1]/NET0131  ;
  assign n33888 = \P1_P1_InstAddrPointer_reg[2]/NET0131  & n33887 ;
  assign n33889 = \P1_P1_InstAddrPointer_reg[3]/NET0131  & n33888 ;
  assign n33890 = \P1_P1_InstAddrPointer_reg[4]/NET0131  & n33889 ;
  assign n33891 = \P1_P1_InstAddrPointer_reg[5]/NET0131  & n33890 ;
  assign n33892 = \P1_P1_InstAddrPointer_reg[6]/NET0131  & n33891 ;
  assign n33893 = \P1_P1_InstAddrPointer_reg[7]/NET0131  & n33892 ;
  assign n33894 = n33832 & n33893 ;
  assign n33895 = ~\P1_P1_InstAddrPointer_reg[10]/NET0131  & ~n33894 ;
  assign n33896 = \P1_P1_InstAddrPointer_reg[10]/NET0131  & n33529 ;
  assign n33897 = \P1_P1_InstAddrPointer_reg[0]/NET0131  & n33896 ;
  assign n33898 = ~n33895 & ~n33897 ;
  assign n33899 = \P1_P1_InstAddrPointer_reg[8]/NET0131  & n33893 ;
  assign n33900 = ~\P1_P1_InstAddrPointer_reg[9]/NET0131  & ~n33899 ;
  assign n33901 = ~n33894 & ~n33900 ;
  assign n33902 = ~\P1_P1_InstAddrPointer_reg[8]/NET0131  & ~n33893 ;
  assign n33903 = ~n33899 & ~n33902 ;
  assign n33904 = ~\P1_P1_InstAddrPointer_reg[7]/NET0131  & ~n33892 ;
  assign n33905 = ~n33893 & ~n33904 ;
  assign n33906 = n29558 & ~n33905 ;
  assign n33907 = ~n29558 & n33905 ;
  assign n33561 = \P1_P1_InstQueue_reg[15][6]/NET0131  & n8291 ;
  assign n33562 = \P1_P1_InstQueue_reg[6][6]/NET0131  & n8307 ;
  assign n33563 = \P1_P1_InstQueue_reg[5][6]/NET0131  & n8295 ;
  assign n33577 = ~n33562 & ~n33563 ;
  assign n33564 = \P1_P1_InstQueue_reg[4][6]/NET0131  & n8323 ;
  assign n33565 = \P1_P1_InstQueue_reg[9][6]/NET0131  & n8305 ;
  assign n33578 = ~n33564 & ~n33565 ;
  assign n33587 = n33577 & n33578 ;
  assign n33588 = ~n33561 & n33587 ;
  assign n33576 = \P1_P1_InstQueue_reg[3][6]/NET0131  & n8314 ;
  assign n33574 = \P1_P1_InstQueue_reg[1][6]/NET0131  & n8309 ;
  assign n33575 = \P1_P1_InstQueue_reg[10][6]/NET0131  & n8325 ;
  assign n33583 = ~n33574 & ~n33575 ;
  assign n33584 = ~n33576 & n33583 ;
  assign n33570 = \P1_P1_InstQueue_reg[7][6]/NET0131  & n8316 ;
  assign n33571 = \P1_P1_InstQueue_reg[8][6]/NET0131  & n8318 ;
  assign n33581 = ~n33570 & ~n33571 ;
  assign n33572 = \P1_P1_InstQueue_reg[0][6]/NET0131  & n8321 ;
  assign n33573 = \P1_P1_InstQueue_reg[12][6]/NET0131  & n8312 ;
  assign n33582 = ~n33572 & ~n33573 ;
  assign n33585 = n33581 & n33582 ;
  assign n33566 = \P1_P1_InstQueue_reg[2][6]/NET0131  & n8299 ;
  assign n33567 = \P1_P1_InstQueue_reg[13][6]/NET0131  & n8329 ;
  assign n33579 = ~n33566 & ~n33567 ;
  assign n33568 = \P1_P1_InstQueue_reg[14][6]/NET0131  & n8327 ;
  assign n33569 = \P1_P1_InstQueue_reg[11][6]/NET0131  & n8303 ;
  assign n33580 = ~n33568 & ~n33569 ;
  assign n33586 = n33579 & n33580 ;
  assign n33589 = n33585 & n33586 ;
  assign n33590 = n33584 & n33589 ;
  assign n33591 = n33588 & n33590 ;
  assign n33908 = ~\P1_P1_InstAddrPointer_reg[6]/NET0131  & ~n33891 ;
  assign n33909 = ~n33892 & ~n33908 ;
  assign n33910 = n33591 & ~n33909 ;
  assign n33911 = ~n33591 & n33909 ;
  assign n33596 = \P1_P1_InstQueue_reg[15][5]/NET0131  & n8291 ;
  assign n33597 = \P1_P1_InstQueue_reg[10][5]/NET0131  & n8325 ;
  assign n33598 = \P1_P1_InstQueue_reg[5][5]/NET0131  & n8295 ;
  assign n33612 = ~n33597 & ~n33598 ;
  assign n33599 = \P1_P1_InstQueue_reg[6][5]/NET0131  & n8307 ;
  assign n33600 = \P1_P1_InstQueue_reg[4][5]/NET0131  & n8323 ;
  assign n33613 = ~n33599 & ~n33600 ;
  assign n33622 = n33612 & n33613 ;
  assign n33623 = ~n33596 & n33622 ;
  assign n33611 = \P1_P1_InstQueue_reg[1][5]/NET0131  & n8309 ;
  assign n33609 = \P1_P1_InstQueue_reg[11][5]/NET0131  & n8303 ;
  assign n33610 = \P1_P1_InstQueue_reg[13][5]/NET0131  & n8329 ;
  assign n33618 = ~n33609 & ~n33610 ;
  assign n33619 = ~n33611 & n33618 ;
  assign n33605 = \P1_P1_InstQueue_reg[7][5]/NET0131  & n8316 ;
  assign n33606 = \P1_P1_InstQueue_reg[0][5]/NET0131  & n8321 ;
  assign n33616 = ~n33605 & ~n33606 ;
  assign n33607 = \P1_P1_InstQueue_reg[8][5]/NET0131  & n8318 ;
  assign n33608 = \P1_P1_InstQueue_reg[12][5]/NET0131  & n8312 ;
  assign n33617 = ~n33607 & ~n33608 ;
  assign n33620 = n33616 & n33617 ;
  assign n33601 = \P1_P1_InstQueue_reg[3][5]/NET0131  & n8314 ;
  assign n33602 = \P1_P1_InstQueue_reg[9][5]/NET0131  & n8305 ;
  assign n33614 = ~n33601 & ~n33602 ;
  assign n33603 = \P1_P1_InstQueue_reg[2][5]/NET0131  & n8299 ;
  assign n33604 = \P1_P1_InstQueue_reg[14][5]/NET0131  & n8327 ;
  assign n33615 = ~n33603 & ~n33604 ;
  assign n33621 = n33614 & n33615 ;
  assign n33624 = n33620 & n33621 ;
  assign n33625 = n33619 & n33624 ;
  assign n33626 = n33623 & n33625 ;
  assign n33912 = ~\P1_P1_InstAddrPointer_reg[5]/NET0131  & ~n33890 ;
  assign n33913 = ~n33891 & ~n33912 ;
  assign n33914 = n33626 & ~n33913 ;
  assign n33915 = ~n33626 & n33913 ;
  assign n33631 = \P1_P1_InstQueue_reg[15][4]/NET0131  & n8291 ;
  assign n33632 = \P1_P1_InstQueue_reg[9][4]/NET0131  & n8305 ;
  assign n33633 = \P1_P1_InstQueue_reg[14][4]/NET0131  & n8327 ;
  assign n33647 = ~n33632 & ~n33633 ;
  assign n33634 = \P1_P1_InstQueue_reg[10][4]/NET0131  & n8325 ;
  assign n33635 = \P1_P1_InstQueue_reg[12][4]/NET0131  & n8312 ;
  assign n33648 = ~n33634 & ~n33635 ;
  assign n33657 = n33647 & n33648 ;
  assign n33658 = ~n33631 & n33657 ;
  assign n33646 = \P1_P1_InstQueue_reg[1][4]/NET0131  & n8309 ;
  assign n33644 = \P1_P1_InstQueue_reg[5][4]/NET0131  & n8295 ;
  assign n33645 = \P1_P1_InstQueue_reg[6][4]/NET0131  & n8307 ;
  assign n33653 = ~n33644 & ~n33645 ;
  assign n33654 = ~n33646 & n33653 ;
  assign n33640 = \P1_P1_InstQueue_reg[7][4]/NET0131  & n8316 ;
  assign n33641 = \P1_P1_InstQueue_reg[0][4]/NET0131  & n8321 ;
  assign n33651 = ~n33640 & ~n33641 ;
  assign n33642 = \P1_P1_InstQueue_reg[8][4]/NET0131  & n8318 ;
  assign n33643 = \P1_P1_InstQueue_reg[4][4]/NET0131  & n8323 ;
  assign n33652 = ~n33642 & ~n33643 ;
  assign n33655 = n33651 & n33652 ;
  assign n33636 = \P1_P1_InstQueue_reg[11][4]/NET0131  & n8303 ;
  assign n33637 = \P1_P1_InstQueue_reg[13][4]/NET0131  & n8329 ;
  assign n33649 = ~n33636 & ~n33637 ;
  assign n33638 = \P1_P1_InstQueue_reg[2][4]/NET0131  & n8299 ;
  assign n33639 = \P1_P1_InstQueue_reg[3][4]/NET0131  & n8314 ;
  assign n33650 = ~n33638 & ~n33639 ;
  assign n33656 = n33649 & n33650 ;
  assign n33659 = n33655 & n33656 ;
  assign n33660 = n33654 & n33659 ;
  assign n33661 = n33658 & n33660 ;
  assign n33916 = ~\P1_P1_InstAddrPointer_reg[4]/NET0131  & ~n33889 ;
  assign n33917 = ~n33890 & ~n33916 ;
  assign n33918 = n33661 & ~n33917 ;
  assign n33919 = ~n33661 & n33917 ;
  assign n33666 = \P1_P1_InstQueue_reg[15][3]/NET0131  & n8291 ;
  assign n33667 = \P1_P1_InstQueue_reg[3][3]/NET0131  & n8314 ;
  assign n33668 = \P1_P1_InstQueue_reg[14][3]/NET0131  & n8327 ;
  assign n33682 = ~n33667 & ~n33668 ;
  assign n33669 = \P1_P1_InstQueue_reg[12][3]/NET0131  & n8312 ;
  assign n33670 = \P1_P1_InstQueue_reg[4][3]/NET0131  & n8323 ;
  assign n33683 = ~n33669 & ~n33670 ;
  assign n33692 = n33682 & n33683 ;
  assign n33693 = ~n33666 & n33692 ;
  assign n33681 = \P1_P1_InstQueue_reg[5][3]/NET0131  & n8295 ;
  assign n33679 = \P1_P1_InstQueue_reg[6][3]/NET0131  & n8307 ;
  assign n33680 = \P1_P1_InstQueue_reg[11][3]/NET0131  & n8303 ;
  assign n33688 = ~n33679 & ~n33680 ;
  assign n33689 = ~n33681 & n33688 ;
  assign n33675 = \P1_P1_InstQueue_reg[7][3]/NET0131  & n8316 ;
  assign n33676 = \P1_P1_InstQueue_reg[0][3]/NET0131  & n8321 ;
  assign n33686 = ~n33675 & ~n33676 ;
  assign n33677 = \P1_P1_InstQueue_reg[8][3]/NET0131  & n8318 ;
  assign n33678 = \P1_P1_InstQueue_reg[13][3]/NET0131  & n8329 ;
  assign n33687 = ~n33677 & ~n33678 ;
  assign n33690 = n33686 & n33687 ;
  assign n33671 = \P1_P1_InstQueue_reg[1][3]/NET0131  & n8309 ;
  assign n33672 = \P1_P1_InstQueue_reg[9][3]/NET0131  & n8305 ;
  assign n33684 = ~n33671 & ~n33672 ;
  assign n33673 = \P1_P1_InstQueue_reg[2][3]/NET0131  & n8299 ;
  assign n33674 = \P1_P1_InstQueue_reg[10][3]/NET0131  & n8325 ;
  assign n33685 = ~n33673 & ~n33674 ;
  assign n33691 = n33684 & n33685 ;
  assign n33694 = n33690 & n33691 ;
  assign n33695 = n33689 & n33694 ;
  assign n33696 = n33693 & n33695 ;
  assign n33920 = ~\P1_P1_InstAddrPointer_reg[3]/NET0131  & ~n33888 ;
  assign n33921 = ~n33889 & ~n33920 ;
  assign n33922 = n33696 & ~n33921 ;
  assign n33923 = ~n33696 & n33921 ;
  assign n33716 = \P1_P1_InstQueue_reg[15][2]/NET0131  & n8291 ;
  assign n33701 = \P1_P1_InstQueue_reg[9][2]/NET0131  & n8305 ;
  assign n33702 = \P1_P1_InstQueue_reg[6][2]/NET0131  & n8307 ;
  assign n33717 = ~n33701 & ~n33702 ;
  assign n33703 = \P1_P1_InstQueue_reg[8][2]/NET0131  & n8318 ;
  assign n33704 = \P1_P1_InstQueue_reg[13][2]/NET0131  & n8329 ;
  assign n33718 = ~n33703 & ~n33704 ;
  assign n33727 = n33717 & n33718 ;
  assign n33728 = ~n33716 & n33727 ;
  assign n33715 = \P1_P1_InstQueue_reg[1][2]/NET0131  & n8309 ;
  assign n33713 = \P1_P1_InstQueue_reg[0][2]/NET0131  & n8321 ;
  assign n33714 = \P1_P1_InstQueue_reg[5][2]/NET0131  & n8295 ;
  assign n33723 = ~n33713 & ~n33714 ;
  assign n33724 = ~n33715 & n33723 ;
  assign n33709 = \P1_P1_InstQueue_reg[14][2]/NET0131  & n8327 ;
  assign n33710 = \P1_P1_InstQueue_reg[11][2]/NET0131  & n8303 ;
  assign n33721 = ~n33709 & ~n33710 ;
  assign n33711 = \P1_P1_InstQueue_reg[2][2]/NET0131  & n8299 ;
  assign n33712 = \P1_P1_InstQueue_reg[3][2]/NET0131  & n8314 ;
  assign n33722 = ~n33711 & ~n33712 ;
  assign n33725 = n33721 & n33722 ;
  assign n33705 = \P1_P1_InstQueue_reg[4][2]/NET0131  & n8323 ;
  assign n33706 = \P1_P1_InstQueue_reg[7][2]/NET0131  & n8316 ;
  assign n33719 = ~n33705 & ~n33706 ;
  assign n33707 = \P1_P1_InstQueue_reg[10][2]/NET0131  & n8325 ;
  assign n33708 = \P1_P1_InstQueue_reg[12][2]/NET0131  & n8312 ;
  assign n33720 = ~n33707 & ~n33708 ;
  assign n33726 = n33719 & n33720 ;
  assign n33729 = n33725 & n33726 ;
  assign n33730 = n33724 & n33729 ;
  assign n33731 = n33728 & n33730 ;
  assign n33924 = ~\P1_P1_InstAddrPointer_reg[2]/NET0131  & ~n33887 ;
  assign n33925 = ~n33888 & ~n33924 ;
  assign n33926 = ~n33731 & n33925 ;
  assign n33927 = n33731 & ~n33925 ;
  assign n33744 = \P1_P1_InstQueue_reg[15][1]/NET0131  & n8291 ;
  assign n33734 = \P1_P1_InstQueue_reg[7][1]/NET0131  & n8316 ;
  assign n33735 = \P1_P1_InstQueue_reg[8][1]/NET0131  & n8318 ;
  assign n33750 = ~n33734 & ~n33735 ;
  assign n33736 = \P1_P1_InstQueue_reg[6][1]/NET0131  & n8307 ;
  assign n33737 = \P1_P1_InstQueue_reg[4][1]/NET0131  & n8323 ;
  assign n33751 = ~n33736 & ~n33737 ;
  assign n33760 = n33750 & n33751 ;
  assign n33761 = ~n33744 & n33760 ;
  assign n33749 = \P1_P1_InstQueue_reg[1][1]/NET0131  & n8309 ;
  assign n33747 = \P1_P1_InstQueue_reg[3][1]/NET0131  & n8314 ;
  assign n33748 = \P1_P1_InstQueue_reg[10][1]/NET0131  & n8325 ;
  assign n33756 = ~n33747 & ~n33748 ;
  assign n33757 = ~n33749 & n33756 ;
  assign n33742 = \P1_P1_InstQueue_reg[12][1]/NET0131  & n8312 ;
  assign n33743 = \P1_P1_InstQueue_reg[13][1]/NET0131  & n8329 ;
  assign n33754 = ~n33742 & ~n33743 ;
  assign n33745 = \P1_P1_InstQueue_reg[14][1]/NET0131  & n8327 ;
  assign n33746 = \P1_P1_InstQueue_reg[11][1]/NET0131  & n8303 ;
  assign n33755 = ~n33745 & ~n33746 ;
  assign n33758 = n33754 & n33755 ;
  assign n33738 = \P1_P1_InstQueue_reg[0][1]/NET0131  & n8321 ;
  assign n33739 = \P1_P1_InstQueue_reg[5][1]/NET0131  & n8295 ;
  assign n33752 = ~n33738 & ~n33739 ;
  assign n33740 = \P1_P1_InstQueue_reg[9][1]/NET0131  & n8305 ;
  assign n33741 = \P1_P1_InstQueue_reg[2][1]/NET0131  & n8299 ;
  assign n33753 = ~n33740 & ~n33741 ;
  assign n33759 = n33752 & n33753 ;
  assign n33762 = n33758 & n33759 ;
  assign n33763 = n33757 & n33762 ;
  assign n33764 = n33761 & n33763 ;
  assign n33765 = ~\P1_P1_InstAddrPointer_reg[1]/NET0131  & ~n33764 ;
  assign n33766 = \P1_P1_InstAddrPointer_reg[1]/NET0131  & n33764 ;
  assign n33777 = \P1_P1_InstQueue_reg[15][0]/NET0131  & n8291 ;
  assign n33767 = \P1_P1_InstQueue_reg[7][0]/NET0131  & n8316 ;
  assign n33768 = \P1_P1_InstQueue_reg[0][0]/NET0131  & n8321 ;
  assign n33783 = ~n33767 & ~n33768 ;
  assign n33769 = \P1_P1_InstQueue_reg[6][0]/NET0131  & n8307 ;
  assign n33770 = \P1_P1_InstQueue_reg[5][0]/NET0131  & n8295 ;
  assign n33784 = ~n33769 & ~n33770 ;
  assign n33793 = n33783 & n33784 ;
  assign n33794 = ~n33777 & n33793 ;
  assign n33782 = \P1_P1_InstQueue_reg[13][0]/NET0131  & n8329 ;
  assign n33780 = \P1_P1_InstQueue_reg[3][0]/NET0131  & n8314 ;
  assign n33781 = \P1_P1_InstQueue_reg[1][0]/NET0131  & n8309 ;
  assign n33789 = ~n33780 & ~n33781 ;
  assign n33790 = ~n33782 & n33789 ;
  assign n33775 = \P1_P1_InstQueue_reg[4][0]/NET0131  & n8323 ;
  assign n33776 = \P1_P1_InstQueue_reg[14][0]/NET0131  & n8327 ;
  assign n33787 = ~n33775 & ~n33776 ;
  assign n33778 = \P1_P1_InstQueue_reg[2][0]/NET0131  & n8299 ;
  assign n33779 = \P1_P1_InstQueue_reg[11][0]/NET0131  & n8303 ;
  assign n33788 = ~n33778 & ~n33779 ;
  assign n33791 = n33787 & n33788 ;
  assign n33771 = \P1_P1_InstQueue_reg[8][0]/NET0131  & n8318 ;
  assign n33772 = \P1_P1_InstQueue_reg[10][0]/NET0131  & n8325 ;
  assign n33785 = ~n33771 & ~n33772 ;
  assign n33773 = \P1_P1_InstQueue_reg[12][0]/NET0131  & n8312 ;
  assign n33774 = \P1_P1_InstQueue_reg[9][0]/NET0131  & n8305 ;
  assign n33786 = ~n33773 & ~n33774 ;
  assign n33792 = n33785 & n33786 ;
  assign n33795 = n33791 & n33792 ;
  assign n33796 = n33790 & n33795 ;
  assign n33797 = n33794 & n33796 ;
  assign n33798 = \P1_P1_InstAddrPointer_reg[0]/NET0131  & ~n33797 ;
  assign n33799 = ~n33766 & n33798 ;
  assign n33800 = ~n33765 & ~n33799 ;
  assign n33928 = ~\P1_P1_InstAddrPointer_reg[0]/NET0131  & \P1_P1_InstAddrPointer_reg[1]/NET0131  ;
  assign n33929 = n33800 & ~n33928 ;
  assign n33930 = ~n33927 & ~n33929 ;
  assign n33931 = ~n33926 & ~n33930 ;
  assign n33932 = ~n33923 & n33931 ;
  assign n33933 = ~n33922 & ~n33932 ;
  assign n33934 = ~n33919 & ~n33933 ;
  assign n33935 = ~n33918 & ~n33934 ;
  assign n33936 = ~n33915 & ~n33935 ;
  assign n33937 = ~n33914 & ~n33936 ;
  assign n33938 = ~n33911 & ~n33937 ;
  assign n33939 = ~n33910 & ~n33938 ;
  assign n33940 = ~n33907 & ~n33939 ;
  assign n33941 = ~n33906 & ~n33940 ;
  assign n33942 = ~n33903 & ~n33941 ;
  assign n33943 = ~n33901 & n33942 ;
  assign n33944 = ~n33898 & n33943 ;
  assign n33945 = ~\P1_P1_InstAddrPointer_reg[11]/NET0131  & ~n33897 ;
  assign n33946 = \P1_P1_InstAddrPointer_reg[11]/NET0131  & n33896 ;
  assign n33947 = \P1_P1_InstAddrPointer_reg[0]/NET0131  & n33946 ;
  assign n33948 = ~n33945 & ~n33947 ;
  assign n33949 = n33944 & ~n33948 ;
  assign n33950 = ~\P1_P1_InstAddrPointer_reg[12]/NET0131  & ~n33947 ;
  assign n33951 = ~n33877 & ~n33950 ;
  assign n33952 = n33949 & ~n33951 ;
  assign n33953 = ~\P1_P1_InstAddrPointer_reg[13]/NET0131  & ~n33877 ;
  assign n33954 = ~n33878 & ~n33953 ;
  assign n33955 = ~\P1_P1_InstAddrPointer_reg[14]/NET0131  & ~n33878 ;
  assign n33956 = ~n33879 & ~n33955 ;
  assign n33957 = ~n33954 & ~n33956 ;
  assign n33958 = n33952 & n33957 ;
  assign n33959 = ~n33886 & n33958 ;
  assign n33960 = ~\P1_P1_InstAddrPointer_reg[16]/NET0131  & ~n33884 ;
  assign n33961 = ~n33880 & ~n33960 ;
  assign n33962 = n33959 & ~n33961 ;
  assign n33963 = ~n33883 & n33962 ;
  assign n33517 = \P1_P1_InstAddrPointer_reg[18]/NET0131  & \P1_P1_InstAddrPointer_reg[19]/NET0131  ;
  assign n33518 = \P1_P1_InstAddrPointer_reg[17]/NET0131  & n33517 ;
  assign n33534 = n33518 & n33533 ;
  assign n33535 = \P1_P1_InstAddrPointer_reg[20]/NET0131  & n33534 ;
  assign n33846 = \P1_P1_InstAddrPointer_reg[21]/NET0131  & n33535 ;
  assign n33870 = \P1_P1_InstAddrPointer_reg[0]/NET0131  & n33846 ;
  assign n33964 = n33518 & n33880 ;
  assign n33965 = \P1_P1_InstAddrPointer_reg[20]/NET0131  & n33964 ;
  assign n33966 = ~\P1_P1_InstAddrPointer_reg[21]/NET0131  & ~n33965 ;
  assign n33967 = ~n33870 & ~n33966 ;
  assign n33968 = \P1_P1_InstAddrPointer_reg[18]/NET0131  & n33823 ;
  assign n33969 = \P1_P1_InstAddrPointer_reg[0]/NET0131  & n33968 ;
  assign n33970 = ~\P1_P1_InstAddrPointer_reg[19]/NET0131  & ~n33969 ;
  assign n33971 = ~n33964 & ~n33970 ;
  assign n33972 = ~\P1_P1_InstAddrPointer_reg[18]/NET0131  & ~n33882 ;
  assign n33973 = ~n33969 & ~n33972 ;
  assign n33974 = ~\P1_P1_InstAddrPointer_reg[20]/NET0131  & ~n33964 ;
  assign n33975 = ~n33965 & ~n33974 ;
  assign n33976 = ~n33973 & ~n33975 ;
  assign n33977 = ~n33971 & n33976 ;
  assign n33978 = ~n33967 & n33977 ;
  assign n33979 = n33963 & n33978 ;
  assign n33871 = ~\P1_P1_InstAddrPointer_reg[22]/NET0131  & ~n33870 ;
  assign n33872 = \P1_P1_InstAddrPointer_reg[22]/NET0131  & n33870 ;
  assign n33873 = ~n33871 & ~n33872 ;
  assign n33874 = \P1_P1_InstAddrPointer_reg[23]/NET0131  & ~n33872 ;
  assign n33875 = ~\P1_P1_InstAddrPointer_reg[23]/NET0131  & n33872 ;
  assign n33876 = ~n33874 & ~n33875 ;
  assign n33980 = ~n33873 & n33876 ;
  assign n33981 = n33979 & n33980 ;
  assign n33515 = \P1_P1_InstAddrPointer_reg[23]/NET0131  & \P1_P1_InstAddrPointer_reg[24]/NET0131  ;
  assign n33982 = n33515 & n33872 ;
  assign n33983 = ~\P1_P1_InstAddrPointer_reg[25]/NET0131  & ~n33982 ;
  assign n33984 = \P1_P1_InstAddrPointer_reg[25]/NET0131  & n33982 ;
  assign n33985 = ~n33983 & ~n33984 ;
  assign n33986 = \P1_P1_InstAddrPointer_reg[24]/NET0131  & ~n33893 ;
  assign n33835 = \P1_P1_InstAddrPointer_reg[23]/NET0131  & n33519 ;
  assign n33836 = n33832 & n33833 ;
  assign n33837 = n33835 & n33836 ;
  assign n33516 = \P1_P1_InstAddrPointer_reg[21]/NET0131  & \P1_P1_InstAddrPointer_reg[22]/NET0131  ;
  assign n33834 = \P1_P1_InstAddrPointer_reg[20]/NET0131  & n33516 ;
  assign n33838 = n33518 & n33521 ;
  assign n33839 = n33834 & n33838 ;
  assign n33840 = n33837 & n33839 ;
  assign n33841 = \P1_P1_InstAddrPointer_reg[24]/NET0131  & ~n33840 ;
  assign n33842 = ~\P1_P1_InstAddrPointer_reg[24]/NET0131  & n33840 ;
  assign n33843 = ~n33841 & ~n33842 ;
  assign n33987 = ~n33843 & n33893 ;
  assign n33988 = ~n33986 & ~n33987 ;
  assign n33989 = ~n33985 & n33988 ;
  assign n33990 = n33981 & n33989 ;
  assign n33991 = \P1_P1_InstAddrPointer_reg[26]/NET0131  & n33984 ;
  assign n33992 = ~\P1_P1_InstAddrPointer_reg[27]/NET0131  & ~n33991 ;
  assign n33539 = \P1_P1_InstAddrPointer_reg[26]/NET0131  & \P1_P1_InstAddrPointer_reg[27]/NET0131  ;
  assign n33993 = n33539 & n33984 ;
  assign n33994 = ~n33992 & ~n33993 ;
  assign n33995 = ~\P1_P1_InstAddrPointer_reg[26]/NET0131  & ~n33984 ;
  assign n33996 = ~n33991 & ~n33995 ;
  assign n33997 = ~n33994 & ~n33996 ;
  assign n33998 = n33990 & n33997 ;
  assign n33999 = ~\P1_P1_InstAddrPointer_reg[28]/NET0131  & ~n33993 ;
  assign n34000 = \P1_P1_InstAddrPointer_reg[28]/NET0131  & n33993 ;
  assign n34001 = ~n33999 & ~n34000 ;
  assign n34002 = n33998 & ~n34001 ;
  assign n34003 = ~\P1_P1_InstAddrPointer_reg[29]/NET0131  & ~n34000 ;
  assign n33536 = n33516 & n33535 ;
  assign n33537 = n33515 & n33536 ;
  assign n33538 = \P1_P1_InstAddrPointer_reg[25]/NET0131  & n33537 ;
  assign n33540 = n33538 & n33539 ;
  assign n33541 = \P1_P1_InstAddrPointer_reg[28]/NET0131  & n33540 ;
  assign n33542 = \P1_P1_InstAddrPointer_reg[29]/NET0131  & n33541 ;
  assign n34004 = \P1_P1_InstAddrPointer_reg[0]/NET0131  & n33542 ;
  assign n34005 = ~n34003 & ~n34004 ;
  assign n34006 = n34002 & ~n34005 ;
  assign n34007 = ~\P1_P1_InstAddrPointer_reg[30]/NET0131  & ~n34004 ;
  assign n33543 = \P1_P1_InstAddrPointer_reg[30]/NET0131  & n33542 ;
  assign n34008 = \P1_P1_InstAddrPointer_reg[0]/NET0131  & n33543 ;
  assign n34009 = ~n34007 & ~n34008 ;
  assign n34010 = n34006 & ~n34009 ;
  assign n34011 = ~\P1_P1_InstAddrPointer_reg[31]/NET0131  & ~n34008 ;
  assign n34012 = \P1_P1_InstAddrPointer_reg[31]/NET0131  & n34008 ;
  assign n34013 = ~n34011 & ~n34012 ;
  assign n34015 = ~n34010 & n34013 ;
  assign n34014 = n34010 & ~n34013 ;
  assign n34016 = ~n29558 & ~n34014 ;
  assign n34017 = ~n34015 & n34016 ;
  assign n33544 = ~\P1_P1_InstAddrPointer_reg[30]/NET0131  & ~n33542 ;
  assign n33545 = ~n33543 & ~n33544 ;
  assign n33546 = ~\P1_P1_InstAddrPointer_reg[28]/NET0131  & ~n33540 ;
  assign n33547 = ~n33541 & ~n33546 ;
  assign n33548 = ~\P1_P1_InstAddrPointer_reg[15]/NET0131  & ~n33531 ;
  assign n33549 = ~n33532 & ~n33548 ;
  assign n33550 = \P1_P1_InstAddrPointer_reg[13]/NET0131  & n33530 ;
  assign n33551 = ~\P1_P1_InstAddrPointer_reg[13]/NET0131  & ~n33530 ;
  assign n33552 = ~n33550 & ~n33551 ;
  assign n33555 = ~\P1_P1_InstAddrPointer_reg[8]/NET0131  & ~n33527 ;
  assign n33556 = ~n33528 & ~n33555 ;
  assign n33557 = ~\P1_P1_InstAddrPointer_reg[7]/NET0131  & ~n33526 ;
  assign n33558 = ~n33527 & ~n33557 ;
  assign n33559 = ~\P1_P1_InstAddrPointer_reg[6]/NET0131  & ~n33525 ;
  assign n33560 = ~n33526 & ~n33559 ;
  assign n33592 = n33560 & ~n33591 ;
  assign n33593 = ~n33560 & n33591 ;
  assign n33594 = ~\P1_P1_InstAddrPointer_reg[5]/NET0131  & ~n33524 ;
  assign n33595 = ~n33525 & ~n33594 ;
  assign n33627 = n33595 & ~n33626 ;
  assign n33628 = ~n33595 & n33626 ;
  assign n33629 = ~\P1_P1_InstAddrPointer_reg[4]/NET0131  & ~n33523 ;
  assign n33630 = ~n33524 & ~n33629 ;
  assign n33662 = n33630 & ~n33661 ;
  assign n33663 = ~n33630 & n33661 ;
  assign n33664 = ~\P1_P1_InstAddrPointer_reg[3]/NET0131  & ~n33522 ;
  assign n33665 = ~n33523 & ~n33664 ;
  assign n33697 = n33665 & ~n33696 ;
  assign n33698 = ~n33665 & n33696 ;
  assign n33699 = ~\P1_P1_InstAddrPointer_reg[1]/NET0131  & ~\P1_P1_InstAddrPointer_reg[2]/NET0131  ;
  assign n33700 = ~n33522 & ~n33699 ;
  assign n33732 = n33700 & ~n33731 ;
  assign n33733 = ~n33700 & n33731 ;
  assign n33801 = ~n33733 & ~n33800 ;
  assign n33802 = ~n33732 & ~n33801 ;
  assign n33803 = ~n33698 & ~n33802 ;
  assign n33804 = ~n33697 & ~n33803 ;
  assign n33805 = ~n33663 & ~n33804 ;
  assign n33806 = ~n33662 & ~n33805 ;
  assign n33807 = ~n33628 & ~n33806 ;
  assign n33808 = ~n33627 & ~n33807 ;
  assign n33809 = ~n33593 & ~n33808 ;
  assign n33810 = ~n33592 & ~n33809 ;
  assign n33811 = n33558 & ~n33810 ;
  assign n33812 = n29558 & ~n33811 ;
  assign n33813 = ~n33558 & n33810 ;
  assign n33814 = ~n33812 & ~n33813 ;
  assign n33815 = n33556 & n33814 ;
  assign n33553 = ~\P1_P1_InstAddrPointer_reg[9]/NET0131  & ~n33528 ;
  assign n33554 = ~n33529 & ~n33553 ;
  assign n33816 = \P1_P1_InstAddrPointer_reg[10]/NET0131  & n33554 ;
  assign n33817 = n33815 & n33816 ;
  assign n33818 = n33520 & n33817 ;
  assign n33819 = n33552 & n33818 ;
  assign n33820 = \P1_P1_InstAddrPointer_reg[14]/NET0131  & n33819 ;
  assign n33821 = n33549 & n33820 ;
  assign n33822 = \P1_P1_InstAddrPointer_reg[16]/NET0131  & n33821 ;
  assign n33824 = ~\P1_P1_InstAddrPointer_reg[17]/NET0131  & ~n33533 ;
  assign n33825 = ~n33823 & ~n33824 ;
  assign n33826 = n33517 & n33825 ;
  assign n33827 = n33822 & n33826 ;
  assign n33828 = ~\P1_P1_InstAddrPointer_reg[20]/NET0131  & ~n33534 ;
  assign n33829 = ~n33535 & ~n33828 ;
  assign n33830 = n33827 & n33829 ;
  assign n33831 = \P1_P1_InstAddrPointer_reg[24]/NET0131  & ~n33527 ;
  assign n33844 = n33527 & ~n33843 ;
  assign n33845 = ~n33831 & ~n33844 ;
  assign n33849 = \P1_P1_InstAddrPointer_reg[23]/NET0131  & n33536 ;
  assign n33850 = ~\P1_P1_InstAddrPointer_reg[23]/NET0131  & ~n33536 ;
  assign n33851 = ~n33849 & ~n33850 ;
  assign n33847 = ~\P1_P1_InstAddrPointer_reg[21]/NET0131  & ~n33535 ;
  assign n33848 = ~n33846 & ~n33847 ;
  assign n33852 = \P1_P1_InstAddrPointer_reg[22]/NET0131  & n33848 ;
  assign n33853 = n33851 & n33852 ;
  assign n33854 = ~n33845 & n33853 ;
  assign n33855 = n33830 & n33854 ;
  assign n33856 = ~\P1_P1_InstAddrPointer_reg[25]/NET0131  & ~n33537 ;
  assign n33857 = ~n33538 & ~n33856 ;
  assign n33858 = n33539 & n33857 ;
  assign n33859 = n33855 & n33858 ;
  assign n33860 = n33547 & n33859 ;
  assign n33861 = \P1_P1_InstAddrPointer_reg[29]/NET0131  & n33860 ;
  assign n33862 = n33545 & n33861 ;
  assign n33867 = ~\P1_P1_InstAddrPointer_reg[31]/NET0131  & n33862 ;
  assign n33863 = \P1_P1_InstAddrPointer_reg[31]/NET0131  & ~n33543 ;
  assign n33864 = ~\P1_P1_InstAddrPointer_reg[31]/NET0131  & n33543 ;
  assign n33865 = ~n33863 & ~n33864 ;
  assign n33866 = ~n33862 & ~n33865 ;
  assign n33868 = n29558 & ~n33866 ;
  assign n33869 = ~n33867 & n33868 ;
  assign n34018 = ~n26249 & ~n33869 ;
  assign n34019 = ~n34017 & n34018 ;
  assign n34020 = ~n33514 & ~n34019 ;
  assign n34021 = n26126 & ~n34020 ;
  assign n34022 = \P1_P1_InstAddrPointer_reg[3]/NET0131  & ~n33924 ;
  assign n34023 = \P1_P1_InstAddrPointer_reg[4]/NET0131  & n34022 ;
  assign n34024 = \P1_P1_InstAddrPointer_reg[5]/NET0131  & n34023 ;
  assign n34025 = \P1_P1_InstAddrPointer_reg[6]/NET0131  & n34024 ;
  assign n34026 = \P1_P1_InstAddrPointer_reg[7]/NET0131  & n34025 ;
  assign n34027 = \P1_P1_InstAddrPointer_reg[8]/NET0131  & n34026 ;
  assign n34028 = \P1_P1_InstAddrPointer_reg[9]/NET0131  & n34027 ;
  assign n34029 = \P1_P1_InstAddrPointer_reg[10]/NET0131  & n34028 ;
  assign n34030 = n33520 & n34029 ;
  assign n34031 = n33519 & n34030 ;
  assign n34032 = \P1_P1_InstAddrPointer_reg[15]/NET0131  & n34031 ;
  assign n34033 = \P1_P1_InstAddrPointer_reg[16]/NET0131  & n34032 ;
  assign n34034 = n33518 & n34033 ;
  assign n34035 = n33834 & n34034 ;
  assign n34036 = n33515 & n34035 ;
  assign n34037 = \P1_P1_InstAddrPointer_reg[25]/NET0131  & n34036 ;
  assign n34038 = \P1_P1_InstAddrPointer_reg[26]/NET0131  & n34037 ;
  assign n34039 = \P1_P1_InstAddrPointer_reg[27]/NET0131  & n34038 ;
  assign n34040 = \P1_P1_InstAddrPointer_reg[28]/NET0131  & n34039 ;
  assign n34041 = ~\P1_P1_InstAddrPointer_reg[28]/NET0131  & ~n34039 ;
  assign n34042 = ~n34040 & ~n34041 ;
  assign n34043 = ~\P1_P1_InstAddrPointer_reg[20]/NET0131  & ~n34034 ;
  assign n34044 = \P1_P1_InstAddrPointer_reg[20]/NET0131  & n34034 ;
  assign n34045 = ~n34043 & ~n34044 ;
  assign n34046 = ~\P1_P1_InstAddrPointer_reg[15]/NET0131  & ~n34031 ;
  assign n34047 = ~n34032 & ~n34046 ;
  assign n34048 = \P1_P1_InstAddrPointer_reg[13]/NET0131  & n34030 ;
  assign n34049 = ~\P1_P1_InstAddrPointer_reg[13]/NET0131  & ~n34030 ;
  assign n34050 = ~n34048 & ~n34049 ;
  assign n34051 = ~\P1_P1_InstAddrPointer_reg[10]/NET0131  & ~n34028 ;
  assign n34052 = ~n34029 & ~n34051 ;
  assign n34053 = ~\P1_P1_InstAddrPointer_reg[8]/NET0131  & ~n34026 ;
  assign n34054 = ~n34027 & ~n34053 ;
  assign n34055 = ~\P1_P1_InstAddrPointer_reg[7]/NET0131  & ~n34025 ;
  assign n34056 = ~n34026 & ~n34055 ;
  assign n34057 = ~n29558 & n34056 ;
  assign n34058 = n29558 & ~n34056 ;
  assign n34059 = ~\P1_P1_InstAddrPointer_reg[6]/NET0131  & ~n34024 ;
  assign n34060 = ~n34025 & ~n34059 ;
  assign n34061 = ~n33591 & n34060 ;
  assign n34062 = n33591 & ~n34060 ;
  assign n34063 = ~\P1_P1_InstAddrPointer_reg[5]/NET0131  & ~n34023 ;
  assign n34064 = ~n34024 & ~n34063 ;
  assign n34065 = ~n33626 & n34064 ;
  assign n34066 = n33626 & ~n34064 ;
  assign n34067 = ~\P1_P1_InstAddrPointer_reg[4]/NET0131  & ~n34022 ;
  assign n34068 = ~n34023 & ~n34067 ;
  assign n34069 = ~n33661 & n34068 ;
  assign n34070 = n33661 & ~n34068 ;
  assign n34071 = ~\P1_P1_InstAddrPointer_reg[3]/NET0131  & n33924 ;
  assign n34072 = ~n34022 & ~n34071 ;
  assign n34073 = ~n33696 & n34072 ;
  assign n34074 = n33696 & ~n34072 ;
  assign n34075 = ~n33731 & ~n33925 ;
  assign n34076 = n33731 & n33925 ;
  assign n34077 = \P1_P1_InstAddrPointer_reg[0]/NET0131  & ~\P1_P1_InstAddrPointer_reg[1]/NET0131  ;
  assign n34078 = ~n33928 & ~n34077 ;
  assign n34079 = ~n33764 & ~n34078 ;
  assign n34080 = n33764 & n34078 ;
  assign n34081 = ~\P1_P1_InstAddrPointer_reg[0]/NET0131  & ~n33797 ;
  assign n34082 = ~n34080 & n34081 ;
  assign n34083 = ~n34079 & ~n34082 ;
  assign n34084 = ~n34076 & ~n34083 ;
  assign n34085 = ~n34075 & ~n34084 ;
  assign n34086 = ~n34074 & ~n34085 ;
  assign n34087 = ~n34073 & ~n34086 ;
  assign n34088 = ~n34070 & ~n34087 ;
  assign n34089 = ~n34069 & ~n34088 ;
  assign n34090 = ~n34066 & ~n34089 ;
  assign n34091 = ~n34065 & ~n34090 ;
  assign n34092 = ~n34062 & ~n34091 ;
  assign n34093 = ~n34061 & ~n34092 ;
  assign n34094 = ~n34058 & ~n34093 ;
  assign n34095 = ~n34057 & ~n34094 ;
  assign n34096 = n34054 & ~n34095 ;
  assign n34097 = \P1_P1_InstAddrPointer_reg[9]/NET0131  & n34096 ;
  assign n34098 = n34052 & n34097 ;
  assign n34099 = n33520 & n34098 ;
  assign n34100 = n34050 & n34099 ;
  assign n34101 = \P1_P1_InstAddrPointer_reg[14]/NET0131  & n34100 ;
  assign n34102 = n34047 & n34101 ;
  assign n34103 = \P1_P1_InstAddrPointer_reg[16]/NET0131  & n34102 ;
  assign n34104 = \P1_P1_InstAddrPointer_reg[17]/NET0131  & n34033 ;
  assign n34105 = ~\P1_P1_InstAddrPointer_reg[17]/NET0131  & ~n34033 ;
  assign n34106 = ~n34104 & ~n34105 ;
  assign n34107 = n34103 & n34106 ;
  assign n34108 = n33517 & n34107 ;
  assign n34109 = n34045 & n34108 ;
  assign n34110 = \P1_P1_InstAddrPointer_reg[21]/NET0131  & n34109 ;
  assign n34111 = \P1_P1_InstAddrPointer_reg[21]/NET0131  & n34044 ;
  assign n34112 = ~\P1_P1_InstAddrPointer_reg[22]/NET0131  & ~n34111 ;
  assign n34113 = ~n34035 & ~n34112 ;
  assign n34114 = n34110 & n34113 ;
  assign n34115 = ~\P1_P1_InstAddrPointer_reg[23]/NET0131  & ~n34035 ;
  assign n34116 = n33840 & n34026 ;
  assign n34117 = ~n34115 & ~n34116 ;
  assign n34118 = n34114 & n34117 ;
  assign n34119 = ~\P1_P1_InstAddrPointer_reg[24]/NET0131  & ~n34116 ;
  assign n34120 = ~n34036 & ~n34119 ;
  assign n34121 = n34118 & n34120 ;
  assign n34122 = ~\P1_P1_InstAddrPointer_reg[25]/NET0131  & ~n34036 ;
  assign n34123 = ~n34037 & ~n34122 ;
  assign n34124 = n33539 & n34123 ;
  assign n34125 = n34121 & n34124 ;
  assign n34126 = n34042 & n34125 ;
  assign n34127 = \P1_P1_InstAddrPointer_reg[29]/NET0131  & n34126 ;
  assign n34128 = \P1_P1_InstAddrPointer_reg[29]/NET0131  & n34040 ;
  assign n34129 = \P1_P1_InstAddrPointer_reg[30]/NET0131  & n34128 ;
  assign n34130 = ~\P1_P1_InstAddrPointer_reg[30]/NET0131  & ~n34128 ;
  assign n34131 = ~n34129 & ~n34130 ;
  assign n34132 = n34127 & n34131 ;
  assign n34134 = \P1_P1_InstAddrPointer_reg[31]/NET0131  & ~n34129 ;
  assign n34135 = ~\P1_P1_InstAddrPointer_reg[31]/NET0131  & n34129 ;
  assign n34136 = ~n34134 & ~n34135 ;
  assign n34137 = ~n34132 & n34136 ;
  assign n34133 = \P1_P1_InstAddrPointer_reg[31]/NET0131  & n34132 ;
  assign n34138 = n26263 & ~n34133 ;
  assign n34139 = ~n34137 & n34138 ;
  assign n34150 = n15428 & n34136 ;
  assign n34151 = ~\P1_P1_InstAddrPointer_reg[31]/NET0131  & ~n15428 ;
  assign n34152 = ~n26123 & ~n34151 ;
  assign n34153 = ~n34150 & n34152 ;
  assign n34143 = ~n15335 & n33865 ;
  assign n34144 = ~n15383 & n26235 ;
  assign n34145 = ~n34143 & ~n34144 ;
  assign n34141 = n15364 & ~n15384 ;
  assign n34142 = ~n26176 & ~n34141 ;
  assign n34146 = ~n26251 & n34142 ;
  assign n34147 = ~n34145 & n34146 ;
  assign n34148 = \P1_P1_InstAddrPointer_reg[31]/NET0131  & ~n34147 ;
  assign n34140 = ~n26189 & ~n33865 ;
  assign n34149 = ~n26151 & n34013 ;
  assign n34154 = ~n34140 & ~n34149 ;
  assign n34155 = ~n34148 & n34154 ;
  assign n34156 = ~n34153 & n34155 ;
  assign n34157 = ~n34139 & n34156 ;
  assign n34158 = ~n34021 & n34157 ;
  assign n34159 = n8355 & ~n34158 ;
  assign n34160 = \P1_P1_rEIP_reg[31]/NET0131  & n8357 ;
  assign n34161 = n8348 & ~n8356 ;
  assign n34162 = ~n8281 & ~n8353 ;
  assign n34163 = ~n8287 & n34162 ;
  assign n34164 = ~n34161 & n34163 ;
  assign n34165 = \P1_P1_InstAddrPointer_reg[31]/NET0131  & ~n34164 ;
  assign n34166 = ~n34160 & ~n34165 ;
  assign n34167 = ~n34159 & n34166 ;
  assign n34168 = \P2_P1_uWord_reg[10]/NET0131  & ~n24913 ;
  assign n34170 = ~\P2_P1_EAX_reg[26]/NET0131  & ~n27397 ;
  assign n34171 = ~n27398 & ~n34170 ;
  assign n34172 = n24898 & n34171 ;
  assign n34173 = ~n21081 & n34172 ;
  assign n34169 = \P2_P1_uWord_reg[10]/NET0131  & ~n25154 ;
  assign n34174 = ~n23830 & ~n34169 ;
  assign n34175 = ~n34173 & n34174 ;
  assign n34176 = n11623 & ~n34175 ;
  assign n34177 = ~n34168 & ~n34176 ;
  assign n34178 = \P1_P1_uWord_reg[10]/NET0131  & ~n24515 ;
  assign n34182 = \P1_P1_uWord_reg[10]/NET0131  & n25363 ;
  assign n34183 = ~n23580 & ~n34182 ;
  assign n34184 = n15334 & ~n34183 ;
  assign n34179 = ~\P1_P1_EAX_reg[26]/NET0131  & ~n25356 ;
  assign n34180 = n24503 & ~n27426 ;
  assign n34181 = ~n34179 & n34180 ;
  assign n34185 = \P1_P1_uWord_reg[10]/NET0131  & n24505 ;
  assign n34186 = ~n34181 & ~n34185 ;
  assign n34187 = ~n34184 & n34186 ;
  assign n34188 = n8355 & ~n34187 ;
  assign n34189 = ~n34178 & ~n34188 ;
  assign n34191 = \P1_P2_InstAddrPointer_reg[30]/NET0131  & n25733 ;
  assign n34195 = ~n31189 & ~n31326 ;
  assign n34196 = ~n30809 & ~n31327 ;
  assign n34197 = ~n34195 & n34196 ;
  assign n34192 = ~n31169 & ~n31174 ;
  assign n34193 = ~n31175 & ~n34192 ;
  assign n34194 = n30809 & ~n34193 ;
  assign n34198 = ~n25733 & ~n34194 ;
  assign n34199 = ~n34197 & n34198 ;
  assign n34200 = ~n34191 & ~n34199 ;
  assign n34201 = n25701 & ~n34200 ;
  assign n34202 = n31357 & ~n31456 ;
  assign n34203 = n25881 & ~n31457 ;
  assign n34204 = ~n34202 & n34203 ;
  assign n34190 = ~n25817 & ~n31189 ;
  assign n34205 = n25887 & ~n31357 ;
  assign n34217 = ~n34190 & ~n34205 ;
  assign n34206 = ~n25752 & ~n25842 ;
  assign n34207 = n31466 & n34206 ;
  assign n34208 = ~n25748 & n34207 ;
  assign n34209 = n25415 & ~n25848 ;
  assign n34210 = n34208 & ~n34209 ;
  assign n34211 = \P1_P2_InstAddrPointer_reg[30]/NET0131  & ~n34210 ;
  assign n34212 = n25773 & n25774 ;
  assign n34213 = ~n25808 & ~n34212 ;
  assign n34214 = ~n25415 & ~n25848 ;
  assign n34215 = n34213 & ~n34214 ;
  assign n34216 = n31174 & ~n34215 ;
  assign n34218 = ~n34211 & ~n34216 ;
  assign n34219 = n34217 & n34218 ;
  assign n34220 = ~n34204 & n34219 ;
  assign n34221 = ~n34201 & n34220 ;
  assign n34222 = n25918 & ~n34221 ;
  assign n34223 = \P1_P2_rEIP_reg[30]/NET0131  & n27967 ;
  assign n34224 = \P1_P2_InstAddrPointer_reg[30]/NET0131  & ~n31487 ;
  assign n34225 = ~n34223 & ~n34224 ;
  assign n34226 = ~n34222 & n34225 ;
  assign n34227 = \P2_P1_InstAddrPointer_reg[30]/NET0131  & n25947 ;
  assign n34231 = ~n31523 & ~n31862 ;
  assign n34232 = ~n31863 & ~n34231 ;
  assign n34233 = n29503 & ~n34232 ;
  assign n34228 = ~n32009 & n32012 ;
  assign n34229 = ~n29503 & ~n32013 ;
  assign n34230 = ~n34228 & n34229 ;
  assign n34234 = ~n25947 & ~n34230 ;
  assign n34235 = ~n34233 & n34234 ;
  assign n34236 = ~n34227 & ~n34235 ;
  assign n34237 = n25945 & ~n34236 ;
  assign n34238 = ~\P2_P1_InstAddrPointer_reg[30]/NET0131  & ~n32150 ;
  assign n34239 = ~n32151 & ~n34238 ;
  assign n34241 = ~n32147 & ~n34239 ;
  assign n34242 = n25964 & ~n32148 ;
  assign n34243 = ~n34241 & n34242 ;
  assign n34247 = ~n25987 & ~n32150 ;
  assign n34248 = n32028 & ~n34247 ;
  assign n34249 = \P2_P1_InstAddrPointer_reg[30]/NET0131  & ~n34248 ;
  assign n34240 = n26068 & n34239 ;
  assign n34244 = ~n26031 & ~n31520 ;
  assign n34245 = n32159 & ~n34244 ;
  assign n34246 = n31523 & ~n34245 ;
  assign n34250 = ~n25995 & n32012 ;
  assign n34251 = ~n34246 & ~n34250 ;
  assign n34252 = ~n34240 & n34251 ;
  assign n34253 = ~n34249 & n34252 ;
  assign n34254 = ~n34243 & n34253 ;
  assign n34255 = ~n34237 & n34254 ;
  assign n34256 = n11623 & ~n34255 ;
  assign n34257 = \P2_P1_rEIP_reg[30]/NET0131  & n11616 ;
  assign n34258 = \P2_P1_InstAddrPointer_reg[30]/NET0131  & ~n32172 ;
  assign n34259 = ~n34257 & ~n34258 ;
  assign n34260 = ~n34256 & n34259 ;
  assign n34302 = ~n32749 & ~n32844 ;
  assign n34303 = n26744 & ~n32845 ;
  assign n34304 = ~n34302 & n34303 ;
  assign n34273 = \P2_P2_InstAddrPointer_reg[30]/NET0131  & n26629 ;
  assign n34277 = ~\P2_P2_InstAddrPointer_reg[14]/NET0131  & ~n32214 ;
  assign n34278 = ~n32196 & ~n34277 ;
  assign n34279 = ~\P2_P2_InstAddrPointer_reg[12]/NET0131  & ~n32579 ;
  assign n34280 = ~n32218 & ~n34279 ;
  assign n34281 = \P2_P2_InstAddrPointer_reg[11]/NET0131  & n32518 ;
  assign n34282 = n34280 & n34281 ;
  assign n34283 = \P2_P2_InstAddrPointer_reg[13]/NET0131  & n34282 ;
  assign n34284 = n34278 & n34283 ;
  assign n34285 = \P2_P2_InstAddrPointer_reg[15]/NET0131  & n34284 ;
  assign n34286 = n32527 & n34285 ;
  assign n34287 = n32531 & n34286 ;
  assign n34288 = \P2_P2_InstAddrPointer_reg[21]/NET0131  & n34287 ;
  assign n34289 = n32545 & n34288 ;
  assign n34290 = n32548 & n34289 ;
  assign n34291 = \P2_P2_InstAddrPointer_reg[26]/NET0131  & n34290 ;
  assign n34292 = n32210 & n34291 ;
  assign n34293 = n32208 & n34292 ;
  assign n34295 = ~n32555 & n34293 ;
  assign n34294 = n32555 & ~n34293 ;
  assign n34296 = n32510 & ~n34294 ;
  assign n34297 = ~n34295 & n34296 ;
  assign n34274 = ~n32708 & n32710 ;
  assign n34275 = ~n32510 & ~n32711 ;
  assign n34276 = ~n34274 & n34275 ;
  assign n34298 = ~n26629 & ~n34276 ;
  assign n34299 = ~n34297 & n34298 ;
  assign n34300 = ~n34273 & ~n34299 ;
  assign n34301 = n26621 & ~n34300 ;
  assign n34264 = ~n26641 & ~n26680 ;
  assign n34265 = ~n26619 & ~n32743 ;
  assign n34266 = ~n34264 & n34265 ;
  assign n34267 = ~n26612 & n34266 ;
  assign n34268 = ~n26583 & ~n32732 ;
  assign n34269 = n34267 & ~n34268 ;
  assign n34270 = \P2_P2_InstAddrPointer_reg[30]/NET0131  & ~n34269 ;
  assign n34263 = ~n26688 & n32710 ;
  assign n34271 = n26757 & n32749 ;
  assign n34272 = ~n26764 & n32555 ;
  assign n34305 = ~n34271 & ~n34272 ;
  assign n34306 = ~n34263 & n34305 ;
  assign n34307 = ~n34270 & n34306 ;
  assign n34308 = ~n34301 & n34307 ;
  assign n34309 = ~n34304 & n34308 ;
  assign n34310 = n26792 & ~n34309 ;
  assign n34261 = \P2_P2_InstAddrPointer_reg[30]/NET0131  & ~n32860 ;
  assign n34262 = \P2_P2_rEIP_reg[30]/NET0131  & n28046 ;
  assign n34311 = ~n34261 & ~n34262 ;
  assign n34312 = ~n34310 & n34311 ;
  assign n34313 = \P2_P3_InstAddrPointer_reg[30]/NET0131  & ~n27283 ;
  assign n34319 = ~n33297 & ~n33321 ;
  assign n34320 = n33300 & ~n34319 ;
  assign n34321 = ~n33323 & ~n34320 ;
  assign n34322 = n33289 & ~n34321 ;
  assign n34323 = n33242 & ~n34322 ;
  assign n34324 = ~n33289 & n34321 ;
  assign n34325 = ~n34323 & ~n34324 ;
  assign n34326 = ~n33330 & ~n34325 ;
  assign n34327 = n33337 & n34326 ;
  assign n34328 = ~n33286 & n34327 ;
  assign n34329 = ~n33342 & n34328 ;
  assign n34330 = n33350 & n34329 ;
  assign n34331 = n33358 & n34330 ;
  assign n34332 = n33380 & n34331 ;
  assign n34333 = ~n33383 & n34332 ;
  assign n34334 = ~n33279 & n34333 ;
  assign n34335 = ~n33388 & n34334 ;
  assign n34336 = ~n33392 & n34335 ;
  assign n34337 = ~n33396 & n34336 ;
  assign n34338 = ~n33400 & n34337 ;
  assign n34339 = ~n33404 & n34338 ;
  assign n34340 = ~n33407 & n34339 ;
  assign n34341 = n33410 & ~n34340 ;
  assign n34342 = ~n33242 & ~n33411 ;
  assign n34343 = ~n34341 & n34342 ;
  assign n34314 = ~\P2_P3_InstAddrPointer_reg[30]/NET0131  & ~n32928 ;
  assign n34315 = ~n32935 & ~n34314 ;
  assign n34316 = ~n33269 & ~n34315 ;
  assign n34317 = ~n33270 & ~n34316 ;
  assign n34318 = n33242 & ~n34317 ;
  assign n34344 = n27283 & ~n34318 ;
  assign n34345 = ~n34343 & n34344 ;
  assign n34346 = ~n34313 & ~n34345 ;
  assign n34347 = n27117 & ~n34346 ;
  assign n34348 = ~\P2_P3_InstAddrPointer_reg[30]/NET0131  & ~n32900 ;
  assign n34349 = ~n32901 & ~n34348 ;
  assign n34351 = ~n33500 & ~n34349 ;
  assign n34352 = n27280 & ~n33501 ;
  assign n34353 = ~n34351 & n34352 ;
  assign n34350 = n27219 & n34349 ;
  assign n34354 = ~n27142 & n33410 ;
  assign n34355 = n27236 & ~n27294 ;
  assign n34356 = \P2_P3_InstAddrPointer_reg[30]/NET0131  & ~n34355 ;
  assign n34357 = ~\P2_P3_InstAddrPointer_reg[30]/NET0131  & ~n27232 ;
  assign n34358 = ~n27180 & ~n34357 ;
  assign n34359 = ~n27057 & ~n27228 ;
  assign n34360 = ~n34358 & n34359 ;
  assign n34361 = n34315 & ~n34360 ;
  assign n34362 = ~n34356 & ~n34361 ;
  assign n34363 = ~n34354 & n34362 ;
  assign n34364 = ~n34350 & n34363 ;
  assign n34365 = ~n34353 & n34364 ;
  assign n34366 = ~n34347 & n34365 ;
  assign n34367 = n27308 & ~n34366 ;
  assign n34368 = \P2_P3_InstAddrPointer_reg[30]/NET0131  & ~n32870 ;
  assign n34369 = \P2_P3_rEIP_reg[30]/NET0131  & n32864 ;
  assign n34370 = ~n34368 & ~n34369 ;
  assign n34371 = ~n34367 & n34370 ;
  assign n34373 = \P1_P1_InstAddrPointer_reg[30]/NET0131  & n26249 ;
  assign n34377 = ~n34006 & n34009 ;
  assign n34378 = ~n29558 & ~n34010 ;
  assign n34379 = ~n34377 & n34378 ;
  assign n34374 = ~n33545 & ~n33861 ;
  assign n34375 = ~n33862 & ~n34374 ;
  assign n34376 = n29558 & ~n34375 ;
  assign n34380 = ~n26249 & ~n34376 ;
  assign n34381 = ~n34379 & n34380 ;
  assign n34382 = ~n34373 & ~n34381 ;
  assign n34383 = n26126 & ~n34382 ;
  assign n34384 = ~n34127 & ~n34131 ;
  assign n34385 = n26263 & ~n34132 ;
  assign n34386 = ~n34384 & n34385 ;
  assign n34387 = ~n15335 & ~n33545 ;
  assign n34388 = ~n26160 & ~n34387 ;
  assign n34389 = n26252 & n34142 ;
  assign n34390 = ~n26200 & n34389 ;
  assign n34391 = ~n34388 & n34390 ;
  assign n34392 = \P1_P1_InstAddrPointer_reg[30]/NET0131  & ~n34391 ;
  assign n34393 = n26192 & n34131 ;
  assign n34372 = ~n26189 & n33545 ;
  assign n34394 = ~n26151 & n34009 ;
  assign n34395 = ~n34372 & ~n34394 ;
  assign n34396 = ~n34393 & n34395 ;
  assign n34397 = ~n34392 & n34396 ;
  assign n34398 = ~n34386 & n34397 ;
  assign n34399 = ~n34383 & n34398 ;
  assign n34400 = n8355 & ~n34399 ;
  assign n34401 = \P1_P1_rEIP_reg[30]/NET0131  & n8357 ;
  assign n34402 = \P1_P1_InstAddrPointer_reg[30]/NET0131  & ~n34164 ;
  assign n34403 = ~n34401 & ~n34402 ;
  assign n34404 = ~n34400 & n34403 ;
  assign n34405 = ~n21062 & ~n24899 ;
  assign n34406 = ~n23161 & ~n34405 ;
  assign n34407 = n11623 & ~n34406 ;
  assign n34408 = n24913 & ~n34407 ;
  assign n34409 = \P2_P1_lWord_reg[7]/NET0131  & ~n34408 ;
  assign n34410 = n11387 & n23167 ;
  assign n34411 = \P2_P1_EAX_reg[7]/NET0131  & n24898 ;
  assign n34412 = ~n34410 & ~n34411 ;
  assign n34413 = n25161 & ~n34412 ;
  assign n34414 = ~n34409 & ~n34413 ;
  assign n34415 = \P2_P1_uWord_reg[9]/NET0131  & ~n24913 ;
  assign n34417 = ~\P2_P1_EAX_reg[25]/NET0131  & ~n27396 ;
  assign n34418 = n24899 & ~n27397 ;
  assign n34419 = ~n34417 & n34418 ;
  assign n34416 = \P2_P1_uWord_reg[9]/NET0131  & ~n25154 ;
  assign n34420 = ~n27889 & ~n34416 ;
  assign n34421 = ~n34419 & n34420 ;
  assign n34422 = n11623 & ~n34421 ;
  assign n34423 = ~n34415 & ~n34422 ;
  assign n34425 = \P1_P1_lWord_reg[7]/NET0131  & n15335 ;
  assign n34426 = ~n24133 & ~n34425 ;
  assign n34427 = n15334 & ~n34426 ;
  assign n34424 = \P1_P1_lWord_reg[7]/NET0131  & n24505 ;
  assign n34428 = \P1_P1_EAX_reg[7]/NET0131  & n24503 ;
  assign n34429 = ~n34424 & ~n34428 ;
  assign n34430 = ~n34427 & n34429 ;
  assign n34431 = n8355 & ~n34430 ;
  assign n34432 = \P1_P1_lWord_reg[7]/NET0131  & ~n24515 ;
  assign n34433 = ~n34431 & ~n34432 ;
  assign n34434 = \P1_P1_uWord_reg[9]/NET0131  & ~n24515 ;
  assign n34436 = n7955 & n15365 ;
  assign n34437 = \P1_P1_uWord_reg[9]/NET0131  & n25363 ;
  assign n34438 = ~n34436 & ~n34437 ;
  assign n34439 = n15334 & ~n34438 ;
  assign n34435 = \P1_P1_uWord_reg[9]/NET0131  & n24505 ;
  assign n34440 = ~\P1_P1_EAX_reg[25]/NET0131  & ~n27424 ;
  assign n34441 = ~n27425 & ~n34440 ;
  assign n34442 = n24503 & n34441 ;
  assign n34443 = ~n34435 & ~n34442 ;
  assign n34444 = ~n34439 & n34443 ;
  assign n34445 = n8355 & ~n34444 ;
  assign n34446 = ~n34434 & ~n34445 ;
  assign n34455 = \P1_buf2_reg[30]/NET0131  & ~n27934 ;
  assign n34456 = \P1_buf1_reg[30]/NET0131  & n27934 ;
  assign n34457 = ~n34455 & ~n34456 ;
  assign n34458 = n27945 & ~n34457 ;
  assign n34459 = \P1_buf2_reg[22]/NET0131  & ~n27934 ;
  assign n34460 = \P1_buf1_reg[22]/NET0131  & n27934 ;
  assign n34461 = ~n34459 & ~n34460 ;
  assign n34462 = n27952 & ~n34461 ;
  assign n34463 = ~n34458 & ~n34462 ;
  assign n34464 = \P1_P2_DataWidth_reg[1]/NET0131  & ~n34463 ;
  assign n34447 = \P1_buf2_reg[6]/NET0131  & ~n27934 ;
  assign n34448 = \P1_buf1_reg[6]/NET0131  & n27934 ;
  assign n34449 = ~n34447 & ~n34448 ;
  assign n34450 = ~n27905 & ~n34449 ;
  assign n34451 = \P1_P2_InstQueue_reg[11][6]/NET0131  & ~n27901 ;
  assign n34452 = ~n27904 & n34451 ;
  assign n34453 = ~n34450 & ~n34452 ;
  assign n34465 = ~n27960 & ~n34453 ;
  assign n34466 = ~n34464 & ~n34465 ;
  assign n34467 = n25928 & ~n34466 ;
  assign n34468 = ~n25571 & n27901 ;
  assign n34469 = ~n34451 & ~n34468 ;
  assign n34470 = n27608 & ~n34469 ;
  assign n34454 = n27898 & ~n34453 ;
  assign n34471 = \P1_P2_InstQueue_reg[11][6]/NET0131  & ~n27972 ;
  assign n34472 = ~n34454 & ~n34471 ;
  assign n34473 = ~n34470 & n34472 ;
  assign n34474 = ~n34467 & n34473 ;
  assign n34486 = \P2_buf2_reg[30]/NET0131  & ~n28013 ;
  assign n34487 = \P2_buf1_reg[30]/NET0131  & n28013 ;
  assign n34488 = ~n34486 & ~n34487 ;
  assign n34489 = n28027 & ~n34488 ;
  assign n34490 = \P2_buf2_reg[22]/NET0131  & ~n28013 ;
  assign n34491 = \P2_buf1_reg[22]/NET0131  & n28013 ;
  assign n34492 = ~n34490 & ~n34491 ;
  assign n34493 = n28034 & ~n34492 ;
  assign n34494 = ~n34489 & ~n34493 ;
  assign n34495 = \P2_P2_DataWidth_reg[1]/NET0131  & ~n34494 ;
  assign n34475 = \P2_buf2_reg[6]/NET0131  & ~n28013 ;
  assign n34476 = \P2_buf1_reg[6]/NET0131  & n28013 ;
  assign n34477 = ~n34475 & ~n34476 ;
  assign n34478 = ~n27984 & ~n34477 ;
  assign n34479 = \P2_P2_InstQueue_reg[11][6]/NET0131  & ~n27980 ;
  assign n34480 = ~n27983 & n34479 ;
  assign n34481 = ~n34478 & ~n34480 ;
  assign n34496 = ~n28042 & ~n34481 ;
  assign n34497 = ~n34495 & ~n34496 ;
  assign n34498 = n26794 & ~n34497 ;
  assign n34483 = ~n26385 & n27980 ;
  assign n34484 = ~n34479 & ~n34483 ;
  assign n34485 = n27613 & ~n34484 ;
  assign n34482 = n27977 & ~n34481 ;
  assign n34499 = \P2_P2_InstQueue_reg[11][6]/NET0131  & ~n28050 ;
  assign n34500 = ~n34482 & ~n34499 ;
  assign n34501 = ~n34485 & n34500 ;
  assign n34502 = ~n34498 & n34501 ;
  assign n34508 = n28065 & ~n34457 ;
  assign n34509 = n28068 & ~n34461 ;
  assign n34510 = ~n34508 & ~n34509 ;
  assign n34511 = \P1_P2_DataWidth_reg[1]/NET0131  & ~n34510 ;
  assign n34503 = ~n28058 & ~n34449 ;
  assign n34504 = \P1_P2_InstQueue_reg[0][6]/NET0131  & ~n28055 ;
  assign n34505 = ~n28057 & n34504 ;
  assign n34506 = ~n34503 & ~n34505 ;
  assign n34512 = ~n28073 & ~n34506 ;
  assign n34513 = ~n34511 & ~n34512 ;
  assign n34514 = n25928 & ~n34513 ;
  assign n34515 = ~n25571 & n28055 ;
  assign n34516 = ~n34504 & ~n34515 ;
  assign n34517 = n27608 & ~n34516 ;
  assign n34507 = n27898 & ~n34506 ;
  assign n34518 = \P1_P2_InstQueue_reg[0][6]/NET0131  & ~n27972 ;
  assign n34519 = ~n34507 & ~n34518 ;
  assign n34520 = ~n34517 & n34519 ;
  assign n34521 = ~n34514 & n34520 ;
  assign n34527 = n28090 & ~n34457 ;
  assign n34528 = n27945 & ~n34461 ;
  assign n34529 = ~n34527 & ~n34528 ;
  assign n34530 = \P1_P2_DataWidth_reg[1]/NET0131  & ~n34529 ;
  assign n34522 = ~n28084 & ~n34449 ;
  assign n34523 = \P1_P2_InstQueue_reg[10][6]/NET0131  & ~n27904 ;
  assign n34524 = ~n27952 & n34523 ;
  assign n34525 = ~n34522 & ~n34524 ;
  assign n34531 = ~n28096 & ~n34525 ;
  assign n34532 = ~n34530 & ~n34531 ;
  assign n34533 = n25928 & ~n34532 ;
  assign n34534 = ~n25571 & n27904 ;
  assign n34535 = ~n34523 & ~n34534 ;
  assign n34536 = n27608 & ~n34535 ;
  assign n34526 = n27898 & ~n34525 ;
  assign n34537 = \P1_P2_InstQueue_reg[10][6]/NET0131  & ~n27972 ;
  assign n34538 = ~n34526 & ~n34537 ;
  assign n34539 = ~n34536 & n34538 ;
  assign n34540 = ~n34533 & n34539 ;
  assign n34546 = n27952 & ~n34457 ;
  assign n34547 = n27904 & ~n34461 ;
  assign n34548 = ~n34546 & ~n34547 ;
  assign n34549 = \P1_P2_DataWidth_reg[1]/NET0131  & ~n34548 ;
  assign n34541 = ~n28109 & ~n34449 ;
  assign n34542 = \P1_P2_InstQueue_reg[12][6]/NET0131  & ~n28108 ;
  assign n34543 = ~n27901 & n34542 ;
  assign n34544 = ~n34541 & ~n34543 ;
  assign n34550 = ~n28119 & ~n34544 ;
  assign n34551 = ~n34549 & ~n34550 ;
  assign n34552 = n25928 & ~n34551 ;
  assign n34553 = ~n25571 & n28108 ;
  assign n34554 = ~n34542 & ~n34553 ;
  assign n34555 = n27608 & ~n34554 ;
  assign n34545 = n27898 & ~n34544 ;
  assign n34556 = \P1_P2_InstQueue_reg[12][6]/NET0131  & ~n27972 ;
  assign n34557 = ~n34545 & ~n34556 ;
  assign n34558 = ~n34555 & n34557 ;
  assign n34559 = ~n34552 & n34558 ;
  assign n34565 = n27904 & ~n34457 ;
  assign n34566 = n27901 & ~n34461 ;
  assign n34567 = ~n34565 & ~n34566 ;
  assign n34568 = \P1_P2_DataWidth_reg[1]/NET0131  & ~n34567 ;
  assign n34560 = ~n28130 & ~n34449 ;
  assign n34561 = \P1_P2_InstQueue_reg[13][6]/NET0131  & ~n28065 ;
  assign n34562 = ~n28108 & n34561 ;
  assign n34563 = ~n34560 & ~n34562 ;
  assign n34569 = ~n28140 & ~n34563 ;
  assign n34570 = ~n34568 & ~n34569 ;
  assign n34571 = n25928 & ~n34570 ;
  assign n34572 = ~n25571 & n28065 ;
  assign n34573 = ~n34561 & ~n34572 ;
  assign n34574 = n27608 & ~n34573 ;
  assign n34564 = n27898 & ~n34563 ;
  assign n34575 = \P1_P2_InstQueue_reg[13][6]/NET0131  & ~n27972 ;
  assign n34576 = ~n34564 & ~n34575 ;
  assign n34577 = ~n34574 & n34576 ;
  assign n34578 = ~n34571 & n34577 ;
  assign n34584 = n27901 & ~n34457 ;
  assign n34585 = n28108 & ~n34461 ;
  assign n34586 = ~n34584 & ~n34585 ;
  assign n34587 = \P1_P2_DataWidth_reg[1]/NET0131  & ~n34586 ;
  assign n34579 = ~n28072 & ~n34449 ;
  assign n34580 = \P1_P2_InstQueue_reg[14][6]/NET0131  & ~n28068 ;
  assign n34581 = ~n28065 & n34580 ;
  assign n34582 = ~n34579 & ~n34581 ;
  assign n34588 = ~n28160 & ~n34582 ;
  assign n34589 = ~n34587 & ~n34588 ;
  assign n34590 = n25928 & ~n34589 ;
  assign n34591 = ~n25571 & n28068 ;
  assign n34592 = ~n34580 & ~n34591 ;
  assign n34593 = n27608 & ~n34592 ;
  assign n34583 = n27898 & ~n34582 ;
  assign n34594 = \P1_P2_InstQueue_reg[14][6]/NET0131  & ~n27972 ;
  assign n34595 = ~n34583 & ~n34594 ;
  assign n34596 = ~n34593 & n34595 ;
  assign n34597 = ~n34590 & n34596 ;
  assign n34603 = n28108 & ~n34457 ;
  assign n34604 = n28065 & ~n34461 ;
  assign n34605 = ~n34603 & ~n34604 ;
  assign n34606 = \P1_P2_DataWidth_reg[1]/NET0131  & ~n34605 ;
  assign n34598 = ~n28171 & ~n34449 ;
  assign n34599 = \P1_P2_InstQueue_reg[15][6]/NET0131  & ~n28057 ;
  assign n34600 = ~n28068 & n34599 ;
  assign n34601 = ~n34598 & ~n34600 ;
  assign n34607 = ~n28181 & ~n34601 ;
  assign n34608 = ~n34606 & ~n34607 ;
  assign n34609 = n25928 & ~n34608 ;
  assign n34610 = ~n25571 & n28057 ;
  assign n34611 = ~n34599 & ~n34610 ;
  assign n34612 = n27608 & ~n34611 ;
  assign n34602 = n27898 & ~n34601 ;
  assign n34613 = \P1_P2_InstQueue_reg[15][6]/NET0131  & ~n27972 ;
  assign n34614 = ~n34602 & ~n34613 ;
  assign n34615 = ~n34612 & n34614 ;
  assign n34616 = ~n34609 & n34615 ;
  assign n34622 = n28068 & ~n34457 ;
  assign n34623 = n28057 & ~n34461 ;
  assign n34624 = ~n34622 & ~n34623 ;
  assign n34625 = \P1_P2_DataWidth_reg[1]/NET0131  & ~n34624 ;
  assign n34617 = ~n28193 & ~n34449 ;
  assign n34618 = \P1_P2_InstQueue_reg[1][6]/NET0131  & ~n28192 ;
  assign n34619 = ~n28055 & n34618 ;
  assign n34620 = ~n34617 & ~n34619 ;
  assign n34626 = ~n28203 & ~n34620 ;
  assign n34627 = ~n34625 & ~n34626 ;
  assign n34628 = n25928 & ~n34627 ;
  assign n34629 = ~n25571 & n28192 ;
  assign n34630 = ~n34618 & ~n34629 ;
  assign n34631 = n27608 & ~n34630 ;
  assign n34621 = n27898 & ~n34620 ;
  assign n34632 = \P1_P2_InstQueue_reg[1][6]/NET0131  & ~n27972 ;
  assign n34633 = ~n34621 & ~n34632 ;
  assign n34634 = ~n34631 & n34633 ;
  assign n34635 = ~n34628 & n34634 ;
  assign n34641 = n28057 & ~n34457 ;
  assign n34642 = n28055 & ~n34461 ;
  assign n34643 = ~n34641 & ~n34642 ;
  assign n34644 = \P1_P2_DataWidth_reg[1]/NET0131  & ~n34643 ;
  assign n34636 = ~n28215 & ~n34449 ;
  assign n34637 = \P1_P2_InstQueue_reg[2][6]/NET0131  & ~n28214 ;
  assign n34638 = ~n28192 & n34637 ;
  assign n34639 = ~n34636 & ~n34638 ;
  assign n34645 = ~n28225 & ~n34639 ;
  assign n34646 = ~n34644 & ~n34645 ;
  assign n34647 = n25928 & ~n34646 ;
  assign n34648 = ~n25571 & n28214 ;
  assign n34649 = ~n34637 & ~n34648 ;
  assign n34650 = n27608 & ~n34649 ;
  assign n34640 = n27898 & ~n34639 ;
  assign n34651 = \P1_P2_InstQueue_reg[2][6]/NET0131  & ~n27972 ;
  assign n34652 = ~n34640 & ~n34651 ;
  assign n34653 = ~n34650 & n34652 ;
  assign n34654 = ~n34647 & n34653 ;
  assign n34660 = n28055 & ~n34457 ;
  assign n34661 = n28192 & ~n34461 ;
  assign n34662 = ~n34660 & ~n34661 ;
  assign n34663 = \P1_P2_DataWidth_reg[1]/NET0131  & ~n34662 ;
  assign n34655 = ~n28237 & ~n34449 ;
  assign n34656 = \P1_P2_InstQueue_reg[3][6]/NET0131  & ~n28236 ;
  assign n34657 = ~n28214 & n34656 ;
  assign n34658 = ~n34655 & ~n34657 ;
  assign n34664 = ~n28247 & ~n34658 ;
  assign n34665 = ~n34663 & ~n34664 ;
  assign n34666 = n25928 & ~n34665 ;
  assign n34667 = ~n25571 & n28236 ;
  assign n34668 = ~n34656 & ~n34667 ;
  assign n34669 = n27608 & ~n34668 ;
  assign n34659 = n27898 & ~n34658 ;
  assign n34670 = \P1_P2_InstQueue_reg[3][6]/NET0131  & ~n27972 ;
  assign n34671 = ~n34659 & ~n34670 ;
  assign n34672 = ~n34669 & n34671 ;
  assign n34673 = ~n34666 & n34672 ;
  assign n34679 = n28192 & ~n34457 ;
  assign n34680 = n28214 & ~n34461 ;
  assign n34681 = ~n34679 & ~n34680 ;
  assign n34682 = \P1_P2_DataWidth_reg[1]/NET0131  & ~n34681 ;
  assign n34674 = ~n28259 & ~n34449 ;
  assign n34675 = \P1_P2_InstQueue_reg[4][6]/NET0131  & ~n28258 ;
  assign n34676 = ~n28236 & n34675 ;
  assign n34677 = ~n34674 & ~n34676 ;
  assign n34683 = ~n28269 & ~n34677 ;
  assign n34684 = ~n34682 & ~n34683 ;
  assign n34685 = n25928 & ~n34684 ;
  assign n34686 = ~n25571 & n28258 ;
  assign n34687 = ~n34675 & ~n34686 ;
  assign n34688 = n27608 & ~n34687 ;
  assign n34678 = n27898 & ~n34677 ;
  assign n34689 = \P1_P2_InstQueue_reg[4][6]/NET0131  & ~n27972 ;
  assign n34690 = ~n34678 & ~n34689 ;
  assign n34691 = ~n34688 & n34690 ;
  assign n34692 = ~n34685 & n34691 ;
  assign n34698 = n28214 & ~n34457 ;
  assign n34699 = n28236 & ~n34461 ;
  assign n34700 = ~n34698 & ~n34699 ;
  assign n34701 = \P1_P2_DataWidth_reg[1]/NET0131  & ~n34700 ;
  assign n34693 = ~n28281 & ~n34449 ;
  assign n34694 = \P1_P2_InstQueue_reg[5][6]/NET0131  & ~n28280 ;
  assign n34695 = ~n28258 & n34694 ;
  assign n34696 = ~n34693 & ~n34695 ;
  assign n34702 = ~n28291 & ~n34696 ;
  assign n34703 = ~n34701 & ~n34702 ;
  assign n34704 = n25928 & ~n34703 ;
  assign n34705 = ~n25571 & n28280 ;
  assign n34706 = ~n34694 & ~n34705 ;
  assign n34707 = n27608 & ~n34706 ;
  assign n34697 = n27898 & ~n34696 ;
  assign n34708 = \P1_P2_InstQueue_reg[5][6]/NET0131  & ~n27972 ;
  assign n34709 = ~n34697 & ~n34708 ;
  assign n34710 = ~n34707 & n34709 ;
  assign n34711 = ~n34704 & n34710 ;
  assign n34717 = n28236 & ~n34457 ;
  assign n34718 = n28258 & ~n34461 ;
  assign n34719 = ~n34717 & ~n34718 ;
  assign n34720 = \P1_P2_DataWidth_reg[1]/NET0131  & ~n34719 ;
  assign n34712 = ~n28303 & ~n34449 ;
  assign n34713 = \P1_P2_InstQueue_reg[6][6]/NET0131  & ~n28302 ;
  assign n34714 = ~n28280 & n34713 ;
  assign n34715 = ~n34712 & ~n34714 ;
  assign n34721 = ~n28313 & ~n34715 ;
  assign n34722 = ~n34720 & ~n34721 ;
  assign n34723 = n25928 & ~n34722 ;
  assign n34724 = ~n25571 & n28302 ;
  assign n34725 = ~n34713 & ~n34724 ;
  assign n34726 = n27608 & ~n34725 ;
  assign n34716 = n27898 & ~n34715 ;
  assign n34727 = \P1_P2_InstQueue_reg[6][6]/NET0131  & ~n27972 ;
  assign n34728 = ~n34716 & ~n34727 ;
  assign n34729 = ~n34726 & n34728 ;
  assign n34730 = ~n34723 & n34729 ;
  assign n34736 = n28258 & ~n34457 ;
  assign n34737 = n28280 & ~n34461 ;
  assign n34738 = ~n34736 & ~n34737 ;
  assign n34739 = \P1_P2_DataWidth_reg[1]/NET0131  & ~n34738 ;
  assign n34731 = ~n28324 & ~n34449 ;
  assign n34732 = \P1_P2_InstQueue_reg[7][6]/NET0131  & ~n28090 ;
  assign n34733 = ~n28302 & n34732 ;
  assign n34734 = ~n34731 & ~n34733 ;
  assign n34740 = ~n28334 & ~n34734 ;
  assign n34741 = ~n34739 & ~n34740 ;
  assign n34742 = n25928 & ~n34741 ;
  assign n34743 = ~n25571 & n28090 ;
  assign n34744 = ~n34732 & ~n34743 ;
  assign n34745 = n27608 & ~n34744 ;
  assign n34735 = n27898 & ~n34734 ;
  assign n34746 = \P1_P2_InstQueue_reg[7][6]/NET0131  & ~n27972 ;
  assign n34747 = ~n34735 & ~n34746 ;
  assign n34748 = ~n34745 & n34747 ;
  assign n34749 = ~n34742 & n34748 ;
  assign n34755 = n28280 & ~n34457 ;
  assign n34756 = n28302 & ~n34461 ;
  assign n34757 = ~n34755 & ~n34756 ;
  assign n34758 = \P1_P2_DataWidth_reg[1]/NET0131  & ~n34757 ;
  assign n34750 = ~n28095 & ~n34449 ;
  assign n34751 = \P1_P2_InstQueue_reg[8][6]/NET0131  & ~n27945 ;
  assign n34752 = ~n28090 & n34751 ;
  assign n34753 = ~n34750 & ~n34752 ;
  assign n34759 = ~n28354 & ~n34753 ;
  assign n34760 = ~n34758 & ~n34759 ;
  assign n34761 = n25928 & ~n34760 ;
  assign n34762 = ~n25571 & n27945 ;
  assign n34763 = ~n34751 & ~n34762 ;
  assign n34764 = n27608 & ~n34763 ;
  assign n34754 = n27898 & ~n34753 ;
  assign n34765 = \P1_P2_InstQueue_reg[8][6]/NET0131  & ~n27972 ;
  assign n34766 = ~n34754 & ~n34765 ;
  assign n34767 = ~n34764 & n34766 ;
  assign n34768 = ~n34761 & n34767 ;
  assign n34774 = n28302 & ~n34457 ;
  assign n34775 = n28090 & ~n34461 ;
  assign n34776 = ~n34774 & ~n34775 ;
  assign n34777 = \P1_P2_DataWidth_reg[1]/NET0131  & ~n34776 ;
  assign n34769 = ~n27959 & ~n34449 ;
  assign n34770 = \P1_P2_InstQueue_reg[9][6]/NET0131  & ~n27952 ;
  assign n34771 = ~n27945 & n34770 ;
  assign n34772 = ~n34769 & ~n34771 ;
  assign n34778 = ~n28374 & ~n34772 ;
  assign n34779 = ~n34777 & ~n34778 ;
  assign n34780 = n25928 & ~n34779 ;
  assign n34781 = ~n25571 & n27952 ;
  assign n34782 = ~n34770 & ~n34781 ;
  assign n34783 = n27608 & ~n34782 ;
  assign n34773 = n27898 & ~n34772 ;
  assign n34784 = \P1_P2_InstQueue_reg[9][6]/NET0131  & ~n27972 ;
  assign n34785 = ~n34773 & ~n34784 ;
  assign n34786 = ~n34783 & n34785 ;
  assign n34787 = ~n34780 & n34786 ;
  assign n34796 = n28398 & ~n34488 ;
  assign n34797 = n28401 & ~n34492 ;
  assign n34798 = ~n34796 & ~n34797 ;
  assign n34799 = \P2_P2_DataWidth_reg[1]/NET0131  & ~n34798 ;
  assign n34788 = ~n28388 & ~n34477 ;
  assign n34789 = \P2_P2_InstQueue_reg[0][6]/NET0131  & ~n28385 ;
  assign n34790 = ~n28387 & n34789 ;
  assign n34791 = ~n34788 & ~n34790 ;
  assign n34800 = ~n28406 & ~n34791 ;
  assign n34801 = ~n34799 & ~n34800 ;
  assign n34802 = n26794 & ~n34801 ;
  assign n34793 = ~n26385 & n28385 ;
  assign n34794 = ~n34789 & ~n34793 ;
  assign n34795 = n27613 & ~n34794 ;
  assign n34792 = n27977 & ~n34791 ;
  assign n34803 = \P2_P2_InstQueue_reg[0][6]/NET0131  & ~n28050 ;
  assign n34804 = ~n34792 & ~n34803 ;
  assign n34805 = ~n34795 & n34804 ;
  assign n34806 = ~n34802 & n34805 ;
  assign n34815 = n28423 & ~n34488 ;
  assign n34816 = n28027 & ~n34492 ;
  assign n34817 = ~n34815 & ~n34816 ;
  assign n34818 = \P2_P2_DataWidth_reg[1]/NET0131  & ~n34817 ;
  assign n34807 = ~n28414 & ~n34477 ;
  assign n34808 = \P2_P2_InstQueue_reg[10][6]/NET0131  & ~n27983 ;
  assign n34809 = ~n28034 & n34808 ;
  assign n34810 = ~n34807 & ~n34809 ;
  assign n34819 = ~n28429 & ~n34810 ;
  assign n34820 = ~n34818 & ~n34819 ;
  assign n34821 = n26794 & ~n34820 ;
  assign n34812 = ~n26385 & n27983 ;
  assign n34813 = ~n34808 & ~n34812 ;
  assign n34814 = n27613 & ~n34813 ;
  assign n34811 = n27977 & ~n34810 ;
  assign n34822 = \P2_P2_InstQueue_reg[10][6]/NET0131  & ~n28050 ;
  assign n34823 = ~n34811 & ~n34822 ;
  assign n34824 = ~n34814 & n34823 ;
  assign n34825 = ~n34821 & n34824 ;
  assign n34834 = n28034 & ~n34488 ;
  assign n34835 = n27983 & ~n34492 ;
  assign n34836 = ~n34834 & ~n34835 ;
  assign n34837 = \P2_P2_DataWidth_reg[1]/NET0131  & ~n34836 ;
  assign n34826 = ~n28439 & ~n34477 ;
  assign n34827 = \P2_P2_InstQueue_reg[12][6]/NET0131  & ~n28438 ;
  assign n34828 = ~n27980 & n34827 ;
  assign n34829 = ~n34826 & ~n34828 ;
  assign n34838 = ~n28452 & ~n34829 ;
  assign n34839 = ~n34837 & ~n34838 ;
  assign n34840 = n26794 & ~n34839 ;
  assign n34831 = ~n26385 & n28438 ;
  assign n34832 = ~n34827 & ~n34831 ;
  assign n34833 = n27613 & ~n34832 ;
  assign n34830 = n27977 & ~n34829 ;
  assign n34841 = \P2_P2_InstQueue_reg[12][6]/NET0131  & ~n28050 ;
  assign n34842 = ~n34830 & ~n34841 ;
  assign n34843 = ~n34833 & n34842 ;
  assign n34844 = ~n34840 & n34843 ;
  assign n34853 = n27983 & ~n34488 ;
  assign n34854 = n27980 & ~n34492 ;
  assign n34855 = ~n34853 & ~n34854 ;
  assign n34856 = \P2_P2_DataWidth_reg[1]/NET0131  & ~n34855 ;
  assign n34845 = ~n28460 & ~n34477 ;
  assign n34846 = \P2_P2_InstQueue_reg[13][6]/NET0131  & ~n28398 ;
  assign n34847 = ~n28438 & n34846 ;
  assign n34848 = ~n34845 & ~n34847 ;
  assign n34857 = ~n28473 & ~n34848 ;
  assign n34858 = ~n34856 & ~n34857 ;
  assign n34859 = n26794 & ~n34858 ;
  assign n34850 = ~n26385 & n28398 ;
  assign n34851 = ~n34846 & ~n34850 ;
  assign n34852 = n27613 & ~n34851 ;
  assign n34849 = n27977 & ~n34848 ;
  assign n34860 = \P2_P2_InstQueue_reg[13][6]/NET0131  & ~n28050 ;
  assign n34861 = ~n34849 & ~n34860 ;
  assign n34862 = ~n34852 & n34861 ;
  assign n34863 = ~n34859 & n34862 ;
  assign n34872 = n27980 & ~n34488 ;
  assign n34873 = n28438 & ~n34492 ;
  assign n34874 = ~n34872 & ~n34873 ;
  assign n34875 = \P2_P2_DataWidth_reg[1]/NET0131  & ~n34874 ;
  assign n34864 = ~n28405 & ~n34477 ;
  assign n34865 = \P2_P2_InstQueue_reg[14][6]/NET0131  & ~n28401 ;
  assign n34866 = ~n28398 & n34865 ;
  assign n34867 = ~n34864 & ~n34866 ;
  assign n34876 = ~n28493 & ~n34867 ;
  assign n34877 = ~n34875 & ~n34876 ;
  assign n34878 = n26794 & ~n34877 ;
  assign n34869 = ~n26385 & n28401 ;
  assign n34870 = ~n34865 & ~n34869 ;
  assign n34871 = n27613 & ~n34870 ;
  assign n34868 = n27977 & ~n34867 ;
  assign n34879 = \P2_P2_InstQueue_reg[14][6]/NET0131  & ~n28050 ;
  assign n34880 = ~n34868 & ~n34879 ;
  assign n34881 = ~n34871 & n34880 ;
  assign n34882 = ~n34878 & n34881 ;
  assign n34891 = n28438 & ~n34488 ;
  assign n34892 = n28398 & ~n34492 ;
  assign n34893 = ~n34891 & ~n34892 ;
  assign n34894 = \P2_P2_DataWidth_reg[1]/NET0131  & ~n34893 ;
  assign n34883 = ~n28501 & ~n34477 ;
  assign n34884 = \P2_P2_InstQueue_reg[15][6]/NET0131  & ~n28387 ;
  assign n34885 = ~n28401 & n34884 ;
  assign n34886 = ~n34883 & ~n34885 ;
  assign n34895 = ~n28514 & ~n34886 ;
  assign n34896 = ~n34894 & ~n34895 ;
  assign n34897 = n26794 & ~n34896 ;
  assign n34888 = ~n26385 & n28387 ;
  assign n34889 = ~n34884 & ~n34888 ;
  assign n34890 = n27613 & ~n34889 ;
  assign n34887 = n27977 & ~n34886 ;
  assign n34898 = \P2_P2_InstQueue_reg[15][6]/NET0131  & ~n28050 ;
  assign n34899 = ~n34887 & ~n34898 ;
  assign n34900 = ~n34890 & n34899 ;
  assign n34901 = ~n34897 & n34900 ;
  assign n34910 = n28401 & ~n34488 ;
  assign n34911 = n28387 & ~n34492 ;
  assign n34912 = ~n34910 & ~n34911 ;
  assign n34913 = \P2_P2_DataWidth_reg[1]/NET0131  & ~n34912 ;
  assign n34902 = ~n28523 & ~n34477 ;
  assign n34903 = \P2_P2_InstQueue_reg[1][6]/NET0131  & ~n28522 ;
  assign n34904 = ~n28385 & n34903 ;
  assign n34905 = ~n34902 & ~n34904 ;
  assign n34914 = ~n28536 & ~n34905 ;
  assign n34915 = ~n34913 & ~n34914 ;
  assign n34916 = n26794 & ~n34915 ;
  assign n34907 = ~n26385 & n28522 ;
  assign n34908 = ~n34903 & ~n34907 ;
  assign n34909 = n27613 & ~n34908 ;
  assign n34906 = n27977 & ~n34905 ;
  assign n34917 = \P2_P2_InstQueue_reg[1][6]/NET0131  & ~n28050 ;
  assign n34918 = ~n34906 & ~n34917 ;
  assign n34919 = ~n34909 & n34918 ;
  assign n34920 = ~n34916 & n34919 ;
  assign n34929 = n28387 & ~n34488 ;
  assign n34930 = n28385 & ~n34492 ;
  assign n34931 = ~n34929 & ~n34930 ;
  assign n34932 = \P2_P2_DataWidth_reg[1]/NET0131  & ~n34931 ;
  assign n34921 = ~n28545 & ~n34477 ;
  assign n34922 = \P2_P2_InstQueue_reg[2][6]/NET0131  & ~n28544 ;
  assign n34923 = ~n28522 & n34922 ;
  assign n34924 = ~n34921 & ~n34923 ;
  assign n34933 = ~n28558 & ~n34924 ;
  assign n34934 = ~n34932 & ~n34933 ;
  assign n34935 = n26794 & ~n34934 ;
  assign n34926 = ~n26385 & n28544 ;
  assign n34927 = ~n34922 & ~n34926 ;
  assign n34928 = n27613 & ~n34927 ;
  assign n34925 = n27977 & ~n34924 ;
  assign n34936 = \P2_P2_InstQueue_reg[2][6]/NET0131  & ~n28050 ;
  assign n34937 = ~n34925 & ~n34936 ;
  assign n34938 = ~n34928 & n34937 ;
  assign n34939 = ~n34935 & n34938 ;
  assign n34948 = n28385 & ~n34488 ;
  assign n34949 = n28522 & ~n34492 ;
  assign n34950 = ~n34948 & ~n34949 ;
  assign n34951 = \P2_P2_DataWidth_reg[1]/NET0131  & ~n34950 ;
  assign n34940 = ~n28567 & ~n34477 ;
  assign n34941 = \P2_P2_InstQueue_reg[3][6]/NET0131  & ~n28566 ;
  assign n34942 = ~n28544 & n34941 ;
  assign n34943 = ~n34940 & ~n34942 ;
  assign n34952 = ~n28580 & ~n34943 ;
  assign n34953 = ~n34951 & ~n34952 ;
  assign n34954 = n26794 & ~n34953 ;
  assign n34945 = ~n26385 & n28566 ;
  assign n34946 = ~n34941 & ~n34945 ;
  assign n34947 = n27613 & ~n34946 ;
  assign n34944 = n27977 & ~n34943 ;
  assign n34955 = \P2_P2_InstQueue_reg[3][6]/NET0131  & ~n28050 ;
  assign n34956 = ~n34944 & ~n34955 ;
  assign n34957 = ~n34947 & n34956 ;
  assign n34958 = ~n34954 & n34957 ;
  assign n34967 = n28522 & ~n34488 ;
  assign n34968 = n28544 & ~n34492 ;
  assign n34969 = ~n34967 & ~n34968 ;
  assign n34970 = \P2_P2_DataWidth_reg[1]/NET0131  & ~n34969 ;
  assign n34959 = ~n28589 & ~n34477 ;
  assign n34960 = \P2_P2_InstQueue_reg[4][6]/NET0131  & ~n28588 ;
  assign n34961 = ~n28566 & n34960 ;
  assign n34962 = ~n34959 & ~n34961 ;
  assign n34971 = ~n28602 & ~n34962 ;
  assign n34972 = ~n34970 & ~n34971 ;
  assign n34973 = n26794 & ~n34972 ;
  assign n34964 = ~n26385 & n28588 ;
  assign n34965 = ~n34960 & ~n34964 ;
  assign n34966 = n27613 & ~n34965 ;
  assign n34963 = n27977 & ~n34962 ;
  assign n34974 = \P2_P2_InstQueue_reg[4][6]/NET0131  & ~n28050 ;
  assign n34975 = ~n34963 & ~n34974 ;
  assign n34976 = ~n34966 & n34975 ;
  assign n34977 = ~n34973 & n34976 ;
  assign n34986 = n28544 & ~n34488 ;
  assign n34987 = n28566 & ~n34492 ;
  assign n34988 = ~n34986 & ~n34987 ;
  assign n34989 = \P2_P2_DataWidth_reg[1]/NET0131  & ~n34988 ;
  assign n34978 = ~n28611 & ~n34477 ;
  assign n34979 = \P2_P2_InstQueue_reg[5][6]/NET0131  & ~n28610 ;
  assign n34980 = ~n28588 & n34979 ;
  assign n34981 = ~n34978 & ~n34980 ;
  assign n34990 = ~n28624 & ~n34981 ;
  assign n34991 = ~n34989 & ~n34990 ;
  assign n34992 = n26794 & ~n34991 ;
  assign n34983 = ~n26385 & n28610 ;
  assign n34984 = ~n34979 & ~n34983 ;
  assign n34985 = n27613 & ~n34984 ;
  assign n34982 = n27977 & ~n34981 ;
  assign n34993 = \P2_P2_InstQueue_reg[5][6]/NET0131  & ~n28050 ;
  assign n34994 = ~n34982 & ~n34993 ;
  assign n34995 = ~n34985 & n34994 ;
  assign n34996 = ~n34992 & n34995 ;
  assign n35005 = n28566 & ~n34488 ;
  assign n35006 = n28588 & ~n34492 ;
  assign n35007 = ~n35005 & ~n35006 ;
  assign n35008 = \P2_P2_DataWidth_reg[1]/NET0131  & ~n35007 ;
  assign n34997 = ~n28633 & ~n34477 ;
  assign n34998 = \P2_P2_InstQueue_reg[6][6]/NET0131  & ~n28632 ;
  assign n34999 = ~n28610 & n34998 ;
  assign n35000 = ~n34997 & ~n34999 ;
  assign n35009 = ~n28646 & ~n35000 ;
  assign n35010 = ~n35008 & ~n35009 ;
  assign n35011 = n26794 & ~n35010 ;
  assign n35002 = ~n26385 & n28632 ;
  assign n35003 = ~n34998 & ~n35002 ;
  assign n35004 = n27613 & ~n35003 ;
  assign n35001 = n27977 & ~n35000 ;
  assign n35012 = \P2_P2_InstQueue_reg[6][6]/NET0131  & ~n28050 ;
  assign n35013 = ~n35001 & ~n35012 ;
  assign n35014 = ~n35004 & n35013 ;
  assign n35015 = ~n35011 & n35014 ;
  assign n35024 = n28588 & ~n34488 ;
  assign n35025 = n28610 & ~n34492 ;
  assign n35026 = ~n35024 & ~n35025 ;
  assign n35027 = \P2_P2_DataWidth_reg[1]/NET0131  & ~n35026 ;
  assign n35016 = ~n28654 & ~n34477 ;
  assign n35017 = \P2_P2_InstQueue_reg[7][6]/NET0131  & ~n28423 ;
  assign n35018 = ~n28632 & n35017 ;
  assign n35019 = ~n35016 & ~n35018 ;
  assign n35028 = ~n28667 & ~n35019 ;
  assign n35029 = ~n35027 & ~n35028 ;
  assign n35030 = n26794 & ~n35029 ;
  assign n35021 = ~n26385 & n28423 ;
  assign n35022 = ~n35017 & ~n35021 ;
  assign n35023 = n27613 & ~n35022 ;
  assign n35020 = n27977 & ~n35019 ;
  assign n35031 = \P2_P2_InstQueue_reg[7][6]/NET0131  & ~n28050 ;
  assign n35032 = ~n35020 & ~n35031 ;
  assign n35033 = ~n35023 & n35032 ;
  assign n35034 = ~n35030 & n35033 ;
  assign n35043 = n28610 & ~n34488 ;
  assign n35044 = n28632 & ~n34492 ;
  assign n35045 = ~n35043 & ~n35044 ;
  assign n35046 = \P2_P2_DataWidth_reg[1]/NET0131  & ~n35045 ;
  assign n35035 = ~n28428 & ~n34477 ;
  assign n35036 = \P2_P2_InstQueue_reg[8][6]/NET0131  & ~n28027 ;
  assign n35037 = ~n28423 & n35036 ;
  assign n35038 = ~n35035 & ~n35037 ;
  assign n35047 = ~n28687 & ~n35038 ;
  assign n35048 = ~n35046 & ~n35047 ;
  assign n35049 = n26794 & ~n35048 ;
  assign n35040 = ~n26385 & n28027 ;
  assign n35041 = ~n35036 & ~n35040 ;
  assign n35042 = n27613 & ~n35041 ;
  assign n35039 = n27977 & ~n35038 ;
  assign n35050 = \P2_P2_InstQueue_reg[8][6]/NET0131  & ~n28050 ;
  assign n35051 = ~n35039 & ~n35050 ;
  assign n35052 = ~n35042 & n35051 ;
  assign n35053 = ~n35049 & n35052 ;
  assign n35062 = n28632 & ~n34488 ;
  assign n35063 = n28423 & ~n34492 ;
  assign n35064 = ~n35062 & ~n35063 ;
  assign n35065 = \P2_P2_DataWidth_reg[1]/NET0131  & ~n35064 ;
  assign n35054 = ~n28041 & ~n34477 ;
  assign n35055 = \P2_P2_InstQueue_reg[9][6]/NET0131  & ~n28034 ;
  assign n35056 = ~n28027 & n35055 ;
  assign n35057 = ~n35054 & ~n35056 ;
  assign n35066 = ~n28707 & ~n35057 ;
  assign n35067 = ~n35065 & ~n35066 ;
  assign n35068 = n26794 & ~n35067 ;
  assign n35059 = ~n26385 & n28034 ;
  assign n35060 = ~n35055 & ~n35059 ;
  assign n35061 = n27613 & ~n35060 ;
  assign n35058 = n27977 & ~n35057 ;
  assign n35069 = \P2_P2_InstQueue_reg[9][6]/NET0131  & ~n28050 ;
  assign n35070 = ~n35058 & ~n35069 ;
  assign n35071 = ~n35061 & n35070 ;
  assign n35072 = ~n35068 & n35071 ;
  assign n35075 = \P1_P2_InstAddrPointer_reg[23]/NET0131  & n25733 ;
  assign n35082 = n31295 & ~n31302 ;
  assign n35081 = ~n31295 & n31302 ;
  assign n35083 = ~n30809 & ~n35081 ;
  assign n35084 = ~n35082 & n35083 ;
  assign n35076 = \P1_P2_InstAddrPointer_reg[22]/NET0131  & n31143 ;
  assign n35077 = ~n31149 & ~n35076 ;
  assign n35078 = \P1_P2_InstAddrPointer_reg[23]/NET0131  & n35076 ;
  assign n35079 = ~n35077 & ~n35078 ;
  assign n35080 = n30809 & ~n35079 ;
  assign n35085 = ~n25733 & ~n35080 ;
  assign n35086 = ~n35084 & n35085 ;
  assign n35087 = ~n35075 & ~n35086 ;
  assign n35088 = n25701 & ~n35087 ;
  assign n35089 = ~\P1_P2_InstAddrPointer_reg[23]/NET0131  & ~n31434 ;
  assign n35090 = ~n31342 & ~n35089 ;
  assign n35091 = ~n31437 & ~n35090 ;
  assign n35092 = n25881 & ~n31438 ;
  assign n35093 = ~n35091 & n35092 ;
  assign n35074 = \P1_P2_InstAddrPointer_reg[23]/NET0131  & ~n34210 ;
  assign n35095 = n25887 & n35090 ;
  assign n35097 = ~n35074 & ~n35095 ;
  assign n35094 = ~n25817 & n31302 ;
  assign n35096 = n31149 & ~n34215 ;
  assign n35098 = ~n35094 & ~n35096 ;
  assign n35099 = n35097 & n35098 ;
  assign n35100 = ~n35093 & n35099 ;
  assign n35101 = ~n35088 & n35100 ;
  assign n35102 = n25918 & ~n35101 ;
  assign n35073 = \P1_P2_InstAddrPointer_reg[23]/NET0131  & ~n31487 ;
  assign n35103 = \P1_P2_rEIP_reg[23]/NET0131  & n27967 ;
  assign n35104 = ~n35073 & ~n35103 ;
  assign n35105 = ~n35102 & n35104 ;
  assign n35109 = \P1_P2_InstAddrPointer_reg[27]/NET0131  & n25733 ;
  assign n35115 = n31310 & n31317 ;
  assign n35117 = ~n31322 & n35115 ;
  assign n35116 = n31322 & ~n35115 ;
  assign n35118 = ~n30809 & ~n35116 ;
  assign n35119 = ~n35117 & n35118 ;
  assign n35110 = n31155 & n31165 ;
  assign n35111 = n31158 & n35110 ;
  assign n35112 = ~n31158 & ~n35110 ;
  assign n35113 = ~n35111 & ~n35112 ;
  assign n35114 = n30809 & ~n35113 ;
  assign n35120 = ~n25733 & ~n35114 ;
  assign n35121 = ~n35119 & n35120 ;
  assign n35122 = ~n35109 & ~n35121 ;
  assign n35123 = n25701 & ~n35122 ;
  assign n35124 = ~\P1_P2_InstAddrPointer_reg[27]/NET0131  & ~n31344 ;
  assign n35125 = ~n31452 & ~n35124 ;
  assign n35126 = n31442 & n31445 ;
  assign n35127 = n31447 & n35126 ;
  assign n35128 = ~n35125 & ~n35127 ;
  assign n35129 = n25881 & ~n31450 ;
  assign n35130 = ~n35128 & n35129 ;
  assign n35134 = ~n25817 & n31322 ;
  assign n35108 = ~n25830 & n31158 ;
  assign n35131 = n25753 & n25779 ;
  assign n35132 = \P1_P2_InstAddrPointer_reg[27]/NET0131  & ~n35131 ;
  assign n35133 = n25887 & n35125 ;
  assign n35135 = ~n35132 & ~n35133 ;
  assign n35136 = ~n35108 & n35135 ;
  assign n35137 = ~n35134 & n35136 ;
  assign n35138 = ~n35130 & n35137 ;
  assign n35139 = ~n35123 & n35138 ;
  assign n35140 = n25918 & ~n35139 ;
  assign n35106 = \P1_P2_rEIP_reg[27]/NET0131  & n27967 ;
  assign n35107 = \P1_P2_InstAddrPointer_reg[27]/NET0131  & ~n31487 ;
  assign n35141 = ~n35106 & ~n35107 ;
  assign n35142 = ~n35140 & n35141 ;
  assign n35161 = \P1_P2_InstAddrPointer_reg[28]/NET0131  & n25733 ;
  assign n35162 = n31320 & ~n35117 ;
  assign n35163 = n31323 & n35115 ;
  assign n35164 = ~n30809 & ~n35163 ;
  assign n35165 = ~n35162 & n35164 ;
  assign n35147 = ~\P1_P2_InstAddrPointer_reg[28]/NET0131  & ~n31156 ;
  assign n35148 = ~n30836 & ~n35147 ;
  assign n35166 = ~n35111 & ~n35148 ;
  assign n35167 = ~n31168 & ~n35166 ;
  assign n35168 = n30809 & ~n35167 ;
  assign n35169 = ~n25733 & ~n35168 ;
  assign n35170 = ~n35165 & n35169 ;
  assign n35171 = ~n35161 & ~n35170 ;
  assign n35172 = n25701 & ~n35171 ;
  assign n35175 = ~\P1_P2_InstAddrPointer_reg[16]/NET0131  & ~n31358 ;
  assign n35176 = ~n31359 & ~n35175 ;
  assign n35177 = \P1_P2_InstAddrPointer_reg[15]/NET0131  & n31420 ;
  assign n35178 = n35176 & n35177 ;
  assign n35179 = n30818 & n31427 ;
  assign n35180 = n35178 & n35179 ;
  assign n35181 = n31363 & n35180 ;
  assign n35173 = ~\P1_P2_InstAddrPointer_reg[21]/NET0131  & ~n31362 ;
  assign n35174 = ~n31433 & ~n35173 ;
  assign n35182 = n30817 & n35174 ;
  assign n35183 = n35181 & n35182 ;
  assign n35184 = n31441 & n35183 ;
  assign n35185 = n31449 & n35184 ;
  assign n35187 = \P1_P2_InstAddrPointer_reg[28]/NET0131  & n35185 ;
  assign n35158 = ~\P1_P2_InstAddrPointer_reg[28]/NET0131  & ~n31452 ;
  assign n35159 = ~n31453 & ~n35158 ;
  assign n35186 = ~n35159 & ~n35185 ;
  assign n35188 = n25881 & ~n35186 ;
  assign n35189 = ~n35187 & n35188 ;
  assign n35145 = ~n25817 & n31320 ;
  assign n35152 = ~n25743 & ~n31452 ;
  assign n35153 = n31467 & ~n35152 ;
  assign n35154 = \P1_P2_InstAddrPointer_reg[28]/NET0131  & ~n35153 ;
  assign n35155 = ~n25763 & n25771 ;
  assign n35156 = ~n25808 & ~n35155 ;
  assign n35157 = n35148 & ~n35156 ;
  assign n35149 = n25773 & ~n35148 ;
  assign n35146 = ~\P1_P2_InstAddrPointer_reg[28]/NET0131  & ~n25773 ;
  assign n35150 = ~n25826 & ~n35146 ;
  assign n35151 = ~n35149 & n35150 ;
  assign n35160 = n25887 & n35159 ;
  assign n35190 = ~n35151 & ~n35160 ;
  assign n35191 = ~n35157 & n35190 ;
  assign n35192 = ~n35154 & n35191 ;
  assign n35193 = ~n35145 & n35192 ;
  assign n35194 = ~n35189 & n35193 ;
  assign n35195 = ~n35172 & n35194 ;
  assign n35196 = n25918 & ~n35195 ;
  assign n35143 = \P1_P2_rEIP_reg[28]/NET0131  & n27967 ;
  assign n35144 = \P1_P2_InstAddrPointer_reg[28]/NET0131  & ~n31487 ;
  assign n35197 = ~n35143 & ~n35144 ;
  assign n35198 = ~n35196 & n35197 ;
  assign n35199 = \P1_P2_InstAddrPointer_reg[29]/NET0131  & n25733 ;
  assign n35217 = n31313 & ~n35163 ;
  assign n35218 = ~n30809 & ~n31326 ;
  assign n35219 = ~n35217 & n35218 ;
  assign n35200 = ~\P1_P2_InstAddrPointer_reg[11]/NET0131  & ~n31118 ;
  assign n35201 = ~n30848 & ~n35200 ;
  assign n35202 = \P1_P2_InstAddrPointer_reg[10]/NET0131  & \P1_P2_InstAddrPointer_reg[12]/NET0131  ;
  assign n35203 = n35201 & n35202 ;
  assign n35204 = n31115 & n35203 ;
  assign n35205 = \P1_P2_InstAddrPointer_reg[13]/NET0131  & n35204 ;
  assign n35206 = \P1_P2_InstAddrPointer_reg[15]/NET0131  & n31125 ;
  assign n35207 = n35205 & n35206 ;
  assign n35208 = n31141 & n35207 ;
  assign n35209 = n30852 & n35208 ;
  assign n35210 = n31151 & n35209 ;
  assign n35211 = n31154 & n35210 ;
  assign n35212 = n31167 & n35211 ;
  assign n35214 = ~n30843 & n35212 ;
  assign n35213 = n30843 & ~n35212 ;
  assign n35215 = n30809 & ~n35213 ;
  assign n35216 = ~n35214 & n35215 ;
  assign n35220 = ~n25733 & ~n35216 ;
  assign n35221 = ~n35219 & n35220 ;
  assign n35222 = ~n35199 & ~n35221 ;
  assign n35223 = n25701 & ~n35222 ;
  assign n35225 = ~n31451 & ~n31455 ;
  assign n35226 = n25881 & ~n31456 ;
  assign n35227 = ~n35225 & n35226 ;
  assign n35224 = ~n25817 & n31313 ;
  assign n35234 = ~n25830 & n30843 ;
  assign n35230 = ~n25752 & ~n25772 ;
  assign n35228 = ~n25415 & ~n30843 ;
  assign n35229 = n25846 & ~n35228 ;
  assign n35231 = n31466 & ~n35229 ;
  assign n35232 = n35230 & n35231 ;
  assign n35233 = \P1_P2_InstAddrPointer_reg[29]/NET0131  & ~n35232 ;
  assign n35236 = n25747 & ~n31455 ;
  assign n35235 = ~\P1_P2_InstAddrPointer_reg[29]/NET0131  & ~n25747 ;
  assign n35237 = ~n25743 & ~n35235 ;
  assign n35238 = ~n35236 & n35237 ;
  assign n35239 = ~n35233 & ~n35238 ;
  assign n35240 = ~n35234 & n35239 ;
  assign n35241 = ~n35224 & n35240 ;
  assign n35242 = ~n35227 & n35241 ;
  assign n35243 = ~n35223 & n35242 ;
  assign n35244 = n25918 & ~n35243 ;
  assign n35245 = \P1_P2_InstAddrPointer_reg[29]/NET0131  & ~n31487 ;
  assign n35246 = \P1_P2_rEIP_reg[29]/NET0131  & n27967 ;
  assign n35247 = ~n35245 & ~n35246 ;
  assign n35248 = ~n35244 & n35247 ;
  assign n35251 = \P2_P1_InstAddrPointer_reg[23]/NET0131  & n25947 ;
  assign n35256 = ~n31849 & ~n31851 ;
  assign n35257 = ~n31852 & ~n35256 ;
  assign n35258 = n29503 & ~n35257 ;
  assign n35252 = n31885 & n31983 ;
  assign n35253 = n31882 & ~n35252 ;
  assign n35254 = ~n29503 & ~n31985 ;
  assign n35255 = ~n35253 & n35254 ;
  assign n35259 = ~n25947 & ~n35255 ;
  assign n35260 = ~n35258 & n35259 ;
  assign n35261 = ~n35251 & ~n35260 ;
  assign n35262 = n25945 & ~n35261 ;
  assign n35263 = n32130 & ~n32133 ;
  assign n35265 = ~n32139 & ~n35263 ;
  assign n35264 = n32139 & n35263 ;
  assign n35266 = n25964 & ~n35264 ;
  assign n35267 = ~n35265 & n35266 ;
  assign n35270 = \P2_P1_InstAddrPointer_reg[23]/NET0131  & ~n32028 ;
  assign n35269 = ~n25995 & n31882 ;
  assign n35250 = n31851 & ~n32159 ;
  assign n35268 = n26068 & n32139 ;
  assign n35271 = ~n35250 & ~n35268 ;
  assign n35272 = ~n35269 & n35271 ;
  assign n35273 = ~n35270 & n35272 ;
  assign n35274 = ~n35267 & n35273 ;
  assign n35275 = ~n35262 & n35274 ;
  assign n35276 = n11623 & ~n35275 ;
  assign n35249 = \P2_P1_rEIP_reg[23]/NET0131  & n11616 ;
  assign n35277 = \P2_P1_InstAddrPointer_reg[23]/NET0131  & ~n32172 ;
  assign n35278 = ~n35249 & ~n35277 ;
  assign n35279 = ~n35276 & n35278 ;
  assign n35281 = \P2_P1_InstAddrPointer_reg[27]/NET0131  & n25947 ;
  assign n35285 = ~n31857 & ~n31859 ;
  assign n35286 = n31857 & n31859 ;
  assign n35287 = ~n35285 & ~n35286 ;
  assign n35288 = n29503 & ~n35287 ;
  assign n35282 = ~n31997 & n32000 ;
  assign n35283 = ~n29503 & ~n32001 ;
  assign n35284 = ~n35282 & n35283 ;
  assign n35289 = ~n25947 & ~n35284 ;
  assign n35290 = ~n35288 & n35289 ;
  assign n35291 = ~n35281 & ~n35290 ;
  assign n35292 = n25945 & ~n35291 ;
  assign n35293 = ~\P2_P1_InstAddrPointer_reg[27]/NET0131  & ~n32038 ;
  assign n35294 = ~n32039 & ~n35293 ;
  assign n35295 = ~n32144 & ~n35294 ;
  assign n35296 = n25964 & ~n32145 ;
  assign n35297 = ~n35295 & n35296 ;
  assign n35300 = \P2_P1_InstAddrPointer_reg[27]/NET0131  & ~n32028 ;
  assign n35299 = ~n25995 & n32000 ;
  assign n35280 = n31859 & ~n32159 ;
  assign n35298 = n26068 & n35294 ;
  assign n35301 = ~n35280 & ~n35298 ;
  assign n35302 = ~n35299 & n35301 ;
  assign n35303 = ~n35300 & n35302 ;
  assign n35304 = ~n35297 & n35303 ;
  assign n35305 = ~n35292 & n35304 ;
  assign n35306 = n11623 & ~n35305 ;
  assign n35307 = \P2_P1_rEIP_reg[27]/NET0131  & n11616 ;
  assign n35308 = \P2_P1_InstAddrPointer_reg[27]/NET0131  & ~n32172 ;
  assign n35309 = ~n35307 & ~n35308 ;
  assign n35310 = ~n35306 & n35309 ;
  assign n35311 = \P2_P1_InstAddrPointer_reg[28]/NET0131  & n25947 ;
  assign n35315 = ~\P2_P1_InstAddrPointer_reg[28]/NET0131  & ~n31518 ;
  assign n35316 = ~n31519 & ~n35315 ;
  assign n35317 = ~n35286 & ~n35316 ;
  assign n35318 = \P2_P1_InstAddrPointer_reg[28]/NET0131  & n35286 ;
  assign n35319 = ~n35317 & ~n35318 ;
  assign n35320 = n29503 & ~n35319 ;
  assign n35312 = ~n32001 & n32004 ;
  assign n35313 = ~n29503 & ~n32005 ;
  assign n35314 = ~n35312 & n35313 ;
  assign n35321 = ~n25947 & ~n35314 ;
  assign n35322 = ~n35320 & n35321 ;
  assign n35323 = ~n35311 & ~n35322 ;
  assign n35324 = n25945 & ~n35323 ;
  assign n35326 = ~n32042 & ~n32145 ;
  assign n35327 = n25964 & ~n32146 ;
  assign n35328 = ~n35326 & n35327 ;
  assign n35332 = ~n25987 & ~n32040 ;
  assign n35333 = n32028 & ~n35332 ;
  assign n35334 = \P2_P1_InstAddrPointer_reg[28]/NET0131  & ~n35333 ;
  assign n35335 = n26068 & n32042 ;
  assign n35325 = ~n25995 & n32004 ;
  assign n35329 = ~n26031 & ~n31518 ;
  assign n35330 = n32159 & ~n35329 ;
  assign n35331 = n35316 & ~n35330 ;
  assign n35336 = ~n35325 & ~n35331 ;
  assign n35337 = ~n35335 & n35336 ;
  assign n35338 = ~n35334 & n35337 ;
  assign n35339 = ~n35328 & n35338 ;
  assign n35340 = ~n35324 & n35339 ;
  assign n35341 = n11623 & ~n35340 ;
  assign n35342 = \P2_P1_rEIP_reg[28]/NET0131  & n11616 ;
  assign n35343 = \P2_P1_InstAddrPointer_reg[28]/NET0131  & ~n32172 ;
  assign n35344 = ~n35342 & ~n35343 ;
  assign n35345 = ~n35341 & n35344 ;
  assign n35346 = \P2_P1_InstAddrPointer_reg[29]/NET0131  & n25947 ;
  assign n35347 = ~\P2_P1_InstAddrPointer_reg[29]/NET0131  & ~n31519 ;
  assign n35348 = ~n31520 & ~n35347 ;
  assign n35349 = ~n35318 & ~n35348 ;
  assign n35350 = ~n31862 & ~n35349 ;
  assign n35351 = n29503 & ~n35350 ;
  assign n35352 = ~n32005 & n32008 ;
  assign n35353 = ~n29503 & ~n32009 ;
  assign n35354 = ~n35352 & n35353 ;
  assign n35355 = ~n25947 & ~n35354 ;
  assign n35356 = ~n35351 & n35355 ;
  assign n35357 = ~n35346 & ~n35356 ;
  assign n35358 = n25945 & ~n35357 ;
  assign n35360 = ~\P2_P1_InstAddrPointer_reg[29]/NET0131  & ~n32040 ;
  assign n35361 = ~n32150 & ~n35360 ;
  assign n35364 = ~\P2_P1_InstAddrPointer_reg[10]/NET0131  & ~n32049 ;
  assign n35365 = ~n32050 & ~n35364 ;
  assign n35366 = n31537 & n35365 ;
  assign n35367 = n32102 & n35366 ;
  assign n35368 = n32054 & n35367 ;
  assign n35369 = n32111 & n35368 ;
  assign n35370 = n32116 & n35369 ;
  assign n35371 = n32126 & n35370 ;
  assign n35372 = n32129 & n35371 ;
  assign n35373 = n32141 & n35372 ;
  assign n35374 = n32044 & n35373 ;
  assign n35362 = ~\P2_P1_InstAddrPointer_reg[26]/NET0131  & ~n32037 ;
  assign n35363 = ~n32038 & ~n35362 ;
  assign n35375 = \P2_P1_InstAddrPointer_reg[28]/NET0131  & n35363 ;
  assign n35376 = n35294 & n35375 ;
  assign n35377 = n35374 & n35376 ;
  assign n35379 = n35361 & n35377 ;
  assign n35378 = ~n35361 & ~n35377 ;
  assign n35380 = n25964 & ~n35378 ;
  assign n35381 = ~n35379 & n35380 ;
  assign n35388 = n26068 & n35361 ;
  assign n35383 = ~n24711 & ~n26054 ;
  assign n35382 = ~n25952 & ~n26057 ;
  assign n35384 = ~n26053 & ~n35382 ;
  assign n35385 = n35383 & n35384 ;
  assign n35386 = ~n35332 & n35385 ;
  assign n35387 = \P2_P1_InstAddrPointer_reg[29]/NET0131  & ~n35386 ;
  assign n35359 = ~n25995 & n32008 ;
  assign n35389 = ~n32159 & n35348 ;
  assign n35390 = ~n35359 & ~n35389 ;
  assign n35391 = ~n35387 & n35390 ;
  assign n35392 = ~n35388 & n35391 ;
  assign n35393 = ~n35381 & n35392 ;
  assign n35394 = ~n35358 & n35393 ;
  assign n35395 = n11623 & ~n35394 ;
  assign n35396 = \P2_P1_InstAddrPointer_reg[29]/NET0131  & ~n32172 ;
  assign n35397 = \P2_P1_rEIP_reg[29]/NET0131  & n11616 ;
  assign n35398 = ~n35396 & ~n35397 ;
  assign n35399 = ~n35395 & n35398 ;
  assign n35402 = \P2_P2_InstAddrPointer_reg[23]/NET0131  & n26629 ;
  assign n35403 = n32533 & ~n32541 ;
  assign n35404 = ~n32543 & ~n35403 ;
  assign n35405 = ~n32541 & n34288 ;
  assign n35406 = n32543 & n35405 ;
  assign n35407 = ~n35404 & ~n35406 ;
  assign n35408 = n32510 & ~n35407 ;
  assign n35409 = n32677 & ~n32689 ;
  assign n35410 = n32687 & n35409 ;
  assign n35411 = n32680 & n35410 ;
  assign n35412 = n32684 & ~n35411 ;
  assign n35413 = ~n32510 & ~n32693 ;
  assign n35414 = ~n35412 & n35413 ;
  assign n35415 = ~n26629 & ~n35414 ;
  assign n35416 = ~n35408 & n35415 ;
  assign n35417 = ~n35402 & ~n35416 ;
  assign n35418 = n26621 & ~n35417 ;
  assign n35419 = ~n32751 & ~n32829 ;
  assign n35420 = n26744 & ~n32830 ;
  assign n35421 = ~n35419 & n35420 ;
  assign n35426 = ~n26688 & n32684 ;
  assign n35423 = ~n26619 & ~n26642 ;
  assign n35424 = n26766 & n35423 ;
  assign n35425 = \P2_P2_InstAddrPointer_reg[23]/NET0131  & ~n35424 ;
  assign n35401 = ~n26764 & n32543 ;
  assign n35422 = n26757 & n32751 ;
  assign n35427 = ~n35401 & ~n35422 ;
  assign n35428 = ~n35425 & n35427 ;
  assign n35429 = ~n35426 & n35428 ;
  assign n35430 = ~n35421 & n35429 ;
  assign n35431 = ~n35418 & n35430 ;
  assign n35432 = n26792 & ~n35431 ;
  assign n35400 = \P2_P2_rEIP_reg[23]/NET0131  & n28046 ;
  assign n35433 = \P2_P2_InstAddrPointer_reg[23]/NET0131  & ~n32860 ;
  assign n35434 = ~n35400 & ~n35433 ;
  assign n35435 = ~n35432 & n35434 ;
  assign n35464 = ~\P2_P2_InstAddrPointer_reg[27]/NET0131  & ~n32730 ;
  assign n35465 = ~n32840 & ~n35464 ;
  assign n35467 = ~n32838 & ~n35465 ;
  assign n35468 = n26744 & ~n32839 ;
  assign n35469 = ~n35467 & n35468 ;
  assign n35438 = \P2_P2_InstAddrPointer_reg[27]/NET0131  & n26629 ;
  assign n35442 = ~n32210 & ~n32550 ;
  assign n35443 = ~n32551 & ~n35442 ;
  assign n35444 = n32510 & ~n35443 ;
  assign n35439 = ~n32698 & n32701 ;
  assign n35440 = ~n32510 & ~n32702 ;
  assign n35441 = ~n35439 & n35440 ;
  assign n35445 = ~n26629 & ~n35441 ;
  assign n35446 = ~n35444 & n35445 ;
  assign n35447 = ~n35438 & ~n35446 ;
  assign n35448 = n26621 & ~n35447 ;
  assign n35462 = ~n26688 & n32701 ;
  assign n35449 = ~n26619 & ~n26728 ;
  assign n35450 = ~n26583 & ~n32840 ;
  assign n35451 = n26766 & ~n35450 ;
  assign n35452 = n35449 & n35451 ;
  assign n35453 = \P2_P2_InstAddrPointer_reg[27]/NET0131  & ~n35452 ;
  assign n35455 = ~n26286 & ~n32210 ;
  assign n35454 = ~\P2_P2_InstAddrPointer_reg[27]/NET0131  & n26286 ;
  assign n35456 = ~n26639 & ~n35454 ;
  assign n35457 = ~n35455 & n35456 ;
  assign n35458 = ~n26645 & n26651 ;
  assign n35459 = n32210 & n35458 ;
  assign n35460 = ~n35457 & ~n35459 ;
  assign n35461 = ~n26640 & ~n35460 ;
  assign n35463 = n26678 & n32210 ;
  assign n35466 = n26757 & n35465 ;
  assign n35470 = ~n35463 & ~n35466 ;
  assign n35471 = ~n35461 & n35470 ;
  assign n35472 = ~n35453 & n35471 ;
  assign n35473 = ~n35462 & n35472 ;
  assign n35474 = ~n35448 & n35473 ;
  assign n35475 = ~n35469 & n35474 ;
  assign n35476 = n26792 & ~n35475 ;
  assign n35436 = \P2_P2_rEIP_reg[27]/NET0131  & n28046 ;
  assign n35437 = \P2_P2_InstAddrPointer_reg[27]/NET0131  & ~n32860 ;
  assign n35477 = ~n35436 & ~n35437 ;
  assign n35478 = ~n35476 & n35477 ;
  assign n35482 = \P2_P2_InstAddrPointer_reg[28]/NET0131  & n26629 ;
  assign n35483 = ~n32702 & n32704 ;
  assign n35484 = ~n32705 & ~n35483 ;
  assign n35485 = ~n32510 & ~n35484 ;
  assign n35479 = ~\P2_P2_InstAddrPointer_reg[28]/NET0131  & ~n32203 ;
  assign n35480 = ~n32204 & ~n35479 ;
  assign n35487 = ~n34292 & ~n35480 ;
  assign n35486 = \P2_P2_InstAddrPointer_reg[28]/NET0131  & n34292 ;
  assign n35488 = n32510 & ~n35486 ;
  assign n35489 = ~n35487 & n35488 ;
  assign n35490 = ~n35485 & ~n35489 ;
  assign n35491 = ~n26629 & ~n35490 ;
  assign n35492 = ~n35482 & ~n35491 ;
  assign n35493 = n26621 & ~n35492 ;
  assign n35495 = ~n32839 & ~n32842 ;
  assign n35494 = \P2_P2_InstAddrPointer_reg[28]/NET0131  & n32839 ;
  assign n35496 = n26744 & ~n35494 ;
  assign n35497 = ~n35495 & n35496 ;
  assign n35501 = ~n26688 & n32704 ;
  assign n35498 = n35424 & ~n35450 ;
  assign n35499 = \P2_P2_InstAddrPointer_reg[28]/NET0131  & ~n35498 ;
  assign n35481 = ~n26764 & n35480 ;
  assign n35500 = n26757 & n32842 ;
  assign n35502 = ~n35481 & ~n35500 ;
  assign n35503 = ~n35499 & n35502 ;
  assign n35504 = ~n35501 & n35503 ;
  assign n35505 = ~n35497 & n35504 ;
  assign n35506 = ~n35493 & n35505 ;
  assign n35507 = n26792 & ~n35506 ;
  assign n35508 = \P2_P2_rEIP_reg[28]/NET0131  & n28046 ;
  assign n35509 = \P2_P2_InstAddrPointer_reg[28]/NET0131  & ~n32860 ;
  assign n35510 = ~n35508 & ~n35509 ;
  assign n35511 = ~n35507 & n35510 ;
  assign n35518 = ~\P2_P2_InstAddrPointer_reg[29]/NET0131  & ~n32731 ;
  assign n35519 = ~n32732 & ~n35518 ;
  assign n35534 = ~n35494 & ~n35519 ;
  assign n35535 = n26744 & ~n32844 ;
  assign n35536 = ~n35534 & n35535 ;
  assign n35522 = \P2_P2_InstAddrPointer_reg[29]/NET0131  & n26629 ;
  assign n35526 = \P2_P2_InstAddrPointer_reg[28]/NET0131  & n32551 ;
  assign n35527 = ~n32207 & ~n35526 ;
  assign n35528 = ~n32552 & ~n35527 ;
  assign n35529 = n32510 & ~n35528 ;
  assign n35523 = ~n32705 & n32707 ;
  assign n35524 = ~n32510 & ~n32708 ;
  assign n35525 = ~n35523 & n35524 ;
  assign n35530 = ~n26629 & ~n35525 ;
  assign n35531 = ~n35529 & n35530 ;
  assign n35532 = ~n35522 & ~n35531 ;
  assign n35533 = n26621 & ~n35532 ;
  assign n35515 = ~n26583 & ~n32731 ;
  assign n35516 = n34267 & ~n35515 ;
  assign n35517 = \P2_P2_InstAddrPointer_reg[29]/NET0131  & ~n35516 ;
  assign n35514 = ~n26688 & n32707 ;
  assign n35520 = n26757 & n35519 ;
  assign n35521 = ~n26764 & n32207 ;
  assign n35537 = ~n35520 & ~n35521 ;
  assign n35538 = ~n35514 & n35537 ;
  assign n35539 = ~n35517 & n35538 ;
  assign n35540 = ~n35533 & n35539 ;
  assign n35541 = ~n35536 & n35540 ;
  assign n35542 = n26792 & ~n35541 ;
  assign n35512 = \P2_P2_InstAddrPointer_reg[29]/NET0131  & ~n32860 ;
  assign n35513 = \P2_P2_rEIP_reg[29]/NET0131  & n28046 ;
  assign n35543 = ~n35512 & ~n35513 ;
  assign n35544 = ~n35542 & n35543 ;
  assign n35547 = n32892 & n32923 ;
  assign n35548 = ~\P2_P3_InstAddrPointer_reg[23]/NET0131  & ~n35547 ;
  assign n35549 = n32893 & n32923 ;
  assign n35550 = ~n35548 & ~n35549 ;
  assign n35551 = \P2_P3_InstAddrPointer_reg[21]/NET0131  & n33263 ;
  assign n35552 = \P2_P3_InstAddrPointer_reg[22]/NET0131  & n35551 ;
  assign n35553 = ~n35550 & ~n35552 ;
  assign n35554 = ~\P2_P3_InstAddrPointer_reg[12]/NET0131  & ~n32917 ;
  assign n35555 = ~n32918 & ~n35554 ;
  assign n35556 = n32884 & n35555 ;
  assign n35557 = n32952 & n35556 ;
  assign n35558 = n33252 & n35557 ;
  assign n35559 = n33259 & n35558 ;
  assign n35560 = n33262 & n35559 ;
  assign n35561 = n32893 & n35560 ;
  assign n35562 = ~n35553 & ~n35561 ;
  assign n35563 = n33242 & ~n35562 ;
  assign n35564 = n33279 & ~n33384 ;
  assign n35565 = ~n33242 & ~n33385 ;
  assign n35566 = ~n35564 & n35565 ;
  assign n35567 = ~n35563 & ~n35566 ;
  assign n35568 = n27283 & ~n35567 ;
  assign n35546 = ~\P2_P3_InstAddrPointer_reg[23]/NET0131  & ~n27283 ;
  assign n35569 = n27117 & ~n35546 ;
  assign n35570 = ~n35568 & n35569 ;
  assign n35574 = ~\P2_P3_InstAddrPointer_reg[22]/NET0131  & ~n33418 ;
  assign n35575 = ~n33419 & ~n35574 ;
  assign n35576 = n33490 & n35575 ;
  assign n35577 = ~n33421 & ~n35576 ;
  assign n35578 = n27280 & ~n33491 ;
  assign n35579 = ~n35577 & n35578 ;
  assign n35587 = ~\P2_P3_InstAddrPointer_reg[23]/NET0131  & ~n27206 ;
  assign n35588 = ~n27111 & ~n35587 ;
  assign n35589 = n33421 & n35588 ;
  assign n35580 = ~n27142 & n33279 ;
  assign n35571 = \P2_P3_InstAddrPointer_reg[23]/NET0131  & ~n27180 ;
  assign n35572 = n27229 & ~n35571 ;
  assign n35573 = n35550 & ~n35572 ;
  assign n35581 = ~n27181 & n27295 ;
  assign n35582 = ~n27253 & n35581 ;
  assign n35583 = n27180 & ~n27256 ;
  assign n35584 = n27192 & ~n35583 ;
  assign n35585 = n35582 & ~n35584 ;
  assign n35586 = \P2_P3_InstAddrPointer_reg[23]/NET0131  & ~n35585 ;
  assign n35590 = ~n35573 & ~n35586 ;
  assign n35591 = ~n35580 & n35590 ;
  assign n35592 = ~n35589 & n35591 ;
  assign n35593 = ~n35579 & n35592 ;
  assign n35594 = ~n35570 & n35593 ;
  assign n35595 = n27308 & ~n35594 ;
  assign n35545 = \P2_P3_rEIP_reg[23]/NET0131  & n32864 ;
  assign n35596 = \P2_P3_InstAddrPointer_reg[23]/NET0131  & ~n32870 ;
  assign n35597 = ~n35545 & ~n35596 ;
  assign n35598 = ~n35595 & n35597 ;
  assign n35604 = \P2_P3_InstAddrPointer_reg[27]/NET0131  & ~n27283 ;
  assign n35608 = \P2_P3_InstAddrPointer_reg[26]/NET0131  & n32925 ;
  assign n35609 = ~\P2_P3_InstAddrPointer_reg[27]/NET0131  & ~n35608 ;
  assign n35610 = ~n32926 & ~n35609 ;
  assign n35611 = n32949 & n33264 ;
  assign n35612 = \P2_P3_InstAddrPointer_reg[26]/NET0131  & n35611 ;
  assign n35613 = ~n35610 & ~n35612 ;
  assign n35614 = ~n33265 & ~n35613 ;
  assign n35615 = n33242 & ~n35614 ;
  assign n35605 = ~n33397 & n33400 ;
  assign n35606 = ~n33242 & ~n33401 ;
  assign n35607 = ~n35605 & n35606 ;
  assign n35616 = n27283 & ~n35607 ;
  assign n35617 = ~n35615 & n35616 ;
  assign n35618 = ~n35604 & ~n35617 ;
  assign n35619 = n27117 & ~n35618 ;
  assign n35601 = ~\P2_P3_InstAddrPointer_reg[27]/NET0131  & ~n32897 ;
  assign n35602 = ~n32898 & ~n35601 ;
  assign n35620 = n33492 & n33494 ;
  assign n35621 = \P2_P3_InstAddrPointer_reg[26]/NET0131  & n35620 ;
  assign n35622 = ~n35602 & ~n35621 ;
  assign n35623 = n27280 & ~n33496 ;
  assign n35624 = ~n35622 & n35623 ;
  assign n35603 = n27219 & n35602 ;
  assign n35625 = ~n27142 & n33400 ;
  assign n35626 = ~n27229 & n35610 ;
  assign n35627 = \P2_P3_InstAddrPointer_reg[27]/NET0131  & ~n34355 ;
  assign n35628 = ~n35626 & ~n35627 ;
  assign n35629 = ~n35625 & n35628 ;
  assign n35630 = ~n35603 & n35629 ;
  assign n35631 = ~n35624 & n35630 ;
  assign n35632 = ~n35619 & n35631 ;
  assign n35633 = n27308 & ~n35632 ;
  assign n35599 = \P2_P3_rEIP_reg[27]/NET0131  & n32864 ;
  assign n35600 = \P2_P3_InstAddrPointer_reg[27]/NET0131  & ~n32870 ;
  assign n35634 = ~n35599 & ~n35600 ;
  assign n35635 = ~n35633 & n35634 ;
  assign n35638 = n33404 & ~n34338 ;
  assign n35639 = ~n33242 & ~n34339 ;
  assign n35640 = ~n35638 & n35639 ;
  assign n35641 = ~\P2_P3_InstAddrPointer_reg[24]/NET0131  & ~n35549 ;
  assign n35642 = ~n32924 & ~n35641 ;
  assign n35643 = n35561 & n35642 ;
  assign n35644 = n32950 & n35643 ;
  assign n35646 = ~n33267 & n35644 ;
  assign n35645 = n33267 & ~n35644 ;
  assign n35647 = n33242 & ~n35645 ;
  assign n35648 = ~n35646 & n35647 ;
  assign n35649 = ~n35640 & ~n35648 ;
  assign n35650 = n27283 & ~n35649 ;
  assign n35637 = ~\P2_P3_InstAddrPointer_reg[28]/NET0131  & ~n27283 ;
  assign n35651 = n27117 & ~n35637 ;
  assign n35652 = ~n35650 & n35651 ;
  assign n35653 = ~\P2_P3_InstAddrPointer_reg[24]/NET0131  & ~n32894 ;
  assign n35654 = ~n32895 & ~n35653 ;
  assign n35657 = \P2_P3_InstAddrPointer_reg[15]/NET0131  & n33481 ;
  assign n35658 = ~\P2_P3_InstAddrPointer_reg[16]/NET0131  & ~n32886 ;
  assign n35659 = ~n32887 & ~n35658 ;
  assign n35660 = n35657 & n35659 ;
  assign n35661 = n33487 & n35660 ;
  assign n35662 = n33424 & n35661 ;
  assign n35655 = ~\P2_P3_InstAddrPointer_reg[21]/NET0131  & ~n32891 ;
  assign n35656 = ~n33418 & ~n35655 ;
  assign n35663 = n33422 & n35656 ;
  assign n35664 = n35662 & n35663 ;
  assign n35665 = n35654 & n35664 ;
  assign n35666 = n33495 & n35665 ;
  assign n35668 = ~n33498 & ~n35666 ;
  assign n35667 = n33498 & n35666 ;
  assign n35669 = n27280 & ~n35667 ;
  assign n35670 = ~n35668 & n35669 ;
  assign n35671 = n27219 & n33498 ;
  assign n35636 = ~n27142 & n33404 ;
  assign n35672 = ~n32941 & n35582 ;
  assign n35673 = \P2_P3_InstAddrPointer_reg[28]/NET0131  & ~n35672 ;
  assign n35674 = ~n27229 & n33267 ;
  assign n35675 = ~n35673 & ~n35674 ;
  assign n35676 = ~n35636 & n35675 ;
  assign n35677 = ~n35671 & n35676 ;
  assign n35678 = ~n35670 & n35677 ;
  assign n35679 = ~n35652 & n35678 ;
  assign n35680 = n27308 & ~n35679 ;
  assign n35681 = \P2_P3_InstAddrPointer_reg[28]/NET0131  & ~n32870 ;
  assign n35682 = \P2_P3_rEIP_reg[28]/NET0131  & n32864 ;
  assign n35683 = ~n35681 & ~n35682 ;
  assign n35684 = ~n35680 & n35683 ;
  assign n35686 = \P2_P3_InstAddrPointer_reg[29]/NET0131  & ~n27283 ;
  assign n35690 = ~\P2_P3_InstAddrPointer_reg[29]/NET0131  & ~n32927 ;
  assign n35691 = ~n32928 & ~n35690 ;
  assign n35692 = ~n33268 & ~n35691 ;
  assign n35693 = ~n33269 & ~n35692 ;
  assign n35694 = n33242 & ~n35693 ;
  assign n35687 = ~n33405 & n33407 ;
  assign n35688 = ~n33242 & ~n33408 ;
  assign n35689 = ~n35687 & n35688 ;
  assign n35695 = n27283 & ~n35689 ;
  assign n35696 = ~n35694 & n35695 ;
  assign n35697 = ~n35686 & ~n35696 ;
  assign n35698 = n27117 & ~n35697 ;
  assign n35699 = ~\P2_P3_InstAddrPointer_reg[29]/NET0131  & ~n32899 ;
  assign n35700 = ~n32900 & ~n35699 ;
  assign n35701 = ~n33499 & ~n35700 ;
  assign n35702 = n27280 & ~n33500 ;
  assign n35703 = ~n35701 & n35702 ;
  assign n35706 = n27219 & n35700 ;
  assign n35704 = ~n27142 & n33407 ;
  assign n35685 = \P2_P3_InstAddrPointer_reg[29]/NET0131  & ~n35672 ;
  assign n35705 = ~n27229 & n35691 ;
  assign n35707 = ~n35685 & ~n35705 ;
  assign n35708 = ~n35704 & n35707 ;
  assign n35709 = ~n35706 & n35708 ;
  assign n35710 = ~n35703 & n35709 ;
  assign n35711 = ~n35698 & n35710 ;
  assign n35712 = n27308 & ~n35711 ;
  assign n35713 = \P2_P3_rEIP_reg[29]/NET0131  & n32864 ;
  assign n35714 = \P2_P3_InstAddrPointer_reg[29]/NET0131  & ~n32870 ;
  assign n35715 = ~n35713 & ~n35714 ;
  assign n35716 = ~n35712 & n35715 ;
  assign n35719 = \P1_P1_InstAddrPointer_reg[23]/NET0131  & n26249 ;
  assign n35724 = n33516 & n33830 ;
  assign n35725 = ~n33851 & ~n35724 ;
  assign n35726 = ~\P1_P1_InstAddrPointer_reg[16]/NET0131  & ~n33532 ;
  assign n35727 = ~n33533 & ~n35726 ;
  assign n35730 = \P1_P1_InstAddrPointer_reg[11]/NET0131  & n33817 ;
  assign n35728 = ~\P1_P1_InstAddrPointer_reg[12]/NET0131  & ~n33946 ;
  assign n35729 = ~n33530 & ~n35728 ;
  assign n35731 = n33519 & n33549 ;
  assign n35732 = n35729 & n35731 ;
  assign n35733 = n35730 & n35732 ;
  assign n35734 = n35727 & n35733 ;
  assign n35735 = n33826 & n35734 ;
  assign n35736 = n33829 & n35735 ;
  assign n35737 = n33853 & n35736 ;
  assign n35738 = ~n35725 & ~n35737 ;
  assign n35739 = n29558 & ~n35738 ;
  assign n35720 = ~n33873 & n33979 ;
  assign n35721 = ~n33876 & ~n35720 ;
  assign n35722 = ~n29558 & ~n33981 ;
  assign n35723 = ~n35721 & n35722 ;
  assign n35740 = ~n26249 & ~n35723 ;
  assign n35741 = ~n35739 & n35740 ;
  assign n35742 = ~n35719 & ~n35741 ;
  assign n35743 = n26126 & ~n35742 ;
  assign n35744 = ~n34114 & ~n34117 ;
  assign n35745 = n26263 & ~n34118 ;
  assign n35746 = ~n35744 & n35745 ;
  assign n35749 = ~n26151 & ~n33876 ;
  assign n35748 = n26192 & n34117 ;
  assign n35718 = \P1_P1_InstAddrPointer_reg[23]/NET0131  & ~n34390 ;
  assign n35747 = ~n26189 & n33851 ;
  assign n35750 = ~n35718 & ~n35747 ;
  assign n35751 = ~n35748 & n35750 ;
  assign n35752 = ~n35749 & n35751 ;
  assign n35753 = ~n35746 & n35752 ;
  assign n35754 = ~n35743 & n35753 ;
  assign n35755 = n8355 & ~n35754 ;
  assign n35717 = \P1_P1_InstAddrPointer_reg[23]/NET0131  & ~n34164 ;
  assign n35756 = \P1_P1_rEIP_reg[23]/NET0131  & n8357 ;
  assign n35757 = ~n35717 & ~n35756 ;
  assign n35758 = ~n35755 & n35757 ;
  assign n35762 = \P1_P1_InstAddrPointer_reg[27]/NET0131  & n26249 ;
  assign n35767 = \P1_P1_InstAddrPointer_reg[26]/NET0131  & n33538 ;
  assign n35768 = ~\P1_P1_InstAddrPointer_reg[27]/NET0131  & ~n35767 ;
  assign n35769 = ~n33540 & ~n35768 ;
  assign n35770 = n33855 & n33857 ;
  assign n35771 = \P1_P1_InstAddrPointer_reg[26]/NET0131  & n35770 ;
  assign n35772 = ~n35769 & ~n35771 ;
  assign n35773 = ~n33859 & ~n35772 ;
  assign n35774 = n29558 & ~n35773 ;
  assign n35763 = n33990 & ~n33996 ;
  assign n35764 = n33994 & ~n35763 ;
  assign n35765 = ~n29558 & ~n33998 ;
  assign n35766 = ~n35764 & n35765 ;
  assign n35775 = ~n26249 & ~n35766 ;
  assign n35776 = ~n35774 & n35775 ;
  assign n35777 = ~n35762 & ~n35776 ;
  assign n35778 = n26126 & ~n35777 ;
  assign n35779 = ~\P1_P1_InstAddrPointer_reg[27]/NET0131  & ~n34038 ;
  assign n35780 = ~n34039 & ~n35779 ;
  assign n35781 = \P1_P1_InstAddrPointer_reg[25]/NET0131  & n34121 ;
  assign n35782 = \P1_P1_InstAddrPointer_reg[26]/NET0131  & n35781 ;
  assign n35783 = ~n35780 & ~n35782 ;
  assign n35784 = n26263 & ~n34125 ;
  assign n35785 = ~n35783 & n35784 ;
  assign n35786 = ~n26151 & n33994 ;
  assign n35788 = n26192 & n35780 ;
  assign n35760 = n26252 & n26256 ;
  assign n35761 = \P1_P1_InstAddrPointer_reg[27]/NET0131  & ~n35760 ;
  assign n35787 = ~n26189 & n35769 ;
  assign n35789 = ~n35761 & ~n35787 ;
  assign n35790 = ~n35788 & n35789 ;
  assign n35791 = ~n35786 & n35790 ;
  assign n35792 = ~n35785 & n35791 ;
  assign n35793 = ~n35778 & n35792 ;
  assign n35794 = n8355 & ~n35793 ;
  assign n35759 = \P1_P1_InstAddrPointer_reg[27]/NET0131  & ~n34164 ;
  assign n35795 = \P1_P1_rEIP_reg[27]/NET0131  & n8357 ;
  assign n35796 = ~n35759 & ~n35795 ;
  assign n35797 = ~n35794 & n35796 ;
  assign n35800 = \P1_P1_InstAddrPointer_reg[28]/NET0131  & n26249 ;
  assign n35807 = ~n33998 & n34001 ;
  assign n35808 = ~n29558 & ~n34002 ;
  assign n35809 = ~n35807 & n35808 ;
  assign n35801 = ~n33845 & n35737 ;
  assign n35802 = n33858 & n35801 ;
  assign n35804 = ~n33547 & n35802 ;
  assign n35803 = n33547 & ~n35802 ;
  assign n35805 = n29558 & ~n35803 ;
  assign n35806 = ~n35804 & n35805 ;
  assign n35810 = ~n26249 & ~n35806 ;
  assign n35811 = ~n35809 & n35810 ;
  assign n35812 = ~n35800 & ~n35811 ;
  assign n35813 = n26126 & ~n35812 ;
  assign n35816 = \P1_P1_InstAddrPointer_reg[15]/NET0131  & n34101 ;
  assign n35817 = ~\P1_P1_InstAddrPointer_reg[16]/NET0131  & ~n34032 ;
  assign n35818 = ~n34033 & ~n35817 ;
  assign n35819 = n35816 & n35818 ;
  assign n35820 = n33517 & n34106 ;
  assign n35821 = n35819 & n35820 ;
  assign n35822 = n34045 & n35821 ;
  assign n35814 = ~\P1_P1_InstAddrPointer_reg[21]/NET0131  & ~n34044 ;
  assign n35815 = ~n34111 & ~n35814 ;
  assign n35823 = \P1_P1_InstAddrPointer_reg[23]/NET0131  & n35815 ;
  assign n35824 = n34113 & n35823 ;
  assign n35825 = n35822 & n35824 ;
  assign n35826 = n34120 & n35825 ;
  assign n35827 = n34124 & n35826 ;
  assign n35829 = ~n34042 & ~n35827 ;
  assign n35828 = n34042 & n35827 ;
  assign n35830 = n26263 & ~n35828 ;
  assign n35831 = ~n35829 & n35830 ;
  assign n35841 = ~n26123 & ~n34040 ;
  assign n35843 = n26177 & ~n26199 ;
  assign n35832 = ~n24504 & n26160 ;
  assign n35842 = n15335 & ~n35832 ;
  assign n35844 = n26252 & ~n35842 ;
  assign n35845 = n35843 & n35844 ;
  assign n35846 = ~n35841 & n35845 ;
  assign n35847 = \P1_P1_InstAddrPointer_reg[28]/NET0131  & ~n35846 ;
  assign n35840 = ~n26151 & n34001 ;
  assign n35799 = n26192 & n34042 ;
  assign n35833 = ~n15335 & ~n26235 ;
  assign n35834 = ~\P1_P1_InstAddrPointer_reg[28]/NET0131  & ~n35833 ;
  assign n35835 = ~n35832 & ~n35834 ;
  assign n35836 = n15365 & n15383 ;
  assign n35837 = ~n26129 & ~n35836 ;
  assign n35838 = ~n35835 & n35837 ;
  assign n35839 = n33547 & ~n35838 ;
  assign n35848 = ~n35799 & ~n35839 ;
  assign n35849 = ~n35840 & n35848 ;
  assign n35850 = ~n35847 & n35849 ;
  assign n35851 = ~n35831 & n35850 ;
  assign n35852 = ~n35813 & n35851 ;
  assign n35853 = n8355 & ~n35852 ;
  assign n35798 = \P1_P1_rEIP_reg[28]/NET0131  & n8357 ;
  assign n35854 = \P1_P1_InstAddrPointer_reg[28]/NET0131  & ~n34164 ;
  assign n35855 = ~n35798 & ~n35854 ;
  assign n35856 = ~n35853 & n35855 ;
  assign n35861 = \P1_P1_InstAddrPointer_reg[29]/NET0131  & n26249 ;
  assign n35867 = ~n34002 & n34005 ;
  assign n35868 = ~n29558 & ~n34006 ;
  assign n35869 = ~n35867 & n35868 ;
  assign n35862 = ~\P1_P1_InstAddrPointer_reg[29]/NET0131  & ~n33541 ;
  assign n35863 = ~n33542 & ~n35862 ;
  assign n35864 = ~n33860 & ~n35863 ;
  assign n35865 = ~n33861 & ~n35864 ;
  assign n35866 = n29558 & ~n35865 ;
  assign n35870 = ~n26249 & ~n35866 ;
  assign n35871 = ~n35869 & n35870 ;
  assign n35872 = ~n35861 & ~n35871 ;
  assign n35873 = n26126 & ~n35872 ;
  assign n35858 = ~\P1_P1_InstAddrPointer_reg[29]/NET0131  & ~n34040 ;
  assign n35859 = ~n34128 & ~n35858 ;
  assign n35874 = ~n34126 & ~n35859 ;
  assign n35875 = n26263 & ~n34127 ;
  assign n35876 = ~n35874 & n35875 ;
  assign n35860 = n26192 & n35859 ;
  assign n35878 = ~n26189 & n35863 ;
  assign n35881 = ~n35860 & ~n35878 ;
  assign n35877 = ~n26151 & n34005 ;
  assign n35879 = n35760 & ~n35841 ;
  assign n35880 = \P1_P1_InstAddrPointer_reg[29]/NET0131  & ~n35879 ;
  assign n35882 = ~n35877 & ~n35880 ;
  assign n35883 = n35881 & n35882 ;
  assign n35884 = ~n35876 & n35883 ;
  assign n35885 = ~n35873 & n35884 ;
  assign n35886 = n8355 & ~n35885 ;
  assign n35857 = \P1_P1_rEIP_reg[29]/NET0131  & n8357 ;
  assign n35887 = \P1_P1_InstAddrPointer_reg[29]/NET0131  & ~n34164 ;
  assign n35888 = ~n35857 & ~n35887 ;
  assign n35889 = ~n35886 & n35888 ;
  assign n35890 = \P2_P1_EAX_reg[5]/NET0131  & ~n27438 ;
  assign n35892 = n11378 & n24708 ;
  assign n35891 = n20728 & ~n31614 ;
  assign n35893 = ~\P2_P1_EAX_reg[5]/NET0131  & ~n21026 ;
  assign n35894 = ~n21027 & ~n35893 ;
  assign n35895 = n21022 & n35894 ;
  assign n35896 = ~n35891 & ~n35895 ;
  assign n35897 = ~n35892 & n35896 ;
  assign n35898 = n11623 & ~n35897 ;
  assign n35899 = ~n35890 & ~n35898 ;
  assign n35900 = \P2_P1_EAX_reg[6]/NET0131  & ~n27438 ;
  assign n35902 = n11383 & n24708 ;
  assign n35901 = n20728 & ~n31579 ;
  assign n35903 = ~\P2_P1_EAX_reg[6]/NET0131  & ~n21027 ;
  assign n35904 = ~n21028 & ~n35903 ;
  assign n35905 = n21022 & n35904 ;
  assign n35906 = ~n35901 & ~n35905 ;
  assign n35907 = ~n35902 & n35906 ;
  assign n35908 = n11623 & ~n35907 ;
  assign n35909 = ~n35900 & ~n35908 ;
  assign n35910 = \P2_P1_uWord_reg[8]/NET0131  & ~n24913 ;
  assign n35911 = ~\P2_P1_EAX_reg[24]/NET0131  & ~n27395 ;
  assign n35912 = ~n27396 & ~n35911 ;
  assign n35913 = n24898 & n35912 ;
  assign n35914 = n21062 & n28717 ;
  assign n35915 = ~n35913 & ~n35914 ;
  assign n35916 = ~n21081 & ~n35915 ;
  assign n35917 = \P2_P1_uWord_reg[8]/NET0131  & ~n25154 ;
  assign n35918 = ~n35916 & ~n35917 ;
  assign n35919 = n11623 & ~n35918 ;
  assign n35920 = ~n35910 & ~n35919 ;
  assign n35921 = \P1_P1_EAX_reg[5]/NET0131  & ~n15326 ;
  assign n35923 = \P1_P1_EAX_reg[5]/NET0131  & ~n15365 ;
  assign n35924 = ~n24439 & ~n35923 ;
  assign n35925 = ~n15384 & ~n35924 ;
  assign n35922 = \P1_P1_EAX_reg[5]/NET0131  & ~n23190 ;
  assign n35926 = n22818 & ~n33626 ;
  assign n35927 = ~\P1_P1_EAX_reg[5]/NET0131  & ~n15391 ;
  assign n35928 = ~n15392 & ~n35927 ;
  assign n35929 = n15377 & n35928 ;
  assign n35930 = ~n35926 & ~n35929 ;
  assign n35931 = ~n35922 & n35930 ;
  assign n35932 = ~n35925 & n35931 ;
  assign n35933 = n8355 & ~n35932 ;
  assign n35934 = ~n35921 & ~n35933 ;
  assign n35935 = \P1_P1_EAX_reg[6]/NET0131  & ~n15326 ;
  assign n35937 = \P1_P1_EAX_reg[6]/NET0131  & ~n15365 ;
  assign n35938 = ~n24167 & ~n35937 ;
  assign n35939 = ~n15384 & ~n35938 ;
  assign n35936 = \P1_P1_EAX_reg[6]/NET0131  & ~n23190 ;
  assign n35940 = n22818 & ~n33591 ;
  assign n35941 = ~\P1_P1_EAX_reg[6]/NET0131  & ~n15392 ;
  assign n35942 = ~n15393 & ~n35941 ;
  assign n35943 = n15377 & n35942 ;
  assign n35944 = ~n35940 & ~n35943 ;
  assign n35945 = ~n35936 & n35944 ;
  assign n35946 = ~n35939 & n35945 ;
  assign n35947 = n8355 & ~n35946 ;
  assign n35948 = ~n35935 & ~n35947 ;
  assign n35949 = \P1_P1_uWord_reg[8]/NET0131  & ~n24515 ;
  assign n35953 = \P1_P1_uWord_reg[8]/NET0131  & n25363 ;
  assign n35954 = ~n23926 & ~n35953 ;
  assign n35955 = n15334 & ~n35954 ;
  assign n35950 = ~\P1_P1_EAX_reg[24]/NET0131  & ~n25355 ;
  assign n35951 = n24503 & ~n27424 ;
  assign n35952 = ~n35950 & n35951 ;
  assign n35956 = \P1_P1_uWord_reg[8]/NET0131  & n24505 ;
  assign n35957 = ~n35952 & ~n35956 ;
  assign n35958 = ~n35955 & n35957 ;
  assign n35959 = n8355 & ~n35958 ;
  assign n35960 = ~n35949 & ~n35959 ;
  assign n35969 = \P1_buf2_reg[26]/NET0131  & ~n27934 ;
  assign n35970 = \P1_buf1_reg[26]/NET0131  & n27934 ;
  assign n35971 = ~n35969 & ~n35970 ;
  assign n35972 = n27945 & ~n35971 ;
  assign n35973 = \P1_buf2_reg[18]/NET0131  & ~n27934 ;
  assign n35974 = \P1_buf1_reg[18]/NET0131  & n27934 ;
  assign n35975 = ~n35973 & ~n35974 ;
  assign n35976 = n27952 & ~n35975 ;
  assign n35977 = ~n35972 & ~n35976 ;
  assign n35978 = \P1_P2_DataWidth_reg[1]/NET0131  & ~n35977 ;
  assign n35961 = \P1_buf2_reg[2]/NET0131  & ~n27934 ;
  assign n35962 = \P1_buf1_reg[2]/NET0131  & n27934 ;
  assign n35963 = ~n35961 & ~n35962 ;
  assign n35964 = ~n27905 & ~n35963 ;
  assign n35965 = \P1_P2_InstQueue_reg[11][2]/NET0131  & ~n27901 ;
  assign n35966 = ~n27904 & n35965 ;
  assign n35967 = ~n35964 & ~n35966 ;
  assign n35979 = ~n27960 & ~n35967 ;
  assign n35980 = ~n35978 & ~n35979 ;
  assign n35981 = n25928 & ~n35980 ;
  assign n35982 = ~n25604 & n27901 ;
  assign n35983 = ~n35965 & ~n35982 ;
  assign n35984 = n27608 & ~n35983 ;
  assign n35968 = n27898 & ~n35967 ;
  assign n35985 = \P1_P2_InstQueue_reg[11][2]/NET0131  & ~n27972 ;
  assign n35986 = ~n35968 & ~n35985 ;
  assign n35987 = ~n35984 & n35986 ;
  assign n35988 = ~n35981 & n35987 ;
  assign n36000 = \P2_buf2_reg[26]/NET0131  & ~n28013 ;
  assign n36001 = \P2_buf1_reg[26]/NET0131  & n28013 ;
  assign n36002 = ~n36000 & ~n36001 ;
  assign n36003 = n28027 & ~n36002 ;
  assign n36004 = \P2_buf2_reg[18]/NET0131  & ~n28013 ;
  assign n36005 = \P2_buf1_reg[18]/NET0131  & n28013 ;
  assign n36006 = ~n36004 & ~n36005 ;
  assign n36007 = n28034 & ~n36006 ;
  assign n36008 = ~n36003 & ~n36007 ;
  assign n36009 = \P2_P2_DataWidth_reg[1]/NET0131  & ~n36008 ;
  assign n35989 = \P2_buf2_reg[2]/NET0131  & ~n28013 ;
  assign n35990 = \P2_buf1_reg[2]/NET0131  & n28013 ;
  assign n35991 = ~n35989 & ~n35990 ;
  assign n35992 = ~n27984 & ~n35991 ;
  assign n35993 = \P2_P2_InstQueue_reg[11][2]/NET0131  & ~n27980 ;
  assign n35994 = ~n27983 & n35993 ;
  assign n35995 = ~n35992 & ~n35994 ;
  assign n36010 = ~n28042 & ~n35995 ;
  assign n36011 = ~n36009 & ~n36010 ;
  assign n36012 = n26794 & ~n36011 ;
  assign n35997 = ~n26481 & n27980 ;
  assign n35998 = ~n35993 & ~n35997 ;
  assign n35999 = n27613 & ~n35998 ;
  assign n35996 = n27977 & ~n35995 ;
  assign n36013 = \P2_P2_InstQueue_reg[11][2]/NET0131  & ~n28050 ;
  assign n36014 = ~n35996 & ~n36013 ;
  assign n36015 = ~n35999 & n36014 ;
  assign n36016 = ~n36012 & n36015 ;
  assign n36022 = n28065 & ~n35971 ;
  assign n36023 = n28068 & ~n35975 ;
  assign n36024 = ~n36022 & ~n36023 ;
  assign n36025 = \P1_P2_DataWidth_reg[1]/NET0131  & ~n36024 ;
  assign n36017 = ~n28058 & ~n35963 ;
  assign n36018 = \P1_P2_InstQueue_reg[0][2]/NET0131  & ~n28055 ;
  assign n36019 = ~n28057 & n36018 ;
  assign n36020 = ~n36017 & ~n36019 ;
  assign n36026 = ~n28073 & ~n36020 ;
  assign n36027 = ~n36025 & ~n36026 ;
  assign n36028 = n25928 & ~n36027 ;
  assign n36029 = ~n25604 & n28055 ;
  assign n36030 = ~n36018 & ~n36029 ;
  assign n36031 = n27608 & ~n36030 ;
  assign n36021 = n27898 & ~n36020 ;
  assign n36032 = \P1_P2_InstQueue_reg[0][2]/NET0131  & ~n27972 ;
  assign n36033 = ~n36021 & ~n36032 ;
  assign n36034 = ~n36031 & n36033 ;
  assign n36035 = ~n36028 & n36034 ;
  assign n36041 = n28090 & ~n35971 ;
  assign n36042 = n27945 & ~n35975 ;
  assign n36043 = ~n36041 & ~n36042 ;
  assign n36044 = \P1_P2_DataWidth_reg[1]/NET0131  & ~n36043 ;
  assign n36036 = ~n28084 & ~n35963 ;
  assign n36037 = \P1_P2_InstQueue_reg[10][2]/NET0131  & ~n27904 ;
  assign n36038 = ~n27952 & n36037 ;
  assign n36039 = ~n36036 & ~n36038 ;
  assign n36045 = ~n28096 & ~n36039 ;
  assign n36046 = ~n36044 & ~n36045 ;
  assign n36047 = n25928 & ~n36046 ;
  assign n36048 = ~n25604 & n27904 ;
  assign n36049 = ~n36037 & ~n36048 ;
  assign n36050 = n27608 & ~n36049 ;
  assign n36040 = n27898 & ~n36039 ;
  assign n36051 = \P1_P2_InstQueue_reg[10][2]/NET0131  & ~n27972 ;
  assign n36052 = ~n36040 & ~n36051 ;
  assign n36053 = ~n36050 & n36052 ;
  assign n36054 = ~n36047 & n36053 ;
  assign n36060 = n27952 & ~n35971 ;
  assign n36061 = n27904 & ~n35975 ;
  assign n36062 = ~n36060 & ~n36061 ;
  assign n36063 = \P1_P2_DataWidth_reg[1]/NET0131  & ~n36062 ;
  assign n36055 = ~n28109 & ~n35963 ;
  assign n36056 = \P1_P2_InstQueue_reg[12][2]/NET0131  & ~n28108 ;
  assign n36057 = ~n27901 & n36056 ;
  assign n36058 = ~n36055 & ~n36057 ;
  assign n36064 = ~n28119 & ~n36058 ;
  assign n36065 = ~n36063 & ~n36064 ;
  assign n36066 = n25928 & ~n36065 ;
  assign n36067 = ~n25604 & n28108 ;
  assign n36068 = ~n36056 & ~n36067 ;
  assign n36069 = n27608 & ~n36068 ;
  assign n36059 = n27898 & ~n36058 ;
  assign n36070 = \P1_P2_InstQueue_reg[12][2]/NET0131  & ~n27972 ;
  assign n36071 = ~n36059 & ~n36070 ;
  assign n36072 = ~n36069 & n36071 ;
  assign n36073 = ~n36066 & n36072 ;
  assign n36079 = n27904 & ~n35971 ;
  assign n36080 = n27901 & ~n35975 ;
  assign n36081 = ~n36079 & ~n36080 ;
  assign n36082 = \P1_P2_DataWidth_reg[1]/NET0131  & ~n36081 ;
  assign n36074 = ~n28130 & ~n35963 ;
  assign n36075 = \P1_P2_InstQueue_reg[13][2]/NET0131  & ~n28065 ;
  assign n36076 = ~n28108 & n36075 ;
  assign n36077 = ~n36074 & ~n36076 ;
  assign n36083 = ~n28140 & ~n36077 ;
  assign n36084 = ~n36082 & ~n36083 ;
  assign n36085 = n25928 & ~n36084 ;
  assign n36086 = ~n25604 & n28065 ;
  assign n36087 = ~n36075 & ~n36086 ;
  assign n36088 = n27608 & ~n36087 ;
  assign n36078 = n27898 & ~n36077 ;
  assign n36089 = \P1_P2_InstQueue_reg[13][2]/NET0131  & ~n27972 ;
  assign n36090 = ~n36078 & ~n36089 ;
  assign n36091 = ~n36088 & n36090 ;
  assign n36092 = ~n36085 & n36091 ;
  assign n36098 = n27901 & ~n35971 ;
  assign n36099 = n28108 & ~n35975 ;
  assign n36100 = ~n36098 & ~n36099 ;
  assign n36101 = \P1_P2_DataWidth_reg[1]/NET0131  & ~n36100 ;
  assign n36093 = ~n28072 & ~n35963 ;
  assign n36094 = \P1_P2_InstQueue_reg[14][2]/NET0131  & ~n28068 ;
  assign n36095 = ~n28065 & n36094 ;
  assign n36096 = ~n36093 & ~n36095 ;
  assign n36102 = ~n28160 & ~n36096 ;
  assign n36103 = ~n36101 & ~n36102 ;
  assign n36104 = n25928 & ~n36103 ;
  assign n36105 = ~n25604 & n28068 ;
  assign n36106 = ~n36094 & ~n36105 ;
  assign n36107 = n27608 & ~n36106 ;
  assign n36097 = n27898 & ~n36096 ;
  assign n36108 = \P1_P2_InstQueue_reg[14][2]/NET0131  & ~n27972 ;
  assign n36109 = ~n36097 & ~n36108 ;
  assign n36110 = ~n36107 & n36109 ;
  assign n36111 = ~n36104 & n36110 ;
  assign n36117 = n28108 & ~n35971 ;
  assign n36118 = n28065 & ~n35975 ;
  assign n36119 = ~n36117 & ~n36118 ;
  assign n36120 = \P1_P2_DataWidth_reg[1]/NET0131  & ~n36119 ;
  assign n36112 = ~n28171 & ~n35963 ;
  assign n36113 = \P1_P2_InstQueue_reg[15][2]/NET0131  & ~n28057 ;
  assign n36114 = ~n28068 & n36113 ;
  assign n36115 = ~n36112 & ~n36114 ;
  assign n36121 = ~n28181 & ~n36115 ;
  assign n36122 = ~n36120 & ~n36121 ;
  assign n36123 = n25928 & ~n36122 ;
  assign n36124 = ~n25604 & n28057 ;
  assign n36125 = ~n36113 & ~n36124 ;
  assign n36126 = n27608 & ~n36125 ;
  assign n36116 = n27898 & ~n36115 ;
  assign n36127 = \P1_P2_InstQueue_reg[15][2]/NET0131  & ~n27972 ;
  assign n36128 = ~n36116 & ~n36127 ;
  assign n36129 = ~n36126 & n36128 ;
  assign n36130 = ~n36123 & n36129 ;
  assign n36136 = n28068 & ~n35971 ;
  assign n36137 = n28057 & ~n35975 ;
  assign n36138 = ~n36136 & ~n36137 ;
  assign n36139 = \P1_P2_DataWidth_reg[1]/NET0131  & ~n36138 ;
  assign n36131 = ~n28193 & ~n35963 ;
  assign n36132 = \P1_P2_InstQueue_reg[1][2]/NET0131  & ~n28192 ;
  assign n36133 = ~n28055 & n36132 ;
  assign n36134 = ~n36131 & ~n36133 ;
  assign n36140 = ~n28203 & ~n36134 ;
  assign n36141 = ~n36139 & ~n36140 ;
  assign n36142 = n25928 & ~n36141 ;
  assign n36143 = ~n25604 & n28192 ;
  assign n36144 = ~n36132 & ~n36143 ;
  assign n36145 = n27608 & ~n36144 ;
  assign n36135 = n27898 & ~n36134 ;
  assign n36146 = \P1_P2_InstQueue_reg[1][2]/NET0131  & ~n27972 ;
  assign n36147 = ~n36135 & ~n36146 ;
  assign n36148 = ~n36145 & n36147 ;
  assign n36149 = ~n36142 & n36148 ;
  assign n36155 = n28057 & ~n35971 ;
  assign n36156 = n28055 & ~n35975 ;
  assign n36157 = ~n36155 & ~n36156 ;
  assign n36158 = \P1_P2_DataWidth_reg[1]/NET0131  & ~n36157 ;
  assign n36150 = ~n28215 & ~n35963 ;
  assign n36151 = \P1_P2_InstQueue_reg[2][2]/NET0131  & ~n28214 ;
  assign n36152 = ~n28192 & n36151 ;
  assign n36153 = ~n36150 & ~n36152 ;
  assign n36159 = ~n28225 & ~n36153 ;
  assign n36160 = ~n36158 & ~n36159 ;
  assign n36161 = n25928 & ~n36160 ;
  assign n36162 = ~n25604 & n28214 ;
  assign n36163 = ~n36151 & ~n36162 ;
  assign n36164 = n27608 & ~n36163 ;
  assign n36154 = n27898 & ~n36153 ;
  assign n36165 = \P1_P2_InstQueue_reg[2][2]/NET0131  & ~n27972 ;
  assign n36166 = ~n36154 & ~n36165 ;
  assign n36167 = ~n36164 & n36166 ;
  assign n36168 = ~n36161 & n36167 ;
  assign n36174 = n28055 & ~n35971 ;
  assign n36175 = n28192 & ~n35975 ;
  assign n36176 = ~n36174 & ~n36175 ;
  assign n36177 = \P1_P2_DataWidth_reg[1]/NET0131  & ~n36176 ;
  assign n36169 = ~n28237 & ~n35963 ;
  assign n36170 = \P1_P2_InstQueue_reg[3][2]/NET0131  & ~n28236 ;
  assign n36171 = ~n28214 & n36170 ;
  assign n36172 = ~n36169 & ~n36171 ;
  assign n36178 = ~n28247 & ~n36172 ;
  assign n36179 = ~n36177 & ~n36178 ;
  assign n36180 = n25928 & ~n36179 ;
  assign n36181 = ~n25604 & n28236 ;
  assign n36182 = ~n36170 & ~n36181 ;
  assign n36183 = n27608 & ~n36182 ;
  assign n36173 = n27898 & ~n36172 ;
  assign n36184 = \P1_P2_InstQueue_reg[3][2]/NET0131  & ~n27972 ;
  assign n36185 = ~n36173 & ~n36184 ;
  assign n36186 = ~n36183 & n36185 ;
  assign n36187 = ~n36180 & n36186 ;
  assign n36193 = n28192 & ~n35971 ;
  assign n36194 = n28214 & ~n35975 ;
  assign n36195 = ~n36193 & ~n36194 ;
  assign n36196 = \P1_P2_DataWidth_reg[1]/NET0131  & ~n36195 ;
  assign n36188 = ~n28259 & ~n35963 ;
  assign n36189 = \P1_P2_InstQueue_reg[4][2]/NET0131  & ~n28258 ;
  assign n36190 = ~n28236 & n36189 ;
  assign n36191 = ~n36188 & ~n36190 ;
  assign n36197 = ~n28269 & ~n36191 ;
  assign n36198 = ~n36196 & ~n36197 ;
  assign n36199 = n25928 & ~n36198 ;
  assign n36200 = ~n25604 & n28258 ;
  assign n36201 = ~n36189 & ~n36200 ;
  assign n36202 = n27608 & ~n36201 ;
  assign n36192 = n27898 & ~n36191 ;
  assign n36203 = \P1_P2_InstQueue_reg[4][2]/NET0131  & ~n27972 ;
  assign n36204 = ~n36192 & ~n36203 ;
  assign n36205 = ~n36202 & n36204 ;
  assign n36206 = ~n36199 & n36205 ;
  assign n36212 = n28214 & ~n35971 ;
  assign n36213 = n28236 & ~n35975 ;
  assign n36214 = ~n36212 & ~n36213 ;
  assign n36215 = \P1_P2_DataWidth_reg[1]/NET0131  & ~n36214 ;
  assign n36207 = ~n28281 & ~n35963 ;
  assign n36208 = \P1_P2_InstQueue_reg[5][2]/NET0131  & ~n28280 ;
  assign n36209 = ~n28258 & n36208 ;
  assign n36210 = ~n36207 & ~n36209 ;
  assign n36216 = ~n28291 & ~n36210 ;
  assign n36217 = ~n36215 & ~n36216 ;
  assign n36218 = n25928 & ~n36217 ;
  assign n36219 = ~n25604 & n28280 ;
  assign n36220 = ~n36208 & ~n36219 ;
  assign n36221 = n27608 & ~n36220 ;
  assign n36211 = n27898 & ~n36210 ;
  assign n36222 = \P1_P2_InstQueue_reg[5][2]/NET0131  & ~n27972 ;
  assign n36223 = ~n36211 & ~n36222 ;
  assign n36224 = ~n36221 & n36223 ;
  assign n36225 = ~n36218 & n36224 ;
  assign n36231 = n28236 & ~n35971 ;
  assign n36232 = n28258 & ~n35975 ;
  assign n36233 = ~n36231 & ~n36232 ;
  assign n36234 = \P1_P2_DataWidth_reg[1]/NET0131  & ~n36233 ;
  assign n36226 = ~n28303 & ~n35963 ;
  assign n36227 = \P1_P2_InstQueue_reg[6][2]/NET0131  & ~n28302 ;
  assign n36228 = ~n28280 & n36227 ;
  assign n36229 = ~n36226 & ~n36228 ;
  assign n36235 = ~n28313 & ~n36229 ;
  assign n36236 = ~n36234 & ~n36235 ;
  assign n36237 = n25928 & ~n36236 ;
  assign n36238 = ~n25604 & n28302 ;
  assign n36239 = ~n36227 & ~n36238 ;
  assign n36240 = n27608 & ~n36239 ;
  assign n36230 = n27898 & ~n36229 ;
  assign n36241 = \P1_P2_InstQueue_reg[6][2]/NET0131  & ~n27972 ;
  assign n36242 = ~n36230 & ~n36241 ;
  assign n36243 = ~n36240 & n36242 ;
  assign n36244 = ~n36237 & n36243 ;
  assign n36250 = n28258 & ~n35971 ;
  assign n36251 = n28280 & ~n35975 ;
  assign n36252 = ~n36250 & ~n36251 ;
  assign n36253 = \P1_P2_DataWidth_reg[1]/NET0131  & ~n36252 ;
  assign n36245 = ~n28324 & ~n35963 ;
  assign n36246 = \P1_P2_InstQueue_reg[7][2]/NET0131  & ~n28090 ;
  assign n36247 = ~n28302 & n36246 ;
  assign n36248 = ~n36245 & ~n36247 ;
  assign n36254 = ~n28334 & ~n36248 ;
  assign n36255 = ~n36253 & ~n36254 ;
  assign n36256 = n25928 & ~n36255 ;
  assign n36257 = ~n25604 & n28090 ;
  assign n36258 = ~n36246 & ~n36257 ;
  assign n36259 = n27608 & ~n36258 ;
  assign n36249 = n27898 & ~n36248 ;
  assign n36260 = \P1_P2_InstQueue_reg[7][2]/NET0131  & ~n27972 ;
  assign n36261 = ~n36249 & ~n36260 ;
  assign n36262 = ~n36259 & n36261 ;
  assign n36263 = ~n36256 & n36262 ;
  assign n36269 = n28280 & ~n35971 ;
  assign n36270 = n28302 & ~n35975 ;
  assign n36271 = ~n36269 & ~n36270 ;
  assign n36272 = \P1_P2_DataWidth_reg[1]/NET0131  & ~n36271 ;
  assign n36264 = ~n28095 & ~n35963 ;
  assign n36265 = \P1_P2_InstQueue_reg[8][2]/NET0131  & ~n27945 ;
  assign n36266 = ~n28090 & n36265 ;
  assign n36267 = ~n36264 & ~n36266 ;
  assign n36273 = ~n28354 & ~n36267 ;
  assign n36274 = ~n36272 & ~n36273 ;
  assign n36275 = n25928 & ~n36274 ;
  assign n36276 = ~n25604 & n27945 ;
  assign n36277 = ~n36265 & ~n36276 ;
  assign n36278 = n27608 & ~n36277 ;
  assign n36268 = n27898 & ~n36267 ;
  assign n36279 = \P1_P2_InstQueue_reg[8][2]/NET0131  & ~n27972 ;
  assign n36280 = ~n36268 & ~n36279 ;
  assign n36281 = ~n36278 & n36280 ;
  assign n36282 = ~n36275 & n36281 ;
  assign n36288 = n28302 & ~n35971 ;
  assign n36289 = n28090 & ~n35975 ;
  assign n36290 = ~n36288 & ~n36289 ;
  assign n36291 = \P1_P2_DataWidth_reg[1]/NET0131  & ~n36290 ;
  assign n36283 = ~n27959 & ~n35963 ;
  assign n36284 = \P1_P2_InstQueue_reg[9][2]/NET0131  & ~n27952 ;
  assign n36285 = ~n27945 & n36284 ;
  assign n36286 = ~n36283 & ~n36285 ;
  assign n36292 = ~n28374 & ~n36286 ;
  assign n36293 = ~n36291 & ~n36292 ;
  assign n36294 = n25928 & ~n36293 ;
  assign n36295 = ~n25604 & n27952 ;
  assign n36296 = ~n36284 & ~n36295 ;
  assign n36297 = n27608 & ~n36296 ;
  assign n36287 = n27898 & ~n36286 ;
  assign n36298 = \P1_P2_InstQueue_reg[9][2]/NET0131  & ~n27972 ;
  assign n36299 = ~n36287 & ~n36298 ;
  assign n36300 = ~n36297 & n36299 ;
  assign n36301 = ~n36294 & n36300 ;
  assign n36310 = n28398 & ~n36002 ;
  assign n36311 = n28401 & ~n36006 ;
  assign n36312 = ~n36310 & ~n36311 ;
  assign n36313 = \P2_P2_DataWidth_reg[1]/NET0131  & ~n36312 ;
  assign n36302 = ~n28388 & ~n35991 ;
  assign n36303 = \P2_P2_InstQueue_reg[0][2]/NET0131  & ~n28385 ;
  assign n36304 = ~n28387 & n36303 ;
  assign n36305 = ~n36302 & ~n36304 ;
  assign n36314 = ~n28406 & ~n36305 ;
  assign n36315 = ~n36313 & ~n36314 ;
  assign n36316 = n26794 & ~n36315 ;
  assign n36307 = ~n26481 & n28385 ;
  assign n36308 = ~n36303 & ~n36307 ;
  assign n36309 = n27613 & ~n36308 ;
  assign n36306 = n27977 & ~n36305 ;
  assign n36317 = \P2_P2_InstQueue_reg[0][2]/NET0131  & ~n28050 ;
  assign n36318 = ~n36306 & ~n36317 ;
  assign n36319 = ~n36309 & n36318 ;
  assign n36320 = ~n36316 & n36319 ;
  assign n36329 = n28423 & ~n36002 ;
  assign n36330 = n28027 & ~n36006 ;
  assign n36331 = ~n36329 & ~n36330 ;
  assign n36332 = \P2_P2_DataWidth_reg[1]/NET0131  & ~n36331 ;
  assign n36321 = ~n28414 & ~n35991 ;
  assign n36322 = \P2_P2_InstQueue_reg[10][2]/NET0131  & ~n27983 ;
  assign n36323 = ~n28034 & n36322 ;
  assign n36324 = ~n36321 & ~n36323 ;
  assign n36333 = ~n28429 & ~n36324 ;
  assign n36334 = ~n36332 & ~n36333 ;
  assign n36335 = n26794 & ~n36334 ;
  assign n36326 = ~n26481 & n27983 ;
  assign n36327 = ~n36322 & ~n36326 ;
  assign n36328 = n27613 & ~n36327 ;
  assign n36325 = n27977 & ~n36324 ;
  assign n36336 = \P2_P2_InstQueue_reg[10][2]/NET0131  & ~n28050 ;
  assign n36337 = ~n36325 & ~n36336 ;
  assign n36338 = ~n36328 & n36337 ;
  assign n36339 = ~n36335 & n36338 ;
  assign n36348 = n28034 & ~n36002 ;
  assign n36349 = n27983 & ~n36006 ;
  assign n36350 = ~n36348 & ~n36349 ;
  assign n36351 = \P2_P2_DataWidth_reg[1]/NET0131  & ~n36350 ;
  assign n36340 = ~n28439 & ~n35991 ;
  assign n36341 = \P2_P2_InstQueue_reg[12][2]/NET0131  & ~n28438 ;
  assign n36342 = ~n27980 & n36341 ;
  assign n36343 = ~n36340 & ~n36342 ;
  assign n36352 = ~n28452 & ~n36343 ;
  assign n36353 = ~n36351 & ~n36352 ;
  assign n36354 = n26794 & ~n36353 ;
  assign n36345 = ~n26481 & n28438 ;
  assign n36346 = ~n36341 & ~n36345 ;
  assign n36347 = n27613 & ~n36346 ;
  assign n36344 = n27977 & ~n36343 ;
  assign n36355 = \P2_P2_InstQueue_reg[12][2]/NET0131  & ~n28050 ;
  assign n36356 = ~n36344 & ~n36355 ;
  assign n36357 = ~n36347 & n36356 ;
  assign n36358 = ~n36354 & n36357 ;
  assign n36367 = n27983 & ~n36002 ;
  assign n36368 = n27980 & ~n36006 ;
  assign n36369 = ~n36367 & ~n36368 ;
  assign n36370 = \P2_P2_DataWidth_reg[1]/NET0131  & ~n36369 ;
  assign n36359 = ~n28460 & ~n35991 ;
  assign n36360 = \P2_P2_InstQueue_reg[13][2]/NET0131  & ~n28398 ;
  assign n36361 = ~n28438 & n36360 ;
  assign n36362 = ~n36359 & ~n36361 ;
  assign n36371 = ~n28473 & ~n36362 ;
  assign n36372 = ~n36370 & ~n36371 ;
  assign n36373 = n26794 & ~n36372 ;
  assign n36364 = ~n26481 & n28398 ;
  assign n36365 = ~n36360 & ~n36364 ;
  assign n36366 = n27613 & ~n36365 ;
  assign n36363 = n27977 & ~n36362 ;
  assign n36374 = \P2_P2_InstQueue_reg[13][2]/NET0131  & ~n28050 ;
  assign n36375 = ~n36363 & ~n36374 ;
  assign n36376 = ~n36366 & n36375 ;
  assign n36377 = ~n36373 & n36376 ;
  assign n36386 = n27980 & ~n36002 ;
  assign n36387 = n28438 & ~n36006 ;
  assign n36388 = ~n36386 & ~n36387 ;
  assign n36389 = \P2_P2_DataWidth_reg[1]/NET0131  & ~n36388 ;
  assign n36378 = ~n28405 & ~n35991 ;
  assign n36379 = \P2_P2_InstQueue_reg[14][2]/NET0131  & ~n28401 ;
  assign n36380 = ~n28398 & n36379 ;
  assign n36381 = ~n36378 & ~n36380 ;
  assign n36390 = ~n28493 & ~n36381 ;
  assign n36391 = ~n36389 & ~n36390 ;
  assign n36392 = n26794 & ~n36391 ;
  assign n36383 = ~n26481 & n28401 ;
  assign n36384 = ~n36379 & ~n36383 ;
  assign n36385 = n27613 & ~n36384 ;
  assign n36382 = n27977 & ~n36381 ;
  assign n36393 = \P2_P2_InstQueue_reg[14][2]/NET0131  & ~n28050 ;
  assign n36394 = ~n36382 & ~n36393 ;
  assign n36395 = ~n36385 & n36394 ;
  assign n36396 = ~n36392 & n36395 ;
  assign n36405 = n28438 & ~n36002 ;
  assign n36406 = n28398 & ~n36006 ;
  assign n36407 = ~n36405 & ~n36406 ;
  assign n36408 = \P2_P2_DataWidth_reg[1]/NET0131  & ~n36407 ;
  assign n36397 = ~n28501 & ~n35991 ;
  assign n36398 = \P2_P2_InstQueue_reg[15][2]/NET0131  & ~n28387 ;
  assign n36399 = ~n28401 & n36398 ;
  assign n36400 = ~n36397 & ~n36399 ;
  assign n36409 = ~n28514 & ~n36400 ;
  assign n36410 = ~n36408 & ~n36409 ;
  assign n36411 = n26794 & ~n36410 ;
  assign n36402 = ~n26481 & n28387 ;
  assign n36403 = ~n36398 & ~n36402 ;
  assign n36404 = n27613 & ~n36403 ;
  assign n36401 = n27977 & ~n36400 ;
  assign n36412 = \P2_P2_InstQueue_reg[15][2]/NET0131  & ~n28050 ;
  assign n36413 = ~n36401 & ~n36412 ;
  assign n36414 = ~n36404 & n36413 ;
  assign n36415 = ~n36411 & n36414 ;
  assign n36424 = n28401 & ~n36002 ;
  assign n36425 = n28387 & ~n36006 ;
  assign n36426 = ~n36424 & ~n36425 ;
  assign n36427 = \P2_P2_DataWidth_reg[1]/NET0131  & ~n36426 ;
  assign n36416 = ~n28523 & ~n35991 ;
  assign n36417 = \P2_P2_InstQueue_reg[1][2]/NET0131  & ~n28522 ;
  assign n36418 = ~n28385 & n36417 ;
  assign n36419 = ~n36416 & ~n36418 ;
  assign n36428 = ~n28536 & ~n36419 ;
  assign n36429 = ~n36427 & ~n36428 ;
  assign n36430 = n26794 & ~n36429 ;
  assign n36421 = ~n26481 & n28522 ;
  assign n36422 = ~n36417 & ~n36421 ;
  assign n36423 = n27613 & ~n36422 ;
  assign n36420 = n27977 & ~n36419 ;
  assign n36431 = \P2_P2_InstQueue_reg[1][2]/NET0131  & ~n28050 ;
  assign n36432 = ~n36420 & ~n36431 ;
  assign n36433 = ~n36423 & n36432 ;
  assign n36434 = ~n36430 & n36433 ;
  assign n36443 = n28387 & ~n36002 ;
  assign n36444 = n28385 & ~n36006 ;
  assign n36445 = ~n36443 & ~n36444 ;
  assign n36446 = \P2_P2_DataWidth_reg[1]/NET0131  & ~n36445 ;
  assign n36435 = ~n28545 & ~n35991 ;
  assign n36436 = \P2_P2_InstQueue_reg[2][2]/NET0131  & ~n28544 ;
  assign n36437 = ~n28522 & n36436 ;
  assign n36438 = ~n36435 & ~n36437 ;
  assign n36447 = ~n28558 & ~n36438 ;
  assign n36448 = ~n36446 & ~n36447 ;
  assign n36449 = n26794 & ~n36448 ;
  assign n36440 = ~n26481 & n28544 ;
  assign n36441 = ~n36436 & ~n36440 ;
  assign n36442 = n27613 & ~n36441 ;
  assign n36439 = n27977 & ~n36438 ;
  assign n36450 = \P2_P2_InstQueue_reg[2][2]/NET0131  & ~n28050 ;
  assign n36451 = ~n36439 & ~n36450 ;
  assign n36452 = ~n36442 & n36451 ;
  assign n36453 = ~n36449 & n36452 ;
  assign n36462 = n28385 & ~n36002 ;
  assign n36463 = n28522 & ~n36006 ;
  assign n36464 = ~n36462 & ~n36463 ;
  assign n36465 = \P2_P2_DataWidth_reg[1]/NET0131  & ~n36464 ;
  assign n36454 = ~n28567 & ~n35991 ;
  assign n36455 = \P2_P2_InstQueue_reg[3][2]/NET0131  & ~n28566 ;
  assign n36456 = ~n28544 & n36455 ;
  assign n36457 = ~n36454 & ~n36456 ;
  assign n36466 = ~n28580 & ~n36457 ;
  assign n36467 = ~n36465 & ~n36466 ;
  assign n36468 = n26794 & ~n36467 ;
  assign n36459 = ~n26481 & n28566 ;
  assign n36460 = ~n36455 & ~n36459 ;
  assign n36461 = n27613 & ~n36460 ;
  assign n36458 = n27977 & ~n36457 ;
  assign n36469 = \P2_P2_InstQueue_reg[3][2]/NET0131  & ~n28050 ;
  assign n36470 = ~n36458 & ~n36469 ;
  assign n36471 = ~n36461 & n36470 ;
  assign n36472 = ~n36468 & n36471 ;
  assign n36481 = n28522 & ~n36002 ;
  assign n36482 = n28544 & ~n36006 ;
  assign n36483 = ~n36481 & ~n36482 ;
  assign n36484 = \P2_P2_DataWidth_reg[1]/NET0131  & ~n36483 ;
  assign n36473 = ~n28589 & ~n35991 ;
  assign n36474 = \P2_P2_InstQueue_reg[4][2]/NET0131  & ~n28588 ;
  assign n36475 = ~n28566 & n36474 ;
  assign n36476 = ~n36473 & ~n36475 ;
  assign n36485 = ~n28602 & ~n36476 ;
  assign n36486 = ~n36484 & ~n36485 ;
  assign n36487 = n26794 & ~n36486 ;
  assign n36478 = ~n26481 & n28588 ;
  assign n36479 = ~n36474 & ~n36478 ;
  assign n36480 = n27613 & ~n36479 ;
  assign n36477 = n27977 & ~n36476 ;
  assign n36488 = \P2_P2_InstQueue_reg[4][2]/NET0131  & ~n28050 ;
  assign n36489 = ~n36477 & ~n36488 ;
  assign n36490 = ~n36480 & n36489 ;
  assign n36491 = ~n36487 & n36490 ;
  assign n36500 = n28544 & ~n36002 ;
  assign n36501 = n28566 & ~n36006 ;
  assign n36502 = ~n36500 & ~n36501 ;
  assign n36503 = \P2_P2_DataWidth_reg[1]/NET0131  & ~n36502 ;
  assign n36492 = ~n28611 & ~n35991 ;
  assign n36493 = \P2_P2_InstQueue_reg[5][2]/NET0131  & ~n28610 ;
  assign n36494 = ~n28588 & n36493 ;
  assign n36495 = ~n36492 & ~n36494 ;
  assign n36504 = ~n28624 & ~n36495 ;
  assign n36505 = ~n36503 & ~n36504 ;
  assign n36506 = n26794 & ~n36505 ;
  assign n36497 = ~n26481 & n28610 ;
  assign n36498 = ~n36493 & ~n36497 ;
  assign n36499 = n27613 & ~n36498 ;
  assign n36496 = n27977 & ~n36495 ;
  assign n36507 = \P2_P2_InstQueue_reg[5][2]/NET0131  & ~n28050 ;
  assign n36508 = ~n36496 & ~n36507 ;
  assign n36509 = ~n36499 & n36508 ;
  assign n36510 = ~n36506 & n36509 ;
  assign n36519 = n28566 & ~n36002 ;
  assign n36520 = n28588 & ~n36006 ;
  assign n36521 = ~n36519 & ~n36520 ;
  assign n36522 = \P2_P2_DataWidth_reg[1]/NET0131  & ~n36521 ;
  assign n36511 = ~n28633 & ~n35991 ;
  assign n36512 = \P2_P2_InstQueue_reg[6][2]/NET0131  & ~n28632 ;
  assign n36513 = ~n28610 & n36512 ;
  assign n36514 = ~n36511 & ~n36513 ;
  assign n36523 = ~n28646 & ~n36514 ;
  assign n36524 = ~n36522 & ~n36523 ;
  assign n36525 = n26794 & ~n36524 ;
  assign n36516 = ~n26481 & n28632 ;
  assign n36517 = ~n36512 & ~n36516 ;
  assign n36518 = n27613 & ~n36517 ;
  assign n36515 = n27977 & ~n36514 ;
  assign n36526 = \P2_P2_InstQueue_reg[6][2]/NET0131  & ~n28050 ;
  assign n36527 = ~n36515 & ~n36526 ;
  assign n36528 = ~n36518 & n36527 ;
  assign n36529 = ~n36525 & n36528 ;
  assign n36538 = n28588 & ~n36002 ;
  assign n36539 = n28610 & ~n36006 ;
  assign n36540 = ~n36538 & ~n36539 ;
  assign n36541 = \P2_P2_DataWidth_reg[1]/NET0131  & ~n36540 ;
  assign n36530 = ~n28654 & ~n35991 ;
  assign n36531 = \P2_P2_InstQueue_reg[7][2]/NET0131  & ~n28423 ;
  assign n36532 = ~n28632 & n36531 ;
  assign n36533 = ~n36530 & ~n36532 ;
  assign n36542 = ~n28667 & ~n36533 ;
  assign n36543 = ~n36541 & ~n36542 ;
  assign n36544 = n26794 & ~n36543 ;
  assign n36535 = ~n26481 & n28423 ;
  assign n36536 = ~n36531 & ~n36535 ;
  assign n36537 = n27613 & ~n36536 ;
  assign n36534 = n27977 & ~n36533 ;
  assign n36545 = \P2_P2_InstQueue_reg[7][2]/NET0131  & ~n28050 ;
  assign n36546 = ~n36534 & ~n36545 ;
  assign n36547 = ~n36537 & n36546 ;
  assign n36548 = ~n36544 & n36547 ;
  assign n36557 = n28610 & ~n36002 ;
  assign n36558 = n28632 & ~n36006 ;
  assign n36559 = ~n36557 & ~n36558 ;
  assign n36560 = \P2_P2_DataWidth_reg[1]/NET0131  & ~n36559 ;
  assign n36549 = ~n28428 & ~n35991 ;
  assign n36550 = \P2_P2_InstQueue_reg[8][2]/NET0131  & ~n28027 ;
  assign n36551 = ~n28423 & n36550 ;
  assign n36552 = ~n36549 & ~n36551 ;
  assign n36561 = ~n28687 & ~n36552 ;
  assign n36562 = ~n36560 & ~n36561 ;
  assign n36563 = n26794 & ~n36562 ;
  assign n36554 = ~n26481 & n28027 ;
  assign n36555 = ~n36550 & ~n36554 ;
  assign n36556 = n27613 & ~n36555 ;
  assign n36553 = n27977 & ~n36552 ;
  assign n36564 = \P2_P2_InstQueue_reg[8][2]/NET0131  & ~n28050 ;
  assign n36565 = ~n36553 & ~n36564 ;
  assign n36566 = ~n36556 & n36565 ;
  assign n36567 = ~n36563 & n36566 ;
  assign n36576 = n28632 & ~n36002 ;
  assign n36577 = n28423 & ~n36006 ;
  assign n36578 = ~n36576 & ~n36577 ;
  assign n36579 = \P2_P2_DataWidth_reg[1]/NET0131  & ~n36578 ;
  assign n36568 = ~n28041 & ~n35991 ;
  assign n36569 = \P2_P2_InstQueue_reg[9][2]/NET0131  & ~n28034 ;
  assign n36570 = ~n28027 & n36569 ;
  assign n36571 = ~n36568 & ~n36570 ;
  assign n36580 = ~n28707 & ~n36571 ;
  assign n36581 = ~n36579 & ~n36580 ;
  assign n36582 = n26794 & ~n36581 ;
  assign n36573 = ~n26481 & n28034 ;
  assign n36574 = ~n36569 & ~n36573 ;
  assign n36575 = n27613 & ~n36574 ;
  assign n36572 = n27977 & ~n36571 ;
  assign n36583 = \P2_P2_InstQueue_reg[9][2]/NET0131  & ~n28050 ;
  assign n36584 = ~n36572 & ~n36583 ;
  assign n36585 = ~n36575 & n36584 ;
  assign n36586 = ~n36582 & n36585 ;
  assign n36587 = \P1_P2_PhyAddrPointer_reg[31]/NET0131  & n25733 ;
  assign n36588 = ~n31333 & ~n36587 ;
  assign n36589 = n25701 & ~n36588 ;
  assign n36590 = ~n25752 & ~n25784 ;
  assign n36591 = \P1_P2_PhyAddrPointer_reg[31]/NET0131  & ~n36590 ;
  assign n36592 = ~n31461 & ~n36591 ;
  assign n36593 = ~n36589 & n36592 ;
  assign n36594 = n25918 & ~n36593 ;
  assign n36597 = \P1_P2_PhyAddrPointer_reg[2]/NET0131  & \P1_P2_PhyAddrPointer_reg[3]/NET0131  ;
  assign n36598 = \P1_P2_PhyAddrPointer_reg[4]/NET0131  & n36597 ;
  assign n36599 = \P1_P2_PhyAddrPointer_reg[5]/NET0131  & n36598 ;
  assign n36600 = \P1_P2_PhyAddrPointer_reg[6]/NET0131  & n36599 ;
  assign n36601 = \P1_P2_PhyAddrPointer_reg[7]/NET0131  & n36600 ;
  assign n36602 = \P1_P2_PhyAddrPointer_reg[8]/NET0131  & n36601 ;
  assign n36603 = \P1_P2_PhyAddrPointer_reg[9]/NET0131  & n36602 ;
  assign n36604 = \P1_P2_PhyAddrPointer_reg[10]/NET0131  & n36603 ;
  assign n36605 = \P1_P2_PhyAddrPointer_reg[11]/NET0131  & n36604 ;
  assign n36606 = \P1_P2_PhyAddrPointer_reg[12]/NET0131  & n36605 ;
  assign n36607 = \P1_P2_PhyAddrPointer_reg[13]/NET0131  & n36606 ;
  assign n36608 = \P1_P2_PhyAddrPointer_reg[14]/NET0131  & n36607 ;
  assign n36609 = \P1_P2_PhyAddrPointer_reg[15]/NET0131  & n36608 ;
  assign n36610 = \P1_P2_PhyAddrPointer_reg[16]/NET0131  & n36609 ;
  assign n36611 = \P1_P2_PhyAddrPointer_reg[17]/NET0131  & n36610 ;
  assign n36612 = \P1_P2_PhyAddrPointer_reg[18]/NET0131  & n36611 ;
  assign n36613 = \P1_P2_PhyAddrPointer_reg[19]/NET0131  & n36612 ;
  assign n36614 = \P1_P2_PhyAddrPointer_reg[20]/NET0131  & n36613 ;
  assign n36615 = \P1_P2_PhyAddrPointer_reg[21]/NET0131  & n36614 ;
  assign n36616 = \P1_P2_PhyAddrPointer_reg[22]/NET0131  & n36615 ;
  assign n36617 = \P1_P2_PhyAddrPointer_reg[23]/NET0131  & n36616 ;
  assign n36618 = \P1_P2_PhyAddrPointer_reg[24]/NET0131  & n36617 ;
  assign n36619 = \P1_P2_PhyAddrPointer_reg[25]/NET0131  & n36618 ;
  assign n36620 = \P1_P2_PhyAddrPointer_reg[26]/NET0131  & n36619 ;
  assign n36621 = \P1_P2_PhyAddrPointer_reg[27]/NET0131  & n36620 ;
  assign n36622 = \P1_P2_PhyAddrPointer_reg[28]/NET0131  & n36621 ;
  assign n36623 = \P1_P2_PhyAddrPointer_reg[29]/NET0131  & n36622 ;
  assign n36624 = \P1_P2_PhyAddrPointer_reg[30]/NET0131  & n36623 ;
  assign n36625 = \P1_P2_PhyAddrPointer_reg[1]/NET0131  & n36624 ;
  assign n36626 = \P1_P2_PhyAddrPointer_reg[31]/NET0131  & ~n36625 ;
  assign n36627 = ~\P1_P2_PhyAddrPointer_reg[31]/NET0131  & n36625 ;
  assign n36628 = ~n36626 & ~n36627 ;
  assign n36629 = \P1_P2_DataWidth_reg[1]/NET0131  & ~n27898 ;
  assign n36630 = ~n28928 & ~n36629 ;
  assign n36631 = ~n36628 & n36630 ;
  assign n36633 = \P1_P2_PhyAddrPointer_reg[31]/NET0131  & n36624 ;
  assign n36632 = ~\P1_P2_PhyAddrPointer_reg[31]/NET0131  & ~n36624 ;
  assign n36634 = n25933 & ~n36632 ;
  assign n36635 = ~n36633 & n36634 ;
  assign n36595 = n27970 & ~n31484 ;
  assign n36596 = \P1_P2_PhyAddrPointer_reg[31]/NET0131  & ~n36595 ;
  assign n36636 = ~n31489 & ~n36596 ;
  assign n36637 = ~n36635 & n36636 ;
  assign n36638 = ~n36631 & n36637 ;
  assign n36639 = ~n36594 & n36638 ;
  assign n36676 = n25945 & n32022 ;
  assign n36677 = ~n25982 & ~n26054 ;
  assign n36678 = ~n26052 & n36677 ;
  assign n36679 = \P2_P1_PhyAddrPointer_reg[31]/NET0131  & ~n36678 ;
  assign n36680 = ~n32157 & ~n36679 ;
  assign n36681 = ~n36676 & n36680 ;
  assign n36682 = n11623 & ~n36681 ;
  assign n36640 = \P2_P1_PhyAddrPointer_reg[23]/NET0131  & \P2_P1_PhyAddrPointer_reg[24]/NET0131  ;
  assign n36641 = \P2_P1_PhyAddrPointer_reg[12]/NET0131  & \P2_P1_PhyAddrPointer_reg[13]/NET0131  ;
  assign n36642 = \P2_P1_PhyAddrPointer_reg[14]/NET0131  & n36641 ;
  assign n36643 = \P2_P1_PhyAddrPointer_reg[2]/NET0131  & \P2_P1_PhyAddrPointer_reg[3]/NET0131  ;
  assign n36644 = \P2_P1_PhyAddrPointer_reg[4]/NET0131  & n36643 ;
  assign n36645 = \P2_P1_PhyAddrPointer_reg[5]/NET0131  & n36644 ;
  assign n36646 = \P2_P1_PhyAddrPointer_reg[6]/NET0131  & n36645 ;
  assign n36647 = \P2_P1_PhyAddrPointer_reg[7]/NET0131  & n36646 ;
  assign n36648 = \P2_P1_PhyAddrPointer_reg[8]/NET0131  & n36647 ;
  assign n36649 = \P2_P1_PhyAddrPointer_reg[9]/NET0131  & n36648 ;
  assign n36650 = \P2_P1_PhyAddrPointer_reg[10]/NET0131  & n36649 ;
  assign n36651 = \P2_P1_PhyAddrPointer_reg[11]/NET0131  & n36650 ;
  assign n36652 = n36642 & n36651 ;
  assign n36653 = \P2_P1_PhyAddrPointer_reg[15]/NET0131  & n36652 ;
  assign n36654 = \P2_P1_PhyAddrPointer_reg[16]/NET0131  & \P2_P1_PhyAddrPointer_reg[17]/NET0131  ;
  assign n36655 = \P2_P1_PhyAddrPointer_reg[18]/NET0131  & \P2_P1_PhyAddrPointer_reg[19]/NET0131  ;
  assign n36656 = n36654 & n36655 ;
  assign n36657 = n36653 & n36656 ;
  assign n36658 = \P2_P1_PhyAddrPointer_reg[20]/NET0131  & n36657 ;
  assign n36659 = \P2_P1_PhyAddrPointer_reg[21]/NET0131  & n36658 ;
  assign n36660 = \P2_P1_PhyAddrPointer_reg[22]/NET0131  & n36659 ;
  assign n36661 = n36640 & n36660 ;
  assign n36662 = \P2_P1_PhyAddrPointer_reg[25]/NET0131  & n36661 ;
  assign n36663 = \P2_P1_PhyAddrPointer_reg[26]/NET0131  & n36662 ;
  assign n36664 = \P2_P1_PhyAddrPointer_reg[27]/NET0131  & n36663 ;
  assign n36665 = \P2_P1_PhyAddrPointer_reg[28]/NET0131  & n36664 ;
  assign n36666 = \P2_P1_PhyAddrPointer_reg[29]/NET0131  & n36665 ;
  assign n36667 = \P2_P1_PhyAddrPointer_reg[30]/NET0131  & n36666 ;
  assign n36668 = \P2_P1_PhyAddrPointer_reg[1]/NET0131  & n36667 ;
  assign n36669 = ~\P2_P1_PhyAddrPointer_reg[31]/NET0131  & ~n36668 ;
  assign n36670 = \P2_P1_PhyAddrPointer_reg[31]/NET0131  & n36667 ;
  assign n36671 = \P2_P1_PhyAddrPointer_reg[1]/NET0131  & n36670 ;
  assign n36672 = ~n36669 & ~n36671 ;
  assign n36673 = \P2_P1_DataWidth_reg[1]/NET0131  & ~n11613 ;
  assign n36674 = ~n12341 & ~n36673 ;
  assign n36675 = n36672 & n36674 ;
  assign n36683 = ~\P2_P1_PhyAddrPointer_reg[31]/NET0131  & ~n36667 ;
  assign n36684 = n27681 & ~n36670 ;
  assign n36685 = ~n36683 & n36684 ;
  assign n36686 = ~n11618 & ~n25942 ;
  assign n36687 = n21097 & n36686 ;
  assign n36688 = \P2_P1_PhyAddrPointer_reg[31]/NET0131  & ~n36687 ;
  assign n36689 = ~n32174 & ~n36688 ;
  assign n36690 = ~n36685 & n36689 ;
  assign n36691 = ~n36675 & n36690 ;
  assign n36692 = ~n36682 & n36691 ;
  assign n36693 = \P1_P1_PhyAddrPointer_reg[31]/NET0131  & n26249 ;
  assign n36694 = ~n34019 & ~n36693 ;
  assign n36695 = n26126 & ~n36694 ;
  assign n36696 = ~n26127 & ~n26251 ;
  assign n36697 = \P1_P1_PhyAddrPointer_reg[31]/NET0131  & ~n36696 ;
  assign n36698 = ~n34139 & ~n36697 ;
  assign n36699 = ~n36695 & n36698 ;
  assign n36700 = n8355 & ~n36699 ;
  assign n36701 = ~n8287 & ~n26280 ;
  assign n36702 = \P1_P1_PhyAddrPointer_reg[2]/NET0131  & \P1_P1_PhyAddrPointer_reg[3]/NET0131  ;
  assign n36703 = \P1_P1_PhyAddrPointer_reg[4]/NET0131  & n36702 ;
  assign n36704 = \P1_P1_PhyAddrPointer_reg[5]/NET0131  & n36703 ;
  assign n36705 = \P1_P1_PhyAddrPointer_reg[6]/NET0131  & n36704 ;
  assign n36706 = \P1_P1_PhyAddrPointer_reg[7]/NET0131  & n36705 ;
  assign n36707 = \P1_P1_PhyAddrPointer_reg[8]/NET0131  & n36706 ;
  assign n36708 = \P1_P1_PhyAddrPointer_reg[9]/NET0131  & n36707 ;
  assign n36709 = \P1_P1_PhyAddrPointer_reg[10]/NET0131  & n36708 ;
  assign n36710 = \P1_P1_PhyAddrPointer_reg[11]/NET0131  & n36709 ;
  assign n36711 = \P1_P1_PhyAddrPointer_reg[12]/NET0131  & n36710 ;
  assign n36712 = \P1_P1_PhyAddrPointer_reg[13]/NET0131  & n36711 ;
  assign n36713 = \P1_P1_PhyAddrPointer_reg[14]/NET0131  & n36712 ;
  assign n36714 = \P1_P1_PhyAddrPointer_reg[15]/NET0131  & n36713 ;
  assign n36715 = \P1_P1_PhyAddrPointer_reg[16]/NET0131  & n36714 ;
  assign n36716 = \P1_P1_PhyAddrPointer_reg[17]/NET0131  & n36715 ;
  assign n36717 = \P1_P1_PhyAddrPointer_reg[18]/NET0131  & n36716 ;
  assign n36718 = \P1_P1_PhyAddrPointer_reg[19]/NET0131  & n36717 ;
  assign n36719 = \P1_P1_PhyAddrPointer_reg[20]/NET0131  & n36718 ;
  assign n36720 = \P1_P1_PhyAddrPointer_reg[21]/NET0131  & n36719 ;
  assign n36721 = \P1_P1_PhyAddrPointer_reg[22]/NET0131  & n36720 ;
  assign n36722 = \P1_P1_PhyAddrPointer_reg[23]/NET0131  & n36721 ;
  assign n36723 = \P1_P1_PhyAddrPointer_reg[24]/NET0131  & n36722 ;
  assign n36724 = \P1_P1_PhyAddrPointer_reg[25]/NET0131  & n36723 ;
  assign n36725 = \P1_P1_PhyAddrPointer_reg[26]/NET0131  & n36724 ;
  assign n36726 = \P1_P1_PhyAddrPointer_reg[27]/NET0131  & n36725 ;
  assign n36727 = \P1_P1_PhyAddrPointer_reg[1]/NET0131  & n36726 ;
  assign n36728 = \P1_P1_PhyAddrPointer_reg[28]/NET0131  & n36727 ;
  assign n36729 = \P1_P1_PhyAddrPointer_reg[29]/NET0131  & n36728 ;
  assign n36730 = \P1_P1_PhyAddrPointer_reg[30]/NET0131  & n36729 ;
  assign n36731 = \P1_P1_PhyAddrPointer_reg[31]/NET0131  & ~n36730 ;
  assign n36732 = ~\P1_P1_PhyAddrPointer_reg[31]/NET0131  & n36730 ;
  assign n36733 = ~n36731 & ~n36732 ;
  assign n36734 = ~n36701 & ~n36733 ;
  assign n36735 = \P1_P1_PhyAddrPointer_reg[28]/NET0131  & n36726 ;
  assign n36736 = \P1_P1_PhyAddrPointer_reg[29]/NET0131  & n36735 ;
  assign n36737 = \P1_P1_PhyAddrPointer_reg[30]/NET0131  & n36736 ;
  assign n36739 = \P1_P1_PhyAddrPointer_reg[31]/NET0131  & n36737 ;
  assign n36738 = ~\P1_P1_PhyAddrPointer_reg[31]/NET0131  & ~n36737 ;
  assign n36740 = n27791 & ~n36738 ;
  assign n36741 = ~n36739 & n36740 ;
  assign n36742 = ~n8359 & ~n26115 ;
  assign n36743 = n15323 & n36742 ;
  assign n36744 = \P1_P1_PhyAddrPointer_reg[31]/NET0131  & ~n36743 ;
  assign n36745 = ~n34160 & ~n36744 ;
  assign n36746 = ~n36741 & n36745 ;
  assign n36747 = ~n36734 & n36746 ;
  assign n36748 = ~n36700 & n36747 ;
  assign n36749 = \P2_P2_PhyAddrPointer_reg[31]/NET0131  & n26629 ;
  assign n36750 = ~n32717 & ~n36749 ;
  assign n36751 = n26621 & ~n36750 ;
  assign n36752 = ~n26619 & ~n26676 ;
  assign n36753 = \P2_P2_PhyAddrPointer_reg[31]/NET0131  & ~n36752 ;
  assign n36754 = ~n36751 & ~n36753 ;
  assign n36755 = ~n32849 & n36754 ;
  assign n36756 = n26792 & ~n36755 ;
  assign n36760 = ~n26795 & ~n27977 ;
  assign n36761 = \P2_P2_PhyAddrPointer_reg[2]/NET0131  & \P2_P2_PhyAddrPointer_reg[3]/NET0131  ;
  assign n36762 = \P2_P2_PhyAddrPointer_reg[4]/NET0131  & n36761 ;
  assign n36763 = \P2_P2_PhyAddrPointer_reg[5]/NET0131  & n36762 ;
  assign n36764 = \P2_P2_PhyAddrPointer_reg[6]/NET0131  & n36763 ;
  assign n36765 = \P2_P2_PhyAddrPointer_reg[7]/NET0131  & n36764 ;
  assign n36766 = \P2_P2_PhyAddrPointer_reg[8]/NET0131  & n36765 ;
  assign n36767 = \P2_P2_PhyAddrPointer_reg[9]/NET0131  & n36766 ;
  assign n36768 = \P2_P2_PhyAddrPointer_reg[10]/NET0131  & n36767 ;
  assign n36769 = \P2_P2_PhyAddrPointer_reg[11]/NET0131  & n36768 ;
  assign n36770 = \P2_P2_PhyAddrPointer_reg[12]/NET0131  & n36769 ;
  assign n36771 = \P2_P2_PhyAddrPointer_reg[13]/NET0131  & n36770 ;
  assign n36772 = \P2_P2_PhyAddrPointer_reg[14]/NET0131  & n36771 ;
  assign n36773 = \P2_P2_PhyAddrPointer_reg[15]/NET0131  & n36772 ;
  assign n36774 = \P2_P2_PhyAddrPointer_reg[16]/NET0131  & n36773 ;
  assign n36775 = \P2_P2_PhyAddrPointer_reg[17]/NET0131  & n36774 ;
  assign n36776 = \P2_P2_PhyAddrPointer_reg[18]/NET0131  & n36775 ;
  assign n36777 = \P2_P2_PhyAddrPointer_reg[19]/NET0131  & n36776 ;
  assign n36778 = \P2_P2_PhyAddrPointer_reg[20]/NET0131  & n36777 ;
  assign n36779 = \P2_P2_PhyAddrPointer_reg[21]/NET0131  & n36778 ;
  assign n36780 = \P2_P2_PhyAddrPointer_reg[22]/NET0131  & n36779 ;
  assign n36781 = \P2_P2_PhyAddrPointer_reg[23]/NET0131  & n36780 ;
  assign n36782 = \P2_P2_PhyAddrPointer_reg[24]/NET0131  & n36781 ;
  assign n36783 = \P2_P2_PhyAddrPointer_reg[25]/NET0131  & n36782 ;
  assign n36784 = \P2_P2_PhyAddrPointer_reg[26]/NET0131  & n36783 ;
  assign n36785 = \P2_P2_PhyAddrPointer_reg[27]/NET0131  & n36784 ;
  assign n36786 = \P2_P2_PhyAddrPointer_reg[28]/NET0131  & n36785 ;
  assign n36787 = \P2_P2_PhyAddrPointer_reg[29]/NET0131  & \P2_P2_PhyAddrPointer_reg[30]/NET0131  ;
  assign n36788 = n36786 & n36787 ;
  assign n36789 = \P2_P2_PhyAddrPointer_reg[1]/NET0131  & n36788 ;
  assign n36790 = ~\P2_P2_PhyAddrPointer_reg[31]/NET0131  & ~n36789 ;
  assign n36791 = \P2_P2_PhyAddrPointer_reg[31]/NET0131  & n36789 ;
  assign n36792 = ~n36790 & ~n36791 ;
  assign n36793 = ~n36760 & n36792 ;
  assign n36795 = ~\P2_P2_PhyAddrPointer_reg[31]/NET0131  & ~n36788 ;
  assign n36794 = \P2_P2_PhyAddrPointer_reg[31]/NET0131  & n36788 ;
  assign n36796 = n26800 & ~n36794 ;
  assign n36797 = ~n36795 & n36796 ;
  assign n36757 = ~n27614 & ~n27635 ;
  assign n36758 = ~n27612 & n36757 ;
  assign n36759 = \P2_P2_PhyAddrPointer_reg[31]/NET0131  & ~n36758 ;
  assign n36798 = ~n32856 & ~n36759 ;
  assign n36799 = ~n36797 & n36798 ;
  assign n36800 = ~n36793 & n36799 ;
  assign n36801 = ~n36756 & n36800 ;
  assign n36802 = \P1_P3_PhyAddrPointer_reg[31]/NET0131  & n9072 ;
  assign n36803 = ~n20356 & ~n36802 ;
  assign n36804 = n9064 & ~n36803 ;
  assign n36805 = ~n9050 & ~n9114 ;
  assign n36806 = \P1_P3_PhyAddrPointer_reg[31]/NET0131  & ~n36805 ;
  assign n36807 = ~n36804 & ~n36806 ;
  assign n36808 = ~n20373 & n36807 ;
  assign n36809 = n9241 & ~n36808 ;
  assign n36810 = ~n9246 & ~n16492 ;
  assign n36811 = n16484 & ~n36810 ;
  assign n36813 = \P1_P3_PhyAddrPointer_reg[31]/NET0131  & n16480 ;
  assign n36812 = ~\P1_P3_PhyAddrPointer_reg[31]/NET0131  & ~n16480 ;
  assign n36814 = n11698 & ~n36812 ;
  assign n36815 = ~n36813 & n36814 ;
  assign n36816 = ~n10036 & n16966 ;
  assign n36817 = \P1_P3_PhyAddrPointer_reg[31]/NET0131  & ~n36816 ;
  assign n36818 = ~n20381 & ~n36817 ;
  assign n36819 = ~n36815 & n36818 ;
  assign n36820 = ~n36811 & n36819 ;
  assign n36821 = ~n36809 & n36820 ;
  assign n36822 = n27283 & n33416 ;
  assign n36823 = ~\P2_P3_PhyAddrPointer_reg[31]/NET0131  & ~n27283 ;
  assign n36824 = n27117 & ~n36823 ;
  assign n36825 = ~n36822 & n36824 ;
  assign n36826 = ~n27118 & ~n27294 ;
  assign n36827 = \P2_P3_PhyAddrPointer_reg[31]/NET0131  & ~n36826 ;
  assign n36828 = ~n33505 & ~n36827 ;
  assign n36829 = ~n36825 & n36828 ;
  assign n36830 = n27308 & ~n36829 ;
  assign n36831 = ~n27316 & ~n32867 ;
  assign n36832 = \P2_P3_PhyAddrPointer_reg[21]/NET0131  & \P2_P3_PhyAddrPointer_reg[22]/NET0131  ;
  assign n36833 = \P2_P3_PhyAddrPointer_reg[23]/NET0131  & n36832 ;
  assign n36834 = \P2_P3_PhyAddrPointer_reg[24]/NET0131  & n36833 ;
  assign n36835 = \P2_P3_PhyAddrPointer_reg[2]/NET0131  & \P2_P3_PhyAddrPointer_reg[3]/NET0131  ;
  assign n36836 = \P2_P3_PhyAddrPointer_reg[4]/NET0131  & n36835 ;
  assign n36837 = \P2_P3_PhyAddrPointer_reg[5]/NET0131  & n36836 ;
  assign n36838 = \P2_P3_PhyAddrPointer_reg[6]/NET0131  & n36837 ;
  assign n36839 = \P2_P3_PhyAddrPointer_reg[7]/NET0131  & n36838 ;
  assign n36840 = \P2_P3_PhyAddrPointer_reg[8]/NET0131  & n36839 ;
  assign n36841 = \P2_P3_PhyAddrPointer_reg[9]/NET0131  & n36840 ;
  assign n36842 = \P2_P3_PhyAddrPointer_reg[10]/NET0131  & n36841 ;
  assign n36843 = \P2_P3_PhyAddrPointer_reg[11]/NET0131  & n36842 ;
  assign n36844 = \P2_P3_PhyAddrPointer_reg[12]/NET0131  & n36843 ;
  assign n36845 = \P2_P3_PhyAddrPointer_reg[13]/NET0131  & n36844 ;
  assign n36846 = \P2_P3_PhyAddrPointer_reg[14]/NET0131  & n36845 ;
  assign n36848 = \P2_P3_PhyAddrPointer_reg[16]/NET0131  & \P2_P3_PhyAddrPointer_reg[17]/NET0131  ;
  assign n36847 = \P2_P3_PhyAddrPointer_reg[15]/NET0131  & \P2_P3_PhyAddrPointer_reg[19]/NET0131  ;
  assign n36849 = \P2_P3_PhyAddrPointer_reg[18]/NET0131  & n36847 ;
  assign n36850 = n36848 & n36849 ;
  assign n36851 = \P2_P3_PhyAddrPointer_reg[20]/NET0131  & n36850 ;
  assign n36852 = n36846 & n36851 ;
  assign n36853 = n36834 & n36852 ;
  assign n36854 = \P2_P3_PhyAddrPointer_reg[25]/NET0131  & n36853 ;
  assign n36855 = \P2_P3_PhyAddrPointer_reg[26]/NET0131  & n36854 ;
  assign n36856 = \P2_P3_PhyAddrPointer_reg[27]/NET0131  & n36855 ;
  assign n36857 = \P2_P3_PhyAddrPointer_reg[1]/NET0131  & n36856 ;
  assign n36858 = \P2_P3_PhyAddrPointer_reg[28]/NET0131  & n36857 ;
  assign n36859 = \P2_P3_PhyAddrPointer_reg[29]/NET0131  & n36858 ;
  assign n36860 = \P2_P3_PhyAddrPointer_reg[30]/NET0131  & n36859 ;
  assign n36861 = \P2_P3_PhyAddrPointer_reg[31]/NET0131  & ~n36860 ;
  assign n36862 = ~\P2_P3_PhyAddrPointer_reg[31]/NET0131  & n36860 ;
  assign n36863 = ~n36861 & ~n36862 ;
  assign n36864 = ~n36831 & ~n36863 ;
  assign n36865 = \P2_P3_PhyAddrPointer_reg[28]/NET0131  & n36856 ;
  assign n36866 = \P2_P3_PhyAddrPointer_reg[29]/NET0131  & n36865 ;
  assign n36867 = \P2_P3_PhyAddrPointer_reg[30]/NET0131  & n36866 ;
  assign n36869 = \P2_P3_PhyAddrPointer_reg[31]/NET0131  & n36867 ;
  assign n36868 = ~\P2_P3_PhyAddrPointer_reg[31]/NET0131  & ~n36867 ;
  assign n36870 = n27325 & ~n36868 ;
  assign n36871 = ~n36869 & n36870 ;
  assign n36872 = ~n27310 & ~n27656 ;
  assign n36873 = ~n27650 & n36872 ;
  assign n36874 = \P2_P3_PhyAddrPointer_reg[31]/NET0131  & ~n36873 ;
  assign n36875 = ~n32865 & ~n36874 ;
  assign n36876 = ~n36871 & n36875 ;
  assign n36877 = ~n36864 & n36876 ;
  assign n36878 = ~n36830 & n36877 ;
  assign n36881 = \P1_P2_InstAddrPointer_reg[24]/NET0131  & n25733 ;
  assign n36889 = ~n31307 & ~n35082 ;
  assign n36888 = n31307 & n35082 ;
  assign n36890 = ~n30809 & ~n36888 ;
  assign n36891 = ~n36889 & n36890 ;
  assign n36882 = n30816 & ~n31305 ;
  assign n36883 = ~\P1_P2_InstAddrPointer_reg[24]/NET0131  & ~n30816 ;
  assign n36884 = ~n36882 & ~n36883 ;
  assign n36885 = ~n35078 & ~n36884 ;
  assign n36886 = ~n31152 & ~n36885 ;
  assign n36887 = n30809 & ~n36886 ;
  assign n36892 = ~n25733 & ~n36887 ;
  assign n36893 = ~n36891 & n36892 ;
  assign n36894 = ~n36881 & ~n36893 ;
  assign n36895 = n25701 & ~n36894 ;
  assign n36906 = ~n31441 & ~n35183 ;
  assign n36907 = n25881 & ~n35184 ;
  assign n36908 = ~n36906 & n36907 ;
  assign n36897 = n25770 & ~n25826 ;
  assign n36898 = n34206 & ~n36897 ;
  assign n36899 = ~n25748 & n36898 ;
  assign n36900 = ~n25847 & ~n25875 ;
  assign n36901 = n25415 & ~n36900 ;
  assign n36902 = n36899 & ~n36901 ;
  assign n36903 = \P1_P2_InstAddrPointer_reg[24]/NET0131  & ~n36902 ;
  assign n36896 = ~n25817 & ~n31307 ;
  assign n36904 = ~n25830 & n36884 ;
  assign n36905 = n25887 & n31441 ;
  assign n36909 = ~n36904 & ~n36905 ;
  assign n36910 = ~n36896 & n36909 ;
  assign n36911 = ~n36903 & n36910 ;
  assign n36912 = ~n36908 & n36911 ;
  assign n36913 = ~n36895 & n36912 ;
  assign n36914 = n25918 & ~n36913 ;
  assign n36879 = \P1_P2_InstAddrPointer_reg[24]/NET0131  & ~n31487 ;
  assign n36880 = \P1_P2_rEIP_reg[24]/NET0131  & n27967 ;
  assign n36915 = ~n36879 & ~n36880 ;
  assign n36916 = ~n36914 & n36915 ;
  assign n36919 = \P2_P1_InstAddrPointer_reg[15]/NET0131  & n25947 ;
  assign n36923 = n31944 & ~n31950 ;
  assign n36924 = ~n31948 & n36923 ;
  assign n36926 = n31956 & ~n36924 ;
  assign n36925 = ~n31956 & n36924 ;
  assign n36927 = ~n29503 & ~n36925 ;
  assign n36928 = ~n36926 & n36927 ;
  assign n36920 = ~n31814 & n31818 ;
  assign n36921 = ~n31819 & ~n36920 ;
  assign n36922 = n29503 & ~n36921 ;
  assign n36929 = ~n25947 & ~n36922 ;
  assign n36930 = ~n36928 & n36929 ;
  assign n36931 = ~n36919 & ~n36930 ;
  assign n36932 = n25945 & ~n36931 ;
  assign n36933 = \P2_P1_InstAddrPointer_reg[14]/NET0131  & n32106 ;
  assign n36935 = ~\P2_P1_InstAddrPointer_reg[15]/NET0131  & ~n32109 ;
  assign n36936 = \P2_P1_InstAddrPointer_reg[15]/NET0131  & n32109 ;
  assign n36937 = ~n36935 & ~n36936 ;
  assign n36938 = ~n36933 & ~n36937 ;
  assign n36934 = \P2_P1_InstAddrPointer_reg[15]/NET0131  & n36933 ;
  assign n36939 = n25964 & ~n36934 ;
  assign n36940 = ~n36938 & n36939 ;
  assign n36918 = ~n31818 & ~n32159 ;
  assign n36944 = n26068 & n36937 ;
  assign n36946 = ~n36918 & ~n36944 ;
  assign n36941 = ~n25987 & ~n32109 ;
  assign n36942 = n35385 & ~n36941 ;
  assign n36943 = \P2_P1_InstAddrPointer_reg[15]/NET0131  & ~n36942 ;
  assign n36945 = ~n25995 & n31956 ;
  assign n36947 = ~n36943 & ~n36945 ;
  assign n36948 = n36946 & n36947 ;
  assign n36949 = ~n36940 & n36948 ;
  assign n36950 = ~n36932 & n36949 ;
  assign n36951 = n11623 & ~n36950 ;
  assign n36917 = \P2_P1_rEIP_reg[15]/NET0131  & n11616 ;
  assign n36952 = \P2_P1_InstAddrPointer_reg[15]/NET0131  & ~n32172 ;
  assign n36953 = ~n36917 & ~n36952 ;
  assign n36954 = ~n36951 & n36953 ;
  assign n36959 = \P2_P1_InstAddrPointer_reg[19]/NET0131  & n25947 ;
  assign n36956 = ~\P2_P1_InstAddrPointer_reg[19]/NET0131  & n31834 ;
  assign n36957 = ~n31835 & ~n36956 ;
  assign n36966 = \P2_P1_InstAddrPointer_reg[18]/NET0131  & n31826 ;
  assign n36967 = n36957 & ~n36966 ;
  assign n36968 = n31826 & n31837 ;
  assign n36969 = ~n36967 & ~n36968 ;
  assign n36970 = n29503 & ~n36969 ;
  assign n36960 = n31960 & n31968 ;
  assign n36961 = ~n31975 & n36960 ;
  assign n36963 = n31972 & ~n36961 ;
  assign n36962 = ~n31972 & n36961 ;
  assign n36964 = ~n29503 & ~n36962 ;
  assign n36965 = ~n36963 & n36964 ;
  assign n36971 = ~n25947 & ~n36965 ;
  assign n36972 = ~n36970 & n36971 ;
  assign n36973 = ~n36959 & ~n36972 ;
  assign n36974 = n25945 & ~n36973 ;
  assign n36975 = ~\P2_P1_InstAddrPointer_reg[19]/NET0131  & ~n32119 ;
  assign n36976 = ~n32121 & ~n36975 ;
  assign n36977 = \P2_P1_InstAddrPointer_reg[18]/NET0131  & n32117 ;
  assign n36979 = ~n36976 & ~n36977 ;
  assign n36978 = n36976 & n36977 ;
  assign n36980 = n25964 & ~n36978 ;
  assign n36981 = ~n36979 & n36980 ;
  assign n36984 = ~n25995 & n31972 ;
  assign n36958 = ~n32159 & ~n36957 ;
  assign n36982 = \P2_P1_InstAddrPointer_reg[19]/NET0131  & ~n35385 ;
  assign n36983 = n26068 & n36976 ;
  assign n36985 = ~n36982 & ~n36983 ;
  assign n36986 = ~n36958 & n36985 ;
  assign n36987 = ~n36984 & n36986 ;
  assign n36988 = ~n36981 & n36987 ;
  assign n36989 = ~n36974 & n36988 ;
  assign n36990 = n11623 & ~n36989 ;
  assign n36955 = \P2_P1_rEIP_reg[19]/NET0131  & n11616 ;
  assign n36991 = \P2_P1_InstAddrPointer_reg[19]/NET0131  & ~n32172 ;
  assign n36992 = ~n36955 & ~n36991 ;
  assign n36993 = ~n36990 & n36992 ;
  assign n36996 = \P2_P1_InstAddrPointer_reg[20]/NET0131  & n25947 ;
  assign n37001 = ~n31833 & ~n36968 ;
  assign n37002 = ~n31839 & ~n37001 ;
  assign n37003 = n29503 & ~n37002 ;
  assign n36997 = n31978 & ~n36962 ;
  assign n36998 = n31980 & n36960 ;
  assign n36999 = ~n29503 & ~n36998 ;
  assign n37000 = ~n36997 & n36999 ;
  assign n37004 = ~n25947 & ~n37000 ;
  assign n37005 = ~n37003 & n37004 ;
  assign n37006 = ~n36996 & ~n37005 ;
  assign n37007 = n25945 & ~n37006 ;
  assign n37008 = ~n32124 & ~n36978 ;
  assign n37009 = n25964 & ~n32127 ;
  assign n37010 = ~n37008 & n37009 ;
  assign n37011 = n25949 & ~n31830 ;
  assign n37012 = n32159 & ~n37011 ;
  assign n37013 = n31833 & ~n37012 ;
  assign n36995 = ~n25995 & n31978 ;
  assign n37014 = n26068 & n32124 ;
  assign n37015 = \P2_P1_InstAddrPointer_reg[20]/NET0131  & ~n35385 ;
  assign n37016 = ~n37014 & ~n37015 ;
  assign n37017 = ~n36995 & n37016 ;
  assign n37018 = ~n37013 & n37017 ;
  assign n37019 = ~n37010 & n37018 ;
  assign n37020 = ~n37007 & n37019 ;
  assign n37021 = n11623 & ~n37020 ;
  assign n36994 = \P2_P1_rEIP_reg[20]/NET0131  & n11616 ;
  assign n37022 = \P2_P1_InstAddrPointer_reg[20]/NET0131  & ~n32172 ;
  assign n37023 = ~n36994 & ~n37022 ;
  assign n37024 = ~n37021 & n37023 ;
  assign n37027 = \P2_P1_InstAddrPointer_reg[22]/NET0131  & n25947 ;
  assign n37031 = ~n31840 & n31848 ;
  assign n37032 = ~n31849 & ~n37031 ;
  assign n37033 = n29503 & ~n37032 ;
  assign n37028 = ~n31885 & ~n31983 ;
  assign n37029 = ~n29503 & ~n35252 ;
  assign n37030 = ~n37028 & n37029 ;
  assign n37034 = ~n25947 & ~n37030 ;
  assign n37035 = ~n37033 & n37034 ;
  assign n37036 = ~n37027 & ~n37035 ;
  assign n37037 = n25945 & ~n37036 ;
  assign n37038 = ~n32130 & n32133 ;
  assign n37039 = n25964 & ~n35263 ;
  assign n37040 = ~n37038 & n37039 ;
  assign n37043 = ~n25995 & ~n31885 ;
  assign n37026 = ~n31848 & ~n32159 ;
  assign n37041 = \P2_P1_InstAddrPointer_reg[22]/NET0131  & ~n35385 ;
  assign n37042 = n26068 & ~n32133 ;
  assign n37044 = ~n37041 & ~n37042 ;
  assign n37045 = ~n37026 & n37044 ;
  assign n37046 = ~n37043 & n37045 ;
  assign n37047 = ~n37040 & n37046 ;
  assign n37048 = ~n37037 & n37047 ;
  assign n37049 = n11623 & ~n37048 ;
  assign n37025 = \P2_P1_rEIP_reg[22]/NET0131  & n11616 ;
  assign n37050 = \P2_P1_InstAddrPointer_reg[22]/NET0131  & ~n32172 ;
  assign n37051 = ~n37025 & ~n37050 ;
  assign n37052 = ~n37049 & n37051 ;
  assign n37055 = \P2_P1_InstAddrPointer_reg[24]/NET0131  & n25947 ;
  assign n37059 = ~\P2_P1_InstAddrPointer_reg[24]/NET0131  & ~n31514 ;
  assign n37060 = ~n31515 & ~n37059 ;
  assign n37061 = ~n31852 & ~n37060 ;
  assign n37062 = ~n31853 & ~n37061 ;
  assign n37063 = n29503 & ~n37062 ;
  assign n37056 = ~n31985 & n31988 ;
  assign n37057 = ~n29503 & ~n31989 ;
  assign n37058 = ~n37056 & n37057 ;
  assign n37064 = ~n25947 & ~n37058 ;
  assign n37065 = ~n37063 & n37064 ;
  assign n37066 = ~n37055 & ~n37065 ;
  assign n37067 = n25945 & ~n37066 ;
  assign n37068 = n32137 & ~n35264 ;
  assign n37069 = n25964 & ~n32142 ;
  assign n37070 = ~n37068 & n37069 ;
  assign n37071 = ~n32159 & n37060 ;
  assign n37054 = ~n25995 & n31988 ;
  assign n37072 = n26068 & ~n32137 ;
  assign n37073 = \P2_P1_InstAddrPointer_reg[24]/NET0131  & ~n35385 ;
  assign n37074 = ~n37072 & ~n37073 ;
  assign n37075 = ~n37054 & n37074 ;
  assign n37076 = ~n37071 & n37075 ;
  assign n37077 = ~n37070 & n37076 ;
  assign n37078 = ~n37067 & n37077 ;
  assign n37079 = n11623 & ~n37078 ;
  assign n37053 = \P2_P1_rEIP_reg[24]/NET0131  & n11616 ;
  assign n37080 = \P2_P1_InstAddrPointer_reg[24]/NET0131  & ~n32172 ;
  assign n37081 = ~n37053 & ~n37080 ;
  assign n37082 = ~n37079 & n37081 ;
  assign n37084 = \P2_P1_InstAddrPointer_reg[26]/NET0131  & n25947 ;
  assign n37088 = ~\P2_P1_InstAddrPointer_reg[26]/NET0131  & ~n31516 ;
  assign n37089 = ~n31517 & ~n37088 ;
  assign n37090 = \P2_P1_InstAddrPointer_reg[25]/NET0131  & n31853 ;
  assign n37091 = ~n37089 & ~n37090 ;
  assign n37092 = ~n31857 & ~n37091 ;
  assign n37093 = n29503 & ~n37092 ;
  assign n37085 = ~n31993 & n31996 ;
  assign n37086 = ~n29503 & ~n31997 ;
  assign n37087 = ~n37085 & n37086 ;
  assign n37094 = ~n25947 & ~n37087 ;
  assign n37095 = ~n37093 & n37094 ;
  assign n37096 = ~n37084 & ~n37095 ;
  assign n37097 = n25945 & ~n37096 ;
  assign n37098 = ~n32143 & ~n35363 ;
  assign n37099 = n25964 & ~n32144 ;
  assign n37100 = ~n37098 & n37099 ;
  assign n37101 = ~n32159 & n37089 ;
  assign n37083 = ~n25995 & n31996 ;
  assign n37102 = n26068 & n35363 ;
  assign n37103 = \P2_P1_InstAddrPointer_reg[26]/NET0131  & ~n35385 ;
  assign n37104 = ~n37102 & ~n37103 ;
  assign n37105 = ~n37083 & n37104 ;
  assign n37106 = ~n37101 & n37105 ;
  assign n37107 = ~n37100 & n37106 ;
  assign n37108 = ~n37097 & n37107 ;
  assign n37109 = n11623 & ~n37108 ;
  assign n37110 = \P2_P1_rEIP_reg[26]/NET0131  & n11616 ;
  assign n37111 = \P2_P1_InstAddrPointer_reg[26]/NET0131  & ~n32172 ;
  assign n37112 = ~n37110 & ~n37111 ;
  assign n37113 = ~n37109 & n37112 ;
  assign n37116 = \P2_P2_InstAddrPointer_reg[15]/NET0131  & n26629 ;
  assign n37117 = n32656 & ~n32659 ;
  assign n37118 = ~n32656 & n32659 ;
  assign n37119 = ~n37117 & ~n37118 ;
  assign n37120 = ~n32510 & ~n37119 ;
  assign n37121 = ~n32213 & ~n32521 ;
  assign n37122 = n32510 & ~n32522 ;
  assign n37123 = ~n37121 & n37122 ;
  assign n37124 = ~n37120 & ~n37123 ;
  assign n37125 = ~n26629 & ~n37124 ;
  assign n37126 = ~n37116 & ~n37125 ;
  assign n37127 = n26621 & ~n37126 ;
  assign n37128 = ~n32812 & ~n32814 ;
  assign n37129 = n26744 & ~n32815 ;
  assign n37130 = ~n37128 & n37129 ;
  assign n37133 = ~n26688 & n32659 ;
  assign n37132 = \P2_P2_InstAddrPointer_reg[15]/NET0131  & ~n35424 ;
  assign n37115 = ~n26764 & n32213 ;
  assign n37131 = n26757 & n32814 ;
  assign n37134 = ~n37115 & ~n37131 ;
  assign n37135 = ~n37132 & n37134 ;
  assign n37136 = ~n37133 & n37135 ;
  assign n37137 = ~n37130 & n37136 ;
  assign n37138 = ~n37127 & n37137 ;
  assign n37139 = n26792 & ~n37138 ;
  assign n37114 = \P2_P2_rEIP_reg[15]/NET0131  & n28046 ;
  assign n37140 = \P2_P2_InstAddrPointer_reg[15]/NET0131  & ~n32860 ;
  assign n37141 = ~n37114 & ~n37140 ;
  assign n37142 = ~n37139 & n37141 ;
  assign n37145 = \P2_P2_InstAddrPointer_reg[19]/NET0131  & n26629 ;
  assign n37150 = ~\P2_P2_InstAddrPointer_reg[19]/NET0131  & ~n32669 ;
  assign n37151 = ~n32529 & ~n37150 ;
  assign n37152 = n32522 & n32526 ;
  assign n37153 = ~n37151 & ~n37152 ;
  assign n37154 = ~n32528 & ~n37153 ;
  assign n37155 = n32510 & ~n37154 ;
  assign n37146 = n32668 & ~n32675 ;
  assign n37147 = n32673 & ~n37146 ;
  assign n37148 = ~n32510 & ~n32677 ;
  assign n37149 = ~n37147 & n37148 ;
  assign n37156 = ~n26629 & ~n37149 ;
  assign n37157 = ~n37155 & n37156 ;
  assign n37158 = ~n37145 & ~n37157 ;
  assign n37159 = n26621 & ~n37158 ;
  assign n37160 = ~n32818 & ~n32822 ;
  assign n37161 = n26744 & ~n32823 ;
  assign n37162 = ~n37160 & n37161 ;
  assign n37144 = ~n26688 & n32673 ;
  assign n37172 = ~n26764 & n37151 ;
  assign n37163 = n26757 & n32819 ;
  assign n37164 = ~\P2_P2_InstAddrPointer_reg[19]/NET0131  & ~n37163 ;
  assign n37165 = ~n26583 & n32822 ;
  assign n37166 = n32742 & ~n37165 ;
  assign n37167 = ~n37164 & ~n37166 ;
  assign n37168 = n26638 & n26640 ;
  assign n37169 = ~n26653 & ~n37168 ;
  assign n37170 = ~n26745 & n37169 ;
  assign n37171 = \P2_P2_InstAddrPointer_reg[19]/NET0131  & ~n37170 ;
  assign n37173 = ~n37167 & ~n37171 ;
  assign n37174 = ~n37172 & n37173 ;
  assign n37175 = ~n37144 & n37174 ;
  assign n37176 = ~n37162 & n37175 ;
  assign n37177 = ~n37159 & n37176 ;
  assign n37178 = n26792 & ~n37177 ;
  assign n37143 = \P2_P2_rEIP_reg[19]/NET0131  & n28046 ;
  assign n37179 = \P2_P2_InstAddrPointer_reg[19]/NET0131  & ~n32860 ;
  assign n37180 = ~n37143 & ~n37179 ;
  assign n37181 = ~n37178 & n37180 ;
  assign n37184 = \P2_P2_InstAddrPointer_reg[20]/NET0131  & n26629 ;
  assign n37188 = ~n32531 & ~n34286 ;
  assign n37189 = ~n34287 & ~n37188 ;
  assign n37190 = n32510 & ~n37189 ;
  assign n37185 = ~n32677 & n32689 ;
  assign n37186 = ~n32510 & ~n35409 ;
  assign n37187 = ~n37185 & n37186 ;
  assign n37191 = ~n26629 & ~n37187 ;
  assign n37192 = ~n37190 & n37191 ;
  assign n37193 = ~n37184 & ~n37192 ;
  assign n37194 = n26621 & ~n37193 ;
  assign n37195 = ~\P2_P2_InstAddrPointer_reg[20]/NET0131  & ~n32821 ;
  assign n37196 = ~n32725 & ~n37195 ;
  assign n37197 = ~n32823 & ~n37196 ;
  assign n37198 = n26744 & ~n32824 ;
  assign n37199 = ~n37197 & n37198 ;
  assign n37183 = ~n26688 & n32689 ;
  assign n37200 = \P2_P2_InstAddrPointer_reg[20]/NET0131  & ~n26679 ;
  assign n37201 = n26700 & ~n37200 ;
  assign n37203 = ~n26286 & n32531 ;
  assign n37202 = \P2_P2_InstAddrPointer_reg[20]/NET0131  & n26286 ;
  assign n37204 = ~n26640 & ~n37202 ;
  assign n37205 = ~n37203 & n37204 ;
  assign n37206 = ~n37201 & ~n37205 ;
  assign n37207 = \P2_P2_InstAddrPointer_reg[20]/NET0131  & ~n32744 ;
  assign n37208 = n26678 & n32531 ;
  assign n37209 = n26757 & n37196 ;
  assign n37210 = ~n37208 & ~n37209 ;
  assign n37211 = ~n37207 & n37210 ;
  assign n37212 = ~n37206 & n37211 ;
  assign n37213 = ~n37183 & n37212 ;
  assign n37214 = ~n37199 & n37213 ;
  assign n37215 = ~n37194 & n37214 ;
  assign n37216 = n26792 & ~n37215 ;
  assign n37182 = \P2_P2_rEIP_reg[20]/NET0131  & n28046 ;
  assign n37217 = \P2_P2_InstAddrPointer_reg[20]/NET0131  & ~n32860 ;
  assign n37218 = ~n37182 & ~n37217 ;
  assign n37219 = ~n37216 & n37218 ;
  assign n37225 = \P2_P2_InstAddrPointer_reg[22]/NET0131  & n26629 ;
  assign n37229 = n32541 & ~n34288 ;
  assign n37230 = ~n35405 & ~n37229 ;
  assign n37231 = n32510 & ~n37230 ;
  assign n37226 = ~n32680 & ~n35410 ;
  assign n37227 = ~n32510 & ~n35411 ;
  assign n37228 = ~n37226 & n37227 ;
  assign n37232 = ~n26629 & ~n37228 ;
  assign n37233 = ~n37231 & n37232 ;
  assign n37234 = ~n37225 & ~n37233 ;
  assign n37235 = n26621 & ~n37234 ;
  assign n37221 = \P2_P2_InstAddrPointer_reg[22]/NET0131  & ~n32722 ;
  assign n37222 = ~n32538 & n32722 ;
  assign n37223 = ~n37221 & ~n37222 ;
  assign n37236 = ~n32828 & n37223 ;
  assign n37237 = n26744 & ~n32829 ;
  assign n37238 = ~n37236 & n37237 ;
  assign n37243 = ~n26688 & ~n32680 ;
  assign n37239 = ~n26693 & n35449 ;
  assign n37240 = ~n26612 & n37239 ;
  assign n37241 = ~n26729 & n37240 ;
  assign n37242 = \P2_P2_InstAddrPointer_reg[22]/NET0131  & ~n37241 ;
  assign n37224 = n26757 & ~n37223 ;
  assign n37244 = ~n26764 & ~n32541 ;
  assign n37245 = ~n37224 & ~n37244 ;
  assign n37246 = ~n37242 & n37245 ;
  assign n37247 = ~n37243 & n37246 ;
  assign n37248 = ~n37238 & n37247 ;
  assign n37249 = ~n37235 & n37248 ;
  assign n37250 = n26792 & ~n37249 ;
  assign n37220 = \P2_P2_rEIP_reg[22]/NET0131  & n28046 ;
  assign n37251 = \P2_P2_InstAddrPointer_reg[22]/NET0131  & ~n32860 ;
  assign n37252 = ~n37220 & ~n37251 ;
  assign n37253 = ~n37250 & n37252 ;
  assign n37256 = \P2_P2_InstAddrPointer_reg[24]/NET0131  & n26629 ;
  assign n37260 = ~\P2_P2_InstAddrPointer_reg[24]/NET0131  & ~n32199 ;
  assign n37261 = ~n32200 & ~n37260 ;
  assign n37262 = ~n35406 & ~n37261 ;
  assign n37263 = ~n34289 & ~n37262 ;
  assign n37264 = n32510 & ~n37263 ;
  assign n37257 = n32578 & ~n32693 ;
  assign n37258 = ~n32510 & ~n32694 ;
  assign n37259 = ~n37257 & n37258 ;
  assign n37265 = ~n26629 & ~n37259 ;
  assign n37266 = ~n37264 & n37265 ;
  assign n37267 = ~n37256 & ~n37266 ;
  assign n37268 = n26621 & ~n37267 ;
  assign n37270 = \P2_P2_InstAddrPointer_reg[24]/NET0131  & n32830 ;
  assign n37269 = ~n32830 & ~n32833 ;
  assign n37271 = n26744 & ~n37269 ;
  assign n37272 = ~n37270 & n37271 ;
  assign n37273 = ~n26688 & n32578 ;
  assign n37274 = ~n26764 & n37261 ;
  assign n37255 = \P2_P2_InstAddrPointer_reg[24]/NET0131  & ~n35424 ;
  assign n37275 = n26757 & n32833 ;
  assign n37276 = ~n37255 & ~n37275 ;
  assign n37277 = ~n37274 & n37276 ;
  assign n37278 = ~n37273 & n37277 ;
  assign n37279 = ~n37272 & n37278 ;
  assign n37280 = ~n37268 & n37279 ;
  assign n37281 = n26792 & ~n37280 ;
  assign n37254 = \P2_P2_rEIP_reg[24]/NET0131  & n28046 ;
  assign n37282 = \P2_P2_InstAddrPointer_reg[24]/NET0131  & ~n32860 ;
  assign n37283 = ~n37254 & ~n37282 ;
  assign n37284 = ~n37281 & n37283 ;
  assign n37305 = ~n32835 & ~n32837 ;
  assign n37306 = n26744 & ~n32838 ;
  assign n37307 = ~n37305 & n37306 ;
  assign n37287 = \P2_P2_InstAddrPointer_reg[26]/NET0131  & n26629 ;
  assign n37291 = ~\P2_P2_InstAddrPointer_reg[26]/NET0131  & ~n32201 ;
  assign n37292 = ~n32202 & ~n37291 ;
  assign n37293 = ~n34290 & ~n37292 ;
  assign n37294 = ~n34291 & ~n37293 ;
  assign n37295 = n32510 & ~n37294 ;
  assign n37288 = ~n32695 & n32697 ;
  assign n37289 = ~n32510 & ~n32698 ;
  assign n37290 = ~n37288 & n37289 ;
  assign n37296 = ~n26629 & ~n37290 ;
  assign n37297 = ~n37295 & n37296 ;
  assign n37298 = ~n37287 & ~n37297 ;
  assign n37299 = n26621 & ~n37298 ;
  assign n37300 = ~n26688 & n32697 ;
  assign n37301 = ~n26583 & n32837 ;
  assign n37302 = n35424 & ~n37301 ;
  assign n37303 = \P2_P2_InstAddrPointer_reg[26]/NET0131  & ~n37302 ;
  assign n37304 = ~n26764 & n37292 ;
  assign n37308 = n26611 & n37301 ;
  assign n37309 = ~n37304 & ~n37308 ;
  assign n37310 = ~n37303 & n37309 ;
  assign n37311 = ~n37300 & n37310 ;
  assign n37312 = ~n37299 & n37311 ;
  assign n37313 = ~n37307 & n37312 ;
  assign n37314 = n26792 & ~n37313 ;
  assign n37285 = \P2_P2_rEIP_reg[26]/NET0131  & n28046 ;
  assign n37286 = \P2_P2_InstAddrPointer_reg[26]/NET0131  & ~n32860 ;
  assign n37315 = ~n37285 & ~n37286 ;
  assign n37316 = ~n37314 & n37315 ;
  assign n37319 = \P1_P2_InstAddrPointer_reg[26]/NET0131  & n25733 ;
  assign n37323 = ~n31310 & ~n31317 ;
  assign n37324 = ~n30809 & ~n35115 ;
  assign n37325 = ~n37323 & n37324 ;
  assign n37320 = ~n31155 & ~n31165 ;
  assign n37321 = ~n35110 & ~n37320 ;
  assign n37322 = n30809 & ~n37321 ;
  assign n37326 = ~n25733 & ~n37322 ;
  assign n37327 = ~n37325 & n37326 ;
  assign n37328 = ~n37319 & ~n37327 ;
  assign n37329 = n25701 & ~n37328 ;
  assign n37330 = ~n31447 & ~n35126 ;
  assign n37331 = n25881 & ~n35127 ;
  assign n37332 = ~n37330 & n37331 ;
  assign n37337 = ~n25817 & ~n31317 ;
  assign n37333 = ~n25743 & ~n31352 ;
  assign n37334 = n35131 & ~n37333 ;
  assign n37335 = \P1_P2_InstAddrPointer_reg[26]/NET0131  & ~n37334 ;
  assign n37318 = ~n25830 & n31165 ;
  assign n37336 = n25887 & n31447 ;
  assign n37338 = ~n37318 & ~n37336 ;
  assign n37339 = ~n37335 & n37338 ;
  assign n37340 = ~n37337 & n37339 ;
  assign n37341 = ~n37332 & n37340 ;
  assign n37342 = ~n37329 & n37341 ;
  assign n37343 = n25918 & ~n37342 ;
  assign n37317 = \P1_P2_InstAddrPointer_reg[26]/NET0131  & ~n31487 ;
  assign n37344 = \P1_P2_rEIP_reg[26]/NET0131  & n27967 ;
  assign n37345 = ~n37317 & ~n37344 ;
  assign n37346 = ~n37343 & n37345 ;
  assign n37349 = \P2_P3_InstAddrPointer_reg[15]/NET0131  & ~n27283 ;
  assign n37354 = ~n32952 & ~n33255 ;
  assign n37355 = ~n33256 & ~n37354 ;
  assign n37356 = n33242 & ~n37355 ;
  assign n37350 = ~n33357 & n34330 ;
  assign n37351 = ~n33351 & n33357 ;
  assign n37352 = ~n33242 & ~n37351 ;
  assign n37353 = ~n37350 & n37352 ;
  assign n37357 = n27283 & ~n37353 ;
  assign n37358 = ~n37356 & n37357 ;
  assign n37359 = ~n37349 & ~n37358 ;
  assign n37360 = n27117 & ~n37359 ;
  assign n37361 = ~n33426 & ~n33481 ;
  assign n37362 = n27280 & ~n33482 ;
  assign n37363 = ~n37361 & n37362 ;
  assign n37366 = ~n27229 & n32952 ;
  assign n37348 = \P2_P3_InstAddrPointer_reg[15]/NET0131  & ~n35672 ;
  assign n37364 = ~n27142 & n33357 ;
  assign n37365 = n27219 & n33426 ;
  assign n37367 = ~n37364 & ~n37365 ;
  assign n37368 = ~n37348 & n37367 ;
  assign n37369 = ~n37366 & n37368 ;
  assign n37370 = ~n37363 & n37369 ;
  assign n37371 = ~n37360 & n37370 ;
  assign n37372 = n27308 & ~n37371 ;
  assign n37347 = \P2_P3_rEIP_reg[15]/NET0131  & n32864 ;
  assign n37373 = \P2_P3_InstAddrPointer_reg[15]/NET0131  & ~n32870 ;
  assign n37374 = ~n37347 & ~n37373 ;
  assign n37375 = ~n37372 & n37374 ;
  assign n37378 = \P2_P3_InstAddrPointer_reg[19]/NET0131  & ~n27283 ;
  assign n37379 = ~\P2_P3_InstAddrPointer_reg[19]/NET0131  & ~n33361 ;
  assign n37380 = ~n32922 & ~n37379 ;
  assign n37381 = ~\P2_P3_InstAddrPointer_reg[18]/NET0131  & ~n33360 ;
  assign n37382 = ~n33361 & ~n37381 ;
  assign n37383 = \P2_P3_InstAddrPointer_reg[16]/NET0131  & n33256 ;
  assign n37384 = \P2_P3_InstAddrPointer_reg[17]/NET0131  & n37383 ;
  assign n37385 = n37382 & n37384 ;
  assign n37386 = ~n37380 & ~n37385 ;
  assign n37387 = ~n33260 & ~n37386 ;
  assign n37388 = n33242 & ~n37387 ;
  assign n37389 = n33359 & n33377 ;
  assign n37391 = n33365 & ~n37389 ;
  assign n37390 = ~n33365 & n37389 ;
  assign n37392 = ~n33242 & ~n37390 ;
  assign n37393 = ~n37391 & n37392 ;
  assign n37394 = n27283 & ~n37393 ;
  assign n37395 = ~n37388 & n37394 ;
  assign n37396 = ~n37378 & ~n37395 ;
  assign n37397 = n27117 & ~n37396 ;
  assign n37398 = \P2_P3_InstAddrPointer_reg[18]/NET0131  & n33484 ;
  assign n37399 = ~\P2_P3_InstAddrPointer_reg[19]/NET0131  & ~n37398 ;
  assign n37400 = ~n32890 & ~n37399 ;
  assign n37401 = n33483 & n33486 ;
  assign n37402 = \P2_P3_InstAddrPointer_reg[18]/NET0131  & n37401 ;
  assign n37403 = ~n37400 & ~n37402 ;
  assign n37404 = n27280 & ~n33488 ;
  assign n37405 = ~n37403 & n37404 ;
  assign n37410 = ~n27142 & n33365 ;
  assign n37406 = ~\P2_P3_InstAddrPointer_reg[19]/NET0131  & ~n27206 ;
  assign n37407 = ~n27111 & ~n37406 ;
  assign n37408 = n37400 & n37407 ;
  assign n37377 = \P2_P3_InstAddrPointer_reg[19]/NET0131  & ~n34355 ;
  assign n37409 = ~n27229 & n37380 ;
  assign n37411 = ~n37377 & ~n37409 ;
  assign n37412 = ~n37408 & n37411 ;
  assign n37413 = ~n37410 & n37412 ;
  assign n37414 = ~n37405 & n37413 ;
  assign n37415 = ~n37397 & n37414 ;
  assign n37416 = n27308 & ~n37415 ;
  assign n37376 = \P2_P3_rEIP_reg[19]/NET0131  & n32864 ;
  assign n37417 = \P2_P3_InstAddrPointer_reg[19]/NET0131  & ~n32870 ;
  assign n37418 = ~n37376 & ~n37417 ;
  assign n37419 = ~n37416 & n37418 ;
  assign n37422 = \P2_P3_InstAddrPointer_reg[20]/NET0131  & ~n27283 ;
  assign n37427 = ~n33262 & ~n35559 ;
  assign n37428 = ~n35560 & ~n37427 ;
  assign n37429 = n33242 & ~n37428 ;
  assign n37424 = n33367 & ~n37390 ;
  assign n37423 = ~n33367 & n37390 ;
  assign n37425 = ~n33242 & ~n37423 ;
  assign n37426 = ~n37424 & n37425 ;
  assign n37430 = n27283 & ~n37426 ;
  assign n37431 = ~n37429 & n37430 ;
  assign n37432 = ~n37422 & ~n37431 ;
  assign n37433 = n27117 & ~n37432 ;
  assign n37434 = ~n33424 & ~n35661 ;
  assign n37435 = n27280 & ~n35662 ;
  assign n37436 = ~n37434 & n37435 ;
  assign n37421 = ~n27229 & n33262 ;
  assign n37437 = ~n27111 & ~n32890 ;
  assign n37438 = n34355 & ~n37437 ;
  assign n37439 = \P2_P3_InstAddrPointer_reg[20]/NET0131  & ~n37438 ;
  assign n37442 = ~n37421 & ~n37439 ;
  assign n37440 = n27219 & n33424 ;
  assign n37441 = ~n27142 & n33367 ;
  assign n37443 = ~n37440 & ~n37441 ;
  assign n37444 = n37442 & n37443 ;
  assign n37445 = ~n37436 & n37444 ;
  assign n37446 = ~n37433 & n37445 ;
  assign n37447 = n27308 & ~n37446 ;
  assign n37420 = \P2_P3_rEIP_reg[20]/NET0131  & n32864 ;
  assign n37448 = \P2_P3_InstAddrPointer_reg[20]/NET0131  & ~n32870 ;
  assign n37449 = ~n37420 & ~n37448 ;
  assign n37450 = ~n37447 & n37449 ;
  assign n37455 = \P2_P3_InstAddrPointer_reg[22]/NET0131  & ~n27283 ;
  assign n37452 = ~\P2_P3_InstAddrPointer_reg[22]/NET0131  & ~n33369 ;
  assign n37453 = ~n35547 & ~n37452 ;
  assign n37459 = ~n35551 & ~n37453 ;
  assign n37460 = ~n35552 & ~n37459 ;
  assign n37461 = n33242 & ~n37460 ;
  assign n37456 = n33383 & ~n34332 ;
  assign n37457 = ~n33242 & ~n34333 ;
  assign n37458 = ~n37456 & n37457 ;
  assign n37462 = n27283 & ~n37458 ;
  assign n37463 = ~n37461 & n37462 ;
  assign n37464 = ~n37455 & ~n37463 ;
  assign n37465 = n27117 & ~n37464 ;
  assign n37466 = ~n33490 & ~n35575 ;
  assign n37467 = n27280 & ~n35576 ;
  assign n37468 = ~n37466 & n37467 ;
  assign n37475 = ~n27142 & n33383 ;
  assign n37469 = ~n27206 & n33418 ;
  assign n37470 = ~n27111 & ~n37469 ;
  assign n37471 = n35575 & n37470 ;
  assign n37454 = ~n27229 & n37453 ;
  assign n37472 = ~n27180 & ~n33369 ;
  assign n37473 = n34355 & ~n37472 ;
  assign n37474 = \P2_P3_InstAddrPointer_reg[22]/NET0131  & ~n37473 ;
  assign n37476 = ~n37454 & ~n37474 ;
  assign n37477 = ~n37471 & n37476 ;
  assign n37478 = ~n37475 & n37477 ;
  assign n37479 = ~n37468 & n37478 ;
  assign n37480 = ~n37465 & n37479 ;
  assign n37481 = n27308 & ~n37480 ;
  assign n37451 = \P2_P3_rEIP_reg[22]/NET0131  & n32864 ;
  assign n37482 = \P2_P3_InstAddrPointer_reg[22]/NET0131  & ~n32870 ;
  assign n37483 = ~n37451 & ~n37482 ;
  assign n37484 = ~n37481 & n37483 ;
  assign n37487 = \P2_P3_InstAddrPointer_reg[24]/NET0131  & ~n27283 ;
  assign n37491 = n33388 & ~n34334 ;
  assign n37492 = ~n33242 & ~n34335 ;
  assign n37493 = ~n37491 & n37492 ;
  assign n37488 = ~n35561 & ~n35642 ;
  assign n37489 = ~n35643 & ~n37488 ;
  assign n37490 = n33242 & ~n37489 ;
  assign n37494 = n27283 & ~n37490 ;
  assign n37495 = ~n37493 & n37494 ;
  assign n37496 = ~n37487 & ~n37495 ;
  assign n37497 = n27117 & ~n37496 ;
  assign n37498 = ~n35654 & ~n35664 ;
  assign n37499 = n27280 & ~n35665 ;
  assign n37500 = ~n37498 & n37499 ;
  assign n37501 = n27219 & n35654 ;
  assign n37486 = ~n27142 & n33388 ;
  assign n37502 = \P2_P3_InstAddrPointer_reg[24]/NET0131  & ~n34355 ;
  assign n37503 = ~n27229 & n35642 ;
  assign n37504 = ~n37502 & ~n37503 ;
  assign n37505 = ~n37486 & n37504 ;
  assign n37506 = ~n37501 & n37505 ;
  assign n37507 = ~n37500 & n37506 ;
  assign n37508 = ~n37497 & n37507 ;
  assign n37509 = n27308 & ~n37508 ;
  assign n37485 = \P2_P3_rEIP_reg[24]/NET0131  & n32864 ;
  assign n37510 = \P2_P3_InstAddrPointer_reg[24]/NET0131  & ~n32870 ;
  assign n37511 = ~n37485 & ~n37510 ;
  assign n37512 = ~n37509 & n37511 ;
  assign n37515 = \P2_P3_InstAddrPointer_reg[26]/NET0131  & ~n27283 ;
  assign n37519 = ~\P2_P3_InstAddrPointer_reg[26]/NET0131  & ~n32925 ;
  assign n37520 = ~n35608 & ~n37519 ;
  assign n37521 = ~n35611 & ~n37520 ;
  assign n37522 = ~n35612 & ~n37521 ;
  assign n37523 = n33242 & ~n37522 ;
  assign n37516 = n33396 & ~n34336 ;
  assign n37517 = ~n33242 & ~n34337 ;
  assign n37518 = ~n37516 & n37517 ;
  assign n37524 = n27283 & ~n37518 ;
  assign n37525 = ~n37523 & n37524 ;
  assign n37526 = ~n37515 & ~n37525 ;
  assign n37527 = n27117 & ~n37526 ;
  assign n37528 = ~\P2_P3_InstAddrPointer_reg[26]/NET0131  & ~n32896 ;
  assign n37529 = ~n32897 & ~n37528 ;
  assign n37530 = ~n35620 & ~n37529 ;
  assign n37531 = n27280 & ~n35621 ;
  assign n37532 = ~n37530 & n37531 ;
  assign n37535 = n27219 & n37529 ;
  assign n37533 = ~n27142 & n33396 ;
  assign n37514 = \P2_P3_InstAddrPointer_reg[26]/NET0131  & ~n34355 ;
  assign n37534 = ~n27229 & n37520 ;
  assign n37536 = ~n37514 & ~n37534 ;
  assign n37537 = ~n37533 & n37536 ;
  assign n37538 = ~n37535 & n37537 ;
  assign n37539 = ~n37532 & n37538 ;
  assign n37540 = ~n37527 & n37539 ;
  assign n37541 = n27308 & ~n37540 ;
  assign n37513 = \P2_P3_rEIP_reg[26]/NET0131  & n32864 ;
  assign n37542 = \P2_P3_InstAddrPointer_reg[26]/NET0131  & ~n32870 ;
  assign n37543 = ~n37513 & ~n37542 ;
  assign n37544 = ~n37541 & n37543 ;
  assign n37547 = \P1_P1_InstAddrPointer_reg[15]/NET0131  & n26249 ;
  assign n37551 = n33886 & ~n33958 ;
  assign n37552 = ~n29558 & ~n33959 ;
  assign n37553 = ~n37551 & n37552 ;
  assign n37548 = ~n33549 & ~n33820 ;
  assign n37549 = ~n33821 & ~n37548 ;
  assign n37550 = n29558 & ~n37549 ;
  assign n37554 = ~n26249 & ~n37550 ;
  assign n37555 = ~n37553 & n37554 ;
  assign n37556 = ~n37547 & ~n37555 ;
  assign n37557 = n26126 & ~n37556 ;
  assign n37558 = ~n34047 & ~n34101 ;
  assign n37559 = n26263 & ~n34102 ;
  assign n37560 = ~n37558 & n37559 ;
  assign n37563 = \P1_P1_InstAddrPointer_reg[15]/NET0131  & ~n34390 ;
  assign n37562 = ~n26189 & n33549 ;
  assign n37546 = ~n26151 & n33886 ;
  assign n37561 = n26192 & n34047 ;
  assign n37564 = ~n37546 & ~n37561 ;
  assign n37565 = ~n37562 & n37564 ;
  assign n37566 = ~n37563 & n37565 ;
  assign n37567 = ~n37560 & n37566 ;
  assign n37568 = ~n37557 & n37567 ;
  assign n37569 = n8355 & ~n37568 ;
  assign n37545 = \P1_P1_rEIP_reg[15]/NET0131  & n8357 ;
  assign n37570 = \P1_P1_InstAddrPointer_reg[15]/NET0131  & ~n34164 ;
  assign n37571 = ~n37545 & ~n37570 ;
  assign n37572 = ~n37569 & n37571 ;
  assign n37578 = \P1_P1_InstAddrPointer_reg[19]/NET0131  & n26249 ;
  assign n37586 = n33963 & ~n33973 ;
  assign n37588 = n33971 & ~n37586 ;
  assign n37587 = ~n33971 & n37586 ;
  assign n37589 = ~n29558 & ~n37587 ;
  assign n37590 = ~n37588 & n37589 ;
  assign n37579 = ~\P1_P1_InstAddrPointer_reg[19]/NET0131  & ~n33968 ;
  assign n37580 = ~n33534 & ~n37579 ;
  assign n37581 = n33822 & n33825 ;
  assign n37582 = \P1_P1_InstAddrPointer_reg[18]/NET0131  & n37581 ;
  assign n37583 = ~n37580 & ~n37582 ;
  assign n37584 = ~n33827 & ~n37583 ;
  assign n37585 = n29558 & ~n37584 ;
  assign n37591 = ~n26249 & ~n37585 ;
  assign n37592 = ~n37590 & n37591 ;
  assign n37593 = ~n37578 & ~n37592 ;
  assign n37594 = n26126 & ~n37593 ;
  assign n37574 = \P1_P1_InstAddrPointer_reg[18]/NET0131  & n34104 ;
  assign n37575 = ~\P1_P1_InstAddrPointer_reg[19]/NET0131  & ~n37574 ;
  assign n37576 = ~n34034 & ~n37575 ;
  assign n37595 = \P1_P1_InstAddrPointer_reg[18]/NET0131  & n34107 ;
  assign n37596 = ~n37576 & ~n37595 ;
  assign n37597 = n26263 & ~n34108 ;
  assign n37598 = ~n37596 & n37597 ;
  assign n37577 = n26192 & n37576 ;
  assign n37605 = ~n26123 & ~n34034 ;
  assign n37606 = n35760 & ~n37605 ;
  assign n37607 = \P1_P1_InstAddrPointer_reg[19]/NET0131  & ~n37606 ;
  assign n37599 = ~n24342 & ~n26129 ;
  assign n37600 = ~\P1_P1_InstAddrPointer_reg[19]/NET0131  & ~n26254 ;
  assign n37601 = ~n26160 & ~n37600 ;
  assign n37602 = n37599 & ~n37601 ;
  assign n37603 = n37580 & ~n37602 ;
  assign n37604 = ~n26151 & n33971 ;
  assign n37608 = ~n37603 & ~n37604 ;
  assign n37609 = ~n37607 & n37608 ;
  assign n37610 = ~n37577 & n37609 ;
  assign n37611 = ~n37598 & n37610 ;
  assign n37612 = ~n37594 & n37611 ;
  assign n37613 = n8355 & ~n37612 ;
  assign n37573 = \P1_P1_rEIP_reg[19]/NET0131  & n8357 ;
  assign n37614 = \P1_P1_InstAddrPointer_reg[19]/NET0131  & ~n34164 ;
  assign n37615 = ~n37573 & ~n37614 ;
  assign n37616 = ~n37613 & n37615 ;
  assign n37619 = \P1_P1_InstAddrPointer_reg[20]/NET0131  & n26249 ;
  assign n37623 = n33975 & ~n37587 ;
  assign n37624 = n33963 & n33977 ;
  assign n37625 = ~n29558 & ~n37624 ;
  assign n37626 = ~n37623 & n37625 ;
  assign n37620 = ~n33829 & ~n35735 ;
  assign n37621 = ~n35736 & ~n37620 ;
  assign n37622 = n29558 & ~n37621 ;
  assign n37627 = ~n26249 & ~n37622 ;
  assign n37628 = ~n37626 & n37627 ;
  assign n37629 = ~n37619 & ~n37628 ;
  assign n37630 = n26126 & ~n37629 ;
  assign n37631 = ~n34045 & ~n35821 ;
  assign n37632 = n26263 & ~n35822 ;
  assign n37633 = ~n37631 & n37632 ;
  assign n37634 = n34390 & ~n37605 ;
  assign n37635 = \P1_P1_InstAddrPointer_reg[20]/NET0131  & ~n37634 ;
  assign n37618 = ~n26189 & n33829 ;
  assign n37636 = n26192 & n34045 ;
  assign n37637 = ~n26151 & n33975 ;
  assign n37638 = ~n37636 & ~n37637 ;
  assign n37639 = ~n37618 & n37638 ;
  assign n37640 = ~n37635 & n37639 ;
  assign n37641 = ~n37633 & n37640 ;
  assign n37642 = ~n37630 & n37641 ;
  assign n37643 = n8355 & ~n37642 ;
  assign n37617 = \P1_P1_rEIP_reg[20]/NET0131  & n8357 ;
  assign n37644 = \P1_P1_InstAddrPointer_reg[20]/NET0131  & ~n34164 ;
  assign n37645 = ~n37617 & ~n37644 ;
  assign n37646 = ~n37643 & n37645 ;
  assign n37649 = \P1_P1_InstAddrPointer_reg[22]/NET0131  & n26249 ;
  assign n37656 = n33873 & ~n33979 ;
  assign n37657 = ~n29558 & ~n35720 ;
  assign n37658 = ~n37656 & n37657 ;
  assign n37650 = \P1_P1_InstAddrPointer_reg[21]/NET0131  & n33830 ;
  assign n37651 = ~\P1_P1_InstAddrPointer_reg[22]/NET0131  & ~n33846 ;
  assign n37652 = ~n33536 & ~n37651 ;
  assign n37653 = ~n37650 & ~n37652 ;
  assign n37654 = ~n35724 & ~n37653 ;
  assign n37655 = n29558 & ~n37654 ;
  assign n37659 = ~n26249 & ~n37655 ;
  assign n37660 = ~n37658 & n37659 ;
  assign n37661 = ~n37649 & ~n37660 ;
  assign n37662 = n26126 & ~n37661 ;
  assign n37663 = ~n34110 & ~n34113 ;
  assign n37664 = n26263 & ~n34114 ;
  assign n37665 = ~n37663 & n37664 ;
  assign n37666 = n26192 & n34113 ;
  assign n37668 = ~n26189 & n37652 ;
  assign n37648 = \P1_P1_InstAddrPointer_reg[22]/NET0131  & ~n35760 ;
  assign n37667 = ~n26151 & n33873 ;
  assign n37669 = ~n37648 & ~n37667 ;
  assign n37670 = ~n37668 & n37669 ;
  assign n37671 = ~n37666 & n37670 ;
  assign n37672 = ~n37665 & n37671 ;
  assign n37673 = ~n37662 & n37672 ;
  assign n37674 = n8355 & ~n37673 ;
  assign n37647 = \P1_P1_rEIP_reg[22]/NET0131  & n8357 ;
  assign n37675 = \P1_P1_InstAddrPointer_reg[22]/NET0131  & ~n34164 ;
  assign n37676 = ~n37647 & ~n37675 ;
  assign n37677 = ~n37674 & n37676 ;
  assign n37680 = \P1_P2_InstAddrPointer_reg[22]/NET0131  & n25733 ;
  assign n37684 = ~n31291 & n31294 ;
  assign n37685 = ~n30809 & ~n31295 ;
  assign n37686 = ~n37684 & n37685 ;
  assign n37681 = ~n31143 & ~n31146 ;
  assign n37682 = ~n35076 & ~n37681 ;
  assign n37683 = n30809 & ~n37682 ;
  assign n37687 = ~n25733 & ~n37683 ;
  assign n37688 = ~n37686 & n37687 ;
  assign n37689 = ~n37680 & ~n37688 ;
  assign n37690 = n25701 & ~n37689 ;
  assign n37691 = ~n31432 & ~n31436 ;
  assign n37692 = n25881 & ~n31437 ;
  assign n37693 = ~n37691 & n37692 ;
  assign n37696 = ~n25817 & n31294 ;
  assign n37679 = ~n25830 & n31146 ;
  assign n37694 = \P1_P2_InstAddrPointer_reg[22]/NET0131  & ~n35131 ;
  assign n37695 = n25887 & n31436 ;
  assign n37697 = ~n37694 & ~n37695 ;
  assign n37698 = ~n37679 & n37697 ;
  assign n37699 = ~n37696 & n37698 ;
  assign n37700 = ~n37693 & n37699 ;
  assign n37701 = ~n37690 & n37700 ;
  assign n37702 = n25918 & ~n37701 ;
  assign n37678 = \P1_P2_rEIP_reg[22]/NET0131  & n27967 ;
  assign n37703 = \P1_P2_InstAddrPointer_reg[22]/NET0131  & ~n31487 ;
  assign n37704 = ~n37678 & ~n37703 ;
  assign n37705 = ~n37702 & n37704 ;
  assign n37708 = \P1_P1_InstAddrPointer_reg[24]/NET0131  & n26249 ;
  assign n37713 = n33981 & n33988 ;
  assign n37712 = ~n33981 & ~n33988 ;
  assign n37714 = ~n29558 & ~n37712 ;
  assign n37715 = ~n37713 & n37714 ;
  assign n37709 = n33845 & ~n35737 ;
  assign n37710 = ~n35801 & ~n37709 ;
  assign n37711 = n29558 & ~n37710 ;
  assign n37716 = ~n26249 & ~n37711 ;
  assign n37717 = ~n37715 & n37716 ;
  assign n37718 = ~n37708 & ~n37717 ;
  assign n37719 = n26126 & ~n37718 ;
  assign n37720 = ~n34120 & ~n35825 ;
  assign n37721 = n26263 & ~n35826 ;
  assign n37722 = ~n37720 & n37721 ;
  assign n37707 = \P1_P1_InstAddrPointer_reg[24]/NET0131  & ~n34390 ;
  assign n37725 = ~n26151 & ~n33988 ;
  assign n37726 = ~n37707 & ~n37725 ;
  assign n37723 = ~n26189 & ~n33845 ;
  assign n37724 = n26192 & n34120 ;
  assign n37727 = ~n37723 & ~n37724 ;
  assign n37728 = n37726 & n37727 ;
  assign n37729 = ~n37722 & n37728 ;
  assign n37730 = ~n37719 & n37729 ;
  assign n37731 = n8355 & ~n37730 ;
  assign n37706 = \P1_P1_rEIP_reg[24]/NET0131  & n8357 ;
  assign n37732 = \P1_P1_InstAddrPointer_reg[24]/NET0131  & ~n34164 ;
  assign n37733 = ~n37706 & ~n37732 ;
  assign n37734 = ~n37731 & n37733 ;
  assign n37750 = ~\P1_P1_InstAddrPointer_reg[26]/NET0131  & ~n34037 ;
  assign n37751 = ~n34038 & ~n37750 ;
  assign n37761 = ~n35781 & ~n37751 ;
  assign n37762 = n26263 & ~n35782 ;
  assign n37763 = ~n37761 & n37762 ;
  assign n37737 = \P1_P1_InstAddrPointer_reg[26]/NET0131  & n26249 ;
  assign n37743 = ~n33990 & n33996 ;
  assign n37744 = ~n29558 & ~n35763 ;
  assign n37745 = ~n37743 & n37744 ;
  assign n37738 = ~\P1_P1_InstAddrPointer_reg[26]/NET0131  & ~n33538 ;
  assign n37739 = ~n35767 & ~n37738 ;
  assign n37740 = ~n35770 & ~n37739 ;
  assign n37741 = ~n35771 & ~n37740 ;
  assign n37742 = n29558 & ~n37741 ;
  assign n37746 = ~n26249 & ~n37742 ;
  assign n37747 = ~n37745 & n37746 ;
  assign n37748 = ~n37737 & ~n37747 ;
  assign n37749 = n26126 & ~n37748 ;
  assign n37752 = ~n26123 & n37751 ;
  assign n37753 = n35760 & ~n37752 ;
  assign n37754 = n26192 & n34037 ;
  assign n37755 = ~\P1_P1_InstAddrPointer_reg[26]/NET0131  & ~n37754 ;
  assign n37756 = ~n37753 & ~n37755 ;
  assign n37757 = ~n26131 & ~n33538 ;
  assign n37758 = n26189 & ~n37757 ;
  assign n37759 = n37739 & ~n37758 ;
  assign n37760 = ~n26151 & n33996 ;
  assign n37764 = ~n37759 & ~n37760 ;
  assign n37765 = ~n37756 & n37764 ;
  assign n37766 = ~n37749 & n37765 ;
  assign n37767 = ~n37763 & n37766 ;
  assign n37768 = n8355 & ~n37767 ;
  assign n37735 = \P1_P1_rEIP_reg[26]/NET0131  & n8357 ;
  assign n37736 = \P1_P1_InstAddrPointer_reg[26]/NET0131  & ~n34164 ;
  assign n37769 = ~n37735 & ~n37736 ;
  assign n37770 = ~n37768 & n37769 ;
  assign n37773 = \P1_P2_InstAddrPointer_reg[15]/NET0131  & n25733 ;
  assign n37779 = ~n31268 & n31271 ;
  assign n37780 = ~n30809 & ~n31272 ;
  assign n37781 = ~n37779 & n37780 ;
  assign n37774 = ~\P1_P2_InstAddrPointer_reg[15]/NET0131  & ~n30844 ;
  assign n37775 = ~n31135 & ~n37774 ;
  assign n37776 = ~n31126 & ~n37775 ;
  assign n37777 = ~n31127 & ~n37776 ;
  assign n37778 = n30809 & ~n37777 ;
  assign n37782 = ~n25733 & ~n37778 ;
  assign n37783 = ~n37781 & n37782 ;
  assign n37784 = ~n37773 & ~n37783 ;
  assign n37785 = n25701 & ~n37784 ;
  assign n37786 = ~n31420 & ~n31422 ;
  assign n37787 = n25881 & ~n31423 ;
  assign n37788 = ~n37786 & n37787 ;
  assign n37789 = n25774 & ~n30844 ;
  assign n37790 = n34208 & ~n37789 ;
  assign n37791 = \P1_P2_InstAddrPointer_reg[15]/NET0131  & ~n37790 ;
  assign n37772 = ~n25817 & n31271 ;
  assign n37792 = ~\P1_P2_InstAddrPointer_reg[15]/NET0131  & n25415 ;
  assign n37793 = ~n25415 & ~n37775 ;
  assign n37794 = ~n37792 & ~n37793 ;
  assign n37795 = ~n36900 & n37794 ;
  assign n37796 = n25808 & n37775 ;
  assign n37797 = n25887 & n31422 ;
  assign n37798 = ~n37796 & ~n37797 ;
  assign n37799 = ~n37795 & n37798 ;
  assign n37800 = ~n37772 & n37799 ;
  assign n37801 = ~n37791 & n37800 ;
  assign n37802 = ~n37788 & n37801 ;
  assign n37803 = ~n37785 & n37802 ;
  assign n37804 = n25918 & ~n37803 ;
  assign n37771 = \P1_P2_rEIP_reg[15]/NET0131  & n27967 ;
  assign n37805 = \P1_P2_InstAddrPointer_reg[15]/NET0131  & ~n31487 ;
  assign n37806 = ~n37771 & ~n37805 ;
  assign n37807 = ~n37804 & n37806 ;
  assign n37810 = \P1_P2_InstAddrPointer_reg[19]/NET0131  & n25733 ;
  assign n37819 = n31275 & ~n31281 ;
  assign n37820 = ~n31286 & n37819 ;
  assign n37821 = n31284 & ~n37820 ;
  assign n37822 = n31287 & n37819 ;
  assign n37823 = ~n30809 & ~n37822 ;
  assign n37824 = ~n37821 & n37823 ;
  assign n37811 = n31127 & n31138 ;
  assign n37812 = ~\P1_P2_InstAddrPointer_reg[18]/NET0131  & ~n31131 ;
  assign n37813 = ~n31132 & ~n37812 ;
  assign n37814 = n37811 & n37813 ;
  assign n37815 = ~n31134 & ~n37814 ;
  assign n37816 = \P1_P2_InstAddrPointer_reg[19]/NET0131  & n37814 ;
  assign n37817 = ~n37815 & ~n37816 ;
  assign n37818 = n30809 & ~n37817 ;
  assign n37825 = ~n25733 & ~n37818 ;
  assign n37826 = ~n37824 & n37825 ;
  assign n37827 = ~n37810 & ~n37826 ;
  assign n37828 = n25701 & ~n37827 ;
  assign n37832 = \P1_P2_InstAddrPointer_reg[18]/NET0131  & n31425 ;
  assign n37833 = ~\P1_P2_InstAddrPointer_reg[19]/NET0131  & ~n37832 ;
  assign n37834 = ~n31360 & ~n37833 ;
  assign n37836 = ~n31429 & ~n37834 ;
  assign n37837 = n25881 & ~n31430 ;
  assign n37838 = ~n37836 & n37837 ;
  assign n37829 = ~n25817 & n31284 ;
  assign n37830 = ~n25830 & n31134 ;
  assign n37831 = \P1_P2_InstAddrPointer_reg[19]/NET0131  & ~n35131 ;
  assign n37835 = n25887 & n37834 ;
  assign n37839 = ~n37831 & ~n37835 ;
  assign n37840 = ~n37830 & n37839 ;
  assign n37841 = ~n37829 & n37840 ;
  assign n37842 = ~n37838 & n37841 ;
  assign n37843 = ~n37828 & n37842 ;
  assign n37844 = n25918 & ~n37843 ;
  assign n37808 = \P1_P2_InstAddrPointer_reg[19]/NET0131  & ~n31487 ;
  assign n37809 = \P1_P2_rEIP_reg[19]/NET0131  & n27967 ;
  assign n37845 = ~n37808 & ~n37809 ;
  assign n37846 = ~n37844 & n37845 ;
  assign n37849 = \P1_P2_InstAddrPointer_reg[20]/NET0131  & n25733 ;
  assign n37853 = n31278 & ~n37822 ;
  assign n37854 = ~n30809 & ~n31290 ;
  assign n37855 = ~n37853 & n37854 ;
  assign n37850 = ~n31130 & ~n37816 ;
  assign n37851 = ~n31142 & ~n37850 ;
  assign n37852 = n30809 & ~n37851 ;
  assign n37856 = ~n25733 & ~n37852 ;
  assign n37857 = ~n37855 & n37856 ;
  assign n37858 = ~n37849 & ~n37857 ;
  assign n37859 = n25701 & ~n37858 ;
  assign n37860 = ~n31363 & ~n35180 ;
  assign n37861 = n25881 & ~n35181 ;
  assign n37862 = ~n37860 & n37861 ;
  assign n37868 = ~n25817 & n31278 ;
  assign n37867 = ~n25830 & n31130 ;
  assign n37848 = n25887 & n31363 ;
  assign n37863 = ~n25743 & n31363 ;
  assign n37864 = n25753 & ~n37863 ;
  assign n37865 = ~n25789 & n37864 ;
  assign n37866 = \P1_P2_InstAddrPointer_reg[20]/NET0131  & ~n37865 ;
  assign n37869 = ~n37848 & ~n37866 ;
  assign n37870 = ~n37867 & n37869 ;
  assign n37871 = ~n37868 & n37870 ;
  assign n37872 = ~n37862 & n37871 ;
  assign n37873 = ~n37859 & n37872 ;
  assign n37874 = n25918 & ~n37873 ;
  assign n37847 = \P1_P2_rEIP_reg[20]/NET0131  & n27967 ;
  assign n37875 = \P1_P2_InstAddrPointer_reg[20]/NET0131  & ~n31487 ;
  assign n37876 = ~n37847 & ~n37875 ;
  assign n37877 = ~n37874 & n37876 ;
  assign n37878 = \P2_P1_lWord_reg[5]/NET0131  & ~n34408 ;
  assign n37879 = n21062 & n24249 ;
  assign n37880 = \P2_P1_EAX_reg[5]/NET0131  & n24899 ;
  assign n37881 = ~n37879 & ~n37880 ;
  assign n37882 = n11623 & ~n37881 ;
  assign n37883 = ~n37878 & ~n37882 ;
  assign n37884 = \P2_P1_lWord_reg[6]/NET0131  & ~n34408 ;
  assign n37885 = \P2_P1_EAX_reg[6]/NET0131  & n24899 ;
  assign n37886 = n21062 & n24298 ;
  assign n37887 = ~n37885 & ~n37886 ;
  assign n37888 = n11623 & ~n37887 ;
  assign n37889 = ~n37884 & ~n37888 ;
  assign n37890 = \P1_P1_EAX_reg[5]/NET0131  & n24502 ;
  assign n37891 = ~n7933 & n23946 ;
  assign n37892 = ~n37890 & ~n37891 ;
  assign n37893 = ~n15364 & ~n37892 ;
  assign n37894 = \P1_P1_lWord_reg[5]/NET0131  & ~n24506 ;
  assign n37895 = ~n37893 & ~n37894 ;
  assign n37896 = n8355 & ~n37895 ;
  assign n37897 = \P1_P1_lWord_reg[5]/NET0131  & ~n24515 ;
  assign n37898 = ~n37896 & ~n37897 ;
  assign n37899 = \P1_P1_EAX_reg[6]/NET0131  & n24502 ;
  assign n37900 = n7906 & n23946 ;
  assign n37901 = ~n37899 & ~n37900 ;
  assign n37902 = ~n15364 & ~n37901 ;
  assign n37903 = \P1_P1_lWord_reg[6]/NET0131  & ~n24506 ;
  assign n37904 = ~n37902 & ~n37903 ;
  assign n37905 = n8355 & ~n37904 ;
  assign n37906 = \P1_P1_lWord_reg[6]/NET0131  & ~n24515 ;
  assign n37907 = ~n37905 & ~n37906 ;
  assign n37908 = \P1_P2_PhyAddrPointer_reg[30]/NET0131  & n25733 ;
  assign n37909 = ~n34199 & ~n37908 ;
  assign n37910 = n25701 & ~n37909 ;
  assign n37911 = \P1_P2_PhyAddrPointer_reg[30]/NET0131  & ~n36590 ;
  assign n37912 = ~n34204 & ~n37911 ;
  assign n37913 = ~n37910 & n37912 ;
  assign n37914 = n25918 & ~n37913 ;
  assign n37921 = \P1_P2_PhyAddrPointer_reg[1]/NET0131  & n36623 ;
  assign n37922 = ~\P1_P2_PhyAddrPointer_reg[30]/NET0131  & ~n37921 ;
  assign n37923 = ~n36625 & ~n37922 ;
  assign n37924 = n27898 & n37923 ;
  assign n37915 = ~\P1_P2_DataWidth_reg[1]/NET0131  & ~\P1_P2_PhyAddrPointer_reg[1]/NET0131  ;
  assign n37916 = n36623 & ~n37915 ;
  assign n37918 = \P1_P2_PhyAddrPointer_reg[30]/NET0131  & n37916 ;
  assign n37917 = ~\P1_P2_PhyAddrPointer_reg[30]/NET0131  & ~n37916 ;
  assign n37919 = n25928 & ~n37917 ;
  assign n37920 = ~n37918 & n37919 ;
  assign n37925 = \P1_P2_PhyAddrPointer_reg[30]/NET0131  & ~n36595 ;
  assign n37926 = ~n34223 & ~n37925 ;
  assign n37927 = ~n37920 & n37926 ;
  assign n37928 = ~n37924 & n37927 ;
  assign n37929 = ~n37914 & n37928 ;
  assign n37930 = \P2_P1_PhyAddrPointer_reg[30]/NET0131  & n25947 ;
  assign n37931 = ~n34235 & ~n37930 ;
  assign n37932 = n25945 & ~n37931 ;
  assign n37933 = \P2_P1_PhyAddrPointer_reg[30]/NET0131  & ~n36677 ;
  assign n37934 = ~n34243 & ~n37933 ;
  assign n37935 = ~n37932 & n37934 ;
  assign n37936 = n11623 & ~n37935 ;
  assign n37940 = \P2_P1_PhyAddrPointer_reg[1]/NET0131  & n36666 ;
  assign n37941 = ~\P2_P1_PhyAddrPointer_reg[30]/NET0131  & ~n37940 ;
  assign n37942 = ~n36668 & ~n37941 ;
  assign n37943 = n36674 & n37942 ;
  assign n37937 = ~\P2_P1_PhyAddrPointer_reg[30]/NET0131  & ~n36666 ;
  assign n37938 = n27681 & ~n36667 ;
  assign n37939 = ~n37937 & n37938 ;
  assign n37944 = \P2_P1_PhyAddrPointer_reg[30]/NET0131  & ~n36687 ;
  assign n37945 = ~n34257 & ~n37944 ;
  assign n37946 = ~n37939 & n37945 ;
  assign n37947 = ~n37943 & n37946 ;
  assign n37948 = ~n37936 & n37947 ;
  assign n37949 = \P1_P1_PhyAddrPointer_reg[30]/NET0131  & n26249 ;
  assign n37950 = ~n34381 & ~n37949 ;
  assign n37951 = n26126 & ~n37950 ;
  assign n37952 = \P1_P1_PhyAddrPointer_reg[30]/NET0131  & ~n36696 ;
  assign n37953 = ~n34386 & ~n37952 ;
  assign n37954 = ~n37951 & n37953 ;
  assign n37955 = n8355 & ~n37954 ;
  assign n37959 = ~\P1_P1_PhyAddrPointer_reg[30]/NET0131  & ~n36729 ;
  assign n37960 = ~n36730 & ~n37959 ;
  assign n37961 = ~n36701 & n37960 ;
  assign n37956 = ~\P1_P1_PhyAddrPointer_reg[30]/NET0131  & ~n36736 ;
  assign n37957 = n27791 & ~n36737 ;
  assign n37958 = ~n37956 & n37957 ;
  assign n37962 = \P1_P1_PhyAddrPointer_reg[30]/NET0131  & ~n36743 ;
  assign n37963 = ~n34401 & ~n37962 ;
  assign n37964 = ~n37958 & n37963 ;
  assign n37965 = ~n37961 & n37964 ;
  assign n37966 = ~n37955 & n37965 ;
  assign n37967 = \P2_P2_PhyAddrPointer_reg[30]/NET0131  & n26629 ;
  assign n37968 = ~n34299 & ~n37967 ;
  assign n37969 = n26621 & ~n37968 ;
  assign n37970 = \P2_P2_PhyAddrPointer_reg[30]/NET0131  & ~n36752 ;
  assign n37971 = ~n34304 & ~n37970 ;
  assign n37972 = ~n37969 & n37971 ;
  assign n37973 = n26792 & ~n37972 ;
  assign n37979 = ~\P2_P2_DataWidth_reg[1]/NET0131  & ~\P2_P2_PhyAddrPointer_reg[1]/NET0131  ;
  assign n37980 = n36786 & ~n37979 ;
  assign n37981 = \P2_P2_PhyAddrPointer_reg[29]/NET0131  & n37980 ;
  assign n37983 = \P2_P2_PhyAddrPointer_reg[30]/NET0131  & n37981 ;
  assign n37982 = ~\P2_P2_PhyAddrPointer_reg[30]/NET0131  & ~n37981 ;
  assign n37984 = n26794 & ~n37982 ;
  assign n37985 = ~n37983 & n37984 ;
  assign n37974 = \P2_P2_PhyAddrPointer_reg[1]/NET0131  & n36786 ;
  assign n37975 = \P2_P2_PhyAddrPointer_reg[29]/NET0131  & n37974 ;
  assign n37976 = ~\P2_P2_PhyAddrPointer_reg[30]/NET0131  & ~n37975 ;
  assign n37977 = ~n36789 & ~n37976 ;
  assign n37978 = n27977 & n37977 ;
  assign n37986 = \P2_P2_PhyAddrPointer_reg[30]/NET0131  & ~n36758 ;
  assign n37987 = ~n34262 & ~n37986 ;
  assign n37988 = ~n37978 & n37987 ;
  assign n37989 = ~n37985 & n37988 ;
  assign n37990 = ~n37973 & n37989 ;
  assign n37992 = ~n9073 & n36805 ;
  assign n37993 = \P1_P3_PhyAddrPointer_reg[30]/NET0131  & ~n37992 ;
  assign n37994 = ~n20327 & ~n37993 ;
  assign n37995 = ~n20317 & n37994 ;
  assign n37996 = n9241 & ~n37995 ;
  assign n37997 = ~\P1_P3_PhyAddrPointer_reg[30]/NET0131  & ~n16479 ;
  assign n37998 = ~n16480 & ~n37997 ;
  assign n37999 = \P1_P3_DataWidth_reg[1]/NET0131  & ~n37998 ;
  assign n38000 = n9245 & ~n37999 ;
  assign n38001 = ~n18330 & n38000 ;
  assign n37991 = n16492 & n18300 ;
  assign n38002 = \P1_P3_PhyAddrPointer_reg[30]/NET0131  & ~n36816 ;
  assign n38003 = ~n20299 & ~n38002 ;
  assign n38004 = ~n37991 & n38003 ;
  assign n38005 = ~n38001 & n38004 ;
  assign n38006 = ~n37996 & n38005 ;
  assign n38007 = \P2_P3_PhyAddrPointer_reg[30]/NET0131  & ~n27283 ;
  assign n38008 = ~n34345 & ~n38007 ;
  assign n38009 = n27117 & ~n38008 ;
  assign n38010 = \P2_P3_PhyAddrPointer_reg[30]/NET0131  & ~n36826 ;
  assign n38011 = ~n34353 & ~n38010 ;
  assign n38012 = ~n38009 & n38011 ;
  assign n38013 = n27308 & ~n38012 ;
  assign n38017 = ~\P2_P3_PhyAddrPointer_reg[30]/NET0131  & ~n36859 ;
  assign n38018 = ~n36860 & ~n38017 ;
  assign n38019 = ~n36831 & n38018 ;
  assign n38014 = ~\P2_P3_PhyAddrPointer_reg[30]/NET0131  & ~n36866 ;
  assign n38015 = n27325 & ~n36867 ;
  assign n38016 = ~n38014 & n38015 ;
  assign n38020 = \P2_P3_PhyAddrPointer_reg[30]/NET0131  & ~n36873 ;
  assign n38021 = ~n34369 & ~n38020 ;
  assign n38022 = ~n38016 & n38021 ;
  assign n38023 = ~n38019 & n38022 ;
  assign n38024 = ~n38013 & n38023 ;
  assign n38026 = \P1_P2_InstAddrPointer_reg[25]/NET0131  & n25733 ;
  assign n38030 = n31300 & ~n36888 ;
  assign n38031 = ~n30809 & ~n31310 ;
  assign n38032 = ~n38030 & n38031 ;
  assign n38027 = ~n31154 & ~n35210 ;
  assign n38028 = ~n35211 & ~n38027 ;
  assign n38029 = n30809 & ~n38028 ;
  assign n38033 = ~n25733 & ~n38029 ;
  assign n38034 = ~n38032 & n38033 ;
  assign n38035 = ~n38026 & ~n38034 ;
  assign n38036 = n25701 & ~n38035 ;
  assign n38037 = ~n31442 & ~n31445 ;
  assign n38038 = n25881 & ~n35126 ;
  assign n38039 = ~n38037 & n38038 ;
  assign n38042 = ~n25817 & n31300 ;
  assign n38025 = \P1_P2_InstAddrPointer_reg[25]/NET0131  & ~n36902 ;
  assign n38040 = n25887 & n31445 ;
  assign n38041 = ~n25830 & n31154 ;
  assign n38043 = ~n38040 & ~n38041 ;
  assign n38044 = ~n38025 & n38043 ;
  assign n38045 = ~n38042 & n38044 ;
  assign n38046 = ~n38039 & n38045 ;
  assign n38047 = ~n38036 & n38046 ;
  assign n38048 = n25918 & ~n38047 ;
  assign n38049 = \P1_P2_InstAddrPointer_reg[25]/NET0131  & ~n31487 ;
  assign n38050 = \P1_P2_rEIP_reg[25]/NET0131  & n27967 ;
  assign n38051 = ~n38049 & ~n38050 ;
  assign n38052 = ~n38048 & n38051 ;
  assign n38057 = \P2_P1_InstAddrPointer_reg[11]/NET0131  & n25947 ;
  assign n38062 = ~n31937 & n31939 ;
  assign n38063 = ~n29503 & ~n31940 ;
  assign n38064 = ~n38062 & n38063 ;
  assign n38054 = ~\P2_P1_InstAddrPointer_reg[11]/NET0131  & ~n31501 ;
  assign n38055 = ~n31502 & ~n38054 ;
  assign n38058 = ~n31811 & ~n38055 ;
  assign n38059 = \P2_P1_InstAddrPointer_reg[11]/NET0131  & n31811 ;
  assign n38060 = ~n38058 & ~n38059 ;
  assign n38061 = n29503 & ~n38060 ;
  assign n38065 = ~n25947 & ~n38061 ;
  assign n38066 = ~n38064 & n38065 ;
  assign n38067 = ~n38057 & ~n38066 ;
  assign n38068 = n25945 & ~n38067 ;
  assign n38069 = ~n32057 & ~n32103 ;
  assign n38070 = n25964 & ~n32104 ;
  assign n38071 = ~n38069 & n38070 ;
  assign n38076 = ~n25995 & n31939 ;
  assign n38056 = ~n32159 & n38055 ;
  assign n38072 = ~\P2_P1_InstAddrPointer_reg[11]/NET0131  & ~n20720 ;
  assign n38073 = n32057 & ~n38072 ;
  assign n38074 = ~n25987 & n38073 ;
  assign n38075 = \P2_P1_InstAddrPointer_reg[11]/NET0131  & ~n35385 ;
  assign n38077 = ~n38074 & ~n38075 ;
  assign n38078 = ~n38056 & n38077 ;
  assign n38079 = ~n38076 & n38078 ;
  assign n38080 = ~n38071 & n38079 ;
  assign n38081 = ~n38068 & n38080 ;
  assign n38082 = n11623 & ~n38081 ;
  assign n38053 = \P2_P1_rEIP_reg[11]/NET0131  & n11616 ;
  assign n38083 = \P2_P1_InstAddrPointer_reg[11]/NET0131  & ~n32172 ;
  assign n38084 = ~n38053 & ~n38083 ;
  assign n38085 = ~n38082 & n38084 ;
  assign n38088 = \P2_P1_InstAddrPointer_reg[14]/NET0131  & n25947 ;
  assign n38094 = n31948 & ~n36923 ;
  assign n38095 = ~n29503 & ~n36924 ;
  assign n38096 = ~n38094 & n38095 ;
  assign n38089 = ~\P2_P1_InstAddrPointer_reg[14]/NET0131  & ~n31539 ;
  assign n38090 = ~n31815 & ~n38089 ;
  assign n38091 = ~n31813 & ~n38090 ;
  assign n38092 = ~n31814 & ~n38091 ;
  assign n38093 = n29503 & ~n38092 ;
  assign n38097 = ~n25947 & ~n38093 ;
  assign n38098 = ~n38096 & n38097 ;
  assign n38099 = ~n38088 & ~n38098 ;
  assign n38100 = n25945 & ~n38099 ;
  assign n38101 = ~n32106 & ~n32110 ;
  assign n38102 = n25964 & ~n36933 ;
  assign n38103 = ~n38101 & n38102 ;
  assign n38104 = ~n32159 & n38090 ;
  assign n38087 = ~n25995 & n31948 ;
  assign n38105 = n26068 & n32110 ;
  assign n38106 = \P2_P1_InstAddrPointer_reg[14]/NET0131  & ~n35385 ;
  assign n38107 = ~n38105 & ~n38106 ;
  assign n38108 = ~n38087 & n38107 ;
  assign n38109 = ~n38104 & n38108 ;
  assign n38110 = ~n38103 & n38109 ;
  assign n38111 = ~n38100 & n38110 ;
  assign n38112 = n11623 & ~n38111 ;
  assign n38086 = \P2_P1_rEIP_reg[14]/NET0131  & n11616 ;
  assign n38113 = \P2_P1_InstAddrPointer_reg[14]/NET0131  & ~n32172 ;
  assign n38114 = ~n38086 & ~n38113 ;
  assign n38115 = ~n38112 & n38114 ;
  assign n38121 = \P2_P1_InstAddrPointer_reg[16]/NET0131  & n25947 ;
  assign n38125 = ~n31953 & ~n36925 ;
  assign n38126 = ~n29503 & ~n31960 ;
  assign n38127 = ~n38125 & n38126 ;
  assign n38122 = ~n31819 & n31824 ;
  assign n38123 = ~n31825 & ~n38122 ;
  assign n38124 = n29503 & ~n38123 ;
  assign n38128 = ~n25947 & ~n38124 ;
  assign n38129 = ~n38127 & n38128 ;
  assign n38130 = ~n38121 & ~n38129 ;
  assign n38131 = n25945 & ~n38130 ;
  assign n38117 = \P2_P1_InstAddrPointer_reg[16]/NET0131  & ~n32055 ;
  assign n38118 = n31822 & n32055 ;
  assign n38119 = ~n38117 & ~n38118 ;
  assign n38132 = ~n36934 & n38119 ;
  assign n38133 = n25964 & ~n32112 ;
  assign n38134 = ~n38132 & n38133 ;
  assign n38136 = ~n25995 & ~n31953 ;
  assign n38135 = ~n31824 & ~n32159 ;
  assign n38120 = n26068 & ~n38119 ;
  assign n38137 = \P2_P1_InstAddrPointer_reg[16]/NET0131  & ~n35385 ;
  assign n38138 = ~n38120 & ~n38137 ;
  assign n38139 = ~n38135 & n38138 ;
  assign n38140 = ~n38136 & n38139 ;
  assign n38141 = ~n38134 & n38140 ;
  assign n38142 = ~n38131 & n38141 ;
  assign n38143 = n11623 & ~n38142 ;
  assign n38116 = \P2_P1_rEIP_reg[16]/NET0131  & n11616 ;
  assign n38144 = \P2_P1_InstAddrPointer_reg[16]/NET0131  & ~n32172 ;
  assign n38145 = ~n38116 & ~n38144 ;
  assign n38146 = ~n38143 & n38145 ;
  assign n38150 = \P2_P1_InstAddrPointer_reg[18]/NET0131  & n25947 ;
  assign n38148 = ~n31834 & ~n31836 ;
  assign n38154 = ~n31826 & ~n38148 ;
  assign n38155 = ~n36966 & ~n38154 ;
  assign n38156 = n29503 & ~n38155 ;
  assign n38151 = n31975 & ~n36960 ;
  assign n38152 = ~n29503 & ~n36961 ;
  assign n38153 = ~n38151 & n38152 ;
  assign n38157 = ~n25947 & ~n38153 ;
  assign n38158 = ~n38156 & n38157 ;
  assign n38159 = ~n38150 & ~n38158 ;
  assign n38160 = n25945 & ~n38159 ;
  assign n38161 = ~n32117 & ~n32120 ;
  assign n38162 = n25964 & ~n36977 ;
  assign n38163 = ~n38161 & n38162 ;
  assign n38166 = ~n25995 & n31975 ;
  assign n38149 = ~n32159 & n38148 ;
  assign n38164 = \P2_P1_InstAddrPointer_reg[18]/NET0131  & ~n35385 ;
  assign n38165 = n26068 & n32120 ;
  assign n38167 = ~n38164 & ~n38165 ;
  assign n38168 = ~n38149 & n38167 ;
  assign n38169 = ~n38166 & n38168 ;
  assign n38170 = ~n38163 & n38169 ;
  assign n38171 = ~n38160 & n38170 ;
  assign n38172 = n11623 & ~n38171 ;
  assign n38147 = \P2_P1_rEIP_reg[18]/NET0131  & n11616 ;
  assign n38173 = \P2_P1_InstAddrPointer_reg[18]/NET0131  & ~n32172 ;
  assign n38174 = ~n38147 & ~n38173 ;
  assign n38175 = ~n38172 & n38174 ;
  assign n38178 = \P2_P1_InstAddrPointer_reg[21]/NET0131  & n25947 ;
  assign n38182 = n31532 & ~n31839 ;
  assign n38183 = ~n31840 & ~n38182 ;
  assign n38184 = n29503 & ~n38183 ;
  assign n38179 = ~n31964 & ~n36998 ;
  assign n38180 = ~n29503 & ~n31983 ;
  assign n38181 = ~n38179 & n38180 ;
  assign n38185 = ~n25947 & ~n38181 ;
  assign n38186 = ~n38184 & n38185 ;
  assign n38187 = ~n38178 & ~n38186 ;
  assign n38188 = n25945 & ~n38187 ;
  assign n38189 = ~n32129 & ~n35371 ;
  assign n38190 = n25964 & ~n35372 ;
  assign n38191 = ~n38189 & n38190 ;
  assign n38194 = ~n25995 & ~n31964 ;
  assign n38177 = ~n31532 & ~n32159 ;
  assign n38192 = \P2_P1_InstAddrPointer_reg[21]/NET0131  & ~n35385 ;
  assign n38193 = n26068 & n32129 ;
  assign n38195 = ~n38192 & ~n38193 ;
  assign n38196 = ~n38177 & n38195 ;
  assign n38197 = ~n38194 & n38196 ;
  assign n38198 = ~n38191 & n38197 ;
  assign n38199 = ~n38188 & n38198 ;
  assign n38200 = n11623 & ~n38199 ;
  assign n38176 = \P2_P1_rEIP_reg[21]/NET0131  & n11616 ;
  assign n38201 = \P2_P1_InstAddrPointer_reg[21]/NET0131  & ~n32172 ;
  assign n38202 = ~n38176 & ~n38201 ;
  assign n38203 = ~n38200 & n38202 ;
  assign n38206 = \P2_P1_InstAddrPointer_reg[25]/NET0131  & n25947 ;
  assign n38210 = ~n31853 & ~n31855 ;
  assign n38211 = ~n37090 & ~n38210 ;
  assign n38212 = n29503 & ~n38211 ;
  assign n38207 = ~n31989 & n31992 ;
  assign n38208 = ~n29503 & ~n31993 ;
  assign n38209 = ~n38207 & n38208 ;
  assign n38213 = ~n25947 & ~n38209 ;
  assign n38214 = ~n38212 & n38213 ;
  assign n38215 = ~n38206 & ~n38214 ;
  assign n38216 = n25945 & ~n38215 ;
  assign n38217 = ~n32044 & ~n35373 ;
  assign n38218 = n25964 & ~n35374 ;
  assign n38219 = ~n38217 & n38218 ;
  assign n38222 = ~n25995 & n31992 ;
  assign n38205 = n31855 & ~n32159 ;
  assign n38220 = \P2_P1_InstAddrPointer_reg[25]/NET0131  & ~n35385 ;
  assign n38221 = n26068 & n32044 ;
  assign n38223 = ~n38220 & ~n38221 ;
  assign n38224 = ~n38205 & n38223 ;
  assign n38225 = ~n38222 & n38224 ;
  assign n38226 = ~n38219 & n38225 ;
  assign n38227 = ~n38216 & n38226 ;
  assign n38228 = n11623 & ~n38227 ;
  assign n38204 = \P2_P1_rEIP_reg[25]/NET0131  & n11616 ;
  assign n38229 = \P2_P1_InstAddrPointer_reg[25]/NET0131  & ~n32172 ;
  assign n38230 = ~n38204 & ~n38229 ;
  assign n38231 = ~n38228 & n38230 ;
  assign n38236 = \P2_P2_InstAddrPointer_reg[11]/NET0131  & n26629 ;
  assign n38233 = ~\P2_P2_InstAddrPointer_reg[11]/NET0131  & ~n32222 ;
  assign n38234 = ~n32579 & ~n38233 ;
  assign n38241 = ~n32518 & ~n38234 ;
  assign n38242 = ~n34281 & ~n38241 ;
  assign n38243 = n32510 & ~n38242 ;
  assign n38237 = n32640 & ~n32643 ;
  assign n38238 = n32645 & ~n38237 ;
  assign n38239 = ~n32510 & ~n32647 ;
  assign n38240 = ~n38238 & n38239 ;
  assign n38244 = ~n26629 & ~n38240 ;
  assign n38245 = ~n38243 & n38244 ;
  assign n38246 = ~n38236 & ~n38245 ;
  assign n38247 = n26621 & ~n38246 ;
  assign n38249 = \P2_P2_InstAddrPointer_reg[11]/NET0131  & n32762 ;
  assign n38250 = ~\P2_P2_InstAddrPointer_reg[11]/NET0131  & ~n32762 ;
  assign n38251 = ~n38249 & ~n38250 ;
  assign n38252 = ~n32806 & ~n38251 ;
  assign n38248 = \P2_P2_InstAddrPointer_reg[11]/NET0131  & n32806 ;
  assign n38253 = n26744 & ~n38248 ;
  assign n38254 = ~n38252 & n38253 ;
  assign n38259 = ~n26688 & n32645 ;
  assign n38255 = ~n26583 & ~n32762 ;
  assign n38256 = n35424 & ~n38255 ;
  assign n38257 = \P2_P2_InstAddrPointer_reg[11]/NET0131  & ~n38256 ;
  assign n38235 = ~n26764 & n38234 ;
  assign n38258 = n26757 & n38251 ;
  assign n38260 = ~n38235 & ~n38258 ;
  assign n38261 = ~n38257 & n38260 ;
  assign n38262 = ~n38259 & n38261 ;
  assign n38263 = ~n38254 & n38262 ;
  assign n38264 = ~n38247 & n38263 ;
  assign n38265 = n26792 & ~n38264 ;
  assign n38232 = \P2_P2_rEIP_reg[11]/NET0131  & n28046 ;
  assign n38266 = \P2_P2_InstAddrPointer_reg[11]/NET0131  & ~n32860 ;
  assign n38267 = ~n38232 & ~n38266 ;
  assign n38268 = ~n38265 & n38267 ;
  assign n38271 = \P2_P2_InstAddrPointer_reg[14]/NET0131  & n26629 ;
  assign n38276 = ~n34278 & ~n34283 ;
  assign n38277 = ~n34284 & ~n38276 ;
  assign n38278 = n32510 & ~n38277 ;
  assign n38272 = n32648 & ~n32654 ;
  assign n38273 = n32652 & ~n38272 ;
  assign n38274 = ~n32510 & ~n32656 ;
  assign n38275 = ~n38273 & n38274 ;
  assign n38279 = ~n26629 & ~n38275 ;
  assign n38280 = ~n38278 & n38279 ;
  assign n38281 = ~n38271 & ~n38280 ;
  assign n38282 = n26621 & ~n38281 ;
  assign n38283 = ~\P2_P2_InstAddrPointer_reg[14]/NET0131  & ~n32723 ;
  assign n38284 = ~n32724 & ~n38283 ;
  assign n38285 = ~n32811 & ~n38284 ;
  assign n38286 = n26744 & ~n32812 ;
  assign n38287 = ~n38285 & n38286 ;
  assign n38270 = ~n26688 & n32652 ;
  assign n38289 = n26697 & ~n32214 ;
  assign n38290 = n35423 & ~n38289 ;
  assign n38291 = \P2_P2_InstAddrPointer_reg[14]/NET0131  & ~n38290 ;
  assign n38288 = ~n26762 & n34278 ;
  assign n38292 = ~\P2_P2_InstAddrPointer_reg[14]/NET0131  & ~n26652 ;
  assign n38293 = n26652 & ~n34278 ;
  assign n38294 = ~n38292 & ~n38293 ;
  assign n38295 = ~n26645 & n38294 ;
  assign n38296 = ~\P2_P2_InstAddrPointer_reg[14]/NET0131  & ~n26611 ;
  assign n38297 = n26611 & ~n38284 ;
  assign n38298 = ~n38296 & ~n38297 ;
  assign n38299 = ~n26583 & n38298 ;
  assign n38300 = ~n38295 & ~n38299 ;
  assign n38301 = ~n38288 & n38300 ;
  assign n38302 = ~n38291 & n38301 ;
  assign n38303 = ~n38270 & n38302 ;
  assign n38304 = ~n38287 & n38303 ;
  assign n38305 = ~n38282 & n38304 ;
  assign n38306 = n26792 & ~n38305 ;
  assign n38269 = \P2_P2_rEIP_reg[14]/NET0131  & n28046 ;
  assign n38307 = \P2_P2_InstAddrPointer_reg[14]/NET0131  & ~n32860 ;
  assign n38308 = ~n38269 & ~n38307 ;
  assign n38309 = ~n38306 & n38308 ;
  assign n38312 = \P2_P2_InstAddrPointer_reg[16]/NET0131  & n26629 ;
  assign n38316 = ~n32525 & ~n34285 ;
  assign n38317 = n32525 & n34285 ;
  assign n38318 = ~n38316 & ~n38317 ;
  assign n38319 = n32510 & ~n38318 ;
  assign n38313 = n32662 & ~n37117 ;
  assign n38314 = ~n32510 & ~n32664 ;
  assign n38315 = ~n38313 & n38314 ;
  assign n38320 = ~n26629 & ~n38315 ;
  assign n38321 = ~n38319 & n38320 ;
  assign n38322 = ~n38312 & ~n38321 ;
  assign n38323 = n26621 & ~n38322 ;
  assign n38324 = ~\P2_P2_InstAddrPointer_reg[16]/NET0131  & ~n32752 ;
  assign n38325 = ~n32753 & ~n38324 ;
  assign n38326 = ~n32815 & ~n38325 ;
  assign n38327 = n26744 & ~n32816 ;
  assign n38328 = ~n38326 & n38327 ;
  assign n38333 = ~n26688 & n32662 ;
  assign n38329 = ~n26583 & ~n32752 ;
  assign n38330 = n35424 & ~n38329 ;
  assign n38331 = \P2_P2_InstAddrPointer_reg[16]/NET0131  & ~n38330 ;
  assign n38311 = ~n26764 & n32525 ;
  assign n38332 = n26757 & n38325 ;
  assign n38334 = ~n38311 & ~n38332 ;
  assign n38335 = ~n38331 & n38334 ;
  assign n38336 = ~n38333 & n38335 ;
  assign n38337 = ~n38328 & n38336 ;
  assign n38338 = ~n38323 & n38337 ;
  assign n38339 = n26792 & ~n38338 ;
  assign n38310 = \P2_P2_rEIP_reg[16]/NET0131  & n28046 ;
  assign n38340 = \P2_P2_InstAddrPointer_reg[16]/NET0131  & ~n32860 ;
  assign n38341 = ~n38310 & ~n38340 ;
  assign n38342 = ~n38339 & n38341 ;
  assign n38345 = \P2_P2_InstAddrPointer_reg[18]/NET0131  & n26629 ;
  assign n38349 = \P2_P2_InstAddrPointer_reg[17]/NET0131  & n32523 ;
  assign n38350 = ~\P2_P2_InstAddrPointer_reg[18]/NET0131  & ~n38349 ;
  assign n38351 = ~n32669 & ~n38350 ;
  assign n38352 = \P2_P2_InstAddrPointer_reg[17]/NET0131  & n38317 ;
  assign n38353 = ~n38351 & ~n38352 ;
  assign n38354 = n32179 & n38317 ;
  assign n38355 = ~n38353 & ~n38354 ;
  assign n38356 = n32510 & ~n38355 ;
  assign n38346 = ~n32668 & n32675 ;
  assign n38347 = ~n32510 & ~n37146 ;
  assign n38348 = ~n38346 & n38347 ;
  assign n38357 = ~n26629 & ~n38348 ;
  assign n38358 = ~n38356 & n38357 ;
  assign n38359 = ~n38345 & ~n38358 ;
  assign n38360 = n26621 & ~n38359 ;
  assign n38361 = ~\P2_P2_InstAddrPointer_reg[18]/NET0131  & ~n32754 ;
  assign n38362 = ~n32819 & ~n38361 ;
  assign n38363 = ~n32817 & ~n38362 ;
  assign n38364 = n26744 & ~n32818 ;
  assign n38365 = ~n38363 & n38364 ;
  assign n38366 = ~n26688 & n32675 ;
  assign n38367 = ~n26764 & n38351 ;
  assign n38344 = \P2_P2_InstAddrPointer_reg[18]/NET0131  & ~n35424 ;
  assign n38368 = n26757 & n38362 ;
  assign n38369 = ~n38344 & ~n38368 ;
  assign n38370 = ~n38367 & n38369 ;
  assign n38371 = ~n38366 & n38370 ;
  assign n38372 = ~n38365 & n38371 ;
  assign n38373 = ~n38360 & n38372 ;
  assign n38374 = n26792 & ~n38373 ;
  assign n38343 = \P2_P2_rEIP_reg[18]/NET0131  & n28046 ;
  assign n38375 = \P2_P2_InstAddrPointer_reg[18]/NET0131  & ~n32860 ;
  assign n38376 = ~n38343 & ~n38375 ;
  assign n38377 = ~n38374 & n38376 ;
  assign n38402 = ~n32824 & ~n32827 ;
  assign n38403 = n26744 & ~n32828 ;
  assign n38404 = ~n38402 & n38403 ;
  assign n38380 = \P2_P2_InstAddrPointer_reg[21]/NET0131  & n26629 ;
  assign n38384 = ~\P2_P2_InstAddrPointer_reg[21]/NET0131  & ~n32197 ;
  assign n38385 = n32187 & n32535 ;
  assign n38386 = ~n38384 & ~n38385 ;
  assign n38387 = ~n32532 & ~n38386 ;
  assign n38388 = ~n32533 & ~n38387 ;
  assign n38389 = n32510 & ~n38388 ;
  assign n38381 = ~n32687 & ~n35409 ;
  assign n38382 = ~n32510 & ~n35410 ;
  assign n38383 = ~n38381 & n38382 ;
  assign n38390 = ~n26629 & ~n38383 ;
  assign n38391 = ~n38389 & n38390 ;
  assign n38392 = ~n38380 & ~n38391 ;
  assign n38393 = n26621 & ~n38392 ;
  assign n38400 = ~n26688 & ~n32687 ;
  assign n38401 = ~n26764 & n38386 ;
  assign n38394 = n26757 & n32725 ;
  assign n38395 = ~\P2_P2_InstAddrPointer_reg[21]/NET0131  & ~n38394 ;
  assign n38396 = ~n26583 & n32827 ;
  assign n38397 = n32742 & ~n38396 ;
  assign n38398 = ~n38395 & ~n38397 ;
  assign n38399 = \P2_P2_InstAddrPointer_reg[21]/NET0131  & ~n37170 ;
  assign n38405 = ~n38398 & ~n38399 ;
  assign n38406 = ~n38401 & n38405 ;
  assign n38407 = ~n38400 & n38406 ;
  assign n38408 = ~n38393 & n38407 ;
  assign n38409 = ~n38404 & n38408 ;
  assign n38410 = n26792 & ~n38409 ;
  assign n38378 = \P2_P2_rEIP_reg[21]/NET0131  & n28046 ;
  assign n38379 = \P2_P2_InstAddrPointer_reg[21]/NET0131  & ~n32860 ;
  assign n38411 = ~n38378 & ~n38379 ;
  assign n38412 = ~n38410 & n38411 ;
  assign n38428 = ~\P2_P2_InstAddrPointer_reg[25]/NET0131  & ~n32832 ;
  assign n38429 = ~n32729 & ~n38428 ;
  assign n38432 = ~n37270 & ~n38429 ;
  assign n38433 = n26744 & ~n32835 ;
  assign n38434 = ~n38432 & n38433 ;
  assign n38415 = \P2_P2_InstAddrPointer_reg[25]/NET0131  & n26629 ;
  assign n38419 = ~n32546 & ~n32548 ;
  assign n38420 = ~n32549 & ~n38419 ;
  assign n38421 = n32510 & ~n38420 ;
  assign n38416 = n32575 & ~n32694 ;
  assign n38417 = ~n32510 & ~n32695 ;
  assign n38418 = ~n38416 & n38417 ;
  assign n38422 = ~n26629 & ~n38418 ;
  assign n38423 = ~n38421 & n38422 ;
  assign n38424 = ~n38415 & ~n38423 ;
  assign n38425 = n26621 & ~n38424 ;
  assign n38427 = \P2_P2_InstAddrPointer_reg[25]/NET0131  & ~n37241 ;
  assign n38426 = ~n26688 & n32575 ;
  assign n38430 = n26757 & n38429 ;
  assign n38431 = ~n26764 & n32548 ;
  assign n38435 = ~n38430 & ~n38431 ;
  assign n38436 = ~n38426 & n38435 ;
  assign n38437 = ~n38427 & n38436 ;
  assign n38438 = ~n38425 & n38437 ;
  assign n38439 = ~n38434 & n38438 ;
  assign n38440 = n26792 & ~n38439 ;
  assign n38413 = \P2_P2_rEIP_reg[25]/NET0131  & n28046 ;
  assign n38414 = \P2_P2_InstAddrPointer_reg[25]/NET0131  & ~n32860 ;
  assign n38441 = ~n38413 & ~n38414 ;
  assign n38442 = ~n38440 & n38441 ;
  assign n38445 = \P1_P1_InstAddrPointer_reg[11]/NET0131  & n26249 ;
  assign n38451 = ~n33944 & n33948 ;
  assign n38452 = ~n29558 & ~n33949 ;
  assign n38453 = ~n38451 & n38452 ;
  assign n38446 = ~\P1_P1_InstAddrPointer_reg[11]/NET0131  & ~n33896 ;
  assign n38447 = ~n33946 & ~n38446 ;
  assign n38448 = ~n33817 & ~n38447 ;
  assign n38449 = ~n35730 & ~n38448 ;
  assign n38450 = n29558 & ~n38449 ;
  assign n38454 = ~n26249 & ~n38450 ;
  assign n38455 = ~n38453 & n38454 ;
  assign n38456 = ~n38445 & ~n38455 ;
  assign n38457 = n26126 & ~n38456 ;
  assign n38459 = ~\P1_P1_InstAddrPointer_reg[11]/NET0131  & ~n34029 ;
  assign n38460 = \P1_P1_InstAddrPointer_reg[11]/NET0131  & n34029 ;
  assign n38461 = ~n38459 & ~n38460 ;
  assign n38462 = ~n34098 & ~n38461 ;
  assign n38458 = \P1_P1_InstAddrPointer_reg[11]/NET0131  & n34098 ;
  assign n38463 = n26263 & ~n38458 ;
  assign n38464 = ~n38462 & n38463 ;
  assign n38467 = ~n15335 & n26162 ;
  assign n38468 = ~n26129 & ~n38467 ;
  assign n38469 = n38447 & ~n38468 ;
  assign n38444 = ~n26151 & n33948 ;
  assign n38465 = n26252 & ~n26255 ;
  assign n38466 = \P1_P1_InstAddrPointer_reg[11]/NET0131  & ~n38465 ;
  assign n38470 = n26192 & n38461 ;
  assign n38471 = ~\P1_P1_InstAddrPointer_reg[11]/NET0131  & ~n15365 ;
  assign n38472 = n15365 & ~n38447 ;
  assign n38473 = ~n38471 & ~n38472 ;
  assign n38474 = ~n15384 & n38473 ;
  assign n38475 = ~n38470 & ~n38474 ;
  assign n38476 = ~n38466 & n38475 ;
  assign n38477 = ~n38444 & n38476 ;
  assign n38478 = ~n38469 & n38477 ;
  assign n38479 = ~n38464 & n38478 ;
  assign n38480 = ~n38457 & n38479 ;
  assign n38481 = n8355 & ~n38480 ;
  assign n38443 = \P1_P1_rEIP_reg[11]/NET0131  & n8357 ;
  assign n38482 = \P1_P1_InstAddrPointer_reg[11]/NET0131  & ~n34164 ;
  assign n38483 = ~n38443 & ~n38482 ;
  assign n38484 = ~n38481 & n38483 ;
  assign n38487 = \P2_P3_InstAddrPointer_reg[11]/NET0131  & ~n27283 ;
  assign n38491 = ~\P2_P3_InstAddrPointer_reg[11]/NET0131  & ~n32916 ;
  assign n38492 = ~n32917 & ~n38491 ;
  assign n38493 = ~n33251 & ~n38492 ;
  assign n38494 = ~n33252 & ~n38493 ;
  assign n38495 = n33242 & ~n38494 ;
  assign n38488 = n33286 & ~n33338 ;
  assign n38489 = ~n33242 & ~n33339 ;
  assign n38490 = ~n38488 & n38489 ;
  assign n38496 = n27283 & ~n38490 ;
  assign n38497 = ~n38495 & n38496 ;
  assign n38498 = ~n38487 & ~n38497 ;
  assign n38499 = n27117 & ~n38498 ;
  assign n38500 = ~\P2_P3_InstAddrPointer_reg[11]/NET0131  & ~n32881 ;
  assign n38501 = ~n32882 & ~n38500 ;
  assign n38502 = ~n33477 & ~n38501 ;
  assign n38503 = n27280 & ~n33478 ;
  assign n38504 = ~n38502 & n38503 ;
  assign n38505 = ~n27180 & ~n32916 ;
  assign n38506 = n27229 & ~n38505 ;
  assign n38507 = n38492 & ~n38506 ;
  assign n38508 = ~n27142 & n33286 ;
  assign n38486 = \P2_P3_InstAddrPointer_reg[11]/NET0131  & ~n34355 ;
  assign n38509 = n27219 & n38501 ;
  assign n38510 = ~n38486 & ~n38509 ;
  assign n38511 = ~n38508 & n38510 ;
  assign n38512 = ~n38507 & n38511 ;
  assign n38513 = ~n38504 & n38512 ;
  assign n38514 = ~n38499 & n38513 ;
  assign n38515 = n27308 & ~n38514 ;
  assign n38485 = \P2_P3_rEIP_reg[11]/NET0131  & n32864 ;
  assign n38516 = \P2_P3_InstAddrPointer_reg[11]/NET0131  & ~n32870 ;
  assign n38517 = ~n38485 & ~n38516 ;
  assign n38518 = ~n38515 & n38517 ;
  assign n38521 = \P2_P3_InstAddrPointer_reg[14]/NET0131  & ~n27283 ;
  assign n38526 = ~\P2_P3_InstAddrPointer_reg[14]/NET0131  & ~n32953 ;
  assign n38527 = ~n32919 & ~n38526 ;
  assign n38528 = ~n33254 & ~n38527 ;
  assign n38529 = ~n33255 & ~n38528 ;
  assign n38530 = n33242 & ~n38529 ;
  assign n38522 = ~n33346 & n34329 ;
  assign n38523 = n33349 & ~n38522 ;
  assign n38524 = ~n33242 & ~n34330 ;
  assign n38525 = ~n38523 & n38524 ;
  assign n38531 = n27283 & ~n38525 ;
  assign n38532 = ~n38530 & n38531 ;
  assign n38533 = ~n38521 & ~n38532 ;
  assign n38534 = n27117 & ~n38533 ;
  assign n38535 = ~\P2_P3_InstAddrPointer_reg[14]/NET0131  & ~n33427 ;
  assign n38536 = ~n32885 & ~n38535 ;
  assign n38537 = ~n33480 & ~n38536 ;
  assign n38538 = n27280 & ~n33481 ;
  assign n38539 = ~n38537 & n38538 ;
  assign n38541 = ~n27229 & n38527 ;
  assign n38542 = \P2_P3_InstAddrPointer_reg[14]/NET0131  & ~n34355 ;
  assign n38520 = ~n27142 & n33349 ;
  assign n38540 = n27219 & n38536 ;
  assign n38543 = ~n38520 & ~n38540 ;
  assign n38544 = ~n38542 & n38543 ;
  assign n38545 = ~n38541 & n38544 ;
  assign n38546 = ~n38539 & n38545 ;
  assign n38547 = ~n38534 & n38546 ;
  assign n38548 = n27308 & ~n38547 ;
  assign n38519 = \P2_P3_rEIP_reg[14]/NET0131  & n32864 ;
  assign n38549 = \P2_P3_InstAddrPointer_reg[14]/NET0131  & ~n32870 ;
  assign n38550 = ~n38519 & ~n38549 ;
  assign n38551 = ~n38548 & n38550 ;
  assign n38553 = \P2_P3_InstAddrPointer_reg[16]/NET0131  & ~n27283 ;
  assign n38558 = ~n33258 & n35558 ;
  assign n38557 = n33258 & ~n35558 ;
  assign n38559 = n33242 & ~n38557 ;
  assign n38560 = ~n38558 & n38559 ;
  assign n38554 = n33355 & ~n37350 ;
  assign n38555 = ~n33242 & ~n34331 ;
  assign n38556 = ~n38554 & n38555 ;
  assign n38561 = n27283 & ~n38556 ;
  assign n38562 = ~n38560 & n38561 ;
  assign n38563 = ~n38553 & ~n38562 ;
  assign n38564 = n27117 & ~n38563 ;
  assign n38568 = ~n35657 & ~n35659 ;
  assign n38569 = n27280 & ~n35660 ;
  assign n38570 = ~n38568 & n38569 ;
  assign n38572 = ~n27229 & n33258 ;
  assign n38565 = ~n27180 & ~n32920 ;
  assign n38566 = n34355 & ~n38565 ;
  assign n38567 = \P2_P3_InstAddrPointer_reg[16]/NET0131  & ~n38566 ;
  assign n38571 = ~n27142 & n33355 ;
  assign n38573 = ~\P2_P3_InstAddrPointer_reg[16]/NET0131  & ~n27206 ;
  assign n38574 = ~n27111 & ~n38573 ;
  assign n38575 = n35659 & n38574 ;
  assign n38576 = ~n38571 & ~n38575 ;
  assign n38577 = ~n38567 & n38576 ;
  assign n38578 = ~n38572 & n38577 ;
  assign n38579 = ~n38570 & n38578 ;
  assign n38580 = ~n38564 & n38579 ;
  assign n38581 = n27308 & ~n38580 ;
  assign n38552 = \P2_P3_rEIP_reg[16]/NET0131  & n32864 ;
  assign n38582 = \P2_P3_InstAddrPointer_reg[16]/NET0131  & ~n32870 ;
  assign n38583 = ~n38552 & ~n38582 ;
  assign n38584 = ~n38581 & n38583 ;
  assign n38587 = \P2_P3_InstAddrPointer_reg[18]/NET0131  & ~n27283 ;
  assign n38592 = ~n37382 & ~n37384 ;
  assign n38593 = ~n37385 & ~n38592 ;
  assign n38594 = n33242 & ~n38593 ;
  assign n38588 = ~n33376 & n34331 ;
  assign n38589 = n33374 & ~n38588 ;
  assign n38590 = ~n33242 & ~n37389 ;
  assign n38591 = ~n38589 & n38590 ;
  assign n38595 = n27283 & ~n38591 ;
  assign n38596 = ~n38594 & n38595 ;
  assign n38597 = ~n38587 & ~n38596 ;
  assign n38598 = n27117 & ~n38597 ;
  assign n38599 = ~\P2_P3_InstAddrPointer_reg[18]/NET0131  & ~n33484 ;
  assign n38600 = ~n37398 & ~n38599 ;
  assign n38601 = ~n37401 & ~n38600 ;
  assign n38602 = n27280 & ~n37402 ;
  assign n38603 = ~n38601 & n38602 ;
  assign n38586 = ~n27229 & n37382 ;
  assign n38606 = \P2_P3_InstAddrPointer_reg[18]/NET0131  & ~n34355 ;
  assign n38607 = ~n38586 & ~n38606 ;
  assign n38604 = n27219 & n38600 ;
  assign n38605 = ~n27142 & n33374 ;
  assign n38608 = ~n38604 & ~n38605 ;
  assign n38609 = n38607 & n38608 ;
  assign n38610 = ~n38603 & n38609 ;
  assign n38611 = ~n38598 & n38610 ;
  assign n38612 = n27308 & ~n38611 ;
  assign n38585 = \P2_P3_rEIP_reg[18]/NET0131  & n32864 ;
  assign n38613 = \P2_P3_InstAddrPointer_reg[18]/NET0131  & ~n32870 ;
  assign n38614 = ~n38585 & ~n38613 ;
  assign n38615 = ~n38612 & n38614 ;
  assign n38618 = \P1_P1_InstAddrPointer_reg[14]/NET0131  & n26249 ;
  assign n38624 = n33952 & ~n33954 ;
  assign n38625 = n33956 & ~n38624 ;
  assign n38626 = ~n29558 & ~n33958 ;
  assign n38627 = ~n38625 & n38626 ;
  assign n38619 = ~\P1_P1_InstAddrPointer_reg[14]/NET0131  & ~n33550 ;
  assign n38620 = ~n33531 & ~n38619 ;
  assign n38621 = ~n33819 & ~n38620 ;
  assign n38622 = ~n33820 & ~n38621 ;
  assign n38623 = n29558 & ~n38622 ;
  assign n38628 = ~n26249 & ~n38623 ;
  assign n38629 = ~n38627 & n38628 ;
  assign n38630 = ~n38618 & ~n38629 ;
  assign n38631 = n26126 & ~n38630 ;
  assign n38632 = ~\P1_P1_InstAddrPointer_reg[14]/NET0131  & ~n34048 ;
  assign n38633 = ~n34031 & ~n38632 ;
  assign n38634 = ~n34100 & ~n38633 ;
  assign n38635 = n26263 & ~n34101 ;
  assign n38636 = ~n38634 & n38635 ;
  assign n38638 = ~n26189 & n38620 ;
  assign n38639 = ~n26151 & n33956 ;
  assign n38617 = \P1_P1_InstAddrPointer_reg[14]/NET0131  & ~n35760 ;
  assign n38637 = n26192 & n38633 ;
  assign n38640 = ~n38617 & ~n38637 ;
  assign n38641 = ~n38639 & n38640 ;
  assign n38642 = ~n38638 & n38641 ;
  assign n38643 = ~n38636 & n38642 ;
  assign n38644 = ~n38631 & n38643 ;
  assign n38645 = n8355 & ~n38644 ;
  assign n38616 = \P1_P1_rEIP_reg[14]/NET0131  & n8357 ;
  assign n38646 = \P1_P1_InstAddrPointer_reg[14]/NET0131  & ~n34164 ;
  assign n38647 = ~n38616 & ~n38646 ;
  assign n38648 = ~n38645 & n38647 ;
  assign n38653 = \P2_P3_InstAddrPointer_reg[21]/NET0131  & ~n27283 ;
  assign n38650 = ~\P2_P3_InstAddrPointer_reg[21]/NET0131  & ~n32923 ;
  assign n38651 = ~n33369 & ~n38650 ;
  assign n38657 = ~n33263 & ~n38651 ;
  assign n38658 = ~n35551 & ~n38657 ;
  assign n38659 = n33242 & ~n38658 ;
  assign n38654 = n33371 & ~n37423 ;
  assign n38655 = ~n33242 & ~n33381 ;
  assign n38656 = ~n38654 & n38655 ;
  assign n38660 = n27283 & ~n38656 ;
  assign n38661 = ~n38659 & n38660 ;
  assign n38662 = ~n38653 & ~n38661 ;
  assign n38663 = n27117 & ~n38662 ;
  assign n38664 = ~n33489 & ~n35656 ;
  assign n38665 = n27280 & ~n33490 ;
  assign n38666 = ~n38664 & n38665 ;
  assign n38668 = n27219 & n35656 ;
  assign n38667 = ~n27142 & n33371 ;
  assign n38652 = ~n27229 & n38651 ;
  assign n38669 = \P2_P3_InstAddrPointer_reg[21]/NET0131  & ~n34355 ;
  assign n38670 = ~n38652 & ~n38669 ;
  assign n38671 = ~n38667 & n38670 ;
  assign n38672 = ~n38668 & n38671 ;
  assign n38673 = ~n38666 & n38672 ;
  assign n38674 = ~n38663 & n38673 ;
  assign n38675 = n27308 & ~n38674 ;
  assign n38649 = \P2_P3_rEIP_reg[21]/NET0131  & n32864 ;
  assign n38676 = \P2_P3_InstAddrPointer_reg[21]/NET0131  & ~n32870 ;
  assign n38677 = ~n38649 & ~n38676 ;
  assign n38678 = ~n38675 & n38677 ;
  assign n38681 = \P2_P3_InstAddrPointer_reg[25]/NET0131  & ~n27283 ;
  assign n38685 = ~n32949 & ~n33264 ;
  assign n38686 = ~n35611 & ~n38685 ;
  assign n38687 = n33242 & ~n38686 ;
  assign n38682 = ~n33389 & n33392 ;
  assign n38683 = ~n33242 & ~n33393 ;
  assign n38684 = ~n38682 & n38683 ;
  assign n38688 = n27283 & ~n38684 ;
  assign n38689 = ~n38687 & n38688 ;
  assign n38690 = ~n38681 & ~n38689 ;
  assign n38691 = n27117 & ~n38690 ;
  assign n38692 = ~n33492 & ~n33494 ;
  assign n38693 = n27280 & ~n35620 ;
  assign n38694 = ~n38692 & n38693 ;
  assign n38702 = ~n27111 & n33494 ;
  assign n38703 = n27206 & n38702 ;
  assign n38704 = ~\P2_P3_InstAddrPointer_reg[25]/NET0131  & ~n38703 ;
  assign n38695 = ~n27192 & n32949 ;
  assign n38696 = \P2_P3_InstAddrPointer_reg[25]/NET0131  & n27192 ;
  assign n38697 = ~n38695 & ~n38696 ;
  assign n38705 = ~n27180 & ~n38697 ;
  assign n38706 = ~n27183 & n35581 ;
  assign n38707 = ~n38702 & n38706 ;
  assign n38708 = ~n38705 & n38707 ;
  assign n38709 = ~n38704 & ~n38708 ;
  assign n38698 = ~n27177 & ~n38697 ;
  assign n38699 = \P2_P3_InstAddrPointer_reg[25]/NET0131  & n27177 ;
  assign n38700 = ~n38698 & ~n38699 ;
  assign n38701 = n27186 & ~n38700 ;
  assign n38710 = ~n27200 & n38698 ;
  assign n38680 = n27057 & n32949 ;
  assign n38711 = ~n27142 & n33392 ;
  assign n38712 = ~n38680 & ~n38711 ;
  assign n38713 = ~n38710 & n38712 ;
  assign n38714 = ~n38701 & n38713 ;
  assign n38715 = ~n38709 & n38714 ;
  assign n38716 = ~n38694 & n38715 ;
  assign n38717 = ~n38691 & n38716 ;
  assign n38718 = n27308 & ~n38717 ;
  assign n38679 = \P2_P3_rEIP_reg[25]/NET0131  & n32864 ;
  assign n38719 = \P2_P3_InstAddrPointer_reg[25]/NET0131  & ~n32870 ;
  assign n38720 = ~n38679 & ~n38719 ;
  assign n38721 = ~n38718 & n38720 ;
  assign n38724 = \P1_P1_InstAddrPointer_reg[16]/NET0131  & n26249 ;
  assign n38728 = ~n33959 & n33961 ;
  assign n38729 = ~n29558 & ~n33962 ;
  assign n38730 = ~n38728 & n38729 ;
  assign n38725 = ~n35727 & ~n35733 ;
  assign n38726 = ~n35734 & ~n38725 ;
  assign n38727 = n29558 & ~n38726 ;
  assign n38731 = ~n26249 & ~n38727 ;
  assign n38732 = ~n38730 & n38731 ;
  assign n38733 = ~n38724 & ~n38732 ;
  assign n38734 = n26126 & ~n38733 ;
  assign n38735 = ~n35816 & ~n35818 ;
  assign n38736 = n26263 & ~n35819 ;
  assign n38737 = ~n38735 & n38736 ;
  assign n38740 = ~n26189 & n35727 ;
  assign n38723 = ~n26151 & n33961 ;
  assign n38738 = n26192 & n35818 ;
  assign n38739 = \P1_P1_InstAddrPointer_reg[16]/NET0131  & ~n35760 ;
  assign n38741 = ~n38738 & ~n38739 ;
  assign n38742 = ~n38723 & n38741 ;
  assign n38743 = ~n38740 & n38742 ;
  assign n38744 = ~n38737 & n38743 ;
  assign n38745 = ~n38734 & n38744 ;
  assign n38746 = n8355 & ~n38745 ;
  assign n38722 = \P1_P1_rEIP_reg[16]/NET0131  & n8357 ;
  assign n38747 = \P1_P1_InstAddrPointer_reg[16]/NET0131  & ~n34164 ;
  assign n38748 = ~n38722 & ~n38747 ;
  assign n38749 = ~n38746 & n38748 ;
  assign n38752 = \P1_P1_InstAddrPointer_reg[18]/NET0131  & n26249 ;
  assign n38758 = ~n33963 & n33973 ;
  assign n38759 = ~n29558 & ~n37586 ;
  assign n38760 = ~n38758 & n38759 ;
  assign n38753 = ~\P1_P1_InstAddrPointer_reg[18]/NET0131  & ~n33823 ;
  assign n38754 = ~n33968 & ~n38753 ;
  assign n38755 = ~n37581 & ~n38754 ;
  assign n38756 = ~n37582 & ~n38755 ;
  assign n38757 = n29558 & ~n38756 ;
  assign n38761 = ~n26249 & ~n38757 ;
  assign n38762 = ~n38760 & n38761 ;
  assign n38763 = ~n38752 & ~n38762 ;
  assign n38764 = n26126 & ~n38763 ;
  assign n38765 = ~\P1_P1_InstAddrPointer_reg[18]/NET0131  & ~n34104 ;
  assign n38766 = ~n37574 & ~n38765 ;
  assign n38767 = ~n34107 & ~n38766 ;
  assign n38768 = n26263 & ~n37595 ;
  assign n38769 = ~n38767 & n38768 ;
  assign n38771 = \P1_P1_InstAddrPointer_reg[18]/NET0131  & ~n34390 ;
  assign n38770 = ~n26189 & n38754 ;
  assign n38751 = ~n26151 & n33973 ;
  assign n38772 = ~\P1_P1_InstAddrPointer_reg[18]/NET0131  & ~n15428 ;
  assign n38773 = ~n26123 & ~n38772 ;
  assign n38774 = n38766 & n38773 ;
  assign n38775 = ~n38751 & ~n38774 ;
  assign n38776 = ~n38770 & n38775 ;
  assign n38777 = ~n38771 & n38776 ;
  assign n38778 = ~n38769 & n38777 ;
  assign n38779 = ~n38764 & n38778 ;
  assign n38780 = n8355 & ~n38779 ;
  assign n38750 = \P1_P1_rEIP_reg[18]/NET0131  & n8357 ;
  assign n38781 = \P1_P1_InstAddrPointer_reg[18]/NET0131  & ~n34164 ;
  assign n38782 = ~n38750 & ~n38781 ;
  assign n38783 = ~n38780 & n38782 ;
  assign n38786 = \P1_P1_InstAddrPointer_reg[21]/NET0131  & n26249 ;
  assign n38790 = n33967 & ~n37624 ;
  assign n38791 = ~n29558 & ~n33979 ;
  assign n38792 = ~n38790 & n38791 ;
  assign n38787 = ~n33830 & ~n33848 ;
  assign n38788 = ~n37650 & ~n38787 ;
  assign n38789 = n29558 & ~n38788 ;
  assign n38793 = ~n26249 & ~n38789 ;
  assign n38794 = ~n38792 & n38793 ;
  assign n38795 = ~n38786 & ~n38794 ;
  assign n38796 = n26126 & ~n38795 ;
  assign n38797 = ~n34109 & ~n35815 ;
  assign n38798 = n26263 & ~n34110 ;
  assign n38799 = ~n38797 & n38798 ;
  assign n38800 = ~\P1_P1_InstAddrPointer_reg[21]/NET0131  & ~n15428 ;
  assign n38801 = ~n26123 & n35815 ;
  assign n38802 = n26252 & ~n38801 ;
  assign n38803 = ~n38800 & ~n38802 ;
  assign n38785 = ~n26189 & n33848 ;
  assign n38804 = ~n15384 & ~n33535 ;
  assign n38805 = n26256 & ~n38804 ;
  assign n38806 = \P1_P1_InstAddrPointer_reg[21]/NET0131  & ~n38805 ;
  assign n38807 = ~n26151 & n33967 ;
  assign n38808 = ~n38806 & ~n38807 ;
  assign n38809 = ~n38785 & n38808 ;
  assign n38810 = ~n38803 & n38809 ;
  assign n38811 = ~n38799 & n38810 ;
  assign n38812 = ~n38796 & n38811 ;
  assign n38813 = n8355 & ~n38812 ;
  assign n38784 = \P1_P1_InstAddrPointer_reg[21]/NET0131  & ~n34164 ;
  assign n38814 = \P1_P1_rEIP_reg[21]/NET0131  & n8357 ;
  assign n38815 = ~n38784 & ~n38814 ;
  assign n38816 = ~n38813 & n38815 ;
  assign n38836 = ~n34121 & ~n34123 ;
  assign n38837 = n26263 & ~n35781 ;
  assign n38838 = ~n38836 & n38837 ;
  assign n38819 = \P1_P1_InstAddrPointer_reg[25]/NET0131  & n26249 ;
  assign n38823 = n33985 & ~n37713 ;
  assign n38824 = ~n29558 & ~n33990 ;
  assign n38825 = ~n38823 & n38824 ;
  assign n38820 = ~n33855 & ~n33857 ;
  assign n38821 = ~n35770 & ~n38820 ;
  assign n38822 = n29558 & ~n38821 ;
  assign n38826 = ~n26249 & ~n38822 ;
  assign n38827 = ~n38825 & n38826 ;
  assign n38828 = ~n38819 & ~n38827 ;
  assign n38829 = n26126 & ~n38828 ;
  assign n38835 = ~n26151 & n33985 ;
  assign n38833 = n26192 & n34123 ;
  assign n38830 = ~n26160 & ~n33537 ;
  assign n38831 = n35760 & ~n38830 ;
  assign n38832 = \P1_P1_InstAddrPointer_reg[25]/NET0131  & ~n38831 ;
  assign n38834 = ~n26189 & n33857 ;
  assign n38839 = ~n38832 & ~n38834 ;
  assign n38840 = ~n38833 & n38839 ;
  assign n38841 = ~n38835 & n38840 ;
  assign n38842 = ~n38829 & n38841 ;
  assign n38843 = ~n38838 & n38842 ;
  assign n38844 = n8355 & ~n38843 ;
  assign n38817 = \P1_P1_rEIP_reg[25]/NET0131  & n8357 ;
  assign n38818 = \P1_P1_InstAddrPointer_reg[25]/NET0131  & ~n34164 ;
  assign n38845 = ~n38817 & ~n38818 ;
  assign n38846 = ~n38844 & n38845 ;
  assign n38849 = \P1_P2_InstAddrPointer_reg[11]/NET0131  & n25733 ;
  assign n38853 = ~n31252 & n31254 ;
  assign n38854 = ~n30809 & ~n31255 ;
  assign n38855 = ~n38853 & n38854 ;
  assign n38850 = ~n31120 & ~n35201 ;
  assign n38851 = ~n31121 & ~n38850 ;
  assign n38852 = n30809 & ~n38851 ;
  assign n38856 = ~n25733 & ~n38852 ;
  assign n38857 = ~n38855 & n38856 ;
  assign n38858 = ~n38849 & ~n38857 ;
  assign n38859 = n25701 & ~n38858 ;
  assign n38861 = ~\P1_P2_InstAddrPointer_reg[11]/NET0131  & n31365 ;
  assign n38862 = \P1_P2_InstAddrPointer_reg[11]/NET0131  & ~n31365 ;
  assign n38863 = ~n38861 & ~n38862 ;
  assign n38864 = ~n31417 & n38863 ;
  assign n38860 = \P1_P2_InstAddrPointer_reg[11]/NET0131  & n31417 ;
  assign n38865 = n25881 & ~n38860 ;
  assign n38866 = ~n38864 & n38865 ;
  assign n38867 = ~n25817 & n31254 ;
  assign n38868 = \P1_P2_InstAddrPointer_reg[11]/NET0131  & ~n25788 ;
  assign n38869 = n25773 & n35201 ;
  assign n38870 = ~n38868 & ~n38869 ;
  assign n38871 = \P1_P2_InstAddrPointer_reg[11]/NET0131  & ~n25763 ;
  assign n38872 = n25828 & ~n38871 ;
  assign n38873 = ~n38870 & ~n38872 ;
  assign n38874 = ~n25743 & ~n31350 ;
  assign n38875 = n25753 & ~n38874 ;
  assign n38876 = \P1_P2_InstAddrPointer_reg[11]/NET0131  & ~n38875 ;
  assign n38848 = n25808 & n35201 ;
  assign n38877 = n25887 & n38861 ;
  assign n38878 = ~n38848 & ~n38877 ;
  assign n38879 = ~n38876 & n38878 ;
  assign n38880 = ~n38873 & n38879 ;
  assign n38881 = ~n38867 & n38880 ;
  assign n38882 = ~n38866 & n38881 ;
  assign n38883 = ~n38859 & n38882 ;
  assign n38884 = n25918 & ~n38883 ;
  assign n38847 = \P1_P2_rEIP_reg[11]/NET0131  & n27967 ;
  assign n38885 = \P1_P2_InstAddrPointer_reg[11]/NET0131  & ~n31487 ;
  assign n38886 = ~n38847 & ~n38885 ;
  assign n38887 = ~n38884 & n38886 ;
  assign n38890 = \P1_P2_InstAddrPointer_reg[14]/NET0131  & n25733 ;
  assign n38894 = ~n31264 & n31267 ;
  assign n38895 = ~n30809 & ~n31268 ;
  assign n38896 = ~n38894 & n38895 ;
  assign n38891 = ~n31122 & ~n31125 ;
  assign n38892 = ~n31126 & ~n38891 ;
  assign n38893 = n30809 & ~n38892 ;
  assign n38897 = ~n25733 & ~n38893 ;
  assign n38898 = ~n38896 & n38897 ;
  assign n38899 = ~n38890 & ~n38898 ;
  assign n38900 = n25701 & ~n38899 ;
  assign n38901 = ~\P1_P2_InstAddrPointer_reg[14]/NET0131  & ~n31351 ;
  assign n38902 = ~n31341 & ~n38901 ;
  assign n38903 = ~n31419 & ~n38902 ;
  assign n38904 = n25881 & ~n31420 ;
  assign n38905 = ~n38903 & n38904 ;
  assign n38910 = ~n25763 & ~n31123 ;
  assign n38911 = n25830 & ~n38910 ;
  assign n38912 = n31125 & ~n38911 ;
  assign n38889 = ~n25817 & n31267 ;
  assign n38906 = n25773 & ~n31125 ;
  assign n38907 = ~n25828 & ~n38906 ;
  assign n38908 = n31467 & ~n38907 ;
  assign n38909 = \P1_P2_InstAddrPointer_reg[14]/NET0131  & ~n38908 ;
  assign n38913 = n25887 & n38902 ;
  assign n38914 = ~n38909 & ~n38913 ;
  assign n38915 = ~n38889 & n38914 ;
  assign n38916 = ~n38912 & n38915 ;
  assign n38917 = ~n38905 & n38916 ;
  assign n38918 = ~n38900 & n38917 ;
  assign n38919 = n25918 & ~n38918 ;
  assign n38888 = \P1_P2_rEIP_reg[14]/NET0131  & n27967 ;
  assign n38920 = \P1_P2_InstAddrPointer_reg[14]/NET0131  & ~n31487 ;
  assign n38921 = ~n38888 & ~n38920 ;
  assign n38922 = ~n38919 & n38921 ;
  assign n38940 = ~n31272 & n31274 ;
  assign n38941 = ~n31275 & ~n38940 ;
  assign n38942 = ~n30809 & ~n38941 ;
  assign n38944 = ~n31127 & ~n31137 ;
  assign n38943 = \P1_P2_InstAddrPointer_reg[16]/NET0131  & n31127 ;
  assign n38945 = n30809 & ~n38943 ;
  assign n38946 = ~n38944 & n38945 ;
  assign n38947 = ~n38942 & ~n38946 ;
  assign n38948 = ~n25733 & n38947 ;
  assign n38939 = ~\P1_P2_InstAddrPointer_reg[16]/NET0131  & n25733 ;
  assign n38949 = n25701 & ~n38939 ;
  assign n38950 = ~n38948 & n38949 ;
  assign n38925 = ~n35176 & ~n35177 ;
  assign n38926 = n25881 & ~n35178 ;
  assign n38927 = ~n38925 & n38926 ;
  assign n38929 = n36899 & ~n38874 ;
  assign n38930 = \P1_P2_InstAddrPointer_reg[16]/NET0131  & ~n38929 ;
  assign n38928 = ~n25817 & n31274 ;
  assign n38931 = ~\P1_P2_InstAddrPointer_reg[16]/NET0131  & n25415 ;
  assign n38932 = ~n25415 & ~n31137 ;
  assign n38933 = ~n38931 & ~n38932 ;
  assign n38934 = ~n36900 & n38933 ;
  assign n38924 = n25808 & n31137 ;
  assign n38935 = n25887 & n31350 ;
  assign n38936 = ~\P1_P2_InstAddrPointer_reg[16]/NET0131  & ~n30846 ;
  assign n38937 = ~n30847 & ~n38936 ;
  assign n38938 = n38935 & n38937 ;
  assign n38951 = ~n38924 & ~n38938 ;
  assign n38952 = ~n38934 & n38951 ;
  assign n38953 = ~n38928 & n38952 ;
  assign n38954 = ~n38930 & n38953 ;
  assign n38955 = ~n38927 & n38954 ;
  assign n38956 = ~n38950 & n38955 ;
  assign n38957 = n25918 & ~n38956 ;
  assign n38923 = \P1_P2_rEIP_reg[16]/NET0131  & n27967 ;
  assign n38958 = \P1_P2_InstAddrPointer_reg[16]/NET0131  & ~n31487 ;
  assign n38959 = ~n38923 & ~n38958 ;
  assign n38960 = ~n38957 & n38959 ;
  assign n38963 = \P1_P2_InstAddrPointer_reg[18]/NET0131  & n25733 ;
  assign n38967 = n31286 & ~n37819 ;
  assign n38968 = ~n30809 & ~n37820 ;
  assign n38969 = ~n38967 & n38968 ;
  assign n38964 = ~n37811 & ~n37813 ;
  assign n38965 = ~n37814 & ~n38964 ;
  assign n38966 = n30809 & ~n38965 ;
  assign n38970 = ~n25733 & ~n38966 ;
  assign n38971 = ~n38969 & n38970 ;
  assign n38972 = ~n38963 & ~n38971 ;
  assign n38973 = n25701 & ~n38972 ;
  assign n38975 = ~\P1_P2_InstAddrPointer_reg[18]/NET0131  & ~n31425 ;
  assign n38976 = ~n37832 & ~n38975 ;
  assign n38980 = \P1_P2_InstAddrPointer_reg[17]/NET0131  & n31424 ;
  assign n38981 = ~n38976 & ~n38980 ;
  assign n38982 = n25881 & ~n31429 ;
  assign n38983 = ~n38981 & n38982 ;
  assign n38974 = ~n34215 & n37813 ;
  assign n38977 = n25887 & n38976 ;
  assign n38984 = ~n38974 & ~n38977 ;
  assign n38978 = \P1_P2_InstAddrPointer_reg[18]/NET0131  & ~n34210 ;
  assign n38979 = ~n25817 & n31286 ;
  assign n38985 = ~n38978 & ~n38979 ;
  assign n38986 = n38984 & n38985 ;
  assign n38987 = ~n38983 & n38986 ;
  assign n38988 = ~n38973 & n38987 ;
  assign n38989 = n25918 & ~n38988 ;
  assign n38961 = \P1_P2_rEIP_reg[18]/NET0131  & n27967 ;
  assign n38962 = \P1_P2_InstAddrPointer_reg[18]/NET0131  & ~n31487 ;
  assign n38990 = ~n38961 & ~n38962 ;
  assign n38991 = ~n38989 & n38990 ;
  assign n38994 = \P1_P2_InstAddrPointer_reg[21]/NET0131  & n25733 ;
  assign n38998 = n31195 & ~n31290 ;
  assign n38999 = ~n30809 & ~n31291 ;
  assign n39000 = ~n38998 & n38999 ;
  assign n38995 = ~n30852 & ~n35208 ;
  assign n38996 = ~n35209 & ~n38995 ;
  assign n38997 = n30809 & ~n38996 ;
  assign n39001 = ~n25733 & ~n38997 ;
  assign n39002 = ~n39000 & n39001 ;
  assign n39003 = ~n38994 & ~n39002 ;
  assign n39004 = n25701 & ~n39003 ;
  assign n39005 = ~n31431 & ~n35174 ;
  assign n39006 = n25881 & ~n31432 ;
  assign n39007 = ~n39005 & n39006 ;
  assign n38993 = ~n25817 & n31195 ;
  assign n39008 = n25887 & n35174 ;
  assign n39011 = ~n38993 & ~n39008 ;
  assign n39009 = n30852 & ~n34215 ;
  assign n39010 = \P1_P2_InstAddrPointer_reg[21]/NET0131  & ~n34210 ;
  assign n39012 = ~n39009 & ~n39010 ;
  assign n39013 = n39011 & n39012 ;
  assign n39014 = ~n39007 & n39013 ;
  assign n39015 = ~n39004 & n39014 ;
  assign n39016 = n25918 & ~n39015 ;
  assign n38992 = \P1_P2_InstAddrPointer_reg[21]/NET0131  & ~n31487 ;
  assign n39017 = \P1_P2_rEIP_reg[21]/NET0131  & n27967 ;
  assign n39018 = ~n38992 & ~n39017 ;
  assign n39019 = ~n39016 & n39018 ;
  assign n39020 = n15736 & n18665 ;
  assign n39032 = \P2_buf2_reg[29]/NET0131  & ~n28013 ;
  assign n39033 = \P2_buf1_reg[29]/NET0131  & n28013 ;
  assign n39034 = ~n39032 & ~n39033 ;
  assign n39035 = n28027 & ~n39034 ;
  assign n39036 = \P2_buf2_reg[21]/NET0131  & ~n28013 ;
  assign n39037 = \P2_buf1_reg[21]/NET0131  & n28013 ;
  assign n39038 = ~n39036 & ~n39037 ;
  assign n39039 = n28034 & ~n39038 ;
  assign n39040 = ~n39035 & ~n39039 ;
  assign n39041 = \P2_P2_DataWidth_reg[1]/NET0131  & ~n39040 ;
  assign n39021 = \P2_buf2_reg[5]/NET0131  & ~n28013 ;
  assign n39022 = \P2_buf1_reg[5]/NET0131  & n28013 ;
  assign n39023 = ~n39021 & ~n39022 ;
  assign n39024 = ~n27984 & ~n39023 ;
  assign n39025 = \P2_P2_InstQueue_reg[11][5]/NET0131  & ~n27980 ;
  assign n39026 = ~n27983 & n39025 ;
  assign n39027 = ~n39024 & ~n39026 ;
  assign n39042 = ~n28042 & ~n39027 ;
  assign n39043 = ~n39041 & ~n39042 ;
  assign n39044 = n26794 & ~n39043 ;
  assign n39029 = ~n26449 & n27980 ;
  assign n39030 = ~n39025 & ~n39029 ;
  assign n39031 = n27613 & ~n39030 ;
  assign n39028 = n27977 & ~n39027 ;
  assign n39045 = \P2_P2_InstQueue_reg[11][5]/NET0131  & ~n28050 ;
  assign n39046 = ~n39028 & ~n39045 ;
  assign n39047 = ~n39031 & n39046 ;
  assign n39048 = ~n39044 & n39047 ;
  assign n39057 = n28398 & ~n39034 ;
  assign n39058 = n28401 & ~n39038 ;
  assign n39059 = ~n39057 & ~n39058 ;
  assign n39060 = \P2_P2_DataWidth_reg[1]/NET0131  & ~n39059 ;
  assign n39049 = ~n28388 & ~n39023 ;
  assign n39050 = \P2_P2_InstQueue_reg[0][5]/NET0131  & ~n28385 ;
  assign n39051 = ~n28387 & n39050 ;
  assign n39052 = ~n39049 & ~n39051 ;
  assign n39061 = ~n28406 & ~n39052 ;
  assign n39062 = ~n39060 & ~n39061 ;
  assign n39063 = n26794 & ~n39062 ;
  assign n39054 = ~n26449 & n28385 ;
  assign n39055 = ~n39050 & ~n39054 ;
  assign n39056 = n27613 & ~n39055 ;
  assign n39053 = n27977 & ~n39052 ;
  assign n39064 = \P2_P2_InstQueue_reg[0][5]/NET0131  & ~n28050 ;
  assign n39065 = ~n39053 & ~n39064 ;
  assign n39066 = ~n39056 & n39065 ;
  assign n39067 = ~n39063 & n39066 ;
  assign n39076 = n28423 & ~n39034 ;
  assign n39077 = n28027 & ~n39038 ;
  assign n39078 = ~n39076 & ~n39077 ;
  assign n39079 = \P2_P2_DataWidth_reg[1]/NET0131  & ~n39078 ;
  assign n39068 = ~n28414 & ~n39023 ;
  assign n39069 = \P2_P2_InstQueue_reg[10][5]/NET0131  & ~n27983 ;
  assign n39070 = ~n28034 & n39069 ;
  assign n39071 = ~n39068 & ~n39070 ;
  assign n39080 = ~n28429 & ~n39071 ;
  assign n39081 = ~n39079 & ~n39080 ;
  assign n39082 = n26794 & ~n39081 ;
  assign n39073 = ~n26449 & n27983 ;
  assign n39074 = ~n39069 & ~n39073 ;
  assign n39075 = n27613 & ~n39074 ;
  assign n39072 = n27977 & ~n39071 ;
  assign n39083 = \P2_P2_InstQueue_reg[10][5]/NET0131  & ~n28050 ;
  assign n39084 = ~n39072 & ~n39083 ;
  assign n39085 = ~n39075 & n39084 ;
  assign n39086 = ~n39082 & n39085 ;
  assign n39095 = n28034 & ~n39034 ;
  assign n39096 = n27983 & ~n39038 ;
  assign n39097 = ~n39095 & ~n39096 ;
  assign n39098 = \P2_P2_DataWidth_reg[1]/NET0131  & ~n39097 ;
  assign n39087 = ~n28439 & ~n39023 ;
  assign n39088 = \P2_P2_InstQueue_reg[12][5]/NET0131  & ~n28438 ;
  assign n39089 = ~n27980 & n39088 ;
  assign n39090 = ~n39087 & ~n39089 ;
  assign n39099 = ~n28452 & ~n39090 ;
  assign n39100 = ~n39098 & ~n39099 ;
  assign n39101 = n26794 & ~n39100 ;
  assign n39092 = ~n26449 & n28438 ;
  assign n39093 = ~n39088 & ~n39092 ;
  assign n39094 = n27613 & ~n39093 ;
  assign n39091 = n27977 & ~n39090 ;
  assign n39102 = \P2_P2_InstQueue_reg[12][5]/NET0131  & ~n28050 ;
  assign n39103 = ~n39091 & ~n39102 ;
  assign n39104 = ~n39094 & n39103 ;
  assign n39105 = ~n39101 & n39104 ;
  assign n39114 = n27983 & ~n39034 ;
  assign n39115 = n27980 & ~n39038 ;
  assign n39116 = ~n39114 & ~n39115 ;
  assign n39117 = \P2_P2_DataWidth_reg[1]/NET0131  & ~n39116 ;
  assign n39106 = ~n28460 & ~n39023 ;
  assign n39107 = \P2_P2_InstQueue_reg[13][5]/NET0131  & ~n28398 ;
  assign n39108 = ~n28438 & n39107 ;
  assign n39109 = ~n39106 & ~n39108 ;
  assign n39118 = ~n28473 & ~n39109 ;
  assign n39119 = ~n39117 & ~n39118 ;
  assign n39120 = n26794 & ~n39119 ;
  assign n39111 = ~n26449 & n28398 ;
  assign n39112 = ~n39107 & ~n39111 ;
  assign n39113 = n27613 & ~n39112 ;
  assign n39110 = n27977 & ~n39109 ;
  assign n39121 = \P2_P2_InstQueue_reg[13][5]/NET0131  & ~n28050 ;
  assign n39122 = ~n39110 & ~n39121 ;
  assign n39123 = ~n39113 & n39122 ;
  assign n39124 = ~n39120 & n39123 ;
  assign n39133 = n27980 & ~n39034 ;
  assign n39134 = n28438 & ~n39038 ;
  assign n39135 = ~n39133 & ~n39134 ;
  assign n39136 = \P2_P2_DataWidth_reg[1]/NET0131  & ~n39135 ;
  assign n39125 = ~n28405 & ~n39023 ;
  assign n39126 = \P2_P2_InstQueue_reg[14][5]/NET0131  & ~n28401 ;
  assign n39127 = ~n28398 & n39126 ;
  assign n39128 = ~n39125 & ~n39127 ;
  assign n39137 = ~n28493 & ~n39128 ;
  assign n39138 = ~n39136 & ~n39137 ;
  assign n39139 = n26794 & ~n39138 ;
  assign n39130 = ~n26449 & n28401 ;
  assign n39131 = ~n39126 & ~n39130 ;
  assign n39132 = n27613 & ~n39131 ;
  assign n39129 = n27977 & ~n39128 ;
  assign n39140 = \P2_P2_InstQueue_reg[14][5]/NET0131  & ~n28050 ;
  assign n39141 = ~n39129 & ~n39140 ;
  assign n39142 = ~n39132 & n39141 ;
  assign n39143 = ~n39139 & n39142 ;
  assign n39152 = n28438 & ~n39034 ;
  assign n39153 = n28398 & ~n39038 ;
  assign n39154 = ~n39152 & ~n39153 ;
  assign n39155 = \P2_P2_DataWidth_reg[1]/NET0131  & ~n39154 ;
  assign n39144 = ~n28501 & ~n39023 ;
  assign n39145 = \P2_P2_InstQueue_reg[15][5]/NET0131  & ~n28387 ;
  assign n39146 = ~n28401 & n39145 ;
  assign n39147 = ~n39144 & ~n39146 ;
  assign n39156 = ~n28514 & ~n39147 ;
  assign n39157 = ~n39155 & ~n39156 ;
  assign n39158 = n26794 & ~n39157 ;
  assign n39149 = ~n26449 & n28387 ;
  assign n39150 = ~n39145 & ~n39149 ;
  assign n39151 = n27613 & ~n39150 ;
  assign n39148 = n27977 & ~n39147 ;
  assign n39159 = \P2_P2_InstQueue_reg[15][5]/NET0131  & ~n28050 ;
  assign n39160 = ~n39148 & ~n39159 ;
  assign n39161 = ~n39151 & n39160 ;
  assign n39162 = ~n39158 & n39161 ;
  assign n39171 = n28401 & ~n39034 ;
  assign n39172 = n28387 & ~n39038 ;
  assign n39173 = ~n39171 & ~n39172 ;
  assign n39174 = \P2_P2_DataWidth_reg[1]/NET0131  & ~n39173 ;
  assign n39163 = ~n28523 & ~n39023 ;
  assign n39164 = \P2_P2_InstQueue_reg[1][5]/NET0131  & ~n28522 ;
  assign n39165 = ~n28385 & n39164 ;
  assign n39166 = ~n39163 & ~n39165 ;
  assign n39175 = ~n28536 & ~n39166 ;
  assign n39176 = ~n39174 & ~n39175 ;
  assign n39177 = n26794 & ~n39176 ;
  assign n39168 = ~n26449 & n28522 ;
  assign n39169 = ~n39164 & ~n39168 ;
  assign n39170 = n27613 & ~n39169 ;
  assign n39167 = n27977 & ~n39166 ;
  assign n39178 = \P2_P2_InstQueue_reg[1][5]/NET0131  & ~n28050 ;
  assign n39179 = ~n39167 & ~n39178 ;
  assign n39180 = ~n39170 & n39179 ;
  assign n39181 = ~n39177 & n39180 ;
  assign n39190 = n28387 & ~n39034 ;
  assign n39191 = n28385 & ~n39038 ;
  assign n39192 = ~n39190 & ~n39191 ;
  assign n39193 = \P2_P2_DataWidth_reg[1]/NET0131  & ~n39192 ;
  assign n39182 = ~n28545 & ~n39023 ;
  assign n39183 = \P2_P2_InstQueue_reg[2][5]/NET0131  & ~n28544 ;
  assign n39184 = ~n28522 & n39183 ;
  assign n39185 = ~n39182 & ~n39184 ;
  assign n39194 = ~n28558 & ~n39185 ;
  assign n39195 = ~n39193 & ~n39194 ;
  assign n39196 = n26794 & ~n39195 ;
  assign n39187 = ~n26449 & n28544 ;
  assign n39188 = ~n39183 & ~n39187 ;
  assign n39189 = n27613 & ~n39188 ;
  assign n39186 = n27977 & ~n39185 ;
  assign n39197 = \P2_P2_InstQueue_reg[2][5]/NET0131  & ~n28050 ;
  assign n39198 = ~n39186 & ~n39197 ;
  assign n39199 = ~n39189 & n39198 ;
  assign n39200 = ~n39196 & n39199 ;
  assign n39209 = n28385 & ~n39034 ;
  assign n39210 = n28522 & ~n39038 ;
  assign n39211 = ~n39209 & ~n39210 ;
  assign n39212 = \P2_P2_DataWidth_reg[1]/NET0131  & ~n39211 ;
  assign n39201 = ~n28567 & ~n39023 ;
  assign n39202 = \P2_P2_InstQueue_reg[3][5]/NET0131  & ~n28566 ;
  assign n39203 = ~n28544 & n39202 ;
  assign n39204 = ~n39201 & ~n39203 ;
  assign n39213 = ~n28580 & ~n39204 ;
  assign n39214 = ~n39212 & ~n39213 ;
  assign n39215 = n26794 & ~n39214 ;
  assign n39206 = ~n26449 & n28566 ;
  assign n39207 = ~n39202 & ~n39206 ;
  assign n39208 = n27613 & ~n39207 ;
  assign n39205 = n27977 & ~n39204 ;
  assign n39216 = \P2_P2_InstQueue_reg[3][5]/NET0131  & ~n28050 ;
  assign n39217 = ~n39205 & ~n39216 ;
  assign n39218 = ~n39208 & n39217 ;
  assign n39219 = ~n39215 & n39218 ;
  assign n39228 = n28522 & ~n39034 ;
  assign n39229 = n28544 & ~n39038 ;
  assign n39230 = ~n39228 & ~n39229 ;
  assign n39231 = \P2_P2_DataWidth_reg[1]/NET0131  & ~n39230 ;
  assign n39220 = ~n28589 & ~n39023 ;
  assign n39221 = \P2_P2_InstQueue_reg[4][5]/NET0131  & ~n28588 ;
  assign n39222 = ~n28566 & n39221 ;
  assign n39223 = ~n39220 & ~n39222 ;
  assign n39232 = ~n28602 & ~n39223 ;
  assign n39233 = ~n39231 & ~n39232 ;
  assign n39234 = n26794 & ~n39233 ;
  assign n39225 = ~n26449 & n28588 ;
  assign n39226 = ~n39221 & ~n39225 ;
  assign n39227 = n27613 & ~n39226 ;
  assign n39224 = n27977 & ~n39223 ;
  assign n39235 = \P2_P2_InstQueue_reg[4][5]/NET0131  & ~n28050 ;
  assign n39236 = ~n39224 & ~n39235 ;
  assign n39237 = ~n39227 & n39236 ;
  assign n39238 = ~n39234 & n39237 ;
  assign n39247 = n28544 & ~n39034 ;
  assign n39248 = n28566 & ~n39038 ;
  assign n39249 = ~n39247 & ~n39248 ;
  assign n39250 = \P2_P2_DataWidth_reg[1]/NET0131  & ~n39249 ;
  assign n39239 = ~n28611 & ~n39023 ;
  assign n39240 = \P2_P2_InstQueue_reg[5][5]/NET0131  & ~n28610 ;
  assign n39241 = ~n28588 & n39240 ;
  assign n39242 = ~n39239 & ~n39241 ;
  assign n39251 = ~n28624 & ~n39242 ;
  assign n39252 = ~n39250 & ~n39251 ;
  assign n39253 = n26794 & ~n39252 ;
  assign n39244 = ~n26449 & n28610 ;
  assign n39245 = ~n39240 & ~n39244 ;
  assign n39246 = n27613 & ~n39245 ;
  assign n39243 = n27977 & ~n39242 ;
  assign n39254 = \P2_P2_InstQueue_reg[5][5]/NET0131  & ~n28050 ;
  assign n39255 = ~n39243 & ~n39254 ;
  assign n39256 = ~n39246 & n39255 ;
  assign n39257 = ~n39253 & n39256 ;
  assign n39266 = n28566 & ~n39034 ;
  assign n39267 = n28588 & ~n39038 ;
  assign n39268 = ~n39266 & ~n39267 ;
  assign n39269 = \P2_P2_DataWidth_reg[1]/NET0131  & ~n39268 ;
  assign n39258 = ~n28633 & ~n39023 ;
  assign n39259 = \P2_P2_InstQueue_reg[6][5]/NET0131  & ~n28632 ;
  assign n39260 = ~n28610 & n39259 ;
  assign n39261 = ~n39258 & ~n39260 ;
  assign n39270 = ~n28646 & ~n39261 ;
  assign n39271 = ~n39269 & ~n39270 ;
  assign n39272 = n26794 & ~n39271 ;
  assign n39263 = ~n26449 & n28632 ;
  assign n39264 = ~n39259 & ~n39263 ;
  assign n39265 = n27613 & ~n39264 ;
  assign n39262 = n27977 & ~n39261 ;
  assign n39273 = \P2_P2_InstQueue_reg[6][5]/NET0131  & ~n28050 ;
  assign n39274 = ~n39262 & ~n39273 ;
  assign n39275 = ~n39265 & n39274 ;
  assign n39276 = ~n39272 & n39275 ;
  assign n39285 = n28588 & ~n39034 ;
  assign n39286 = n28610 & ~n39038 ;
  assign n39287 = ~n39285 & ~n39286 ;
  assign n39288 = \P2_P2_DataWidth_reg[1]/NET0131  & ~n39287 ;
  assign n39277 = ~n28654 & ~n39023 ;
  assign n39278 = \P2_P2_InstQueue_reg[7][5]/NET0131  & ~n28423 ;
  assign n39279 = ~n28632 & n39278 ;
  assign n39280 = ~n39277 & ~n39279 ;
  assign n39289 = ~n28667 & ~n39280 ;
  assign n39290 = ~n39288 & ~n39289 ;
  assign n39291 = n26794 & ~n39290 ;
  assign n39282 = ~n26449 & n28423 ;
  assign n39283 = ~n39278 & ~n39282 ;
  assign n39284 = n27613 & ~n39283 ;
  assign n39281 = n27977 & ~n39280 ;
  assign n39292 = \P2_P2_InstQueue_reg[7][5]/NET0131  & ~n28050 ;
  assign n39293 = ~n39281 & ~n39292 ;
  assign n39294 = ~n39284 & n39293 ;
  assign n39295 = ~n39291 & n39294 ;
  assign n39304 = n28610 & ~n39034 ;
  assign n39305 = n28632 & ~n39038 ;
  assign n39306 = ~n39304 & ~n39305 ;
  assign n39307 = \P2_P2_DataWidth_reg[1]/NET0131  & ~n39306 ;
  assign n39296 = ~n28428 & ~n39023 ;
  assign n39297 = \P2_P2_InstQueue_reg[8][5]/NET0131  & ~n28027 ;
  assign n39298 = ~n28423 & n39297 ;
  assign n39299 = ~n39296 & ~n39298 ;
  assign n39308 = ~n28687 & ~n39299 ;
  assign n39309 = ~n39307 & ~n39308 ;
  assign n39310 = n26794 & ~n39309 ;
  assign n39301 = ~n26449 & n28027 ;
  assign n39302 = ~n39297 & ~n39301 ;
  assign n39303 = n27613 & ~n39302 ;
  assign n39300 = n27977 & ~n39299 ;
  assign n39311 = \P2_P2_InstQueue_reg[8][5]/NET0131  & ~n28050 ;
  assign n39312 = ~n39300 & ~n39311 ;
  assign n39313 = ~n39303 & n39312 ;
  assign n39314 = ~n39310 & n39313 ;
  assign n39323 = n28632 & ~n39034 ;
  assign n39324 = n28423 & ~n39038 ;
  assign n39325 = ~n39323 & ~n39324 ;
  assign n39326 = \P2_P2_DataWidth_reg[1]/NET0131  & ~n39325 ;
  assign n39315 = ~n28041 & ~n39023 ;
  assign n39316 = \P2_P2_InstQueue_reg[9][5]/NET0131  & ~n28034 ;
  assign n39317 = ~n28027 & n39316 ;
  assign n39318 = ~n39315 & ~n39317 ;
  assign n39327 = ~n28707 & ~n39318 ;
  assign n39328 = ~n39326 & ~n39327 ;
  assign n39329 = n26794 & ~n39328 ;
  assign n39320 = ~n26449 & n28034 ;
  assign n39321 = ~n39316 & ~n39320 ;
  assign n39322 = n27613 & ~n39321 ;
  assign n39319 = n27977 & ~n39318 ;
  assign n39330 = \P2_P2_InstQueue_reg[9][5]/NET0131  & ~n28050 ;
  assign n39331 = ~n39319 & ~n39330 ;
  assign n39332 = ~n39322 & n39331 ;
  assign n39333 = ~n39329 & n39332 ;
  assign n39339 = n25701 & n37783 ;
  assign n39340 = ~n25734 & n36590 ;
  assign n39341 = \P1_P2_PhyAddrPointer_reg[15]/NET0131  & ~n39340 ;
  assign n39342 = ~n37788 & ~n39341 ;
  assign n39343 = ~n39339 & n39342 ;
  assign n39344 = n25918 & ~n39343 ;
  assign n39334 = \P1_P2_PhyAddrPointer_reg[1]/NET0131  & n36608 ;
  assign n39335 = ~\P1_P2_PhyAddrPointer_reg[15]/NET0131  & ~n39334 ;
  assign n39336 = \P1_P2_PhyAddrPointer_reg[1]/NET0131  & n36609 ;
  assign n39337 = ~n39335 & ~n39336 ;
  assign n39345 = ~\P1_P2_DataWidth_reg[1]/NET0131  & ~n39337 ;
  assign n39346 = ~\P1_P2_PhyAddrPointer_reg[15]/NET0131  & ~n36608 ;
  assign n39347 = ~n36609 & ~n39346 ;
  assign n39348 = \P1_P2_DataWidth_reg[1]/NET0131  & ~n39347 ;
  assign n39349 = n25928 & ~n39348 ;
  assign n39350 = ~n39345 & n39349 ;
  assign n39338 = n27898 & n39337 ;
  assign n39351 = ~n25417 & ~n25921 ;
  assign n39352 = ~n27607 & n39351 ;
  assign n39353 = \P1_P2_PhyAddrPointer_reg[15]/NET0131  & ~n39352 ;
  assign n39354 = ~n37771 & ~n39353 ;
  assign n39355 = ~n39338 & n39354 ;
  assign n39356 = ~n39350 & n39355 ;
  assign n39357 = ~n39344 & n39356 ;
  assign n39358 = n25701 & n35086 ;
  assign n39359 = \P1_P2_PhyAddrPointer_reg[23]/NET0131  & ~n39340 ;
  assign n39360 = ~n35093 & ~n39359 ;
  assign n39361 = ~n39358 & n39360 ;
  assign n39362 = n25918 & ~n39361 ;
  assign n39369 = \P1_P2_PhyAddrPointer_reg[1]/NET0131  & n36613 ;
  assign n39370 = \P1_P2_PhyAddrPointer_reg[20]/NET0131  & n39369 ;
  assign n39371 = \P1_P2_PhyAddrPointer_reg[21]/NET0131  & n39370 ;
  assign n39372 = \P1_P2_PhyAddrPointer_reg[22]/NET0131  & n39371 ;
  assign n39373 = ~\P1_P2_PhyAddrPointer_reg[23]/NET0131  & ~n39372 ;
  assign n39374 = \P1_P2_PhyAddrPointer_reg[1]/NET0131  & n36617 ;
  assign n39375 = ~n39373 & ~n39374 ;
  assign n39376 = n27898 & n39375 ;
  assign n39363 = n36615 & ~n37915 ;
  assign n39364 = \P1_P2_PhyAddrPointer_reg[22]/NET0131  & n39363 ;
  assign n39366 = \P1_P2_PhyAddrPointer_reg[23]/NET0131  & n39364 ;
  assign n39365 = ~\P1_P2_PhyAddrPointer_reg[23]/NET0131  & ~n39364 ;
  assign n39367 = n25928 & ~n39365 ;
  assign n39368 = ~n39366 & n39367 ;
  assign n39377 = \P1_P2_PhyAddrPointer_reg[23]/NET0131  & ~n36595 ;
  assign n39378 = ~n35103 & ~n39377 ;
  assign n39379 = ~n39368 & n39378 ;
  assign n39380 = ~n39376 & n39379 ;
  assign n39381 = ~n39362 & n39380 ;
  assign n39389 = n25701 & n35121 ;
  assign n39390 = \P1_P2_PhyAddrPointer_reg[27]/NET0131  & ~n39340 ;
  assign n39391 = ~n35130 & ~n39390 ;
  assign n39392 = ~n39389 & n39391 ;
  assign n39393 = n25918 & ~n39392 ;
  assign n39382 = \P1_P2_PhyAddrPointer_reg[24]/NET0131  & n39374 ;
  assign n39383 = \P1_P2_PhyAddrPointer_reg[25]/NET0131  & n39382 ;
  assign n39384 = \P1_P2_PhyAddrPointer_reg[26]/NET0131  & n39383 ;
  assign n39385 = ~\P1_P2_PhyAddrPointer_reg[27]/NET0131  & ~n39384 ;
  assign n39386 = \P1_P2_PhyAddrPointer_reg[1]/NET0131  & n36621 ;
  assign n39387 = ~n39385 & ~n39386 ;
  assign n39394 = ~\P1_P2_DataWidth_reg[1]/NET0131  & ~n39387 ;
  assign n39395 = ~\P1_P2_PhyAddrPointer_reg[27]/NET0131  & ~n36620 ;
  assign n39396 = ~n36621 & ~n39395 ;
  assign n39397 = \P1_P2_DataWidth_reg[1]/NET0131  & ~n39396 ;
  assign n39398 = n25928 & ~n39397 ;
  assign n39399 = ~n39394 & n39398 ;
  assign n39388 = n27898 & n39387 ;
  assign n39400 = \P1_P2_PhyAddrPointer_reg[27]/NET0131  & ~n36595 ;
  assign n39401 = ~n35106 & ~n39400 ;
  assign n39402 = ~n39388 & n39401 ;
  assign n39403 = ~n39399 & n39402 ;
  assign n39404 = ~n39393 & n39403 ;
  assign n39414 = \P1_P2_PhyAddrPointer_reg[28]/NET0131  & n25733 ;
  assign n39415 = ~n35170 & ~n39414 ;
  assign n39416 = n25701 & ~n39415 ;
  assign n39417 = \P1_P2_PhyAddrPointer_reg[28]/NET0131  & ~n36590 ;
  assign n39418 = ~n35189 & ~n39417 ;
  assign n39419 = ~n39416 & n39418 ;
  assign n39420 = n25918 & ~n39419 ;
  assign n39410 = ~\P1_P2_PhyAddrPointer_reg[28]/NET0131  & ~n39386 ;
  assign n39411 = \P1_P2_PhyAddrPointer_reg[1]/NET0131  & n36622 ;
  assign n39412 = ~n39410 & ~n39411 ;
  assign n39413 = n36630 & n39412 ;
  assign n39405 = n25933 & ~n36621 ;
  assign n39406 = n36595 & ~n39405 ;
  assign n39407 = \P1_P2_PhyAddrPointer_reg[28]/NET0131  & ~n39406 ;
  assign n39408 = ~\P1_P2_PhyAddrPointer_reg[28]/NET0131  & n25933 ;
  assign n39409 = n36621 & n39408 ;
  assign n39421 = ~n35143 & ~n39409 ;
  assign n39422 = ~n39407 & n39421 ;
  assign n39423 = ~n39413 & n39422 ;
  assign n39424 = ~n39420 & n39423 ;
  assign n39425 = \P1_P2_PhyAddrPointer_reg[29]/NET0131  & n25733 ;
  assign n39426 = ~n35221 & ~n39425 ;
  assign n39427 = n25701 & ~n39426 ;
  assign n39428 = \P1_P2_PhyAddrPointer_reg[29]/NET0131  & ~n36590 ;
  assign n39429 = ~n35227 & ~n39428 ;
  assign n39430 = ~n39427 & n39429 ;
  assign n39431 = n25918 & ~n39430 ;
  assign n39437 = ~\P1_P2_PhyAddrPointer_reg[29]/NET0131  & ~n39411 ;
  assign n39438 = ~n37921 & ~n39437 ;
  assign n39439 = n36630 & n39438 ;
  assign n39432 = n25933 & ~n36622 ;
  assign n39433 = n36595 & ~n39432 ;
  assign n39434 = \P1_P2_PhyAddrPointer_reg[29]/NET0131  & ~n39433 ;
  assign n39435 = ~\P1_P2_PhyAddrPointer_reg[29]/NET0131  & n25933 ;
  assign n39436 = n36622 & n39435 ;
  assign n39440 = ~n35246 & ~n39436 ;
  assign n39441 = ~n39434 & n39440 ;
  assign n39442 = ~n39439 & n39441 ;
  assign n39443 = ~n39431 & n39442 ;
  assign n39446 = n25945 & n36930 ;
  assign n39447 = \P2_P1_PhyAddrPointer_reg[15]/NET0131  & ~n36678 ;
  assign n39448 = ~n36940 & ~n39447 ;
  assign n39449 = ~n39446 & n39448 ;
  assign n39450 = n11623 & ~n39449 ;
  assign n39453 = \P2_P1_PhyAddrPointer_reg[10]/NET0131  & \P2_P1_PhyAddrPointer_reg[11]/NET0131  ;
  assign n39454 = \P2_P1_PhyAddrPointer_reg[1]/NET0131  & n36648 ;
  assign n39455 = \P2_P1_PhyAddrPointer_reg[9]/NET0131  & n39454 ;
  assign n39456 = n39453 & n39455 ;
  assign n39457 = n36641 & n39456 ;
  assign n39458 = \P2_P1_PhyAddrPointer_reg[14]/NET0131  & n39457 ;
  assign n39459 = ~\P2_P1_PhyAddrPointer_reg[15]/NET0131  & ~n39458 ;
  assign n39460 = \P2_P1_PhyAddrPointer_reg[1]/NET0131  & n36653 ;
  assign n39461 = ~n39459 & ~n39460 ;
  assign n39462 = n36674 & n39461 ;
  assign n39444 = n27681 & ~n36653 ;
  assign n39451 = n36687 & ~n39444 ;
  assign n39452 = \P2_P1_PhyAddrPointer_reg[15]/NET0131  & ~n39451 ;
  assign n39445 = n36652 & n39444 ;
  assign n39463 = ~n36917 & ~n39445 ;
  assign n39464 = ~n39452 & n39463 ;
  assign n39465 = ~n39462 & n39464 ;
  assign n39466 = ~n39450 & n39465 ;
  assign n39467 = \P2_P1_PhyAddrPointer_reg[23]/NET0131  & n25947 ;
  assign n39468 = ~n35260 & ~n39467 ;
  assign n39469 = n25945 & ~n39468 ;
  assign n39470 = \P2_P1_PhyAddrPointer_reg[23]/NET0131  & ~n36677 ;
  assign n39471 = ~n35267 & ~n39470 ;
  assign n39472 = ~n39469 & n39471 ;
  assign n39473 = n11623 & ~n39472 ;
  assign n39480 = \P2_P1_PhyAddrPointer_reg[1]/NET0131  & n36660 ;
  assign n39481 = ~\P2_P1_PhyAddrPointer_reg[23]/NET0131  & ~n39480 ;
  assign n39482 = \P2_P1_PhyAddrPointer_reg[23]/NET0131  & n39480 ;
  assign n39483 = ~n39481 & ~n39482 ;
  assign n39484 = n11613 & n39483 ;
  assign n39474 = ~\P2_P1_DataWidth_reg[1]/NET0131  & ~\P2_P1_PhyAddrPointer_reg[1]/NET0131  ;
  assign n39475 = n36660 & ~n39474 ;
  assign n39477 = \P2_P1_PhyAddrPointer_reg[23]/NET0131  & n39475 ;
  assign n39476 = ~\P2_P1_PhyAddrPointer_reg[23]/NET0131  & ~n39475 ;
  assign n39478 = n11609 & ~n39476 ;
  assign n39479 = ~n39477 & n39478 ;
  assign n39485 = \P2_P1_PhyAddrPointer_reg[23]/NET0131  & ~n36687 ;
  assign n39486 = ~n35249 & ~n39485 ;
  assign n39487 = ~n39479 & n39486 ;
  assign n39488 = ~n39484 & n39487 ;
  assign n39489 = ~n39473 & n39488 ;
  assign n39491 = n25945 & n35290 ;
  assign n39492 = \P2_P1_PhyAddrPointer_reg[27]/NET0131  & ~n36678 ;
  assign n39493 = ~n35297 & ~n39492 ;
  assign n39494 = ~n39491 & n39493 ;
  assign n39495 = n11623 & ~n39494 ;
  assign n39496 = n36640 & n39480 ;
  assign n39497 = \P2_P1_PhyAddrPointer_reg[25]/NET0131  & n39496 ;
  assign n39498 = \P2_P1_PhyAddrPointer_reg[26]/NET0131  & n39497 ;
  assign n39499 = ~\P2_P1_PhyAddrPointer_reg[27]/NET0131  & ~n39498 ;
  assign n39500 = \P2_P1_PhyAddrPointer_reg[27]/NET0131  & n39498 ;
  assign n39501 = ~n39499 & ~n39500 ;
  assign n39502 = n36674 & n39501 ;
  assign n39503 = ~\P2_P1_PhyAddrPointer_reg[27]/NET0131  & ~n36663 ;
  assign n39504 = n27681 & ~n36664 ;
  assign n39505 = ~n39503 & n39504 ;
  assign n39490 = \P2_P1_PhyAddrPointer_reg[27]/NET0131  & ~n36687 ;
  assign n39506 = ~n35307 & ~n39490 ;
  assign n39507 = ~n39505 & n39506 ;
  assign n39508 = ~n39502 & n39507 ;
  assign n39509 = ~n39495 & n39508 ;
  assign n39510 = \P2_P1_PhyAddrPointer_reg[28]/NET0131  & n25947 ;
  assign n39511 = ~n35322 & ~n39510 ;
  assign n39512 = n25945 & ~n39511 ;
  assign n39513 = \P2_P1_PhyAddrPointer_reg[28]/NET0131  & ~n36677 ;
  assign n39514 = ~n35328 & ~n39513 ;
  assign n39515 = ~n39512 & n39514 ;
  assign n39516 = n11623 & ~n39515 ;
  assign n39521 = ~\P2_P1_PhyAddrPointer_reg[28]/NET0131  & ~n39500 ;
  assign n39522 = \P2_P1_PhyAddrPointer_reg[1]/NET0131  & n36665 ;
  assign n39523 = ~n39521 & ~n39522 ;
  assign n39524 = n36674 & n39523 ;
  assign n39517 = n36687 & ~n39504 ;
  assign n39518 = \P2_P1_PhyAddrPointer_reg[28]/NET0131  & ~n39517 ;
  assign n39519 = ~\P2_P1_PhyAddrPointer_reg[28]/NET0131  & n27681 ;
  assign n39520 = n36664 & n39519 ;
  assign n39525 = ~n35342 & ~n39520 ;
  assign n39526 = ~n39518 & n39525 ;
  assign n39527 = ~n39524 & n39526 ;
  assign n39528 = ~n39516 & n39527 ;
  assign n39529 = \P2_P1_PhyAddrPointer_reg[29]/NET0131  & n25947 ;
  assign n39530 = ~n35356 & ~n39529 ;
  assign n39531 = n25945 & ~n39530 ;
  assign n39532 = \P2_P1_PhyAddrPointer_reg[29]/NET0131  & ~n36677 ;
  assign n39533 = ~n35381 & ~n39532 ;
  assign n39534 = ~n39531 & n39533 ;
  assign n39535 = n11623 & ~n39534 ;
  assign n39539 = ~\P2_P1_PhyAddrPointer_reg[29]/NET0131  & ~n39522 ;
  assign n39540 = ~n37940 & ~n39539 ;
  assign n39541 = n36674 & n39540 ;
  assign n39536 = ~\P2_P1_PhyAddrPointer_reg[29]/NET0131  & ~n36665 ;
  assign n39537 = n27681 & ~n36666 ;
  assign n39538 = ~n39536 & n39537 ;
  assign n39542 = \P2_P1_PhyAddrPointer_reg[29]/NET0131  & ~n36687 ;
  assign n39543 = ~n35397 & ~n39542 ;
  assign n39544 = ~n39538 & n39543 ;
  assign n39545 = ~n39541 & n39544 ;
  assign n39546 = ~n39535 & n39545 ;
  assign n39547 = \P1_P1_PhyAddrPointer_reg[15]/NET0131  & n26249 ;
  assign n39548 = ~n37555 & ~n39547 ;
  assign n39549 = n26126 & ~n39548 ;
  assign n39550 = \P1_P1_PhyAddrPointer_reg[15]/NET0131  & ~n36696 ;
  assign n39551 = ~n37560 & ~n39550 ;
  assign n39552 = ~n39549 & n39551 ;
  assign n39553 = n8355 & ~n39552 ;
  assign n39557 = \P1_P1_PhyAddrPointer_reg[1]/NET0131  & n36711 ;
  assign n39558 = \P1_P1_PhyAddrPointer_reg[13]/NET0131  & n39557 ;
  assign n39559 = \P1_P1_PhyAddrPointer_reg[14]/NET0131  & n39558 ;
  assign n39560 = ~\P1_P1_PhyAddrPointer_reg[15]/NET0131  & ~n39559 ;
  assign n39561 = \P1_P1_PhyAddrPointer_reg[15]/NET0131  & n39559 ;
  assign n39562 = ~n39560 & ~n39561 ;
  assign n39563 = ~n36701 & n39562 ;
  assign n39554 = ~\P1_P1_PhyAddrPointer_reg[15]/NET0131  & ~n36713 ;
  assign n39555 = n27791 & ~n36714 ;
  assign n39556 = ~n39554 & n39555 ;
  assign n39564 = \P1_P1_PhyAddrPointer_reg[15]/NET0131  & ~n36743 ;
  assign n39565 = ~n37545 & ~n39564 ;
  assign n39566 = ~n39556 & n39565 ;
  assign n39567 = ~n39563 & n39566 ;
  assign n39568 = ~n39553 & n39567 ;
  assign n39581 = \P1_P1_PhyAddrPointer_reg[23]/NET0131  & n26249 ;
  assign n39582 = ~n35741 & ~n39581 ;
  assign n39583 = n26126 & ~n39582 ;
  assign n39584 = \P1_P1_PhyAddrPointer_reg[23]/NET0131  & ~n36696 ;
  assign n39585 = ~n35746 & ~n39584 ;
  assign n39586 = ~n39583 & n39585 ;
  assign n39587 = n8355 & ~n39586 ;
  assign n39576 = \P1_P1_PhyAddrPointer_reg[1]/NET0131  & n36721 ;
  assign n39577 = ~\P1_P1_PhyAddrPointer_reg[23]/NET0131  & ~n39576 ;
  assign n39578 = \P1_P1_PhyAddrPointer_reg[1]/NET0131  & n36722 ;
  assign n39579 = ~n39577 & ~n39578 ;
  assign n39580 = n8287 & n39579 ;
  assign n39569 = ~\P1_P1_DataWidth_reg[1]/NET0131  & ~\P1_P1_PhyAddrPointer_reg[1]/NET0131  ;
  assign n39570 = n36721 & ~n39569 ;
  assign n39571 = n8282 & ~n39570 ;
  assign n39572 = n36743 & ~n39571 ;
  assign n39573 = \P1_P1_PhyAddrPointer_reg[23]/NET0131  & ~n39572 ;
  assign n39574 = ~\P1_P1_PhyAddrPointer_reg[23]/NET0131  & n8282 ;
  assign n39575 = n39570 & n39574 ;
  assign n39588 = ~n35756 & ~n39575 ;
  assign n39589 = ~n39573 & n39588 ;
  assign n39590 = ~n39580 & n39589 ;
  assign n39591 = ~n39587 & n39590 ;
  assign n39592 = \P1_P1_PhyAddrPointer_reg[27]/NET0131  & n26249 ;
  assign n39593 = ~n35776 & ~n39592 ;
  assign n39594 = n26126 & ~n39593 ;
  assign n39595 = \P1_P1_PhyAddrPointer_reg[27]/NET0131  & ~n36696 ;
  assign n39596 = ~n35785 & ~n39595 ;
  assign n39597 = ~n39594 & n39596 ;
  assign n39598 = n8355 & ~n39597 ;
  assign n39602 = \P1_P1_PhyAddrPointer_reg[1]/NET0131  & n36725 ;
  assign n39603 = ~\P1_P1_PhyAddrPointer_reg[27]/NET0131  & ~n39602 ;
  assign n39604 = ~n36727 & ~n39603 ;
  assign n39605 = ~n36701 & n39604 ;
  assign n39599 = ~\P1_P1_PhyAddrPointer_reg[27]/NET0131  & ~n36725 ;
  assign n39600 = n27791 & ~n36726 ;
  assign n39601 = ~n39599 & n39600 ;
  assign n39606 = \P1_P1_PhyAddrPointer_reg[27]/NET0131  & ~n36743 ;
  assign n39607 = ~n35795 & ~n39606 ;
  assign n39608 = ~n39601 & n39607 ;
  assign n39609 = ~n39605 & n39608 ;
  assign n39610 = ~n39598 & n39609 ;
  assign n39611 = \P1_P1_PhyAddrPointer_reg[28]/NET0131  & n26249 ;
  assign n39612 = ~n35811 & ~n39611 ;
  assign n39613 = n26126 & ~n39612 ;
  assign n39614 = \P1_P1_PhyAddrPointer_reg[28]/NET0131  & ~n36696 ;
  assign n39615 = ~n35831 & ~n39614 ;
  assign n39616 = ~n39613 & n39615 ;
  assign n39617 = n8355 & ~n39616 ;
  assign n39621 = ~\P1_P1_PhyAddrPointer_reg[28]/NET0131  & ~n36727 ;
  assign n39622 = ~n36728 & ~n39621 ;
  assign n39623 = ~n36701 & n39622 ;
  assign n39618 = ~\P1_P1_PhyAddrPointer_reg[28]/NET0131  & ~n36726 ;
  assign n39619 = n27791 & ~n36735 ;
  assign n39620 = ~n39618 & n39619 ;
  assign n39624 = \P1_P1_PhyAddrPointer_reg[28]/NET0131  & ~n36743 ;
  assign n39625 = ~n35798 & ~n39624 ;
  assign n39626 = ~n39620 & n39625 ;
  assign n39627 = ~n39623 & n39626 ;
  assign n39628 = ~n39617 & n39627 ;
  assign n39629 = \P1_P1_PhyAddrPointer_reg[29]/NET0131  & n26249 ;
  assign n39630 = ~n35871 & ~n39629 ;
  assign n39631 = n26126 & ~n39630 ;
  assign n39632 = \P1_P1_PhyAddrPointer_reg[29]/NET0131  & ~n36696 ;
  assign n39633 = ~n35876 & ~n39632 ;
  assign n39634 = ~n39631 & n39633 ;
  assign n39635 = n8355 & ~n39634 ;
  assign n39639 = ~\P1_P1_PhyAddrPointer_reg[29]/NET0131  & ~n36728 ;
  assign n39640 = ~n36729 & ~n39639 ;
  assign n39641 = ~n36701 & n39640 ;
  assign n39636 = ~\P1_P1_PhyAddrPointer_reg[29]/NET0131  & ~n36735 ;
  assign n39637 = n27791 & ~n36736 ;
  assign n39638 = ~n39636 & n39637 ;
  assign n39642 = \P1_P1_PhyAddrPointer_reg[29]/NET0131  & ~n36743 ;
  assign n39643 = ~n35857 & ~n39642 ;
  assign n39644 = ~n39638 & n39643 ;
  assign n39645 = ~n39641 & n39644 ;
  assign n39646 = ~n39635 & n39645 ;
  assign n39654 = \P2_P2_PhyAddrPointer_reg[15]/NET0131  & n26629 ;
  assign n39655 = ~n37125 & ~n39654 ;
  assign n39656 = n26621 & ~n39655 ;
  assign n39657 = \P2_P2_PhyAddrPointer_reg[15]/NET0131  & ~n36752 ;
  assign n39658 = ~n37130 & ~n39657 ;
  assign n39659 = ~n39656 & n39658 ;
  assign n39660 = n26792 & ~n39659 ;
  assign n39647 = \P2_P2_PhyAddrPointer_reg[1]/NET0131  & n36770 ;
  assign n39648 = \P2_P2_PhyAddrPointer_reg[13]/NET0131  & n39647 ;
  assign n39649 = \P2_P2_PhyAddrPointer_reg[14]/NET0131  & n39648 ;
  assign n39650 = ~\P2_P2_PhyAddrPointer_reg[15]/NET0131  & ~n39649 ;
  assign n39651 = \P2_P2_PhyAddrPointer_reg[15]/NET0131  & n39649 ;
  assign n39652 = ~n39650 & ~n39651 ;
  assign n39661 = ~\P2_P2_DataWidth_reg[1]/NET0131  & ~n39652 ;
  assign n39662 = ~\P2_P2_PhyAddrPointer_reg[15]/NET0131  & ~n36772 ;
  assign n39663 = ~n36773 & ~n39662 ;
  assign n39664 = \P2_P2_DataWidth_reg[1]/NET0131  & ~n39663 ;
  assign n39665 = n26794 & ~n39664 ;
  assign n39666 = ~n39661 & n39665 ;
  assign n39653 = n27977 & n39652 ;
  assign n39667 = \P2_P2_PhyAddrPointer_reg[15]/NET0131  & ~n36758 ;
  assign n39668 = ~n37114 & ~n39667 ;
  assign n39669 = ~n39653 & n39668 ;
  assign n39670 = ~n39666 & n39669 ;
  assign n39671 = ~n39660 & n39670 ;
  assign n39672 = \P2_P2_PhyAddrPointer_reg[23]/NET0131  & n26629 ;
  assign n39673 = ~n35416 & ~n39672 ;
  assign n39674 = n26621 & ~n39673 ;
  assign n39675 = \P2_P2_PhyAddrPointer_reg[23]/NET0131  & ~n36752 ;
  assign n39676 = ~n35421 & ~n39675 ;
  assign n39677 = ~n39674 & n39676 ;
  assign n39678 = n26792 & ~n39677 ;
  assign n39682 = \P2_P2_PhyAddrPointer_reg[1]/NET0131  & n36780 ;
  assign n39683 = ~\P2_P2_PhyAddrPointer_reg[23]/NET0131  & ~n39682 ;
  assign n39684 = \P2_P2_PhyAddrPointer_reg[23]/NET0131  & n39682 ;
  assign n39685 = ~n39683 & ~n39684 ;
  assign n39686 = ~n36760 & n39685 ;
  assign n39679 = ~\P2_P2_PhyAddrPointer_reg[23]/NET0131  & ~n36780 ;
  assign n39680 = n26800 & ~n36781 ;
  assign n39681 = ~n39679 & n39680 ;
  assign n39687 = \P2_P2_PhyAddrPointer_reg[23]/NET0131  & ~n36758 ;
  assign n39688 = ~n35400 & ~n39687 ;
  assign n39689 = ~n39681 & n39688 ;
  assign n39690 = ~n39686 & n39689 ;
  assign n39691 = ~n39678 & n39690 ;
  assign n39692 = \P2_P2_PhyAddrPointer_reg[27]/NET0131  & n26629 ;
  assign n39693 = ~n35446 & ~n39692 ;
  assign n39694 = n26621 & ~n39693 ;
  assign n39695 = \P2_P2_PhyAddrPointer_reg[27]/NET0131  & ~n36752 ;
  assign n39696 = ~n39694 & ~n39695 ;
  assign n39697 = ~n35469 & n39696 ;
  assign n39698 = n26792 & ~n39697 ;
  assign n39702 = \P2_P2_PhyAddrPointer_reg[1]/NET0131  & n36783 ;
  assign n39703 = \P2_P2_PhyAddrPointer_reg[26]/NET0131  & n39702 ;
  assign n39704 = ~\P2_P2_PhyAddrPointer_reg[27]/NET0131  & ~n39703 ;
  assign n39705 = \P2_P2_PhyAddrPointer_reg[27]/NET0131  & n39703 ;
  assign n39706 = ~n39704 & ~n39705 ;
  assign n39707 = ~n36760 & n39706 ;
  assign n39699 = ~\P2_P2_PhyAddrPointer_reg[27]/NET0131  & ~n36784 ;
  assign n39700 = n26800 & ~n36785 ;
  assign n39701 = ~n39699 & n39700 ;
  assign n39708 = \P2_P2_PhyAddrPointer_reg[27]/NET0131  & ~n36758 ;
  assign n39709 = ~n35436 & ~n39708 ;
  assign n39710 = ~n39701 & n39709 ;
  assign n39711 = ~n39707 & n39710 ;
  assign n39712 = ~n39698 & n39711 ;
  assign n39713 = \P2_P2_PhyAddrPointer_reg[28]/NET0131  & n26629 ;
  assign n39714 = ~n35491 & ~n39713 ;
  assign n39715 = n26621 & ~n39714 ;
  assign n39716 = \P2_P2_PhyAddrPointer_reg[28]/NET0131  & ~n36752 ;
  assign n39717 = ~n35497 & ~n39716 ;
  assign n39718 = ~n39715 & n39717 ;
  assign n39719 = n26792 & ~n39718 ;
  assign n39723 = ~\P2_P2_PhyAddrPointer_reg[28]/NET0131  & ~n39705 ;
  assign n39724 = ~n37974 & ~n39723 ;
  assign n39725 = ~n36760 & n39724 ;
  assign n39720 = ~\P2_P2_PhyAddrPointer_reg[28]/NET0131  & ~n36785 ;
  assign n39721 = n26800 & ~n36786 ;
  assign n39722 = ~n39720 & n39721 ;
  assign n39726 = \P2_P2_PhyAddrPointer_reg[28]/NET0131  & ~n36758 ;
  assign n39727 = ~n35508 & ~n39726 ;
  assign n39728 = ~n39722 & n39727 ;
  assign n39729 = ~n39725 & n39728 ;
  assign n39730 = ~n39719 & n39729 ;
  assign n39731 = \P2_P2_PhyAddrPointer_reg[29]/NET0131  & n26629 ;
  assign n39732 = ~n35531 & ~n39731 ;
  assign n39733 = n26621 & ~n39732 ;
  assign n39734 = \P2_P2_PhyAddrPointer_reg[29]/NET0131  & ~n36752 ;
  assign n39735 = ~n35536 & ~n39734 ;
  assign n39736 = ~n39733 & n39735 ;
  assign n39737 = n26792 & ~n39736 ;
  assign n39741 = ~\P2_P2_PhyAddrPointer_reg[29]/NET0131  & ~n37974 ;
  assign n39742 = ~n37975 & ~n39741 ;
  assign n39743 = n27977 & n39742 ;
  assign n39738 = ~\P2_P2_PhyAddrPointer_reg[29]/NET0131  & ~n37980 ;
  assign n39739 = n26794 & ~n37981 ;
  assign n39740 = ~n39738 & n39739 ;
  assign n39744 = \P2_P2_PhyAddrPointer_reg[29]/NET0131  & ~n36758 ;
  assign n39745 = ~n35513 & ~n39744 ;
  assign n39746 = ~n39740 & n39745 ;
  assign n39747 = ~n39743 & n39746 ;
  assign n39748 = ~n39737 & n39747 ;
  assign n39749 = n9192 & ~n19543 ;
  assign n39750 = \P1_P3_PhyAddrPointer_reg[15]/NET0131  & ~n37992 ;
  assign n39751 = ~n19558 & ~n39750 ;
  assign n39752 = ~n39749 & n39751 ;
  assign n39753 = n9241 & ~n39752 ;
  assign n39757 = n17429 & ~n36810 ;
  assign n39754 = ~\P1_P3_PhyAddrPointer_reg[15]/NET0131  & ~n16464 ;
  assign n39755 = n11698 & ~n16465 ;
  assign n39756 = ~n39754 & n39755 ;
  assign n39758 = \P1_P3_PhyAddrPointer_reg[15]/NET0131  & ~n36816 ;
  assign n39759 = ~n19526 & ~n39758 ;
  assign n39760 = ~n39756 & n39759 ;
  assign n39761 = ~n39757 & n39760 ;
  assign n39762 = ~n39753 & n39761 ;
  assign n39769 = \P1_P3_PhyAddrPointer_reg[23]/NET0131  & n9072 ;
  assign n39770 = ~n19971 & ~n39769 ;
  assign n39771 = n9064 & ~n39770 ;
  assign n39772 = \P1_P3_PhyAddrPointer_reg[23]/NET0131  & ~n36805 ;
  assign n39773 = ~n19981 & ~n39772 ;
  assign n39774 = ~n39771 & n39773 ;
  assign n39775 = n9241 & ~n39774 ;
  assign n39768 = n16711 & ~n36810 ;
  assign n39763 = n11698 & ~n16472 ;
  assign n39764 = n36816 & ~n39763 ;
  assign n39765 = \P1_P3_PhyAddrPointer_reg[23]/NET0131  & ~n39764 ;
  assign n39766 = ~\P1_P3_PhyAddrPointer_reg[23]/NET0131  & n11698 ;
  assign n39767 = n16472 & n39766 ;
  assign n39776 = ~n19948 & ~n39767 ;
  assign n39777 = ~n39765 & n39776 ;
  assign n39778 = ~n39768 & n39777 ;
  assign n39779 = ~n39775 & n39778 ;
  assign n39786 = \P1_P3_PhyAddrPointer_reg[27]/NET0131  & n9072 ;
  assign n39787 = ~n20163 & ~n39786 ;
  assign n39788 = n9064 & ~n39787 ;
  assign n39789 = \P1_P3_PhyAddrPointer_reg[27]/NET0131  & ~n36805 ;
  assign n39790 = ~n20169 & ~n39789 ;
  assign n39791 = ~n39788 & n39790 ;
  assign n39792 = n9241 & ~n39791 ;
  assign n39785 = n16836 & ~n36810 ;
  assign n39780 = n11698 & ~n16476 ;
  assign n39781 = n36816 & ~n39780 ;
  assign n39782 = \P1_P3_PhyAddrPointer_reg[27]/NET0131  & ~n39781 ;
  assign n39783 = ~\P1_P3_PhyAddrPointer_reg[27]/NET0131  & n11698 ;
  assign n39784 = n16476 & n39783 ;
  assign n39793 = ~n20130 & ~n39784 ;
  assign n39794 = ~n39782 & n39793 ;
  assign n39795 = ~n39785 & n39794 ;
  assign n39796 = ~n39792 & n39795 ;
  assign n39797 = \P1_P3_PhyAddrPointer_reg[28]/NET0131  & n9072 ;
  assign n39798 = ~n20198 & ~n39797 ;
  assign n39799 = n9064 & ~n39798 ;
  assign n39800 = \P1_P3_PhyAddrPointer_reg[28]/NET0131  & ~n36805 ;
  assign n39801 = ~n39799 & ~n39800 ;
  assign n39802 = ~n20211 & n39801 ;
  assign n39803 = n9241 & ~n39802 ;
  assign n39807 = n16900 & ~n36810 ;
  assign n39804 = ~\P1_P3_PhyAddrPointer_reg[28]/NET0131  & ~n16477 ;
  assign n39805 = n11698 & ~n16478 ;
  assign n39806 = ~n39804 & n39805 ;
  assign n39808 = \P1_P3_PhyAddrPointer_reg[28]/NET0131  & ~n36816 ;
  assign n39809 = ~n20178 & ~n39808 ;
  assign n39810 = ~n39806 & n39809 ;
  assign n39811 = ~n39807 & n39810 ;
  assign n39812 = ~n39803 & n39811 ;
  assign n39813 = \P1_P3_PhyAddrPointer_reg[29]/NET0131  & n9072 ;
  assign n39814 = ~n20239 & ~n39813 ;
  assign n39815 = n9064 & ~n39814 ;
  assign n39816 = \P1_P3_PhyAddrPointer_reg[29]/NET0131  & ~n36805 ;
  assign n39817 = ~n20255 & ~n39816 ;
  assign n39818 = ~n39815 & n39817 ;
  assign n39819 = n9241 & ~n39818 ;
  assign n39823 = n18264 & ~n36810 ;
  assign n39820 = ~\P1_P3_PhyAddrPointer_reg[29]/NET0131  & ~n16478 ;
  assign n39821 = n11698 & ~n16479 ;
  assign n39822 = ~n39820 & n39821 ;
  assign n39824 = \P1_P3_PhyAddrPointer_reg[29]/NET0131  & ~n36816 ;
  assign n39825 = ~n20221 & ~n39824 ;
  assign n39826 = ~n39822 & n39825 ;
  assign n39827 = ~n39823 & n39826 ;
  assign n39828 = ~n39819 & n39827 ;
  assign n39830 = \P2_P3_PhyAddrPointer_reg[15]/NET0131  & ~n27283 ;
  assign n39831 = ~n37358 & ~n39830 ;
  assign n39832 = n27117 & ~n39831 ;
  assign n39833 = \P2_P3_PhyAddrPointer_reg[15]/NET0131  & ~n36826 ;
  assign n39834 = ~n37363 & ~n39833 ;
  assign n39835 = ~n39832 & n39834 ;
  assign n39836 = n27308 & ~n39835 ;
  assign n39837 = \P2_P3_PhyAddrPointer_reg[12]/NET0131  & \P2_P3_PhyAddrPointer_reg[13]/NET0131  ;
  assign n39838 = \P2_P3_PhyAddrPointer_reg[1]/NET0131  & n36840 ;
  assign n39839 = \P2_P3_PhyAddrPointer_reg[9]/NET0131  & n39838 ;
  assign n39840 = \P2_P3_PhyAddrPointer_reg[10]/NET0131  & n39839 ;
  assign n39841 = \P2_P3_PhyAddrPointer_reg[11]/NET0131  & n39840 ;
  assign n39842 = n39837 & n39841 ;
  assign n39843 = \P2_P3_PhyAddrPointer_reg[14]/NET0131  & n39842 ;
  assign n39844 = ~\P2_P3_PhyAddrPointer_reg[15]/NET0131  & ~n39843 ;
  assign n39845 = \P2_P3_PhyAddrPointer_reg[15]/NET0131  & n36846 ;
  assign n39846 = \P2_P3_PhyAddrPointer_reg[1]/NET0131  & n39845 ;
  assign n39847 = ~n39844 & ~n39846 ;
  assign n39848 = ~n36831 & n39847 ;
  assign n39849 = ~\P2_P3_PhyAddrPointer_reg[15]/NET0131  & ~n36846 ;
  assign n39850 = n27325 & ~n39845 ;
  assign n39851 = ~n39849 & n39850 ;
  assign n39829 = \P2_P3_PhyAddrPointer_reg[15]/NET0131  & ~n36873 ;
  assign n39852 = ~n37347 & ~n39829 ;
  assign n39853 = ~n39851 & n39852 ;
  assign n39854 = ~n39848 & n39853 ;
  assign n39855 = ~n39836 & n39854 ;
  assign n39856 = n27284 & n35567 ;
  assign n39857 = ~n27293 & n36826 ;
  assign n39858 = \P2_P3_PhyAddrPointer_reg[23]/NET0131  & ~n39857 ;
  assign n39859 = ~n35579 & ~n39858 ;
  assign n39860 = ~n39856 & n39859 ;
  assign n39861 = n27308 & ~n39860 ;
  assign n39863 = \P2_P3_PhyAddrPointer_reg[21]/NET0131  & n36852 ;
  assign n39870 = \P2_P3_PhyAddrPointer_reg[1]/NET0131  & n39863 ;
  assign n39871 = \P2_P3_PhyAddrPointer_reg[22]/NET0131  & n39870 ;
  assign n39872 = ~\P2_P3_PhyAddrPointer_reg[23]/NET0131  & ~n39871 ;
  assign n39873 = n36851 & n39843 ;
  assign n39874 = n36833 & n39873 ;
  assign n39875 = ~n39872 & ~n39874 ;
  assign n39876 = n32867 & n39875 ;
  assign n39862 = ~\P2_P3_DataWidth_reg[1]/NET0131  & ~\P2_P3_PhyAddrPointer_reg[1]/NET0131  ;
  assign n39864 = \P2_P3_PhyAddrPointer_reg[22]/NET0131  & ~n39862 ;
  assign n39865 = n39863 & n39864 ;
  assign n39867 = ~\P2_P3_PhyAddrPointer_reg[23]/NET0131  & ~n39865 ;
  assign n39866 = \P2_P3_PhyAddrPointer_reg[23]/NET0131  & n39865 ;
  assign n39868 = n27315 & ~n39866 ;
  assign n39869 = ~n39867 & n39868 ;
  assign n39877 = \P2_P3_PhyAddrPointer_reg[23]/NET0131  & ~n36873 ;
  assign n39878 = ~n35545 & ~n39877 ;
  assign n39879 = ~n39869 & n39878 ;
  assign n39880 = ~n39876 & n39879 ;
  assign n39881 = ~n39861 & n39880 ;
  assign n39890 = \P2_P3_PhyAddrPointer_reg[27]/NET0131  & ~n27283 ;
  assign n39891 = ~n35617 & ~n39890 ;
  assign n39892 = n27117 & ~n39891 ;
  assign n39893 = \P2_P3_PhyAddrPointer_reg[27]/NET0131  & ~n36826 ;
  assign n39894 = ~n35624 & ~n39893 ;
  assign n39895 = ~n39892 & n39894 ;
  assign n39896 = n27308 & ~n39895 ;
  assign n39885 = \P2_P3_PhyAddrPointer_reg[1]/NET0131  & n36855 ;
  assign n39886 = ~\P2_P3_PhyAddrPointer_reg[27]/NET0131  & ~n39885 ;
  assign n39887 = ~n36857 & ~n39886 ;
  assign n39888 = ~n36831 & n39887 ;
  assign n39882 = ~\P2_P3_PhyAddrPointer_reg[27]/NET0131  & ~n36855 ;
  assign n39883 = n27325 & ~n36856 ;
  assign n39884 = ~n39882 & n39883 ;
  assign n39889 = \P2_P3_PhyAddrPointer_reg[27]/NET0131  & ~n36873 ;
  assign n39897 = ~n35599 & ~n39889 ;
  assign n39898 = ~n39884 & n39897 ;
  assign n39899 = ~n39888 & n39898 ;
  assign n39900 = ~n39896 & n39899 ;
  assign n39901 = n27284 & n35649 ;
  assign n39902 = \P2_P3_PhyAddrPointer_reg[28]/NET0131  & ~n39857 ;
  assign n39903 = ~n35670 & ~n39902 ;
  assign n39904 = ~n39901 & n39903 ;
  assign n39905 = n27308 & ~n39904 ;
  assign n39909 = ~\P2_P3_PhyAddrPointer_reg[28]/NET0131  & ~n36857 ;
  assign n39910 = ~n36858 & ~n39909 ;
  assign n39911 = ~n36831 & n39910 ;
  assign n39906 = ~\P2_P3_PhyAddrPointer_reg[28]/NET0131  & ~n36856 ;
  assign n39907 = n27325 & ~n36865 ;
  assign n39908 = ~n39906 & n39907 ;
  assign n39912 = \P2_P3_PhyAddrPointer_reg[28]/NET0131  & ~n36873 ;
  assign n39913 = ~n35682 & ~n39912 ;
  assign n39914 = ~n39908 & n39913 ;
  assign n39915 = ~n39911 & n39914 ;
  assign n39916 = ~n39905 & n39915 ;
  assign n39917 = \P2_P3_PhyAddrPointer_reg[29]/NET0131  & ~n27283 ;
  assign n39918 = ~n35696 & ~n39917 ;
  assign n39919 = n27117 & ~n39918 ;
  assign n39920 = \P2_P3_PhyAddrPointer_reg[29]/NET0131  & ~n36826 ;
  assign n39921 = ~n35703 & ~n39920 ;
  assign n39922 = ~n39919 & n39921 ;
  assign n39923 = n27308 & ~n39922 ;
  assign n39927 = ~\P2_P3_PhyAddrPointer_reg[29]/NET0131  & ~n36858 ;
  assign n39928 = ~n36859 & ~n39927 ;
  assign n39929 = ~n36831 & n39928 ;
  assign n39924 = ~\P2_P3_PhyAddrPointer_reg[29]/NET0131  & ~n36865 ;
  assign n39925 = n27325 & ~n36866 ;
  assign n39926 = ~n39924 & n39925 ;
  assign n39930 = \P2_P3_PhyAddrPointer_reg[29]/NET0131  & ~n36873 ;
  assign n39931 = ~n35713 & ~n39930 ;
  assign n39932 = ~n39926 & n39931 ;
  assign n39933 = ~n39929 & n39932 ;
  assign n39934 = ~n39923 & n39933 ;
  assign n39937 = \P2_P1_InstAddrPointer_reg[10]/NET0131  & n25947 ;
  assign n39941 = ~n31934 & n31936 ;
  assign n39942 = ~n29503 & ~n31937 ;
  assign n39943 = ~n39941 & n39942 ;
  assign n39938 = ~n31807 & ~n31810 ;
  assign n39939 = ~n31811 & ~n39938 ;
  assign n39940 = n29503 & ~n39939 ;
  assign n39944 = ~n25947 & ~n39940 ;
  assign n39945 = ~n39943 & n39944 ;
  assign n39946 = ~n39937 & ~n39945 ;
  assign n39947 = n25945 & ~n39946 ;
  assign n39948 = ~n32102 & ~n35365 ;
  assign n39949 = n25964 & ~n32103 ;
  assign n39950 = ~n39948 & n39949 ;
  assign n39953 = ~n25995 & n31936 ;
  assign n39936 = n31810 & ~n32159 ;
  assign n39951 = \P2_P1_InstAddrPointer_reg[10]/NET0131  & ~n35385 ;
  assign n39952 = n26068 & n35365 ;
  assign n39954 = ~n39951 & ~n39952 ;
  assign n39955 = ~n39936 & n39954 ;
  assign n39956 = ~n39953 & n39955 ;
  assign n39957 = ~n39950 & n39956 ;
  assign n39958 = ~n39947 & n39957 ;
  assign n39959 = n11623 & ~n39958 ;
  assign n39935 = \P2_P1_rEIP_reg[10]/NET0131  & n11616 ;
  assign n39960 = \P2_P1_InstAddrPointer_reg[10]/NET0131  & ~n32172 ;
  assign n39961 = ~n39935 & ~n39960 ;
  assign n39962 = ~n39959 & n39961 ;
  assign n39965 = \P2_P1_InstAddrPointer_reg[12]/NET0131  & n25947 ;
  assign n39971 = ~n31940 & n31943 ;
  assign n39972 = ~n29503 & ~n31944 ;
  assign n39973 = ~n39971 & n39972 ;
  assign n39966 = ~\P2_P1_InstAddrPointer_reg[12]/NET0131  & ~n31502 ;
  assign n39967 = ~n31538 & ~n39966 ;
  assign n39968 = ~n38059 & ~n39967 ;
  assign n39969 = ~n31812 & ~n39968 ;
  assign n39970 = n29503 & ~n39969 ;
  assign n39974 = ~n25947 & ~n39970 ;
  assign n39975 = ~n39973 & n39974 ;
  assign n39976 = ~n39965 & ~n39975 ;
  assign n39977 = n25945 & ~n39976 ;
  assign n39978 = ~\P2_P1_InstAddrPointer_reg[12]/NET0131  & ~n32055 ;
  assign n39979 = ~n32051 & ~n39978 ;
  assign n39980 = ~n32104 & ~n39979 ;
  assign n39981 = n25964 & ~n32105 ;
  assign n39982 = ~n39980 & n39981 ;
  assign n39964 = ~n25995 & n31943 ;
  assign n39986 = n26068 & n39979 ;
  assign n39988 = ~n39964 & ~n39986 ;
  assign n39983 = ~n25987 & ~n32055 ;
  assign n39984 = n35385 & ~n39983 ;
  assign n39985 = \P2_P1_InstAddrPointer_reg[12]/NET0131  & ~n39984 ;
  assign n39987 = ~n32159 & n39967 ;
  assign n39989 = ~n39985 & ~n39987 ;
  assign n39990 = n39988 & n39989 ;
  assign n39991 = ~n39982 & n39990 ;
  assign n39992 = ~n39977 & n39991 ;
  assign n39993 = n11623 & ~n39992 ;
  assign n39963 = \P2_P1_rEIP_reg[12]/NET0131  & n11616 ;
  assign n39994 = \P2_P1_InstAddrPointer_reg[12]/NET0131  & ~n32172 ;
  assign n39995 = ~n39963 & ~n39994 ;
  assign n39996 = ~n39993 & n39995 ;
  assign n39999 = \P2_P1_InstAddrPointer_reg[13]/NET0131  & n25947 ;
  assign n40003 = ~n31944 & n31950 ;
  assign n40004 = ~n29503 & ~n36923 ;
  assign n40005 = ~n40003 & n40004 ;
  assign n40000 = ~n31541 & ~n31812 ;
  assign n40001 = ~n31813 & ~n40000 ;
  assign n40002 = n29503 & ~n40001 ;
  assign n40006 = ~n25947 & ~n40002 ;
  assign n40007 = ~n40005 & n40006 ;
  assign n40008 = ~n39999 & ~n40007 ;
  assign n40009 = n25945 & ~n40008 ;
  assign n40010 = ~n32054 & ~n35367 ;
  assign n40011 = n25964 & ~n35368 ;
  assign n40012 = ~n40010 & n40011 ;
  assign n40015 = ~n25995 & n31950 ;
  assign n39998 = n31541 & ~n32159 ;
  assign n40013 = \P2_P1_InstAddrPointer_reg[13]/NET0131  & ~n35385 ;
  assign n40014 = n26068 & n32054 ;
  assign n40016 = ~n40013 & ~n40014 ;
  assign n40017 = ~n39998 & n40016 ;
  assign n40018 = ~n40015 & n40017 ;
  assign n40019 = ~n40012 & n40018 ;
  assign n40020 = ~n40009 & n40019 ;
  assign n40021 = n11623 & ~n40020 ;
  assign n39997 = \P2_P1_rEIP_reg[13]/NET0131  & n11616 ;
  assign n40022 = \P2_P1_InstAddrPointer_reg[13]/NET0131  & ~n32172 ;
  assign n40023 = ~n39997 & ~n40022 ;
  assign n40024 = ~n40021 & n40023 ;
  assign n40027 = \P2_P1_InstAddrPointer_reg[17]/NET0131  & n25947 ;
  assign n40031 = ~n31536 & ~n31825 ;
  assign n40032 = ~n31826 & ~n40031 ;
  assign n40033 = n29503 & ~n40032 ;
  assign n40028 = ~n31960 & ~n31968 ;
  assign n40029 = ~n29503 & ~n36960 ;
  assign n40030 = ~n40028 & n40029 ;
  assign n40034 = ~n25947 & ~n40030 ;
  assign n40035 = ~n40033 & n40034 ;
  assign n40036 = ~n40027 & ~n40035 ;
  assign n40037 = n25945 & ~n40036 ;
  assign n40038 = ~n32116 & ~n35369 ;
  assign n40039 = n25964 & ~n35370 ;
  assign n40040 = ~n40038 & n40039 ;
  assign n40043 = ~n25995 & ~n31968 ;
  assign n40026 = n31536 & ~n32159 ;
  assign n40041 = \P2_P1_InstAddrPointer_reg[17]/NET0131  & ~n35385 ;
  assign n40042 = n26068 & n32116 ;
  assign n40044 = ~n40041 & ~n40042 ;
  assign n40045 = ~n40026 & n40044 ;
  assign n40046 = ~n40043 & n40045 ;
  assign n40047 = ~n40040 & n40046 ;
  assign n40048 = ~n40037 & n40047 ;
  assign n40049 = n11623 & ~n40048 ;
  assign n40025 = \P2_P1_rEIP_reg[17]/NET0131  & n11616 ;
  assign n40050 = \P2_P1_InstAddrPointer_reg[17]/NET0131  & ~n32172 ;
  assign n40051 = ~n40025 & ~n40050 ;
  assign n40052 = ~n40049 & n40051 ;
  assign n40055 = \P2_P1_InstAddrPointer_reg[8]/NET0131  & n25947 ;
  assign n40061 = ~n31799 & ~n31803 ;
  assign n40062 = n29503 & ~n40061 ;
  assign n40063 = ~n31806 & n40062 ;
  assign n40056 = ~n29503 & ~n31892 ;
  assign n40057 = ~n31927 & n40056 ;
  assign n40058 = ~n31890 & n40057 ;
  assign n40059 = ~n29503 & n31890 ;
  assign n40060 = n31929 & n40059 ;
  assign n40064 = ~n40058 & ~n40060 ;
  assign n40065 = ~n40063 & n40064 ;
  assign n40066 = ~n25947 & ~n40065 ;
  assign n40067 = ~n40055 & ~n40066 ;
  assign n40068 = n25945 & ~n40067 ;
  assign n40069 = ~n32059 & n32100 ;
  assign n40070 = n25964 & ~n32101 ;
  assign n40071 = ~n40069 & n40070 ;
  assign n40074 = ~n25995 & n31890 ;
  assign n40054 = n31803 & ~n32159 ;
  assign n40072 = \P2_P1_InstAddrPointer_reg[8]/NET0131  & ~n35385 ;
  assign n40073 = n26068 & n32059 ;
  assign n40075 = ~n40072 & ~n40073 ;
  assign n40076 = ~n40054 & n40075 ;
  assign n40077 = ~n40074 & n40076 ;
  assign n40078 = ~n40071 & n40077 ;
  assign n40079 = ~n40068 & n40078 ;
  assign n40080 = n11623 & ~n40079 ;
  assign n40053 = \P2_P1_rEIP_reg[8]/NET0131  & n11616 ;
  assign n40081 = \P2_P1_InstAddrPointer_reg[8]/NET0131  & ~n32172 ;
  assign n40082 = ~n40053 & ~n40081 ;
  assign n40083 = ~n40080 & n40082 ;
  assign n40086 = \P1_P2_InstAddrPointer_reg[8]/NET0131  & n25733 ;
  assign n40090 = n31211 & ~n31249 ;
  assign n40091 = ~n30809 & ~n31250 ;
  assign n40092 = ~n40090 & n40091 ;
  assign n40087 = ~n30855 & n31113 ;
  assign n40088 = ~n31114 & ~n40087 ;
  assign n40089 = n30809 & ~n40088 ;
  assign n40093 = ~n25733 & ~n40089 ;
  assign n40094 = ~n40092 & n40093 ;
  assign n40095 = ~n40086 & ~n40094 ;
  assign n40096 = n25701 & ~n40095 ;
  assign n40097 = ~n31370 & n31411 ;
  assign n40098 = n25881 & ~n31412 ;
  assign n40099 = ~n40097 & n40098 ;
  assign n40102 = ~n25817 & n31211 ;
  assign n40085 = ~n25830 & n30855 ;
  assign n40100 = \P1_P2_InstAddrPointer_reg[8]/NET0131  & ~n35131 ;
  assign n40101 = n25887 & n31370 ;
  assign n40103 = ~n40100 & ~n40101 ;
  assign n40104 = ~n40085 & n40103 ;
  assign n40105 = ~n40102 & n40104 ;
  assign n40106 = ~n40099 & n40105 ;
  assign n40107 = ~n40096 & n40106 ;
  assign n40108 = n25918 & ~n40107 ;
  assign n40084 = \P1_P2_rEIP_reg[8]/NET0131  & n27967 ;
  assign n40109 = \P1_P2_InstAddrPointer_reg[8]/NET0131  & ~n31487 ;
  assign n40110 = ~n40084 & ~n40109 ;
  assign n40111 = ~n40108 & n40110 ;
  assign n40114 = \P2_P2_InstAddrPointer_reg[10]/NET0131  & n26629 ;
  assign n40118 = ~n32224 & ~n32517 ;
  assign n40119 = ~n32518 & ~n40118 ;
  assign n40120 = n32510 & ~n40119 ;
  assign n40115 = ~n32640 & n32643 ;
  assign n40116 = ~n32510 & ~n38237 ;
  assign n40117 = ~n40115 & n40116 ;
  assign n40121 = ~n26629 & ~n40117 ;
  assign n40122 = ~n40120 & n40121 ;
  assign n40123 = ~n40114 & ~n40122 ;
  assign n40124 = n26621 & ~n40123 ;
  assign n40125 = ~n32763 & ~n32805 ;
  assign n40126 = n26744 & ~n32806 ;
  assign n40127 = ~n40125 & n40126 ;
  assign n40130 = ~n26688 & n32643 ;
  assign n40113 = \P2_P2_InstAddrPointer_reg[10]/NET0131  & ~n37241 ;
  assign n40128 = ~n26764 & n32224 ;
  assign n40129 = n26757 & n32763 ;
  assign n40131 = ~n40128 & ~n40129 ;
  assign n40132 = ~n40113 & n40131 ;
  assign n40133 = ~n40130 & n40132 ;
  assign n40134 = ~n40127 & n40133 ;
  assign n40135 = ~n40124 & n40134 ;
  assign n40136 = n26792 & ~n40135 ;
  assign n40112 = \P2_P2_rEIP_reg[10]/NET0131  & n28046 ;
  assign n40137 = \P2_P2_InstAddrPointer_reg[10]/NET0131  & ~n32860 ;
  assign n40138 = ~n40112 & ~n40137 ;
  assign n40139 = ~n40136 & n40138 ;
  assign n40142 = \P2_P2_InstAddrPointer_reg[12]/NET0131  & n26629 ;
  assign n40146 = ~n34280 & ~n34281 ;
  assign n40147 = ~n34282 & ~n40146 ;
  assign n40148 = n32510 & ~n40147 ;
  assign n40143 = n32583 & ~n32647 ;
  assign n40144 = ~n32510 & ~n32648 ;
  assign n40145 = ~n40143 & n40144 ;
  assign n40149 = ~n26629 & ~n40145 ;
  assign n40150 = ~n40148 & n40149 ;
  assign n40151 = ~n40142 & ~n40150 ;
  assign n40152 = n26621 & ~n40151 ;
  assign n40155 = ~\P2_P2_InstAddrPointer_reg[12]/NET0131  & ~n38249 ;
  assign n40156 = ~n38248 & n40155 ;
  assign n40153 = ~n32762 & ~n32806 ;
  assign n40154 = n32188 & ~n40153 ;
  assign n40157 = n26744 & ~n40154 ;
  assign n40158 = ~n40156 & n40157 ;
  assign n40159 = ~n26688 & n32583 ;
  assign n40160 = ~n26583 & ~n32808 ;
  assign n40161 = n35424 & ~n40160 ;
  assign n40162 = \P2_P2_InstAddrPointer_reg[12]/NET0131  & ~n40161 ;
  assign n40141 = ~n26764 & n34280 ;
  assign n40163 = ~n32808 & ~n40155 ;
  assign n40164 = n26757 & n40163 ;
  assign n40165 = ~n40141 & ~n40164 ;
  assign n40166 = ~n40162 & n40165 ;
  assign n40167 = ~n40159 & n40166 ;
  assign n40168 = ~n40158 & n40167 ;
  assign n40169 = ~n40152 & n40168 ;
  assign n40170 = n26792 & ~n40169 ;
  assign n40140 = \P2_P2_rEIP_reg[12]/NET0131  & n28046 ;
  assign n40171 = \P2_P2_InstAddrPointer_reg[12]/NET0131  & ~n32860 ;
  assign n40172 = ~n40140 & ~n40171 ;
  assign n40173 = ~n40170 & n40172 ;
  assign n40176 = \P2_P2_InstAddrPointer_reg[13]/NET0131  & n26629 ;
  assign n40180 = ~n32220 & ~n32519 ;
  assign n40181 = ~n32520 & ~n40180 ;
  assign n40182 = n32510 & ~n40181 ;
  assign n40177 = ~n32648 & n32654 ;
  assign n40178 = ~n32510 & ~n38272 ;
  assign n40179 = ~n40177 & n40178 ;
  assign n40183 = ~n26629 & ~n40179 ;
  assign n40184 = ~n40182 & n40183 ;
  assign n40185 = ~n40176 & ~n40184 ;
  assign n40186 = n26621 & ~n40185 ;
  assign n40187 = ~n32807 & ~n32810 ;
  assign n40188 = n26744 & ~n32811 ;
  assign n40189 = ~n40187 & n40188 ;
  assign n40192 = ~n26688 & n32654 ;
  assign n40175 = \P2_P2_InstAddrPointer_reg[13]/NET0131  & ~n37241 ;
  assign n40190 = ~n26764 & n32220 ;
  assign n40191 = n26757 & n32810 ;
  assign n40193 = ~n40190 & ~n40191 ;
  assign n40194 = ~n40175 & n40193 ;
  assign n40195 = ~n40192 & n40194 ;
  assign n40196 = ~n40189 & n40195 ;
  assign n40197 = ~n40186 & n40196 ;
  assign n40198 = n26792 & ~n40197 ;
  assign n40174 = \P2_P2_rEIP_reg[13]/NET0131  & n28046 ;
  assign n40199 = \P2_P2_InstAddrPointer_reg[13]/NET0131  & ~n32860 ;
  assign n40200 = ~n40174 & ~n40199 ;
  assign n40201 = ~n40198 & n40200 ;
  assign n40206 = \P2_P2_InstAddrPointer_reg[17]/NET0131  & n26629 ;
  assign n40207 = \P2_P2_InstAddrPointer_reg[16]/NET0131  & n32522 ;
  assign n40209 = ~\P2_P2_InstAddrPointer_reg[17]/NET0131  & n40207 ;
  assign n40203 = ~\P2_P2_InstAddrPointer_reg[17]/NET0131  & ~n32523 ;
  assign n40204 = ~n38349 & ~n40203 ;
  assign n40208 = n40204 & ~n40207 ;
  assign n40210 = n32510 & ~n40208 ;
  assign n40211 = ~n40209 & n40210 ;
  assign n40212 = ~n32664 & n32667 ;
  assign n40213 = ~n32510 & ~n32668 ;
  assign n40214 = ~n40212 & n40213 ;
  assign n40215 = ~n26629 & ~n40214 ;
  assign n40216 = ~n40211 & n40215 ;
  assign n40217 = ~n40206 & ~n40216 ;
  assign n40218 = n26621 & ~n40217 ;
  assign n40219 = ~n32756 & ~n32816 ;
  assign n40220 = n26744 & ~n32817 ;
  assign n40221 = ~n40219 & n40220 ;
  assign n40222 = ~n26688 & n32667 ;
  assign n40223 = \P2_P2_InstAddrPointer_reg[17]/NET0131  & ~n37240 ;
  assign n40225 = ~\P2_P2_InstAddrPointer_reg[17]/NET0131  & n26286 ;
  assign n40226 = ~n26286 & ~n40204 ;
  assign n40227 = ~n40225 & ~n40226 ;
  assign n40228 = ~n26700 & n40227 ;
  assign n40205 = n26678 & n40204 ;
  assign n40224 = n26757 & n32756 ;
  assign n40229 = ~n40205 & ~n40224 ;
  assign n40230 = ~n40228 & n40229 ;
  assign n40231 = ~n40223 & n40230 ;
  assign n40232 = ~n40222 & n40231 ;
  assign n40233 = ~n40221 & n40232 ;
  assign n40234 = ~n40218 & n40233 ;
  assign n40235 = n26792 & ~n40234 ;
  assign n40202 = \P2_P2_rEIP_reg[17]/NET0131  & n28046 ;
  assign n40236 = \P2_P2_InstAddrPointer_reg[17]/NET0131  & ~n32860 ;
  assign n40237 = ~n40202 & ~n40236 ;
  assign n40238 = ~n40235 & n40237 ;
  assign n40242 = \P2_P2_InstAddrPointer_reg[8]/NET0131  & n26629 ;
  assign n40243 = ~n32632 & n32635 ;
  assign n40244 = ~n32636 & ~n40243 ;
  assign n40245 = ~n32510 & ~n40244 ;
  assign n40247 = ~n32479 & ~n32513 ;
  assign n40246 = \P2_P2_InstAddrPointer_reg[8]/NET0131  & n32479 ;
  assign n40248 = n32510 & ~n40246 ;
  assign n40249 = ~n40247 & n40248 ;
  assign n40250 = ~n40245 & ~n40249 ;
  assign n40251 = ~n26629 & ~n40250 ;
  assign n40252 = ~n40242 & ~n40251 ;
  assign n40253 = n26621 & ~n40252 ;
  assign n40254 = ~n32765 & n32803 ;
  assign n40255 = n26744 & ~n32804 ;
  assign n40256 = ~n40254 & n40255 ;
  assign n40241 = ~n26688 & n32635 ;
  assign n40258 = ~\P2_P2_InstAddrPointer_reg[8]/NET0131  & n26286 ;
  assign n40259 = ~n26286 & ~n32513 ;
  assign n40260 = ~n40258 & ~n40259 ;
  assign n40261 = ~n26700 & n40260 ;
  assign n40257 = \P2_P2_InstAddrPointer_reg[8]/NET0131  & ~n37239 ;
  assign n40262 = ~\P2_P2_InstAddrPointer_reg[8]/NET0131  & ~n26611 ;
  assign n40263 = n26611 & ~n32765 ;
  assign n40264 = ~n40262 & ~n40263 ;
  assign n40265 = ~n26583 & n40264 ;
  assign n40266 = n26678 & n32513 ;
  assign n40267 = ~n40265 & ~n40266 ;
  assign n40268 = ~n40257 & n40267 ;
  assign n40269 = ~n40261 & n40268 ;
  assign n40270 = ~n40241 & n40269 ;
  assign n40271 = ~n40256 & n40270 ;
  assign n40272 = ~n40253 & n40271 ;
  assign n40273 = n26792 & ~n40272 ;
  assign n40239 = \P2_P2_rEIP_reg[8]/NET0131  & n28046 ;
  assign n40240 = \P2_P2_InstAddrPointer_reg[8]/NET0131  & ~n32860 ;
  assign n40274 = ~n40239 & ~n40240 ;
  assign n40275 = ~n40273 & n40274 ;
  assign n40278 = \P1_P1_InstAddrPointer_reg[10]/NET0131  & n26249 ;
  assign n40282 = ~\P1_P1_InstAddrPointer_reg[10]/NET0131  & ~n33529 ;
  assign n40283 = ~n33896 & ~n40282 ;
  assign n40284 = \P1_P1_InstAddrPointer_reg[9]/NET0131  & n33815 ;
  assign n40285 = ~n40283 & ~n40284 ;
  assign n40286 = ~n33817 & ~n40285 ;
  assign n40287 = n29558 & ~n40286 ;
  assign n40279 = n33898 & ~n33943 ;
  assign n40280 = ~n29558 & ~n33944 ;
  assign n40281 = ~n40279 & n40280 ;
  assign n40288 = ~n26249 & ~n40281 ;
  assign n40289 = ~n40287 & n40288 ;
  assign n40290 = ~n40278 & ~n40289 ;
  assign n40291 = n26126 & ~n40290 ;
  assign n40292 = ~n34052 & ~n34097 ;
  assign n40293 = n26263 & ~n34098 ;
  assign n40294 = ~n40292 & n40293 ;
  assign n40296 = ~n26189 & n40283 ;
  assign n40297 = ~n26151 & n33898 ;
  assign n40277 = \P1_P1_InstAddrPointer_reg[10]/NET0131  & ~n35760 ;
  assign n40295 = n26192 & n34052 ;
  assign n40298 = ~n40277 & ~n40295 ;
  assign n40299 = ~n40297 & n40298 ;
  assign n40300 = ~n40296 & n40299 ;
  assign n40301 = ~n40294 & n40300 ;
  assign n40302 = ~n40291 & n40301 ;
  assign n40303 = n8355 & ~n40302 ;
  assign n40276 = \P1_P1_rEIP_reg[10]/NET0131  & n8357 ;
  assign n40304 = \P1_P1_InstAddrPointer_reg[10]/NET0131  & ~n34164 ;
  assign n40305 = ~n40276 & ~n40304 ;
  assign n40306 = ~n40303 & n40305 ;
  assign n40312 = \P1_P1_InstAddrPointer_reg[12]/NET0131  & n26249 ;
  assign n40316 = ~n33949 & n33951 ;
  assign n40317 = ~n29558 & ~n33952 ;
  assign n40318 = ~n40316 & n40317 ;
  assign n40313 = ~n35729 & ~n35730 ;
  assign n40314 = ~n33818 & ~n40313 ;
  assign n40315 = n29558 & ~n40314 ;
  assign n40319 = ~n26249 & ~n40315 ;
  assign n40320 = ~n40318 & n40319 ;
  assign n40321 = ~n40312 & ~n40320 ;
  assign n40322 = n26126 & ~n40321 ;
  assign n40308 = ~\P1_P1_InstAddrPointer_reg[12]/NET0131  & ~n38460 ;
  assign n40309 = ~n34030 & ~n40308 ;
  assign n40323 = ~n38458 & ~n40309 ;
  assign n40324 = n26263 & ~n34099 ;
  assign n40325 = ~n40323 & n40324 ;
  assign n40328 = ~n26189 & n35729 ;
  assign n40329 = ~n26151 & n33951 ;
  assign n40310 = ~n26123 & n40309 ;
  assign n40311 = n15428 & n40310 ;
  assign n40326 = n35760 & ~n40310 ;
  assign n40327 = \P1_P1_InstAddrPointer_reg[12]/NET0131  & ~n40326 ;
  assign n40330 = ~n40311 & ~n40327 ;
  assign n40331 = ~n40329 & n40330 ;
  assign n40332 = ~n40328 & n40331 ;
  assign n40333 = ~n40325 & n40332 ;
  assign n40334 = ~n40322 & n40333 ;
  assign n40335 = n8355 & ~n40334 ;
  assign n40307 = \P1_P1_rEIP_reg[12]/NET0131  & n8357 ;
  assign n40336 = \P1_P1_InstAddrPointer_reg[12]/NET0131  & ~n34164 ;
  assign n40337 = ~n40307 & ~n40336 ;
  assign n40338 = ~n40335 & n40337 ;
  assign n40341 = \P2_P3_InstAddrPointer_reg[10]/NET0131  & ~n27283 ;
  assign n40346 = ~n33248 & ~n33250 ;
  assign n40347 = ~n33251 & ~n40346 ;
  assign n40348 = n33242 & ~n40347 ;
  assign n40342 = ~n33334 & n34326 ;
  assign n40343 = n33336 & ~n40342 ;
  assign n40344 = ~n33242 & ~n34327 ;
  assign n40345 = ~n40343 & n40344 ;
  assign n40349 = n27283 & ~n40345 ;
  assign n40350 = ~n40348 & n40349 ;
  assign n40351 = ~n40341 & ~n40350 ;
  assign n40352 = n27117 & ~n40351 ;
  assign n40353 = ~n33474 & ~n33476 ;
  assign n40354 = n27280 & ~n33477 ;
  assign n40355 = ~n40353 & n40354 ;
  assign n40358 = ~n27229 & n33250 ;
  assign n40357 = ~n27142 & n33336 ;
  assign n40340 = \P2_P3_InstAddrPointer_reg[10]/NET0131  & ~n34355 ;
  assign n40356 = n27219 & n33476 ;
  assign n40359 = ~n40340 & ~n40356 ;
  assign n40360 = ~n40357 & n40359 ;
  assign n40361 = ~n40358 & n40360 ;
  assign n40362 = ~n40355 & n40361 ;
  assign n40363 = ~n40352 & n40362 ;
  assign n40364 = n27308 & ~n40363 ;
  assign n40339 = \P2_P3_rEIP_reg[10]/NET0131  & n32864 ;
  assign n40365 = \P2_P3_InstAddrPointer_reg[10]/NET0131  & ~n32870 ;
  assign n40366 = ~n40339 & ~n40365 ;
  assign n40367 = ~n40364 & n40366 ;
  assign n40370 = \P1_P1_InstAddrPointer_reg[13]/NET0131  & n26249 ;
  assign n40374 = ~n33952 & n33954 ;
  assign n40375 = ~n29558 & ~n38624 ;
  assign n40376 = ~n40374 & n40375 ;
  assign n40371 = ~n33552 & ~n33818 ;
  assign n40372 = ~n33819 & ~n40371 ;
  assign n40373 = n29558 & ~n40372 ;
  assign n40377 = ~n26249 & ~n40373 ;
  assign n40378 = ~n40376 & n40377 ;
  assign n40379 = ~n40370 & ~n40378 ;
  assign n40380 = n26126 & ~n40379 ;
  assign n40381 = ~n34050 & ~n34099 ;
  assign n40382 = n26263 & ~n34100 ;
  assign n40383 = ~n40381 & n40382 ;
  assign n40386 = ~n26189 & n33552 ;
  assign n40369 = ~n26151 & n33954 ;
  assign n40384 = n26192 & n34050 ;
  assign n40385 = \P1_P1_InstAddrPointer_reg[13]/NET0131  & ~n35760 ;
  assign n40387 = ~n40384 & ~n40385 ;
  assign n40388 = ~n40369 & n40387 ;
  assign n40389 = ~n40386 & n40388 ;
  assign n40390 = ~n40383 & n40389 ;
  assign n40391 = ~n40380 & n40390 ;
  assign n40392 = n8355 & ~n40391 ;
  assign n40368 = \P1_P1_rEIP_reg[13]/NET0131  & n8357 ;
  assign n40393 = \P1_P1_InstAddrPointer_reg[13]/NET0131  & ~n34164 ;
  assign n40394 = ~n40368 & ~n40393 ;
  assign n40395 = ~n40392 & n40394 ;
  assign n40398 = \P2_P3_InstAddrPointer_reg[12]/NET0131  & ~n27283 ;
  assign n40402 = ~n33252 & ~n35555 ;
  assign n40403 = ~n33253 & ~n40402 ;
  assign n40404 = n33242 & ~n40403 ;
  assign n40399 = n33342 & ~n34328 ;
  assign n40400 = ~n33242 & ~n34329 ;
  assign n40401 = ~n40399 & n40400 ;
  assign n40405 = n27283 & ~n40401 ;
  assign n40406 = ~n40404 & n40405 ;
  assign n40407 = ~n40398 & ~n40406 ;
  assign n40408 = n27117 & ~n40407 ;
  assign n40409 = ~\P2_P3_InstAddrPointer_reg[12]/NET0131  & ~n32882 ;
  assign n40410 = ~n32883 & ~n40409 ;
  assign n40411 = ~n33478 & ~n40410 ;
  assign n40412 = n27280 & ~n33479 ;
  assign n40413 = ~n40411 & n40412 ;
  assign n40414 = ~n27257 & ~n32917 ;
  assign n40415 = n35672 & ~n40414 ;
  assign n40416 = \P2_P3_InstAddrPointer_reg[12]/NET0131  & ~n40415 ;
  assign n40397 = ~n27229 & n35555 ;
  assign n40417 = n27219 & n40410 ;
  assign n40418 = ~n27142 & n33342 ;
  assign n40419 = ~n40417 & ~n40418 ;
  assign n40420 = ~n40397 & n40419 ;
  assign n40421 = ~n40416 & n40420 ;
  assign n40422 = ~n40413 & n40421 ;
  assign n40423 = ~n40408 & n40422 ;
  assign n40424 = n27308 & ~n40423 ;
  assign n40396 = \P2_P3_rEIP_reg[12]/NET0131  & n32864 ;
  assign n40425 = \P2_P3_InstAddrPointer_reg[12]/NET0131  & ~n32870 ;
  assign n40426 = ~n40396 & ~n40425 ;
  assign n40427 = ~n40424 & n40426 ;
  assign n40430 = \P2_P3_InstAddrPointer_reg[13]/NET0131  & ~n27283 ;
  assign n40434 = ~n32955 & ~n33253 ;
  assign n40435 = ~n33254 & ~n40434 ;
  assign n40436 = n33242 & ~n40435 ;
  assign n40431 = ~n33343 & n33346 ;
  assign n40432 = ~n33242 & ~n40431 ;
  assign n40433 = ~n38522 & n40432 ;
  assign n40437 = n27283 & ~n40433 ;
  assign n40438 = ~n40436 & n40437 ;
  assign n40439 = ~n40430 & ~n40438 ;
  assign n40440 = n27117 & ~n40439 ;
  assign n40441 = ~n33429 & ~n33479 ;
  assign n40442 = n27280 & ~n33480 ;
  assign n40443 = ~n40441 & n40442 ;
  assign n40446 = ~n27229 & n32955 ;
  assign n40445 = ~n27142 & n33346 ;
  assign n40429 = \P2_P3_InstAddrPointer_reg[13]/NET0131  & ~n34355 ;
  assign n40444 = n27219 & n33429 ;
  assign n40447 = ~n40429 & ~n40444 ;
  assign n40448 = ~n40445 & n40447 ;
  assign n40449 = ~n40446 & n40448 ;
  assign n40450 = ~n40443 & n40449 ;
  assign n40451 = ~n40440 & n40450 ;
  assign n40452 = n27308 & ~n40451 ;
  assign n40428 = \P2_P3_rEIP_reg[13]/NET0131  & n32864 ;
  assign n40453 = \P2_P3_InstAddrPointer_reg[13]/NET0131  & ~n32870 ;
  assign n40454 = ~n40428 & ~n40453 ;
  assign n40455 = ~n40452 & n40454 ;
  assign n40458 = \P2_P3_InstAddrPointer_reg[17]/NET0131  & ~n27283 ;
  assign n40462 = ~\P2_P3_InstAddrPointer_reg[17]/NET0131  & ~n32921 ;
  assign n40463 = ~n33360 & ~n40462 ;
  assign n40464 = ~n37383 & ~n40463 ;
  assign n40465 = ~n37384 & ~n40464 ;
  assign n40466 = n33242 & ~n40465 ;
  assign n40459 = ~n33359 & n33376 ;
  assign n40460 = ~n33242 & ~n40459 ;
  assign n40461 = ~n38588 & n40460 ;
  assign n40467 = n27283 & ~n40461 ;
  assign n40468 = ~n40466 & n40467 ;
  assign n40469 = ~n40458 & ~n40468 ;
  assign n40470 = n27117 & ~n40469 ;
  assign n40471 = ~n33483 & ~n33486 ;
  assign n40472 = n27280 & ~n37401 ;
  assign n40473 = ~n40471 & n40472 ;
  assign n40474 = ~n27226 & ~n32921 ;
  assign n40475 = n27229 & ~n40474 ;
  assign n40476 = n40463 & ~n40475 ;
  assign n40477 = ~n27111 & ~n32887 ;
  assign n40478 = n34355 & ~n40477 ;
  assign n40479 = \P2_P3_InstAddrPointer_reg[17]/NET0131  & ~n40478 ;
  assign n40457 = n27219 & n33486 ;
  assign n40480 = ~n27142 & n33376 ;
  assign n40481 = ~n40457 & ~n40480 ;
  assign n40482 = ~n40479 & n40481 ;
  assign n40483 = ~n40476 & n40482 ;
  assign n40484 = ~n40473 & n40483 ;
  assign n40485 = ~n40470 & n40484 ;
  assign n40486 = n27308 & ~n40485 ;
  assign n40456 = \P2_P3_rEIP_reg[17]/NET0131  & n32864 ;
  assign n40487 = \P2_P3_InstAddrPointer_reg[17]/NET0131  & ~n32870 ;
  assign n40488 = ~n40456 & ~n40487 ;
  assign n40489 = ~n40486 & n40488 ;
  assign n40492 = \P2_P3_InstAddrPointer_reg[8]/NET0131  & ~n27283 ;
  assign n40496 = n33244 & ~n33246 ;
  assign n40497 = ~n33247 & ~n40496 ;
  assign n40498 = n33242 & ~n40497 ;
  assign n40493 = n33330 & n34325 ;
  assign n40494 = ~n33242 & ~n34326 ;
  assign n40495 = ~n40493 & n40494 ;
  assign n40499 = n27283 & ~n40495 ;
  assign n40500 = ~n40498 & n40499 ;
  assign n40501 = ~n40492 & ~n40500 ;
  assign n40502 = n27117 & ~n40501 ;
  assign n40503 = ~n33431 & n33472 ;
  assign n40504 = n27280 & ~n33473 ;
  assign n40505 = ~n40503 & n40504 ;
  assign n40508 = ~n27229 & n33246 ;
  assign n40507 = ~n27142 & n33330 ;
  assign n40491 = \P2_P3_InstAddrPointer_reg[8]/NET0131  & ~n34355 ;
  assign n40506 = n27219 & n33431 ;
  assign n40509 = ~n40491 & ~n40506 ;
  assign n40510 = ~n40507 & n40509 ;
  assign n40511 = ~n40508 & n40510 ;
  assign n40512 = ~n40505 & n40511 ;
  assign n40513 = ~n40502 & n40512 ;
  assign n40514 = n27308 & ~n40513 ;
  assign n40490 = \P2_P3_rEIP_reg[8]/NET0131  & n32864 ;
  assign n40515 = \P2_P3_InstAddrPointer_reg[8]/NET0131  & ~n32870 ;
  assign n40516 = ~n40490 & ~n40515 ;
  assign n40517 = ~n40514 & n40516 ;
  assign n40520 = \P1_P1_InstAddrPointer_reg[17]/NET0131  & n26249 ;
  assign n40524 = n33883 & ~n33962 ;
  assign n40525 = ~n29558 & ~n33963 ;
  assign n40526 = ~n40524 & n40525 ;
  assign n40521 = ~n33822 & ~n33825 ;
  assign n40522 = ~n37581 & ~n40521 ;
  assign n40523 = n29558 & ~n40522 ;
  assign n40527 = ~n26249 & ~n40523 ;
  assign n40528 = ~n40526 & n40527 ;
  assign n40529 = ~n40520 & ~n40528 ;
  assign n40530 = n26126 & ~n40529 ;
  assign n40531 = ~n34103 & ~n34106 ;
  assign n40532 = n26263 & ~n34107 ;
  assign n40533 = ~n40531 & n40532 ;
  assign n40519 = ~n26151 & n33883 ;
  assign n40534 = ~n15384 & ~n33533 ;
  assign n40535 = ~n24345 & ~n40534 ;
  assign n40536 = n26252 & n40535 ;
  assign n40537 = \P1_P1_InstAddrPointer_reg[17]/NET0131  & ~n40536 ;
  assign n40540 = n26254 & ~n33825 ;
  assign n40539 = ~\P1_P1_InstAddrPointer_reg[17]/NET0131  & ~n26254 ;
  assign n40541 = ~n26160 & ~n40539 ;
  assign n40542 = ~n40540 & n40541 ;
  assign n40546 = ~n40537 & ~n40542 ;
  assign n40538 = n33825 & ~n37599 ;
  assign n40543 = ~n15428 & n34033 ;
  assign n40544 = ~n26123 & ~n40543 ;
  assign n40545 = n34106 & n40544 ;
  assign n40547 = ~n40538 & ~n40545 ;
  assign n40548 = n40546 & n40547 ;
  assign n40549 = ~n40519 & n40548 ;
  assign n40550 = ~n40533 & n40549 ;
  assign n40551 = ~n40530 & n40550 ;
  assign n40552 = n8355 & ~n40551 ;
  assign n40518 = \P1_P1_rEIP_reg[17]/NET0131  & n8357 ;
  assign n40553 = \P1_P1_InstAddrPointer_reg[17]/NET0131  & ~n34164 ;
  assign n40554 = ~n40518 & ~n40553 ;
  assign n40555 = ~n40552 & n40554 ;
  assign n40558 = \P1_P2_InstAddrPointer_reg[10]/NET0131  & n25733 ;
  assign n40562 = n31207 & ~n31251 ;
  assign n40563 = ~n30809 & ~n31252 ;
  assign n40564 = ~n40562 & n40563 ;
  assign n40559 = ~n31115 & ~n31119 ;
  assign n40560 = ~n31120 & ~n40559 ;
  assign n40561 = n30809 & ~n40560 ;
  assign n40565 = ~n25733 & ~n40561 ;
  assign n40566 = ~n40564 & n40565 ;
  assign n40567 = ~n40558 & ~n40566 ;
  assign n40568 = n25701 & ~n40567 ;
  assign n40569 = ~n31413 & ~n31416 ;
  assign n40570 = n25881 & ~n31417 ;
  assign n40571 = ~n40569 & n40570 ;
  assign n40557 = ~n25817 & n31207 ;
  assign n40572 = \P1_P2_InstAddrPointer_reg[10]/NET0131  & ~n25763 ;
  assign n40573 = n25848 & ~n40572 ;
  assign n40574 = ~n25415 & ~n31119 ;
  assign n40575 = ~\P1_P2_InstAddrPointer_reg[10]/NET0131  & n25415 ;
  assign n40576 = ~n40574 & ~n40575 ;
  assign n40577 = ~n40573 & n40576 ;
  assign n40578 = \P1_P2_InstAddrPointer_reg[10]/NET0131  & ~n34207 ;
  assign n40579 = n31119 & ~n34213 ;
  assign n40580 = ~\P1_P2_InstAddrPointer_reg[10]/NET0131  & ~n25747 ;
  assign n40581 = n25747 & ~n31416 ;
  assign n40582 = ~n40580 & ~n40581 ;
  assign n40583 = ~n25743 & n40582 ;
  assign n40584 = ~n40579 & ~n40583 ;
  assign n40585 = ~n40578 & n40584 ;
  assign n40586 = ~n40577 & n40585 ;
  assign n40587 = ~n40557 & n40586 ;
  assign n40588 = ~n40571 & n40587 ;
  assign n40589 = ~n40568 & n40588 ;
  assign n40590 = n25918 & ~n40589 ;
  assign n40556 = \P1_P2_rEIP_reg[10]/NET0131  & n27967 ;
  assign n40591 = \P1_P2_InstAddrPointer_reg[10]/NET0131  & ~n31487 ;
  assign n40592 = ~n40556 & ~n40591 ;
  assign n40593 = ~n40590 & n40592 ;
  assign n40599 = \P1_P2_InstAddrPointer_reg[12]/NET0131  & n25733 ;
  assign n40604 = ~n31255 & n31259 ;
  assign n40605 = ~n30809 & ~n31260 ;
  assign n40606 = ~n40604 & n40605 ;
  assign n40601 = ~\P1_P2_InstAddrPointer_reg[12]/NET0131  & n31121 ;
  assign n40595 = \P1_P2_InstAddrPointer_reg[12]/NET0131  & n30848 ;
  assign n40596 = ~\P1_P2_InstAddrPointer_reg[12]/NET0131  & ~n30848 ;
  assign n40597 = ~n40595 & ~n40596 ;
  assign n40600 = ~n31121 & n40597 ;
  assign n40602 = n30809 & ~n40600 ;
  assign n40603 = ~n40601 & n40602 ;
  assign n40607 = ~n25733 & ~n40603 ;
  assign n40608 = ~n40606 & n40607 ;
  assign n40609 = ~n40599 & ~n40608 ;
  assign n40610 = n25701 & ~n40609 ;
  assign n40611 = ~n31350 & ~n38860 ;
  assign n40613 = ~\P1_P2_InstAddrPointer_reg[12]/NET0131  & n40611 ;
  assign n40612 = \P1_P2_InstAddrPointer_reg[12]/NET0131  & ~n40611 ;
  assign n40614 = n25881 & ~n40612 ;
  assign n40615 = ~n40613 & n40614 ;
  assign n40616 = ~n25817 & n31259 ;
  assign n40618 = n35131 & ~n38874 ;
  assign n40619 = \P1_P2_InstAddrPointer_reg[12]/NET0131  & ~n40618 ;
  assign n40598 = ~n25830 & n40597 ;
  assign n40617 = ~\P1_P2_InstAddrPointer_reg[12]/NET0131  & n38935 ;
  assign n40620 = ~n40598 & ~n40617 ;
  assign n40621 = ~n40619 & n40620 ;
  assign n40622 = ~n40616 & n40621 ;
  assign n40623 = ~n40615 & n40622 ;
  assign n40624 = ~n40610 & n40623 ;
  assign n40625 = n25918 & ~n40624 ;
  assign n40594 = \P1_P2_rEIP_reg[12]/NET0131  & n27967 ;
  assign n40626 = \P1_P2_InstAddrPointer_reg[12]/NET0131  & ~n31487 ;
  assign n40627 = ~n40594 & ~n40626 ;
  assign n40628 = ~n40625 & n40627 ;
  assign n40631 = \P1_P2_InstAddrPointer_reg[13]/NET0131  & n25733 ;
  assign n40637 = ~n31260 & n31263 ;
  assign n40638 = ~n30809 & ~n31264 ;
  assign n40639 = ~n40637 & n40638 ;
  assign n40632 = ~\P1_P2_InstAddrPointer_reg[13]/NET0131  & ~n40595 ;
  assign n40633 = ~n31123 & ~n40632 ;
  assign n40634 = ~n35204 & ~n40633 ;
  assign n40635 = ~n35205 & ~n40634 ;
  assign n40636 = n30809 & ~n40635 ;
  assign n40640 = ~n25733 & ~n40636 ;
  assign n40641 = ~n40639 & n40640 ;
  assign n40642 = ~n40631 & ~n40641 ;
  assign n40643 = n25701 & ~n40642 ;
  assign n40644 = ~n31368 & ~n31418 ;
  assign n40645 = n25881 & ~n31419 ;
  assign n40646 = ~n40644 & n40645 ;
  assign n40647 = ~n25817 & n31263 ;
  assign n40648 = ~n25830 & n40633 ;
  assign n40630 = n25887 & n31368 ;
  assign n40649 = \P1_P2_InstAddrPointer_reg[13]/NET0131  & ~n35131 ;
  assign n40650 = ~n40630 & ~n40649 ;
  assign n40651 = ~n40648 & n40650 ;
  assign n40652 = ~n40647 & n40651 ;
  assign n40653 = ~n40646 & n40652 ;
  assign n40654 = ~n40643 & n40653 ;
  assign n40655 = n25918 & ~n40654 ;
  assign n40629 = \P1_P2_rEIP_reg[13]/NET0131  & n27967 ;
  assign n40656 = \P1_P2_InstAddrPointer_reg[13]/NET0131  & ~n31487 ;
  assign n40657 = ~n40629 & ~n40656 ;
  assign n40658 = ~n40655 & n40657 ;
  assign n40661 = \P1_P1_InstAddrPointer_reg[8]/NET0131  & n26249 ;
  assign n40665 = ~n33556 & ~n33814 ;
  assign n40666 = n29558 & ~n33815 ;
  assign n40667 = ~n40665 & n40666 ;
  assign n40662 = ~n29558 & ~n33905 ;
  assign n40663 = ~n33939 & n40662 ;
  assign n40664 = ~n33903 & n40663 ;
  assign n40668 = ~n29558 & n33903 ;
  assign n40669 = n33941 & n40668 ;
  assign n40670 = ~n40664 & ~n40669 ;
  assign n40671 = ~n40667 & n40670 ;
  assign n40672 = ~n26249 & ~n40671 ;
  assign n40673 = ~n40661 & ~n40672 ;
  assign n40674 = n26126 & ~n40673 ;
  assign n40675 = ~n34054 & n34095 ;
  assign n40676 = n26263 & ~n34096 ;
  assign n40677 = ~n40675 & n40676 ;
  assign n40680 = ~n26189 & n33556 ;
  assign n40660 = ~n26151 & n33903 ;
  assign n40678 = n26192 & n34054 ;
  assign n40679 = \P1_P1_InstAddrPointer_reg[8]/NET0131  & ~n35760 ;
  assign n40681 = ~n40678 & ~n40679 ;
  assign n40682 = ~n40660 & n40681 ;
  assign n40683 = ~n40680 & n40682 ;
  assign n40684 = ~n40677 & n40683 ;
  assign n40685 = ~n40674 & n40684 ;
  assign n40686 = n8355 & ~n40685 ;
  assign n40659 = \P1_P1_rEIP_reg[8]/NET0131  & n8357 ;
  assign n40687 = \P1_P1_InstAddrPointer_reg[8]/NET0131  & ~n34164 ;
  assign n40688 = ~n40659 & ~n40687 ;
  assign n40689 = ~n40686 & n40688 ;
  assign n40692 = \P1_P2_InstAddrPointer_reg[17]/NET0131  & n25733 ;
  assign n40700 = ~n31275 & n31281 ;
  assign n40701 = ~n30809 & ~n37819 ;
  assign n40702 = ~n40700 & n40701 ;
  assign n40693 = n31137 & n35207 ;
  assign n40695 = ~\P1_P2_InstAddrPointer_reg[17]/NET0131  & ~n30849 ;
  assign n40696 = ~n31131 & ~n40695 ;
  assign n40697 = ~n40693 & n40696 ;
  assign n40694 = ~\P1_P2_InstAddrPointer_reg[17]/NET0131  & n40693 ;
  assign n40698 = n30809 & ~n40694 ;
  assign n40699 = ~n40697 & n40698 ;
  assign n40703 = ~n25733 & ~n40699 ;
  assign n40704 = ~n40702 & n40703 ;
  assign n40705 = ~n40692 & ~n40704 ;
  assign n40706 = n25701 & ~n40705 ;
  assign n40711 = ~n31424 & ~n31427 ;
  assign n40712 = n25881 & ~n38980 ;
  assign n40713 = ~n40711 & n40712 ;
  assign n40708 = \P1_P2_InstAddrPointer_reg[17]/NET0131  & ~n36902 ;
  assign n40707 = ~n25817 & n31281 ;
  assign n40709 = n25887 & n31427 ;
  assign n40710 = ~n25830 & n40696 ;
  assign n40714 = ~n40709 & ~n40710 ;
  assign n40715 = ~n40707 & n40714 ;
  assign n40716 = ~n40708 & n40715 ;
  assign n40717 = ~n40713 & n40716 ;
  assign n40718 = ~n40706 & n40717 ;
  assign n40719 = n25918 & ~n40718 ;
  assign n40690 = \P1_P2_rEIP_reg[17]/NET0131  & n27967 ;
  assign n40691 = \P1_P2_InstAddrPointer_reg[17]/NET0131  & ~n31487 ;
  assign n40720 = ~n40690 & ~n40691 ;
  assign n40721 = ~n40719 & n40720 ;
  assign n40722 = ~\P2_P1_EAX_reg[23]/NET0131  & ~n27394 ;
  assign n40723 = ~n27395 & ~n40722 ;
  assign n40724 = n24898 & n40723 ;
  assign n40725 = ~n34410 & ~n40724 ;
  assign n40726 = ~n21081 & ~n40725 ;
  assign n40727 = \P2_P1_uWord_reg[7]/NET0131  & ~n25154 ;
  assign n40728 = ~n40726 & ~n40727 ;
  assign n40729 = n11623 & ~n40728 ;
  assign n40730 = \P2_P1_uWord_reg[7]/NET0131  & ~n24913 ;
  assign n40731 = ~n40729 & ~n40730 ;
  assign n40732 = \P1_P1_uWord_reg[7]/NET0131  & ~n24515 ;
  assign n40734 = \P1_P1_uWord_reg[7]/NET0131  & n25363 ;
  assign n40735 = ~n24133 & ~n40734 ;
  assign n40736 = n15334 & ~n40735 ;
  assign n40733 = \P1_P1_uWord_reg[7]/NET0131  & n24505 ;
  assign n40737 = ~\P1_P1_EAX_reg[23]/NET0131  & ~n25354 ;
  assign n40738 = ~n25355 & ~n40737 ;
  assign n40739 = n24503 & n40738 ;
  assign n40740 = ~n40733 & ~n40739 ;
  assign n40741 = ~n40736 & n40740 ;
  assign n40742 = n8355 & ~n40741 ;
  assign n40743 = ~n40732 & ~n40742 ;
  assign n40752 = \P1_buf2_reg[25]/NET0131  & ~n27934 ;
  assign n40753 = \P1_buf1_reg[25]/NET0131  & n27934 ;
  assign n40754 = ~n40752 & ~n40753 ;
  assign n40755 = n27945 & ~n40754 ;
  assign n40756 = \P1_buf2_reg[17]/NET0131  & ~n27934 ;
  assign n40757 = \P1_buf1_reg[17]/NET0131  & n27934 ;
  assign n40758 = ~n40756 & ~n40757 ;
  assign n40759 = n27952 & ~n40758 ;
  assign n40760 = ~n40755 & ~n40759 ;
  assign n40761 = \P1_P2_DataWidth_reg[1]/NET0131  & ~n40760 ;
  assign n40744 = \P1_buf2_reg[1]/NET0131  & ~n27934 ;
  assign n40745 = \P1_buf1_reg[1]/NET0131  & n27934 ;
  assign n40746 = ~n40744 & ~n40745 ;
  assign n40747 = ~n27905 & ~n40746 ;
  assign n40748 = \P1_P2_InstQueue_reg[11][1]/NET0131  & ~n27901 ;
  assign n40749 = ~n27904 & n40748 ;
  assign n40750 = ~n40747 & ~n40749 ;
  assign n40762 = ~n27960 & ~n40750 ;
  assign n40763 = ~n40761 & ~n40762 ;
  assign n40764 = n25928 & ~n40763 ;
  assign n40765 = ~n25635 & n27901 ;
  assign n40766 = ~n40748 & ~n40765 ;
  assign n40767 = n27608 & ~n40766 ;
  assign n40751 = n27898 & ~n40750 ;
  assign n40768 = \P1_P2_InstQueue_reg[11][1]/NET0131  & ~n27972 ;
  assign n40769 = ~n40751 & ~n40768 ;
  assign n40770 = ~n40767 & n40769 ;
  assign n40771 = ~n40764 & n40770 ;
  assign n40783 = \P2_buf2_reg[25]/NET0131  & ~n28013 ;
  assign n40784 = \P2_buf1_reg[25]/NET0131  & n28013 ;
  assign n40785 = ~n40783 & ~n40784 ;
  assign n40786 = n28027 & ~n40785 ;
  assign n40787 = \P2_buf2_reg[17]/NET0131  & ~n28013 ;
  assign n40788 = \P2_buf1_reg[17]/NET0131  & n28013 ;
  assign n40789 = ~n40787 & ~n40788 ;
  assign n40790 = n28034 & ~n40789 ;
  assign n40791 = ~n40786 & ~n40790 ;
  assign n40792 = \P2_P2_DataWidth_reg[1]/NET0131  & ~n40791 ;
  assign n40772 = \P2_buf2_reg[1]/NET0131  & ~n28013 ;
  assign n40773 = \P2_buf1_reg[1]/NET0131  & n28013 ;
  assign n40774 = ~n40772 & ~n40773 ;
  assign n40775 = ~n27984 & ~n40774 ;
  assign n40776 = \P2_P2_InstQueue_reg[11][1]/NET0131  & ~n27980 ;
  assign n40777 = ~n27983 & n40776 ;
  assign n40778 = ~n40775 & ~n40777 ;
  assign n40793 = ~n28042 & ~n40778 ;
  assign n40794 = ~n40792 & ~n40793 ;
  assign n40795 = n26794 & ~n40794 ;
  assign n40780 = ~n26512 & n27980 ;
  assign n40781 = ~n40776 & ~n40780 ;
  assign n40782 = n27613 & ~n40781 ;
  assign n40779 = n27977 & ~n40778 ;
  assign n40796 = \P2_P2_InstQueue_reg[11][1]/NET0131  & ~n28050 ;
  assign n40797 = ~n40779 & ~n40796 ;
  assign n40798 = ~n40782 & n40797 ;
  assign n40799 = ~n40795 & n40798 ;
  assign n40805 = n28065 & ~n40754 ;
  assign n40806 = n28068 & ~n40758 ;
  assign n40807 = ~n40805 & ~n40806 ;
  assign n40808 = \P1_P2_DataWidth_reg[1]/NET0131  & ~n40807 ;
  assign n40800 = ~n28058 & ~n40746 ;
  assign n40801 = \P1_P2_InstQueue_reg[0][1]/NET0131  & ~n28055 ;
  assign n40802 = ~n28057 & n40801 ;
  assign n40803 = ~n40800 & ~n40802 ;
  assign n40809 = ~n28073 & ~n40803 ;
  assign n40810 = ~n40808 & ~n40809 ;
  assign n40811 = n25928 & ~n40810 ;
  assign n40812 = ~n25635 & n28055 ;
  assign n40813 = ~n40801 & ~n40812 ;
  assign n40814 = n27608 & ~n40813 ;
  assign n40804 = n27898 & ~n40803 ;
  assign n40815 = \P1_P2_InstQueue_reg[0][1]/NET0131  & ~n27972 ;
  assign n40816 = ~n40804 & ~n40815 ;
  assign n40817 = ~n40814 & n40816 ;
  assign n40818 = ~n40811 & n40817 ;
  assign n40824 = n28090 & ~n40754 ;
  assign n40825 = n27945 & ~n40758 ;
  assign n40826 = ~n40824 & ~n40825 ;
  assign n40827 = \P1_P2_DataWidth_reg[1]/NET0131  & ~n40826 ;
  assign n40819 = ~n28084 & ~n40746 ;
  assign n40820 = \P1_P2_InstQueue_reg[10][1]/NET0131  & ~n27904 ;
  assign n40821 = ~n27952 & n40820 ;
  assign n40822 = ~n40819 & ~n40821 ;
  assign n40828 = ~n28096 & ~n40822 ;
  assign n40829 = ~n40827 & ~n40828 ;
  assign n40830 = n25928 & ~n40829 ;
  assign n40831 = ~n25635 & n27904 ;
  assign n40832 = ~n40820 & ~n40831 ;
  assign n40833 = n27608 & ~n40832 ;
  assign n40823 = n27898 & ~n40822 ;
  assign n40834 = \P1_P2_InstQueue_reg[10][1]/NET0131  & ~n27972 ;
  assign n40835 = ~n40823 & ~n40834 ;
  assign n40836 = ~n40833 & n40835 ;
  assign n40837 = ~n40830 & n40836 ;
  assign n40843 = n27952 & ~n40754 ;
  assign n40844 = n27904 & ~n40758 ;
  assign n40845 = ~n40843 & ~n40844 ;
  assign n40846 = \P1_P2_DataWidth_reg[1]/NET0131  & ~n40845 ;
  assign n40838 = ~n28109 & ~n40746 ;
  assign n40839 = \P1_P2_InstQueue_reg[12][1]/NET0131  & ~n28108 ;
  assign n40840 = ~n27901 & n40839 ;
  assign n40841 = ~n40838 & ~n40840 ;
  assign n40847 = ~n28119 & ~n40841 ;
  assign n40848 = ~n40846 & ~n40847 ;
  assign n40849 = n25928 & ~n40848 ;
  assign n40850 = ~n25635 & n28108 ;
  assign n40851 = ~n40839 & ~n40850 ;
  assign n40852 = n27608 & ~n40851 ;
  assign n40842 = n27898 & ~n40841 ;
  assign n40853 = \P1_P2_InstQueue_reg[12][1]/NET0131  & ~n27972 ;
  assign n40854 = ~n40842 & ~n40853 ;
  assign n40855 = ~n40852 & n40854 ;
  assign n40856 = ~n40849 & n40855 ;
  assign n40862 = n27904 & ~n40754 ;
  assign n40863 = n27901 & ~n40758 ;
  assign n40864 = ~n40862 & ~n40863 ;
  assign n40865 = \P1_P2_DataWidth_reg[1]/NET0131  & ~n40864 ;
  assign n40857 = ~n28130 & ~n40746 ;
  assign n40858 = \P1_P2_InstQueue_reg[13][1]/NET0131  & ~n28065 ;
  assign n40859 = ~n28108 & n40858 ;
  assign n40860 = ~n40857 & ~n40859 ;
  assign n40866 = ~n28140 & ~n40860 ;
  assign n40867 = ~n40865 & ~n40866 ;
  assign n40868 = n25928 & ~n40867 ;
  assign n40869 = ~n25635 & n28065 ;
  assign n40870 = ~n40858 & ~n40869 ;
  assign n40871 = n27608 & ~n40870 ;
  assign n40861 = n27898 & ~n40860 ;
  assign n40872 = \P1_P2_InstQueue_reg[13][1]/NET0131  & ~n27972 ;
  assign n40873 = ~n40861 & ~n40872 ;
  assign n40874 = ~n40871 & n40873 ;
  assign n40875 = ~n40868 & n40874 ;
  assign n40881 = n27901 & ~n40754 ;
  assign n40882 = n28108 & ~n40758 ;
  assign n40883 = ~n40881 & ~n40882 ;
  assign n40884 = \P1_P2_DataWidth_reg[1]/NET0131  & ~n40883 ;
  assign n40876 = ~n28072 & ~n40746 ;
  assign n40877 = \P1_P2_InstQueue_reg[14][1]/NET0131  & ~n28068 ;
  assign n40878 = ~n28065 & n40877 ;
  assign n40879 = ~n40876 & ~n40878 ;
  assign n40885 = ~n28160 & ~n40879 ;
  assign n40886 = ~n40884 & ~n40885 ;
  assign n40887 = n25928 & ~n40886 ;
  assign n40888 = ~n25635 & n28068 ;
  assign n40889 = ~n40877 & ~n40888 ;
  assign n40890 = n27608 & ~n40889 ;
  assign n40880 = n27898 & ~n40879 ;
  assign n40891 = \P1_P2_InstQueue_reg[14][1]/NET0131  & ~n27972 ;
  assign n40892 = ~n40880 & ~n40891 ;
  assign n40893 = ~n40890 & n40892 ;
  assign n40894 = ~n40887 & n40893 ;
  assign n40900 = n28108 & ~n40754 ;
  assign n40901 = n28065 & ~n40758 ;
  assign n40902 = ~n40900 & ~n40901 ;
  assign n40903 = \P1_P2_DataWidth_reg[1]/NET0131  & ~n40902 ;
  assign n40895 = ~n28171 & ~n40746 ;
  assign n40896 = \P1_P2_InstQueue_reg[15][1]/NET0131  & ~n28057 ;
  assign n40897 = ~n28068 & n40896 ;
  assign n40898 = ~n40895 & ~n40897 ;
  assign n40904 = ~n28181 & ~n40898 ;
  assign n40905 = ~n40903 & ~n40904 ;
  assign n40906 = n25928 & ~n40905 ;
  assign n40907 = ~n25635 & n28057 ;
  assign n40908 = ~n40896 & ~n40907 ;
  assign n40909 = n27608 & ~n40908 ;
  assign n40899 = n27898 & ~n40898 ;
  assign n40910 = \P1_P2_InstQueue_reg[15][1]/NET0131  & ~n27972 ;
  assign n40911 = ~n40899 & ~n40910 ;
  assign n40912 = ~n40909 & n40911 ;
  assign n40913 = ~n40906 & n40912 ;
  assign n40919 = n28068 & ~n40754 ;
  assign n40920 = n28057 & ~n40758 ;
  assign n40921 = ~n40919 & ~n40920 ;
  assign n40922 = \P1_P2_DataWidth_reg[1]/NET0131  & ~n40921 ;
  assign n40914 = ~n28193 & ~n40746 ;
  assign n40915 = \P1_P2_InstQueue_reg[1][1]/NET0131  & ~n28192 ;
  assign n40916 = ~n28055 & n40915 ;
  assign n40917 = ~n40914 & ~n40916 ;
  assign n40923 = ~n28203 & ~n40917 ;
  assign n40924 = ~n40922 & ~n40923 ;
  assign n40925 = n25928 & ~n40924 ;
  assign n40926 = ~n25635 & n28192 ;
  assign n40927 = ~n40915 & ~n40926 ;
  assign n40928 = n27608 & ~n40927 ;
  assign n40918 = n27898 & ~n40917 ;
  assign n40929 = \P1_P2_InstQueue_reg[1][1]/NET0131  & ~n27972 ;
  assign n40930 = ~n40918 & ~n40929 ;
  assign n40931 = ~n40928 & n40930 ;
  assign n40932 = ~n40925 & n40931 ;
  assign n40938 = n28057 & ~n40754 ;
  assign n40939 = n28055 & ~n40758 ;
  assign n40940 = ~n40938 & ~n40939 ;
  assign n40941 = \P1_P2_DataWidth_reg[1]/NET0131  & ~n40940 ;
  assign n40933 = ~n28215 & ~n40746 ;
  assign n40934 = \P1_P2_InstQueue_reg[2][1]/NET0131  & ~n28214 ;
  assign n40935 = ~n28192 & n40934 ;
  assign n40936 = ~n40933 & ~n40935 ;
  assign n40942 = ~n28225 & ~n40936 ;
  assign n40943 = ~n40941 & ~n40942 ;
  assign n40944 = n25928 & ~n40943 ;
  assign n40945 = ~n25635 & n28214 ;
  assign n40946 = ~n40934 & ~n40945 ;
  assign n40947 = n27608 & ~n40946 ;
  assign n40937 = n27898 & ~n40936 ;
  assign n40948 = \P1_P2_InstQueue_reg[2][1]/NET0131  & ~n27972 ;
  assign n40949 = ~n40937 & ~n40948 ;
  assign n40950 = ~n40947 & n40949 ;
  assign n40951 = ~n40944 & n40950 ;
  assign n40957 = n28055 & ~n40754 ;
  assign n40958 = n28192 & ~n40758 ;
  assign n40959 = ~n40957 & ~n40958 ;
  assign n40960 = \P1_P2_DataWidth_reg[1]/NET0131  & ~n40959 ;
  assign n40952 = ~n28237 & ~n40746 ;
  assign n40953 = \P1_P2_InstQueue_reg[3][1]/NET0131  & ~n28236 ;
  assign n40954 = ~n28214 & n40953 ;
  assign n40955 = ~n40952 & ~n40954 ;
  assign n40961 = ~n28247 & ~n40955 ;
  assign n40962 = ~n40960 & ~n40961 ;
  assign n40963 = n25928 & ~n40962 ;
  assign n40964 = ~n25635 & n28236 ;
  assign n40965 = ~n40953 & ~n40964 ;
  assign n40966 = n27608 & ~n40965 ;
  assign n40956 = n27898 & ~n40955 ;
  assign n40967 = \P1_P2_InstQueue_reg[3][1]/NET0131  & ~n27972 ;
  assign n40968 = ~n40956 & ~n40967 ;
  assign n40969 = ~n40966 & n40968 ;
  assign n40970 = ~n40963 & n40969 ;
  assign n40976 = n28192 & ~n40754 ;
  assign n40977 = n28214 & ~n40758 ;
  assign n40978 = ~n40976 & ~n40977 ;
  assign n40979 = \P1_P2_DataWidth_reg[1]/NET0131  & ~n40978 ;
  assign n40971 = ~n28259 & ~n40746 ;
  assign n40972 = \P1_P2_InstQueue_reg[4][1]/NET0131  & ~n28258 ;
  assign n40973 = ~n28236 & n40972 ;
  assign n40974 = ~n40971 & ~n40973 ;
  assign n40980 = ~n28269 & ~n40974 ;
  assign n40981 = ~n40979 & ~n40980 ;
  assign n40982 = n25928 & ~n40981 ;
  assign n40983 = ~n25635 & n28258 ;
  assign n40984 = ~n40972 & ~n40983 ;
  assign n40985 = n27608 & ~n40984 ;
  assign n40975 = n27898 & ~n40974 ;
  assign n40986 = \P1_P2_InstQueue_reg[4][1]/NET0131  & ~n27972 ;
  assign n40987 = ~n40975 & ~n40986 ;
  assign n40988 = ~n40985 & n40987 ;
  assign n40989 = ~n40982 & n40988 ;
  assign n40995 = n28214 & ~n40754 ;
  assign n40996 = n28236 & ~n40758 ;
  assign n40997 = ~n40995 & ~n40996 ;
  assign n40998 = \P1_P2_DataWidth_reg[1]/NET0131  & ~n40997 ;
  assign n40990 = ~n28281 & ~n40746 ;
  assign n40991 = \P1_P2_InstQueue_reg[5][1]/NET0131  & ~n28280 ;
  assign n40992 = ~n28258 & n40991 ;
  assign n40993 = ~n40990 & ~n40992 ;
  assign n40999 = ~n28291 & ~n40993 ;
  assign n41000 = ~n40998 & ~n40999 ;
  assign n41001 = n25928 & ~n41000 ;
  assign n41002 = ~n25635 & n28280 ;
  assign n41003 = ~n40991 & ~n41002 ;
  assign n41004 = n27608 & ~n41003 ;
  assign n40994 = n27898 & ~n40993 ;
  assign n41005 = \P1_P2_InstQueue_reg[5][1]/NET0131  & ~n27972 ;
  assign n41006 = ~n40994 & ~n41005 ;
  assign n41007 = ~n41004 & n41006 ;
  assign n41008 = ~n41001 & n41007 ;
  assign n41014 = n28236 & ~n40754 ;
  assign n41015 = n28258 & ~n40758 ;
  assign n41016 = ~n41014 & ~n41015 ;
  assign n41017 = \P1_P2_DataWidth_reg[1]/NET0131  & ~n41016 ;
  assign n41009 = ~n28303 & ~n40746 ;
  assign n41010 = \P1_P2_InstQueue_reg[6][1]/NET0131  & ~n28302 ;
  assign n41011 = ~n28280 & n41010 ;
  assign n41012 = ~n41009 & ~n41011 ;
  assign n41018 = ~n28313 & ~n41012 ;
  assign n41019 = ~n41017 & ~n41018 ;
  assign n41020 = n25928 & ~n41019 ;
  assign n41021 = ~n25635 & n28302 ;
  assign n41022 = ~n41010 & ~n41021 ;
  assign n41023 = n27608 & ~n41022 ;
  assign n41013 = n27898 & ~n41012 ;
  assign n41024 = \P1_P2_InstQueue_reg[6][1]/NET0131  & ~n27972 ;
  assign n41025 = ~n41013 & ~n41024 ;
  assign n41026 = ~n41023 & n41025 ;
  assign n41027 = ~n41020 & n41026 ;
  assign n41033 = n28258 & ~n40754 ;
  assign n41034 = n28280 & ~n40758 ;
  assign n41035 = ~n41033 & ~n41034 ;
  assign n41036 = \P1_P2_DataWidth_reg[1]/NET0131  & ~n41035 ;
  assign n41028 = ~n28324 & ~n40746 ;
  assign n41029 = \P1_P2_InstQueue_reg[7][1]/NET0131  & ~n28090 ;
  assign n41030 = ~n28302 & n41029 ;
  assign n41031 = ~n41028 & ~n41030 ;
  assign n41037 = ~n28334 & ~n41031 ;
  assign n41038 = ~n41036 & ~n41037 ;
  assign n41039 = n25928 & ~n41038 ;
  assign n41040 = ~n25635 & n28090 ;
  assign n41041 = ~n41029 & ~n41040 ;
  assign n41042 = n27608 & ~n41041 ;
  assign n41032 = n27898 & ~n41031 ;
  assign n41043 = \P1_P2_InstQueue_reg[7][1]/NET0131  & ~n27972 ;
  assign n41044 = ~n41032 & ~n41043 ;
  assign n41045 = ~n41042 & n41044 ;
  assign n41046 = ~n41039 & n41045 ;
  assign n41052 = n28280 & ~n40754 ;
  assign n41053 = n28302 & ~n40758 ;
  assign n41054 = ~n41052 & ~n41053 ;
  assign n41055 = \P1_P2_DataWidth_reg[1]/NET0131  & ~n41054 ;
  assign n41047 = ~n28095 & ~n40746 ;
  assign n41048 = \P1_P2_InstQueue_reg[8][1]/NET0131  & ~n27945 ;
  assign n41049 = ~n28090 & n41048 ;
  assign n41050 = ~n41047 & ~n41049 ;
  assign n41056 = ~n28354 & ~n41050 ;
  assign n41057 = ~n41055 & ~n41056 ;
  assign n41058 = n25928 & ~n41057 ;
  assign n41059 = ~n25635 & n27945 ;
  assign n41060 = ~n41048 & ~n41059 ;
  assign n41061 = n27608 & ~n41060 ;
  assign n41051 = n27898 & ~n41050 ;
  assign n41062 = \P1_P2_InstQueue_reg[8][1]/NET0131  & ~n27972 ;
  assign n41063 = ~n41051 & ~n41062 ;
  assign n41064 = ~n41061 & n41063 ;
  assign n41065 = ~n41058 & n41064 ;
  assign n41071 = n28302 & ~n40754 ;
  assign n41072 = n28090 & ~n40758 ;
  assign n41073 = ~n41071 & ~n41072 ;
  assign n41074 = \P1_P2_DataWidth_reg[1]/NET0131  & ~n41073 ;
  assign n41066 = ~n27959 & ~n40746 ;
  assign n41067 = \P1_P2_InstQueue_reg[9][1]/NET0131  & ~n27952 ;
  assign n41068 = ~n27945 & n41067 ;
  assign n41069 = ~n41066 & ~n41068 ;
  assign n41075 = ~n28374 & ~n41069 ;
  assign n41076 = ~n41074 & ~n41075 ;
  assign n41077 = n25928 & ~n41076 ;
  assign n41078 = ~n25635 & n27952 ;
  assign n41079 = ~n41067 & ~n41078 ;
  assign n41080 = n27608 & ~n41079 ;
  assign n41070 = n27898 & ~n41069 ;
  assign n41081 = \P1_P2_InstQueue_reg[9][1]/NET0131  & ~n27972 ;
  assign n41082 = ~n41070 & ~n41081 ;
  assign n41083 = ~n41080 & n41082 ;
  assign n41084 = ~n41077 & n41083 ;
  assign n41093 = n28398 & ~n40785 ;
  assign n41094 = n28401 & ~n40789 ;
  assign n41095 = ~n41093 & ~n41094 ;
  assign n41096 = \P2_P2_DataWidth_reg[1]/NET0131  & ~n41095 ;
  assign n41085 = ~n28388 & ~n40774 ;
  assign n41086 = \P2_P2_InstQueue_reg[0][1]/NET0131  & ~n28385 ;
  assign n41087 = ~n28387 & n41086 ;
  assign n41088 = ~n41085 & ~n41087 ;
  assign n41097 = ~n28406 & ~n41088 ;
  assign n41098 = ~n41096 & ~n41097 ;
  assign n41099 = n26794 & ~n41098 ;
  assign n41090 = ~n26512 & n28385 ;
  assign n41091 = ~n41086 & ~n41090 ;
  assign n41092 = n27613 & ~n41091 ;
  assign n41089 = n27977 & ~n41088 ;
  assign n41100 = \P2_P2_InstQueue_reg[0][1]/NET0131  & ~n28050 ;
  assign n41101 = ~n41089 & ~n41100 ;
  assign n41102 = ~n41092 & n41101 ;
  assign n41103 = ~n41099 & n41102 ;
  assign n41112 = n28423 & ~n40785 ;
  assign n41113 = n28027 & ~n40789 ;
  assign n41114 = ~n41112 & ~n41113 ;
  assign n41115 = \P2_P2_DataWidth_reg[1]/NET0131  & ~n41114 ;
  assign n41104 = ~n28414 & ~n40774 ;
  assign n41105 = \P2_P2_InstQueue_reg[10][1]/NET0131  & ~n27983 ;
  assign n41106 = ~n28034 & n41105 ;
  assign n41107 = ~n41104 & ~n41106 ;
  assign n41116 = ~n28429 & ~n41107 ;
  assign n41117 = ~n41115 & ~n41116 ;
  assign n41118 = n26794 & ~n41117 ;
  assign n41109 = ~n26512 & n27983 ;
  assign n41110 = ~n41105 & ~n41109 ;
  assign n41111 = n27613 & ~n41110 ;
  assign n41108 = n27977 & ~n41107 ;
  assign n41119 = \P2_P2_InstQueue_reg[10][1]/NET0131  & ~n28050 ;
  assign n41120 = ~n41108 & ~n41119 ;
  assign n41121 = ~n41111 & n41120 ;
  assign n41122 = ~n41118 & n41121 ;
  assign n41131 = n28034 & ~n40785 ;
  assign n41132 = n27983 & ~n40789 ;
  assign n41133 = ~n41131 & ~n41132 ;
  assign n41134 = \P2_P2_DataWidth_reg[1]/NET0131  & ~n41133 ;
  assign n41123 = ~n28439 & ~n40774 ;
  assign n41124 = \P2_P2_InstQueue_reg[12][1]/NET0131  & ~n28438 ;
  assign n41125 = ~n27980 & n41124 ;
  assign n41126 = ~n41123 & ~n41125 ;
  assign n41135 = ~n28452 & ~n41126 ;
  assign n41136 = ~n41134 & ~n41135 ;
  assign n41137 = n26794 & ~n41136 ;
  assign n41128 = ~n26512 & n28438 ;
  assign n41129 = ~n41124 & ~n41128 ;
  assign n41130 = n27613 & ~n41129 ;
  assign n41127 = n27977 & ~n41126 ;
  assign n41138 = \P2_P2_InstQueue_reg[12][1]/NET0131  & ~n28050 ;
  assign n41139 = ~n41127 & ~n41138 ;
  assign n41140 = ~n41130 & n41139 ;
  assign n41141 = ~n41137 & n41140 ;
  assign n41150 = n27983 & ~n40785 ;
  assign n41151 = n27980 & ~n40789 ;
  assign n41152 = ~n41150 & ~n41151 ;
  assign n41153 = \P2_P2_DataWidth_reg[1]/NET0131  & ~n41152 ;
  assign n41142 = ~n28460 & ~n40774 ;
  assign n41143 = \P2_P2_InstQueue_reg[13][1]/NET0131  & ~n28398 ;
  assign n41144 = ~n28438 & n41143 ;
  assign n41145 = ~n41142 & ~n41144 ;
  assign n41154 = ~n28473 & ~n41145 ;
  assign n41155 = ~n41153 & ~n41154 ;
  assign n41156 = n26794 & ~n41155 ;
  assign n41147 = ~n26512 & n28398 ;
  assign n41148 = ~n41143 & ~n41147 ;
  assign n41149 = n27613 & ~n41148 ;
  assign n41146 = n27977 & ~n41145 ;
  assign n41157 = \P2_P2_InstQueue_reg[13][1]/NET0131  & ~n28050 ;
  assign n41158 = ~n41146 & ~n41157 ;
  assign n41159 = ~n41149 & n41158 ;
  assign n41160 = ~n41156 & n41159 ;
  assign n41169 = n27980 & ~n40785 ;
  assign n41170 = n28438 & ~n40789 ;
  assign n41171 = ~n41169 & ~n41170 ;
  assign n41172 = \P2_P2_DataWidth_reg[1]/NET0131  & ~n41171 ;
  assign n41161 = ~n28405 & ~n40774 ;
  assign n41162 = \P2_P2_InstQueue_reg[14][1]/NET0131  & ~n28401 ;
  assign n41163 = ~n28398 & n41162 ;
  assign n41164 = ~n41161 & ~n41163 ;
  assign n41173 = ~n28493 & ~n41164 ;
  assign n41174 = ~n41172 & ~n41173 ;
  assign n41175 = n26794 & ~n41174 ;
  assign n41166 = ~n26512 & n28401 ;
  assign n41167 = ~n41162 & ~n41166 ;
  assign n41168 = n27613 & ~n41167 ;
  assign n41165 = n27977 & ~n41164 ;
  assign n41176 = \P2_P2_InstQueue_reg[14][1]/NET0131  & ~n28050 ;
  assign n41177 = ~n41165 & ~n41176 ;
  assign n41178 = ~n41168 & n41177 ;
  assign n41179 = ~n41175 & n41178 ;
  assign n41188 = n28438 & ~n40785 ;
  assign n41189 = n28398 & ~n40789 ;
  assign n41190 = ~n41188 & ~n41189 ;
  assign n41191 = \P2_P2_DataWidth_reg[1]/NET0131  & ~n41190 ;
  assign n41180 = ~n28501 & ~n40774 ;
  assign n41181 = \P2_P2_InstQueue_reg[15][1]/NET0131  & ~n28387 ;
  assign n41182 = ~n28401 & n41181 ;
  assign n41183 = ~n41180 & ~n41182 ;
  assign n41192 = ~n28514 & ~n41183 ;
  assign n41193 = ~n41191 & ~n41192 ;
  assign n41194 = n26794 & ~n41193 ;
  assign n41185 = ~n26512 & n28387 ;
  assign n41186 = ~n41181 & ~n41185 ;
  assign n41187 = n27613 & ~n41186 ;
  assign n41184 = n27977 & ~n41183 ;
  assign n41195 = \P2_P2_InstQueue_reg[15][1]/NET0131  & ~n28050 ;
  assign n41196 = ~n41184 & ~n41195 ;
  assign n41197 = ~n41187 & n41196 ;
  assign n41198 = ~n41194 & n41197 ;
  assign n41207 = n28401 & ~n40785 ;
  assign n41208 = n28387 & ~n40789 ;
  assign n41209 = ~n41207 & ~n41208 ;
  assign n41210 = \P2_P2_DataWidth_reg[1]/NET0131  & ~n41209 ;
  assign n41199 = ~n28523 & ~n40774 ;
  assign n41200 = \P2_P2_InstQueue_reg[1][1]/NET0131  & ~n28522 ;
  assign n41201 = ~n28385 & n41200 ;
  assign n41202 = ~n41199 & ~n41201 ;
  assign n41211 = ~n28536 & ~n41202 ;
  assign n41212 = ~n41210 & ~n41211 ;
  assign n41213 = n26794 & ~n41212 ;
  assign n41204 = ~n26512 & n28522 ;
  assign n41205 = ~n41200 & ~n41204 ;
  assign n41206 = n27613 & ~n41205 ;
  assign n41203 = n27977 & ~n41202 ;
  assign n41214 = \P2_P2_InstQueue_reg[1][1]/NET0131  & ~n28050 ;
  assign n41215 = ~n41203 & ~n41214 ;
  assign n41216 = ~n41206 & n41215 ;
  assign n41217 = ~n41213 & n41216 ;
  assign n41226 = n28387 & ~n40785 ;
  assign n41227 = n28385 & ~n40789 ;
  assign n41228 = ~n41226 & ~n41227 ;
  assign n41229 = \P2_P2_DataWidth_reg[1]/NET0131  & ~n41228 ;
  assign n41218 = ~n28545 & ~n40774 ;
  assign n41219 = \P2_P2_InstQueue_reg[2][1]/NET0131  & ~n28544 ;
  assign n41220 = ~n28522 & n41219 ;
  assign n41221 = ~n41218 & ~n41220 ;
  assign n41230 = ~n28558 & ~n41221 ;
  assign n41231 = ~n41229 & ~n41230 ;
  assign n41232 = n26794 & ~n41231 ;
  assign n41223 = ~n26512 & n28544 ;
  assign n41224 = ~n41219 & ~n41223 ;
  assign n41225 = n27613 & ~n41224 ;
  assign n41222 = n27977 & ~n41221 ;
  assign n41233 = \P2_P2_InstQueue_reg[2][1]/NET0131  & ~n28050 ;
  assign n41234 = ~n41222 & ~n41233 ;
  assign n41235 = ~n41225 & n41234 ;
  assign n41236 = ~n41232 & n41235 ;
  assign n41245 = n28385 & ~n40785 ;
  assign n41246 = n28522 & ~n40789 ;
  assign n41247 = ~n41245 & ~n41246 ;
  assign n41248 = \P2_P2_DataWidth_reg[1]/NET0131  & ~n41247 ;
  assign n41237 = ~n28567 & ~n40774 ;
  assign n41238 = \P2_P2_InstQueue_reg[3][1]/NET0131  & ~n28566 ;
  assign n41239 = ~n28544 & n41238 ;
  assign n41240 = ~n41237 & ~n41239 ;
  assign n41249 = ~n28580 & ~n41240 ;
  assign n41250 = ~n41248 & ~n41249 ;
  assign n41251 = n26794 & ~n41250 ;
  assign n41242 = ~n26512 & n28566 ;
  assign n41243 = ~n41238 & ~n41242 ;
  assign n41244 = n27613 & ~n41243 ;
  assign n41241 = n27977 & ~n41240 ;
  assign n41252 = \P2_P2_InstQueue_reg[3][1]/NET0131  & ~n28050 ;
  assign n41253 = ~n41241 & ~n41252 ;
  assign n41254 = ~n41244 & n41253 ;
  assign n41255 = ~n41251 & n41254 ;
  assign n41264 = n28522 & ~n40785 ;
  assign n41265 = n28544 & ~n40789 ;
  assign n41266 = ~n41264 & ~n41265 ;
  assign n41267 = \P2_P2_DataWidth_reg[1]/NET0131  & ~n41266 ;
  assign n41256 = ~n28589 & ~n40774 ;
  assign n41257 = \P2_P2_InstQueue_reg[4][1]/NET0131  & ~n28588 ;
  assign n41258 = ~n28566 & n41257 ;
  assign n41259 = ~n41256 & ~n41258 ;
  assign n41268 = ~n28602 & ~n41259 ;
  assign n41269 = ~n41267 & ~n41268 ;
  assign n41270 = n26794 & ~n41269 ;
  assign n41261 = ~n26512 & n28588 ;
  assign n41262 = ~n41257 & ~n41261 ;
  assign n41263 = n27613 & ~n41262 ;
  assign n41260 = n27977 & ~n41259 ;
  assign n41271 = \P2_P2_InstQueue_reg[4][1]/NET0131  & ~n28050 ;
  assign n41272 = ~n41260 & ~n41271 ;
  assign n41273 = ~n41263 & n41272 ;
  assign n41274 = ~n41270 & n41273 ;
  assign n41283 = n28544 & ~n40785 ;
  assign n41284 = n28566 & ~n40789 ;
  assign n41285 = ~n41283 & ~n41284 ;
  assign n41286 = \P2_P2_DataWidth_reg[1]/NET0131  & ~n41285 ;
  assign n41275 = ~n28611 & ~n40774 ;
  assign n41276 = \P2_P2_InstQueue_reg[5][1]/NET0131  & ~n28610 ;
  assign n41277 = ~n28588 & n41276 ;
  assign n41278 = ~n41275 & ~n41277 ;
  assign n41287 = ~n28624 & ~n41278 ;
  assign n41288 = ~n41286 & ~n41287 ;
  assign n41289 = n26794 & ~n41288 ;
  assign n41280 = ~n26512 & n28610 ;
  assign n41281 = ~n41276 & ~n41280 ;
  assign n41282 = n27613 & ~n41281 ;
  assign n41279 = n27977 & ~n41278 ;
  assign n41290 = \P2_P2_InstQueue_reg[5][1]/NET0131  & ~n28050 ;
  assign n41291 = ~n41279 & ~n41290 ;
  assign n41292 = ~n41282 & n41291 ;
  assign n41293 = ~n41289 & n41292 ;
  assign n41302 = n28566 & ~n40785 ;
  assign n41303 = n28588 & ~n40789 ;
  assign n41304 = ~n41302 & ~n41303 ;
  assign n41305 = \P2_P2_DataWidth_reg[1]/NET0131  & ~n41304 ;
  assign n41294 = ~n28633 & ~n40774 ;
  assign n41295 = \P2_P2_InstQueue_reg[6][1]/NET0131  & ~n28632 ;
  assign n41296 = ~n28610 & n41295 ;
  assign n41297 = ~n41294 & ~n41296 ;
  assign n41306 = ~n28646 & ~n41297 ;
  assign n41307 = ~n41305 & ~n41306 ;
  assign n41308 = n26794 & ~n41307 ;
  assign n41299 = ~n26512 & n28632 ;
  assign n41300 = ~n41295 & ~n41299 ;
  assign n41301 = n27613 & ~n41300 ;
  assign n41298 = n27977 & ~n41297 ;
  assign n41309 = \P2_P2_InstQueue_reg[6][1]/NET0131  & ~n28050 ;
  assign n41310 = ~n41298 & ~n41309 ;
  assign n41311 = ~n41301 & n41310 ;
  assign n41312 = ~n41308 & n41311 ;
  assign n41321 = n28588 & ~n40785 ;
  assign n41322 = n28610 & ~n40789 ;
  assign n41323 = ~n41321 & ~n41322 ;
  assign n41324 = \P2_P2_DataWidth_reg[1]/NET0131  & ~n41323 ;
  assign n41313 = ~n28654 & ~n40774 ;
  assign n41314 = \P2_P2_InstQueue_reg[7][1]/NET0131  & ~n28423 ;
  assign n41315 = ~n28632 & n41314 ;
  assign n41316 = ~n41313 & ~n41315 ;
  assign n41325 = ~n28667 & ~n41316 ;
  assign n41326 = ~n41324 & ~n41325 ;
  assign n41327 = n26794 & ~n41326 ;
  assign n41318 = ~n26512 & n28423 ;
  assign n41319 = ~n41314 & ~n41318 ;
  assign n41320 = n27613 & ~n41319 ;
  assign n41317 = n27977 & ~n41316 ;
  assign n41328 = \P2_P2_InstQueue_reg[7][1]/NET0131  & ~n28050 ;
  assign n41329 = ~n41317 & ~n41328 ;
  assign n41330 = ~n41320 & n41329 ;
  assign n41331 = ~n41327 & n41330 ;
  assign n41340 = n28610 & ~n40785 ;
  assign n41341 = n28632 & ~n40789 ;
  assign n41342 = ~n41340 & ~n41341 ;
  assign n41343 = \P2_P2_DataWidth_reg[1]/NET0131  & ~n41342 ;
  assign n41332 = ~n28428 & ~n40774 ;
  assign n41333 = \P2_P2_InstQueue_reg[8][1]/NET0131  & ~n28027 ;
  assign n41334 = ~n28423 & n41333 ;
  assign n41335 = ~n41332 & ~n41334 ;
  assign n41344 = ~n28687 & ~n41335 ;
  assign n41345 = ~n41343 & ~n41344 ;
  assign n41346 = n26794 & ~n41345 ;
  assign n41337 = ~n26512 & n28027 ;
  assign n41338 = ~n41333 & ~n41337 ;
  assign n41339 = n27613 & ~n41338 ;
  assign n41336 = n27977 & ~n41335 ;
  assign n41347 = \P2_P2_InstQueue_reg[8][1]/NET0131  & ~n28050 ;
  assign n41348 = ~n41336 & ~n41347 ;
  assign n41349 = ~n41339 & n41348 ;
  assign n41350 = ~n41346 & n41349 ;
  assign n41359 = n28632 & ~n40785 ;
  assign n41360 = n28423 & ~n40789 ;
  assign n41361 = ~n41359 & ~n41360 ;
  assign n41362 = \P2_P2_DataWidth_reg[1]/NET0131  & ~n41361 ;
  assign n41351 = ~n28041 & ~n40774 ;
  assign n41352 = \P2_P2_InstQueue_reg[9][1]/NET0131  & ~n28034 ;
  assign n41353 = ~n28027 & n41352 ;
  assign n41354 = ~n41351 & ~n41353 ;
  assign n41363 = ~n28707 & ~n41354 ;
  assign n41364 = ~n41362 & ~n41363 ;
  assign n41365 = n26794 & ~n41364 ;
  assign n41356 = ~n26512 & n28034 ;
  assign n41357 = ~n41352 & ~n41356 ;
  assign n41358 = n27613 & ~n41357 ;
  assign n41355 = n27977 & ~n41354 ;
  assign n41366 = \P2_P2_InstQueue_reg[9][1]/NET0131  & ~n28050 ;
  assign n41367 = ~n41355 & ~n41366 ;
  assign n41368 = ~n41358 & n41367 ;
  assign n41369 = ~n41365 & n41368 ;
  assign n41375 = \P1_P2_PhyAddrPointer_reg[11]/NET0131  & n25733 ;
  assign n41376 = ~n38857 & ~n41375 ;
  assign n41377 = n25701 & ~n41376 ;
  assign n41378 = \P1_P2_PhyAddrPointer_reg[11]/NET0131  & ~n36590 ;
  assign n41379 = ~n38866 & ~n41378 ;
  assign n41380 = ~n41377 & n41379 ;
  assign n41381 = n25918 & ~n41380 ;
  assign n41370 = \P1_P2_PhyAddrPointer_reg[1]/NET0131  & n36604 ;
  assign n41371 = ~\P1_P2_PhyAddrPointer_reg[11]/NET0131  & ~n41370 ;
  assign n41372 = \P1_P2_PhyAddrPointer_reg[1]/NET0131  & n36605 ;
  assign n41373 = ~n41371 & ~n41372 ;
  assign n41382 = ~\P1_P2_DataWidth_reg[1]/NET0131  & ~n41373 ;
  assign n41383 = ~\P1_P2_PhyAddrPointer_reg[11]/NET0131  & ~n36604 ;
  assign n41384 = ~n36605 & ~n41383 ;
  assign n41385 = \P1_P2_DataWidth_reg[1]/NET0131  & ~n41384 ;
  assign n41386 = n25928 & ~n41385 ;
  assign n41387 = ~n41382 & n41386 ;
  assign n41374 = n27898 & n41373 ;
  assign n41388 = \P1_P2_PhyAddrPointer_reg[11]/NET0131  & ~n39352 ;
  assign n41389 = ~n38847 & ~n41388 ;
  assign n41390 = ~n41374 & n41389 ;
  assign n41391 = ~n41387 & n41390 ;
  assign n41392 = ~n41381 & n41391 ;
  assign n41397 = n25701 & n38898 ;
  assign n41398 = \P1_P2_PhyAddrPointer_reg[14]/NET0131  & ~n39340 ;
  assign n41399 = ~n38905 & ~n41398 ;
  assign n41400 = ~n41397 & n41399 ;
  assign n41401 = n25918 & ~n41400 ;
  assign n41393 = \P1_P2_PhyAddrPointer_reg[1]/NET0131  & n36607 ;
  assign n41394 = ~\P1_P2_PhyAddrPointer_reg[14]/NET0131  & ~n41393 ;
  assign n41395 = ~n39334 & ~n41394 ;
  assign n41402 = ~\P1_P2_DataWidth_reg[1]/NET0131  & ~n41395 ;
  assign n41403 = ~\P1_P2_PhyAddrPointer_reg[14]/NET0131  & ~n36607 ;
  assign n41404 = ~n36608 & ~n41403 ;
  assign n41405 = \P1_P2_DataWidth_reg[1]/NET0131  & ~n41404 ;
  assign n41406 = n25928 & ~n41405 ;
  assign n41407 = ~n41402 & n41406 ;
  assign n41396 = n27898 & n41395 ;
  assign n41408 = \P1_P2_PhyAddrPointer_reg[14]/NET0131  & ~n39352 ;
  assign n41409 = ~n38888 & ~n41408 ;
  assign n41410 = ~n41396 & n41409 ;
  assign n41411 = ~n41407 & n41410 ;
  assign n41412 = ~n41401 & n41411 ;
  assign n41423 = \P1_P2_PhyAddrPointer_reg[19]/NET0131  & n25733 ;
  assign n41424 = ~n37826 & ~n41423 ;
  assign n41425 = n25701 & ~n41424 ;
  assign n41426 = \P1_P2_PhyAddrPointer_reg[19]/NET0131  & ~n36590 ;
  assign n41427 = ~n37838 & ~n41426 ;
  assign n41428 = ~n41425 & n41427 ;
  assign n41429 = n25918 & ~n41428 ;
  assign n41419 = n36612 & ~n37915 ;
  assign n41420 = ~\P1_P2_PhyAddrPointer_reg[19]/NET0131  & ~n41419 ;
  assign n41418 = n36613 & ~n37915 ;
  assign n41421 = n25928 & ~n41418 ;
  assign n41422 = ~n41420 & n41421 ;
  assign n41414 = \P1_P2_PhyAddrPointer_reg[1]/NET0131  & n36612 ;
  assign n41415 = ~\P1_P2_PhyAddrPointer_reg[19]/NET0131  & ~n41414 ;
  assign n41416 = ~n39369 & ~n41415 ;
  assign n41417 = n27898 & n41416 ;
  assign n41413 = \P1_P2_PhyAddrPointer_reg[19]/NET0131  & ~n36595 ;
  assign n41430 = ~n37809 & ~n41413 ;
  assign n41431 = ~n41417 & n41430 ;
  assign n41432 = ~n41422 & n41431 ;
  assign n41433 = ~n41429 & n41432 ;
  assign n41434 = n25701 & n37857 ;
  assign n41435 = \P1_P2_PhyAddrPointer_reg[20]/NET0131  & ~n39340 ;
  assign n41436 = ~n37862 & ~n41435 ;
  assign n41437 = ~n41434 & n41436 ;
  assign n41438 = n25918 & ~n41437 ;
  assign n41442 = ~\P1_P2_PhyAddrPointer_reg[20]/NET0131  & ~n39369 ;
  assign n41443 = ~n39370 & ~n41442 ;
  assign n41444 = n36630 & n41443 ;
  assign n41439 = ~\P1_P2_PhyAddrPointer_reg[20]/NET0131  & ~n36613 ;
  assign n41440 = n25933 & ~n36614 ;
  assign n41441 = ~n41439 & n41440 ;
  assign n41445 = \P1_P2_PhyAddrPointer_reg[20]/NET0131  & ~n36595 ;
  assign n41446 = ~n37847 & ~n41445 ;
  assign n41447 = ~n41441 & n41446 ;
  assign n41448 = ~n41444 & n41447 ;
  assign n41449 = ~n41438 & n41448 ;
  assign n41450 = n25701 & n37688 ;
  assign n41451 = \P1_P2_PhyAddrPointer_reg[22]/NET0131  & ~n39340 ;
  assign n41452 = ~n37693 & ~n41451 ;
  assign n41453 = ~n41450 & n41452 ;
  assign n41454 = n25918 & ~n41453 ;
  assign n41458 = ~\P1_P2_PhyAddrPointer_reg[22]/NET0131  & ~n39371 ;
  assign n41459 = ~n39372 & ~n41458 ;
  assign n41460 = n36630 & n41459 ;
  assign n41455 = ~\P1_P2_PhyAddrPointer_reg[22]/NET0131  & ~n36615 ;
  assign n41456 = n25933 & ~n36616 ;
  assign n41457 = ~n41455 & n41456 ;
  assign n41461 = \P1_P2_PhyAddrPointer_reg[22]/NET0131  & ~n36595 ;
  assign n41462 = ~n37678 & ~n41461 ;
  assign n41463 = ~n41457 & n41462 ;
  assign n41464 = ~n41460 & n41463 ;
  assign n41465 = ~n41454 & n41464 ;
  assign n41467 = n25701 & n36893 ;
  assign n41468 = \P1_P2_PhyAddrPointer_reg[24]/NET0131  & ~n39340 ;
  assign n41469 = ~n36908 & ~n41468 ;
  assign n41470 = ~n41467 & n41469 ;
  assign n41471 = n25918 & ~n41470 ;
  assign n41476 = ~\P1_P2_PhyAddrPointer_reg[24]/NET0131  & ~n39374 ;
  assign n41477 = ~n39382 & ~n41476 ;
  assign n41478 = n27898 & n41477 ;
  assign n41473 = \P1_P2_PhyAddrPointer_reg[24]/NET0131  & n39366 ;
  assign n41472 = ~\P1_P2_PhyAddrPointer_reg[24]/NET0131  & ~n39366 ;
  assign n41474 = n25928 & ~n41472 ;
  assign n41475 = ~n41473 & n41474 ;
  assign n41466 = \P1_P2_PhyAddrPointer_reg[24]/NET0131  & ~n36595 ;
  assign n41479 = ~n36880 & ~n41466 ;
  assign n41480 = ~n41475 & n41479 ;
  assign n41481 = ~n41478 & n41480 ;
  assign n41482 = ~n41471 & n41481 ;
  assign n41483 = \P1_P2_PhyAddrPointer_reg[26]/NET0131  & n25733 ;
  assign n41484 = ~n37327 & ~n41483 ;
  assign n41485 = n25701 & ~n41484 ;
  assign n41486 = \P1_P2_PhyAddrPointer_reg[26]/NET0131  & ~n36590 ;
  assign n41487 = ~n37332 & ~n41486 ;
  assign n41488 = ~n41485 & n41487 ;
  assign n41489 = n25918 & ~n41488 ;
  assign n41493 = ~\P1_P2_PhyAddrPointer_reg[26]/NET0131  & ~n39383 ;
  assign n41494 = ~n39384 & ~n41493 ;
  assign n41495 = n36630 & n41494 ;
  assign n41490 = ~\P1_P2_PhyAddrPointer_reg[26]/NET0131  & ~n36619 ;
  assign n41491 = n25933 & ~n36620 ;
  assign n41492 = ~n41490 & n41491 ;
  assign n41496 = \P1_P2_PhyAddrPointer_reg[26]/NET0131  & ~n36595 ;
  assign n41497 = ~n37344 & ~n41496 ;
  assign n41498 = ~n41492 & n41497 ;
  assign n41499 = ~n41495 & n41498 ;
  assign n41500 = ~n41489 & n41499 ;
  assign n41502 = \P2_P1_PhyAddrPointer_reg[11]/NET0131  & n25947 ;
  assign n41503 = ~n38066 & ~n41502 ;
  assign n41504 = n25945 & ~n41503 ;
  assign n41505 = \P2_P1_PhyAddrPointer_reg[11]/NET0131  & ~n36677 ;
  assign n41506 = ~n38071 & ~n41505 ;
  assign n41507 = ~n41504 & n41506 ;
  assign n41508 = n11623 & ~n41507 ;
  assign n41512 = \P2_P1_PhyAddrPointer_reg[10]/NET0131  & n39455 ;
  assign n41513 = ~\P2_P1_PhyAddrPointer_reg[11]/NET0131  & ~n41512 ;
  assign n41514 = ~n39456 & ~n41513 ;
  assign n41515 = n36674 & n41514 ;
  assign n41509 = ~\P2_P1_PhyAddrPointer_reg[11]/NET0131  & ~n36650 ;
  assign n41510 = n27681 & ~n36651 ;
  assign n41511 = ~n41509 & n41510 ;
  assign n41501 = \P2_P1_PhyAddrPointer_reg[11]/NET0131  & ~n36687 ;
  assign n41516 = ~n38053 & ~n41501 ;
  assign n41517 = ~n41511 & n41516 ;
  assign n41518 = ~n41515 & n41517 ;
  assign n41519 = ~n41508 & n41518 ;
  assign n41520 = \P2_P1_PhyAddrPointer_reg[14]/NET0131  & n25947 ;
  assign n41521 = ~n38098 & ~n41520 ;
  assign n41522 = n25945 & ~n41521 ;
  assign n41523 = \P2_P1_PhyAddrPointer_reg[14]/NET0131  & ~n36677 ;
  assign n41524 = ~n38103 & ~n41523 ;
  assign n41525 = ~n41522 & n41524 ;
  assign n41526 = n11623 & ~n41525 ;
  assign n41532 = ~\P2_P1_PhyAddrPointer_reg[14]/NET0131  & ~n39457 ;
  assign n41533 = ~n39458 & ~n41532 ;
  assign n41534 = n36674 & n41533 ;
  assign n41527 = \P2_P1_PhyAddrPointer_reg[12]/NET0131  & n36651 ;
  assign n41528 = \P2_P1_PhyAddrPointer_reg[13]/NET0131  & n41527 ;
  assign n41529 = ~\P2_P1_PhyAddrPointer_reg[14]/NET0131  & ~n41528 ;
  assign n41530 = n27681 & ~n36652 ;
  assign n41531 = ~n41529 & n41530 ;
  assign n41535 = \P2_P1_PhyAddrPointer_reg[14]/NET0131  & ~n36687 ;
  assign n41536 = ~n38086 & ~n41535 ;
  assign n41537 = ~n41531 & n41536 ;
  assign n41538 = ~n41534 & n41537 ;
  assign n41539 = ~n41526 & n41538 ;
  assign n41555 = \P2_P1_PhyAddrPointer_reg[19]/NET0131  & n25947 ;
  assign n41556 = ~n36972 & ~n41555 ;
  assign n41557 = n25945 & ~n41556 ;
  assign n41558 = \P2_P1_PhyAddrPointer_reg[19]/NET0131  & ~n36677 ;
  assign n41559 = ~n36981 & ~n41558 ;
  assign n41560 = ~n41557 & n41559 ;
  assign n41561 = n11623 & ~n41560 ;
  assign n41540 = \P2_P1_PhyAddrPointer_reg[16]/NET0131  & n36653 ;
  assign n41541 = \P2_P1_PhyAddrPointer_reg[17]/NET0131  & n41540 ;
  assign n41549 = \P2_P1_PhyAddrPointer_reg[1]/NET0131  & n41541 ;
  assign n41550 = \P2_P1_PhyAddrPointer_reg[18]/NET0131  & n41549 ;
  assign n41551 = ~\P2_P1_PhyAddrPointer_reg[19]/NET0131  & ~n41550 ;
  assign n41552 = \P2_P1_PhyAddrPointer_reg[1]/NET0131  & n36657 ;
  assign n41553 = ~n41551 & ~n41552 ;
  assign n41554 = n11613 & n41553 ;
  assign n41542 = ~n39474 & n41541 ;
  assign n41543 = \P2_P1_PhyAddrPointer_reg[18]/NET0131  & n41542 ;
  assign n41544 = n11609 & ~n41543 ;
  assign n41545 = n36687 & ~n41544 ;
  assign n41546 = \P2_P1_PhyAddrPointer_reg[19]/NET0131  & ~n41545 ;
  assign n41547 = ~\P2_P1_PhyAddrPointer_reg[19]/NET0131  & n11609 ;
  assign n41548 = n41543 & n41547 ;
  assign n41562 = ~n36955 & ~n41548 ;
  assign n41563 = ~n41546 & n41562 ;
  assign n41564 = ~n41554 & n41563 ;
  assign n41565 = ~n41561 & n41564 ;
  assign n41566 = n25945 & n37005 ;
  assign n41567 = \P2_P1_PhyAddrPointer_reg[20]/NET0131  & ~n36678 ;
  assign n41568 = ~n37010 & ~n41567 ;
  assign n41569 = ~n41566 & n41568 ;
  assign n41570 = n11623 & ~n41569 ;
  assign n41576 = ~\P2_P1_PhyAddrPointer_reg[20]/NET0131  & ~n41552 ;
  assign n41577 = \P2_P1_PhyAddrPointer_reg[20]/NET0131  & n41552 ;
  assign n41578 = ~n41576 & ~n41577 ;
  assign n41579 = n11613 & n41578 ;
  assign n41571 = n36657 & ~n39474 ;
  assign n41573 = \P2_P1_PhyAddrPointer_reg[20]/NET0131  & n41571 ;
  assign n41572 = ~\P2_P1_PhyAddrPointer_reg[20]/NET0131  & ~n41571 ;
  assign n41574 = n11609 & ~n41572 ;
  assign n41575 = ~n41573 & n41574 ;
  assign n41580 = \P2_P1_PhyAddrPointer_reg[20]/NET0131  & ~n36687 ;
  assign n41581 = ~n36994 & ~n41580 ;
  assign n41582 = ~n41575 & n41581 ;
  assign n41583 = ~n41579 & n41582 ;
  assign n41584 = ~n41570 & n41583 ;
  assign n41585 = \P2_P1_PhyAddrPointer_reg[22]/NET0131  & n25947 ;
  assign n41586 = ~n37035 & ~n41585 ;
  assign n41587 = n25945 & ~n41586 ;
  assign n41588 = \P2_P1_PhyAddrPointer_reg[22]/NET0131  & ~n36677 ;
  assign n41589 = ~n37040 & ~n41588 ;
  assign n41590 = ~n41587 & n41589 ;
  assign n41591 = n11623 & ~n41590 ;
  assign n41595 = \P2_P1_PhyAddrPointer_reg[21]/NET0131  & n41577 ;
  assign n41596 = ~\P2_P1_PhyAddrPointer_reg[22]/NET0131  & ~n41595 ;
  assign n41597 = ~n39480 & ~n41596 ;
  assign n41598 = n36674 & n41597 ;
  assign n41592 = ~\P2_P1_PhyAddrPointer_reg[22]/NET0131  & ~n36659 ;
  assign n41593 = n27681 & ~n36660 ;
  assign n41594 = ~n41592 & n41593 ;
  assign n41599 = \P2_P1_PhyAddrPointer_reg[22]/NET0131  & ~n36687 ;
  assign n41600 = ~n37025 & ~n41599 ;
  assign n41601 = ~n41594 & n41600 ;
  assign n41602 = ~n41598 & n41601 ;
  assign n41603 = ~n41591 & n41602 ;
  assign n41605 = \P2_P1_PhyAddrPointer_reg[24]/NET0131  & n25947 ;
  assign n41606 = ~n37065 & ~n41605 ;
  assign n41607 = n25945 & ~n41606 ;
  assign n41608 = \P2_P1_PhyAddrPointer_reg[24]/NET0131  & ~n36677 ;
  assign n41609 = ~n37070 & ~n41608 ;
  assign n41610 = ~n41607 & n41609 ;
  assign n41611 = n11623 & ~n41610 ;
  assign n41612 = ~\P2_P1_PhyAddrPointer_reg[24]/NET0131  & ~n39482 ;
  assign n41613 = ~n39496 & ~n41612 ;
  assign n41614 = n11613 & n41613 ;
  assign n41616 = ~\P2_P1_PhyAddrPointer_reg[24]/NET0131  & ~n39477 ;
  assign n41615 = n36661 & ~n39474 ;
  assign n41617 = n11609 & ~n41615 ;
  assign n41618 = ~n41616 & n41617 ;
  assign n41604 = \P2_P1_PhyAddrPointer_reg[24]/NET0131  & ~n36687 ;
  assign n41619 = ~n37053 & ~n41604 ;
  assign n41620 = ~n41618 & n41619 ;
  assign n41621 = ~n41614 & n41620 ;
  assign n41622 = ~n41611 & n41621 ;
  assign n41639 = \P2_P1_PhyAddrPointer_reg[26]/NET0131  & n25947 ;
  assign n41640 = ~n37095 & ~n41639 ;
  assign n41641 = n25945 & ~n41640 ;
  assign n41642 = \P2_P1_PhyAddrPointer_reg[26]/NET0131  & ~n36677 ;
  assign n41643 = ~n37100 & ~n41642 ;
  assign n41644 = ~n41641 & n41643 ;
  assign n41645 = n11623 & ~n41644 ;
  assign n41623 = \P2_P1_PhyAddrPointer_reg[26]/NET0131  & ~n39455 ;
  assign n41624 = \P2_P1_PhyAddrPointer_reg[15]/NET0131  & \P2_P1_PhyAddrPointer_reg[20]/NET0131  ;
  assign n41627 = n36640 & n41624 ;
  assign n41628 = n39453 & n41627 ;
  assign n41625 = \P2_P1_PhyAddrPointer_reg[21]/NET0131  & \P2_P1_PhyAddrPointer_reg[22]/NET0131  ;
  assign n41626 = \P2_P1_PhyAddrPointer_reg[25]/NET0131  & n41625 ;
  assign n41629 = n36642 & n41626 ;
  assign n41630 = n36656 & n41629 ;
  assign n41631 = n41628 & n41630 ;
  assign n41632 = \P2_P1_PhyAddrPointer_reg[26]/NET0131  & n41631 ;
  assign n41633 = ~\P2_P1_PhyAddrPointer_reg[26]/NET0131  & ~n41631 ;
  assign n41634 = ~n41632 & ~n41633 ;
  assign n41635 = n36649 & n41634 ;
  assign n41636 = \P2_P1_PhyAddrPointer_reg[1]/NET0131  & n41635 ;
  assign n41637 = ~n41623 & ~n41636 ;
  assign n41649 = ~\P2_P1_DataWidth_reg[1]/NET0131  & n41637 ;
  assign n41646 = \P2_P1_PhyAddrPointer_reg[26]/NET0131  & ~n36649 ;
  assign n41647 = \P2_P1_DataWidth_reg[1]/NET0131  & ~n41635 ;
  assign n41648 = ~n41646 & n41647 ;
  assign n41650 = n11609 & ~n41648 ;
  assign n41651 = ~n41649 & n41650 ;
  assign n41638 = n11613 & ~n41637 ;
  assign n41652 = \P2_P1_PhyAddrPointer_reg[26]/NET0131  & ~n36687 ;
  assign n41653 = ~n37110 & ~n41652 ;
  assign n41654 = ~n41638 & n41653 ;
  assign n41655 = ~n41651 & n41654 ;
  assign n41656 = ~n41645 & n41655 ;
  assign n41657 = n26126 & n38455 ;
  assign n41658 = ~n26250 & n36696 ;
  assign n41659 = \P1_P1_PhyAddrPointer_reg[11]/NET0131  & ~n41658 ;
  assign n41660 = ~n38464 & ~n41659 ;
  assign n41661 = ~n41657 & n41660 ;
  assign n41662 = n8355 & ~n41661 ;
  assign n41666 = \P1_P1_PhyAddrPointer_reg[1]/NET0131  & n36707 ;
  assign n41667 = \P1_P1_PhyAddrPointer_reg[9]/NET0131  & n41666 ;
  assign n41668 = \P1_P1_PhyAddrPointer_reg[10]/NET0131  & n41667 ;
  assign n41669 = ~\P1_P1_PhyAddrPointer_reg[11]/NET0131  & ~n41668 ;
  assign n41670 = \P1_P1_PhyAddrPointer_reg[11]/NET0131  & n41668 ;
  assign n41671 = ~n41669 & ~n41670 ;
  assign n41672 = ~n36701 & n41671 ;
  assign n41663 = ~\P1_P1_PhyAddrPointer_reg[11]/NET0131  & ~n36709 ;
  assign n41664 = n27791 & ~n36710 ;
  assign n41665 = ~n41663 & n41664 ;
  assign n41673 = \P1_P1_PhyAddrPointer_reg[11]/NET0131  & ~n36743 ;
  assign n41674 = ~n38443 & ~n41673 ;
  assign n41675 = ~n41665 & n41674 ;
  assign n41676 = ~n41672 & n41675 ;
  assign n41677 = ~n41662 & n41676 ;
  assign n41681 = \P1_P1_PhyAddrPointer_reg[14]/NET0131  & n26249 ;
  assign n41682 = ~n38629 & ~n41681 ;
  assign n41683 = n26126 & ~n41682 ;
  assign n41684 = \P1_P1_PhyAddrPointer_reg[14]/NET0131  & ~n36696 ;
  assign n41685 = ~n38636 & ~n41684 ;
  assign n41686 = ~n41683 & n41685 ;
  assign n41687 = n8355 & ~n41686 ;
  assign n41678 = ~\P1_P1_PhyAddrPointer_reg[14]/NET0131  & ~n39558 ;
  assign n41679 = ~n39559 & ~n41678 ;
  assign n41688 = \P1_P1_DataWidth_reg[1]/NET0131  & ~n41667 ;
  assign n41690 = n36712 & n41688 ;
  assign n41691 = ~n41679 & ~n41690 ;
  assign n41689 = n36713 & n41688 ;
  assign n41692 = n8282 & ~n41689 ;
  assign n41693 = ~n41691 & n41692 ;
  assign n41680 = n8287 & n41679 ;
  assign n41694 = \P1_P1_PhyAddrPointer_reg[14]/NET0131  & ~n36743 ;
  assign n41695 = ~n38616 & ~n41694 ;
  assign n41696 = ~n41680 & n41695 ;
  assign n41697 = ~n41693 & n41696 ;
  assign n41698 = ~n41687 & n41697 ;
  assign n41699 = \P1_P1_PhyAddrPointer_reg[19]/NET0131  & n26249 ;
  assign n41700 = ~n37592 & ~n41699 ;
  assign n41701 = n26126 & ~n41700 ;
  assign n41702 = \P1_P1_PhyAddrPointer_reg[19]/NET0131  & ~n36696 ;
  assign n41703 = ~n37598 & ~n41702 ;
  assign n41704 = ~n41701 & n41703 ;
  assign n41705 = n8355 & ~n41704 ;
  assign n41711 = \P1_P1_PhyAddrPointer_reg[1]/NET0131  & n36715 ;
  assign n41712 = \P1_P1_PhyAddrPointer_reg[17]/NET0131  & n41711 ;
  assign n41713 = \P1_P1_PhyAddrPointer_reg[18]/NET0131  & n41712 ;
  assign n41714 = ~\P1_P1_PhyAddrPointer_reg[19]/NET0131  & ~n41713 ;
  assign n41715 = \P1_P1_PhyAddrPointer_reg[19]/NET0131  & n41713 ;
  assign n41716 = ~n41714 & ~n41715 ;
  assign n41717 = n8287 & n41716 ;
  assign n41706 = n36717 & ~n39569 ;
  assign n41708 = ~\P1_P1_PhyAddrPointer_reg[19]/NET0131  & ~n41706 ;
  assign n41707 = \P1_P1_PhyAddrPointer_reg[19]/NET0131  & n41706 ;
  assign n41709 = n8282 & ~n41707 ;
  assign n41710 = ~n41708 & n41709 ;
  assign n41718 = \P1_P1_PhyAddrPointer_reg[19]/NET0131  & ~n36743 ;
  assign n41719 = ~n37573 & ~n41718 ;
  assign n41720 = ~n41710 & n41719 ;
  assign n41721 = ~n41717 & n41720 ;
  assign n41722 = ~n41705 & n41721 ;
  assign n41724 = \P1_P1_PhyAddrPointer_reg[20]/NET0131  & n26249 ;
  assign n41725 = ~n37628 & ~n41724 ;
  assign n41726 = n26126 & ~n41725 ;
  assign n41727 = \P1_P1_PhyAddrPointer_reg[20]/NET0131  & ~n36696 ;
  assign n41728 = ~n37633 & ~n41727 ;
  assign n41729 = ~n41726 & n41728 ;
  assign n41730 = n8355 & ~n41729 ;
  assign n41736 = ~\P1_P1_PhyAddrPointer_reg[20]/NET0131  & ~n41707 ;
  assign n41735 = n36719 & ~n39569 ;
  assign n41737 = n8282 & ~n41735 ;
  assign n41738 = ~n41736 & n41737 ;
  assign n41731 = ~\P1_P1_PhyAddrPointer_reg[20]/NET0131  & ~n41715 ;
  assign n41732 = \P1_P1_PhyAddrPointer_reg[1]/NET0131  & n36719 ;
  assign n41733 = ~n41731 & ~n41732 ;
  assign n41734 = n8287 & n41733 ;
  assign n41723 = \P1_P1_PhyAddrPointer_reg[20]/NET0131  & ~n36743 ;
  assign n41739 = ~n37617 & ~n41723 ;
  assign n41740 = ~n41734 & n41739 ;
  assign n41741 = ~n41738 & n41740 ;
  assign n41742 = ~n41730 & n41741 ;
  assign n41747 = \P1_P1_PhyAddrPointer_reg[22]/NET0131  & n26249 ;
  assign n41748 = ~n37660 & ~n41747 ;
  assign n41749 = n26126 & ~n41748 ;
  assign n41750 = \P1_P1_PhyAddrPointer_reg[22]/NET0131  & ~n36696 ;
  assign n41751 = ~n37665 & ~n41750 ;
  assign n41752 = ~n41749 & n41751 ;
  assign n41753 = n8355 & ~n41752 ;
  assign n41754 = \P1_P1_PhyAddrPointer_reg[21]/NET0131  & n41735 ;
  assign n41755 = ~\P1_P1_PhyAddrPointer_reg[22]/NET0131  & ~n41754 ;
  assign n41756 = n39571 & ~n41755 ;
  assign n41743 = \P1_P1_PhyAddrPointer_reg[1]/NET0131  & n36720 ;
  assign n41744 = ~\P1_P1_PhyAddrPointer_reg[22]/NET0131  & ~n41743 ;
  assign n41745 = ~n39576 & ~n41744 ;
  assign n41746 = n8287 & n41745 ;
  assign n41757 = \P1_P1_PhyAddrPointer_reg[22]/NET0131  & ~n36743 ;
  assign n41758 = ~n37647 & ~n41757 ;
  assign n41759 = ~n41746 & n41758 ;
  assign n41760 = ~n41756 & n41759 ;
  assign n41761 = ~n41753 & n41760 ;
  assign n41763 = \P1_P1_PhyAddrPointer_reg[24]/NET0131  & n26249 ;
  assign n41764 = ~n37717 & ~n41763 ;
  assign n41765 = n26126 & ~n41764 ;
  assign n41766 = \P1_P1_PhyAddrPointer_reg[24]/NET0131  & ~n36696 ;
  assign n41767 = ~n37722 & ~n41766 ;
  assign n41768 = ~n41765 & n41767 ;
  assign n41769 = n8355 & ~n41768 ;
  assign n41774 = n36722 & ~n39569 ;
  assign n41776 = \P1_P1_PhyAddrPointer_reg[24]/NET0131  & n41774 ;
  assign n41775 = ~\P1_P1_PhyAddrPointer_reg[24]/NET0131  & ~n41774 ;
  assign n41777 = n8282 & ~n41775 ;
  assign n41778 = ~n41776 & n41777 ;
  assign n41770 = ~\P1_P1_PhyAddrPointer_reg[24]/NET0131  & ~n39578 ;
  assign n41771 = \P1_P1_PhyAddrPointer_reg[1]/NET0131  & n36723 ;
  assign n41772 = ~n41770 & ~n41771 ;
  assign n41773 = n8287 & n41772 ;
  assign n41762 = \P1_P1_PhyAddrPointer_reg[24]/NET0131  & ~n36743 ;
  assign n41779 = ~n37706 & ~n41762 ;
  assign n41780 = ~n41773 & n41779 ;
  assign n41781 = ~n41778 & n41780 ;
  assign n41782 = ~n41769 & n41781 ;
  assign n41792 = \P1_P1_PhyAddrPointer_reg[26]/NET0131  & n26249 ;
  assign n41793 = ~n37747 & ~n41792 ;
  assign n41794 = n26126 & ~n41793 ;
  assign n41795 = \P1_P1_PhyAddrPointer_reg[26]/NET0131  & ~n36696 ;
  assign n41796 = ~n37763 & ~n41795 ;
  assign n41797 = ~n41794 & n41796 ;
  assign n41798 = n8355 & ~n41797 ;
  assign n41788 = \P1_P1_PhyAddrPointer_reg[1]/NET0131  & n36724 ;
  assign n41789 = ~\P1_P1_PhyAddrPointer_reg[26]/NET0131  & ~n41788 ;
  assign n41790 = ~n39602 & ~n41789 ;
  assign n41791 = ~n36701 & n41790 ;
  assign n41783 = n27791 & ~n36724 ;
  assign n41784 = n36743 & ~n41783 ;
  assign n41785 = \P1_P1_PhyAddrPointer_reg[26]/NET0131  & ~n41784 ;
  assign n41786 = ~\P1_P1_PhyAddrPointer_reg[26]/NET0131  & n27791 ;
  assign n41787 = n36724 & n41786 ;
  assign n41799 = ~n37735 & ~n41787 ;
  assign n41800 = ~n41785 & n41799 ;
  assign n41801 = ~n41791 & n41800 ;
  assign n41802 = ~n41798 & n41801 ;
  assign n41803 = \P2_P2_PhyAddrPointer_reg[11]/NET0131  & n26629 ;
  assign n41804 = ~n38245 & ~n41803 ;
  assign n41805 = n26621 & ~n41804 ;
  assign n41806 = \P2_P2_PhyAddrPointer_reg[11]/NET0131  & ~n36752 ;
  assign n41807 = ~n38254 & ~n41806 ;
  assign n41808 = ~n41805 & n41807 ;
  assign n41809 = n26792 & ~n41808 ;
  assign n41813 = \P2_P2_PhyAddrPointer_reg[1]/NET0131  & n36765 ;
  assign n41814 = \P2_P2_PhyAddrPointer_reg[8]/NET0131  & n41813 ;
  assign n41815 = \P2_P2_PhyAddrPointer_reg[9]/NET0131  & n41814 ;
  assign n41816 = \P2_P2_PhyAddrPointer_reg[10]/NET0131  & n41815 ;
  assign n41817 = ~\P2_P2_PhyAddrPointer_reg[11]/NET0131  & ~n41816 ;
  assign n41818 = \P2_P2_PhyAddrPointer_reg[11]/NET0131  & n41816 ;
  assign n41819 = ~n41817 & ~n41818 ;
  assign n41820 = ~n36760 & n41819 ;
  assign n41810 = ~\P2_P2_PhyAddrPointer_reg[11]/NET0131  & ~n36768 ;
  assign n41811 = n26800 & ~n36769 ;
  assign n41812 = ~n41810 & n41811 ;
  assign n41821 = \P2_P2_PhyAddrPointer_reg[11]/NET0131  & ~n36758 ;
  assign n41822 = ~n38232 & ~n41821 ;
  assign n41823 = ~n41812 & n41822 ;
  assign n41824 = ~n41820 & n41823 ;
  assign n41825 = ~n41809 & n41824 ;
  assign n41829 = \P2_P2_PhyAddrPointer_reg[14]/NET0131  & n26629 ;
  assign n41830 = ~n38280 & ~n41829 ;
  assign n41831 = n26621 & ~n41830 ;
  assign n41832 = \P2_P2_PhyAddrPointer_reg[14]/NET0131  & ~n36752 ;
  assign n41833 = ~n38287 & ~n41832 ;
  assign n41834 = ~n41831 & n41833 ;
  assign n41835 = n26792 & ~n41834 ;
  assign n41826 = ~\P2_P2_PhyAddrPointer_reg[14]/NET0131  & ~n39648 ;
  assign n41827 = ~n39649 & ~n41826 ;
  assign n41836 = ~\P2_P2_DataWidth_reg[1]/NET0131  & ~n41827 ;
  assign n41837 = ~\P2_P2_PhyAddrPointer_reg[14]/NET0131  & ~n36771 ;
  assign n41838 = ~n36772 & ~n41837 ;
  assign n41839 = \P2_P2_DataWidth_reg[1]/NET0131  & ~n41838 ;
  assign n41840 = n26794 & ~n41839 ;
  assign n41841 = ~n41836 & n41840 ;
  assign n41828 = n27977 & n41827 ;
  assign n41842 = \P2_P2_PhyAddrPointer_reg[14]/NET0131  & ~n36758 ;
  assign n41843 = ~n38269 & ~n41842 ;
  assign n41844 = ~n41828 & n41843 ;
  assign n41845 = ~n41841 & n41844 ;
  assign n41846 = ~n41835 & n41845 ;
  assign n41847 = \P2_P2_PhyAddrPointer_reg[19]/NET0131  & n26629 ;
  assign n41848 = ~n37157 & ~n41847 ;
  assign n41849 = n26621 & ~n41848 ;
  assign n41850 = \P2_P2_PhyAddrPointer_reg[19]/NET0131  & ~n36752 ;
  assign n41851 = ~n37162 & ~n41850 ;
  assign n41852 = ~n41849 & n41851 ;
  assign n41853 = n26792 & ~n41852 ;
  assign n41857 = \P2_P2_PhyAddrPointer_reg[1]/NET0131  & n36775 ;
  assign n41858 = \P2_P2_PhyAddrPointer_reg[18]/NET0131  & n41857 ;
  assign n41859 = ~\P2_P2_PhyAddrPointer_reg[19]/NET0131  & ~n41858 ;
  assign n41860 = \P2_P2_PhyAddrPointer_reg[19]/NET0131  & n41858 ;
  assign n41861 = ~n41859 & ~n41860 ;
  assign n41862 = ~n36760 & n41861 ;
  assign n41854 = ~\P2_P2_PhyAddrPointer_reg[19]/NET0131  & ~n36776 ;
  assign n41855 = n26800 & ~n36777 ;
  assign n41856 = ~n41854 & n41855 ;
  assign n41863 = \P2_P2_PhyAddrPointer_reg[19]/NET0131  & ~n36758 ;
  assign n41864 = ~n37143 & ~n41863 ;
  assign n41865 = ~n41856 & n41864 ;
  assign n41866 = ~n41862 & n41865 ;
  assign n41867 = ~n41853 & n41866 ;
  assign n41872 = n26621 & n37192 ;
  assign n41873 = ~n26630 & n36752 ;
  assign n41874 = \P2_P2_PhyAddrPointer_reg[20]/NET0131  & ~n41873 ;
  assign n41875 = ~n37199 & ~n41874 ;
  assign n41876 = ~n41872 & n41875 ;
  assign n41877 = n26792 & ~n41876 ;
  assign n41880 = n36778 & ~n37979 ;
  assign n41878 = n36777 & ~n37979 ;
  assign n41879 = ~\P2_P2_PhyAddrPointer_reg[20]/NET0131  & ~n41878 ;
  assign n41881 = n26794 & ~n41879 ;
  assign n41882 = ~n41880 & n41881 ;
  assign n41868 = ~\P2_P2_PhyAddrPointer_reg[20]/NET0131  & ~n41860 ;
  assign n41869 = \P2_P2_PhyAddrPointer_reg[1]/NET0131  & n36778 ;
  assign n41870 = ~n41868 & ~n41869 ;
  assign n41871 = n27977 & n41870 ;
  assign n41883 = \P2_P2_PhyAddrPointer_reg[20]/NET0131  & ~n36758 ;
  assign n41884 = ~n37182 & ~n41883 ;
  assign n41885 = ~n41871 & n41884 ;
  assign n41886 = ~n41882 & n41885 ;
  assign n41887 = ~n41877 & n41886 ;
  assign n41888 = \P2_P2_PhyAddrPointer_reg[22]/NET0131  & n26629 ;
  assign n41889 = ~n37233 & ~n41888 ;
  assign n41890 = n26621 & ~n41889 ;
  assign n41891 = \P2_P2_PhyAddrPointer_reg[22]/NET0131  & ~n36752 ;
  assign n41892 = ~n37238 & ~n41891 ;
  assign n41893 = ~n41890 & n41892 ;
  assign n41894 = n26792 & ~n41893 ;
  assign n41898 = \P2_P2_PhyAddrPointer_reg[1]/NET0131  & n36779 ;
  assign n41899 = ~\P2_P2_PhyAddrPointer_reg[22]/NET0131  & ~n41898 ;
  assign n41900 = ~n39682 & ~n41899 ;
  assign n41901 = ~n36760 & n41900 ;
  assign n41895 = ~\P2_P2_PhyAddrPointer_reg[22]/NET0131  & ~n36779 ;
  assign n41896 = n26800 & ~n36780 ;
  assign n41897 = ~n41895 & n41896 ;
  assign n41902 = \P2_P2_PhyAddrPointer_reg[22]/NET0131  & ~n36758 ;
  assign n41903 = ~n37220 & ~n41902 ;
  assign n41904 = ~n41897 & n41903 ;
  assign n41905 = ~n41901 & n41904 ;
  assign n41906 = ~n41894 & n41905 ;
  assign n41907 = n26621 & n37266 ;
  assign n41908 = \P2_P2_PhyAddrPointer_reg[24]/NET0131  & ~n41873 ;
  assign n41909 = ~n37272 & ~n41908 ;
  assign n41910 = ~n41907 & n41909 ;
  assign n41911 = n26792 & ~n41910 ;
  assign n41915 = ~\P2_P2_PhyAddrPointer_reg[24]/NET0131  & ~n39684 ;
  assign n41916 = \P2_P2_PhyAddrPointer_reg[24]/NET0131  & n39684 ;
  assign n41917 = ~n41915 & ~n41916 ;
  assign n41918 = ~n36760 & n41917 ;
  assign n41912 = ~\P2_P2_PhyAddrPointer_reg[24]/NET0131  & ~n36781 ;
  assign n41913 = n26800 & ~n36782 ;
  assign n41914 = ~n41912 & n41913 ;
  assign n41919 = \P2_P2_PhyAddrPointer_reg[24]/NET0131  & ~n36758 ;
  assign n41920 = ~n37254 & ~n41919 ;
  assign n41921 = ~n41914 & n41920 ;
  assign n41922 = ~n41918 & n41921 ;
  assign n41923 = ~n41911 & n41922 ;
  assign n41924 = \P2_P2_PhyAddrPointer_reg[26]/NET0131  & n26629 ;
  assign n41925 = ~n37297 & ~n41924 ;
  assign n41926 = n26621 & ~n41925 ;
  assign n41927 = \P2_P2_PhyAddrPointer_reg[26]/NET0131  & ~n36752 ;
  assign n41928 = ~n37307 & ~n41927 ;
  assign n41929 = ~n41926 & n41928 ;
  assign n41930 = n26792 & ~n41929 ;
  assign n41934 = ~\P2_P2_PhyAddrPointer_reg[26]/NET0131  & ~n39702 ;
  assign n41935 = ~n39703 & ~n41934 ;
  assign n41936 = ~n36760 & n41935 ;
  assign n41931 = ~\P2_P2_PhyAddrPointer_reg[26]/NET0131  & ~n36783 ;
  assign n41932 = n26800 & ~n36784 ;
  assign n41933 = ~n41931 & n41932 ;
  assign n41937 = \P2_P2_PhyAddrPointer_reg[26]/NET0131  & ~n36758 ;
  assign n41938 = ~n37285 & ~n41937 ;
  assign n41939 = ~n41933 & n41938 ;
  assign n41940 = ~n41936 & n41939 ;
  assign n41941 = ~n41930 & n41940 ;
  assign n41942 = \P1_P3_PhyAddrPointer_reg[11]/NET0131  & n9072 ;
  assign n41943 = ~n19406 & ~n41942 ;
  assign n41944 = n9064 & ~n41943 ;
  assign n41945 = \P1_P3_PhyAddrPointer_reg[11]/NET0131  & ~n36805 ;
  assign n41946 = ~n19415 & ~n41945 ;
  assign n41947 = ~n41944 & n41946 ;
  assign n41948 = n9241 & ~n41947 ;
  assign n41952 = n17681 & ~n36810 ;
  assign n41949 = ~\P1_P3_PhyAddrPointer_reg[11]/NET0131  & ~n16460 ;
  assign n41950 = n11698 & ~n16461 ;
  assign n41951 = ~n41949 & n41950 ;
  assign n41953 = \P1_P3_PhyAddrPointer_reg[11]/NET0131  & ~n36816 ;
  assign n41954 = ~n19387 & ~n41953 ;
  assign n41955 = ~n41951 & n41954 ;
  assign n41956 = ~n41952 & n41955 ;
  assign n41957 = ~n41948 & n41956 ;
  assign n41959 = \P1_P3_PhyAddrPointer_reg[14]/NET0131  & n9072 ;
  assign n41960 = ~n19497 & ~n41959 ;
  assign n41961 = n9064 & ~n41960 ;
  assign n41962 = \P1_P3_PhyAddrPointer_reg[14]/NET0131  & ~n36805 ;
  assign n41963 = ~n19506 & ~n41962 ;
  assign n41964 = ~n41961 & n41963 ;
  assign n41965 = n9241 & ~n41964 ;
  assign n41966 = ~\P1_P3_DataWidth_reg[1]/NET0131  & ~n17793 ;
  assign n41967 = ~\P1_P3_PhyAddrPointer_reg[14]/NET0131  & ~n16463 ;
  assign n41968 = ~n16464 & ~n41967 ;
  assign n41969 = \P1_P3_DataWidth_reg[1]/NET0131  & ~n41968 ;
  assign n41970 = n9245 & ~n41969 ;
  assign n41971 = ~n41966 & n41970 ;
  assign n41958 = n16492 & n17793 ;
  assign n41972 = \P1_P3_PhyAddrPointer_reg[14]/NET0131  & ~n36816 ;
  assign n41973 = ~n19478 & ~n41972 ;
  assign n41974 = ~n41958 & n41973 ;
  assign n41975 = ~n41971 & n41974 ;
  assign n41976 = ~n41965 & n41975 ;
  assign n41977 = \P1_P3_PhyAddrPointer_reg[19]/NET0131  & n9072 ;
  assign n41978 = ~n19778 & ~n41977 ;
  assign n41979 = n9064 & ~n41978 ;
  assign n41980 = \P1_P3_PhyAddrPointer_reg[19]/NET0131  & ~n36805 ;
  assign n41981 = ~n19789 & ~n41980 ;
  assign n41982 = ~n41979 & n41981 ;
  assign n41983 = n9241 & ~n41982 ;
  assign n41987 = n16544 & ~n36810 ;
  assign n41984 = ~\P1_P3_PhyAddrPointer_reg[19]/NET0131  & ~n16468 ;
  assign n41985 = n11698 & ~n16469 ;
  assign n41986 = ~n41984 & n41985 ;
  assign n41988 = \P1_P3_PhyAddrPointer_reg[19]/NET0131  & ~n36816 ;
  assign n41989 = ~n19756 & ~n41988 ;
  assign n41990 = ~n41986 & n41989 ;
  assign n41991 = ~n41987 & n41990 ;
  assign n41992 = ~n41983 & n41991 ;
  assign n41993 = \P1_P3_PhyAddrPointer_reg[20]/NET0131  & n9072 ;
  assign n41994 = ~n19821 & ~n41993 ;
  assign n41995 = n9064 & ~n41994 ;
  assign n41996 = \P1_P3_PhyAddrPointer_reg[20]/NET0131  & ~n36805 ;
  assign n41997 = ~n19830 & ~n41996 ;
  assign n41998 = ~n41995 & n41997 ;
  assign n41999 = n9241 & ~n41998 ;
  assign n42006 = n16492 & n16542 ;
  assign n42000 = ~\P1_P3_DataWidth_reg[1]/NET0131  & ~\P1_P3_PhyAddrPointer_reg[1]/NET0131  ;
  assign n42001 = n16469 & ~n42000 ;
  assign n42003 = \P1_P3_PhyAddrPointer_reg[20]/NET0131  & n42001 ;
  assign n42002 = ~\P1_P3_PhyAddrPointer_reg[20]/NET0131  & ~n42001 ;
  assign n42004 = n9245 & ~n42002 ;
  assign n42005 = ~n42003 & n42004 ;
  assign n42007 = \P1_P3_PhyAddrPointer_reg[20]/NET0131  & ~n36816 ;
  assign n42008 = ~n19802 & ~n42007 ;
  assign n42009 = ~n42005 & n42008 ;
  assign n42010 = ~n42006 & n42009 ;
  assign n42011 = ~n41999 & n42010 ;
  assign n42013 = \P1_P3_PhyAddrPointer_reg[22]/NET0131  & n9072 ;
  assign n42014 = ~n19925 & ~n42013 ;
  assign n42015 = n9064 & ~n42014 ;
  assign n42016 = \P1_P3_PhyAddrPointer_reg[22]/NET0131  & ~n36805 ;
  assign n42017 = ~n19935 & ~n42016 ;
  assign n42018 = ~n42015 & n42017 ;
  assign n42019 = n9241 & ~n42018 ;
  assign n42020 = ~\P1_P3_DataWidth_reg[1]/NET0131  & ~n16670 ;
  assign n42021 = ~\P1_P3_PhyAddrPointer_reg[22]/NET0131  & ~n16471 ;
  assign n42022 = ~n16472 & ~n42021 ;
  assign n42023 = \P1_P3_DataWidth_reg[1]/NET0131  & ~n42022 ;
  assign n42024 = n9245 & ~n42023 ;
  assign n42025 = ~n42020 & n42024 ;
  assign n42012 = n16492 & n16670 ;
  assign n42026 = \P1_P3_PhyAddrPointer_reg[22]/NET0131  & ~n36816 ;
  assign n42027 = ~n19898 & ~n42026 ;
  assign n42028 = ~n42012 & n42027 ;
  assign n42029 = ~n42025 & n42028 ;
  assign n42030 = ~n42019 & n42029 ;
  assign n42031 = \P1_P3_PhyAddrPointer_reg[24]/NET0131  & n9072 ;
  assign n42032 = ~n20012 & ~n42031 ;
  assign n42033 = n9064 & ~n42032 ;
  assign n42034 = \P1_P3_PhyAddrPointer_reg[24]/NET0131  & ~n36805 ;
  assign n42035 = ~n20021 & ~n42034 ;
  assign n42036 = ~n42033 & n42035 ;
  assign n42037 = n9241 & ~n42036 ;
  assign n42041 = n16749 & ~n36810 ;
  assign n42038 = ~\P1_P3_PhyAddrPointer_reg[24]/NET0131  & ~n16473 ;
  assign n42039 = n11698 & ~n16474 ;
  assign n42040 = ~n42038 & n42039 ;
  assign n42042 = \P1_P3_PhyAddrPointer_reg[24]/NET0131  & ~n36816 ;
  assign n42043 = ~n19994 & ~n42042 ;
  assign n42044 = ~n42040 & n42043 ;
  assign n42045 = ~n42041 & n42044 ;
  assign n42046 = ~n42037 & n42045 ;
  assign n42048 = \P1_P3_PhyAddrPointer_reg[26]/NET0131  & n9072 ;
  assign n42049 = ~n20103 & ~n42048 ;
  assign n42050 = n9064 & ~n42049 ;
  assign n42051 = \P1_P3_PhyAddrPointer_reg[26]/NET0131  & ~n36805 ;
  assign n42052 = ~n20121 & ~n42051 ;
  assign n42053 = ~n42050 & n42052 ;
  assign n42054 = n9241 & ~n42053 ;
  assign n42055 = n16799 & ~n36810 ;
  assign n42056 = ~\P1_P3_PhyAddrPointer_reg[26]/NET0131  & ~n16475 ;
  assign n42057 = n39780 & ~n42056 ;
  assign n42047 = \P1_P3_PhyAddrPointer_reg[26]/NET0131  & ~n36816 ;
  assign n42058 = ~n20082 & ~n42047 ;
  assign n42059 = ~n42057 & n42058 ;
  assign n42060 = ~n42055 & n42059 ;
  assign n42061 = ~n42054 & n42060 ;
  assign n42062 = \P2_P3_PhyAddrPointer_reg[11]/NET0131  & ~n27283 ;
  assign n42063 = ~n38497 & ~n42062 ;
  assign n42064 = n27117 & ~n42063 ;
  assign n42065 = \P2_P3_PhyAddrPointer_reg[11]/NET0131  & ~n36826 ;
  assign n42066 = ~n38504 & ~n42065 ;
  assign n42067 = ~n42064 & n42066 ;
  assign n42068 = n27308 & ~n42067 ;
  assign n42072 = ~\P2_P3_PhyAddrPointer_reg[11]/NET0131  & ~n39840 ;
  assign n42073 = ~n39841 & ~n42072 ;
  assign n42074 = ~n36831 & n42073 ;
  assign n42069 = ~\P2_P3_PhyAddrPointer_reg[11]/NET0131  & ~n36842 ;
  assign n42070 = n27325 & ~n36843 ;
  assign n42071 = ~n42069 & n42070 ;
  assign n42075 = \P2_P3_PhyAddrPointer_reg[11]/NET0131  & ~n36873 ;
  assign n42076 = ~n38485 & ~n42075 ;
  assign n42077 = ~n42071 & n42076 ;
  assign n42078 = ~n42074 & n42077 ;
  assign n42079 = ~n42068 & n42078 ;
  assign n42088 = \P2_P3_PhyAddrPointer_reg[14]/NET0131  & ~n27283 ;
  assign n42089 = ~n38532 & ~n42088 ;
  assign n42090 = n27117 & ~n42089 ;
  assign n42091 = \P2_P3_PhyAddrPointer_reg[14]/NET0131  & ~n36826 ;
  assign n42092 = ~n38539 & ~n42091 ;
  assign n42093 = ~n42090 & n42092 ;
  assign n42094 = n27308 & ~n42093 ;
  assign n42085 = ~\P2_P3_PhyAddrPointer_reg[14]/NET0131  & ~n39842 ;
  assign n42086 = ~n39843 & ~n42085 ;
  assign n42087 = ~n36831 & n42086 ;
  assign n42080 = n27325 & ~n36845 ;
  assign n42081 = n36873 & ~n42080 ;
  assign n42082 = \P2_P3_PhyAddrPointer_reg[14]/NET0131  & ~n42081 ;
  assign n42083 = ~\P2_P3_PhyAddrPointer_reg[14]/NET0131  & n27325 ;
  assign n42084 = n36845 & n42083 ;
  assign n42095 = ~n38519 & ~n42084 ;
  assign n42096 = ~n42082 & n42095 ;
  assign n42097 = ~n42087 & n42096 ;
  assign n42098 = ~n42094 & n42097 ;
  assign n42099 = \P2_P3_PhyAddrPointer_reg[19]/NET0131  & ~n27283 ;
  assign n42100 = ~n37395 & ~n42099 ;
  assign n42101 = n27117 & ~n42100 ;
  assign n42102 = \P2_P3_PhyAddrPointer_reg[19]/NET0131  & ~n36826 ;
  assign n42103 = ~n37405 & ~n42102 ;
  assign n42104 = ~n42101 & n42103 ;
  assign n42105 = n27308 & ~n42104 ;
  assign n42113 = n36850 & n39843 ;
  assign n42106 = n36848 & n39845 ;
  assign n42107 = \P2_P3_PhyAddrPointer_reg[18]/NET0131  & n42106 ;
  assign n42114 = \P2_P3_PhyAddrPointer_reg[1]/NET0131  & n42107 ;
  assign n42115 = ~\P2_P3_PhyAddrPointer_reg[19]/NET0131  & ~n42114 ;
  assign n42116 = ~n42113 & ~n42115 ;
  assign n42117 = n32867 & n42116 ;
  assign n42108 = ~n39862 & n42107 ;
  assign n42110 = ~\P2_P3_PhyAddrPointer_reg[19]/NET0131  & ~n42108 ;
  assign n42109 = \P2_P3_PhyAddrPointer_reg[19]/NET0131  & n42108 ;
  assign n42111 = n27315 & ~n42109 ;
  assign n42112 = ~n42110 & n42111 ;
  assign n42118 = \P2_P3_PhyAddrPointer_reg[19]/NET0131  & ~n36873 ;
  assign n42119 = ~n37376 & ~n42118 ;
  assign n42120 = ~n42112 & n42119 ;
  assign n42121 = ~n42117 & n42120 ;
  assign n42122 = ~n42105 & n42121 ;
  assign n42126 = n27117 & n37431 ;
  assign n42127 = \P2_P3_PhyAddrPointer_reg[20]/NET0131  & ~n39857 ;
  assign n42128 = ~n37436 & ~n42127 ;
  assign n42129 = ~n42126 & n42128 ;
  assign n42130 = n27308 & ~n42129 ;
  assign n42132 = \P2_P3_PhyAddrPointer_reg[20]/NET0131  & n42109 ;
  assign n42131 = ~\P2_P3_PhyAddrPointer_reg[20]/NET0131  & ~n42109 ;
  assign n42133 = n27315 & ~n42131 ;
  assign n42134 = ~n42132 & n42133 ;
  assign n42123 = ~\P2_P3_PhyAddrPointer_reg[20]/NET0131  & ~n42113 ;
  assign n42124 = ~n39873 & ~n42123 ;
  assign n42125 = n32867 & n42124 ;
  assign n42135 = \P2_P3_PhyAddrPointer_reg[20]/NET0131  & ~n36873 ;
  assign n42136 = ~n37420 & ~n42135 ;
  assign n42137 = ~n42125 & n42136 ;
  assign n42138 = ~n42134 & n42137 ;
  assign n42139 = ~n42130 & n42138 ;
  assign n42148 = \P2_P3_PhyAddrPointer_reg[22]/NET0131  & ~n27283 ;
  assign n42149 = ~n37463 & ~n42148 ;
  assign n42150 = n27117 & ~n42149 ;
  assign n42151 = \P2_P3_PhyAddrPointer_reg[22]/NET0131  & ~n36826 ;
  assign n42152 = ~n37468 & ~n42151 ;
  assign n42153 = ~n42150 & n42152 ;
  assign n42154 = n27308 & ~n42153 ;
  assign n42145 = ~\P2_P3_PhyAddrPointer_reg[22]/NET0131  & ~n39870 ;
  assign n42146 = ~n39871 & ~n42145 ;
  assign n42147 = ~n36831 & n42146 ;
  assign n42140 = n27325 & ~n39863 ;
  assign n42141 = n36873 & ~n42140 ;
  assign n42142 = \P2_P3_PhyAddrPointer_reg[22]/NET0131  & ~n42141 ;
  assign n42143 = ~\P2_P3_PhyAddrPointer_reg[22]/NET0131  & n27325 ;
  assign n42144 = n39863 & n42143 ;
  assign n42155 = ~n37451 & ~n42144 ;
  assign n42156 = ~n42142 & n42155 ;
  assign n42157 = ~n42147 & n42156 ;
  assign n42158 = ~n42154 & n42157 ;
  assign n42163 = \P2_P3_PhyAddrPointer_reg[24]/NET0131  & ~n27283 ;
  assign n42164 = ~n37495 & ~n42163 ;
  assign n42165 = n27117 & ~n42164 ;
  assign n42166 = \P2_P3_PhyAddrPointer_reg[24]/NET0131  & ~n36826 ;
  assign n42167 = ~n37500 & ~n42166 ;
  assign n42168 = ~n42165 & n42167 ;
  assign n42169 = n27308 & ~n42168 ;
  assign n42171 = \P2_P3_PhyAddrPointer_reg[24]/NET0131  & n39866 ;
  assign n42170 = ~\P2_P3_PhyAddrPointer_reg[24]/NET0131  & ~n39866 ;
  assign n42172 = n27315 & ~n42170 ;
  assign n42173 = ~n42171 & n42172 ;
  assign n42159 = ~\P2_P3_PhyAddrPointer_reg[24]/NET0131  & ~n39874 ;
  assign n42160 = \P2_P3_PhyAddrPointer_reg[1]/NET0131  & n36853 ;
  assign n42161 = ~n42159 & ~n42160 ;
  assign n42162 = n32867 & n42161 ;
  assign n42174 = \P2_P3_PhyAddrPointer_reg[24]/NET0131  & ~n36873 ;
  assign n42175 = ~n37485 & ~n42174 ;
  assign n42176 = ~n42162 & n42175 ;
  assign n42177 = ~n42173 & n42176 ;
  assign n42178 = ~n42169 & n42177 ;
  assign n42179 = \P2_P3_PhyAddrPointer_reg[26]/NET0131  & ~n27283 ;
  assign n42180 = ~n37525 & ~n42179 ;
  assign n42181 = n27117 & ~n42180 ;
  assign n42182 = \P2_P3_PhyAddrPointer_reg[26]/NET0131  & ~n36826 ;
  assign n42183 = ~n37532 & ~n42182 ;
  assign n42184 = ~n42181 & n42183 ;
  assign n42185 = n27308 & ~n42184 ;
  assign n42186 = ~\P2_P3_PhyAddrPointer_reg[26]/NET0131  & ~n36854 ;
  assign n42187 = n27325 & ~n36855 ;
  assign n42188 = ~n42186 & n42187 ;
  assign n42189 = \P2_P3_PhyAddrPointer_reg[25]/NET0131  & n36834 ;
  assign n42190 = n39873 & n42189 ;
  assign n42191 = ~\P2_P3_PhyAddrPointer_reg[26]/NET0131  & ~n42190 ;
  assign n42192 = \P2_P3_PhyAddrPointer_reg[26]/NET0131  & n42190 ;
  assign n42193 = ~n42191 & ~n42192 ;
  assign n42194 = ~n36831 & n42193 ;
  assign n42195 = \P2_P3_PhyAddrPointer_reg[26]/NET0131  & ~n36873 ;
  assign n42196 = ~n37513 & ~n42195 ;
  assign n42197 = ~n42194 & n42196 ;
  assign n42198 = ~n42188 & n42197 ;
  assign n42199 = ~n42185 & n42198 ;
  assign n42202 = \P2_P1_InstAddrPointer_reg[7]/NET0131  & n25947 ;
  assign n42203 = n31800 & ~n31804 ;
  assign n42204 = n31894 & n31927 ;
  assign n42205 = ~n40057 & ~n42204 ;
  assign n42206 = ~n42203 & n42205 ;
  assign n42207 = ~n25947 & ~n42206 ;
  assign n42208 = ~n42202 & ~n42207 ;
  assign n42209 = n25945 & ~n42208 ;
  assign n42210 = ~n32062 & ~n32063 ;
  assign n42212 = ~n32098 & n42210 ;
  assign n42211 = n32098 & ~n42210 ;
  assign n42213 = n25964 & ~n42211 ;
  assign n42214 = ~n42212 & n42213 ;
  assign n42217 = ~n25995 & n31892 ;
  assign n42201 = n31546 & ~n32159 ;
  assign n42215 = \P2_P1_InstAddrPointer_reg[7]/NET0131  & ~n35385 ;
  assign n42216 = n26068 & n32061 ;
  assign n42218 = ~n42215 & ~n42216 ;
  assign n42219 = ~n42201 & n42218 ;
  assign n42220 = ~n42217 & n42219 ;
  assign n42221 = ~n42214 & n42220 ;
  assign n42222 = ~n42209 & n42221 ;
  assign n42223 = n11623 & ~n42222 ;
  assign n42200 = \P2_P1_rEIP_reg[7]/NET0131  & n11616 ;
  assign n42224 = \P2_P1_InstAddrPointer_reg[7]/NET0131  & ~n32172 ;
  assign n42225 = ~n42200 & ~n42224 ;
  assign n42226 = ~n42223 & n42225 ;
  assign n42231 = \P2_P1_InstAddrPointer_reg[9]/NET0131  & n25947 ;
  assign n42237 = ~n31930 & n31933 ;
  assign n42238 = ~n29503 & ~n31934 ;
  assign n42239 = ~n42237 & n42238 ;
  assign n42232 = ~\P2_P1_InstAddrPointer_reg[9]/NET0131  & ~n31802 ;
  assign n42233 = ~n31808 & ~n42232 ;
  assign n42234 = ~n31806 & ~n42233 ;
  assign n42235 = ~n31807 & ~n42234 ;
  assign n42236 = n29503 & ~n42235 ;
  assign n42240 = ~n25947 & ~n42236 ;
  assign n42241 = ~n42239 & n42240 ;
  assign n42242 = ~n42231 & ~n42241 ;
  assign n42243 = n25945 & ~n42242 ;
  assign n42228 = ~\P2_P1_InstAddrPointer_reg[9]/NET0131  & ~n32048 ;
  assign n42229 = ~n32049 & ~n42228 ;
  assign n42244 = ~n32101 & ~n42229 ;
  assign n42245 = n25964 & ~n32102 ;
  assign n42246 = ~n42244 & n42245 ;
  assign n42248 = ~n25995 & n31933 ;
  assign n42247 = ~n32159 & n42233 ;
  assign n42230 = n26068 & n42229 ;
  assign n42249 = \P2_P1_InstAddrPointer_reg[9]/NET0131  & ~n35385 ;
  assign n42250 = ~n42230 & ~n42249 ;
  assign n42251 = ~n42247 & n42250 ;
  assign n42252 = ~n42248 & n42251 ;
  assign n42253 = ~n42246 & n42252 ;
  assign n42254 = ~n42243 & n42253 ;
  assign n42255 = n11623 & ~n42254 ;
  assign n42227 = \P2_P1_rEIP_reg[9]/NET0131  & n11616 ;
  assign n42256 = \P2_P1_InstAddrPointer_reg[9]/NET0131  & ~n32172 ;
  assign n42257 = ~n42227 & ~n42256 ;
  assign n42258 = ~n42255 & n42257 ;
  assign n42263 = \P1_P2_InstAddrPointer_reg[9]/NET0131  & n25733 ;
  assign n42267 = n31209 & ~n31250 ;
  assign n42268 = ~n30809 & ~n31251 ;
  assign n42269 = ~n42267 & n42268 ;
  assign n42260 = ~\P1_P2_InstAddrPointer_reg[9]/NET0131  & ~n30853 ;
  assign n42261 = ~n31116 & ~n42260 ;
  assign n42264 = ~n31114 & ~n42261 ;
  assign n42265 = ~n31115 & ~n42264 ;
  assign n42266 = n30809 & ~n42265 ;
  assign n42270 = ~n25733 & ~n42266 ;
  assign n42271 = ~n42269 & n42270 ;
  assign n42272 = ~n42263 & ~n42271 ;
  assign n42273 = n25701 & ~n42272 ;
  assign n42274 = ~\P1_P2_InstAddrPointer_reg[9]/NET0131  & ~n31364 ;
  assign n42275 = ~n31414 & ~n42274 ;
  assign n42276 = ~n31412 & ~n42275 ;
  assign n42277 = n25881 & ~n31413 ;
  assign n42278 = ~n42276 & n42277 ;
  assign n42283 = ~n25817 & n31209 ;
  assign n42279 = ~n25743 & ~n31364 ;
  assign n42280 = n35131 & ~n42279 ;
  assign n42281 = \P1_P2_InstAddrPointer_reg[9]/NET0131  & ~n42280 ;
  assign n42262 = ~n25830 & n42261 ;
  assign n42282 = n25887 & n42275 ;
  assign n42284 = ~n42262 & ~n42282 ;
  assign n42285 = ~n42281 & n42284 ;
  assign n42286 = ~n42283 & n42285 ;
  assign n42287 = ~n42278 & n42286 ;
  assign n42288 = ~n42273 & n42287 ;
  assign n42289 = n25918 & ~n42288 ;
  assign n42259 = \P1_P2_rEIP_reg[9]/NET0131  & n27967 ;
  assign n42290 = \P1_P2_InstAddrPointer_reg[9]/NET0131  & ~n31487 ;
  assign n42291 = ~n42259 & ~n42290 ;
  assign n42292 = ~n42289 & n42291 ;
  assign n42296 = \P2_P2_InstAddrPointer_reg[7]/NET0131  & n26629 ;
  assign n42298 = ~n32479 & ~n32514 ;
  assign n42299 = n32510 & ~n42298 ;
  assign n42297 = ~n32629 & n32631 ;
  assign n42300 = ~n26629 & ~n42297 ;
  assign n42301 = ~n42299 & n42300 ;
  assign n42302 = ~n42296 & ~n42301 ;
  assign n42303 = n26621 & ~n42302 ;
  assign n42304 = ~n32768 & ~n32769 ;
  assign n42306 = ~n32801 & n42304 ;
  assign n42305 = n32801 & ~n42304 ;
  assign n42307 = n26744 & ~n42305 ;
  assign n42308 = ~n42306 & n42307 ;
  assign n42311 = ~n26688 & n32592 ;
  assign n42310 = \P2_P2_InstAddrPointer_reg[7]/NET0131  & ~n35424 ;
  assign n42295 = ~n26764 & n32226 ;
  assign n42309 = n26757 & n32767 ;
  assign n42312 = ~n42295 & ~n42309 ;
  assign n42313 = ~n42310 & n42312 ;
  assign n42314 = ~n42311 & n42313 ;
  assign n42315 = ~n42308 & n42314 ;
  assign n42316 = ~n42303 & n42315 ;
  assign n42317 = n26792 & ~n42316 ;
  assign n42293 = \P2_P2_rEIP_reg[7]/NET0131  & n28046 ;
  assign n42294 = \P2_P2_InstAddrPointer_reg[7]/NET0131  & ~n32860 ;
  assign n42318 = ~n42293 & ~n42294 ;
  assign n42319 = ~n42317 & n42318 ;
  assign n42323 = ~\P2_P2_InstAddrPointer_reg[9]/NET0131  & ~n32217 ;
  assign n42324 = ~n32221 & ~n42323 ;
  assign n42325 = ~n32516 & ~n42324 ;
  assign n42326 = ~n32517 & ~n42325 ;
  assign n42327 = n32510 & ~n42326 ;
  assign n42328 = ~n32636 & n32639 ;
  assign n42329 = ~n32510 & ~n32640 ;
  assign n42330 = ~n42328 & n42329 ;
  assign n42331 = ~n42327 & ~n42330 ;
  assign n42332 = ~n26629 & ~n42331 ;
  assign n42322 = ~\P2_P2_InstAddrPointer_reg[9]/NET0131  & n26629 ;
  assign n42333 = n26621 & ~n42322 ;
  assign n42334 = ~n42332 & n42333 ;
  assign n42335 = ~\P2_P2_InstAddrPointer_reg[9]/NET0131  & ~n32759 ;
  assign n42336 = ~n32760 & ~n42335 ;
  assign n42337 = ~n32804 & ~n42336 ;
  assign n42338 = n26744 & ~n32805 ;
  assign n42339 = ~n42337 & n42338 ;
  assign n42340 = ~n26688 & n32639 ;
  assign n42341 = ~n26764 & n42324 ;
  assign n42321 = \P2_P2_InstAddrPointer_reg[9]/NET0131  & ~n35424 ;
  assign n42342 = n26757 & n42336 ;
  assign n42343 = ~n42321 & ~n42342 ;
  assign n42344 = ~n42341 & n42343 ;
  assign n42345 = ~n42340 & n42344 ;
  assign n42346 = ~n42339 & n42345 ;
  assign n42347 = ~n42334 & n42346 ;
  assign n42348 = n26792 & ~n42347 ;
  assign n42320 = \P2_P2_rEIP_reg[9]/NET0131  & n28046 ;
  assign n42349 = \P2_P2_InstAddrPointer_reg[9]/NET0131  & ~n32860 ;
  assign n42350 = ~n42320 & ~n42349 ;
  assign n42351 = ~n42348 & n42350 ;
  assign n42354 = \P2_P3_InstAddrPointer_reg[7]/NET0131  & ~n27283 ;
  assign n42356 = ~n33210 & ~n33211 ;
  assign n42357 = n33242 & ~n42356 ;
  assign n42355 = n33327 & ~n33328 ;
  assign n42358 = n27283 & ~n42355 ;
  assign n42359 = ~n42357 & n42358 ;
  assign n42360 = ~n42354 & ~n42359 ;
  assign n42361 = n27117 & ~n42360 ;
  assign n42362 = ~n33434 & ~n33435 ;
  assign n42364 = ~n33470 & n42362 ;
  assign n42363 = n33470 & ~n42362 ;
  assign n42365 = n27280 & ~n42363 ;
  assign n42366 = ~n42364 & n42365 ;
  assign n42369 = ~n27229 & n32957 ;
  assign n42368 = ~n27142 & n33289 ;
  assign n42353 = \P2_P3_InstAddrPointer_reg[7]/NET0131  & ~n34355 ;
  assign n42367 = n27219 & n33433 ;
  assign n42370 = ~n42353 & ~n42367 ;
  assign n42371 = ~n42368 & n42370 ;
  assign n42372 = ~n42369 & n42371 ;
  assign n42373 = ~n42366 & n42372 ;
  assign n42374 = ~n42361 & n42373 ;
  assign n42375 = n27308 & ~n42374 ;
  assign n42352 = \P2_P3_rEIP_reg[7]/NET0131  & n32864 ;
  assign n42376 = \P2_P3_InstAddrPointer_reg[7]/NET0131  & ~n32870 ;
  assign n42377 = ~n42352 & ~n42376 ;
  assign n42378 = ~n42375 & n42377 ;
  assign n42382 = \P2_P3_InstAddrPointer_reg[9]/NET0131  & ~n27283 ;
  assign n42386 = ~\P2_P3_InstAddrPointer_reg[9]/NET0131  & ~n32914 ;
  assign n42387 = ~n32915 & ~n42386 ;
  assign n42388 = ~n33247 & ~n42387 ;
  assign n42389 = ~n33248 & ~n42388 ;
  assign n42390 = n33242 & ~n42389 ;
  assign n42383 = ~n33332 & n33334 ;
  assign n42384 = ~n33242 & ~n42383 ;
  assign n42385 = ~n40342 & n42384 ;
  assign n42391 = n27283 & ~n42385 ;
  assign n42392 = ~n42390 & n42391 ;
  assign n42393 = ~n42382 & ~n42392 ;
  assign n42394 = n27117 & ~n42393 ;
  assign n42395 = ~\P2_P3_InstAddrPointer_reg[9]/NET0131  & ~n32879 ;
  assign n42396 = ~n32880 & ~n42395 ;
  assign n42397 = ~n33473 & ~n42396 ;
  assign n42398 = n27280 & ~n33474 ;
  assign n42399 = ~n42397 & n42398 ;
  assign n42401 = ~n27229 & n42387 ;
  assign n42400 = ~n27142 & n33334 ;
  assign n42380 = n27235 & ~n27294 ;
  assign n42381 = \P2_P3_InstAddrPointer_reg[9]/NET0131  & ~n42380 ;
  assign n42402 = ~\P2_P3_InstAddrPointer_reg[9]/NET0131  & ~n27206 ;
  assign n42403 = n27206 & ~n42396 ;
  assign n42404 = ~n42402 & ~n42403 ;
  assign n42405 = ~n27111 & n42404 ;
  assign n42406 = ~n42381 & ~n42405 ;
  assign n42407 = ~n42400 & n42406 ;
  assign n42408 = ~n42401 & n42407 ;
  assign n42409 = ~n42399 & n42408 ;
  assign n42410 = ~n42394 & n42409 ;
  assign n42411 = n27308 & ~n42410 ;
  assign n42379 = \P2_P3_rEIP_reg[9]/NET0131  & n32864 ;
  assign n42412 = \P2_P3_InstAddrPointer_reg[9]/NET0131  & ~n32870 ;
  assign n42413 = ~n42379 & ~n42412 ;
  assign n42414 = ~n42411 & n42413 ;
  assign n42417 = \P1_P2_InstAddrPointer_reg[7]/NET0131  & n25733 ;
  assign n42420 = ~n31246 & n31248 ;
  assign n42418 = ~n31110 & ~n31111 ;
  assign n42419 = n30809 & ~n42418 ;
  assign n42421 = ~n25733 & ~n42419 ;
  assign n42422 = ~n42420 & n42421 ;
  assign n42423 = ~n42417 & ~n42422 ;
  assign n42424 = n25701 & ~n42423 ;
  assign n42425 = ~n31373 & ~n31374 ;
  assign n42427 = ~n31409 & n42425 ;
  assign n42426 = n31409 & ~n42425 ;
  assign n42428 = n25881 & ~n42426 ;
  assign n42429 = ~n42427 & n42428 ;
  assign n42416 = ~n25817 & n31213 ;
  assign n42430 = n25887 & n31372 ;
  assign n42433 = ~n42416 & ~n42430 ;
  assign n42431 = \P1_P2_InstAddrPointer_reg[7]/NET0131  & ~n34210 ;
  assign n42432 = n31109 & ~n34215 ;
  assign n42434 = ~n42431 & ~n42432 ;
  assign n42435 = n42433 & n42434 ;
  assign n42436 = ~n42429 & n42435 ;
  assign n42437 = ~n42424 & n42436 ;
  assign n42438 = n25918 & ~n42437 ;
  assign n42415 = \P1_P2_rEIP_reg[7]/NET0131  & n27967 ;
  assign n42439 = \P1_P2_InstAddrPointer_reg[7]/NET0131  & ~n31487 ;
  assign n42440 = ~n42415 & ~n42439 ;
  assign n42441 = ~n42438 & n42440 ;
  assign n42444 = \P1_P1_InstAddrPointer_reg[7]/NET0131  & n26249 ;
  assign n42445 = n33812 & ~n33813 ;
  assign n42446 = n33907 & n33939 ;
  assign n42447 = ~n40663 & ~n42446 ;
  assign n42448 = ~n42445 & n42447 ;
  assign n42449 = ~n26249 & ~n42448 ;
  assign n42450 = ~n42444 & ~n42449 ;
  assign n42451 = n26126 & ~n42450 ;
  assign n42452 = ~n34057 & ~n34058 ;
  assign n42454 = ~n34093 & n42452 ;
  assign n42453 = n34093 & ~n42452 ;
  assign n42455 = n26263 & ~n42453 ;
  assign n42456 = ~n42454 & n42455 ;
  assign n42443 = ~n26151 & n33905 ;
  assign n42462 = n26254 & ~n33558 ;
  assign n42461 = ~\P1_P1_InstAddrPointer_reg[7]/NET0131  & ~n26254 ;
  assign n42463 = ~n26160 & ~n42461 ;
  assign n42464 = ~n42462 & n42463 ;
  assign n42465 = ~\P1_P1_InstAddrPointer_reg[7]/NET0131  & ~n15365 ;
  assign n42466 = n15365 & ~n33558 ;
  assign n42467 = ~n42465 & ~n42466 ;
  assign n42468 = ~n15384 & n42467 ;
  assign n42457 = ~\P1_P1_InstAddrPointer_reg[7]/NET0131  & ~n15428 ;
  assign n42458 = n15428 & ~n34056 ;
  assign n42459 = ~n42457 & ~n42458 ;
  assign n42460 = ~n26123 & n42459 ;
  assign n42469 = \P1_P1_InstAddrPointer_reg[7]/NET0131  & n26251 ;
  assign n42470 = n26129 & n33558 ;
  assign n42471 = ~n42469 & ~n42470 ;
  assign n42472 = ~n42460 & n42471 ;
  assign n42473 = ~n42468 & n42472 ;
  assign n42474 = ~n42464 & n42473 ;
  assign n42475 = ~n42443 & n42474 ;
  assign n42476 = ~n42456 & n42475 ;
  assign n42477 = ~n42451 & n42476 ;
  assign n42478 = n8355 & ~n42477 ;
  assign n42442 = \P1_P1_rEIP_reg[7]/NET0131  & n8357 ;
  assign n42479 = \P1_P1_InstAddrPointer_reg[7]/NET0131  & ~n34164 ;
  assign n42480 = ~n42442 & ~n42479 ;
  assign n42481 = ~n42478 & n42480 ;
  assign n42484 = \P1_P1_InstAddrPointer_reg[9]/NET0131  & n26249 ;
  assign n42488 = ~n33554 & ~n33815 ;
  assign n42489 = ~n40284 & ~n42488 ;
  assign n42490 = n29558 & ~n42489 ;
  assign n42485 = n33901 & ~n33942 ;
  assign n42486 = ~n29558 & ~n33943 ;
  assign n42487 = ~n42485 & n42486 ;
  assign n42491 = ~n26249 & ~n42487 ;
  assign n42492 = ~n42490 & n42491 ;
  assign n42493 = ~n42484 & ~n42492 ;
  assign n42494 = n26126 & ~n42493 ;
  assign n42495 = ~\P1_P1_InstAddrPointer_reg[9]/NET0131  & ~n34027 ;
  assign n42496 = ~n34028 & ~n42495 ;
  assign n42497 = ~n34096 & ~n42496 ;
  assign n42498 = n26263 & ~n34097 ;
  assign n42499 = ~n42497 & n42498 ;
  assign n42504 = ~n26189 & n33554 ;
  assign n42500 = ~n26123 & ~n34027 ;
  assign n42501 = n35760 & ~n42500 ;
  assign n42502 = \P1_P1_InstAddrPointer_reg[9]/NET0131  & ~n42501 ;
  assign n42483 = ~n26151 & n33901 ;
  assign n42503 = n26192 & n42496 ;
  assign n42505 = ~n42483 & ~n42503 ;
  assign n42506 = ~n42502 & n42505 ;
  assign n42507 = ~n42504 & n42506 ;
  assign n42508 = ~n42499 & n42507 ;
  assign n42509 = ~n42494 & n42508 ;
  assign n42510 = n8355 & ~n42509 ;
  assign n42482 = \P1_P1_rEIP_reg[9]/NET0131  & n8357 ;
  assign n42511 = \P1_P1_InstAddrPointer_reg[9]/NET0131  & ~n34164 ;
  assign n42512 = ~n42482 & ~n42511 ;
  assign n42513 = ~n42510 & n42512 ;
  assign n42514 = \P2_P1_EAX_reg[4]/NET0131  & ~n27438 ;
  assign n42516 = ~n21069 & n24887 ;
  assign n42515 = n20728 & ~n31649 ;
  assign n42517 = ~\P2_P1_EAX_reg[4]/NET0131  & ~n21025 ;
  assign n42518 = ~n21026 & ~n42517 ;
  assign n42519 = n21022 & n42518 ;
  assign n42520 = ~n42515 & ~n42519 ;
  assign n42521 = ~n42516 & n42520 ;
  assign n42522 = n11623 & ~n42521 ;
  assign n42523 = ~n42514 & ~n42522 ;
  assign n42524 = \P1_P1_EAX_reg[4]/NET0131  & ~n15326 ;
  assign n42526 = \P1_P1_EAX_reg[4]/NET0131  & ~n15365 ;
  assign n42527 = ~n24696 & ~n42526 ;
  assign n42528 = ~n15384 & ~n42527 ;
  assign n42525 = \P1_P1_EAX_reg[4]/NET0131  & ~n23190 ;
  assign n42529 = n22818 & ~n33661 ;
  assign n42530 = ~\P1_P1_EAX_reg[4]/NET0131  & ~n15390 ;
  assign n42531 = ~n15391 & ~n42530 ;
  assign n42532 = n15377 & n42531 ;
  assign n42533 = ~n42529 & ~n42532 ;
  assign n42534 = ~n42525 & n42533 ;
  assign n42535 = ~n42528 & n42534 ;
  assign n42536 = n8355 & ~n42535 ;
  assign n42537 = ~n42524 & ~n42536 ;
  assign n42833 = \P2_P3_EAX_reg[0]/NET0131  & \P2_P3_EAX_reg[1]/NET0131  ;
  assign n42834 = \P2_P3_EAX_reg[2]/NET0131  & n42833 ;
  assign n42835 = \P2_P3_EAX_reg[3]/NET0131  & n42834 ;
  assign n42836 = \P2_P3_EAX_reg[4]/NET0131  & n42835 ;
  assign n42837 = \P2_P3_EAX_reg[5]/NET0131  & n42836 ;
  assign n42838 = \P2_P3_EAX_reg[6]/NET0131  & n42837 ;
  assign n42839 = \P2_P3_EAX_reg[7]/NET0131  & n42838 ;
  assign n42840 = \P2_P3_EAX_reg[8]/NET0131  & n42839 ;
  assign n42841 = \P2_P3_EAX_reg[9]/NET0131  & n42840 ;
  assign n42842 = \P2_P3_EAX_reg[10]/NET0131  & n42841 ;
  assign n42843 = \P2_P3_EAX_reg[11]/NET0131  & n42842 ;
  assign n42844 = \P2_P3_EAX_reg[12]/NET0131  & n42843 ;
  assign n42845 = \P2_P3_EAX_reg[13]/NET0131  & n42844 ;
  assign n42846 = \P2_P3_EAX_reg[14]/NET0131  & n42845 ;
  assign n42847 = \P2_P3_EAX_reg[15]/NET0131  & n42846 ;
  assign n42848 = \P2_P3_EAX_reg[16]/NET0131  & n42847 ;
  assign n42849 = \P2_P3_EAX_reg[17]/NET0131  & n42848 ;
  assign n42850 = \P2_P3_EAX_reg[18]/NET0131  & n42849 ;
  assign n42851 = \P2_P3_EAX_reg[21]/NET0131  & \P2_P3_EAX_reg[22]/NET0131  ;
  assign n42852 = \P2_P3_EAX_reg[23]/NET0131  & n42851 ;
  assign n42853 = \P2_P3_EAX_reg[20]/NET0131  & \P2_P3_EAX_reg[24]/NET0131  ;
  assign n42854 = \P2_P3_EAX_reg[19]/NET0131  & n42853 ;
  assign n42855 = n42852 & n42854 ;
  assign n42856 = n42850 & n42855 ;
  assign n42857 = \P2_P3_EAX_reg[25]/NET0131  & n42856 ;
  assign n42858 = \P2_P3_EAX_reg[26]/NET0131  & n42857 ;
  assign n42859 = \P2_P3_EAX_reg[27]/NET0131  & n42858 ;
  assign n42860 = \P2_P3_EAX_reg[28]/NET0131  & n42859 ;
  assign n42861 = \P2_P3_EAX_reg[29]/NET0131  & n42860 ;
  assign n42862 = \P2_P3_EAX_reg[30]/NET0131  & n42861 ;
  assign n42864 = \P2_P3_EAX_reg[31]/NET0131  & n42862 ;
  assign n42539 = n27055 & n27131 ;
  assign n42863 = ~\P2_P3_EAX_reg[31]/NET0131  & ~n42862 ;
  assign n42865 = n42539 & ~n42863 ;
  assign n42866 = ~n42864 & n42865 ;
  assign n42538 = n27110 & n27206 ;
  assign n42540 = n27226 & ~n42539 ;
  assign n42541 = ~n27110 & ~n42540 ;
  assign n42542 = ~n42538 & ~n42541 ;
  assign n42543 = ~n27234 & ~n42542 ;
  assign n42544 = \P2_P3_EAX_reg[31]/NET0131  & ~n42543 ;
  assign n42554 = \P2_P3_InstQueue_reg[10][7]/NET0131  & n26839 ;
  assign n42545 = \P2_P3_InstQueue_reg[8][7]/NET0131  & n26822 ;
  assign n42546 = \P2_P3_InstQueue_reg[7][7]/NET0131  & n26815 ;
  assign n42561 = ~n42545 & ~n42546 ;
  assign n42570 = ~n42554 & n42561 ;
  assign n42555 = \P2_P3_InstQueue_reg[2][7]/NET0131  & n26837 ;
  assign n42558 = \P2_P3_InstQueue_reg[1][7]/NET0131  & n26845 ;
  assign n42571 = ~n42555 & ~n42558 ;
  assign n42572 = n42570 & n42571 ;
  assign n42560 = \P2_P3_InstQueue_reg[3][7]/NET0131  & n26812 ;
  assign n42557 = \P2_P3_InstQueue_reg[11][7]/NET0131  & n26827 ;
  assign n42559 = \P2_P3_InstQueue_reg[0][7]/NET0131  & n26825 ;
  assign n42566 = ~n42557 & ~n42559 ;
  assign n42567 = ~n42560 & n42566 ;
  assign n42551 = \P2_P3_InstQueue_reg[5][7]/NET0131  & n26843 ;
  assign n42552 = \P2_P3_InstQueue_reg[12][7]/NET0131  & n26833 ;
  assign n42564 = ~n42551 & ~n42552 ;
  assign n42553 = \P2_P3_InstQueue_reg[6][7]/NET0131  & n26847 ;
  assign n42556 = \P2_P3_InstQueue_reg[9][7]/NET0131  & n26841 ;
  assign n42565 = ~n42553 & ~n42556 ;
  assign n42568 = n42564 & n42565 ;
  assign n42547 = \P2_P3_InstQueue_reg[14][7]/NET0131  & n26849 ;
  assign n42548 = \P2_P3_InstQueue_reg[13][7]/NET0131  & n26819 ;
  assign n42562 = ~n42547 & ~n42548 ;
  assign n42549 = \P2_P3_InstQueue_reg[4][7]/NET0131  & n26831 ;
  assign n42550 = \P2_P3_InstQueue_reg[15][7]/NET0131  & n26829 ;
  assign n42563 = ~n42549 & ~n42550 ;
  assign n42569 = n42562 & n42563 ;
  assign n42573 = n42568 & n42569 ;
  assign n42574 = n42567 & n42573 ;
  assign n42575 = n42572 & n42574 ;
  assign n42585 = \P2_P3_InstQueue_reg[3][0]/NET0131  & n26837 ;
  assign n42576 = \P2_P3_InstQueue_reg[5][0]/NET0131  & n26831 ;
  assign n42577 = \P2_P3_InstQueue_reg[7][0]/NET0131  & n26847 ;
  assign n42592 = ~n42576 & ~n42577 ;
  assign n42601 = ~n42585 & n42592 ;
  assign n42586 = \P2_P3_InstQueue_reg[11][0]/NET0131  & n26839 ;
  assign n42589 = \P2_P3_InstQueue_reg[2][0]/NET0131  & n26845 ;
  assign n42602 = ~n42586 & ~n42589 ;
  assign n42603 = n42601 & n42602 ;
  assign n42591 = \P2_P3_InstQueue_reg[1][0]/NET0131  & n26825 ;
  assign n42588 = \P2_P3_InstQueue_reg[12][0]/NET0131  & n26827 ;
  assign n42590 = \P2_P3_InstQueue_reg[15][0]/NET0131  & n26849 ;
  assign n42597 = ~n42588 & ~n42590 ;
  assign n42598 = ~n42591 & n42597 ;
  assign n42582 = \P2_P3_InstQueue_reg[6][0]/NET0131  & n26843 ;
  assign n42583 = \P2_P3_InstQueue_reg[14][0]/NET0131  & n26819 ;
  assign n42595 = ~n42582 & ~n42583 ;
  assign n42584 = \P2_P3_InstQueue_reg[0][0]/NET0131  & n26829 ;
  assign n42587 = \P2_P3_InstQueue_reg[10][0]/NET0131  & n26841 ;
  assign n42596 = ~n42584 & ~n42587 ;
  assign n42599 = n42595 & n42596 ;
  assign n42578 = \P2_P3_InstQueue_reg[8][0]/NET0131  & n26815 ;
  assign n42579 = \P2_P3_InstQueue_reg[9][0]/NET0131  & n26822 ;
  assign n42593 = ~n42578 & ~n42579 ;
  assign n42580 = \P2_P3_InstQueue_reg[13][0]/NET0131  & n26833 ;
  assign n42581 = \P2_P3_InstQueue_reg[4][0]/NET0131  & n26812 ;
  assign n42594 = ~n42580 & ~n42581 ;
  assign n42600 = n42593 & n42594 ;
  assign n42604 = n42599 & n42600 ;
  assign n42605 = n42598 & n42604 ;
  assign n42606 = n42603 & n42605 ;
  assign n42607 = ~n42575 & ~n42606 ;
  assign n42617 = \P2_P3_InstQueue_reg[3][1]/NET0131  & n26837 ;
  assign n42608 = \P2_P3_InstQueue_reg[5][1]/NET0131  & n26831 ;
  assign n42609 = \P2_P3_InstQueue_reg[7][1]/NET0131  & n26847 ;
  assign n42624 = ~n42608 & ~n42609 ;
  assign n42633 = ~n42617 & n42624 ;
  assign n42618 = \P2_P3_InstQueue_reg[11][1]/NET0131  & n26839 ;
  assign n42621 = \P2_P3_InstQueue_reg[2][1]/NET0131  & n26845 ;
  assign n42634 = ~n42618 & ~n42621 ;
  assign n42635 = n42633 & n42634 ;
  assign n42623 = \P2_P3_InstQueue_reg[1][1]/NET0131  & n26825 ;
  assign n42620 = \P2_P3_InstQueue_reg[12][1]/NET0131  & n26827 ;
  assign n42622 = \P2_P3_InstQueue_reg[15][1]/NET0131  & n26849 ;
  assign n42629 = ~n42620 & ~n42622 ;
  assign n42630 = ~n42623 & n42629 ;
  assign n42614 = \P2_P3_InstQueue_reg[6][1]/NET0131  & n26843 ;
  assign n42615 = \P2_P3_InstQueue_reg[14][1]/NET0131  & n26819 ;
  assign n42627 = ~n42614 & ~n42615 ;
  assign n42616 = \P2_P3_InstQueue_reg[0][1]/NET0131  & n26829 ;
  assign n42619 = \P2_P3_InstQueue_reg[10][1]/NET0131  & n26841 ;
  assign n42628 = ~n42616 & ~n42619 ;
  assign n42631 = n42627 & n42628 ;
  assign n42610 = \P2_P3_InstQueue_reg[8][1]/NET0131  & n26815 ;
  assign n42611 = \P2_P3_InstQueue_reg[9][1]/NET0131  & n26822 ;
  assign n42625 = ~n42610 & ~n42611 ;
  assign n42612 = \P2_P3_InstQueue_reg[13][1]/NET0131  & n26833 ;
  assign n42613 = \P2_P3_InstQueue_reg[4][1]/NET0131  & n26812 ;
  assign n42626 = ~n42612 & ~n42613 ;
  assign n42632 = n42625 & n42626 ;
  assign n42636 = n42631 & n42632 ;
  assign n42637 = n42630 & n42636 ;
  assign n42638 = n42635 & n42637 ;
  assign n42639 = n42607 & ~n42638 ;
  assign n42648 = \P2_P3_InstQueue_reg[2][2]/NET0131  & n26845 ;
  assign n42640 = \P2_P3_InstQueue_reg[13][2]/NET0131  & n26833 ;
  assign n42641 = \P2_P3_InstQueue_reg[1][2]/NET0131  & n26825 ;
  assign n42656 = ~n42640 & ~n42641 ;
  assign n42665 = ~n42648 & n42656 ;
  assign n42650 = \P2_P3_InstQueue_reg[3][2]/NET0131  & n26837 ;
  assign n42651 = \P2_P3_InstQueue_reg[11][2]/NET0131  & n26839 ;
  assign n42666 = ~n42650 & ~n42651 ;
  assign n42667 = n42665 & n42666 ;
  assign n42655 = \P2_P3_InstQueue_reg[8][2]/NET0131  & n26815 ;
  assign n42653 = \P2_P3_InstQueue_reg[14][2]/NET0131  & n26819 ;
  assign n42654 = \P2_P3_InstQueue_reg[5][2]/NET0131  & n26831 ;
  assign n42661 = ~n42653 & ~n42654 ;
  assign n42662 = ~n42655 & n42661 ;
  assign n42646 = \P2_P3_InstQueue_reg[15][2]/NET0131  & n26849 ;
  assign n42647 = \P2_P3_InstQueue_reg[7][2]/NET0131  & n26847 ;
  assign n42659 = ~n42646 & ~n42647 ;
  assign n42649 = \P2_P3_InstQueue_reg[10][2]/NET0131  & n26841 ;
  assign n42652 = \P2_P3_InstQueue_reg[4][2]/NET0131  & n26812 ;
  assign n42660 = ~n42649 & ~n42652 ;
  assign n42663 = n42659 & n42660 ;
  assign n42642 = \P2_P3_InstQueue_reg[6][2]/NET0131  & n26843 ;
  assign n42643 = \P2_P3_InstQueue_reg[0][2]/NET0131  & n26829 ;
  assign n42657 = ~n42642 & ~n42643 ;
  assign n42644 = \P2_P3_InstQueue_reg[9][2]/NET0131  & n26822 ;
  assign n42645 = \P2_P3_InstQueue_reg[12][2]/NET0131  & n26827 ;
  assign n42658 = ~n42644 & ~n42645 ;
  assign n42664 = n42657 & n42658 ;
  assign n42668 = n42663 & n42664 ;
  assign n42669 = n42662 & n42668 ;
  assign n42670 = n42667 & n42669 ;
  assign n42671 = n42639 & ~n42670 ;
  assign n42681 = \P2_P3_InstQueue_reg[3][3]/NET0131  & n26837 ;
  assign n42672 = \P2_P3_InstQueue_reg[1][3]/NET0131  & n26825 ;
  assign n42673 = \P2_P3_InstQueue_reg[7][3]/NET0131  & n26847 ;
  assign n42688 = ~n42672 & ~n42673 ;
  assign n42697 = ~n42681 & n42688 ;
  assign n42682 = \P2_P3_InstQueue_reg[11][3]/NET0131  & n26839 ;
  assign n42685 = \P2_P3_InstQueue_reg[2][3]/NET0131  & n26845 ;
  assign n42698 = ~n42682 & ~n42685 ;
  assign n42699 = n42697 & n42698 ;
  assign n42687 = \P2_P3_InstQueue_reg[5][3]/NET0131  & n26831 ;
  assign n42684 = \P2_P3_InstQueue_reg[12][3]/NET0131  & n26827 ;
  assign n42686 = \P2_P3_InstQueue_reg[15][3]/NET0131  & n26849 ;
  assign n42693 = ~n42684 & ~n42686 ;
  assign n42694 = ~n42687 & n42693 ;
  assign n42678 = \P2_P3_InstQueue_reg[6][3]/NET0131  & n26843 ;
  assign n42679 = \P2_P3_InstQueue_reg[14][3]/NET0131  & n26819 ;
  assign n42691 = ~n42678 & ~n42679 ;
  assign n42680 = \P2_P3_InstQueue_reg[0][3]/NET0131  & n26829 ;
  assign n42683 = \P2_P3_InstQueue_reg[10][3]/NET0131  & n26841 ;
  assign n42692 = ~n42680 & ~n42683 ;
  assign n42695 = n42691 & n42692 ;
  assign n42674 = \P2_P3_InstQueue_reg[8][3]/NET0131  & n26815 ;
  assign n42675 = \P2_P3_InstQueue_reg[9][3]/NET0131  & n26822 ;
  assign n42689 = ~n42674 & ~n42675 ;
  assign n42676 = \P2_P3_InstQueue_reg[13][3]/NET0131  & n26833 ;
  assign n42677 = \P2_P3_InstQueue_reg[4][3]/NET0131  & n26812 ;
  assign n42690 = ~n42676 & ~n42677 ;
  assign n42696 = n42689 & n42690 ;
  assign n42700 = n42695 & n42696 ;
  assign n42701 = n42694 & n42700 ;
  assign n42702 = n42699 & n42701 ;
  assign n42703 = n42671 & ~n42702 ;
  assign n42712 = \P2_P3_InstQueue_reg[2][4]/NET0131  & n26845 ;
  assign n42704 = \P2_P3_InstQueue_reg[13][4]/NET0131  & n26833 ;
  assign n42705 = \P2_P3_InstQueue_reg[1][4]/NET0131  & n26825 ;
  assign n42720 = ~n42704 & ~n42705 ;
  assign n42729 = ~n42712 & n42720 ;
  assign n42714 = \P2_P3_InstQueue_reg[3][4]/NET0131  & n26837 ;
  assign n42715 = \P2_P3_InstQueue_reg[11][4]/NET0131  & n26839 ;
  assign n42730 = ~n42714 & ~n42715 ;
  assign n42731 = n42729 & n42730 ;
  assign n42719 = \P2_P3_InstQueue_reg[8][4]/NET0131  & n26815 ;
  assign n42717 = \P2_P3_InstQueue_reg[14][4]/NET0131  & n26819 ;
  assign n42718 = \P2_P3_InstQueue_reg[5][4]/NET0131  & n26831 ;
  assign n42725 = ~n42717 & ~n42718 ;
  assign n42726 = ~n42719 & n42725 ;
  assign n42710 = \P2_P3_InstQueue_reg[15][4]/NET0131  & n26849 ;
  assign n42711 = \P2_P3_InstQueue_reg[7][4]/NET0131  & n26847 ;
  assign n42723 = ~n42710 & ~n42711 ;
  assign n42713 = \P2_P3_InstQueue_reg[10][4]/NET0131  & n26841 ;
  assign n42716 = \P2_P3_InstQueue_reg[4][4]/NET0131  & n26812 ;
  assign n42724 = ~n42713 & ~n42716 ;
  assign n42727 = n42723 & n42724 ;
  assign n42706 = \P2_P3_InstQueue_reg[6][4]/NET0131  & n26843 ;
  assign n42707 = \P2_P3_InstQueue_reg[0][4]/NET0131  & n26829 ;
  assign n42721 = ~n42706 & ~n42707 ;
  assign n42708 = \P2_P3_InstQueue_reg[9][4]/NET0131  & n26822 ;
  assign n42709 = \P2_P3_InstQueue_reg[12][4]/NET0131  & n26827 ;
  assign n42722 = ~n42708 & ~n42709 ;
  assign n42728 = n42721 & n42722 ;
  assign n42732 = n42727 & n42728 ;
  assign n42733 = n42726 & n42732 ;
  assign n42734 = n42731 & n42733 ;
  assign n42735 = n42703 & ~n42734 ;
  assign n42745 = \P2_P3_InstQueue_reg[3][5]/NET0131  & n26837 ;
  assign n42736 = \P2_P3_InstQueue_reg[8][5]/NET0131  & n26815 ;
  assign n42737 = \P2_P3_InstQueue_reg[7][5]/NET0131  & n26847 ;
  assign n42752 = ~n42736 & ~n42737 ;
  assign n42761 = ~n42745 & n42752 ;
  assign n42746 = \P2_P3_InstQueue_reg[11][5]/NET0131  & n26839 ;
  assign n42749 = \P2_P3_InstQueue_reg[2][5]/NET0131  & n26845 ;
  assign n42762 = ~n42746 & ~n42749 ;
  assign n42763 = n42761 & n42762 ;
  assign n42751 = \P2_P3_InstQueue_reg[9][5]/NET0131  & n26822 ;
  assign n42748 = \P2_P3_InstQueue_reg[6][5]/NET0131  & n26843 ;
  assign n42750 = \P2_P3_InstQueue_reg[15][5]/NET0131  & n26849 ;
  assign n42757 = ~n42748 & ~n42750 ;
  assign n42758 = ~n42751 & n42757 ;
  assign n42742 = \P2_P3_InstQueue_reg[5][5]/NET0131  & n26831 ;
  assign n42743 = \P2_P3_InstQueue_reg[4][5]/NET0131  & n26812 ;
  assign n42755 = ~n42742 & ~n42743 ;
  assign n42744 = \P2_P3_InstQueue_reg[14][5]/NET0131  & n26819 ;
  assign n42747 = \P2_P3_InstQueue_reg[10][5]/NET0131  & n26841 ;
  assign n42756 = ~n42744 & ~n42747 ;
  assign n42759 = n42755 & n42756 ;
  assign n42738 = \P2_P3_InstQueue_reg[0][5]/NET0131  & n26829 ;
  assign n42739 = \P2_P3_InstQueue_reg[1][5]/NET0131  & n26825 ;
  assign n42753 = ~n42738 & ~n42739 ;
  assign n42740 = \P2_P3_InstQueue_reg[13][5]/NET0131  & n26833 ;
  assign n42741 = \P2_P3_InstQueue_reg[12][5]/NET0131  & n26827 ;
  assign n42754 = ~n42740 & ~n42741 ;
  assign n42760 = n42753 & n42754 ;
  assign n42764 = n42759 & n42760 ;
  assign n42765 = n42758 & n42764 ;
  assign n42766 = n42763 & n42765 ;
  assign n42767 = n42735 & ~n42766 ;
  assign n42776 = \P2_P3_InstQueue_reg[2][6]/NET0131  & n26845 ;
  assign n42768 = \P2_P3_InstQueue_reg[5][6]/NET0131  & n26831 ;
  assign n42769 = \P2_P3_InstQueue_reg[9][6]/NET0131  & n26822 ;
  assign n42784 = ~n42768 & ~n42769 ;
  assign n42793 = ~n42776 & n42784 ;
  assign n42778 = \P2_P3_InstQueue_reg[3][6]/NET0131  & n26837 ;
  assign n42779 = \P2_P3_InstQueue_reg[11][6]/NET0131  & n26839 ;
  assign n42794 = ~n42778 & ~n42779 ;
  assign n42795 = n42793 & n42794 ;
  assign n42783 = \P2_P3_InstQueue_reg[1][6]/NET0131  & n26825 ;
  assign n42781 = \P2_P3_InstQueue_reg[15][6]/NET0131  & n26849 ;
  assign n42782 = \P2_P3_InstQueue_reg[7][6]/NET0131  & n26847 ;
  assign n42789 = ~n42781 & ~n42782 ;
  assign n42790 = ~n42783 & n42789 ;
  assign n42774 = \P2_P3_InstQueue_reg[13][6]/NET0131  & n26833 ;
  assign n42775 = \P2_P3_InstQueue_reg[4][6]/NET0131  & n26812 ;
  assign n42787 = ~n42774 & ~n42775 ;
  assign n42777 = \P2_P3_InstQueue_reg[10][6]/NET0131  & n26841 ;
  assign n42780 = \P2_P3_InstQueue_reg[14][6]/NET0131  & n26819 ;
  assign n42788 = ~n42777 & ~n42780 ;
  assign n42791 = n42787 & n42788 ;
  assign n42770 = \P2_P3_InstQueue_reg[6][6]/NET0131  & n26843 ;
  assign n42771 = \P2_P3_InstQueue_reg[8][6]/NET0131  & n26815 ;
  assign n42785 = ~n42770 & ~n42771 ;
  assign n42772 = \P2_P3_InstQueue_reg[0][6]/NET0131  & n26829 ;
  assign n42773 = \P2_P3_InstQueue_reg[12][6]/NET0131  & n26827 ;
  assign n42786 = ~n42772 & ~n42773 ;
  assign n42792 = n42785 & n42786 ;
  assign n42796 = n42791 & n42792 ;
  assign n42797 = n42790 & n42796 ;
  assign n42798 = n42795 & n42797 ;
  assign n42799 = n42767 & ~n42798 ;
  assign n42809 = \P2_P3_InstQueue_reg[3][7]/NET0131  & n26837 ;
  assign n42800 = \P2_P3_InstQueue_reg[15][7]/NET0131  & n26849 ;
  assign n42801 = \P2_P3_InstQueue_reg[7][7]/NET0131  & n26847 ;
  assign n42816 = ~n42800 & ~n42801 ;
  assign n42825 = ~n42809 & n42816 ;
  assign n42810 = \P2_P3_InstQueue_reg[11][7]/NET0131  & n26839 ;
  assign n42813 = \P2_P3_InstQueue_reg[2][7]/NET0131  & n26845 ;
  assign n42826 = ~n42810 & ~n42813 ;
  assign n42827 = n42825 & n42826 ;
  assign n42815 = \P2_P3_InstQueue_reg[9][7]/NET0131  & n26822 ;
  assign n42812 = \P2_P3_InstQueue_reg[6][7]/NET0131  & n26843 ;
  assign n42814 = \P2_P3_InstQueue_reg[8][7]/NET0131  & n26815 ;
  assign n42821 = ~n42812 & ~n42814 ;
  assign n42822 = ~n42815 & n42821 ;
  assign n42806 = \P2_P3_InstQueue_reg[5][7]/NET0131  & n26831 ;
  assign n42807 = \P2_P3_InstQueue_reg[0][7]/NET0131  & n26829 ;
  assign n42819 = ~n42806 & ~n42807 ;
  assign n42808 = \P2_P3_InstQueue_reg[14][7]/NET0131  & n26819 ;
  assign n42811 = \P2_P3_InstQueue_reg[10][7]/NET0131  & n26841 ;
  assign n42820 = ~n42808 & ~n42811 ;
  assign n42823 = n42819 & n42820 ;
  assign n42802 = \P2_P3_InstQueue_reg[4][7]/NET0131  & n26812 ;
  assign n42803 = \P2_P3_InstQueue_reg[1][7]/NET0131  & n26825 ;
  assign n42817 = ~n42802 & ~n42803 ;
  assign n42804 = \P2_P3_InstQueue_reg[12][7]/NET0131  & n26827 ;
  assign n42805 = \P2_P3_InstQueue_reg[13][7]/NET0131  & n26833 ;
  assign n42818 = ~n42804 & ~n42805 ;
  assign n42824 = n42817 & n42818 ;
  assign n42828 = n42823 & n42824 ;
  assign n42829 = n42822 & n42828 ;
  assign n42830 = n42827 & n42829 ;
  assign n42831 = n42799 & ~n42830 ;
  assign n42832 = n42538 & n42831 ;
  assign n42867 = ~n42544 & ~n42832 ;
  assign n42868 = ~n42866 & n42867 ;
  assign n42869 = n27308 & ~n42868 ;
  assign n42870 = ~n27650 & ~n27657 ;
  assign n42871 = ~n27310 & ~n27317 ;
  assign n42872 = n42870 & n42871 ;
  assign n42873 = \P2_P3_EAX_reg[31]/NET0131  & ~n42872 ;
  assign n42874 = ~n42869 & ~n42873 ;
  assign n43171 = \P1_P2_EAX_reg[0]/NET0131  & \P1_P2_EAX_reg[1]/NET0131  ;
  assign n43172 = \P1_P2_EAX_reg[2]/NET0131  & n43171 ;
  assign n43173 = \P1_P2_EAX_reg[3]/NET0131  & n43172 ;
  assign n43174 = \P1_P2_EAX_reg[4]/NET0131  & n43173 ;
  assign n43175 = \P1_P2_EAX_reg[5]/NET0131  & n43174 ;
  assign n43176 = \P1_P2_EAX_reg[6]/NET0131  & n43175 ;
  assign n43177 = \P1_P2_EAX_reg[7]/NET0131  & n43176 ;
  assign n43178 = \P1_P2_EAX_reg[8]/NET0131  & n43177 ;
  assign n43179 = \P1_P2_EAX_reg[9]/NET0131  & n43178 ;
  assign n43180 = \P1_P2_EAX_reg[10]/NET0131  & n43179 ;
  assign n43181 = \P1_P2_EAX_reg[11]/NET0131  & n43180 ;
  assign n43182 = \P1_P2_EAX_reg[12]/NET0131  & n43181 ;
  assign n43183 = \P1_P2_EAX_reg[13]/NET0131  & n43182 ;
  assign n43184 = \P1_P2_EAX_reg[14]/NET0131  & n43183 ;
  assign n43185 = \P1_P2_EAX_reg[15]/NET0131  & n43184 ;
  assign n43186 = \P1_P2_EAX_reg[16]/NET0131  & n43185 ;
  assign n43187 = \P1_P2_EAX_reg[17]/NET0131  & n43186 ;
  assign n43188 = \P1_P2_EAX_reg[18]/NET0131  & n43187 ;
  assign n43189 = \P1_P2_EAX_reg[19]/NET0131  & n43188 ;
  assign n43190 = \P1_P2_EAX_reg[20]/NET0131  & n43189 ;
  assign n43191 = \P1_P2_EAX_reg[21]/NET0131  & n43190 ;
  assign n43192 = \P1_P2_EAX_reg[22]/NET0131  & n43191 ;
  assign n43193 = \P1_P2_EAX_reg[23]/NET0131  & n43192 ;
  assign n43194 = \P1_P2_EAX_reg[24]/NET0131  & n43193 ;
  assign n43195 = \P1_P2_EAX_reg[25]/NET0131  & n43194 ;
  assign n43196 = \P1_P2_EAX_reg[26]/NET0131  & n43195 ;
  assign n43197 = \P1_P2_EAX_reg[27]/NET0131  & n43196 ;
  assign n43198 = \P1_P2_EAX_reg[28]/NET0131  & n43197 ;
  assign n43199 = \P1_P2_EAX_reg[29]/NET0131  & n43198 ;
  assign n43200 = \P1_P2_EAX_reg[30]/NET0131  & n43199 ;
  assign n43202 = \P1_P2_EAX_reg[31]/NET0131  & n43200 ;
  assign n43164 = n25793 & n25796 ;
  assign n43201 = ~\P1_P2_EAX_reg[31]/NET0131  & ~n43200 ;
  assign n43203 = n43164 & ~n43201 ;
  assign n43204 = ~n43202 & n43203 ;
  assign n42875 = n25742 & n25747 ;
  assign n42887 = \P1_P2_InstQueue_reg[9][7]/NET0131  & n25453 ;
  assign n42880 = \P1_P2_InstQueue_reg[10][7]/NET0131  & n25435 ;
  assign n42876 = \P1_P2_InstQueue_reg[4][7]/NET0131  & n25428 ;
  assign n42877 = \P1_P2_InstQueue_reg[0][7]/NET0131  & n25442 ;
  assign n42892 = ~n42876 & ~n42877 ;
  assign n42902 = ~n42880 & n42892 ;
  assign n42903 = ~n42887 & n42902 ;
  assign n42888 = \P1_P2_InstQueue_reg[13][7]/NET0131  & n25440 ;
  assign n42889 = \P1_P2_InstQueue_reg[3][7]/NET0131  & n25425 ;
  assign n42897 = ~n42888 & ~n42889 ;
  assign n42890 = \P1_P2_InstQueue_reg[6][7]/NET0131  & n25437 ;
  assign n42891 = \P1_P2_InstQueue_reg[8][7]/NET0131  & n25449 ;
  assign n42898 = ~n42890 & ~n42891 ;
  assign n42899 = n42897 & n42898 ;
  assign n42883 = \P1_P2_InstQueue_reg[11][7]/NET0131  & n25455 ;
  assign n42884 = \P1_P2_InstQueue_reg[7][7]/NET0131  & n25461 ;
  assign n42895 = ~n42883 & ~n42884 ;
  assign n42885 = \P1_P2_InstQueue_reg[2][7]/NET0131  & n25446 ;
  assign n42886 = \P1_P2_InstQueue_reg[15][7]/NET0131  & n25422 ;
  assign n42896 = ~n42885 & ~n42886 ;
  assign n42900 = n42895 & n42896 ;
  assign n42878 = \P1_P2_InstQueue_reg[14][7]/NET0131  & n25459 ;
  assign n42879 = \P1_P2_InstQueue_reg[1][7]/NET0131  & n25431 ;
  assign n42893 = ~n42878 & ~n42879 ;
  assign n42881 = \P1_P2_InstQueue_reg[12][7]/NET0131  & n25457 ;
  assign n42882 = \P1_P2_InstQueue_reg[5][7]/NET0131  & n25444 ;
  assign n42894 = ~n42881 & ~n42882 ;
  assign n42901 = n42893 & n42894 ;
  assign n42904 = n42900 & n42901 ;
  assign n42905 = n42899 & n42904 ;
  assign n42906 = n42903 & n42905 ;
  assign n42918 = \P1_P2_InstQueue_reg[10][0]/NET0131  & n25453 ;
  assign n42911 = \P1_P2_InstQueue_reg[11][0]/NET0131  & n25435 ;
  assign n42907 = \P1_P2_InstQueue_reg[5][0]/NET0131  & n25428 ;
  assign n42908 = \P1_P2_InstQueue_reg[4][0]/NET0131  & n25425 ;
  assign n42923 = ~n42907 & ~n42908 ;
  assign n42933 = ~n42911 & n42923 ;
  assign n42934 = ~n42918 & n42933 ;
  assign n42919 = \P1_P2_InstQueue_reg[12][0]/NET0131  & n25455 ;
  assign n42920 = \P1_P2_InstQueue_reg[0][0]/NET0131  & n25422 ;
  assign n42928 = ~n42919 & ~n42920 ;
  assign n42921 = \P1_P2_InstQueue_reg[7][0]/NET0131  & n25437 ;
  assign n42922 = \P1_P2_InstQueue_reg[14][0]/NET0131  & n25440 ;
  assign n42929 = ~n42921 & ~n42922 ;
  assign n42930 = n42928 & n42929 ;
  assign n42914 = \P1_P2_InstQueue_reg[8][0]/NET0131  & n25461 ;
  assign n42915 = \P1_P2_InstQueue_reg[1][0]/NET0131  & n25442 ;
  assign n42926 = ~n42914 & ~n42915 ;
  assign n42916 = \P1_P2_InstQueue_reg[3][0]/NET0131  & n25446 ;
  assign n42917 = \P1_P2_InstQueue_reg[13][0]/NET0131  & n25457 ;
  assign n42927 = ~n42916 & ~n42917 ;
  assign n42931 = n42926 & n42927 ;
  assign n42909 = \P1_P2_InstQueue_reg[6][0]/NET0131  & n25444 ;
  assign n42910 = \P1_P2_InstQueue_reg[2][0]/NET0131  & n25431 ;
  assign n42924 = ~n42909 & ~n42910 ;
  assign n42912 = \P1_P2_InstQueue_reg[15][0]/NET0131  & n25459 ;
  assign n42913 = \P1_P2_InstQueue_reg[9][0]/NET0131  & n25449 ;
  assign n42925 = ~n42912 & ~n42913 ;
  assign n42932 = n42924 & n42925 ;
  assign n42935 = n42931 & n42932 ;
  assign n42936 = n42930 & n42935 ;
  assign n42937 = n42934 & n42936 ;
  assign n42938 = ~n42906 & ~n42937 ;
  assign n42950 = \P1_P2_InstQueue_reg[10][1]/NET0131  & n25453 ;
  assign n42943 = \P1_P2_InstQueue_reg[11][1]/NET0131  & n25435 ;
  assign n42939 = \P1_P2_InstQueue_reg[1][1]/NET0131  & n25442 ;
  assign n42940 = \P1_P2_InstQueue_reg[4][1]/NET0131  & n25425 ;
  assign n42955 = ~n42939 & ~n42940 ;
  assign n42965 = ~n42943 & n42955 ;
  assign n42966 = ~n42950 & n42965 ;
  assign n42951 = \P1_P2_InstQueue_reg[14][1]/NET0131  & n25440 ;
  assign n42952 = \P1_P2_InstQueue_reg[0][1]/NET0131  & n25422 ;
  assign n42960 = ~n42951 & ~n42952 ;
  assign n42953 = \P1_P2_InstQueue_reg[6][1]/NET0131  & n25444 ;
  assign n42954 = \P1_P2_InstQueue_reg[5][1]/NET0131  & n25428 ;
  assign n42961 = ~n42953 & ~n42954 ;
  assign n42962 = n42960 & n42961 ;
  assign n42946 = \P1_P2_InstQueue_reg[8][1]/NET0131  & n25461 ;
  assign n42947 = \P1_P2_InstQueue_reg[7][1]/NET0131  & n25437 ;
  assign n42958 = ~n42946 & ~n42947 ;
  assign n42948 = \P1_P2_InstQueue_reg[3][1]/NET0131  & n25446 ;
  assign n42949 = \P1_P2_InstQueue_reg[13][1]/NET0131  & n25457 ;
  assign n42959 = ~n42948 & ~n42949 ;
  assign n42963 = n42958 & n42959 ;
  assign n42941 = \P1_P2_InstQueue_reg[12][1]/NET0131  & n25455 ;
  assign n42942 = \P1_P2_InstQueue_reg[2][1]/NET0131  & n25431 ;
  assign n42956 = ~n42941 & ~n42942 ;
  assign n42944 = \P1_P2_InstQueue_reg[9][1]/NET0131  & n25449 ;
  assign n42945 = \P1_P2_InstQueue_reg[15][1]/NET0131  & n25459 ;
  assign n42957 = ~n42944 & ~n42945 ;
  assign n42964 = n42956 & n42957 ;
  assign n42967 = n42963 & n42964 ;
  assign n42968 = n42962 & n42967 ;
  assign n42969 = n42966 & n42968 ;
  assign n42970 = n42938 & ~n42969 ;
  assign n42982 = \P1_P2_InstQueue_reg[10][2]/NET0131  & n25453 ;
  assign n42975 = \P1_P2_InstQueue_reg[11][2]/NET0131  & n25435 ;
  assign n42971 = \P1_P2_InstQueue_reg[1][2]/NET0131  & n25442 ;
  assign n42972 = \P1_P2_InstQueue_reg[4][2]/NET0131  & n25425 ;
  assign n42987 = ~n42971 & ~n42972 ;
  assign n42997 = ~n42975 & n42987 ;
  assign n42998 = ~n42982 & n42997 ;
  assign n42983 = \P1_P2_InstQueue_reg[14][2]/NET0131  & n25440 ;
  assign n42984 = \P1_P2_InstQueue_reg[0][2]/NET0131  & n25422 ;
  assign n42992 = ~n42983 & ~n42984 ;
  assign n42985 = \P1_P2_InstQueue_reg[6][2]/NET0131  & n25444 ;
  assign n42986 = \P1_P2_InstQueue_reg[5][2]/NET0131  & n25428 ;
  assign n42993 = ~n42985 & ~n42986 ;
  assign n42994 = n42992 & n42993 ;
  assign n42978 = \P1_P2_InstQueue_reg[8][2]/NET0131  & n25461 ;
  assign n42979 = \P1_P2_InstQueue_reg[7][2]/NET0131  & n25437 ;
  assign n42990 = ~n42978 & ~n42979 ;
  assign n42980 = \P1_P2_InstQueue_reg[3][2]/NET0131  & n25446 ;
  assign n42981 = \P1_P2_InstQueue_reg[13][2]/NET0131  & n25457 ;
  assign n42991 = ~n42980 & ~n42981 ;
  assign n42995 = n42990 & n42991 ;
  assign n42973 = \P1_P2_InstQueue_reg[12][2]/NET0131  & n25455 ;
  assign n42974 = \P1_P2_InstQueue_reg[2][2]/NET0131  & n25431 ;
  assign n42988 = ~n42973 & ~n42974 ;
  assign n42976 = \P1_P2_InstQueue_reg[9][2]/NET0131  & n25449 ;
  assign n42977 = \P1_P2_InstQueue_reg[15][2]/NET0131  & n25459 ;
  assign n42989 = ~n42976 & ~n42977 ;
  assign n42996 = n42988 & n42989 ;
  assign n42999 = n42995 & n42996 ;
  assign n43000 = n42994 & n42999 ;
  assign n43001 = n42998 & n43000 ;
  assign n43002 = n42970 & ~n43001 ;
  assign n43014 = \P1_P2_InstQueue_reg[10][3]/NET0131  & n25453 ;
  assign n43007 = \P1_P2_InstQueue_reg[11][3]/NET0131  & n25435 ;
  assign n43003 = \P1_P2_InstQueue_reg[1][3]/NET0131  & n25442 ;
  assign n43004 = \P1_P2_InstQueue_reg[4][3]/NET0131  & n25425 ;
  assign n43019 = ~n43003 & ~n43004 ;
  assign n43029 = ~n43007 & n43019 ;
  assign n43030 = ~n43014 & n43029 ;
  assign n43015 = \P1_P2_InstQueue_reg[14][3]/NET0131  & n25440 ;
  assign n43016 = \P1_P2_InstQueue_reg[0][3]/NET0131  & n25422 ;
  assign n43024 = ~n43015 & ~n43016 ;
  assign n43017 = \P1_P2_InstQueue_reg[6][3]/NET0131  & n25444 ;
  assign n43018 = \P1_P2_InstQueue_reg[5][3]/NET0131  & n25428 ;
  assign n43025 = ~n43017 & ~n43018 ;
  assign n43026 = n43024 & n43025 ;
  assign n43010 = \P1_P2_InstQueue_reg[8][3]/NET0131  & n25461 ;
  assign n43011 = \P1_P2_InstQueue_reg[7][3]/NET0131  & n25437 ;
  assign n43022 = ~n43010 & ~n43011 ;
  assign n43012 = \P1_P2_InstQueue_reg[3][3]/NET0131  & n25446 ;
  assign n43013 = \P1_P2_InstQueue_reg[13][3]/NET0131  & n25457 ;
  assign n43023 = ~n43012 & ~n43013 ;
  assign n43027 = n43022 & n43023 ;
  assign n43005 = \P1_P2_InstQueue_reg[12][3]/NET0131  & n25455 ;
  assign n43006 = \P1_P2_InstQueue_reg[2][3]/NET0131  & n25431 ;
  assign n43020 = ~n43005 & ~n43006 ;
  assign n43008 = \P1_P2_InstQueue_reg[9][3]/NET0131  & n25449 ;
  assign n43009 = \P1_P2_InstQueue_reg[15][3]/NET0131  & n25459 ;
  assign n43021 = ~n43008 & ~n43009 ;
  assign n43028 = n43020 & n43021 ;
  assign n43031 = n43027 & n43028 ;
  assign n43032 = n43026 & n43031 ;
  assign n43033 = n43030 & n43032 ;
  assign n43034 = n43002 & ~n43033 ;
  assign n43046 = \P1_P2_InstQueue_reg[10][4]/NET0131  & n25453 ;
  assign n43039 = \P1_P2_InstQueue_reg[11][4]/NET0131  & n25435 ;
  assign n43035 = \P1_P2_InstQueue_reg[1][4]/NET0131  & n25442 ;
  assign n43036 = \P1_P2_InstQueue_reg[4][4]/NET0131  & n25425 ;
  assign n43051 = ~n43035 & ~n43036 ;
  assign n43061 = ~n43039 & n43051 ;
  assign n43062 = ~n43046 & n43061 ;
  assign n43047 = \P1_P2_InstQueue_reg[14][4]/NET0131  & n25440 ;
  assign n43048 = \P1_P2_InstQueue_reg[0][4]/NET0131  & n25422 ;
  assign n43056 = ~n43047 & ~n43048 ;
  assign n43049 = \P1_P2_InstQueue_reg[6][4]/NET0131  & n25444 ;
  assign n43050 = \P1_P2_InstQueue_reg[5][4]/NET0131  & n25428 ;
  assign n43057 = ~n43049 & ~n43050 ;
  assign n43058 = n43056 & n43057 ;
  assign n43042 = \P1_P2_InstQueue_reg[8][4]/NET0131  & n25461 ;
  assign n43043 = \P1_P2_InstQueue_reg[7][4]/NET0131  & n25437 ;
  assign n43054 = ~n43042 & ~n43043 ;
  assign n43044 = \P1_P2_InstQueue_reg[3][4]/NET0131  & n25446 ;
  assign n43045 = \P1_P2_InstQueue_reg[13][4]/NET0131  & n25457 ;
  assign n43055 = ~n43044 & ~n43045 ;
  assign n43059 = n43054 & n43055 ;
  assign n43037 = \P1_P2_InstQueue_reg[12][4]/NET0131  & n25455 ;
  assign n43038 = \P1_P2_InstQueue_reg[2][4]/NET0131  & n25431 ;
  assign n43052 = ~n43037 & ~n43038 ;
  assign n43040 = \P1_P2_InstQueue_reg[9][4]/NET0131  & n25449 ;
  assign n43041 = \P1_P2_InstQueue_reg[15][4]/NET0131  & n25459 ;
  assign n43053 = ~n43040 & ~n43041 ;
  assign n43060 = n43052 & n43053 ;
  assign n43063 = n43059 & n43060 ;
  assign n43064 = n43058 & n43063 ;
  assign n43065 = n43062 & n43064 ;
  assign n43066 = n43034 & ~n43065 ;
  assign n43078 = \P1_P2_InstQueue_reg[10][5]/NET0131  & n25453 ;
  assign n43071 = \P1_P2_InstQueue_reg[11][5]/NET0131  & n25435 ;
  assign n43067 = \P1_P2_InstQueue_reg[5][5]/NET0131  & n25428 ;
  assign n43068 = \P1_P2_InstQueue_reg[12][5]/NET0131  & n25455 ;
  assign n43083 = ~n43067 & ~n43068 ;
  assign n43093 = ~n43071 & n43083 ;
  assign n43094 = ~n43078 & n43093 ;
  assign n43079 = \P1_P2_InstQueue_reg[0][5]/NET0131  & n25422 ;
  assign n43080 = \P1_P2_InstQueue_reg[8][5]/NET0131  & n25461 ;
  assign n43088 = ~n43079 & ~n43080 ;
  assign n43081 = \P1_P2_InstQueue_reg[13][5]/NET0131  & n25457 ;
  assign n43082 = \P1_P2_InstQueue_reg[9][5]/NET0131  & n25449 ;
  assign n43089 = ~n43081 & ~n43082 ;
  assign n43090 = n43088 & n43089 ;
  assign n43074 = \P1_P2_InstQueue_reg[14][5]/NET0131  & n25440 ;
  assign n43075 = \P1_P2_InstQueue_reg[6][5]/NET0131  & n25444 ;
  assign n43086 = ~n43074 & ~n43075 ;
  assign n43076 = \P1_P2_InstQueue_reg[3][5]/NET0131  & n25446 ;
  assign n43077 = \P1_P2_InstQueue_reg[7][5]/NET0131  & n25437 ;
  assign n43087 = ~n43076 & ~n43077 ;
  assign n43091 = n43086 & n43087 ;
  assign n43069 = \P1_P2_InstQueue_reg[4][5]/NET0131  & n25425 ;
  assign n43070 = \P1_P2_InstQueue_reg[2][5]/NET0131  & n25431 ;
  assign n43084 = ~n43069 & ~n43070 ;
  assign n43072 = \P1_P2_InstQueue_reg[15][5]/NET0131  & n25459 ;
  assign n43073 = \P1_P2_InstQueue_reg[1][5]/NET0131  & n25442 ;
  assign n43085 = ~n43072 & ~n43073 ;
  assign n43092 = n43084 & n43085 ;
  assign n43095 = n43091 & n43092 ;
  assign n43096 = n43090 & n43095 ;
  assign n43097 = n43094 & n43096 ;
  assign n43098 = n43066 & ~n43097 ;
  assign n43110 = \P1_P2_InstQueue_reg[10][6]/NET0131  & n25453 ;
  assign n43103 = \P1_P2_InstQueue_reg[11][6]/NET0131  & n25435 ;
  assign n43099 = \P1_P2_InstQueue_reg[9][6]/NET0131  & n25449 ;
  assign n43100 = \P1_P2_InstQueue_reg[14][6]/NET0131  & n25440 ;
  assign n43115 = ~n43099 & ~n43100 ;
  assign n43125 = ~n43103 & n43115 ;
  assign n43126 = ~n43110 & n43125 ;
  assign n43111 = \P1_P2_InstQueue_reg[0][6]/NET0131  & n25422 ;
  assign n43112 = \P1_P2_InstQueue_reg[8][6]/NET0131  & n25461 ;
  assign n43120 = ~n43111 & ~n43112 ;
  assign n43113 = \P1_P2_InstQueue_reg[15][6]/NET0131  & n25459 ;
  assign n43114 = \P1_P2_InstQueue_reg[4][6]/NET0131  & n25425 ;
  assign n43121 = ~n43113 & ~n43114 ;
  assign n43122 = n43120 & n43121 ;
  assign n43106 = \P1_P2_InstQueue_reg[5][6]/NET0131  & n25428 ;
  assign n43107 = \P1_P2_InstQueue_reg[12][6]/NET0131  & n25455 ;
  assign n43118 = ~n43106 & ~n43107 ;
  assign n43108 = \P1_P2_InstQueue_reg[3][6]/NET0131  & n25446 ;
  assign n43109 = \P1_P2_InstQueue_reg[13][6]/NET0131  & n25457 ;
  assign n43119 = ~n43108 & ~n43109 ;
  assign n43123 = n43118 & n43119 ;
  assign n43101 = \P1_P2_InstQueue_reg[7][6]/NET0131  & n25437 ;
  assign n43102 = \P1_P2_InstQueue_reg[2][6]/NET0131  & n25431 ;
  assign n43116 = ~n43101 & ~n43102 ;
  assign n43104 = \P1_P2_InstQueue_reg[1][6]/NET0131  & n25442 ;
  assign n43105 = \P1_P2_InstQueue_reg[6][6]/NET0131  & n25444 ;
  assign n43117 = ~n43104 & ~n43105 ;
  assign n43124 = n43116 & n43117 ;
  assign n43127 = n43123 & n43124 ;
  assign n43128 = n43122 & n43127 ;
  assign n43129 = n43126 & n43128 ;
  assign n43130 = n43098 & ~n43129 ;
  assign n43142 = \P1_P2_InstQueue_reg[10][7]/NET0131  & n25453 ;
  assign n43135 = \P1_P2_InstQueue_reg[11][7]/NET0131  & n25435 ;
  assign n43131 = \P1_P2_InstQueue_reg[9][7]/NET0131  & n25449 ;
  assign n43132 = \P1_P2_InstQueue_reg[14][7]/NET0131  & n25440 ;
  assign n43147 = ~n43131 & ~n43132 ;
  assign n43157 = ~n43135 & n43147 ;
  assign n43158 = ~n43142 & n43157 ;
  assign n43143 = \P1_P2_InstQueue_reg[4][7]/NET0131  & n25425 ;
  assign n43144 = \P1_P2_InstQueue_reg[1][7]/NET0131  & n25442 ;
  assign n43152 = ~n43143 & ~n43144 ;
  assign n43145 = \P1_P2_InstQueue_reg[15][7]/NET0131  & n25459 ;
  assign n43146 = \P1_P2_InstQueue_reg[6][7]/NET0131  & n25444 ;
  assign n43153 = ~n43145 & ~n43146 ;
  assign n43154 = n43152 & n43153 ;
  assign n43138 = \P1_P2_InstQueue_reg[12][7]/NET0131  & n25455 ;
  assign n43139 = \P1_P2_InstQueue_reg[13][7]/NET0131  & n25457 ;
  assign n43150 = ~n43138 & ~n43139 ;
  assign n43140 = \P1_P2_InstQueue_reg[3][7]/NET0131  & n25446 ;
  assign n43141 = \P1_P2_InstQueue_reg[0][7]/NET0131  & n25422 ;
  assign n43151 = ~n43140 & ~n43141 ;
  assign n43155 = n43150 & n43151 ;
  assign n43133 = \P1_P2_InstQueue_reg[5][7]/NET0131  & n25428 ;
  assign n43134 = \P1_P2_InstQueue_reg[2][7]/NET0131  & n25431 ;
  assign n43148 = ~n43133 & ~n43134 ;
  assign n43136 = \P1_P2_InstQueue_reg[7][7]/NET0131  & n25437 ;
  assign n43137 = \P1_P2_InstQueue_reg[8][7]/NET0131  & n25461 ;
  assign n43149 = ~n43136 & ~n43137 ;
  assign n43156 = n43148 & n43149 ;
  assign n43159 = n43155 & n43156 ;
  assign n43160 = n43154 & n43159 ;
  assign n43161 = n43158 & n43160 ;
  assign n43162 = n43130 & ~n43161 ;
  assign n43163 = n42875 & n43162 ;
  assign n43165 = n25826 & ~n43164 ;
  assign n43166 = ~n25742 & ~n43165 ;
  assign n43167 = ~n42875 & ~n43166 ;
  assign n43168 = ~n25777 & ~n43167 ;
  assign n43169 = ~n25775 & n43168 ;
  assign n43170 = \P1_P2_EAX_reg[31]/NET0131  & ~n43169 ;
  assign n43205 = ~n43163 & ~n43170 ;
  assign n43206 = ~n43204 & n43205 ;
  assign n43207 = n25918 & ~n43206 ;
  assign n43208 = ~n25416 & n27606 ;
  assign n43209 = ~n25417 & ~n27609 ;
  assign n43210 = ~n25928 & n43209 ;
  assign n43211 = ~n25935 & n43210 ;
  assign n43212 = ~n43208 & n43211 ;
  assign n43213 = \P1_P2_EAX_reg[31]/NET0131  & ~n43212 ;
  assign n43214 = ~n43207 & ~n43213 ;
  assign n43216 = n25903 & n25918 ;
  assign n43217 = ~n25924 & ~n25935 ;
  assign n43218 = n27969 & n43217 ;
  assign n43219 = \P1_P2_InstQueueRd_Addr_reg[0]/NET0131  & ~n43218 ;
  assign n43215 = ~\P1_P2_InstQueueRd_Addr_reg[0]/NET0131  & n27608 ;
  assign n43220 = \P1_P2_Flush_reg/NET0131  & \P1_P2_InstAddrPointer_reg[0]/NET0131  ;
  assign n43221 = ~\P1_P2_Flush_reg/NET0131  & ~\P1_P2_InstQueueRd_Addr_reg[0]/NET0131  ;
  assign n43222 = ~n43220 & ~n43221 ;
  assign n43223 = n27609 & n43222 ;
  assign n43224 = ~n43215 & ~n43223 ;
  assign n43225 = ~n43219 & n43224 ;
  assign n43226 = ~n43216 & n43225 ;
  assign n43228 = n11623 & n26092 ;
  assign n43229 = ~n11608 & ~n25940 ;
  assign n43230 = ~n11625 & n43229 ;
  assign n43231 = n11619 & n43230 ;
  assign n43232 = \P2_P1_InstQueueRd_Addr_reg[0]/NET0131  & ~n43231 ;
  assign n43227 = ~\P2_P1_InstQueueRd_Addr_reg[0]/NET0131  & n11692 ;
  assign n43233 = \P2_P1_Flush_reg/NET0131  & \P2_P1_InstAddrPointer_reg[0]/NET0131  ;
  assign n43234 = ~\P2_P1_Flush_reg/NET0131  & ~\P2_P1_InstQueueRd_Addr_reg[0]/NET0131  ;
  assign n43235 = ~n43233 & ~n43234 ;
  assign n43236 = n21096 & n43235 ;
  assign n43237 = ~n43227 & ~n43236 ;
  assign n43238 = ~n43232 & n43237 ;
  assign n43239 = ~n43228 & n43238 ;
  assign n43241 = n26775 & n26792 ;
  assign n43242 = ~n26285 & ~n27635 ;
  assign n43243 = ~n26290 & ~n43242 ;
  assign n43244 = n28047 & ~n43243 ;
  assign n43245 = \P2_P2_InstQueueRd_Addr_reg[0]/NET0131  & ~n43244 ;
  assign n43240 = ~\P2_P2_InstQueueRd_Addr_reg[0]/NET0131  & n27613 ;
  assign n43246 = \P2_P2_Flush_reg/NET0131  & \P2_P2_InstAddrPointer_reg[0]/NET0131  ;
  assign n43247 = ~\P2_P2_Flush_reg/NET0131  & ~\P2_P2_InstQueueRd_Addr_reg[0]/NET0131  ;
  assign n43248 = ~n43246 & ~n43247 ;
  assign n43249 = n27615 & n43248 ;
  assign n43250 = ~n43240 & ~n43249 ;
  assign n43251 = ~n43245 & n43250 ;
  assign n43252 = ~n43241 & n43251 ;
  assign n43254 = n9225 & n9241 ;
  assign n43256 = ~\P1_P3_State2_reg[0]/NET0131  & n10036 ;
  assign n43257 = ~n10031 & ~n43256 ;
  assign n43255 = ~n9247 & ~n17426 ;
  assign n43258 = n18340 & n43255 ;
  assign n43259 = n43257 & n43258 ;
  assign n43260 = \P1_P3_InstQueueRd_Addr_reg[0]/NET0131  & ~n43259 ;
  assign n43253 = ~\P1_P3_InstQueueRd_Addr_reg[0]/NET0131  & n10046 ;
  assign n43261 = ~\P1_P3_Flush_reg/NET0131  & ~\P1_P3_InstQueueRd_Addr_reg[0]/NET0131  ;
  assign n43262 = ~n15306 & ~n43261 ;
  assign n43263 = n10037 & n43262 ;
  assign n43264 = ~n43253 & ~n43263 ;
  assign n43265 = ~n43260 & n43264 ;
  assign n43266 = ~n43254 & n43265 ;
  assign n43268 = n27245 & n27308 ;
  assign n43269 = ~n27311 & ~n32864 ;
  assign n43270 = ~n27651 & n43269 ;
  assign n43271 = ~n27314 & ~n27318 ;
  assign n43272 = n43270 & n43271 ;
  assign n43273 = \P2_P3_InstQueueRd_Addr_reg[0]/NET0131  & ~n43272 ;
  assign n43267 = ~\P2_P3_InstQueueRd_Addr_reg[0]/NET0131  & n27788 ;
  assign n43274 = \P2_P3_Flush_reg/NET0131  & \P2_P3_InstAddrPointer_reg[0]/NET0131  ;
  assign n43275 = ~\P2_P3_Flush_reg/NET0131  & ~\P2_P3_InstQueueRd_Addr_reg[0]/NET0131  ;
  assign n43276 = ~n43274 & ~n43275 ;
  assign n43277 = n27657 & n43276 ;
  assign n43278 = ~n43267 & ~n43277 ;
  assign n43279 = ~n43273 & n43278 ;
  assign n43280 = ~n43268 & n43279 ;
  assign n43282 = n8355 & n26212 ;
  assign n43283 = ~n8281 & ~n26113 ;
  assign n43284 = n8362 & n43283 ;
  assign n43285 = \P1_P1_InstQueueRd_Addr_reg[0]/NET0131  & ~n43284 ;
  assign n43281 = ~\P1_P1_InstQueueRd_Addr_reg[0]/NET0131  & n8350 ;
  assign n43286 = \P1_P1_Flush_reg/NET0131  & \P1_P1_InstAddrPointer_reg[0]/NET0131  ;
  assign n43287 = ~\P1_P1_Flush_reg/NET0131  & ~\P1_P1_InstQueueRd_Addr_reg[0]/NET0131  ;
  assign n43288 = ~n43286 & ~n43287 ;
  assign n43289 = n15322 & n43288 ;
  assign n43290 = ~n43281 & ~n43289 ;
  assign n43291 = ~n43285 & n43290 ;
  assign n43292 = ~n43282 & n43291 ;
  assign n43297 = n25701 & n40608 ;
  assign n43298 = \P1_P2_PhyAddrPointer_reg[12]/NET0131  & ~n39340 ;
  assign n43299 = ~n40615 & ~n43298 ;
  assign n43300 = ~n43297 & n43299 ;
  assign n43301 = n25918 & ~n43300 ;
  assign n43302 = n36605 & ~n37915 ;
  assign n43304 = \P1_P2_PhyAddrPointer_reg[12]/NET0131  & n43302 ;
  assign n43303 = ~\P1_P2_PhyAddrPointer_reg[12]/NET0131  & ~n43302 ;
  assign n43305 = n25928 & ~n43303 ;
  assign n43306 = ~n43304 & n43305 ;
  assign n43293 = \P1_P2_PhyAddrPointer_reg[1]/NET0131  & n36606 ;
  assign n43294 = ~\P1_P2_PhyAddrPointer_reg[12]/NET0131  & ~n41372 ;
  assign n43295 = ~n43293 & ~n43294 ;
  assign n43296 = n27898 & n43295 ;
  assign n43307 = \P1_P2_PhyAddrPointer_reg[12]/NET0131  & ~n39352 ;
  assign n43308 = ~n40594 & ~n43307 ;
  assign n43309 = ~n43296 & n43308 ;
  assign n43310 = ~n43306 & n43309 ;
  assign n43311 = ~n43301 & n43310 ;
  assign n43312 = \P1_P2_PhyAddrPointer_reg[13]/NET0131  & n25733 ;
  assign n43313 = ~n40641 & ~n43312 ;
  assign n43314 = n25701 & ~n43313 ;
  assign n43315 = \P1_P2_PhyAddrPointer_reg[13]/NET0131  & ~n36590 ;
  assign n43316 = ~n40646 & ~n43315 ;
  assign n43317 = ~n43314 & n43316 ;
  assign n43318 = n25918 & ~n43317 ;
  assign n43322 = ~\P1_P2_PhyAddrPointer_reg[13]/NET0131  & ~n43293 ;
  assign n43323 = ~n41393 & ~n43322 ;
  assign n43324 = n36630 & n43323 ;
  assign n43319 = ~\P1_P2_PhyAddrPointer_reg[13]/NET0131  & ~n36606 ;
  assign n43320 = n25933 & ~n36607 ;
  assign n43321 = ~n43319 & n43320 ;
  assign n43325 = \P1_P2_PhyAddrPointer_reg[13]/NET0131  & ~n39352 ;
  assign n43326 = ~n40629 & ~n43325 ;
  assign n43327 = ~n43321 & n43326 ;
  assign n43328 = ~n43324 & n43327 ;
  assign n43329 = ~n43318 & n43328 ;
  assign n43334 = n25874 & ~n38947 ;
  assign n43335 = \P1_P2_PhyAddrPointer_reg[16]/NET0131  & ~n39340 ;
  assign n43336 = ~n38927 & ~n43335 ;
  assign n43337 = ~n43334 & n43336 ;
  assign n43338 = n25918 & ~n43337 ;
  assign n43330 = ~\P1_P2_PhyAddrPointer_reg[16]/NET0131  & ~n39336 ;
  assign n43331 = \P1_P2_PhyAddrPointer_reg[1]/NET0131  & n36610 ;
  assign n43332 = ~n43330 & ~n43331 ;
  assign n43339 = ~\P1_P2_DataWidth_reg[1]/NET0131  & ~n43332 ;
  assign n43340 = ~\P1_P2_PhyAddrPointer_reg[16]/NET0131  & ~n36609 ;
  assign n43341 = ~n36610 & ~n43340 ;
  assign n43342 = \P1_P2_DataWidth_reg[1]/NET0131  & ~n43341 ;
  assign n43343 = n25928 & ~n43342 ;
  assign n43344 = ~n43339 & n43343 ;
  assign n43333 = n27898 & n43332 ;
  assign n43345 = \P1_P2_PhyAddrPointer_reg[16]/NET0131  & ~n36595 ;
  assign n43346 = ~n38923 & ~n43345 ;
  assign n43347 = ~n43333 & n43346 ;
  assign n43348 = ~n43344 & n43347 ;
  assign n43349 = ~n43338 & n43348 ;
  assign n43350 = n25701 & n40704 ;
  assign n43351 = \P1_P2_PhyAddrPointer_reg[17]/NET0131  & ~n39340 ;
  assign n43352 = ~n40713 & ~n43351 ;
  assign n43353 = ~n43350 & n43352 ;
  assign n43354 = n25918 & ~n43353 ;
  assign n43358 = ~\P1_P2_PhyAddrPointer_reg[17]/NET0131  & ~n43331 ;
  assign n43359 = \P1_P2_PhyAddrPointer_reg[1]/NET0131  & n36611 ;
  assign n43360 = ~n43358 & ~n43359 ;
  assign n43361 = n36630 & n43360 ;
  assign n43355 = ~\P1_P2_PhyAddrPointer_reg[17]/NET0131  & ~n36610 ;
  assign n43356 = n25933 & ~n36611 ;
  assign n43357 = ~n43355 & n43356 ;
  assign n43362 = \P1_P2_PhyAddrPointer_reg[17]/NET0131  & ~n39352 ;
  assign n43363 = ~n40690 & ~n43362 ;
  assign n43364 = ~n43357 & n43363 ;
  assign n43365 = ~n43361 & n43364 ;
  assign n43366 = ~n43354 & n43365 ;
  assign n43374 = \P1_P2_PhyAddrPointer_reg[18]/NET0131  & n25733 ;
  assign n43375 = ~n38971 & ~n43374 ;
  assign n43376 = n25701 & ~n43375 ;
  assign n43377 = \P1_P2_PhyAddrPointer_reg[18]/NET0131  & ~n36590 ;
  assign n43378 = ~n38983 & ~n43377 ;
  assign n43379 = ~n43376 & n43378 ;
  assign n43380 = n25918 & ~n43379 ;
  assign n43370 = ~\P1_P2_PhyAddrPointer_reg[18]/NET0131  & ~n43359 ;
  assign n43371 = ~n41414 & ~n43370 ;
  assign n43372 = n36630 & n43371 ;
  assign n43367 = ~\P1_P2_PhyAddrPointer_reg[18]/NET0131  & ~n36611 ;
  assign n43368 = n25933 & ~n36612 ;
  assign n43369 = ~n43367 & n43368 ;
  assign n43373 = \P1_P2_PhyAddrPointer_reg[18]/NET0131  & ~n36595 ;
  assign n43381 = ~n38961 & ~n43373 ;
  assign n43382 = ~n43369 & n43381 ;
  assign n43383 = ~n43372 & n43382 ;
  assign n43384 = ~n43380 & n43383 ;
  assign n43385 = \P1_P2_PhyAddrPointer_reg[21]/NET0131  & n25733 ;
  assign n43386 = ~n39002 & ~n43385 ;
  assign n43387 = n25701 & ~n43386 ;
  assign n43388 = \P1_P2_PhyAddrPointer_reg[21]/NET0131  & ~n36590 ;
  assign n43389 = ~n39007 & ~n43388 ;
  assign n43390 = ~n43387 & n43389 ;
  assign n43391 = n25918 & ~n43390 ;
  assign n43396 = ~\P1_P2_PhyAddrPointer_reg[21]/NET0131  & ~n39370 ;
  assign n43397 = ~n39371 & ~n43396 ;
  assign n43398 = n27898 & n43397 ;
  assign n43392 = \P1_P2_PhyAddrPointer_reg[20]/NET0131  & n41418 ;
  assign n43393 = ~\P1_P2_PhyAddrPointer_reg[21]/NET0131  & ~n43392 ;
  assign n43394 = n25928 & ~n39363 ;
  assign n43395 = ~n43393 & n43394 ;
  assign n43399 = \P1_P2_PhyAddrPointer_reg[21]/NET0131  & ~n36595 ;
  assign n43400 = ~n39017 & ~n43399 ;
  assign n43401 = ~n43395 & n43400 ;
  assign n43402 = ~n43398 & n43401 ;
  assign n43403 = ~n43391 & n43402 ;
  assign n43404 = \P1_P2_PhyAddrPointer_reg[25]/NET0131  & n25733 ;
  assign n43405 = ~n38034 & ~n43404 ;
  assign n43406 = n25701 & ~n43405 ;
  assign n43407 = \P1_P2_PhyAddrPointer_reg[25]/NET0131  & ~n36590 ;
  assign n43408 = ~n38039 & ~n43407 ;
  assign n43409 = ~n43406 & n43408 ;
  assign n43410 = n25918 & ~n43409 ;
  assign n43414 = ~\P1_P2_PhyAddrPointer_reg[25]/NET0131  & ~n39382 ;
  assign n43415 = ~n39383 & ~n43414 ;
  assign n43416 = n36630 & n43415 ;
  assign n43411 = ~\P1_P2_PhyAddrPointer_reg[25]/NET0131  & ~n36618 ;
  assign n43412 = n25933 & ~n36619 ;
  assign n43413 = ~n43411 & n43412 ;
  assign n43417 = \P1_P2_PhyAddrPointer_reg[25]/NET0131  & ~n36595 ;
  assign n43418 = ~n38050 & ~n43417 ;
  assign n43419 = ~n43413 & n43418 ;
  assign n43420 = ~n43416 & n43419 ;
  assign n43421 = ~n43410 & n43420 ;
  assign n43422 = \P2_P1_PhyAddrPointer_reg[12]/NET0131  & n25947 ;
  assign n43423 = ~n39975 & ~n43422 ;
  assign n43424 = n25945 & ~n43423 ;
  assign n43425 = \P2_P1_PhyAddrPointer_reg[12]/NET0131  & ~n36677 ;
  assign n43426 = ~n39982 & ~n43425 ;
  assign n43427 = ~n43424 & n43426 ;
  assign n43428 = n11623 & ~n43427 ;
  assign n43434 = ~\P2_P1_PhyAddrPointer_reg[12]/NET0131  & ~n39456 ;
  assign n43435 = \P2_P1_PhyAddrPointer_reg[1]/NET0131  & n41527 ;
  assign n43436 = ~n43434 & ~n43435 ;
  assign n43437 = n11613 & n43436 ;
  assign n43429 = n36651 & ~n39474 ;
  assign n43431 = \P2_P1_PhyAddrPointer_reg[12]/NET0131  & n43429 ;
  assign n43430 = ~\P2_P1_PhyAddrPointer_reg[12]/NET0131  & ~n43429 ;
  assign n43432 = n11609 & ~n43430 ;
  assign n43433 = ~n43431 & n43432 ;
  assign n43438 = \P2_P1_PhyAddrPointer_reg[12]/NET0131  & ~n36687 ;
  assign n43439 = ~n39963 & ~n43438 ;
  assign n43440 = ~n43433 & n43439 ;
  assign n43441 = ~n43437 & n43440 ;
  assign n43442 = ~n43428 & n43441 ;
  assign n43446 = \P2_P1_PhyAddrPointer_reg[13]/NET0131  & n25947 ;
  assign n43447 = ~n40007 & ~n43446 ;
  assign n43448 = n25945 & ~n43447 ;
  assign n43449 = \P2_P1_PhyAddrPointer_reg[13]/NET0131  & ~n36677 ;
  assign n43450 = ~n40012 & ~n43449 ;
  assign n43451 = ~n43448 & n43450 ;
  assign n43452 = n11623 & ~n43451 ;
  assign n43443 = ~\P2_P1_PhyAddrPointer_reg[13]/NET0131  & ~n43435 ;
  assign n43444 = ~n39457 & ~n43443 ;
  assign n43456 = ~\P2_P1_DataWidth_reg[1]/NET0131  & ~n43444 ;
  assign n43453 = ~\P2_P1_PhyAddrPointer_reg[13]/NET0131  & ~n41527 ;
  assign n43454 = ~n41528 & ~n43453 ;
  assign n43455 = \P2_P1_DataWidth_reg[1]/NET0131  & ~n43454 ;
  assign n43457 = n11609 & ~n43455 ;
  assign n43458 = ~n43456 & n43457 ;
  assign n43445 = n11613 & n43444 ;
  assign n43459 = \P2_P1_PhyAddrPointer_reg[13]/NET0131  & ~n36687 ;
  assign n43460 = ~n39997 & ~n43459 ;
  assign n43461 = ~n43445 & n43460 ;
  assign n43462 = ~n43458 & n43461 ;
  assign n43463 = ~n43452 & n43462 ;
  assign n43464 = \P2_P1_PhyAddrPointer_reg[16]/NET0131  & n25947 ;
  assign n43465 = ~n38129 & ~n43464 ;
  assign n43466 = n25945 & ~n43465 ;
  assign n43467 = \P2_P1_PhyAddrPointer_reg[16]/NET0131  & ~n36677 ;
  assign n43468 = ~n38134 & ~n43467 ;
  assign n43469 = ~n43466 & n43468 ;
  assign n43470 = n11623 & ~n43469 ;
  assign n43474 = ~\P2_P1_PhyAddrPointer_reg[16]/NET0131  & ~n39460 ;
  assign n43475 = \P2_P1_PhyAddrPointer_reg[1]/NET0131  & n41540 ;
  assign n43476 = ~n43474 & ~n43475 ;
  assign n43477 = n36674 & n43476 ;
  assign n43473 = \P2_P1_PhyAddrPointer_reg[16]/NET0131  & ~n39451 ;
  assign n43471 = ~\P2_P1_PhyAddrPointer_reg[16]/NET0131  & n27681 ;
  assign n43472 = n36653 & n43471 ;
  assign n43478 = ~n38116 & ~n43472 ;
  assign n43479 = ~n43473 & n43478 ;
  assign n43480 = ~n43477 & n43479 ;
  assign n43481 = ~n43470 & n43480 ;
  assign n43482 = \P2_P1_PhyAddrPointer_reg[17]/NET0131  & n25947 ;
  assign n43483 = ~n40035 & ~n43482 ;
  assign n43484 = n25945 & ~n43483 ;
  assign n43485 = \P2_P1_PhyAddrPointer_reg[17]/NET0131  & ~n36677 ;
  assign n43486 = ~n40040 & ~n43485 ;
  assign n43487 = ~n43484 & n43486 ;
  assign n43488 = n11623 & ~n43487 ;
  assign n43492 = ~\P2_P1_PhyAddrPointer_reg[17]/NET0131  & ~n43475 ;
  assign n43493 = ~n41549 & ~n43492 ;
  assign n43494 = n36674 & n43493 ;
  assign n43489 = ~\P2_P1_PhyAddrPointer_reg[17]/NET0131  & ~n41540 ;
  assign n43490 = n27681 & ~n41541 ;
  assign n43491 = ~n43489 & n43490 ;
  assign n43495 = \P2_P1_PhyAddrPointer_reg[17]/NET0131  & ~n36687 ;
  assign n43496 = ~n40025 & ~n43495 ;
  assign n43497 = ~n43491 & n43496 ;
  assign n43498 = ~n43494 & n43497 ;
  assign n43499 = ~n43488 & n43498 ;
  assign n43503 = \P2_P1_PhyAddrPointer_reg[18]/NET0131  & n25947 ;
  assign n43504 = ~n38158 & ~n43503 ;
  assign n43505 = n25945 & ~n43504 ;
  assign n43506 = \P2_P1_PhyAddrPointer_reg[18]/NET0131  & ~n36677 ;
  assign n43507 = ~n38163 & ~n43506 ;
  assign n43508 = ~n43505 & n43507 ;
  assign n43509 = n11623 & ~n43508 ;
  assign n43510 = ~\P2_P1_PhyAddrPointer_reg[18]/NET0131  & ~n41542 ;
  assign n43511 = n41544 & ~n43510 ;
  assign n43500 = ~\P2_P1_PhyAddrPointer_reg[18]/NET0131  & ~n41549 ;
  assign n43501 = ~n41550 & ~n43500 ;
  assign n43502 = n11613 & n43501 ;
  assign n43512 = \P2_P1_PhyAddrPointer_reg[18]/NET0131  & ~n36687 ;
  assign n43513 = ~n38147 & ~n43512 ;
  assign n43514 = ~n43502 & n43513 ;
  assign n43515 = ~n43511 & n43514 ;
  assign n43516 = ~n43509 & n43515 ;
  assign n43523 = \P1_P2_PhyAddrPointer_reg[8]/NET0131  & n25733 ;
  assign n43524 = ~n40094 & ~n43523 ;
  assign n43525 = n25701 & ~n43524 ;
  assign n43526 = \P1_P2_PhyAddrPointer_reg[8]/NET0131  & ~n36590 ;
  assign n43527 = ~n40099 & ~n43526 ;
  assign n43528 = ~n43525 & n43527 ;
  assign n43529 = n25918 & ~n43528 ;
  assign n43517 = \P1_P2_PhyAddrPointer_reg[1]/NET0131  & n36600 ;
  assign n43518 = \P1_P2_PhyAddrPointer_reg[7]/NET0131  & n43517 ;
  assign n43519 = ~\P1_P2_PhyAddrPointer_reg[8]/NET0131  & ~n43518 ;
  assign n43520 = \P1_P2_PhyAddrPointer_reg[8]/NET0131  & n43518 ;
  assign n43521 = ~n43519 & ~n43520 ;
  assign n43530 = ~\P1_P2_DataWidth_reg[1]/NET0131  & ~n43521 ;
  assign n43531 = ~\P1_P2_PhyAddrPointer_reg[8]/NET0131  & ~n36601 ;
  assign n43532 = ~n36602 & ~n43531 ;
  assign n43533 = \P1_P2_DataWidth_reg[1]/NET0131  & ~n43532 ;
  assign n43534 = n25928 & ~n43533 ;
  assign n43535 = ~n43530 & n43534 ;
  assign n43522 = n27898 & n43521 ;
  assign n43536 = \P1_P2_PhyAddrPointer_reg[8]/NET0131  & ~n39352 ;
  assign n43537 = ~n40084 & ~n43536 ;
  assign n43538 = ~n43522 & n43537 ;
  assign n43539 = ~n43535 & n43538 ;
  assign n43540 = ~n43529 & n43539 ;
  assign n43542 = \P2_P1_PhyAddrPointer_reg[21]/NET0131  & n25947 ;
  assign n43543 = ~n38186 & ~n43542 ;
  assign n43544 = n25945 & ~n43543 ;
  assign n43545 = \P2_P1_PhyAddrPointer_reg[21]/NET0131  & ~n36677 ;
  assign n43546 = ~n38191 & ~n43545 ;
  assign n43547 = ~n43544 & n43546 ;
  assign n43548 = n11623 & ~n43547 ;
  assign n43552 = ~\P2_P1_PhyAddrPointer_reg[21]/NET0131  & ~n41577 ;
  assign n43553 = ~n41595 & ~n43552 ;
  assign n43554 = n36674 & n43553 ;
  assign n43549 = ~\P2_P1_PhyAddrPointer_reg[21]/NET0131  & ~n36658 ;
  assign n43550 = n27681 & ~n36659 ;
  assign n43551 = ~n43549 & n43550 ;
  assign n43541 = \P2_P1_PhyAddrPointer_reg[21]/NET0131  & ~n36687 ;
  assign n43555 = ~n38176 & ~n43541 ;
  assign n43556 = ~n43551 & n43555 ;
  assign n43557 = ~n43554 & n43556 ;
  assign n43558 = ~n43548 & n43557 ;
  assign n43566 = \P2_P1_PhyAddrPointer_reg[25]/NET0131  & n25947 ;
  assign n43567 = ~n38214 & ~n43566 ;
  assign n43568 = n25945 & ~n43567 ;
  assign n43569 = \P2_P1_PhyAddrPointer_reg[25]/NET0131  & ~n36677 ;
  assign n43570 = ~n38219 & ~n43569 ;
  assign n43571 = ~n43568 & n43570 ;
  assign n43572 = n11623 & ~n43571 ;
  assign n43562 = ~\P2_P1_PhyAddrPointer_reg[25]/NET0131  & ~n39496 ;
  assign n43563 = ~n39497 & ~n43562 ;
  assign n43564 = n36674 & n43563 ;
  assign n43559 = ~\P2_P1_PhyAddrPointer_reg[25]/NET0131  & ~n36661 ;
  assign n43560 = n27681 & ~n36662 ;
  assign n43561 = ~n43559 & n43560 ;
  assign n43565 = \P2_P1_PhyAddrPointer_reg[25]/NET0131  & ~n36687 ;
  assign n43573 = ~n38204 & ~n43565 ;
  assign n43574 = ~n43561 & n43573 ;
  assign n43575 = ~n43564 & n43574 ;
  assign n43576 = ~n43572 & n43575 ;
  assign n43583 = n25945 & n40066 ;
  assign n43582 = \P2_P1_PhyAddrPointer_reg[8]/NET0131  & ~n36678 ;
  assign n43584 = ~n40071 & ~n43582 ;
  assign n43585 = ~n43583 & n43584 ;
  assign n43586 = n11623 & ~n43585 ;
  assign n43587 = n36647 & ~n39474 ;
  assign n43589 = \P2_P1_PhyAddrPointer_reg[8]/NET0131  & n43587 ;
  assign n43588 = ~\P2_P1_PhyAddrPointer_reg[8]/NET0131  & ~n43587 ;
  assign n43590 = n11609 & ~n43588 ;
  assign n43591 = ~n43589 & n43590 ;
  assign n43577 = \P2_P1_PhyAddrPointer_reg[1]/NET0131  & n36646 ;
  assign n43578 = \P2_P1_PhyAddrPointer_reg[7]/NET0131  & n43577 ;
  assign n43579 = ~\P2_P1_PhyAddrPointer_reg[8]/NET0131  & ~n43578 ;
  assign n43580 = ~n39454 & ~n43579 ;
  assign n43581 = n11613 & n43580 ;
  assign n43592 = \P2_P1_PhyAddrPointer_reg[8]/NET0131  & ~n36687 ;
  assign n43593 = ~n40053 & ~n43592 ;
  assign n43594 = ~n43581 & n43593 ;
  assign n43595 = ~n43591 & n43594 ;
  assign n43596 = ~n43586 & n43595 ;
  assign n43600 = n26126 & n40320 ;
  assign n43601 = \P1_P1_PhyAddrPointer_reg[12]/NET0131  & ~n41658 ;
  assign n43602 = ~n40325 & ~n43601 ;
  assign n43603 = ~n43600 & n43602 ;
  assign n43604 = n8355 & ~n43603 ;
  assign n43607 = n36711 & ~n39569 ;
  assign n43605 = n36710 & ~n39569 ;
  assign n43606 = ~\P1_P1_PhyAddrPointer_reg[12]/NET0131  & ~n43605 ;
  assign n43608 = n8282 & ~n43606 ;
  assign n43609 = ~n43607 & n43608 ;
  assign n43597 = ~\P1_P1_PhyAddrPointer_reg[12]/NET0131  & ~n41670 ;
  assign n43598 = ~n39557 & ~n43597 ;
  assign n43599 = n8287 & n43598 ;
  assign n43610 = \P1_P1_PhyAddrPointer_reg[12]/NET0131  & ~n36743 ;
  assign n43611 = ~n40307 & ~n43610 ;
  assign n43612 = ~n43599 & n43611 ;
  assign n43613 = ~n43609 & n43612 ;
  assign n43614 = ~n43604 & n43613 ;
  assign n43618 = \P1_P1_PhyAddrPointer_reg[13]/NET0131  & n26249 ;
  assign n43619 = ~n40378 & ~n43618 ;
  assign n43620 = n26126 & ~n43619 ;
  assign n43621 = \P1_P1_PhyAddrPointer_reg[13]/NET0131  & ~n36696 ;
  assign n43622 = ~n40383 & ~n43621 ;
  assign n43623 = ~n43620 & n43622 ;
  assign n43624 = n8355 & ~n43623 ;
  assign n43615 = ~\P1_P1_PhyAddrPointer_reg[13]/NET0131  & ~n39557 ;
  assign n43616 = ~n39558 & ~n43615 ;
  assign n43625 = ~\P1_P1_DataWidth_reg[1]/NET0131  & ~n43616 ;
  assign n43626 = ~\P1_P1_PhyAddrPointer_reg[13]/NET0131  & ~n36711 ;
  assign n43627 = ~n36712 & ~n43626 ;
  assign n43628 = \P1_P1_DataWidth_reg[1]/NET0131  & ~n43627 ;
  assign n43629 = n8282 & ~n43628 ;
  assign n43630 = ~n43625 & n43629 ;
  assign n43617 = n8287 & n43616 ;
  assign n43631 = \P1_P1_PhyAddrPointer_reg[13]/NET0131  & ~n36743 ;
  assign n43632 = ~n40368 & ~n43631 ;
  assign n43633 = ~n43617 & n43632 ;
  assign n43634 = ~n43630 & n43633 ;
  assign n43635 = ~n43624 & n43634 ;
  assign n43636 = \P1_P1_PhyAddrPointer_reg[16]/NET0131  & n26249 ;
  assign n43637 = ~n38732 & ~n43636 ;
  assign n43638 = n26126 & ~n43637 ;
  assign n43639 = \P1_P1_PhyAddrPointer_reg[16]/NET0131  & ~n36696 ;
  assign n43640 = ~n38737 & ~n43639 ;
  assign n43641 = ~n43638 & n43640 ;
  assign n43642 = n8355 & ~n43641 ;
  assign n43646 = ~\P1_P1_PhyAddrPointer_reg[16]/NET0131  & ~n39561 ;
  assign n43647 = ~n41711 & ~n43646 ;
  assign n43648 = ~n36701 & n43647 ;
  assign n43643 = ~\P1_P1_PhyAddrPointer_reg[16]/NET0131  & ~n36714 ;
  assign n43644 = n27791 & ~n36715 ;
  assign n43645 = ~n43643 & n43644 ;
  assign n43649 = \P1_P1_PhyAddrPointer_reg[16]/NET0131  & ~n36743 ;
  assign n43650 = ~n38722 & ~n43649 ;
  assign n43651 = ~n43645 & n43650 ;
  assign n43652 = ~n43648 & n43651 ;
  assign n43653 = ~n43642 & n43652 ;
  assign n43654 = \P1_P1_PhyAddrPointer_reg[17]/NET0131  & n26249 ;
  assign n43655 = ~n40528 & ~n43654 ;
  assign n43656 = n26126 & ~n43655 ;
  assign n43657 = \P1_P1_PhyAddrPointer_reg[17]/NET0131  & ~n36696 ;
  assign n43658 = ~n40533 & ~n43657 ;
  assign n43659 = ~n43656 & n43658 ;
  assign n43660 = n8355 & ~n43659 ;
  assign n43664 = ~\P1_P1_PhyAddrPointer_reg[17]/NET0131  & ~n41711 ;
  assign n43665 = ~n41712 & ~n43664 ;
  assign n43666 = ~n36701 & n43665 ;
  assign n43661 = ~\P1_P1_PhyAddrPointer_reg[17]/NET0131  & ~n36715 ;
  assign n43662 = n27791 & ~n36716 ;
  assign n43663 = ~n43661 & n43662 ;
  assign n43667 = \P1_P1_PhyAddrPointer_reg[17]/NET0131  & ~n36743 ;
  assign n43668 = ~n40518 & ~n43667 ;
  assign n43669 = ~n43663 & n43668 ;
  assign n43670 = ~n43666 & n43669 ;
  assign n43671 = ~n43660 & n43670 ;
  assign n43672 = \P1_P1_PhyAddrPointer_reg[18]/NET0131  & n26249 ;
  assign n43673 = ~n38762 & ~n43672 ;
  assign n43674 = n26126 & ~n43673 ;
  assign n43675 = \P1_P1_PhyAddrPointer_reg[18]/NET0131  & ~n36696 ;
  assign n43676 = ~n38769 & ~n43675 ;
  assign n43677 = ~n43674 & n43676 ;
  assign n43678 = n8355 & ~n43677 ;
  assign n43682 = ~\P1_P1_PhyAddrPointer_reg[18]/NET0131  & ~n41712 ;
  assign n43683 = ~n41713 & ~n43682 ;
  assign n43684 = ~n36701 & n43683 ;
  assign n43679 = ~\P1_P1_PhyAddrPointer_reg[18]/NET0131  & ~n36716 ;
  assign n43680 = n27791 & ~n36717 ;
  assign n43681 = ~n43679 & n43680 ;
  assign n43685 = \P1_P1_PhyAddrPointer_reg[18]/NET0131  & ~n36743 ;
  assign n43686 = ~n38750 & ~n43685 ;
  assign n43687 = ~n43681 & n43686 ;
  assign n43688 = ~n43684 & n43687 ;
  assign n43689 = ~n43678 & n43688 ;
  assign n43690 = \P1_P1_PhyAddrPointer_reg[21]/NET0131  & n26249 ;
  assign n43691 = ~n38794 & ~n43690 ;
  assign n43692 = n26126 & ~n43691 ;
  assign n43693 = \P1_P1_PhyAddrPointer_reg[21]/NET0131  & ~n36696 ;
  assign n43694 = ~n38799 & ~n43693 ;
  assign n43695 = ~n43692 & n43694 ;
  assign n43696 = n8355 & ~n43695 ;
  assign n43700 = ~\P1_P1_PhyAddrPointer_reg[21]/NET0131  & ~n41732 ;
  assign n43701 = ~n41743 & ~n43700 ;
  assign n43702 = ~n36701 & n43701 ;
  assign n43697 = ~\P1_P1_PhyAddrPointer_reg[21]/NET0131  & ~n36719 ;
  assign n43698 = n27791 & ~n36720 ;
  assign n43699 = ~n43697 & n43698 ;
  assign n43703 = \P1_P1_PhyAddrPointer_reg[21]/NET0131  & ~n36743 ;
  assign n43704 = ~n38814 & ~n43703 ;
  assign n43705 = ~n43699 & n43704 ;
  assign n43706 = ~n43702 & n43705 ;
  assign n43707 = ~n43696 & n43706 ;
  assign n43709 = \P1_P1_PhyAddrPointer_reg[25]/NET0131  & n26249 ;
  assign n43710 = ~n38827 & ~n43709 ;
  assign n43711 = n26126 & ~n43710 ;
  assign n43712 = \P1_P1_PhyAddrPointer_reg[25]/NET0131  & ~n36696 ;
  assign n43713 = ~n38838 & ~n43712 ;
  assign n43714 = ~n43711 & n43713 ;
  assign n43715 = n8355 & ~n43714 ;
  assign n43716 = ~\P1_P1_PhyAddrPointer_reg[25]/NET0131  & ~n41771 ;
  assign n43717 = ~n41788 & ~n43716 ;
  assign n43718 = ~n36701 & n43717 ;
  assign n43719 = ~\P1_P1_PhyAddrPointer_reg[25]/NET0131  & ~n36723 ;
  assign n43720 = n41783 & ~n43719 ;
  assign n43708 = \P1_P1_PhyAddrPointer_reg[25]/NET0131  & ~n36743 ;
  assign n43721 = ~n38817 & ~n43708 ;
  assign n43722 = ~n43720 & n43721 ;
  assign n43723 = ~n43718 & n43722 ;
  assign n43724 = ~n43715 & n43723 ;
  assign n43725 = \P1_P1_PhyAddrPointer_reg[8]/NET0131  & n26249 ;
  assign n43726 = ~n40672 & ~n43725 ;
  assign n43727 = n26126 & ~n43726 ;
  assign n43728 = \P1_P1_PhyAddrPointer_reg[8]/NET0131  & ~n36696 ;
  assign n43729 = ~n40677 & ~n43728 ;
  assign n43730 = ~n43727 & n43729 ;
  assign n43731 = n8355 & ~n43730 ;
  assign n43737 = \P1_P1_PhyAddrPointer_reg[1]/NET0131  & n36705 ;
  assign n43738 = \P1_P1_PhyAddrPointer_reg[7]/NET0131  & n43737 ;
  assign n43739 = ~\P1_P1_PhyAddrPointer_reg[8]/NET0131  & ~n43738 ;
  assign n43740 = ~n41666 & ~n43739 ;
  assign n43741 = n8287 & n43740 ;
  assign n43732 = n36706 & ~n39569 ;
  assign n43734 = \P1_P1_PhyAddrPointer_reg[8]/NET0131  & n43732 ;
  assign n43733 = ~\P1_P1_PhyAddrPointer_reg[8]/NET0131  & ~n43732 ;
  assign n43735 = n8282 & ~n43733 ;
  assign n43736 = ~n43734 & n43735 ;
  assign n43742 = \P1_P1_PhyAddrPointer_reg[8]/NET0131  & ~n36743 ;
  assign n43743 = ~n40659 & ~n43742 ;
  assign n43744 = ~n43736 & n43743 ;
  assign n43745 = ~n43741 & n43744 ;
  assign n43746 = ~n43731 & n43745 ;
  assign n43747 = \P2_P2_PhyAddrPointer_reg[12]/NET0131  & n26629 ;
  assign n43748 = ~n40150 & ~n43747 ;
  assign n43749 = n26621 & ~n43748 ;
  assign n43750 = \P2_P2_PhyAddrPointer_reg[12]/NET0131  & ~n36752 ;
  assign n43751 = ~n40158 & ~n43750 ;
  assign n43752 = ~n43749 & n43751 ;
  assign n43753 = n26792 & ~n43752 ;
  assign n43757 = ~\P2_P2_PhyAddrPointer_reg[12]/NET0131  & ~n41818 ;
  assign n43758 = ~n39647 & ~n43757 ;
  assign n43759 = ~n36760 & n43758 ;
  assign n43754 = ~\P2_P2_PhyAddrPointer_reg[12]/NET0131  & ~n36769 ;
  assign n43755 = n26800 & ~n36770 ;
  assign n43756 = ~n43754 & n43755 ;
  assign n43760 = \P2_P2_PhyAddrPointer_reg[12]/NET0131  & ~n36758 ;
  assign n43761 = ~n40140 & ~n43760 ;
  assign n43762 = ~n43756 & n43761 ;
  assign n43763 = ~n43759 & n43762 ;
  assign n43764 = ~n43753 & n43763 ;
  assign n43768 = \P2_P2_PhyAddrPointer_reg[13]/NET0131  & n26629 ;
  assign n43769 = ~n40184 & ~n43768 ;
  assign n43770 = n26621 & ~n43769 ;
  assign n43771 = \P2_P2_PhyAddrPointer_reg[13]/NET0131  & ~n36752 ;
  assign n43772 = ~n40189 & ~n43771 ;
  assign n43773 = ~n43770 & n43772 ;
  assign n43774 = n26792 & ~n43773 ;
  assign n43765 = ~\P2_P2_PhyAddrPointer_reg[13]/NET0131  & ~n39647 ;
  assign n43766 = ~n39648 & ~n43765 ;
  assign n43775 = ~\P2_P2_DataWidth_reg[1]/NET0131  & ~n43766 ;
  assign n43776 = ~\P2_P2_PhyAddrPointer_reg[13]/NET0131  & ~n36770 ;
  assign n43777 = ~n36771 & ~n43776 ;
  assign n43778 = \P2_P2_DataWidth_reg[1]/NET0131  & ~n43777 ;
  assign n43779 = n26794 & ~n43778 ;
  assign n43780 = ~n43775 & n43779 ;
  assign n43767 = n27977 & n43766 ;
  assign n43781 = \P2_P2_PhyAddrPointer_reg[13]/NET0131  & ~n36758 ;
  assign n43782 = ~n40174 & ~n43781 ;
  assign n43783 = ~n43767 & n43782 ;
  assign n43784 = ~n43780 & n43783 ;
  assign n43785 = ~n43774 & n43784 ;
  assign n43786 = n26621 & n38321 ;
  assign n43787 = \P2_P2_PhyAddrPointer_reg[16]/NET0131  & ~n41873 ;
  assign n43788 = ~n38328 & ~n43787 ;
  assign n43789 = ~n43786 & n43788 ;
  assign n43790 = n26792 & ~n43789 ;
  assign n43794 = ~\P2_P2_PhyAddrPointer_reg[16]/NET0131  & ~n39651 ;
  assign n43795 = \P2_P2_PhyAddrPointer_reg[16]/NET0131  & n39651 ;
  assign n43796 = ~n43794 & ~n43795 ;
  assign n43797 = ~n36760 & n43796 ;
  assign n43791 = ~\P2_P2_PhyAddrPointer_reg[16]/NET0131  & ~n36773 ;
  assign n43792 = n26800 & ~n36774 ;
  assign n43793 = ~n43791 & n43792 ;
  assign n43798 = \P2_P2_PhyAddrPointer_reg[16]/NET0131  & ~n36758 ;
  assign n43799 = ~n38310 & ~n43798 ;
  assign n43800 = ~n43793 & n43799 ;
  assign n43801 = ~n43797 & n43800 ;
  assign n43802 = ~n43790 & n43801 ;
  assign n43803 = \P2_P2_PhyAddrPointer_reg[17]/NET0131  & n26629 ;
  assign n43804 = ~n40216 & ~n43803 ;
  assign n43805 = n26621 & ~n43804 ;
  assign n43806 = \P2_P2_PhyAddrPointer_reg[17]/NET0131  & ~n36752 ;
  assign n43807 = ~n40221 & ~n43806 ;
  assign n43808 = ~n43805 & n43807 ;
  assign n43809 = n26792 & ~n43808 ;
  assign n43813 = ~\P2_P2_PhyAddrPointer_reg[17]/NET0131  & ~n43795 ;
  assign n43814 = ~n41857 & ~n43813 ;
  assign n43815 = ~n36760 & n43814 ;
  assign n43810 = ~\P2_P2_PhyAddrPointer_reg[17]/NET0131  & ~n36774 ;
  assign n43811 = n26800 & ~n36775 ;
  assign n43812 = ~n43810 & n43811 ;
  assign n43816 = \P2_P2_PhyAddrPointer_reg[17]/NET0131  & ~n36758 ;
  assign n43817 = ~n40202 & ~n43816 ;
  assign n43818 = ~n43812 & n43817 ;
  assign n43819 = ~n43815 & n43818 ;
  assign n43820 = ~n43809 & n43819 ;
  assign n43821 = \P2_P2_PhyAddrPointer_reg[18]/NET0131  & n26629 ;
  assign n43822 = ~n38358 & ~n43821 ;
  assign n43823 = n26621 & ~n43822 ;
  assign n43824 = \P2_P2_PhyAddrPointer_reg[18]/NET0131  & ~n36752 ;
  assign n43825 = ~n38365 & ~n43824 ;
  assign n43826 = ~n43823 & n43825 ;
  assign n43827 = n26792 & ~n43826 ;
  assign n43831 = ~\P2_P2_PhyAddrPointer_reg[18]/NET0131  & ~n41857 ;
  assign n43832 = ~n41858 & ~n43831 ;
  assign n43833 = ~n36760 & n43832 ;
  assign n43828 = ~\P2_P2_PhyAddrPointer_reg[18]/NET0131  & ~n36775 ;
  assign n43829 = n26800 & ~n36776 ;
  assign n43830 = ~n43828 & n43829 ;
  assign n43834 = \P2_P2_PhyAddrPointer_reg[18]/NET0131  & ~n36758 ;
  assign n43835 = ~n38343 & ~n43834 ;
  assign n43836 = ~n43830 & n43835 ;
  assign n43837 = ~n43833 & n43836 ;
  assign n43838 = ~n43827 & n43837 ;
  assign n43839 = \P2_P2_PhyAddrPointer_reg[21]/NET0131  & n26629 ;
  assign n43840 = ~n38391 & ~n43839 ;
  assign n43841 = n26621 & ~n43840 ;
  assign n43842 = \P2_P2_PhyAddrPointer_reg[21]/NET0131  & ~n36752 ;
  assign n43843 = ~n38404 & ~n43842 ;
  assign n43844 = ~n43841 & n43843 ;
  assign n43845 = n26792 & ~n43844 ;
  assign n43849 = ~\P2_P2_PhyAddrPointer_reg[21]/NET0131  & ~n41869 ;
  assign n43850 = ~n41898 & ~n43849 ;
  assign n43851 = ~n36760 & n43850 ;
  assign n43846 = ~\P2_P2_PhyAddrPointer_reg[21]/NET0131  & ~n36778 ;
  assign n43847 = n26800 & ~n36779 ;
  assign n43848 = ~n43846 & n43847 ;
  assign n43852 = \P2_P2_PhyAddrPointer_reg[21]/NET0131  & ~n36758 ;
  assign n43853 = ~n38378 & ~n43852 ;
  assign n43854 = ~n43848 & n43853 ;
  assign n43855 = ~n43851 & n43854 ;
  assign n43856 = ~n43845 & n43855 ;
  assign n43857 = \P2_P2_PhyAddrPointer_reg[25]/NET0131  & n26629 ;
  assign n43858 = ~n38423 & ~n43857 ;
  assign n43859 = n26621 & ~n43858 ;
  assign n43860 = \P2_P2_PhyAddrPointer_reg[25]/NET0131  & ~n36752 ;
  assign n43861 = ~n43859 & ~n43860 ;
  assign n43862 = ~n38434 & n43861 ;
  assign n43863 = n26792 & ~n43862 ;
  assign n43867 = ~\P2_P2_PhyAddrPointer_reg[25]/NET0131  & ~n41916 ;
  assign n43868 = ~n39702 & ~n43867 ;
  assign n43869 = ~n36760 & n43868 ;
  assign n43864 = ~\P2_P2_PhyAddrPointer_reg[25]/NET0131  & ~n36782 ;
  assign n43865 = n26800 & ~n36783 ;
  assign n43866 = ~n43864 & n43865 ;
  assign n43870 = \P2_P2_PhyAddrPointer_reg[25]/NET0131  & ~n36758 ;
  assign n43871 = ~n38413 & ~n43870 ;
  assign n43872 = ~n43866 & n43871 ;
  assign n43873 = ~n43869 & n43872 ;
  assign n43874 = ~n43863 & n43873 ;
  assign n43876 = n26621 & n40251 ;
  assign n43875 = \P2_P2_PhyAddrPointer_reg[8]/NET0131  & ~n41873 ;
  assign n43877 = ~n40256 & ~n43875 ;
  assign n43878 = ~n43876 & n43877 ;
  assign n43879 = n26792 & ~n43878 ;
  assign n43883 = ~\P2_P2_PhyAddrPointer_reg[8]/NET0131  & ~n41813 ;
  assign n43884 = ~n41814 & ~n43883 ;
  assign n43885 = ~n36760 & n43884 ;
  assign n43880 = ~\P2_P2_PhyAddrPointer_reg[8]/NET0131  & ~n36765 ;
  assign n43881 = n26800 & ~n36766 ;
  assign n43882 = ~n43880 & n43881 ;
  assign n43886 = \P2_P2_PhyAddrPointer_reg[8]/NET0131  & ~n36758 ;
  assign n43887 = ~n40239 & ~n43886 ;
  assign n43888 = ~n43882 & n43887 ;
  assign n43889 = ~n43885 & n43888 ;
  assign n43890 = ~n43879 & n43889 ;
  assign n43892 = \P1_P3_PhyAddrPointer_reg[12]/NET0131  & n9072 ;
  assign n43893 = ~n19579 & ~n43892 ;
  assign n43894 = n9064 & ~n43893 ;
  assign n43895 = \P1_P3_PhyAddrPointer_reg[12]/NET0131  & ~n36805 ;
  assign n43896 = ~n19586 & ~n43895 ;
  assign n43897 = ~n43894 & n43896 ;
  assign n43898 = n9241 & ~n43897 ;
  assign n43899 = ~\P1_P3_DataWidth_reg[1]/NET0131  & ~n17719 ;
  assign n43900 = ~\P1_P3_PhyAddrPointer_reg[12]/NET0131  & ~n16461 ;
  assign n43901 = ~n16462 & ~n43900 ;
  assign n43902 = \P1_P3_DataWidth_reg[1]/NET0131  & ~n43901 ;
  assign n43903 = n9245 & ~n43902 ;
  assign n43904 = ~n43899 & n43903 ;
  assign n43891 = n16492 & n17719 ;
  assign n43905 = \P1_P3_PhyAddrPointer_reg[12]/NET0131  & ~n36816 ;
  assign n43906 = ~n19567 & ~n43905 ;
  assign n43907 = ~n43891 & n43906 ;
  assign n43908 = ~n43904 & n43907 ;
  assign n43909 = ~n43898 & n43908 ;
  assign n43911 = n9192 & ~n19452 ;
  assign n43912 = \P1_P3_PhyAddrPointer_reg[13]/NET0131  & ~n37992 ;
  assign n43913 = ~n19465 & ~n43912 ;
  assign n43914 = ~n43911 & n43913 ;
  assign n43915 = n9241 & ~n43914 ;
  assign n43916 = ~\P1_P3_DataWidth_reg[1]/NET0131  & ~n17754 ;
  assign n43917 = ~\P1_P3_PhyAddrPointer_reg[13]/NET0131  & ~n16462 ;
  assign n43918 = ~n16463 & ~n43917 ;
  assign n43919 = \P1_P3_DataWidth_reg[1]/NET0131  & ~n43918 ;
  assign n43920 = n9245 & ~n43919 ;
  assign n43921 = ~n43916 & n43920 ;
  assign n43910 = n16492 & n17754 ;
  assign n43922 = \P1_P3_PhyAddrPointer_reg[13]/NET0131  & ~n36816 ;
  assign n43923 = ~n19429 & ~n43922 ;
  assign n43924 = ~n43910 & n43923 ;
  assign n43925 = ~n43921 & n43924 ;
  assign n43926 = ~n43915 & n43925 ;
  assign n43928 = \P1_P3_PhyAddrPointer_reg[16]/NET0131  & n9072 ;
  assign n43929 = ~n19629 & ~n43928 ;
  assign n43930 = n9064 & ~n43929 ;
  assign n43931 = \P1_P3_PhyAddrPointer_reg[16]/NET0131  & ~n36805 ;
  assign n43932 = ~n19638 & ~n43931 ;
  assign n43933 = ~n43930 & n43932 ;
  assign n43934 = n9241 & ~n43933 ;
  assign n43935 = ~\P1_P3_DataWidth_reg[1]/NET0131  & ~n17830 ;
  assign n43936 = ~\P1_P3_PhyAddrPointer_reg[16]/NET0131  & ~n16465 ;
  assign n43937 = ~n16466 & ~n43936 ;
  assign n43938 = \P1_P3_DataWidth_reg[1]/NET0131  & ~n43937 ;
  assign n43939 = n9245 & ~n43938 ;
  assign n43940 = ~n43935 & n43939 ;
  assign n43927 = n16492 & n17830 ;
  assign n43941 = \P1_P3_PhyAddrPointer_reg[16]/NET0131  & ~n36816 ;
  assign n43942 = ~n19608 & ~n43941 ;
  assign n43943 = ~n43927 & n43942 ;
  assign n43944 = ~n43940 & n43943 ;
  assign n43945 = ~n43934 & n43944 ;
  assign n43946 = \P1_P3_PhyAddrPointer_reg[17]/NET0131  & n9072 ;
  assign n43947 = ~n19687 & ~n43946 ;
  assign n43948 = n9064 & ~n43947 ;
  assign n43949 = \P1_P3_PhyAddrPointer_reg[17]/NET0131  & ~n36805 ;
  assign n43950 = ~n19693 & ~n43949 ;
  assign n43951 = ~n43948 & n43950 ;
  assign n43952 = n9241 & ~n43951 ;
  assign n43956 = n16546 & ~n36810 ;
  assign n43953 = ~\P1_P3_PhyAddrPointer_reg[17]/NET0131  & ~n16466 ;
  assign n43954 = n11698 & ~n16467 ;
  assign n43955 = ~n43953 & n43954 ;
  assign n43957 = \P1_P3_PhyAddrPointer_reg[17]/NET0131  & ~n36816 ;
  assign n43958 = ~n19665 & ~n43957 ;
  assign n43959 = ~n43955 & n43958 ;
  assign n43960 = ~n43956 & n43959 ;
  assign n43961 = ~n43952 & n43960 ;
  assign n43962 = \P1_P3_PhyAddrPointer_reg[18]/NET0131  & n9072 ;
  assign n43963 = ~n19726 & ~n43962 ;
  assign n43964 = n9064 & ~n43963 ;
  assign n43965 = \P1_P3_PhyAddrPointer_reg[18]/NET0131  & ~n36805 ;
  assign n43966 = ~n19735 & ~n43965 ;
  assign n43967 = ~n43964 & n43966 ;
  assign n43968 = n9241 & ~n43967 ;
  assign n43972 = n16553 & ~n36810 ;
  assign n43969 = ~\P1_P3_PhyAddrPointer_reg[18]/NET0131  & ~n16467 ;
  assign n43970 = n11698 & ~n16468 ;
  assign n43971 = ~n43969 & n43970 ;
  assign n43973 = \P1_P3_PhyAddrPointer_reg[18]/NET0131  & ~n36816 ;
  assign n43974 = ~n19706 & ~n43973 ;
  assign n43975 = ~n43971 & n43974 ;
  assign n43976 = ~n43972 & n43975 ;
  assign n43977 = ~n43968 & n43976 ;
  assign n43978 = n9064 & n19875 ;
  assign n43979 = \P1_P3_PhyAddrPointer_reg[21]/NET0131  & ~n37992 ;
  assign n43980 = ~n19885 & ~n43979 ;
  assign n43981 = ~n43978 & n43980 ;
  assign n43982 = n9241 & ~n43981 ;
  assign n43986 = n16630 & ~n36810 ;
  assign n43983 = ~\P1_P3_PhyAddrPointer_reg[21]/NET0131  & ~n16470 ;
  assign n43984 = n11698 & ~n16471 ;
  assign n43985 = ~n43983 & n43984 ;
  assign n43987 = \P1_P3_PhyAddrPointer_reg[21]/NET0131  & ~n36816 ;
  assign n43988 = ~n19845 & ~n43987 ;
  assign n43989 = ~n43985 & n43988 ;
  assign n43990 = ~n43986 & n43989 ;
  assign n43991 = ~n43982 & n43990 ;
  assign n43992 = \P1_P3_PhyAddrPointer_reg[25]/NET0131  & n9072 ;
  assign n43993 = ~n20063 & ~n43992 ;
  assign n43994 = n9064 & ~n43993 ;
  assign n43995 = \P1_P3_PhyAddrPointer_reg[25]/NET0131  & ~n36805 ;
  assign n43996 = ~n20069 & ~n43995 ;
  assign n43997 = ~n43994 & n43996 ;
  assign n43998 = n9241 & ~n43997 ;
  assign n44002 = n16794 & ~n36810 ;
  assign n43999 = ~\P1_P3_PhyAddrPointer_reg[25]/NET0131  & ~n16474 ;
  assign n44000 = n11698 & ~n16475 ;
  assign n44001 = ~n43999 & n44000 ;
  assign n44003 = \P1_P3_PhyAddrPointer_reg[25]/NET0131  & ~n36816 ;
  assign n44004 = ~n20039 & ~n44003 ;
  assign n44005 = ~n44001 & n44004 ;
  assign n44006 = ~n44002 & n44005 ;
  assign n44007 = ~n43998 & n44006 ;
  assign n44008 = \P1_P3_PhyAddrPointer_reg[8]/NET0131  & n9072 ;
  assign n44009 = ~n20597 & ~n44008 ;
  assign n44010 = n9064 & ~n44009 ;
  assign n44011 = \P1_P3_PhyAddrPointer_reg[8]/NET0131  & ~n36805 ;
  assign n44012 = ~n20602 & ~n44011 ;
  assign n44013 = ~n44010 & n44012 ;
  assign n44014 = n9241 & ~n44013 ;
  assign n44018 = n17938 & ~n36810 ;
  assign n44015 = ~\P1_P3_PhyAddrPointer_reg[8]/NET0131  & ~n16457 ;
  assign n44016 = n11698 & ~n16458 ;
  assign n44017 = ~n44015 & n44016 ;
  assign n44019 = \P1_P3_PhyAddrPointer_reg[8]/NET0131  & ~n36816 ;
  assign n44020 = ~n20587 & ~n44019 ;
  assign n44021 = ~n44017 & n44020 ;
  assign n44022 = ~n44018 & n44021 ;
  assign n44023 = ~n44014 & n44022 ;
  assign n44025 = \P2_P3_PhyAddrPointer_reg[12]/NET0131  & ~n27283 ;
  assign n44026 = ~n40406 & ~n44025 ;
  assign n44027 = n27117 & ~n44026 ;
  assign n44028 = \P2_P3_PhyAddrPointer_reg[12]/NET0131  & ~n36826 ;
  assign n44029 = ~n40413 & ~n44028 ;
  assign n44030 = ~n44027 & n44029 ;
  assign n44031 = n27308 & ~n44030 ;
  assign n44036 = n36841 & ~n39862 ;
  assign n44037 = \P2_P3_PhyAddrPointer_reg[10]/NET0131  & n44036 ;
  assign n44038 = \P2_P3_PhyAddrPointer_reg[11]/NET0131  & n44037 ;
  assign n44040 = ~\P2_P3_PhyAddrPointer_reg[12]/NET0131  & ~n44038 ;
  assign n44039 = \P2_P3_PhyAddrPointer_reg[12]/NET0131  & n44038 ;
  assign n44041 = n27315 & ~n44039 ;
  assign n44042 = ~n44040 & n44041 ;
  assign n44032 = ~\P2_P3_PhyAddrPointer_reg[12]/NET0131  & ~n39841 ;
  assign n44033 = \P2_P3_PhyAddrPointer_reg[12]/NET0131  & n39841 ;
  assign n44034 = ~n44032 & ~n44033 ;
  assign n44035 = n32867 & n44034 ;
  assign n44024 = \P2_P3_PhyAddrPointer_reg[12]/NET0131  & ~n36873 ;
  assign n44043 = ~n40396 & ~n44024 ;
  assign n44044 = ~n44035 & n44043 ;
  assign n44045 = ~n44042 & n44044 ;
  assign n44046 = ~n44031 & n44045 ;
  assign n44048 = \P2_P3_PhyAddrPointer_reg[13]/NET0131  & ~n27283 ;
  assign n44049 = ~n40438 & ~n44048 ;
  assign n44050 = n27117 & ~n44049 ;
  assign n44051 = \P2_P3_PhyAddrPointer_reg[13]/NET0131  & ~n36826 ;
  assign n44052 = ~n40443 & ~n44051 ;
  assign n44053 = ~n44050 & n44052 ;
  assign n44054 = n27308 & ~n44053 ;
  assign n44055 = ~\P2_P3_PhyAddrPointer_reg[13]/NET0131  & ~n44033 ;
  assign n44056 = ~n39842 & ~n44055 ;
  assign n44057 = ~n36831 & n44056 ;
  assign n44058 = ~\P2_P3_PhyAddrPointer_reg[13]/NET0131  & ~n36844 ;
  assign n44059 = n42080 & ~n44058 ;
  assign n44047 = \P2_P3_PhyAddrPointer_reg[13]/NET0131  & ~n36873 ;
  assign n44060 = ~n40428 & ~n44047 ;
  assign n44061 = ~n44059 & n44060 ;
  assign n44062 = ~n44057 & n44061 ;
  assign n44063 = ~n44054 & n44062 ;
  assign n44072 = \P2_P3_PhyAddrPointer_reg[16]/NET0131  & ~n27283 ;
  assign n44073 = ~n38562 & ~n44072 ;
  assign n44074 = n27117 & ~n44073 ;
  assign n44075 = \P2_P3_PhyAddrPointer_reg[16]/NET0131  & ~n36826 ;
  assign n44076 = ~n38570 & ~n44075 ;
  assign n44077 = ~n44074 & n44076 ;
  assign n44078 = n27308 & ~n44077 ;
  assign n44068 = ~\P2_P3_PhyAddrPointer_reg[16]/NET0131  & ~n39846 ;
  assign n44069 = \P2_P3_PhyAddrPointer_reg[16]/NET0131  & n39846 ;
  assign n44070 = ~n44068 & ~n44069 ;
  assign n44071 = ~n36831 & n44070 ;
  assign n44064 = n36873 & ~n39850 ;
  assign n44065 = \P2_P3_PhyAddrPointer_reg[16]/NET0131  & ~n44064 ;
  assign n44066 = ~\P2_P3_PhyAddrPointer_reg[16]/NET0131  & n27325 ;
  assign n44067 = n39845 & n44066 ;
  assign n44079 = ~n38552 & ~n44067 ;
  assign n44080 = ~n44065 & n44079 ;
  assign n44081 = ~n44071 & n44080 ;
  assign n44082 = ~n44078 & n44081 ;
  assign n44083 = \P2_P3_PhyAddrPointer_reg[17]/NET0131  & ~n27283 ;
  assign n44084 = ~n40468 & ~n44083 ;
  assign n44085 = n27117 & ~n44084 ;
  assign n44086 = \P2_P3_PhyAddrPointer_reg[17]/NET0131  & ~n36826 ;
  assign n44087 = ~n40473 & ~n44086 ;
  assign n44088 = ~n44085 & n44087 ;
  assign n44089 = n27308 & ~n44088 ;
  assign n44094 = ~\P2_P3_PhyAddrPointer_reg[17]/NET0131  & ~n44069 ;
  assign n44095 = n36848 & n39846 ;
  assign n44096 = ~n44094 & ~n44095 ;
  assign n44097 = ~n36831 & n44096 ;
  assign n44090 = \P2_P3_PhyAddrPointer_reg[16]/NET0131  & n39845 ;
  assign n44091 = ~\P2_P3_PhyAddrPointer_reg[17]/NET0131  & ~n44090 ;
  assign n44092 = n27325 & ~n42106 ;
  assign n44093 = ~n44091 & n44092 ;
  assign n44098 = \P2_P3_PhyAddrPointer_reg[17]/NET0131  & ~n36873 ;
  assign n44099 = ~n40456 & ~n44098 ;
  assign n44100 = ~n44093 & n44099 ;
  assign n44101 = ~n44097 & n44100 ;
  assign n44102 = ~n44089 & n44101 ;
  assign n44104 = \P2_P3_PhyAddrPointer_reg[18]/NET0131  & ~n27283 ;
  assign n44105 = ~n38596 & ~n44104 ;
  assign n44106 = n27117 & ~n44105 ;
  assign n44107 = \P2_P3_PhyAddrPointer_reg[18]/NET0131  & ~n36826 ;
  assign n44108 = ~n38603 & ~n44107 ;
  assign n44109 = ~n44106 & n44108 ;
  assign n44110 = n27308 & ~n44109 ;
  assign n44114 = ~\P2_P3_PhyAddrPointer_reg[18]/NET0131  & ~n44095 ;
  assign n44115 = ~n42114 & ~n44114 ;
  assign n44116 = ~n36831 & n44115 ;
  assign n44111 = ~\P2_P3_PhyAddrPointer_reg[18]/NET0131  & ~n42106 ;
  assign n44112 = n27325 & ~n42107 ;
  assign n44113 = ~n44111 & n44112 ;
  assign n44103 = \P2_P3_PhyAddrPointer_reg[18]/NET0131  & ~n36873 ;
  assign n44117 = ~n38585 & ~n44103 ;
  assign n44118 = ~n44113 & n44117 ;
  assign n44119 = ~n44116 & n44118 ;
  assign n44120 = ~n44110 & n44119 ;
  assign n44122 = \P2_P3_PhyAddrPointer_reg[21]/NET0131  & ~n27283 ;
  assign n44123 = ~n38661 & ~n44122 ;
  assign n44124 = n27117 & ~n44123 ;
  assign n44125 = \P2_P3_PhyAddrPointer_reg[21]/NET0131  & ~n36826 ;
  assign n44126 = ~n38666 & ~n44125 ;
  assign n44127 = ~n44124 & n44126 ;
  assign n44128 = n27308 & ~n44127 ;
  assign n44129 = ~\P2_P3_PhyAddrPointer_reg[21]/NET0131  & ~n39873 ;
  assign n44130 = ~n39870 & ~n44129 ;
  assign n44131 = ~n36831 & n44130 ;
  assign n44132 = ~\P2_P3_PhyAddrPointer_reg[21]/NET0131  & ~n36852 ;
  assign n44133 = n42140 & ~n44132 ;
  assign n44121 = \P2_P3_PhyAddrPointer_reg[21]/NET0131  & ~n36873 ;
  assign n44134 = ~n38649 & ~n44121 ;
  assign n44135 = ~n44133 & n44134 ;
  assign n44136 = ~n44131 & n44135 ;
  assign n44137 = ~n44128 & n44136 ;
  assign n44139 = \P2_P3_PhyAddrPointer_reg[25]/NET0131  & ~n27283 ;
  assign n44140 = ~n38689 & ~n44139 ;
  assign n44141 = n27117 & ~n44140 ;
  assign n44142 = \P2_P3_PhyAddrPointer_reg[25]/NET0131  & ~n36826 ;
  assign n44143 = ~n38694 & ~n44142 ;
  assign n44144 = ~n44141 & n44143 ;
  assign n44145 = n27308 & ~n44144 ;
  assign n44149 = ~\P2_P3_PhyAddrPointer_reg[25]/NET0131  & ~n42160 ;
  assign n44150 = ~n42190 & ~n44149 ;
  assign n44151 = ~n36831 & n44150 ;
  assign n44146 = ~\P2_P3_PhyAddrPointer_reg[25]/NET0131  & ~n36853 ;
  assign n44147 = n27325 & ~n36854 ;
  assign n44148 = ~n44146 & n44147 ;
  assign n44138 = \P2_P3_PhyAddrPointer_reg[25]/NET0131  & ~n36873 ;
  assign n44152 = ~n38679 & ~n44138 ;
  assign n44153 = ~n44148 & n44152 ;
  assign n44154 = ~n44151 & n44153 ;
  assign n44155 = ~n44145 & n44154 ;
  assign n44161 = \P2_P3_PhyAddrPointer_reg[8]/NET0131  & ~n27283 ;
  assign n44162 = ~n40500 & ~n44161 ;
  assign n44163 = n27117 & ~n44162 ;
  assign n44164 = \P2_P3_PhyAddrPointer_reg[8]/NET0131  & ~n36826 ;
  assign n44165 = ~n40505 & ~n44164 ;
  assign n44166 = ~n44163 & n44165 ;
  assign n44167 = n27308 & ~n44166 ;
  assign n44168 = n36839 & ~n39862 ;
  assign n44170 = \P2_P3_PhyAddrPointer_reg[8]/NET0131  & n44168 ;
  assign n44169 = ~\P2_P3_PhyAddrPointer_reg[8]/NET0131  & ~n44168 ;
  assign n44171 = n27315 & ~n44169 ;
  assign n44172 = ~n44170 & n44171 ;
  assign n44156 = \P2_P3_PhyAddrPointer_reg[1]/NET0131  & n36838 ;
  assign n44157 = \P2_P3_PhyAddrPointer_reg[7]/NET0131  & n44156 ;
  assign n44158 = ~\P2_P3_PhyAddrPointer_reg[8]/NET0131  & ~n44157 ;
  assign n44159 = ~n39838 & ~n44158 ;
  assign n44160 = n32867 & n44159 ;
  assign n44173 = \P2_P3_PhyAddrPointer_reg[8]/NET0131  & ~n36873 ;
  assign n44174 = ~n40490 & ~n44173 ;
  assign n44175 = ~n44160 & n44174 ;
  assign n44176 = ~n44172 & n44175 ;
  assign n44177 = ~n44167 & n44176 ;
  assign n44193 = ~n25830 & n30927 ;
  assign n44182 = ~n25743 & ~n31336 ;
  assign n44183 = n35131 & ~n44182 ;
  assign n44184 = \P1_P2_InstAddrPointer_reg[4]/NET0131  & ~n44183 ;
  assign n44180 = n25887 & n31384 ;
  assign n44196 = ~n31385 & n31404 ;
  assign n44194 = ~n31385 & ~n31386 ;
  assign n44195 = n31403 & ~n44194 ;
  assign n44197 = n25881 & ~n44195 ;
  assign n44198 = ~n44196 & n44197 ;
  assign n44199 = ~n44180 & ~n44198 ;
  assign n44200 = ~n44184 & n44199 ;
  assign n44201 = ~n44193 & n44200 ;
  assign n44181 = ~n25817 & n31223 ;
  assign n44185 = \P1_P2_InstAddrPointer_reg[4]/NET0131  & n25733 ;
  assign n44188 = ~n30959 & n31102 ;
  assign n44186 = ~n30959 & ~n30960 ;
  assign n44187 = n31101 & ~n44186 ;
  assign n44189 = ~n25733 & ~n44187 ;
  assign n44190 = ~n44188 & n44189 ;
  assign n44191 = ~n44185 & ~n44190 ;
  assign n44192 = n25701 & ~n44191 ;
  assign n44202 = ~n44181 & ~n44192 ;
  assign n44203 = n44201 & n44202 ;
  assign n44204 = n25918 & ~n44203 ;
  assign n44178 = \P1_P2_rEIP_reg[4]/NET0131  & n27967 ;
  assign n44179 = \P1_P2_InstAddrPointer_reg[4]/NET0131  & ~n31487 ;
  assign n44205 = ~n44178 & ~n44179 ;
  assign n44206 = ~n44204 & n44205 ;
  assign n44210 = \P1_P2_InstAddrPointer_reg[6]/NET0131  & n25733 ;
  assign n44213 = ~n30889 & n31106 ;
  assign n44211 = ~n30889 & ~n30890 ;
  assign n44212 = n31105 & ~n44211 ;
  assign n44214 = ~n25733 & ~n44212 ;
  assign n44215 = ~n44213 & n44214 ;
  assign n44216 = ~n44210 & ~n44215 ;
  assign n44217 = n25701 & ~n44216 ;
  assign n44223 = ~n31377 & n31408 ;
  assign n44221 = ~n31377 & ~n31378 ;
  assign n44222 = n31407 & ~n44221 ;
  assign n44224 = n25881 & ~n44222 ;
  assign n44225 = ~n44223 & n44224 ;
  assign n44218 = ~n25817 & n31215 ;
  assign n44219 = ~n25830 & n30857 ;
  assign n44209 = n25887 & n31376 ;
  assign n44220 = \P1_P2_InstAddrPointer_reg[6]/NET0131  & ~n35131 ;
  assign n44226 = ~n44209 & ~n44220 ;
  assign n44227 = ~n44219 & n44226 ;
  assign n44228 = ~n44218 & n44227 ;
  assign n44229 = ~n44225 & n44228 ;
  assign n44230 = ~n44217 & n44229 ;
  assign n44231 = n25918 & ~n44230 ;
  assign n44207 = \P1_P2_rEIP_reg[6]/NET0131  & n27967 ;
  assign n44208 = \P1_P2_InstAddrPointer_reg[6]/NET0131  & ~n31487 ;
  assign n44232 = ~n44207 & ~n44208 ;
  assign n44233 = ~n44231 & n44232 ;
  assign n44240 = \P2_P1_InstAddrPointer_reg[4]/NET0131  & n25947 ;
  assign n44243 = ~n31650 & n31793 ;
  assign n44241 = ~n31650 & ~n31651 ;
  assign n44242 = n31792 & ~n44241 ;
  assign n44244 = ~n25947 & ~n44242 ;
  assign n44245 = ~n44243 & n44244 ;
  assign n44246 = ~n44240 & ~n44245 ;
  assign n44247 = n25945 & ~n44246 ;
  assign n44236 = n31618 & ~n32159 ;
  assign n44238 = \P2_P1_InstAddrPointer_reg[4]/NET0131  & ~n35385 ;
  assign n44239 = n26068 & n32073 ;
  assign n44253 = ~n44238 & ~n44239 ;
  assign n44254 = ~n44236 & n44253 ;
  assign n44237 = ~n25995 & n31905 ;
  assign n44248 = ~n32074 & ~n32075 ;
  assign n44250 = ~n32092 & n44248 ;
  assign n44249 = n32092 & ~n44248 ;
  assign n44251 = n25964 & ~n44249 ;
  assign n44252 = ~n44250 & n44251 ;
  assign n44255 = ~n44237 & ~n44252 ;
  assign n44256 = n44254 & n44255 ;
  assign n44257 = ~n44247 & n44256 ;
  assign n44258 = n11623 & ~n44257 ;
  assign n44234 = \P2_P1_rEIP_reg[4]/NET0131  & n11616 ;
  assign n44235 = \P2_P1_InstAddrPointer_reg[4]/NET0131  & ~n32172 ;
  assign n44259 = ~n44234 & ~n44235 ;
  assign n44260 = ~n44258 & n44259 ;
  assign n44264 = \P2_P1_InstAddrPointer_reg[6]/NET0131  & n25947 ;
  assign n44267 = ~n31580 & n31797 ;
  assign n44265 = ~n31580 & ~n31581 ;
  assign n44266 = ~n31796 & ~n44265 ;
  assign n44268 = ~n25947 & ~n44266 ;
  assign n44269 = ~n44267 & n44268 ;
  assign n44270 = ~n44264 & ~n44269 ;
  assign n44271 = n25945 & ~n44270 ;
  assign n44275 = ~n32066 & ~n32067 ;
  assign n44277 = ~n32096 & n44275 ;
  assign n44276 = n32096 & ~n44275 ;
  assign n44278 = n25964 & ~n44276 ;
  assign n44279 = ~n44277 & n44278 ;
  assign n44273 = n31548 & ~n32159 ;
  assign n44272 = ~n25995 & n31896 ;
  assign n44263 = n26068 & n32065 ;
  assign n44274 = \P2_P1_InstAddrPointer_reg[6]/NET0131  & ~n35385 ;
  assign n44280 = ~n44263 & ~n44274 ;
  assign n44281 = ~n44272 & n44280 ;
  assign n44282 = ~n44273 & n44281 ;
  assign n44283 = ~n44279 & n44282 ;
  assign n44284 = ~n44271 & n44283 ;
  assign n44285 = n11623 & ~n44284 ;
  assign n44261 = \P2_P1_rEIP_reg[6]/NET0131  & n11616 ;
  assign n44262 = \P2_P1_InstAddrPointer_reg[6]/NET0131  & ~n32172 ;
  assign n44286 = ~n44261 & ~n44262 ;
  assign n44287 = ~n44285 & n44286 ;
  assign n44300 = ~n26688 & n32618 ;
  assign n44292 = \P2_P2_InstAddrPointer_reg[4]/NET0131  & n26629 ;
  assign n44295 = ~n32330 & n32473 ;
  assign n44293 = ~n32330 & ~n32331 ;
  assign n44294 = n32472 & ~n44293 ;
  assign n44296 = ~n26629 & ~n44294 ;
  assign n44297 = ~n44295 & n44296 ;
  assign n44298 = ~n44292 & ~n44297 ;
  assign n44299 = n26621 & ~n44298 ;
  assign n44290 = \P2_P2_InstAddrPointer_reg[4]/NET0131  & ~n35424 ;
  assign n44291 = n26757 & n32779 ;
  assign n44307 = ~n44290 & ~n44291 ;
  assign n44301 = ~n26764 & n32298 ;
  assign n44304 = ~n32780 & n32796 ;
  assign n44302 = ~n32780 & ~n32781 ;
  assign n44303 = ~n32795 & ~n44302 ;
  assign n44305 = n26744 & ~n44303 ;
  assign n44306 = ~n44304 & n44305 ;
  assign n44308 = ~n44301 & ~n44306 ;
  assign n44309 = n44307 & n44308 ;
  assign n44310 = ~n44299 & n44309 ;
  assign n44311 = ~n44300 & n44310 ;
  assign n44312 = n26792 & ~n44311 ;
  assign n44288 = \P2_P2_rEIP_reg[4]/NET0131  & n28046 ;
  assign n44289 = \P2_P2_InstAddrPointer_reg[4]/NET0131  & ~n32860 ;
  assign n44313 = ~n44288 & ~n44289 ;
  assign n44314 = ~n44312 & n44313 ;
  assign n44319 = \P2_P2_InstAddrPointer_reg[6]/NET0131  & n26629 ;
  assign n44325 = ~n32260 & ~n32261 ;
  assign n44327 = n32476 & n44325 ;
  assign n44326 = ~n32476 & ~n44325 ;
  assign n44328 = n32510 & ~n44326 ;
  assign n44329 = ~n44327 & n44328 ;
  assign n44320 = ~n32595 & ~n32596 ;
  assign n44322 = ~n32626 & n44320 ;
  assign n44321 = n32626 & ~n44320 ;
  assign n44323 = ~n32510 & ~n44321 ;
  assign n44324 = ~n44322 & n44323 ;
  assign n44330 = ~n26629 & ~n44324 ;
  assign n44331 = ~n44329 & n44330 ;
  assign n44332 = ~n44319 & ~n44331 ;
  assign n44333 = n26621 & ~n44332 ;
  assign n44338 = ~n32772 & n32800 ;
  assign n44336 = ~n32772 & ~n32773 ;
  assign n44337 = n32799 & ~n44336 ;
  assign n44339 = n26744 & ~n44337 ;
  assign n44340 = ~n44338 & n44339 ;
  assign n44317 = ~n26688 & n32594 ;
  assign n44335 = \P2_P2_InstAddrPointer_reg[6]/NET0131  & ~n35424 ;
  assign n44318 = ~n26764 & n32228 ;
  assign n44334 = n26757 & n32771 ;
  assign n44341 = ~n44318 & ~n44334 ;
  assign n44342 = ~n44335 & n44341 ;
  assign n44343 = ~n44317 & n44342 ;
  assign n44344 = ~n44340 & n44343 ;
  assign n44345 = ~n44333 & n44344 ;
  assign n44346 = n26792 & ~n44345 ;
  assign n44315 = \P2_P2_rEIP_reg[6]/NET0131  & n28046 ;
  assign n44316 = \P2_P2_InstAddrPointer_reg[6]/NET0131  & ~n32860 ;
  assign n44347 = ~n44315 & ~n44316 ;
  assign n44348 = ~n44346 & n44347 ;
  assign n44357 = \P2_P3_InstAddrPointer_reg[4]/NET0131  & ~n27283 ;
  assign n44363 = ~n33304 & ~n33305 ;
  assign n44365 = ~n33319 & n44363 ;
  assign n44364 = n33319 & ~n44363 ;
  assign n44366 = ~n33242 & ~n44364 ;
  assign n44367 = ~n44365 & n44366 ;
  assign n44358 = ~n33061 & ~n33062 ;
  assign n44360 = n33203 & n44358 ;
  assign n44359 = ~n33203 & ~n44358 ;
  assign n44361 = n33242 & ~n44359 ;
  assign n44362 = ~n44360 & n44361 ;
  assign n44368 = n27283 & ~n44362 ;
  assign n44369 = ~n44367 & n44368 ;
  assign n44370 = ~n44357 & ~n44369 ;
  assign n44371 = n27117 & ~n44370 ;
  assign n44374 = ~n33446 & n33465 ;
  assign n44372 = ~n33446 & ~n33447 ;
  assign n44373 = n33464 & ~n44372 ;
  assign n44375 = n27280 & ~n44373 ;
  assign n44376 = ~n44374 & n44375 ;
  assign n44354 = n27219 & n33445 ;
  assign n44356 = ~n27142 & n33303 ;
  assign n44377 = ~n44354 & ~n44356 ;
  assign n44378 = ~n44376 & n44377 ;
  assign n44351 = ~n27111 & ~n32874 ;
  assign n44352 = n34355 & ~n44351 ;
  assign n44353 = \P2_P3_InstAddrPointer_reg[4]/NET0131  & ~n44352 ;
  assign n44355 = ~n27229 & n33029 ;
  assign n44379 = ~n44353 & ~n44355 ;
  assign n44380 = n44378 & n44379 ;
  assign n44381 = ~n44371 & n44380 ;
  assign n44382 = n27308 & ~n44381 ;
  assign n44349 = \P2_P3_rEIP_reg[4]/NET0131  & n32864 ;
  assign n44350 = \P2_P3_InstAddrPointer_reg[4]/NET0131  & ~n32870 ;
  assign n44383 = ~n44349 & ~n44350 ;
  assign n44384 = ~n44382 & n44383 ;
  assign n44386 = \P2_P3_InstAddrPointer_reg[6]/NET0131  & ~n27283 ;
  assign n44389 = ~n32991 & n33208 ;
  assign n44387 = ~n32991 & ~n32992 ;
  assign n44388 = n33207 & ~n44387 ;
  assign n44390 = n27283 & ~n44388 ;
  assign n44391 = ~n44389 & n44390 ;
  assign n44392 = ~n44386 & ~n44391 ;
  assign n44393 = n27117 & ~n44392 ;
  assign n44400 = ~n33438 & n33469 ;
  assign n44398 = ~n33438 & ~n33439 ;
  assign n44399 = n33468 & ~n44398 ;
  assign n44401 = n27280 & ~n44399 ;
  assign n44402 = ~n44400 & n44401 ;
  assign n44394 = ~n27229 & n32959 ;
  assign n44397 = ~n27142 & n33292 ;
  assign n44395 = \P2_P3_InstAddrPointer_reg[6]/NET0131  & ~n34355 ;
  assign n44396 = n27219 & n33437 ;
  assign n44403 = ~n44395 & ~n44396 ;
  assign n44404 = ~n44397 & n44403 ;
  assign n44405 = ~n44394 & n44404 ;
  assign n44406 = ~n44402 & n44405 ;
  assign n44407 = ~n44393 & n44406 ;
  assign n44408 = n27308 & ~n44407 ;
  assign n44385 = \P2_P3_rEIP_reg[6]/NET0131  & n32864 ;
  assign n44409 = \P2_P3_InstAddrPointer_reg[6]/NET0131  & ~n32870 ;
  assign n44410 = ~n44385 & ~n44409 ;
  assign n44411 = ~n44408 & n44410 ;
  assign n44423 = \P1_P1_InstAddrPointer_reg[4]/NET0131  & n26249 ;
  assign n44429 = ~n33918 & ~n33919 ;
  assign n44431 = ~n33933 & n44429 ;
  assign n44430 = n33933 & ~n44429 ;
  assign n44432 = ~n29558 & ~n44430 ;
  assign n44433 = ~n44431 & n44432 ;
  assign n44424 = ~n33662 & ~n33663 ;
  assign n44426 = n33804 & n44424 ;
  assign n44425 = ~n33804 & ~n44424 ;
  assign n44427 = n29558 & ~n44425 ;
  assign n44428 = ~n44426 & n44427 ;
  assign n44434 = ~n26249 & ~n44428 ;
  assign n44435 = ~n44433 & n44434 ;
  assign n44436 = ~n44423 & ~n44435 ;
  assign n44437 = n26126 & ~n44436 ;
  assign n44415 = ~n26189 & n33630 ;
  assign n44422 = ~n26151 & n33917 ;
  assign n44419 = ~n34069 & n34088 ;
  assign n44417 = ~n34069 & ~n34070 ;
  assign n44418 = n34087 & ~n44417 ;
  assign n44420 = n26263 & ~n44418 ;
  assign n44421 = ~n44419 & n44420 ;
  assign n44414 = \P1_P1_InstAddrPointer_reg[4]/NET0131  & ~n35760 ;
  assign n44416 = n26192 & n34068 ;
  assign n44438 = ~n44414 & ~n44416 ;
  assign n44439 = ~n44421 & n44438 ;
  assign n44440 = ~n44422 & n44439 ;
  assign n44441 = ~n44415 & n44440 ;
  assign n44442 = ~n44437 & n44441 ;
  assign n44443 = n8355 & ~n44442 ;
  assign n44412 = \P1_P1_rEIP_reg[4]/NET0131  & n8357 ;
  assign n44413 = \P1_P1_InstAddrPointer_reg[4]/NET0131  & ~n34164 ;
  assign n44444 = ~n44412 & ~n44413 ;
  assign n44445 = ~n44443 & n44444 ;
  assign n44448 = \P1_P1_InstAddrPointer_reg[6]/NET0131  & n26249 ;
  assign n44454 = ~n33910 & ~n33911 ;
  assign n44456 = ~n33937 & n44454 ;
  assign n44455 = n33937 & ~n44454 ;
  assign n44457 = ~n29558 & ~n44455 ;
  assign n44458 = ~n44456 & n44457 ;
  assign n44449 = ~n33592 & ~n33593 ;
  assign n44451 = n33808 & n44449 ;
  assign n44450 = ~n33808 & ~n44449 ;
  assign n44452 = n29558 & ~n44450 ;
  assign n44453 = ~n44451 & n44452 ;
  assign n44459 = ~n26249 & ~n44453 ;
  assign n44460 = ~n44458 & n44459 ;
  assign n44461 = ~n44448 & ~n44460 ;
  assign n44462 = n26126 & ~n44461 ;
  assign n44465 = ~n34061 & n34092 ;
  assign n44463 = ~n34061 & ~n34062 ;
  assign n44464 = n34091 & ~n44463 ;
  assign n44466 = n26263 & ~n44464 ;
  assign n44467 = ~n44465 & n44466 ;
  assign n44470 = ~n26189 & n33560 ;
  assign n44447 = ~n26151 & n33909 ;
  assign n44468 = n26192 & n34060 ;
  assign n44469 = \P1_P1_InstAddrPointer_reg[6]/NET0131  & ~n35760 ;
  assign n44471 = ~n44468 & ~n44469 ;
  assign n44472 = ~n44447 & n44471 ;
  assign n44473 = ~n44470 & n44472 ;
  assign n44474 = ~n44467 & n44473 ;
  assign n44475 = ~n44462 & n44474 ;
  assign n44476 = n8355 & ~n44475 ;
  assign n44446 = \P1_P1_rEIP_reg[6]/NET0131  & n8357 ;
  assign n44477 = \P1_P1_InstAddrPointer_reg[6]/NET0131  & ~n34164 ;
  assign n44478 = ~n44446 & ~n44477 ;
  assign n44479 = ~n44476 & n44478 ;
  assign n44480 = \P2_P1_lWord_reg[4]/NET0131  & ~n34408 ;
  assign n44481 = \P2_P1_EAX_reg[4]/NET0131  & n24899 ;
  assign n44482 = n21062 & n24887 ;
  assign n44483 = ~n44481 & ~n44482 ;
  assign n44484 = n11623 & ~n44483 ;
  assign n44485 = ~n44480 & ~n44484 ;
  assign n44486 = \P2_P1_uWord_reg[5]/NET0131  & ~n24913 ;
  assign n44487 = \P2_P1_uWord_reg[5]/NET0131  & n34405 ;
  assign n44488 = \P2_P1_uWord_reg[5]/NET0131  & ~n22337 ;
  assign n44489 = ~n24249 & ~n44488 ;
  assign n44490 = n21062 & ~n44489 ;
  assign n44491 = ~\P2_P1_EAX_reg[21]/NET0131  & ~n27392 ;
  assign n44492 = ~n27393 & ~n44491 ;
  assign n44493 = n24899 & n44492 ;
  assign n44494 = ~n44490 & ~n44493 ;
  assign n44495 = ~n44487 & n44494 ;
  assign n44496 = n11623 & ~n44495 ;
  assign n44497 = ~n44486 & ~n44496 ;
  assign n44498 = \P2_P1_uWord_reg[6]/NET0131  & ~n24913 ;
  assign n44499 = \P2_P1_uWord_reg[6]/NET0131  & ~n34406 ;
  assign n44500 = ~\P2_P1_EAX_reg[22]/NET0131  & ~n27393 ;
  assign n44501 = ~n27394 & ~n44500 ;
  assign n44502 = n24899 & n44501 ;
  assign n44503 = ~n37886 & ~n44502 ;
  assign n44504 = ~n44499 & n44503 ;
  assign n44505 = n11623 & ~n44504 ;
  assign n44506 = ~n44498 & ~n44505 ;
  assign n44507 = ~n27612 & ~n27615 ;
  assign n44508 = n43242 & n44507 ;
  assign n44509 = \P2_P2_EAX_reg[27]/NET0131  & ~n44508 ;
  assign n44705 = \P2_P2_EAX_reg[0]/NET0131  & \P2_P2_EAX_reg[1]/NET0131  ;
  assign n44706 = \P2_P2_EAX_reg[2]/NET0131  & n44705 ;
  assign n44707 = \P2_P2_EAX_reg[3]/NET0131  & n44706 ;
  assign n44708 = \P2_P2_EAX_reg[4]/NET0131  & n44707 ;
  assign n44709 = \P2_P2_EAX_reg[5]/NET0131  & n44708 ;
  assign n44710 = \P2_P2_EAX_reg[6]/NET0131  & n44709 ;
  assign n44711 = \P2_P2_EAX_reg[7]/NET0131  & n44710 ;
  assign n44712 = \P2_P2_EAX_reg[8]/NET0131  & n44711 ;
  assign n44713 = \P2_P2_EAX_reg[9]/NET0131  & n44712 ;
  assign n44714 = \P2_P2_EAX_reg[10]/NET0131  & n44713 ;
  assign n44715 = \P2_P2_EAX_reg[11]/NET0131  & n44714 ;
  assign n44716 = \P2_P2_EAX_reg[12]/NET0131  & n44715 ;
  assign n44717 = \P2_P2_EAX_reg[13]/NET0131  & n44716 ;
  assign n44718 = \P2_P2_EAX_reg[14]/NET0131  & n44717 ;
  assign n44719 = \P2_P2_EAX_reg[15]/NET0131  & n44718 ;
  assign n44720 = \P2_P2_EAX_reg[16]/NET0131  & n44719 ;
  assign n44721 = \P2_P2_EAX_reg[17]/NET0131  & n44720 ;
  assign n44722 = \P2_P2_EAX_reg[18]/NET0131  & n44721 ;
  assign n44723 = \P2_P2_EAX_reg[19]/NET0131  & n44722 ;
  assign n44724 = \P2_P2_EAX_reg[20]/NET0131  & n44723 ;
  assign n44725 = \P2_P2_EAX_reg[21]/NET0131  & n44724 ;
  assign n44726 = \P2_P2_EAX_reg[22]/NET0131  & n44725 ;
  assign n44727 = \P2_P2_EAX_reg[23]/NET0131  & n44726 ;
  assign n44728 = \P2_P2_EAX_reg[24]/NET0131  & n44727 ;
  assign n44729 = \P2_P2_EAX_reg[25]/NET0131  & n44728 ;
  assign n44730 = \P2_P2_EAX_reg[26]/NET0131  & n44729 ;
  assign n44731 = \P2_P2_EAX_reg[27]/NET0131  & n44730 ;
  assign n44732 = n26660 & n26669 ;
  assign n44733 = ~n44731 & n44732 ;
  assign n44510 = n26582 & n26611 ;
  assign n44734 = n26639 & ~n44732 ;
  assign n44735 = ~n26582 & ~n44734 ;
  assign n44736 = ~n44510 & ~n44735 ;
  assign n44737 = ~n44733 & ~n44736 ;
  assign n44738 = \P2_P2_EAX_reg[27]/NET0131  & ~n44737 ;
  assign n44739 = n44730 & n44733 ;
  assign n44522 = \P2_P2_InstQueue_reg[1][7]/NET0131  & n26330 ;
  assign n44520 = \P2_P2_InstQueue_reg[2][7]/NET0131  & n26325 ;
  assign n44511 = \P2_P2_InstQueue_reg[9][7]/NET0131  & n26300 ;
  assign n44512 = \P2_P2_InstQueue_reg[0][7]/NET0131  & n26336 ;
  assign n44527 = ~n44511 & ~n44512 ;
  assign n44537 = ~n44520 & n44527 ;
  assign n44538 = ~n44522 & n44537 ;
  assign n44523 = \P2_P2_InstQueue_reg[8][7]/NET0131  & n26318 ;
  assign n44524 = \P2_P2_InstQueue_reg[11][7]/NET0131  & n26334 ;
  assign n44532 = ~n44523 & ~n44524 ;
  assign n44525 = \P2_P2_InstQueue_reg[4][7]/NET0131  & n26338 ;
  assign n44526 = \P2_P2_InstQueue_reg[3][7]/NET0131  & n26322 ;
  assign n44533 = ~n44525 & ~n44526 ;
  assign n44534 = n44532 & n44533 ;
  assign n44517 = \P2_P2_InstQueue_reg[15][7]/NET0131  & n26313 ;
  assign n44518 = \P2_P2_InstQueue_reg[13][7]/NET0131  & n26320 ;
  assign n44530 = ~n44517 & ~n44518 ;
  assign n44519 = \P2_P2_InstQueue_reg[7][7]/NET0131  & n26307 ;
  assign n44521 = \P2_P2_InstQueue_reg[10][7]/NET0131  & n26327 ;
  assign n44531 = ~n44519 & ~n44521 ;
  assign n44535 = n44530 & n44531 ;
  assign n44513 = \P2_P2_InstQueue_reg[5][7]/NET0131  & n26316 ;
  assign n44514 = \P2_P2_InstQueue_reg[6][7]/NET0131  & n26332 ;
  assign n44528 = ~n44513 & ~n44514 ;
  assign n44515 = \P2_P2_InstQueue_reg[14][7]/NET0131  & n26310 ;
  assign n44516 = \P2_P2_InstQueue_reg[12][7]/NET0131  & n26304 ;
  assign n44529 = ~n44515 & ~n44516 ;
  assign n44536 = n44528 & n44529 ;
  assign n44539 = n44535 & n44536 ;
  assign n44540 = n44534 & n44539 ;
  assign n44541 = n44538 & n44540 ;
  assign n44553 = \P2_P2_InstQueue_reg[2][0]/NET0131  & n26330 ;
  assign n44551 = \P2_P2_InstQueue_reg[3][0]/NET0131  & n26325 ;
  assign n44542 = \P2_P2_InstQueue_reg[10][0]/NET0131  & n26300 ;
  assign n44543 = \P2_P2_InstQueue_reg[13][0]/NET0131  & n26304 ;
  assign n44558 = ~n44542 & ~n44543 ;
  assign n44568 = ~n44551 & n44558 ;
  assign n44569 = ~n44553 & n44568 ;
  assign n44554 = \P2_P2_InstQueue_reg[9][0]/NET0131  & n26318 ;
  assign n44555 = \P2_P2_InstQueue_reg[4][0]/NET0131  & n26322 ;
  assign n44563 = ~n44554 & ~n44555 ;
  assign n44556 = \P2_P2_InstQueue_reg[6][0]/NET0131  & n26316 ;
  assign n44557 = \P2_P2_InstQueue_reg[15][0]/NET0131  & n26310 ;
  assign n44564 = ~n44556 & ~n44557 ;
  assign n44565 = n44563 & n44564 ;
  assign n44548 = \P2_P2_InstQueue_reg[8][0]/NET0131  & n26307 ;
  assign n44549 = \P2_P2_InstQueue_reg[1][0]/NET0131  & n26336 ;
  assign n44561 = ~n44548 & ~n44549 ;
  assign n44550 = \P2_P2_InstQueue_reg[7][0]/NET0131  & n26332 ;
  assign n44552 = \P2_P2_InstQueue_reg[11][0]/NET0131  & n26327 ;
  assign n44562 = ~n44550 & ~n44552 ;
  assign n44566 = n44561 & n44562 ;
  assign n44544 = \P2_P2_InstQueue_reg[14][0]/NET0131  & n26320 ;
  assign n44545 = \P2_P2_InstQueue_reg[12][0]/NET0131  & n26334 ;
  assign n44559 = ~n44544 & ~n44545 ;
  assign n44546 = \P2_P2_InstQueue_reg[5][0]/NET0131  & n26338 ;
  assign n44547 = \P2_P2_InstQueue_reg[0][0]/NET0131  & n26313 ;
  assign n44560 = ~n44546 & ~n44547 ;
  assign n44567 = n44559 & n44560 ;
  assign n44570 = n44566 & n44567 ;
  assign n44571 = n44565 & n44570 ;
  assign n44572 = n44569 & n44571 ;
  assign n44573 = ~n44541 & ~n44572 ;
  assign n44585 = \P2_P2_InstQueue_reg[2][1]/NET0131  & n26330 ;
  assign n44583 = \P2_P2_InstQueue_reg[3][1]/NET0131  & n26325 ;
  assign n44574 = \P2_P2_InstQueue_reg[10][1]/NET0131  & n26300 ;
  assign n44575 = \P2_P2_InstQueue_reg[13][1]/NET0131  & n26304 ;
  assign n44590 = ~n44574 & ~n44575 ;
  assign n44600 = ~n44583 & n44590 ;
  assign n44601 = ~n44585 & n44600 ;
  assign n44586 = \P2_P2_InstQueue_reg[9][1]/NET0131  & n26318 ;
  assign n44587 = \P2_P2_InstQueue_reg[4][1]/NET0131  & n26322 ;
  assign n44595 = ~n44586 & ~n44587 ;
  assign n44588 = \P2_P2_InstQueue_reg[6][1]/NET0131  & n26316 ;
  assign n44589 = \P2_P2_InstQueue_reg[15][1]/NET0131  & n26310 ;
  assign n44596 = ~n44588 & ~n44589 ;
  assign n44597 = n44595 & n44596 ;
  assign n44580 = \P2_P2_InstQueue_reg[8][1]/NET0131  & n26307 ;
  assign n44581 = \P2_P2_InstQueue_reg[1][1]/NET0131  & n26336 ;
  assign n44593 = ~n44580 & ~n44581 ;
  assign n44582 = \P2_P2_InstQueue_reg[7][1]/NET0131  & n26332 ;
  assign n44584 = \P2_P2_InstQueue_reg[11][1]/NET0131  & n26327 ;
  assign n44594 = ~n44582 & ~n44584 ;
  assign n44598 = n44593 & n44594 ;
  assign n44576 = \P2_P2_InstQueue_reg[14][1]/NET0131  & n26320 ;
  assign n44577 = \P2_P2_InstQueue_reg[12][1]/NET0131  & n26334 ;
  assign n44591 = ~n44576 & ~n44577 ;
  assign n44578 = \P2_P2_InstQueue_reg[5][1]/NET0131  & n26338 ;
  assign n44579 = \P2_P2_InstQueue_reg[0][1]/NET0131  & n26313 ;
  assign n44592 = ~n44578 & ~n44579 ;
  assign n44599 = n44591 & n44592 ;
  assign n44602 = n44598 & n44599 ;
  assign n44603 = n44597 & n44602 ;
  assign n44604 = n44601 & n44603 ;
  assign n44605 = n44573 & ~n44604 ;
  assign n44617 = \P2_P2_InstQueue_reg[2][2]/NET0131  & n26330 ;
  assign n44615 = \P2_P2_InstQueue_reg[3][2]/NET0131  & n26325 ;
  assign n44606 = \P2_P2_InstQueue_reg[10][2]/NET0131  & n26300 ;
  assign n44607 = \P2_P2_InstQueue_reg[9][2]/NET0131  & n26318 ;
  assign n44622 = ~n44606 & ~n44607 ;
  assign n44632 = ~n44615 & n44622 ;
  assign n44633 = ~n44617 & n44632 ;
  assign n44618 = \P2_P2_InstQueue_reg[5][2]/NET0131  & n26338 ;
  assign n44619 = \P2_P2_InstQueue_reg[4][2]/NET0131  & n26322 ;
  assign n44627 = ~n44618 & ~n44619 ;
  assign n44620 = \P2_P2_InstQueue_reg[6][2]/NET0131  & n26316 ;
  assign n44621 = \P2_P2_InstQueue_reg[1][2]/NET0131  & n26336 ;
  assign n44628 = ~n44620 & ~n44621 ;
  assign n44629 = n44627 & n44628 ;
  assign n44612 = \P2_P2_InstQueue_reg[0][2]/NET0131  & n26313 ;
  assign n44613 = \P2_P2_InstQueue_reg[14][2]/NET0131  & n26320 ;
  assign n44625 = ~n44612 & ~n44613 ;
  assign n44614 = \P2_P2_InstQueue_reg[12][2]/NET0131  & n26334 ;
  assign n44616 = \P2_P2_InstQueue_reg[11][2]/NET0131  & n26327 ;
  assign n44626 = ~n44614 & ~n44616 ;
  assign n44630 = n44625 & n44626 ;
  assign n44608 = \P2_P2_InstQueue_reg[15][2]/NET0131  & n26310 ;
  assign n44609 = \P2_P2_InstQueue_reg[7][2]/NET0131  & n26332 ;
  assign n44623 = ~n44608 & ~n44609 ;
  assign n44610 = \P2_P2_InstQueue_reg[13][2]/NET0131  & n26304 ;
  assign n44611 = \P2_P2_InstQueue_reg[8][2]/NET0131  & n26307 ;
  assign n44624 = ~n44610 & ~n44611 ;
  assign n44631 = n44623 & n44624 ;
  assign n44634 = n44630 & n44631 ;
  assign n44635 = n44629 & n44634 ;
  assign n44636 = n44633 & n44635 ;
  assign n44637 = n44605 & ~n44636 ;
  assign n44649 = \P2_P2_InstQueue_reg[2][3]/NET0131  & n26330 ;
  assign n44647 = \P2_P2_InstQueue_reg[3][3]/NET0131  & n26325 ;
  assign n44638 = \P2_P2_InstQueue_reg[10][3]/NET0131  & n26300 ;
  assign n44639 = \P2_P2_InstQueue_reg[9][3]/NET0131  & n26318 ;
  assign n44654 = ~n44638 & ~n44639 ;
  assign n44664 = ~n44647 & n44654 ;
  assign n44665 = ~n44649 & n44664 ;
  assign n44650 = \P2_P2_InstQueue_reg[5][3]/NET0131  & n26338 ;
  assign n44651 = \P2_P2_InstQueue_reg[4][3]/NET0131  & n26322 ;
  assign n44659 = ~n44650 & ~n44651 ;
  assign n44652 = \P2_P2_InstQueue_reg[6][3]/NET0131  & n26316 ;
  assign n44653 = \P2_P2_InstQueue_reg[1][3]/NET0131  & n26336 ;
  assign n44660 = ~n44652 & ~n44653 ;
  assign n44661 = n44659 & n44660 ;
  assign n44644 = \P2_P2_InstQueue_reg[0][3]/NET0131  & n26313 ;
  assign n44645 = \P2_P2_InstQueue_reg[14][3]/NET0131  & n26320 ;
  assign n44657 = ~n44644 & ~n44645 ;
  assign n44646 = \P2_P2_InstQueue_reg[12][3]/NET0131  & n26334 ;
  assign n44648 = \P2_P2_InstQueue_reg[11][3]/NET0131  & n26327 ;
  assign n44658 = ~n44646 & ~n44648 ;
  assign n44662 = n44657 & n44658 ;
  assign n44640 = \P2_P2_InstQueue_reg[15][3]/NET0131  & n26310 ;
  assign n44641 = \P2_P2_InstQueue_reg[7][3]/NET0131  & n26332 ;
  assign n44655 = ~n44640 & ~n44641 ;
  assign n44642 = \P2_P2_InstQueue_reg[13][3]/NET0131  & n26304 ;
  assign n44643 = \P2_P2_InstQueue_reg[8][3]/NET0131  & n26307 ;
  assign n44656 = ~n44642 & ~n44643 ;
  assign n44663 = n44655 & n44656 ;
  assign n44666 = n44662 & n44663 ;
  assign n44667 = n44661 & n44666 ;
  assign n44668 = n44665 & n44667 ;
  assign n44669 = n44637 & ~n44668 ;
  assign n44681 = \P2_P2_InstQueue_reg[2][4]/NET0131  & n26330 ;
  assign n44679 = \P2_P2_InstQueue_reg[3][4]/NET0131  & n26325 ;
  assign n44670 = \P2_P2_InstQueue_reg[10][4]/NET0131  & n26300 ;
  assign n44671 = \P2_P2_InstQueue_reg[13][4]/NET0131  & n26304 ;
  assign n44686 = ~n44670 & ~n44671 ;
  assign n44696 = ~n44679 & n44686 ;
  assign n44697 = ~n44681 & n44696 ;
  assign n44682 = \P2_P2_InstQueue_reg[9][4]/NET0131  & n26318 ;
  assign n44683 = \P2_P2_InstQueue_reg[4][4]/NET0131  & n26322 ;
  assign n44691 = ~n44682 & ~n44683 ;
  assign n44684 = \P2_P2_InstQueue_reg[6][4]/NET0131  & n26316 ;
  assign n44685 = \P2_P2_InstQueue_reg[15][4]/NET0131  & n26310 ;
  assign n44692 = ~n44684 & ~n44685 ;
  assign n44693 = n44691 & n44692 ;
  assign n44676 = \P2_P2_InstQueue_reg[8][4]/NET0131  & n26307 ;
  assign n44677 = \P2_P2_InstQueue_reg[1][4]/NET0131  & n26336 ;
  assign n44689 = ~n44676 & ~n44677 ;
  assign n44678 = \P2_P2_InstQueue_reg[7][4]/NET0131  & n26332 ;
  assign n44680 = \P2_P2_InstQueue_reg[11][4]/NET0131  & n26327 ;
  assign n44690 = ~n44678 & ~n44680 ;
  assign n44694 = n44689 & n44690 ;
  assign n44672 = \P2_P2_InstQueue_reg[14][4]/NET0131  & n26320 ;
  assign n44673 = \P2_P2_InstQueue_reg[12][4]/NET0131  & n26334 ;
  assign n44687 = ~n44672 & ~n44673 ;
  assign n44674 = \P2_P2_InstQueue_reg[5][4]/NET0131  & n26338 ;
  assign n44675 = \P2_P2_InstQueue_reg[0][4]/NET0131  & n26313 ;
  assign n44688 = ~n44674 & ~n44675 ;
  assign n44695 = n44687 & n44688 ;
  assign n44698 = n44694 & n44695 ;
  assign n44699 = n44693 & n44698 ;
  assign n44700 = n44697 & n44699 ;
  assign n44701 = ~n44669 & n44700 ;
  assign n44702 = n44669 & ~n44700 ;
  assign n44703 = ~n44701 & ~n44702 ;
  assign n44704 = n44510 & n44703 ;
  assign n44740 = \P2_P2_EAX_reg[27]/NET0131  & ~n26641 ;
  assign n44741 = ~\P2_buf2_reg[11]/NET0131  & ~n28013 ;
  assign n44742 = ~\P2_buf1_reg[11]/NET0131  & n28013 ;
  assign n44743 = ~n44741 & ~n44742 ;
  assign n44744 = n26641 & n44743 ;
  assign n44745 = ~n44740 & ~n44744 ;
  assign n44746 = n26633 & ~n44745 ;
  assign n44747 = n26641 & ~n29899 ;
  assign n44748 = ~n44740 & ~n44747 ;
  assign n44749 = n26638 & ~n44748 ;
  assign n44750 = ~n44746 & ~n44749 ;
  assign n44751 = ~n44704 & n44750 ;
  assign n44752 = ~n44739 & n44751 ;
  assign n44753 = ~n44738 & n44752 ;
  assign n44754 = n26792 & ~n44753 ;
  assign n44755 = ~n44509 & ~n44754 ;
  assign n44756 = \P1_P1_EAX_reg[4]/NET0131  & n24502 ;
  assign n44757 = ~n7940 & n23946 ;
  assign n44758 = ~n44756 & ~n44757 ;
  assign n44759 = ~n15364 & ~n44758 ;
  assign n44760 = \P1_P1_lWord_reg[4]/NET0131  & ~n24506 ;
  assign n44761 = ~n44759 & ~n44760 ;
  assign n44762 = n8355 & ~n44761 ;
  assign n44763 = \P1_P1_lWord_reg[4]/NET0131  & ~n24515 ;
  assign n44764 = ~n44762 & ~n44763 ;
  assign n44765 = \P1_P1_uWord_reg[5]/NET0131  & ~n24515 ;
  assign n44769 = \P1_P1_uWord_reg[5]/NET0131  & n25363 ;
  assign n44770 = ~n24439 & ~n44769 ;
  assign n44771 = n15334 & ~n44770 ;
  assign n44766 = ~\P1_P1_EAX_reg[21]/NET0131  & ~n25352 ;
  assign n44767 = ~n25353 & ~n44766 ;
  assign n44768 = n24503 & n44767 ;
  assign n44772 = \P1_P1_uWord_reg[5]/NET0131  & n24505 ;
  assign n44773 = ~n44768 & ~n44772 ;
  assign n44774 = ~n44771 & n44773 ;
  assign n44775 = n8355 & ~n44774 ;
  assign n44776 = ~n44765 & ~n44775 ;
  assign n44777 = \P1_P1_uWord_reg[6]/NET0131  & ~n24515 ;
  assign n44781 = \P1_P1_uWord_reg[6]/NET0131  & n25363 ;
  assign n44782 = ~n24167 & ~n44781 ;
  assign n44783 = n15334 & ~n44782 ;
  assign n44778 = ~\P1_P1_EAX_reg[22]/NET0131  & ~n25353 ;
  assign n44779 = n24503 & ~n25354 ;
  assign n44780 = ~n44778 & n44779 ;
  assign n44784 = \P1_P1_uWord_reg[6]/NET0131  & n24505 ;
  assign n44785 = ~n44780 & ~n44784 ;
  assign n44786 = ~n44783 & n44785 ;
  assign n44787 = n8355 & ~n44786 ;
  assign n44788 = ~n44777 & ~n44787 ;
  assign n44792 = ~\P2_P3_EAX_reg[27]/NET0131  & ~n42858 ;
  assign n44793 = n42539 & ~n42859 ;
  assign n44794 = ~n44792 & n44793 ;
  assign n44795 = \P2_P3_EAX_reg[27]/NET0131  & n42542 ;
  assign n44789 = ~n42703 & n42734 ;
  assign n44790 = ~n42735 & ~n44789 ;
  assign n44791 = n42538 & n44790 ;
  assign n44796 = \P2_P3_EAX_reg[27]/NET0131  & ~n27227 ;
  assign n44797 = \P2_buf2_reg[27]/NET0131  & n27227 ;
  assign n44798 = ~n44796 & ~n44797 ;
  assign n44799 = n27186 & ~n44798 ;
  assign n44800 = \P2_buf2_reg[11]/NET0131  & n27227 ;
  assign n44801 = ~n44796 & ~n44800 ;
  assign n44802 = n27122 & ~n44801 ;
  assign n44803 = ~n44799 & ~n44802 ;
  assign n44804 = ~n44791 & n44803 ;
  assign n44805 = ~n44795 & n44804 ;
  assign n44806 = ~n44794 & n44805 ;
  assign n44807 = n27308 & ~n44806 ;
  assign n44808 = \P2_P3_EAX_reg[27]/NET0131  & ~n42872 ;
  assign n44809 = ~n44807 & ~n44808 ;
  assign n44810 = ~\P1_P2_EAX_reg[27]/NET0131  & ~n43196 ;
  assign n44811 = n43164 & ~n43197 ;
  assign n44812 = ~n44810 & n44811 ;
  assign n44820 = \P1_P2_EAX_reg[27]/NET0131  & n43167 ;
  assign n44821 = ~n43034 & n43065 ;
  assign n44822 = ~n43066 & ~n44821 ;
  assign n44823 = n42875 & n44822 ;
  assign n44813 = \P1_P2_EAX_reg[27]/NET0131  & ~n25773 ;
  assign n44814 = ~\P1_buf2_reg[11]/NET0131  & ~n27934 ;
  assign n44815 = ~\P1_buf1_reg[11]/NET0131  & n27934 ;
  assign n44816 = ~n44814 & ~n44815 ;
  assign n44817 = n25773 & n44816 ;
  assign n44818 = ~n44813 & ~n44817 ;
  assign n44819 = n25776 & ~n44818 ;
  assign n44824 = n25773 & ~n29840 ;
  assign n44825 = ~n44813 & ~n44824 ;
  assign n44826 = n25774 & ~n44825 ;
  assign n44827 = ~n44819 & ~n44826 ;
  assign n44828 = ~n44823 & n44827 ;
  assign n44829 = ~n44820 & n44828 ;
  assign n44830 = ~n44812 & n44829 ;
  assign n44831 = n25918 & ~n44830 ;
  assign n44832 = \P1_P2_EAX_reg[27]/NET0131  & ~n43212 ;
  assign n44833 = ~n44831 & ~n44832 ;
  assign n44835 = ~n25836 & n25918 ;
  assign n44836 = \P1_P2_InstAddrPointer_reg[1]/NET0131  & ~\P1_P2_InstAddrPointer_reg[31]/NET0131  ;
  assign n44837 = \P1_P2_InstAddrPointer_reg[31]/NET0131  & ~n31394 ;
  assign n44838 = ~n44836 & ~n44837 ;
  assign n44839 = n43220 & ~n44838 ;
  assign n44840 = ~n27670 & ~n44839 ;
  assign n44841 = n27609 & ~n44840 ;
  assign n44834 = \P1_P2_InstQueueRd_Addr_reg[2]/NET0131  & ~n43218 ;
  assign n44842 = n25819 & n27608 ;
  assign n44843 = ~n44834 & ~n44842 ;
  assign n44844 = ~n44841 & n44843 ;
  assign n44845 = ~n44835 & n44844 ;
  assign n44847 = n11623 & ~n26047 ;
  assign n44848 = \P2_P1_InstAddrPointer_reg[1]/NET0131  & ~\P2_P1_InstAddrPointer_reg[31]/NET0131  ;
  assign n44849 = \P2_P1_InstAddrPointer_reg[31]/NET0131  & ~n32083 ;
  assign n44850 = ~n44848 & ~n44849 ;
  assign n44851 = n43233 & ~n44850 ;
  assign n44852 = ~n27483 & ~n44851 ;
  assign n44853 = n21096 & ~n44852 ;
  assign n44846 = \P2_P1_InstQueueRd_Addr_reg[2]/NET0131  & ~n43231 ;
  assign n44854 = n11692 & n26028 ;
  assign n44855 = ~n44846 & ~n44854 ;
  assign n44856 = ~n44853 & n44855 ;
  assign n44857 = ~n44847 & n44856 ;
  assign n44859 = \P1_P2_PhyAddrPointer_reg[10]/NET0131  & n25733 ;
  assign n44860 = ~n40566 & ~n44859 ;
  assign n44861 = n25701 & ~n44860 ;
  assign n44862 = \P1_P2_PhyAddrPointer_reg[10]/NET0131  & ~n36590 ;
  assign n44863 = ~n40571 & ~n44862 ;
  assign n44864 = ~n44861 & n44863 ;
  assign n44865 = n25918 & ~n44864 ;
  assign n44871 = n36603 & ~n37915 ;
  assign n44872 = ~\P1_P2_PhyAddrPointer_reg[10]/NET0131  & ~n44871 ;
  assign n44870 = n36604 & ~n37915 ;
  assign n44873 = n25928 & ~n44870 ;
  assign n44874 = ~n44872 & n44873 ;
  assign n44866 = \P1_P2_PhyAddrPointer_reg[1]/NET0131  & n36603 ;
  assign n44867 = ~\P1_P2_PhyAddrPointer_reg[10]/NET0131  & ~n44866 ;
  assign n44868 = ~n41370 & ~n44867 ;
  assign n44869 = n27898 & n44868 ;
  assign n44858 = \P1_P2_PhyAddrPointer_reg[10]/NET0131  & ~n36595 ;
  assign n44875 = ~n40556 & ~n44858 ;
  assign n44876 = ~n44869 & n44875 ;
  assign n44877 = ~n44874 & n44876 ;
  assign n44878 = ~n44865 & n44877 ;
  assign n44880 = n8355 & ~n26185 ;
  assign n44881 = \P1_P1_InstAddrPointer_reg[1]/NET0131  & ~\P1_P1_InstAddrPointer_reg[31]/NET0131  ;
  assign n44882 = \P1_P1_InstAddrPointer_reg[31]/NET0131  & ~n34078 ;
  assign n44883 = ~n44881 & ~n44882 ;
  assign n44884 = n43286 & ~n44883 ;
  assign n44885 = ~n27620 & ~n44884 ;
  assign n44886 = n15322 & ~n44885 ;
  assign n44879 = \P1_P1_InstQueueRd_Addr_reg[2]/NET0131  & ~n43284 ;
  assign n44887 = n8350 & n26119 ;
  assign n44888 = ~n44879 & ~n44887 ;
  assign n44889 = ~n44886 & n44888 ;
  assign n44890 = ~n44880 & n44889 ;
  assign n44894 = \P2_P1_PhyAddrPointer_reg[10]/NET0131  & n25947 ;
  assign n44895 = ~n39945 & ~n44894 ;
  assign n44896 = n25945 & ~n44895 ;
  assign n44897 = \P2_P1_PhyAddrPointer_reg[10]/NET0131  & ~n36677 ;
  assign n44898 = ~n39950 & ~n44897 ;
  assign n44899 = ~n44896 & n44898 ;
  assign n44900 = n11623 & ~n44899 ;
  assign n44902 = n36649 & ~n39474 ;
  assign n44903 = ~\P2_P1_PhyAddrPointer_reg[10]/NET0131  & ~n44902 ;
  assign n44901 = n36650 & ~n39474 ;
  assign n44904 = n11609 & ~n44901 ;
  assign n44905 = ~n44903 & n44904 ;
  assign n44891 = ~\P2_P1_PhyAddrPointer_reg[10]/NET0131  & ~n39455 ;
  assign n44892 = ~n41512 & ~n44891 ;
  assign n44893 = n11613 & n44892 ;
  assign n44906 = \P2_P1_PhyAddrPointer_reg[10]/NET0131  & ~n36687 ;
  assign n44907 = ~n39935 & ~n44906 ;
  assign n44908 = ~n44893 & n44907 ;
  assign n44909 = ~n44905 & n44908 ;
  assign n44910 = ~n44900 & n44909 ;
  assign n44914 = n25701 & n42422 ;
  assign n44915 = \P1_P2_PhyAddrPointer_reg[7]/NET0131  & ~n39340 ;
  assign n44916 = ~n42429 & ~n44915 ;
  assign n44917 = ~n44914 & n44916 ;
  assign n44918 = n25918 & ~n44917 ;
  assign n44911 = ~\P1_P2_PhyAddrPointer_reg[7]/NET0131  & ~n43517 ;
  assign n44912 = ~n43518 & ~n44911 ;
  assign n44919 = ~\P1_P2_DataWidth_reg[1]/NET0131  & ~n44912 ;
  assign n44920 = ~\P1_P2_PhyAddrPointer_reg[7]/NET0131  & ~n36600 ;
  assign n44921 = ~n36601 & ~n44920 ;
  assign n44922 = \P1_P2_DataWidth_reg[1]/NET0131  & ~n44921 ;
  assign n44923 = n25928 & ~n44922 ;
  assign n44924 = ~n44919 & n44923 ;
  assign n44913 = n27898 & n44912 ;
  assign n44925 = \P1_P2_PhyAddrPointer_reg[7]/NET0131  & ~n39352 ;
  assign n44926 = ~n42415 & ~n44925 ;
  assign n44927 = ~n44913 & n44926 ;
  assign n44928 = ~n44924 & n44927 ;
  assign n44929 = ~n44918 & n44928 ;
  assign n44933 = \P1_P2_PhyAddrPointer_reg[9]/NET0131  & n25733 ;
  assign n44934 = ~n42271 & ~n44933 ;
  assign n44935 = n25701 & ~n44934 ;
  assign n44936 = \P1_P2_PhyAddrPointer_reg[9]/NET0131  & ~n36590 ;
  assign n44937 = ~n42278 & ~n44936 ;
  assign n44938 = ~n44935 & n44937 ;
  assign n44939 = n25918 & ~n44938 ;
  assign n44930 = ~\P1_P2_PhyAddrPointer_reg[9]/NET0131  & ~n43520 ;
  assign n44931 = ~n44866 & ~n44930 ;
  assign n44940 = ~\P1_P2_DataWidth_reg[1]/NET0131  & ~n44931 ;
  assign n44941 = ~\P1_P2_PhyAddrPointer_reg[9]/NET0131  & ~n36602 ;
  assign n44942 = ~n36603 & ~n44941 ;
  assign n44943 = \P1_P2_DataWidth_reg[1]/NET0131  & ~n44942 ;
  assign n44944 = n25928 & ~n44943 ;
  assign n44945 = ~n44940 & n44944 ;
  assign n44932 = n27898 & n44931 ;
  assign n44946 = \P1_P2_PhyAddrPointer_reg[9]/NET0131  & ~n39352 ;
  assign n44947 = ~n42259 & ~n44946 ;
  assign n44948 = ~n44932 & n44947 ;
  assign n44949 = ~n44945 & n44948 ;
  assign n44950 = ~n44939 & n44949 ;
  assign n44951 = \P2_P1_PhyAddrPointer_reg[7]/NET0131  & n25947 ;
  assign n44952 = ~n42207 & ~n44951 ;
  assign n44953 = n25945 & ~n44952 ;
  assign n44954 = \P2_P1_PhyAddrPointer_reg[7]/NET0131  & ~n36677 ;
  assign n44955 = ~n42214 & ~n44954 ;
  assign n44956 = ~n44953 & n44955 ;
  assign n44957 = n11623 & ~n44956 ;
  assign n44961 = ~\P2_P1_PhyAddrPointer_reg[7]/NET0131  & ~n43577 ;
  assign n44962 = ~n43578 & ~n44961 ;
  assign n44963 = n36674 & n44962 ;
  assign n44964 = \P2_P1_PhyAddrPointer_reg[7]/NET0131  & ~n36687 ;
  assign n44958 = ~\P2_P1_PhyAddrPointer_reg[7]/NET0131  & ~n36646 ;
  assign n44959 = n27681 & ~n36647 ;
  assign n44960 = ~n44958 & n44959 ;
  assign n44965 = ~n42200 & ~n44960 ;
  assign n44966 = ~n44964 & n44965 ;
  assign n44967 = ~n44963 & n44966 ;
  assign n44968 = ~n44957 & n44967 ;
  assign n44969 = \P2_P1_PhyAddrPointer_reg[9]/NET0131  & n25947 ;
  assign n44970 = ~n42241 & ~n44969 ;
  assign n44971 = n25945 & ~n44970 ;
  assign n44972 = \P2_P1_PhyAddrPointer_reg[9]/NET0131  & ~n36677 ;
  assign n44973 = ~n42246 & ~n44972 ;
  assign n44974 = ~n44971 & n44973 ;
  assign n44975 = n11623 & ~n44974 ;
  assign n44979 = ~\P2_P1_PhyAddrPointer_reg[9]/NET0131  & ~n39454 ;
  assign n44980 = ~n39455 & ~n44979 ;
  assign n44981 = n36674 & n44980 ;
  assign n44976 = ~\P2_P1_PhyAddrPointer_reg[9]/NET0131  & ~n36648 ;
  assign n44977 = n27681 & ~n36649 ;
  assign n44978 = ~n44976 & n44977 ;
  assign n44982 = \P2_P1_PhyAddrPointer_reg[9]/NET0131  & ~n36687 ;
  assign n44983 = ~n42227 & ~n44982 ;
  assign n44984 = ~n44978 & n44983 ;
  assign n44985 = ~n44981 & n44984 ;
  assign n44986 = ~n44975 & n44985 ;
  assign n44988 = \P1_P1_PhyAddrPointer_reg[10]/NET0131  & n26249 ;
  assign n44989 = ~n40289 & ~n44988 ;
  assign n44990 = n26126 & ~n44989 ;
  assign n44991 = \P1_P1_PhyAddrPointer_reg[10]/NET0131  & ~n36696 ;
  assign n44992 = ~n40294 & ~n44991 ;
  assign n44993 = ~n44990 & n44992 ;
  assign n44994 = n8355 & ~n44993 ;
  assign n44998 = \P1_P1_PhyAddrPointer_reg[9]/NET0131  & n43734 ;
  assign n45000 = \P1_P1_PhyAddrPointer_reg[10]/NET0131  & n44998 ;
  assign n44999 = ~\P1_P1_PhyAddrPointer_reg[10]/NET0131  & ~n44998 ;
  assign n45001 = n8282 & ~n44999 ;
  assign n45002 = ~n45000 & n45001 ;
  assign n44995 = ~\P1_P1_PhyAddrPointer_reg[10]/NET0131  & ~n41667 ;
  assign n44996 = ~n41668 & ~n44995 ;
  assign n44997 = n8287 & n44996 ;
  assign n44987 = \P1_P1_PhyAddrPointer_reg[10]/NET0131  & ~n36743 ;
  assign n45003 = ~n40276 & ~n44987 ;
  assign n45004 = ~n44997 & n45003 ;
  assign n45005 = ~n45002 & n45004 ;
  assign n45006 = ~n44994 & n45005 ;
  assign n45007 = \P1_P1_PhyAddrPointer_reg[7]/NET0131  & n26249 ;
  assign n45008 = ~n42449 & ~n45007 ;
  assign n45009 = n26126 & ~n45008 ;
  assign n45010 = \P1_P1_PhyAddrPointer_reg[7]/NET0131  & ~n36696 ;
  assign n45011 = ~n42456 & ~n45010 ;
  assign n45012 = ~n45009 & n45011 ;
  assign n45013 = n8355 & ~n45012 ;
  assign n45017 = ~\P1_P1_PhyAddrPointer_reg[7]/NET0131  & ~n43737 ;
  assign n45018 = ~n43738 & ~n45017 ;
  assign n45019 = ~n36701 & n45018 ;
  assign n45020 = \P1_P1_PhyAddrPointer_reg[7]/NET0131  & ~n36743 ;
  assign n45014 = ~\P1_P1_PhyAddrPointer_reg[7]/NET0131  & ~n36705 ;
  assign n45015 = n27791 & ~n36706 ;
  assign n45016 = ~n45014 & n45015 ;
  assign n45021 = ~n42442 & ~n45016 ;
  assign n45022 = ~n45020 & n45021 ;
  assign n45023 = ~n45019 & n45022 ;
  assign n45024 = ~n45013 & n45023 ;
  assign n45025 = \P1_P1_PhyAddrPointer_reg[9]/NET0131  & n26249 ;
  assign n45026 = ~n42492 & ~n45025 ;
  assign n45027 = n26126 & ~n45026 ;
  assign n45028 = \P1_P1_PhyAddrPointer_reg[9]/NET0131  & ~n36696 ;
  assign n45029 = ~n42499 & ~n45028 ;
  assign n45030 = ~n45027 & n45029 ;
  assign n45031 = n8355 & ~n45030 ;
  assign n45035 = ~\P1_P1_PhyAddrPointer_reg[9]/NET0131  & ~n41666 ;
  assign n45036 = ~n41667 & ~n45035 ;
  assign n45037 = ~n36701 & n45036 ;
  assign n45032 = ~\P1_P1_PhyAddrPointer_reg[9]/NET0131  & ~n36707 ;
  assign n45033 = n27791 & ~n36708 ;
  assign n45034 = ~n45032 & n45033 ;
  assign n45038 = \P1_P1_PhyAddrPointer_reg[9]/NET0131  & ~n36743 ;
  assign n45039 = ~n42482 & ~n45038 ;
  assign n45040 = ~n45034 & n45039 ;
  assign n45041 = ~n45037 & n45040 ;
  assign n45042 = ~n45031 & n45041 ;
  assign n45048 = ~n26718 & n26792 ;
  assign n45049 = \P2_P2_InstAddrPointer_reg[31]/NET0131  & ~n32608 ;
  assign n45050 = ~\P2_P2_InstAddrPointer_reg[1]/NET0131  & ~\P2_P2_InstAddrPointer_reg[31]/NET0131  ;
  assign n45051 = ~n45049 & ~n45050 ;
  assign n45052 = n43246 & n45051 ;
  assign n45053 = ~n27639 & ~n45052 ;
  assign n45054 = n27615 & ~n45053 ;
  assign n45043 = ~n26802 & ~n27637 ;
  assign n45044 = ~n26292 & ~n28046 ;
  assign n45045 = ~n26295 & n45044 ;
  assign n45046 = n45043 & n45045 ;
  assign n45047 = \P2_P2_InstQueueRd_Addr_reg[2]/NET0131  & ~n45046 ;
  assign n45055 = n26690 & n27613 ;
  assign n45056 = ~n45047 & ~n45055 ;
  assign n45057 = ~n45054 & n45056 ;
  assign n45058 = ~n45048 & n45057 ;
  assign n45062 = \P2_P2_PhyAddrPointer_reg[10]/NET0131  & n26629 ;
  assign n45063 = ~n40122 & ~n45062 ;
  assign n45064 = n26621 & ~n45063 ;
  assign n45065 = \P2_P2_PhyAddrPointer_reg[10]/NET0131  & ~n36752 ;
  assign n45066 = ~n40127 & ~n45065 ;
  assign n45067 = ~n45064 & n45066 ;
  assign n45068 = n26792 & ~n45067 ;
  assign n45071 = n36768 & ~n37979 ;
  assign n45069 = n36767 & ~n37979 ;
  assign n45070 = ~\P2_P2_PhyAddrPointer_reg[10]/NET0131  & ~n45069 ;
  assign n45072 = n26794 & ~n45070 ;
  assign n45073 = ~n45071 & n45072 ;
  assign n45059 = ~\P2_P2_PhyAddrPointer_reg[10]/NET0131  & ~n41815 ;
  assign n45060 = ~n41816 & ~n45059 ;
  assign n45061 = n27977 & n45060 ;
  assign n45074 = \P2_P2_PhyAddrPointer_reg[10]/NET0131  & ~n36758 ;
  assign n45075 = ~n40112 & ~n45074 ;
  assign n45076 = ~n45061 & n45075 ;
  assign n45077 = ~n45073 & n45076 ;
  assign n45078 = ~n45068 & n45077 ;
  assign n45084 = \P2_P2_PhyAddrPointer_reg[7]/NET0131  & n26629 ;
  assign n45085 = ~n42301 & ~n45084 ;
  assign n45086 = n26621 & ~n45085 ;
  assign n45087 = \P2_P2_PhyAddrPointer_reg[7]/NET0131  & ~n36752 ;
  assign n45088 = ~n42308 & ~n45087 ;
  assign n45089 = ~n45086 & n45088 ;
  assign n45090 = n26792 & ~n45089 ;
  assign n45079 = \P2_P2_PhyAddrPointer_reg[1]/NET0131  & n36763 ;
  assign n45080 = \P2_P2_PhyAddrPointer_reg[6]/NET0131  & n45079 ;
  assign n45081 = ~\P2_P2_PhyAddrPointer_reg[7]/NET0131  & ~n45080 ;
  assign n45082 = ~n41813 & ~n45081 ;
  assign n45091 = ~\P2_P2_DataWidth_reg[1]/NET0131  & ~n45082 ;
  assign n45092 = ~\P2_P2_PhyAddrPointer_reg[7]/NET0131  & ~n36764 ;
  assign n45093 = ~n36765 & ~n45092 ;
  assign n45094 = \P2_P2_DataWidth_reg[1]/NET0131  & ~n45093 ;
  assign n45095 = n26794 & ~n45094 ;
  assign n45096 = ~n45091 & n45095 ;
  assign n45083 = n27977 & n45082 ;
  assign n45097 = \P2_P2_PhyAddrPointer_reg[7]/NET0131  & ~n36758 ;
  assign n45098 = ~n42293 & ~n45097 ;
  assign n45099 = ~n45083 & n45098 ;
  assign n45100 = ~n45096 & n45099 ;
  assign n45101 = ~n45090 & n45100 ;
  assign n45105 = n26749 & n42331 ;
  assign n45106 = \P2_P2_PhyAddrPointer_reg[9]/NET0131  & ~n41873 ;
  assign n45107 = ~n42339 & ~n45106 ;
  assign n45108 = ~n45105 & n45107 ;
  assign n45109 = n26792 & ~n45108 ;
  assign n45102 = ~\P2_P2_PhyAddrPointer_reg[9]/NET0131  & ~n41814 ;
  assign n45103 = ~n41815 & ~n45102 ;
  assign n45110 = ~\P2_P2_DataWidth_reg[1]/NET0131  & ~n45103 ;
  assign n45111 = ~\P2_P2_PhyAddrPointer_reg[9]/NET0131  & ~n36766 ;
  assign n45112 = ~n36767 & ~n45111 ;
  assign n45113 = \P2_P2_DataWidth_reg[1]/NET0131  & ~n45112 ;
  assign n45114 = n26794 & ~n45113 ;
  assign n45115 = ~n45110 & n45114 ;
  assign n45104 = n27977 & n45103 ;
  assign n45116 = \P2_P2_PhyAddrPointer_reg[9]/NET0131  & ~n36758 ;
  assign n45117 = ~n42320 & ~n45116 ;
  assign n45118 = ~n45104 & n45117 ;
  assign n45119 = ~n45115 & n45118 ;
  assign n45120 = ~n45109 & n45119 ;
  assign n45122 = ~n27269 & n27308 ;
  assign n45123 = \P2_P3_InstAddrPointer_reg[1]/NET0131  & ~\P2_P3_InstAddrPointer_reg[31]/NET0131  ;
  assign n45124 = \P2_P3_InstAddrPointer_reg[31]/NET0131  & ~n33455 ;
  assign n45125 = ~n45123 & ~n45124 ;
  assign n45126 = n43274 & ~n45125 ;
  assign n45127 = ~n27658 & ~n45126 ;
  assign n45128 = n27657 & ~n45127 ;
  assign n45121 = \P2_P3_InstQueueRd_Addr_reg[2]/NET0131  & ~n43272 ;
  assign n45129 = n27251 & n27788 ;
  assign n45130 = ~n45121 & ~n45129 ;
  assign n45131 = ~n45128 & n45130 ;
  assign n45132 = ~n45122 & n45131 ;
  assign n45134 = \P1_P3_PhyAddrPointer_reg[10]/NET0131  & n9072 ;
  assign n45135 = ~n19311 & ~n45134 ;
  assign n45136 = n9064 & ~n45135 ;
  assign n45137 = \P1_P3_PhyAddrPointer_reg[10]/NET0131  & ~n36805 ;
  assign n45138 = ~n19367 & ~n45137 ;
  assign n45139 = ~n45136 & n45138 ;
  assign n45140 = n9241 & ~n45139 ;
  assign n45141 = ~\P1_P3_DataWidth_reg[1]/NET0131  & ~n17665 ;
  assign n45142 = ~\P1_P3_PhyAddrPointer_reg[10]/NET0131  & ~n16459 ;
  assign n45143 = ~n16460 & ~n45142 ;
  assign n45144 = \P1_P3_DataWidth_reg[1]/NET0131  & ~n45143 ;
  assign n45145 = n9245 & ~n45144 ;
  assign n45146 = ~n45141 & n45145 ;
  assign n45133 = n16492 & n17665 ;
  assign n45147 = \P1_P3_PhyAddrPointer_reg[10]/NET0131  & ~n36816 ;
  assign n45148 = ~n19190 & ~n45147 ;
  assign n45149 = ~n45133 & n45148 ;
  assign n45150 = ~n45146 & n45149 ;
  assign n45151 = ~n45140 & n45150 ;
  assign n45152 = \P1_P3_PhyAddrPointer_reg[7]/NET0131  & n9072 ;
  assign n45153 = ~n20554 & ~n45152 ;
  assign n45154 = n9064 & ~n45153 ;
  assign n45155 = \P1_P3_PhyAddrPointer_reg[7]/NET0131  & ~n36805 ;
  assign n45156 = ~n20561 & ~n45155 ;
  assign n45157 = ~n45154 & n45156 ;
  assign n45158 = n9241 & ~n45157 ;
  assign n45162 = n17607 & ~n36810 ;
  assign n45159 = ~\P1_P3_PhyAddrPointer_reg[7]/NET0131  & ~n16456 ;
  assign n45160 = n11698 & ~n16457 ;
  assign n45161 = ~n45159 & n45160 ;
  assign n45163 = \P1_P3_PhyAddrPointer_reg[7]/NET0131  & ~n36816 ;
  assign n45164 = ~n20547 & ~n45163 ;
  assign n45165 = ~n45161 & n45164 ;
  assign n45166 = ~n45162 & n45165 ;
  assign n45167 = ~n45158 & n45166 ;
  assign n45168 = \P2_P3_PhyAddrPointer_reg[10]/NET0131  & ~n27283 ;
  assign n45169 = ~n40350 & ~n45168 ;
  assign n45170 = n27117 & ~n45169 ;
  assign n45171 = \P2_P3_PhyAddrPointer_reg[10]/NET0131  & ~n36826 ;
  assign n45172 = ~n40355 & ~n45171 ;
  assign n45173 = ~n45170 & n45172 ;
  assign n45174 = n27308 & ~n45173 ;
  assign n45178 = ~\P2_P3_PhyAddrPointer_reg[10]/NET0131  & ~n39839 ;
  assign n45179 = ~n39840 & ~n45178 ;
  assign n45180 = n32867 & n45179 ;
  assign n45175 = ~\P2_P3_PhyAddrPointer_reg[10]/NET0131  & ~n44036 ;
  assign n45176 = n27315 & ~n44037 ;
  assign n45177 = ~n45175 & n45176 ;
  assign n45181 = \P2_P3_PhyAddrPointer_reg[10]/NET0131  & ~n36873 ;
  assign n45182 = ~n40339 & ~n45181 ;
  assign n45183 = ~n45177 & n45182 ;
  assign n45184 = ~n45180 & n45183 ;
  assign n45185 = ~n45174 & n45184 ;
  assign n45187 = \P1_P3_PhyAddrPointer_reg[9]/NET0131  & n9072 ;
  assign n45188 = ~n20631 & ~n45187 ;
  assign n45189 = n9064 & ~n45188 ;
  assign n45190 = \P1_P3_PhyAddrPointer_reg[9]/NET0131  & ~n36805 ;
  assign n45191 = ~n20636 & ~n45190 ;
  assign n45192 = ~n45189 & n45191 ;
  assign n45193 = n9241 & ~n45192 ;
  assign n45194 = ~\P1_P3_DataWidth_reg[1]/NET0131  & ~n17900 ;
  assign n45195 = ~\P1_P3_PhyAddrPointer_reg[9]/NET0131  & ~n16458 ;
  assign n45196 = ~n16459 & ~n45195 ;
  assign n45197 = \P1_P3_DataWidth_reg[1]/NET0131  & ~n45196 ;
  assign n45198 = n9245 & ~n45197 ;
  assign n45199 = ~n45194 & n45198 ;
  assign n45186 = n16492 & n17900 ;
  assign n45200 = \P1_P3_PhyAddrPointer_reg[9]/NET0131  & ~n36816 ;
  assign n45201 = ~n20617 & ~n45200 ;
  assign n45202 = ~n45186 & n45201 ;
  assign n45203 = ~n45199 & n45202 ;
  assign n45204 = ~n45193 & n45203 ;
  assign n45208 = \P2_P3_PhyAddrPointer_reg[7]/NET0131  & ~n27283 ;
  assign n45209 = ~n42359 & ~n45208 ;
  assign n45210 = n27117 & ~n45209 ;
  assign n45211 = \P2_P3_PhyAddrPointer_reg[7]/NET0131  & ~n36826 ;
  assign n45212 = ~n42366 & ~n45211 ;
  assign n45213 = ~n45210 & n45212 ;
  assign n45214 = n27308 & ~n45213 ;
  assign n45205 = ~\P2_P3_PhyAddrPointer_reg[7]/NET0131  & ~n44156 ;
  assign n45206 = ~n44157 & ~n45205 ;
  assign n45215 = ~\P2_P3_DataWidth_reg[1]/NET0131  & ~n45206 ;
  assign n45216 = ~\P2_P3_PhyAddrPointer_reg[7]/NET0131  & ~n36838 ;
  assign n45217 = ~n36839 & ~n45216 ;
  assign n45218 = \P2_P3_DataWidth_reg[1]/NET0131  & ~n45217 ;
  assign n45219 = n27315 & ~n45218 ;
  assign n45220 = ~n45215 & n45219 ;
  assign n45207 = n32867 & n45206 ;
  assign n45221 = \P2_P3_PhyAddrPointer_reg[7]/NET0131  & ~n36873 ;
  assign n45222 = ~n42352 & ~n45221 ;
  assign n45223 = ~n45207 & n45222 ;
  assign n45224 = ~n45220 & n45223 ;
  assign n45225 = ~n45214 & n45224 ;
  assign n45226 = \P2_P3_PhyAddrPointer_reg[9]/NET0131  & ~n27283 ;
  assign n45227 = ~n42392 & ~n45226 ;
  assign n45228 = n27117 & ~n45227 ;
  assign n45229 = \P2_P3_PhyAddrPointer_reg[9]/NET0131  & ~n36826 ;
  assign n45230 = ~n42399 & ~n45229 ;
  assign n45231 = ~n45228 & n45230 ;
  assign n45232 = n27308 & ~n45231 ;
  assign n45236 = ~\P2_P3_PhyAddrPointer_reg[9]/NET0131  & ~n39838 ;
  assign n45237 = ~n39839 & ~n45236 ;
  assign n45238 = ~n36831 & n45237 ;
  assign n45233 = ~\P2_P3_PhyAddrPointer_reg[9]/NET0131  & ~n36840 ;
  assign n45234 = n27325 & ~n36841 ;
  assign n45235 = ~n45233 & n45234 ;
  assign n45239 = \P2_P3_PhyAddrPointer_reg[9]/NET0131  & ~n36873 ;
  assign n45240 = ~n42379 & ~n45239 ;
  assign n45241 = ~n45235 & n45240 ;
  assign n45242 = ~n45238 & n45241 ;
  assign n45243 = ~n45232 & n45242 ;
  assign n45245 = n8355 & ~n26244 ;
  assign n45246 = ~\P1_P1_Flush_reg/NET0131  & \P1_P1_InstQueueRd_Addr_reg[3]/NET0131  ;
  assign n45247 = ~n44884 & ~n45246 ;
  assign n45248 = n15322 & ~n45247 ;
  assign n45244 = \P1_P1_InstQueueRd_Addr_reg[3]/NET0131  & ~n43284 ;
  assign n45249 = n8350 & ~n26238 ;
  assign n45250 = ~n45244 & ~n45249 ;
  assign n45251 = ~n45248 & n45250 ;
  assign n45252 = ~n45245 & n45251 ;
  assign n45262 = ~\P2_P1_InstAddrPointer_reg[0]/NET0131  & n26069 ;
  assign n45263 = \P2_P1_InstAddrPointer_reg[0]/NET0131  & ~n25984 ;
  assign n45264 = n26088 & n45263 ;
  assign n45265 = n26055 & n45264 ;
  assign n45266 = ~n45262 & ~n45265 ;
  assign n45255 = \P2_P1_InstAddrPointer_reg[0]/NET0131  & n31785 ;
  assign n45256 = ~n32086 & ~n45255 ;
  assign n45257 = n25964 & n45256 ;
  assign n45258 = \P2_P1_InstAddrPointer_reg[0]/NET0131  & n25947 ;
  assign n45259 = ~n25947 & ~n45256 ;
  assign n45260 = ~n45258 & ~n45259 ;
  assign n45261 = n25945 & ~n45260 ;
  assign n45267 = ~n45257 & ~n45261 ;
  assign n45268 = ~n45266 & n45267 ;
  assign n45269 = n11623 & ~n45268 ;
  assign n45253 = \P2_P1_rEIP_reg[0]/NET0131  & n11616 ;
  assign n45254 = \P2_P1_InstAddrPointer_reg[0]/NET0131  & ~n32172 ;
  assign n45270 = ~n45253 & ~n45254 ;
  assign n45271 = ~n45269 & n45270 ;
  assign n45291 = ~\P2_P1_InstAddrPointer_reg[0]/NET0131  & ~n25987 ;
  assign n45292 = n26069 & ~n45291 ;
  assign n45293 = ~n32083 & ~n45292 ;
  assign n45276 = ~n31753 & ~n31754 ;
  assign n45277 = n45255 & ~n45276 ;
  assign n45274 = ~n32084 & ~n32085 ;
  assign n45275 = ~n45255 & n45274 ;
  assign n45278 = ~n29503 & ~n45275 ;
  assign n45279 = ~n45277 & n45278 ;
  assign n45281 = n31786 & n45276 ;
  assign n45280 = ~n31786 & ~n45276 ;
  assign n45282 = n29503 & ~n45280 ;
  assign n45283 = ~n45281 & n45282 ;
  assign n45284 = ~n45279 & ~n45283 ;
  assign n45285 = n25948 & ~n45284 ;
  assign n45286 = ~n32086 & ~n45274 ;
  assign n45287 = n32086 & ~n45276 ;
  assign n45288 = ~n45286 & ~n45287 ;
  assign n45289 = n25964 & n45288 ;
  assign n45290 = ~n45285 & ~n45289 ;
  assign n45294 = ~\P2_P1_InstAddrPointer_reg[1]/NET0131  & n32159 ;
  assign n45295 = ~n21068 & ~n24901 ;
  assign n45296 = ~n26030 & n45295 ;
  assign n45297 = n21073 & ~n45296 ;
  assign n45298 = \P2_P1_InstAddrPointer_reg[1]/NET0131  & ~n21082 ;
  assign n45299 = ~n26037 & n45298 ;
  assign n45300 = n26056 & n45299 ;
  assign n45301 = ~n45297 & n45300 ;
  assign n45302 = ~n45294 & ~n45301 ;
  assign n45303 = n45290 & ~n45302 ;
  assign n45304 = ~n45293 & n45303 ;
  assign n45305 = n11623 & ~n45304 ;
  assign n45272 = \P2_P1_rEIP_reg[1]/NET0131  & n11616 ;
  assign n45273 = \P2_P1_InstAddrPointer_reg[1]/NET0131  & ~n32172 ;
  assign n45306 = ~n45272 & ~n45273 ;
  assign n45307 = ~n45305 & n45306 ;
  assign n45320 = \P2_P1_InstAddrPointer_reg[2]/NET0131  & n25947 ;
  assign n45326 = ~n31914 & ~n31915 ;
  assign n45328 = n31917 & n45326 ;
  assign n45327 = ~n31917 & ~n45326 ;
  assign n45329 = ~n29503 & ~n45327 ;
  assign n45330 = ~n45328 & n45329 ;
  assign n45321 = ~n31720 & ~n31721 ;
  assign n45323 = n31788 & n45321 ;
  assign n45322 = ~n31788 & ~n45321 ;
  assign n45324 = n29503 & ~n45322 ;
  assign n45325 = ~n45323 & n45324 ;
  assign n45331 = ~n25947 & ~n45325 ;
  assign n45332 = ~n45330 & n45331 ;
  assign n45333 = ~n45320 & ~n45332 ;
  assign n45334 = n25945 & ~n45333 ;
  assign n45310 = ~n25995 & n31913 ;
  assign n45335 = ~n24708 & ~n25984 ;
  assign n45336 = n31688 & ~n45335 ;
  assign n45311 = \P2_P1_InstAddrPointer_reg[2]/NET0131  & ~n35383 ;
  assign n45338 = n32088 & n45326 ;
  assign n45337 = ~n32088 & ~n45326 ;
  assign n45339 = n25964 & ~n45337 ;
  assign n45340 = ~n45338 & n45339 ;
  assign n45312 = ~\P2_P1_InstAddrPointer_reg[2]/NET0131  & ~n20720 ;
  assign n45313 = n20720 & n31913 ;
  assign n45314 = ~n45312 & ~n45313 ;
  assign n45315 = ~n25987 & n45314 ;
  assign n45316 = ~\P2_P1_InstAddrPointer_reg[2]/NET0131  & ~n26057 ;
  assign n45317 = n26057 & ~n31688 ;
  assign n45318 = ~n45316 & ~n45317 ;
  assign n45319 = ~n25952 & n45318 ;
  assign n45341 = ~n45315 & ~n45319 ;
  assign n45342 = ~n45340 & n45341 ;
  assign n45343 = ~n45311 & n45342 ;
  assign n45344 = ~n45336 & n45343 ;
  assign n45345 = ~n45310 & n45344 ;
  assign n45346 = ~n45334 & n45345 ;
  assign n45347 = n11623 & ~n45346 ;
  assign n45308 = \P2_P1_rEIP_reg[2]/NET0131  & n11616 ;
  assign n45309 = \P2_P1_InstAddrPointer_reg[2]/NET0131  & ~n32172 ;
  assign n45348 = ~n45308 & ~n45309 ;
  assign n45349 = ~n45347 & n45348 ;
  assign n45369 = \P2_P1_InstAddrPointer_reg[3]/NET0131  & n25947 ;
  assign n45375 = ~n31910 & ~n31911 ;
  assign n45377 = n31919 & n45375 ;
  assign n45376 = ~n31919 & ~n45375 ;
  assign n45378 = ~n29503 & ~n45376 ;
  assign n45379 = ~n45377 & n45378 ;
  assign n45370 = ~n31685 & ~n31686 ;
  assign n45372 = n31790 & n45370 ;
  assign n45371 = ~n31790 & ~n45370 ;
  assign n45373 = n29503 & ~n45371 ;
  assign n45374 = ~n45372 & n45373 ;
  assign n45380 = ~n25947 & ~n45374 ;
  assign n45381 = ~n45379 & n45380 ;
  assign n45382 = ~n45369 & ~n45381 ;
  assign n45383 = n25945 & ~n45382 ;
  assign n45361 = ~\P2_P1_InstAddrPointer_reg[3]/NET0131  & ~n26006 ;
  assign n45362 = ~n25952 & ~n45361 ;
  assign n45363 = ~n25949 & ~n45362 ;
  assign n45364 = ~n21073 & n31653 ;
  assign n45365 = ~n21073 & ~n26037 ;
  assign n45366 = \P2_P1_InstAddrPointer_reg[3]/NET0131  & ~n45365 ;
  assign n45367 = ~n45364 & ~n45366 ;
  assign n45368 = ~n45363 & ~n45367 ;
  assign n45352 = ~n25995 & n31909 ;
  assign n45359 = \P2_P1_InstAddrPointer_reg[3]/NET0131  & ~n32025 ;
  assign n45354 = ~n32078 & ~n32079 ;
  assign n45356 = ~n32090 & n45354 ;
  assign n45355 = n32090 & ~n45354 ;
  assign n45357 = n25964 & ~n45355 ;
  assign n45358 = ~n45356 & n45357 ;
  assign n45353 = n25984 & n31653 ;
  assign n45360 = n26068 & n32077 ;
  assign n45384 = ~n45353 & ~n45360 ;
  assign n45385 = ~n45358 & n45384 ;
  assign n45386 = ~n45359 & n45385 ;
  assign n45387 = ~n45352 & n45386 ;
  assign n45388 = ~n45368 & n45387 ;
  assign n45389 = ~n45383 & n45388 ;
  assign n45390 = n11623 & ~n45389 ;
  assign n45350 = \P2_P1_rEIP_reg[3]/NET0131  & n11616 ;
  assign n45351 = \P2_P1_InstAddrPointer_reg[3]/NET0131  & ~n32172 ;
  assign n45391 = ~n45350 & ~n45351 ;
  assign n45392 = ~n45390 & n45391 ;
  assign n45397 = \P2_P1_InstAddrPointer_reg[5]/NET0131  & n25947 ;
  assign n45403 = ~n31902 & ~n31903 ;
  assign n45404 = n31923 & ~n45403 ;
  assign n45405 = ~n31923 & n45403 ;
  assign n45406 = ~n45404 & ~n45405 ;
  assign n45407 = ~n29503 & ~n45406 ;
  assign n45398 = ~n31615 & ~n31616 ;
  assign n45400 = n31794 & n45398 ;
  assign n45399 = ~n31794 & ~n45398 ;
  assign n45401 = n29503 & ~n45399 ;
  assign n45402 = ~n45400 & n45401 ;
  assign n45408 = ~n25947 & ~n45402 ;
  assign n45409 = ~n45407 & n45408 ;
  assign n45410 = ~n45397 & ~n45409 ;
  assign n45411 = n25945 & ~n45410 ;
  assign n45416 = ~n32070 & n32095 ;
  assign n45414 = ~n32070 & ~n32071 ;
  assign n45415 = n32094 & ~n45414 ;
  assign n45417 = n25964 & ~n45415 ;
  assign n45418 = ~n45416 & n45417 ;
  assign n45413 = n31583 & ~n32159 ;
  assign n45412 = ~n25995 & n31901 ;
  assign n45395 = \P2_P1_InstAddrPointer_reg[5]/NET0131  & ~n35385 ;
  assign n45396 = n26068 & n32069 ;
  assign n45419 = ~n45395 & ~n45396 ;
  assign n45420 = ~n45412 & n45419 ;
  assign n45421 = ~n45413 & n45420 ;
  assign n45422 = ~n45418 & n45421 ;
  assign n45423 = ~n45411 & n45422 ;
  assign n45424 = n11623 & ~n45423 ;
  assign n45393 = \P2_P1_rEIP_reg[5]/NET0131  & n11616 ;
  assign n45394 = \P2_P1_InstAddrPointer_reg[5]/NET0131  & ~n32172 ;
  assign n45425 = ~n45393 & ~n45394 ;
  assign n45426 = ~n45424 & n45425 ;
  assign n45428 = n11623 & ~n26023 ;
  assign n45429 = ~\P2_P1_Flush_reg/NET0131  & \P2_P1_InstQueueRd_Addr_reg[3]/NET0131  ;
  assign n45430 = ~n44851 & ~n45429 ;
  assign n45431 = n21096 & ~n45430 ;
  assign n45427 = \P2_P1_InstQueueRd_Addr_reg[3]/NET0131  & ~n43231 ;
  assign n45432 = n11692 & ~n25968 ;
  assign n45433 = ~n45427 & ~n45432 ;
  assign n45434 = ~n45431 & n45433 ;
  assign n45435 = ~n45428 & n45434 ;
  assign n45446 = \P1_P2_InstAddrPointer_reg[5]/NET0131  & n25733 ;
  assign n45452 = ~n31220 & ~n31221 ;
  assign n45453 = n31241 & ~n45452 ;
  assign n45454 = ~n31241 & n45452 ;
  assign n45455 = ~n45453 & ~n45454 ;
  assign n45456 = ~n30809 & ~n45455 ;
  assign n45447 = ~n30924 & ~n30925 ;
  assign n45449 = n31103 & n45447 ;
  assign n45448 = ~n31103 & ~n45447 ;
  assign n45450 = n30809 & ~n45448 ;
  assign n45451 = ~n45449 & n45450 ;
  assign n45457 = ~n25733 & ~n45451 ;
  assign n45458 = ~n45456 & n45457 ;
  assign n45459 = ~n45446 & ~n45458 ;
  assign n45460 = n25701 & ~n45459 ;
  assign n45440 = ~n31381 & ~n31382 ;
  assign n45442 = ~n31405 & n45440 ;
  assign n45441 = n31405 & ~n45440 ;
  assign n45443 = n25881 & ~n45441 ;
  assign n45444 = ~n45442 & n45443 ;
  assign n45439 = ~n25817 & n31219 ;
  assign n45438 = ~n25830 & n30892 ;
  assign n45445 = n25887 & n31380 ;
  assign n45461 = \P1_P2_InstAddrPointer_reg[5]/NET0131  & ~n35131 ;
  assign n45462 = ~n45445 & ~n45461 ;
  assign n45463 = ~n45438 & n45462 ;
  assign n45464 = ~n45439 & n45463 ;
  assign n45465 = ~n45444 & n45464 ;
  assign n45466 = ~n45460 & n45465 ;
  assign n45467 = n25918 & ~n45466 ;
  assign n45436 = \P1_P2_rEIP_reg[5]/NET0131  & n27967 ;
  assign n45437 = \P1_P2_InstAddrPointer_reg[5]/NET0131  & ~n31487 ;
  assign n45468 = ~n45436 & ~n45437 ;
  assign n45469 = ~n45467 & n45468 ;
  assign n45481 = ~\P2_P2_InstAddrPointer_reg[0]/NET0131  & ~n26687 ;
  assign n45477 = ~\P2_P2_InstAddrPointer_reg[0]/NET0131  & n26758 ;
  assign n45478 = \P2_P2_InstAddrPointer_reg[0]/NET0131  & n26620 ;
  assign n45479 = n26681 & n45478 ;
  assign n45480 = ~n45477 & ~n45479 ;
  assign n45472 = \P2_P2_InstAddrPointer_reg[0]/NET0131  & n26629 ;
  assign n45473 = ~n32610 & ~n32789 ;
  assign n45474 = ~n26629 & ~n45473 ;
  assign n45475 = ~n45472 & ~n45474 ;
  assign n45476 = n26621 & ~n45475 ;
  assign n45482 = n26744 & n45473 ;
  assign n45483 = ~n45476 & ~n45482 ;
  assign n45484 = ~n45480 & n45483 ;
  assign n45485 = ~n45481 & n45484 ;
  assign n45486 = n26792 & ~n45485 ;
  assign n45470 = \P2_P2_rEIP_reg[0]/NET0131  & n28046 ;
  assign n45471 = \P2_P2_InstAddrPointer_reg[0]/NET0131  & ~n32860 ;
  assign n45487 = ~n45470 & ~n45471 ;
  assign n45488 = ~n45486 & n45487 ;
  assign n45523 = ~n26688 & n32608 ;
  assign n45503 = ~n26630 & n35449 ;
  assign n45504 = \P2_P2_InstAddrPointer_reg[1]/NET0131  & ~n45503 ;
  assign n45508 = ~n32609 & ~n32788 ;
  assign n45509 = ~n32610 & n45508 ;
  assign n45506 = ~n32433 & ~n32434 ;
  assign n45507 = n32610 & ~n45506 ;
  assign n45510 = ~n32510 & ~n45507 ;
  assign n45511 = ~n45509 & n45510 ;
  assign n45513 = n32466 & n45506 ;
  assign n45512 = ~n32466 & ~n45506 ;
  assign n45514 = n32510 & ~n45512 ;
  assign n45515 = ~n45513 & n45514 ;
  assign n45516 = ~n45511 & ~n45515 ;
  assign n45517 = n26749 & ~n45516 ;
  assign n45518 = ~n32789 & ~n45508 ;
  assign n45519 = n32789 & ~n45506 ;
  assign n45520 = ~n45518 & ~n45519 ;
  assign n45521 = n26744 & n45520 ;
  assign n45522 = ~n45517 & ~n45521 ;
  assign n45493 = ~\P2_P2_InstAddrPointer_reg[1]/NET0131  & ~n26286 ;
  assign n45494 = \P2_P2_InstAddrPointer_reg[1]/NET0131  & n26286 ;
  assign n45495 = ~n45493 & ~n45494 ;
  assign n45505 = n26697 & ~n45495 ;
  assign n45492 = ~\P2_P2_InstAddrPointer_reg[1]/NET0131  & ~n26692 ;
  assign n45496 = n26692 & n45495 ;
  assign n45497 = ~n45492 & ~n45496 ;
  assign n45498 = ~n26645 & n45497 ;
  assign n45491 = ~\P2_P2_InstAddrPointer_reg[1]/NET0131  & n26678 ;
  assign n45499 = ~\P2_P2_InstAddrPointer_reg[1]/NET0131  & ~n26611 ;
  assign n45500 = n26611 & ~n32608 ;
  assign n45501 = ~n45499 & ~n45500 ;
  assign n45502 = ~n26583 & n45501 ;
  assign n45524 = ~n45491 & ~n45502 ;
  assign n45525 = ~n45498 & n45524 ;
  assign n45526 = ~n45505 & n45525 ;
  assign n45527 = n45522 & n45526 ;
  assign n45528 = ~n45504 & n45527 ;
  assign n45529 = ~n45523 & n45528 ;
  assign n45530 = n26792 & ~n45529 ;
  assign n45489 = \P2_P2_rEIP_reg[1]/NET0131  & n28046 ;
  assign n45490 = \P2_P2_InstAddrPointer_reg[1]/NET0131  & ~n32860 ;
  assign n45531 = ~n45489 & ~n45490 ;
  assign n45532 = ~n45530 & n45531 ;
  assign n45552 = ~n26688 & n32604 ;
  assign n45536 = ~n26764 & n32368 ;
  assign n45535 = \P2_P2_InstAddrPointer_reg[2]/NET0131  & ~n34266 ;
  assign n45538 = ~n32400 & ~n32401 ;
  assign n45540 = n32468 & n45538 ;
  assign n45539 = ~n32468 & ~n45538 ;
  assign n45541 = n32510 & ~n45539 ;
  assign n45542 = ~n45540 & n45541 ;
  assign n45543 = ~n32605 & ~n32606 ;
  assign n45545 = ~n32612 & n45543 ;
  assign n45544 = n32612 & ~n45543 ;
  assign n45546 = ~n32510 & ~n45544 ;
  assign n45547 = ~n45545 & n45546 ;
  assign n45548 = ~n45542 & ~n45547 ;
  assign n45549 = ~n26629 & ~n45548 ;
  assign n45537 = ~\P2_P2_InstAddrPointer_reg[2]/NET0131  & n26629 ;
  assign n45550 = n26621 & ~n45537 ;
  assign n45551 = ~n45549 & n45550 ;
  assign n45554 = ~n32791 & n45543 ;
  assign n45553 = n32791 & ~n45543 ;
  assign n45555 = n26744 & ~n45553 ;
  assign n45556 = ~n45554 & n45555 ;
  assign n45557 = ~\P2_P2_InstAddrPointer_reg[2]/NET0131  & ~n26611 ;
  assign n45558 = n26611 & n32604 ;
  assign n45559 = ~n45557 & ~n45558 ;
  assign n45560 = ~n26583 & n45559 ;
  assign n45561 = ~n45556 & ~n45560 ;
  assign n45562 = ~n45551 & n45561 ;
  assign n45563 = ~n45535 & n45562 ;
  assign n45564 = ~n45536 & n45563 ;
  assign n45565 = ~n45552 & n45564 ;
  assign n45566 = n26792 & ~n45565 ;
  assign n45533 = \P2_P2_rEIP_reg[2]/NET0131  & n28046 ;
  assign n45534 = \P2_P2_InstAddrPointer_reg[2]/NET0131  & ~n32860 ;
  assign n45567 = ~n45533 & ~n45534 ;
  assign n45568 = ~n45566 & n45567 ;
  assign n45571 = ~n26688 & n32601 ;
  assign n45598 = ~n26583 & n32783 ;
  assign n45599 = n26611 & n45598 ;
  assign n45600 = ~\P2_P2_InstAddrPointer_reg[3]/NET0131  & ~n45599 ;
  assign n45601 = ~n26645 & n32333 ;
  assign n45602 = ~n45598 & ~n45601 ;
  assign n45603 = n32742 & n45602 ;
  assign n45604 = n37169 & n45603 ;
  assign n45605 = ~n45600 & ~n45604 ;
  assign n45584 = ~n32365 & ~n32366 ;
  assign n45585 = n32470 & ~n45584 ;
  assign n45586 = ~n32470 & n45584 ;
  assign n45587 = ~n45585 & ~n45586 ;
  assign n45588 = n32510 & ~n45587 ;
  assign n45589 = ~n32602 & ~n32616 ;
  assign n45591 = n32614 & n45589 ;
  assign n45590 = ~n32614 & ~n45589 ;
  assign n45592 = ~n32510 & ~n45590 ;
  assign n45593 = ~n45591 & n45592 ;
  assign n45594 = ~n45588 & ~n45593 ;
  assign n45595 = ~n26629 & ~n45594 ;
  assign n45583 = ~\P2_P2_InstAddrPointer_reg[3]/NET0131  & n26629 ;
  assign n45596 = n26621 & ~n45583 ;
  assign n45597 = ~n45595 & n45596 ;
  assign n45576 = ~n26678 & ~n26763 ;
  assign n45577 = n32333 & ~n45576 ;
  assign n45572 = ~n26286 & ~n32333 ;
  assign n45573 = ~\P2_P2_InstAddrPointer_reg[3]/NET0131  & n26286 ;
  assign n45574 = ~n45572 & ~n45573 ;
  assign n45575 = n26697 & n45574 ;
  assign n45578 = ~n32784 & ~n32785 ;
  assign n45580 = n32793 & n45578 ;
  assign n45579 = ~n32793 & ~n45578 ;
  assign n45581 = n26744 & ~n45579 ;
  assign n45582 = ~n45580 & n45581 ;
  assign n45606 = ~n45575 & ~n45582 ;
  assign n45607 = ~n45577 & n45606 ;
  assign n45608 = ~n45597 & n45607 ;
  assign n45609 = ~n45605 & n45608 ;
  assign n45610 = ~n45571 & n45609 ;
  assign n45611 = n26792 & ~n45610 ;
  assign n45569 = \P2_P2_rEIP_reg[3]/NET0131  & n28046 ;
  assign n45570 = \P2_P2_InstAddrPointer_reg[3]/NET0131  & ~n32860 ;
  assign n45612 = ~n45569 & ~n45570 ;
  assign n45613 = ~n45611 & n45612 ;
  assign n45619 = \P2_P2_InstAddrPointer_reg[5]/NET0131  & n26629 ;
  assign n45620 = ~n32295 & ~n32296 ;
  assign n45621 = ~n32474 & ~n45620 ;
  assign n45622 = n32474 & n45620 ;
  assign n45623 = ~n45621 & ~n45622 ;
  assign n45624 = ~n26629 & ~n45623 ;
  assign n45625 = ~n45619 & ~n45624 ;
  assign n45626 = n26621 & ~n45625 ;
  assign n45628 = ~n32776 & ~n32777 ;
  assign n45630 = ~n32797 & n45628 ;
  assign n45629 = n32797 & ~n45628 ;
  assign n45631 = n26744 & ~n45629 ;
  assign n45632 = ~n45630 & n45631 ;
  assign n45627 = ~n26688 & n32598 ;
  assign n45618 = \P2_P2_InstAddrPointer_reg[5]/NET0131  & ~n35424 ;
  assign n45616 = n26757 & n32775 ;
  assign n45617 = ~n26764 & n32263 ;
  assign n45633 = ~n45616 & ~n45617 ;
  assign n45634 = ~n45618 & n45633 ;
  assign n45635 = ~n45627 & n45634 ;
  assign n45636 = ~n45632 & n45635 ;
  assign n45637 = ~n45626 & n45636 ;
  assign n45638 = n26792 & ~n45637 ;
  assign n45614 = \P2_P2_rEIP_reg[5]/NET0131  & n28046 ;
  assign n45615 = \P2_P2_InstAddrPointer_reg[5]/NET0131  & ~n32860 ;
  assign n45639 = ~n45614 & ~n45615 ;
  assign n45640 = ~n45638 & n45639 ;
  assign n45642 = ~n26742 & n26792 ;
  assign n45643 = ~\P2_P2_Flush_reg/NET0131  & \P2_P2_InstQueueRd_Addr_reg[3]/NET0131  ;
  assign n45644 = ~n45052 & ~n45643 ;
  assign n45645 = n27615 & ~n45644 ;
  assign n45641 = \P2_P2_InstQueueRd_Addr_reg[3]/NET0131  & ~n45046 ;
  assign n45646 = ~n26721 & n27613 ;
  assign n45647 = ~n45641 & ~n45646 ;
  assign n45648 = ~n45645 & n45647 ;
  assign n45649 = ~n45642 & n45648 ;
  assign n45662 = ~\P1_P3_InstAddrPointer_reg[0]/NET0131  & n9133 ;
  assign n45663 = \P1_P3_InstAddrPointer_reg[0]/NET0131  & ~n9050 ;
  assign n45664 = n9119 & n45663 ;
  assign n45665 = ~n45662 & ~n45664 ;
  assign n45657 = ~\P1_P3_InstAddrPointer_reg[0]/NET0131  & ~n9049 ;
  assign n45658 = \P1_P3_InstAddrPointer_reg[0]/NET0131  & n9049 ;
  assign n45659 = ~n45657 & ~n45658 ;
  assign n45660 = ~n9061 & n45659 ;
  assign n45652 = \P1_P3_InstAddrPointer_reg[0]/NET0131  & n9072 ;
  assign n45653 = ~n18410 & ~n18423 ;
  assign n45654 = ~n9072 & ~n45653 ;
  assign n45655 = ~n45652 & ~n45654 ;
  assign n45656 = n9064 & ~n45655 ;
  assign n45661 = n9191 & n45653 ;
  assign n45666 = ~n45656 & ~n45661 ;
  assign n45667 = ~n45660 & n45666 ;
  assign n45668 = ~n45665 & n45667 ;
  assign n45669 = n9241 & ~n45668 ;
  assign n45650 = \P1_P3_rEIP_reg[0]/NET0131  & n17426 ;
  assign n45651 = \P1_P3_InstAddrPointer_reg[0]/NET0131  & ~n18343 ;
  assign n45670 = ~n45650 & ~n45651 ;
  assign n45671 = ~n45669 & n45670 ;
  assign n45685 = ~\P1_P1_InstAddrPointer_reg[0]/NET0131  & n26151 ;
  assign n45686 = \P1_P1_InstAddrPointer_reg[0]/NET0131  & ~n26251 ;
  assign n45687 = n26132 & n45686 ;
  assign n45688 = ~n45685 & ~n45687 ;
  assign n45680 = ~\P1_P1_InstAddrPointer_reg[0]/NET0131  & ~n15428 ;
  assign n45681 = \P1_P1_InstAddrPointer_reg[0]/NET0131  & n15428 ;
  assign n45682 = ~n45680 & ~n45681 ;
  assign n45683 = ~n26123 & n45682 ;
  assign n45674 = \P1_P1_InstAddrPointer_reg[0]/NET0131  & n26249 ;
  assign n45675 = \P1_P1_InstAddrPointer_reg[0]/NET0131  & n33797 ;
  assign n45676 = ~n34081 & ~n45675 ;
  assign n45677 = ~n26249 & ~n45676 ;
  assign n45678 = ~n45674 & ~n45677 ;
  assign n45679 = n26126 & ~n45678 ;
  assign n45684 = n26263 & n45676 ;
  assign n45689 = ~n45679 & ~n45684 ;
  assign n45690 = ~n45683 & n45689 ;
  assign n45691 = ~n45688 & n45690 ;
  assign n45692 = n8355 & ~n45691 ;
  assign n45672 = \P1_P1_rEIP_reg[0]/NET0131  & n8357 ;
  assign n45673 = \P1_P1_InstAddrPointer_reg[0]/NET0131  & ~n34164 ;
  assign n45693 = ~n45672 & ~n45673 ;
  assign n45694 = ~n45692 & n45693 ;
  assign n45704 = ~\P2_P3_InstAddrPointer_reg[0]/NET0131  & n27220 ;
  assign n45705 = \P2_P3_InstAddrPointer_reg[0]/NET0131  & n27127 ;
  assign n45706 = n27295 & n45705 ;
  assign n45707 = ~n45704 & ~n45706 ;
  assign n45698 = \P2_P3_InstAddrPointer_reg[0]/NET0131  & n33196 ;
  assign n45699 = ~n33458 & ~n45698 ;
  assign n45700 = n27283 & n45699 ;
  assign n45697 = ~\P2_P3_InstAddrPointer_reg[0]/NET0131  & ~n27283 ;
  assign n45701 = n27117 & ~n45697 ;
  assign n45702 = ~n45700 & n45701 ;
  assign n45703 = n27280 & n45699 ;
  assign n45708 = ~n45702 & ~n45703 ;
  assign n45709 = ~n45707 & n45708 ;
  assign n45710 = n27308 & ~n45709 ;
  assign n45695 = \P2_P3_rEIP_reg[0]/NET0131  & n32864 ;
  assign n45696 = \P2_P3_InstAddrPointer_reg[0]/NET0131  & ~n32870 ;
  assign n45711 = ~n45695 & ~n45696 ;
  assign n45712 = ~n45710 & n45711 ;
  assign n45739 = ~\P2_P3_InstAddrPointer_reg[1]/NET0131  & ~n27057 ;
  assign n45740 = n27186 & ~n27227 ;
  assign n45741 = \P2_P3_InstAddrPointer_reg[1]/NET0131  & ~n45740 ;
  assign n45742 = n38706 & n45741 ;
  assign n45743 = ~n45739 & ~n45742 ;
  assign n45715 = ~n27220 & ~n33455 ;
  assign n45731 = \P2_P3_InstAddrPointer_reg[1]/NET0131  & ~n27192 ;
  assign n45732 = ~\P2_P3_InstAddrPointer_reg[1]/NET0131  & n27192 ;
  assign n45733 = ~n45731 & ~n45732 ;
  assign n45734 = ~n27257 & n45733 ;
  assign n45719 = ~n33164 & ~n33165 ;
  assign n45720 = n45698 & ~n45719 ;
  assign n45717 = ~n33456 & ~n33457 ;
  assign n45718 = ~n45698 & n45717 ;
  assign n45721 = ~n33242 & ~n45718 ;
  assign n45722 = ~n45720 & n45721 ;
  assign n45724 = n33197 & n45719 ;
  assign n45723 = ~n33197 & ~n45719 ;
  assign n45725 = n33242 & ~n45723 ;
  assign n45726 = ~n45724 & n45725 ;
  assign n45727 = ~n45722 & ~n45726 ;
  assign n45728 = n27283 & n45727 ;
  assign n45716 = ~\P2_P3_InstAddrPointer_reg[1]/NET0131  & ~n27283 ;
  assign n45729 = n27117 & ~n45716 ;
  assign n45730 = ~n45728 & n45729 ;
  assign n45735 = ~n33458 & ~n45717 ;
  assign n45736 = n33458 & ~n45719 ;
  assign n45737 = ~n45735 & ~n45736 ;
  assign n45738 = n27280 & n45737 ;
  assign n45744 = ~n45730 & ~n45738 ;
  assign n45745 = ~n45734 & n45744 ;
  assign n45746 = ~n45715 & n45745 ;
  assign n45747 = ~n45743 & n45746 ;
  assign n45748 = n27308 & ~n45747 ;
  assign n45713 = \P2_P3_rEIP_reg[1]/NET0131  & n32864 ;
  assign n45714 = \P2_P3_InstAddrPointer_reg[1]/NET0131  & ~n32870 ;
  assign n45749 = ~n45713 & ~n45714 ;
  assign n45750 = ~n45748 & n45749 ;
  assign n45753 = ~n33131 & ~n33132 ;
  assign n45754 = n33199 & ~n45753 ;
  assign n45755 = ~n33199 & n45753 ;
  assign n45756 = ~n45754 & ~n45755 ;
  assign n45757 = n33242 & ~n45756 ;
  assign n45758 = ~n33312 & ~n33313 ;
  assign n45760 = n33315 & n45758 ;
  assign n45759 = ~n33315 & ~n45758 ;
  assign n45761 = ~n33242 & ~n45759 ;
  assign n45762 = ~n45760 & n45761 ;
  assign n45763 = ~n45757 & ~n45762 ;
  assign n45764 = n27283 & ~n45763 ;
  assign n45765 = n27117 & ~n45764 ;
  assign n45766 = n27227 & ~n27275 ;
  assign n45767 = ~n27126 & ~n45766 ;
  assign n45768 = ~n27294 & ~n45767 ;
  assign n45769 = ~n45765 & n45768 ;
  assign n45770 = \P2_P3_InstAddrPointer_reg[2]/NET0131  & ~n45769 ;
  assign n45775 = ~n27229 & n33099 ;
  assign n45780 = ~n27142 & n33311 ;
  assign n45781 = n27284 & n45763 ;
  assign n45772 = n33460 & n45758 ;
  assign n45771 = ~n33460 & ~n45758 ;
  assign n45773 = n27280 & ~n45771 ;
  assign n45774 = ~n45772 & n45773 ;
  assign n45776 = ~\P2_P3_InstAddrPointer_reg[2]/NET0131  & ~n27206 ;
  assign n45777 = n27206 & n33311 ;
  assign n45778 = ~n45776 & ~n45777 ;
  assign n45779 = ~n27111 & n45778 ;
  assign n45782 = ~n45774 & ~n45779 ;
  assign n45783 = ~n45781 & n45782 ;
  assign n45784 = ~n45780 & n45783 ;
  assign n45785 = ~n45775 & n45784 ;
  assign n45786 = ~n45770 & n45785 ;
  assign n45787 = n27308 & ~n45786 ;
  assign n45751 = \P2_P3_rEIP_reg[2]/NET0131  & n32864 ;
  assign n45752 = \P2_P3_InstAddrPointer_reg[2]/NET0131  & ~n32870 ;
  assign n45788 = ~n45751 & ~n45752 ;
  assign n45789 = ~n45787 & n45788 ;
  assign n45792 = \P2_P3_InstAddrPointer_reg[3]/NET0131  & ~n27283 ;
  assign n45798 = ~n33309 & ~n33310 ;
  assign n45799 = n33317 & ~n45798 ;
  assign n45800 = ~n33317 & n45798 ;
  assign n45801 = ~n45799 & ~n45800 ;
  assign n45802 = ~n33242 & ~n45801 ;
  assign n45793 = ~n33096 & ~n33097 ;
  assign n45795 = n33201 & n45793 ;
  assign n45794 = ~n33201 & ~n45793 ;
  assign n45796 = n33242 & ~n45794 ;
  assign n45797 = ~n45795 & n45796 ;
  assign n45803 = n27283 & ~n45797 ;
  assign n45804 = ~n45802 & n45803 ;
  assign n45805 = ~n45792 & ~n45804 ;
  assign n45806 = n27117 & ~n45805 ;
  assign n45821 = n27122 & n27227 ;
  assign n45822 = n27225 & ~n45821 ;
  assign n45823 = n33064 & ~n45822 ;
  assign n45807 = ~n27142 & n33308 ;
  assign n45824 = n27122 & ~n27227 ;
  assign n45825 = ~n27294 & ~n45824 ;
  assign n45826 = ~n27233 & n45825 ;
  assign n45827 = \P2_P3_InstAddrPointer_reg[3]/NET0131  & ~n45826 ;
  assign n45816 = ~n33450 & ~n33451 ;
  assign n45818 = ~n33462 & n45816 ;
  assign n45817 = n33462 & ~n45816 ;
  assign n45819 = n27280 & ~n45817 ;
  assign n45820 = ~n45818 & n45819 ;
  assign n45808 = ~\P2_P3_InstAddrPointer_reg[3]/NET0131  & ~n27206 ;
  assign n45809 = n27206 & ~n33449 ;
  assign n45810 = ~n45808 & ~n45809 ;
  assign n45811 = ~n27111 & n45810 ;
  assign n45813 = n27227 & ~n33064 ;
  assign n45812 = ~\P2_P3_InstAddrPointer_reg[3]/NET0131  & ~n27227 ;
  assign n45814 = n27186 & ~n45812 ;
  assign n45815 = ~n45813 & n45814 ;
  assign n45828 = ~n45811 & ~n45815 ;
  assign n45829 = ~n45820 & n45828 ;
  assign n45830 = ~n45827 & n45829 ;
  assign n45831 = ~n45807 & n45830 ;
  assign n45832 = ~n45823 & n45831 ;
  assign n45833 = ~n45806 & n45832 ;
  assign n45834 = n27308 & ~n45833 ;
  assign n45790 = \P2_P3_rEIP_reg[3]/NET0131  & n32864 ;
  assign n45791 = \P2_P3_InstAddrPointer_reg[3]/NET0131  & ~n32870 ;
  assign n45835 = ~n45790 & ~n45791 ;
  assign n45836 = ~n45834 & n45835 ;
  assign n45847 = \P2_P3_InstAddrPointer_reg[5]/NET0131  & ~n27283 ;
  assign n45848 = ~n33026 & ~n33027 ;
  assign n45850 = ~n33205 & n45848 ;
  assign n45849 = n33205 & ~n45848 ;
  assign n45851 = n27283 & ~n45849 ;
  assign n45852 = ~n45850 & n45851 ;
  assign n45853 = ~n45847 & ~n45852 ;
  assign n45854 = n27117 & ~n45853 ;
  assign n45856 = ~n33442 & ~n33443 ;
  assign n45858 = ~n33466 & n45856 ;
  assign n45857 = n33466 & ~n45856 ;
  assign n45859 = n27280 & ~n45857 ;
  assign n45860 = ~n45858 & n45859 ;
  assign n45846 = ~n27229 & n32994 ;
  assign n45855 = ~n27142 & n33296 ;
  assign n45839 = ~\P2_P3_InstAddrPointer_reg[5]/NET0131  & ~n27206 ;
  assign n45840 = n27206 & ~n33441 ;
  assign n45841 = ~n45839 & ~n45840 ;
  assign n45842 = ~n27111 & n45841 ;
  assign n45843 = ~n27226 & ~n32910 ;
  assign n45844 = n42380 & ~n45843 ;
  assign n45845 = \P2_P3_InstAddrPointer_reg[5]/NET0131  & ~n45844 ;
  assign n45861 = ~n45842 & ~n45845 ;
  assign n45862 = ~n45855 & n45861 ;
  assign n45863 = ~n45846 & n45862 ;
  assign n45864 = ~n45860 & n45863 ;
  assign n45865 = ~n45854 & n45864 ;
  assign n45866 = n27308 & ~n45865 ;
  assign n45837 = \P2_P3_rEIP_reg[5]/NET0131  & n32864 ;
  assign n45838 = \P2_P3_InstAddrPointer_reg[5]/NET0131  & ~n32870 ;
  assign n45867 = ~n45837 & ~n45838 ;
  assign n45868 = ~n45866 & n45867 ;
  assign n45870 = ~n27217 & n27308 ;
  assign n45871 = ~\P2_P3_Flush_reg/NET0131  & \P2_P3_InstQueueRd_Addr_reg[3]/NET0131  ;
  assign n45872 = ~n45126 & ~n45871 ;
  assign n45873 = n27657 & ~n45872 ;
  assign n45869 = \P2_P3_InstQueueRd_Addr_reg[3]/NET0131  & ~n43272 ;
  assign n45874 = ~n27060 & n27788 ;
  assign n45875 = ~n45869 & ~n45874 ;
  assign n45876 = ~n45873 & n45875 ;
  assign n45877 = ~n45870 & n45876 ;
  assign n45899 = ~\P1_P1_InstAddrPointer_reg[1]/NET0131  & ~n26189 ;
  assign n45879 = ~n26193 & ~n34078 ;
  assign n45880 = ~n26250 & n35760 ;
  assign n45881 = \P1_P1_InstAddrPointer_reg[1]/NET0131  & ~n45880 ;
  assign n45884 = ~n33765 & ~n33766 ;
  assign n45885 = n45675 & ~n45884 ;
  assign n45882 = ~n34079 & ~n34080 ;
  assign n45883 = ~n45675 & n45882 ;
  assign n45886 = ~n29558 & ~n45883 ;
  assign n45887 = ~n45885 & n45886 ;
  assign n45889 = n33798 & n45884 ;
  assign n45888 = ~n33798 & ~n45884 ;
  assign n45890 = n29558 & ~n45888 ;
  assign n45891 = ~n45889 & n45890 ;
  assign n45892 = ~n45887 & ~n45891 ;
  assign n45893 = n26262 & ~n45892 ;
  assign n45894 = ~n34081 & ~n45882 ;
  assign n45895 = n34081 & ~n45884 ;
  assign n45896 = ~n45894 & ~n45895 ;
  assign n45897 = n26263 & n45896 ;
  assign n45898 = ~n45893 & ~n45897 ;
  assign n45900 = ~n45881 & n45898 ;
  assign n45901 = ~n45879 & n45900 ;
  assign n45902 = ~n45899 & n45901 ;
  assign n45903 = n8355 & ~n45902 ;
  assign n45878 = \P1_P1_rEIP_reg[1]/NET0131  & n8357 ;
  assign n45904 = \P1_P1_InstAddrPointer_reg[1]/NET0131  & ~n34164 ;
  assign n45905 = ~n45878 & ~n45904 ;
  assign n45906 = ~n45903 & n45905 ;
  assign n45908 = ~n25868 & n25918 ;
  assign n45909 = ~\P1_P2_Flush_reg/NET0131  & \P1_P2_InstQueueRd_Addr_reg[3]/NET0131  ;
  assign n45910 = ~n44839 & ~n45909 ;
  assign n45911 = n27609 & ~n45910 ;
  assign n45907 = \P1_P2_InstQueueRd_Addr_reg[3]/NET0131  & ~n43218 ;
  assign n45912 = ~n25858 & n27608 ;
  assign n45913 = ~n45907 & ~n45912 ;
  assign n45914 = ~n45911 & n45913 ;
  assign n45915 = ~n45908 & n45914 ;
  assign n45944 = ~\P1_P2_InstAddrPointer_reg[1]/NET0131  & ~n25763 ;
  assign n45945 = n25830 & ~n45944 ;
  assign n45946 = n30997 & ~n45945 ;
  assign n45918 = ~n25817 & n31231 ;
  assign n45942 = ~n25752 & n25779 ;
  assign n45943 = \P1_P2_InstAddrPointer_reg[2]/NET0131  & ~n45942 ;
  assign n45928 = \P1_P2_InstAddrPointer_reg[2]/NET0131  & n25733 ;
  assign n45919 = ~n31232 & ~n31233 ;
  assign n45935 = n31235 & n45919 ;
  assign n45934 = ~n31235 & ~n45919 ;
  assign n45936 = ~n30809 & ~n45934 ;
  assign n45937 = ~n45935 & n45936 ;
  assign n45929 = ~n31029 & ~n31030 ;
  assign n45931 = n31097 & n45929 ;
  assign n45930 = ~n31097 & ~n45929 ;
  assign n45932 = n30809 & ~n45930 ;
  assign n45933 = ~n45931 & n45932 ;
  assign n45938 = ~n25733 & ~n45933 ;
  assign n45939 = ~n45937 & n45938 ;
  assign n45940 = ~n45928 & ~n45939 ;
  assign n45941 = n25701 & ~n45940 ;
  assign n45921 = n31399 & n45919 ;
  assign n45920 = ~n31399 & ~n45919 ;
  assign n45922 = n25881 & ~n45920 ;
  assign n45923 = ~n45921 & n45922 ;
  assign n45924 = ~\P1_P2_InstAddrPointer_reg[2]/NET0131  & ~n25747 ;
  assign n45925 = n25747 & n31231 ;
  assign n45926 = ~n45924 & ~n45925 ;
  assign n45927 = ~n25743 & n45926 ;
  assign n45947 = ~n45923 & ~n45927 ;
  assign n45948 = ~n45941 & n45947 ;
  assign n45949 = ~n45943 & n45948 ;
  assign n45950 = ~n45918 & n45949 ;
  assign n45951 = ~n45946 & n45950 ;
  assign n45952 = n25918 & ~n45951 ;
  assign n45916 = \P1_P2_rEIP_reg[2]/NET0131  & n27967 ;
  assign n45917 = \P1_P2_InstAddrPointer_reg[2]/NET0131  & ~n31487 ;
  assign n45953 = ~n45916 & ~n45917 ;
  assign n45954 = ~n45952 & n45953 ;
  assign n45957 = ~\P1_P2_InstAddrPointer_reg[0]/NET0131  & n25901 ;
  assign n45958 = \P1_P2_InstAddrPointer_reg[0]/NET0131  & n25753 ;
  assign n45959 = n25809 & n45958 ;
  assign n45960 = ~n45957 & ~n45959 ;
  assign n45961 = \P1_P2_InstAddrPointer_reg[0]/NET0131  & n25733 ;
  assign n45962 = \P1_P2_InstAddrPointer_reg[0]/NET0131  & n31094 ;
  assign n45963 = ~n31397 & ~n45962 ;
  assign n45964 = ~n25733 & ~n45963 ;
  assign n45965 = ~n45961 & ~n45964 ;
  assign n45966 = n25701 & ~n45965 ;
  assign n45967 = n25881 & n45963 ;
  assign n45968 = ~n45966 & ~n45967 ;
  assign n45969 = ~n45960 & n45968 ;
  assign n45970 = n25918 & ~n45969 ;
  assign n45955 = \P1_P2_rEIP_reg[0]/NET0131  & n27967 ;
  assign n45956 = \P1_P2_InstAddrPointer_reg[0]/NET0131  & ~n31487 ;
  assign n45971 = ~n45955 & ~n45956 ;
  assign n45972 = ~n45970 & n45971 ;
  assign n45995 = ~n26189 & n33700 ;
  assign n45996 = ~n26251 & ~n26255 ;
  assign n45997 = ~n34141 & n45996 ;
  assign n45998 = ~n26197 & ~n26250 ;
  assign n45999 = ~n26266 & n45998 ;
  assign n46000 = n45997 & n45999 ;
  assign n46001 = \P1_P1_InstAddrPointer_reg[2]/NET0131  & ~n46000 ;
  assign n45975 = ~n26151 & n33925 ;
  assign n45976 = ~n33926 & ~n33927 ;
  assign n45977 = n34083 & n45976 ;
  assign n45978 = ~n34083 & ~n45976 ;
  assign n45979 = ~n45977 & ~n45978 ;
  assign n45980 = n26124 & n45979 ;
  assign n45981 = ~n26123 & ~n33925 ;
  assign n45982 = ~n45980 & ~n45981 ;
  assign n45983 = n15428 & ~n45982 ;
  assign n45990 = n33929 & n45976 ;
  assign n45989 = ~n33929 & ~n45976 ;
  assign n45991 = ~n29558 & ~n45989 ;
  assign n45992 = ~n45990 & n45991 ;
  assign n45984 = ~n33732 & ~n33733 ;
  assign n45986 = n33800 & n45984 ;
  assign n45985 = ~n33800 & ~n45984 ;
  assign n45987 = n29558 & ~n45985 ;
  assign n45988 = ~n45986 & n45987 ;
  assign n45993 = n26262 & ~n45988 ;
  assign n45994 = ~n45992 & n45993 ;
  assign n46002 = ~n45983 & ~n45994 ;
  assign n46003 = ~n45975 & n46002 ;
  assign n46004 = ~n46001 & n46003 ;
  assign n46005 = ~n45995 & n46004 ;
  assign n46006 = n8355 & ~n46005 ;
  assign n45973 = \P1_P1_rEIP_reg[2]/NET0131  & n8357 ;
  assign n45974 = \P1_P1_InstAddrPointer_reg[2]/NET0131  & ~n34164 ;
  assign n46007 = ~n45973 & ~n45974 ;
  assign n46008 = ~n46006 & n46007 ;
  assign n46012 = \P1_P1_InstAddrPointer_reg[3]/NET0131  & n26249 ;
  assign n46018 = ~n33922 & ~n33923 ;
  assign n46019 = n33931 & ~n46018 ;
  assign n46020 = ~n33931 & n46018 ;
  assign n46021 = ~n46019 & ~n46020 ;
  assign n46022 = ~n29558 & ~n46021 ;
  assign n46013 = ~n33697 & ~n33698 ;
  assign n46015 = n33802 & n46013 ;
  assign n46014 = ~n33802 & ~n46013 ;
  assign n46016 = n29558 & ~n46014 ;
  assign n46017 = ~n46015 & n46016 ;
  assign n46023 = ~n26249 & ~n46017 ;
  assign n46024 = ~n46022 & n46023 ;
  assign n46025 = ~n46012 & ~n46024 ;
  assign n46026 = n26126 & ~n46025 ;
  assign n46031 = ~n26189 & n33665 ;
  assign n46011 = ~n26151 & n33921 ;
  assign n46032 = ~n26251 & n26256 ;
  assign n46033 = \P1_P1_InstAddrPointer_reg[3]/NET0131  & ~n46032 ;
  assign n46027 = n15428 & ~n34072 ;
  assign n46028 = ~\P1_P1_InstAddrPointer_reg[3]/NET0131  & ~n15428 ;
  assign n46029 = ~n46027 & ~n46028 ;
  assign n46030 = ~n26123 & n46029 ;
  assign n46034 = ~n34073 & ~n34074 ;
  assign n46036 = ~n34085 & n46034 ;
  assign n46035 = n34085 & ~n46034 ;
  assign n46037 = n26263 & ~n46035 ;
  assign n46038 = ~n46036 & n46037 ;
  assign n46039 = ~n46030 & ~n46038 ;
  assign n46040 = ~n46033 & n46039 ;
  assign n46041 = ~n46011 & n46040 ;
  assign n46042 = ~n46031 & n46041 ;
  assign n46043 = ~n46026 & n46042 ;
  assign n46044 = n8355 & ~n46043 ;
  assign n46009 = \P1_P1_rEIP_reg[3]/NET0131  & n8357 ;
  assign n46010 = \P1_P1_InstAddrPointer_reg[3]/NET0131  & ~n34164 ;
  assign n46045 = ~n46009 & ~n46010 ;
  assign n46046 = ~n46044 & n46045 ;
  assign n46050 = ~n25830 & n30811 ;
  assign n46051 = ~\P1_P2_InstAddrPointer_reg[3]/NET0131  & ~n46050 ;
  assign n46049 = n25779 & n30812 ;
  assign n46052 = ~n25809 & ~n46049 ;
  assign n46053 = ~n46051 & n46052 ;
  assign n46069 = ~n25817 & n31227 ;
  assign n46055 = ~n31228 & ~n31229 ;
  assign n46057 = n31237 & n46055 ;
  assign n46056 = ~n31237 & ~n46055 ;
  assign n46058 = ~n30809 & ~n46056 ;
  assign n46059 = ~n46057 & n46058 ;
  assign n46060 = ~n30994 & ~n30995 ;
  assign n46062 = n31099 & n46060 ;
  assign n46061 = ~n31099 & ~n46060 ;
  assign n46063 = n30809 & ~n46061 ;
  assign n46064 = ~n46062 & n46063 ;
  assign n46065 = ~n46059 & ~n46064 ;
  assign n46066 = ~n25733 & ~n46065 ;
  assign n46054 = ~\P1_P2_InstAddrPointer_reg[3]/NET0131  & n25733 ;
  assign n46067 = n25701 & ~n46054 ;
  assign n46068 = ~n46066 & n46067 ;
  assign n46070 = ~\P1_P2_InstAddrPointer_reg[3]/NET0131  & ~n25747 ;
  assign n46071 = ~n25743 & n31388 ;
  assign n46072 = n25753 & ~n46071 ;
  assign n46073 = ~n46070 & ~n46072 ;
  assign n46074 = ~n31389 & ~n31390 ;
  assign n46076 = ~n31401 & n46074 ;
  assign n46075 = n31401 & ~n46074 ;
  assign n46077 = n25881 & ~n46075 ;
  assign n46078 = ~n46076 & n46077 ;
  assign n46079 = ~n46073 & ~n46078 ;
  assign n46080 = ~n46068 & n46079 ;
  assign n46081 = ~n46069 & n46080 ;
  assign n46082 = ~n46053 & n46081 ;
  assign n46083 = n25918 & ~n46082 ;
  assign n46047 = \P1_P2_rEIP_reg[3]/NET0131  & n27967 ;
  assign n46048 = \P1_P2_InstAddrPointer_reg[3]/NET0131  & ~n31487 ;
  assign n46084 = ~n46047 & ~n46048 ;
  assign n46085 = ~n46083 & n46084 ;
  assign n46102 = \P1_P1_InstAddrPointer_reg[5]/NET0131  & n26249 ;
  assign n46108 = ~n33914 & ~n33915 ;
  assign n46110 = ~n33935 & n46108 ;
  assign n46109 = n33935 & ~n46108 ;
  assign n46111 = ~n29558 & ~n46109 ;
  assign n46112 = ~n46110 & n46111 ;
  assign n46103 = ~n33627 & ~n33628 ;
  assign n46105 = n33806 & n46103 ;
  assign n46104 = ~n33806 & ~n46103 ;
  assign n46106 = n29558 & ~n46104 ;
  assign n46107 = ~n46105 & n46106 ;
  assign n46113 = ~n26249 & ~n46107 ;
  assign n46114 = ~n46112 & n46113 ;
  assign n46115 = ~n46102 & ~n46114 ;
  assign n46116 = n26126 & ~n46115 ;
  assign n46092 = ~n34065 & ~n34066 ;
  assign n46094 = ~n34089 & n46092 ;
  assign n46093 = n34089 & ~n46092 ;
  assign n46095 = n26263 & ~n46093 ;
  assign n46096 = ~n46094 & n46095 ;
  assign n46091 = ~n26189 & n33595 ;
  assign n46101 = ~n26151 & n33913 ;
  assign n46087 = ~n15383 & ~n24504 ;
  assign n46088 = n15335 & ~n46087 ;
  assign n46089 = n45997 & ~n46088 ;
  assign n46090 = \P1_P1_InstAddrPointer_reg[5]/NET0131  & ~n46089 ;
  assign n46097 = ~\P1_P1_InstAddrPointer_reg[5]/NET0131  & ~n15428 ;
  assign n46098 = n15428 & ~n34064 ;
  assign n46099 = ~n46097 & ~n46098 ;
  assign n46100 = ~n26123 & n46099 ;
  assign n46117 = ~n46090 & ~n46100 ;
  assign n46118 = ~n46101 & n46117 ;
  assign n46119 = ~n46091 & n46118 ;
  assign n46120 = ~n46096 & n46119 ;
  assign n46121 = ~n46116 & n46120 ;
  assign n46122 = n8355 & ~n46121 ;
  assign n46086 = \P1_P1_rEIP_reg[5]/NET0131  & n8357 ;
  assign n46123 = \P1_P1_InstAddrPointer_reg[5]/NET0131  & ~n34164 ;
  assign n46124 = ~n46086 & ~n46123 ;
  assign n46125 = ~n46122 & n46124 ;
  assign n46136 = ~n25817 & ~n31394 ;
  assign n46154 = ~\P1_P2_InstAddrPointer_reg[1]/NET0131  & ~n25808 ;
  assign n46155 = \P1_P2_InstAddrPointer_reg[1]/NET0131  & ~n25734 ;
  assign n46156 = n36898 & n46155 ;
  assign n46157 = ~n46154 & ~n46156 ;
  assign n46128 = \P1_P2_InstAddrPointer_reg[1]/NET0131  & ~n25415 ;
  assign n46129 = ~\P1_P2_InstAddrPointer_reg[1]/NET0131  & n25415 ;
  assign n46130 = ~n46128 & ~n46129 ;
  assign n46131 = ~n36900 & n46130 ;
  assign n46132 = ~\P1_P2_InstAddrPointer_reg[1]/NET0131  & ~n25747 ;
  assign n46133 = n25747 & n31394 ;
  assign n46134 = ~n46132 & ~n46133 ;
  assign n46135 = ~n25743 & n46134 ;
  assign n46139 = ~n31062 & ~n31063 ;
  assign n46140 = n45962 & ~n46139 ;
  assign n46137 = ~n31395 & ~n31396 ;
  assign n46138 = ~n45962 & n46137 ;
  assign n46141 = ~n30809 & ~n46138 ;
  assign n46142 = ~n46140 & n46141 ;
  assign n46144 = n31095 & n46139 ;
  assign n46143 = ~n31095 & ~n46139 ;
  assign n46145 = n30809 & ~n46143 ;
  assign n46146 = ~n46144 & n46145 ;
  assign n46147 = ~n46142 & ~n46146 ;
  assign n46148 = n25874 & ~n46147 ;
  assign n46149 = ~n31397 & ~n46137 ;
  assign n46150 = n31397 & ~n46139 ;
  assign n46151 = ~n46149 & ~n46150 ;
  assign n46152 = n25881 & n46151 ;
  assign n46153 = ~n46148 & ~n46152 ;
  assign n46158 = ~n46135 & n46153 ;
  assign n46159 = ~n46131 & n46158 ;
  assign n46160 = ~n46157 & n46159 ;
  assign n46161 = ~n46136 & n46160 ;
  assign n46162 = n25918 & ~n46161 ;
  assign n46126 = \P1_P2_rEIP_reg[1]/NET0131  & n27967 ;
  assign n46127 = \P1_P2_InstAddrPointer_reg[1]/NET0131  & ~n31487 ;
  assign n46163 = ~n46126 & ~n46127 ;
  assign n46164 = ~n46162 & n46163 ;
  assign n46166 = ~n25898 & n25918 ;
  assign n46167 = ~\P1_P2_Flush_reg/NET0131  & \P1_P2_InstQueueRd_Addr_reg[1]/NET0131  ;
  assign n46168 = n43220 & n44838 ;
  assign n46169 = ~n46167 & ~n46168 ;
  assign n46170 = n27609 & ~n46169 ;
  assign n46165 = \P1_P2_InstQueueRd_Addr_reg[1]/NET0131  & ~n43218 ;
  assign n46171 = ~n25885 & n27608 ;
  assign n46172 = ~n46165 & ~n46171 ;
  assign n46173 = ~n46170 & n46172 ;
  assign n46174 = ~n46166 & n46173 ;
  assign n46176 = n11623 & ~n26084 ;
  assign n46177 = ~\P2_P1_Flush_reg/NET0131  & \P2_P1_InstQueueRd_Addr_reg[1]/NET0131  ;
  assign n46178 = n43233 & n44850 ;
  assign n46179 = ~n46177 & ~n46178 ;
  assign n46180 = n21096 & ~n46179 ;
  assign n46175 = \P2_P1_InstQueueRd_Addr_reg[1]/NET0131  & ~n43231 ;
  assign n46181 = n11692 & n26070 ;
  assign n46182 = ~n46175 & ~n46181 ;
  assign n46183 = ~n46180 & n46182 ;
  assign n46184 = ~n46176 & n46183 ;
  assign n46186 = ~n26770 & n26792 ;
  assign n46187 = ~\P2_P2_Flush_reg/NET0131  & \P2_P2_InstQueueRd_Addr_reg[1]/NET0131  ;
  assign n46188 = n43246 & ~n45051 ;
  assign n46189 = ~n46187 & ~n46188 ;
  assign n46190 = n27615 & ~n46189 ;
  assign n46185 = \P2_P2_InstQueueRd_Addr_reg[1]/NET0131  & ~n45046 ;
  assign n46191 = n26756 & n27613 ;
  assign n46192 = ~n46185 & ~n46191 ;
  assign n46193 = ~n46190 & n46192 ;
  assign n46194 = ~n46186 & n46193 ;
  assign n46196 = ~n27240 & n27308 ;
  assign n46197 = ~\P2_P3_Flush_reg/NET0131  & \P2_P3_InstQueueRd_Addr_reg[1]/NET0131  ;
  assign n46198 = n43274 & n45125 ;
  assign n46199 = ~n46197 & ~n46198 ;
  assign n46200 = n27657 & ~n46199 ;
  assign n46195 = \P2_P3_InstQueueRd_Addr_reg[1]/NET0131  & ~n43272 ;
  assign n46201 = n27221 & n27788 ;
  assign n46202 = ~n46195 & ~n46201 ;
  assign n46203 = ~n46200 & n46202 ;
  assign n46204 = ~n46196 & n46203 ;
  assign n46206 = n8355 & ~n26206 ;
  assign n46207 = ~\P1_P1_Flush_reg/NET0131  & \P1_P1_InstQueueRd_Addr_reg[1]/NET0131  ;
  assign n46208 = n43286 & n44883 ;
  assign n46209 = ~n46207 & ~n46208 ;
  assign n46210 = n15322 & ~n46209 ;
  assign n46205 = \P1_P1_InstQueueRd_Addr_reg[1]/NET0131  & ~n43284 ;
  assign n46211 = n8350 & n26191 ;
  assign n46212 = ~n46205 & ~n46211 ;
  assign n46213 = ~n46210 & n46212 ;
  assign n46214 = ~n46206 & n46213 ;
  assign n46215 = \P2_P1_EAX_reg[3]/NET0131  & ~n27438 ;
  assign n46217 = ~n21069 & n24487 ;
  assign n46216 = n20728 & ~n31684 ;
  assign n46218 = ~\P2_P1_EAX_reg[3]/NET0131  & ~n21024 ;
  assign n46219 = ~n21025 & ~n46218 ;
  assign n46220 = n21022 & n46219 ;
  assign n46221 = ~n46216 & ~n46220 ;
  assign n46222 = ~n46217 & n46221 ;
  assign n46223 = n11623 & ~n46222 ;
  assign n46224 = ~n46215 & ~n46223 ;
  assign n46230 = \P2_P1_EBX_reg[0]/NET0131  & \P2_P1_EBX_reg[1]/NET0131  ;
  assign n46231 = \P2_P1_EBX_reg[2]/NET0131  & n46230 ;
  assign n46232 = \P2_P1_EBX_reg[3]/NET0131  & n46231 ;
  assign n46233 = \P2_P1_EBX_reg[4]/NET0131  & n46232 ;
  assign n46234 = \P2_P1_EBX_reg[5]/NET0131  & n46233 ;
  assign n46235 = \P2_P1_EBX_reg[6]/NET0131  & n46234 ;
  assign n46236 = \P2_P1_EBX_reg[7]/NET0131  & n46235 ;
  assign n46237 = \P2_P1_EBX_reg[8]/NET0131  & n46236 ;
  assign n46238 = \P2_P1_EBX_reg[9]/NET0131  & n46237 ;
  assign n46239 = \P2_P1_EBX_reg[10]/NET0131  & n46238 ;
  assign n46240 = \P2_P1_EBX_reg[11]/NET0131  & n46239 ;
  assign n46241 = \P2_P1_EBX_reg[12]/NET0131  & n46240 ;
  assign n46242 = \P2_P1_EBX_reg[13]/NET0131  & n46241 ;
  assign n46243 = \P2_P1_EBX_reg[14]/NET0131  & n46242 ;
  assign n46244 = \P2_P1_EBX_reg[15]/NET0131  & n46243 ;
  assign n46245 = \P2_P1_EBX_reg[16]/NET0131  & n46244 ;
  assign n46246 = \P2_P1_EBX_reg[17]/NET0131  & n46245 ;
  assign n46247 = \P2_P1_EBX_reg[18]/NET0131  & n46246 ;
  assign n46248 = \P2_P1_EBX_reg[19]/NET0131  & n46247 ;
  assign n46249 = \P2_P1_EBX_reg[20]/NET0131  & n46248 ;
  assign n46250 = \P2_P1_EBX_reg[21]/NET0131  & n46249 ;
  assign n46251 = \P2_P1_EBX_reg[22]/NET0131  & n46250 ;
  assign n46252 = \P2_P1_EBX_reg[23]/NET0131  & n46251 ;
  assign n46253 = \P2_P1_EBX_reg[24]/NET0131  & n46252 ;
  assign n46254 = \P2_P1_EBX_reg[25]/NET0131  & n46253 ;
  assign n46255 = \P2_P1_EBX_reg[26]/NET0131  & n46254 ;
  assign n46257 = \P2_P1_EBX_reg[27]/NET0131  & n46255 ;
  assign n46256 = ~\P2_P1_EBX_reg[27]/NET0131  & ~n46255 ;
  assign n46258 = n25981 & ~n46256 ;
  assign n46259 = ~n46257 & n46258 ;
  assign n46225 = n20720 & n25986 ;
  assign n46226 = n25981 & ~n25986 ;
  assign n46227 = ~n46225 & ~n46226 ;
  assign n46228 = \P2_P1_EBX_reg[27]/NET0131  & n46227 ;
  assign n46229 = n23855 & n46225 ;
  assign n46260 = ~n46228 & ~n46229 ;
  assign n46261 = ~n46259 & n46260 ;
  assign n46262 = n11623 & ~n46261 ;
  assign n46263 = \P2_P1_EBX_reg[27]/NET0131  & ~n21100 ;
  assign n46264 = ~n46262 & ~n46263 ;
  assign n46267 = \P2_P1_EBX_reg[28]/NET0131  & n46257 ;
  assign n46268 = \P2_P1_EBX_reg[29]/NET0131  & n46267 ;
  assign n46269 = \P2_P1_EBX_reg[30]/NET0131  & n46268 ;
  assign n46271 = \P2_P1_EBX_reg[31]/NET0131  & n46269 ;
  assign n46270 = ~\P2_P1_EBX_reg[31]/NET0131  & ~n46269 ;
  assign n46272 = n25981 & ~n46270 ;
  assign n46273 = ~n46271 & n46272 ;
  assign n46265 = n21015 & n46225 ;
  assign n46266 = \P2_P1_EBX_reg[31]/NET0131  & n46227 ;
  assign n46274 = ~n46265 & ~n46266 ;
  assign n46275 = ~n46273 & n46274 ;
  assign n46276 = n11623 & ~n46275 ;
  assign n46277 = \P2_P1_EBX_reg[31]/NET0131  & ~n21100 ;
  assign n46278 = ~n46276 & ~n46277 ;
  assign n46279 = \P2_P2_EAX_reg[30]/NET0131  & ~n44508 ;
  assign n46390 = \P2_P2_EAX_reg[28]/NET0131  & n44731 ;
  assign n46391 = \P2_P2_EAX_reg[29]/NET0131  & n46390 ;
  assign n46393 = ~\P2_P2_EAX_reg[30]/NET0131  & ~n46391 ;
  assign n46392 = \P2_P2_EAX_reg[30]/NET0131  & n46391 ;
  assign n46394 = n44732 & ~n46392 ;
  assign n46395 = ~n46393 & n46394 ;
  assign n46299 = \P2_P2_InstQueue_reg[2][5]/NET0131  & n26330 ;
  assign n46297 = \P2_P2_InstQueue_reg[3][5]/NET0131  & n26325 ;
  assign n46288 = \P2_P2_InstQueue_reg[10][5]/NET0131  & n26300 ;
  assign n46289 = \P2_P2_InstQueue_reg[9][5]/NET0131  & n26318 ;
  assign n46304 = ~n46288 & ~n46289 ;
  assign n46314 = ~n46297 & n46304 ;
  assign n46315 = ~n46299 & n46314 ;
  assign n46300 = \P2_P2_InstQueue_reg[13][5]/NET0131  & n26304 ;
  assign n46301 = \P2_P2_InstQueue_reg[6][5]/NET0131  & n26316 ;
  assign n46309 = ~n46300 & ~n46301 ;
  assign n46302 = \P2_P2_InstQueue_reg[12][5]/NET0131  & n26334 ;
  assign n46303 = \P2_P2_InstQueue_reg[4][5]/NET0131  & n26322 ;
  assign n46310 = ~n46302 & ~n46303 ;
  assign n46311 = n46309 & n46310 ;
  assign n46294 = \P2_P2_InstQueue_reg[8][5]/NET0131  & n26307 ;
  assign n46295 = \P2_P2_InstQueue_reg[0][5]/NET0131  & n26313 ;
  assign n46307 = ~n46294 & ~n46295 ;
  assign n46296 = \P2_P2_InstQueue_reg[5][5]/NET0131  & n26338 ;
  assign n46298 = \P2_P2_InstQueue_reg[11][5]/NET0131  & n26327 ;
  assign n46308 = ~n46296 & ~n46298 ;
  assign n46312 = n46307 & n46308 ;
  assign n46290 = \P2_P2_InstQueue_reg[7][5]/NET0131  & n26332 ;
  assign n46291 = \P2_P2_InstQueue_reg[14][5]/NET0131  & n26320 ;
  assign n46305 = ~n46290 & ~n46291 ;
  assign n46292 = \P2_P2_InstQueue_reg[1][5]/NET0131  & n26336 ;
  assign n46293 = \P2_P2_InstQueue_reg[15][5]/NET0131  & n26310 ;
  assign n46306 = ~n46292 & ~n46293 ;
  assign n46313 = n46305 & n46306 ;
  assign n46316 = n46312 & n46313 ;
  assign n46317 = n46311 & n46316 ;
  assign n46318 = n46315 & n46317 ;
  assign n46319 = n44702 & ~n46318 ;
  assign n46331 = \P2_P2_InstQueue_reg[2][6]/NET0131  & n26330 ;
  assign n46329 = \P2_P2_InstQueue_reg[3][6]/NET0131  & n26325 ;
  assign n46320 = \P2_P2_InstQueue_reg[10][6]/NET0131  & n26300 ;
  assign n46321 = \P2_P2_InstQueue_reg[9][6]/NET0131  & n26318 ;
  assign n46336 = ~n46320 & ~n46321 ;
  assign n46346 = ~n46329 & n46336 ;
  assign n46347 = ~n46331 & n46346 ;
  assign n46332 = \P2_P2_InstQueue_reg[13][6]/NET0131  & n26304 ;
  assign n46333 = \P2_P2_InstQueue_reg[6][6]/NET0131  & n26316 ;
  assign n46341 = ~n46332 & ~n46333 ;
  assign n46334 = \P2_P2_InstQueue_reg[12][6]/NET0131  & n26334 ;
  assign n46335 = \P2_P2_InstQueue_reg[4][6]/NET0131  & n26322 ;
  assign n46342 = ~n46334 & ~n46335 ;
  assign n46343 = n46341 & n46342 ;
  assign n46326 = \P2_P2_InstQueue_reg[8][6]/NET0131  & n26307 ;
  assign n46327 = \P2_P2_InstQueue_reg[0][6]/NET0131  & n26313 ;
  assign n46339 = ~n46326 & ~n46327 ;
  assign n46328 = \P2_P2_InstQueue_reg[5][6]/NET0131  & n26338 ;
  assign n46330 = \P2_P2_InstQueue_reg[11][6]/NET0131  & n26327 ;
  assign n46340 = ~n46328 & ~n46330 ;
  assign n46344 = n46339 & n46340 ;
  assign n46322 = \P2_P2_InstQueue_reg[7][6]/NET0131  & n26332 ;
  assign n46323 = \P2_P2_InstQueue_reg[14][6]/NET0131  & n26320 ;
  assign n46337 = ~n46322 & ~n46323 ;
  assign n46324 = \P2_P2_InstQueue_reg[1][6]/NET0131  & n26336 ;
  assign n46325 = \P2_P2_InstQueue_reg[15][6]/NET0131  & n26310 ;
  assign n46338 = ~n46324 & ~n46325 ;
  assign n46345 = n46337 & n46338 ;
  assign n46348 = n46344 & n46345 ;
  assign n46349 = n46343 & n46348 ;
  assign n46350 = n46347 & n46349 ;
  assign n46351 = n46319 & ~n46350 ;
  assign n46363 = \P2_P2_InstQueue_reg[2][7]/NET0131  & n26330 ;
  assign n46361 = \P2_P2_InstQueue_reg[3][7]/NET0131  & n26325 ;
  assign n46352 = \P2_P2_InstQueue_reg[10][7]/NET0131  & n26300 ;
  assign n46353 = \P2_P2_InstQueue_reg[13][7]/NET0131  & n26304 ;
  assign n46368 = ~n46352 & ~n46353 ;
  assign n46378 = ~n46361 & n46368 ;
  assign n46379 = ~n46363 & n46378 ;
  assign n46364 = \P2_P2_InstQueue_reg[9][7]/NET0131  & n26318 ;
  assign n46365 = \P2_P2_InstQueue_reg[4][7]/NET0131  & n26322 ;
  assign n46373 = ~n46364 & ~n46365 ;
  assign n46366 = \P2_P2_InstQueue_reg[6][7]/NET0131  & n26316 ;
  assign n46367 = \P2_P2_InstQueue_reg[15][7]/NET0131  & n26310 ;
  assign n46374 = ~n46366 & ~n46367 ;
  assign n46375 = n46373 & n46374 ;
  assign n46358 = \P2_P2_InstQueue_reg[8][7]/NET0131  & n26307 ;
  assign n46359 = \P2_P2_InstQueue_reg[1][7]/NET0131  & n26336 ;
  assign n46371 = ~n46358 & ~n46359 ;
  assign n46360 = \P2_P2_InstQueue_reg[7][7]/NET0131  & n26332 ;
  assign n46362 = \P2_P2_InstQueue_reg[11][7]/NET0131  & n26327 ;
  assign n46372 = ~n46360 & ~n46362 ;
  assign n46376 = n46371 & n46372 ;
  assign n46354 = \P2_P2_InstQueue_reg[14][7]/NET0131  & n26320 ;
  assign n46355 = \P2_P2_InstQueue_reg[12][7]/NET0131  & n26334 ;
  assign n46369 = ~n46354 & ~n46355 ;
  assign n46356 = \P2_P2_InstQueue_reg[5][7]/NET0131  & n26338 ;
  assign n46357 = \P2_P2_InstQueue_reg[0][7]/NET0131  & n26313 ;
  assign n46370 = ~n46356 & ~n46357 ;
  assign n46377 = n46369 & n46370 ;
  assign n46380 = n46376 & n46377 ;
  assign n46381 = n46375 & n46380 ;
  assign n46382 = n46379 & n46381 ;
  assign n46383 = ~n46351 & n46382 ;
  assign n46384 = n46351 & ~n46382 ;
  assign n46385 = ~n46383 & ~n46384 ;
  assign n46386 = n44510 & n46385 ;
  assign n46287 = \P2_P2_EAX_reg[30]/NET0131  & n44736 ;
  assign n46280 = \P2_P2_EAX_reg[30]/NET0131  & ~n26641 ;
  assign n46281 = \P2_buf2_reg[14]/NET0131  & ~n28013 ;
  assign n46282 = \P2_buf1_reg[14]/NET0131  & n28013 ;
  assign n46283 = ~n46281 & ~n46282 ;
  assign n46284 = n26641 & ~n46283 ;
  assign n46285 = ~n46280 & ~n46284 ;
  assign n46286 = n26633 & ~n46285 ;
  assign n46387 = n26641 & ~n34488 ;
  assign n46388 = ~n46280 & ~n46387 ;
  assign n46389 = n26638 & ~n46388 ;
  assign n46396 = ~n46286 & ~n46389 ;
  assign n46397 = ~n46287 & n46396 ;
  assign n46398 = ~n46386 & n46397 ;
  assign n46399 = ~n46395 & n46398 ;
  assign n46400 = n26792 & ~n46399 ;
  assign n46401 = ~n46279 & ~n46400 ;
  assign n46408 = \P2_P2_EAX_reg[31]/NET0131  & n46392 ;
  assign n46407 = ~\P2_P2_EAX_reg[31]/NET0131  & ~n46392 ;
  assign n46409 = n44732 & ~n46407 ;
  assign n46410 = ~n46408 & n46409 ;
  assign n46402 = ~n26642 & ~n44736 ;
  assign n46403 = \P2_P2_EAX_reg[31]/NET0131  & ~n46402 ;
  assign n46404 = \P2_P2_EAX_reg[31]/NET0131  & ~n44735 ;
  assign n46405 = ~n44510 & ~n46404 ;
  assign n46406 = n46384 & ~n46405 ;
  assign n46411 = ~n46403 & ~n46406 ;
  assign n46412 = ~n46410 & n46411 ;
  assign n46413 = n26792 & ~n46412 ;
  assign n46414 = \P2_P2_EAX_reg[31]/NET0131  & ~n44508 ;
  assign n46415 = ~n46413 & ~n46414 ;
  assign n46420 = \P2_P2_EBX_reg[0]/NET0131  & \P2_P2_EBX_reg[1]/NET0131  ;
  assign n46421 = \P2_P2_EBX_reg[2]/NET0131  & n46420 ;
  assign n46422 = \P2_P2_EBX_reg[3]/NET0131  & n46421 ;
  assign n46423 = \P2_P2_EBX_reg[4]/NET0131  & n46422 ;
  assign n46424 = \P2_P2_EBX_reg[5]/NET0131  & n46423 ;
  assign n46425 = \P2_P2_EBX_reg[6]/NET0131  & n46424 ;
  assign n46426 = \P2_P2_EBX_reg[7]/NET0131  & n46425 ;
  assign n46427 = \P2_P2_EBX_reg[8]/NET0131  & n46426 ;
  assign n46428 = \P2_P2_EBX_reg[9]/NET0131  & n46427 ;
  assign n46429 = \P2_P2_EBX_reg[10]/NET0131  & n46428 ;
  assign n46430 = \P2_P2_EBX_reg[11]/NET0131  & n46429 ;
  assign n46431 = \P2_P2_EBX_reg[12]/NET0131  & n46430 ;
  assign n46432 = \P2_P2_EBX_reg[13]/NET0131  & n46431 ;
  assign n46433 = \P2_P2_EBX_reg[14]/NET0131  & n46432 ;
  assign n46434 = \P2_P2_EBX_reg[15]/NET0131  & n46433 ;
  assign n46435 = \P2_P2_EBX_reg[16]/NET0131  & n46434 ;
  assign n46436 = \P2_P2_EBX_reg[17]/NET0131  & n46435 ;
  assign n46437 = \P2_P2_EBX_reg[18]/NET0131  & n46436 ;
  assign n46438 = \P2_P2_EBX_reg[19]/NET0131  & n46437 ;
  assign n46439 = \P2_P2_EBX_reg[20]/NET0131  & n46438 ;
  assign n46440 = \P2_P2_EBX_reg[21]/NET0131  & n46439 ;
  assign n46441 = \P2_P2_EBX_reg[22]/NET0131  & n46440 ;
  assign n46442 = \P2_P2_EBX_reg[23]/NET0131  & n46441 ;
  assign n46443 = \P2_P2_EBX_reg[24]/NET0131  & n46442 ;
  assign n46444 = \P2_P2_EBX_reg[25]/NET0131  & n46443 ;
  assign n46445 = \P2_P2_EBX_reg[26]/NET0131  & n46444 ;
  assign n46447 = \P2_P2_EBX_reg[27]/NET0131  & n46445 ;
  assign n46446 = ~\P2_P2_EBX_reg[27]/NET0131  & ~n46445 ;
  assign n46448 = n26662 & ~n46446 ;
  assign n46449 = ~n46447 & n46448 ;
  assign n46416 = n26578 & n26611 ;
  assign n46417 = ~n26662 & ~n46416 ;
  assign n46418 = \P2_P2_EBX_reg[27]/NET0131  & n46417 ;
  assign n46419 = n44703 & n46416 ;
  assign n46450 = ~n46418 & ~n46419 ;
  assign n46451 = ~n46449 & n46450 ;
  assign n46452 = n26792 & ~n46451 ;
  assign n46453 = \P2_P2_EBX_reg[27]/NET0131  & ~n44508 ;
  assign n46454 = ~n46452 & ~n46453 ;
  assign n46455 = \P2_P2_EBX_reg[31]/NET0131  & ~n44508 ;
  assign n46458 = \P2_P2_EBX_reg[28]/NET0131  & n46447 ;
  assign n46459 = \P2_P2_EBX_reg[29]/NET0131  & n46458 ;
  assign n46460 = \P2_P2_EBX_reg[30]/NET0131  & n46459 ;
  assign n46462 = \P2_P2_EBX_reg[31]/NET0131  & n46460 ;
  assign n46461 = ~\P2_P2_EBX_reg[31]/NET0131  & ~n46460 ;
  assign n46463 = n26662 & ~n46461 ;
  assign n46464 = ~n46462 & n46463 ;
  assign n46456 = n46384 & n46416 ;
  assign n46457 = \P2_P2_EBX_reg[31]/NET0131  & n46417 ;
  assign n46465 = ~n46456 & ~n46457 ;
  assign n46466 = ~n46464 & n46465 ;
  assign n46467 = n26792 & ~n46466 ;
  assign n46468 = ~n46455 & ~n46467 ;
  assign n46469 = \P1_P1_EAX_reg[3]/NET0131  & ~n27551 ;
  assign n46471 = ~n15384 & n24648 ;
  assign n46470 = n22818 & ~n33696 ;
  assign n46472 = ~\P1_P1_EAX_reg[3]/NET0131  & ~n15389 ;
  assign n46473 = ~n15390 & ~n46472 ;
  assign n46474 = n15377 & n46473 ;
  assign n46475 = ~n46470 & ~n46474 ;
  assign n46476 = ~n46471 & n46475 ;
  assign n46477 = n8355 & ~n46476 ;
  assign n46478 = ~n46469 & ~n46477 ;
  assign n46483 = \P1_P3_EBX_reg[2]/NET0131  & n19132 ;
  assign n46484 = \P1_P3_EBX_reg[3]/NET0131  & n46483 ;
  assign n46485 = \P1_P3_EBX_reg[4]/NET0131  & n46484 ;
  assign n46486 = \P1_P3_EBX_reg[5]/NET0131  & n46485 ;
  assign n46487 = \P1_P3_EBX_reg[6]/NET0131  & n46486 ;
  assign n46488 = \P1_P3_EBX_reg[7]/NET0131  & n46487 ;
  assign n46489 = \P1_P3_EBX_reg[8]/NET0131  & n46488 ;
  assign n46490 = \P1_P3_EBX_reg[9]/NET0131  & n46489 ;
  assign n46491 = \P1_P3_EBX_reg[10]/NET0131  & n46490 ;
  assign n46492 = \P1_P3_EBX_reg[11]/NET0131  & n46491 ;
  assign n46493 = \P1_P3_EBX_reg[12]/NET0131  & n46492 ;
  assign n46494 = \P1_P3_EBX_reg[13]/NET0131  & n46493 ;
  assign n46495 = \P1_P3_EBX_reg[14]/NET0131  & n46494 ;
  assign n46496 = \P1_P3_EBX_reg[15]/NET0131  & n46495 ;
  assign n46497 = \P1_P3_EBX_reg[16]/NET0131  & n46496 ;
  assign n46498 = \P1_P3_EBX_reg[17]/NET0131  & n46497 ;
  assign n46499 = \P1_P3_EBX_reg[18]/NET0131  & n46498 ;
  assign n46500 = \P1_P3_EBX_reg[19]/NET0131  & n46499 ;
  assign n46501 = \P1_P3_EBX_reg[20]/NET0131  & n46500 ;
  assign n46502 = \P1_P3_EBX_reg[21]/NET0131  & n46501 ;
  assign n46503 = \P1_P3_EBX_reg[22]/NET0131  & n46502 ;
  assign n46504 = \P1_P3_EBX_reg[23]/NET0131  & n46503 ;
  assign n46505 = \P1_P3_EBX_reg[24]/NET0131  & n46504 ;
  assign n46506 = \P1_P3_EBX_reg[25]/NET0131  & n46505 ;
  assign n46507 = \P1_P3_EBX_reg[26]/NET0131  & n46506 ;
  assign n46509 = \P1_P3_EBX_reg[27]/NET0131  & n46507 ;
  assign n46508 = ~\P1_P3_EBX_reg[27]/NET0131  & ~n46507 ;
  assign n46510 = n9108 & ~n46508 ;
  assign n46511 = ~n46509 & n46510 ;
  assign n46479 = n9049 & n9057 ;
  assign n46480 = ~n9108 & ~n46479 ;
  assign n46481 = \P1_P3_EBX_reg[27]/NET0131  & n46480 ;
  assign n46482 = n22404 & n46479 ;
  assign n46512 = ~n46481 & ~n46482 ;
  assign n46513 = ~n46511 & n46512 ;
  assign n46514 = n9241 & ~n46513 ;
  assign n46515 = \P1_P3_EBX_reg[27]/NET0131  & ~n16968 ;
  assign n46516 = ~n46514 & ~n46515 ;
  assign n46517 = \P1_P3_EBX_reg[31]/NET0131  & ~n16968 ;
  assign n46520 = \P1_P3_EBX_reg[28]/NET0131  & n46509 ;
  assign n46521 = \P1_P3_EBX_reg[29]/NET0131  & n46520 ;
  assign n46522 = \P1_P3_EBX_reg[30]/NET0131  & n46521 ;
  assign n46524 = \P1_P3_EBX_reg[31]/NET0131  & n46522 ;
  assign n46523 = ~\P1_P3_EBX_reg[31]/NET0131  & ~n46522 ;
  assign n46525 = n9108 & ~n46523 ;
  assign n46526 = ~n46524 & n46525 ;
  assign n46518 = \P1_P3_EBX_reg[31]/NET0131  & n46480 ;
  assign n46519 = n21717 & n46479 ;
  assign n46527 = ~n46518 & ~n46519 ;
  assign n46528 = ~n46526 & n46527 ;
  assign n46529 = n9241 & ~n46528 ;
  assign n46530 = ~n46517 & ~n46529 ;
  assign n46537 = \P1_P1_EBX_reg[0]/NET0131  & \P1_P1_EBX_reg[1]/NET0131  ;
  assign n46538 = \P1_P1_EBX_reg[2]/NET0131  & n46537 ;
  assign n46539 = \P1_P1_EBX_reg[3]/NET0131  & n46538 ;
  assign n46540 = \P1_P1_EBX_reg[4]/NET0131  & n46539 ;
  assign n46541 = \P1_P1_EBX_reg[5]/NET0131  & n46540 ;
  assign n46542 = \P1_P1_EBX_reg[6]/NET0131  & n46541 ;
  assign n46543 = \P1_P1_EBX_reg[7]/NET0131  & n46542 ;
  assign n46544 = \P1_P1_EBX_reg[8]/NET0131  & n46543 ;
  assign n46545 = \P1_P1_EBX_reg[9]/NET0131  & n46544 ;
  assign n46546 = \P1_P1_EBX_reg[10]/NET0131  & n46545 ;
  assign n46547 = \P1_P1_EBX_reg[11]/NET0131  & n46546 ;
  assign n46548 = \P1_P1_EBX_reg[12]/NET0131  & n46547 ;
  assign n46549 = \P1_P1_EBX_reg[13]/NET0131  & n46548 ;
  assign n46550 = \P1_P1_EBX_reg[14]/NET0131  & n46549 ;
  assign n46551 = \P1_P1_EBX_reg[15]/NET0131  & n46550 ;
  assign n46552 = \P1_P1_EBX_reg[16]/NET0131  & n46551 ;
  assign n46553 = \P1_P1_EBX_reg[17]/NET0131  & n46552 ;
  assign n46554 = \P1_P1_EBX_reg[18]/NET0131  & n46553 ;
  assign n46555 = \P1_P1_EBX_reg[19]/NET0131  & n46554 ;
  assign n46556 = \P1_P1_EBX_reg[20]/NET0131  & n46555 ;
  assign n46557 = \P1_P1_EBX_reg[21]/NET0131  & n46556 ;
  assign n46558 = \P1_P1_EBX_reg[22]/NET0131  & n46557 ;
  assign n46559 = \P1_P1_EBX_reg[23]/NET0131  & n46558 ;
  assign n46560 = \P1_P1_EBX_reg[24]/NET0131  & n46559 ;
  assign n46561 = \P1_P1_EBX_reg[25]/NET0131  & n46560 ;
  assign n46562 = \P1_P1_EBX_reg[26]/NET0131  & n46561 ;
  assign n46564 = \P1_P1_EBX_reg[27]/NET0131  & n46562 ;
  assign n46563 = ~\P1_P1_EBX_reg[27]/NET0131  & ~n46562 ;
  assign n46565 = n26146 & ~n46563 ;
  assign n46566 = ~n46564 & n46565 ;
  assign n46531 = ~n26122 & ~n26146 ;
  assign n46532 = ~n15428 & n26122 ;
  assign n46533 = ~n46531 & ~n46532 ;
  assign n46534 = \P1_P1_EBX_reg[27]/NET0131  & ~n46533 ;
  assign n46535 = n15428 & n26122 ;
  assign n46536 = n23964 & n46535 ;
  assign n46567 = ~n46534 & ~n46536 ;
  assign n46568 = ~n46566 & n46567 ;
  assign n46569 = n8355 & ~n46568 ;
  assign n46570 = \P1_P1_EBX_reg[27]/NET0131  & ~n15326 ;
  assign n46571 = ~n46569 & ~n46570 ;
  assign n46572 = \P1_P1_EBX_reg[31]/NET0131  & ~n15326 ;
  assign n46575 = \P1_P1_EBX_reg[28]/NET0131  & n46564 ;
  assign n46576 = \P1_P1_EBX_reg[29]/NET0131  & n46575 ;
  assign n46577 = \P1_P1_EBX_reg[30]/NET0131  & n46576 ;
  assign n46579 = \P1_P1_EBX_reg[31]/NET0131  & n46577 ;
  assign n46578 = ~\P1_P1_EBX_reg[31]/NET0131  & ~n46577 ;
  assign n46580 = n26146 & ~n46578 ;
  assign n46581 = ~n46579 & n46580 ;
  assign n46573 = n15716 & n46535 ;
  assign n46574 = \P1_P1_EBX_reg[31]/NET0131  & ~n46533 ;
  assign n46582 = ~n46573 & ~n46574 ;
  assign n46583 = ~n46581 & n46582 ;
  assign n46584 = n8355 & ~n46583 ;
  assign n46585 = ~n46572 & ~n46584 ;
  assign n46586 = \P2_P3_EAX_reg[30]/NET0131  & ~n42872 ;
  assign n46590 = \P2_P3_EAX_reg[26]/NET0131  & \P2_P3_EAX_reg[27]/NET0131  ;
  assign n46591 = \P2_P3_EAX_reg[19]/NET0131  & n42850 ;
  assign n46592 = \P2_P3_EAX_reg[25]/NET0131  & n42853 ;
  assign n46593 = n42852 & n46592 ;
  assign n46594 = n46591 & n46593 ;
  assign n46595 = n46590 & n46594 ;
  assign n46596 = \P2_P3_EAX_reg[28]/NET0131  & n46595 ;
  assign n46597 = \P2_P3_EAX_reg[29]/NET0131  & n46596 ;
  assign n46599 = \P2_P3_EAX_reg[30]/NET0131  & n46597 ;
  assign n46598 = ~\P2_P3_EAX_reg[30]/NET0131  & ~n46597 ;
  assign n46600 = n42539 & ~n46598 ;
  assign n46601 = ~n46599 & n46600 ;
  assign n46605 = \P2_P3_EAX_reg[30]/NET0131  & ~n42543 ;
  assign n46602 = ~n42799 & n42830 ;
  assign n46603 = ~n42831 & ~n46602 ;
  assign n46604 = n42538 & n46603 ;
  assign n46587 = n27122 & ~n27177 ;
  assign n46588 = \P2_buf2_reg[14]/NET0131  & ~n27192 ;
  assign n46589 = n46587 & n46588 ;
  assign n46606 = n27186 & n27227 ;
  assign n46607 = \P2_buf2_reg[30]/NET0131  & n46606 ;
  assign n46608 = ~n46589 & ~n46607 ;
  assign n46609 = ~n46604 & n46608 ;
  assign n46610 = ~n46605 & n46609 ;
  assign n46611 = ~n46601 & n46610 ;
  assign n46612 = n27308 & ~n46611 ;
  assign n46613 = ~n46586 & ~n46612 ;
  assign n46618 = \P2_P3_EBX_reg[0]/NET0131  & \P2_P3_EBX_reg[1]/NET0131  ;
  assign n46619 = \P2_P3_EBX_reg[2]/NET0131  & n46618 ;
  assign n46620 = \P2_P3_EBX_reg[3]/NET0131  & n46619 ;
  assign n46621 = \P2_P3_EBX_reg[4]/NET0131  & n46620 ;
  assign n46622 = \P2_P3_EBX_reg[5]/NET0131  & n46621 ;
  assign n46623 = \P2_P3_EBX_reg[6]/NET0131  & n46622 ;
  assign n46624 = \P2_P3_EBX_reg[7]/NET0131  & n46623 ;
  assign n46625 = \P2_P3_EBX_reg[8]/NET0131  & n46624 ;
  assign n46626 = \P2_P3_EBX_reg[9]/NET0131  & n46625 ;
  assign n46627 = \P2_P3_EBX_reg[10]/NET0131  & n46626 ;
  assign n46628 = \P2_P3_EBX_reg[11]/NET0131  & n46627 ;
  assign n46629 = \P2_P3_EBX_reg[12]/NET0131  & n46628 ;
  assign n46630 = \P2_P3_EBX_reg[13]/NET0131  & n46629 ;
  assign n46631 = \P2_P3_EBX_reg[14]/NET0131  & n46630 ;
  assign n46632 = \P2_P3_EBX_reg[15]/NET0131  & n46631 ;
  assign n46633 = \P2_P3_EBX_reg[16]/NET0131  & n46632 ;
  assign n46634 = \P2_P3_EBX_reg[17]/NET0131  & n46633 ;
  assign n46635 = \P2_P3_EBX_reg[18]/NET0131  & n46634 ;
  assign n46636 = \P2_P3_EBX_reg[19]/NET0131  & n46635 ;
  assign n46637 = \P2_P3_EBX_reg[20]/NET0131  & n46636 ;
  assign n46638 = \P2_P3_EBX_reg[21]/NET0131  & n46637 ;
  assign n46639 = \P2_P3_EBX_reg[22]/NET0131  & n46638 ;
  assign n46640 = \P2_P3_EBX_reg[23]/NET0131  & n46639 ;
  assign n46641 = \P2_P3_EBX_reg[24]/NET0131  & n46640 ;
  assign n46642 = \P2_P3_EBX_reg[25]/NET0131  & n46641 ;
  assign n46643 = \P2_P3_EBX_reg[26]/NET0131  & n46642 ;
  assign n46645 = \P2_P3_EBX_reg[27]/NET0131  & n46643 ;
  assign n46644 = ~\P2_P3_EBX_reg[27]/NET0131  & ~n46643 ;
  assign n46646 = n27133 & ~n46644 ;
  assign n46647 = ~n46645 & n46646 ;
  assign n46614 = n27108 & n27206 ;
  assign n46615 = ~n27133 & ~n46614 ;
  assign n46616 = \P2_P3_EBX_reg[27]/NET0131  & n46615 ;
  assign n46617 = n44790 & n46614 ;
  assign n46648 = ~n46616 & ~n46617 ;
  assign n46649 = ~n46647 & n46648 ;
  assign n46650 = n27308 & ~n46649 ;
  assign n46651 = \P2_P3_EBX_reg[27]/NET0131  & ~n42872 ;
  assign n46652 = ~n46650 & ~n46651 ;
  assign n46655 = \P2_P3_EBX_reg[28]/NET0131  & n46645 ;
  assign n46656 = \P2_P3_EBX_reg[29]/NET0131  & n46655 ;
  assign n46657 = \P2_P3_EBX_reg[30]/NET0131  & n46656 ;
  assign n46659 = \P2_P3_EBX_reg[31]/NET0131  & n46657 ;
  assign n46658 = ~\P2_P3_EBX_reg[31]/NET0131  & ~n46657 ;
  assign n46660 = n27133 & ~n46658 ;
  assign n46661 = ~n46659 & n46660 ;
  assign n46653 = n42831 & n46614 ;
  assign n46654 = \P2_P3_EBX_reg[31]/NET0131  & n46615 ;
  assign n46662 = ~n46653 & ~n46654 ;
  assign n46663 = ~n46661 & n46662 ;
  assign n46664 = n27308 & ~n46663 ;
  assign n46665 = \P2_P3_EBX_reg[31]/NET0131  & ~n42872 ;
  assign n46666 = ~n46664 & ~n46665 ;
  assign n46667 = \P1_P2_EAX_reg[30]/NET0131  & ~n43212 ;
  assign n46668 = n43164 & ~n43199 ;
  assign n46669 = ~n43167 & ~n46668 ;
  assign n46670 = \P1_P2_EAX_reg[30]/NET0131  & ~n46669 ;
  assign n46671 = n43164 & n43198 ;
  assign n46672 = \P1_P2_EAX_reg[29]/NET0131  & ~\P1_P2_EAX_reg[30]/NET0131  ;
  assign n46673 = n46671 & n46672 ;
  assign n46674 = ~n43130 & n43161 ;
  assign n46675 = ~n43162 & ~n46674 ;
  assign n46676 = n42875 & n46675 ;
  assign n46677 = \P1_P2_EAX_reg[30]/NET0131  & ~n25773 ;
  assign n46678 = n25773 & ~n34457 ;
  assign n46679 = ~n46677 & ~n46678 ;
  assign n46680 = n25774 & ~n46679 ;
  assign n46682 = ~\P1_buf1_reg[14]/NET0131  & n27934 ;
  assign n46681 = ~\P1_buf2_reg[14]/NET0131  & ~n27934 ;
  assign n46683 = ~n25415 & ~n46681 ;
  assign n46684 = ~n46682 & n46683 ;
  assign n46685 = ~n25770 & n46684 ;
  assign n46686 = ~n46677 & ~n46685 ;
  assign n46687 = n25776 & ~n46686 ;
  assign n46688 = ~n46680 & ~n46687 ;
  assign n46689 = ~n46676 & n46688 ;
  assign n46690 = ~n46673 & n46689 ;
  assign n46691 = ~n46670 & n46690 ;
  assign n46692 = n25918 & ~n46691 ;
  assign n46693 = ~n46667 & ~n46692 ;
  assign n46698 = \P1_P2_EBX_reg[0]/NET0131  & \P1_P2_EBX_reg[1]/NET0131  ;
  assign n46699 = \P1_P2_EBX_reg[2]/NET0131  & n46698 ;
  assign n46700 = \P1_P2_EBX_reg[3]/NET0131  & n46699 ;
  assign n46701 = \P1_P2_EBX_reg[4]/NET0131  & n46700 ;
  assign n46702 = \P1_P2_EBX_reg[5]/NET0131  & n46701 ;
  assign n46703 = \P1_P2_EBX_reg[6]/NET0131  & n46702 ;
  assign n46704 = \P1_P2_EBX_reg[7]/NET0131  & n46703 ;
  assign n46705 = \P1_P2_EBX_reg[8]/NET0131  & n46704 ;
  assign n46706 = \P1_P2_EBX_reg[9]/NET0131  & n46705 ;
  assign n46707 = \P1_P2_EBX_reg[10]/NET0131  & n46706 ;
  assign n46708 = \P1_P2_EBX_reg[11]/NET0131  & n46707 ;
  assign n46709 = \P1_P2_EBX_reg[12]/NET0131  & n46708 ;
  assign n46710 = \P1_P2_EBX_reg[13]/NET0131  & n46709 ;
  assign n46711 = \P1_P2_EBX_reg[14]/NET0131  & n46710 ;
  assign n46712 = \P1_P2_EBX_reg[15]/NET0131  & n46711 ;
  assign n46713 = \P1_P2_EBX_reg[16]/NET0131  & n46712 ;
  assign n46714 = \P1_P2_EBX_reg[17]/NET0131  & n46713 ;
  assign n46715 = \P1_P2_EBX_reg[18]/NET0131  & n46714 ;
  assign n46716 = \P1_P2_EBX_reg[19]/NET0131  & n46715 ;
  assign n46717 = \P1_P2_EBX_reg[20]/NET0131  & n46716 ;
  assign n46718 = \P1_P2_EBX_reg[21]/NET0131  & n46717 ;
  assign n46719 = \P1_P2_EBX_reg[22]/NET0131  & n46718 ;
  assign n46720 = \P1_P2_EBX_reg[23]/NET0131  & n46719 ;
  assign n46721 = \P1_P2_EBX_reg[24]/NET0131  & n46720 ;
  assign n46722 = \P1_P2_EBX_reg[25]/NET0131  & n46721 ;
  assign n46723 = \P1_P2_EBX_reg[26]/NET0131  & n46722 ;
  assign n46725 = ~\P1_P2_EBX_reg[27]/NET0131  & ~n46723 ;
  assign n46724 = \P1_P2_EBX_reg[27]/NET0131  & n46723 ;
  assign n46726 = n25803 & ~n46724 ;
  assign n46727 = ~n46725 & n46726 ;
  assign n46694 = n25738 & n25747 ;
  assign n46695 = ~n25803 & ~n46694 ;
  assign n46696 = \P1_P2_EBX_reg[27]/NET0131  & n46695 ;
  assign n46697 = n44822 & n46694 ;
  assign n46728 = ~n46696 & ~n46697 ;
  assign n46729 = ~n46727 & n46728 ;
  assign n46730 = n25918 & ~n46729 ;
  assign n46731 = \P1_P2_EBX_reg[27]/NET0131  & ~n43212 ;
  assign n46732 = ~n46730 & ~n46731 ;
  assign n46733 = \P1_P2_EBX_reg[31]/NET0131  & ~n43212 ;
  assign n46736 = \P1_P2_EBX_reg[28]/NET0131  & n46724 ;
  assign n46737 = \P1_P2_EBX_reg[29]/NET0131  & n46736 ;
  assign n46738 = \P1_P2_EBX_reg[30]/NET0131  & n46737 ;
  assign n46740 = \P1_P2_EBX_reg[31]/NET0131  & n46738 ;
  assign n46739 = ~\P1_P2_EBX_reg[31]/NET0131  & ~n46738 ;
  assign n46741 = n25803 & ~n46739 ;
  assign n46742 = ~n46740 & n46741 ;
  assign n46734 = n43162 & n46694 ;
  assign n46735 = \P1_P2_EBX_reg[31]/NET0131  & n46695 ;
  assign n46743 = ~n46734 & ~n46735 ;
  assign n46744 = ~n46742 & n46743 ;
  assign n46745 = n25918 & ~n46744 ;
  assign n46746 = ~n46733 & ~n46745 ;
  assign n46755 = \P1_buf2_reg[24]/NET0131  & ~n27934 ;
  assign n46756 = \P1_buf1_reg[24]/NET0131  & n27934 ;
  assign n46757 = ~n46755 & ~n46756 ;
  assign n46758 = n27945 & ~n46757 ;
  assign n46759 = \P1_buf2_reg[16]/NET0131  & ~n27934 ;
  assign n46760 = \P1_buf1_reg[16]/NET0131  & n27934 ;
  assign n46761 = ~n46759 & ~n46760 ;
  assign n46762 = n27952 & ~n46761 ;
  assign n46763 = ~n46758 & ~n46762 ;
  assign n46764 = \P1_P2_DataWidth_reg[1]/NET0131  & ~n46763 ;
  assign n46747 = \P1_buf2_reg[0]/NET0131  & ~n27934 ;
  assign n46748 = \P1_buf1_reg[0]/NET0131  & n27934 ;
  assign n46749 = ~n46747 & ~n46748 ;
  assign n46750 = ~n27905 & ~n46749 ;
  assign n46751 = \P1_P2_InstQueue_reg[11][0]/NET0131  & ~n27901 ;
  assign n46752 = ~n27904 & n46751 ;
  assign n46753 = ~n46750 & ~n46752 ;
  assign n46765 = ~n27960 & ~n46753 ;
  assign n46766 = ~n46764 & ~n46765 ;
  assign n46767 = n25928 & ~n46766 ;
  assign n46768 = ~n25667 & n27901 ;
  assign n46769 = ~n46751 & ~n46768 ;
  assign n46770 = n27608 & ~n46769 ;
  assign n46754 = n27898 & ~n46753 ;
  assign n46771 = \P1_P2_InstQueue_reg[11][0]/NET0131  & ~n27972 ;
  assign n46772 = ~n46754 & ~n46771 ;
  assign n46773 = ~n46770 & n46772 ;
  assign n46774 = ~n46767 & n46773 ;
  assign n46786 = \P2_buf2_reg[24]/NET0131  & ~n28013 ;
  assign n46787 = \P2_buf1_reg[24]/NET0131  & n28013 ;
  assign n46788 = ~n46786 & ~n46787 ;
  assign n46789 = n28027 & ~n46788 ;
  assign n46790 = \P2_buf2_reg[16]/NET0131  & ~n28013 ;
  assign n46791 = \P2_buf1_reg[16]/NET0131  & n28013 ;
  assign n46792 = ~n46790 & ~n46791 ;
  assign n46793 = n28034 & ~n46792 ;
  assign n46794 = ~n46789 & ~n46793 ;
  assign n46795 = \P2_P2_DataWidth_reg[1]/NET0131  & ~n46794 ;
  assign n46775 = \P2_buf2_reg[0]/NET0131  & ~n28013 ;
  assign n46776 = \P2_buf1_reg[0]/NET0131  & n28013 ;
  assign n46777 = ~n46775 & ~n46776 ;
  assign n46778 = ~n27984 & ~n46777 ;
  assign n46779 = \P2_P2_InstQueue_reg[11][0]/NET0131  & ~n27980 ;
  assign n46780 = ~n27983 & n46779 ;
  assign n46781 = ~n46778 & ~n46780 ;
  assign n46796 = ~n28042 & ~n46781 ;
  assign n46797 = ~n46795 & ~n46796 ;
  assign n46798 = n26794 & ~n46797 ;
  assign n46783 = ~n26544 & n27980 ;
  assign n46784 = ~n46779 & ~n46783 ;
  assign n46785 = n27613 & ~n46784 ;
  assign n46782 = n27977 & ~n46781 ;
  assign n46799 = \P2_P2_InstQueue_reg[11][0]/NET0131  & ~n28050 ;
  assign n46800 = ~n46782 & ~n46799 ;
  assign n46801 = ~n46785 & n46800 ;
  assign n46802 = ~n46798 & n46801 ;
  assign n46808 = n28065 & ~n46757 ;
  assign n46809 = n28068 & ~n46761 ;
  assign n46810 = ~n46808 & ~n46809 ;
  assign n46811 = \P1_P2_DataWidth_reg[1]/NET0131  & ~n46810 ;
  assign n46803 = ~n28058 & ~n46749 ;
  assign n46804 = \P1_P2_InstQueue_reg[0][0]/NET0131  & ~n28055 ;
  assign n46805 = ~n28057 & n46804 ;
  assign n46806 = ~n46803 & ~n46805 ;
  assign n46812 = ~n28073 & ~n46806 ;
  assign n46813 = ~n46811 & ~n46812 ;
  assign n46814 = n25928 & ~n46813 ;
  assign n46815 = ~n25667 & n28055 ;
  assign n46816 = ~n46804 & ~n46815 ;
  assign n46817 = n27608 & ~n46816 ;
  assign n46807 = n27898 & ~n46806 ;
  assign n46818 = \P1_P2_InstQueue_reg[0][0]/NET0131  & ~n27972 ;
  assign n46819 = ~n46807 & ~n46818 ;
  assign n46820 = ~n46817 & n46819 ;
  assign n46821 = ~n46814 & n46820 ;
  assign n46827 = n28090 & ~n46757 ;
  assign n46828 = n27945 & ~n46761 ;
  assign n46829 = ~n46827 & ~n46828 ;
  assign n46830 = \P1_P2_DataWidth_reg[1]/NET0131  & ~n46829 ;
  assign n46822 = ~n28084 & ~n46749 ;
  assign n46823 = \P1_P2_InstQueue_reg[10][0]/NET0131  & ~n27904 ;
  assign n46824 = ~n27952 & n46823 ;
  assign n46825 = ~n46822 & ~n46824 ;
  assign n46831 = ~n28096 & ~n46825 ;
  assign n46832 = ~n46830 & ~n46831 ;
  assign n46833 = n25928 & ~n46832 ;
  assign n46834 = ~n25667 & n27904 ;
  assign n46835 = ~n46823 & ~n46834 ;
  assign n46836 = n27608 & ~n46835 ;
  assign n46826 = n27898 & ~n46825 ;
  assign n46837 = \P1_P2_InstQueue_reg[10][0]/NET0131  & ~n27972 ;
  assign n46838 = ~n46826 & ~n46837 ;
  assign n46839 = ~n46836 & n46838 ;
  assign n46840 = ~n46833 & n46839 ;
  assign n46846 = n27952 & ~n46757 ;
  assign n46847 = n27904 & ~n46761 ;
  assign n46848 = ~n46846 & ~n46847 ;
  assign n46849 = \P1_P2_DataWidth_reg[1]/NET0131  & ~n46848 ;
  assign n46841 = ~n28109 & ~n46749 ;
  assign n46842 = \P1_P2_InstQueue_reg[12][0]/NET0131  & ~n28108 ;
  assign n46843 = ~n27901 & n46842 ;
  assign n46844 = ~n46841 & ~n46843 ;
  assign n46850 = ~n28119 & ~n46844 ;
  assign n46851 = ~n46849 & ~n46850 ;
  assign n46852 = n25928 & ~n46851 ;
  assign n46853 = ~n25667 & n28108 ;
  assign n46854 = ~n46842 & ~n46853 ;
  assign n46855 = n27608 & ~n46854 ;
  assign n46845 = n27898 & ~n46844 ;
  assign n46856 = \P1_P2_InstQueue_reg[12][0]/NET0131  & ~n27972 ;
  assign n46857 = ~n46845 & ~n46856 ;
  assign n46858 = ~n46855 & n46857 ;
  assign n46859 = ~n46852 & n46858 ;
  assign n46865 = n27904 & ~n46757 ;
  assign n46866 = n27901 & ~n46761 ;
  assign n46867 = ~n46865 & ~n46866 ;
  assign n46868 = \P1_P2_DataWidth_reg[1]/NET0131  & ~n46867 ;
  assign n46860 = ~n28130 & ~n46749 ;
  assign n46861 = \P1_P2_InstQueue_reg[13][0]/NET0131  & ~n28065 ;
  assign n46862 = ~n28108 & n46861 ;
  assign n46863 = ~n46860 & ~n46862 ;
  assign n46869 = ~n28140 & ~n46863 ;
  assign n46870 = ~n46868 & ~n46869 ;
  assign n46871 = n25928 & ~n46870 ;
  assign n46872 = ~n25667 & n28065 ;
  assign n46873 = ~n46861 & ~n46872 ;
  assign n46874 = n27608 & ~n46873 ;
  assign n46864 = n27898 & ~n46863 ;
  assign n46875 = \P1_P2_InstQueue_reg[13][0]/NET0131  & ~n27972 ;
  assign n46876 = ~n46864 & ~n46875 ;
  assign n46877 = ~n46874 & n46876 ;
  assign n46878 = ~n46871 & n46877 ;
  assign n46884 = n27901 & ~n46757 ;
  assign n46885 = n28108 & ~n46761 ;
  assign n46886 = ~n46884 & ~n46885 ;
  assign n46887 = \P1_P2_DataWidth_reg[1]/NET0131  & ~n46886 ;
  assign n46879 = ~n28072 & ~n46749 ;
  assign n46880 = \P1_P2_InstQueue_reg[14][0]/NET0131  & ~n28068 ;
  assign n46881 = ~n28065 & n46880 ;
  assign n46882 = ~n46879 & ~n46881 ;
  assign n46888 = ~n28160 & ~n46882 ;
  assign n46889 = ~n46887 & ~n46888 ;
  assign n46890 = n25928 & ~n46889 ;
  assign n46891 = ~n25667 & n28068 ;
  assign n46892 = ~n46880 & ~n46891 ;
  assign n46893 = n27608 & ~n46892 ;
  assign n46883 = n27898 & ~n46882 ;
  assign n46894 = \P1_P2_InstQueue_reg[14][0]/NET0131  & ~n27972 ;
  assign n46895 = ~n46883 & ~n46894 ;
  assign n46896 = ~n46893 & n46895 ;
  assign n46897 = ~n46890 & n46896 ;
  assign n46903 = n28108 & ~n46757 ;
  assign n46904 = n28065 & ~n46761 ;
  assign n46905 = ~n46903 & ~n46904 ;
  assign n46906 = \P1_P2_DataWidth_reg[1]/NET0131  & ~n46905 ;
  assign n46898 = ~n28171 & ~n46749 ;
  assign n46899 = \P1_P2_InstQueue_reg[15][0]/NET0131  & ~n28057 ;
  assign n46900 = ~n28068 & n46899 ;
  assign n46901 = ~n46898 & ~n46900 ;
  assign n46907 = ~n28181 & ~n46901 ;
  assign n46908 = ~n46906 & ~n46907 ;
  assign n46909 = n25928 & ~n46908 ;
  assign n46910 = ~n25667 & n28057 ;
  assign n46911 = ~n46899 & ~n46910 ;
  assign n46912 = n27608 & ~n46911 ;
  assign n46902 = n27898 & ~n46901 ;
  assign n46913 = \P1_P2_InstQueue_reg[15][0]/NET0131  & ~n27972 ;
  assign n46914 = ~n46902 & ~n46913 ;
  assign n46915 = ~n46912 & n46914 ;
  assign n46916 = ~n46909 & n46915 ;
  assign n46922 = n28068 & ~n46757 ;
  assign n46923 = n28057 & ~n46761 ;
  assign n46924 = ~n46922 & ~n46923 ;
  assign n46925 = \P1_P2_DataWidth_reg[1]/NET0131  & ~n46924 ;
  assign n46917 = ~n28193 & ~n46749 ;
  assign n46918 = \P1_P2_InstQueue_reg[1][0]/NET0131  & ~n28192 ;
  assign n46919 = ~n28055 & n46918 ;
  assign n46920 = ~n46917 & ~n46919 ;
  assign n46926 = ~n28203 & ~n46920 ;
  assign n46927 = ~n46925 & ~n46926 ;
  assign n46928 = n25928 & ~n46927 ;
  assign n46929 = ~n25667 & n28192 ;
  assign n46930 = ~n46918 & ~n46929 ;
  assign n46931 = n27608 & ~n46930 ;
  assign n46921 = n27898 & ~n46920 ;
  assign n46932 = \P1_P2_InstQueue_reg[1][0]/NET0131  & ~n27972 ;
  assign n46933 = ~n46921 & ~n46932 ;
  assign n46934 = ~n46931 & n46933 ;
  assign n46935 = ~n46928 & n46934 ;
  assign n46941 = n28057 & ~n46757 ;
  assign n46942 = n28055 & ~n46761 ;
  assign n46943 = ~n46941 & ~n46942 ;
  assign n46944 = \P1_P2_DataWidth_reg[1]/NET0131  & ~n46943 ;
  assign n46936 = ~n28215 & ~n46749 ;
  assign n46937 = \P1_P2_InstQueue_reg[2][0]/NET0131  & ~n28214 ;
  assign n46938 = ~n28192 & n46937 ;
  assign n46939 = ~n46936 & ~n46938 ;
  assign n46945 = ~n28225 & ~n46939 ;
  assign n46946 = ~n46944 & ~n46945 ;
  assign n46947 = n25928 & ~n46946 ;
  assign n46948 = ~n25667 & n28214 ;
  assign n46949 = ~n46937 & ~n46948 ;
  assign n46950 = n27608 & ~n46949 ;
  assign n46940 = n27898 & ~n46939 ;
  assign n46951 = \P1_P2_InstQueue_reg[2][0]/NET0131  & ~n27972 ;
  assign n46952 = ~n46940 & ~n46951 ;
  assign n46953 = ~n46950 & n46952 ;
  assign n46954 = ~n46947 & n46953 ;
  assign n46960 = n28055 & ~n46757 ;
  assign n46961 = n28192 & ~n46761 ;
  assign n46962 = ~n46960 & ~n46961 ;
  assign n46963 = \P1_P2_DataWidth_reg[1]/NET0131  & ~n46962 ;
  assign n46955 = ~n28237 & ~n46749 ;
  assign n46956 = \P1_P2_InstQueue_reg[3][0]/NET0131  & ~n28236 ;
  assign n46957 = ~n28214 & n46956 ;
  assign n46958 = ~n46955 & ~n46957 ;
  assign n46964 = ~n28247 & ~n46958 ;
  assign n46965 = ~n46963 & ~n46964 ;
  assign n46966 = n25928 & ~n46965 ;
  assign n46967 = ~n25667 & n28236 ;
  assign n46968 = ~n46956 & ~n46967 ;
  assign n46969 = n27608 & ~n46968 ;
  assign n46959 = n27898 & ~n46958 ;
  assign n46970 = \P1_P2_InstQueue_reg[3][0]/NET0131  & ~n27972 ;
  assign n46971 = ~n46959 & ~n46970 ;
  assign n46972 = ~n46969 & n46971 ;
  assign n46973 = ~n46966 & n46972 ;
  assign n46979 = n28192 & ~n46757 ;
  assign n46980 = n28214 & ~n46761 ;
  assign n46981 = ~n46979 & ~n46980 ;
  assign n46982 = \P1_P2_DataWidth_reg[1]/NET0131  & ~n46981 ;
  assign n46974 = ~n28259 & ~n46749 ;
  assign n46975 = \P1_P2_InstQueue_reg[4][0]/NET0131  & ~n28258 ;
  assign n46976 = ~n28236 & n46975 ;
  assign n46977 = ~n46974 & ~n46976 ;
  assign n46983 = ~n28269 & ~n46977 ;
  assign n46984 = ~n46982 & ~n46983 ;
  assign n46985 = n25928 & ~n46984 ;
  assign n46986 = ~n25667 & n28258 ;
  assign n46987 = ~n46975 & ~n46986 ;
  assign n46988 = n27608 & ~n46987 ;
  assign n46978 = n27898 & ~n46977 ;
  assign n46989 = \P1_P2_InstQueue_reg[4][0]/NET0131  & ~n27972 ;
  assign n46990 = ~n46978 & ~n46989 ;
  assign n46991 = ~n46988 & n46990 ;
  assign n46992 = ~n46985 & n46991 ;
  assign n46998 = n28214 & ~n46757 ;
  assign n46999 = n28236 & ~n46761 ;
  assign n47000 = ~n46998 & ~n46999 ;
  assign n47001 = \P1_P2_DataWidth_reg[1]/NET0131  & ~n47000 ;
  assign n46993 = ~n28281 & ~n46749 ;
  assign n46994 = \P1_P2_InstQueue_reg[5][0]/NET0131  & ~n28280 ;
  assign n46995 = ~n28258 & n46994 ;
  assign n46996 = ~n46993 & ~n46995 ;
  assign n47002 = ~n28291 & ~n46996 ;
  assign n47003 = ~n47001 & ~n47002 ;
  assign n47004 = n25928 & ~n47003 ;
  assign n47005 = ~n25667 & n28280 ;
  assign n47006 = ~n46994 & ~n47005 ;
  assign n47007 = n27608 & ~n47006 ;
  assign n46997 = n27898 & ~n46996 ;
  assign n47008 = \P1_P2_InstQueue_reg[5][0]/NET0131  & ~n27972 ;
  assign n47009 = ~n46997 & ~n47008 ;
  assign n47010 = ~n47007 & n47009 ;
  assign n47011 = ~n47004 & n47010 ;
  assign n47017 = n28236 & ~n46757 ;
  assign n47018 = n28258 & ~n46761 ;
  assign n47019 = ~n47017 & ~n47018 ;
  assign n47020 = \P1_P2_DataWidth_reg[1]/NET0131  & ~n47019 ;
  assign n47012 = ~n28303 & ~n46749 ;
  assign n47013 = \P1_P2_InstQueue_reg[6][0]/NET0131  & ~n28302 ;
  assign n47014 = ~n28280 & n47013 ;
  assign n47015 = ~n47012 & ~n47014 ;
  assign n47021 = ~n28313 & ~n47015 ;
  assign n47022 = ~n47020 & ~n47021 ;
  assign n47023 = n25928 & ~n47022 ;
  assign n47024 = ~n25667 & n28302 ;
  assign n47025 = ~n47013 & ~n47024 ;
  assign n47026 = n27608 & ~n47025 ;
  assign n47016 = n27898 & ~n47015 ;
  assign n47027 = \P1_P2_InstQueue_reg[6][0]/NET0131  & ~n27972 ;
  assign n47028 = ~n47016 & ~n47027 ;
  assign n47029 = ~n47026 & n47028 ;
  assign n47030 = ~n47023 & n47029 ;
  assign n47036 = n28258 & ~n46757 ;
  assign n47037 = n28280 & ~n46761 ;
  assign n47038 = ~n47036 & ~n47037 ;
  assign n47039 = \P1_P2_DataWidth_reg[1]/NET0131  & ~n47038 ;
  assign n47031 = ~n28324 & ~n46749 ;
  assign n47032 = \P1_P2_InstQueue_reg[7][0]/NET0131  & ~n28090 ;
  assign n47033 = ~n28302 & n47032 ;
  assign n47034 = ~n47031 & ~n47033 ;
  assign n47040 = ~n28334 & ~n47034 ;
  assign n47041 = ~n47039 & ~n47040 ;
  assign n47042 = n25928 & ~n47041 ;
  assign n47043 = ~n25667 & n28090 ;
  assign n47044 = ~n47032 & ~n47043 ;
  assign n47045 = n27608 & ~n47044 ;
  assign n47035 = n27898 & ~n47034 ;
  assign n47046 = \P1_P2_InstQueue_reg[7][0]/NET0131  & ~n27972 ;
  assign n47047 = ~n47035 & ~n47046 ;
  assign n47048 = ~n47045 & n47047 ;
  assign n47049 = ~n47042 & n47048 ;
  assign n47055 = n28280 & ~n46757 ;
  assign n47056 = n28302 & ~n46761 ;
  assign n47057 = ~n47055 & ~n47056 ;
  assign n47058 = \P1_P2_DataWidth_reg[1]/NET0131  & ~n47057 ;
  assign n47050 = ~n28095 & ~n46749 ;
  assign n47051 = \P1_P2_InstQueue_reg[8][0]/NET0131  & ~n27945 ;
  assign n47052 = ~n28090 & n47051 ;
  assign n47053 = ~n47050 & ~n47052 ;
  assign n47059 = ~n28354 & ~n47053 ;
  assign n47060 = ~n47058 & ~n47059 ;
  assign n47061 = n25928 & ~n47060 ;
  assign n47062 = ~n25667 & n27945 ;
  assign n47063 = ~n47051 & ~n47062 ;
  assign n47064 = n27608 & ~n47063 ;
  assign n47054 = n27898 & ~n47053 ;
  assign n47065 = \P1_P2_InstQueue_reg[8][0]/NET0131  & ~n27972 ;
  assign n47066 = ~n47054 & ~n47065 ;
  assign n47067 = ~n47064 & n47066 ;
  assign n47068 = ~n47061 & n47067 ;
  assign n47074 = n28302 & ~n46757 ;
  assign n47075 = n28090 & ~n46761 ;
  assign n47076 = ~n47074 & ~n47075 ;
  assign n47077 = \P1_P2_DataWidth_reg[1]/NET0131  & ~n47076 ;
  assign n47069 = ~n27959 & ~n46749 ;
  assign n47070 = \P1_P2_InstQueue_reg[9][0]/NET0131  & ~n27952 ;
  assign n47071 = ~n27945 & n47070 ;
  assign n47072 = ~n47069 & ~n47071 ;
  assign n47078 = ~n28374 & ~n47072 ;
  assign n47079 = ~n47077 & ~n47078 ;
  assign n47080 = n25928 & ~n47079 ;
  assign n47081 = ~n25667 & n27952 ;
  assign n47082 = ~n47070 & ~n47081 ;
  assign n47083 = n27608 & ~n47082 ;
  assign n47073 = n27898 & ~n47072 ;
  assign n47084 = \P1_P2_InstQueue_reg[9][0]/NET0131  & ~n27972 ;
  assign n47085 = ~n47073 & ~n47084 ;
  assign n47086 = ~n47083 & n47085 ;
  assign n47087 = ~n47080 & n47086 ;
  assign n47096 = n28398 & ~n46788 ;
  assign n47097 = n28401 & ~n46792 ;
  assign n47098 = ~n47096 & ~n47097 ;
  assign n47099 = \P2_P2_DataWidth_reg[1]/NET0131  & ~n47098 ;
  assign n47088 = ~n28388 & ~n46777 ;
  assign n47089 = \P2_P2_InstQueue_reg[0][0]/NET0131  & ~n28385 ;
  assign n47090 = ~n28387 & n47089 ;
  assign n47091 = ~n47088 & ~n47090 ;
  assign n47100 = ~n28406 & ~n47091 ;
  assign n47101 = ~n47099 & ~n47100 ;
  assign n47102 = n26794 & ~n47101 ;
  assign n47093 = ~n26544 & n28385 ;
  assign n47094 = ~n47089 & ~n47093 ;
  assign n47095 = n27613 & ~n47094 ;
  assign n47092 = n27977 & ~n47091 ;
  assign n47103 = \P2_P2_InstQueue_reg[0][0]/NET0131  & ~n28050 ;
  assign n47104 = ~n47092 & ~n47103 ;
  assign n47105 = ~n47095 & n47104 ;
  assign n47106 = ~n47102 & n47105 ;
  assign n47115 = n28423 & ~n46788 ;
  assign n47116 = n28027 & ~n46792 ;
  assign n47117 = ~n47115 & ~n47116 ;
  assign n47118 = \P2_P2_DataWidth_reg[1]/NET0131  & ~n47117 ;
  assign n47107 = ~n28414 & ~n46777 ;
  assign n47108 = \P2_P2_InstQueue_reg[10][0]/NET0131  & ~n27983 ;
  assign n47109 = ~n28034 & n47108 ;
  assign n47110 = ~n47107 & ~n47109 ;
  assign n47119 = ~n28429 & ~n47110 ;
  assign n47120 = ~n47118 & ~n47119 ;
  assign n47121 = n26794 & ~n47120 ;
  assign n47112 = ~n26544 & n27983 ;
  assign n47113 = ~n47108 & ~n47112 ;
  assign n47114 = n27613 & ~n47113 ;
  assign n47111 = n27977 & ~n47110 ;
  assign n47122 = \P2_P2_InstQueue_reg[10][0]/NET0131  & ~n28050 ;
  assign n47123 = ~n47111 & ~n47122 ;
  assign n47124 = ~n47114 & n47123 ;
  assign n47125 = ~n47121 & n47124 ;
  assign n47134 = n28034 & ~n46788 ;
  assign n47135 = n27983 & ~n46792 ;
  assign n47136 = ~n47134 & ~n47135 ;
  assign n47137 = \P2_P2_DataWidth_reg[1]/NET0131  & ~n47136 ;
  assign n47126 = ~n28439 & ~n46777 ;
  assign n47127 = \P2_P2_InstQueue_reg[12][0]/NET0131  & ~n28438 ;
  assign n47128 = ~n27980 & n47127 ;
  assign n47129 = ~n47126 & ~n47128 ;
  assign n47138 = ~n28452 & ~n47129 ;
  assign n47139 = ~n47137 & ~n47138 ;
  assign n47140 = n26794 & ~n47139 ;
  assign n47131 = ~n26544 & n28438 ;
  assign n47132 = ~n47127 & ~n47131 ;
  assign n47133 = n27613 & ~n47132 ;
  assign n47130 = n27977 & ~n47129 ;
  assign n47141 = \P2_P2_InstQueue_reg[12][0]/NET0131  & ~n28050 ;
  assign n47142 = ~n47130 & ~n47141 ;
  assign n47143 = ~n47133 & n47142 ;
  assign n47144 = ~n47140 & n47143 ;
  assign n47153 = n27983 & ~n46788 ;
  assign n47154 = n27980 & ~n46792 ;
  assign n47155 = ~n47153 & ~n47154 ;
  assign n47156 = \P2_P2_DataWidth_reg[1]/NET0131  & ~n47155 ;
  assign n47145 = ~n28460 & ~n46777 ;
  assign n47146 = \P2_P2_InstQueue_reg[13][0]/NET0131  & ~n28398 ;
  assign n47147 = ~n28438 & n47146 ;
  assign n47148 = ~n47145 & ~n47147 ;
  assign n47157 = ~n28473 & ~n47148 ;
  assign n47158 = ~n47156 & ~n47157 ;
  assign n47159 = n26794 & ~n47158 ;
  assign n47150 = ~n26544 & n28398 ;
  assign n47151 = ~n47146 & ~n47150 ;
  assign n47152 = n27613 & ~n47151 ;
  assign n47149 = n27977 & ~n47148 ;
  assign n47160 = \P2_P2_InstQueue_reg[13][0]/NET0131  & ~n28050 ;
  assign n47161 = ~n47149 & ~n47160 ;
  assign n47162 = ~n47152 & n47161 ;
  assign n47163 = ~n47159 & n47162 ;
  assign n47172 = n27980 & ~n46788 ;
  assign n47173 = n28438 & ~n46792 ;
  assign n47174 = ~n47172 & ~n47173 ;
  assign n47175 = \P2_P2_DataWidth_reg[1]/NET0131  & ~n47174 ;
  assign n47164 = ~n28405 & ~n46777 ;
  assign n47165 = \P2_P2_InstQueue_reg[14][0]/NET0131  & ~n28401 ;
  assign n47166 = ~n28398 & n47165 ;
  assign n47167 = ~n47164 & ~n47166 ;
  assign n47176 = ~n28493 & ~n47167 ;
  assign n47177 = ~n47175 & ~n47176 ;
  assign n47178 = n26794 & ~n47177 ;
  assign n47169 = ~n26544 & n28401 ;
  assign n47170 = ~n47165 & ~n47169 ;
  assign n47171 = n27613 & ~n47170 ;
  assign n47168 = n27977 & ~n47167 ;
  assign n47179 = \P2_P2_InstQueue_reg[14][0]/NET0131  & ~n28050 ;
  assign n47180 = ~n47168 & ~n47179 ;
  assign n47181 = ~n47171 & n47180 ;
  assign n47182 = ~n47178 & n47181 ;
  assign n47191 = n28438 & ~n46788 ;
  assign n47192 = n28398 & ~n46792 ;
  assign n47193 = ~n47191 & ~n47192 ;
  assign n47194 = \P2_P2_DataWidth_reg[1]/NET0131  & ~n47193 ;
  assign n47183 = ~n28501 & ~n46777 ;
  assign n47184 = \P2_P2_InstQueue_reg[15][0]/NET0131  & ~n28387 ;
  assign n47185 = ~n28401 & n47184 ;
  assign n47186 = ~n47183 & ~n47185 ;
  assign n47195 = ~n28514 & ~n47186 ;
  assign n47196 = ~n47194 & ~n47195 ;
  assign n47197 = n26794 & ~n47196 ;
  assign n47188 = ~n26544 & n28387 ;
  assign n47189 = ~n47184 & ~n47188 ;
  assign n47190 = n27613 & ~n47189 ;
  assign n47187 = n27977 & ~n47186 ;
  assign n47198 = \P2_P2_InstQueue_reg[15][0]/NET0131  & ~n28050 ;
  assign n47199 = ~n47187 & ~n47198 ;
  assign n47200 = ~n47190 & n47199 ;
  assign n47201 = ~n47197 & n47200 ;
  assign n47210 = n28401 & ~n46788 ;
  assign n47211 = n28387 & ~n46792 ;
  assign n47212 = ~n47210 & ~n47211 ;
  assign n47213 = \P2_P2_DataWidth_reg[1]/NET0131  & ~n47212 ;
  assign n47202 = ~n28523 & ~n46777 ;
  assign n47203 = \P2_P2_InstQueue_reg[1][0]/NET0131  & ~n28522 ;
  assign n47204 = ~n28385 & n47203 ;
  assign n47205 = ~n47202 & ~n47204 ;
  assign n47214 = ~n28536 & ~n47205 ;
  assign n47215 = ~n47213 & ~n47214 ;
  assign n47216 = n26794 & ~n47215 ;
  assign n47207 = ~n26544 & n28522 ;
  assign n47208 = ~n47203 & ~n47207 ;
  assign n47209 = n27613 & ~n47208 ;
  assign n47206 = n27977 & ~n47205 ;
  assign n47217 = \P2_P2_InstQueue_reg[1][0]/NET0131  & ~n28050 ;
  assign n47218 = ~n47206 & ~n47217 ;
  assign n47219 = ~n47209 & n47218 ;
  assign n47220 = ~n47216 & n47219 ;
  assign n47229 = n28387 & ~n46788 ;
  assign n47230 = n28385 & ~n46792 ;
  assign n47231 = ~n47229 & ~n47230 ;
  assign n47232 = \P2_P2_DataWidth_reg[1]/NET0131  & ~n47231 ;
  assign n47221 = ~n28545 & ~n46777 ;
  assign n47222 = \P2_P2_InstQueue_reg[2][0]/NET0131  & ~n28544 ;
  assign n47223 = ~n28522 & n47222 ;
  assign n47224 = ~n47221 & ~n47223 ;
  assign n47233 = ~n28558 & ~n47224 ;
  assign n47234 = ~n47232 & ~n47233 ;
  assign n47235 = n26794 & ~n47234 ;
  assign n47226 = ~n26544 & n28544 ;
  assign n47227 = ~n47222 & ~n47226 ;
  assign n47228 = n27613 & ~n47227 ;
  assign n47225 = n27977 & ~n47224 ;
  assign n47236 = \P2_P2_InstQueue_reg[2][0]/NET0131  & ~n28050 ;
  assign n47237 = ~n47225 & ~n47236 ;
  assign n47238 = ~n47228 & n47237 ;
  assign n47239 = ~n47235 & n47238 ;
  assign n47248 = n28385 & ~n46788 ;
  assign n47249 = n28522 & ~n46792 ;
  assign n47250 = ~n47248 & ~n47249 ;
  assign n47251 = \P2_P2_DataWidth_reg[1]/NET0131  & ~n47250 ;
  assign n47240 = ~n28567 & ~n46777 ;
  assign n47241 = \P2_P2_InstQueue_reg[3][0]/NET0131  & ~n28566 ;
  assign n47242 = ~n28544 & n47241 ;
  assign n47243 = ~n47240 & ~n47242 ;
  assign n47252 = ~n28580 & ~n47243 ;
  assign n47253 = ~n47251 & ~n47252 ;
  assign n47254 = n26794 & ~n47253 ;
  assign n47245 = ~n26544 & n28566 ;
  assign n47246 = ~n47241 & ~n47245 ;
  assign n47247 = n27613 & ~n47246 ;
  assign n47244 = n27977 & ~n47243 ;
  assign n47255 = \P2_P2_InstQueue_reg[3][0]/NET0131  & ~n28050 ;
  assign n47256 = ~n47244 & ~n47255 ;
  assign n47257 = ~n47247 & n47256 ;
  assign n47258 = ~n47254 & n47257 ;
  assign n47267 = n28522 & ~n46788 ;
  assign n47268 = n28544 & ~n46792 ;
  assign n47269 = ~n47267 & ~n47268 ;
  assign n47270 = \P2_P2_DataWidth_reg[1]/NET0131  & ~n47269 ;
  assign n47259 = ~n28589 & ~n46777 ;
  assign n47260 = \P2_P2_InstQueue_reg[4][0]/NET0131  & ~n28588 ;
  assign n47261 = ~n28566 & n47260 ;
  assign n47262 = ~n47259 & ~n47261 ;
  assign n47271 = ~n28602 & ~n47262 ;
  assign n47272 = ~n47270 & ~n47271 ;
  assign n47273 = n26794 & ~n47272 ;
  assign n47264 = ~n26544 & n28588 ;
  assign n47265 = ~n47260 & ~n47264 ;
  assign n47266 = n27613 & ~n47265 ;
  assign n47263 = n27977 & ~n47262 ;
  assign n47274 = \P2_P2_InstQueue_reg[4][0]/NET0131  & ~n28050 ;
  assign n47275 = ~n47263 & ~n47274 ;
  assign n47276 = ~n47266 & n47275 ;
  assign n47277 = ~n47273 & n47276 ;
  assign n47286 = n28544 & ~n46788 ;
  assign n47287 = n28566 & ~n46792 ;
  assign n47288 = ~n47286 & ~n47287 ;
  assign n47289 = \P2_P2_DataWidth_reg[1]/NET0131  & ~n47288 ;
  assign n47278 = ~n28611 & ~n46777 ;
  assign n47279 = \P2_P2_InstQueue_reg[5][0]/NET0131  & ~n28610 ;
  assign n47280 = ~n28588 & n47279 ;
  assign n47281 = ~n47278 & ~n47280 ;
  assign n47290 = ~n28624 & ~n47281 ;
  assign n47291 = ~n47289 & ~n47290 ;
  assign n47292 = n26794 & ~n47291 ;
  assign n47283 = ~n26544 & n28610 ;
  assign n47284 = ~n47279 & ~n47283 ;
  assign n47285 = n27613 & ~n47284 ;
  assign n47282 = n27977 & ~n47281 ;
  assign n47293 = \P2_P2_InstQueue_reg[5][0]/NET0131  & ~n28050 ;
  assign n47294 = ~n47282 & ~n47293 ;
  assign n47295 = ~n47285 & n47294 ;
  assign n47296 = ~n47292 & n47295 ;
  assign n47305 = n28566 & ~n46788 ;
  assign n47306 = n28588 & ~n46792 ;
  assign n47307 = ~n47305 & ~n47306 ;
  assign n47308 = \P2_P2_DataWidth_reg[1]/NET0131  & ~n47307 ;
  assign n47297 = ~n28633 & ~n46777 ;
  assign n47298 = \P2_P2_InstQueue_reg[6][0]/NET0131  & ~n28632 ;
  assign n47299 = ~n28610 & n47298 ;
  assign n47300 = ~n47297 & ~n47299 ;
  assign n47309 = ~n28646 & ~n47300 ;
  assign n47310 = ~n47308 & ~n47309 ;
  assign n47311 = n26794 & ~n47310 ;
  assign n47302 = ~n26544 & n28632 ;
  assign n47303 = ~n47298 & ~n47302 ;
  assign n47304 = n27613 & ~n47303 ;
  assign n47301 = n27977 & ~n47300 ;
  assign n47312 = \P2_P2_InstQueue_reg[6][0]/NET0131  & ~n28050 ;
  assign n47313 = ~n47301 & ~n47312 ;
  assign n47314 = ~n47304 & n47313 ;
  assign n47315 = ~n47311 & n47314 ;
  assign n47324 = n28588 & ~n46788 ;
  assign n47325 = n28610 & ~n46792 ;
  assign n47326 = ~n47324 & ~n47325 ;
  assign n47327 = \P2_P2_DataWidth_reg[1]/NET0131  & ~n47326 ;
  assign n47316 = ~n28654 & ~n46777 ;
  assign n47317 = \P2_P2_InstQueue_reg[7][0]/NET0131  & ~n28423 ;
  assign n47318 = ~n28632 & n47317 ;
  assign n47319 = ~n47316 & ~n47318 ;
  assign n47328 = ~n28667 & ~n47319 ;
  assign n47329 = ~n47327 & ~n47328 ;
  assign n47330 = n26794 & ~n47329 ;
  assign n47321 = ~n26544 & n28423 ;
  assign n47322 = ~n47317 & ~n47321 ;
  assign n47323 = n27613 & ~n47322 ;
  assign n47320 = n27977 & ~n47319 ;
  assign n47331 = \P2_P2_InstQueue_reg[7][0]/NET0131  & ~n28050 ;
  assign n47332 = ~n47320 & ~n47331 ;
  assign n47333 = ~n47323 & n47332 ;
  assign n47334 = ~n47330 & n47333 ;
  assign n47343 = n28610 & ~n46788 ;
  assign n47344 = n28632 & ~n46792 ;
  assign n47345 = ~n47343 & ~n47344 ;
  assign n47346 = \P2_P2_DataWidth_reg[1]/NET0131  & ~n47345 ;
  assign n47335 = ~n28428 & ~n46777 ;
  assign n47336 = \P2_P2_InstQueue_reg[8][0]/NET0131  & ~n28027 ;
  assign n47337 = ~n28423 & n47336 ;
  assign n47338 = ~n47335 & ~n47337 ;
  assign n47347 = ~n28687 & ~n47338 ;
  assign n47348 = ~n47346 & ~n47347 ;
  assign n47349 = n26794 & ~n47348 ;
  assign n47340 = ~n26544 & n28027 ;
  assign n47341 = ~n47336 & ~n47340 ;
  assign n47342 = n27613 & ~n47341 ;
  assign n47339 = n27977 & ~n47338 ;
  assign n47350 = \P2_P2_InstQueue_reg[8][0]/NET0131  & ~n28050 ;
  assign n47351 = ~n47339 & ~n47350 ;
  assign n47352 = ~n47342 & n47351 ;
  assign n47353 = ~n47349 & n47352 ;
  assign n47362 = n28632 & ~n46788 ;
  assign n47363 = n28423 & ~n46792 ;
  assign n47364 = ~n47362 & ~n47363 ;
  assign n47365 = \P2_P2_DataWidth_reg[1]/NET0131  & ~n47364 ;
  assign n47354 = ~n28041 & ~n46777 ;
  assign n47355 = \P2_P2_InstQueue_reg[9][0]/NET0131  & ~n28034 ;
  assign n47356 = ~n28027 & n47355 ;
  assign n47357 = ~n47354 & ~n47356 ;
  assign n47366 = ~n28707 & ~n47357 ;
  assign n47367 = ~n47365 & ~n47366 ;
  assign n47368 = n26794 & ~n47367 ;
  assign n47359 = ~n26544 & n28034 ;
  assign n47360 = ~n47355 & ~n47359 ;
  assign n47361 = n27613 & ~n47360 ;
  assign n47358 = n27977 & ~n47357 ;
  assign n47369 = \P2_P2_InstQueue_reg[9][0]/NET0131  & ~n28050 ;
  assign n47370 = ~n47358 & ~n47369 ;
  assign n47371 = ~n47361 & n47370 ;
  assign n47372 = ~n47368 & n47371 ;
  assign n47373 = \P1_P2_PhyAddrPointer_reg[4]/NET0131  & n25733 ;
  assign n47374 = ~n44190 & ~n47373 ;
  assign n47375 = n25701 & ~n47374 ;
  assign n47376 = \P1_P2_PhyAddrPointer_reg[4]/NET0131  & ~n36590 ;
  assign n47377 = ~n44198 & ~n47376 ;
  assign n47378 = ~n47375 & n47377 ;
  assign n47379 = n25918 & ~n47378 ;
  assign n47384 = \P1_P2_PhyAddrPointer_reg[1]/NET0131  & \P1_P2_PhyAddrPointer_reg[2]/NET0131  ;
  assign n47385 = \P1_P2_PhyAddrPointer_reg[3]/NET0131  & n47384 ;
  assign n47386 = ~\P1_P2_PhyAddrPointer_reg[4]/NET0131  & ~n47385 ;
  assign n47387 = \P1_P2_PhyAddrPointer_reg[1]/NET0131  & n36598 ;
  assign n47388 = ~n47386 & ~n47387 ;
  assign n47389 = n36630 & n47388 ;
  assign n47383 = \P1_P2_PhyAddrPointer_reg[4]/NET0131  & ~n39352 ;
  assign n47380 = ~\P1_P2_PhyAddrPointer_reg[4]/NET0131  & ~n36597 ;
  assign n47381 = ~n36598 & ~n47380 ;
  assign n47382 = n25933 & n47381 ;
  assign n47390 = ~n44178 & ~n47382 ;
  assign n47391 = ~n47383 & n47390 ;
  assign n47392 = ~n47389 & n47391 ;
  assign n47393 = ~n47379 & n47392 ;
  assign n47394 = \P2_P1_PhyAddrPointer_reg[4]/NET0131  & n25947 ;
  assign n47395 = ~n44245 & ~n47394 ;
  assign n47396 = n25945 & ~n47395 ;
  assign n47397 = \P2_P1_PhyAddrPointer_reg[4]/NET0131  & ~n36677 ;
  assign n47398 = ~n44252 & ~n47397 ;
  assign n47399 = ~n47396 & n47398 ;
  assign n47400 = n11623 & ~n47399 ;
  assign n47404 = ~n11617 & ~n25942 ;
  assign n47405 = n27787 & n47404 ;
  assign n47406 = \P2_P1_PhyAddrPointer_reg[4]/NET0131  & ~n47405 ;
  assign n47407 = \P2_P1_PhyAddrPointer_reg[1]/NET0131  & \P2_P1_PhyAddrPointer_reg[2]/NET0131  ;
  assign n47408 = \P2_P1_PhyAddrPointer_reg[3]/NET0131  & n47407 ;
  assign n47409 = ~\P2_P1_PhyAddrPointer_reg[4]/NET0131  & ~n47408 ;
  assign n47410 = \P2_P1_PhyAddrPointer_reg[1]/NET0131  & n36644 ;
  assign n47411 = ~n47409 & ~n47410 ;
  assign n47412 = n36674 & n47411 ;
  assign n47401 = ~\P2_P1_PhyAddrPointer_reg[4]/NET0131  & ~n36643 ;
  assign n47402 = ~n36644 & ~n47401 ;
  assign n47403 = n27681 & n47402 ;
  assign n47413 = ~n44234 & ~n47403 ;
  assign n47414 = ~n47412 & n47413 ;
  assign n47415 = ~n47406 & n47414 ;
  assign n47416 = ~n47400 & n47415 ;
  assign n47417 = \P1_P1_PhyAddrPointer_reg[4]/NET0131  & n26249 ;
  assign n47418 = ~n44435 & ~n47417 ;
  assign n47419 = n26126 & ~n47418 ;
  assign n47420 = \P1_P1_PhyAddrPointer_reg[4]/NET0131  & ~n36696 ;
  assign n47421 = ~n44421 & ~n47420 ;
  assign n47422 = ~n47419 & n47421 ;
  assign n47423 = n8355 & ~n47422 ;
  assign n47427 = ~n8358 & ~n26115 ;
  assign n47428 = n27611 & n47427 ;
  assign n47429 = \P1_P1_PhyAddrPointer_reg[4]/NET0131  & ~n47428 ;
  assign n47430 = \P1_P1_PhyAddrPointer_reg[1]/NET0131  & \P1_P1_PhyAddrPointer_reg[2]/NET0131  ;
  assign n47431 = \P1_P1_PhyAddrPointer_reg[3]/NET0131  & n47430 ;
  assign n47432 = ~\P1_P1_PhyAddrPointer_reg[4]/NET0131  & ~n47431 ;
  assign n47433 = \P1_P1_PhyAddrPointer_reg[1]/NET0131  & n36703 ;
  assign n47434 = ~n47432 & ~n47433 ;
  assign n47435 = ~n36701 & n47434 ;
  assign n47424 = ~\P1_P1_PhyAddrPointer_reg[4]/NET0131  & ~n36702 ;
  assign n47425 = ~n36703 & ~n47424 ;
  assign n47426 = n27791 & n47425 ;
  assign n47436 = ~n44412 & ~n47426 ;
  assign n47437 = ~n47435 & n47436 ;
  assign n47438 = ~n47429 & n47437 ;
  assign n47439 = ~n47423 & n47438 ;
  assign n47440 = \P2_P2_PhyAddrPointer_reg[4]/NET0131  & n26629 ;
  assign n47441 = ~n44297 & ~n47440 ;
  assign n47442 = n26621 & ~n47441 ;
  assign n47443 = \P2_P2_PhyAddrPointer_reg[4]/NET0131  & ~n36752 ;
  assign n47444 = ~n44306 & ~n47443 ;
  assign n47445 = ~n47442 & n47444 ;
  assign n47446 = n26792 & ~n47445 ;
  assign n47451 = \P2_P2_PhyAddrPointer_reg[1]/NET0131  & \P2_P2_PhyAddrPointer_reg[2]/NET0131  ;
  assign n47452 = \P2_P2_PhyAddrPointer_reg[3]/NET0131  & n47451 ;
  assign n47453 = ~\P2_P2_PhyAddrPointer_reg[4]/NET0131  & ~n47452 ;
  assign n47454 = \P2_P2_PhyAddrPointer_reg[4]/NET0131  & n47452 ;
  assign n47455 = ~n47453 & ~n47454 ;
  assign n47456 = ~n36760 & n47455 ;
  assign n47450 = \P2_P2_PhyAddrPointer_reg[4]/NET0131  & ~n36758 ;
  assign n47447 = ~\P2_P2_PhyAddrPointer_reg[4]/NET0131  & ~n36761 ;
  assign n47448 = ~n36762 & ~n47447 ;
  assign n47449 = n26800 & n47448 ;
  assign n47457 = ~n44288 & ~n47449 ;
  assign n47458 = ~n47450 & n47457 ;
  assign n47459 = ~n47456 & n47458 ;
  assign n47460 = ~n47446 & n47459 ;
  assign n47461 = \P1_P3_PhyAddrPointer_reg[4]/NET0131  & n9072 ;
  assign n47462 = ~n20438 & ~n47461 ;
  assign n47463 = n9064 & ~n47462 ;
  assign n47464 = \P1_P3_PhyAddrPointer_reg[4]/NET0131  & ~n36805 ;
  assign n47465 = ~n20452 & ~n47464 ;
  assign n47466 = ~n47463 & n47465 ;
  assign n47467 = n9241 & ~n47466 ;
  assign n47472 = n17534 & ~n36810 ;
  assign n47471 = \P1_P3_PhyAddrPointer_reg[4]/NET0131  & ~n36816 ;
  assign n47468 = ~\P1_P3_PhyAddrPointer_reg[4]/NET0131  & ~n16453 ;
  assign n47469 = ~n16454 & ~n47468 ;
  assign n47470 = n11698 & n47469 ;
  assign n47473 = ~n20430 & ~n47470 ;
  assign n47474 = ~n47471 & n47473 ;
  assign n47475 = ~n47472 & n47474 ;
  assign n47476 = ~n47467 & n47475 ;
  assign n47483 = \P2_P3_PhyAddrPointer_reg[4]/NET0131  & ~n27283 ;
  assign n47484 = ~n44369 & ~n47483 ;
  assign n47485 = n27117 & ~n47484 ;
  assign n47486 = \P2_P3_PhyAddrPointer_reg[4]/NET0131  & ~n36826 ;
  assign n47487 = ~n44376 & ~n47486 ;
  assign n47488 = ~n47485 & n47487 ;
  assign n47489 = n27308 & ~n47488 ;
  assign n47477 = \P2_P3_PhyAddrPointer_reg[1]/NET0131  & \P2_P3_PhyAddrPointer_reg[2]/NET0131  ;
  assign n47478 = \P2_P3_PhyAddrPointer_reg[3]/NET0131  & n47477 ;
  assign n47479 = ~\P2_P3_PhyAddrPointer_reg[4]/NET0131  & ~n47478 ;
  assign n47480 = \P2_P3_PhyAddrPointer_reg[1]/NET0131  & n36836 ;
  assign n47481 = ~n47479 & ~n47480 ;
  assign n47490 = ~\P2_P3_DataWidth_reg[1]/NET0131  & ~n47481 ;
  assign n47491 = ~\P2_P3_PhyAddrPointer_reg[4]/NET0131  & ~n36835 ;
  assign n47492 = ~n36836 & ~n47491 ;
  assign n47493 = \P2_P3_DataWidth_reg[1]/NET0131  & ~n47492 ;
  assign n47494 = n27315 & ~n47493 ;
  assign n47495 = ~n47490 & n47494 ;
  assign n47496 = \P2_P3_PhyAddrPointer_reg[4]/NET0131  & ~n36873 ;
  assign n47482 = n32867 & n47481 ;
  assign n47497 = ~n44349 & ~n47482 ;
  assign n47498 = ~n47496 & n47497 ;
  assign n47499 = ~n47495 & n47498 ;
  assign n47500 = ~n47489 & n47499 ;
  assign n47503 = ~\P2_P1_EBX_reg[30]/NET0131  & ~n46268 ;
  assign n47504 = n25981 & ~n46269 ;
  assign n47505 = ~n47503 & n47504 ;
  assign n47501 = n22335 & n46225 ;
  assign n47502 = \P2_P1_EBX_reg[30]/NET0131  & n46227 ;
  assign n47506 = ~n47501 & ~n47502 ;
  assign n47507 = ~n47505 & n47506 ;
  assign n47508 = n11623 & ~n47507 ;
  assign n47509 = \P2_P1_EBX_reg[30]/NET0131  & ~n21100 ;
  assign n47510 = ~n47508 & ~n47509 ;
  assign n47513 = ~\P1_P2_EBX_reg[30]/NET0131  & ~n46737 ;
  assign n47514 = n25803 & ~n46738 ;
  assign n47515 = ~n47513 & n47514 ;
  assign n47511 = n46675 & n46694 ;
  assign n47512 = \P1_P2_EBX_reg[30]/NET0131  & n46695 ;
  assign n47516 = ~n47511 & ~n47512 ;
  assign n47517 = ~n47515 & n47516 ;
  assign n47518 = n25918 & ~n47517 ;
  assign n47519 = \P1_P2_EBX_reg[30]/NET0131  & ~n43212 ;
  assign n47520 = ~n47518 & ~n47519 ;
  assign n47521 = \P2_P1_lWord_reg[3]/NET0131  & ~n34408 ;
  assign n47522 = \P2_P1_EAX_reg[3]/NET0131  & n24899 ;
  assign n47523 = n21062 & n24487 ;
  assign n47524 = ~n47522 & ~n47523 ;
  assign n47525 = n11623 & ~n47524 ;
  assign n47526 = ~n47521 & ~n47525 ;
  assign n47527 = ~n27607 & n27970 ;
  assign n47528 = n28928 & n47527 ;
  assign n47529 = n27968 & n47528 ;
  assign n47530 = \P1_P2_uWord_reg[12]/NET0131  & ~n47529 ;
  assign n47533 = ~\P1_P2_EAX_reg[13]/NET0131  & ~\P1_P2_EAX_reg[14]/NET0131  ;
  assign n47534 = ~\P1_P2_EAX_reg[15]/NET0131  & ~\P1_P2_EAX_reg[1]/NET0131  ;
  assign n47541 = n47533 & n47534 ;
  assign n47531 = ~\P1_P2_EAX_reg[0]/NET0131  & ~\P1_P2_EAX_reg[10]/NET0131  ;
  assign n47532 = ~\P1_P2_EAX_reg[11]/NET0131  & ~\P1_P2_EAX_reg[12]/NET0131  ;
  assign n47542 = n47531 & n47532 ;
  assign n47543 = n47541 & n47542 ;
  assign n47537 = ~\P1_P2_EAX_reg[6]/NET0131  & ~\P1_P2_EAX_reg[7]/NET0131  ;
  assign n47538 = ~\P1_P2_EAX_reg[8]/NET0131  & ~\P1_P2_EAX_reg[9]/NET0131  ;
  assign n47539 = n47537 & n47538 ;
  assign n47535 = ~\P1_P2_EAX_reg[2]/NET0131  & ~\P1_P2_EAX_reg[3]/NET0131  ;
  assign n47536 = ~\P1_P2_EAX_reg[4]/NET0131  & ~\P1_P2_EAX_reg[5]/NET0131  ;
  assign n47540 = n47535 & n47536 ;
  assign n47544 = n47539 & n47540 ;
  assign n47545 = n47543 & n47544 ;
  assign n47546 = \P1_P2_EAX_reg[31]/NET0131  & ~n47545 ;
  assign n47547 = \P1_P2_EAX_reg[16]/NET0131  & n47546 ;
  assign n47548 = \P1_P2_EAX_reg[17]/NET0131  & n47547 ;
  assign n47549 = \P1_P2_EAX_reg[18]/NET0131  & n47548 ;
  assign n47550 = \P1_P2_EAX_reg[19]/NET0131  & n47549 ;
  assign n47551 = \P1_P2_EAX_reg[20]/NET0131  & n47550 ;
  assign n47552 = \P1_P2_EAX_reg[21]/NET0131  & n47551 ;
  assign n47553 = \P1_P2_EAX_reg[22]/NET0131  & n47552 ;
  assign n47554 = \P1_P2_EAX_reg[23]/NET0131  & n47553 ;
  assign n47555 = \P1_P2_EAX_reg[24]/NET0131  & n47554 ;
  assign n47556 = \P1_P2_EAX_reg[25]/NET0131  & n47555 ;
  assign n47557 = \P1_P2_EAX_reg[26]/NET0131  & n47556 ;
  assign n47558 = \P1_P2_EAX_reg[27]/NET0131  & n47557 ;
  assign n47559 = ~\P1_P2_EAX_reg[28]/NET0131  & ~n47558 ;
  assign n47560 = \P1_P2_EAX_reg[28]/NET0131  & n47558 ;
  assign n47561 = ~n47559 & ~n47560 ;
  assign n47562 = n25757 & n47561 ;
  assign n47564 = ~\P1_buf1_reg[12]/NET0131  & n27934 ;
  assign n47563 = ~\P1_buf2_reg[12]/NET0131  & ~n27934 ;
  assign n47565 = ~n25415 & ~n47563 ;
  assign n47566 = ~n47564 & n47565 ;
  assign n47567 = n25776 & n47566 ;
  assign n47568 = ~n47562 & ~n47567 ;
  assign n47569 = ~n25770 & ~n47568 ;
  assign n47570 = n25757 & ~n25770 ;
  assign n47571 = ~n25846 & ~n47570 ;
  assign n47572 = ~n31470 & ~n47571 ;
  assign n47573 = \P1_P2_uWord_reg[12]/NET0131  & ~n47572 ;
  assign n47574 = ~n47569 & ~n47573 ;
  assign n47575 = n25918 & ~n47574 ;
  assign n47576 = ~n47530 & ~n47575 ;
  assign n47577 = \P2_P2_EAX_reg[26]/NET0131  & ~n44508 ;
  assign n47581 = ~n44729 & n44732 ;
  assign n47582 = ~n44736 & ~n47581 ;
  assign n47583 = \P2_P2_EAX_reg[26]/NET0131  & ~n47582 ;
  assign n47594 = ~\P2_P2_EAX_reg[26]/NET0131  & n44732 ;
  assign n47595 = n44729 & n47594 ;
  assign n47584 = \P2_P2_EAX_reg[26]/NET0131  & ~n26641 ;
  assign n47588 = \P2_buf2_reg[10]/NET0131  & ~n28013 ;
  assign n47589 = \P2_buf1_reg[10]/NET0131  & n28013 ;
  assign n47590 = ~n47588 & ~n47589 ;
  assign n47591 = n26641 & ~n47590 ;
  assign n47592 = ~n47584 & ~n47591 ;
  assign n47593 = n26633 & ~n47592 ;
  assign n47578 = ~n44637 & n44668 ;
  assign n47579 = ~n44669 & ~n47578 ;
  assign n47580 = n44510 & n47579 ;
  assign n47585 = n26641 & ~n36002 ;
  assign n47586 = ~n47584 & ~n47585 ;
  assign n47587 = n26638 & ~n47586 ;
  assign n47596 = ~n47580 & ~n47587 ;
  assign n47597 = ~n47593 & n47596 ;
  assign n47598 = ~n47595 & n47597 ;
  assign n47599 = ~n47583 & n47598 ;
  assign n47600 = n26792 & ~n47599 ;
  assign n47601 = ~n47577 & ~n47600 ;
  assign n47604 = ~\P2_P2_EBX_reg[30]/NET0131  & ~n46459 ;
  assign n47605 = n26662 & ~n46460 ;
  assign n47606 = ~n47604 & n47605 ;
  assign n47602 = n46385 & n46416 ;
  assign n47603 = \P2_P2_EBX_reg[30]/NET0131  & n46417 ;
  assign n47607 = ~n47602 & ~n47603 ;
  assign n47608 = ~n47606 & n47607 ;
  assign n47609 = n26792 & ~n47608 ;
  assign n47610 = \P2_P2_EBX_reg[30]/NET0131  & ~n44508 ;
  assign n47611 = ~n47609 & ~n47610 ;
  assign n47612 = \P1_P1_EAX_reg[3]/NET0131  & n24502 ;
  assign n47613 = ~n7913 & n23946 ;
  assign n47614 = ~n47612 & ~n47613 ;
  assign n47615 = ~n15364 & ~n47614 ;
  assign n47616 = \P1_P1_lWord_reg[3]/NET0131  & ~n24506 ;
  assign n47617 = ~n47615 & ~n47616 ;
  assign n47618 = n8355 & ~n47617 ;
  assign n47619 = \P1_P1_lWord_reg[3]/NET0131  & ~n24515 ;
  assign n47620 = ~n47618 & ~n47619 ;
  assign n47623 = ~\P1_P3_EBX_reg[30]/NET0131  & ~n46521 ;
  assign n47624 = n9108 & ~n46522 ;
  assign n47625 = ~n47623 & n47624 ;
  assign n47621 = n21719 & n46479 ;
  assign n47622 = \P1_P3_EBX_reg[30]/NET0131  & n46480 ;
  assign n47626 = ~n47621 & ~n47622 ;
  assign n47627 = ~n47625 & n47626 ;
  assign n47628 = n9241 & ~n47627 ;
  assign n47629 = \P1_P3_EBX_reg[30]/NET0131  & ~n16968 ;
  assign n47630 = ~n47628 & ~n47629 ;
  assign n47633 = ~\P1_P1_EBX_reg[30]/NET0131  & ~n46576 ;
  assign n47634 = n26146 & ~n46577 ;
  assign n47635 = ~n47633 & n47634 ;
  assign n47631 = \P1_P1_EBX_reg[30]/NET0131  & ~n46533 ;
  assign n47632 = n22856 & n46535 ;
  assign n47636 = ~n47631 & ~n47632 ;
  assign n47637 = ~n47635 & n47636 ;
  assign n47638 = n8355 & ~n47637 ;
  assign n47639 = \P1_P1_EBX_reg[30]/NET0131  & ~n15326 ;
  assign n47640 = ~n47638 & ~n47639 ;
  assign n47641 = ~n43243 & n44507 ;
  assign n47642 = n45044 & n47641 ;
  assign n47643 = \P2_P2_uWord_reg[12]/NET0131  & ~n47642 ;
  assign n47646 = ~\P2_P2_EAX_reg[13]/NET0131  & ~\P2_P2_EAX_reg[14]/NET0131  ;
  assign n47647 = ~\P2_P2_EAX_reg[15]/NET0131  & ~\P2_P2_EAX_reg[1]/NET0131  ;
  assign n47654 = n47646 & n47647 ;
  assign n47644 = ~\P2_P2_EAX_reg[0]/NET0131  & ~\P2_P2_EAX_reg[10]/NET0131  ;
  assign n47645 = ~\P2_P2_EAX_reg[11]/NET0131  & ~\P2_P2_EAX_reg[12]/NET0131  ;
  assign n47655 = n47644 & n47645 ;
  assign n47656 = n47654 & n47655 ;
  assign n47650 = ~\P2_P2_EAX_reg[6]/NET0131  & ~\P2_P2_EAX_reg[7]/NET0131  ;
  assign n47651 = ~\P2_P2_EAX_reg[8]/NET0131  & ~\P2_P2_EAX_reg[9]/NET0131  ;
  assign n47652 = n47650 & n47651 ;
  assign n47648 = ~\P2_P2_EAX_reg[2]/NET0131  & ~\P2_P2_EAX_reg[3]/NET0131  ;
  assign n47649 = ~\P2_P2_EAX_reg[4]/NET0131  & ~\P2_P2_EAX_reg[5]/NET0131  ;
  assign n47653 = n47648 & n47649 ;
  assign n47657 = n47652 & n47653 ;
  assign n47658 = n47656 & n47657 ;
  assign n47659 = \P2_P2_EAX_reg[31]/NET0131  & ~n47658 ;
  assign n47660 = \P2_P2_EAX_reg[16]/NET0131  & n47659 ;
  assign n47661 = \P2_P2_EAX_reg[17]/NET0131  & n47660 ;
  assign n47662 = \P2_P2_EAX_reg[18]/NET0131  & n47661 ;
  assign n47663 = \P2_P2_EAX_reg[19]/NET0131  & n47662 ;
  assign n47664 = \P2_P2_EAX_reg[20]/NET0131  & n47663 ;
  assign n47665 = \P2_P2_EAX_reg[21]/NET0131  & n47664 ;
  assign n47666 = \P2_P2_EAX_reg[22]/NET0131  & n47665 ;
  assign n47667 = \P2_P2_EAX_reg[23]/NET0131  & n47666 ;
  assign n47668 = \P2_P2_EAX_reg[24]/NET0131  & n47667 ;
  assign n47669 = \P2_P2_EAX_reg[25]/NET0131  & n47668 ;
  assign n47670 = \P2_P2_EAX_reg[26]/NET0131  & n47669 ;
  assign n47671 = \P2_P2_EAX_reg[27]/NET0131  & n47670 ;
  assign n47672 = ~\P2_P2_EAX_reg[28]/NET0131  & ~n47671 ;
  assign n47673 = \P2_P2_EAX_reg[28]/NET0131  & n47671 ;
  assign n47674 = ~n47672 & ~n47673 ;
  assign n47675 = n26643 & n47674 ;
  assign n47676 = ~n26286 & n26633 ;
  assign n47677 = \P2_buf2_reg[12]/NET0131  & ~n28013 ;
  assign n47678 = \P2_buf1_reg[12]/NET0131  & n28013 ;
  assign n47679 = ~n47677 & ~n47678 ;
  assign n47680 = n47676 & ~n47679 ;
  assign n47681 = ~n47675 & ~n47680 ;
  assign n47682 = ~n26640 & ~n47681 ;
  assign n47683 = n26286 & n26633 ;
  assign n47684 = n26633 & ~n26640 ;
  assign n47685 = ~n26786 & ~n47684 ;
  assign n47686 = ~n47683 & ~n47685 ;
  assign n47687 = \P2_P2_uWord_reg[12]/NET0131  & ~n47686 ;
  assign n47688 = ~n47682 & ~n47687 ;
  assign n47689 = n26792 & ~n47688 ;
  assign n47690 = ~n47643 & ~n47689 ;
  assign n47693 = ~\P2_P3_EAX_reg[26]/NET0131  & ~n46594 ;
  assign n47692 = \P2_P3_EAX_reg[26]/NET0131  & n46594 ;
  assign n47694 = n42539 & ~n47692 ;
  assign n47695 = ~n47693 & n47694 ;
  assign n47691 = \P2_P3_EAX_reg[26]/NET0131  & ~n42543 ;
  assign n47696 = \P2_buf2_reg[10]/NET0131  & n27122 ;
  assign n47697 = \P2_buf2_reg[26]/NET0131  & n27186 ;
  assign n47698 = ~n47696 & ~n47697 ;
  assign n47699 = n27227 & ~n47698 ;
  assign n47700 = ~n42671 & n42702 ;
  assign n47701 = ~n42703 & ~n47700 ;
  assign n47702 = n42538 & n47701 ;
  assign n47703 = ~n47699 & ~n47702 ;
  assign n47704 = ~n47691 & n47703 ;
  assign n47705 = ~n47695 & n47704 ;
  assign n47706 = n27308 & ~n47705 ;
  assign n47707 = \P2_P3_EAX_reg[26]/NET0131  & ~n42872 ;
  assign n47708 = ~n47706 & ~n47707 ;
  assign n47711 = ~\P2_P3_EBX_reg[30]/NET0131  & ~n46656 ;
  assign n47712 = n27133 & ~n46657 ;
  assign n47713 = ~n47711 & n47712 ;
  assign n47709 = n46603 & n46614 ;
  assign n47710 = \P2_P3_EBX_reg[30]/NET0131  & n46615 ;
  assign n47714 = ~n47709 & ~n47710 ;
  assign n47715 = ~n47713 & n47714 ;
  assign n47716 = n27308 & ~n47715 ;
  assign n47717 = \P2_P3_EBX_reg[30]/NET0131  & ~n42872 ;
  assign n47718 = ~n47716 & ~n47717 ;
  assign n47719 = \P1_P2_EAX_reg[26]/NET0131  & ~n43212 ;
  assign n47724 = ~\P1_P2_EAX_reg[26]/NET0131  & ~n43195 ;
  assign n47725 = n43164 & ~n43196 ;
  assign n47726 = ~n47724 & n47725 ;
  assign n47727 = \P1_P2_EAX_reg[26]/NET0131  & n43167 ;
  assign n47720 = ~n43002 & n43033 ;
  assign n47721 = n25747 & ~n43034 ;
  assign n47722 = ~n47720 & n47721 ;
  assign n47723 = n25742 & n47722 ;
  assign n47728 = \P1_P2_EAX_reg[26]/NET0131  & ~n25773 ;
  assign n47730 = ~\P1_buf1_reg[10]/NET0131  & n27934 ;
  assign n47729 = ~\P1_buf2_reg[10]/NET0131  & ~n27934 ;
  assign n47731 = ~n25415 & ~n47729 ;
  assign n47732 = ~n47730 & n47731 ;
  assign n47733 = ~n25770 & n47732 ;
  assign n47734 = ~n47728 & ~n47733 ;
  assign n47735 = n25776 & ~n47734 ;
  assign n47736 = n25773 & ~n35971 ;
  assign n47737 = ~n47728 & ~n47736 ;
  assign n47738 = n25774 & ~n47737 ;
  assign n47739 = ~n47735 & ~n47738 ;
  assign n47740 = ~n47723 & n47739 ;
  assign n47741 = ~n47727 & n47740 ;
  assign n47742 = ~n47726 & n47741 ;
  assign n47743 = n25918 & ~n47742 ;
  assign n47744 = ~n47719 & ~n47743 ;
  assign n47745 = n42870 & n43271 ;
  assign n47746 = n43269 & n47745 ;
  assign n47747 = n27121 & ~n27177 ;
  assign n47748 = ~n46587 & ~n47747 ;
  assign n47749 = n27122 & n27192 ;
  assign n47750 = ~n47748 & ~n47749 ;
  assign n47751 = n27308 & ~n47750 ;
  assign n47752 = n47746 & ~n47751 ;
  assign n47753 = \P2_P3_uWord_reg[12]/NET0131  & ~n47752 ;
  assign n47754 = ~n27177 & n27308 ;
  assign n47755 = \P2_buf2_reg[12]/NET0131  & ~n27192 ;
  assign n47756 = n27122 & n47755 ;
  assign n47759 = ~\P2_P3_EAX_reg[13]/NET0131  & ~\P2_P3_EAX_reg[14]/NET0131  ;
  assign n47760 = ~\P2_P3_EAX_reg[15]/NET0131  & ~\P2_P3_EAX_reg[1]/NET0131  ;
  assign n47767 = n47759 & n47760 ;
  assign n47757 = ~\P2_P3_EAX_reg[0]/NET0131  & ~\P2_P3_EAX_reg[10]/NET0131  ;
  assign n47758 = ~\P2_P3_EAX_reg[11]/NET0131  & ~\P2_P3_EAX_reg[12]/NET0131  ;
  assign n47768 = n47757 & n47758 ;
  assign n47769 = n47767 & n47768 ;
  assign n47763 = ~\P2_P3_EAX_reg[6]/NET0131  & ~\P2_P3_EAX_reg[7]/NET0131  ;
  assign n47764 = ~\P2_P3_EAX_reg[8]/NET0131  & ~\P2_P3_EAX_reg[9]/NET0131  ;
  assign n47765 = n47763 & n47764 ;
  assign n47761 = ~\P2_P3_EAX_reg[2]/NET0131  & ~\P2_P3_EAX_reg[3]/NET0131  ;
  assign n47762 = ~\P2_P3_EAX_reg[4]/NET0131  & ~\P2_P3_EAX_reg[5]/NET0131  ;
  assign n47766 = n47761 & n47762 ;
  assign n47770 = n47765 & n47766 ;
  assign n47771 = n47769 & n47770 ;
  assign n47772 = \P2_P3_EAX_reg[31]/NET0131  & ~n47771 ;
  assign n47773 = \P2_P3_EAX_reg[16]/NET0131  & n47772 ;
  assign n47774 = \P2_P3_EAX_reg[17]/NET0131  & n47773 ;
  assign n47775 = \P2_P3_EAX_reg[18]/NET0131  & n47774 ;
  assign n47776 = \P2_P3_EAX_reg[19]/NET0131  & n47775 ;
  assign n47777 = n46593 & n47776 ;
  assign n47778 = n46590 & n47777 ;
  assign n47779 = \P2_P3_EAX_reg[28]/NET0131  & n47778 ;
  assign n47780 = ~\P2_P3_EAX_reg[28]/NET0131  & ~n47778 ;
  assign n47781 = ~n47779 & ~n47780 ;
  assign n47782 = n27121 & n47781 ;
  assign n47783 = ~n47756 & ~n47782 ;
  assign n47784 = n47754 & ~n47783 ;
  assign n47785 = ~n47753 & ~n47784 ;
  assign n47795 = n25874 & n46065 ;
  assign n47796 = \P1_P2_PhyAddrPointer_reg[3]/NET0131  & ~n39340 ;
  assign n47797 = ~n46078 & ~n47796 ;
  assign n47798 = ~n47795 & n47797 ;
  assign n47799 = n25918 & ~n47798 ;
  assign n47786 = \P1_P2_PhyAddrPointer_reg[2]/NET0131  & ~n37915 ;
  assign n47787 = n25928 & ~n47786 ;
  assign n47788 = n36595 & ~n47787 ;
  assign n47789 = \P1_P2_PhyAddrPointer_reg[3]/NET0131  & ~n47788 ;
  assign n47793 = ~\P1_P2_PhyAddrPointer_reg[3]/NET0131  & n47786 ;
  assign n47794 = n25928 & n47793 ;
  assign n47790 = ~\P1_P2_PhyAddrPointer_reg[3]/NET0131  & ~n47384 ;
  assign n47791 = ~n47385 & ~n47790 ;
  assign n47792 = n27898 & n47791 ;
  assign n47800 = ~n46047 & ~n47792 ;
  assign n47801 = ~n47794 & n47800 ;
  assign n47802 = ~n47789 & n47801 ;
  assign n47803 = ~n47799 & n47802 ;
  assign n47808 = \P1_P2_PhyAddrPointer_reg[5]/NET0131  & n25733 ;
  assign n47809 = ~n45458 & ~n47808 ;
  assign n47810 = n25701 & ~n47809 ;
  assign n47811 = \P1_P2_PhyAddrPointer_reg[5]/NET0131  & ~n36590 ;
  assign n47812 = ~n45444 & ~n47811 ;
  assign n47813 = ~n47810 & n47812 ;
  assign n47814 = n25918 & ~n47813 ;
  assign n47804 = \P1_P2_PhyAddrPointer_reg[1]/NET0131  & n36599 ;
  assign n47805 = ~\P1_P2_PhyAddrPointer_reg[5]/NET0131  & ~n47387 ;
  assign n47806 = ~n47804 & ~n47805 ;
  assign n47815 = ~\P1_P2_DataWidth_reg[1]/NET0131  & ~n47806 ;
  assign n47816 = ~\P1_P2_PhyAddrPointer_reg[5]/NET0131  & ~n36598 ;
  assign n47817 = ~n36599 & ~n47816 ;
  assign n47818 = \P1_P2_DataWidth_reg[1]/NET0131  & ~n47817 ;
  assign n47819 = n25928 & ~n47818 ;
  assign n47820 = ~n47815 & n47819 ;
  assign n47807 = n27898 & n47806 ;
  assign n47821 = \P1_P2_PhyAddrPointer_reg[5]/NET0131  & ~n39352 ;
  assign n47822 = ~n45436 & ~n47821 ;
  assign n47823 = ~n47807 & n47822 ;
  assign n47824 = ~n47820 & n47823 ;
  assign n47825 = ~n47814 & n47824 ;
  assign n47828 = \P1_P2_PhyAddrPointer_reg[6]/NET0131  & n25733 ;
  assign n47829 = ~n44215 & ~n47828 ;
  assign n47830 = n25701 & ~n47829 ;
  assign n47831 = \P1_P2_PhyAddrPointer_reg[6]/NET0131  & ~n36590 ;
  assign n47832 = ~n44225 & ~n47831 ;
  assign n47833 = ~n47830 & n47832 ;
  assign n47834 = n25918 & ~n47833 ;
  assign n47826 = n25933 & ~n36600 ;
  assign n47838 = n36595 & ~n47826 ;
  assign n47839 = \P1_P2_PhyAddrPointer_reg[6]/NET0131  & ~n47838 ;
  assign n47835 = ~\P1_P2_PhyAddrPointer_reg[6]/NET0131  & ~n47804 ;
  assign n47836 = ~n43517 & ~n47835 ;
  assign n47837 = n36630 & n47836 ;
  assign n47827 = n36599 & n47826 ;
  assign n47840 = ~n44207 & ~n47827 ;
  assign n47841 = ~n47837 & n47840 ;
  assign n47842 = ~n47839 & n47841 ;
  assign n47843 = ~n47834 & n47842 ;
  assign n47855 = \P2_P1_PhyAddrPointer_reg[3]/NET0131  & n25947 ;
  assign n47856 = ~n45381 & ~n47855 ;
  assign n47857 = n25945 & ~n47856 ;
  assign n47858 = \P2_P1_PhyAddrPointer_reg[3]/NET0131  & ~n36677 ;
  assign n47859 = ~n45358 & ~n47858 ;
  assign n47860 = ~n47857 & n47859 ;
  assign n47861 = n11623 & ~n47860 ;
  assign n47844 = n27787 & n36686 ;
  assign n47845 = \P2_P1_PhyAddrPointer_reg[3]/NET0131  & ~n47844 ;
  assign n47846 = \P2_P1_PhyAddrPointer_reg[2]/NET0131  & ~n39474 ;
  assign n47847 = ~\P2_P1_PhyAddrPointer_reg[3]/NET0131  & ~n47846 ;
  assign n47848 = n36643 & ~n39474 ;
  assign n47849 = n11609 & ~n47848 ;
  assign n47850 = ~n47847 & n47849 ;
  assign n47854 = \P2_P1_PhyAddrPointer_reg[3]/NET0131  & n11625 ;
  assign n47851 = ~\P2_P1_PhyAddrPointer_reg[3]/NET0131  & ~n47407 ;
  assign n47852 = ~n47408 & ~n47851 ;
  assign n47853 = n11613 & n47852 ;
  assign n47862 = ~n45350 & ~n47853 ;
  assign n47863 = ~n47854 & n47862 ;
  assign n47864 = ~n47850 & n47863 ;
  assign n47865 = ~n47845 & n47864 ;
  assign n47866 = ~n47861 & n47865 ;
  assign n47867 = \P2_P1_PhyAddrPointer_reg[5]/NET0131  & n25947 ;
  assign n47868 = ~n45409 & ~n47867 ;
  assign n47869 = n25945 & ~n47868 ;
  assign n47870 = \P2_P1_PhyAddrPointer_reg[5]/NET0131  & ~n36677 ;
  assign n47871 = ~n45418 & ~n47870 ;
  assign n47872 = ~n47869 & n47871 ;
  assign n47873 = n11623 & ~n47872 ;
  assign n47877 = \P2_P1_PhyAddrPointer_reg[5]/NET0131  & ~n36687 ;
  assign n47878 = \P2_P1_PhyAddrPointer_reg[1]/NET0131  & n36645 ;
  assign n47879 = ~\P2_P1_PhyAddrPointer_reg[5]/NET0131  & ~n47410 ;
  assign n47880 = ~n47878 & ~n47879 ;
  assign n47881 = n36674 & n47880 ;
  assign n47874 = ~\P2_P1_PhyAddrPointer_reg[5]/NET0131  & ~n36644 ;
  assign n47875 = n27681 & ~n36645 ;
  assign n47876 = ~n47874 & n47875 ;
  assign n47882 = ~n45393 & ~n47876 ;
  assign n47883 = ~n47881 & n47882 ;
  assign n47884 = ~n47877 & n47883 ;
  assign n47885 = ~n47873 & n47884 ;
  assign n47893 = \P2_P1_PhyAddrPointer_reg[6]/NET0131  & n25947 ;
  assign n47894 = ~n44269 & ~n47893 ;
  assign n47895 = n25945 & ~n47894 ;
  assign n47896 = \P2_P1_PhyAddrPointer_reg[6]/NET0131  & ~n36677 ;
  assign n47897 = ~n44279 & ~n47896 ;
  assign n47898 = ~n47895 & n47897 ;
  assign n47899 = n11623 & ~n47898 ;
  assign n47886 = n36687 & ~n47875 ;
  assign n47887 = \P2_P1_PhyAddrPointer_reg[6]/NET0131  & ~n47886 ;
  assign n47890 = ~\P2_P1_PhyAddrPointer_reg[6]/NET0131  & ~n47878 ;
  assign n47891 = ~n43577 & ~n47890 ;
  assign n47892 = n36674 & n47891 ;
  assign n47888 = ~\P2_P1_PhyAddrPointer_reg[6]/NET0131  & n36645 ;
  assign n47889 = n27681 & n47888 ;
  assign n47900 = ~n44261 & ~n47889 ;
  assign n47901 = ~n47892 & n47900 ;
  assign n47902 = ~n47887 & n47901 ;
  assign n47903 = ~n47899 & n47902 ;
  assign n47915 = \P1_P1_PhyAddrPointer_reg[3]/NET0131  & n26249 ;
  assign n47916 = ~n46024 & ~n47915 ;
  assign n47917 = n26126 & ~n47916 ;
  assign n47918 = \P1_P1_PhyAddrPointer_reg[3]/NET0131  & ~n36696 ;
  assign n47919 = ~n46038 & ~n47918 ;
  assign n47920 = ~n47917 & n47919 ;
  assign n47921 = n8355 & ~n47920 ;
  assign n47904 = n27611 & n36742 ;
  assign n47905 = \P1_P1_PhyAddrPointer_reg[3]/NET0131  & ~n47904 ;
  assign n47906 = \P1_P1_PhyAddrPointer_reg[2]/NET0131  & ~n39569 ;
  assign n47907 = ~\P1_P1_PhyAddrPointer_reg[3]/NET0131  & ~n47906 ;
  assign n47908 = n36702 & ~n39569 ;
  assign n47909 = n8282 & ~n47908 ;
  assign n47910 = ~n47907 & n47909 ;
  assign n47914 = \P1_P1_PhyAddrPointer_reg[3]/NET0131  & n8361 ;
  assign n47911 = ~\P1_P1_PhyAddrPointer_reg[3]/NET0131  & ~n47430 ;
  assign n47912 = ~n47431 & ~n47911 ;
  assign n47913 = n8287 & n47912 ;
  assign n47922 = ~n46009 & ~n47913 ;
  assign n47923 = ~n47914 & n47922 ;
  assign n47924 = ~n47910 & n47923 ;
  assign n47925 = ~n47905 & n47924 ;
  assign n47926 = ~n47921 & n47925 ;
  assign n47927 = \P1_P1_PhyAddrPointer_reg[5]/NET0131  & n26249 ;
  assign n47928 = ~n46114 & ~n47927 ;
  assign n47929 = n26126 & ~n47928 ;
  assign n47930 = \P1_P1_PhyAddrPointer_reg[5]/NET0131  & ~n36696 ;
  assign n47931 = ~n46096 & ~n47930 ;
  assign n47932 = ~n47929 & n47931 ;
  assign n47933 = n8355 & ~n47932 ;
  assign n47937 = \P1_P1_PhyAddrPointer_reg[5]/NET0131  & ~n36743 ;
  assign n47938 = \P1_P1_PhyAddrPointer_reg[1]/NET0131  & n36704 ;
  assign n47939 = ~\P1_P1_PhyAddrPointer_reg[5]/NET0131  & ~n47433 ;
  assign n47940 = ~n47938 & ~n47939 ;
  assign n47941 = ~n36701 & n47940 ;
  assign n47934 = ~\P1_P1_PhyAddrPointer_reg[5]/NET0131  & ~n36703 ;
  assign n47935 = n27791 & ~n36704 ;
  assign n47936 = ~n47934 & n47935 ;
  assign n47942 = ~n46086 & ~n47936 ;
  assign n47943 = ~n47941 & n47942 ;
  assign n47944 = ~n47937 & n47943 ;
  assign n47945 = ~n47933 & n47944 ;
  assign n47953 = \P1_P1_PhyAddrPointer_reg[6]/NET0131  & n26249 ;
  assign n47954 = ~n44460 & ~n47953 ;
  assign n47955 = n26126 & ~n47954 ;
  assign n47956 = \P1_P1_PhyAddrPointer_reg[6]/NET0131  & ~n36696 ;
  assign n47957 = ~n44467 & ~n47956 ;
  assign n47958 = ~n47955 & n47957 ;
  assign n47959 = n8355 & ~n47958 ;
  assign n47946 = n36743 & ~n47935 ;
  assign n47947 = \P1_P1_PhyAddrPointer_reg[6]/NET0131  & ~n47946 ;
  assign n47950 = ~\P1_P1_PhyAddrPointer_reg[6]/NET0131  & ~n47938 ;
  assign n47951 = ~n43737 & ~n47950 ;
  assign n47952 = ~n36701 & n47951 ;
  assign n47948 = ~\P1_P1_PhyAddrPointer_reg[6]/NET0131  & n36704 ;
  assign n47949 = n27791 & n47948 ;
  assign n47960 = ~n44446 & ~n47949 ;
  assign n47961 = ~n47952 & n47960 ;
  assign n47962 = ~n47947 & n47961 ;
  assign n47963 = ~n47959 & n47962 ;
  assign n47967 = n26749 & n45594 ;
  assign n47968 = \P2_P2_PhyAddrPointer_reg[3]/NET0131  & ~n41873 ;
  assign n47969 = ~n45582 & ~n47968 ;
  assign n47970 = ~n47967 & n47969 ;
  assign n47971 = n26792 & ~n47970 ;
  assign n47974 = \P2_P2_PhyAddrPointer_reg[2]/NET0131  & ~n37979 ;
  assign n47975 = ~\P2_P2_PhyAddrPointer_reg[3]/NET0131  & ~n47974 ;
  assign n47973 = n36761 & ~n37979 ;
  assign n47976 = n26794 & ~n47973 ;
  assign n47977 = ~n47975 & n47976 ;
  assign n47972 = \P2_P2_PhyAddrPointer_reg[3]/NET0131  & ~n36758 ;
  assign n47964 = ~\P2_P2_PhyAddrPointer_reg[3]/NET0131  & ~n47451 ;
  assign n47965 = ~n47452 & ~n47964 ;
  assign n47966 = n27977 & n47965 ;
  assign n47978 = ~n45569 & ~n47966 ;
  assign n47979 = ~n47972 & n47978 ;
  assign n47980 = ~n47977 & n47979 ;
  assign n47981 = ~n47971 & n47980 ;
  assign n47985 = \P2_P2_PhyAddrPointer_reg[5]/NET0131  & n26629 ;
  assign n47986 = ~n45624 & ~n47985 ;
  assign n47987 = n26621 & ~n47986 ;
  assign n47988 = \P2_P2_PhyAddrPointer_reg[5]/NET0131  & ~n36752 ;
  assign n47989 = ~n45632 & ~n47988 ;
  assign n47990 = ~n47987 & n47989 ;
  assign n47991 = n26792 & ~n47990 ;
  assign n47982 = ~\P2_P2_PhyAddrPointer_reg[5]/NET0131  & ~n47454 ;
  assign n47983 = ~n45079 & ~n47982 ;
  assign n47992 = ~\P2_P2_DataWidth_reg[1]/NET0131  & ~n47983 ;
  assign n47993 = ~\P2_P2_PhyAddrPointer_reg[5]/NET0131  & ~n36762 ;
  assign n47994 = ~n36763 & ~n47993 ;
  assign n47995 = \P2_P2_DataWidth_reg[1]/NET0131  & ~n47994 ;
  assign n47996 = n26794 & ~n47995 ;
  assign n47997 = ~n47992 & n47996 ;
  assign n47984 = n27977 & n47983 ;
  assign n47998 = \P2_P2_PhyAddrPointer_reg[5]/NET0131  & ~n36758 ;
  assign n47999 = ~n45614 & ~n47998 ;
  assign n48000 = ~n47984 & n47999 ;
  assign n48001 = ~n47997 & n48000 ;
  assign n48002 = ~n47991 & n48001 ;
  assign n48006 = n26621 & n44331 ;
  assign n48007 = \P2_P2_PhyAddrPointer_reg[6]/NET0131  & ~n41873 ;
  assign n48008 = ~n44340 & ~n48007 ;
  assign n48009 = ~n48006 & n48008 ;
  assign n48010 = n26792 & ~n48009 ;
  assign n48003 = ~\P2_P2_PhyAddrPointer_reg[6]/NET0131  & ~n45079 ;
  assign n48004 = ~n45080 & ~n48003 ;
  assign n48011 = ~\P2_P2_DataWidth_reg[1]/NET0131  & ~n48004 ;
  assign n48012 = ~\P2_P2_PhyAddrPointer_reg[6]/NET0131  & ~n36763 ;
  assign n48013 = ~n36764 & ~n48012 ;
  assign n48014 = \P2_P2_DataWidth_reg[1]/NET0131  & ~n48013 ;
  assign n48015 = n26794 & ~n48014 ;
  assign n48016 = ~n48011 & n48015 ;
  assign n48005 = n27977 & n48004 ;
  assign n48017 = \P2_P2_PhyAddrPointer_reg[6]/NET0131  & ~n36758 ;
  assign n48018 = ~n44315 & ~n48017 ;
  assign n48019 = ~n48005 & n48018 ;
  assign n48020 = ~n48016 & n48019 ;
  assign n48021 = ~n48010 & n48020 ;
  assign n48029 = n9192 & n20399 ;
  assign n48030 = \P1_P3_PhyAddrPointer_reg[3]/NET0131  & ~n37992 ;
  assign n48031 = ~n20419 & ~n48030 ;
  assign n48032 = ~n48029 & n48031 ;
  assign n48033 = n9241 & ~n48032 ;
  assign n48025 = \P1_P3_PhyAddrPointer_reg[2]/NET0131  & ~n42000 ;
  assign n48026 = ~\P1_P3_PhyAddrPointer_reg[3]/NET0131  & ~n48025 ;
  assign n48024 = n16453 & ~n42000 ;
  assign n48027 = n9245 & ~n48024 ;
  assign n48028 = ~n48026 & n48027 ;
  assign n48023 = \P1_P3_PhyAddrPointer_reg[3]/NET0131  & ~n36816 ;
  assign n48022 = n16451 & n16492 ;
  assign n48034 = ~n20384 & ~n48022 ;
  assign n48035 = ~n48023 & n48034 ;
  assign n48036 = ~n48028 & n48035 ;
  assign n48037 = ~n48033 & n48036 ;
  assign n48039 = n9064 & n20488 ;
  assign n48040 = \P1_P3_PhyAddrPointer_reg[5]/NET0131  & ~n37992 ;
  assign n48041 = ~n20474 & ~n48040 ;
  assign n48042 = ~n48039 & n48041 ;
  assign n48043 = n9241 & ~n48042 ;
  assign n48044 = ~\P1_P3_DataWidth_reg[1]/NET0131  & ~n21734 ;
  assign n48045 = ~\P1_P3_PhyAddrPointer_reg[5]/NET0131  & ~n16454 ;
  assign n48046 = ~n16455 & ~n48045 ;
  assign n48047 = \P1_P3_DataWidth_reg[1]/NET0131  & ~n48046 ;
  assign n48048 = n9245 & ~n48047 ;
  assign n48049 = ~n48044 & n48048 ;
  assign n48038 = n16492 & n21734 ;
  assign n48050 = \P1_P3_PhyAddrPointer_reg[5]/NET0131  & ~n36816 ;
  assign n48051 = ~n20466 & ~n48050 ;
  assign n48052 = ~n48038 & n48051 ;
  assign n48053 = ~n48049 & n48052 ;
  assign n48054 = ~n48043 & n48053 ;
  assign n48056 = n9064 & n20514 ;
  assign n48057 = \P1_P3_PhyAddrPointer_reg[6]/NET0131  & ~n37992 ;
  assign n48058 = ~n20522 & ~n48057 ;
  assign n48059 = ~n48056 & n48058 ;
  assign n48060 = n9241 & ~n48059 ;
  assign n48061 = \P1_P3_DataWidth_reg[1]/NET0131  & ~\P1_P3_PhyAddrPointer_reg[1]/NET0131  ;
  assign n48063 = n16455 & n48061 ;
  assign n48064 = ~n17571 & ~n48063 ;
  assign n48062 = n16456 & n48061 ;
  assign n48065 = n9245 & ~n48062 ;
  assign n48066 = ~n48064 & n48065 ;
  assign n48055 = n16492 & n17571 ;
  assign n48067 = \P1_P3_PhyAddrPointer_reg[6]/NET0131  & ~n36816 ;
  assign n48068 = ~n20500 & ~n48067 ;
  assign n48069 = ~n48055 & n48068 ;
  assign n48070 = ~n48066 & n48069 ;
  assign n48071 = ~n48060 & n48070 ;
  assign n48072 = \P2_P3_PhyAddrPointer_reg[3]/NET0131  & ~n27283 ;
  assign n48073 = ~n45804 & ~n48072 ;
  assign n48074 = n27117 & ~n48073 ;
  assign n48075 = \P2_P3_PhyAddrPointer_reg[3]/NET0131  & ~n36826 ;
  assign n48076 = ~n45820 & ~n48075 ;
  assign n48077 = ~n48074 & n48076 ;
  assign n48078 = n27308 & ~n48077 ;
  assign n48089 = \P2_P3_PhyAddrPointer_reg[3]/NET0131  & n27651 ;
  assign n48086 = ~\P2_P3_PhyAddrPointer_reg[3]/NET0131  & ~n47477 ;
  assign n48087 = ~n47478 & ~n48086 ;
  assign n48088 = n32867 & n48087 ;
  assign n48090 = ~n45790 & ~n48088 ;
  assign n48091 = ~n48089 & n48090 ;
  assign n48079 = \P2_P3_PhyAddrPointer_reg[2]/NET0131  & ~n39862 ;
  assign n48080 = ~\P2_P3_PhyAddrPointer_reg[3]/NET0131  & ~n48079 ;
  assign n48081 = n36835 & ~n39862 ;
  assign n48082 = n27315 & ~n48081 ;
  assign n48083 = ~n48080 & n48082 ;
  assign n48084 = ~n27788 & n36872 ;
  assign n48085 = \P2_P3_PhyAddrPointer_reg[3]/NET0131  & ~n48084 ;
  assign n48092 = ~n48083 & ~n48085 ;
  assign n48093 = n48091 & n48092 ;
  assign n48094 = ~n48078 & n48093 ;
  assign n48095 = \P2_P3_PhyAddrPointer_reg[5]/NET0131  & ~n27283 ;
  assign n48096 = ~n45852 & ~n48095 ;
  assign n48097 = n27117 & ~n48096 ;
  assign n48098 = \P2_P3_PhyAddrPointer_reg[5]/NET0131  & ~n36826 ;
  assign n48099 = ~n45860 & ~n48098 ;
  assign n48100 = ~n48097 & n48099 ;
  assign n48101 = n27308 & ~n48100 ;
  assign n48105 = \P2_P3_PhyAddrPointer_reg[1]/NET0131  & n36837 ;
  assign n48106 = ~\P2_P3_PhyAddrPointer_reg[5]/NET0131  & ~n47480 ;
  assign n48107 = ~n48105 & ~n48106 ;
  assign n48108 = ~n36831 & n48107 ;
  assign n48109 = \P2_P3_PhyAddrPointer_reg[5]/NET0131  & ~n36873 ;
  assign n48102 = ~\P2_P3_PhyAddrPointer_reg[5]/NET0131  & ~n36836 ;
  assign n48103 = ~n36837 & ~n48102 ;
  assign n48104 = n27325 & n48103 ;
  assign n48110 = ~n45837 & ~n48104 ;
  assign n48111 = ~n48109 & n48110 ;
  assign n48112 = ~n48108 & n48111 ;
  assign n48113 = ~n48101 & n48112 ;
  assign n48115 = \P2_P3_PhyAddrPointer_reg[6]/NET0131  & ~n27283 ;
  assign n48116 = ~n44391 & ~n48115 ;
  assign n48117 = n27117 & ~n48116 ;
  assign n48118 = \P2_P3_PhyAddrPointer_reg[6]/NET0131  & ~n36826 ;
  assign n48119 = ~n44402 & ~n48118 ;
  assign n48120 = ~n48117 & n48119 ;
  assign n48121 = n27308 & ~n48120 ;
  assign n48126 = n36837 & ~n39862 ;
  assign n48127 = ~\P2_P3_PhyAddrPointer_reg[6]/NET0131  & ~n48126 ;
  assign n48125 = n36838 & ~n39862 ;
  assign n48128 = n27315 & ~n48125 ;
  assign n48129 = ~n48127 & n48128 ;
  assign n48122 = ~\P2_P3_PhyAddrPointer_reg[6]/NET0131  & ~n48105 ;
  assign n48123 = ~n44156 & ~n48122 ;
  assign n48124 = n32867 & n48123 ;
  assign n48114 = \P2_P3_PhyAddrPointer_reg[6]/NET0131  & ~n36873 ;
  assign n48130 = ~n44385 & ~n48114 ;
  assign n48131 = ~n48124 & n48130 ;
  assign n48132 = ~n48129 & n48131 ;
  assign n48133 = ~n48121 & n48132 ;
  assign n48139 = ~\P2_P1_EBX_reg[26]/NET0131  & ~n46254 ;
  assign n48140 = n25981 & ~n46255 ;
  assign n48141 = ~n48139 & n48140 ;
  assign n48134 = \P2_P1_EBX_reg[26]/NET0131  & ~n20720 ;
  assign n48135 = ~n23823 & ~n48134 ;
  assign n48136 = n25986 & ~n48135 ;
  assign n48137 = ~n25981 & ~n25986 ;
  assign n48138 = \P2_P1_EBX_reg[26]/NET0131  & n48137 ;
  assign n48142 = ~n48136 & ~n48138 ;
  assign n48143 = ~n48141 & n48142 ;
  assign n48144 = n11623 & ~n48143 ;
  assign n48145 = \P2_P1_EBX_reg[26]/NET0131  & ~n21100 ;
  assign n48146 = ~n48144 & ~n48145 ;
  assign n48147 = \P2_P2_EAX_reg[15]/NET0131  & ~n44508 ;
  assign n48183 = ~n32741 & ~n44736 ;
  assign n48184 = \P2_P2_EAX_reg[15]/NET0131  & ~n48183 ;
  assign n48180 = ~\P2_P2_EAX_reg[15]/NET0131  & ~n44718 ;
  assign n48181 = ~n44719 & n44732 ;
  assign n48182 = ~n48180 & n48181 ;
  assign n48159 = \P2_P2_InstQueue_reg[0][7]/NET0131  & n26330 ;
  assign n48157 = \P2_P2_InstQueue_reg[1][7]/NET0131  & n26325 ;
  assign n48148 = \P2_P2_InstQueue_reg[8][7]/NET0131  & n26300 ;
  assign n48149 = \P2_P2_InstQueue_reg[12][7]/NET0131  & n26320 ;
  assign n48164 = ~n48148 & ~n48149 ;
  assign n48174 = ~n48157 & n48164 ;
  assign n48175 = ~n48159 & n48174 ;
  assign n48160 = \P2_P2_InstQueue_reg[15][7]/NET0131  & n26336 ;
  assign n48161 = \P2_P2_InstQueue_reg[7][7]/NET0131  & n26318 ;
  assign n48169 = ~n48160 & ~n48161 ;
  assign n48162 = \P2_P2_InstQueue_reg[4][7]/NET0131  & n26316 ;
  assign n48163 = \P2_P2_InstQueue_reg[3][7]/NET0131  & n26338 ;
  assign n48170 = ~n48162 & ~n48163 ;
  assign n48171 = n48169 & n48170 ;
  assign n48154 = \P2_P2_InstQueue_reg[11][7]/NET0131  & n26304 ;
  assign n48155 = \P2_P2_InstQueue_reg[5][7]/NET0131  & n26332 ;
  assign n48167 = ~n48154 & ~n48155 ;
  assign n48156 = \P2_P2_InstQueue_reg[6][7]/NET0131  & n26307 ;
  assign n48158 = \P2_P2_InstQueue_reg[9][7]/NET0131  & n26327 ;
  assign n48168 = ~n48156 & ~n48158 ;
  assign n48172 = n48167 & n48168 ;
  assign n48150 = \P2_P2_InstQueue_reg[2][7]/NET0131  & n26322 ;
  assign n48151 = \P2_P2_InstQueue_reg[13][7]/NET0131  & n26310 ;
  assign n48165 = ~n48150 & ~n48151 ;
  assign n48152 = \P2_P2_InstQueue_reg[10][7]/NET0131  & n26334 ;
  assign n48153 = \P2_P2_InstQueue_reg[14][7]/NET0131  & n26313 ;
  assign n48166 = ~n48152 & ~n48153 ;
  assign n48173 = n48165 & n48166 ;
  assign n48176 = n48172 & n48173 ;
  assign n48177 = n48171 & n48176 ;
  assign n48178 = n48175 & n48177 ;
  assign n48179 = n44510 & ~n48178 ;
  assign n48185 = ~n26638 & ~n47684 ;
  assign n48186 = ~\P2_P2_EAX_reg[15]/NET0131  & ~n26641 ;
  assign n48187 = \P2_buf2_reg[15]/NET0131  & ~n28013 ;
  assign n48188 = \P2_buf1_reg[15]/NET0131  & n28013 ;
  assign n48189 = ~n48187 & ~n48188 ;
  assign n48190 = n26641 & n48189 ;
  assign n48191 = ~n48186 & ~n48190 ;
  assign n48192 = ~n48185 & n48191 ;
  assign n48193 = ~n48179 & ~n48192 ;
  assign n48194 = ~n48182 & n48193 ;
  assign n48195 = ~n48184 & n48194 ;
  assign n48196 = n26792 & ~n48195 ;
  assign n48197 = ~n48147 & ~n48196 ;
  assign n48212 = ~\P2_P2_EAX_reg[29]/NET0131  & ~n46390 ;
  assign n48213 = n44732 & ~n46391 ;
  assign n48214 = ~n48212 & n48213 ;
  assign n48202 = \P2_P2_EAX_reg[29]/NET0131  & n44736 ;
  assign n48203 = ~n46319 & n46350 ;
  assign n48204 = ~n46351 & ~n48203 ;
  assign n48205 = n44510 & n48204 ;
  assign n48198 = \P2_P2_EAX_reg[29]/NET0131  & ~n26641 ;
  assign n48199 = n26641 & ~n39034 ;
  assign n48200 = ~n48198 & ~n48199 ;
  assign n48201 = n26638 & ~n48200 ;
  assign n48206 = \P2_buf2_reg[13]/NET0131  & ~n28013 ;
  assign n48207 = \P2_buf1_reg[13]/NET0131  & n28013 ;
  assign n48208 = ~n48206 & ~n48207 ;
  assign n48209 = n26641 & ~n48208 ;
  assign n48210 = ~n48198 & ~n48209 ;
  assign n48211 = n26633 & ~n48210 ;
  assign n48215 = ~n48201 & ~n48211 ;
  assign n48216 = ~n48205 & n48215 ;
  assign n48217 = ~n48202 & n48216 ;
  assign n48218 = ~n48214 & n48217 ;
  assign n48219 = n26792 & ~n48218 ;
  assign n48220 = \P2_P2_EAX_reg[29]/NET0131  & ~n44508 ;
  assign n48221 = ~n48219 & ~n48220 ;
  assign n48224 = ~\P2_P2_EBX_reg[26]/NET0131  & ~n46444 ;
  assign n48225 = n26662 & ~n46445 ;
  assign n48226 = ~n48224 & n48225 ;
  assign n48222 = n46416 & n47579 ;
  assign n48223 = \P2_P2_EBX_reg[26]/NET0131  & n46417 ;
  assign n48227 = ~n48222 & ~n48223 ;
  assign n48228 = ~n48226 & n48227 ;
  assign n48229 = n26792 & ~n48228 ;
  assign n48230 = \P2_P2_EBX_reg[26]/NET0131  & ~n44508 ;
  assign n48231 = ~n48229 & ~n48230 ;
  assign n48234 = ~\P1_P3_EBX_reg[26]/NET0131  & ~n46506 ;
  assign n48235 = n9108 & ~n46507 ;
  assign n48236 = ~n48234 & n48235 ;
  assign n48232 = n22379 & n46479 ;
  assign n48233 = \P1_P3_EBX_reg[26]/NET0131  & n46480 ;
  assign n48237 = ~n48232 & ~n48233 ;
  assign n48238 = ~n48236 & n48237 ;
  assign n48239 = n9241 & ~n48238 ;
  assign n48240 = \P1_P3_EBX_reg[26]/NET0131  & ~n16968 ;
  assign n48241 = ~n48239 & ~n48240 ;
  assign n48246 = ~\P1_P1_EBX_reg[26]/NET0131  & ~n46561 ;
  assign n48247 = n26146 & ~n46562 ;
  assign n48248 = ~n48246 & n48247 ;
  assign n48242 = \P1_P1_EBX_reg[26]/NET0131  & ~n15428 ;
  assign n48243 = ~n23577 & ~n48242 ;
  assign n48244 = n26122 & ~n48243 ;
  assign n48245 = \P1_P1_EBX_reg[26]/NET0131  & n46531 ;
  assign n48249 = ~n48244 & ~n48245 ;
  assign n48250 = ~n48248 & n48249 ;
  assign n48251 = n8355 & ~n48250 ;
  assign n48252 = \P1_P1_EBX_reg[26]/NET0131  & ~n15326 ;
  assign n48253 = ~n48251 & ~n48252 ;
  assign n48254 = \P2_P3_EAX_reg[29]/NET0131  & ~n42872 ;
  assign n48265 = ~\P2_P3_EAX_reg[29]/NET0131  & ~n42860 ;
  assign n48266 = n42539 & ~n42861 ;
  assign n48267 = ~n48265 & n48266 ;
  assign n48259 = ~n42542 & ~n45824 ;
  assign n48260 = \P2_P3_EAX_reg[29]/NET0131  & ~n48259 ;
  assign n48261 = ~n42767 & n42798 ;
  assign n48262 = ~n42799 & ~n48261 ;
  assign n48263 = n42538 & n48262 ;
  assign n48256 = ~\P2_buf2_reg[29]/NET0131  & n27227 ;
  assign n48255 = ~\P2_P3_EAX_reg[29]/NET0131  & ~n27227 ;
  assign n48257 = n27186 & ~n48255 ;
  assign n48258 = ~n48256 & n48257 ;
  assign n48264 = \P2_buf2_reg[13]/NET0131  & n45821 ;
  assign n48268 = ~n48258 & ~n48264 ;
  assign n48269 = ~n48263 & n48268 ;
  assign n48270 = ~n48260 & n48269 ;
  assign n48271 = ~n48267 & n48270 ;
  assign n48272 = n27308 & ~n48271 ;
  assign n48273 = ~n48254 & ~n48272 ;
  assign n48276 = ~\P2_P3_EBX_reg[26]/NET0131  & ~n46642 ;
  assign n48277 = n27133 & ~n46643 ;
  assign n48278 = ~n48276 & n48277 ;
  assign n48274 = \P2_P3_EBX_reg[26]/NET0131  & n46615 ;
  assign n48275 = n46614 & n47701 ;
  assign n48279 = ~n48274 & ~n48275 ;
  assign n48280 = ~n48278 & n48279 ;
  assign n48281 = n27308 & ~n48280 ;
  assign n48282 = \P2_P3_EBX_reg[26]/NET0131  & ~n42872 ;
  assign n48283 = ~n48281 & ~n48282 ;
  assign n48284 = \P1_P2_EAX_reg[15]/NET0131  & ~n43212 ;
  assign n48290 = n43164 & ~n43184 ;
  assign n48291 = ~n43167 & ~n48290 ;
  assign n48292 = n25778 & n48291 ;
  assign n48293 = \P1_P2_EAX_reg[15]/NET0131  & ~n48292 ;
  assign n48286 = ~\P1_buf1_reg[15]/NET0131  & n27934 ;
  assign n48285 = ~\P1_buf2_reg[15]/NET0131  & ~n27934 ;
  assign n48287 = ~n25415 & ~n48285 ;
  assign n48288 = ~n48286 & n48287 ;
  assign n48289 = n25875 & n48288 ;
  assign n48305 = \P1_P2_InstQueue_reg[8][7]/NET0131  & n25453 ;
  assign n48298 = \P1_P2_InstQueue_reg[9][7]/NET0131  & n25435 ;
  assign n48294 = \P1_P2_InstQueue_reg[3][7]/NET0131  & n25428 ;
  assign n48295 = \P1_P2_InstQueue_reg[11][7]/NET0131  & n25457 ;
  assign n48310 = ~n48294 & ~n48295 ;
  assign n48320 = ~n48298 & n48310 ;
  assign n48321 = ~n48305 & n48320 ;
  assign n48306 = \P1_P2_InstQueue_reg[15][7]/NET0131  & n25442 ;
  assign n48307 = \P1_P2_InstQueue_reg[2][7]/NET0131  & n25425 ;
  assign n48315 = ~n48306 & ~n48307 ;
  assign n48308 = \P1_P2_InstQueue_reg[5][7]/NET0131  & n25437 ;
  assign n48309 = \P1_P2_InstQueue_reg[4][7]/NET0131  & n25444 ;
  assign n48316 = ~n48308 & ~n48309 ;
  assign n48317 = n48315 & n48316 ;
  assign n48301 = \P1_P2_InstQueue_reg[12][7]/NET0131  & n25440 ;
  assign n48302 = \P1_P2_InstQueue_reg[10][7]/NET0131  & n25455 ;
  assign n48313 = ~n48301 & ~n48302 ;
  assign n48303 = \P1_P2_InstQueue_reg[1][7]/NET0131  & n25446 ;
  assign n48304 = \P1_P2_InstQueue_reg[14][7]/NET0131  & n25422 ;
  assign n48314 = ~n48303 & ~n48304 ;
  assign n48318 = n48313 & n48314 ;
  assign n48296 = \P1_P2_InstQueue_reg[6][7]/NET0131  & n25461 ;
  assign n48297 = \P1_P2_InstQueue_reg[0][7]/NET0131  & n25431 ;
  assign n48311 = ~n48296 & ~n48297 ;
  assign n48299 = \P1_P2_InstQueue_reg[13][7]/NET0131  & n25459 ;
  assign n48300 = \P1_P2_InstQueue_reg[7][7]/NET0131  & n25449 ;
  assign n48312 = ~n48299 & ~n48300 ;
  assign n48319 = n48311 & n48312 ;
  assign n48322 = n48318 & n48319 ;
  assign n48323 = n48317 & n48322 ;
  assign n48324 = n48321 & n48323 ;
  assign n48325 = n42875 & ~n48324 ;
  assign n48326 = ~\P1_P2_EAX_reg[15]/NET0131  & n43164 ;
  assign n48327 = n43184 & n48326 ;
  assign n48328 = ~n48325 & ~n48327 ;
  assign n48329 = ~n48289 & n48328 ;
  assign n48330 = ~n48293 & n48329 ;
  assign n48331 = n25918 & ~n48330 ;
  assign n48332 = ~n48284 & ~n48331 ;
  assign n48333 = \P1_P2_EAX_reg[29]/NET0131  & ~n43212 ;
  assign n48334 = n43164 & ~n43198 ;
  assign n48335 = ~n43167 & ~n48334 ;
  assign n48336 = \P1_P2_EAX_reg[29]/NET0131  & ~n48335 ;
  assign n48350 = ~\P1_P2_EAX_reg[29]/NET0131  & n46671 ;
  assign n48341 = ~n43098 & n43129 ;
  assign n48342 = ~n43130 & ~n48341 ;
  assign n48343 = n42875 & n48342 ;
  assign n48337 = \P1_P2_EAX_reg[29]/NET0131  & ~n25773 ;
  assign n48338 = n25773 & ~n29868 ;
  assign n48339 = ~n48337 & ~n48338 ;
  assign n48340 = n25774 & ~n48339 ;
  assign n48344 = ~\P1_buf2_reg[13]/NET0131  & ~n27934 ;
  assign n48345 = ~\P1_buf1_reg[13]/NET0131  & n27934 ;
  assign n48346 = ~n48344 & ~n48345 ;
  assign n48347 = n25773 & n48346 ;
  assign n48348 = ~n48337 & ~n48347 ;
  assign n48349 = n25776 & ~n48348 ;
  assign n48351 = ~n48340 & ~n48349 ;
  assign n48352 = ~n48343 & n48351 ;
  assign n48353 = ~n48350 & n48352 ;
  assign n48354 = ~n48336 & n48353 ;
  assign n48355 = n25918 & ~n48354 ;
  assign n48356 = ~n48333 & ~n48355 ;
  assign n48362 = ~\P1_P2_EBX_reg[26]/NET0131  & ~n46722 ;
  assign n48363 = n25803 & ~n46723 ;
  assign n48364 = ~n48362 & n48363 ;
  assign n48357 = \P1_P2_EBX_reg[26]/NET0131  & ~n25747 ;
  assign n48358 = ~n47722 & ~n48357 ;
  assign n48359 = n25738 & ~n48358 ;
  assign n48360 = ~n25738 & ~n25803 ;
  assign n48361 = \P1_P2_EBX_reg[26]/NET0131  & n48360 ;
  assign n48365 = ~n48359 & ~n48361 ;
  assign n48366 = ~n48364 & n48365 ;
  assign n48367 = n25918 & ~n48366 ;
  assign n48368 = \P1_P2_EBX_reg[26]/NET0131  & ~n43212 ;
  assign n48369 = ~n48367 & ~n48368 ;
  assign n48455 = ~\P1_P2_PhyAddrPointer_reg[0]/NET0131  & n43518 ;
  assign n48456 = n36604 & n48455 ;
  assign n48457 = n39370 & n48456 ;
  assign n48458 = \P1_P2_PhyAddrPointer_reg[21]/NET0131  & n48457 ;
  assign n48459 = n37921 & n48458 ;
  assign n48460 = ~n36628 & ~n48459 ;
  assign n48462 = ~n37923 & n48460 ;
  assign n48461 = n37923 & ~n48460 ;
  assign n48463 = ~\P1_P2_DataWidth_reg[1]/NET0131  & ~n48461 ;
  assign n48464 = ~n48462 & n48463 ;
  assign n48454 = \P1_P2_DataWidth_reg[1]/NET0131  & ~\P1_P2_rEIP_reg[30]/NET0131  ;
  assign n48465 = n25928 & ~n48454 ;
  assign n48466 = ~n48464 & n48465 ;
  assign n48407 = ~\P1_P2_EBX_reg[0]/NET0131  & ~\P1_P2_EBX_reg[1]/NET0131  ;
  assign n48408 = ~\P1_P2_EBX_reg[2]/NET0131  & n48407 ;
  assign n48409 = ~\P1_P2_EBX_reg[3]/NET0131  & n48408 ;
  assign n48410 = ~\P1_P2_EBX_reg[4]/NET0131  & n48409 ;
  assign n48411 = ~\P1_P2_EBX_reg[5]/NET0131  & n48410 ;
  assign n48412 = ~\P1_P2_EBX_reg[6]/NET0131  & n48411 ;
  assign n48413 = ~\P1_P2_EBX_reg[7]/NET0131  & n48412 ;
  assign n48414 = ~\P1_P2_EBX_reg[8]/NET0131  & n48413 ;
  assign n48415 = ~\P1_P2_EBX_reg[9]/NET0131  & n48414 ;
  assign n48416 = ~\P1_P2_EBX_reg[10]/NET0131  & n48415 ;
  assign n48417 = ~\P1_P2_EBX_reg[11]/NET0131  & n48416 ;
  assign n48418 = ~\P1_P2_EBX_reg[12]/NET0131  & n48417 ;
  assign n48419 = ~\P1_P2_EBX_reg[13]/NET0131  & n48418 ;
  assign n48420 = ~\P1_P2_EBX_reg[14]/NET0131  & n48419 ;
  assign n48421 = ~\P1_P2_EBX_reg[15]/NET0131  & n48420 ;
  assign n48422 = ~\P1_P2_EBX_reg[16]/NET0131  & n48421 ;
  assign n48423 = ~\P1_P2_EBX_reg[17]/NET0131  & n48422 ;
  assign n48424 = ~\P1_P2_EBX_reg[18]/NET0131  & n48423 ;
  assign n48425 = ~\P1_P2_EBX_reg[19]/NET0131  & n48424 ;
  assign n48426 = ~\P1_P2_EBX_reg[20]/NET0131  & n48425 ;
  assign n48427 = ~\P1_P2_EBX_reg[21]/NET0131  & n48426 ;
  assign n48428 = ~\P1_P2_EBX_reg[22]/NET0131  & n48427 ;
  assign n48429 = ~\P1_P2_EBX_reg[23]/NET0131  & n48428 ;
  assign n48430 = ~\P1_P2_EBX_reg[24]/NET0131  & n48429 ;
  assign n48431 = ~\P1_P2_EBX_reg[25]/NET0131  & n48430 ;
  assign n48432 = ~\P1_P2_EBX_reg[26]/NET0131  & n48431 ;
  assign n48433 = ~\P1_P2_EBX_reg[27]/NET0131  & n48432 ;
  assign n48434 = ~\P1_P2_EBX_reg[28]/NET0131  & n48433 ;
  assign n48435 = ~\P1_P2_EBX_reg[29]/NET0131  & n48434 ;
  assign n48436 = \P1_P2_EBX_reg[31]/NET0131  & ~n48435 ;
  assign n48438 = ~\P1_P2_EBX_reg[30]/NET0131  & n48436 ;
  assign n48373 = ~\P1_P2_DataWidth_reg[1]/NET0131  & ~n25415 ;
  assign n48437 = \P1_P2_EBX_reg[30]/NET0131  & ~n48436 ;
  assign n48439 = ~n48373 & ~n48437 ;
  assign n48440 = ~n48438 & n48439 ;
  assign n48374 = \P1_P2_rEIP_reg[23]/NET0131  & \P1_P2_rEIP_reg[24]/NET0131  ;
  assign n48375 = \P1_P2_rEIP_reg[25]/NET0131  & n48374 ;
  assign n48376 = \P1_P2_rEIP_reg[26]/NET0131  & n48375 ;
  assign n48377 = \P1_P2_rEIP_reg[19]/NET0131  & \P1_P2_rEIP_reg[20]/NET0131  ;
  assign n48378 = \P1_P2_rEIP_reg[21]/NET0131  & n48377 ;
  assign n48379 = \P1_P2_rEIP_reg[22]/NET0131  & n48378 ;
  assign n48380 = \P1_P2_rEIP_reg[1]/NET0131  & \P1_P2_rEIP_reg[2]/NET0131  ;
  assign n48381 = \P1_P2_rEIP_reg[3]/NET0131  & n48380 ;
  assign n48382 = \P1_P2_rEIP_reg[4]/NET0131  & n48381 ;
  assign n48383 = \P1_P2_rEIP_reg[5]/NET0131  & n48382 ;
  assign n48384 = \P1_P2_rEIP_reg[6]/NET0131  & n48383 ;
  assign n48385 = \P1_P2_rEIP_reg[7]/NET0131  & n48384 ;
  assign n48386 = \P1_P2_rEIP_reg[8]/NET0131  & n48385 ;
  assign n48387 = \P1_P2_rEIP_reg[16]/NET0131  & \P1_P2_rEIP_reg[17]/NET0131  ;
  assign n48388 = \P1_P2_rEIP_reg[18]/NET0131  & n48387 ;
  assign n48389 = \P1_P2_rEIP_reg[15]/NET0131  & n48388 ;
  assign n48390 = \P1_P2_rEIP_reg[12]/NET0131  & \P1_P2_rEIP_reg[13]/NET0131  ;
  assign n48391 = \P1_P2_rEIP_reg[14]/NET0131  & n48390 ;
  assign n48392 = \P1_P2_rEIP_reg[10]/NET0131  & \P1_P2_rEIP_reg[11]/NET0131  ;
  assign n48393 = \P1_P2_rEIP_reg[9]/NET0131  & n48392 ;
  assign n48394 = n48391 & n48393 ;
  assign n48395 = n48389 & n48394 ;
  assign n48396 = n48386 & n48395 ;
  assign n48397 = n48379 & n48396 ;
  assign n48398 = n48376 & n48397 ;
  assign n48399 = \P1_P2_rEIP_reg[27]/NET0131  & n48398 ;
  assign n48400 = \P1_P2_rEIP_reg[28]/NET0131  & \P1_P2_rEIP_reg[29]/NET0131  ;
  assign n48401 = n48399 & n48400 ;
  assign n48402 = ~\P1_P2_rEIP_reg[30]/NET0131  & ~n48401 ;
  assign n48403 = \P1_P2_rEIP_reg[30]/NET0131  & n48400 ;
  assign n48404 = n48399 & n48403 ;
  assign n48405 = ~n48402 & ~n48404 ;
  assign n48406 = n48373 & ~n48405 ;
  assign n48441 = n25846 & ~n48406 ;
  assign n48442 = ~n48440 & n48441 ;
  assign n48371 = ~n25770 & ~n25786 ;
  assign n48372 = \P1_P2_rEIP_reg[30]/NET0131  & ~n48371 ;
  assign n48443 = ~n25768 & n48373 ;
  assign n48445 = ~n48405 & n48443 ;
  assign n48444 = ~\P1_P2_EBX_reg[30]/NET0131  & ~n48443 ;
  assign n48446 = n47570 & ~n48444 ;
  assign n48447 = ~n48445 & n48446 ;
  assign n48448 = ~n48372 & ~n48447 ;
  assign n48449 = ~n48442 & n48448 ;
  assign n48450 = n25918 & ~n48449 ;
  assign n48370 = \P1_P2_PhyAddrPointer_reg[30]/NET0131  & n27675 ;
  assign n48451 = ~n27608 & ~n27898 ;
  assign n48452 = n39351 & n48451 ;
  assign n48453 = \P1_P2_rEIP_reg[30]/NET0131  & ~n48452 ;
  assign n48467 = ~n48370 & ~n48453 ;
  assign n48468 = ~n48450 & n48467 ;
  assign n48469 = ~n48466 & n48468 ;
  assign n48471 = ~n26158 & n35952 ;
  assign n48472 = \P1_P1_Datao_reg[24]/NET0131  & ~n26162 ;
  assign n48473 = ~n48471 & ~n48472 ;
  assign n48474 = n8355 & ~n48473 ;
  assign n48470 = \P1_P1_uWord_reg[8]/NET0131  & n27790 ;
  assign n48477 = ~n8282 & ~n15324 ;
  assign n48475 = ~n8286 & ~n8348 ;
  assign n48476 = ~n8354 & ~n48475 ;
  assign n48478 = ~n15322 & ~n48476 ;
  assign n48479 = n48477 & n48478 ;
  assign n48480 = \P1_P1_Datao_reg[24]/NET0131  & ~n48479 ;
  assign n48481 = ~n48470 & ~n48480 ;
  assign n48482 = ~n48474 & n48481 ;
  assign n48484 = ~n26158 & n27597 ;
  assign n48485 = \P1_P1_Datao_reg[28]/NET0131  & ~n26162 ;
  assign n48486 = ~n48484 & ~n48485 ;
  assign n48487 = n8355 & ~n48486 ;
  assign n48483 = \P1_P1_uWord_reg[12]/NET0131  & n27790 ;
  assign n48488 = \P1_P1_Datao_reg[28]/NET0131  & ~n48479 ;
  assign n48489 = ~n48483 & ~n48488 ;
  assign n48490 = ~n48487 & n48489 ;
  assign n48493 = n26644 & n26650 ;
  assign n48494 = n26698 & ~n48493 ;
  assign n48495 = ~\P2_P2_EAX_reg[24]/NET0131  & ~n47667 ;
  assign n48496 = ~n47668 & ~n48495 ;
  assign n48497 = ~n26650 & ~n48496 ;
  assign n48498 = n26786 & ~n48497 ;
  assign n48499 = n48494 & ~n48498 ;
  assign n48500 = \P2_P2_Datao_reg[24]/NET0131  & ~n48499 ;
  assign n48501 = n26643 & n48496 ;
  assign n48502 = n26692 & n48501 ;
  assign n48503 = ~n48500 & ~n48502 ;
  assign n48504 = n26792 & ~n48503 ;
  assign n48491 = ~\P2_P2_State2_reg[0]/NET0131  & n27614 ;
  assign n48492 = \P2_P2_uWord_reg[8]/NET0131  & n48491 ;
  assign n48505 = \P2_P2_State2_reg[1]/NET0131  & \P2_P2_State2_reg[3]/NET0131  ;
  assign n48506 = \P2_P2_State2_reg[2]/NET0131  & ~n27977 ;
  assign n48507 = ~n48505 & ~n48506 ;
  assign n48508 = ~n27615 & ~n48507 ;
  assign n48509 = \P2_P2_Datao_reg[24]/NET0131  & ~n48508 ;
  assign n48510 = ~n48492 & ~n48509 ;
  assign n48511 = ~n48504 & n48510 ;
  assign n48513 = ~n26650 & ~n47674 ;
  assign n48514 = n26786 & ~n48513 ;
  assign n48515 = n48494 & ~n48514 ;
  assign n48516 = \P2_P2_Datao_reg[28]/NET0131  & ~n48515 ;
  assign n48517 = n26692 & n47675 ;
  assign n48518 = ~n48516 & ~n48517 ;
  assign n48519 = n26792 & ~n48518 ;
  assign n48512 = \P2_P2_uWord_reg[12]/NET0131  & n48491 ;
  assign n48520 = \P2_P2_Datao_reg[28]/NET0131  & ~n48508 ;
  assign n48521 = ~n48512 & ~n48520 ;
  assign n48522 = ~n48519 & n48521 ;
  assign n48525 = \P2_P3_Datao_reg[24]/NET0131  & ~n27223 ;
  assign n48526 = \P2_P3_EAX_reg[20]/NET0131  & n47776 ;
  assign n48527 = \P2_P3_EAX_reg[21]/NET0131  & n48526 ;
  assign n48528 = \P2_P3_EAX_reg[22]/NET0131  & n48527 ;
  assign n48529 = \P2_P3_EAX_reg[23]/NET0131  & n48528 ;
  assign n48530 = ~\P2_P3_EAX_reg[24]/NET0131  & ~n48529 ;
  assign n48531 = n42855 & n47775 ;
  assign n48532 = n27121 & ~n48531 ;
  assign n48533 = ~n48530 & n48532 ;
  assign n48534 = n27178 & n48533 ;
  assign n48535 = ~n48525 & ~n48534 ;
  assign n48536 = n27308 & ~n48535 ;
  assign n48523 = ~\P2_P3_State2_reg[0]/NET0131  & n27656 ;
  assign n48524 = \P2_P3_uWord_reg[8]/NET0131  & n48523 ;
  assign n48538 = \P2_P3_State2_reg[1]/NET0131  & n27306 ;
  assign n48537 = n27317 & ~n27653 ;
  assign n48539 = ~n27649 & ~n48537 ;
  assign n48540 = ~n48538 & n48539 ;
  assign n48541 = \P2_P3_Datao_reg[24]/NET0131  & ~n48540 ;
  assign n48542 = ~n48524 & ~n48541 ;
  assign n48543 = ~n48536 & n48542 ;
  assign n48545 = \P2_P3_Datao_reg[28]/NET0131  & ~n27223 ;
  assign n48546 = n27303 & n47781 ;
  assign n48547 = ~n48545 & ~n48546 ;
  assign n48548 = n27308 & ~n48547 ;
  assign n48544 = \P2_P3_uWord_reg[12]/NET0131  & n48523 ;
  assign n48549 = \P2_P3_Datao_reg[28]/NET0131  & ~n48540 ;
  assign n48550 = ~n48544 & ~n48549 ;
  assign n48551 = ~n48548 & n48550 ;
  assign n48553 = n25762 & n25768 ;
  assign n48554 = n25877 & ~n48553 ;
  assign n48555 = ~\P1_P2_EAX_reg[24]/NET0131  & ~n47554 ;
  assign n48556 = ~n47555 & ~n48555 ;
  assign n48557 = ~n25768 & ~n48556 ;
  assign n48558 = n47570 & ~n48557 ;
  assign n48559 = n48554 & ~n48558 ;
  assign n48560 = \P1_P2_Datao_reg[24]/NET0131  & ~n48559 ;
  assign n48561 = n25757 & n48556 ;
  assign n48562 = n25841 & n48561 ;
  assign n48563 = ~n48560 & ~n48562 ;
  assign n48564 = n25918 & ~n48563 ;
  assign n48552 = \P1_P2_uWord_reg[8]/NET0131  & n25922 ;
  assign n48565 = ~n27898 & ~n43208 ;
  assign n48566 = n43210 & n48565 ;
  assign n48567 = \P1_P2_Datao_reg[24]/NET0131  & ~n48566 ;
  assign n48568 = ~n48552 & ~n48567 ;
  assign n48569 = ~n48564 & n48568 ;
  assign n48571 = ~n25768 & ~n47561 ;
  assign n48572 = n47570 & ~n48571 ;
  assign n48573 = n48554 & ~n48572 ;
  assign n48574 = \P1_P2_Datao_reg[28]/NET0131  & ~n48573 ;
  assign n48575 = n25841 & n47562 ;
  assign n48576 = ~n48574 & ~n48575 ;
  assign n48577 = n25918 & ~n48576 ;
  assign n48570 = \P1_P2_uWord_reg[12]/NET0131  & n25922 ;
  assign n48578 = \P1_P2_Datao_reg[28]/NET0131  & ~n48566 ;
  assign n48579 = ~n48570 & ~n48578 ;
  assign n48580 = ~n48577 & n48579 ;
  assign n48583 = n25951 & n25958 ;
  assign n48584 = n25953 & ~n48583 ;
  assign n48585 = ~n25958 & ~n35912 ;
  assign n48586 = n24899 & ~n48585 ;
  assign n48587 = n48584 & ~n48586 ;
  assign n48588 = \P2_P1_Datao_reg[24]/NET0131  & ~n48587 ;
  assign n48589 = n26006 & n35913 ;
  assign n48590 = ~n48588 & ~n48589 ;
  assign n48591 = n11623 & ~n48590 ;
  assign n48581 = ~\P2_P1_State2_reg[0]/NET0131  & n11621 ;
  assign n48582 = \P2_P1_uWord_reg[8]/NET0131  & n48581 ;
  assign n48592 = \P2_P1_State2_reg[1]/NET0131  & n11622 ;
  assign n48593 = ~n11615 & ~n48592 ;
  assign n48594 = n12341 & n48593 ;
  assign n48595 = \P2_P1_Datao_reg[24]/NET0131  & ~n48594 ;
  assign n48596 = ~n48582 & ~n48595 ;
  assign n48597 = ~n48591 & n48596 ;
  assign n48599 = ~n25958 & ~n27732 ;
  assign n48600 = n24899 & ~n48599 ;
  assign n48601 = n48584 & ~n48600 ;
  assign n48602 = \P2_P1_Datao_reg[28]/NET0131  & ~n48601 ;
  assign n48603 = n26006 & n27733 ;
  assign n48604 = ~n48602 & ~n48603 ;
  assign n48605 = n11623 & ~n48604 ;
  assign n48598 = \P2_P1_uWord_reg[12]/NET0131  & n48581 ;
  assign n48606 = \P2_P1_Datao_reg[28]/NET0131  & ~n48594 ;
  assign n48607 = ~n48598 & ~n48606 ;
  assign n48608 = ~n48605 & n48607 ;
  assign n48611 = ~\P1_P2_EBX_reg[29]/NET0131  & ~n46736 ;
  assign n48612 = n25803 & ~n46737 ;
  assign n48613 = ~n48611 & n48612 ;
  assign n48609 = n46694 & n48342 ;
  assign n48610 = \P1_P2_EBX_reg[29]/NET0131  & n46695 ;
  assign n48614 = ~n48609 & ~n48610 ;
  assign n48615 = ~n48613 & n48614 ;
  assign n48616 = n25918 & ~n48615 ;
  assign n48617 = \P1_P2_EBX_reg[29]/NET0131  & ~n43212 ;
  assign n48618 = ~n48616 & ~n48617 ;
  assign n48619 = \P2_P1_EAX_reg[2]/NET0131  & ~n27438 ;
  assign n48621 = ~n21069 & n24838 ;
  assign n48620 = n20728 & ~n31719 ;
  assign n48622 = ~\P2_P1_EAX_reg[2]/NET0131  & ~n21023 ;
  assign n48623 = ~n21024 & ~n48622 ;
  assign n48624 = n21022 & n48623 ;
  assign n48625 = ~n48620 & ~n48624 ;
  assign n48626 = ~n48621 & n48625 ;
  assign n48627 = n11623 & ~n48626 ;
  assign n48628 = ~n48619 & ~n48627 ;
  assign n48631 = ~\P2_P1_EBX_reg[29]/NET0131  & ~n46267 ;
  assign n48632 = n25981 & ~n46268 ;
  assign n48633 = ~n48631 & n48632 ;
  assign n48629 = n23165 & n46225 ;
  assign n48630 = \P2_P1_EBX_reg[29]/NET0131  & n46227 ;
  assign n48634 = ~n48629 & ~n48630 ;
  assign n48635 = ~n48633 & n48634 ;
  assign n48636 = n11623 & ~n48635 ;
  assign n48637 = \P2_P1_EBX_reg[29]/NET0131  & ~n21100 ;
  assign n48638 = ~n48636 & ~n48637 ;
  assign n48639 = \P2_P1_uWord_reg[4]/NET0131  & ~n25156 ;
  assign n48640 = ~\P2_P1_EAX_reg[20]/NET0131  & ~n27391 ;
  assign n48641 = ~n27392 & ~n48640 ;
  assign n48642 = n24899 & n48641 ;
  assign n48643 = ~n44482 & ~n48642 ;
  assign n48644 = n11623 & ~n48643 ;
  assign n48645 = ~n48639 & ~n48644 ;
  assign n48646 = \P1_P1_EAX_reg[2]/NET0131  & ~n27551 ;
  assign n48648 = n7947 & n24342 ;
  assign n48647 = n22818 & ~n33731 ;
  assign n48649 = ~\P1_P1_EAX_reg[2]/NET0131  & ~n15388 ;
  assign n48650 = ~n15389 & ~n48649 ;
  assign n48651 = n15377 & n48650 ;
  assign n48652 = ~n48647 & ~n48651 ;
  assign n48653 = ~n48648 & n48652 ;
  assign n48654 = n8355 & ~n48653 ;
  assign n48655 = ~n48646 & ~n48654 ;
  assign n48656 = \P1_P2_uWord_reg[8]/NET0131  & ~n47529 ;
  assign n48657 = \P1_buf2_reg[8]/NET0131  & ~n27934 ;
  assign n48658 = \P1_buf1_reg[8]/NET0131  & n27934 ;
  assign n48659 = ~n48657 & ~n48658 ;
  assign n48660 = n25776 & ~n48659 ;
  assign n48661 = ~n25415 & n48660 ;
  assign n48662 = ~n48561 & ~n48661 ;
  assign n48663 = ~n25770 & ~n48662 ;
  assign n48664 = \P1_P2_uWord_reg[8]/NET0131  & ~n47572 ;
  assign n48665 = ~n48663 & ~n48664 ;
  assign n48666 = n25918 & ~n48665 ;
  assign n48667 = ~n48656 & ~n48666 ;
  assign n48668 = n26792 & ~n46402 ;
  assign n48669 = n44508 & ~n48668 ;
  assign n48670 = \P2_P2_EAX_reg[10]/NET0131  & ~n48669 ;
  assign n48703 = ~n26639 & n47591 ;
  assign n48682 = \P2_P2_InstQueue_reg[0][2]/NET0131  & n26330 ;
  assign n48680 = \P2_P2_InstQueue_reg[1][2]/NET0131  & n26325 ;
  assign n48671 = \P2_P2_InstQueue_reg[8][2]/NET0131  & n26300 ;
  assign n48672 = \P2_P2_InstQueue_reg[12][2]/NET0131  & n26320 ;
  assign n48687 = ~n48671 & ~n48672 ;
  assign n48697 = ~n48680 & n48687 ;
  assign n48698 = ~n48682 & n48697 ;
  assign n48683 = \P2_P2_InstQueue_reg[15][2]/NET0131  & n26336 ;
  assign n48684 = \P2_P2_InstQueue_reg[7][2]/NET0131  & n26318 ;
  assign n48692 = ~n48683 & ~n48684 ;
  assign n48685 = \P2_P2_InstQueue_reg[4][2]/NET0131  & n26316 ;
  assign n48686 = \P2_P2_InstQueue_reg[3][2]/NET0131  & n26338 ;
  assign n48693 = ~n48685 & ~n48686 ;
  assign n48694 = n48692 & n48693 ;
  assign n48677 = \P2_P2_InstQueue_reg[11][2]/NET0131  & n26304 ;
  assign n48678 = \P2_P2_InstQueue_reg[5][2]/NET0131  & n26332 ;
  assign n48690 = ~n48677 & ~n48678 ;
  assign n48679 = \P2_P2_InstQueue_reg[6][2]/NET0131  & n26307 ;
  assign n48681 = \P2_P2_InstQueue_reg[9][2]/NET0131  & n26327 ;
  assign n48691 = ~n48679 & ~n48681 ;
  assign n48695 = n48690 & n48691 ;
  assign n48673 = \P2_P2_InstQueue_reg[2][2]/NET0131  & n26322 ;
  assign n48674 = \P2_P2_InstQueue_reg[13][2]/NET0131  & n26310 ;
  assign n48688 = ~n48673 & ~n48674 ;
  assign n48675 = \P2_P2_InstQueue_reg[10][2]/NET0131  & n26334 ;
  assign n48676 = \P2_P2_InstQueue_reg[14][2]/NET0131  & n26313 ;
  assign n48689 = ~n48675 & ~n48676 ;
  assign n48696 = n48688 & n48689 ;
  assign n48699 = n48695 & n48696 ;
  assign n48700 = n48694 & n48699 ;
  assign n48701 = n48698 & n48700 ;
  assign n48702 = n44510 & ~n48701 ;
  assign n48704 = ~\P2_P2_EAX_reg[10]/NET0131  & ~n44713 ;
  assign n48705 = ~n44714 & ~n48704 ;
  assign n48706 = n44732 & n48705 ;
  assign n48707 = ~n48702 & ~n48706 ;
  assign n48708 = ~n48703 & n48707 ;
  assign n48709 = n26792 & ~n48708 ;
  assign n48710 = ~n48670 & ~n48709 ;
  assign n48711 = \P2_P2_EAX_reg[11]/NET0131  & ~n48669 ;
  assign n48744 = ~n26639 & n44744 ;
  assign n48723 = \P2_P2_InstQueue_reg[0][3]/NET0131  & n26330 ;
  assign n48721 = \P2_P2_InstQueue_reg[1][3]/NET0131  & n26325 ;
  assign n48712 = \P2_P2_InstQueue_reg[8][3]/NET0131  & n26300 ;
  assign n48713 = \P2_P2_InstQueue_reg[3][3]/NET0131  & n26338 ;
  assign n48728 = ~n48712 & ~n48713 ;
  assign n48738 = ~n48721 & n48728 ;
  assign n48739 = ~n48723 & n48738 ;
  assign n48724 = \P2_P2_InstQueue_reg[10][3]/NET0131  & n26334 ;
  assign n48725 = \P2_P2_InstQueue_reg[15][3]/NET0131  & n26336 ;
  assign n48733 = ~n48724 & ~n48725 ;
  assign n48726 = \P2_P2_InstQueue_reg[14][3]/NET0131  & n26313 ;
  assign n48727 = \P2_P2_InstQueue_reg[2][3]/NET0131  & n26322 ;
  assign n48734 = ~n48726 & ~n48727 ;
  assign n48735 = n48733 & n48734 ;
  assign n48718 = \P2_P2_InstQueue_reg[13][3]/NET0131  & n26310 ;
  assign n48719 = \P2_P2_InstQueue_reg[5][3]/NET0131  & n26332 ;
  assign n48731 = ~n48718 & ~n48719 ;
  assign n48720 = \P2_P2_InstQueue_reg[7][3]/NET0131  & n26318 ;
  assign n48722 = \P2_P2_InstQueue_reg[9][3]/NET0131  & n26327 ;
  assign n48732 = ~n48720 & ~n48722 ;
  assign n48736 = n48731 & n48732 ;
  assign n48714 = \P2_P2_InstQueue_reg[6][3]/NET0131  & n26307 ;
  assign n48715 = \P2_P2_InstQueue_reg[4][3]/NET0131  & n26316 ;
  assign n48729 = ~n48714 & ~n48715 ;
  assign n48716 = \P2_P2_InstQueue_reg[11][3]/NET0131  & n26304 ;
  assign n48717 = \P2_P2_InstQueue_reg[12][3]/NET0131  & n26320 ;
  assign n48730 = ~n48716 & ~n48717 ;
  assign n48737 = n48729 & n48730 ;
  assign n48740 = n48736 & n48737 ;
  assign n48741 = n48735 & n48740 ;
  assign n48742 = n48739 & n48741 ;
  assign n48743 = n44510 & ~n48742 ;
  assign n48745 = ~\P2_P2_EAX_reg[11]/NET0131  & ~n44714 ;
  assign n48746 = ~n44715 & ~n48745 ;
  assign n48747 = n44732 & n48746 ;
  assign n48748 = ~n48743 & ~n48747 ;
  assign n48749 = ~n48744 & n48748 ;
  assign n48750 = n26792 & ~n48749 ;
  assign n48751 = ~n48711 & ~n48750 ;
  assign n48752 = \P2_P2_EAX_reg[12]/NET0131  & ~n44508 ;
  assign n48753 = ~n44716 & n44732 ;
  assign n48755 = ~n44736 & ~n48753 ;
  assign n48756 = \P2_P2_EAX_reg[12]/NET0131  & ~n48755 ;
  assign n48789 = n26641 & ~n47679 ;
  assign n48790 = \P2_P2_EAX_reg[12]/NET0131  & ~n26641 ;
  assign n48791 = ~n48789 & ~n48790 ;
  assign n48792 = ~n26639 & ~n48791 ;
  assign n48754 = n44715 & n48753 ;
  assign n48768 = \P2_P2_InstQueue_reg[0][4]/NET0131  & n26330 ;
  assign n48766 = \P2_P2_InstQueue_reg[1][4]/NET0131  & n26325 ;
  assign n48757 = \P2_P2_InstQueue_reg[8][4]/NET0131  & n26300 ;
  assign n48758 = \P2_P2_InstQueue_reg[7][4]/NET0131  & n26318 ;
  assign n48773 = ~n48757 & ~n48758 ;
  assign n48783 = ~n48766 & n48773 ;
  assign n48784 = ~n48768 & n48783 ;
  assign n48769 = \P2_P2_InstQueue_reg[3][4]/NET0131  & n26338 ;
  assign n48770 = \P2_P2_InstQueue_reg[6][4]/NET0131  & n26307 ;
  assign n48778 = ~n48769 & ~n48770 ;
  assign n48771 = \P2_P2_InstQueue_reg[10][4]/NET0131  & n26334 ;
  assign n48772 = \P2_P2_InstQueue_reg[2][4]/NET0131  & n26322 ;
  assign n48779 = ~n48771 & ~n48772 ;
  assign n48780 = n48778 & n48779 ;
  assign n48763 = \P2_P2_InstQueue_reg[4][4]/NET0131  & n26316 ;
  assign n48764 = \P2_P2_InstQueue_reg[11][4]/NET0131  & n26304 ;
  assign n48776 = ~n48763 & ~n48764 ;
  assign n48765 = \P2_P2_InstQueue_reg[15][4]/NET0131  & n26336 ;
  assign n48767 = \P2_P2_InstQueue_reg[9][4]/NET0131  & n26327 ;
  assign n48777 = ~n48765 & ~n48767 ;
  assign n48781 = n48776 & n48777 ;
  assign n48759 = \P2_P2_InstQueue_reg[5][4]/NET0131  & n26332 ;
  assign n48760 = \P2_P2_InstQueue_reg[12][4]/NET0131  & n26320 ;
  assign n48774 = ~n48759 & ~n48760 ;
  assign n48761 = \P2_P2_InstQueue_reg[14][4]/NET0131  & n26313 ;
  assign n48762 = \P2_P2_InstQueue_reg[13][4]/NET0131  & n26310 ;
  assign n48775 = ~n48761 & ~n48762 ;
  assign n48782 = n48774 & n48775 ;
  assign n48785 = n48781 & n48782 ;
  assign n48786 = n48780 & n48785 ;
  assign n48787 = n48784 & n48786 ;
  assign n48788 = n44510 & ~n48787 ;
  assign n48793 = ~n48754 & ~n48788 ;
  assign n48794 = ~n48792 & n48793 ;
  assign n48795 = ~n48756 & n48794 ;
  assign n48796 = n26792 & ~n48795 ;
  assign n48797 = ~n48752 & ~n48796 ;
  assign n48798 = \P2_P2_EAX_reg[13]/NET0131  & ~n44508 ;
  assign n48801 = \P2_P2_EAX_reg[13]/NET0131  & ~n48755 ;
  assign n48834 = \P2_P2_EAX_reg[13]/NET0131  & ~n26641 ;
  assign n48835 = ~n48209 & ~n48834 ;
  assign n48836 = ~n26639 & ~n48835 ;
  assign n48799 = ~\P2_P2_EAX_reg[13]/NET0131  & n44716 ;
  assign n48800 = n44732 & n48799 ;
  assign n48813 = \P2_P2_InstQueue_reg[0][5]/NET0131  & n26330 ;
  assign n48811 = \P2_P2_InstQueue_reg[1][5]/NET0131  & n26325 ;
  assign n48802 = \P2_P2_InstQueue_reg[8][5]/NET0131  & n26300 ;
  assign n48803 = \P2_P2_InstQueue_reg[12][5]/NET0131  & n26320 ;
  assign n48818 = ~n48802 & ~n48803 ;
  assign n48828 = ~n48811 & n48818 ;
  assign n48829 = ~n48813 & n48828 ;
  assign n48814 = \P2_P2_InstQueue_reg[15][5]/NET0131  & n26336 ;
  assign n48815 = \P2_P2_InstQueue_reg[7][5]/NET0131  & n26318 ;
  assign n48823 = ~n48814 & ~n48815 ;
  assign n48816 = \P2_P2_InstQueue_reg[4][5]/NET0131  & n26316 ;
  assign n48817 = \P2_P2_InstQueue_reg[3][5]/NET0131  & n26338 ;
  assign n48824 = ~n48816 & ~n48817 ;
  assign n48825 = n48823 & n48824 ;
  assign n48808 = \P2_P2_InstQueue_reg[11][5]/NET0131  & n26304 ;
  assign n48809 = \P2_P2_InstQueue_reg[5][5]/NET0131  & n26332 ;
  assign n48821 = ~n48808 & ~n48809 ;
  assign n48810 = \P2_P2_InstQueue_reg[6][5]/NET0131  & n26307 ;
  assign n48812 = \P2_P2_InstQueue_reg[9][5]/NET0131  & n26327 ;
  assign n48822 = ~n48810 & ~n48812 ;
  assign n48826 = n48821 & n48822 ;
  assign n48804 = \P2_P2_InstQueue_reg[2][5]/NET0131  & n26322 ;
  assign n48805 = \P2_P2_InstQueue_reg[13][5]/NET0131  & n26310 ;
  assign n48819 = ~n48804 & ~n48805 ;
  assign n48806 = \P2_P2_InstQueue_reg[10][5]/NET0131  & n26334 ;
  assign n48807 = \P2_P2_InstQueue_reg[14][5]/NET0131  & n26313 ;
  assign n48820 = ~n48806 & ~n48807 ;
  assign n48827 = n48819 & n48820 ;
  assign n48830 = n48826 & n48827 ;
  assign n48831 = n48825 & n48830 ;
  assign n48832 = n48829 & n48831 ;
  assign n48833 = n44510 & ~n48832 ;
  assign n48837 = ~n48800 & ~n48833 ;
  assign n48838 = ~n48836 & n48837 ;
  assign n48839 = ~n48801 & n48838 ;
  assign n48840 = n26792 & ~n48839 ;
  assign n48841 = ~n48798 & ~n48840 ;
  assign n48842 = \P2_P2_EAX_reg[14]/NET0131  & ~n44508 ;
  assign n48843 = ~n44718 & n44732 ;
  assign n48845 = ~n44736 & ~n48843 ;
  assign n48846 = \P2_P2_EAX_reg[14]/NET0131  & ~n48845 ;
  assign n48844 = n44717 & n48843 ;
  assign n48858 = \P2_P2_InstQueue_reg[0][6]/NET0131  & n26330 ;
  assign n48856 = \P2_P2_InstQueue_reg[1][6]/NET0131  & n26325 ;
  assign n48847 = \P2_P2_InstQueue_reg[8][6]/NET0131  & n26300 ;
  assign n48848 = \P2_P2_InstQueue_reg[4][6]/NET0131  & n26316 ;
  assign n48863 = ~n48847 & ~n48848 ;
  assign n48873 = ~n48856 & n48863 ;
  assign n48874 = ~n48858 & n48873 ;
  assign n48859 = \P2_P2_InstQueue_reg[6][6]/NET0131  & n26307 ;
  assign n48860 = \P2_P2_InstQueue_reg[15][6]/NET0131  & n26336 ;
  assign n48868 = ~n48859 & ~n48860 ;
  assign n48861 = \P2_P2_InstQueue_reg[10][6]/NET0131  & n26334 ;
  assign n48862 = \P2_P2_InstQueue_reg[14][6]/NET0131  & n26313 ;
  assign n48869 = ~n48861 & ~n48862 ;
  assign n48870 = n48868 & n48869 ;
  assign n48853 = \P2_P2_InstQueue_reg[12][6]/NET0131  & n26320 ;
  assign n48854 = \P2_P2_InstQueue_reg[11][6]/NET0131  & n26304 ;
  assign n48866 = ~n48853 & ~n48854 ;
  assign n48855 = \P2_P2_InstQueue_reg[2][6]/NET0131  & n26322 ;
  assign n48857 = \P2_P2_InstQueue_reg[9][6]/NET0131  & n26327 ;
  assign n48867 = ~n48855 & ~n48857 ;
  assign n48871 = n48866 & n48867 ;
  assign n48849 = \P2_P2_InstQueue_reg[5][6]/NET0131  & n26332 ;
  assign n48850 = \P2_P2_InstQueue_reg[7][6]/NET0131  & n26318 ;
  assign n48864 = ~n48849 & ~n48850 ;
  assign n48851 = \P2_P2_InstQueue_reg[3][6]/NET0131  & n26338 ;
  assign n48852 = \P2_P2_InstQueue_reg[13][6]/NET0131  & n26310 ;
  assign n48865 = ~n48851 & ~n48852 ;
  assign n48872 = n48864 & n48865 ;
  assign n48875 = n48871 & n48872 ;
  assign n48876 = n48870 & n48875 ;
  assign n48877 = n48874 & n48876 ;
  assign n48878 = n44510 & ~n48877 ;
  assign n48879 = \P2_P2_EAX_reg[14]/NET0131  & ~n26641 ;
  assign n48880 = ~n46284 & ~n48879 ;
  assign n48881 = ~n26639 & ~n48880 ;
  assign n48882 = ~n48878 & ~n48881 ;
  assign n48883 = ~n48844 & n48882 ;
  assign n48884 = ~n48846 & n48883 ;
  assign n48885 = n26792 & ~n48884 ;
  assign n48886 = ~n48842 & ~n48885 ;
  assign n48887 = \P2_P2_EAX_reg[7]/NET0131  & ~n48669 ;
  assign n48889 = n26641 & ~n28951 ;
  assign n48890 = ~n26639 & n48889 ;
  assign n48888 = ~n32510 & n44510 ;
  assign n48891 = ~\P2_P2_EAX_reg[7]/NET0131  & ~n44710 ;
  assign n48892 = ~n44711 & ~n48891 ;
  assign n48893 = n44732 & n48892 ;
  assign n48894 = ~n48888 & ~n48893 ;
  assign n48895 = ~n48890 & n48894 ;
  assign n48896 = n26792 & ~n48895 ;
  assign n48897 = ~n48887 & ~n48896 ;
  assign n48898 = \P2_P2_EAX_reg[8]/NET0131  & ~n48669 ;
  assign n48899 = \P2_buf2_reg[8]/NET0131  & ~n28013 ;
  assign n48900 = \P2_buf1_reg[8]/NET0131  & n28013 ;
  assign n48901 = ~n48899 & ~n48900 ;
  assign n48902 = n26641 & ~n48901 ;
  assign n48903 = ~n26639 & n48902 ;
  assign n48915 = \P2_P2_InstQueue_reg[0][0]/NET0131  & n26330 ;
  assign n48913 = \P2_P2_InstQueue_reg[1][0]/NET0131  & n26325 ;
  assign n48904 = \P2_P2_InstQueue_reg[8][0]/NET0131  & n26300 ;
  assign n48905 = \P2_P2_InstQueue_reg[15][0]/NET0131  & n26336 ;
  assign n48920 = ~n48904 & ~n48905 ;
  assign n48930 = ~n48913 & n48920 ;
  assign n48931 = ~n48915 & n48930 ;
  assign n48916 = \P2_P2_InstQueue_reg[14][0]/NET0131  & n26313 ;
  assign n48917 = \P2_P2_InstQueue_reg[11][0]/NET0131  & n26304 ;
  assign n48925 = ~n48916 & ~n48917 ;
  assign n48918 = \P2_P2_InstQueue_reg[7][0]/NET0131  & n26318 ;
  assign n48919 = \P2_P2_InstQueue_reg[13][0]/NET0131  & n26310 ;
  assign n48926 = ~n48918 & ~n48919 ;
  assign n48927 = n48925 & n48926 ;
  assign n48910 = \P2_P2_InstQueue_reg[10][0]/NET0131  & n26334 ;
  assign n48911 = \P2_P2_InstQueue_reg[2][0]/NET0131  & n26322 ;
  assign n48923 = ~n48910 & ~n48911 ;
  assign n48912 = \P2_P2_InstQueue_reg[6][0]/NET0131  & n26307 ;
  assign n48914 = \P2_P2_InstQueue_reg[9][0]/NET0131  & n26327 ;
  assign n48924 = ~n48912 & ~n48914 ;
  assign n48928 = n48923 & n48924 ;
  assign n48906 = \P2_P2_InstQueue_reg[12][0]/NET0131  & n26320 ;
  assign n48907 = \P2_P2_InstQueue_reg[5][0]/NET0131  & n26332 ;
  assign n48921 = ~n48906 & ~n48907 ;
  assign n48908 = \P2_P2_InstQueue_reg[3][0]/NET0131  & n26338 ;
  assign n48909 = \P2_P2_InstQueue_reg[4][0]/NET0131  & n26316 ;
  assign n48922 = ~n48908 & ~n48909 ;
  assign n48929 = n48921 & n48922 ;
  assign n48932 = n48928 & n48929 ;
  assign n48933 = n48927 & n48932 ;
  assign n48934 = n48931 & n48933 ;
  assign n48935 = n44510 & ~n48934 ;
  assign n48936 = ~\P2_P2_EAX_reg[8]/NET0131  & ~n44711 ;
  assign n48937 = ~n44712 & ~n48936 ;
  assign n48938 = n44732 & n48937 ;
  assign n48939 = ~n48935 & ~n48938 ;
  assign n48940 = ~n48903 & n48939 ;
  assign n48941 = n26792 & ~n48940 ;
  assign n48942 = ~n48898 & ~n48941 ;
  assign n48943 = \P2_P2_EAX_reg[9]/NET0131  & ~n48669 ;
  assign n48944 = \P2_buf2_reg[9]/NET0131  & ~n28013 ;
  assign n48945 = \P2_buf1_reg[9]/NET0131  & n28013 ;
  assign n48946 = ~n48944 & ~n48945 ;
  assign n48947 = n26641 & ~n48946 ;
  assign n48948 = ~n26639 & n48947 ;
  assign n48960 = \P2_P2_InstQueue_reg[0][1]/NET0131  & n26330 ;
  assign n48958 = \P2_P2_InstQueue_reg[1][1]/NET0131  & n26325 ;
  assign n48949 = \P2_P2_InstQueue_reg[8][1]/NET0131  & n26300 ;
  assign n48950 = \P2_P2_InstQueue_reg[3][1]/NET0131  & n26338 ;
  assign n48965 = ~n48949 & ~n48950 ;
  assign n48975 = ~n48958 & n48965 ;
  assign n48976 = ~n48960 & n48975 ;
  assign n48961 = \P2_P2_InstQueue_reg[4][1]/NET0131  & n26316 ;
  assign n48962 = \P2_P2_InstQueue_reg[15][1]/NET0131  & n26336 ;
  assign n48970 = ~n48961 & ~n48962 ;
  assign n48963 = \P2_P2_InstQueue_reg[14][1]/NET0131  & n26313 ;
  assign n48964 = \P2_P2_InstQueue_reg[13][1]/NET0131  & n26310 ;
  assign n48971 = ~n48963 & ~n48964 ;
  assign n48972 = n48970 & n48971 ;
  assign n48955 = \P2_P2_InstQueue_reg[11][1]/NET0131  & n26304 ;
  assign n48956 = \P2_P2_InstQueue_reg[7][1]/NET0131  & n26318 ;
  assign n48968 = ~n48955 & ~n48956 ;
  assign n48957 = \P2_P2_InstQueue_reg[6][1]/NET0131  & n26307 ;
  assign n48959 = \P2_P2_InstQueue_reg[9][1]/NET0131  & n26327 ;
  assign n48969 = ~n48957 & ~n48959 ;
  assign n48973 = n48968 & n48969 ;
  assign n48951 = \P2_P2_InstQueue_reg[10][1]/NET0131  & n26334 ;
  assign n48952 = \P2_P2_InstQueue_reg[5][1]/NET0131  & n26332 ;
  assign n48966 = ~n48951 & ~n48952 ;
  assign n48953 = \P2_P2_InstQueue_reg[12][1]/NET0131  & n26320 ;
  assign n48954 = \P2_P2_InstQueue_reg[2][1]/NET0131  & n26322 ;
  assign n48967 = ~n48953 & ~n48954 ;
  assign n48974 = n48966 & n48967 ;
  assign n48977 = n48973 & n48974 ;
  assign n48978 = n48972 & n48977 ;
  assign n48979 = n48976 & n48978 ;
  assign n48980 = n44510 & ~n48979 ;
  assign n48981 = ~\P2_P2_EAX_reg[9]/NET0131  & ~n44712 ;
  assign n48982 = ~n44713 & ~n48981 ;
  assign n48983 = n44732 & n48982 ;
  assign n48984 = ~n48980 & ~n48983 ;
  assign n48985 = ~n48948 & n48984 ;
  assign n48986 = n26792 & ~n48985 ;
  assign n48987 = ~n48943 & ~n48986 ;
  assign n48990 = ~\P2_P2_EBX_reg[29]/NET0131  & ~n46458 ;
  assign n48991 = n26662 & ~n46459 ;
  assign n48992 = ~n48990 & n48991 ;
  assign n48988 = \P2_P2_EBX_reg[29]/NET0131  & n46417 ;
  assign n48989 = n46416 & n48204 ;
  assign n48993 = ~n48988 & ~n48989 ;
  assign n48994 = ~n48992 & n48993 ;
  assign n48995 = n26792 & ~n48994 ;
  assign n48996 = \P2_P2_EBX_reg[29]/NET0131  & ~n44508 ;
  assign n48997 = ~n48995 & ~n48996 ;
  assign n49000 = ~\P1_P3_EBX_reg[29]/NET0131  & ~n46520 ;
  assign n49001 = n9108 & ~n46521 ;
  assign n49002 = ~n49000 & n49001 ;
  assign n48998 = \P1_P3_EBX_reg[29]/NET0131  & n46480 ;
  assign n48999 = n21665 & n46479 ;
  assign n49003 = ~n48998 & ~n48999 ;
  assign n49004 = ~n49002 & n49003 ;
  assign n49005 = n9241 & ~n49004 ;
  assign n49006 = \P1_P3_EBX_reg[29]/NET0131  & ~n16968 ;
  assign n49007 = ~n49005 & ~n49006 ;
  assign n49008 = \P1_P1_uWord_reg[4]/NET0131  & ~n24515 ;
  assign n49010 = \P1_P1_uWord_reg[4]/NET0131  & n15335 ;
  assign n49011 = ~n24696 & ~n49010 ;
  assign n49012 = n15334 & ~n49011 ;
  assign n49009 = \P1_P1_uWord_reg[4]/NET0131  & n24505 ;
  assign n49013 = ~\P1_P1_EAX_reg[20]/NET0131  & ~n25351 ;
  assign n49014 = ~n25352 & ~n49013 ;
  assign n49015 = n24503 & n49014 ;
  assign n49016 = ~n49009 & ~n49015 ;
  assign n49017 = ~n49012 & n49016 ;
  assign n49018 = n8355 & ~n49017 ;
  assign n49019 = ~n49008 & ~n49018 ;
  assign n49022 = ~\P1_P1_EBX_reg[29]/NET0131  & ~n46575 ;
  assign n49023 = n26146 & ~n46576 ;
  assign n49024 = ~n49022 & n49023 ;
  assign n49020 = n23181 & n46535 ;
  assign n49021 = \P1_P1_EBX_reg[29]/NET0131  & ~n46533 ;
  assign n49025 = ~n49020 & ~n49021 ;
  assign n49026 = ~n49024 & n49025 ;
  assign n49027 = n8355 & ~n49026 ;
  assign n49028 = \P1_P1_EBX_reg[29]/NET0131  & ~n15326 ;
  assign n49029 = ~n49027 & ~n49028 ;
  assign n49030 = \P2_P2_uWord_reg[8]/NET0131  & ~n47642 ;
  assign n49031 = n47676 & ~n48901 ;
  assign n49032 = ~n48501 & ~n49031 ;
  assign n49033 = ~n26640 & ~n49032 ;
  assign n49034 = \P2_P2_uWord_reg[8]/NET0131  & ~n47686 ;
  assign n49035 = ~n49033 & ~n49034 ;
  assign n49036 = n26792 & ~n49035 ;
  assign n49037 = ~n49030 & ~n49036 ;
  assign n49038 = n27308 & ~n42543 ;
  assign n49039 = n42872 & ~n49038 ;
  assign n49040 = \P2_P3_EAX_reg[10]/NET0131  & ~n49039 ;
  assign n49076 = \P2_buf2_reg[10]/NET0131  & n27228 ;
  assign n49041 = ~\P2_P3_EAX_reg[10]/NET0131  & ~n42841 ;
  assign n49042 = n42539 & ~n42842 ;
  assign n49043 = ~n49041 & n49042 ;
  assign n49052 = \P2_P3_InstQueue_reg[0][2]/NET0131  & n26845 ;
  assign n49044 = \P2_P3_InstQueue_reg[6][2]/NET0131  & n26815 ;
  assign n49045 = \P2_P3_InstQueue_reg[7][2]/NET0131  & n26822 ;
  assign n49060 = ~n49044 & ~n49045 ;
  assign n49069 = ~n49052 & n49060 ;
  assign n49054 = \P2_P3_InstQueue_reg[1][2]/NET0131  & n26837 ;
  assign n49055 = \P2_P3_InstQueue_reg[9][2]/NET0131  & n26839 ;
  assign n49070 = ~n49054 & ~n49055 ;
  assign n49071 = n49069 & n49070 ;
  assign n49059 = \P2_P3_InstQueue_reg[3][2]/NET0131  & n26831 ;
  assign n49057 = \P2_P3_InstQueue_reg[5][2]/NET0131  & n26847 ;
  assign n49058 = \P2_P3_InstQueue_reg[2][2]/NET0131  & n26812 ;
  assign n49065 = ~n49057 & ~n49058 ;
  assign n49066 = ~n49059 & n49065 ;
  assign n49050 = \P2_P3_InstQueue_reg[12][2]/NET0131  & n26819 ;
  assign n49051 = \P2_P3_InstQueue_reg[15][2]/NET0131  & n26825 ;
  assign n49063 = ~n49050 & ~n49051 ;
  assign n49053 = \P2_P3_InstQueue_reg[8][2]/NET0131  & n26841 ;
  assign n49056 = \P2_P3_InstQueue_reg[13][2]/NET0131  & n26849 ;
  assign n49064 = ~n49053 & ~n49056 ;
  assign n49067 = n49063 & n49064 ;
  assign n49046 = \P2_P3_InstQueue_reg[4][2]/NET0131  & n26843 ;
  assign n49047 = \P2_P3_InstQueue_reg[14][2]/NET0131  & n26829 ;
  assign n49061 = ~n49046 & ~n49047 ;
  assign n49048 = \P2_P3_InstQueue_reg[11][2]/NET0131  & n26833 ;
  assign n49049 = \P2_P3_InstQueue_reg[10][2]/NET0131  & n26827 ;
  assign n49062 = ~n49048 & ~n49049 ;
  assign n49068 = n49061 & n49062 ;
  assign n49072 = n49067 & n49068 ;
  assign n49073 = n49066 & n49072 ;
  assign n49074 = n49071 & n49073 ;
  assign n49075 = n42538 & ~n49074 ;
  assign n49077 = ~n49043 & ~n49075 ;
  assign n49078 = ~n49076 & n49077 ;
  assign n49079 = n27308 & ~n49078 ;
  assign n49080 = ~n49040 & ~n49079 ;
  assign n49081 = \P2_P3_EAX_reg[11]/NET0131  & ~n42872 ;
  assign n49084 = ~n42542 & ~n49042 ;
  assign n49085 = \P2_P3_EAX_reg[11]/NET0131  & ~n49084 ;
  assign n49118 = \P2_P3_EAX_reg[11]/NET0131  & ~n27227 ;
  assign n49119 = ~n44800 & ~n49118 ;
  assign n49120 = ~n27226 & ~n49119 ;
  assign n49082 = n42539 & ~n42843 ;
  assign n49083 = n42842 & n49082 ;
  assign n49094 = \P2_P3_InstQueue_reg[0][3]/NET0131  & n26845 ;
  assign n49086 = \P2_P3_InstQueue_reg[6][3]/NET0131  & n26815 ;
  assign n49087 = \P2_P3_InstQueue_reg[5][3]/NET0131  & n26847 ;
  assign n49102 = ~n49086 & ~n49087 ;
  assign n49111 = ~n49094 & n49102 ;
  assign n49096 = \P2_P3_InstQueue_reg[1][3]/NET0131  & n26837 ;
  assign n49097 = \P2_P3_InstQueue_reg[9][3]/NET0131  & n26839 ;
  assign n49112 = ~n49096 & ~n49097 ;
  assign n49113 = n49111 & n49112 ;
  assign n49101 = \P2_P3_InstQueue_reg[14][3]/NET0131  & n26829 ;
  assign n49099 = \P2_P3_InstQueue_reg[15][3]/NET0131  & n26825 ;
  assign n49100 = \P2_P3_InstQueue_reg[2][3]/NET0131  & n26812 ;
  assign n49107 = ~n49099 & ~n49100 ;
  assign n49108 = ~n49101 & n49107 ;
  assign n49092 = \P2_P3_InstQueue_reg[3][3]/NET0131  & n26831 ;
  assign n49093 = \P2_P3_InstQueue_reg[7][3]/NET0131  & n26822 ;
  assign n49105 = ~n49092 & ~n49093 ;
  assign n49095 = \P2_P3_InstQueue_reg[8][3]/NET0131  & n26841 ;
  assign n49098 = \P2_P3_InstQueue_reg[11][3]/NET0131  & n26833 ;
  assign n49106 = ~n49095 & ~n49098 ;
  assign n49109 = n49105 & n49106 ;
  assign n49088 = \P2_P3_InstQueue_reg[4][3]/NET0131  & n26843 ;
  assign n49089 = \P2_P3_InstQueue_reg[10][3]/NET0131  & n26827 ;
  assign n49103 = ~n49088 & ~n49089 ;
  assign n49090 = \P2_P3_InstQueue_reg[12][3]/NET0131  & n26819 ;
  assign n49091 = \P2_P3_InstQueue_reg[13][3]/NET0131  & n26849 ;
  assign n49104 = ~n49090 & ~n49091 ;
  assign n49110 = n49103 & n49104 ;
  assign n49114 = n49109 & n49110 ;
  assign n49115 = n49108 & n49114 ;
  assign n49116 = n49113 & n49115 ;
  assign n49117 = n42538 & ~n49116 ;
  assign n49121 = ~n49083 & ~n49117 ;
  assign n49122 = ~n49120 & n49121 ;
  assign n49123 = ~n49085 & n49122 ;
  assign n49124 = n27308 & ~n49123 ;
  assign n49125 = ~n49081 & ~n49124 ;
  assign n49126 = \P2_P3_EAX_reg[12]/NET0131  & ~n42872 ;
  assign n49128 = n42543 & ~n49082 ;
  assign n49129 = \P2_P3_EAX_reg[12]/NET0131  & ~n49128 ;
  assign n49127 = \P2_buf2_reg[12]/NET0131  & n27228 ;
  assign n49130 = n42539 & ~n42844 ;
  assign n49131 = n42843 & n49130 ;
  assign n49140 = \P2_P3_InstQueue_reg[0][4]/NET0131  & n26845 ;
  assign n49132 = \P2_P3_InstQueue_reg[6][4]/NET0131  & n26815 ;
  assign n49133 = \P2_P3_InstQueue_reg[7][4]/NET0131  & n26822 ;
  assign n49148 = ~n49132 & ~n49133 ;
  assign n49157 = ~n49140 & n49148 ;
  assign n49142 = \P2_P3_InstQueue_reg[1][4]/NET0131  & n26837 ;
  assign n49143 = \P2_P3_InstQueue_reg[9][4]/NET0131  & n26839 ;
  assign n49158 = ~n49142 & ~n49143 ;
  assign n49159 = n49157 & n49158 ;
  assign n49147 = \P2_P3_InstQueue_reg[3][4]/NET0131  & n26831 ;
  assign n49145 = \P2_P3_InstQueue_reg[5][4]/NET0131  & n26847 ;
  assign n49146 = \P2_P3_InstQueue_reg[2][4]/NET0131  & n26812 ;
  assign n49153 = ~n49145 & ~n49146 ;
  assign n49154 = ~n49147 & n49153 ;
  assign n49138 = \P2_P3_InstQueue_reg[12][4]/NET0131  & n26819 ;
  assign n49139 = \P2_P3_InstQueue_reg[15][4]/NET0131  & n26825 ;
  assign n49151 = ~n49138 & ~n49139 ;
  assign n49141 = \P2_P3_InstQueue_reg[8][4]/NET0131  & n26841 ;
  assign n49144 = \P2_P3_InstQueue_reg[13][4]/NET0131  & n26849 ;
  assign n49152 = ~n49141 & ~n49144 ;
  assign n49155 = n49151 & n49152 ;
  assign n49134 = \P2_P3_InstQueue_reg[4][4]/NET0131  & n26843 ;
  assign n49135 = \P2_P3_InstQueue_reg[14][4]/NET0131  & n26829 ;
  assign n49149 = ~n49134 & ~n49135 ;
  assign n49136 = \P2_P3_InstQueue_reg[11][4]/NET0131  & n26833 ;
  assign n49137 = \P2_P3_InstQueue_reg[10][4]/NET0131  & n26827 ;
  assign n49150 = ~n49136 & ~n49137 ;
  assign n49156 = n49149 & n49150 ;
  assign n49160 = n49155 & n49156 ;
  assign n49161 = n49154 & n49160 ;
  assign n49162 = n49159 & n49161 ;
  assign n49163 = n42538 & ~n49162 ;
  assign n49164 = ~n49131 & ~n49163 ;
  assign n49165 = ~n49127 & n49164 ;
  assign n49166 = ~n49129 & n49165 ;
  assign n49167 = n27308 & ~n49166 ;
  assign n49168 = ~n49126 & ~n49167 ;
  assign n49169 = \P2_P3_EAX_reg[13]/NET0131  & ~n42872 ;
  assign n49170 = ~n42542 & ~n49130 ;
  assign n49171 = \P2_P3_EAX_reg[13]/NET0131  & ~n49170 ;
  assign n49206 = \P2_buf2_reg[13]/NET0131  & n27227 ;
  assign n49207 = \P2_P3_EAX_reg[13]/NET0131  & ~n27227 ;
  assign n49208 = ~n49206 & ~n49207 ;
  assign n49209 = ~n27226 & ~n49208 ;
  assign n49172 = ~\P2_P3_EAX_reg[13]/NET0131  & n42539 ;
  assign n49173 = n42844 & n49172 ;
  assign n49182 = \P2_P3_InstQueue_reg[0][5]/NET0131  & n26845 ;
  assign n49174 = \P2_P3_InstQueue_reg[6][5]/NET0131  & n26815 ;
  assign n49175 = \P2_P3_InstQueue_reg[7][5]/NET0131  & n26822 ;
  assign n49190 = ~n49174 & ~n49175 ;
  assign n49199 = ~n49182 & n49190 ;
  assign n49184 = \P2_P3_InstQueue_reg[1][5]/NET0131  & n26837 ;
  assign n49185 = \P2_P3_InstQueue_reg[9][5]/NET0131  & n26839 ;
  assign n49200 = ~n49184 & ~n49185 ;
  assign n49201 = n49199 & n49200 ;
  assign n49189 = \P2_P3_InstQueue_reg[3][5]/NET0131  & n26831 ;
  assign n49187 = \P2_P3_InstQueue_reg[5][5]/NET0131  & n26847 ;
  assign n49188 = \P2_P3_InstQueue_reg[2][5]/NET0131  & n26812 ;
  assign n49195 = ~n49187 & ~n49188 ;
  assign n49196 = ~n49189 & n49195 ;
  assign n49180 = \P2_P3_InstQueue_reg[12][5]/NET0131  & n26819 ;
  assign n49181 = \P2_P3_InstQueue_reg[15][5]/NET0131  & n26825 ;
  assign n49193 = ~n49180 & ~n49181 ;
  assign n49183 = \P2_P3_InstQueue_reg[8][5]/NET0131  & n26841 ;
  assign n49186 = \P2_P3_InstQueue_reg[13][5]/NET0131  & n26849 ;
  assign n49194 = ~n49183 & ~n49186 ;
  assign n49197 = n49193 & n49194 ;
  assign n49176 = \P2_P3_InstQueue_reg[4][5]/NET0131  & n26843 ;
  assign n49177 = \P2_P3_InstQueue_reg[14][5]/NET0131  & n26829 ;
  assign n49191 = ~n49176 & ~n49177 ;
  assign n49178 = \P2_P3_InstQueue_reg[11][5]/NET0131  & n26833 ;
  assign n49179 = \P2_P3_InstQueue_reg[10][5]/NET0131  & n26827 ;
  assign n49192 = ~n49178 & ~n49179 ;
  assign n49198 = n49191 & n49192 ;
  assign n49202 = n49197 & n49198 ;
  assign n49203 = n49196 & n49202 ;
  assign n49204 = n49201 & n49203 ;
  assign n49205 = n42538 & ~n49204 ;
  assign n49210 = ~n49173 & ~n49205 ;
  assign n49211 = ~n49209 & n49210 ;
  assign n49212 = ~n49171 & n49211 ;
  assign n49213 = n27308 & ~n49212 ;
  assign n49214 = ~n49169 & ~n49213 ;
  assign n49215 = \P2_P3_EAX_reg[14]/NET0131  & ~n42872 ;
  assign n49216 = n42539 & ~n42846 ;
  assign n49218 = ~n42542 & ~n49216 ;
  assign n49219 = \P2_P3_EAX_reg[14]/NET0131  & ~n49218 ;
  assign n49217 = n42845 & n49216 ;
  assign n49228 = \P2_P3_InstQueue_reg[0][6]/NET0131  & n26845 ;
  assign n49220 = \P2_P3_InstQueue_reg[6][6]/NET0131  & n26815 ;
  assign n49221 = \P2_P3_InstQueue_reg[5][6]/NET0131  & n26847 ;
  assign n49236 = ~n49220 & ~n49221 ;
  assign n49245 = ~n49228 & n49236 ;
  assign n49230 = \P2_P3_InstQueue_reg[1][6]/NET0131  & n26837 ;
  assign n49231 = \P2_P3_InstQueue_reg[9][6]/NET0131  & n26839 ;
  assign n49246 = ~n49230 & ~n49231 ;
  assign n49247 = n49245 & n49246 ;
  assign n49235 = \P2_P3_InstQueue_reg[14][6]/NET0131  & n26829 ;
  assign n49233 = \P2_P3_InstQueue_reg[7][6]/NET0131  & n26822 ;
  assign n49234 = \P2_P3_InstQueue_reg[2][6]/NET0131  & n26812 ;
  assign n49241 = ~n49233 & ~n49234 ;
  assign n49242 = ~n49235 & n49241 ;
  assign n49226 = \P2_P3_InstQueue_reg[3][6]/NET0131  & n26831 ;
  assign n49227 = \P2_P3_InstQueue_reg[15][6]/NET0131  & n26825 ;
  assign n49239 = ~n49226 & ~n49227 ;
  assign n49229 = \P2_P3_InstQueue_reg[8][6]/NET0131  & n26841 ;
  assign n49232 = \P2_P3_InstQueue_reg[11][6]/NET0131  & n26833 ;
  assign n49240 = ~n49229 & ~n49232 ;
  assign n49243 = n49239 & n49240 ;
  assign n49222 = \P2_P3_InstQueue_reg[4][6]/NET0131  & n26843 ;
  assign n49223 = \P2_P3_InstQueue_reg[13][6]/NET0131  & n26849 ;
  assign n49237 = ~n49222 & ~n49223 ;
  assign n49224 = \P2_P3_InstQueue_reg[12][6]/NET0131  & n26819 ;
  assign n49225 = \P2_P3_InstQueue_reg[10][6]/NET0131  & n26827 ;
  assign n49238 = ~n49224 & ~n49225 ;
  assign n49244 = n49237 & n49238 ;
  assign n49248 = n49243 & n49244 ;
  assign n49249 = n49242 & n49248 ;
  assign n49250 = n49247 & n49249 ;
  assign n49251 = n42538 & ~n49250 ;
  assign n49252 = \P2_P3_EAX_reg[14]/NET0131  & ~n27227 ;
  assign n49253 = ~n27177 & n46588 ;
  assign n49254 = ~n49252 & ~n49253 ;
  assign n49255 = ~n27226 & ~n49254 ;
  assign n49256 = ~n49251 & ~n49255 ;
  assign n49257 = ~n49217 & n49256 ;
  assign n49258 = ~n49219 & n49257 ;
  assign n49259 = n27308 & ~n49258 ;
  assign n49260 = ~n49215 & ~n49259 ;
  assign n49261 = \P2_P3_EAX_reg[15]/NET0131  & ~n42872 ;
  assign n49264 = \P2_P3_EAX_reg[15]/NET0131  & ~n49218 ;
  assign n49262 = ~\P2_P3_EAX_reg[15]/NET0131  & n42539 ;
  assign n49263 = n42846 & n49262 ;
  assign n49273 = \P2_P3_InstQueue_reg[0][7]/NET0131  & n26845 ;
  assign n49265 = \P2_P3_InstQueue_reg[6][7]/NET0131  & n26815 ;
  assign n49266 = \P2_P3_InstQueue_reg[7][7]/NET0131  & n26822 ;
  assign n49281 = ~n49265 & ~n49266 ;
  assign n49290 = ~n49273 & n49281 ;
  assign n49275 = \P2_P3_InstQueue_reg[1][7]/NET0131  & n26837 ;
  assign n49276 = \P2_P3_InstQueue_reg[9][7]/NET0131  & n26839 ;
  assign n49291 = ~n49275 & ~n49276 ;
  assign n49292 = n49290 & n49291 ;
  assign n49280 = \P2_P3_InstQueue_reg[3][7]/NET0131  & n26831 ;
  assign n49278 = \P2_P3_InstQueue_reg[5][7]/NET0131  & n26847 ;
  assign n49279 = \P2_P3_InstQueue_reg[2][7]/NET0131  & n26812 ;
  assign n49286 = ~n49278 & ~n49279 ;
  assign n49287 = ~n49280 & n49286 ;
  assign n49271 = \P2_P3_InstQueue_reg[12][7]/NET0131  & n26819 ;
  assign n49272 = \P2_P3_InstQueue_reg[15][7]/NET0131  & n26825 ;
  assign n49284 = ~n49271 & ~n49272 ;
  assign n49274 = \P2_P3_InstQueue_reg[8][7]/NET0131  & n26841 ;
  assign n49277 = \P2_P3_InstQueue_reg[13][7]/NET0131  & n26849 ;
  assign n49285 = ~n49274 & ~n49277 ;
  assign n49288 = n49284 & n49285 ;
  assign n49267 = \P2_P3_InstQueue_reg[4][7]/NET0131  & n26843 ;
  assign n49268 = \P2_P3_InstQueue_reg[14][7]/NET0131  & n26829 ;
  assign n49282 = ~n49267 & ~n49268 ;
  assign n49269 = \P2_P3_InstQueue_reg[11][7]/NET0131  & n26833 ;
  assign n49270 = \P2_P3_InstQueue_reg[10][7]/NET0131  & n26827 ;
  assign n49283 = ~n49269 & ~n49270 ;
  assign n49289 = n49282 & n49283 ;
  assign n49293 = n49288 & n49289 ;
  assign n49294 = n49287 & n49293 ;
  assign n49295 = n49292 & n49294 ;
  assign n49296 = n42538 & ~n49295 ;
  assign n49297 = \P2_P3_EAX_reg[15]/NET0131  & ~n27227 ;
  assign n49298 = \P2_buf2_reg[15]/NET0131  & n27227 ;
  assign n49299 = ~n49297 & ~n49298 ;
  assign n49300 = ~n27226 & ~n49299 ;
  assign n49301 = ~n49296 & ~n49300 ;
  assign n49302 = ~n49263 & n49301 ;
  assign n49303 = ~n49264 & n49302 ;
  assign n49304 = n27308 & ~n49303 ;
  assign n49305 = ~n49261 & ~n49304 ;
  assign n49306 = \P2_P3_EAX_reg[7]/NET0131  & ~n49039 ;
  assign n49308 = \P2_buf2_reg[7]/NET0131  & n27228 ;
  assign n49307 = ~n33242 & n42538 ;
  assign n49309 = ~\P2_P3_EAX_reg[7]/NET0131  & ~n42838 ;
  assign n49310 = ~n42839 & ~n49309 ;
  assign n49311 = n42539 & n49310 ;
  assign n49312 = ~n49307 & ~n49311 ;
  assign n49313 = ~n49308 & n49312 ;
  assign n49314 = n27308 & ~n49313 ;
  assign n49315 = ~n49306 & ~n49314 ;
  assign n49316 = \P2_P3_EAX_reg[8]/NET0131  & ~n49039 ;
  assign n49349 = \P2_buf2_reg[8]/NET0131  & n27228 ;
  assign n49325 = \P2_P3_InstQueue_reg[0][0]/NET0131  & n26845 ;
  assign n49317 = \P2_P3_InstQueue_reg[5][0]/NET0131  & n26847 ;
  assign n49318 = \P2_P3_InstQueue_reg[15][0]/NET0131  & n26825 ;
  assign n49333 = ~n49317 & ~n49318 ;
  assign n49342 = ~n49325 & n49333 ;
  assign n49327 = \P2_P3_InstQueue_reg[1][0]/NET0131  & n26837 ;
  assign n49328 = \P2_P3_InstQueue_reg[9][0]/NET0131  & n26839 ;
  assign n49343 = ~n49327 & ~n49328 ;
  assign n49344 = n49342 & n49343 ;
  assign n49332 = \P2_P3_InstQueue_reg[3][0]/NET0131  & n26831 ;
  assign n49330 = \P2_P3_InstQueue_reg[11][0]/NET0131  & n26833 ;
  assign n49331 = \P2_P3_InstQueue_reg[2][0]/NET0131  & n26812 ;
  assign n49338 = ~n49330 & ~n49331 ;
  assign n49339 = ~n49332 & n49338 ;
  assign n49323 = \P2_P3_InstQueue_reg[12][0]/NET0131  & n26819 ;
  assign n49324 = \P2_P3_InstQueue_reg[7][0]/NET0131  & n26822 ;
  assign n49336 = ~n49323 & ~n49324 ;
  assign n49326 = \P2_P3_InstQueue_reg[8][0]/NET0131  & n26841 ;
  assign n49329 = \P2_P3_InstQueue_reg[10][0]/NET0131  & n26827 ;
  assign n49337 = ~n49326 & ~n49329 ;
  assign n49340 = n49336 & n49337 ;
  assign n49319 = \P2_P3_InstQueue_reg[4][0]/NET0131  & n26843 ;
  assign n49320 = \P2_P3_InstQueue_reg[6][0]/NET0131  & n26815 ;
  assign n49334 = ~n49319 & ~n49320 ;
  assign n49321 = \P2_P3_InstQueue_reg[14][0]/NET0131  & n26829 ;
  assign n49322 = \P2_P3_InstQueue_reg[13][0]/NET0131  & n26849 ;
  assign n49335 = ~n49321 & ~n49322 ;
  assign n49341 = n49334 & n49335 ;
  assign n49345 = n49340 & n49341 ;
  assign n49346 = n49339 & n49345 ;
  assign n49347 = n49344 & n49346 ;
  assign n49348 = n42538 & ~n49347 ;
  assign n49350 = ~\P2_P3_EAX_reg[8]/NET0131  & ~n42839 ;
  assign n49351 = ~n42840 & ~n49350 ;
  assign n49352 = n42539 & n49351 ;
  assign n49353 = ~n49348 & ~n49352 ;
  assign n49354 = ~n49349 & n49353 ;
  assign n49355 = n27308 & ~n49354 ;
  assign n49356 = ~n49316 & ~n49355 ;
  assign n49357 = \P2_P3_EAX_reg[9]/NET0131  & ~n49039 ;
  assign n49358 = \P2_buf2_reg[9]/NET0131  & n27228 ;
  assign n49367 = \P2_P3_InstQueue_reg[0][1]/NET0131  & n26845 ;
  assign n49359 = \P2_P3_InstQueue_reg[6][1]/NET0131  & n26815 ;
  assign n49360 = \P2_P3_InstQueue_reg[7][1]/NET0131  & n26822 ;
  assign n49375 = ~n49359 & ~n49360 ;
  assign n49384 = ~n49367 & n49375 ;
  assign n49369 = \P2_P3_InstQueue_reg[1][1]/NET0131  & n26837 ;
  assign n49370 = \P2_P3_InstQueue_reg[9][1]/NET0131  & n26839 ;
  assign n49385 = ~n49369 & ~n49370 ;
  assign n49386 = n49384 & n49385 ;
  assign n49374 = \P2_P3_InstQueue_reg[3][1]/NET0131  & n26831 ;
  assign n49372 = \P2_P3_InstQueue_reg[11][1]/NET0131  & n26833 ;
  assign n49373 = \P2_P3_InstQueue_reg[2][1]/NET0131  & n26812 ;
  assign n49380 = ~n49372 & ~n49373 ;
  assign n49381 = ~n49374 & n49380 ;
  assign n49365 = \P2_P3_InstQueue_reg[12][1]/NET0131  & n26819 ;
  assign n49366 = \P2_P3_InstQueue_reg[15][1]/NET0131  & n26825 ;
  assign n49378 = ~n49365 & ~n49366 ;
  assign n49368 = \P2_P3_InstQueue_reg[8][1]/NET0131  & n26841 ;
  assign n49371 = \P2_P3_InstQueue_reg[13][1]/NET0131  & n26849 ;
  assign n49379 = ~n49368 & ~n49371 ;
  assign n49382 = n49378 & n49379 ;
  assign n49361 = \P2_P3_InstQueue_reg[4][1]/NET0131  & n26843 ;
  assign n49362 = \P2_P3_InstQueue_reg[14][1]/NET0131  & n26829 ;
  assign n49376 = ~n49361 & ~n49362 ;
  assign n49363 = \P2_P3_InstQueue_reg[5][1]/NET0131  & n26847 ;
  assign n49364 = \P2_P3_InstQueue_reg[10][1]/NET0131  & n26827 ;
  assign n49377 = ~n49363 & ~n49364 ;
  assign n49383 = n49376 & n49377 ;
  assign n49387 = n49382 & n49383 ;
  assign n49388 = n49381 & n49387 ;
  assign n49389 = n49386 & n49388 ;
  assign n49390 = n42538 & ~n49389 ;
  assign n49391 = ~\P2_P3_EAX_reg[9]/NET0131  & ~n42840 ;
  assign n49392 = ~n42841 & ~n49391 ;
  assign n49393 = n42539 & n49392 ;
  assign n49394 = ~n49390 & ~n49393 ;
  assign n49395 = ~n49358 & n49394 ;
  assign n49396 = n27308 & ~n49395 ;
  assign n49397 = ~n49357 & ~n49396 ;
  assign n49400 = ~\P2_P3_EBX_reg[29]/NET0131  & ~n46655 ;
  assign n49401 = n27133 & ~n46656 ;
  assign n49402 = ~n49400 & n49401 ;
  assign n49398 = \P2_P3_EBX_reg[29]/NET0131  & n46615 ;
  assign n49399 = n46614 & n48262 ;
  assign n49403 = ~n49398 & ~n49399 ;
  assign n49404 = ~n49402 & n49403 ;
  assign n49405 = n27308 & ~n49404 ;
  assign n49406 = \P2_P3_EBX_reg[29]/NET0131  & ~n42872 ;
  assign n49407 = ~n49405 & ~n49406 ;
  assign n49408 = \P1_P2_EAX_reg[10]/NET0131  & ~n43212 ;
  assign n49410 = n43164 & ~n43180 ;
  assign n49411 = n43169 & ~n49410 ;
  assign n49412 = \P1_P2_EAX_reg[10]/NET0131  & ~n49411 ;
  assign n49409 = ~n25826 & n47733 ;
  assign n49424 = \P1_P2_InstQueue_reg[8][2]/NET0131  & n25453 ;
  assign n49417 = \P1_P2_InstQueue_reg[9][2]/NET0131  & n25435 ;
  assign n49413 = \P1_P2_InstQueue_reg[12][2]/NET0131  & n25440 ;
  assign n49414 = \P1_P2_InstQueue_reg[2][2]/NET0131  & n25425 ;
  assign n49429 = ~n49413 & ~n49414 ;
  assign n49439 = ~n49417 & n49429 ;
  assign n49440 = ~n49424 & n49439 ;
  assign n49425 = \P1_P2_InstQueue_reg[15][2]/NET0131  & n25442 ;
  assign n49426 = \P1_P2_InstQueue_reg[11][2]/NET0131  & n25457 ;
  assign n49434 = ~n49425 & ~n49426 ;
  assign n49427 = \P1_P2_InstQueue_reg[6][2]/NET0131  & n25461 ;
  assign n49428 = \P1_P2_InstQueue_reg[3][2]/NET0131  & n25428 ;
  assign n49435 = ~n49427 & ~n49428 ;
  assign n49436 = n49434 & n49435 ;
  assign n49420 = \P1_P2_InstQueue_reg[10][2]/NET0131  & n25455 ;
  assign n49421 = \P1_P2_InstQueue_reg[7][2]/NET0131  & n25449 ;
  assign n49432 = ~n49420 & ~n49421 ;
  assign n49422 = \P1_P2_InstQueue_reg[1][2]/NET0131  & n25446 ;
  assign n49423 = \P1_P2_InstQueue_reg[14][2]/NET0131  & n25422 ;
  assign n49433 = ~n49422 & ~n49423 ;
  assign n49437 = n49432 & n49433 ;
  assign n49415 = \P1_P2_InstQueue_reg[4][2]/NET0131  & n25444 ;
  assign n49416 = \P1_P2_InstQueue_reg[0][2]/NET0131  & n25431 ;
  assign n49430 = ~n49415 & ~n49416 ;
  assign n49418 = \P1_P2_InstQueue_reg[13][2]/NET0131  & n25459 ;
  assign n49419 = \P1_P2_InstQueue_reg[5][2]/NET0131  & n25437 ;
  assign n49431 = ~n49418 & ~n49419 ;
  assign n49438 = n49430 & n49431 ;
  assign n49441 = n49437 & n49438 ;
  assign n49442 = n49436 & n49441 ;
  assign n49443 = n49440 & n49442 ;
  assign n49444 = n42875 & ~n49443 ;
  assign n49445 = n43179 & n49410 ;
  assign n49446 = ~n49444 & ~n49445 ;
  assign n49447 = ~n49409 & n49446 ;
  assign n49448 = ~n49412 & n49447 ;
  assign n49449 = n25918 & ~n49448 ;
  assign n49450 = ~n49408 & ~n49449 ;
  assign n49451 = \P1_P2_EAX_reg[11]/NET0131  & ~n43212 ;
  assign n49453 = \P1_P2_EAX_reg[11]/NET0131  & ~n49411 ;
  assign n49452 = ~n25826 & n44817 ;
  assign n49465 = \P1_P2_InstQueue_reg[8][3]/NET0131  & n25453 ;
  assign n49458 = \P1_P2_InstQueue_reg[9][3]/NET0131  & n25435 ;
  assign n49454 = \P1_P2_InstQueue_reg[2][3]/NET0131  & n25425 ;
  assign n49455 = \P1_P2_InstQueue_reg[3][3]/NET0131  & n25428 ;
  assign n49470 = ~n49454 & ~n49455 ;
  assign n49480 = ~n49458 & n49470 ;
  assign n49481 = ~n49465 & n49480 ;
  assign n49466 = \P1_P2_InstQueue_reg[4][3]/NET0131  & n25444 ;
  assign n49467 = \P1_P2_InstQueue_reg[12][3]/NET0131  & n25440 ;
  assign n49475 = ~n49466 & ~n49467 ;
  assign n49468 = \P1_P2_InstQueue_reg[15][3]/NET0131  & n25442 ;
  assign n49469 = \P1_P2_InstQueue_reg[11][3]/NET0131  & n25457 ;
  assign n49476 = ~n49468 & ~n49469 ;
  assign n49477 = n49475 & n49476 ;
  assign n49461 = \P1_P2_InstQueue_reg[14][3]/NET0131  & n25422 ;
  assign n49462 = \P1_P2_InstQueue_reg[5][3]/NET0131  & n25437 ;
  assign n49473 = ~n49461 & ~n49462 ;
  assign n49463 = \P1_P2_InstQueue_reg[1][3]/NET0131  & n25446 ;
  assign n49464 = \P1_P2_InstQueue_reg[7][3]/NET0131  & n25449 ;
  assign n49474 = ~n49463 & ~n49464 ;
  assign n49478 = n49473 & n49474 ;
  assign n49456 = \P1_P2_InstQueue_reg[10][3]/NET0131  & n25455 ;
  assign n49457 = \P1_P2_InstQueue_reg[0][3]/NET0131  & n25431 ;
  assign n49471 = ~n49456 & ~n49457 ;
  assign n49459 = \P1_P2_InstQueue_reg[6][3]/NET0131  & n25461 ;
  assign n49460 = \P1_P2_InstQueue_reg[13][3]/NET0131  & n25459 ;
  assign n49472 = ~n49459 & ~n49460 ;
  assign n49479 = n49471 & n49472 ;
  assign n49482 = n49478 & n49479 ;
  assign n49483 = n49477 & n49482 ;
  assign n49484 = n49481 & n49483 ;
  assign n49485 = n42875 & ~n49484 ;
  assign n49486 = ~\P1_P2_EAX_reg[11]/NET0131  & n43180 ;
  assign n49487 = n43164 & n49486 ;
  assign n49488 = ~n49485 & ~n49487 ;
  assign n49489 = ~n49452 & n49488 ;
  assign n49490 = ~n49453 & n49489 ;
  assign n49491 = n25918 & ~n49490 ;
  assign n49492 = ~n49451 & ~n49491 ;
  assign n49493 = \P1_P2_EAX_reg[12]/NET0131  & ~n43212 ;
  assign n49494 = n43164 & ~n43182 ;
  assign n49496 = ~n43167 & ~n49494 ;
  assign n49497 = \P1_P2_EAX_reg[12]/NET0131  & ~n49496 ;
  assign n49530 = \P1_P2_EAX_reg[12]/NET0131  & ~n25773 ;
  assign n49531 = ~n25770 & n47566 ;
  assign n49532 = ~n49530 & ~n49531 ;
  assign n49533 = ~n25826 & ~n49532 ;
  assign n49495 = n43181 & n49494 ;
  assign n49509 = \P1_P2_InstQueue_reg[8][4]/NET0131  & n25453 ;
  assign n49502 = \P1_P2_InstQueue_reg[9][4]/NET0131  & n25435 ;
  assign n49498 = \P1_P2_InstQueue_reg[15][4]/NET0131  & n25442 ;
  assign n49499 = \P1_P2_InstQueue_reg[3][4]/NET0131  & n25428 ;
  assign n49514 = ~n49498 & ~n49499 ;
  assign n49524 = ~n49502 & n49514 ;
  assign n49525 = ~n49509 & n49524 ;
  assign n49510 = \P1_P2_InstQueue_reg[2][4]/NET0131  & n25425 ;
  assign n49511 = \P1_P2_InstQueue_reg[4][4]/NET0131  & n25444 ;
  assign n49519 = ~n49510 & ~n49511 ;
  assign n49512 = \P1_P2_InstQueue_reg[12][4]/NET0131  & n25440 ;
  assign n49513 = \P1_P2_InstQueue_reg[7][4]/NET0131  & n25449 ;
  assign n49520 = ~n49512 & ~n49513 ;
  assign n49521 = n49519 & n49520 ;
  assign n49505 = \P1_P2_InstQueue_reg[6][4]/NET0131  & n25461 ;
  assign n49506 = \P1_P2_InstQueue_reg[10][4]/NET0131  & n25455 ;
  assign n49517 = ~n49505 & ~n49506 ;
  assign n49507 = \P1_P2_InstQueue_reg[1][4]/NET0131  & n25446 ;
  assign n49508 = \P1_P2_InstQueue_reg[14][4]/NET0131  & n25422 ;
  assign n49518 = ~n49507 & ~n49508 ;
  assign n49522 = n49517 & n49518 ;
  assign n49500 = \P1_P2_InstQueue_reg[11][4]/NET0131  & n25457 ;
  assign n49501 = \P1_P2_InstQueue_reg[0][4]/NET0131  & n25431 ;
  assign n49515 = ~n49500 & ~n49501 ;
  assign n49503 = \P1_P2_InstQueue_reg[13][4]/NET0131  & n25459 ;
  assign n49504 = \P1_P2_InstQueue_reg[5][4]/NET0131  & n25437 ;
  assign n49516 = ~n49503 & ~n49504 ;
  assign n49523 = n49515 & n49516 ;
  assign n49526 = n49522 & n49523 ;
  assign n49527 = n49521 & n49526 ;
  assign n49528 = n49525 & n49527 ;
  assign n49529 = n42875 & ~n49528 ;
  assign n49534 = ~n49495 & ~n49529 ;
  assign n49535 = ~n49533 & n49534 ;
  assign n49536 = ~n49497 & n49535 ;
  assign n49537 = n25918 & ~n49536 ;
  assign n49538 = ~n49493 & ~n49537 ;
  assign n49539 = \P1_P2_EAX_reg[13]/NET0131  & ~n43212 ;
  assign n49542 = \P1_P2_EAX_reg[13]/NET0131  & ~n49496 ;
  assign n49575 = \P1_P2_EAX_reg[13]/NET0131  & ~n25773 ;
  assign n49576 = ~n48347 & ~n49575 ;
  assign n49577 = ~n25826 & ~n49576 ;
  assign n49540 = ~\P1_P2_EAX_reg[13]/NET0131  & n43164 ;
  assign n49541 = n43182 & n49540 ;
  assign n49554 = \P1_P2_InstQueue_reg[8][5]/NET0131  & n25453 ;
  assign n49547 = \P1_P2_InstQueue_reg[9][5]/NET0131  & n25435 ;
  assign n49543 = \P1_P2_InstQueue_reg[7][5]/NET0131  & n25449 ;
  assign n49544 = \P1_P2_InstQueue_reg[4][5]/NET0131  & n25444 ;
  assign n49559 = ~n49543 & ~n49544 ;
  assign n49569 = ~n49547 & n49559 ;
  assign n49570 = ~n49554 & n49569 ;
  assign n49555 = \P1_P2_InstQueue_reg[11][5]/NET0131  & n25457 ;
  assign n49556 = \P1_P2_InstQueue_reg[10][5]/NET0131  & n25455 ;
  assign n49564 = ~n49555 & ~n49556 ;
  assign n49557 = \P1_P2_InstQueue_reg[3][5]/NET0131  & n25428 ;
  assign n49558 = \P1_P2_InstQueue_reg[14][5]/NET0131  & n25422 ;
  assign n49565 = ~n49557 & ~n49558 ;
  assign n49566 = n49564 & n49565 ;
  assign n49550 = \P1_P2_InstQueue_reg[6][5]/NET0131  & n25461 ;
  assign n49551 = \P1_P2_InstQueue_reg[5][5]/NET0131  & n25437 ;
  assign n49562 = ~n49550 & ~n49551 ;
  assign n49552 = \P1_P2_InstQueue_reg[1][5]/NET0131  & n25446 ;
  assign n49553 = \P1_P2_InstQueue_reg[15][5]/NET0131  & n25442 ;
  assign n49563 = ~n49552 & ~n49553 ;
  assign n49567 = n49562 & n49563 ;
  assign n49545 = \P1_P2_InstQueue_reg[12][5]/NET0131  & n25440 ;
  assign n49546 = \P1_P2_InstQueue_reg[0][5]/NET0131  & n25431 ;
  assign n49560 = ~n49545 & ~n49546 ;
  assign n49548 = \P1_P2_InstQueue_reg[2][5]/NET0131  & n25425 ;
  assign n49549 = \P1_P2_InstQueue_reg[13][5]/NET0131  & n25459 ;
  assign n49561 = ~n49548 & ~n49549 ;
  assign n49568 = n49560 & n49561 ;
  assign n49571 = n49567 & n49568 ;
  assign n49572 = n49566 & n49571 ;
  assign n49573 = n49570 & n49572 ;
  assign n49574 = n42875 & ~n49573 ;
  assign n49578 = ~n49541 & ~n49574 ;
  assign n49579 = ~n49577 & n49578 ;
  assign n49580 = ~n49542 & n49579 ;
  assign n49581 = n25918 & ~n49580 ;
  assign n49582 = ~n49539 & ~n49581 ;
  assign n49583 = \P1_P2_EAX_reg[14]/NET0131  & ~n43212 ;
  assign n49585 = \P1_P2_EAX_reg[14]/NET0131  & ~n48291 ;
  assign n49584 = n43183 & n48290 ;
  assign n49597 = \P1_P2_InstQueue_reg[8][6]/NET0131  & n25453 ;
  assign n49590 = \P1_P2_InstQueue_reg[9][6]/NET0131  & n25435 ;
  assign n49586 = \P1_P2_InstQueue_reg[2][6]/NET0131  & n25425 ;
  assign n49587 = \P1_P2_InstQueue_reg[15][6]/NET0131  & n25442 ;
  assign n49602 = ~n49586 & ~n49587 ;
  assign n49612 = ~n49590 & n49602 ;
  assign n49613 = ~n49597 & n49612 ;
  assign n49598 = \P1_P2_InstQueue_reg[12][6]/NET0131  & n25440 ;
  assign n49599 = \P1_P2_InstQueue_reg[10][6]/NET0131  & n25455 ;
  assign n49607 = ~n49598 & ~n49599 ;
  assign n49600 = \P1_P2_InstQueue_reg[13][6]/NET0131  & n25459 ;
  assign n49601 = \P1_P2_InstQueue_reg[14][6]/NET0131  & n25422 ;
  assign n49608 = ~n49600 & ~n49601 ;
  assign n49609 = n49607 & n49608 ;
  assign n49593 = \P1_P2_InstQueue_reg[7][6]/NET0131  & n25449 ;
  assign n49594 = \P1_P2_InstQueue_reg[11][6]/NET0131  & n25457 ;
  assign n49605 = ~n49593 & ~n49594 ;
  assign n49595 = \P1_P2_InstQueue_reg[1][6]/NET0131  & n25446 ;
  assign n49596 = \P1_P2_InstQueue_reg[6][6]/NET0131  & n25461 ;
  assign n49606 = ~n49595 & ~n49596 ;
  assign n49610 = n49605 & n49606 ;
  assign n49588 = \P1_P2_InstQueue_reg[4][6]/NET0131  & n25444 ;
  assign n49589 = \P1_P2_InstQueue_reg[0][6]/NET0131  & n25431 ;
  assign n49603 = ~n49588 & ~n49589 ;
  assign n49591 = \P1_P2_InstQueue_reg[5][6]/NET0131  & n25437 ;
  assign n49592 = \P1_P2_InstQueue_reg[3][6]/NET0131  & n25428 ;
  assign n49604 = ~n49591 & ~n49592 ;
  assign n49611 = n49603 & n49604 ;
  assign n49614 = n49610 & n49611 ;
  assign n49615 = n49609 & n49614 ;
  assign n49616 = n49613 & n49615 ;
  assign n49617 = n42875 & ~n49616 ;
  assign n49618 = \P1_P2_EAX_reg[14]/NET0131  & ~n25773 ;
  assign n49619 = ~n46685 & ~n49618 ;
  assign n49620 = ~n25826 & ~n49619 ;
  assign n49621 = ~n49617 & ~n49620 ;
  assign n49622 = ~n49584 & n49621 ;
  assign n49623 = ~n49585 & n49622 ;
  assign n49624 = n25918 & ~n49623 ;
  assign n49625 = ~n49583 & ~n49624 ;
  assign n49626 = n25918 & ~n43169 ;
  assign n49627 = n43212 & ~n49626 ;
  assign n49628 = \P1_P2_EAX_reg[7]/NET0131  & ~n49627 ;
  assign n49630 = ~n25415 & n25875 ;
  assign n49631 = ~n28931 & n49630 ;
  assign n49629 = ~n30809 & n42875 ;
  assign n49632 = ~\P1_P2_EAX_reg[7]/NET0131  & ~n43176 ;
  assign n49633 = ~n43177 & ~n49632 ;
  assign n49634 = n43164 & n49633 ;
  assign n49635 = ~n49629 & ~n49634 ;
  assign n49636 = ~n49631 & n49635 ;
  assign n49637 = n25918 & ~n49636 ;
  assign n49638 = ~n49628 & ~n49637 ;
  assign n49639 = \P2_P3_uWord_reg[8]/NET0131  & ~n47752 ;
  assign n49640 = \P2_buf2_reg[8]/NET0131  & n27122 ;
  assign n49641 = ~n27192 & n49640 ;
  assign n49642 = ~n48533 & ~n49641 ;
  assign n49643 = n47754 & ~n49642 ;
  assign n49644 = ~n49639 & ~n49643 ;
  assign n49645 = \P1_P2_EAX_reg[8]/NET0131  & ~n49627 ;
  assign n49678 = ~n48659 & n49630 ;
  assign n49657 = \P1_P2_InstQueue_reg[8][0]/NET0131  & n25453 ;
  assign n49650 = \P1_P2_InstQueue_reg[9][0]/NET0131  & n25435 ;
  assign n49646 = \P1_P2_InstQueue_reg[6][0]/NET0131  & n25461 ;
  assign n49647 = \P1_P2_InstQueue_reg[3][0]/NET0131  & n25428 ;
  assign n49662 = ~n49646 & ~n49647 ;
  assign n49672 = ~n49650 & n49662 ;
  assign n49673 = ~n49657 & n49672 ;
  assign n49658 = \P1_P2_InstQueue_reg[11][0]/NET0131  & n25457 ;
  assign n49659 = \P1_P2_InstQueue_reg[10][0]/NET0131  & n25455 ;
  assign n49667 = ~n49658 & ~n49659 ;
  assign n49660 = \P1_P2_InstQueue_reg[7][0]/NET0131  & n25449 ;
  assign n49661 = \P1_P2_InstQueue_reg[14][0]/NET0131  & n25422 ;
  assign n49668 = ~n49660 & ~n49661 ;
  assign n49669 = n49667 & n49668 ;
  assign n49653 = \P1_P2_InstQueue_reg[15][0]/NET0131  & n25442 ;
  assign n49654 = \P1_P2_InstQueue_reg[4][0]/NET0131  & n25444 ;
  assign n49665 = ~n49653 & ~n49654 ;
  assign n49655 = \P1_P2_InstQueue_reg[1][0]/NET0131  & n25446 ;
  assign n49656 = \P1_P2_InstQueue_reg[12][0]/NET0131  & n25440 ;
  assign n49666 = ~n49655 & ~n49656 ;
  assign n49670 = n49665 & n49666 ;
  assign n49648 = \P1_P2_InstQueue_reg[2][0]/NET0131  & n25425 ;
  assign n49649 = \P1_P2_InstQueue_reg[0][0]/NET0131  & n25431 ;
  assign n49663 = ~n49648 & ~n49649 ;
  assign n49651 = \P1_P2_InstQueue_reg[13][0]/NET0131  & n25459 ;
  assign n49652 = \P1_P2_InstQueue_reg[5][0]/NET0131  & n25437 ;
  assign n49664 = ~n49651 & ~n49652 ;
  assign n49671 = n49663 & n49664 ;
  assign n49674 = n49670 & n49671 ;
  assign n49675 = n49669 & n49674 ;
  assign n49676 = n49673 & n49675 ;
  assign n49677 = n42875 & ~n49676 ;
  assign n49679 = ~\P1_P2_EAX_reg[8]/NET0131  & ~n43177 ;
  assign n49680 = ~n43178 & ~n49679 ;
  assign n49681 = n43164 & n49680 ;
  assign n49682 = ~n49677 & ~n49681 ;
  assign n49683 = ~n49678 & n49682 ;
  assign n49684 = n25918 & ~n49683 ;
  assign n49685 = ~n49645 & ~n49684 ;
  assign n49686 = \P1_P2_EAX_reg[9]/NET0131  & ~n49627 ;
  assign n49719 = \P1_buf2_reg[9]/NET0131  & ~n27934 ;
  assign n49720 = \P1_buf1_reg[9]/NET0131  & n27934 ;
  assign n49721 = ~n49719 & ~n49720 ;
  assign n49722 = n49630 & ~n49721 ;
  assign n49698 = \P1_P2_InstQueue_reg[8][1]/NET0131  & n25453 ;
  assign n49691 = \P1_P2_InstQueue_reg[9][1]/NET0131  & n25435 ;
  assign n49687 = \P1_P2_InstQueue_reg[15][1]/NET0131  & n25442 ;
  assign n49688 = \P1_P2_InstQueue_reg[3][1]/NET0131  & n25428 ;
  assign n49703 = ~n49687 & ~n49688 ;
  assign n49713 = ~n49691 & n49703 ;
  assign n49714 = ~n49698 & n49713 ;
  assign n49699 = \P1_P2_InstQueue_reg[14][1]/NET0131  & n25422 ;
  assign n49700 = \P1_P2_InstQueue_reg[4][1]/NET0131  & n25444 ;
  assign n49708 = ~n49699 & ~n49700 ;
  assign n49701 = \P1_P2_InstQueue_reg[5][1]/NET0131  & n25437 ;
  assign n49702 = \P1_P2_InstQueue_reg[2][1]/NET0131  & n25425 ;
  assign n49709 = ~n49701 & ~n49702 ;
  assign n49710 = n49708 & n49709 ;
  assign n49694 = \P1_P2_InstQueue_reg[10][1]/NET0131  & n25455 ;
  assign n49695 = \P1_P2_InstQueue_reg[7][1]/NET0131  & n25449 ;
  assign n49706 = ~n49694 & ~n49695 ;
  assign n49696 = \P1_P2_InstQueue_reg[1][1]/NET0131  & n25446 ;
  assign n49697 = \P1_P2_InstQueue_reg[6][1]/NET0131  & n25461 ;
  assign n49707 = ~n49696 & ~n49697 ;
  assign n49711 = n49706 & n49707 ;
  assign n49689 = \P1_P2_InstQueue_reg[11][1]/NET0131  & n25457 ;
  assign n49690 = \P1_P2_InstQueue_reg[0][1]/NET0131  & n25431 ;
  assign n49704 = ~n49689 & ~n49690 ;
  assign n49692 = \P1_P2_InstQueue_reg[13][1]/NET0131  & n25459 ;
  assign n49693 = \P1_P2_InstQueue_reg[12][1]/NET0131  & n25440 ;
  assign n49705 = ~n49692 & ~n49693 ;
  assign n49712 = n49704 & n49705 ;
  assign n49715 = n49711 & n49712 ;
  assign n49716 = n49710 & n49715 ;
  assign n49717 = n49714 & n49716 ;
  assign n49718 = n42875 & ~n49717 ;
  assign n49723 = ~\P1_P2_EAX_reg[9]/NET0131  & ~n43178 ;
  assign n49724 = ~n43179 & ~n49723 ;
  assign n49725 = n43164 & n49724 ;
  assign n49726 = ~n49718 & ~n49725 ;
  assign n49727 = ~n49722 & n49726 ;
  assign n49728 = n25918 & ~n49727 ;
  assign n49729 = ~n49686 & ~n49728 ;
  assign n49730 = ~\P1_P3_InstQueueWr_Addr_reg[0]/NET0131  & ~\P1_P3_InstQueueWr_Addr_reg[1]/NET0131  ;
  assign n49731 = ~\P1_P3_InstQueueWr_Addr_reg[2]/NET0131  & n49730 ;
  assign n49732 = ~\P1_P3_InstQueueWr_Addr_reg[3]/NET0131  & n49731 ;
  assign n49753 = n8891 & n49732 ;
  assign n49752 = ~\P1_P3_InstQueue_reg[0][4]/NET0131  & ~n49732 ;
  assign n49754 = n10046 & ~n49752 ;
  assign n49755 = ~n49753 & n49754 ;
  assign n49733 = \P1_P3_InstQueueWr_Addr_reg[0]/NET0131  & \P1_P3_InstQueueWr_Addr_reg[1]/NET0131  ;
  assign n49734 = \P1_P3_InstQueueWr_Addr_reg[2]/NET0131  & n49733 ;
  assign n49735 = \P1_P3_InstQueueWr_Addr_reg[3]/NET0131  & n49734 ;
  assign n49736 = ~n49732 & ~n49735 ;
  assign n49737 = \P1_P3_InstQueueWr_Addr_reg[0]/NET0131  & ~\P1_P3_InstQueueWr_Addr_reg[1]/NET0131  ;
  assign n49738 = \P1_P3_InstQueueWr_Addr_reg[2]/NET0131  & n49737 ;
  assign n49739 = \P1_P3_InstQueueWr_Addr_reg[3]/NET0131  & n49738 ;
  assign n49740 = ~\P1_P3_InstQueueWr_Addr_reg[0]/NET0131  & \P1_P3_InstQueueWr_Addr_reg[1]/NET0131  ;
  assign n49741 = \P1_P3_InstQueueWr_Addr_reg[2]/NET0131  & n49740 ;
  assign n49742 = \P1_P3_InstQueueWr_Addr_reg[3]/NET0131  & n49741 ;
  assign n49743 = ~n49739 & ~n49742 ;
  assign n49744 = n9245 & n49743 ;
  assign n49745 = n36810 & ~n49744 ;
  assign n49746 = n49736 & ~n49745 ;
  assign n49747 = ~n9241 & ~n10036 ;
  assign n49748 = ~n21771 & n49747 ;
  assign n49749 = ~n10031 & n49748 ;
  assign n49750 = ~n49746 & n49749 ;
  assign n49751 = \P1_P3_InstQueue_reg[0][4]/NET0131  & ~n49750 ;
  assign n49756 = \P1_buf2_reg[28]/NET0131  & n49739 ;
  assign n49757 = \P1_buf2_reg[20]/NET0131  & n49742 ;
  assign n49758 = ~n49756 & ~n49757 ;
  assign n49759 = n11698 & ~n49758 ;
  assign n49760 = ~n49736 & ~n49745 ;
  assign n49761 = \P1_buf2_reg[4]/NET0131  & n49760 ;
  assign n49762 = ~n49759 & ~n49761 ;
  assign n49763 = ~n49751 & n49762 ;
  assign n49764 = ~n49755 & n49763 ;
  assign n49765 = ~\P1_P3_InstQueueWr_Addr_reg[2]/NET0131  & n49740 ;
  assign n49766 = \P1_P3_InstQueueWr_Addr_reg[3]/NET0131  & n49765 ;
  assign n49779 = n8891 & n49766 ;
  assign n49778 = ~\P1_P3_InstQueue_reg[10][4]/NET0131  & ~n49766 ;
  assign n49780 = n10046 & ~n49778 ;
  assign n49781 = ~n49779 & n49780 ;
  assign n49767 = ~\P1_P3_InstQueueWr_Addr_reg[2]/NET0131  & n49737 ;
  assign n49768 = \P1_P3_InstQueueWr_Addr_reg[3]/NET0131  & n49767 ;
  assign n49769 = ~n49766 & ~n49768 ;
  assign n49770 = ~\P1_P3_InstQueueWr_Addr_reg[3]/NET0131  & n49734 ;
  assign n49771 = \P1_P3_InstQueueWr_Addr_reg[3]/NET0131  & n49731 ;
  assign n49772 = ~n49770 & ~n49771 ;
  assign n49773 = n9245 & n49772 ;
  assign n49774 = n36810 & ~n49773 ;
  assign n49775 = n49769 & ~n49774 ;
  assign n49776 = n49749 & ~n49775 ;
  assign n49777 = \P1_P3_InstQueue_reg[10][4]/NET0131  & ~n49776 ;
  assign n49782 = \P1_buf2_reg[28]/NET0131  & n49770 ;
  assign n49783 = \P1_buf2_reg[20]/NET0131  & n49771 ;
  assign n49784 = ~n49782 & ~n49783 ;
  assign n49785 = n11698 & ~n49784 ;
  assign n49786 = ~n49769 & ~n49774 ;
  assign n49787 = \P1_buf2_reg[4]/NET0131  & n49786 ;
  assign n49788 = ~n49785 & ~n49787 ;
  assign n49789 = ~n49777 & n49788 ;
  assign n49790 = ~n49781 & n49789 ;
  assign n49791 = ~\P1_P3_InstQueueWr_Addr_reg[2]/NET0131  & n49733 ;
  assign n49792 = \P1_P3_InstQueueWr_Addr_reg[3]/NET0131  & n49791 ;
  assign n49801 = n8891 & n49792 ;
  assign n49800 = ~\P1_P3_InstQueue_reg[11][4]/NET0131  & ~n49792 ;
  assign n49802 = n10046 & ~n49800 ;
  assign n49803 = ~n49801 & n49802 ;
  assign n49793 = ~n49766 & ~n49792 ;
  assign n49794 = ~n49768 & ~n49771 ;
  assign n49795 = n9245 & n49794 ;
  assign n49796 = n36810 & ~n49795 ;
  assign n49797 = n49793 & ~n49796 ;
  assign n49798 = n49749 & ~n49797 ;
  assign n49799 = \P1_P3_InstQueue_reg[11][4]/NET0131  & ~n49798 ;
  assign n49804 = \P1_buf2_reg[28]/NET0131  & n49771 ;
  assign n49805 = \P1_buf2_reg[20]/NET0131  & n49768 ;
  assign n49806 = ~n49804 & ~n49805 ;
  assign n49807 = n11698 & ~n49806 ;
  assign n49808 = ~n49793 & ~n49796 ;
  assign n49809 = \P1_buf2_reg[4]/NET0131  & n49808 ;
  assign n49810 = ~n49807 & ~n49809 ;
  assign n49811 = ~n49799 & n49810 ;
  assign n49812 = ~n49803 & n49811 ;
  assign n49813 = \P1_P3_InstQueueWr_Addr_reg[2]/NET0131  & n49730 ;
  assign n49814 = \P1_P3_InstQueueWr_Addr_reg[3]/NET0131  & n49813 ;
  assign n49822 = n8891 & n49814 ;
  assign n49821 = ~\P1_P3_InstQueue_reg[12][4]/NET0131  & ~n49814 ;
  assign n49823 = n10046 & ~n49821 ;
  assign n49824 = ~n49822 & n49823 ;
  assign n49815 = ~n49792 & ~n49814 ;
  assign n49816 = n9245 & n49769 ;
  assign n49817 = n36810 & ~n49816 ;
  assign n49818 = n49815 & ~n49817 ;
  assign n49819 = n49749 & ~n49818 ;
  assign n49820 = \P1_P3_InstQueue_reg[12][4]/NET0131  & ~n49819 ;
  assign n49825 = \P1_buf2_reg[28]/NET0131  & n49768 ;
  assign n49826 = \P1_buf2_reg[20]/NET0131  & n49766 ;
  assign n49827 = ~n49825 & ~n49826 ;
  assign n49828 = n11698 & ~n49827 ;
  assign n49829 = ~n49815 & ~n49817 ;
  assign n49830 = \P1_buf2_reg[4]/NET0131  & n49829 ;
  assign n49831 = ~n49828 & ~n49830 ;
  assign n49832 = ~n49820 & n49831 ;
  assign n49833 = ~n49824 & n49832 ;
  assign n49841 = n8891 & n49739 ;
  assign n49840 = ~\P1_P3_InstQueue_reg[13][4]/NET0131  & ~n49739 ;
  assign n49842 = n10046 & ~n49840 ;
  assign n49843 = ~n49841 & n49842 ;
  assign n49834 = ~n49739 & ~n49814 ;
  assign n49835 = n9245 & n49793 ;
  assign n49836 = n36810 & ~n49835 ;
  assign n49837 = n49834 & ~n49836 ;
  assign n49838 = n49749 & ~n49837 ;
  assign n49839 = \P1_P3_InstQueue_reg[13][4]/NET0131  & ~n49838 ;
  assign n49844 = \P1_buf2_reg[28]/NET0131  & n49766 ;
  assign n49845 = \P1_buf2_reg[20]/NET0131  & n49792 ;
  assign n49846 = ~n49844 & ~n49845 ;
  assign n49847 = n11698 & ~n49846 ;
  assign n49848 = ~n49834 & ~n49836 ;
  assign n49849 = \P1_buf2_reg[4]/NET0131  & n49848 ;
  assign n49850 = ~n49847 & ~n49849 ;
  assign n49851 = ~n49839 & n49850 ;
  assign n49852 = ~n49843 & n49851 ;
  assign n49859 = n8891 & n49742 ;
  assign n49858 = ~\P1_P3_InstQueue_reg[14][4]/NET0131  & ~n49742 ;
  assign n49860 = n10046 & ~n49858 ;
  assign n49861 = ~n49859 & n49860 ;
  assign n49853 = n9245 & n49815 ;
  assign n49854 = n36810 & ~n49853 ;
  assign n49855 = n49743 & ~n49854 ;
  assign n49856 = n49749 & ~n49855 ;
  assign n49857 = \P1_P3_InstQueue_reg[14][4]/NET0131  & ~n49856 ;
  assign n49862 = \P1_buf2_reg[28]/NET0131  & n49792 ;
  assign n49863 = \P1_buf2_reg[20]/NET0131  & n49814 ;
  assign n49864 = ~n49862 & ~n49863 ;
  assign n49865 = n11698 & ~n49864 ;
  assign n49866 = ~n49743 & ~n49854 ;
  assign n49867 = \P1_buf2_reg[4]/NET0131  & n49866 ;
  assign n49868 = ~n49865 & ~n49867 ;
  assign n49869 = ~n49857 & n49868 ;
  assign n49870 = ~n49861 & n49869 ;
  assign n49878 = n8891 & n49735 ;
  assign n49877 = ~\P1_P3_InstQueue_reg[15][4]/NET0131  & ~n49735 ;
  assign n49879 = n10046 & ~n49877 ;
  assign n49880 = ~n49878 & n49879 ;
  assign n49871 = ~n49735 & ~n49742 ;
  assign n49872 = n9245 & n49834 ;
  assign n49873 = n36810 & ~n49872 ;
  assign n49874 = n49871 & ~n49873 ;
  assign n49875 = n49749 & ~n49874 ;
  assign n49876 = \P1_P3_InstQueue_reg[15][4]/NET0131  & ~n49875 ;
  assign n49881 = \P1_buf2_reg[28]/NET0131  & n49814 ;
  assign n49882 = \P1_buf2_reg[20]/NET0131  & n49739 ;
  assign n49883 = ~n49881 & ~n49882 ;
  assign n49884 = n11698 & ~n49883 ;
  assign n49885 = ~n49871 & ~n49873 ;
  assign n49886 = \P1_buf2_reg[4]/NET0131  & n49885 ;
  assign n49887 = ~n49884 & ~n49886 ;
  assign n49888 = ~n49876 & n49887 ;
  assign n49889 = ~n49880 & n49888 ;
  assign n49890 = ~\P1_P3_InstQueueWr_Addr_reg[3]/NET0131  & n49767 ;
  assign n49898 = n8891 & n49890 ;
  assign n49897 = ~\P1_P3_InstQueue_reg[1][4]/NET0131  & ~n49890 ;
  assign n49899 = n10046 & ~n49897 ;
  assign n49900 = ~n49898 & n49899 ;
  assign n49891 = ~n49732 & ~n49890 ;
  assign n49892 = n9245 & n49871 ;
  assign n49893 = n36810 & ~n49892 ;
  assign n49894 = n49891 & ~n49893 ;
  assign n49895 = n49749 & ~n49894 ;
  assign n49896 = \P1_P3_InstQueue_reg[1][4]/NET0131  & ~n49895 ;
  assign n49901 = \P1_buf2_reg[28]/NET0131  & n49742 ;
  assign n49902 = \P1_buf2_reg[20]/NET0131  & n49735 ;
  assign n49903 = ~n49901 & ~n49902 ;
  assign n49904 = n11698 & ~n49903 ;
  assign n49905 = ~n49891 & ~n49893 ;
  assign n49906 = \P1_buf2_reg[4]/NET0131  & n49905 ;
  assign n49907 = ~n49904 & ~n49906 ;
  assign n49908 = ~n49896 & n49907 ;
  assign n49909 = ~n49900 & n49908 ;
  assign n49910 = ~\P1_P3_InstQueueWr_Addr_reg[3]/NET0131  & n49765 ;
  assign n49918 = n8891 & n49910 ;
  assign n49917 = ~\P1_P3_InstQueue_reg[2][4]/NET0131  & ~n49910 ;
  assign n49919 = n10046 & ~n49917 ;
  assign n49920 = ~n49918 & n49919 ;
  assign n49911 = ~n49890 & ~n49910 ;
  assign n49912 = n9245 & n49736 ;
  assign n49913 = n36810 & ~n49912 ;
  assign n49914 = n49911 & ~n49913 ;
  assign n49915 = n49749 & ~n49914 ;
  assign n49916 = \P1_P3_InstQueue_reg[2][4]/NET0131  & ~n49915 ;
  assign n49921 = \P1_buf2_reg[28]/NET0131  & n49735 ;
  assign n49922 = \P1_buf2_reg[20]/NET0131  & n49732 ;
  assign n49923 = ~n49921 & ~n49922 ;
  assign n49924 = n11698 & ~n49923 ;
  assign n49925 = ~n49911 & ~n49913 ;
  assign n49926 = \P1_buf2_reg[4]/NET0131  & n49925 ;
  assign n49927 = ~n49924 & ~n49926 ;
  assign n49928 = ~n49916 & n49927 ;
  assign n49929 = ~n49920 & n49928 ;
  assign n49930 = ~\P1_P3_InstQueueWr_Addr_reg[3]/NET0131  & n49791 ;
  assign n49938 = n8891 & n49930 ;
  assign n49937 = ~\P1_P3_InstQueue_reg[3][4]/NET0131  & ~n49930 ;
  assign n49939 = n10046 & ~n49937 ;
  assign n49940 = ~n49938 & n49939 ;
  assign n49931 = ~n49910 & ~n49930 ;
  assign n49932 = n9245 & n49891 ;
  assign n49933 = n36810 & ~n49932 ;
  assign n49934 = n49931 & ~n49933 ;
  assign n49935 = n49749 & ~n49934 ;
  assign n49936 = \P1_P3_InstQueue_reg[3][4]/NET0131  & ~n49935 ;
  assign n49941 = \P1_buf2_reg[28]/NET0131  & n49732 ;
  assign n49942 = \P1_buf2_reg[20]/NET0131  & n49890 ;
  assign n49943 = ~n49941 & ~n49942 ;
  assign n49944 = n11698 & ~n49943 ;
  assign n49945 = ~n49931 & ~n49933 ;
  assign n49946 = \P1_buf2_reg[4]/NET0131  & n49945 ;
  assign n49947 = ~n49944 & ~n49946 ;
  assign n49948 = ~n49936 & n49947 ;
  assign n49949 = ~n49940 & n49948 ;
  assign n49950 = ~\P1_P3_InstQueueWr_Addr_reg[3]/NET0131  & n49813 ;
  assign n49958 = n8891 & n49950 ;
  assign n49957 = ~\P1_P3_InstQueue_reg[4][4]/NET0131  & ~n49950 ;
  assign n49959 = n10046 & ~n49957 ;
  assign n49960 = ~n49958 & n49959 ;
  assign n49951 = ~n49930 & ~n49950 ;
  assign n49952 = n9245 & n49911 ;
  assign n49953 = n36810 & ~n49952 ;
  assign n49954 = n49951 & ~n49953 ;
  assign n49955 = n49749 & ~n49954 ;
  assign n49956 = \P1_P3_InstQueue_reg[4][4]/NET0131  & ~n49955 ;
  assign n49961 = \P1_buf2_reg[28]/NET0131  & n49890 ;
  assign n49962 = \P1_buf2_reg[20]/NET0131  & n49910 ;
  assign n49963 = ~n49961 & ~n49962 ;
  assign n49964 = n11698 & ~n49963 ;
  assign n49965 = ~n49951 & ~n49953 ;
  assign n49966 = \P1_buf2_reg[4]/NET0131  & n49965 ;
  assign n49967 = ~n49964 & ~n49966 ;
  assign n49968 = ~n49956 & n49967 ;
  assign n49969 = ~n49960 & n49968 ;
  assign n49970 = ~\P1_P3_InstQueueWr_Addr_reg[3]/NET0131  & n49738 ;
  assign n49978 = n8891 & n49970 ;
  assign n49977 = ~\P1_P3_InstQueue_reg[5][4]/NET0131  & ~n49970 ;
  assign n49979 = n10046 & ~n49977 ;
  assign n49980 = ~n49978 & n49979 ;
  assign n49971 = ~n49950 & ~n49970 ;
  assign n49972 = n9245 & n49931 ;
  assign n49973 = n36810 & ~n49972 ;
  assign n49974 = n49971 & ~n49973 ;
  assign n49975 = n49749 & ~n49974 ;
  assign n49976 = \P1_P3_InstQueue_reg[5][4]/NET0131  & ~n49975 ;
  assign n49981 = \P1_buf2_reg[28]/NET0131  & n49910 ;
  assign n49982 = \P1_buf2_reg[20]/NET0131  & n49930 ;
  assign n49983 = ~n49981 & ~n49982 ;
  assign n49984 = n11698 & ~n49983 ;
  assign n49985 = ~n49971 & ~n49973 ;
  assign n49986 = \P1_buf2_reg[4]/NET0131  & n49985 ;
  assign n49987 = ~n49984 & ~n49986 ;
  assign n49988 = ~n49976 & n49987 ;
  assign n49989 = ~n49980 & n49988 ;
  assign n49990 = ~\P1_P3_InstQueueWr_Addr_reg[3]/NET0131  & n49741 ;
  assign n49998 = n8891 & n49990 ;
  assign n49997 = ~\P1_P3_InstQueue_reg[6][4]/NET0131  & ~n49990 ;
  assign n49999 = n10046 & ~n49997 ;
  assign n50000 = ~n49998 & n49999 ;
  assign n49991 = ~n49970 & ~n49990 ;
  assign n49992 = n9245 & n49951 ;
  assign n49993 = n36810 & ~n49992 ;
  assign n49994 = n49991 & ~n49993 ;
  assign n49995 = n49749 & ~n49994 ;
  assign n49996 = \P1_P3_InstQueue_reg[6][4]/NET0131  & ~n49995 ;
  assign n50001 = \P1_buf2_reg[28]/NET0131  & n49930 ;
  assign n50002 = \P1_buf2_reg[20]/NET0131  & n49950 ;
  assign n50003 = ~n50001 & ~n50002 ;
  assign n50004 = n11698 & ~n50003 ;
  assign n50005 = ~n49991 & ~n49993 ;
  assign n50006 = \P1_buf2_reg[4]/NET0131  & n50005 ;
  assign n50007 = ~n50004 & ~n50006 ;
  assign n50008 = ~n49996 & n50007 ;
  assign n50009 = ~n50000 & n50008 ;
  assign n50019 = ~\P2_P3_InstQueueWr_Addr_reg[0]/NET0131  & ~\P2_P3_InstQueueWr_Addr_reg[1]/NET0131  ;
  assign n50020 = ~\P2_P3_InstQueueWr_Addr_reg[2]/NET0131  & n50019 ;
  assign n50021 = ~\P2_P3_InstQueueWr_Addr_reg[3]/NET0131  & n50020 ;
  assign n50033 = n27091 & n50021 ;
  assign n50032 = ~\P2_P3_InstQueue_reg[0][4]/NET0131  & ~n50021 ;
  assign n50034 = n27788 & ~n50032 ;
  assign n50035 = ~n50033 & n50034 ;
  assign n50010 = \P2_P3_InstQueueWr_Addr_reg[0]/NET0131  & ~\P2_P3_InstQueueWr_Addr_reg[1]/NET0131  ;
  assign n50011 = \P2_P3_InstQueueWr_Addr_reg[2]/NET0131  & n50010 ;
  assign n50012 = \P2_P3_InstQueueWr_Addr_reg[3]/NET0131  & n50011 ;
  assign n50013 = ~\P2_P3_InstQueueWr_Addr_reg[0]/NET0131  & \P2_P3_InstQueueWr_Addr_reg[1]/NET0131  ;
  assign n50014 = \P2_P3_InstQueueWr_Addr_reg[2]/NET0131  & n50013 ;
  assign n50015 = \P2_P3_InstQueueWr_Addr_reg[3]/NET0131  & n50014 ;
  assign n50016 = ~n50012 & ~n50015 ;
  assign n50017 = n27315 & n50016 ;
  assign n50018 = n36831 & ~n50017 ;
  assign n50022 = \P2_P3_InstQueueWr_Addr_reg[0]/NET0131  & \P2_P3_InstQueueWr_Addr_reg[1]/NET0131  ;
  assign n50023 = \P2_P3_InstQueueWr_Addr_reg[2]/NET0131  & n50022 ;
  assign n50024 = \P2_P3_InstQueueWr_Addr_reg[3]/NET0131  & n50023 ;
  assign n50025 = ~n50021 & ~n50024 ;
  assign n50026 = ~n50018 & n50025 ;
  assign n50027 = ~n27308 & ~n27656 ;
  assign n50028 = ~n27326 & n50027 ;
  assign n50029 = n43270 & n50028 ;
  assign n50030 = ~n50026 & n50029 ;
  assign n50031 = \P2_P3_InstQueue_reg[0][4]/NET0131  & ~n50030 ;
  assign n50036 = \P2_buf2_reg[28]/NET0131  & n50012 ;
  assign n50037 = \P2_buf2_reg[20]/NET0131  & n50015 ;
  assign n50038 = ~n50036 & ~n50037 ;
  assign n50039 = n27325 & ~n50038 ;
  assign n50040 = ~n50018 & ~n50025 ;
  assign n50041 = \P2_buf2_reg[4]/NET0131  & n50040 ;
  assign n50042 = ~n50039 & ~n50041 ;
  assign n50043 = ~n50031 & n50042 ;
  assign n50044 = ~n50035 & n50043 ;
  assign n50050 = ~\P2_P3_InstQueueWr_Addr_reg[2]/NET0131  & n50013 ;
  assign n50051 = \P2_P3_InstQueueWr_Addr_reg[3]/NET0131  & n50050 ;
  assign n50059 = n27091 & n50051 ;
  assign n50058 = ~\P2_P3_InstQueue_reg[10][4]/NET0131  & ~n50051 ;
  assign n50060 = n27788 & ~n50058 ;
  assign n50061 = ~n50059 & n50060 ;
  assign n50045 = \P2_P3_InstQueueWr_Addr_reg[3]/NET0131  & n50020 ;
  assign n50046 = ~\P2_P3_InstQueueWr_Addr_reg[3]/NET0131  & n50023 ;
  assign n50047 = ~n50045 & ~n50046 ;
  assign n50048 = n27315 & n50047 ;
  assign n50049 = n36831 & ~n50048 ;
  assign n50052 = ~\P2_P3_InstQueueWr_Addr_reg[2]/NET0131  & n50010 ;
  assign n50053 = \P2_P3_InstQueueWr_Addr_reg[3]/NET0131  & n50052 ;
  assign n50054 = ~n50051 & ~n50053 ;
  assign n50055 = ~n50049 & n50054 ;
  assign n50056 = n50029 & ~n50055 ;
  assign n50057 = \P2_P3_InstQueue_reg[10][4]/NET0131  & ~n50056 ;
  assign n50062 = \P2_buf2_reg[20]/NET0131  & n50045 ;
  assign n50063 = \P2_buf2_reg[28]/NET0131  & n50046 ;
  assign n50064 = ~n50062 & ~n50063 ;
  assign n50065 = n27325 & ~n50064 ;
  assign n50066 = ~n50049 & ~n50054 ;
  assign n50067 = \P2_buf2_reg[4]/NET0131  & n50066 ;
  assign n50068 = ~n50065 & ~n50067 ;
  assign n50069 = ~n50057 & n50068 ;
  assign n50070 = ~n50061 & n50069 ;
  assign n50078 = n8891 & n49770 ;
  assign n50077 = ~\P1_P3_InstQueue_reg[7][4]/NET0131  & ~n49770 ;
  assign n50079 = n10046 & ~n50077 ;
  assign n50080 = ~n50078 & n50079 ;
  assign n50071 = ~n49770 & ~n49990 ;
  assign n50072 = n9245 & n49971 ;
  assign n50073 = n36810 & ~n50072 ;
  assign n50074 = n50071 & ~n50073 ;
  assign n50075 = n49749 & ~n50074 ;
  assign n50076 = \P1_P3_InstQueue_reg[7][4]/NET0131  & ~n50075 ;
  assign n50081 = \P1_buf2_reg[28]/NET0131  & n49950 ;
  assign n50082 = \P1_buf2_reg[20]/NET0131  & n49970 ;
  assign n50083 = ~n50081 & ~n50082 ;
  assign n50084 = n11698 & ~n50083 ;
  assign n50085 = ~n50071 & ~n50073 ;
  assign n50086 = \P1_buf2_reg[4]/NET0131  & n50085 ;
  assign n50087 = ~n50084 & ~n50086 ;
  assign n50088 = ~n50076 & n50087 ;
  assign n50089 = ~n50080 & n50088 ;
  assign n50093 = ~\P2_P3_InstQueueWr_Addr_reg[2]/NET0131  & n50022 ;
  assign n50094 = \P2_P3_InstQueueWr_Addr_reg[3]/NET0131  & n50093 ;
  assign n50100 = n27091 & n50094 ;
  assign n50099 = ~\P2_P3_InstQueue_reg[11][4]/NET0131  & ~n50094 ;
  assign n50101 = n27788 & ~n50099 ;
  assign n50102 = ~n50100 & n50101 ;
  assign n50090 = ~n50045 & ~n50053 ;
  assign n50091 = n27315 & n50090 ;
  assign n50092 = n36831 & ~n50091 ;
  assign n50095 = ~n50051 & ~n50094 ;
  assign n50096 = ~n50092 & n50095 ;
  assign n50097 = n50029 & ~n50096 ;
  assign n50098 = \P2_P3_InstQueue_reg[11][4]/NET0131  & ~n50097 ;
  assign n50103 = \P2_buf2_reg[28]/NET0131  & n50045 ;
  assign n50104 = \P2_buf2_reg[20]/NET0131  & n50053 ;
  assign n50105 = ~n50103 & ~n50104 ;
  assign n50106 = n27325 & ~n50105 ;
  assign n50107 = ~n50092 & ~n50095 ;
  assign n50108 = \P2_buf2_reg[4]/NET0131  & n50107 ;
  assign n50109 = ~n50106 & ~n50108 ;
  assign n50110 = ~n50098 & n50109 ;
  assign n50111 = ~n50102 & n50110 ;
  assign n50114 = \P2_P3_InstQueueWr_Addr_reg[2]/NET0131  & n50019 ;
  assign n50115 = \P2_P3_InstQueueWr_Addr_reg[3]/NET0131  & n50114 ;
  assign n50121 = n27091 & n50115 ;
  assign n50120 = ~\P2_P3_InstQueue_reg[12][4]/NET0131  & ~n50115 ;
  assign n50122 = n27788 & ~n50120 ;
  assign n50123 = ~n50121 & n50122 ;
  assign n50112 = n27315 & n50054 ;
  assign n50113 = n36831 & ~n50112 ;
  assign n50116 = ~n50094 & ~n50115 ;
  assign n50117 = ~n50113 & n50116 ;
  assign n50118 = n50029 & ~n50117 ;
  assign n50119 = \P2_P3_InstQueue_reg[12][4]/NET0131  & ~n50118 ;
  assign n50124 = \P2_buf2_reg[28]/NET0131  & n50053 ;
  assign n50125 = \P2_buf2_reg[20]/NET0131  & n50051 ;
  assign n50126 = ~n50124 & ~n50125 ;
  assign n50127 = n27325 & ~n50126 ;
  assign n50128 = ~n50113 & ~n50116 ;
  assign n50129 = \P2_buf2_reg[4]/NET0131  & n50128 ;
  assign n50130 = ~n50127 & ~n50129 ;
  assign n50131 = ~n50119 & n50130 ;
  assign n50132 = ~n50123 & n50131 ;
  assign n50139 = n8891 & n49771 ;
  assign n50138 = ~\P1_P3_InstQueue_reg[8][4]/NET0131  & ~n49771 ;
  assign n50140 = n10046 & ~n50138 ;
  assign n50141 = ~n50139 & n50140 ;
  assign n50133 = n9245 & n49991 ;
  assign n50134 = n36810 & ~n50133 ;
  assign n50135 = n49772 & ~n50134 ;
  assign n50136 = n49749 & ~n50135 ;
  assign n50137 = \P1_P3_InstQueue_reg[8][4]/NET0131  & ~n50136 ;
  assign n50142 = \P1_buf2_reg[28]/NET0131  & n49970 ;
  assign n50143 = \P1_buf2_reg[20]/NET0131  & n49990 ;
  assign n50144 = ~n50142 & ~n50143 ;
  assign n50145 = n11698 & ~n50144 ;
  assign n50146 = ~n49772 & ~n50134 ;
  assign n50147 = \P1_buf2_reg[4]/NET0131  & n50146 ;
  assign n50148 = ~n50145 & ~n50147 ;
  assign n50149 = ~n50137 & n50148 ;
  assign n50150 = ~n50141 & n50149 ;
  assign n50158 = n27091 & n50012 ;
  assign n50157 = ~\P2_P3_InstQueue_reg[13][4]/NET0131  & ~n50012 ;
  assign n50159 = n27788 & ~n50157 ;
  assign n50160 = ~n50158 & n50159 ;
  assign n50151 = n27315 & n50095 ;
  assign n50152 = n36831 & ~n50151 ;
  assign n50153 = ~n50012 & ~n50115 ;
  assign n50154 = ~n50152 & n50153 ;
  assign n50155 = n50029 & ~n50154 ;
  assign n50156 = \P2_P3_InstQueue_reg[13][4]/NET0131  & ~n50155 ;
  assign n50161 = \P2_buf2_reg[28]/NET0131  & n50051 ;
  assign n50162 = \P2_buf2_reg[20]/NET0131  & n50094 ;
  assign n50163 = ~n50161 & ~n50162 ;
  assign n50164 = n27325 & ~n50163 ;
  assign n50165 = ~n50152 & ~n50153 ;
  assign n50166 = \P2_buf2_reg[4]/NET0131  & n50165 ;
  assign n50167 = ~n50164 & ~n50166 ;
  assign n50168 = ~n50156 & n50167 ;
  assign n50169 = ~n50160 & n50168 ;
  assign n50176 = n27091 & n50015 ;
  assign n50175 = ~\P2_P3_InstQueue_reg[14][4]/NET0131  & ~n50015 ;
  assign n50177 = n27788 & ~n50175 ;
  assign n50178 = ~n50176 & n50177 ;
  assign n50170 = n27315 & n50116 ;
  assign n50171 = n36831 & ~n50170 ;
  assign n50172 = n50016 & ~n50171 ;
  assign n50173 = n50029 & ~n50172 ;
  assign n50174 = \P2_P3_InstQueue_reg[14][4]/NET0131  & ~n50173 ;
  assign n50179 = \P2_buf2_reg[28]/NET0131  & n50094 ;
  assign n50180 = \P2_buf2_reg[20]/NET0131  & n50115 ;
  assign n50181 = ~n50179 & ~n50180 ;
  assign n50182 = n27325 & ~n50181 ;
  assign n50183 = ~n50016 & ~n50171 ;
  assign n50184 = \P2_buf2_reg[4]/NET0131  & n50183 ;
  assign n50185 = ~n50182 & ~n50184 ;
  assign n50186 = ~n50174 & n50185 ;
  assign n50187 = ~n50178 & n50186 ;
  assign n50194 = n8891 & n49768 ;
  assign n50193 = ~\P1_P3_InstQueue_reg[9][4]/NET0131  & ~n49768 ;
  assign n50195 = n10046 & ~n50193 ;
  assign n50196 = ~n50194 & n50195 ;
  assign n50188 = n9245 & n50071 ;
  assign n50189 = n36810 & ~n50188 ;
  assign n50190 = n49794 & ~n50189 ;
  assign n50191 = n49749 & ~n50190 ;
  assign n50192 = \P1_P3_InstQueue_reg[9][4]/NET0131  & ~n50191 ;
  assign n50197 = \P1_buf2_reg[28]/NET0131  & n49990 ;
  assign n50198 = \P1_buf2_reg[20]/NET0131  & n49770 ;
  assign n50199 = ~n50197 & ~n50198 ;
  assign n50200 = n11698 & ~n50199 ;
  assign n50201 = ~n49794 & ~n50189 ;
  assign n50202 = \P1_buf2_reg[4]/NET0131  & n50201 ;
  assign n50203 = ~n50200 & ~n50202 ;
  assign n50204 = ~n50192 & n50203 ;
  assign n50205 = ~n50196 & n50204 ;
  assign n50213 = n27091 & n50024 ;
  assign n50212 = ~\P2_P3_InstQueue_reg[15][4]/NET0131  & ~n50024 ;
  assign n50214 = n27788 & ~n50212 ;
  assign n50215 = ~n50213 & n50214 ;
  assign n50206 = n27315 & n50153 ;
  assign n50207 = n36831 & ~n50206 ;
  assign n50208 = ~n50015 & ~n50024 ;
  assign n50209 = ~n50207 & n50208 ;
  assign n50210 = n50029 & ~n50209 ;
  assign n50211 = \P2_P3_InstQueue_reg[15][4]/NET0131  & ~n50210 ;
  assign n50216 = \P2_buf2_reg[28]/NET0131  & n50115 ;
  assign n50217 = \P2_buf2_reg[20]/NET0131  & n50012 ;
  assign n50218 = ~n50216 & ~n50217 ;
  assign n50219 = n27325 & ~n50218 ;
  assign n50220 = ~n50207 & ~n50208 ;
  assign n50221 = \P2_buf2_reg[4]/NET0131  & n50220 ;
  assign n50222 = ~n50219 & ~n50221 ;
  assign n50223 = ~n50211 & n50222 ;
  assign n50224 = ~n50215 & n50223 ;
  assign n50227 = ~\P2_P3_InstQueueWr_Addr_reg[3]/NET0131  & n50052 ;
  assign n50233 = n27091 & n50227 ;
  assign n50232 = ~\P2_P3_InstQueue_reg[1][4]/NET0131  & ~n50227 ;
  assign n50234 = n27788 & ~n50232 ;
  assign n50235 = ~n50233 & n50234 ;
  assign n50225 = n27315 & n50208 ;
  assign n50226 = n36831 & ~n50225 ;
  assign n50228 = ~n50021 & ~n50227 ;
  assign n50229 = ~n50226 & n50228 ;
  assign n50230 = n50029 & ~n50229 ;
  assign n50231 = \P2_P3_InstQueue_reg[1][4]/NET0131  & ~n50230 ;
  assign n50236 = \P2_buf2_reg[28]/NET0131  & n50015 ;
  assign n50237 = \P2_buf2_reg[20]/NET0131  & n50024 ;
  assign n50238 = ~n50236 & ~n50237 ;
  assign n50239 = n27325 & ~n50238 ;
  assign n50240 = ~n50226 & ~n50228 ;
  assign n50241 = \P2_buf2_reg[4]/NET0131  & n50240 ;
  assign n50242 = ~n50239 & ~n50241 ;
  assign n50243 = ~n50231 & n50242 ;
  assign n50244 = ~n50235 & n50243 ;
  assign n50247 = ~\P2_P3_InstQueueWr_Addr_reg[3]/NET0131  & n50050 ;
  assign n50253 = n27091 & n50247 ;
  assign n50252 = ~\P2_P3_InstQueue_reg[2][4]/NET0131  & ~n50247 ;
  assign n50254 = n27788 & ~n50252 ;
  assign n50255 = ~n50253 & n50254 ;
  assign n50245 = n27315 & n50025 ;
  assign n50246 = n36831 & ~n50245 ;
  assign n50248 = ~n50227 & ~n50247 ;
  assign n50249 = ~n50246 & n50248 ;
  assign n50250 = n50029 & ~n50249 ;
  assign n50251 = \P2_P3_InstQueue_reg[2][4]/NET0131  & ~n50250 ;
  assign n50256 = \P2_buf2_reg[20]/NET0131  & n50021 ;
  assign n50257 = \P2_buf2_reg[28]/NET0131  & n50024 ;
  assign n50258 = ~n50256 & ~n50257 ;
  assign n50259 = n27325 & ~n50258 ;
  assign n50260 = ~n50246 & ~n50248 ;
  assign n50261 = \P2_buf2_reg[4]/NET0131  & n50260 ;
  assign n50262 = ~n50259 & ~n50261 ;
  assign n50263 = ~n50251 & n50262 ;
  assign n50264 = ~n50255 & n50263 ;
  assign n50267 = ~\P2_P3_InstQueueWr_Addr_reg[3]/NET0131  & n50093 ;
  assign n50273 = n27091 & n50267 ;
  assign n50272 = ~\P2_P3_InstQueue_reg[3][4]/NET0131  & ~n50267 ;
  assign n50274 = n27788 & ~n50272 ;
  assign n50275 = ~n50273 & n50274 ;
  assign n50265 = n27315 & n50228 ;
  assign n50266 = n36831 & ~n50265 ;
  assign n50268 = ~n50247 & ~n50267 ;
  assign n50269 = ~n50266 & n50268 ;
  assign n50270 = n50029 & ~n50269 ;
  assign n50271 = \P2_P3_InstQueue_reg[3][4]/NET0131  & ~n50270 ;
  assign n50276 = \P2_buf2_reg[28]/NET0131  & n50021 ;
  assign n50277 = \P2_buf2_reg[20]/NET0131  & n50227 ;
  assign n50278 = ~n50276 & ~n50277 ;
  assign n50279 = n27325 & ~n50278 ;
  assign n50280 = ~n50266 & ~n50268 ;
  assign n50281 = \P2_buf2_reg[4]/NET0131  & n50280 ;
  assign n50282 = ~n50279 & ~n50281 ;
  assign n50283 = ~n50271 & n50282 ;
  assign n50284 = ~n50275 & n50283 ;
  assign n50287 = ~\P2_P3_InstQueueWr_Addr_reg[3]/NET0131  & n50114 ;
  assign n50293 = n27091 & n50287 ;
  assign n50292 = ~\P2_P3_InstQueue_reg[4][4]/NET0131  & ~n50287 ;
  assign n50294 = n27788 & ~n50292 ;
  assign n50295 = ~n50293 & n50294 ;
  assign n50285 = n27315 & n50248 ;
  assign n50286 = n36831 & ~n50285 ;
  assign n50288 = ~n50267 & ~n50287 ;
  assign n50289 = ~n50286 & n50288 ;
  assign n50290 = n50029 & ~n50289 ;
  assign n50291 = \P2_P3_InstQueue_reg[4][4]/NET0131  & ~n50290 ;
  assign n50296 = \P2_buf2_reg[28]/NET0131  & n50227 ;
  assign n50297 = \P2_buf2_reg[20]/NET0131  & n50247 ;
  assign n50298 = ~n50296 & ~n50297 ;
  assign n50299 = n27325 & ~n50298 ;
  assign n50300 = ~n50286 & ~n50288 ;
  assign n50301 = \P2_buf2_reg[4]/NET0131  & n50300 ;
  assign n50302 = ~n50299 & ~n50301 ;
  assign n50303 = ~n50291 & n50302 ;
  assign n50304 = ~n50295 & n50303 ;
  assign n50307 = ~\P2_P3_InstQueueWr_Addr_reg[3]/NET0131  & n50011 ;
  assign n50313 = n27091 & n50307 ;
  assign n50312 = ~\P2_P3_InstQueue_reg[5][4]/NET0131  & ~n50307 ;
  assign n50314 = n27788 & ~n50312 ;
  assign n50315 = ~n50313 & n50314 ;
  assign n50305 = n27315 & n50268 ;
  assign n50306 = n36831 & ~n50305 ;
  assign n50308 = ~n50287 & ~n50307 ;
  assign n50309 = ~n50306 & n50308 ;
  assign n50310 = n50029 & ~n50309 ;
  assign n50311 = \P2_P3_InstQueue_reg[5][4]/NET0131  & ~n50310 ;
  assign n50316 = \P2_buf2_reg[28]/NET0131  & n50247 ;
  assign n50317 = \P2_buf2_reg[20]/NET0131  & n50267 ;
  assign n50318 = ~n50316 & ~n50317 ;
  assign n50319 = n27325 & ~n50318 ;
  assign n50320 = ~n50306 & ~n50308 ;
  assign n50321 = \P2_buf2_reg[4]/NET0131  & n50320 ;
  assign n50322 = ~n50319 & ~n50321 ;
  assign n50323 = ~n50311 & n50322 ;
  assign n50324 = ~n50315 & n50323 ;
  assign n50327 = ~\P2_P3_InstQueueWr_Addr_reg[3]/NET0131  & n50014 ;
  assign n50333 = n27091 & n50327 ;
  assign n50332 = ~\P2_P3_InstQueue_reg[6][4]/NET0131  & ~n50327 ;
  assign n50334 = n27788 & ~n50332 ;
  assign n50335 = ~n50333 & n50334 ;
  assign n50325 = n27315 & n50288 ;
  assign n50326 = n36831 & ~n50325 ;
  assign n50328 = ~n50307 & ~n50327 ;
  assign n50329 = ~n50326 & n50328 ;
  assign n50330 = n50029 & ~n50329 ;
  assign n50331 = \P2_P3_InstQueue_reg[6][4]/NET0131  & ~n50330 ;
  assign n50336 = \P2_buf2_reg[28]/NET0131  & n50267 ;
  assign n50337 = \P2_buf2_reg[20]/NET0131  & n50287 ;
  assign n50338 = ~n50336 & ~n50337 ;
  assign n50339 = n27325 & ~n50338 ;
  assign n50340 = ~n50326 & ~n50328 ;
  assign n50341 = \P2_buf2_reg[4]/NET0131  & n50340 ;
  assign n50342 = ~n50339 & ~n50341 ;
  assign n50343 = ~n50331 & n50342 ;
  assign n50344 = ~n50335 & n50343 ;
  assign n50352 = n27091 & n50046 ;
  assign n50351 = ~\P2_P3_InstQueue_reg[7][4]/NET0131  & ~n50046 ;
  assign n50353 = n27788 & ~n50351 ;
  assign n50354 = ~n50352 & n50353 ;
  assign n50345 = n27315 & n50308 ;
  assign n50346 = n36831 & ~n50345 ;
  assign n50347 = ~n50046 & ~n50327 ;
  assign n50348 = ~n50346 & n50347 ;
  assign n50349 = n50029 & ~n50348 ;
  assign n50350 = \P2_P3_InstQueue_reg[7][4]/NET0131  & ~n50349 ;
  assign n50355 = \P2_buf2_reg[28]/NET0131  & n50287 ;
  assign n50356 = \P2_buf2_reg[20]/NET0131  & n50307 ;
  assign n50357 = ~n50355 & ~n50356 ;
  assign n50358 = n27325 & ~n50357 ;
  assign n50359 = ~n50346 & ~n50347 ;
  assign n50360 = \P2_buf2_reg[4]/NET0131  & n50359 ;
  assign n50361 = ~n50358 & ~n50360 ;
  assign n50362 = ~n50350 & n50361 ;
  assign n50363 = ~n50354 & n50362 ;
  assign n50370 = n27091 & n50045 ;
  assign n50369 = ~\P2_P3_InstQueue_reg[8][4]/NET0131  & ~n50045 ;
  assign n50371 = n27788 & ~n50369 ;
  assign n50372 = ~n50370 & n50371 ;
  assign n50364 = n27315 & n50328 ;
  assign n50365 = n36831 & ~n50364 ;
  assign n50366 = n50047 & ~n50365 ;
  assign n50367 = n50029 & ~n50366 ;
  assign n50368 = \P2_P3_InstQueue_reg[8][4]/NET0131  & ~n50367 ;
  assign n50373 = \P2_buf2_reg[28]/NET0131  & n50307 ;
  assign n50374 = \P2_buf2_reg[20]/NET0131  & n50327 ;
  assign n50375 = ~n50373 & ~n50374 ;
  assign n50376 = n27325 & ~n50375 ;
  assign n50377 = ~n50047 & ~n50365 ;
  assign n50378 = \P2_buf2_reg[4]/NET0131  & n50377 ;
  assign n50379 = ~n50376 & ~n50378 ;
  assign n50380 = ~n50368 & n50379 ;
  assign n50381 = ~n50372 & n50380 ;
  assign n50388 = n27091 & n50053 ;
  assign n50387 = ~\P2_P3_InstQueue_reg[9][4]/NET0131  & ~n50053 ;
  assign n50389 = n27788 & ~n50387 ;
  assign n50390 = ~n50388 & n50389 ;
  assign n50382 = n27315 & n50347 ;
  assign n50383 = n36831 & ~n50382 ;
  assign n50384 = n50090 & ~n50383 ;
  assign n50385 = n50029 & ~n50384 ;
  assign n50386 = \P2_P3_InstQueue_reg[9][4]/NET0131  & ~n50385 ;
  assign n50391 = \P2_buf2_reg[28]/NET0131  & n50327 ;
  assign n50392 = \P2_buf2_reg[20]/NET0131  & n50046 ;
  assign n50393 = ~n50391 & ~n50392 ;
  assign n50394 = n27325 & ~n50393 ;
  assign n50395 = ~n50090 & ~n50383 ;
  assign n50396 = \P2_buf2_reg[4]/NET0131  & n50395 ;
  assign n50397 = ~n50394 & ~n50396 ;
  assign n50398 = ~n50386 & n50397 ;
  assign n50399 = ~n50390 & n50398 ;
  assign n50402 = \P2_P1_PhyAddrPointer_reg[0]/NET0131  & n36672 ;
  assign n50403 = \P2_P1_PhyAddrPointer_reg[1]/NET0131  & ~n50402 ;
  assign n50404 = ~\P2_P1_PhyAddrPointer_reg[1]/NET0131  & n50402 ;
  assign n50405 = ~n50403 & ~n50404 ;
  assign n50406 = ~\P2_P1_DataWidth_reg[1]/NET0131  & ~n50405 ;
  assign n50401 = \P2_P1_DataWidth_reg[1]/NET0131  & ~\P2_P1_rEIP_reg[1]/NET0131  ;
  assign n50407 = n11609 & ~n50401 ;
  assign n50408 = ~n50406 & n50407 ;
  assign n50414 = ~n21081 & ~n26088 ;
  assign n50415 = \P2_P1_rEIP_reg[1]/NET0131  & ~n50414 ;
  assign n50423 = ~\P2_P1_EBX_reg[0]/NET0131  & ~\P2_P1_EBX_reg[1]/NET0131  ;
  assign n50424 = ~n46230 & ~n50423 ;
  assign n50425 = \P2_P1_EBX_reg[31]/NET0131  & ~n50424 ;
  assign n50421 = ~\P2_P1_EBX_reg[1]/NET0131  & ~\P2_P1_EBX_reg[31]/NET0131  ;
  assign n50422 = ~\P2_P1_DataWidth_reg[1]/NET0131  & ~n21073 ;
  assign n50426 = ~n50421 & ~n50422 ;
  assign n50427 = ~n50425 & n50426 ;
  assign n50417 = ~\P2_P1_DataWidth_reg[1]/NET0131  & ~\P2_P1_rEIP_reg[1]/NET0131  ;
  assign n50428 = ~n21073 & n50417 ;
  assign n50429 = ~n50427 & ~n50428 ;
  assign n50430 = n24901 & ~n50429 ;
  assign n50413 = n21087 & n26070 ;
  assign n50416 = \P2_P1_EBX_reg[1]/NET0131  & ~n26103 ;
  assign n50418 = n25959 & n50417 ;
  assign n50419 = ~n50416 & ~n50418 ;
  assign n50420 = n24899 & ~n50419 ;
  assign n50431 = ~n50413 & ~n50420 ;
  assign n50432 = ~n50430 & n50431 ;
  assign n50433 = ~n50415 & n50432 ;
  assign n50434 = n11623 & ~n50433 ;
  assign n50400 = \P2_P1_PhyAddrPointer_reg[1]/NET0131  & n11625 ;
  assign n50409 = ~n11621 & ~n21098 ;
  assign n50410 = ~n11613 & ~n11692 ;
  assign n50411 = n50409 & n50410 ;
  assign n50412 = \P2_P1_rEIP_reg[1]/NET0131  & ~n50411 ;
  assign n50435 = ~n50400 & ~n50412 ;
  assign n50436 = ~n50434 & n50435 ;
  assign n50437 = ~n50408 & n50436 ;
  assign n50439 = \P1_P2_PhyAddrPointer_reg[0]/NET0131  & ~n36628 ;
  assign n50440 = \P1_P2_PhyAddrPointer_reg[1]/NET0131  & ~n50439 ;
  assign n50441 = ~\P1_P2_PhyAddrPointer_reg[1]/NET0131  & \P1_P2_PhyAddrPointer_reg[31]/NET0131  ;
  assign n50442 = \P1_P2_PhyAddrPointer_reg[0]/NET0131  & n50441 ;
  assign n50443 = ~n50440 & ~n50442 ;
  assign n50444 = ~\P1_P2_DataWidth_reg[1]/NET0131  & ~n50443 ;
  assign n50445 = \P1_P2_DataWidth_reg[1]/NET0131  & ~\P1_P2_rEIP_reg[1]/NET0131  ;
  assign n50446 = n25928 & ~n50445 ;
  assign n50447 = ~n50444 & n50446 ;
  assign n50449 = \P1_P2_rEIP_reg[1]/NET0131  & ~n48371 ;
  assign n50457 = ~n46698 & ~n48407 ;
  assign n50458 = \P1_P2_EBX_reg[31]/NET0131  & ~n50457 ;
  assign n50456 = ~\P1_P2_EBX_reg[1]/NET0131  & ~\P1_P2_EBX_reg[31]/NET0131  ;
  assign n50459 = ~n48373 & ~n50456 ;
  assign n50460 = ~n50458 & n50459 ;
  assign n50452 = ~\P1_P2_DataWidth_reg[1]/NET0131  & ~\P1_P2_rEIP_reg[1]/NET0131  ;
  assign n50461 = ~n25415 & n50452 ;
  assign n50462 = ~n50460 & ~n50461 ;
  assign n50463 = n25776 & ~n50462 ;
  assign n50450 = n25761 & ~n25885 ;
  assign n50451 = \P1_P2_EBX_reg[1]/NET0131  & ~n48443 ;
  assign n50453 = n25769 & n50452 ;
  assign n50454 = ~n50451 & ~n50453 ;
  assign n50455 = n25757 & ~n50454 ;
  assign n50464 = ~n50450 & ~n50455 ;
  assign n50465 = ~n50463 & n50464 ;
  assign n50466 = ~n25770 & ~n50465 ;
  assign n50467 = ~n50449 & ~n50466 ;
  assign n50468 = n25918 & ~n50467 ;
  assign n50438 = \P1_P2_PhyAddrPointer_reg[1]/NET0131  & n27675 ;
  assign n50448 = \P1_P2_rEIP_reg[1]/NET0131  & ~n48452 ;
  assign n50469 = ~n50438 & ~n50448 ;
  assign n50470 = ~n50468 & n50469 ;
  assign n50471 = ~n50447 & n50470 ;
  assign n50474 = ~\P2_P1_PhyAddrPointer_reg[1]/NET0131  & ~\P2_P1_PhyAddrPointer_reg[2]/NET0131  ;
  assign n50475 = ~n47407 & ~n50474 ;
  assign n50476 = ~\P2_P1_PhyAddrPointer_reg[0]/NET0131  & \P2_P1_PhyAddrPointer_reg[1]/NET0131  ;
  assign n50477 = n36672 & ~n50476 ;
  assign n50478 = ~n50475 & ~n50477 ;
  assign n50479 = n36672 & ~n50478 ;
  assign n50481 = ~n47852 & n50479 ;
  assign n50480 = n47852 & ~n50479 ;
  assign n50482 = ~\P2_P1_DataWidth_reg[1]/NET0131  & ~n50480 ;
  assign n50483 = ~n50481 & n50482 ;
  assign n50473 = \P2_P1_DataWidth_reg[1]/NET0131  & ~\P2_P1_rEIP_reg[3]/NET0131  ;
  assign n50484 = n11609 & ~n50473 ;
  assign n50485 = ~n50483 & n50484 ;
  assign n50486 = \P2_P1_rEIP_reg[3]/NET0131  & ~n50414 ;
  assign n50502 = \P2_P1_EBX_reg[3]/NET0131  & ~n26103 ;
  assign n50494 = \P2_P1_rEIP_reg[1]/NET0131  & \P2_P1_rEIP_reg[2]/NET0131  ;
  assign n50496 = ~\P2_P1_rEIP_reg[3]/NET0131  & ~n50494 ;
  assign n50495 = \P2_P1_rEIP_reg[3]/NET0131  & n50494 ;
  assign n50497 = ~\P2_P1_DataWidth_reg[1]/NET0131  & ~n50495 ;
  assign n50498 = ~n50496 & n50497 ;
  assign n50503 = n25959 & n50498 ;
  assign n50504 = ~n50502 & ~n50503 ;
  assign n50505 = n24898 & ~n50504 ;
  assign n50487 = n21067 & ~n25968 ;
  assign n50488 = ~\P2_P1_EBX_reg[2]/NET0131  & n50423 ;
  assign n50489 = \P2_P1_EBX_reg[31]/NET0131  & ~n50488 ;
  assign n50491 = \P2_P1_EBX_reg[3]/NET0131  & n50489 ;
  assign n50490 = ~\P2_P1_EBX_reg[3]/NET0131  & ~n50489 ;
  assign n50492 = ~n50422 & ~n50490 ;
  assign n50493 = ~n50491 & n50492 ;
  assign n50499 = ~n21073 & n50498 ;
  assign n50500 = ~n50493 & ~n50499 ;
  assign n50501 = n21062 & ~n50500 ;
  assign n50506 = ~n50487 & ~n50501 ;
  assign n50507 = ~n50505 & n50506 ;
  assign n50508 = ~n21081 & ~n50507 ;
  assign n50509 = ~n50486 & ~n50508 ;
  assign n50510 = n11623 & ~n50509 ;
  assign n50472 = \P2_P1_rEIP_reg[3]/NET0131  & ~n50411 ;
  assign n50511 = ~n47854 & ~n50472 ;
  assign n50512 = ~n50510 & n50511 ;
  assign n50513 = ~n50485 & n50512 ;
  assign n50516 = ~\P1_P2_PhyAddrPointer_reg[0]/NET0131  & n47384 ;
  assign n50517 = ~n36628 & ~n50516 ;
  assign n50519 = n47791 & ~n50517 ;
  assign n50518 = ~n47791 & n50517 ;
  assign n50520 = ~\P1_P2_DataWidth_reg[1]/NET0131  & ~n50518 ;
  assign n50521 = ~n50519 & n50520 ;
  assign n50515 = \P1_P2_DataWidth_reg[1]/NET0131  & ~\P1_P2_rEIP_reg[3]/NET0131  ;
  assign n50522 = n25928 & ~n50515 ;
  assign n50523 = ~n50521 & n50522 ;
  assign n50524 = \P1_P2_rEIP_reg[3]/NET0131  & ~n48371 ;
  assign n50533 = \P1_P2_EBX_reg[31]/NET0131  & ~n48408 ;
  assign n50535 = \P1_P2_EBX_reg[3]/NET0131  & n50533 ;
  assign n50534 = ~\P1_P2_EBX_reg[3]/NET0131  & ~n50533 ;
  assign n50536 = ~n48373 & ~n50534 ;
  assign n50537 = ~n50535 & n50536 ;
  assign n50527 = ~\P1_P2_rEIP_reg[3]/NET0131  & ~n48380 ;
  assign n50528 = ~\P1_P2_DataWidth_reg[1]/NET0131  & ~n48381 ;
  assign n50529 = ~n50527 & n50528 ;
  assign n50538 = ~n25415 & n50529 ;
  assign n50539 = ~n50537 & ~n50538 ;
  assign n50540 = n25776 & ~n50539 ;
  assign n50525 = n25761 & ~n25858 ;
  assign n50526 = \P1_P2_EBX_reg[3]/NET0131  & ~n48443 ;
  assign n50530 = n25769 & n50529 ;
  assign n50531 = ~n50526 & ~n50530 ;
  assign n50532 = n25757 & ~n50531 ;
  assign n50541 = ~n50525 & ~n50532 ;
  assign n50542 = ~n50540 & n50541 ;
  assign n50543 = ~n25770 & ~n50542 ;
  assign n50544 = ~n50524 & ~n50543 ;
  assign n50545 = n25918 & ~n50544 ;
  assign n50514 = \P1_P2_PhyAddrPointer_reg[3]/NET0131  & n27675 ;
  assign n50546 = \P1_P2_rEIP_reg[3]/NET0131  & ~n48452 ;
  assign n50547 = ~n50514 & ~n50546 ;
  assign n50548 = ~n50545 & n50547 ;
  assign n50549 = ~n50523 & n50548 ;
  assign n50552 = \P1_P1_PhyAddrPointer_reg[0]/NET0131  & ~n36733 ;
  assign n50554 = \P1_P1_PhyAddrPointer_reg[1]/NET0131  & n50552 ;
  assign n50553 = ~\P1_P1_PhyAddrPointer_reg[1]/NET0131  & ~n50552 ;
  assign n50555 = ~\P1_P1_DataWidth_reg[1]/NET0131  & ~n50553 ;
  assign n50556 = ~n50554 & n50555 ;
  assign n50551 = \P1_P1_DataWidth_reg[1]/NET0131  & ~\P1_P1_rEIP_reg[1]/NET0131  ;
  assign n50557 = n8282 & ~n50551 ;
  assign n50558 = ~n50556 & n50557 ;
  assign n50559 = ~n15364 & ~n26131 ;
  assign n50560 = \P1_P1_rEIP_reg[1]/NET0131  & ~n50559 ;
  assign n50572 = \P1_P1_EBX_reg[1]/NET0131  & ~n26275 ;
  assign n50568 = ~\P1_P1_DataWidth_reg[1]/NET0131  & ~\P1_P1_rEIP_reg[1]/NET0131  ;
  assign n50573 = n26264 & n50568 ;
  assign n50574 = ~n50572 & ~n50573 ;
  assign n50575 = n24502 & ~n50574 ;
  assign n50561 = n15382 & n26191 ;
  assign n50562 = ~\P1_P1_EBX_reg[0]/NET0131  & ~\P1_P1_EBX_reg[1]/NET0131  ;
  assign n50563 = ~n46537 & ~n50562 ;
  assign n50564 = \P1_P1_EBX_reg[31]/NET0131  & ~n50563 ;
  assign n50565 = ~\P1_P1_EBX_reg[1]/NET0131  & ~\P1_P1_EBX_reg[31]/NET0131  ;
  assign n50566 = ~n26274 & ~n50565 ;
  assign n50567 = ~n50564 & n50566 ;
  assign n50569 = ~n15335 & n50568 ;
  assign n50570 = ~n50567 & ~n50569 ;
  assign n50571 = n15334 & ~n50570 ;
  assign n50576 = ~n50561 & ~n50571 ;
  assign n50577 = ~n50575 & n50576 ;
  assign n50578 = ~n15364 & ~n50577 ;
  assign n50579 = ~n50560 & ~n50578 ;
  assign n50580 = n8355 & ~n50579 ;
  assign n50550 = \P1_P1_PhyAddrPointer_reg[1]/NET0131  & n8361 ;
  assign n50581 = ~n8353 & ~n15324 ;
  assign n50582 = ~n8287 & ~n8350 ;
  assign n50583 = n50581 & n50582 ;
  assign n50584 = \P1_P1_rEIP_reg[1]/NET0131  & ~n50583 ;
  assign n50585 = ~n50550 & ~n50584 ;
  assign n50586 = ~n50580 & n50585 ;
  assign n50587 = ~n50558 & n50586 ;
  assign n50590 = ~\P1_P1_PhyAddrPointer_reg[0]/NET0131  & n47430 ;
  assign n50591 = ~n36733 & ~n50590 ;
  assign n50593 = ~n47912 & n50591 ;
  assign n50592 = n47912 & ~n50591 ;
  assign n50594 = ~\P1_P1_DataWidth_reg[1]/NET0131  & ~n50592 ;
  assign n50595 = ~n50593 & n50594 ;
  assign n50589 = \P1_P1_DataWidth_reg[1]/NET0131  & ~\P1_P1_rEIP_reg[3]/NET0131  ;
  assign n50596 = n8282 & ~n50589 ;
  assign n50597 = ~n50595 & n50596 ;
  assign n50598 = \P1_P1_rEIP_reg[3]/NET0131  & ~n50559 ;
  assign n50609 = ~\P1_P1_EBX_reg[2]/NET0131  & n50562 ;
  assign n50610 = \P1_P1_EBX_reg[31]/NET0131  & ~n50609 ;
  assign n50612 = \P1_P1_EBX_reg[3]/NET0131  & n50610 ;
  assign n50611 = ~\P1_P1_EBX_reg[3]/NET0131  & ~n50610 ;
  assign n50613 = ~n26274 & ~n50611 ;
  assign n50614 = ~n50612 & n50613 ;
  assign n50600 = \P1_P1_rEIP_reg[1]/NET0131  & \P1_P1_rEIP_reg[2]/NET0131  ;
  assign n50602 = ~\P1_P1_rEIP_reg[3]/NET0131  & ~n50600 ;
  assign n50601 = \P1_P1_rEIP_reg[3]/NET0131  & n50600 ;
  assign n50603 = ~\P1_P1_DataWidth_reg[1]/NET0131  & ~n50601 ;
  assign n50604 = ~n50602 & n50603 ;
  assign n50615 = ~n15335 & n50604 ;
  assign n50616 = ~n50614 & ~n50615 ;
  assign n50617 = n15334 & ~n50616 ;
  assign n50599 = \P1_P1_EBX_reg[3]/NET0131  & ~n26275 ;
  assign n50605 = n26264 & n50604 ;
  assign n50606 = ~n50599 & ~n50605 ;
  assign n50607 = n24502 & ~n50606 ;
  assign n50608 = n15382 & ~n26238 ;
  assign n50618 = ~n50607 & ~n50608 ;
  assign n50619 = ~n50617 & n50618 ;
  assign n50620 = ~n15364 & ~n50619 ;
  assign n50621 = ~n50598 & ~n50620 ;
  assign n50622 = n8355 & ~n50621 ;
  assign n50588 = \P1_P1_rEIP_reg[3]/NET0131  & ~n50583 ;
  assign n50623 = ~n47914 & ~n50588 ;
  assign n50624 = ~n50622 & n50623 ;
  assign n50625 = ~n50597 & n50624 ;
  assign n50628 = \P2_P2_PhyAddrPointer_reg[0]/NET0131  & n36792 ;
  assign n50630 = \P2_P2_PhyAddrPointer_reg[1]/NET0131  & n50628 ;
  assign n50629 = ~\P2_P2_PhyAddrPointer_reg[1]/NET0131  & ~n50628 ;
  assign n50631 = ~\P2_P2_DataWidth_reg[1]/NET0131  & ~n50629 ;
  assign n50632 = ~n50630 & n50631 ;
  assign n50627 = \P2_P2_DataWidth_reg[1]/NET0131  & ~\P2_P2_rEIP_reg[1]/NET0131  ;
  assign n50633 = n26794 & ~n50627 ;
  assign n50634 = ~n50632 & n50633 ;
  assign n50640 = ~n26640 & ~n26680 ;
  assign n50641 = \P2_P2_rEIP_reg[1]/NET0131  & ~n50640 ;
  assign n50650 = ~\P2_P2_EBX_reg[0]/NET0131  & ~\P2_P2_EBX_reg[1]/NET0131  ;
  assign n50651 = ~n46420 & ~n50650 ;
  assign n50652 = \P2_P2_EBX_reg[31]/NET0131  & ~n50651 ;
  assign n50648 = ~\P2_P2_EBX_reg[1]/NET0131  & ~\P2_P2_EBX_reg[31]/NET0131  ;
  assign n50649 = ~\P2_P2_DataWidth_reg[1]/NET0131  & ~n26286 ;
  assign n50653 = ~n50648 & ~n50649 ;
  assign n50654 = ~n50652 & n50653 ;
  assign n50644 = ~\P2_P2_DataWidth_reg[1]/NET0131  & ~\P2_P2_rEIP_reg[1]/NET0131  ;
  assign n50655 = ~n26286 & n50644 ;
  assign n50656 = ~n50654 & ~n50655 ;
  assign n50657 = n47684 & ~n50656 ;
  assign n50638 = n26637 & ~n26640 ;
  assign n50639 = n26756 & n50638 ;
  assign n50642 = ~\P2_P2_DataWidth_reg[1]/NET0131  & n26651 ;
  assign n50643 = \P2_P2_EBX_reg[1]/NET0131  & ~n50642 ;
  assign n50645 = n26651 & n50644 ;
  assign n50646 = ~n50643 & ~n50645 ;
  assign n50647 = n26786 & ~n50646 ;
  assign n50658 = ~n50639 & ~n50647 ;
  assign n50659 = ~n50657 & n50658 ;
  assign n50660 = ~n50641 & n50659 ;
  assign n50661 = n26792 & ~n50660 ;
  assign n50626 = \P2_P2_PhyAddrPointer_reg[1]/NET0131  & n27637 ;
  assign n50635 = ~n27613 & ~n27977 ;
  assign n50636 = n36757 & n50635 ;
  assign n50637 = \P2_P2_rEIP_reg[1]/NET0131  & ~n50636 ;
  assign n50662 = ~n50626 & ~n50637 ;
  assign n50663 = ~n50661 & n50662 ;
  assign n50664 = ~n50634 & n50663 ;
  assign n50667 = ~\P2_P2_PhyAddrPointer_reg[0]/NET0131  & n47451 ;
  assign n50668 = n36792 & ~n50667 ;
  assign n50670 = n47965 & ~n50668 ;
  assign n50669 = ~n47965 & n50668 ;
  assign n50671 = ~\P2_P2_DataWidth_reg[1]/NET0131  & ~n50669 ;
  assign n50672 = ~n50670 & n50671 ;
  assign n50666 = \P2_P2_DataWidth_reg[1]/NET0131  & ~\P2_P2_rEIP_reg[3]/NET0131  ;
  assign n50673 = n26794 & ~n50666 ;
  assign n50674 = ~n50672 & n50673 ;
  assign n50677 = \P2_P2_rEIP_reg[3]/NET0131  & ~n50640 ;
  assign n50678 = ~\P2_P2_EBX_reg[2]/NET0131  & n50650 ;
  assign n50679 = \P2_P2_EBX_reg[31]/NET0131  & ~n50678 ;
  assign n50681 = \P2_P2_EBX_reg[3]/NET0131  & n50679 ;
  assign n50680 = ~\P2_P2_EBX_reg[3]/NET0131  & ~n50679 ;
  assign n50682 = ~n50649 & ~n50680 ;
  assign n50683 = ~n50681 & n50682 ;
  assign n50684 = \P2_P2_rEIP_reg[1]/NET0131  & \P2_P2_rEIP_reg[2]/NET0131  ;
  assign n50686 = ~\P2_P2_rEIP_reg[3]/NET0131  & ~n50684 ;
  assign n50685 = \P2_P2_rEIP_reg[3]/NET0131  & n50684 ;
  assign n50687 = ~\P2_P2_DataWidth_reg[1]/NET0131  & ~n50685 ;
  assign n50688 = ~n50686 & n50687 ;
  assign n50689 = ~n26286 & n50688 ;
  assign n50690 = ~n50683 & ~n50689 ;
  assign n50691 = n47684 & ~n50690 ;
  assign n50676 = ~n26721 & n50638 ;
  assign n50692 = \P2_P2_EBX_reg[3]/NET0131  & ~n50642 ;
  assign n50693 = n26651 & n50688 ;
  assign n50694 = ~n50692 & ~n50693 ;
  assign n50695 = n26786 & ~n50694 ;
  assign n50696 = ~n50676 & ~n50695 ;
  assign n50697 = ~n50691 & n50696 ;
  assign n50698 = ~n50677 & n50697 ;
  assign n50699 = n26792 & ~n50698 ;
  assign n50665 = \P2_P2_rEIP_reg[3]/NET0131  & ~n50636 ;
  assign n50675 = \P2_P2_PhyAddrPointer_reg[3]/NET0131  & n27637 ;
  assign n50700 = ~n50665 & ~n50675 ;
  assign n50701 = ~n50699 & n50700 ;
  assign n50702 = ~n50674 & n50701 ;
  assign n50706 = ~\P2_P3_PhyAddrPointer_reg[1]/NET0131  & ~\P2_P3_PhyAddrPointer_reg[2]/NET0131  ;
  assign n50707 = ~n47477 & ~n50706 ;
  assign n50708 = ~\P2_P3_PhyAddrPointer_reg[0]/NET0131  & \P2_P3_PhyAddrPointer_reg[1]/NET0131  ;
  assign n50709 = ~n36863 & ~n50708 ;
  assign n50710 = ~n50707 & ~n50709 ;
  assign n50711 = ~n36863 & ~n50710 ;
  assign n50713 = ~n48087 & n50711 ;
  assign n50712 = n48087 & ~n50711 ;
  assign n50714 = ~\P2_P3_DataWidth_reg[1]/NET0131  & ~n50712 ;
  assign n50715 = ~n50713 & n50714 ;
  assign n50705 = \P2_P3_DataWidth_reg[1]/NET0131  & ~\P2_P3_rEIP_reg[3]/NET0131  ;
  assign n50716 = n27315 & ~n50705 ;
  assign n50717 = ~n50715 & n50716 ;
  assign n50718 = \P2_P3_rEIP_reg[3]/NET0131  & ~n27277 ;
  assign n50720 = ~\P2_P3_EBX_reg[0]/NET0131  & ~\P2_P3_EBX_reg[1]/NET0131  ;
  assign n50721 = ~\P2_P3_EBX_reg[2]/NET0131  & n50720 ;
  assign n50722 = \P2_P3_EBX_reg[31]/NET0131  & ~n50721 ;
  assign n50723 = \P2_P3_EBX_reg[3]/NET0131  & n50722 ;
  assign n50724 = ~\P2_P3_EBX_reg[3]/NET0131  & ~n50722 ;
  assign n50725 = ~n50723 & ~n50724 ;
  assign n50726 = ~n27302 & n50725 ;
  assign n50727 = \P2_P3_rEIP_reg[1]/NET0131  & \P2_P3_rEIP_reg[2]/NET0131  ;
  assign n50729 = ~\P2_P3_rEIP_reg[3]/NET0131  & ~n50727 ;
  assign n50728 = \P2_P3_rEIP_reg[3]/NET0131  & n50727 ;
  assign n50730 = ~\P2_P3_DataWidth_reg[1]/NET0131  & ~n50728 ;
  assign n50731 = ~n50729 & n50730 ;
  assign n50732 = ~n27192 & n50731 ;
  assign n50733 = ~n50726 & ~n50732 ;
  assign n50734 = n27122 & ~n50733 ;
  assign n50719 = ~n27060 & n27124 ;
  assign n50735 = ~n27148 & n27302 ;
  assign n50736 = \P2_P3_EBX_reg[3]/NET0131  & ~n50735 ;
  assign n50737 = ~n27148 & ~n27192 ;
  assign n50738 = n50731 & n50737 ;
  assign n50739 = ~n50736 & ~n50738 ;
  assign n50740 = n27121 & ~n50739 ;
  assign n50741 = ~n50719 & ~n50740 ;
  assign n50742 = ~n50734 & n50741 ;
  assign n50743 = ~n27177 & ~n50742 ;
  assign n50744 = ~n50718 & ~n50743 ;
  assign n50745 = n27308 & ~n50744 ;
  assign n50703 = ~n32867 & n48084 ;
  assign n50704 = \P2_P3_rEIP_reg[3]/NET0131  & ~n50703 ;
  assign n50746 = ~n48089 & ~n50704 ;
  assign n50747 = ~n50745 & n50746 ;
  assign n50748 = ~n50717 & n50747 ;
  assign n50751 = ~\P2_P1_PhyAddrPointer_reg[0]/NET0131  & n39457 ;
  assign n50752 = \P2_P1_PhyAddrPointer_reg[14]/NET0131  & n50751 ;
  assign n50753 = \P2_P1_PhyAddrPointer_reg[15]/NET0131  & n50752 ;
  assign n50754 = n36656 & n50753 ;
  assign n50755 = n36672 & ~n50754 ;
  assign n50757 = ~n41578 & n50755 ;
  assign n50756 = n41578 & ~n50755 ;
  assign n50758 = ~\P2_P1_DataWidth_reg[1]/NET0131  & ~n50756 ;
  assign n50759 = ~n50757 & n50758 ;
  assign n50750 = \P2_P1_DataWidth_reg[1]/NET0131  & ~\P2_P1_rEIP_reg[20]/NET0131  ;
  assign n50760 = n11609 & ~n50750 ;
  assign n50761 = ~n50759 & n50760 ;
  assign n50762 = \P2_P1_rEIP_reg[20]/NET0131  & ~n50414 ;
  assign n50784 = ~\P2_P1_EBX_reg[20]/NET0131  & ~n26103 ;
  assign n50785 = n24898 & ~n50784 ;
  assign n50789 = ~\P2_P1_EBX_reg[3]/NET0131  & n50488 ;
  assign n50790 = ~\P2_P1_EBX_reg[4]/NET0131  & n50789 ;
  assign n50791 = ~\P2_P1_EBX_reg[5]/NET0131  & n50790 ;
  assign n50792 = ~\P2_P1_EBX_reg[6]/NET0131  & n50791 ;
  assign n50793 = ~\P2_P1_EBX_reg[7]/NET0131  & n50792 ;
  assign n50794 = ~\P2_P1_EBX_reg[8]/NET0131  & n50793 ;
  assign n50795 = ~\P2_P1_EBX_reg[9]/NET0131  & n50794 ;
  assign n50796 = ~\P2_P1_EBX_reg[10]/NET0131  & n50795 ;
  assign n50797 = ~\P2_P1_EBX_reg[11]/NET0131  & n50796 ;
  assign n50798 = ~\P2_P1_EBX_reg[12]/NET0131  & n50797 ;
  assign n50799 = ~\P2_P1_EBX_reg[13]/NET0131  & n50798 ;
  assign n50800 = ~\P2_P1_EBX_reg[14]/NET0131  & n50799 ;
  assign n50801 = ~\P2_P1_EBX_reg[15]/NET0131  & n50800 ;
  assign n50802 = ~\P2_P1_EBX_reg[16]/NET0131  & n50801 ;
  assign n50803 = ~\P2_P1_EBX_reg[17]/NET0131  & n50802 ;
  assign n50804 = ~\P2_P1_EBX_reg[18]/NET0131  & n50803 ;
  assign n50805 = ~\P2_P1_EBX_reg[19]/NET0131  & n50804 ;
  assign n50806 = \P2_P1_EBX_reg[31]/NET0131  & ~n50805 ;
  assign n50808 = ~\P2_P1_EBX_reg[20]/NET0131  & n50806 ;
  assign n50807 = \P2_P1_EBX_reg[20]/NET0131  & ~n50806 ;
  assign n50809 = ~n50422 & ~n50807 ;
  assign n50810 = ~n50808 & n50809 ;
  assign n50811 = n21062 & ~n50810 ;
  assign n50812 = ~n50785 & ~n50811 ;
  assign n50763 = \P2_P1_rEIP_reg[15]/NET0131  & \P2_P1_rEIP_reg[16]/NET0131  ;
  assign n50764 = \P2_P1_rEIP_reg[17]/NET0131  & n50763 ;
  assign n50765 = \P2_P1_rEIP_reg[12]/NET0131  & \P2_P1_rEIP_reg[13]/NET0131  ;
  assign n50766 = \P2_P1_rEIP_reg[4]/NET0131  & n50495 ;
  assign n50767 = \P2_P1_rEIP_reg[5]/NET0131  & n50766 ;
  assign n50768 = \P2_P1_rEIP_reg[6]/NET0131  & n50767 ;
  assign n50769 = \P2_P1_rEIP_reg[7]/NET0131  & n50768 ;
  assign n50770 = \P2_P1_rEIP_reg[8]/NET0131  & n50769 ;
  assign n50771 = \P2_P1_rEIP_reg[9]/NET0131  & n50770 ;
  assign n50772 = \P2_P1_rEIP_reg[10]/NET0131  & \P2_P1_rEIP_reg[11]/NET0131  ;
  assign n50773 = n50771 & n50772 ;
  assign n50774 = n50765 & n50773 ;
  assign n50775 = \P2_P1_rEIP_reg[14]/NET0131  & n50774 ;
  assign n50776 = n50764 & n50775 ;
  assign n50777 = \P2_P1_rEIP_reg[18]/NET0131  & n50776 ;
  assign n50778 = \P2_P1_rEIP_reg[19]/NET0131  & n50777 ;
  assign n50779 = ~\P2_P1_rEIP_reg[20]/NET0131  & ~n50778 ;
  assign n50780 = \P2_P1_rEIP_reg[18]/NET0131  & \P2_P1_rEIP_reg[19]/NET0131  ;
  assign n50781 = \P2_P1_rEIP_reg[20]/NET0131  & n50780 ;
  assign n50782 = n50776 & n50781 ;
  assign n50783 = ~n50779 & ~n50782 ;
  assign n50786 = n25958 & n50785 ;
  assign n50787 = n50422 & ~n50786 ;
  assign n50788 = ~n50783 & n50787 ;
  assign n50813 = ~n21081 & ~n50788 ;
  assign n50814 = ~n50812 & n50813 ;
  assign n50815 = ~n50762 & ~n50814 ;
  assign n50816 = n11623 & ~n50815 ;
  assign n50749 = \P2_P1_PhyAddrPointer_reg[20]/NET0131  & n11625 ;
  assign n50817 = \P2_P1_rEIP_reg[20]/NET0131  & ~n50411 ;
  assign n50818 = ~n50749 & ~n50817 ;
  assign n50819 = ~n50816 & n50818 ;
  assign n50820 = ~n50761 & n50819 ;
  assign n50823 = ~\P2_P1_PhyAddrPointer_reg[0]/NET0131  & n39455 ;
  assign n50824 = n39453 & n50823 ;
  assign n50825 = n36658 & n50824 ;
  assign n50826 = n36672 & ~n50825 ;
  assign n50828 = n43553 & ~n50826 ;
  assign n50827 = ~n43553 & n50826 ;
  assign n50829 = ~\P2_P1_DataWidth_reg[1]/NET0131  & ~n50827 ;
  assign n50830 = ~n50828 & n50829 ;
  assign n50822 = \P2_P1_DataWidth_reg[1]/NET0131  & ~\P2_P1_rEIP_reg[21]/NET0131  ;
  assign n50831 = n11609 & ~n50822 ;
  assign n50832 = ~n50830 & n50831 ;
  assign n50838 = ~\P2_P1_EBX_reg[20]/NET0131  & n50805 ;
  assign n50839 = \P2_P1_EBX_reg[31]/NET0131  & ~n50838 ;
  assign n50841 = ~\P2_P1_EBX_reg[21]/NET0131  & n50839 ;
  assign n50840 = \P2_P1_EBX_reg[21]/NET0131  & ~n50839 ;
  assign n50842 = ~n50422 & ~n50840 ;
  assign n50843 = ~n50841 & n50842 ;
  assign n50834 = ~\P2_P1_rEIP_reg[21]/NET0131  & ~n50782 ;
  assign n50835 = \P2_P1_rEIP_reg[21]/NET0131  & n50782 ;
  assign n50836 = ~n50834 & ~n50835 ;
  assign n50837 = n50422 & ~n50836 ;
  assign n50844 = n24901 & ~n50837 ;
  assign n50845 = ~n50843 & n50844 ;
  assign n50833 = \P2_P1_rEIP_reg[21]/NET0131  & ~n50414 ;
  assign n50847 = n26103 & ~n50836 ;
  assign n50846 = ~\P2_P1_EBX_reg[21]/NET0131  & ~n26103 ;
  assign n50848 = n24899 & ~n50846 ;
  assign n50849 = ~n50847 & n50848 ;
  assign n50850 = ~n50833 & ~n50849 ;
  assign n50851 = ~n50845 & n50850 ;
  assign n50852 = n11623 & ~n50851 ;
  assign n50821 = \P2_P1_PhyAddrPointer_reg[21]/NET0131  & n11625 ;
  assign n50853 = \P2_P1_rEIP_reg[21]/NET0131  & ~n50411 ;
  assign n50854 = ~n50821 & ~n50853 ;
  assign n50855 = ~n50852 & n50854 ;
  assign n50856 = ~n50832 & n50855 ;
  assign n50859 = n41550 & n50824 ;
  assign n50860 = n41595 & n50859 ;
  assign n50861 = n36672 & ~n50860 ;
  assign n50863 = ~n41597 & n50861 ;
  assign n50862 = n41597 & ~n50861 ;
  assign n50864 = ~\P2_P1_DataWidth_reg[1]/NET0131  & ~n50862 ;
  assign n50865 = ~n50863 & n50864 ;
  assign n50858 = \P2_P1_DataWidth_reg[1]/NET0131  & ~\P2_P1_rEIP_reg[22]/NET0131  ;
  assign n50866 = n11609 & ~n50858 ;
  assign n50867 = ~n50865 & n50866 ;
  assign n50873 = ~\P2_P1_EBX_reg[21]/NET0131  & n50838 ;
  assign n50874 = \P2_P1_EBX_reg[31]/NET0131  & ~n50873 ;
  assign n50876 = ~\P2_P1_EBX_reg[22]/NET0131  & n50874 ;
  assign n50875 = \P2_P1_EBX_reg[22]/NET0131  & ~n50874 ;
  assign n50877 = ~n50422 & ~n50875 ;
  assign n50878 = ~n50876 & n50877 ;
  assign n50869 = ~\P2_P1_rEIP_reg[22]/NET0131  & ~n50835 ;
  assign n50870 = \P2_P1_rEIP_reg[22]/NET0131  & n50835 ;
  assign n50871 = ~n50869 & ~n50870 ;
  assign n50872 = n50422 & ~n50871 ;
  assign n50879 = n24901 & ~n50872 ;
  assign n50880 = ~n50878 & n50879 ;
  assign n50868 = \P2_P1_rEIP_reg[22]/NET0131  & ~n50414 ;
  assign n50882 = n26103 & ~n50871 ;
  assign n50881 = ~\P2_P1_EBX_reg[22]/NET0131  & ~n26103 ;
  assign n50883 = n24899 & ~n50881 ;
  assign n50884 = ~n50882 & n50883 ;
  assign n50885 = ~n50868 & ~n50884 ;
  assign n50886 = ~n50880 & n50885 ;
  assign n50887 = n11623 & ~n50886 ;
  assign n50857 = \P2_P1_PhyAddrPointer_reg[22]/NET0131  & n11625 ;
  assign n50888 = \P2_P1_rEIP_reg[22]/NET0131  & ~n50411 ;
  assign n50889 = ~n50857 & ~n50888 ;
  assign n50890 = ~n50887 & n50889 ;
  assign n50891 = ~n50867 & n50890 ;
  assign n50915 = n39480 & n50859 ;
  assign n50916 = n36672 & ~n50915 ;
  assign n50918 = ~n39483 & n50916 ;
  assign n50917 = n39483 & ~n50916 ;
  assign n50919 = ~\P2_P1_DataWidth_reg[1]/NET0131  & ~n50917 ;
  assign n50920 = ~n50918 & n50919 ;
  assign n50914 = \P2_P1_DataWidth_reg[1]/NET0131  & ~\P2_P1_rEIP_reg[23]/NET0131  ;
  assign n50921 = n11609 & ~n50914 ;
  assign n50922 = ~n50920 & n50921 ;
  assign n50898 = ~\P2_P1_EBX_reg[22]/NET0131  & n50873 ;
  assign n50899 = \P2_P1_EBX_reg[31]/NET0131  & ~n50898 ;
  assign n50901 = ~\P2_P1_EBX_reg[23]/NET0131  & n50899 ;
  assign n50900 = \P2_P1_EBX_reg[23]/NET0131  & ~n50899 ;
  assign n50902 = ~n50422 & ~n50900 ;
  assign n50903 = ~n50901 & n50902 ;
  assign n50894 = ~\P2_P1_rEIP_reg[23]/NET0131  & ~n50870 ;
  assign n50895 = \P2_P1_rEIP_reg[23]/NET0131  & n50870 ;
  assign n50896 = ~n50894 & ~n50895 ;
  assign n50897 = n50422 & ~n50896 ;
  assign n50904 = n24901 & ~n50897 ;
  assign n50905 = ~n50903 & n50904 ;
  assign n50893 = \P2_P1_rEIP_reg[23]/NET0131  & ~n50414 ;
  assign n50907 = n26103 & ~n50896 ;
  assign n50906 = ~\P2_P1_EBX_reg[23]/NET0131  & ~n26103 ;
  assign n50908 = n24899 & ~n50906 ;
  assign n50909 = ~n50907 & n50908 ;
  assign n50910 = ~n50893 & ~n50909 ;
  assign n50911 = ~n50905 & n50910 ;
  assign n50912 = n11623 & ~n50911 ;
  assign n50892 = \P2_P1_PhyAddrPointer_reg[23]/NET0131  & n11625 ;
  assign n50913 = \P2_P1_rEIP_reg[23]/NET0131  & ~n50411 ;
  assign n50923 = ~n50892 & ~n50913 ;
  assign n50924 = ~n50912 & n50923 ;
  assign n50925 = ~n50922 & n50924 ;
  assign n50949 = n39482 & n50859 ;
  assign n50950 = n36672 & ~n50949 ;
  assign n50952 = n41613 & ~n50950 ;
  assign n50951 = ~n41613 & n50950 ;
  assign n50953 = ~\P2_P1_DataWidth_reg[1]/NET0131  & ~n50951 ;
  assign n50954 = ~n50952 & n50953 ;
  assign n50948 = \P2_P1_DataWidth_reg[1]/NET0131  & ~\P2_P1_rEIP_reg[24]/NET0131  ;
  assign n50955 = n11609 & ~n50948 ;
  assign n50956 = ~n50954 & n50955 ;
  assign n50933 = ~\P2_P1_EBX_reg[23]/NET0131  & n50898 ;
  assign n50934 = \P2_P1_EBX_reg[31]/NET0131  & ~n50933 ;
  assign n50936 = ~\P2_P1_EBX_reg[24]/NET0131  & n50934 ;
  assign n50935 = \P2_P1_EBX_reg[24]/NET0131  & ~n50934 ;
  assign n50937 = ~n50422 & ~n50935 ;
  assign n50938 = ~n50936 & n50937 ;
  assign n50929 = ~\P2_P1_rEIP_reg[24]/NET0131  & ~n50895 ;
  assign n50930 = \P2_P1_rEIP_reg[24]/NET0131  & n50895 ;
  assign n50931 = ~n50929 & ~n50930 ;
  assign n50932 = n50422 & ~n50931 ;
  assign n50939 = n24901 & ~n50932 ;
  assign n50940 = ~n50938 & n50939 ;
  assign n50928 = \P2_P1_rEIP_reg[24]/NET0131  & ~n50414 ;
  assign n50942 = n26103 & ~n50931 ;
  assign n50941 = ~\P2_P1_EBX_reg[24]/NET0131  & ~n26103 ;
  assign n50943 = n24899 & ~n50941 ;
  assign n50944 = ~n50942 & n50943 ;
  assign n50945 = ~n50928 & ~n50944 ;
  assign n50946 = ~n50940 & n50945 ;
  assign n50947 = n11623 & ~n50946 ;
  assign n50926 = \P2_P1_PhyAddrPointer_reg[24]/NET0131  & n11625 ;
  assign n50927 = \P2_P1_rEIP_reg[24]/NET0131  & ~n50411 ;
  assign n50957 = ~n50926 & ~n50927 ;
  assign n50958 = ~n50947 & n50957 ;
  assign n50959 = ~n50956 & n50958 ;
  assign n50983 = ~\P2_P1_EBX_reg[24]/NET0131  & n50933 ;
  assign n50984 = \P2_P1_EBX_reg[31]/NET0131  & ~n50983 ;
  assign n50986 = ~\P2_P1_EBX_reg[25]/NET0131  & n50984 ;
  assign n50985 = \P2_P1_EBX_reg[25]/NET0131  & ~n50984 ;
  assign n50987 = ~n50422 & ~n50985 ;
  assign n50988 = ~n50986 & n50987 ;
  assign n50977 = \P2_P1_rEIP_reg[25]/NET0131  & ~n50770 ;
  assign n50967 = \P2_P1_rEIP_reg[24]/NET0131  & \P2_P1_rEIP_reg[9]/NET0131  ;
  assign n50968 = n50772 & n50967 ;
  assign n50969 = n50764 & n50968 ;
  assign n50966 = \P2_P1_rEIP_reg[14]/NET0131  & n50765 ;
  assign n50964 = \P2_P1_rEIP_reg[21]/NET0131  & \P2_P1_rEIP_reg[22]/NET0131  ;
  assign n50965 = \P2_P1_rEIP_reg[23]/NET0131  & n50964 ;
  assign n50970 = n50781 & n50965 ;
  assign n50971 = n50966 & n50970 ;
  assign n50972 = n50969 & n50971 ;
  assign n50973 = \P2_P1_rEIP_reg[25]/NET0131  & ~n50972 ;
  assign n50974 = ~\P2_P1_rEIP_reg[25]/NET0131  & n50972 ;
  assign n50975 = ~n50973 & ~n50974 ;
  assign n50976 = n50770 & ~n50975 ;
  assign n50978 = n50422 & ~n50976 ;
  assign n50979 = ~n50977 & n50978 ;
  assign n50989 = n24901 & ~n50979 ;
  assign n50990 = ~n50988 & n50989 ;
  assign n50962 = \P2_P1_rEIP_reg[25]/NET0131  & ~n50414 ;
  assign n50963 = ~\P2_P1_EBX_reg[25]/NET0131  & ~n26103 ;
  assign n50980 = ~n25958 & n50979 ;
  assign n50981 = ~n50963 & ~n50980 ;
  assign n50982 = n24899 & n50981 ;
  assign n50991 = ~n50962 & ~n50982 ;
  assign n50992 = ~n50990 & n50991 ;
  assign n50993 = n11623 & ~n50992 ;
  assign n50995 = n39496 & n50859 ;
  assign n50996 = n36672 & ~n50995 ;
  assign n50998 = ~n43563 & n50996 ;
  assign n50997 = n43563 & ~n50996 ;
  assign n50999 = ~\P2_P1_DataWidth_reg[1]/NET0131  & ~n50997 ;
  assign n51000 = ~n50998 & n50999 ;
  assign n50994 = \P2_P1_DataWidth_reg[1]/NET0131  & ~\P2_P1_rEIP_reg[25]/NET0131  ;
  assign n51001 = n11609 & ~n50994 ;
  assign n51002 = ~n51000 & n51001 ;
  assign n50960 = \P2_P1_PhyAddrPointer_reg[25]/NET0131  & n11625 ;
  assign n50961 = \P2_P1_rEIP_reg[25]/NET0131  & ~n50411 ;
  assign n51003 = ~n50960 & ~n50961 ;
  assign n51004 = ~n51002 & n51003 ;
  assign n51005 = ~n50993 & n51004 ;
  assign n51015 = ~\P2_P1_EBX_reg[25]/NET0131  & n50983 ;
  assign n51016 = \P2_P1_EBX_reg[31]/NET0131  & ~n51015 ;
  assign n51018 = ~\P2_P1_EBX_reg[26]/NET0131  & n51016 ;
  assign n51017 = \P2_P1_EBX_reg[26]/NET0131  & ~n51016 ;
  assign n51019 = ~n50422 & ~n51017 ;
  assign n51020 = ~n51018 & n51019 ;
  assign n51009 = \P2_P1_rEIP_reg[24]/NET0131  & \P2_P1_rEIP_reg[25]/NET0131  ;
  assign n51010 = n50895 & n51009 ;
  assign n51011 = ~\P2_P1_rEIP_reg[26]/NET0131  & ~n51010 ;
  assign n51012 = \P2_P1_rEIP_reg[26]/NET0131  & n51010 ;
  assign n51013 = ~n51011 & ~n51012 ;
  assign n51014 = n50422 & ~n51013 ;
  assign n51021 = n24901 & ~n51014 ;
  assign n51022 = ~n51020 & n51021 ;
  assign n51008 = \P2_P1_rEIP_reg[26]/NET0131  & ~n50414 ;
  assign n51024 = n26103 & ~n51013 ;
  assign n51023 = ~\P2_P1_EBX_reg[26]/NET0131  & ~n26103 ;
  assign n51025 = n24899 & ~n51023 ;
  assign n51026 = ~n51024 & n51025 ;
  assign n51027 = ~n51008 & ~n51026 ;
  assign n51028 = ~n51022 & n51027 ;
  assign n51029 = n11623 & ~n51028 ;
  assign n51031 = n36662 & n50824 ;
  assign n51032 = n36672 & ~n51031 ;
  assign n51034 = n41637 & n51032 ;
  assign n51033 = ~n41637 & ~n51032 ;
  assign n51035 = ~\P2_P1_DataWidth_reg[1]/NET0131  & ~n51033 ;
  assign n51036 = ~n51034 & n51035 ;
  assign n51030 = \P2_P1_DataWidth_reg[1]/NET0131  & ~\P2_P1_rEIP_reg[26]/NET0131  ;
  assign n51037 = n11609 & ~n51030 ;
  assign n51038 = ~n51036 & n51037 ;
  assign n51006 = \P2_P1_PhyAddrPointer_reg[26]/NET0131  & n11625 ;
  assign n51007 = \P2_P1_rEIP_reg[26]/NET0131  & ~n50411 ;
  assign n51039 = ~n51006 & ~n51007 ;
  assign n51040 = ~n51038 & n51039 ;
  assign n51041 = ~n51029 & n51040 ;
  assign n51057 = ~\P2_P1_EBX_reg[26]/NET0131  & n51015 ;
  assign n51058 = \P2_P1_EBX_reg[31]/NET0131  & ~n51057 ;
  assign n51060 = ~\P2_P1_EBX_reg[27]/NET0131  & n51058 ;
  assign n51059 = \P2_P1_EBX_reg[27]/NET0131  & ~n51058 ;
  assign n51061 = ~n50422 & ~n51059 ;
  assign n51062 = ~n51060 & n51061 ;
  assign n51053 = ~\P2_P1_rEIP_reg[27]/NET0131  & ~n51012 ;
  assign n51054 = \P2_P1_rEIP_reg[27]/NET0131  & n51012 ;
  assign n51055 = ~n51053 & ~n51054 ;
  assign n51056 = n50422 & ~n51055 ;
  assign n51063 = n24901 & ~n51056 ;
  assign n51064 = ~n51062 & n51063 ;
  assign n51052 = \P2_P1_rEIP_reg[27]/NET0131  & ~n50414 ;
  assign n51066 = n26103 & ~n51055 ;
  assign n51065 = ~\P2_P1_EBX_reg[27]/NET0131  & ~n26103 ;
  assign n51067 = n24899 & ~n51065 ;
  assign n51068 = ~n51066 & n51067 ;
  assign n51069 = ~n51052 & ~n51068 ;
  assign n51070 = ~n51064 & n51069 ;
  assign n51071 = n11623 & ~n51070 ;
  assign n51044 = n41637 & n51031 ;
  assign n51045 = n36672 & ~n51044 ;
  assign n51047 = n39501 & ~n51045 ;
  assign n51046 = ~n39501 & n51045 ;
  assign n51048 = ~\P2_P1_DataWidth_reg[1]/NET0131  & ~n51046 ;
  assign n51049 = ~n51047 & n51048 ;
  assign n51043 = \P2_P1_DataWidth_reg[1]/NET0131  & ~\P2_P1_rEIP_reg[27]/NET0131  ;
  assign n51050 = n11609 & ~n51043 ;
  assign n51051 = ~n51049 & n51050 ;
  assign n51042 = \P2_P1_PhyAddrPointer_reg[27]/NET0131  & n11625 ;
  assign n51072 = \P2_P1_rEIP_reg[27]/NET0131  & ~n50411 ;
  assign n51073 = ~n51042 & ~n51072 ;
  assign n51074 = ~n51051 & n51073 ;
  assign n51075 = ~n51071 & n51074 ;
  assign n51087 = ~\P2_P1_EBX_reg[27]/NET0131  & n51057 ;
  assign n51088 = \P2_P1_EBX_reg[31]/NET0131  & ~n51087 ;
  assign n51090 = \P2_P1_EBX_reg[28]/NET0131  & ~n51088 ;
  assign n51089 = ~\P2_P1_EBX_reg[28]/NET0131  & n51088 ;
  assign n51091 = ~n50422 & ~n51089 ;
  assign n51092 = ~n51090 & n51091 ;
  assign n51079 = ~\P2_P1_rEIP_reg[28]/NET0131  & ~n51054 ;
  assign n51080 = \P2_P1_rEIP_reg[27]/NET0131  & \P2_P1_rEIP_reg[28]/NET0131  ;
  assign n51081 = n51012 & n51080 ;
  assign n51082 = ~n51079 & ~n51081 ;
  assign n51083 = n50422 & ~n51082 ;
  assign n51093 = n24901 & ~n51083 ;
  assign n51094 = ~n51092 & n51093 ;
  assign n51077 = \P2_P1_rEIP_reg[28]/NET0131  & ~n50414 ;
  assign n51084 = ~n25958 & n51083 ;
  assign n51078 = ~\P2_P1_EBX_reg[28]/NET0131  & ~n26103 ;
  assign n51085 = n24899 & ~n51078 ;
  assign n51086 = ~n51084 & n51085 ;
  assign n51095 = ~n51077 & ~n51086 ;
  assign n51096 = ~n51094 & n51095 ;
  assign n51097 = n11623 & ~n51096 ;
  assign n51100 = ~n39501 & n51044 ;
  assign n51101 = n36672 & ~n51100 ;
  assign n51103 = n39523 & ~n51101 ;
  assign n51102 = ~n39523 & n51101 ;
  assign n51104 = ~\P2_P1_DataWidth_reg[1]/NET0131  & ~n51102 ;
  assign n51105 = ~n51103 & n51104 ;
  assign n51099 = \P2_P1_DataWidth_reg[1]/NET0131  & ~\P2_P1_rEIP_reg[28]/NET0131  ;
  assign n51106 = n11609 & ~n51099 ;
  assign n51107 = ~n51105 & n51106 ;
  assign n51076 = \P2_P1_PhyAddrPointer_reg[28]/NET0131  & n11625 ;
  assign n51098 = \P2_P1_rEIP_reg[28]/NET0131  & ~n50411 ;
  assign n51108 = ~n51076 & ~n51098 ;
  assign n51109 = ~n51107 & n51108 ;
  assign n51110 = ~n51097 & n51109 ;
  assign n51117 = ~\P2_P1_EBX_reg[28]/NET0131  & n51087 ;
  assign n51118 = \P2_P1_EBX_reg[31]/NET0131  & ~n51117 ;
  assign n51120 = \P2_P1_EBX_reg[29]/NET0131  & ~n51118 ;
  assign n51119 = ~\P2_P1_EBX_reg[29]/NET0131  & n51118 ;
  assign n51121 = ~n50422 & ~n51119 ;
  assign n51122 = ~n51120 & n51121 ;
  assign n51113 = ~\P2_P1_rEIP_reg[29]/NET0131  & ~n51081 ;
  assign n51114 = \P2_P1_rEIP_reg[29]/NET0131  & n51081 ;
  assign n51115 = ~n51113 & ~n51114 ;
  assign n51116 = n50422 & ~n51115 ;
  assign n51123 = n24901 & ~n51116 ;
  assign n51124 = ~n51122 & n51123 ;
  assign n51112 = \P2_P1_rEIP_reg[29]/NET0131  & ~n50414 ;
  assign n51126 = n26103 & ~n51115 ;
  assign n51125 = ~\P2_P1_EBX_reg[29]/NET0131  & ~n26103 ;
  assign n51127 = n24899 & ~n51125 ;
  assign n51128 = ~n51126 & n51127 ;
  assign n51129 = ~n51112 & ~n51128 ;
  assign n51130 = ~n51124 & n51129 ;
  assign n51131 = n11623 & ~n51130 ;
  assign n51134 = ~n39523 & n51100 ;
  assign n51135 = n36672 & ~n51134 ;
  assign n51137 = n39540 & ~n51135 ;
  assign n51136 = ~n39540 & n51135 ;
  assign n51138 = ~\P2_P1_DataWidth_reg[1]/NET0131  & ~n51136 ;
  assign n51139 = ~n51137 & n51138 ;
  assign n51133 = \P2_P1_DataWidth_reg[1]/NET0131  & ~\P2_P1_rEIP_reg[29]/NET0131  ;
  assign n51140 = n11609 & ~n51133 ;
  assign n51141 = ~n51139 & n51140 ;
  assign n51111 = \P2_P1_PhyAddrPointer_reg[29]/NET0131  & n11625 ;
  assign n51132 = \P2_P1_rEIP_reg[29]/NET0131  & ~n50411 ;
  assign n51142 = ~n51111 & ~n51132 ;
  assign n51143 = ~n51141 & n51142 ;
  assign n51144 = ~n51131 & n51143 ;
  assign n51146 = n50475 & n50477 ;
  assign n51147 = ~n50478 & ~n51146 ;
  assign n51148 = ~\P2_P1_DataWidth_reg[1]/NET0131  & ~n51147 ;
  assign n51149 = \P2_P1_DataWidth_reg[1]/NET0131  & ~\P2_P1_rEIP_reg[2]/NET0131  ;
  assign n51150 = n11609 & ~n51149 ;
  assign n51151 = ~n51148 & n51150 ;
  assign n51153 = \P2_P1_rEIP_reg[2]/NET0131  & ~n50414 ;
  assign n51155 = ~\P2_P1_rEIP_reg[1]/NET0131  & ~\P2_P1_rEIP_reg[2]/NET0131  ;
  assign n51156 = ~\P2_P1_DataWidth_reg[1]/NET0131  & ~n50494 ;
  assign n51157 = ~n51155 & n51156 ;
  assign n51162 = ~n21073 & n51157 ;
  assign n51163 = \P2_P1_EBX_reg[31]/NET0131  & ~n50423 ;
  assign n51165 = \P2_P1_EBX_reg[2]/NET0131  & n51163 ;
  assign n51164 = ~\P2_P1_EBX_reg[2]/NET0131  & ~n51163 ;
  assign n51166 = ~n50422 & ~n51164 ;
  assign n51167 = ~n51165 & n51166 ;
  assign n51168 = ~n51162 & ~n51167 ;
  assign n51169 = n21062 & ~n51168 ;
  assign n51154 = \P2_P1_EBX_reg[2]/NET0131  & ~n26103 ;
  assign n51158 = n25959 & n51157 ;
  assign n51159 = ~n51154 & ~n51158 ;
  assign n51160 = n24898 & ~n51159 ;
  assign n51161 = n21067 & n26028 ;
  assign n51170 = ~n51160 & ~n51161 ;
  assign n51171 = ~n51169 & n51170 ;
  assign n51172 = ~n21081 & ~n51171 ;
  assign n51173 = ~n51153 & ~n51172 ;
  assign n51174 = n11623 & ~n51173 ;
  assign n51145 = \P2_P1_PhyAddrPointer_reg[2]/NET0131  & n11625 ;
  assign n51152 = \P2_P1_rEIP_reg[2]/NET0131  & ~n50411 ;
  assign n51175 = ~n51145 & ~n51152 ;
  assign n51176 = ~n51174 & n51175 ;
  assign n51177 = ~n51151 & n51176 ;
  assign n51180 = ~\P1_P2_PhyAddrPointer_reg[19]/NET0131  & ~n36628 ;
  assign n51181 = ~n36628 & ~n48456 ;
  assign n51182 = ~n36628 & ~n41414 ;
  assign n51183 = ~n51181 & ~n51182 ;
  assign n51184 = ~n51180 & n51183 ;
  assign n51186 = n41443 & n51184 ;
  assign n51185 = ~n41443 & ~n51184 ;
  assign n51187 = ~\P1_P2_DataWidth_reg[1]/NET0131  & ~n51185 ;
  assign n51188 = ~n51186 & n51187 ;
  assign n51179 = \P1_P2_DataWidth_reg[1]/NET0131  & ~\P1_P2_rEIP_reg[20]/NET0131  ;
  assign n51189 = n25928 & ~n51179 ;
  assign n51190 = ~n51188 & n51189 ;
  assign n51213 = \P1_P2_EBX_reg[31]/NET0131  & ~n48425 ;
  assign n51215 = ~\P1_P2_EBX_reg[20]/NET0131  & n51213 ;
  assign n51214 = \P1_P2_EBX_reg[20]/NET0131  & ~n51213 ;
  assign n51216 = ~n48373 & ~n51214 ;
  assign n51217 = ~n51215 & n51216 ;
  assign n51198 = \P1_P2_rEIP_reg[15]/NET0131  & n48391 ;
  assign n51199 = \P1_P2_rEIP_reg[8]/NET0131  & n48393 ;
  assign n51200 = n51198 & n51199 ;
  assign n51201 = n48385 & n51200 ;
  assign n51202 = n48388 & n51201 ;
  assign n51203 = \P1_P2_rEIP_reg[19]/NET0131  & n51202 ;
  assign n51205 = ~\P1_P2_rEIP_reg[20]/NET0131  & n51203 ;
  assign n51204 = \P1_P2_rEIP_reg[20]/NET0131  & ~n51203 ;
  assign n51206 = n48373 & ~n51204 ;
  assign n51207 = ~n51205 & n51206 ;
  assign n51218 = n25846 & ~n51207 ;
  assign n51219 = ~n51217 & n51218 ;
  assign n51191 = n25757 & ~n25761 ;
  assign n51192 = ~n48371 & ~n51191 ;
  assign n51193 = \P1_P2_rEIP_reg[20]/NET0131  & n51192 ;
  assign n51197 = ~\P1_P2_EBX_reg[20]/NET0131  & ~n48373 ;
  assign n51208 = n25841 & ~n51197 ;
  assign n51209 = ~n51207 & n51208 ;
  assign n51194 = n25768 & ~n25770 ;
  assign n51195 = \P1_P2_EBX_reg[20]/NET0131  & n51194 ;
  assign n51196 = \P1_P2_rEIP_reg[20]/NET0131  & n25770 ;
  assign n51210 = ~n51195 & ~n51196 ;
  assign n51211 = ~n51209 & n51210 ;
  assign n51212 = n25757 & ~n51211 ;
  assign n51220 = ~n51193 & ~n51212 ;
  assign n51221 = ~n51219 & n51220 ;
  assign n51222 = n25918 & ~n51221 ;
  assign n51178 = \P1_P2_PhyAddrPointer_reg[20]/NET0131  & n27675 ;
  assign n51223 = \P1_P2_rEIP_reg[20]/NET0131  & ~n48452 ;
  assign n51224 = ~n51178 & ~n51223 ;
  assign n51225 = ~n51222 & n51224 ;
  assign n51226 = ~n51190 & n51225 ;
  assign n51229 = ~n36628 & ~n48457 ;
  assign n51231 = n43397 & ~n51229 ;
  assign n51230 = ~n43397 & n51229 ;
  assign n51232 = ~\P1_P2_DataWidth_reg[1]/NET0131  & ~n51230 ;
  assign n51233 = ~n51231 & n51232 ;
  assign n51228 = \P1_P2_DataWidth_reg[1]/NET0131  & ~\P1_P2_rEIP_reg[21]/NET0131  ;
  assign n51234 = n25928 & ~n51228 ;
  assign n51235 = ~n51233 & n51234 ;
  assign n51248 = \P1_P2_EBX_reg[31]/NET0131  & ~n48426 ;
  assign n51250 = \P1_P2_EBX_reg[21]/NET0131  & ~n51248 ;
  assign n51249 = ~\P1_P2_EBX_reg[21]/NET0131  & n51248 ;
  assign n51251 = ~n48373 & ~n51249 ;
  assign n51252 = ~n51250 & n51251 ;
  assign n51237 = n48378 & n48396 ;
  assign n51238 = \P1_P2_rEIP_reg[18]/NET0131  & n48377 ;
  assign n51239 = \P1_P2_rEIP_reg[9]/NET0131  & n48386 ;
  assign n51240 = n48392 & n51239 ;
  assign n51241 = \P1_P2_rEIP_reg[16]/NET0131  & n51198 ;
  assign n51242 = n51240 & n51241 ;
  assign n51243 = \P1_P2_rEIP_reg[17]/NET0131  & n51242 ;
  assign n51244 = n51238 & n51243 ;
  assign n51245 = ~\P1_P2_rEIP_reg[21]/NET0131  & ~n51244 ;
  assign n51246 = ~n51237 & ~n51245 ;
  assign n51247 = n48373 & ~n51246 ;
  assign n51253 = n25846 & ~n51247 ;
  assign n51254 = ~n51252 & n51253 ;
  assign n51236 = \P1_P2_rEIP_reg[21]/NET0131  & ~n48371 ;
  assign n51256 = n48443 & ~n51246 ;
  assign n51255 = ~\P1_P2_EBX_reg[21]/NET0131  & ~n48443 ;
  assign n51257 = n47570 & ~n51255 ;
  assign n51258 = ~n51256 & n51257 ;
  assign n51259 = ~n51236 & ~n51258 ;
  assign n51260 = ~n51254 & n51259 ;
  assign n51261 = n25918 & ~n51260 ;
  assign n51227 = \P1_P2_PhyAddrPointer_reg[21]/NET0131  & n27675 ;
  assign n51262 = \P1_P2_rEIP_reg[21]/NET0131  & ~n48452 ;
  assign n51263 = ~n51227 & ~n51262 ;
  assign n51264 = ~n51261 & n51263 ;
  assign n51265 = ~n51235 & n51264 ;
  assign n51268 = ~n36628 & ~n48458 ;
  assign n51270 = ~n41459 & n51268 ;
  assign n51269 = n41459 & ~n51268 ;
  assign n51271 = ~\P1_P2_DataWidth_reg[1]/NET0131  & ~n51269 ;
  assign n51272 = ~n51270 & n51271 ;
  assign n51267 = \P1_P2_DataWidth_reg[1]/NET0131  & ~\P1_P2_rEIP_reg[22]/NET0131  ;
  assign n51273 = n25928 & ~n51267 ;
  assign n51274 = ~n51272 & n51273 ;
  assign n51279 = \P1_P2_EBX_reg[31]/NET0131  & ~n48427 ;
  assign n51281 = ~\P1_P2_EBX_reg[22]/NET0131  & n51279 ;
  assign n51280 = \P1_P2_EBX_reg[22]/NET0131  & ~n51279 ;
  assign n51282 = ~n48373 & ~n51280 ;
  assign n51283 = ~n51281 & n51282 ;
  assign n51276 = ~\P1_P2_rEIP_reg[22]/NET0131  & ~n51237 ;
  assign n51277 = ~n48397 & ~n51276 ;
  assign n51278 = n48373 & ~n51277 ;
  assign n51284 = n25846 & ~n51278 ;
  assign n51285 = ~n51283 & n51284 ;
  assign n51275 = \P1_P2_rEIP_reg[22]/NET0131  & ~n48371 ;
  assign n51286 = ~\P1_P2_EBX_reg[22]/NET0131  & ~n48443 ;
  assign n51287 = n48443 & ~n51277 ;
  assign n51288 = ~n51286 & ~n51287 ;
  assign n51289 = n47570 & n51288 ;
  assign n51290 = ~n51275 & ~n51289 ;
  assign n51291 = ~n51285 & n51290 ;
  assign n51292 = n25918 & ~n51291 ;
  assign n51266 = \P1_P2_PhyAddrPointer_reg[22]/NET0131  & n27675 ;
  assign n51293 = \P1_P2_rEIP_reg[22]/NET0131  & ~n48452 ;
  assign n51294 = ~n51266 & ~n51293 ;
  assign n51295 = ~n51292 & n51294 ;
  assign n51296 = ~n51274 & n51295 ;
  assign n51299 = ~n36616 & ~n36628 ;
  assign n51300 = ~n51229 & ~n51299 ;
  assign n51302 = ~n39375 & ~n51300 ;
  assign n51301 = n39375 & n51300 ;
  assign n51303 = ~\P1_P2_DataWidth_reg[1]/NET0131  & ~n51301 ;
  assign n51304 = ~n51302 & n51303 ;
  assign n51298 = \P1_P2_DataWidth_reg[1]/NET0131  & ~\P1_P2_rEIP_reg[23]/NET0131  ;
  assign n51305 = n25928 & ~n51298 ;
  assign n51306 = ~n51304 & n51305 ;
  assign n51323 = \P1_P2_EBX_reg[31]/NET0131  & ~n48428 ;
  assign n51325 = ~\P1_P2_EBX_reg[23]/NET0131  & n51323 ;
  assign n51324 = \P1_P2_EBX_reg[23]/NET0131  & ~n51323 ;
  assign n51326 = ~n48373 & ~n51324 ;
  assign n51327 = ~n51325 & n51326 ;
  assign n51310 = n48379 & n51202 ;
  assign n51311 = ~\P1_P2_rEIP_reg[23]/NET0131  & ~n51310 ;
  assign n51312 = \P1_P2_rEIP_reg[23]/NET0131  & n48388 ;
  assign n51313 = n48379 & n51312 ;
  assign n51314 = n51201 & n51313 ;
  assign n51315 = ~n51311 & ~n51314 ;
  assign n51316 = n48373 & ~n51315 ;
  assign n51328 = n25846 & ~n51316 ;
  assign n51329 = ~n51327 & n51328 ;
  assign n51307 = \P1_P2_rEIP_reg[23]/NET0131  & n51192 ;
  assign n51317 = ~\P1_P2_EBX_reg[23]/NET0131  & ~n48373 ;
  assign n51318 = n25841 & ~n51317 ;
  assign n51319 = ~n51316 & n51318 ;
  assign n51308 = \P1_P2_EBX_reg[23]/NET0131  & n51194 ;
  assign n51309 = \P1_P2_rEIP_reg[23]/NET0131  & n25770 ;
  assign n51320 = ~n51308 & ~n51309 ;
  assign n51321 = ~n51319 & n51320 ;
  assign n51322 = n25757 & ~n51321 ;
  assign n51330 = ~n51307 & ~n51322 ;
  assign n51331 = ~n51329 & n51330 ;
  assign n51332 = n25918 & ~n51331 ;
  assign n51297 = \P1_P2_PhyAddrPointer_reg[23]/NET0131  & n27675 ;
  assign n51333 = \P1_P2_rEIP_reg[23]/NET0131  & ~n48452 ;
  assign n51334 = ~n51297 & ~n51333 ;
  assign n51335 = ~n51332 & n51334 ;
  assign n51336 = ~n51306 & n51335 ;
  assign n51339 = ~n36617 & ~n36628 ;
  assign n51340 = ~n51229 & ~n51339 ;
  assign n51342 = n41477 & n51340 ;
  assign n51341 = ~n41477 & ~n51340 ;
  assign n51343 = ~\P1_P2_DataWidth_reg[1]/NET0131  & ~n51341 ;
  assign n51344 = ~n51342 & n51343 ;
  assign n51338 = \P1_P2_DataWidth_reg[1]/NET0131  & ~\P1_P2_rEIP_reg[24]/NET0131  ;
  assign n51345 = n25928 & ~n51338 ;
  assign n51346 = ~n51344 & n51345 ;
  assign n51349 = n51200 & n51313 ;
  assign n51350 = ~\P1_P2_rEIP_reg[24]/NET0131  & n51349 ;
  assign n51351 = \P1_P2_rEIP_reg[24]/NET0131  & ~n51349 ;
  assign n51352 = ~n51350 & ~n51351 ;
  assign n51353 = n48385 & n51352 ;
  assign n51348 = ~\P1_P2_rEIP_reg[24]/NET0131  & ~n48385 ;
  assign n51354 = n48373 & ~n51348 ;
  assign n51355 = ~n51353 & n51354 ;
  assign n51356 = \P1_P2_EBX_reg[31]/NET0131  & ~n48429 ;
  assign n51358 = \P1_P2_EBX_reg[24]/NET0131  & n51356 ;
  assign n51357 = ~\P1_P2_EBX_reg[24]/NET0131  & ~n51356 ;
  assign n51359 = ~n48373 & ~n51357 ;
  assign n51360 = ~n51358 & n51359 ;
  assign n51361 = ~n51355 & ~n51360 ;
  assign n51362 = n25846 & ~n51361 ;
  assign n51347 = \P1_P2_rEIP_reg[24]/NET0131  & n51192 ;
  assign n51365 = \P1_P2_EBX_reg[24]/NET0131  & ~n48373 ;
  assign n51366 = ~n51355 & ~n51365 ;
  assign n51367 = n25841 & ~n51366 ;
  assign n51363 = \P1_P2_rEIP_reg[24]/NET0131  & n25770 ;
  assign n51364 = \P1_P2_EBX_reg[24]/NET0131  & n51194 ;
  assign n51368 = ~n51363 & ~n51364 ;
  assign n51369 = ~n51367 & n51368 ;
  assign n51370 = n25757 & ~n51369 ;
  assign n51371 = ~n51347 & ~n51370 ;
  assign n51372 = ~n51362 & n51371 ;
  assign n51373 = n25918 & ~n51372 ;
  assign n51337 = \P1_P2_PhyAddrPointer_reg[24]/NET0131  & n27675 ;
  assign n51374 = \P1_P2_rEIP_reg[24]/NET0131  & ~n48452 ;
  assign n51375 = ~n51337 & ~n51374 ;
  assign n51376 = ~n51373 & n51375 ;
  assign n51377 = ~n51346 & n51376 ;
  assign n51380 = ~n41459 & ~n43397 ;
  assign n51381 = ~n39375 & n51380 ;
  assign n51382 = ~n41477 & n51381 ;
  assign n51383 = ~\P1_P2_PhyAddrPointer_reg[0]/NET0131  & n43520 ;
  assign n51384 = n36605 & n51383 ;
  assign n51385 = ~n43295 & n51384 ;
  assign n51386 = ~n43323 & n51385 ;
  assign n51387 = ~n41395 & n51386 ;
  assign n51388 = ~n39337 & n51387 ;
  assign n51389 = ~n43332 & n51388 ;
  assign n51390 = ~n43360 & n51389 ;
  assign n51391 = ~n43371 & n51390 ;
  assign n51392 = ~n41416 & n51391 ;
  assign n51393 = ~n41443 & n51392 ;
  assign n51394 = n51382 & n51393 ;
  assign n51395 = ~n36628 & ~n51394 ;
  assign n51397 = n43415 & ~n51395 ;
  assign n51396 = ~n43415 & n51395 ;
  assign n51398 = ~\P1_P2_DataWidth_reg[1]/NET0131  & ~n51396 ;
  assign n51399 = ~n51397 & n51398 ;
  assign n51379 = \P1_P2_DataWidth_reg[1]/NET0131  & ~\P1_P2_rEIP_reg[25]/NET0131  ;
  assign n51400 = n25928 & ~n51379 ;
  assign n51401 = ~n51399 & n51400 ;
  assign n51416 = \P1_P2_EBX_reg[31]/NET0131  & ~n48430 ;
  assign n51418 = ~\P1_P2_EBX_reg[25]/NET0131  & n51416 ;
  assign n51417 = \P1_P2_EBX_reg[25]/NET0131  & ~n51416 ;
  assign n51419 = ~n48373 & ~n51417 ;
  assign n51420 = ~n51418 & n51419 ;
  assign n51410 = \P1_P2_rEIP_reg[25]/NET0131  & ~n48386 ;
  assign n51404 = n48374 & n48379 ;
  assign n51405 = n48395 & n51404 ;
  assign n51406 = ~\P1_P2_rEIP_reg[25]/NET0131  & ~n51405 ;
  assign n51407 = \P1_P2_rEIP_reg[25]/NET0131  & n51405 ;
  assign n51408 = ~n51406 & ~n51407 ;
  assign n51409 = n48386 & n51408 ;
  assign n51411 = n48373 & ~n51409 ;
  assign n51412 = ~n51410 & n51411 ;
  assign n51421 = n25846 & ~n51412 ;
  assign n51422 = ~n51420 & n51421 ;
  assign n51402 = \P1_P2_rEIP_reg[25]/NET0131  & ~n48371 ;
  assign n51403 = ~\P1_P2_EBX_reg[25]/NET0131  & ~n48443 ;
  assign n51413 = ~n25768 & n51412 ;
  assign n51414 = ~n51403 & ~n51413 ;
  assign n51415 = n47570 & n51414 ;
  assign n51423 = ~n51402 & ~n51415 ;
  assign n51424 = ~n51422 & n51423 ;
  assign n51425 = n25918 & ~n51424 ;
  assign n51378 = \P1_P2_PhyAddrPointer_reg[25]/NET0131  & n27675 ;
  assign n51426 = \P1_P2_rEIP_reg[25]/NET0131  & ~n48452 ;
  assign n51427 = ~n51378 & ~n51426 ;
  assign n51428 = ~n51425 & n51427 ;
  assign n51429 = ~n51401 & n51428 ;
  assign n51432 = ~n36619 & ~n36628 ;
  assign n51433 = ~n51268 & ~n51432 ;
  assign n51435 = n41494 & n51433 ;
  assign n51434 = ~n41494 & ~n51433 ;
  assign n51436 = ~\P1_P2_DataWidth_reg[1]/NET0131  & ~n51434 ;
  assign n51437 = ~n51435 & n51436 ;
  assign n51431 = \P1_P2_DataWidth_reg[1]/NET0131  & ~\P1_P2_rEIP_reg[26]/NET0131  ;
  assign n51438 = n25928 & ~n51431 ;
  assign n51439 = ~n51437 & n51438 ;
  assign n51441 = n48386 & n51407 ;
  assign n51442 = ~\P1_P2_rEIP_reg[26]/NET0131  & ~n51441 ;
  assign n51443 = ~\P1_P2_DataWidth_reg[1]/NET0131  & ~n51442 ;
  assign n51444 = ~n48398 & n51443 ;
  assign n51445 = ~n25415 & n51444 ;
  assign n51446 = \P1_P2_EBX_reg[31]/NET0131  & ~n48431 ;
  assign n51448 = \P1_P2_EBX_reg[26]/NET0131  & n51446 ;
  assign n51447 = ~\P1_P2_EBX_reg[26]/NET0131  & ~n51446 ;
  assign n51449 = ~n48373 & ~n51447 ;
  assign n51450 = ~n51448 & n51449 ;
  assign n51451 = ~n51445 & ~n51450 ;
  assign n51452 = n25846 & ~n51451 ;
  assign n51440 = \P1_P2_rEIP_reg[26]/NET0131  & ~n48371 ;
  assign n51453 = \P1_P2_EBX_reg[26]/NET0131  & ~n48443 ;
  assign n51454 = n25769 & n51444 ;
  assign n51455 = ~n51453 & ~n51454 ;
  assign n51456 = n47570 & ~n51455 ;
  assign n51457 = ~n51440 & ~n51456 ;
  assign n51458 = ~n51452 & n51457 ;
  assign n51459 = n25918 & ~n51458 ;
  assign n51430 = \P1_P2_PhyAddrPointer_reg[26]/NET0131  & n27675 ;
  assign n51460 = \P1_P2_rEIP_reg[26]/NET0131  & ~n48452 ;
  assign n51461 = ~n51430 & ~n51460 ;
  assign n51462 = ~n51459 & n51461 ;
  assign n51463 = ~n51439 & n51462 ;
  assign n51466 = ~n36620 & ~n36628 ;
  assign n51467 = ~n51268 & ~n51466 ;
  assign n51469 = n39387 & n51467 ;
  assign n51468 = ~n39387 & ~n51467 ;
  assign n51470 = ~\P1_P2_DataWidth_reg[1]/NET0131  & ~n51468 ;
  assign n51471 = ~n51469 & n51470 ;
  assign n51465 = \P1_P2_DataWidth_reg[1]/NET0131  & ~\P1_P2_rEIP_reg[27]/NET0131  ;
  assign n51472 = n25928 & ~n51465 ;
  assign n51473 = ~n51471 & n51472 ;
  assign n51485 = \P1_P2_EBX_reg[31]/NET0131  & ~n48432 ;
  assign n51487 = ~\P1_P2_EBX_reg[27]/NET0131  & n51485 ;
  assign n51486 = \P1_P2_EBX_reg[27]/NET0131  & ~n51485 ;
  assign n51488 = ~n48373 & ~n51486 ;
  assign n51489 = ~n51487 & n51488 ;
  assign n51475 = ~\P1_P2_rEIP_reg[27]/NET0131  & ~n48398 ;
  assign n51476 = ~n48399 & ~n51475 ;
  assign n51484 = n48373 & ~n51476 ;
  assign n51490 = n25846 & ~n51484 ;
  assign n51491 = ~n51489 & n51490 ;
  assign n51477 = n48443 & n51476 ;
  assign n51474 = \P1_P2_EBX_reg[27]/NET0131  & ~n48443 ;
  assign n51478 = ~n25770 & ~n51474 ;
  assign n51479 = ~n51477 & n51478 ;
  assign n51480 = n25757 & ~n51479 ;
  assign n51481 = ~n25770 & n51480 ;
  assign n51482 = ~n51192 & ~n51480 ;
  assign n51483 = \P1_P2_rEIP_reg[27]/NET0131  & ~n51482 ;
  assign n51492 = ~n51481 & ~n51483 ;
  assign n51493 = ~n51491 & n51492 ;
  assign n51494 = n25918 & ~n51493 ;
  assign n51464 = \P1_P2_PhyAddrPointer_reg[27]/NET0131  & n27675 ;
  assign n51495 = \P1_P2_rEIP_reg[27]/NET0131  & ~n48452 ;
  assign n51496 = ~n51464 & ~n51495 ;
  assign n51497 = ~n51494 & n51496 ;
  assign n51498 = ~n51473 & n51497 ;
  assign n51501 = ~n36621 & ~n36628 ;
  assign n51502 = ~n51268 & ~n51501 ;
  assign n51504 = n39412 & n51502 ;
  assign n51503 = ~n39412 & ~n51502 ;
  assign n51505 = ~\P1_P2_DataWidth_reg[1]/NET0131  & ~n51503 ;
  assign n51506 = ~n51504 & n51505 ;
  assign n51500 = \P1_P2_DataWidth_reg[1]/NET0131  & ~\P1_P2_rEIP_reg[28]/NET0131  ;
  assign n51507 = n25928 & ~n51500 ;
  assign n51508 = ~n51506 & n51507 ;
  assign n51509 = \P1_P2_EBX_reg[31]/NET0131  & ~n48433 ;
  assign n51511 = \P1_P2_EBX_reg[28]/NET0131  & n51509 ;
  assign n51510 = ~\P1_P2_EBX_reg[28]/NET0131  & ~n51509 ;
  assign n51512 = ~n48373 & ~n51510 ;
  assign n51513 = ~n51511 & n51512 ;
  assign n51514 = \P1_P2_rEIP_reg[24]/NET0131  & \P1_P2_rEIP_reg[25]/NET0131  ;
  assign n51515 = \P1_P2_rEIP_reg[26]/NET0131  & \P1_P2_rEIP_reg[27]/NET0131  ;
  assign n51516 = n51514 & n51515 ;
  assign n51517 = n51198 & n51516 ;
  assign n51518 = n51313 & n51517 ;
  assign n51519 = n51240 & n51518 ;
  assign n51521 = \P1_P2_rEIP_reg[28]/NET0131  & n51519 ;
  assign n51520 = ~\P1_P2_rEIP_reg[28]/NET0131  & ~n51519 ;
  assign n51522 = n48373 & ~n51520 ;
  assign n51523 = ~n51521 & n51522 ;
  assign n51524 = ~n51513 & ~n51523 ;
  assign n51525 = n25846 & ~n51524 ;
  assign n51527 = n48443 & ~n51521 ;
  assign n51526 = \P1_P2_EBX_reg[28]/NET0131  & ~n48443 ;
  assign n51528 = ~n25770 & ~n51526 ;
  assign n51529 = ~n51527 & n51528 ;
  assign n51530 = n25757 & ~n51529 ;
  assign n51531 = ~n51192 & ~n51530 ;
  assign n51532 = \P1_P2_rEIP_reg[28]/NET0131  & ~n51531 ;
  assign n51533 = n48443 & ~n51519 ;
  assign n51534 = n47570 & ~n51533 ;
  assign n51535 = ~n51529 & n51534 ;
  assign n51536 = ~n51532 & ~n51535 ;
  assign n51537 = ~n51525 & n51536 ;
  assign n51538 = n25918 & ~n51537 ;
  assign n51499 = \P1_P2_PhyAddrPointer_reg[28]/NET0131  & n27675 ;
  assign n51539 = \P1_P2_rEIP_reg[28]/NET0131  & ~n48452 ;
  assign n51540 = ~n51499 & ~n51539 ;
  assign n51541 = ~n51538 & n51540 ;
  assign n51542 = ~n51508 & n51541 ;
  assign n51545 = ~n43415 & n48457 ;
  assign n51546 = n51382 & n51545 ;
  assign n51547 = ~n41494 & n51546 ;
  assign n51548 = ~n39387 & n51547 ;
  assign n51549 = ~n39412 & n51548 ;
  assign n51550 = ~n36628 & ~n51549 ;
  assign n51552 = n39438 & ~n51550 ;
  assign n51551 = ~n39438 & n51550 ;
  assign n51553 = ~\P1_P2_DataWidth_reg[1]/NET0131  & ~n51551 ;
  assign n51554 = ~n51552 & n51553 ;
  assign n51544 = \P1_P2_DataWidth_reg[1]/NET0131  & ~\P1_P2_rEIP_reg[29]/NET0131  ;
  assign n51555 = n25928 & ~n51544 ;
  assign n51556 = ~n51554 & n51555 ;
  assign n51570 = \P1_P2_EBX_reg[31]/NET0131  & ~n48434 ;
  assign n51572 = ~\P1_P2_EBX_reg[29]/NET0131  & n51570 ;
  assign n51571 = \P1_P2_EBX_reg[29]/NET0131  & ~n51570 ;
  assign n51573 = ~n48373 & ~n51571 ;
  assign n51574 = ~n51572 & n51573 ;
  assign n51560 = \P1_P2_rEIP_reg[28]/NET0131  & n48399 ;
  assign n51561 = ~\P1_P2_rEIP_reg[29]/NET0131  & ~n51560 ;
  assign n51562 = ~n48401 & ~n51561 ;
  assign n51563 = n48373 & ~n51562 ;
  assign n51575 = n25846 & ~n51563 ;
  assign n51576 = ~n51574 & n51575 ;
  assign n51557 = \P1_P2_rEIP_reg[29]/NET0131  & n51192 ;
  assign n51564 = ~\P1_P2_EBX_reg[29]/NET0131  & ~n48373 ;
  assign n51565 = n25841 & ~n51564 ;
  assign n51566 = ~n51563 & n51565 ;
  assign n51558 = \P1_P2_EBX_reg[29]/NET0131  & n51194 ;
  assign n51559 = \P1_P2_rEIP_reg[29]/NET0131  & n25770 ;
  assign n51567 = ~n51558 & ~n51559 ;
  assign n51568 = ~n51566 & n51567 ;
  assign n51569 = n25757 & ~n51568 ;
  assign n51577 = ~n51557 & ~n51569 ;
  assign n51578 = ~n51576 & n51577 ;
  assign n51579 = n25918 & ~n51578 ;
  assign n51543 = \P1_P2_PhyAddrPointer_reg[29]/NET0131  & n27675 ;
  assign n51580 = \P1_P2_rEIP_reg[29]/NET0131  & ~n48452 ;
  assign n51581 = ~n51543 & ~n51580 ;
  assign n51582 = ~n51579 & n51581 ;
  assign n51583 = ~n51556 & n51582 ;
  assign n51586 = ~\P1_P2_PhyAddrPointer_reg[1]/NET0131  & ~\P1_P2_PhyAddrPointer_reg[2]/NET0131  ;
  assign n51587 = ~n47384 & ~n51586 ;
  assign n51588 = ~n50439 & ~n50441 ;
  assign n51590 = ~n51587 & ~n51588 ;
  assign n51589 = n51587 & n51588 ;
  assign n51591 = ~\P1_P2_DataWidth_reg[1]/NET0131  & ~n51589 ;
  assign n51592 = ~n51590 & n51591 ;
  assign n51585 = \P1_P2_DataWidth_reg[1]/NET0131  & ~\P1_P2_rEIP_reg[2]/NET0131  ;
  assign n51593 = n25928 & ~n51585 ;
  assign n51594 = ~n51592 & n51593 ;
  assign n51596 = \P1_P2_rEIP_reg[2]/NET0131  & ~n48371 ;
  assign n51599 = ~\P1_P2_rEIP_reg[1]/NET0131  & ~\P1_P2_rEIP_reg[2]/NET0131  ;
  assign n51600 = ~\P1_P2_DataWidth_reg[1]/NET0131  & ~n48380 ;
  assign n51601 = ~n51599 & n51600 ;
  assign n51605 = ~n25415 & n51601 ;
  assign n51606 = \P1_P2_EBX_reg[31]/NET0131  & ~n48407 ;
  assign n51608 = \P1_P2_EBX_reg[2]/NET0131  & n51606 ;
  assign n51607 = ~\P1_P2_EBX_reg[2]/NET0131  & ~n51606 ;
  assign n51609 = ~n48373 & ~n51607 ;
  assign n51610 = ~n51608 & n51609 ;
  assign n51611 = ~n51605 & ~n51610 ;
  assign n51612 = n25776 & ~n51611 ;
  assign n51597 = n25761 & n25819 ;
  assign n51598 = \P1_P2_EBX_reg[2]/NET0131  & ~n48443 ;
  assign n51602 = n25769 & n51601 ;
  assign n51603 = ~n51598 & ~n51602 ;
  assign n51604 = n25757 & ~n51603 ;
  assign n51613 = ~n51597 & ~n51604 ;
  assign n51614 = ~n51612 & n51613 ;
  assign n51615 = ~n25770 & ~n51614 ;
  assign n51616 = ~n51596 & ~n51615 ;
  assign n51617 = n25918 & ~n51616 ;
  assign n51584 = \P1_P2_PhyAddrPointer_reg[2]/NET0131  & n27675 ;
  assign n51595 = \P1_P2_rEIP_reg[2]/NET0131  & ~n48452 ;
  assign n51618 = ~n51584 & ~n51595 ;
  assign n51619 = ~n51617 & n51618 ;
  assign n51620 = ~n51594 & n51619 ;
  assign n51631 = \P1_P2_rEIP_reg[31]/NET0131  & n48404 ;
  assign n51630 = ~\P1_P2_rEIP_reg[31]/NET0131  & ~n48404 ;
  assign n51632 = n48373 & ~n51630 ;
  assign n51633 = ~n51631 & n51632 ;
  assign n51640 = ~\P1_P2_EBX_reg[30]/NET0131  & n48435 ;
  assign n51641 = ~n51633 & ~n51640 ;
  assign n51629 = \P1_P2_EBX_reg[31]/NET0131  & ~n48373 ;
  assign n51634 = ~n51629 & ~n51633 ;
  assign n51642 = n25846 & ~n51634 ;
  assign n51643 = ~n51641 & n51642 ;
  assign n51627 = \P1_P2_rEIP_reg[31]/NET0131  & n51192 ;
  assign n51635 = n25841 & ~n51634 ;
  assign n51628 = \P1_P2_EBX_reg[31]/NET0131  & n51194 ;
  assign n51636 = \P1_P2_rEIP_reg[31]/NET0131  & n25770 ;
  assign n51637 = ~n51628 & ~n51636 ;
  assign n51638 = ~n51635 & n51637 ;
  assign n51639 = n25757 & ~n51638 ;
  assign n51644 = ~n51627 & ~n51639 ;
  assign n51645 = ~n51643 & n51644 ;
  assign n51646 = n25918 & ~n51645 ;
  assign n51622 = \P1_P2_DataWidth_reg[1]/NET0131  & \P1_P2_rEIP_reg[31]/NET0131  ;
  assign n51623 = ~\P1_P2_DataWidth_reg[1]/NET0131  & n48459 ;
  assign n51624 = n36627 & n51623 ;
  assign n51625 = ~n51622 & ~n51624 ;
  assign n51626 = n25928 & ~n51625 ;
  assign n51621 = \P1_P2_PhyAddrPointer_reg[31]/NET0131  & n27675 ;
  assign n51647 = \P1_P2_rEIP_reg[31]/NET0131  & ~n48452 ;
  assign n51648 = ~n51621 & ~n51647 ;
  assign n51649 = ~n51626 & n51648 ;
  assign n51650 = ~n51646 & n51649 ;
  assign n51653 = ~\P1_P1_PhyAddrPointer_reg[0]/NET0131  & n41711 ;
  assign n51654 = ~n36733 & ~n51653 ;
  assign n51655 = ~n36718 & ~n36733 ;
  assign n51656 = ~n51654 & ~n51655 ;
  assign n51658 = n41733 & n51656 ;
  assign n51657 = ~n41733 & ~n51656 ;
  assign n51659 = ~\P1_P1_DataWidth_reg[1]/NET0131  & ~n51657 ;
  assign n51660 = ~n51658 & n51659 ;
  assign n51652 = \P1_P1_DataWidth_reg[1]/NET0131  & ~\P1_P1_rEIP_reg[20]/NET0131  ;
  assign n51661 = n8282 & ~n51652 ;
  assign n51662 = ~n51660 & n51661 ;
  assign n51663 = \P1_P1_rEIP_reg[20]/NET0131  & ~n50559 ;
  assign n51665 = \P1_P1_rEIP_reg[17]/NET0131  & \P1_P1_rEIP_reg[18]/NET0131  ;
  assign n51666 = \P1_P1_rEIP_reg[19]/NET0131  & n51665 ;
  assign n51667 = \P1_P1_rEIP_reg[12]/NET0131  & \P1_P1_rEIP_reg[13]/NET0131  ;
  assign n51668 = \P1_P1_rEIP_reg[4]/NET0131  & n50601 ;
  assign n51669 = \P1_P1_rEIP_reg[5]/NET0131  & n51668 ;
  assign n51670 = \P1_P1_rEIP_reg[6]/NET0131  & n51669 ;
  assign n51671 = \P1_P1_rEIP_reg[7]/NET0131  & n51670 ;
  assign n51672 = \P1_P1_rEIP_reg[8]/NET0131  & n51671 ;
  assign n51673 = \P1_P1_rEIP_reg[9]/NET0131  & n51672 ;
  assign n51674 = \P1_P1_rEIP_reg[10]/NET0131  & n51673 ;
  assign n51675 = \P1_P1_rEIP_reg[11]/NET0131  & n51674 ;
  assign n51676 = n51667 & n51675 ;
  assign n51677 = \P1_P1_rEIP_reg[14]/NET0131  & n51676 ;
  assign n51678 = \P1_P1_rEIP_reg[15]/NET0131  & n51677 ;
  assign n51679 = \P1_P1_rEIP_reg[16]/NET0131  & n51678 ;
  assign n51680 = n51666 & n51679 ;
  assign n51681 = ~\P1_P1_rEIP_reg[20]/NET0131  & ~n51680 ;
  assign n51682 = \P1_P1_rEIP_reg[20]/NET0131  & n51680 ;
  assign n51683 = ~n51681 & ~n51682 ;
  assign n51684 = n26275 & ~n51683 ;
  assign n51664 = ~\P1_P1_EBX_reg[20]/NET0131  & ~n26275 ;
  assign n51685 = n24502 & ~n51664 ;
  assign n51686 = ~n51684 & n51685 ;
  assign n51688 = ~\P1_P1_EBX_reg[3]/NET0131  & n50609 ;
  assign n51689 = ~\P1_P1_EBX_reg[4]/NET0131  & n51688 ;
  assign n51690 = ~\P1_P1_EBX_reg[5]/NET0131  & n51689 ;
  assign n51691 = ~\P1_P1_EBX_reg[6]/NET0131  & n51690 ;
  assign n51692 = ~\P1_P1_EBX_reg[7]/NET0131  & n51691 ;
  assign n51693 = ~\P1_P1_EBX_reg[8]/NET0131  & n51692 ;
  assign n51694 = ~\P1_P1_EBX_reg[9]/NET0131  & n51693 ;
  assign n51695 = ~\P1_P1_EBX_reg[10]/NET0131  & n51694 ;
  assign n51696 = ~\P1_P1_EBX_reg[11]/NET0131  & n51695 ;
  assign n51697 = ~\P1_P1_EBX_reg[12]/NET0131  & n51696 ;
  assign n51698 = ~\P1_P1_EBX_reg[13]/NET0131  & n51697 ;
  assign n51699 = ~\P1_P1_EBX_reg[14]/NET0131  & n51698 ;
  assign n51700 = ~\P1_P1_EBX_reg[15]/NET0131  & n51699 ;
  assign n51701 = ~\P1_P1_EBX_reg[16]/NET0131  & n51700 ;
  assign n51702 = ~\P1_P1_EBX_reg[17]/NET0131  & n51701 ;
  assign n51703 = ~\P1_P1_EBX_reg[18]/NET0131  & n51702 ;
  assign n51704 = ~\P1_P1_EBX_reg[19]/NET0131  & n51703 ;
  assign n51705 = \P1_P1_EBX_reg[31]/NET0131  & ~n51704 ;
  assign n51707 = ~\P1_P1_EBX_reg[20]/NET0131  & n51705 ;
  assign n51706 = \P1_P1_EBX_reg[20]/NET0131  & ~n51705 ;
  assign n51708 = ~n26274 & ~n51706 ;
  assign n51709 = ~n51707 & n51708 ;
  assign n51687 = n26274 & ~n51683 ;
  assign n51710 = n15334 & ~n51687 ;
  assign n51711 = ~n51709 & n51710 ;
  assign n51712 = ~n51686 & ~n51711 ;
  assign n51713 = ~n15364 & ~n51712 ;
  assign n51714 = ~n51663 & ~n51713 ;
  assign n51715 = n8355 & ~n51714 ;
  assign n51651 = \P1_P1_PhyAddrPointer_reg[20]/NET0131  & n8361 ;
  assign n51716 = \P1_P1_rEIP_reg[20]/NET0131  & ~n50583 ;
  assign n51717 = ~n51651 & ~n51716 ;
  assign n51718 = ~n51715 & n51717 ;
  assign n51719 = ~n51662 & n51718 ;
  assign n51722 = ~n36719 & ~n36733 ;
  assign n51723 = ~n51654 & ~n51722 ;
  assign n51725 = ~n43701 & ~n51723 ;
  assign n51724 = n43701 & n51723 ;
  assign n51726 = ~\P1_P1_DataWidth_reg[1]/NET0131  & ~n51724 ;
  assign n51727 = ~n51725 & n51726 ;
  assign n51721 = \P1_P1_DataWidth_reg[1]/NET0131  & ~\P1_P1_rEIP_reg[21]/NET0131  ;
  assign n51728 = n8282 & ~n51721 ;
  assign n51729 = ~n51727 & n51728 ;
  assign n51730 = \P1_P1_rEIP_reg[21]/NET0131  & ~n50559 ;
  assign n51732 = ~\P1_P1_rEIP_reg[21]/NET0131  & ~n51682 ;
  assign n51733 = \P1_P1_rEIP_reg[15]/NET0131  & \P1_P1_rEIP_reg[16]/NET0131  ;
  assign n51734 = \P1_P1_rEIP_reg[20]/NET0131  & \P1_P1_rEIP_reg[21]/NET0131  ;
  assign n51735 = n51733 & n51734 ;
  assign n51736 = n51666 & n51735 ;
  assign n51737 = n51677 & n51736 ;
  assign n51738 = ~n51732 & ~n51737 ;
  assign n51739 = n26275 & ~n51738 ;
  assign n51731 = ~\P1_P1_EBX_reg[21]/NET0131  & ~n26275 ;
  assign n51740 = n24502 & ~n51731 ;
  assign n51741 = ~n51739 & n51740 ;
  assign n51743 = ~\P1_P1_EBX_reg[20]/NET0131  & n51704 ;
  assign n51744 = \P1_P1_EBX_reg[31]/NET0131  & ~n51743 ;
  assign n51746 = ~\P1_P1_EBX_reg[21]/NET0131  & n51744 ;
  assign n51745 = \P1_P1_EBX_reg[21]/NET0131  & ~n51744 ;
  assign n51747 = ~n26274 & ~n51745 ;
  assign n51748 = ~n51746 & n51747 ;
  assign n51742 = n26274 & ~n51738 ;
  assign n51749 = n15334 & ~n51742 ;
  assign n51750 = ~n51748 & n51749 ;
  assign n51751 = ~n51741 & ~n51750 ;
  assign n51752 = ~n15364 & ~n51751 ;
  assign n51753 = ~n51730 & ~n51752 ;
  assign n51754 = n8355 & ~n51753 ;
  assign n51720 = \P1_P1_PhyAddrPointer_reg[21]/NET0131  & n8361 ;
  assign n51755 = \P1_P1_rEIP_reg[21]/NET0131  & ~n50583 ;
  assign n51756 = ~n51720 & ~n51755 ;
  assign n51757 = ~n51754 & n51756 ;
  assign n51758 = ~n51729 & n51757 ;
  assign n51761 = ~n36720 & ~n36733 ;
  assign n51762 = \P1_P1_PhyAddrPointer_reg[17]/NET0131  & n51653 ;
  assign n51763 = ~n36733 & ~n51762 ;
  assign n51764 = ~n51761 & ~n51763 ;
  assign n51766 = n41745 & n51764 ;
  assign n51765 = ~n41745 & ~n51764 ;
  assign n51767 = ~\P1_P1_DataWidth_reg[1]/NET0131  & ~n51765 ;
  assign n51768 = ~n51766 & n51767 ;
  assign n51760 = \P1_P1_DataWidth_reg[1]/NET0131  & ~\P1_P1_rEIP_reg[22]/NET0131  ;
  assign n51769 = n8282 & ~n51760 ;
  assign n51770 = ~n51768 & n51769 ;
  assign n51771 = \P1_P1_rEIP_reg[22]/NET0131  & ~n50559 ;
  assign n51773 = ~\P1_P1_rEIP_reg[22]/NET0131  & ~n51737 ;
  assign n51774 = \P1_P1_rEIP_reg[22]/NET0131  & n51737 ;
  assign n51775 = ~n51773 & ~n51774 ;
  assign n51776 = n26275 & ~n51775 ;
  assign n51772 = ~\P1_P1_EBX_reg[22]/NET0131  & ~n26275 ;
  assign n51777 = n24502 & ~n51772 ;
  assign n51778 = ~n51776 & n51777 ;
  assign n51780 = ~\P1_P1_EBX_reg[21]/NET0131  & n51743 ;
  assign n51781 = \P1_P1_EBX_reg[31]/NET0131  & ~n51780 ;
  assign n51783 = ~\P1_P1_EBX_reg[22]/NET0131  & n51781 ;
  assign n51782 = \P1_P1_EBX_reg[22]/NET0131  & ~n51781 ;
  assign n51784 = ~n26274 & ~n51782 ;
  assign n51785 = ~n51783 & n51784 ;
  assign n51779 = n26274 & ~n51775 ;
  assign n51786 = n15334 & ~n51779 ;
  assign n51787 = ~n51785 & n51786 ;
  assign n51788 = ~n51778 & ~n51787 ;
  assign n51789 = ~n15364 & ~n51788 ;
  assign n51790 = ~n51771 & ~n51789 ;
  assign n51791 = n8355 & ~n51790 ;
  assign n51759 = \P1_P1_PhyAddrPointer_reg[22]/NET0131  & n8361 ;
  assign n51792 = \P1_P1_rEIP_reg[22]/NET0131  & ~n50583 ;
  assign n51793 = ~n51759 & ~n51792 ;
  assign n51794 = ~n51791 & n51793 ;
  assign n51795 = ~n51770 & n51794 ;
  assign n51798 = ~n36721 & ~n36733 ;
  assign n51799 = ~n51654 & ~n51798 ;
  assign n51801 = n39579 & n51799 ;
  assign n51800 = ~n39579 & ~n51799 ;
  assign n51802 = ~\P1_P1_DataWidth_reg[1]/NET0131  & ~n51800 ;
  assign n51803 = ~n51801 & n51802 ;
  assign n51797 = \P1_P1_DataWidth_reg[1]/NET0131  & ~\P1_P1_rEIP_reg[23]/NET0131  ;
  assign n51804 = n8282 & ~n51797 ;
  assign n51805 = ~n51803 & n51804 ;
  assign n51806 = \P1_P1_rEIP_reg[23]/NET0131  & ~n50559 ;
  assign n51811 = ~\P1_P1_EBX_reg[22]/NET0131  & n51780 ;
  assign n51812 = \P1_P1_EBX_reg[31]/NET0131  & ~n51811 ;
  assign n51814 = ~\P1_P1_EBX_reg[23]/NET0131  & n51812 ;
  assign n51813 = \P1_P1_EBX_reg[23]/NET0131  & ~n51812 ;
  assign n51815 = ~n26274 & ~n51813 ;
  assign n51816 = ~n51814 & n51815 ;
  assign n51807 = ~\P1_P1_rEIP_reg[23]/NET0131  & ~n51774 ;
  assign n51808 = \P1_P1_rEIP_reg[23]/NET0131  & n51774 ;
  assign n51809 = ~n51807 & ~n51808 ;
  assign n51810 = n26274 & ~n51809 ;
  assign n51817 = n15334 & ~n51810 ;
  assign n51818 = ~n51816 & n51817 ;
  assign n51820 = n26275 & ~n51809 ;
  assign n51819 = ~\P1_P1_EBX_reg[23]/NET0131  & ~n26275 ;
  assign n51821 = n24502 & ~n51819 ;
  assign n51822 = ~n51820 & n51821 ;
  assign n51823 = ~n51818 & ~n51822 ;
  assign n51824 = ~n15364 & ~n51823 ;
  assign n51825 = ~n51806 & ~n51824 ;
  assign n51826 = n8355 & ~n51825 ;
  assign n51796 = \P1_P1_PhyAddrPointer_reg[23]/NET0131  & n8361 ;
  assign n51827 = \P1_P1_rEIP_reg[23]/NET0131  & ~n50583 ;
  assign n51828 = ~n51796 & ~n51827 ;
  assign n51829 = ~n51826 & n51828 ;
  assign n51830 = ~n51805 & n51829 ;
  assign n51833 = n36722 & n51653 ;
  assign n51834 = ~n36733 & ~n51833 ;
  assign n51836 = n41772 & ~n51834 ;
  assign n51835 = ~n41772 & n51834 ;
  assign n51837 = ~\P1_P1_DataWidth_reg[1]/NET0131  & ~n51835 ;
  assign n51838 = ~n51836 & n51837 ;
  assign n51832 = \P1_P1_DataWidth_reg[1]/NET0131  & ~\P1_P1_rEIP_reg[24]/NET0131  ;
  assign n51839 = n8282 & ~n51832 ;
  assign n51840 = ~n51838 & n51839 ;
  assign n51841 = \P1_P1_rEIP_reg[24]/NET0131  & ~n50559 ;
  assign n51843 = ~\P1_P1_rEIP_reg[24]/NET0131  & ~n51808 ;
  assign n51844 = \P1_P1_rEIP_reg[22]/NET0131  & n51736 ;
  assign n51845 = \P1_P1_rEIP_reg[23]/NET0131  & n51844 ;
  assign n51846 = \P1_P1_rEIP_reg[24]/NET0131  & n51845 ;
  assign n51847 = n51677 & n51846 ;
  assign n51848 = ~n51843 & ~n51847 ;
  assign n51849 = n26275 & ~n51848 ;
  assign n51842 = ~\P1_P1_EBX_reg[24]/NET0131  & ~n26275 ;
  assign n51850 = n24502 & ~n51842 ;
  assign n51851 = ~n51849 & n51850 ;
  assign n51853 = ~\P1_P1_EBX_reg[23]/NET0131  & n51811 ;
  assign n51854 = \P1_P1_EBX_reg[31]/NET0131  & ~n51853 ;
  assign n51856 = ~\P1_P1_EBX_reg[24]/NET0131  & n51854 ;
  assign n51855 = \P1_P1_EBX_reg[24]/NET0131  & ~n51854 ;
  assign n51857 = ~n26274 & ~n51855 ;
  assign n51858 = ~n51856 & n51857 ;
  assign n51852 = n26274 & ~n51848 ;
  assign n51859 = n15334 & ~n51852 ;
  assign n51860 = ~n51858 & n51859 ;
  assign n51861 = ~n51851 & ~n51860 ;
  assign n51862 = ~n15364 & ~n51861 ;
  assign n51863 = ~n51841 & ~n51862 ;
  assign n51864 = n8355 & ~n51863 ;
  assign n51831 = \P1_P1_PhyAddrPointer_reg[24]/NET0131  & n8361 ;
  assign n51865 = \P1_P1_rEIP_reg[24]/NET0131  & ~n50583 ;
  assign n51866 = ~n51831 & ~n51865 ;
  assign n51867 = ~n51864 & n51866 ;
  assign n51868 = ~n51840 & n51867 ;
  assign n51893 = n36723 & n51653 ;
  assign n51894 = ~n36733 & ~n51893 ;
  assign n51895 = ~n43717 & ~n51894 ;
  assign n51896 = n43717 & n51894 ;
  assign n51897 = ~n51895 & ~n51896 ;
  assign n51898 = ~\P1_P1_DataWidth_reg[1]/NET0131  & ~n51897 ;
  assign n51892 = \P1_P1_DataWidth_reg[1]/NET0131  & ~\P1_P1_rEIP_reg[25]/NET0131  ;
  assign n51899 = n8282 & ~n51892 ;
  assign n51900 = ~n51898 & n51899 ;
  assign n51876 = ~\P1_P1_EBX_reg[24]/NET0131  & n51853 ;
  assign n51877 = \P1_P1_EBX_reg[31]/NET0131  & ~n51876 ;
  assign n51879 = ~\P1_P1_EBX_reg[25]/NET0131  & n51877 ;
  assign n51878 = \P1_P1_EBX_reg[25]/NET0131  & ~n51877 ;
  assign n51880 = ~n26274 & ~n51878 ;
  assign n51881 = ~n51879 & n51880 ;
  assign n51871 = ~\P1_P1_rEIP_reg[25]/NET0131  & ~n51847 ;
  assign n51872 = \P1_P1_rEIP_reg[24]/NET0131  & \P1_P1_rEIP_reg[25]/NET0131  ;
  assign n51873 = n51808 & n51872 ;
  assign n51874 = ~n51871 & ~n51873 ;
  assign n51875 = n26274 & ~n51874 ;
  assign n51882 = n24504 & ~n51875 ;
  assign n51883 = ~n51881 & n51882 ;
  assign n51870 = \P1_P1_rEIP_reg[25]/NET0131  & ~n50559 ;
  assign n51885 = n26275 & ~n51874 ;
  assign n51884 = ~\P1_P1_EBX_reg[25]/NET0131  & ~n26275 ;
  assign n51886 = n24503 & ~n51884 ;
  assign n51887 = ~n51885 & n51886 ;
  assign n51888 = ~n51870 & ~n51887 ;
  assign n51889 = ~n51883 & n51888 ;
  assign n51890 = n8355 & ~n51889 ;
  assign n51869 = \P1_P1_PhyAddrPointer_reg[25]/NET0131  & n8361 ;
  assign n51891 = \P1_P1_rEIP_reg[25]/NET0131  & ~n50583 ;
  assign n51901 = ~n51869 & ~n51891 ;
  assign n51902 = ~n51890 & n51901 ;
  assign n51903 = ~n51900 & n51902 ;
  assign n51906 = \P1_P1_PhyAddrPointer_reg[25]/NET0131  & n51893 ;
  assign n51907 = ~n36733 & ~n51906 ;
  assign n51909 = n41790 & ~n51907 ;
  assign n51908 = ~n41790 & n51907 ;
  assign n51910 = ~\P1_P1_DataWidth_reg[1]/NET0131  & ~n51908 ;
  assign n51911 = ~n51909 & n51910 ;
  assign n51905 = \P1_P1_DataWidth_reg[1]/NET0131  & ~\P1_P1_rEIP_reg[26]/NET0131  ;
  assign n51912 = n8282 & ~n51905 ;
  assign n51913 = ~n51911 & n51912 ;
  assign n51919 = ~\P1_P1_EBX_reg[25]/NET0131  & n51876 ;
  assign n51920 = \P1_P1_EBX_reg[31]/NET0131  & ~n51919 ;
  assign n51922 = ~\P1_P1_EBX_reg[26]/NET0131  & n51920 ;
  assign n51921 = \P1_P1_EBX_reg[26]/NET0131  & ~n51920 ;
  assign n51923 = ~n26274 & ~n51921 ;
  assign n51924 = ~n51922 & n51923 ;
  assign n51915 = ~\P1_P1_rEIP_reg[26]/NET0131  & ~n51873 ;
  assign n51916 = \P1_P1_rEIP_reg[26]/NET0131  & n51873 ;
  assign n51917 = ~n51915 & ~n51916 ;
  assign n51918 = n26274 & ~n51917 ;
  assign n51925 = n24504 & ~n51918 ;
  assign n51926 = ~n51924 & n51925 ;
  assign n51914 = \P1_P1_rEIP_reg[26]/NET0131  & ~n50559 ;
  assign n51928 = n26275 & ~n51917 ;
  assign n51927 = ~\P1_P1_EBX_reg[26]/NET0131  & ~n26275 ;
  assign n51929 = n24503 & ~n51927 ;
  assign n51930 = ~n51928 & n51929 ;
  assign n51931 = ~n51914 & ~n51930 ;
  assign n51932 = ~n51926 & n51931 ;
  assign n51933 = n8355 & ~n51932 ;
  assign n51904 = \P1_P1_PhyAddrPointer_reg[26]/NET0131  & n8361 ;
  assign n51934 = \P1_P1_rEIP_reg[26]/NET0131  & ~n50583 ;
  assign n51935 = ~n51904 & ~n51934 ;
  assign n51936 = ~n51933 & n51935 ;
  assign n51937 = ~n51913 & n51936 ;
  assign n51940 = ~n36733 & ~n39602 ;
  assign n51941 = ~n51894 & ~n51940 ;
  assign n51943 = n39604 & n51941 ;
  assign n51942 = ~n39604 & ~n51941 ;
  assign n51944 = ~\P1_P1_DataWidth_reg[1]/NET0131  & ~n51942 ;
  assign n51945 = ~n51943 & n51944 ;
  assign n51939 = \P1_P1_DataWidth_reg[1]/NET0131  & ~\P1_P1_rEIP_reg[27]/NET0131  ;
  assign n51946 = n8282 & ~n51939 ;
  assign n51947 = ~n51945 & n51946 ;
  assign n51955 = ~\P1_P1_EBX_reg[26]/NET0131  & n51919 ;
  assign n51956 = \P1_P1_EBX_reg[31]/NET0131  & ~n51955 ;
  assign n51958 = ~\P1_P1_EBX_reg[27]/NET0131  & n51956 ;
  assign n51957 = \P1_P1_EBX_reg[27]/NET0131  & ~n51956 ;
  assign n51959 = ~n26274 & ~n51957 ;
  assign n51960 = ~n51958 & n51959 ;
  assign n51949 = ~\P1_P1_rEIP_reg[27]/NET0131  & ~n51916 ;
  assign n51950 = \P1_P1_rEIP_reg[26]/NET0131  & n51872 ;
  assign n51951 = \P1_P1_rEIP_reg[27]/NET0131  & n51950 ;
  assign n51952 = n51808 & n51951 ;
  assign n51953 = ~n51949 & ~n51952 ;
  assign n51954 = n26274 & ~n51953 ;
  assign n51961 = n24504 & ~n51954 ;
  assign n51962 = ~n51960 & n51961 ;
  assign n51948 = \P1_P1_rEIP_reg[27]/NET0131  & ~n50559 ;
  assign n51964 = n26275 & ~n51953 ;
  assign n51963 = ~\P1_P1_EBX_reg[27]/NET0131  & ~n26275 ;
  assign n51965 = n24503 & ~n51963 ;
  assign n51966 = ~n51964 & n51965 ;
  assign n51967 = ~n51948 & ~n51966 ;
  assign n51968 = ~n51962 & n51967 ;
  assign n51969 = n8355 & ~n51968 ;
  assign n51938 = \P1_P1_PhyAddrPointer_reg[27]/NET0131  & n8361 ;
  assign n51970 = \P1_P1_rEIP_reg[27]/NET0131  & ~n50583 ;
  assign n51971 = ~n51938 & ~n51970 ;
  assign n51972 = ~n51969 & n51971 ;
  assign n51973 = ~n51947 & n51972 ;
  assign n51976 = ~n36727 & ~n36733 ;
  assign n51977 = ~n51894 & ~n51976 ;
  assign n51979 = n39622 & n51977 ;
  assign n51978 = ~n39622 & ~n51977 ;
  assign n51980 = ~\P1_P1_DataWidth_reg[1]/NET0131  & ~n51978 ;
  assign n51981 = ~n51979 & n51980 ;
  assign n51975 = \P1_P1_DataWidth_reg[1]/NET0131  & ~\P1_P1_rEIP_reg[28]/NET0131  ;
  assign n51982 = n8282 & ~n51975 ;
  assign n51983 = ~n51981 & n51982 ;
  assign n51993 = ~\P1_P1_EBX_reg[27]/NET0131  & n51955 ;
  assign n51994 = \P1_P1_EBX_reg[31]/NET0131  & ~n51993 ;
  assign n51996 = ~\P1_P1_EBX_reg[28]/NET0131  & n51994 ;
  assign n51995 = \P1_P1_EBX_reg[28]/NET0131  & ~n51994 ;
  assign n51997 = ~n26274 & ~n51995 ;
  assign n51998 = ~n51996 & n51997 ;
  assign n51986 = \P1_P1_rEIP_reg[28]/NET0131  & n51952 ;
  assign n51987 = ~\P1_P1_rEIP_reg[28]/NET0131  & ~n51952 ;
  assign n51988 = ~n51986 & ~n51987 ;
  assign n51989 = n26274 & ~n51988 ;
  assign n51999 = n24504 & ~n51989 ;
  assign n52000 = ~n51998 & n51999 ;
  assign n51984 = \P1_P1_rEIP_reg[28]/NET0131  & ~n50559 ;
  assign n51990 = ~n26158 & n51989 ;
  assign n51985 = ~\P1_P1_EBX_reg[28]/NET0131  & ~n26275 ;
  assign n51991 = n24503 & ~n51985 ;
  assign n51992 = ~n51990 & n51991 ;
  assign n52001 = ~n51984 & ~n51992 ;
  assign n52002 = ~n52000 & n52001 ;
  assign n52003 = n8355 & ~n52002 ;
  assign n51974 = \P1_P1_PhyAddrPointer_reg[28]/NET0131  & n8361 ;
  assign n52004 = \P1_P1_rEIP_reg[28]/NET0131  & ~n50583 ;
  assign n52005 = ~n51974 & ~n52004 ;
  assign n52006 = ~n52003 & n52005 ;
  assign n52007 = ~n51983 & n52006 ;
  assign n52010 = ~n36728 & ~n36733 ;
  assign n52011 = ~n51894 & ~n52010 ;
  assign n52013 = ~n39640 & ~n52011 ;
  assign n52012 = n39640 & n52011 ;
  assign n52014 = ~\P1_P1_DataWidth_reg[1]/NET0131  & ~n52012 ;
  assign n52015 = ~n52013 & n52014 ;
  assign n52009 = \P1_P1_DataWidth_reg[1]/NET0131  & ~\P1_P1_rEIP_reg[29]/NET0131  ;
  assign n52016 = n8282 & ~n52009 ;
  assign n52017 = ~n52015 & n52016 ;
  assign n52025 = ~\P1_P1_EBX_reg[28]/NET0131  & n51993 ;
  assign n52026 = \P1_P1_EBX_reg[31]/NET0131  & ~n52025 ;
  assign n52028 = \P1_P1_EBX_reg[29]/NET0131  & ~n52026 ;
  assign n52027 = ~\P1_P1_EBX_reg[29]/NET0131  & n52026 ;
  assign n52029 = ~n26274 & ~n52027 ;
  assign n52030 = ~n52028 & n52029 ;
  assign n52019 = ~\P1_P1_rEIP_reg[29]/NET0131  & ~n51986 ;
  assign n52020 = \P1_P1_rEIP_reg[27]/NET0131  & \P1_P1_rEIP_reg[28]/NET0131  ;
  assign n52021 = \P1_P1_rEIP_reg[29]/NET0131  & n52020 ;
  assign n52022 = n51916 & n52021 ;
  assign n52023 = ~n52019 & ~n52022 ;
  assign n52024 = n26274 & ~n52023 ;
  assign n52031 = n24504 & ~n52024 ;
  assign n52032 = ~n52030 & n52031 ;
  assign n52018 = \P1_P1_rEIP_reg[29]/NET0131  & ~n50559 ;
  assign n52034 = n26275 & ~n52023 ;
  assign n52033 = ~\P1_P1_EBX_reg[29]/NET0131  & ~n26275 ;
  assign n52035 = n24503 & ~n52033 ;
  assign n52036 = ~n52034 & n52035 ;
  assign n52037 = ~n52018 & ~n52036 ;
  assign n52038 = ~n52032 & n52037 ;
  assign n52039 = n8355 & ~n52038 ;
  assign n52008 = \P1_P1_PhyAddrPointer_reg[29]/NET0131  & n8361 ;
  assign n52040 = \P1_P1_rEIP_reg[29]/NET0131  & ~n50583 ;
  assign n52041 = ~n52008 & ~n52040 ;
  assign n52042 = ~n52039 & n52041 ;
  assign n52043 = ~n52017 & n52042 ;
  assign n52046 = ~\P1_P1_PhyAddrPointer_reg[0]/NET0131  & \P1_P1_PhyAddrPointer_reg[1]/NET0131  ;
  assign n52047 = ~n36733 & ~n52046 ;
  assign n52048 = ~\P1_P1_PhyAddrPointer_reg[1]/NET0131  & ~\P1_P1_PhyAddrPointer_reg[2]/NET0131  ;
  assign n52049 = ~n47430 & ~n52048 ;
  assign n52051 = ~n52047 & n52049 ;
  assign n52050 = n52047 & ~n52049 ;
  assign n52052 = ~\P1_P1_DataWidth_reg[1]/NET0131  & ~n52050 ;
  assign n52053 = ~n52051 & n52052 ;
  assign n52045 = \P1_P1_DataWidth_reg[1]/NET0131  & ~\P1_P1_rEIP_reg[2]/NET0131  ;
  assign n52054 = n8282 & ~n52045 ;
  assign n52055 = ~n52053 & n52054 ;
  assign n52056 = \P1_P1_rEIP_reg[2]/NET0131  & ~n50559 ;
  assign n52069 = \P1_P1_EBX_reg[2]/NET0131  & ~n26275 ;
  assign n52058 = ~\P1_P1_rEIP_reg[1]/NET0131  & ~\P1_P1_rEIP_reg[2]/NET0131  ;
  assign n52059 = ~\P1_P1_DataWidth_reg[1]/NET0131  & ~n50600 ;
  assign n52060 = ~n52058 & n52059 ;
  assign n52070 = n26264 & n52060 ;
  assign n52071 = ~n52069 & ~n52070 ;
  assign n52072 = n24502 & ~n52071 ;
  assign n52057 = n15382 & n26119 ;
  assign n52061 = ~n15335 & n52060 ;
  assign n52062 = \P1_P1_EBX_reg[31]/NET0131  & ~n50562 ;
  assign n52064 = \P1_P1_EBX_reg[2]/NET0131  & n52062 ;
  assign n52063 = ~\P1_P1_EBX_reg[2]/NET0131  & ~n52062 ;
  assign n52065 = ~n26274 & ~n52063 ;
  assign n52066 = ~n52064 & n52065 ;
  assign n52067 = ~n52061 & ~n52066 ;
  assign n52068 = n15334 & ~n52067 ;
  assign n52073 = ~n52057 & ~n52068 ;
  assign n52074 = ~n52072 & n52073 ;
  assign n52075 = ~n15364 & ~n52074 ;
  assign n52076 = ~n52056 & ~n52075 ;
  assign n52077 = n8355 & ~n52076 ;
  assign n52044 = \P1_P1_PhyAddrPointer_reg[2]/NET0131  & n8361 ;
  assign n52078 = \P1_P1_rEIP_reg[2]/NET0131  & ~n50583 ;
  assign n52079 = ~n52044 & ~n52078 ;
  assign n52080 = ~n52077 & n52079 ;
  assign n52081 = ~n52055 & n52080 ;
  assign n52084 = ~\P2_P2_PhyAddrPointer_reg[0]/NET0131  & n39648 ;
  assign n52085 = \P2_P2_PhyAddrPointer_reg[14]/NET0131  & n52084 ;
  assign n52086 = n36777 & n52085 ;
  assign n52087 = n36792 & ~n52086 ;
  assign n52089 = n41870 & ~n52087 ;
  assign n52088 = ~n41870 & n52087 ;
  assign n52090 = ~\P2_P2_DataWidth_reg[1]/NET0131  & ~n52088 ;
  assign n52091 = ~n52089 & n52090 ;
  assign n52083 = \P2_P2_DataWidth_reg[1]/NET0131  & ~\P2_P2_rEIP_reg[20]/NET0131  ;
  assign n52092 = n26794 & ~n52083 ;
  assign n52093 = ~n52091 & n52092 ;
  assign n52115 = ~\P2_P2_EBX_reg[3]/NET0131  & n50678 ;
  assign n52116 = ~\P2_P2_EBX_reg[4]/NET0131  & n52115 ;
  assign n52117 = ~\P2_P2_EBX_reg[5]/NET0131  & n52116 ;
  assign n52118 = ~\P2_P2_EBX_reg[6]/NET0131  & n52117 ;
  assign n52119 = ~\P2_P2_EBX_reg[7]/NET0131  & n52118 ;
  assign n52120 = ~\P2_P2_EBX_reg[8]/NET0131  & n52119 ;
  assign n52121 = ~\P2_P2_EBX_reg[9]/NET0131  & n52120 ;
  assign n52122 = ~\P2_P2_EBX_reg[10]/NET0131  & n52121 ;
  assign n52123 = ~\P2_P2_EBX_reg[11]/NET0131  & n52122 ;
  assign n52124 = ~\P2_P2_EBX_reg[12]/NET0131  & n52123 ;
  assign n52125 = ~\P2_P2_EBX_reg[13]/NET0131  & n52124 ;
  assign n52126 = ~\P2_P2_EBX_reg[14]/NET0131  & n52125 ;
  assign n52127 = ~\P2_P2_EBX_reg[15]/NET0131  & n52126 ;
  assign n52128 = ~\P2_P2_EBX_reg[16]/NET0131  & n52127 ;
  assign n52129 = ~\P2_P2_EBX_reg[17]/NET0131  & n52128 ;
  assign n52130 = ~\P2_P2_EBX_reg[18]/NET0131  & n52129 ;
  assign n52131 = ~\P2_P2_EBX_reg[19]/NET0131  & n52130 ;
  assign n52132 = \P2_P2_EBX_reg[31]/NET0131  & ~n52131 ;
  assign n52134 = ~\P2_P2_EBX_reg[20]/NET0131  & n52132 ;
  assign n52133 = \P2_P2_EBX_reg[20]/NET0131  & ~n52132 ;
  assign n52135 = ~n50649 & ~n52133 ;
  assign n52136 = ~n52134 & n52135 ;
  assign n52095 = \P2_P2_rEIP_reg[4]/NET0131  & n50685 ;
  assign n52096 = \P2_P2_rEIP_reg[5]/NET0131  & n52095 ;
  assign n52097 = \P2_P2_rEIP_reg[6]/NET0131  & n52096 ;
  assign n52098 = \P2_P2_rEIP_reg[7]/NET0131  & n52097 ;
  assign n52099 = \P2_P2_rEIP_reg[8]/NET0131  & n52098 ;
  assign n52100 = \P2_P2_rEIP_reg[15]/NET0131  & \P2_P2_rEIP_reg[16]/NET0131  ;
  assign n52101 = \P2_P2_rEIP_reg[17]/NET0131  & n52100 ;
  assign n52102 = \P2_P2_rEIP_reg[18]/NET0131  & \P2_P2_rEIP_reg[19]/NET0131  ;
  assign n52103 = n52101 & n52102 ;
  assign n52105 = \P2_P2_rEIP_reg[10]/NET0131  & \P2_P2_rEIP_reg[11]/NET0131  ;
  assign n52104 = \P2_P2_rEIP_reg[12]/NET0131  & \P2_P2_rEIP_reg[13]/NET0131  ;
  assign n52106 = \P2_P2_rEIP_reg[14]/NET0131  & \P2_P2_rEIP_reg[9]/NET0131  ;
  assign n52107 = n52104 & n52106 ;
  assign n52108 = n52105 & n52107 ;
  assign n52109 = n52103 & n52108 ;
  assign n52110 = n52099 & n52109 ;
  assign n52111 = ~\P2_P2_rEIP_reg[20]/NET0131  & ~n52110 ;
  assign n52112 = \P2_P2_rEIP_reg[20]/NET0131  & n52110 ;
  assign n52113 = ~n52111 & ~n52112 ;
  assign n52114 = n50649 & ~n52113 ;
  assign n52137 = n47684 & ~n52114 ;
  assign n52138 = ~n52136 & n52137 ;
  assign n52094 = \P2_P2_rEIP_reg[20]/NET0131  & ~n50640 ;
  assign n52139 = ~\P2_P2_EBX_reg[20]/NET0131  & ~n50642 ;
  assign n52140 = n50642 & ~n52113 ;
  assign n52141 = ~n52139 & ~n52140 ;
  assign n52142 = n26786 & n52141 ;
  assign n52143 = ~n52094 & ~n52142 ;
  assign n52144 = ~n52138 & n52143 ;
  assign n52145 = n26792 & ~n52144 ;
  assign n52082 = \P2_P2_PhyAddrPointer_reg[20]/NET0131  & n27637 ;
  assign n52146 = \P2_P2_rEIP_reg[20]/NET0131  & ~n50636 ;
  assign n52147 = ~n52082 & ~n52146 ;
  assign n52148 = ~n52145 & n52147 ;
  assign n52149 = ~n52093 & n52148 ;
  assign n52152 = ~\P2_P2_PhyAddrPointer_reg[0]/NET0131  & n47452 ;
  assign n52153 = n36772 & n52152 ;
  assign n52154 = n36778 & n52153 ;
  assign n52155 = n36792 & ~n52154 ;
  assign n52157 = n43850 & ~n52155 ;
  assign n52156 = ~n43850 & n52155 ;
  assign n52158 = ~\P2_P2_DataWidth_reg[1]/NET0131  & ~n52156 ;
  assign n52159 = ~n52157 & n52158 ;
  assign n52151 = \P2_P2_DataWidth_reg[1]/NET0131  & ~\P2_P2_rEIP_reg[21]/NET0131  ;
  assign n52160 = n26794 & ~n52151 ;
  assign n52161 = ~n52159 & n52160 ;
  assign n52168 = ~\P2_P2_EBX_reg[20]/NET0131  & n52131 ;
  assign n52169 = \P2_P2_EBX_reg[31]/NET0131  & ~n52168 ;
  assign n52171 = ~\P2_P2_EBX_reg[21]/NET0131  & n52169 ;
  assign n52170 = \P2_P2_EBX_reg[21]/NET0131  & ~n52169 ;
  assign n52172 = ~n50649 & ~n52170 ;
  assign n52173 = ~n52171 & n52172 ;
  assign n52163 = ~\P2_P2_rEIP_reg[21]/NET0131  & ~n52112 ;
  assign n52164 = \P2_P2_rEIP_reg[20]/NET0131  & \P2_P2_rEIP_reg[21]/NET0131  ;
  assign n52165 = n52110 & n52164 ;
  assign n52166 = ~n52163 & ~n52165 ;
  assign n52167 = n50649 & ~n52166 ;
  assign n52174 = n47684 & ~n52167 ;
  assign n52175 = ~n52173 & n52174 ;
  assign n52162 = \P2_P2_rEIP_reg[21]/NET0131  & ~n50640 ;
  assign n52177 = n50642 & ~n52166 ;
  assign n52176 = ~\P2_P2_EBX_reg[21]/NET0131  & ~n50642 ;
  assign n52178 = n26786 & ~n52176 ;
  assign n52179 = ~n52177 & n52178 ;
  assign n52180 = ~n52162 & ~n52179 ;
  assign n52181 = ~n52175 & n52180 ;
  assign n52182 = n26792 & ~n52181 ;
  assign n52150 = \P2_P2_PhyAddrPointer_reg[21]/NET0131  & n27637 ;
  assign n52183 = \P2_P2_rEIP_reg[21]/NET0131  & ~n50636 ;
  assign n52184 = ~n52150 & ~n52183 ;
  assign n52185 = ~n52182 & n52184 ;
  assign n52186 = ~n52161 & n52185 ;
  assign n52189 = n36779 & n52085 ;
  assign n52190 = n36792 & ~n52189 ;
  assign n52192 = ~n41900 & n52190 ;
  assign n52191 = n41900 & ~n52190 ;
  assign n52193 = ~\P2_P2_DataWidth_reg[1]/NET0131  & ~n52191 ;
  assign n52194 = ~n52192 & n52193 ;
  assign n52188 = \P2_P2_DataWidth_reg[1]/NET0131  & ~\P2_P2_rEIP_reg[22]/NET0131  ;
  assign n52195 = n26794 & ~n52188 ;
  assign n52196 = ~n52194 & n52195 ;
  assign n52202 = ~\P2_P2_EBX_reg[21]/NET0131  & n52168 ;
  assign n52203 = \P2_P2_EBX_reg[31]/NET0131  & ~n52202 ;
  assign n52205 = ~\P2_P2_EBX_reg[22]/NET0131  & n52203 ;
  assign n52204 = \P2_P2_EBX_reg[22]/NET0131  & ~n52203 ;
  assign n52206 = ~n50649 & ~n52204 ;
  assign n52207 = ~n52205 & n52206 ;
  assign n52198 = \P2_P2_rEIP_reg[22]/NET0131  & n52165 ;
  assign n52199 = ~\P2_P2_rEIP_reg[22]/NET0131  & ~n52165 ;
  assign n52200 = ~n52198 & ~n52199 ;
  assign n52201 = n50649 & ~n52200 ;
  assign n52208 = n47684 & ~n52201 ;
  assign n52209 = ~n52207 & n52208 ;
  assign n52197 = \P2_P2_rEIP_reg[22]/NET0131  & ~n50640 ;
  assign n52211 = n50642 & ~n52200 ;
  assign n52210 = ~\P2_P2_EBX_reg[22]/NET0131  & ~n50642 ;
  assign n52212 = n26786 & ~n52210 ;
  assign n52213 = ~n52211 & n52212 ;
  assign n52214 = ~n52197 & ~n52213 ;
  assign n52215 = ~n52209 & n52214 ;
  assign n52216 = n26792 & ~n52215 ;
  assign n52187 = \P2_P2_PhyAddrPointer_reg[22]/NET0131  & n27637 ;
  assign n52217 = \P2_P2_rEIP_reg[22]/NET0131  & ~n50636 ;
  assign n52218 = ~n52187 & ~n52217 ;
  assign n52219 = ~n52216 & n52218 ;
  assign n52220 = ~n52196 & n52219 ;
  assign n52223 = \P2_P2_PhyAddrPointer_reg[22]/NET0131  & n52189 ;
  assign n52224 = n36792 & ~n52223 ;
  assign n52226 = n39685 & ~n52224 ;
  assign n52225 = ~n39685 & n52224 ;
  assign n52227 = ~\P2_P2_DataWidth_reg[1]/NET0131  & ~n52225 ;
  assign n52228 = ~n52226 & n52227 ;
  assign n52222 = \P2_P2_DataWidth_reg[1]/NET0131  & ~\P2_P2_rEIP_reg[23]/NET0131  ;
  assign n52229 = n26794 & ~n52222 ;
  assign n52230 = ~n52228 & n52229 ;
  assign n52231 = \P2_P2_rEIP_reg[23]/NET0131  & ~n50640 ;
  assign n52233 = ~\P2_P2_rEIP_reg[23]/NET0131  & ~n52198 ;
  assign n52234 = \P2_P2_rEIP_reg[23]/NET0131  & n52198 ;
  assign n52235 = ~n52233 & ~n52234 ;
  assign n52236 = n50642 & ~n52235 ;
  assign n52232 = ~\P2_P2_EBX_reg[23]/NET0131  & ~n50642 ;
  assign n52237 = n26643 & ~n52232 ;
  assign n52238 = ~n52236 & n52237 ;
  assign n52240 = ~\P2_P2_EBX_reg[22]/NET0131  & n52202 ;
  assign n52241 = \P2_P2_EBX_reg[31]/NET0131  & ~n52240 ;
  assign n52243 = \P2_P2_EBX_reg[23]/NET0131  & ~n52241 ;
  assign n52242 = ~\P2_P2_EBX_reg[23]/NET0131  & n52241 ;
  assign n52244 = ~n50649 & ~n52242 ;
  assign n52245 = ~n52243 & n52244 ;
  assign n52239 = n50649 & ~n52235 ;
  assign n52246 = n26633 & ~n52239 ;
  assign n52247 = ~n52245 & n52246 ;
  assign n52248 = ~n52238 & ~n52247 ;
  assign n52249 = ~n26640 & ~n52248 ;
  assign n52250 = ~n52231 & ~n52249 ;
  assign n52251 = n26792 & ~n52250 ;
  assign n52221 = \P2_P2_PhyAddrPointer_reg[23]/NET0131  & n27637 ;
  assign n52252 = \P2_P2_rEIP_reg[23]/NET0131  & ~n50636 ;
  assign n52253 = ~n52221 & ~n52252 ;
  assign n52254 = ~n52251 & n52253 ;
  assign n52255 = ~n52230 & n52254 ;
  assign n52258 = \P2_P2_PhyAddrPointer_reg[23]/NET0131  & n52223 ;
  assign n52259 = n36792 & ~n52258 ;
  assign n52261 = n41917 & ~n52259 ;
  assign n52260 = ~n41917 & n52259 ;
  assign n52262 = ~\P2_P2_DataWidth_reg[1]/NET0131  & ~n52260 ;
  assign n52263 = ~n52261 & n52262 ;
  assign n52257 = \P2_P2_DataWidth_reg[1]/NET0131  & ~\P2_P2_rEIP_reg[24]/NET0131  ;
  assign n52264 = n26794 & ~n52257 ;
  assign n52265 = ~n52263 & n52264 ;
  assign n52266 = \P2_P2_rEIP_reg[24]/NET0131  & ~n50640 ;
  assign n52268 = ~\P2_P2_rEIP_reg[24]/NET0131  & ~n52234 ;
  assign n52269 = \P2_P2_rEIP_reg[22]/NET0131  & \P2_P2_rEIP_reg[23]/NET0131  ;
  assign n52270 = \P2_P2_rEIP_reg[24]/NET0131  & n52269 ;
  assign n52271 = n52165 & n52270 ;
  assign n52272 = ~n52268 & ~n52271 ;
  assign n52273 = n50642 & ~n52272 ;
  assign n52267 = ~\P2_P2_EBX_reg[24]/NET0131  & ~n50642 ;
  assign n52274 = n26643 & ~n52267 ;
  assign n52275 = ~n52273 & n52274 ;
  assign n52277 = ~\P2_P2_EBX_reg[23]/NET0131  & n52240 ;
  assign n52278 = \P2_P2_EBX_reg[31]/NET0131  & ~n52277 ;
  assign n52280 = \P2_P2_EBX_reg[24]/NET0131  & ~n52278 ;
  assign n52279 = ~\P2_P2_EBX_reg[24]/NET0131  & n52278 ;
  assign n52281 = ~n50649 & ~n52279 ;
  assign n52282 = ~n52280 & n52281 ;
  assign n52276 = n50649 & ~n52272 ;
  assign n52283 = n26633 & ~n52276 ;
  assign n52284 = ~n52282 & n52283 ;
  assign n52285 = ~n52275 & ~n52284 ;
  assign n52286 = ~n26640 & ~n52285 ;
  assign n52287 = ~n52266 & ~n52286 ;
  assign n52288 = n26792 & ~n52287 ;
  assign n52256 = \P2_P2_PhyAddrPointer_reg[24]/NET0131  & n27637 ;
  assign n52289 = \P2_P2_rEIP_reg[24]/NET0131  & ~n50636 ;
  assign n52290 = ~n52256 & ~n52289 ;
  assign n52291 = ~n52288 & n52290 ;
  assign n52292 = ~n52265 & n52291 ;
  assign n52295 = n36782 & n52153 ;
  assign n52296 = n36792 & ~n52295 ;
  assign n52298 = n43868 & ~n52296 ;
  assign n52297 = ~n43868 & n52296 ;
  assign n52299 = ~\P2_P2_DataWidth_reg[1]/NET0131  & ~n52297 ;
  assign n52300 = ~n52298 & n52299 ;
  assign n52294 = \P2_P2_DataWidth_reg[1]/NET0131  & ~\P2_P2_rEIP_reg[25]/NET0131  ;
  assign n52301 = n26794 & ~n52294 ;
  assign n52302 = ~n52300 & n52301 ;
  assign n52303 = \P2_P2_rEIP_reg[25]/NET0131  & ~n50640 ;
  assign n52305 = n52109 & n52164 ;
  assign n52306 = n52270 & n52305 ;
  assign n52307 = \P2_P2_rEIP_reg[25]/NET0131  & n52306 ;
  assign n52308 = n52099 & n52307 ;
  assign n52309 = ~\P2_P2_rEIP_reg[25]/NET0131  & ~n52271 ;
  assign n52310 = ~n52308 & ~n52309 ;
  assign n52311 = n50642 & ~n52310 ;
  assign n52304 = ~\P2_P2_EBX_reg[25]/NET0131  & ~n50642 ;
  assign n52312 = n26643 & ~n52304 ;
  assign n52313 = ~n52311 & n52312 ;
  assign n52315 = ~\P2_P2_EBX_reg[24]/NET0131  & n52277 ;
  assign n52316 = \P2_P2_EBX_reg[31]/NET0131  & ~n52315 ;
  assign n52318 = \P2_P2_EBX_reg[25]/NET0131  & ~n52316 ;
  assign n52317 = ~\P2_P2_EBX_reg[25]/NET0131  & n52316 ;
  assign n52319 = ~n50649 & ~n52317 ;
  assign n52320 = ~n52318 & n52319 ;
  assign n52314 = n50649 & ~n52310 ;
  assign n52321 = n26633 & ~n52314 ;
  assign n52322 = ~n52320 & n52321 ;
  assign n52323 = ~n52313 & ~n52322 ;
  assign n52324 = ~n26640 & ~n52323 ;
  assign n52325 = ~n52303 & ~n52324 ;
  assign n52326 = n26792 & ~n52325 ;
  assign n52293 = \P2_P2_PhyAddrPointer_reg[25]/NET0131  & n27637 ;
  assign n52327 = \P2_P2_rEIP_reg[25]/NET0131  & ~n50636 ;
  assign n52328 = ~n52293 & ~n52327 ;
  assign n52329 = ~n52326 & n52328 ;
  assign n52330 = ~n52302 & n52329 ;
  assign n52333 = n36783 & n52085 ;
  assign n52334 = n36792 & ~n52333 ;
  assign n52336 = ~n41935 & n52334 ;
  assign n52335 = n41935 & ~n52334 ;
  assign n52337 = ~\P2_P2_DataWidth_reg[1]/NET0131  & ~n52335 ;
  assign n52338 = ~n52336 & n52337 ;
  assign n52332 = \P2_P2_DataWidth_reg[1]/NET0131  & ~\P2_P2_rEIP_reg[26]/NET0131  ;
  assign n52339 = n26794 & ~n52332 ;
  assign n52340 = ~n52338 & n52339 ;
  assign n52341 = ~\P2_P2_EBX_reg[26]/NET0131  & ~n50642 ;
  assign n52342 = ~\P2_P2_rEIP_reg[26]/NET0131  & ~n52308 ;
  assign n52343 = \P2_P2_rEIP_reg[26]/NET0131  & n52308 ;
  assign n52344 = ~n52342 & ~n52343 ;
  assign n52345 = n50649 & ~n52344 ;
  assign n52346 = ~n26650 & n52345 ;
  assign n52347 = ~n52341 & ~n52346 ;
  assign n52348 = ~n26640 & ~n52347 ;
  assign n52349 = n26643 & ~n52348 ;
  assign n52350 = ~n26633 & ~n26637 ;
  assign n52351 = ~n26680 & n52350 ;
  assign n52352 = ~n50640 & ~n52351 ;
  assign n52353 = ~n52349 & ~n52352 ;
  assign n52354 = \P2_P2_rEIP_reg[26]/NET0131  & ~n52353 ;
  assign n52355 = ~\P2_P2_EBX_reg[25]/NET0131  & n52315 ;
  assign n52356 = \P2_P2_EBX_reg[31]/NET0131  & ~n52355 ;
  assign n52358 = \P2_P2_EBX_reg[26]/NET0131  & ~n52356 ;
  assign n52357 = ~\P2_P2_EBX_reg[26]/NET0131  & n52356 ;
  assign n52359 = ~n50649 & ~n52357 ;
  assign n52360 = ~n52358 & n52359 ;
  assign n52361 = n26633 & ~n52345 ;
  assign n52362 = ~n52360 & n52361 ;
  assign n52363 = ~n52349 & ~n52362 ;
  assign n52364 = ~n26640 & ~n52363 ;
  assign n52365 = ~n52354 & ~n52364 ;
  assign n52366 = n26792 & ~n52365 ;
  assign n52331 = \P2_P2_PhyAddrPointer_reg[26]/NET0131  & n27637 ;
  assign n52367 = \P2_P2_rEIP_reg[26]/NET0131  & ~n50636 ;
  assign n52368 = ~n52331 & ~n52367 ;
  assign n52369 = ~n52366 & n52368 ;
  assign n52370 = ~n52340 & n52369 ;
  assign n52381 = ~\P2_P2_EBX_reg[27]/NET0131  & ~n50642 ;
  assign n52382 = \P2_P2_rEIP_reg[27]/NET0131  & n52343 ;
  assign n52383 = ~\P2_P2_rEIP_reg[27]/NET0131  & ~n52343 ;
  assign n52384 = ~n52382 & ~n52383 ;
  assign n52385 = n50649 & ~n52384 ;
  assign n52386 = ~n26650 & n52385 ;
  assign n52387 = ~n52381 & ~n52386 ;
  assign n52388 = ~n26640 & ~n52387 ;
  assign n52389 = n26643 & ~n52388 ;
  assign n52390 = ~n52352 & ~n52389 ;
  assign n52391 = \P2_P2_rEIP_reg[27]/NET0131  & ~n52390 ;
  assign n52392 = ~\P2_P2_EBX_reg[26]/NET0131  & n52355 ;
  assign n52393 = \P2_P2_EBX_reg[31]/NET0131  & ~n52392 ;
  assign n52395 = \P2_P2_EBX_reg[27]/NET0131  & ~n52393 ;
  assign n52394 = ~\P2_P2_EBX_reg[27]/NET0131  & n52393 ;
  assign n52396 = ~n50649 & ~n52394 ;
  assign n52397 = ~n52395 & n52396 ;
  assign n52398 = n26633 & ~n52385 ;
  assign n52399 = ~n52397 & n52398 ;
  assign n52400 = ~n52389 & ~n52399 ;
  assign n52401 = ~n26640 & ~n52400 ;
  assign n52402 = ~n52391 & ~n52401 ;
  assign n52403 = n26792 & ~n52402 ;
  assign n52373 = \P2_P2_PhyAddrPointer_reg[26]/NET0131  & n52333 ;
  assign n52374 = n36792 & ~n52373 ;
  assign n52376 = n39706 & ~n52374 ;
  assign n52375 = ~n39706 & n52374 ;
  assign n52377 = ~\P2_P2_DataWidth_reg[1]/NET0131  & ~n52375 ;
  assign n52378 = ~n52376 & n52377 ;
  assign n52372 = \P2_P2_DataWidth_reg[1]/NET0131  & ~\P2_P2_rEIP_reg[27]/NET0131  ;
  assign n52379 = n26794 & ~n52372 ;
  assign n52380 = ~n52378 & n52379 ;
  assign n52371 = \P2_P2_PhyAddrPointer_reg[27]/NET0131  & n27637 ;
  assign n52404 = \P2_P2_rEIP_reg[27]/NET0131  & ~n50636 ;
  assign n52405 = ~n52371 & ~n52404 ;
  assign n52406 = ~n52380 & n52405 ;
  assign n52407 = ~n52403 & n52406 ;
  assign n52409 = \P2_P2_rEIP_reg[28]/NET0131  & ~n50640 ;
  assign n52411 = ~\P2_P2_rEIP_reg[28]/NET0131  & ~n52382 ;
  assign n52412 = \P2_P2_rEIP_reg[28]/NET0131  & n52382 ;
  assign n52413 = ~n52411 & ~n52412 ;
  assign n52414 = n50649 & ~n52413 ;
  assign n52415 = ~n26650 & n52414 ;
  assign n52410 = ~\P2_P2_EBX_reg[28]/NET0131  & ~n50642 ;
  assign n52416 = n26643 & ~n52410 ;
  assign n52417 = ~n52415 & n52416 ;
  assign n52418 = ~\P2_P2_EBX_reg[27]/NET0131  & n52392 ;
  assign n52419 = \P2_P2_EBX_reg[31]/NET0131  & ~n52418 ;
  assign n52421 = \P2_P2_EBX_reg[28]/NET0131  & ~n52419 ;
  assign n52420 = ~\P2_P2_EBX_reg[28]/NET0131  & n52419 ;
  assign n52422 = ~n50649 & ~n52420 ;
  assign n52423 = ~n52421 & n52422 ;
  assign n52424 = n26633 & ~n52414 ;
  assign n52425 = ~n52423 & n52424 ;
  assign n52426 = ~n52417 & ~n52425 ;
  assign n52427 = ~n26640 & ~n52426 ;
  assign n52428 = ~n52409 & ~n52427 ;
  assign n52429 = n26792 & ~n52428 ;
  assign n52432 = \P2_P2_PhyAddrPointer_reg[27]/NET0131  & n52373 ;
  assign n52433 = n36792 & ~n52432 ;
  assign n52435 = ~n39724 & n52433 ;
  assign n52434 = n39724 & ~n52433 ;
  assign n52436 = ~\P2_P2_DataWidth_reg[1]/NET0131  & ~n52434 ;
  assign n52437 = ~n52435 & n52436 ;
  assign n52431 = \P2_P2_DataWidth_reg[1]/NET0131  & ~\P2_P2_rEIP_reg[28]/NET0131  ;
  assign n52438 = n26794 & ~n52431 ;
  assign n52439 = ~n52437 & n52438 ;
  assign n52408 = \P2_P2_PhyAddrPointer_reg[28]/NET0131  & n27637 ;
  assign n52430 = \P2_P2_rEIP_reg[28]/NET0131  & ~n50636 ;
  assign n52440 = ~n52408 & ~n52430 ;
  assign n52441 = ~n52439 & n52440 ;
  assign n52442 = ~n52429 & n52441 ;
  assign n52445 = ~\P2_P2_EBX_reg[29]/NET0131  & ~n50642 ;
  assign n52446 = \P2_P2_rEIP_reg[29]/NET0131  & n52412 ;
  assign n52447 = ~\P2_P2_rEIP_reg[29]/NET0131  & ~n52412 ;
  assign n52448 = ~n52446 & ~n52447 ;
  assign n52449 = n50649 & ~n52448 ;
  assign n52450 = ~n26650 & n52449 ;
  assign n52451 = ~n52445 & ~n52450 ;
  assign n52452 = ~n26640 & ~n52451 ;
  assign n52453 = n26643 & ~n52452 ;
  assign n52454 = ~n52352 & ~n52453 ;
  assign n52455 = \P2_P2_rEIP_reg[29]/NET0131  & ~n52454 ;
  assign n52456 = ~\P2_P2_EBX_reg[28]/NET0131  & n52418 ;
  assign n52457 = \P2_P2_EBX_reg[31]/NET0131  & ~n52456 ;
  assign n52459 = ~\P2_P2_EBX_reg[29]/NET0131  & n52457 ;
  assign n52458 = \P2_P2_EBX_reg[29]/NET0131  & ~n52457 ;
  assign n52460 = ~n50649 & ~n52458 ;
  assign n52461 = ~n52459 & n52460 ;
  assign n52462 = n26633 & ~n52449 ;
  assign n52463 = ~n52461 & n52462 ;
  assign n52464 = ~n52453 & ~n52463 ;
  assign n52465 = ~n26640 & ~n52464 ;
  assign n52466 = ~n52455 & ~n52465 ;
  assign n52467 = n26792 & ~n52466 ;
  assign n52469 = ~n39706 & ~n41935 ;
  assign n52470 = ~n39724 & n52469 ;
  assign n52471 = n36761 & n52333 ;
  assign n52472 = n52470 & n52471 ;
  assign n52473 = n36792 & ~n52472 ;
  assign n52475 = n39742 & ~n52473 ;
  assign n52474 = ~n39742 & n52473 ;
  assign n52476 = ~\P2_P2_DataWidth_reg[1]/NET0131  & ~n52474 ;
  assign n52477 = ~n52475 & n52476 ;
  assign n52468 = \P2_P2_DataWidth_reg[1]/NET0131  & ~\P2_P2_rEIP_reg[29]/NET0131  ;
  assign n52478 = n26794 & ~n52468 ;
  assign n52479 = ~n52477 & n52478 ;
  assign n52443 = \P2_P2_PhyAddrPointer_reg[29]/NET0131  & n27637 ;
  assign n52444 = \P2_P2_rEIP_reg[29]/NET0131  & ~n50636 ;
  assign n52480 = ~n52443 & ~n52444 ;
  assign n52481 = ~n52479 & n52480 ;
  assign n52482 = ~n52467 & n52481 ;
  assign n52485 = ~\P2_P2_PhyAddrPointer_reg[0]/NET0131  & \P2_P2_PhyAddrPointer_reg[1]/NET0131  ;
  assign n52486 = n36792 & ~n52485 ;
  assign n52487 = ~\P2_P2_PhyAddrPointer_reg[1]/NET0131  & ~\P2_P2_PhyAddrPointer_reg[2]/NET0131  ;
  assign n52488 = ~n47451 & ~n52487 ;
  assign n52490 = ~n52486 & n52488 ;
  assign n52489 = n52486 & ~n52488 ;
  assign n52491 = ~\P2_P2_DataWidth_reg[1]/NET0131  & ~n52489 ;
  assign n52492 = ~n52490 & n52491 ;
  assign n52484 = \P2_P2_DataWidth_reg[1]/NET0131  & ~\P2_P2_rEIP_reg[2]/NET0131  ;
  assign n52493 = n26794 & ~n52484 ;
  assign n52494 = ~n52492 & n52493 ;
  assign n52497 = \P2_P2_rEIP_reg[2]/NET0131  & ~n50640 ;
  assign n52498 = ~\P2_P2_rEIP_reg[1]/NET0131  & ~\P2_P2_rEIP_reg[2]/NET0131  ;
  assign n52499 = ~\P2_P2_DataWidth_reg[1]/NET0131  & ~n50684 ;
  assign n52500 = ~n52498 & n52499 ;
  assign n52501 = ~n26286 & n52500 ;
  assign n52502 = \P2_P2_EBX_reg[31]/NET0131  & ~n50650 ;
  assign n52504 = \P2_P2_EBX_reg[2]/NET0131  & n52502 ;
  assign n52503 = ~\P2_P2_EBX_reg[2]/NET0131  & ~n52502 ;
  assign n52505 = ~n50649 & ~n52503 ;
  assign n52506 = ~n52504 & n52505 ;
  assign n52507 = ~n52501 & ~n52506 ;
  assign n52508 = n47684 & ~n52507 ;
  assign n52496 = n26690 & n50638 ;
  assign n52509 = \P2_P2_EBX_reg[2]/NET0131  & ~n50642 ;
  assign n52510 = n26651 & n52500 ;
  assign n52511 = ~n52509 & ~n52510 ;
  assign n52512 = n26786 & ~n52511 ;
  assign n52513 = ~n52496 & ~n52512 ;
  assign n52514 = ~n52508 & n52513 ;
  assign n52515 = ~n52497 & n52514 ;
  assign n52516 = n26792 & ~n52515 ;
  assign n52483 = \P2_P2_PhyAddrPointer_reg[2]/NET0131  & n27637 ;
  assign n52495 = \P2_P2_rEIP_reg[2]/NET0131  & ~n50636 ;
  assign n52517 = ~n52483 & ~n52495 ;
  assign n52518 = ~n52516 & n52517 ;
  assign n52519 = ~n52494 & n52518 ;
  assign n52576 = n36844 & n50708 ;
  assign n52577 = n42107 & n52576 ;
  assign n52578 = n36847 & n52577 ;
  assign n52579 = ~n36863 & ~n52578 ;
  assign n52581 = n42124 & ~n52579 ;
  assign n52580 = ~n42124 & n52579 ;
  assign n52582 = ~\P2_P3_DataWidth_reg[1]/NET0131  & ~n52580 ;
  assign n52583 = ~n52581 & n52582 ;
  assign n52575 = \P2_P3_DataWidth_reg[1]/NET0131  & ~\P2_P3_rEIP_reg[20]/NET0131  ;
  assign n52584 = n27315 & ~n52575 ;
  assign n52585 = ~n52583 & n52584 ;
  assign n52521 = \P2_P3_rEIP_reg[20]/NET0131  & ~n27277 ;
  assign n52522 = ~\P2_P3_EBX_reg[20]/NET0131  & ~n50735 ;
  assign n52523 = n27121 & ~n52522 ;
  assign n52524 = ~\P2_P3_EBX_reg[3]/NET0131  & n50721 ;
  assign n52525 = ~\P2_P3_EBX_reg[4]/NET0131  & n52524 ;
  assign n52526 = ~\P2_P3_EBX_reg[5]/NET0131  & n52525 ;
  assign n52527 = ~\P2_P3_EBX_reg[6]/NET0131  & n52526 ;
  assign n52528 = ~\P2_P3_EBX_reg[7]/NET0131  & n52527 ;
  assign n52529 = ~\P2_P3_EBX_reg[8]/NET0131  & n52528 ;
  assign n52530 = ~\P2_P3_EBX_reg[9]/NET0131  & n52529 ;
  assign n52531 = ~\P2_P3_EBX_reg[10]/NET0131  & n52530 ;
  assign n52532 = ~\P2_P3_EBX_reg[11]/NET0131  & n52531 ;
  assign n52533 = ~\P2_P3_EBX_reg[12]/NET0131  & n52532 ;
  assign n52534 = ~\P2_P3_EBX_reg[13]/NET0131  & n52533 ;
  assign n52535 = ~\P2_P3_EBX_reg[14]/NET0131  & n52534 ;
  assign n52536 = ~\P2_P3_EBX_reg[15]/NET0131  & n52535 ;
  assign n52537 = ~\P2_P3_EBX_reg[16]/NET0131  & n52536 ;
  assign n52538 = ~\P2_P3_EBX_reg[17]/NET0131  & n52537 ;
  assign n52539 = ~\P2_P3_EBX_reg[18]/NET0131  & n52538 ;
  assign n52540 = ~\P2_P3_EBX_reg[19]/NET0131  & n52539 ;
  assign n52541 = \P2_P3_EBX_reg[31]/NET0131  & ~n52540 ;
  assign n52543 = ~\P2_P3_EBX_reg[20]/NET0131  & n52541 ;
  assign n52542 = \P2_P3_EBX_reg[20]/NET0131  & ~n52541 ;
  assign n52544 = ~n27302 & ~n52542 ;
  assign n52545 = ~n52543 & n52544 ;
  assign n52546 = n27122 & ~n52545 ;
  assign n52547 = ~n52523 & ~n52546 ;
  assign n52549 = \P2_P3_rEIP_reg[4]/NET0131  & n50728 ;
  assign n52550 = \P2_P3_rEIP_reg[5]/NET0131  & n52549 ;
  assign n52551 = \P2_P3_rEIP_reg[6]/NET0131  & n52550 ;
  assign n52552 = \P2_P3_rEIP_reg[7]/NET0131  & n52551 ;
  assign n52553 = \P2_P3_rEIP_reg[8]/NET0131  & n52552 ;
  assign n52554 = \P2_P3_rEIP_reg[9]/NET0131  & n52553 ;
  assign n52555 = \P2_P3_rEIP_reg[10]/NET0131  & n52554 ;
  assign n52556 = \P2_P3_rEIP_reg[11]/NET0131  & n52555 ;
  assign n52557 = \P2_P3_rEIP_reg[12]/NET0131  & n52556 ;
  assign n52558 = \P2_P3_rEIP_reg[13]/NET0131  & n52557 ;
  assign n52559 = \P2_P3_rEIP_reg[14]/NET0131  & n52558 ;
  assign n52560 = \P2_P3_rEIP_reg[15]/NET0131  & n52559 ;
  assign n52561 = \P2_P3_rEIP_reg[16]/NET0131  & n52560 ;
  assign n52562 = \P2_P3_rEIP_reg[17]/NET0131  & n52561 ;
  assign n52563 = \P2_P3_rEIP_reg[18]/NET0131  & n52562 ;
  assign n52564 = \P2_P3_rEIP_reg[19]/NET0131  & n52563 ;
  assign n52565 = ~\P2_P3_rEIP_reg[20]/NET0131  & ~n52564 ;
  assign n52566 = \P2_P3_rEIP_reg[20]/NET0131  & n52564 ;
  assign n52567 = ~n52565 & ~n52566 ;
  assign n52548 = n27148 & n52523 ;
  assign n52568 = n27302 & ~n52548 ;
  assign n52569 = ~n52567 & n52568 ;
  assign n52570 = ~n27177 & ~n52569 ;
  assign n52571 = ~n52547 & n52570 ;
  assign n52572 = ~n52521 & ~n52571 ;
  assign n52573 = n27308 & ~n52572 ;
  assign n52520 = \P2_P3_PhyAddrPointer_reg[20]/NET0131  & n27651 ;
  assign n52574 = \P2_P3_rEIP_reg[20]/NET0131  & ~n50703 ;
  assign n52586 = ~n52520 & ~n52574 ;
  assign n52587 = ~n52573 & n52586 ;
  assign n52588 = ~n52585 & n52587 ;
  assign n52613 = ~\P2_P3_PhyAddrPointer_reg[20]/NET0131  & ~n36863 ;
  assign n52614 = ~n52579 & ~n52613 ;
  assign n52616 = n44130 & n52614 ;
  assign n52615 = ~n44130 & ~n52614 ;
  assign n52617 = ~\P2_P3_DataWidth_reg[1]/NET0131  & ~n52615 ;
  assign n52618 = ~n52616 & n52617 ;
  assign n52612 = \P2_P3_DataWidth_reg[1]/NET0131  & ~\P2_P3_rEIP_reg[21]/NET0131  ;
  assign n52619 = n27315 & ~n52612 ;
  assign n52620 = ~n52618 & n52619 ;
  assign n52590 = \P2_P3_rEIP_reg[21]/NET0131  & ~n27277 ;
  assign n52592 = ~\P2_P3_rEIP_reg[21]/NET0131  & ~n52566 ;
  assign n52593 = \P2_P3_rEIP_reg[21]/NET0131  & n52566 ;
  assign n52594 = ~n52592 & ~n52593 ;
  assign n52595 = n50735 & ~n52594 ;
  assign n52591 = ~\P2_P3_EBX_reg[21]/NET0131  & ~n50735 ;
  assign n52596 = n27121 & ~n52591 ;
  assign n52597 = ~n52595 & n52596 ;
  assign n52599 = ~\P2_P3_EBX_reg[20]/NET0131  & n52540 ;
  assign n52600 = \P2_P3_EBX_reg[31]/NET0131  & ~n52599 ;
  assign n52601 = ~\P2_P3_EBX_reg[21]/NET0131  & ~n52600 ;
  assign n52602 = \P2_P3_EBX_reg[21]/NET0131  & n52600 ;
  assign n52603 = ~n52601 & ~n52602 ;
  assign n52604 = ~n27302 & ~n52603 ;
  assign n52598 = n27302 & ~n52594 ;
  assign n52605 = n27122 & ~n52598 ;
  assign n52606 = ~n52604 & n52605 ;
  assign n52607 = ~n52597 & ~n52606 ;
  assign n52608 = ~n27177 & ~n52607 ;
  assign n52609 = ~n52590 & ~n52608 ;
  assign n52610 = n27308 & ~n52609 ;
  assign n52589 = \P2_P3_PhyAddrPointer_reg[21]/NET0131  & n27651 ;
  assign n52611 = \P2_P3_rEIP_reg[21]/NET0131  & ~n50703 ;
  assign n52621 = ~n52589 & ~n52611 ;
  assign n52622 = ~n52610 & n52621 ;
  assign n52623 = ~n52620 & n52622 ;
  assign n52647 = n39870 & n52577 ;
  assign n52648 = ~n36863 & ~n52647 ;
  assign n52650 = ~n42146 & n52648 ;
  assign n52649 = n42146 & ~n52648 ;
  assign n52651 = ~\P2_P3_DataWidth_reg[1]/NET0131  & ~n52649 ;
  assign n52652 = ~n52650 & n52651 ;
  assign n52646 = \P2_P3_DataWidth_reg[1]/NET0131  & ~\P2_P3_rEIP_reg[22]/NET0131  ;
  assign n52653 = n27315 & ~n52646 ;
  assign n52654 = ~n52652 & n52653 ;
  assign n52635 = ~\P2_P3_EBX_reg[21]/NET0131  & n52599 ;
  assign n52636 = \P2_P3_EBX_reg[31]/NET0131  & ~n52635 ;
  assign n52638 = ~\P2_P3_EBX_reg[22]/NET0131  & n52636 ;
  assign n52637 = \P2_P3_EBX_reg[22]/NET0131  & ~n52636 ;
  assign n52639 = ~n27302 & ~n52637 ;
  assign n52640 = ~n52638 & n52639 ;
  assign n52627 = ~\P2_P3_rEIP_reg[22]/NET0131  & ~n52593 ;
  assign n52628 = \P2_P3_rEIP_reg[22]/NET0131  & n52593 ;
  assign n52629 = ~n52627 & ~n52628 ;
  assign n52634 = n27302 & ~n52629 ;
  assign n52641 = n46587 & ~n52634 ;
  assign n52642 = ~n52640 & n52641 ;
  assign n52630 = n50735 & ~n52629 ;
  assign n52626 = ~\P2_P3_EBX_reg[22]/NET0131  & ~n50735 ;
  assign n52631 = n47747 & ~n52626 ;
  assign n52632 = ~n52630 & n52631 ;
  assign n52633 = \P2_P3_rEIP_reg[22]/NET0131  & ~n27277 ;
  assign n52643 = ~n52632 & ~n52633 ;
  assign n52644 = ~n52642 & n52643 ;
  assign n52645 = n27308 & ~n52644 ;
  assign n52624 = \P2_P3_PhyAddrPointer_reg[22]/NET0131  & n27651 ;
  assign n52625 = \P2_P3_rEIP_reg[22]/NET0131  & ~n50703 ;
  assign n52655 = ~n52624 & ~n52625 ;
  assign n52656 = ~n52645 & n52655 ;
  assign n52657 = ~n52654 & n52656 ;
  assign n52660 = ~\P2_P3_EBX_reg[22]/NET0131  & n52635 ;
  assign n52661 = \P2_P3_EBX_reg[31]/NET0131  & ~n52660 ;
  assign n52663 = \P2_P3_EBX_reg[23]/NET0131  & n52661 ;
  assign n52662 = ~\P2_P3_EBX_reg[23]/NET0131  & ~n52661 ;
  assign n52664 = ~n27302 & ~n52662 ;
  assign n52665 = ~n52663 & n52664 ;
  assign n52667 = ~\P2_P3_rEIP_reg[23]/NET0131  & ~n52628 ;
  assign n52666 = \P2_P3_rEIP_reg[23]/NET0131  & n52628 ;
  assign n52668 = ~\P2_P3_DataWidth_reg[1]/NET0131  & ~n52666 ;
  assign n52669 = ~n52667 & n52668 ;
  assign n52670 = ~n27192 & n52669 ;
  assign n52671 = ~n52665 & ~n52670 ;
  assign n52672 = n46587 & ~n52671 ;
  assign n52659 = \P2_P3_rEIP_reg[23]/NET0131  & ~n27277 ;
  assign n52673 = \P2_P3_EBX_reg[23]/NET0131  & ~n50735 ;
  assign n52674 = n50737 & n52669 ;
  assign n52675 = ~n52673 & ~n52674 ;
  assign n52676 = n47747 & ~n52675 ;
  assign n52677 = ~n52659 & ~n52676 ;
  assign n52678 = ~n52672 & n52677 ;
  assign n52679 = n27308 & ~n52678 ;
  assign n52682 = n39871 & n52577 ;
  assign n52683 = ~n36863 & ~n52682 ;
  assign n52685 = n39875 & ~n52683 ;
  assign n52684 = ~n39875 & n52683 ;
  assign n52686 = ~\P2_P3_DataWidth_reg[1]/NET0131  & ~n52684 ;
  assign n52687 = ~n52685 & n52686 ;
  assign n52681 = \P2_P3_DataWidth_reg[1]/NET0131  & ~\P2_P3_rEIP_reg[23]/NET0131  ;
  assign n52688 = n27315 & ~n52681 ;
  assign n52689 = ~n52687 & n52688 ;
  assign n52658 = \P2_P3_PhyAddrPointer_reg[23]/NET0131  & n27651 ;
  assign n52680 = \P2_P3_rEIP_reg[23]/NET0131  & ~n50703 ;
  assign n52690 = ~n52658 & ~n52680 ;
  assign n52691 = ~n52689 & n52690 ;
  assign n52692 = ~n52679 & n52691 ;
  assign n52703 = ~\P2_P3_EBX_reg[23]/NET0131  & n52660 ;
  assign n52704 = \P2_P3_EBX_reg[31]/NET0131  & ~n52703 ;
  assign n52706 = ~\P2_P3_EBX_reg[24]/NET0131  & n52704 ;
  assign n52705 = \P2_P3_EBX_reg[24]/NET0131  & ~n52704 ;
  assign n52707 = ~n27302 & ~n52705 ;
  assign n52708 = ~n52706 & n52707 ;
  assign n52696 = ~\P2_P3_rEIP_reg[24]/NET0131  & ~n52666 ;
  assign n52697 = \P2_P3_rEIP_reg[24]/NET0131  & n52666 ;
  assign n52698 = ~n52696 & ~n52697 ;
  assign n52702 = n27302 & ~n52698 ;
  assign n52709 = n46587 & ~n52702 ;
  assign n52710 = ~n52708 & n52709 ;
  assign n52694 = \P2_P3_rEIP_reg[24]/NET0131  & ~n27277 ;
  assign n52699 = n50735 & ~n52698 ;
  assign n52695 = ~\P2_P3_EBX_reg[24]/NET0131  & ~n50735 ;
  assign n52700 = n47747 & ~n52695 ;
  assign n52701 = ~n52699 & n52700 ;
  assign n52711 = ~n52694 & ~n52701 ;
  assign n52712 = ~n52710 & n52711 ;
  assign n52713 = n27308 & ~n52712 ;
  assign n52716 = ~n36833 & ~n36863 ;
  assign n52717 = ~n52648 & ~n52716 ;
  assign n52719 = n42161 & n52717 ;
  assign n52718 = ~n42161 & ~n52717 ;
  assign n52720 = ~\P2_P3_DataWidth_reg[1]/NET0131  & ~n52718 ;
  assign n52721 = ~n52719 & n52720 ;
  assign n52715 = \P2_P3_DataWidth_reg[1]/NET0131  & ~\P2_P3_rEIP_reg[24]/NET0131  ;
  assign n52722 = n27315 & ~n52715 ;
  assign n52723 = ~n52721 & n52722 ;
  assign n52693 = \P2_P3_PhyAddrPointer_reg[24]/NET0131  & n27651 ;
  assign n52714 = \P2_P3_rEIP_reg[24]/NET0131  & ~n50703 ;
  assign n52724 = ~n52693 & ~n52714 ;
  assign n52725 = ~n52723 & n52724 ;
  assign n52726 = ~n52713 & n52725 ;
  assign n52729 = ~\P2_P3_EBX_reg[24]/NET0131  & n52703 ;
  assign n52730 = ~\P2_P3_EBX_reg[25]/NET0131  & n52729 ;
  assign n52731 = \P2_P3_EBX_reg[31]/NET0131  & ~n52730 ;
  assign n52733 = \P2_P3_EBX_reg[26]/NET0131  & n52731 ;
  assign n52732 = ~\P2_P3_EBX_reg[26]/NET0131  & ~n52731 ;
  assign n52734 = ~n27302 & ~n52732 ;
  assign n52735 = ~n52733 & n52734 ;
  assign n52736 = \P2_P3_rEIP_reg[25]/NET0131  & n52697 ;
  assign n52738 = \P2_P3_rEIP_reg[26]/NET0131  & n52736 ;
  assign n52737 = ~\P2_P3_rEIP_reg[26]/NET0131  & ~n52736 ;
  assign n52739 = ~\P2_P3_DataWidth_reg[1]/NET0131  & ~n52737 ;
  assign n52740 = ~n52738 & n52739 ;
  assign n52741 = ~n27192 & n52740 ;
  assign n52742 = ~n52735 & ~n52741 ;
  assign n52743 = n46587 & ~n52742 ;
  assign n52728 = \P2_P3_rEIP_reg[26]/NET0131  & ~n27277 ;
  assign n52744 = \P2_P3_EBX_reg[26]/NET0131  & ~n50735 ;
  assign n52745 = n50737 & n52740 ;
  assign n52746 = ~n52744 & ~n52745 ;
  assign n52747 = n47747 & ~n52746 ;
  assign n52748 = ~n52728 & ~n52747 ;
  assign n52749 = ~n52743 & n52748 ;
  assign n52750 = n27308 & ~n52749 ;
  assign n52753 = n36854 & n52647 ;
  assign n52754 = ~n36863 & ~n52753 ;
  assign n52756 = n42193 & ~n52754 ;
  assign n52755 = ~n42193 & n52754 ;
  assign n52757 = ~\P2_P3_DataWidth_reg[1]/NET0131  & ~n52755 ;
  assign n52758 = ~n52756 & n52757 ;
  assign n52752 = \P2_P3_DataWidth_reg[1]/NET0131  & ~\P2_P3_rEIP_reg[26]/NET0131  ;
  assign n52759 = n27315 & ~n52752 ;
  assign n52760 = ~n52758 & n52759 ;
  assign n52727 = \P2_P3_PhyAddrPointer_reg[26]/NET0131  & n27651 ;
  assign n52751 = \P2_P3_rEIP_reg[26]/NET0131  & ~n50703 ;
  assign n52761 = ~n52727 & ~n52751 ;
  assign n52762 = ~n52760 & n52761 ;
  assign n52763 = ~n52750 & n52762 ;
  assign n52774 = ~\P2_P3_EBX_reg[26]/NET0131  & n52730 ;
  assign n52775 = \P2_P3_EBX_reg[31]/NET0131  & ~n52774 ;
  assign n52776 = ~\P2_P3_EBX_reg[27]/NET0131  & ~n52775 ;
  assign n52777 = \P2_P3_EBX_reg[27]/NET0131  & n52775 ;
  assign n52778 = ~n52776 & ~n52777 ;
  assign n52779 = ~n27302 & ~n52778 ;
  assign n52767 = ~\P2_P3_rEIP_reg[27]/NET0131  & ~n52738 ;
  assign n52768 = \P2_P3_rEIP_reg[27]/NET0131  & n52738 ;
  assign n52769 = ~n52767 & ~n52768 ;
  assign n52773 = n27302 & ~n52769 ;
  assign n52780 = n46587 & ~n52773 ;
  assign n52781 = ~n52779 & n52780 ;
  assign n52765 = \P2_P3_rEIP_reg[27]/NET0131  & ~n27277 ;
  assign n52770 = n50735 & ~n52769 ;
  assign n52766 = ~\P2_P3_EBX_reg[27]/NET0131  & ~n50735 ;
  assign n52771 = n47747 & ~n52766 ;
  assign n52772 = ~n52770 & n52771 ;
  assign n52782 = ~n52765 & ~n52772 ;
  assign n52783 = ~n52781 & n52782 ;
  assign n52784 = n27308 & ~n52783 ;
  assign n52787 = ~n42193 & n52753 ;
  assign n52788 = ~n36863 & ~n52787 ;
  assign n52790 = n39887 & ~n52788 ;
  assign n52789 = ~n39887 & n52788 ;
  assign n52791 = ~\P2_P3_DataWidth_reg[1]/NET0131  & ~n52789 ;
  assign n52792 = ~n52790 & n52791 ;
  assign n52786 = \P2_P3_DataWidth_reg[1]/NET0131  & ~\P2_P3_rEIP_reg[27]/NET0131  ;
  assign n52793 = n27315 & ~n52786 ;
  assign n52794 = ~n52792 & n52793 ;
  assign n52764 = \P2_P3_PhyAddrPointer_reg[27]/NET0131  & n27651 ;
  assign n52785 = \P2_P3_rEIP_reg[27]/NET0131  & ~n50703 ;
  assign n52795 = ~n52764 & ~n52785 ;
  assign n52796 = ~n52794 & n52795 ;
  assign n52797 = ~n52784 & n52796 ;
  assign n52803 = ~\P2_P3_EBX_reg[27]/NET0131  & n52774 ;
  assign n52804 = \P2_P3_EBX_reg[31]/NET0131  & ~n52803 ;
  assign n52806 = ~\P2_P3_EBX_reg[28]/NET0131  & n52804 ;
  assign n52805 = \P2_P3_EBX_reg[28]/NET0131  & ~n52804 ;
  assign n52807 = ~n27302 & ~n52805 ;
  assign n52808 = ~n52806 & n52807 ;
  assign n52799 = ~\P2_P3_rEIP_reg[28]/NET0131  & ~n52768 ;
  assign n52800 = \P2_P3_rEIP_reg[28]/NET0131  & n52768 ;
  assign n52801 = ~n52799 & ~n52800 ;
  assign n52802 = n27302 & ~n52801 ;
  assign n52809 = n46587 & ~n52802 ;
  assign n52810 = ~n52808 & n52809 ;
  assign n52811 = \P2_P3_rEIP_reg[28]/NET0131  & ~n27277 ;
  assign n52813 = ~n27148 & n52802 ;
  assign n52812 = ~\P2_P3_EBX_reg[28]/NET0131  & ~n50735 ;
  assign n52814 = n47747 & ~n52812 ;
  assign n52815 = ~n52813 & n52814 ;
  assign n52816 = ~n52811 & ~n52815 ;
  assign n52817 = ~n52810 & n52816 ;
  assign n52818 = n27308 & ~n52817 ;
  assign n52821 = ~n39887 & n52787 ;
  assign n52822 = ~n36863 & ~n52821 ;
  assign n52824 = n39910 & ~n52822 ;
  assign n52823 = ~n39910 & n52822 ;
  assign n52825 = ~\P2_P3_DataWidth_reg[1]/NET0131  & ~n52823 ;
  assign n52826 = ~n52824 & n52825 ;
  assign n52820 = \P2_P3_DataWidth_reg[1]/NET0131  & ~\P2_P3_rEIP_reg[28]/NET0131  ;
  assign n52827 = n27315 & ~n52820 ;
  assign n52828 = ~n52826 & n52827 ;
  assign n52798 = \P2_P3_PhyAddrPointer_reg[28]/NET0131  & n27651 ;
  assign n52819 = \P2_P3_rEIP_reg[28]/NET0131  & ~n50703 ;
  assign n52829 = ~n52798 & ~n52819 ;
  assign n52830 = ~n52828 & n52829 ;
  assign n52831 = ~n52818 & n52830 ;
  assign n52833 = n50707 & n50709 ;
  assign n52834 = ~n50710 & ~n52833 ;
  assign n52835 = ~\P2_P3_DataWidth_reg[1]/NET0131  & ~n52834 ;
  assign n52836 = \P2_P3_DataWidth_reg[1]/NET0131  & ~\P2_P3_rEIP_reg[2]/NET0131  ;
  assign n52837 = n27315 & ~n52836 ;
  assign n52838 = ~n52835 & n52837 ;
  assign n52840 = \P2_P3_rEIP_reg[2]/NET0131  & ~n27277 ;
  assign n52842 = ~\P2_P3_rEIP_reg[1]/NET0131  & ~\P2_P3_rEIP_reg[2]/NET0131  ;
  assign n52843 = ~\P2_P3_DataWidth_reg[1]/NET0131  & ~n50727 ;
  assign n52844 = ~n52842 & n52843 ;
  assign n52845 = ~n27192 & n52844 ;
  assign n52846 = \P2_P3_EBX_reg[31]/NET0131  & ~n50720 ;
  assign n52847 = ~\P2_P3_EBX_reg[2]/NET0131  & ~n52846 ;
  assign n52848 = \P2_P3_EBX_reg[2]/NET0131  & n52846 ;
  assign n52849 = ~n52847 & ~n52848 ;
  assign n52850 = ~n27302 & n52849 ;
  assign n52851 = ~n52845 & ~n52850 ;
  assign n52852 = n27122 & ~n52851 ;
  assign n52841 = n27124 & n27251 ;
  assign n52853 = \P2_P3_EBX_reg[2]/NET0131  & ~n50735 ;
  assign n52854 = n50737 & n52844 ;
  assign n52855 = ~n52853 & ~n52854 ;
  assign n52856 = n27121 & ~n52855 ;
  assign n52857 = ~n52841 & ~n52856 ;
  assign n52858 = ~n52852 & n52857 ;
  assign n52859 = ~n27177 & ~n52858 ;
  assign n52860 = ~n52840 & ~n52859 ;
  assign n52861 = n27308 & ~n52860 ;
  assign n52832 = \P2_P3_PhyAddrPointer_reg[2]/NET0131  & n27651 ;
  assign n52839 = \P2_P3_rEIP_reg[2]/NET0131  & ~n50703 ;
  assign n52862 = ~n52832 & ~n52839 ;
  assign n52863 = ~n52861 & n52862 ;
  assign n52864 = ~n52838 & n52863 ;
  assign n52866 = n25701 & n45939 ;
  assign n52867 = \P1_P2_PhyAddrPointer_reg[2]/NET0131  & ~n39340 ;
  assign n52868 = ~n45923 & ~n52867 ;
  assign n52869 = ~n52866 & n52868 ;
  assign n52870 = n25918 & ~n52869 ;
  assign n52871 = \P1_P2_PhyAddrPointer_reg[2]/NET0131  & ~n36595 ;
  assign n52872 = ~\P1_P2_DataWidth_reg[1]/NET0131  & n51586 ;
  assign n52873 = n47787 & ~n52872 ;
  assign n52865 = n27898 & n51587 ;
  assign n52874 = ~n45916 & ~n52865 ;
  assign n52875 = ~n52873 & n52874 ;
  assign n52876 = ~n52871 & n52875 ;
  assign n52877 = ~n52870 & n52876 ;
  assign n52883 = \P1_P2_RequestPending_reg/NET0131  & ~n48371 ;
  assign n52884 = n25415 & ~n25786 ;
  assign n52885 = ~n25787 & ~n25914 ;
  assign n52886 = ~n52884 & n52885 ;
  assign n52887 = ~n25770 & ~n52886 ;
  assign n52888 = ~n52883 & ~n52887 ;
  assign n52889 = n25918 & ~n52888 ;
  assign n52878 = n25415 & n25922 ;
  assign n52879 = ~n27607 & ~n27609 ;
  assign n52880 = ~n52878 & n52879 ;
  assign n52881 = \P1_P2_RequestPending_reg/NET0131  & ~n52880 ;
  assign n52882 = ~n25417 & ~n27967 ;
  assign n52890 = ~n52881 & n52882 ;
  assign n52891 = ~n52889 & n52890 ;
  assign n52893 = n25945 & n45332 ;
  assign n52894 = \P2_P1_PhyAddrPointer_reg[2]/NET0131  & ~n36678 ;
  assign n52895 = ~n45340 & ~n52894 ;
  assign n52896 = ~n52893 & n52895 ;
  assign n52897 = n11623 & ~n52896 ;
  assign n52898 = \P2_P1_PhyAddrPointer_reg[2]/NET0131  & ~n47405 ;
  assign n52892 = n36674 & n50475 ;
  assign n52899 = ~\P2_P1_PhyAddrPointer_reg[2]/NET0131  & n27681 ;
  assign n52900 = ~n45308 & ~n52899 ;
  assign n52901 = ~n52892 & n52900 ;
  assign n52902 = ~n52898 & n52901 ;
  assign n52903 = ~n52897 & n52902 ;
  assign n52909 = \P2_P1_RequestPending_reg/NET0131  & n26088 ;
  assign n52910 = \P2_P1_DataWidth_reg[1]/NET0131  & n26057 ;
  assign n52911 = n25951 & ~n26057 ;
  assign n52912 = ~n24898 & ~n52911 ;
  assign n52913 = ~n24711 & n52912 ;
  assign n52914 = ~n52910 & ~n52913 ;
  assign n52915 = ~n52909 & ~n52914 ;
  assign n52908 = ~\P2_P1_RequestPending_reg/NET0131  & n21081 ;
  assign n52916 = n11623 & ~n52908 ;
  assign n52917 = ~n52915 & n52916 ;
  assign n52904 = n11611 & n27487 ;
  assign n52905 = n21097 & ~n52904 ;
  assign n52906 = \P2_P1_RequestPending_reg/NET0131  & ~n52905 ;
  assign n52907 = ~n11616 & ~n21098 ;
  assign n52918 = ~n52906 & n52907 ;
  assign n52919 = ~n52917 & n52918 ;
  assign n52921 = \P1_P1_PhyAddrPointer_reg[2]/NET0131  & ~n41658 ;
  assign n52922 = n26263 & n45979 ;
  assign n52923 = ~n45994 & ~n52922 ;
  assign n52924 = ~n52921 & n52923 ;
  assign n52925 = n8355 & ~n52924 ;
  assign n52926 = \P1_P1_PhyAddrPointer_reg[2]/NET0131  & ~n47428 ;
  assign n52920 = ~n36701 & n52049 ;
  assign n52927 = ~\P1_P1_PhyAddrPointer_reg[2]/NET0131  & n27791 ;
  assign n52928 = ~n45973 & ~n52927 ;
  assign n52929 = ~n52920 & n52928 ;
  assign n52930 = ~n52926 & n52929 ;
  assign n52931 = ~n52925 & n52930 ;
  assign n52939 = ~n26131 & ~n34141 ;
  assign n52940 = \P1_P1_RequestPending_reg/NET0131  & ~n52939 ;
  assign n52937 = ~\P1_P1_RequestPending_reg/NET0131  & n15364 ;
  assign n52938 = n26255 & ~n52937 ;
  assign n52936 = ~\P1_P1_DataWidth_reg[1]/NET0131  & n24503 ;
  assign n52941 = ~n26266 & ~n52936 ;
  assign n52942 = ~n52938 & n52941 ;
  assign n52943 = ~n52940 & n52942 ;
  assign n52944 = n8355 & ~n52943 ;
  assign n52932 = n8356 & n27624 ;
  assign n52933 = n15323 & ~n52932 ;
  assign n52934 = \P1_P1_RequestPending_reg/NET0131  & ~n52933 ;
  assign n52935 = ~n8357 & ~n15324 ;
  assign n52945 = ~n52934 & n52935 ;
  assign n52946 = ~n52944 & n52945 ;
  assign n52949 = \P2_P2_PhyAddrPointer_reg[2]/NET0131  & ~n41873 ;
  assign n52948 = n26749 & n45548 ;
  assign n52950 = ~n45556 & ~n52948 ;
  assign n52951 = ~n52949 & n52950 ;
  assign n52952 = n26792 & ~n52951 ;
  assign n52953 = ~n26291 & ~n27614 ;
  assign n52954 = ~n26296 & n52953 ;
  assign n52955 = ~n27613 & n52954 ;
  assign n52956 = \P2_P2_PhyAddrPointer_reg[2]/NET0131  & ~n52955 ;
  assign n52947 = ~n36760 & n52488 ;
  assign n52957 = ~\P2_P2_PhyAddrPointer_reg[2]/NET0131  & n26800 ;
  assign n52958 = ~n45533 & ~n52957 ;
  assign n52959 = ~n52947 & n52958 ;
  assign n52960 = ~n52956 & n52959 ;
  assign n52961 = ~n52952 & n52960 ;
  assign n52966 = ~\P2_P2_RequestPending_reg/NET0131  & n26640 ;
  assign n52967 = ~n26654 & ~n52966 ;
  assign n52965 = \P2_P2_RequestPending_reg/NET0131  & n26680 ;
  assign n52968 = ~n26787 & ~n52965 ;
  assign n52969 = ~n52967 & n52968 ;
  assign n52970 = n26792 & ~n52969 ;
  assign n52962 = ~n26289 & n44507 ;
  assign n52963 = \P2_P2_RequestPending_reg/NET0131  & ~n52962 ;
  assign n52964 = ~n27635 & ~n28046 ;
  assign n52971 = ~n52963 & n52964 ;
  assign n52972 = ~n52970 & n52971 ;
  assign n52974 = \P1_P3_PhyAddrPointer_reg[2]/NET0131  & ~n37992 ;
  assign n52975 = n9191 & n20269 ;
  assign n52976 = ~n20290 & ~n52975 ;
  assign n52977 = ~n52974 & n52976 ;
  assign n52978 = n9241 & ~n52977 ;
  assign n52979 = n16913 & ~n36810 ;
  assign n52980 = \P1_P3_PhyAddrPointer_reg[2]/NET0131  & ~n36816 ;
  assign n52973 = ~\P1_P3_PhyAddrPointer_reg[2]/NET0131  & n11698 ;
  assign n52981 = ~n20264 & ~n52973 ;
  assign n52982 = ~n52980 & n52981 ;
  assign n52983 = ~n52979 & n52982 ;
  assign n52984 = ~n52978 & n52983 ;
  assign n52986 = \P2_P3_PhyAddrPointer_reg[2]/NET0131  & ~n39857 ;
  assign n52987 = ~n45774 & ~n52986 ;
  assign n52988 = ~n45781 & n52987 ;
  assign n52989 = n27308 & ~n52988 ;
  assign n52990 = ~n36831 & n50707 ;
  assign n52991 = \P2_P3_PhyAddrPointer_reg[2]/NET0131  & ~n36873 ;
  assign n52985 = ~\P2_P3_PhyAddrPointer_reg[2]/NET0131  & n27325 ;
  assign n52992 = ~n45751 & ~n52985 ;
  assign n52993 = ~n52991 & n52992 ;
  assign n52994 = ~n52990 & n52993 ;
  assign n52995 = ~n52989 & n52994 ;
  assign n52998 = ~\P2_P3_RequestPending_reg/NET0131  & n27177 ;
  assign n52999 = ~n27235 & ~n52998 ;
  assign n52997 = ~\P2_P3_DataWidth_reg[1]/NET0131  & n47747 ;
  assign n53000 = \P2_P3_RequestPending_reg/NET0131  & n27126 ;
  assign n53001 = ~n52997 & ~n53000 ;
  assign n53002 = ~n52999 & n53001 ;
  assign n53003 = n27308 & ~n53002 ;
  assign n52996 = ~n27310 & ~n32864 ;
  assign n53004 = n27317 & n27654 ;
  assign n53005 = n42870 & ~n53004 ;
  assign n53006 = \P2_P3_RequestPending_reg/NET0131  & ~n53005 ;
  assign n53007 = n52996 & ~n53006 ;
  assign n53008 = ~n53003 & n53007 ;
  assign n53010 = n26158 & n26159 ;
  assign n53011 = n26161 & ~n53010 ;
  assign n53012 = ~n26158 & ~n49014 ;
  assign n53013 = n24503 & ~n53012 ;
  assign n53014 = n53011 & ~n53013 ;
  assign n53015 = \P1_P1_Datao_reg[20]/NET0131  & ~n53014 ;
  assign n53016 = ~n26158 & n49015 ;
  assign n53017 = ~n53015 & ~n53016 ;
  assign n53018 = n8355 & ~n53017 ;
  assign n53009 = \P1_P1_uWord_reg[4]/NET0131  & n27790 ;
  assign n53019 = \P1_P1_Datao_reg[20]/NET0131  & ~n48479 ;
  assign n53020 = ~n53009 & ~n53019 ;
  assign n53021 = ~n53018 & n53020 ;
  assign n53023 = ~\P2_P2_EAX_reg[20]/NET0131  & ~n47663 ;
  assign n53024 = ~n47664 & ~n53023 ;
  assign n53025 = ~n26650 & ~n53024 ;
  assign n53026 = n26786 & ~n53025 ;
  assign n53027 = n48494 & ~n53026 ;
  assign n53028 = \P2_P2_Datao_reg[20]/NET0131  & ~n53027 ;
  assign n53029 = n26786 & n53024 ;
  assign n53030 = ~n26650 & n53029 ;
  assign n53031 = ~n53028 & ~n53030 ;
  assign n53032 = n26792 & ~n53031 ;
  assign n53022 = \P2_P2_uWord_reg[4]/NET0131  & n48491 ;
  assign n53033 = \P2_P2_Datao_reg[20]/NET0131  & ~n48508 ;
  assign n53034 = ~n53022 & ~n53033 ;
  assign n53035 = ~n53032 & n53034 ;
  assign n53037 = \P2_P3_Datao_reg[20]/NET0131  & ~n27223 ;
  assign n53038 = ~\P2_P3_EAX_reg[20]/NET0131  & ~n47776 ;
  assign n53039 = ~n48526 & ~n53038 ;
  assign n53040 = n47747 & n53039 ;
  assign n53041 = ~n27148 & n53040 ;
  assign n53042 = ~n53037 & ~n53041 ;
  assign n53043 = n27308 & ~n53042 ;
  assign n53036 = \P2_P3_uWord_reg[4]/NET0131  & n48523 ;
  assign n53044 = \P2_P3_Datao_reg[20]/NET0131  & ~n48540 ;
  assign n53045 = ~n53036 & ~n53044 ;
  assign n53046 = ~n53043 & n53045 ;
  assign n53048 = ~\P1_P2_EAX_reg[20]/NET0131  & ~n47550 ;
  assign n53049 = ~n47551 & ~n53048 ;
  assign n53050 = ~n25768 & ~n53049 ;
  assign n53051 = n47570 & ~n53050 ;
  assign n53052 = n48554 & ~n53051 ;
  assign n53053 = \P1_P2_Datao_reg[20]/NET0131  & ~n53052 ;
  assign n53054 = n47570 & n53049 ;
  assign n53055 = ~n25768 & n53054 ;
  assign n53056 = ~n53053 & ~n53055 ;
  assign n53057 = n25918 & ~n53056 ;
  assign n53047 = \P1_P2_uWord_reg[4]/NET0131  & n25922 ;
  assign n53058 = \P1_P2_Datao_reg[20]/NET0131  & ~n48566 ;
  assign n53059 = ~n53047 & ~n53058 ;
  assign n53060 = ~n53057 & n53059 ;
  assign n53062 = ~n25958 & ~n48641 ;
  assign n53063 = n24899 & ~n53062 ;
  assign n53064 = n48584 & ~n53063 ;
  assign n53065 = \P2_P1_Datao_reg[20]/NET0131  & ~n53064 ;
  assign n53066 = ~n25958 & n48642 ;
  assign n53067 = ~n53065 & ~n53066 ;
  assign n53068 = n11623 & ~n53067 ;
  assign n53061 = \P2_P1_uWord_reg[4]/NET0131  & n48581 ;
  assign n53069 = \P2_P1_Datao_reg[20]/NET0131  & ~n48594 ;
  assign n53070 = ~n53061 & ~n53069 ;
  assign n53071 = ~n53068 & n53070 ;
  assign n53072 = \P2_P1_EAX_reg[1]/NET0131  & ~n21100 ;
  assign n53073 = ~\P2_P1_EAX_reg[0]/NET0131  & n21022 ;
  assign n53074 = ~n21072 & ~n53073 ;
  assign n53075 = \P2_P1_EAX_reg[1]/NET0131  & ~n53074 ;
  assign n53079 = \P2_P1_EAX_reg[1]/NET0131  & ~n22337 ;
  assign n53080 = ~n25140 & ~n53079 ;
  assign n53081 = ~n21069 & ~n53080 ;
  assign n53076 = \P2_P1_EAX_reg[0]/NET0131  & ~\P2_P1_EAX_reg[1]/NET0131  ;
  assign n53077 = n21022 & n53076 ;
  assign n53078 = n20728 & ~n31752 ;
  assign n53082 = ~n53077 & ~n53078 ;
  assign n53083 = ~n53081 & n53082 ;
  assign n53084 = ~n53075 & n53083 ;
  assign n53085 = n11623 & ~n53084 ;
  assign n53086 = ~n53072 & ~n53085 ;
  assign n53087 = \P1_P1_EAX_reg[1]/NET0131  & ~n15326 ;
  assign n53089 = ~\P1_P1_EAX_reg[0]/NET0131  & n15377 ;
  assign n53090 = n24346 & ~n53089 ;
  assign n53091 = \P1_P1_EAX_reg[1]/NET0131  & ~n53090 ;
  assign n53088 = n7920 & n24342 ;
  assign n53092 = n22818 & ~n33764 ;
  assign n53093 = \P1_P1_EAX_reg[0]/NET0131  & ~\P1_P1_EAX_reg[1]/NET0131  ;
  assign n53094 = n15377 & n53093 ;
  assign n53095 = ~n53092 & ~n53094 ;
  assign n53096 = ~n53088 & n53095 ;
  assign n53097 = ~n53091 & n53096 ;
  assign n53098 = n8355 & ~n53097 ;
  assign n53099 = ~n53087 & ~n53098 ;
  assign n53100 = \P1_P1_EAX_reg[0]/NET0131  & ~n27551 ;
  assign n53102 = ~n7924 & n24342 ;
  assign n53101 = n22818 & ~n33797 ;
  assign n53103 = ~n53089 & ~n53101 ;
  assign n53104 = ~n53102 & n53103 ;
  assign n53105 = n8355 & ~n53104 ;
  assign n53106 = ~n53100 & ~n53105 ;
  assign n53107 = \P2_P1_lWord_reg[2]/NET0131  & ~n34408 ;
  assign n53108 = \P2_P1_EAX_reg[2]/NET0131  & n24899 ;
  assign n53109 = n21062 & n24838 ;
  assign n53110 = ~n53108 & ~n53109 ;
  assign n53111 = n11623 & ~n53110 ;
  assign n53112 = ~n53107 & ~n53111 ;
  assign n53113 = n25918 & ~n47572 ;
  assign n53114 = n47529 & ~n53113 ;
  assign n53115 = \P1_P2_uWord_reg[4]/NET0131  & ~n53114 ;
  assign n53116 = n25773 & n25776 ;
  assign n53117 = ~n27937 & n53116 ;
  assign n53118 = ~n53054 & ~n53117 ;
  assign n53119 = n25918 & ~n53118 ;
  assign n53120 = ~n53115 & ~n53119 ;
  assign n53121 = \P2_P2_EAX_reg[0]/NET0131  & ~n48669 ;
  assign n53124 = n26761 & ~n46777 ;
  assign n53122 = ~\P2_P2_EAX_reg[0]/NET0131  & n44732 ;
  assign n53123 = ~n32465 & n44510 ;
  assign n53125 = ~n53122 & ~n53123 ;
  assign n53126 = ~n53124 & n53125 ;
  assign n53127 = n26792 & ~n53126 ;
  assign n53128 = ~n53121 & ~n53127 ;
  assign n53129 = \P2_P2_EAX_reg[1]/NET0131  & ~n44508 ;
  assign n53132 = n46402 & ~n53122 ;
  assign n53133 = \P2_P2_EAX_reg[1]/NET0131  & ~n53132 ;
  assign n53130 = n26641 & ~n40774 ;
  assign n53131 = ~n26639 & n53130 ;
  assign n53134 = ~n32432 & n44510 ;
  assign n53135 = \P2_P2_EAX_reg[0]/NET0131  & ~\P2_P2_EAX_reg[1]/NET0131  ;
  assign n53136 = n44732 & n53135 ;
  assign n53137 = ~n53134 & ~n53136 ;
  assign n53138 = ~n53131 & n53137 ;
  assign n53139 = ~n53133 & n53138 ;
  assign n53140 = n26792 & ~n53139 ;
  assign n53141 = ~n53129 & ~n53140 ;
  assign n53142 = \P2_P2_EAX_reg[25]/NET0131  & ~n44508 ;
  assign n53146 = \P2_P2_EAX_reg[25]/NET0131  & ~n47582 ;
  assign n53147 = n44728 & n47581 ;
  assign n53148 = \P2_P2_EAX_reg[25]/NET0131  & ~n26641 ;
  assign n53152 = ~n48947 & ~n53148 ;
  assign n53153 = n26633 & ~n53152 ;
  assign n53143 = ~n44605 & n44636 ;
  assign n53144 = ~n44637 & ~n53143 ;
  assign n53145 = n44510 & n53144 ;
  assign n53149 = n26641 & ~n40785 ;
  assign n53150 = ~n53148 & ~n53149 ;
  assign n53151 = n26638 & ~n53150 ;
  assign n53154 = ~n53145 & ~n53151 ;
  assign n53155 = ~n53153 & n53154 ;
  assign n53156 = ~n53147 & n53155 ;
  assign n53157 = ~n53146 & n53156 ;
  assign n53158 = n26792 & ~n53157 ;
  assign n53159 = ~n53142 & ~n53158 ;
  assign n53160 = \P2_P2_EAX_reg[2]/NET0131  & ~n48669 ;
  assign n53162 = n26761 & ~n35991 ;
  assign n53161 = ~n32399 & n44510 ;
  assign n53163 = ~\P2_P2_EAX_reg[2]/NET0131  & ~n44705 ;
  assign n53164 = ~n44706 & ~n53163 ;
  assign n53165 = n44732 & n53164 ;
  assign n53166 = ~n53161 & ~n53165 ;
  assign n53167 = ~n53162 & n53166 ;
  assign n53168 = n26792 & ~n53167 ;
  assign n53169 = ~n53160 & ~n53168 ;
  assign n53170 = \P2_P2_EAX_reg[3]/NET0131  & ~n48669 ;
  assign n53172 = n26761 & ~n29888 ;
  assign n53171 = ~n32364 & n44510 ;
  assign n53173 = ~\P2_P2_EAX_reg[3]/NET0131  & ~n44706 ;
  assign n53174 = ~n44707 & ~n53173 ;
  assign n53175 = n44732 & n53174 ;
  assign n53176 = ~n53171 & ~n53175 ;
  assign n53177 = ~n53172 & n53176 ;
  assign n53178 = n26792 & ~n53177 ;
  assign n53179 = ~n53170 & ~n53178 ;
  assign n53180 = \P2_P2_EAX_reg[4]/NET0131  & ~n48669 ;
  assign n53182 = n26641 & ~n28016 ;
  assign n53183 = ~n26639 & n53182 ;
  assign n53181 = ~n32329 & n44510 ;
  assign n53184 = ~\P2_P2_EAX_reg[4]/NET0131  & ~n44707 ;
  assign n53185 = ~n44708 & ~n53184 ;
  assign n53186 = n44732 & n53185 ;
  assign n53187 = ~n53181 & ~n53186 ;
  assign n53188 = ~n53183 & n53187 ;
  assign n53189 = n26792 & ~n53188 ;
  assign n53190 = ~n53180 & ~n53189 ;
  assign n53191 = \P2_P2_EAX_reg[5]/NET0131  & ~n44508 ;
  assign n53192 = ~n44709 & n44732 ;
  assign n53194 = ~n44736 & ~n53192 ;
  assign n53195 = \P2_P2_EAX_reg[5]/NET0131  & ~n53194 ;
  assign n53197 = \P2_P2_EAX_reg[5]/NET0131  & ~n26641 ;
  assign n53198 = n26641 & ~n39023 ;
  assign n53199 = ~n53197 & ~n53198 ;
  assign n53200 = ~n26639 & ~n53199 ;
  assign n53193 = n44708 & n53192 ;
  assign n53196 = ~n32294 & n44510 ;
  assign n53201 = ~n53193 & ~n53196 ;
  assign n53202 = ~n53200 & n53201 ;
  assign n53203 = ~n53195 & n53202 ;
  assign n53204 = n26792 & ~n53203 ;
  assign n53205 = ~n53191 & ~n53204 ;
  assign n53206 = \P2_P2_EAX_reg[6]/NET0131  & ~n44508 ;
  assign n53209 = \P2_P2_EAX_reg[6]/NET0131  & ~n53194 ;
  assign n53211 = \P2_P2_EAX_reg[6]/NET0131  & ~n26641 ;
  assign n53212 = n26641 & ~n34477 ;
  assign n53213 = ~n53211 & ~n53212 ;
  assign n53214 = ~n26639 & ~n53213 ;
  assign n53207 = ~\P2_P2_EAX_reg[6]/NET0131  & n44709 ;
  assign n53208 = n44732 & n53207 ;
  assign n53210 = ~n32259 & n44510 ;
  assign n53215 = ~n53208 & ~n53210 ;
  assign n53216 = ~n53214 & n53215 ;
  assign n53217 = ~n53209 & n53216 ;
  assign n53218 = n26792 & ~n53217 ;
  assign n53219 = ~n53206 & ~n53218 ;
  assign n53220 = n7947 & n23946 ;
  assign n53221 = \P1_P1_EAX_reg[2]/NET0131  & n24502 ;
  assign n53222 = ~n53220 & ~n53221 ;
  assign n53223 = ~n15364 & ~n53222 ;
  assign n53224 = \P1_P1_lWord_reg[2]/NET0131  & ~n24506 ;
  assign n53225 = ~n53223 & ~n53224 ;
  assign n53226 = n8355 & ~n53225 ;
  assign n53227 = \P1_P1_lWord_reg[2]/NET0131  & ~n24515 ;
  assign n53228 = ~n53226 & ~n53227 ;
  assign n53229 = \P2_P1_EAX_reg[0]/NET0131  & ~n27438 ;
  assign n53231 = n11379 & n24708 ;
  assign n53230 = n20728 & ~n31785 ;
  assign n53232 = ~n53073 & ~n53230 ;
  assign n53233 = ~n53231 & n53232 ;
  assign n53234 = n11623 & ~n53233 ;
  assign n53235 = ~n53229 & ~n53234 ;
  assign n53236 = \P2_P2_uWord_reg[4]/NET0131  & ~n47642 ;
  assign n53240 = \P2_P2_uWord_reg[4]/NET0131  & n47685 ;
  assign n53237 = \P2_P2_uWord_reg[4]/NET0131  & n26286 ;
  assign n53238 = ~n53182 & ~n53237 ;
  assign n53239 = n26633 & ~n53238 ;
  assign n53241 = ~n53029 & ~n53239 ;
  assign n53242 = ~n53240 & n53241 ;
  assign n53243 = n26792 & ~n53242 ;
  assign n53244 = ~n53236 & ~n53243 ;
  assign n53245 = \P2_P3_EAX_reg[0]/NET0131  & ~n49039 ;
  assign n53248 = \P2_buf2_reg[0]/NET0131  & n27227 ;
  assign n53249 = ~n27226 & n53248 ;
  assign n53246 = ~n33196 & n42538 ;
  assign n53247 = ~\P2_P3_EAX_reg[0]/NET0131  & n42539 ;
  assign n53250 = ~n53246 & ~n53247 ;
  assign n53251 = ~n53249 & n53250 ;
  assign n53252 = n27308 & ~n53251 ;
  assign n53253 = ~n53245 & ~n53252 ;
  assign n53254 = \P2_P3_EAX_reg[1]/NET0131  & ~n42872 ;
  assign n53256 = n42543 & ~n53247 ;
  assign n53257 = \P2_P3_EAX_reg[1]/NET0131  & ~n53256 ;
  assign n53255 = \P2_buf2_reg[1]/NET0131  & n27228 ;
  assign n53258 = ~n33163 & n42538 ;
  assign n53259 = \P2_P3_EAX_reg[0]/NET0131  & ~\P2_P3_EAX_reg[1]/NET0131  ;
  assign n53260 = n42539 & n53259 ;
  assign n53261 = ~n53258 & ~n53260 ;
  assign n53262 = ~n53255 & n53261 ;
  assign n53263 = ~n53257 & n53262 ;
  assign n53264 = n27308 & ~n53263 ;
  assign n53265 = ~n53254 & ~n53264 ;
  assign n53267 = ~\P2_P3_EAX_reg[25]/NET0131  & ~n42856 ;
  assign n53268 = n42539 & ~n42857 ;
  assign n53269 = ~n53267 & n53268 ;
  assign n53266 = \P2_P3_EAX_reg[25]/NET0131  & ~n42543 ;
  assign n53270 = \P2_buf2_reg[9]/NET0131  & n27122 ;
  assign n53271 = \P2_buf2_reg[25]/NET0131  & n27186 ;
  assign n53272 = ~n53270 & ~n53271 ;
  assign n53273 = n27227 & ~n53272 ;
  assign n53274 = ~n42639 & n42670 ;
  assign n53275 = ~n42671 & ~n53274 ;
  assign n53276 = n42538 & n53275 ;
  assign n53277 = ~n53273 & ~n53276 ;
  assign n53278 = ~n53266 & n53277 ;
  assign n53279 = ~n53269 & n53278 ;
  assign n53280 = n27308 & ~n53279 ;
  assign n53281 = \P2_P3_EAX_reg[25]/NET0131  & ~n42872 ;
  assign n53282 = ~n53280 & ~n53281 ;
  assign n53283 = \P2_P3_EAX_reg[2]/NET0131  & ~n49039 ;
  assign n53285 = \P2_buf2_reg[2]/NET0131  & n27228 ;
  assign n53284 = ~n33130 & n42538 ;
  assign n53286 = ~\P2_P3_EAX_reg[2]/NET0131  & ~n42833 ;
  assign n53287 = ~n42834 & ~n53286 ;
  assign n53288 = n42539 & n53287 ;
  assign n53289 = ~n53284 & ~n53288 ;
  assign n53290 = ~n53285 & n53289 ;
  assign n53291 = n27308 & ~n53290 ;
  assign n53292 = ~n53283 & ~n53291 ;
  assign n53293 = \P2_P3_EAX_reg[3]/NET0131  & ~n49039 ;
  assign n53295 = \P2_buf2_reg[3]/NET0131  & n27228 ;
  assign n53294 = ~n33095 & n42538 ;
  assign n53296 = ~\P2_P3_EAX_reg[3]/NET0131  & ~n42834 ;
  assign n53297 = ~n42835 & ~n53296 ;
  assign n53298 = n42539 & n53297 ;
  assign n53299 = ~n53294 & ~n53298 ;
  assign n53300 = ~n53295 & n53299 ;
  assign n53301 = n27308 & ~n53300 ;
  assign n53302 = ~n53293 & ~n53301 ;
  assign n53303 = \P2_P3_EAX_reg[4]/NET0131  & ~n49039 ;
  assign n53305 = \P2_buf2_reg[4]/NET0131  & n27228 ;
  assign n53304 = ~n33060 & n42538 ;
  assign n53306 = ~\P2_P3_EAX_reg[4]/NET0131  & ~n42835 ;
  assign n53307 = ~n42836 & ~n53306 ;
  assign n53308 = n42539 & n53307 ;
  assign n53309 = ~n53304 & ~n53308 ;
  assign n53310 = ~n53305 & n53309 ;
  assign n53311 = n27308 & ~n53310 ;
  assign n53312 = ~n53303 & ~n53311 ;
  assign n53313 = \P2_P3_EAX_reg[5]/NET0131  & ~n42872 ;
  assign n53316 = n42539 & ~n42837 ;
  assign n53317 = n42543 & ~n53316 ;
  assign n53318 = \P2_P3_EAX_reg[5]/NET0131  & ~n53317 ;
  assign n53314 = \P2_buf2_reg[5]/NET0131  & ~n27192 ;
  assign n53315 = n27256 & n53314 ;
  assign n53319 = ~n33025 & n42538 ;
  assign n53320 = n42836 & n53316 ;
  assign n53321 = ~n53319 & ~n53320 ;
  assign n53322 = ~n53315 & n53321 ;
  assign n53323 = ~n53318 & n53322 ;
  assign n53324 = n27308 & ~n53323 ;
  assign n53325 = ~n53313 & ~n53324 ;
  assign n53326 = \P2_P3_EAX_reg[6]/NET0131  & ~n42872 ;
  assign n53327 = ~n42542 & ~n53316 ;
  assign n53328 = \P2_P3_EAX_reg[6]/NET0131  & ~n53327 ;
  assign n53332 = \P2_P3_EAX_reg[6]/NET0131  & ~n27227 ;
  assign n53333 = \P2_buf2_reg[6]/NET0131  & n27227 ;
  assign n53334 = ~n53332 & ~n53333 ;
  assign n53335 = ~n27226 & ~n53334 ;
  assign n53329 = ~\P2_P3_EAX_reg[6]/NET0131  & n42837 ;
  assign n53330 = n42539 & n53329 ;
  assign n53331 = ~n32990 & n42538 ;
  assign n53336 = ~n53330 & ~n53331 ;
  assign n53337 = ~n53335 & n53336 ;
  assign n53338 = ~n53328 & n53337 ;
  assign n53339 = n27308 & ~n53338 ;
  assign n53340 = ~n53326 & ~n53339 ;
  assign n53341 = \P1_P2_EAX_reg[0]/NET0131  & ~n49627 ;
  assign n53344 = ~n46749 & n49630 ;
  assign n53342 = ~\P1_P2_EAX_reg[0]/NET0131  & n43164 ;
  assign n53343 = ~n31094 & n42875 ;
  assign n53345 = ~n53342 & ~n53343 ;
  assign n53346 = ~n53344 & n53345 ;
  assign n53347 = n25918 & ~n53346 ;
  assign n53348 = ~n53341 & ~n53347 ;
  assign n53349 = \P1_P2_EAX_reg[1]/NET0131  & ~n43212 ;
  assign n53350 = ~n43167 & ~n53342 ;
  assign n53351 = \P1_P2_EAX_reg[1]/NET0131  & ~n53350 ;
  assign n53355 = \P1_P2_EAX_reg[1]/NET0131  & ~n25773 ;
  assign n53356 = n25773 & ~n40746 ;
  assign n53357 = ~n53355 & ~n53356 ;
  assign n53358 = ~n25826 & ~n53357 ;
  assign n53352 = \P1_P2_EAX_reg[0]/NET0131  & ~\P1_P2_EAX_reg[1]/NET0131  ;
  assign n53353 = n43164 & n53352 ;
  assign n53354 = ~n31061 & n42875 ;
  assign n53359 = ~n53353 & ~n53354 ;
  assign n53360 = ~n53358 & n53359 ;
  assign n53361 = ~n53351 & n53360 ;
  assign n53362 = n25918 & ~n53361 ;
  assign n53363 = ~n53349 & ~n53362 ;
  assign n53365 = ~\P1_P2_EAX_reg[25]/NET0131  & ~n43194 ;
  assign n53366 = n43164 & ~n43195 ;
  assign n53367 = ~n53365 & n53366 ;
  assign n53364 = \P1_P2_EAX_reg[25]/NET0131  & ~n43169 ;
  assign n53368 = n25774 & ~n40754 ;
  assign n53369 = n25776 & ~n49721 ;
  assign n53370 = ~n53368 & ~n53369 ;
  assign n53371 = n25773 & ~n53370 ;
  assign n53372 = ~n42970 & n43001 ;
  assign n53373 = ~n43002 & ~n53372 ;
  assign n53374 = n42875 & n53373 ;
  assign n53375 = ~n53371 & ~n53374 ;
  assign n53376 = ~n53364 & n53375 ;
  assign n53377 = ~n53367 & n53376 ;
  assign n53378 = n25918 & ~n53377 ;
  assign n53379 = \P1_P2_EAX_reg[25]/NET0131  & ~n43212 ;
  assign n53380 = ~n53378 & ~n53379 ;
  assign n53381 = \P1_P2_EAX_reg[2]/NET0131  & ~n49627 ;
  assign n53383 = n25773 & ~n35963 ;
  assign n53384 = ~n25826 & n53383 ;
  assign n53382 = ~n31028 & n42875 ;
  assign n53385 = ~\P1_P2_EAX_reg[2]/NET0131  & ~n43171 ;
  assign n53386 = ~n43172 & ~n53385 ;
  assign n53387 = n43164 & n53386 ;
  assign n53388 = ~n53382 & ~n53387 ;
  assign n53389 = ~n53384 & n53388 ;
  assign n53390 = n25918 & ~n53389 ;
  assign n53391 = ~n53381 & ~n53390 ;
  assign n53392 = \P1_P2_EAX_reg[3]/NET0131  & ~n49627 ;
  assign n53394 = n25773 & ~n29832 ;
  assign n53395 = ~n25826 & n53394 ;
  assign n53393 = ~n30993 & n42875 ;
  assign n53396 = ~\P1_P2_EAX_reg[3]/NET0131  & ~n43172 ;
  assign n53397 = ~n43173 & ~n53396 ;
  assign n53398 = n43164 & n53397 ;
  assign n53399 = ~n53393 & ~n53398 ;
  assign n53400 = ~n53395 & n53399 ;
  assign n53401 = n25918 & ~n53400 ;
  assign n53402 = ~n53392 & ~n53401 ;
  assign n53403 = \P1_P2_EAX_reg[4]/NET0131  & ~n49627 ;
  assign n53405 = ~n27937 & n49630 ;
  assign n53404 = ~n30958 & n42875 ;
  assign n53406 = ~\P1_P2_EAX_reg[4]/NET0131  & ~n43173 ;
  assign n53407 = ~n43174 & ~n53406 ;
  assign n53408 = n43164 & n53407 ;
  assign n53409 = ~n53404 & ~n53408 ;
  assign n53410 = ~n53405 & n53409 ;
  assign n53411 = n25918 & ~n53410 ;
  assign n53412 = ~n53403 & ~n53411 ;
  assign n53413 = \P1_P2_EAX_reg[5]/NET0131  & ~n49627 ;
  assign n53415 = ~n29860 & n49630 ;
  assign n53414 = ~n30923 & n42875 ;
  assign n53416 = ~\P1_P2_EAX_reg[5]/NET0131  & ~n43174 ;
  assign n53417 = ~n43175 & ~n53416 ;
  assign n53418 = n43164 & n53417 ;
  assign n53419 = ~n53414 & ~n53418 ;
  assign n53420 = ~n53415 & n53419 ;
  assign n53421 = n25918 & ~n53420 ;
  assign n53422 = ~n53413 & ~n53421 ;
  assign n53423 = \P1_P2_EAX_reg[6]/NET0131  & ~n49627 ;
  assign n53425 = ~n34449 & n49630 ;
  assign n53424 = ~n30888 & n42875 ;
  assign n53426 = ~\P1_P2_EAX_reg[6]/NET0131  & ~n43175 ;
  assign n53427 = ~n43176 & ~n53426 ;
  assign n53428 = n43164 & n53427 ;
  assign n53429 = ~n53424 & ~n53428 ;
  assign n53430 = ~n53425 & n53429 ;
  assign n53431 = n25918 & ~n53430 ;
  assign n53432 = ~n53423 & ~n53431 ;
  assign n53433 = \P2_P3_uWord_reg[4]/NET0131  & ~n47752 ;
  assign n53434 = \P2_buf2_reg[4]/NET0131  & n27227 ;
  assign n53435 = n27122 & n53434 ;
  assign n53436 = ~n53040 & ~n53435 ;
  assign n53437 = n27308 & ~n53436 ;
  assign n53438 = ~n53433 & ~n53437 ;
  assign n53440 = n25761 & ~n25770 ;
  assign n53441 = \P1_P2_MemoryFetch_reg/NET0131  & ~n53440 ;
  assign n53442 = n47571 & ~n53441 ;
  assign n53443 = n25918 & ~n53442 ;
  assign n53439 = \P1_P2_MemoryFetch_reg/NET0131  & ~n47528 ;
  assign n53444 = n27968 & ~n53439 ;
  assign n53445 = ~n53443 & n53444 ;
  assign n53447 = \P2_P1_MemoryFetch_reg/NET0131  & ~n21087 ;
  assign n53448 = n24902 & ~n53447 ;
  assign n53449 = n11623 & ~n53448 ;
  assign n53446 = \P2_P1_MemoryFetch_reg/NET0131  & ~n24912 ;
  assign n53450 = n11619 & ~n53446 ;
  assign n53451 = ~n53449 & n53450 ;
  assign n53453 = \P1_P2_ReadRequest_reg/NET0131  & ~n25877 ;
  assign n53454 = ~n25875 & ~n53453 ;
  assign n53455 = n25918 & ~n53454 ;
  assign n53452 = \P1_P2_ReadRequest_reg/NET0131  & ~n47528 ;
  assign n53456 = n27968 & ~n53452 ;
  assign n53457 = ~n53455 & n53456 ;
  assign n53459 = \P2_P1_ReadRequest_reg/NET0131  & ~n25953 ;
  assign n53460 = ~n25949 & ~n53459 ;
  assign n53461 = n11623 & ~n53460 ;
  assign n53458 = \P2_P1_ReadRequest_reg/NET0131  & ~n24912 ;
  assign n53462 = n11619 & ~n53458 ;
  assign n53463 = ~n53461 & n53462 ;
  assign n53467 = n36672 & ~n50752 ;
  assign n53469 = ~n39461 & n53467 ;
  assign n53468 = n39461 & ~n53467 ;
  assign n53470 = ~\P2_P1_DataWidth_reg[1]/NET0131  & ~n53468 ;
  assign n53471 = ~n53469 & n53470 ;
  assign n53466 = \P2_P1_DataWidth_reg[1]/NET0131  & ~\P2_P1_rEIP_reg[15]/NET0131  ;
  assign n53472 = n11609 & ~n53466 ;
  assign n53473 = ~n53471 & n53472 ;
  assign n53478 = \P2_P1_EBX_reg[31]/NET0131  & ~n50800 ;
  assign n53480 = ~\P2_P1_EBX_reg[15]/NET0131  & n53478 ;
  assign n53479 = \P2_P1_EBX_reg[15]/NET0131  & ~n53478 ;
  assign n53481 = ~n50422 & ~n53479 ;
  assign n53482 = ~n53480 & n53481 ;
  assign n53474 = \P2_P1_rEIP_reg[15]/NET0131  & n50775 ;
  assign n53475 = ~\P2_P1_rEIP_reg[15]/NET0131  & ~n50775 ;
  assign n53476 = ~n53474 & ~n53475 ;
  assign n53477 = n50422 & ~n53476 ;
  assign n53483 = n24901 & ~n53477 ;
  assign n53484 = ~n53482 & n53483 ;
  assign n53485 = \P2_P1_rEIP_reg[15]/NET0131  & ~n50414 ;
  assign n53487 = ~n25958 & n53477 ;
  assign n53486 = ~\P2_P1_EBX_reg[15]/NET0131  & ~n26103 ;
  assign n53488 = n24899 & ~n53486 ;
  assign n53489 = ~n53487 & n53488 ;
  assign n53490 = ~n53485 & ~n53489 ;
  assign n53491 = ~n53484 & n53490 ;
  assign n53492 = n11623 & ~n53491 ;
  assign n53464 = n25941 & n27787 ;
  assign n53465 = \P2_P1_rEIP_reg[15]/NET0131  & ~n53464 ;
  assign n53493 = \P2_P1_PhyAddrPointer_reg[15]/NET0131  & n11625 ;
  assign n53494 = ~n11616 & ~n53493 ;
  assign n53495 = ~n53465 & n53494 ;
  assign n53496 = ~n53492 & n53495 ;
  assign n53497 = ~n53473 & n53496 ;
  assign n53500 = ~\P2_P1_PhyAddrPointer_reg[0]/NET0131  & n43475 ;
  assign n53501 = n36672 & ~n53500 ;
  assign n53503 = ~n43493 & n53501 ;
  assign n53502 = n43493 & ~n53501 ;
  assign n53504 = ~\P2_P1_DataWidth_reg[1]/NET0131  & ~n53502 ;
  assign n53505 = ~n53503 & n53504 ;
  assign n53499 = \P2_P1_DataWidth_reg[1]/NET0131  & ~\P2_P1_rEIP_reg[17]/NET0131  ;
  assign n53506 = n11609 & ~n53499 ;
  assign n53507 = ~n53505 & n53506 ;
  assign n53510 = n50763 & n50775 ;
  assign n53511 = ~\P2_P1_rEIP_reg[17]/NET0131  & ~n53510 ;
  assign n53512 = n50422 & ~n50776 ;
  assign n53513 = ~n53511 & n53512 ;
  assign n53517 = \P2_P1_EBX_reg[31]/NET0131  & ~n50802 ;
  assign n53519 = ~\P2_P1_EBX_reg[17]/NET0131  & ~n53517 ;
  assign n53518 = \P2_P1_EBX_reg[17]/NET0131  & n53517 ;
  assign n53520 = ~n50422 & ~n53518 ;
  assign n53521 = ~n53519 & n53520 ;
  assign n53522 = ~n53513 & ~n53521 ;
  assign n53523 = n24901 & ~n53522 ;
  assign n53508 = \P2_P1_rEIP_reg[17]/NET0131  & ~n50414 ;
  assign n53509 = \P2_P1_EBX_reg[17]/NET0131  & ~n26103 ;
  assign n53514 = ~n25958 & n53513 ;
  assign n53515 = ~n53509 & ~n53514 ;
  assign n53516 = n24899 & ~n53515 ;
  assign n53524 = ~n53508 & ~n53516 ;
  assign n53525 = ~n53523 & n53524 ;
  assign n53526 = n11623 & ~n53525 ;
  assign n53498 = \P2_P1_rEIP_reg[17]/NET0131  & ~n53464 ;
  assign n53527 = \P2_P1_PhyAddrPointer_reg[17]/NET0131  & n11625 ;
  assign n53528 = ~n11616 & ~n53527 ;
  assign n53529 = ~n53498 & n53528 ;
  assign n53530 = ~n53526 & n53529 ;
  assign n53531 = ~n53507 & n53530 ;
  assign n53534 = n36654 & n50753 ;
  assign n53535 = n36672 & ~n53534 ;
  assign n53537 = ~n43501 & n53535 ;
  assign n53536 = n43501 & ~n53535 ;
  assign n53538 = ~\P2_P1_DataWidth_reg[1]/NET0131  & ~n53536 ;
  assign n53539 = ~n53537 & n53538 ;
  assign n53533 = \P2_P1_DataWidth_reg[1]/NET0131  & ~\P2_P1_rEIP_reg[18]/NET0131  ;
  assign n53540 = n11609 & ~n53533 ;
  assign n53541 = ~n53539 & n53540 ;
  assign n53550 = \P2_P1_EBX_reg[31]/NET0131  & ~n50803 ;
  assign n53552 = ~\P2_P1_EBX_reg[18]/NET0131  & n53550 ;
  assign n53551 = \P2_P1_EBX_reg[18]/NET0131  & ~n53550 ;
  assign n53553 = ~n50422 & ~n53551 ;
  assign n53554 = ~n53552 & n53553 ;
  assign n53544 = ~\P2_P1_rEIP_reg[18]/NET0131  & ~n50776 ;
  assign n53545 = ~n50777 & ~n53544 ;
  assign n53546 = n50422 & ~n53545 ;
  assign n53555 = n24901 & ~n53546 ;
  assign n53556 = ~n53554 & n53555 ;
  assign n53542 = \P2_P1_rEIP_reg[18]/NET0131  & ~n50414 ;
  assign n53547 = ~n25958 & n53546 ;
  assign n53543 = ~\P2_P1_EBX_reg[18]/NET0131  & ~n26103 ;
  assign n53548 = n24899 & ~n53543 ;
  assign n53549 = ~n53547 & n53548 ;
  assign n53557 = ~n53542 & ~n53549 ;
  assign n53558 = ~n53556 & n53557 ;
  assign n53559 = n11623 & ~n53558 ;
  assign n53532 = \P2_P1_rEIP_reg[18]/NET0131  & ~n53464 ;
  assign n53560 = \P2_P1_PhyAddrPointer_reg[18]/NET0131  & n11625 ;
  assign n53561 = ~n11616 & ~n53560 ;
  assign n53562 = ~n53532 & n53561 ;
  assign n53563 = ~n53559 & n53562 ;
  assign n53564 = ~n53541 & n53563 ;
  assign n53569 = ~\P1_P2_PhyAddrPointer_reg[14]/NET0131  & ~n36628 ;
  assign n53570 = ~n36628 & ~n41393 ;
  assign n53571 = ~n51181 & ~n53570 ;
  assign n53572 = ~n53569 & n53571 ;
  assign n53574 = n39337 & n53572 ;
  assign n53573 = ~n39337 & ~n53572 ;
  assign n53575 = ~\P1_P2_DataWidth_reg[1]/NET0131  & ~n53573 ;
  assign n53576 = ~n53574 & n53575 ;
  assign n53568 = \P1_P2_DataWidth_reg[1]/NET0131  & ~\P1_P2_rEIP_reg[15]/NET0131  ;
  assign n53577 = n25928 & ~n53568 ;
  assign n53578 = ~n53576 & n53577 ;
  assign n53583 = \P1_P2_EBX_reg[31]/NET0131  & ~n48420 ;
  assign n53585 = ~\P1_P2_EBX_reg[15]/NET0131  & n53583 ;
  assign n53584 = \P1_P2_EBX_reg[15]/NET0131  & ~n53583 ;
  assign n53586 = ~n48373 & ~n53584 ;
  assign n53587 = ~n53585 & n53586 ;
  assign n53579 = n48386 & n48394 ;
  assign n53580 = ~\P1_P2_rEIP_reg[15]/NET0131  & ~n53579 ;
  assign n53581 = ~n51201 & ~n53580 ;
  assign n53582 = n48373 & ~n53581 ;
  assign n53588 = n25776 & ~n53582 ;
  assign n53589 = ~n53587 & n53588 ;
  assign n53590 = ~\P1_P2_EBX_reg[15]/NET0131  & ~n48443 ;
  assign n53591 = n48443 & ~n53581 ;
  assign n53592 = ~n53590 & ~n53591 ;
  assign n53593 = n25757 & n53592 ;
  assign n53594 = ~n53589 & ~n53593 ;
  assign n53595 = ~n25770 & ~n53594 ;
  assign n53596 = \P1_P2_rEIP_reg[15]/NET0131  & ~n48371 ;
  assign n53597 = ~n53595 & ~n53596 ;
  assign n53598 = n25918 & ~n53597 ;
  assign n53565 = ~n25935 & ~n27608 ;
  assign n53566 = n43209 & n53565 ;
  assign n53567 = \P1_P2_rEIP_reg[15]/NET0131  & ~n53566 ;
  assign n53599 = \P1_P2_PhyAddrPointer_reg[15]/NET0131  & n27675 ;
  assign n53600 = ~n27967 & ~n53599 ;
  assign n53601 = ~n53567 & n53600 ;
  assign n53602 = ~n53598 & n53601 ;
  assign n53603 = ~n53578 & n53602 ;
  assign n53606 = ~n36628 & ~n51389 ;
  assign n53608 = ~n43360 & n53606 ;
  assign n53607 = n43360 & ~n53606 ;
  assign n53609 = ~\P1_P2_DataWidth_reg[1]/NET0131  & ~n53607 ;
  assign n53610 = ~n53608 & n53609 ;
  assign n53605 = \P1_P2_DataWidth_reg[1]/NET0131  & ~\P1_P2_rEIP_reg[17]/NET0131  ;
  assign n53611 = n25928 & ~n53605 ;
  assign n53612 = ~n53610 & n53611 ;
  assign n53617 = \P1_P2_EBX_reg[31]/NET0131  & ~n48422 ;
  assign n53619 = ~\P1_P2_EBX_reg[17]/NET0131  & n53617 ;
  assign n53618 = \P1_P2_EBX_reg[17]/NET0131  & ~n53617 ;
  assign n53620 = ~n48373 & ~n53618 ;
  assign n53621 = ~n53619 & n53620 ;
  assign n53614 = ~\P1_P2_rEIP_reg[17]/NET0131  & ~n51242 ;
  assign n53615 = ~n51243 & ~n53614 ;
  assign n53616 = n48373 & ~n53615 ;
  assign n53622 = n25846 & ~n53616 ;
  assign n53623 = ~n53621 & n53622 ;
  assign n53613 = \P1_P2_rEIP_reg[17]/NET0131  & ~n48371 ;
  assign n53624 = n48443 & ~n53615 ;
  assign n53625 = ~\P1_P2_EBX_reg[17]/NET0131  & ~n48443 ;
  assign n53626 = n47570 & ~n53625 ;
  assign n53627 = ~n53624 & n53626 ;
  assign n53628 = ~n53613 & ~n53627 ;
  assign n53629 = ~n53623 & n53628 ;
  assign n53630 = n25918 & ~n53629 ;
  assign n53604 = \P1_P2_rEIP_reg[17]/NET0131  & ~n53566 ;
  assign n53631 = \P1_P2_PhyAddrPointer_reg[17]/NET0131  & n27675 ;
  assign n53632 = ~n27967 & ~n53631 ;
  assign n53633 = ~n53604 & n53632 ;
  assign n53634 = ~n53630 & n53633 ;
  assign n53635 = ~n53612 & n53634 ;
  assign n53638 = ~n36628 & ~n43359 ;
  assign n53639 = ~n51181 & ~n53638 ;
  assign n53641 = ~n43371 & ~n53639 ;
  assign n53640 = n43371 & n53639 ;
  assign n53642 = ~\P1_P2_DataWidth_reg[1]/NET0131  & ~n53640 ;
  assign n53643 = ~n53641 & n53642 ;
  assign n53637 = \P1_P2_DataWidth_reg[1]/NET0131  & ~\P1_P2_rEIP_reg[18]/NET0131  ;
  assign n53644 = n25928 & ~n53637 ;
  assign n53645 = ~n53643 & n53644 ;
  assign n53650 = \P1_P2_EBX_reg[31]/NET0131  & ~n48423 ;
  assign n53652 = ~\P1_P2_EBX_reg[18]/NET0131  & n53650 ;
  assign n53651 = \P1_P2_EBX_reg[18]/NET0131  & ~n53650 ;
  assign n53653 = ~n48373 & ~n53651 ;
  assign n53654 = ~n53652 & n53653 ;
  assign n53647 = ~\P1_P2_rEIP_reg[18]/NET0131  & ~n51243 ;
  assign n53648 = ~n48396 & ~n53647 ;
  assign n53649 = n48373 & ~n53648 ;
  assign n53655 = n25846 & ~n53649 ;
  assign n53656 = ~n53654 & n53655 ;
  assign n53646 = \P1_P2_rEIP_reg[18]/NET0131  & ~n48371 ;
  assign n53658 = n48443 & ~n53648 ;
  assign n53657 = ~\P1_P2_EBX_reg[18]/NET0131  & ~n48443 ;
  assign n53659 = n47570 & ~n53657 ;
  assign n53660 = ~n53658 & n53659 ;
  assign n53661 = ~n53646 & ~n53660 ;
  assign n53662 = ~n53656 & n53661 ;
  assign n53663 = n25918 & ~n53662 ;
  assign n53636 = \P1_P2_rEIP_reg[18]/NET0131  & ~n53566 ;
  assign n53664 = \P1_P2_PhyAddrPointer_reg[18]/NET0131  & n27675 ;
  assign n53665 = ~n27967 & ~n53664 ;
  assign n53666 = ~n53636 & n53665 ;
  assign n53667 = ~n53663 & n53666 ;
  assign n53668 = ~n53645 & n53667 ;
  assign n53671 = n36643 & n50476 ;
  assign n53672 = n36672 & ~n53671 ;
  assign n53674 = n47411 & ~n53672 ;
  assign n53673 = ~n47411 & n53672 ;
  assign n53675 = ~\P2_P1_DataWidth_reg[1]/NET0131  & ~n53673 ;
  assign n53676 = ~n53674 & n53675 ;
  assign n53670 = \P2_P1_DataWidth_reg[1]/NET0131  & ~\P2_P1_rEIP_reg[4]/NET0131  ;
  assign n53677 = n11609 & ~n53670 ;
  assign n53678 = ~n53676 & n53677 ;
  assign n53679 = \P2_P1_rEIP_reg[4]/NET0131  & ~n50414 ;
  assign n53680 = \P2_P1_EBX_reg[31]/NET0131  & ~n50789 ;
  assign n53682 = ~\P2_P1_EBX_reg[4]/NET0131  & n53680 ;
  assign n53681 = \P2_P1_EBX_reg[4]/NET0131  & ~n53680 ;
  assign n53683 = ~n50422 & ~n53681 ;
  assign n53684 = ~n53682 & n53683 ;
  assign n53685 = ~\P2_P1_rEIP_reg[4]/NET0131  & ~n50495 ;
  assign n53686 = ~n50766 & ~n53685 ;
  assign n53687 = n50422 & ~n53686 ;
  assign n53688 = ~n53684 & ~n53687 ;
  assign n53689 = n24901 & n53688 ;
  assign n53690 = ~\P2_P1_EBX_reg[4]/NET0131  & ~n26103 ;
  assign n53691 = n26103 & ~n53686 ;
  assign n53692 = ~n53690 & ~n53691 ;
  assign n53693 = n24899 & n53692 ;
  assign n53694 = ~n53689 & ~n53693 ;
  assign n53695 = ~n53679 & n53694 ;
  assign n53696 = n11623 & ~n53695 ;
  assign n53669 = \P2_P1_rEIP_reg[4]/NET0131  & ~n53464 ;
  assign n53697 = \P2_P1_PhyAddrPointer_reg[4]/NET0131  & n11625 ;
  assign n53698 = ~n11616 & ~n53697 ;
  assign n53699 = ~n53669 & n53698 ;
  assign n53700 = ~n53696 & n53699 ;
  assign n53701 = ~n53678 & n53700 ;
  assign n53703 = \P1_P1_MemoryFetch_reg/NET0131  & ~n15724 ;
  assign n53704 = n24505 & ~n53703 ;
  assign n53705 = n8355 & ~n53704 ;
  assign n53702 = \P1_P1_MemoryFetch_reg/NET0131  & ~n24514 ;
  assign n53706 = n8360 & ~n53702 ;
  assign n53707 = ~n53705 & n53706 ;
  assign n53710 = ~\P2_P1_PhyAddrPointer_reg[0]/NET0131  & n47878 ;
  assign n53711 = n36672 & ~n53710 ;
  assign n53713 = n47891 & ~n53711 ;
  assign n53712 = ~n47891 & n53711 ;
  assign n53714 = ~\P2_P1_DataWidth_reg[1]/NET0131  & ~n53712 ;
  assign n53715 = ~n53713 & n53714 ;
  assign n53709 = \P2_P1_DataWidth_reg[1]/NET0131  & ~\P2_P1_rEIP_reg[6]/NET0131  ;
  assign n53716 = n11609 & ~n53709 ;
  assign n53717 = ~n53715 & n53716 ;
  assign n53718 = \P2_P1_rEIP_reg[6]/NET0131  & ~n50414 ;
  assign n53719 = ~\P2_P1_EBX_reg[6]/NET0131  & ~n26103 ;
  assign n53720 = ~\P2_P1_rEIP_reg[6]/NET0131  & ~n50767 ;
  assign n53721 = ~n50768 & ~n53720 ;
  assign n53722 = n26103 & ~n53721 ;
  assign n53723 = ~n53719 & ~n53722 ;
  assign n53724 = n24899 & n53723 ;
  assign n53725 = n50422 & ~n53721 ;
  assign n53726 = \P2_P1_EBX_reg[31]/NET0131  & ~n50791 ;
  assign n53728 = ~\P2_P1_EBX_reg[6]/NET0131  & n53726 ;
  assign n53727 = \P2_P1_EBX_reg[6]/NET0131  & ~n53726 ;
  assign n53729 = ~n50422 & ~n53727 ;
  assign n53730 = ~n53728 & n53729 ;
  assign n53731 = ~n53725 & ~n53730 ;
  assign n53732 = n24901 & n53731 ;
  assign n53733 = ~n53724 & ~n53732 ;
  assign n53734 = ~n53718 & n53733 ;
  assign n53735 = n11623 & ~n53734 ;
  assign n53708 = \P2_P1_rEIP_reg[6]/NET0131  & ~n53464 ;
  assign n53736 = \P2_P1_PhyAddrPointer_reg[6]/NET0131  & n11625 ;
  assign n53737 = ~n11616 & ~n53736 ;
  assign n53738 = ~n53708 & n53737 ;
  assign n53739 = ~n53735 & n53738 ;
  assign n53740 = ~n53717 & n53739 ;
  assign n53743 = \P2_P1_PhyAddrPointer_reg[6]/NET0131  & n53710 ;
  assign n53744 = n36672 & ~n53743 ;
  assign n53746 = n44962 & ~n53744 ;
  assign n53745 = ~n44962 & n53744 ;
  assign n53747 = ~\P2_P1_DataWidth_reg[1]/NET0131  & ~n53745 ;
  assign n53748 = ~n53746 & n53747 ;
  assign n53742 = \P2_P1_DataWidth_reg[1]/NET0131  & ~\P2_P1_rEIP_reg[7]/NET0131  ;
  assign n53749 = n11609 & ~n53742 ;
  assign n53750 = ~n53748 & n53749 ;
  assign n53751 = \P2_P1_rEIP_reg[7]/NET0131  & ~n50414 ;
  assign n53752 = ~\P2_P1_EBX_reg[7]/NET0131  & ~n26103 ;
  assign n53753 = ~\P2_P1_rEIP_reg[7]/NET0131  & ~n50768 ;
  assign n53754 = ~n50769 & ~n53753 ;
  assign n53755 = n26103 & ~n53754 ;
  assign n53756 = ~n53752 & ~n53755 ;
  assign n53757 = n24899 & n53756 ;
  assign n53758 = n50422 & ~n53754 ;
  assign n53759 = \P2_P1_EBX_reg[31]/NET0131  & ~n50792 ;
  assign n53761 = \P2_P1_EBX_reg[7]/NET0131  & ~n53759 ;
  assign n53760 = ~\P2_P1_EBX_reg[7]/NET0131  & n53759 ;
  assign n53762 = ~n50422 & ~n53760 ;
  assign n53763 = ~n53761 & n53762 ;
  assign n53764 = ~n53758 & ~n53763 ;
  assign n53765 = n24901 & n53764 ;
  assign n53766 = ~n53757 & ~n53765 ;
  assign n53767 = ~n53751 & n53766 ;
  assign n53768 = n11623 & ~n53767 ;
  assign n53741 = \P2_P1_rEIP_reg[7]/NET0131  & ~n53464 ;
  assign n53769 = \P2_P1_PhyAddrPointer_reg[7]/NET0131  & n11625 ;
  assign n53770 = ~n11616 & ~n53769 ;
  assign n53771 = ~n53741 & n53770 ;
  assign n53772 = ~n53768 & n53771 ;
  assign n53773 = ~n53750 & n53772 ;
  assign n53776 = \P1_P2_PhyAddrPointer_reg[3]/NET0131  & n50516 ;
  assign n53777 = ~n36628 & ~n53776 ;
  assign n53779 = ~n47388 & n53777 ;
  assign n53778 = n47388 & ~n53777 ;
  assign n53780 = ~\P1_P2_DataWidth_reg[1]/NET0131  & ~n53778 ;
  assign n53781 = ~n53779 & n53780 ;
  assign n53775 = \P1_P2_DataWidth_reg[1]/NET0131  & ~\P1_P2_rEIP_reg[4]/NET0131  ;
  assign n53782 = n25928 & ~n53775 ;
  assign n53783 = ~n53781 & n53782 ;
  assign n53784 = \P1_P2_rEIP_reg[4]/NET0131  & ~n48371 ;
  assign n53785 = ~\P1_P2_rEIP_reg[4]/NET0131  & ~n48381 ;
  assign n53786 = ~n48382 & ~n53785 ;
  assign n53787 = n48443 & ~n53786 ;
  assign n53788 = ~\P1_P2_EBX_reg[4]/NET0131  & ~n48443 ;
  assign n53789 = ~n53787 & ~n53788 ;
  assign n53790 = n25757 & n53789 ;
  assign n53791 = n48373 & ~n53786 ;
  assign n53792 = \P1_P2_EBX_reg[31]/NET0131  & ~n48409 ;
  assign n53794 = \P1_P2_EBX_reg[4]/NET0131  & ~n53792 ;
  assign n53793 = ~\P1_P2_EBX_reg[4]/NET0131  & n53792 ;
  assign n53795 = ~n48373 & ~n53793 ;
  assign n53796 = ~n53794 & n53795 ;
  assign n53797 = ~n53791 & ~n53796 ;
  assign n53798 = n25776 & n53797 ;
  assign n53799 = ~n53790 & ~n53798 ;
  assign n53800 = ~n25770 & ~n53799 ;
  assign n53801 = ~n53784 & ~n53800 ;
  assign n53802 = n25918 & ~n53801 ;
  assign n53774 = \P1_P2_rEIP_reg[4]/NET0131  & ~n53566 ;
  assign n53803 = \P1_P2_PhyAddrPointer_reg[4]/NET0131  & n27675 ;
  assign n53804 = ~n27967 & ~n53803 ;
  assign n53805 = ~n53774 & n53804 ;
  assign n53806 = ~n53802 & n53805 ;
  assign n53807 = ~n53783 & n53806 ;
  assign n53810 = ~\P1_P2_PhyAddrPointer_reg[0]/NET0131  & n47387 ;
  assign n53811 = \P1_P2_PhyAddrPointer_reg[5]/NET0131  & n53810 ;
  assign n53812 = ~n36628 & ~n53811 ;
  assign n53814 = n47836 & ~n53812 ;
  assign n53813 = ~n47836 & n53812 ;
  assign n53815 = ~\P1_P2_DataWidth_reg[1]/NET0131  & ~n53813 ;
  assign n53816 = ~n53814 & n53815 ;
  assign n53809 = \P1_P2_DataWidth_reg[1]/NET0131  & ~\P1_P2_rEIP_reg[6]/NET0131  ;
  assign n53817 = n25928 & ~n53809 ;
  assign n53818 = ~n53816 & n53817 ;
  assign n53819 = \P1_P2_rEIP_reg[6]/NET0131  & ~n48371 ;
  assign n53820 = ~\P1_P2_rEIP_reg[6]/NET0131  & ~n48383 ;
  assign n53821 = ~n48384 & ~n53820 ;
  assign n53822 = n48443 & ~n53821 ;
  assign n53823 = ~\P1_P2_EBX_reg[6]/NET0131  & ~n48443 ;
  assign n53824 = ~n53822 & ~n53823 ;
  assign n53825 = n25757 & n53824 ;
  assign n53826 = n48373 & ~n53821 ;
  assign n53827 = \P1_P2_EBX_reg[31]/NET0131  & ~n48411 ;
  assign n53829 = ~\P1_P2_EBX_reg[6]/NET0131  & n53827 ;
  assign n53828 = \P1_P2_EBX_reg[6]/NET0131  & ~n53827 ;
  assign n53830 = ~n48373 & ~n53828 ;
  assign n53831 = ~n53829 & n53830 ;
  assign n53832 = ~n53826 & ~n53831 ;
  assign n53833 = n25776 & n53832 ;
  assign n53834 = ~n53825 & ~n53833 ;
  assign n53835 = ~n25770 & ~n53834 ;
  assign n53836 = ~n53819 & ~n53835 ;
  assign n53837 = n25918 & ~n53836 ;
  assign n53808 = \P1_P2_rEIP_reg[6]/NET0131  & ~n53566 ;
  assign n53838 = \P1_P2_PhyAddrPointer_reg[6]/NET0131  & n27675 ;
  assign n53839 = ~n27967 & ~n53838 ;
  assign n53840 = ~n53808 & n53839 ;
  assign n53841 = ~n53837 & n53840 ;
  assign n53842 = ~n53818 & n53841 ;
  assign n53845 = ~\P1_P2_PhyAddrPointer_reg[6]/NET0131  & ~n36628 ;
  assign n53846 = ~n53812 & ~n53845 ;
  assign n53848 = n44912 & n53846 ;
  assign n53847 = ~n44912 & ~n53846 ;
  assign n53849 = ~\P1_P2_DataWidth_reg[1]/NET0131  & ~n53847 ;
  assign n53850 = ~n53848 & n53849 ;
  assign n53844 = \P1_P2_DataWidth_reg[1]/NET0131  & ~\P1_P2_rEIP_reg[7]/NET0131  ;
  assign n53851 = n25928 & ~n53844 ;
  assign n53852 = ~n53850 & n53851 ;
  assign n53853 = \P1_P2_rEIP_reg[7]/NET0131  & ~n48371 ;
  assign n53854 = ~\P1_P2_rEIP_reg[7]/NET0131  & ~n48384 ;
  assign n53855 = ~n48385 & ~n53854 ;
  assign n53856 = n48443 & ~n53855 ;
  assign n53857 = ~\P1_P2_EBX_reg[7]/NET0131  & ~n48443 ;
  assign n53858 = ~n53856 & ~n53857 ;
  assign n53859 = n25757 & n53858 ;
  assign n53860 = n48373 & ~n53855 ;
  assign n53861 = \P1_P2_EBX_reg[31]/NET0131  & ~n48412 ;
  assign n53863 = ~\P1_P2_EBX_reg[7]/NET0131  & n53861 ;
  assign n53862 = \P1_P2_EBX_reg[7]/NET0131  & ~n53861 ;
  assign n53864 = ~n48373 & ~n53862 ;
  assign n53865 = ~n53863 & n53864 ;
  assign n53866 = ~n53860 & ~n53865 ;
  assign n53867 = n25776 & n53866 ;
  assign n53868 = ~n53859 & ~n53867 ;
  assign n53869 = ~n25770 & ~n53868 ;
  assign n53870 = ~n53853 & ~n53869 ;
  assign n53871 = n25918 & ~n53870 ;
  assign n53843 = \P1_P2_rEIP_reg[7]/NET0131  & ~n53566 ;
  assign n53872 = \P1_P2_PhyAddrPointer_reg[7]/NET0131  & n27675 ;
  assign n53873 = ~n27967 & ~n53872 ;
  assign n53874 = ~n53843 & n53873 ;
  assign n53875 = ~n53871 & n53874 ;
  assign n53876 = ~n53852 & n53875 ;
  assign n53878 = \P1_P1_ReadRequest_reg/NET0131  & ~n26161 ;
  assign n53879 = ~n24341 & ~n53878 ;
  assign n53880 = n8355 & ~n53879 ;
  assign n53877 = \P1_P1_ReadRequest_reg/NET0131  & ~n24514 ;
  assign n53881 = n8360 & ~n53877 ;
  assign n53882 = ~n53880 & n53881 ;
  assign n53886 = n36713 & n52046 ;
  assign n53887 = ~n36733 & ~n53886 ;
  assign n53889 = ~n39562 & n53887 ;
  assign n53888 = n39562 & ~n53887 ;
  assign n53890 = ~\P1_P1_DataWidth_reg[1]/NET0131  & ~n53888 ;
  assign n53891 = ~n53889 & n53890 ;
  assign n53885 = \P1_P1_DataWidth_reg[1]/NET0131  & ~\P1_P1_rEIP_reg[15]/NET0131  ;
  assign n53892 = n8282 & ~n53885 ;
  assign n53893 = ~n53891 & n53892 ;
  assign n53894 = \P1_P1_rEIP_reg[15]/NET0131  & ~n50559 ;
  assign n53896 = ~\P1_P1_rEIP_reg[15]/NET0131  & ~n51677 ;
  assign n53897 = ~n51678 & ~n53896 ;
  assign n53898 = n26275 & ~n53897 ;
  assign n53895 = ~\P1_P1_EBX_reg[15]/NET0131  & ~n26275 ;
  assign n53899 = n24502 & ~n53895 ;
  assign n53900 = ~n53898 & n53899 ;
  assign n53902 = \P1_P1_EBX_reg[31]/NET0131  & ~n51699 ;
  assign n53904 = ~\P1_P1_EBX_reg[15]/NET0131  & n53902 ;
  assign n53903 = \P1_P1_EBX_reg[15]/NET0131  & ~n53902 ;
  assign n53905 = ~n26274 & ~n53903 ;
  assign n53906 = ~n53904 & n53905 ;
  assign n53901 = n26274 & ~n53897 ;
  assign n53907 = n15334 & ~n53901 ;
  assign n53908 = ~n53906 & n53907 ;
  assign n53909 = ~n53900 & ~n53908 ;
  assign n53910 = ~n15364 & ~n53909 ;
  assign n53911 = ~n53894 & ~n53910 ;
  assign n53912 = n8355 & ~n53911 ;
  assign n53883 = n26114 & n27611 ;
  assign n53884 = \P1_P1_rEIP_reg[15]/NET0131  & ~n53883 ;
  assign n53913 = \P1_P1_PhyAddrPointer_reg[15]/NET0131  & n8361 ;
  assign n53914 = ~n8357 & ~n53913 ;
  assign n53915 = ~n53884 & n53914 ;
  assign n53916 = ~n53912 & n53915 ;
  assign n53917 = ~n53893 & n53916 ;
  assign n53921 = n43665 & ~n51654 ;
  assign n53920 = ~n43665 & n51654 ;
  assign n53922 = ~\P1_P1_DataWidth_reg[1]/NET0131  & ~n53920 ;
  assign n53923 = ~n53921 & n53922 ;
  assign n53919 = \P1_P1_DataWidth_reg[1]/NET0131  & ~\P1_P1_rEIP_reg[17]/NET0131  ;
  assign n53924 = n8282 & ~n53919 ;
  assign n53925 = ~n53923 & n53924 ;
  assign n53926 = \P1_P1_rEIP_reg[17]/NET0131  & ~n50559 ;
  assign n53928 = \P1_P1_rEIP_reg[17]/NET0131  & n51679 ;
  assign n53929 = ~\P1_P1_rEIP_reg[17]/NET0131  & ~n51679 ;
  assign n53930 = ~n53928 & ~n53929 ;
  assign n53931 = n26275 & ~n53930 ;
  assign n53927 = ~\P1_P1_EBX_reg[17]/NET0131  & ~n26275 ;
  assign n53932 = n24502 & ~n53927 ;
  assign n53933 = ~n53931 & n53932 ;
  assign n53935 = \P1_P1_EBX_reg[31]/NET0131  & ~n51701 ;
  assign n53937 = ~\P1_P1_EBX_reg[17]/NET0131  & n53935 ;
  assign n53936 = \P1_P1_EBX_reg[17]/NET0131  & ~n53935 ;
  assign n53938 = ~n26274 & ~n53936 ;
  assign n53939 = ~n53937 & n53938 ;
  assign n53934 = n26274 & ~n53930 ;
  assign n53940 = n15334 & ~n53934 ;
  assign n53941 = ~n53939 & n53940 ;
  assign n53942 = ~n53933 & ~n53941 ;
  assign n53943 = ~n15364 & ~n53942 ;
  assign n53944 = ~n53926 & ~n53943 ;
  assign n53945 = n8355 & ~n53944 ;
  assign n53918 = \P1_P1_rEIP_reg[17]/NET0131  & ~n53883 ;
  assign n53946 = \P1_P1_PhyAddrPointer_reg[17]/NET0131  & n8361 ;
  assign n53947 = ~n8357 & ~n53946 ;
  assign n53948 = ~n53918 & n53947 ;
  assign n53949 = ~n53945 & n53948 ;
  assign n53950 = ~n53925 & n53949 ;
  assign n53954 = ~n43683 & n51763 ;
  assign n53953 = n43683 & ~n51763 ;
  assign n53955 = ~\P1_P1_DataWidth_reg[1]/NET0131  & ~n53953 ;
  assign n53956 = ~n53954 & n53955 ;
  assign n53952 = \P1_P1_DataWidth_reg[1]/NET0131  & ~\P1_P1_rEIP_reg[18]/NET0131  ;
  assign n53957 = n8282 & ~n53952 ;
  assign n53958 = ~n53956 & n53957 ;
  assign n53959 = \P1_P1_rEIP_reg[18]/NET0131  & ~n50559 ;
  assign n53961 = ~\P1_P1_rEIP_reg[18]/NET0131  & ~n53928 ;
  assign n53962 = n51665 & n51679 ;
  assign n53963 = ~n53961 & ~n53962 ;
  assign n53964 = n26274 & ~n53963 ;
  assign n53965 = ~n26158 & n53964 ;
  assign n53960 = ~\P1_P1_EBX_reg[18]/NET0131  & ~n26275 ;
  assign n53966 = n24502 & ~n53960 ;
  assign n53967 = ~n53965 & n53966 ;
  assign n53968 = \P1_P1_EBX_reg[31]/NET0131  & ~n51702 ;
  assign n53970 = ~\P1_P1_EBX_reg[18]/NET0131  & n53968 ;
  assign n53969 = \P1_P1_EBX_reg[18]/NET0131  & ~n53968 ;
  assign n53971 = ~n26274 & ~n53969 ;
  assign n53972 = ~n53970 & n53971 ;
  assign n53973 = n15334 & ~n53964 ;
  assign n53974 = ~n53972 & n53973 ;
  assign n53975 = ~n53967 & ~n53974 ;
  assign n53976 = ~n15364 & ~n53975 ;
  assign n53977 = ~n53959 & ~n53976 ;
  assign n53978 = n8355 & ~n53977 ;
  assign n53951 = \P1_P1_rEIP_reg[18]/NET0131  & ~n53883 ;
  assign n53979 = \P1_P1_PhyAddrPointer_reg[18]/NET0131  & n8361 ;
  assign n53980 = ~n8357 & ~n53979 ;
  assign n53981 = ~n53951 & n53980 ;
  assign n53982 = ~n53978 & n53981 ;
  assign n53983 = ~n53958 & n53982 ;
  assign n53986 = \P1_P1_PhyAddrPointer_reg[3]/NET0131  & n50590 ;
  assign n53987 = ~n36733 & ~n53986 ;
  assign n53989 = n47434 & ~n53987 ;
  assign n53988 = ~n47434 & n53987 ;
  assign n53990 = ~\P1_P1_DataWidth_reg[1]/NET0131  & ~n53988 ;
  assign n53991 = ~n53989 & n53990 ;
  assign n53985 = \P1_P1_DataWidth_reg[1]/NET0131  & ~\P1_P1_rEIP_reg[4]/NET0131  ;
  assign n53992 = n8282 & ~n53985 ;
  assign n53993 = ~n53991 & n53992 ;
  assign n53994 = \P1_P1_rEIP_reg[4]/NET0131  & ~n50559 ;
  assign n53995 = ~\P1_P1_rEIP_reg[4]/NET0131  & ~n50601 ;
  assign n53996 = ~n51668 & ~n53995 ;
  assign n53997 = n26275 & ~n53996 ;
  assign n53998 = ~\P1_P1_EBX_reg[4]/NET0131  & ~n26275 ;
  assign n53999 = ~n53997 & ~n53998 ;
  assign n54000 = n24502 & n53999 ;
  assign n54001 = n26274 & ~n53996 ;
  assign n54002 = \P1_P1_EBX_reg[31]/NET0131  & ~n51688 ;
  assign n54004 = \P1_P1_EBX_reg[4]/NET0131  & ~n54002 ;
  assign n54003 = ~\P1_P1_EBX_reg[4]/NET0131  & n54002 ;
  assign n54005 = ~n26274 & ~n54003 ;
  assign n54006 = ~n54004 & n54005 ;
  assign n54007 = ~n54001 & ~n54006 ;
  assign n54008 = n15334 & n54007 ;
  assign n54009 = ~n54000 & ~n54008 ;
  assign n54010 = ~n15364 & ~n54009 ;
  assign n54011 = ~n53994 & ~n54010 ;
  assign n54012 = n8355 & ~n54011 ;
  assign n53984 = \P1_P1_rEIP_reg[4]/NET0131  & ~n53883 ;
  assign n54013 = \P1_P1_PhyAddrPointer_reg[4]/NET0131  & n8361 ;
  assign n54014 = ~n8357 & ~n54013 ;
  assign n54015 = ~n53984 & n54014 ;
  assign n54016 = ~n54012 & n54015 ;
  assign n54017 = ~n53993 & n54016 ;
  assign n54020 = n36704 & n52046 ;
  assign n54021 = ~n36733 & ~n54020 ;
  assign n54023 = n47951 & ~n54021 ;
  assign n54022 = ~n47951 & n54021 ;
  assign n54024 = ~\P1_P1_DataWidth_reg[1]/NET0131  & ~n54022 ;
  assign n54025 = ~n54023 & n54024 ;
  assign n54019 = \P1_P1_DataWidth_reg[1]/NET0131  & ~\P1_P1_rEIP_reg[6]/NET0131  ;
  assign n54026 = n8282 & ~n54019 ;
  assign n54027 = ~n54025 & n54026 ;
  assign n54028 = \P1_P1_rEIP_reg[6]/NET0131  & ~n50559 ;
  assign n54029 = ~\P1_P1_EBX_reg[6]/NET0131  & ~n26275 ;
  assign n54030 = ~\P1_P1_rEIP_reg[6]/NET0131  & ~n51669 ;
  assign n54031 = ~n51670 & ~n54030 ;
  assign n54032 = n26274 & ~n54031 ;
  assign n54033 = ~n26158 & n54032 ;
  assign n54034 = ~n54029 & ~n54033 ;
  assign n54035 = n24502 & n54034 ;
  assign n54036 = \P1_P1_EBX_reg[31]/NET0131  & ~n51690 ;
  assign n54038 = ~\P1_P1_EBX_reg[6]/NET0131  & n54036 ;
  assign n54037 = \P1_P1_EBX_reg[6]/NET0131  & ~n54036 ;
  assign n54039 = ~n26274 & ~n54037 ;
  assign n54040 = ~n54038 & n54039 ;
  assign n54041 = ~n54032 & ~n54040 ;
  assign n54042 = n15334 & n54041 ;
  assign n54043 = ~n54035 & ~n54042 ;
  assign n54044 = ~n15364 & ~n54043 ;
  assign n54045 = ~n54028 & ~n54044 ;
  assign n54046 = n8355 & ~n54045 ;
  assign n54018 = \P1_P1_rEIP_reg[6]/NET0131  & ~n53883 ;
  assign n54047 = \P1_P1_PhyAddrPointer_reg[6]/NET0131  & n8361 ;
  assign n54048 = ~n8357 & ~n54047 ;
  assign n54049 = ~n54018 & n54048 ;
  assign n54050 = ~n54046 & n54049 ;
  assign n54051 = ~n54027 & n54050 ;
  assign n54053 = \P2_P2_MemoryFetch_reg/NET0131  & ~n50638 ;
  assign n54054 = n47685 & ~n54053 ;
  assign n54055 = n26792 & ~n54054 ;
  assign n54052 = \P2_P2_MemoryFetch_reg/NET0131  & ~n47641 ;
  assign n54056 = n45044 & ~n54052 ;
  assign n54057 = ~n54055 & n54056 ;
  assign n54080 = n36705 & n52046 ;
  assign n54081 = ~n36733 & ~n54080 ;
  assign n54082 = ~n45018 & ~n54081 ;
  assign n54083 = n45018 & n54081 ;
  assign n54084 = ~n54082 & ~n54083 ;
  assign n54085 = ~\P1_P1_DataWidth_reg[1]/NET0131  & ~n54084 ;
  assign n54079 = \P1_P1_DataWidth_reg[1]/NET0131  & ~\P1_P1_rEIP_reg[7]/NET0131  ;
  assign n54086 = n8282 & ~n54079 ;
  assign n54087 = ~n54085 & n54086 ;
  assign n54059 = \P1_P1_rEIP_reg[7]/NET0131  & ~n50559 ;
  assign n54060 = ~\P1_P1_rEIP_reg[7]/NET0131  & ~n51670 ;
  assign n54061 = ~n51671 & ~n54060 ;
  assign n54062 = n26275 & ~n54061 ;
  assign n54063 = ~\P1_P1_EBX_reg[7]/NET0131  & ~n26275 ;
  assign n54064 = ~n54062 & ~n54063 ;
  assign n54065 = n24502 & n54064 ;
  assign n54066 = n26274 & ~n54061 ;
  assign n54067 = \P1_P1_EBX_reg[31]/NET0131  & ~n51691 ;
  assign n54069 = \P1_P1_EBX_reg[7]/NET0131  & ~n54067 ;
  assign n54068 = ~\P1_P1_EBX_reg[7]/NET0131  & n54067 ;
  assign n54070 = ~n26274 & ~n54068 ;
  assign n54071 = ~n54069 & n54070 ;
  assign n54072 = ~n54066 & ~n54071 ;
  assign n54073 = n15334 & n54072 ;
  assign n54074 = ~n54065 & ~n54073 ;
  assign n54075 = ~n15364 & ~n54074 ;
  assign n54076 = ~n54059 & ~n54075 ;
  assign n54077 = n8355 & ~n54076 ;
  assign n54058 = \P1_P1_rEIP_reg[7]/NET0131  & ~n53883 ;
  assign n54078 = \P1_P1_PhyAddrPointer_reg[7]/NET0131  & n8361 ;
  assign n54088 = ~n8357 & ~n54078 ;
  assign n54089 = ~n54058 & n54088 ;
  assign n54090 = ~n54077 & n54089 ;
  assign n54091 = ~n54087 & n54090 ;
  assign n54093 = \P2_P2_ReadRequest_reg/NET0131  & ~n26698 ;
  assign n54094 = ~n26697 & ~n54093 ;
  assign n54095 = n26792 & ~n54094 ;
  assign n54092 = \P2_P2_ReadRequest_reg/NET0131  & ~n47641 ;
  assign n54096 = n45044 & ~n54092 ;
  assign n54097 = ~n54095 & n54096 ;
  assign n54102 = n36792 & ~n52085 ;
  assign n54104 = n39652 & ~n54102 ;
  assign n54103 = ~n39652 & n54102 ;
  assign n54105 = ~\P2_P2_DataWidth_reg[1]/NET0131  & ~n54103 ;
  assign n54106 = ~n54104 & n54105 ;
  assign n54101 = \P2_P2_DataWidth_reg[1]/NET0131  & ~\P2_P2_rEIP_reg[15]/NET0131  ;
  assign n54107 = n26794 & ~n54101 ;
  assign n54108 = ~n54106 & n54107 ;
  assign n54109 = \P2_P2_rEIP_reg[15]/NET0131  & ~n50640 ;
  assign n54111 = n52099 & n52108 ;
  assign n54112 = \P2_P2_rEIP_reg[15]/NET0131  & n54111 ;
  assign n54113 = ~\P2_P2_rEIP_reg[15]/NET0131  & ~n54111 ;
  assign n54114 = ~n54112 & ~n54113 ;
  assign n54115 = n50642 & ~n54114 ;
  assign n54110 = ~\P2_P2_EBX_reg[15]/NET0131  & ~n50642 ;
  assign n54116 = n26643 & ~n54110 ;
  assign n54117 = ~n54115 & n54116 ;
  assign n54119 = \P2_P2_EBX_reg[31]/NET0131  & ~n52126 ;
  assign n54121 = \P2_P2_EBX_reg[15]/NET0131  & ~n54119 ;
  assign n54120 = ~\P2_P2_EBX_reg[15]/NET0131  & n54119 ;
  assign n54122 = ~n50649 & ~n54120 ;
  assign n54123 = ~n54121 & n54122 ;
  assign n54118 = n50649 & ~n54114 ;
  assign n54124 = n26633 & ~n54118 ;
  assign n54125 = ~n54123 & n54124 ;
  assign n54126 = ~n54117 & ~n54125 ;
  assign n54127 = ~n26640 & ~n54126 ;
  assign n54128 = ~n54109 & ~n54127 ;
  assign n54129 = n26792 & ~n54128 ;
  assign n54098 = n27616 & ~n27635 ;
  assign n54099 = ~n26802 & n54098 ;
  assign n54100 = \P2_P2_rEIP_reg[15]/NET0131  & ~n54099 ;
  assign n54130 = \P2_P2_PhyAddrPointer_reg[15]/NET0131  & n27637 ;
  assign n54131 = ~n28046 & ~n54130 ;
  assign n54132 = ~n54100 & n54131 ;
  assign n54133 = ~n54129 & n54132 ;
  assign n54134 = ~n54108 & n54133 ;
  assign n54137 = n36774 & n52152 ;
  assign n54138 = n36792 & ~n54137 ;
  assign n54140 = ~n43814 & n54138 ;
  assign n54139 = n43814 & ~n54138 ;
  assign n54141 = ~\P2_P2_DataWidth_reg[1]/NET0131  & ~n54139 ;
  assign n54142 = ~n54140 & n54141 ;
  assign n54136 = \P2_P2_DataWidth_reg[1]/NET0131  & ~\P2_P2_rEIP_reg[17]/NET0131  ;
  assign n54143 = n26794 & ~n54136 ;
  assign n54144 = ~n54142 & n54143 ;
  assign n54145 = \P2_P2_rEIP_reg[17]/NET0131  & ~n50640 ;
  assign n54150 = ~\P2_P2_EBX_reg[17]/NET0131  & ~n50642 ;
  assign n54151 = n26643 & ~n54150 ;
  assign n54155 = \P2_P2_EBX_reg[31]/NET0131  & ~n52128 ;
  assign n54157 = ~\P2_P2_EBX_reg[17]/NET0131  & n54155 ;
  assign n54156 = \P2_P2_EBX_reg[17]/NET0131  & ~n54155 ;
  assign n54158 = ~n50649 & ~n54156 ;
  assign n54159 = ~n54157 & n54158 ;
  assign n54160 = n26633 & ~n54159 ;
  assign n54161 = ~n54151 & ~n54160 ;
  assign n54152 = n26650 & n54151 ;
  assign n54146 = n52100 & n54111 ;
  assign n54147 = ~\P2_P2_rEIP_reg[17]/NET0131  & ~n54146 ;
  assign n54148 = n52101 & n54111 ;
  assign n54149 = ~n54147 & ~n54148 ;
  assign n54153 = n50649 & ~n54149 ;
  assign n54154 = ~n54152 & n54153 ;
  assign n54162 = ~n26640 & ~n54154 ;
  assign n54163 = ~n54161 & n54162 ;
  assign n54164 = ~n54145 & ~n54163 ;
  assign n54165 = n26792 & ~n54164 ;
  assign n54135 = \P2_P2_rEIP_reg[17]/NET0131  & ~n54099 ;
  assign n54166 = \P2_P2_PhyAddrPointer_reg[17]/NET0131  & n27637 ;
  assign n54167 = ~n28046 & ~n54166 ;
  assign n54168 = ~n54135 & n54167 ;
  assign n54169 = ~n54165 & n54168 ;
  assign n54170 = ~n54144 & n54169 ;
  assign n54173 = n36775 & n52085 ;
  assign n54174 = n36792 & ~n54173 ;
  assign n54176 = ~n43832 & n54174 ;
  assign n54175 = n43832 & ~n54174 ;
  assign n54177 = ~\P2_P2_DataWidth_reg[1]/NET0131  & ~n54175 ;
  assign n54178 = ~n54176 & n54177 ;
  assign n54172 = \P2_P2_DataWidth_reg[1]/NET0131  & ~\P2_P2_rEIP_reg[18]/NET0131  ;
  assign n54179 = n26794 & ~n54172 ;
  assign n54180 = ~n54178 & n54179 ;
  assign n54181 = \P2_P2_rEIP_reg[18]/NET0131  & ~n50640 ;
  assign n54182 = ~\P2_P2_rEIP_reg[18]/NET0131  & ~n54148 ;
  assign n54183 = \P2_P2_rEIP_reg[18]/NET0131  & n54148 ;
  assign n54184 = ~n54182 & ~n54183 ;
  assign n54185 = n50649 & ~n54184 ;
  assign n54186 = ~n26650 & n54185 ;
  assign n54187 = ~\P2_P2_EBX_reg[18]/NET0131  & ~n50642 ;
  assign n54188 = n26643 & ~n54187 ;
  assign n54189 = ~n54186 & n54188 ;
  assign n54190 = \P2_P2_EBX_reg[31]/NET0131  & ~n52129 ;
  assign n54192 = ~\P2_P2_EBX_reg[18]/NET0131  & n54190 ;
  assign n54191 = \P2_P2_EBX_reg[18]/NET0131  & ~n54190 ;
  assign n54193 = ~n50649 & ~n54191 ;
  assign n54194 = ~n54192 & n54193 ;
  assign n54195 = n26633 & ~n54185 ;
  assign n54196 = ~n54194 & n54195 ;
  assign n54197 = ~n54189 & ~n54196 ;
  assign n54198 = ~n26640 & ~n54197 ;
  assign n54199 = ~n54181 & ~n54198 ;
  assign n54200 = n26792 & ~n54199 ;
  assign n54171 = \P2_P2_rEIP_reg[18]/NET0131  & ~n54099 ;
  assign n54201 = \P2_P2_PhyAddrPointer_reg[18]/NET0131  & n27637 ;
  assign n54202 = ~n28046 & ~n54201 ;
  assign n54203 = ~n54171 & n54202 ;
  assign n54204 = ~n54200 & n54203 ;
  assign n54205 = ~n54180 & n54204 ;
  assign n54208 = n36792 & ~n52152 ;
  assign n54210 = n47455 & ~n54208 ;
  assign n54209 = ~n47455 & n54208 ;
  assign n54211 = ~\P2_P2_DataWidth_reg[1]/NET0131  & ~n54209 ;
  assign n54212 = ~n54210 & n54211 ;
  assign n54207 = \P2_P2_DataWidth_reg[1]/NET0131  & ~\P2_P2_rEIP_reg[4]/NET0131  ;
  assign n54213 = n26794 & ~n54207 ;
  assign n54214 = ~n54212 & n54213 ;
  assign n54215 = \P2_P2_rEIP_reg[4]/NET0131  & ~n50640 ;
  assign n54216 = \P2_P2_EBX_reg[31]/NET0131  & ~n52115 ;
  assign n54218 = ~\P2_P2_EBX_reg[4]/NET0131  & n54216 ;
  assign n54217 = \P2_P2_EBX_reg[4]/NET0131  & ~n54216 ;
  assign n54219 = ~n50649 & ~n54217 ;
  assign n54220 = ~n54218 & n54219 ;
  assign n54221 = ~\P2_P2_rEIP_reg[4]/NET0131  & ~n50685 ;
  assign n54222 = ~n52095 & ~n54221 ;
  assign n54223 = n50649 & ~n54222 ;
  assign n54224 = ~n54220 & ~n54223 ;
  assign n54225 = n47684 & n54224 ;
  assign n54226 = ~\P2_P2_EBX_reg[4]/NET0131  & ~n50642 ;
  assign n54227 = n50642 & ~n54222 ;
  assign n54228 = ~n54226 & ~n54227 ;
  assign n54229 = n26786 & n54228 ;
  assign n54230 = ~n54225 & ~n54229 ;
  assign n54231 = ~n54215 & n54230 ;
  assign n54232 = n26792 & ~n54231 ;
  assign n54206 = \P2_P2_rEIP_reg[4]/NET0131  & ~n54099 ;
  assign n54233 = \P2_P2_PhyAddrPointer_reg[4]/NET0131  & n27637 ;
  assign n54234 = ~n28046 & ~n54233 ;
  assign n54235 = ~n54206 & n54234 ;
  assign n54236 = ~n54232 & n54235 ;
  assign n54237 = ~n54214 & n54236 ;
  assign n54240 = ~\P2_P2_PhyAddrPointer_reg[0]/NET0131  & n45079 ;
  assign n54241 = n36792 & ~n54240 ;
  assign n54243 = n48004 & ~n54241 ;
  assign n54242 = ~n48004 & n54241 ;
  assign n54244 = ~\P2_P2_DataWidth_reg[1]/NET0131  & ~n54242 ;
  assign n54245 = ~n54243 & n54244 ;
  assign n54239 = \P2_P2_DataWidth_reg[1]/NET0131  & ~\P2_P2_rEIP_reg[6]/NET0131  ;
  assign n54246 = n26794 & ~n54239 ;
  assign n54247 = ~n54245 & n54246 ;
  assign n54248 = \P2_P2_rEIP_reg[6]/NET0131  & ~n50640 ;
  assign n54249 = \P2_P2_EBX_reg[31]/NET0131  & ~n52117 ;
  assign n54251 = ~\P2_P2_EBX_reg[6]/NET0131  & n54249 ;
  assign n54250 = \P2_P2_EBX_reg[6]/NET0131  & ~n54249 ;
  assign n54252 = ~n50649 & ~n54250 ;
  assign n54253 = ~n54251 & n54252 ;
  assign n54254 = ~\P2_P2_rEIP_reg[6]/NET0131  & ~n52096 ;
  assign n54255 = ~n52097 & ~n54254 ;
  assign n54256 = n50649 & ~n54255 ;
  assign n54257 = ~n54253 & ~n54256 ;
  assign n54258 = n47684 & n54257 ;
  assign n54259 = ~\P2_P2_EBX_reg[6]/NET0131  & ~n50642 ;
  assign n54260 = n50642 & ~n54255 ;
  assign n54261 = ~n54259 & ~n54260 ;
  assign n54262 = n26786 & n54261 ;
  assign n54263 = ~n54258 & ~n54262 ;
  assign n54264 = ~n54248 & n54263 ;
  assign n54265 = n26792 & ~n54264 ;
  assign n54238 = \P2_P2_rEIP_reg[6]/NET0131  & ~n54099 ;
  assign n54266 = \P2_P2_PhyAddrPointer_reg[6]/NET0131  & n27637 ;
  assign n54267 = ~n28046 & ~n54266 ;
  assign n54268 = ~n54238 & n54267 ;
  assign n54269 = ~n54265 & n54268 ;
  assign n54270 = ~n54247 & n54269 ;
  assign n54273 = n36764 & n52485 ;
  assign n54274 = n36792 & ~n54273 ;
  assign n54276 = ~n45082 & n54274 ;
  assign n54275 = n45082 & ~n54274 ;
  assign n54277 = ~\P2_P2_DataWidth_reg[1]/NET0131  & ~n54275 ;
  assign n54278 = ~n54276 & n54277 ;
  assign n54272 = \P2_P2_DataWidth_reg[1]/NET0131  & ~\P2_P2_rEIP_reg[7]/NET0131  ;
  assign n54279 = n26794 & ~n54272 ;
  assign n54280 = ~n54278 & n54279 ;
  assign n54281 = \P2_P2_rEIP_reg[7]/NET0131  & ~n50640 ;
  assign n54282 = ~\P2_P2_EBX_reg[7]/NET0131  & ~n50642 ;
  assign n54283 = ~\P2_P2_rEIP_reg[7]/NET0131  & ~n52097 ;
  assign n54284 = ~n52098 & ~n54283 ;
  assign n54285 = n50642 & ~n54284 ;
  assign n54286 = ~n54282 & ~n54285 ;
  assign n54287 = n26786 & n54286 ;
  assign n54288 = n50649 & ~n54284 ;
  assign n54289 = \P2_P2_EBX_reg[31]/NET0131  & ~n52118 ;
  assign n54291 = \P2_P2_EBX_reg[7]/NET0131  & ~n54289 ;
  assign n54290 = ~\P2_P2_EBX_reg[7]/NET0131  & n54289 ;
  assign n54292 = ~n50649 & ~n54290 ;
  assign n54293 = ~n54291 & n54292 ;
  assign n54294 = ~n54288 & ~n54293 ;
  assign n54295 = n47684 & n54294 ;
  assign n54296 = ~n54287 & ~n54295 ;
  assign n54297 = ~n54281 & n54296 ;
  assign n54298 = n26792 & ~n54297 ;
  assign n54271 = \P2_P2_rEIP_reg[7]/NET0131  & ~n54099 ;
  assign n54299 = \P2_P2_PhyAddrPointer_reg[7]/NET0131  & n27637 ;
  assign n54300 = ~n28046 & ~n54299 ;
  assign n54301 = ~n54271 & n54300 ;
  assign n54302 = ~n54298 & n54301 ;
  assign n54303 = ~n54280 & n54302 ;
  assign n54311 = \P1_P3_InstQueue_reg[0][7]/NET0131  & ~n49750 ;
  assign n54306 = n8797 & n49732 ;
  assign n54305 = ~\P1_P3_InstQueue_reg[0][7]/NET0131  & ~n49732 ;
  assign n54307 = n10046 & ~n54305 ;
  assign n54308 = ~n54306 & n54307 ;
  assign n54304 = \P1_buf2_reg[7]/NET0131  & n49760 ;
  assign n54309 = \P1_buf2_reg[23]/NET0131  & n11698 ;
  assign n54310 = n49742 & n54309 ;
  assign n54312 = ~n54304 & ~n54310 ;
  assign n54313 = ~n54308 & n54312 ;
  assign n54314 = ~n54311 & n54313 ;
  assign n54321 = \P1_P3_InstQueue_reg[10][7]/NET0131  & ~n49776 ;
  assign n54317 = n8797 & n49766 ;
  assign n54316 = ~\P1_P3_InstQueue_reg[10][7]/NET0131  & ~n49766 ;
  assign n54318 = n10046 & ~n54316 ;
  assign n54319 = ~n54317 & n54318 ;
  assign n54315 = \P1_buf2_reg[7]/NET0131  & n49786 ;
  assign n54320 = n49771 & n54309 ;
  assign n54322 = ~n54315 & ~n54320 ;
  assign n54323 = ~n54319 & n54322 ;
  assign n54324 = ~n54321 & n54323 ;
  assign n54331 = \P1_P3_InstQueue_reg[11][7]/NET0131  & ~n49798 ;
  assign n54327 = n8797 & n49792 ;
  assign n54326 = ~\P1_P3_InstQueue_reg[11][7]/NET0131  & ~n49792 ;
  assign n54328 = n10046 & ~n54326 ;
  assign n54329 = ~n54327 & n54328 ;
  assign n54325 = \P1_buf2_reg[7]/NET0131  & n49808 ;
  assign n54330 = n49768 & n54309 ;
  assign n54332 = ~n54325 & ~n54330 ;
  assign n54333 = ~n54329 & n54332 ;
  assign n54334 = ~n54331 & n54333 ;
  assign n54341 = \P1_P3_InstQueue_reg[12][7]/NET0131  & ~n49819 ;
  assign n54337 = n8797 & n49814 ;
  assign n54336 = ~\P1_P3_InstQueue_reg[12][7]/NET0131  & ~n49814 ;
  assign n54338 = n10046 & ~n54336 ;
  assign n54339 = ~n54337 & n54338 ;
  assign n54335 = \P1_buf2_reg[7]/NET0131  & n49829 ;
  assign n54340 = n49766 & n54309 ;
  assign n54342 = ~n54335 & ~n54340 ;
  assign n54343 = ~n54339 & n54342 ;
  assign n54344 = ~n54341 & n54343 ;
  assign n54351 = \P1_P3_InstQueue_reg[13][7]/NET0131  & ~n49838 ;
  assign n54347 = n8797 & n49739 ;
  assign n54346 = ~\P1_P3_InstQueue_reg[13][7]/NET0131  & ~n49739 ;
  assign n54348 = n10046 & ~n54346 ;
  assign n54349 = ~n54347 & n54348 ;
  assign n54345 = \P1_buf2_reg[7]/NET0131  & n49848 ;
  assign n54350 = n49792 & n54309 ;
  assign n54352 = ~n54345 & ~n54350 ;
  assign n54353 = ~n54349 & n54352 ;
  assign n54354 = ~n54351 & n54353 ;
  assign n54361 = \P1_P3_InstQueue_reg[14][7]/NET0131  & ~n49856 ;
  assign n54357 = n8797 & n49742 ;
  assign n54356 = ~\P1_P3_InstQueue_reg[14][7]/NET0131  & ~n49742 ;
  assign n54358 = n10046 & ~n54356 ;
  assign n54359 = ~n54357 & n54358 ;
  assign n54355 = \P1_buf2_reg[7]/NET0131  & n49866 ;
  assign n54360 = n49814 & n54309 ;
  assign n54362 = ~n54355 & ~n54360 ;
  assign n54363 = ~n54359 & n54362 ;
  assign n54364 = ~n54361 & n54363 ;
  assign n54371 = \P1_P3_InstQueue_reg[15][7]/NET0131  & ~n49875 ;
  assign n54367 = n8797 & n49735 ;
  assign n54366 = ~\P1_P3_InstQueue_reg[15][7]/NET0131  & ~n49735 ;
  assign n54368 = n10046 & ~n54366 ;
  assign n54369 = ~n54367 & n54368 ;
  assign n54365 = \P1_buf2_reg[7]/NET0131  & n49885 ;
  assign n54370 = n49739 & n54309 ;
  assign n54372 = ~n54365 & ~n54370 ;
  assign n54373 = ~n54369 & n54372 ;
  assign n54374 = ~n54371 & n54373 ;
  assign n54381 = \P1_P3_InstQueue_reg[1][7]/NET0131  & ~n49895 ;
  assign n54377 = n8797 & n49890 ;
  assign n54376 = ~\P1_P3_InstQueue_reg[1][7]/NET0131  & ~n49890 ;
  assign n54378 = n10046 & ~n54376 ;
  assign n54379 = ~n54377 & n54378 ;
  assign n54375 = \P1_buf2_reg[7]/NET0131  & n49905 ;
  assign n54380 = n49735 & n54309 ;
  assign n54382 = ~n54375 & ~n54380 ;
  assign n54383 = ~n54379 & n54382 ;
  assign n54384 = ~n54381 & n54383 ;
  assign n54391 = \P1_P3_InstQueue_reg[2][7]/NET0131  & ~n49915 ;
  assign n54387 = n8797 & n49910 ;
  assign n54386 = ~\P1_P3_InstQueue_reg[2][7]/NET0131  & ~n49910 ;
  assign n54388 = n10046 & ~n54386 ;
  assign n54389 = ~n54387 & n54388 ;
  assign n54385 = \P1_buf2_reg[7]/NET0131  & n49925 ;
  assign n54390 = n49732 & n54309 ;
  assign n54392 = ~n54385 & ~n54390 ;
  assign n54393 = ~n54389 & n54392 ;
  assign n54394 = ~n54391 & n54393 ;
  assign n54401 = \P1_P3_InstQueue_reg[3][7]/NET0131  & ~n49935 ;
  assign n54397 = n8797 & n49930 ;
  assign n54396 = ~\P1_P3_InstQueue_reg[3][7]/NET0131  & ~n49930 ;
  assign n54398 = n10046 & ~n54396 ;
  assign n54399 = ~n54397 & n54398 ;
  assign n54395 = \P1_buf2_reg[7]/NET0131  & n49945 ;
  assign n54400 = n49890 & n54309 ;
  assign n54402 = ~n54395 & ~n54400 ;
  assign n54403 = ~n54399 & n54402 ;
  assign n54404 = ~n54401 & n54403 ;
  assign n54411 = \P1_P3_InstQueue_reg[4][7]/NET0131  & ~n49955 ;
  assign n54407 = n8797 & n49950 ;
  assign n54406 = ~\P1_P3_InstQueue_reg[4][7]/NET0131  & ~n49950 ;
  assign n54408 = n10046 & ~n54406 ;
  assign n54409 = ~n54407 & n54408 ;
  assign n54405 = \P1_buf2_reg[7]/NET0131  & n49965 ;
  assign n54410 = n49910 & n54309 ;
  assign n54412 = ~n54405 & ~n54410 ;
  assign n54413 = ~n54409 & n54412 ;
  assign n54414 = ~n54411 & n54413 ;
  assign n54421 = \P1_P3_InstQueue_reg[5][7]/NET0131  & ~n49975 ;
  assign n54417 = n8797 & n49970 ;
  assign n54416 = ~\P1_P3_InstQueue_reg[5][7]/NET0131  & ~n49970 ;
  assign n54418 = n10046 & ~n54416 ;
  assign n54419 = ~n54417 & n54418 ;
  assign n54415 = \P1_buf2_reg[7]/NET0131  & n49985 ;
  assign n54420 = n49930 & n54309 ;
  assign n54422 = ~n54415 & ~n54420 ;
  assign n54423 = ~n54419 & n54422 ;
  assign n54424 = ~n54421 & n54423 ;
  assign n54427 = n26896 & n50021 ;
  assign n54426 = ~\P2_P3_InstQueue_reg[0][7]/NET0131  & ~n50021 ;
  assign n54428 = n27788 & ~n54426 ;
  assign n54429 = ~n54427 & n54428 ;
  assign n54432 = \P2_P3_InstQueue_reg[0][7]/NET0131  & ~n50030 ;
  assign n54425 = \P2_buf2_reg[7]/NET0131  & n50040 ;
  assign n54430 = \P2_buf2_reg[23]/NET0131  & n27325 ;
  assign n54431 = n50015 & n54430 ;
  assign n54433 = ~n54425 & ~n54431 ;
  assign n54434 = ~n54432 & n54433 ;
  assign n54435 = ~n54429 & n54434 ;
  assign n54442 = \P1_P3_InstQueue_reg[6][7]/NET0131  & ~n49995 ;
  assign n54438 = n8797 & n49990 ;
  assign n54437 = ~\P1_P3_InstQueue_reg[6][7]/NET0131  & ~n49990 ;
  assign n54439 = n10046 & ~n54437 ;
  assign n54440 = ~n54438 & n54439 ;
  assign n54436 = \P1_buf2_reg[7]/NET0131  & n50005 ;
  assign n54441 = n49950 & n54309 ;
  assign n54443 = ~n54436 & ~n54441 ;
  assign n54444 = ~n54440 & n54443 ;
  assign n54445 = ~n54442 & n54444 ;
  assign n54448 = n26896 & n50051 ;
  assign n54447 = ~\P2_P3_InstQueue_reg[10][7]/NET0131  & ~n50051 ;
  assign n54449 = n27788 & ~n54447 ;
  assign n54450 = ~n54448 & n54449 ;
  assign n54452 = \P2_P3_InstQueue_reg[10][7]/NET0131  & ~n50056 ;
  assign n54446 = \P2_buf2_reg[7]/NET0131  & n50066 ;
  assign n54451 = n50045 & n54430 ;
  assign n54453 = ~n54446 & ~n54451 ;
  assign n54454 = ~n54452 & n54453 ;
  assign n54455 = ~n54450 & n54454 ;
  assign n54462 = \P1_P3_InstQueue_reg[7][7]/NET0131  & ~n50075 ;
  assign n54458 = n8797 & n49770 ;
  assign n54457 = ~\P1_P3_InstQueue_reg[7][7]/NET0131  & ~n49770 ;
  assign n54459 = n10046 & ~n54457 ;
  assign n54460 = ~n54458 & n54459 ;
  assign n54456 = \P1_buf2_reg[7]/NET0131  & n50085 ;
  assign n54461 = n49970 & n54309 ;
  assign n54463 = ~n54456 & ~n54461 ;
  assign n54464 = ~n54460 & n54463 ;
  assign n54465 = ~n54462 & n54464 ;
  assign n54468 = n26896 & n50094 ;
  assign n54467 = ~\P2_P3_InstQueue_reg[11][7]/NET0131  & ~n50094 ;
  assign n54469 = n27788 & ~n54467 ;
  assign n54470 = ~n54468 & n54469 ;
  assign n54472 = \P2_P3_InstQueue_reg[11][7]/NET0131  & ~n50097 ;
  assign n54466 = \P2_buf2_reg[7]/NET0131  & n50107 ;
  assign n54471 = n50053 & n54430 ;
  assign n54473 = ~n54466 & ~n54471 ;
  assign n54474 = ~n54472 & n54473 ;
  assign n54475 = ~n54470 & n54474 ;
  assign n54478 = n26896 & n50115 ;
  assign n54477 = ~\P2_P3_InstQueue_reg[12][7]/NET0131  & ~n50115 ;
  assign n54479 = n27788 & ~n54477 ;
  assign n54480 = ~n54478 & n54479 ;
  assign n54482 = \P2_P3_InstQueue_reg[12][7]/NET0131  & ~n50118 ;
  assign n54476 = \P2_buf2_reg[7]/NET0131  & n50128 ;
  assign n54481 = n50051 & n54430 ;
  assign n54483 = ~n54476 & ~n54481 ;
  assign n54484 = ~n54482 & n54483 ;
  assign n54485 = ~n54480 & n54484 ;
  assign n54492 = \P1_P3_InstQueue_reg[8][7]/NET0131  & ~n50136 ;
  assign n54488 = n8797 & n49771 ;
  assign n54487 = ~\P1_P3_InstQueue_reg[8][7]/NET0131  & ~n49771 ;
  assign n54489 = n10046 & ~n54487 ;
  assign n54490 = ~n54488 & n54489 ;
  assign n54486 = \P1_buf2_reg[7]/NET0131  & n50146 ;
  assign n54491 = n49990 & n54309 ;
  assign n54493 = ~n54486 & ~n54491 ;
  assign n54494 = ~n54490 & n54493 ;
  assign n54495 = ~n54492 & n54494 ;
  assign n54498 = n26896 & n50012 ;
  assign n54497 = ~\P2_P3_InstQueue_reg[13][7]/NET0131  & ~n50012 ;
  assign n54499 = n27788 & ~n54497 ;
  assign n54500 = ~n54498 & n54499 ;
  assign n54502 = \P2_P3_InstQueue_reg[13][7]/NET0131  & ~n50155 ;
  assign n54496 = \P2_buf2_reg[7]/NET0131  & n50165 ;
  assign n54501 = n50094 & n54430 ;
  assign n54503 = ~n54496 & ~n54501 ;
  assign n54504 = ~n54502 & n54503 ;
  assign n54505 = ~n54500 & n54504 ;
  assign n54508 = n26896 & n50015 ;
  assign n54507 = ~\P2_P3_InstQueue_reg[14][7]/NET0131  & ~n50015 ;
  assign n54509 = n27788 & ~n54507 ;
  assign n54510 = ~n54508 & n54509 ;
  assign n54512 = \P2_P3_InstQueue_reg[14][7]/NET0131  & ~n50173 ;
  assign n54506 = \P2_buf2_reg[7]/NET0131  & n50183 ;
  assign n54511 = n50115 & n54430 ;
  assign n54513 = ~n54506 & ~n54511 ;
  assign n54514 = ~n54512 & n54513 ;
  assign n54515 = ~n54510 & n54514 ;
  assign n54522 = \P1_P3_InstQueue_reg[9][7]/NET0131  & ~n50191 ;
  assign n54518 = n8797 & n49768 ;
  assign n54517 = ~\P1_P3_InstQueue_reg[9][7]/NET0131  & ~n49768 ;
  assign n54519 = n10046 & ~n54517 ;
  assign n54520 = ~n54518 & n54519 ;
  assign n54516 = \P1_buf2_reg[7]/NET0131  & n50201 ;
  assign n54521 = n49770 & n54309 ;
  assign n54523 = ~n54516 & ~n54521 ;
  assign n54524 = ~n54520 & n54523 ;
  assign n54525 = ~n54522 & n54524 ;
  assign n54528 = n26896 & n50024 ;
  assign n54527 = ~\P2_P3_InstQueue_reg[15][7]/NET0131  & ~n50024 ;
  assign n54529 = n27788 & ~n54527 ;
  assign n54530 = ~n54528 & n54529 ;
  assign n54532 = \P2_P3_InstQueue_reg[15][7]/NET0131  & ~n50210 ;
  assign n54526 = \P2_buf2_reg[7]/NET0131  & n50220 ;
  assign n54531 = n50012 & n54430 ;
  assign n54533 = ~n54526 & ~n54531 ;
  assign n54534 = ~n54532 & n54533 ;
  assign n54535 = ~n54530 & n54534 ;
  assign n54538 = \P1_P3_MemoryFetch_reg/NET0131  & ~n16498 ;
  assign n54539 = n22899 & ~n54538 ;
  assign n54540 = n9241 & ~n54539 ;
  assign n54536 = ~n10030 & n18341 ;
  assign n54537 = \P1_P3_MemoryFetch_reg/NET0131  & ~n54536 ;
  assign n54541 = n43255 & ~n54537 ;
  assign n54542 = ~n54540 & n54541 ;
  assign n54545 = n26896 & n50227 ;
  assign n54544 = ~\P2_P3_InstQueue_reg[1][7]/NET0131  & ~n50227 ;
  assign n54546 = n27788 & ~n54544 ;
  assign n54547 = ~n54545 & n54546 ;
  assign n54549 = \P2_P3_InstQueue_reg[1][7]/NET0131  & ~n50230 ;
  assign n54543 = \P2_buf2_reg[7]/NET0131  & n50240 ;
  assign n54548 = n50024 & n54430 ;
  assign n54550 = ~n54543 & ~n54548 ;
  assign n54551 = ~n54549 & n54550 ;
  assign n54552 = ~n54547 & n54551 ;
  assign n54555 = n26896 & n50247 ;
  assign n54554 = ~\P2_P3_InstQueue_reg[2][7]/NET0131  & ~n50247 ;
  assign n54556 = n27788 & ~n54554 ;
  assign n54557 = ~n54555 & n54556 ;
  assign n54559 = \P2_P3_InstQueue_reg[2][7]/NET0131  & ~n50250 ;
  assign n54553 = \P2_buf2_reg[7]/NET0131  & n50260 ;
  assign n54558 = n50021 & n54430 ;
  assign n54560 = ~n54553 & ~n54558 ;
  assign n54561 = ~n54559 & n54560 ;
  assign n54562 = ~n54557 & n54561 ;
  assign n54565 = n26896 & n50267 ;
  assign n54564 = ~\P2_P3_InstQueue_reg[3][7]/NET0131  & ~n50267 ;
  assign n54566 = n27788 & ~n54564 ;
  assign n54567 = ~n54565 & n54566 ;
  assign n54569 = \P2_P3_InstQueue_reg[3][7]/NET0131  & ~n50270 ;
  assign n54563 = \P2_buf2_reg[7]/NET0131  & n50280 ;
  assign n54568 = n50227 & n54430 ;
  assign n54570 = ~n54563 & ~n54568 ;
  assign n54571 = ~n54569 & n54570 ;
  assign n54572 = ~n54567 & n54571 ;
  assign n54575 = n26896 & n50287 ;
  assign n54574 = ~\P2_P3_InstQueue_reg[4][7]/NET0131  & ~n50287 ;
  assign n54576 = n27788 & ~n54574 ;
  assign n54577 = ~n54575 & n54576 ;
  assign n54579 = \P2_P3_InstQueue_reg[4][7]/NET0131  & ~n50290 ;
  assign n54573 = \P2_buf2_reg[7]/NET0131  & n50300 ;
  assign n54578 = n50247 & n54430 ;
  assign n54580 = ~n54573 & ~n54578 ;
  assign n54581 = ~n54579 & n54580 ;
  assign n54582 = ~n54577 & n54581 ;
  assign n54585 = n26896 & n50307 ;
  assign n54584 = ~\P2_P3_InstQueue_reg[5][7]/NET0131  & ~n50307 ;
  assign n54586 = n27788 & ~n54584 ;
  assign n54587 = ~n54585 & n54586 ;
  assign n54589 = \P2_P3_InstQueue_reg[5][7]/NET0131  & ~n50310 ;
  assign n54583 = \P2_buf2_reg[7]/NET0131  & n50320 ;
  assign n54588 = n50267 & n54430 ;
  assign n54590 = ~n54583 & ~n54588 ;
  assign n54591 = ~n54589 & n54590 ;
  assign n54592 = ~n54587 & n54591 ;
  assign n54595 = n26896 & n50327 ;
  assign n54594 = ~\P2_P3_InstQueue_reg[6][7]/NET0131  & ~n50327 ;
  assign n54596 = n27788 & ~n54594 ;
  assign n54597 = ~n54595 & n54596 ;
  assign n54599 = \P2_P3_InstQueue_reg[6][7]/NET0131  & ~n50330 ;
  assign n54593 = \P2_buf2_reg[7]/NET0131  & n50340 ;
  assign n54598 = n50287 & n54430 ;
  assign n54600 = ~n54593 & ~n54598 ;
  assign n54601 = ~n54599 & n54600 ;
  assign n54602 = ~n54597 & n54601 ;
  assign n54605 = n26896 & n50046 ;
  assign n54604 = ~\P2_P3_InstQueue_reg[7][7]/NET0131  & ~n50046 ;
  assign n54606 = n27788 & ~n54604 ;
  assign n54607 = ~n54605 & n54606 ;
  assign n54609 = \P2_P3_InstQueue_reg[7][7]/NET0131  & ~n50349 ;
  assign n54603 = \P2_buf2_reg[7]/NET0131  & n50359 ;
  assign n54608 = n50307 & n54430 ;
  assign n54610 = ~n54603 & ~n54608 ;
  assign n54611 = ~n54609 & n54610 ;
  assign n54612 = ~n54607 & n54611 ;
  assign n54615 = n26896 & n50045 ;
  assign n54614 = ~\P2_P3_InstQueue_reg[8][7]/NET0131  & ~n50045 ;
  assign n54616 = n27788 & ~n54614 ;
  assign n54617 = ~n54615 & n54616 ;
  assign n54619 = \P2_P3_InstQueue_reg[8][7]/NET0131  & ~n50367 ;
  assign n54613 = \P2_buf2_reg[7]/NET0131  & n50377 ;
  assign n54618 = n50327 & n54430 ;
  assign n54620 = ~n54613 & ~n54618 ;
  assign n54621 = ~n54619 & n54620 ;
  assign n54622 = ~n54617 & n54621 ;
  assign n54625 = n26896 & n50053 ;
  assign n54624 = ~\P2_P3_InstQueue_reg[9][7]/NET0131  & ~n50053 ;
  assign n54626 = n27788 & ~n54624 ;
  assign n54627 = ~n54625 & n54626 ;
  assign n54629 = \P2_P3_InstQueue_reg[9][7]/NET0131  & ~n50385 ;
  assign n54623 = \P2_buf2_reg[7]/NET0131  & n50395 ;
  assign n54628 = n50046 & n54430 ;
  assign n54630 = ~n54623 & ~n54628 ;
  assign n54631 = ~n54629 & n54630 ;
  assign n54632 = ~n54627 & n54631 ;
  assign n54634 = n27124 & ~n27177 ;
  assign n54635 = \P2_P3_MemoryFetch_reg/NET0131  & ~n54634 ;
  assign n54636 = n47748 & ~n54635 ;
  assign n54637 = n27308 & ~n54636 ;
  assign n54633 = \P2_P3_MemoryFetch_reg/NET0131  & ~n47745 ;
  assign n54638 = n43269 & ~n54633 ;
  assign n54639 = ~n54637 & n54638 ;
  assign n54641 = \P1_P3_ReadRequest_reg/NET0131  & ~n21775 ;
  assign n54642 = ~n9147 & ~n54641 ;
  assign n54643 = n9241 & ~n54642 ;
  assign n54640 = \P1_P3_ReadRequest_reg/NET0131  & ~n54536 ;
  assign n54644 = n43255 & ~n54640 ;
  assign n54645 = ~n54643 & n54644 ;
  assign n54647 = ~n27177 & ~n27180 ;
  assign n54648 = \P2_P3_ReadRequest_reg/NET0131  & ~n54647 ;
  assign n54649 = ~n27256 & ~n54648 ;
  assign n54650 = n27308 & ~n54649 ;
  assign n54646 = \P2_P3_ReadRequest_reg/NET0131  & ~n47745 ;
  assign n54651 = n43269 & ~n54646 ;
  assign n54652 = ~n54650 & n54651 ;
  assign n54656 = \P2_P3_PhyAddrPointer_reg[14]/NET0131  & n39837 ;
  assign n54657 = n52576 & n54656 ;
  assign n54658 = ~n36863 & ~n54657 ;
  assign n54660 = ~n39847 & n54658 ;
  assign n54659 = n39847 & ~n54658 ;
  assign n54661 = ~\P2_P3_DataWidth_reg[1]/NET0131  & ~n54659 ;
  assign n54662 = ~n54660 & n54661 ;
  assign n54655 = \P2_P3_DataWidth_reg[1]/NET0131  & ~\P2_P3_rEIP_reg[15]/NET0131  ;
  assign n54663 = n27315 & ~n54655 ;
  assign n54664 = ~n54662 & n54663 ;
  assign n54669 = \P2_P3_EBX_reg[31]/NET0131  & ~n52535 ;
  assign n54670 = ~\P2_P3_EBX_reg[15]/NET0131  & ~n54669 ;
  assign n54671 = \P2_P3_EBX_reg[15]/NET0131  & n54669 ;
  assign n54672 = ~n54670 & ~n54671 ;
  assign n54673 = ~n27302 & ~n54672 ;
  assign n54666 = ~\P2_P3_rEIP_reg[15]/NET0131  & ~n52559 ;
  assign n54667 = ~n52560 & ~n54666 ;
  assign n54668 = n27302 & ~n54667 ;
  assign n54674 = n46587 & ~n54668 ;
  assign n54675 = ~n54673 & n54674 ;
  assign n54665 = \P2_P3_rEIP_reg[15]/NET0131  & ~n27277 ;
  assign n54677 = n50735 & ~n54667 ;
  assign n54676 = ~\P2_P3_EBX_reg[15]/NET0131  & ~n50735 ;
  assign n54678 = n47747 & ~n54676 ;
  assign n54679 = ~n54677 & n54678 ;
  assign n54680 = ~n54665 & ~n54679 ;
  assign n54681 = ~n54675 & n54680 ;
  assign n54682 = n27308 & ~n54681 ;
  assign n54653 = n27319 & n27789 ;
  assign n54654 = \P2_P3_rEIP_reg[15]/NET0131  & ~n54653 ;
  assign n54683 = \P2_P3_PhyAddrPointer_reg[15]/NET0131  & n27651 ;
  assign n54684 = ~n32864 & ~n54683 ;
  assign n54685 = ~n54654 & n54684 ;
  assign n54686 = ~n54682 & n54685 ;
  assign n54687 = ~n54664 & n54686 ;
  assign n54690 = n44090 & n52576 ;
  assign n54691 = ~n36863 & ~n54690 ;
  assign n54693 = n44096 & ~n54691 ;
  assign n54692 = ~n44096 & n54691 ;
  assign n54694 = ~\P2_P3_DataWidth_reg[1]/NET0131  & ~n54692 ;
  assign n54695 = ~n54693 & n54694 ;
  assign n54689 = \P2_P3_DataWidth_reg[1]/NET0131  & ~\P2_P3_rEIP_reg[17]/NET0131  ;
  assign n54696 = n27315 & ~n54689 ;
  assign n54697 = ~n54695 & n54696 ;
  assign n54698 = \P2_P3_rEIP_reg[17]/NET0131  & ~n27277 ;
  assign n54700 = ~\P2_P3_rEIP_reg[17]/NET0131  & ~n52561 ;
  assign n54701 = ~n52562 & ~n54700 ;
  assign n54702 = n50735 & ~n54701 ;
  assign n54699 = ~\P2_P3_EBX_reg[17]/NET0131  & ~n50735 ;
  assign n54703 = n27121 & ~n54699 ;
  assign n54704 = ~n54702 & n54703 ;
  assign n54706 = \P2_P3_EBX_reg[31]/NET0131  & ~n52537 ;
  assign n54707 = ~\P2_P3_EBX_reg[17]/NET0131  & ~n54706 ;
  assign n54708 = \P2_P3_EBX_reg[17]/NET0131  & n54706 ;
  assign n54709 = ~n54707 & ~n54708 ;
  assign n54710 = ~n27302 & ~n54709 ;
  assign n54705 = n27302 & ~n54701 ;
  assign n54711 = n27122 & ~n54705 ;
  assign n54712 = ~n54710 & n54711 ;
  assign n54713 = ~n54704 & ~n54712 ;
  assign n54714 = ~n27177 & ~n54713 ;
  assign n54715 = ~n54698 & ~n54714 ;
  assign n54716 = n27308 & ~n54715 ;
  assign n54688 = \P2_P3_rEIP_reg[17]/NET0131  & ~n54653 ;
  assign n54717 = \P2_P3_PhyAddrPointer_reg[17]/NET0131  & n27651 ;
  assign n54718 = ~n32864 & ~n54717 ;
  assign n54719 = ~n54688 & n54718 ;
  assign n54720 = ~n54716 & n54719 ;
  assign n54721 = ~n54697 & n54720 ;
  assign n54743 = ~n36863 & ~n52576 ;
  assign n54744 = ~n36863 & ~n42106 ;
  assign n54745 = ~n54743 & ~n54744 ;
  assign n54747 = ~n44115 & ~n54745 ;
  assign n54746 = n44115 & n54745 ;
  assign n54748 = ~\P2_P3_DataWidth_reg[1]/NET0131  & ~n54746 ;
  assign n54749 = ~n54747 & n54748 ;
  assign n54742 = \P2_P3_DataWidth_reg[1]/NET0131  & ~\P2_P3_rEIP_reg[18]/NET0131  ;
  assign n54750 = n27315 & ~n54742 ;
  assign n54751 = ~n54749 & n54750 ;
  assign n54723 = \P2_P3_rEIP_reg[18]/NET0131  & ~n27277 ;
  assign n54725 = ~\P2_P3_rEIP_reg[18]/NET0131  & ~n52562 ;
  assign n54726 = ~n52563 & ~n54725 ;
  assign n54727 = n50735 & ~n54726 ;
  assign n54724 = ~\P2_P3_EBX_reg[18]/NET0131  & ~n50735 ;
  assign n54728 = n27121 & ~n54724 ;
  assign n54729 = ~n54727 & n54728 ;
  assign n54731 = \P2_P3_EBX_reg[31]/NET0131  & ~n52538 ;
  assign n54733 = ~\P2_P3_EBX_reg[18]/NET0131  & n54731 ;
  assign n54732 = \P2_P3_EBX_reg[18]/NET0131  & ~n54731 ;
  assign n54734 = ~n27302 & ~n54732 ;
  assign n54735 = ~n54733 & n54734 ;
  assign n54730 = n27302 & ~n54726 ;
  assign n54736 = n27122 & ~n54730 ;
  assign n54737 = ~n54735 & n54736 ;
  assign n54738 = ~n54729 & ~n54737 ;
  assign n54739 = ~n27177 & ~n54738 ;
  assign n54740 = ~n54723 & ~n54739 ;
  assign n54741 = n27308 & ~n54740 ;
  assign n54722 = \P2_P3_rEIP_reg[18]/NET0131  & ~n54653 ;
  assign n54752 = \P2_P3_PhyAddrPointer_reg[18]/NET0131  & n27651 ;
  assign n54753 = ~n32864 & ~n54752 ;
  assign n54754 = ~n54722 & n54753 ;
  assign n54755 = ~n54741 & n54754 ;
  assign n54756 = ~n54751 & n54755 ;
  assign n54759 = ~n36835 & ~n36863 ;
  assign n54760 = ~n50709 & ~n54759 ;
  assign n54762 = ~n47481 & ~n54760 ;
  assign n54761 = n47481 & n54760 ;
  assign n54763 = ~\P2_P3_DataWidth_reg[1]/NET0131  & ~n54761 ;
  assign n54764 = ~n54762 & n54763 ;
  assign n54758 = \P2_P3_DataWidth_reg[1]/NET0131  & ~\P2_P3_rEIP_reg[4]/NET0131  ;
  assign n54765 = n27315 & ~n54758 ;
  assign n54766 = ~n54764 & n54765 ;
  assign n54767 = \P2_P3_rEIP_reg[4]/NET0131  & ~n27277 ;
  assign n54768 = ~\P2_P3_EBX_reg[4]/NET0131  & ~n50735 ;
  assign n54769 = ~\P2_P3_rEIP_reg[4]/NET0131  & ~n50728 ;
  assign n54770 = ~n52549 & ~n54769 ;
  assign n54771 = n50735 & ~n54770 ;
  assign n54772 = ~n54768 & ~n54771 ;
  assign n54773 = n47747 & n54772 ;
  assign n54774 = n27302 & ~n54770 ;
  assign n54775 = \P2_P3_EBX_reg[31]/NET0131  & ~n52524 ;
  assign n54777 = ~\P2_P3_EBX_reg[4]/NET0131  & n54775 ;
  assign n54776 = \P2_P3_EBX_reg[4]/NET0131  & ~n54775 ;
  assign n54778 = ~n27302 & ~n54776 ;
  assign n54779 = ~n54777 & n54778 ;
  assign n54780 = ~n54774 & ~n54779 ;
  assign n54781 = n46587 & n54780 ;
  assign n54782 = ~n54773 & ~n54781 ;
  assign n54783 = ~n54767 & n54782 ;
  assign n54784 = n27308 & ~n54783 ;
  assign n54757 = \P2_P3_rEIP_reg[4]/NET0131  & ~n54653 ;
  assign n54785 = \P2_P3_PhyAddrPointer_reg[4]/NET0131  & n27651 ;
  assign n54786 = ~n32864 & ~n54785 ;
  assign n54787 = ~n54757 & n54786 ;
  assign n54788 = ~n54784 & n54787 ;
  assign n54789 = ~n54766 & n54788 ;
  assign n54792 = n36837 & n50708 ;
  assign n54793 = ~n36863 & ~n54792 ;
  assign n54795 = ~n48123 & n54793 ;
  assign n54794 = n48123 & ~n54793 ;
  assign n54796 = ~\P2_P3_DataWidth_reg[1]/NET0131  & ~n54794 ;
  assign n54797 = ~n54795 & n54796 ;
  assign n54791 = \P2_P3_DataWidth_reg[1]/NET0131  & ~\P2_P3_rEIP_reg[6]/NET0131  ;
  assign n54798 = n27315 & ~n54791 ;
  assign n54799 = ~n54797 & n54798 ;
  assign n54800 = \P2_P3_rEIP_reg[6]/NET0131  & ~n27277 ;
  assign n54801 = ~\P2_P3_rEIP_reg[6]/NET0131  & ~n52550 ;
  assign n54802 = ~n52551 & ~n54801 ;
  assign n54803 = n27302 & ~n54802 ;
  assign n54804 = ~n27148 & n54803 ;
  assign n54805 = ~\P2_P3_EBX_reg[6]/NET0131  & ~n50735 ;
  assign n54806 = ~n54804 & ~n54805 ;
  assign n54807 = n47747 & n54806 ;
  assign n54808 = \P2_P3_EBX_reg[31]/NET0131  & ~n52526 ;
  assign n54810 = ~\P2_P3_EBX_reg[6]/NET0131  & n54808 ;
  assign n54809 = \P2_P3_EBX_reg[6]/NET0131  & ~n54808 ;
  assign n54811 = ~n27302 & ~n54809 ;
  assign n54812 = ~n54810 & n54811 ;
  assign n54813 = ~n54803 & ~n54812 ;
  assign n54814 = n46587 & n54813 ;
  assign n54815 = ~n54807 & ~n54814 ;
  assign n54816 = ~n54800 & n54815 ;
  assign n54817 = n27308 & ~n54816 ;
  assign n54790 = \P2_P3_rEIP_reg[6]/NET0131  & ~n54653 ;
  assign n54818 = \P2_P3_PhyAddrPointer_reg[6]/NET0131  & n27651 ;
  assign n54819 = ~n32864 & ~n54818 ;
  assign n54820 = ~n54790 & n54819 ;
  assign n54821 = ~n54817 & n54820 ;
  assign n54822 = ~n54799 & n54821 ;
  assign n54825 = ~\P2_P3_PhyAddrPointer_reg[0]/NET0131  & n44156 ;
  assign n54826 = ~n36863 & ~n54825 ;
  assign n54828 = ~n45206 & n54826 ;
  assign n54827 = n45206 & ~n54826 ;
  assign n54829 = ~\P2_P3_DataWidth_reg[1]/NET0131  & ~n54827 ;
  assign n54830 = ~n54828 & n54829 ;
  assign n54824 = \P2_P3_DataWidth_reg[1]/NET0131  & ~\P2_P3_rEIP_reg[7]/NET0131  ;
  assign n54831 = n27315 & ~n54824 ;
  assign n54832 = ~n54830 & n54831 ;
  assign n54833 = \P2_P3_rEIP_reg[7]/NET0131  & ~n27277 ;
  assign n54834 = \P2_P3_EBX_reg[31]/NET0131  & ~n52527 ;
  assign n54835 = ~\P2_P3_EBX_reg[7]/NET0131  & ~n54834 ;
  assign n54836 = \P2_P3_EBX_reg[7]/NET0131  & n54834 ;
  assign n54837 = ~n54835 & ~n54836 ;
  assign n54838 = ~n27302 & ~n54837 ;
  assign n54839 = ~\P2_P3_rEIP_reg[7]/NET0131  & ~n52551 ;
  assign n54840 = ~n52552 & ~n54839 ;
  assign n54841 = n27302 & ~n54840 ;
  assign n54842 = ~n54838 & ~n54841 ;
  assign n54843 = n46587 & n54842 ;
  assign n54844 = n50735 & ~n54840 ;
  assign n54845 = ~\P2_P3_EBX_reg[7]/NET0131  & ~n50735 ;
  assign n54846 = ~n54844 & ~n54845 ;
  assign n54847 = n47747 & n54846 ;
  assign n54848 = ~n54843 & ~n54847 ;
  assign n54849 = ~n54833 & n54848 ;
  assign n54850 = n27308 & ~n54849 ;
  assign n54823 = \P2_P3_rEIP_reg[7]/NET0131  & ~n54653 ;
  assign n54851 = \P2_P3_PhyAddrPointer_reg[7]/NET0131  & n27651 ;
  assign n54852 = ~n32864 & ~n54851 ;
  assign n54853 = ~n54823 & n54852 ;
  assign n54854 = ~n54850 & n54853 ;
  assign n54855 = ~n54832 & n54854 ;
  assign n54858 = n36672 & ~n50823 ;
  assign n54860 = n44892 & ~n54858 ;
  assign n54859 = ~n44892 & n54858 ;
  assign n54861 = ~\P2_P1_DataWidth_reg[1]/NET0131  & ~n54859 ;
  assign n54862 = ~n54860 & n54861 ;
  assign n54857 = \P2_P1_DataWidth_reg[1]/NET0131  & ~\P2_P1_rEIP_reg[10]/NET0131  ;
  assign n54863 = n11609 & ~n54857 ;
  assign n54864 = ~n54862 & n54863 ;
  assign n54865 = \P2_P1_rEIP_reg[10]/NET0131  & ~n50414 ;
  assign n54867 = \P2_P1_rEIP_reg[10]/NET0131  & n50771 ;
  assign n54868 = ~\P2_P1_rEIP_reg[10]/NET0131  & ~n50771 ;
  assign n54869 = ~n54867 & ~n54868 ;
  assign n54870 = n50422 & ~n54869 ;
  assign n54871 = ~n25958 & n54870 ;
  assign n54866 = ~\P2_P1_EBX_reg[10]/NET0131  & ~n26103 ;
  assign n54872 = n24898 & ~n54866 ;
  assign n54873 = ~n54871 & n54872 ;
  assign n54874 = \P2_P1_EBX_reg[31]/NET0131  & ~n50795 ;
  assign n54876 = ~\P2_P1_EBX_reg[10]/NET0131  & n54874 ;
  assign n54875 = \P2_P1_EBX_reg[10]/NET0131  & ~n54874 ;
  assign n54877 = ~n50422 & ~n54875 ;
  assign n54878 = ~n54876 & n54877 ;
  assign n54879 = n21062 & ~n54870 ;
  assign n54880 = ~n54878 & n54879 ;
  assign n54881 = ~n54873 & ~n54880 ;
  assign n54882 = ~n21081 & ~n54881 ;
  assign n54883 = ~n54865 & ~n54882 ;
  assign n54884 = n11623 & ~n54883 ;
  assign n54856 = \P2_P1_rEIP_reg[10]/NET0131  & ~n53464 ;
  assign n54885 = \P2_P1_PhyAddrPointer_reg[10]/NET0131  & n11625 ;
  assign n54886 = ~n11616 & ~n54885 ;
  assign n54887 = ~n54856 & n54886 ;
  assign n54888 = ~n54884 & n54887 ;
  assign n54889 = ~n54864 & n54888 ;
  assign n54892 = ~n36628 & ~n48455 ;
  assign n54893 = ~n36628 & ~n44866 ;
  assign n54894 = ~n54892 & ~n54893 ;
  assign n54896 = n44868 & n54894 ;
  assign n54895 = ~n44868 & ~n54894 ;
  assign n54897 = ~\P1_P2_DataWidth_reg[1]/NET0131  & ~n54895 ;
  assign n54898 = ~n54896 & n54897 ;
  assign n54891 = \P1_P2_DataWidth_reg[1]/NET0131  & ~\P1_P2_rEIP_reg[10]/NET0131  ;
  assign n54899 = n25928 & ~n54891 ;
  assign n54900 = ~n54898 & n54899 ;
  assign n54901 = \P1_P2_rEIP_reg[10]/NET0131  & ~n48371 ;
  assign n54902 = \P1_P2_rEIP_reg[10]/NET0131  & n51239 ;
  assign n54903 = ~\P1_P2_rEIP_reg[10]/NET0131  & ~n51239 ;
  assign n54904 = ~n54902 & ~n54903 ;
  assign n54905 = n48443 & ~n54904 ;
  assign n54906 = ~\P1_P2_EBX_reg[10]/NET0131  & ~n48443 ;
  assign n54907 = ~n54905 & ~n54906 ;
  assign n54908 = n25757 & n54907 ;
  assign n54910 = \P1_P2_EBX_reg[31]/NET0131  & ~n48415 ;
  assign n54912 = ~\P1_P2_EBX_reg[10]/NET0131  & n54910 ;
  assign n54911 = \P1_P2_EBX_reg[10]/NET0131  & ~n54910 ;
  assign n54913 = ~n48373 & ~n54911 ;
  assign n54914 = ~n54912 & n54913 ;
  assign n54909 = n48373 & ~n54904 ;
  assign n54915 = n25776 & ~n54909 ;
  assign n54916 = ~n54914 & n54915 ;
  assign n54917 = ~n54908 & ~n54916 ;
  assign n54918 = ~n25770 & ~n54917 ;
  assign n54919 = ~n54901 & ~n54918 ;
  assign n54920 = n25918 & ~n54919 ;
  assign n54890 = \P1_P2_rEIP_reg[10]/NET0131  & ~n53566 ;
  assign n54921 = \P1_P2_PhyAddrPointer_reg[10]/NET0131  & n27675 ;
  assign n54922 = ~n27967 & ~n54921 ;
  assign n54923 = ~n54890 & n54922 ;
  assign n54924 = ~n54920 & n54923 ;
  assign n54925 = ~n54900 & n54924 ;
  assign n54928 = n36650 & n50476 ;
  assign n54929 = n36672 & ~n54928 ;
  assign n54931 = n41514 & ~n54929 ;
  assign n54930 = ~n41514 & n54929 ;
  assign n54932 = ~\P2_P1_DataWidth_reg[1]/NET0131  & ~n54930 ;
  assign n54933 = ~n54931 & n54932 ;
  assign n54927 = \P2_P1_DataWidth_reg[1]/NET0131  & ~\P2_P1_rEIP_reg[11]/NET0131  ;
  assign n54934 = n11609 & ~n54927 ;
  assign n54935 = ~n54933 & n54934 ;
  assign n54936 = \P2_P1_rEIP_reg[11]/NET0131  & ~n50414 ;
  assign n54938 = ~\P2_P1_rEIP_reg[11]/NET0131  & ~n54867 ;
  assign n54939 = ~n50773 & ~n54938 ;
  assign n54940 = n50422 & ~n54939 ;
  assign n54941 = ~n25958 & n54940 ;
  assign n54937 = ~\P2_P1_EBX_reg[11]/NET0131  & ~n26103 ;
  assign n54942 = n24898 & ~n54937 ;
  assign n54943 = ~n54941 & n54942 ;
  assign n54944 = \P2_P1_EBX_reg[31]/NET0131  & ~n50796 ;
  assign n54946 = \P2_P1_EBX_reg[11]/NET0131  & ~n54944 ;
  assign n54945 = ~\P2_P1_EBX_reg[11]/NET0131  & n54944 ;
  assign n54947 = ~n50422 & ~n54945 ;
  assign n54948 = ~n54946 & n54947 ;
  assign n54949 = n21062 & ~n54940 ;
  assign n54950 = ~n54948 & n54949 ;
  assign n54951 = ~n54943 & ~n54950 ;
  assign n54952 = ~n21081 & ~n54951 ;
  assign n54953 = ~n54936 & ~n54952 ;
  assign n54954 = n11623 & ~n54953 ;
  assign n54926 = \P2_P1_rEIP_reg[11]/NET0131  & ~n53464 ;
  assign n54955 = \P2_P1_PhyAddrPointer_reg[11]/NET0131  & n11625 ;
  assign n54956 = ~n11616 & ~n54955 ;
  assign n54957 = ~n54926 & n54956 ;
  assign n54958 = ~n54954 & n54957 ;
  assign n54959 = ~n54935 & n54958 ;
  assign n54962 = n36672 & ~n50824 ;
  assign n54964 = ~n43436 & n54962 ;
  assign n54963 = n43436 & ~n54962 ;
  assign n54965 = ~\P2_P1_DataWidth_reg[1]/NET0131  & ~n54963 ;
  assign n54966 = ~n54964 & n54965 ;
  assign n54961 = \P2_P1_DataWidth_reg[1]/NET0131  & ~\P2_P1_rEIP_reg[12]/NET0131  ;
  assign n54967 = n11609 & ~n54961 ;
  assign n54968 = ~n54966 & n54967 ;
  assign n54978 = \P2_P1_EBX_reg[31]/NET0131  & ~n50797 ;
  assign n54980 = ~\P2_P1_EBX_reg[12]/NET0131  & n54978 ;
  assign n54979 = \P2_P1_EBX_reg[12]/NET0131  & ~n54978 ;
  assign n54981 = ~n50422 & ~n54979 ;
  assign n54982 = ~n54980 & n54981 ;
  assign n54971 = \P2_P1_rEIP_reg[12]/NET0131  & n50773 ;
  assign n54972 = ~\P2_P1_rEIP_reg[12]/NET0131  & ~n50773 ;
  assign n54973 = ~n54971 & ~n54972 ;
  assign n54977 = n50422 & ~n54973 ;
  assign n54983 = n24901 & ~n54977 ;
  assign n54984 = ~n54982 & n54983 ;
  assign n54969 = \P2_P1_rEIP_reg[12]/NET0131  & ~n50414 ;
  assign n54970 = ~\P2_P1_EBX_reg[12]/NET0131  & ~n26103 ;
  assign n54974 = n26103 & ~n54973 ;
  assign n54975 = ~n54970 & ~n54974 ;
  assign n54976 = n24899 & n54975 ;
  assign n54985 = ~n54969 & ~n54976 ;
  assign n54986 = ~n54984 & n54985 ;
  assign n54987 = n11623 & ~n54986 ;
  assign n54960 = \P2_P1_rEIP_reg[12]/NET0131  & ~n53464 ;
  assign n54988 = \P2_P1_PhyAddrPointer_reg[12]/NET0131  & n11625 ;
  assign n54989 = ~n11616 & ~n54988 ;
  assign n54990 = ~n54960 & n54989 ;
  assign n54991 = ~n54987 & n54990 ;
  assign n54992 = ~n54968 & n54991 ;
  assign n54996 = n41373 & ~n51181 ;
  assign n54995 = ~n41373 & n51181 ;
  assign n54997 = ~\P1_P2_DataWidth_reg[1]/NET0131  & ~n54995 ;
  assign n54998 = ~n54996 & n54997 ;
  assign n54994 = \P1_P2_DataWidth_reg[1]/NET0131  & ~\P1_P2_rEIP_reg[11]/NET0131  ;
  assign n54999 = n25928 & ~n54994 ;
  assign n55000 = ~n54998 & n54999 ;
  assign n55001 = \P1_P2_rEIP_reg[11]/NET0131  & ~n48371 ;
  assign n55003 = ~\P1_P2_rEIP_reg[11]/NET0131  & ~n54902 ;
  assign n55004 = ~n51240 & ~n55003 ;
  assign n55005 = n48373 & ~n55004 ;
  assign n55006 = ~n25768 & n55005 ;
  assign n55002 = ~\P1_P2_EBX_reg[11]/NET0131  & ~n48443 ;
  assign n55007 = n25757 & ~n55002 ;
  assign n55008 = ~n55006 & n55007 ;
  assign n55009 = \P1_P2_EBX_reg[31]/NET0131  & ~n48416 ;
  assign n55011 = ~\P1_P2_EBX_reg[11]/NET0131  & n55009 ;
  assign n55010 = \P1_P2_EBX_reg[11]/NET0131  & ~n55009 ;
  assign n55012 = ~n48373 & ~n55010 ;
  assign n55013 = ~n55011 & n55012 ;
  assign n55014 = n25776 & ~n55005 ;
  assign n55015 = ~n55013 & n55014 ;
  assign n55016 = ~n55008 & ~n55015 ;
  assign n55017 = ~n25770 & ~n55016 ;
  assign n55018 = ~n55001 & ~n55017 ;
  assign n55019 = n25918 & ~n55018 ;
  assign n54993 = \P1_P2_rEIP_reg[11]/NET0131  & ~n53566 ;
  assign n55020 = \P1_P2_PhyAddrPointer_reg[11]/NET0131  & n27675 ;
  assign n55021 = ~n27967 & ~n55020 ;
  assign n55022 = ~n54993 & n55021 ;
  assign n55023 = ~n55019 & n55022 ;
  assign n55024 = ~n55000 & n55023 ;
  assign n55027 = n41527 & n50476 ;
  assign n55028 = n36672 & ~n55027 ;
  assign n55030 = n43444 & ~n55028 ;
  assign n55029 = ~n43444 & n55028 ;
  assign n55031 = ~\P2_P1_DataWidth_reg[1]/NET0131  & ~n55029 ;
  assign n55032 = ~n55030 & n55031 ;
  assign n55026 = \P2_P1_DataWidth_reg[1]/NET0131  & ~\P2_P1_rEIP_reg[13]/NET0131  ;
  assign n55033 = n11609 & ~n55026 ;
  assign n55034 = ~n55032 & n55033 ;
  assign n55043 = \P2_P1_EBX_reg[31]/NET0131  & ~n50798 ;
  assign n55045 = ~\P2_P1_EBX_reg[13]/NET0131  & n55043 ;
  assign n55044 = \P2_P1_EBX_reg[13]/NET0131  & ~n55043 ;
  assign n55046 = ~n50422 & ~n55044 ;
  assign n55047 = ~n55045 & n55046 ;
  assign n55037 = ~\P2_P1_rEIP_reg[13]/NET0131  & ~n54971 ;
  assign n55038 = ~n50774 & ~n55037 ;
  assign n55042 = n50422 & ~n55038 ;
  assign n55048 = n24901 & ~n55042 ;
  assign n55049 = ~n55047 & n55048 ;
  assign n55035 = \P2_P1_rEIP_reg[13]/NET0131  & ~n50414 ;
  assign n55039 = n26103 & ~n55038 ;
  assign n55036 = ~\P2_P1_EBX_reg[13]/NET0131  & ~n26103 ;
  assign n55040 = n24899 & ~n55036 ;
  assign n55041 = ~n55039 & n55040 ;
  assign n55050 = ~n55035 & ~n55041 ;
  assign n55051 = ~n55049 & n55050 ;
  assign n55052 = n11623 & ~n55051 ;
  assign n55025 = \P2_P1_rEIP_reg[13]/NET0131  & ~n53464 ;
  assign n55053 = \P2_P1_PhyAddrPointer_reg[13]/NET0131  & n11625 ;
  assign n55054 = ~n11616 & ~n55053 ;
  assign n55055 = ~n55025 & n55054 ;
  assign n55056 = ~n55052 & n55055 ;
  assign n55057 = ~n55034 & n55056 ;
  assign n55060 = n36672 & ~n50751 ;
  assign n55062 = n41533 & ~n55060 ;
  assign n55061 = ~n41533 & n55060 ;
  assign n55063 = ~\P2_P1_DataWidth_reg[1]/NET0131  & ~n55061 ;
  assign n55064 = ~n55062 & n55063 ;
  assign n55059 = \P2_P1_DataWidth_reg[1]/NET0131  & ~\P2_P1_rEIP_reg[14]/NET0131  ;
  assign n55065 = n11609 & ~n55059 ;
  assign n55066 = ~n55064 & n55065 ;
  assign n55067 = \P2_P1_rEIP_reg[14]/NET0131  & ~n50414 ;
  assign n55069 = ~\P2_P1_rEIP_reg[14]/NET0131  & ~n50774 ;
  assign n55070 = ~n50775 & ~n55069 ;
  assign n55071 = n26103 & ~n55070 ;
  assign n55068 = ~\P2_P1_EBX_reg[14]/NET0131  & ~n26103 ;
  assign n55072 = n24898 & ~n55068 ;
  assign n55073 = ~n55071 & n55072 ;
  assign n55075 = \P2_P1_EBX_reg[31]/NET0131  & ~n50799 ;
  assign n55077 = ~\P2_P1_EBX_reg[14]/NET0131  & n55075 ;
  assign n55076 = \P2_P1_EBX_reg[14]/NET0131  & ~n55075 ;
  assign n55078 = ~n50422 & ~n55076 ;
  assign n55079 = ~n55077 & n55078 ;
  assign n55074 = n50422 & ~n55070 ;
  assign n55080 = n21062 & ~n55074 ;
  assign n55081 = ~n55079 & n55080 ;
  assign n55082 = ~n55073 & ~n55081 ;
  assign n55083 = ~n21081 & ~n55082 ;
  assign n55084 = ~n55067 & ~n55083 ;
  assign n55085 = n11623 & ~n55084 ;
  assign n55058 = \P2_P1_rEIP_reg[14]/NET0131  & ~n53464 ;
  assign n55086 = \P2_P1_PhyAddrPointer_reg[14]/NET0131  & n11625 ;
  assign n55087 = ~n11616 & ~n55086 ;
  assign n55088 = ~n55058 & n55087 ;
  assign n55089 = ~n55085 & n55088 ;
  assign n55090 = ~n55066 & n55089 ;
  assign n55093 = ~n36628 & ~n41372 ;
  assign n55094 = ~n54892 & ~n55093 ;
  assign n55096 = n43295 & n55094 ;
  assign n55095 = ~n43295 & ~n55094 ;
  assign n55097 = ~\P1_P2_DataWidth_reg[1]/NET0131  & ~n55095 ;
  assign n55098 = ~n55096 & n55097 ;
  assign n55092 = \P1_P2_DataWidth_reg[1]/NET0131  & ~\P1_P2_rEIP_reg[12]/NET0131  ;
  assign n55099 = n25928 & ~n55092 ;
  assign n55100 = ~n55098 & n55099 ;
  assign n55101 = \P1_P2_rEIP_reg[12]/NET0131  & ~n48371 ;
  assign n55103 = \P1_P2_rEIP_reg[12]/NET0131  & n51240 ;
  assign n55104 = ~\P1_P2_rEIP_reg[12]/NET0131  & ~n51240 ;
  assign n55105 = ~n55103 & ~n55104 ;
  assign n55106 = n48373 & ~n55105 ;
  assign n55107 = ~n25768 & n55106 ;
  assign n55102 = ~\P1_P2_EBX_reg[12]/NET0131  & ~n48443 ;
  assign n55108 = n25757 & ~n55102 ;
  assign n55109 = ~n55107 & n55108 ;
  assign n55110 = \P1_P2_EBX_reg[31]/NET0131  & ~n48417 ;
  assign n55112 = \P1_P2_EBX_reg[12]/NET0131  & ~n55110 ;
  assign n55111 = ~\P1_P2_EBX_reg[12]/NET0131  & n55110 ;
  assign n55113 = ~n48373 & ~n55111 ;
  assign n55114 = ~n55112 & n55113 ;
  assign n55115 = n25776 & ~n55106 ;
  assign n55116 = ~n55114 & n55115 ;
  assign n55117 = ~n55109 & ~n55116 ;
  assign n55118 = ~n25770 & ~n55117 ;
  assign n55119 = ~n55101 & ~n55118 ;
  assign n55120 = n25918 & ~n55119 ;
  assign n55091 = \P1_P2_rEIP_reg[12]/NET0131  & ~n53566 ;
  assign n55121 = \P1_P2_PhyAddrPointer_reg[12]/NET0131  & n27675 ;
  assign n55122 = ~n27967 & ~n55121 ;
  assign n55123 = ~n55091 & n55122 ;
  assign n55124 = ~n55120 & n55123 ;
  assign n55125 = ~n55100 & n55124 ;
  assign n55128 = n36672 & ~n50753 ;
  assign n55130 = ~n43476 & n55128 ;
  assign n55129 = n43476 & ~n55128 ;
  assign n55131 = ~\P2_P1_DataWidth_reg[1]/NET0131  & ~n55129 ;
  assign n55132 = ~n55130 & n55131 ;
  assign n55127 = \P2_P1_DataWidth_reg[1]/NET0131  & ~\P2_P1_rEIP_reg[16]/NET0131  ;
  assign n55133 = n11609 & ~n55127 ;
  assign n55134 = ~n55132 & n55133 ;
  assign n55135 = \P2_P1_rEIP_reg[16]/NET0131  & ~n50414 ;
  assign n55138 = ~\P2_P1_EBX_reg[16]/NET0131  & ~n26103 ;
  assign n55139 = n24898 & ~n55138 ;
  assign n55143 = \P2_P1_EBX_reg[31]/NET0131  & ~n50801 ;
  assign n55145 = ~\P2_P1_EBX_reg[16]/NET0131  & n55143 ;
  assign n55144 = \P2_P1_EBX_reg[16]/NET0131  & ~n55143 ;
  assign n55146 = ~n50422 & ~n55144 ;
  assign n55147 = ~n55145 & n55146 ;
  assign n55148 = n21062 & ~n55147 ;
  assign n55149 = ~n55139 & ~n55148 ;
  assign n55140 = n25958 & n55139 ;
  assign n55136 = ~\P2_P1_rEIP_reg[16]/NET0131  & ~n53474 ;
  assign n55137 = ~n53510 & ~n55136 ;
  assign n55141 = n50422 & ~n55137 ;
  assign n55142 = ~n55140 & n55141 ;
  assign n55150 = ~n21081 & ~n55142 ;
  assign n55151 = ~n55149 & n55150 ;
  assign n55152 = ~n55135 & ~n55151 ;
  assign n55153 = n11623 & ~n55152 ;
  assign n55126 = \P2_P1_rEIP_reg[16]/NET0131  & ~n53464 ;
  assign n55154 = \P2_P1_PhyAddrPointer_reg[16]/NET0131  & n11625 ;
  assign n55155 = ~n11616 & ~n55154 ;
  assign n55156 = ~n55126 & n55155 ;
  assign n55157 = ~n55153 & n55156 ;
  assign n55158 = ~n55134 & n55157 ;
  assign n55161 = ~n36628 & ~n43293 ;
  assign n55162 = ~n51181 & ~n55161 ;
  assign n55164 = n43323 & n55162 ;
  assign n55163 = ~n43323 & ~n55162 ;
  assign n55165 = ~\P1_P2_DataWidth_reg[1]/NET0131  & ~n55163 ;
  assign n55166 = ~n55164 & n55165 ;
  assign n55160 = \P1_P2_DataWidth_reg[1]/NET0131  & ~\P1_P2_rEIP_reg[13]/NET0131  ;
  assign n55167 = n25928 & ~n55160 ;
  assign n55168 = ~n55166 & n55167 ;
  assign n55169 = \P1_P2_rEIP_reg[13]/NET0131  & ~n48371 ;
  assign n55171 = ~\P1_P2_rEIP_reg[13]/NET0131  & ~n55103 ;
  assign n55172 = \P1_P2_rEIP_reg[13]/NET0131  & n55103 ;
  assign n55173 = ~n55171 & ~n55172 ;
  assign n55174 = n48443 & ~n55173 ;
  assign n55170 = ~\P1_P2_EBX_reg[13]/NET0131  & ~n48443 ;
  assign n55175 = n25757 & ~n55170 ;
  assign n55176 = ~n55174 & n55175 ;
  assign n55178 = \P1_P2_EBX_reg[31]/NET0131  & ~n48418 ;
  assign n55179 = ~\P1_P2_EBX_reg[13]/NET0131  & ~n55178 ;
  assign n55180 = \P1_P2_EBX_reg[13]/NET0131  & n55178 ;
  assign n55181 = ~n55179 & ~n55180 ;
  assign n55182 = ~n48373 & ~n55181 ;
  assign n55177 = n48373 & ~n55173 ;
  assign n55183 = n25776 & ~n55177 ;
  assign n55184 = ~n55182 & n55183 ;
  assign n55185 = ~n55176 & ~n55184 ;
  assign n55186 = ~n25770 & ~n55185 ;
  assign n55187 = ~n55169 & ~n55186 ;
  assign n55188 = n25918 & ~n55187 ;
  assign n55159 = \P1_P2_rEIP_reg[13]/NET0131  & ~n53566 ;
  assign n55189 = \P1_P2_PhyAddrPointer_reg[13]/NET0131  & n27675 ;
  assign n55190 = ~n27967 & ~n55189 ;
  assign n55191 = ~n55159 & n55190 ;
  assign n55192 = ~n55188 & n55191 ;
  assign n55193 = ~n55168 & n55192 ;
  assign n55196 = n36672 & ~n50859 ;
  assign n55198 = ~n41553 & n55196 ;
  assign n55197 = n41553 & ~n55196 ;
  assign n55199 = ~\P2_P1_DataWidth_reg[1]/NET0131  & ~n55197 ;
  assign n55200 = ~n55198 & n55199 ;
  assign n55195 = \P2_P1_DataWidth_reg[1]/NET0131  & ~\P2_P1_rEIP_reg[19]/NET0131  ;
  assign n55201 = n11609 & ~n55195 ;
  assign n55202 = ~n55200 & n55201 ;
  assign n55211 = \P2_P1_EBX_reg[31]/NET0131  & ~n50804 ;
  assign n55213 = ~\P2_P1_EBX_reg[19]/NET0131  & n55211 ;
  assign n55212 = \P2_P1_EBX_reg[19]/NET0131  & ~n55211 ;
  assign n55214 = ~n50422 & ~n55212 ;
  assign n55215 = ~n55213 & n55214 ;
  assign n55205 = ~\P2_P1_rEIP_reg[19]/NET0131  & ~n50777 ;
  assign n55206 = ~n50778 & ~n55205 ;
  assign n55207 = n50422 & ~n55206 ;
  assign n55216 = n24901 & ~n55207 ;
  assign n55217 = ~n55215 & n55216 ;
  assign n55203 = \P2_P1_rEIP_reg[19]/NET0131  & ~n50414 ;
  assign n55208 = ~n25958 & n55207 ;
  assign n55204 = ~\P2_P1_EBX_reg[19]/NET0131  & ~n26103 ;
  assign n55209 = n24899 & ~n55204 ;
  assign n55210 = ~n55208 & n55209 ;
  assign n55218 = ~n55203 & ~n55210 ;
  assign n55219 = ~n55217 & n55218 ;
  assign n55220 = n11623 & ~n55219 ;
  assign n55194 = \P2_P1_rEIP_reg[19]/NET0131  & ~n53464 ;
  assign n55221 = \P2_P1_PhyAddrPointer_reg[19]/NET0131  & n11625 ;
  assign n55222 = ~n11616 & ~n55221 ;
  assign n55223 = ~n55194 & n55222 ;
  assign n55224 = ~n55220 & n55223 ;
  assign n55225 = ~n55202 & n55224 ;
  assign n55229 = n41395 & n53571 ;
  assign n55228 = ~n41395 & ~n53571 ;
  assign n55230 = ~\P1_P2_DataWidth_reg[1]/NET0131  & ~n55228 ;
  assign n55231 = ~n55229 & n55230 ;
  assign n55227 = \P1_P2_DataWidth_reg[1]/NET0131  & ~\P1_P2_rEIP_reg[14]/NET0131  ;
  assign n55232 = n25928 & ~n55227 ;
  assign n55233 = ~n55231 & n55232 ;
  assign n55234 = \P1_P2_rEIP_reg[14]/NET0131  & ~n48371 ;
  assign n55236 = ~\P1_P2_rEIP_reg[14]/NET0131  & ~n55172 ;
  assign n55237 = ~n53579 & ~n55236 ;
  assign n55238 = n48373 & ~n55237 ;
  assign n55239 = ~n25768 & n55238 ;
  assign n55235 = ~\P1_P2_EBX_reg[14]/NET0131  & ~n48443 ;
  assign n55240 = n25757 & ~n55235 ;
  assign n55241 = ~n55239 & n55240 ;
  assign n55242 = \P1_P2_EBX_reg[31]/NET0131  & ~n48419 ;
  assign n55244 = ~\P1_P2_EBX_reg[14]/NET0131  & n55242 ;
  assign n55243 = \P1_P2_EBX_reg[14]/NET0131  & ~n55242 ;
  assign n55245 = ~n48373 & ~n55243 ;
  assign n55246 = ~n55244 & n55245 ;
  assign n55247 = n25776 & ~n55238 ;
  assign n55248 = ~n55246 & n55247 ;
  assign n55249 = ~n55241 & ~n55248 ;
  assign n55250 = ~n25770 & ~n55249 ;
  assign n55251 = ~n55234 & ~n55250 ;
  assign n55252 = n25918 & ~n55251 ;
  assign n55226 = \P1_P2_rEIP_reg[14]/NET0131  & ~n53566 ;
  assign n55253 = \P1_P2_PhyAddrPointer_reg[14]/NET0131  & n27675 ;
  assign n55254 = ~n27967 & ~n55253 ;
  assign n55255 = ~n55226 & n55254 ;
  assign n55256 = ~n55252 & n55255 ;
  assign n55257 = ~n55233 & n55256 ;
  assign n55260 = ~n36628 & ~n39336 ;
  assign n55261 = ~n51181 & ~n55260 ;
  assign n55263 = n43332 & n55261 ;
  assign n55262 = ~n43332 & ~n55261 ;
  assign n55264 = ~\P1_P2_DataWidth_reg[1]/NET0131  & ~n55262 ;
  assign n55265 = ~n55263 & n55264 ;
  assign n55259 = \P1_P2_DataWidth_reg[1]/NET0131  & ~\P1_P2_rEIP_reg[16]/NET0131  ;
  assign n55266 = n25928 & ~n55259 ;
  assign n55267 = ~n55265 & n55266 ;
  assign n55281 = \P1_P2_EBX_reg[31]/NET0131  & ~n48421 ;
  assign n55283 = ~\P1_P2_EBX_reg[16]/NET0131  & n55281 ;
  assign n55282 = \P1_P2_EBX_reg[16]/NET0131  & ~n55281 ;
  assign n55284 = ~n48373 & ~n55282 ;
  assign n55285 = ~n55283 & n55284 ;
  assign n55273 = ~\P1_P2_rEIP_reg[16]/NET0131  & n51201 ;
  assign n55272 = \P1_P2_rEIP_reg[16]/NET0131  & ~n51201 ;
  assign n55274 = n48373 & ~n55272 ;
  assign n55275 = ~n55273 & n55274 ;
  assign n55286 = n25846 & ~n55275 ;
  assign n55287 = ~n55285 & n55286 ;
  assign n55268 = \P1_P2_rEIP_reg[16]/NET0131  & n51192 ;
  assign n55271 = ~\P1_P2_EBX_reg[16]/NET0131  & ~n48373 ;
  assign n55276 = ~n55271 & ~n55275 ;
  assign n55277 = n25841 & n55276 ;
  assign n55269 = \P1_P2_EBX_reg[16]/NET0131  & n51194 ;
  assign n55270 = \P1_P2_rEIP_reg[16]/NET0131  & n25770 ;
  assign n55278 = ~n55269 & ~n55270 ;
  assign n55279 = ~n55277 & n55278 ;
  assign n55280 = n25757 & ~n55279 ;
  assign n55288 = ~n55268 & ~n55280 ;
  assign n55289 = ~n55287 & n55288 ;
  assign n55290 = n25918 & ~n55289 ;
  assign n55258 = \P1_P2_rEIP_reg[16]/NET0131  & ~n53566 ;
  assign n55291 = \P1_P2_PhyAddrPointer_reg[16]/NET0131  & n27675 ;
  assign n55292 = ~n27967 & ~n55291 ;
  assign n55293 = ~n55258 & n55292 ;
  assign n55294 = ~n55290 & n55293 ;
  assign n55295 = ~n55267 & n55294 ;
  assign n55299 = n41416 & n51183 ;
  assign n55298 = ~n41416 & ~n51183 ;
  assign n55300 = ~\P1_P2_DataWidth_reg[1]/NET0131  & ~n55298 ;
  assign n55301 = ~n55299 & n55300 ;
  assign n55297 = \P1_P2_DataWidth_reg[1]/NET0131  & ~\P1_P2_rEIP_reg[19]/NET0131  ;
  assign n55302 = n25928 & ~n55297 ;
  assign n55303 = ~n55301 & n55302 ;
  assign n55308 = \P1_P2_EBX_reg[31]/NET0131  & ~n48424 ;
  assign n55310 = \P1_P2_EBX_reg[19]/NET0131  & ~n55308 ;
  assign n55309 = ~\P1_P2_EBX_reg[19]/NET0131  & n55308 ;
  assign n55311 = ~n48373 & ~n55309 ;
  assign n55312 = ~n55310 & n55311 ;
  assign n55305 = ~\P1_P2_rEIP_reg[19]/NET0131  & ~n51202 ;
  assign n55306 = ~n51203 & ~n55305 ;
  assign n55307 = n48373 & ~n55306 ;
  assign n55313 = n25846 & ~n55307 ;
  assign n55314 = ~n55312 & n55313 ;
  assign n55304 = \P1_P2_rEIP_reg[19]/NET0131  & ~n48371 ;
  assign n55315 = n48443 & ~n55306 ;
  assign n55316 = ~\P1_P2_EBX_reg[19]/NET0131  & ~n48443 ;
  assign n55317 = ~n55315 & ~n55316 ;
  assign n55318 = n47570 & n55317 ;
  assign n55319 = ~n55304 & ~n55318 ;
  assign n55320 = ~n55314 & n55319 ;
  assign n55321 = n25918 & ~n55320 ;
  assign n55296 = \P1_P2_rEIP_reg[19]/NET0131  & ~n53566 ;
  assign n55322 = \P1_P2_PhyAddrPointer_reg[19]/NET0131  & n27675 ;
  assign n55323 = ~n27967 & ~n55322 ;
  assign n55324 = ~n55296 & n55323 ;
  assign n55325 = ~n55321 & n55324 ;
  assign n55326 = ~n55303 & n55325 ;
  assign n55329 = n36647 & n50476 ;
  assign n55330 = n36672 & ~n55329 ;
  assign n55332 = n43580 & ~n55330 ;
  assign n55331 = ~n43580 & n55330 ;
  assign n55333 = ~\P2_P1_DataWidth_reg[1]/NET0131  & ~n55331 ;
  assign n55334 = ~n55332 & n55333 ;
  assign n55328 = \P2_P1_DataWidth_reg[1]/NET0131  & ~\P2_P1_rEIP_reg[8]/NET0131  ;
  assign n55335 = n11609 & ~n55328 ;
  assign n55336 = ~n55334 & n55335 ;
  assign n55337 = \P2_P1_rEIP_reg[8]/NET0131  & ~n50414 ;
  assign n55338 = ~\P2_P1_EBX_reg[8]/NET0131  & ~n26103 ;
  assign n55339 = ~\P2_P1_rEIP_reg[8]/NET0131  & ~n50769 ;
  assign n55340 = ~n50770 & ~n55339 ;
  assign n55341 = n26103 & ~n55340 ;
  assign n55342 = ~n55338 & ~n55341 ;
  assign n55343 = n24899 & n55342 ;
  assign n55344 = n50422 & ~n55340 ;
  assign n55345 = \P2_P1_EBX_reg[31]/NET0131  & ~n50793 ;
  assign n55347 = ~\P2_P1_EBX_reg[8]/NET0131  & n55345 ;
  assign n55346 = \P2_P1_EBX_reg[8]/NET0131  & ~n55345 ;
  assign n55348 = ~n50422 & ~n55346 ;
  assign n55349 = ~n55347 & n55348 ;
  assign n55350 = ~n55344 & ~n55349 ;
  assign n55351 = n24901 & n55350 ;
  assign n55352 = ~n55343 & ~n55351 ;
  assign n55353 = ~n55337 & n55352 ;
  assign n55354 = n11623 & ~n55353 ;
  assign n55327 = \P2_P1_rEIP_reg[8]/NET0131  & ~n53464 ;
  assign n55355 = \P2_P1_PhyAddrPointer_reg[8]/NET0131  & n11625 ;
  assign n55356 = ~n11616 & ~n55355 ;
  assign n55357 = ~n55327 & n55356 ;
  assign n55358 = ~n55354 & n55357 ;
  assign n55359 = ~n55336 & n55358 ;
  assign n55362 = ~\P2_P1_PhyAddrPointer_reg[0]/NET0131  & n39454 ;
  assign n55363 = n36672 & ~n55362 ;
  assign n55365 = n44980 & ~n55363 ;
  assign n55364 = ~n44980 & n55363 ;
  assign n55366 = ~\P2_P1_DataWidth_reg[1]/NET0131  & ~n55364 ;
  assign n55367 = ~n55365 & n55366 ;
  assign n55361 = \P2_P1_DataWidth_reg[1]/NET0131  & ~\P2_P1_rEIP_reg[9]/NET0131  ;
  assign n55368 = n11609 & ~n55361 ;
  assign n55369 = ~n55367 & n55368 ;
  assign n55370 = \P2_P1_rEIP_reg[9]/NET0131  & ~n50414 ;
  assign n55371 = ~\P2_P1_EBX_reg[9]/NET0131  & ~n26103 ;
  assign n55372 = ~\P2_P1_rEIP_reg[9]/NET0131  & ~n50770 ;
  assign n55373 = ~n50771 & ~n55372 ;
  assign n55374 = n26103 & ~n55373 ;
  assign n55375 = ~n55371 & ~n55374 ;
  assign n55376 = n24899 & n55375 ;
  assign n55377 = n50422 & ~n55373 ;
  assign n55378 = \P2_P1_EBX_reg[31]/NET0131  & ~n50794 ;
  assign n55380 = ~\P2_P1_EBX_reg[9]/NET0131  & n55378 ;
  assign n55379 = \P2_P1_EBX_reg[9]/NET0131  & ~n55378 ;
  assign n55381 = ~n50422 & ~n55379 ;
  assign n55382 = ~n55380 & n55381 ;
  assign n55383 = ~n55377 & ~n55382 ;
  assign n55384 = n24901 & n55383 ;
  assign n55385 = ~n55376 & ~n55384 ;
  assign n55386 = ~n55370 & n55385 ;
  assign n55387 = n11623 & ~n55386 ;
  assign n55360 = \P2_P1_rEIP_reg[9]/NET0131  & ~n53464 ;
  assign n55388 = \P2_P1_PhyAddrPointer_reg[9]/NET0131  & n11625 ;
  assign n55389 = ~n11616 & ~n55388 ;
  assign n55390 = ~n55360 & n55389 ;
  assign n55391 = ~n55387 & n55390 ;
  assign n55392 = ~n55369 & n55391 ;
  assign n55396 = ~n43521 & n54892 ;
  assign n55395 = n43521 & ~n54892 ;
  assign n55397 = ~\P1_P2_DataWidth_reg[1]/NET0131  & ~n55395 ;
  assign n55398 = ~n55396 & n55397 ;
  assign n55394 = \P1_P2_DataWidth_reg[1]/NET0131  & ~\P1_P2_rEIP_reg[8]/NET0131  ;
  assign n55399 = n25928 & ~n55394 ;
  assign n55400 = ~n55398 & n55399 ;
  assign n55401 = \P1_P2_rEIP_reg[8]/NET0131  & ~n48371 ;
  assign n55402 = ~\P1_P2_rEIP_reg[8]/NET0131  & ~n48385 ;
  assign n55403 = ~n48386 & ~n55402 ;
  assign n55404 = n48443 & ~n55403 ;
  assign n55405 = ~\P1_P2_EBX_reg[8]/NET0131  & ~n48443 ;
  assign n55406 = ~n55404 & ~n55405 ;
  assign n55407 = n25757 & n55406 ;
  assign n55408 = n48373 & ~n55403 ;
  assign n55409 = \P1_P2_EBX_reg[31]/NET0131  & ~n48413 ;
  assign n55411 = ~\P1_P2_EBX_reg[8]/NET0131  & n55409 ;
  assign n55410 = \P1_P2_EBX_reg[8]/NET0131  & ~n55409 ;
  assign n55412 = ~n48373 & ~n55410 ;
  assign n55413 = ~n55411 & n55412 ;
  assign n55414 = ~n55408 & ~n55413 ;
  assign n55415 = n25776 & n55414 ;
  assign n55416 = ~n55407 & ~n55415 ;
  assign n55417 = ~n25770 & ~n55416 ;
  assign n55418 = ~n55401 & ~n55417 ;
  assign n55419 = n25918 & ~n55418 ;
  assign n55393 = \P1_P2_rEIP_reg[8]/NET0131  & ~n53566 ;
  assign n55420 = \P1_P2_PhyAddrPointer_reg[8]/NET0131  & n27675 ;
  assign n55421 = ~n27967 & ~n55420 ;
  assign n55422 = ~n55393 & n55421 ;
  assign n55423 = ~n55419 & n55422 ;
  assign n55424 = ~n55400 & n55423 ;
  assign n55427 = ~n36628 & ~n51383 ;
  assign n55429 = n44931 & ~n55427 ;
  assign n55428 = ~n44931 & n55427 ;
  assign n55430 = ~\P1_P2_DataWidth_reg[1]/NET0131  & ~n55428 ;
  assign n55431 = ~n55429 & n55430 ;
  assign n55426 = \P1_P2_DataWidth_reg[1]/NET0131  & ~\P1_P2_rEIP_reg[9]/NET0131  ;
  assign n55432 = n25928 & ~n55426 ;
  assign n55433 = ~n55431 & n55432 ;
  assign n55434 = \P1_P2_rEIP_reg[9]/NET0131  & ~n48371 ;
  assign n55435 = ~\P1_P2_rEIP_reg[9]/NET0131  & ~n48386 ;
  assign n55436 = ~n51239 & ~n55435 ;
  assign n55437 = n48443 & ~n55436 ;
  assign n55438 = ~\P1_P2_EBX_reg[9]/NET0131  & ~n48443 ;
  assign n55439 = ~n55437 & ~n55438 ;
  assign n55440 = n25757 & n55439 ;
  assign n55442 = \P1_P2_EBX_reg[31]/NET0131  & ~n48414 ;
  assign n55444 = \P1_P2_EBX_reg[9]/NET0131  & ~n55442 ;
  assign n55443 = ~\P1_P2_EBX_reg[9]/NET0131  & n55442 ;
  assign n55445 = ~n48373 & ~n55443 ;
  assign n55446 = ~n55444 & n55445 ;
  assign n55441 = n48373 & ~n55436 ;
  assign n55447 = n25776 & ~n55441 ;
  assign n55448 = ~n55446 & n55447 ;
  assign n55449 = ~n55440 & ~n55448 ;
  assign n55450 = ~n25770 & ~n55449 ;
  assign n55451 = ~n55434 & ~n55450 ;
  assign n55452 = n25918 & ~n55451 ;
  assign n55425 = \P1_P2_rEIP_reg[9]/NET0131  & ~n53566 ;
  assign n55453 = \P1_P2_PhyAddrPointer_reg[9]/NET0131  & n27675 ;
  assign n55454 = ~n27967 & ~n55453 ;
  assign n55455 = ~n55425 & n55454 ;
  assign n55456 = ~n55452 & n55455 ;
  assign n55457 = ~n55433 & n55456 ;
  assign n55460 = ~n36708 & ~n36733 ;
  assign n55461 = ~n52047 & ~n55460 ;
  assign n55463 = n44996 & n55461 ;
  assign n55462 = ~n44996 & ~n55461 ;
  assign n55464 = ~\P1_P1_DataWidth_reg[1]/NET0131  & ~n55462 ;
  assign n55465 = ~n55463 & n55464 ;
  assign n55459 = \P1_P1_DataWidth_reg[1]/NET0131  & ~\P1_P1_rEIP_reg[10]/NET0131  ;
  assign n55466 = n8282 & ~n55459 ;
  assign n55467 = ~n55465 & n55466 ;
  assign n55468 = \P1_P1_rEIP_reg[10]/NET0131  & ~n50559 ;
  assign n55470 = ~\P1_P1_rEIP_reg[10]/NET0131  & ~n51673 ;
  assign n55471 = ~n51674 & ~n55470 ;
  assign n55472 = n26275 & ~n55471 ;
  assign n55469 = ~\P1_P1_EBX_reg[10]/NET0131  & ~n26275 ;
  assign n55473 = n24502 & ~n55469 ;
  assign n55474 = ~n55472 & n55473 ;
  assign n55476 = \P1_P1_EBX_reg[31]/NET0131  & ~n51694 ;
  assign n55478 = ~\P1_P1_EBX_reg[10]/NET0131  & n55476 ;
  assign n55477 = \P1_P1_EBX_reg[10]/NET0131  & ~n55476 ;
  assign n55479 = ~n26274 & ~n55477 ;
  assign n55480 = ~n55478 & n55479 ;
  assign n55475 = n26274 & ~n55471 ;
  assign n55481 = n15334 & ~n55475 ;
  assign n55482 = ~n55480 & n55481 ;
  assign n55483 = ~n55474 & ~n55482 ;
  assign n55484 = ~n15364 & ~n55483 ;
  assign n55485 = ~n55468 & ~n55484 ;
  assign n55486 = n8355 & ~n55485 ;
  assign n55458 = \P1_P1_rEIP_reg[10]/NET0131  & ~n53883 ;
  assign n55487 = \P1_P1_PhyAddrPointer_reg[10]/NET0131  & n8361 ;
  assign n55488 = ~n8357 & ~n55487 ;
  assign n55489 = ~n55458 & n55488 ;
  assign n55490 = ~n55486 & n55489 ;
  assign n55491 = ~n55467 & n55490 ;
  assign n55494 = ~n36709 & ~n36733 ;
  assign n55495 = ~n52047 & ~n55494 ;
  assign n55497 = n41671 & n55495 ;
  assign n55496 = ~n41671 & ~n55495 ;
  assign n55498 = ~\P1_P1_DataWidth_reg[1]/NET0131  & ~n55496 ;
  assign n55499 = ~n55497 & n55498 ;
  assign n55493 = \P1_P1_DataWidth_reg[1]/NET0131  & ~\P1_P1_rEIP_reg[11]/NET0131  ;
  assign n55500 = n8282 & ~n55493 ;
  assign n55501 = ~n55499 & n55500 ;
  assign n55502 = \P1_P1_rEIP_reg[11]/NET0131  & ~n50559 ;
  assign n55503 = ~\P1_P1_rEIP_reg[11]/NET0131  & ~n51674 ;
  assign n55504 = ~n51675 & ~n55503 ;
  assign n55505 = n26274 & ~n55504 ;
  assign n55506 = ~n26158 & n55505 ;
  assign n55507 = ~\P1_P1_EBX_reg[11]/NET0131  & ~n26275 ;
  assign n55508 = n24502 & ~n55507 ;
  assign n55509 = ~n55506 & n55508 ;
  assign n55510 = \P1_P1_EBX_reg[31]/NET0131  & ~n51695 ;
  assign n55512 = \P1_P1_EBX_reg[11]/NET0131  & ~n55510 ;
  assign n55511 = ~\P1_P1_EBX_reg[11]/NET0131  & n55510 ;
  assign n55513 = ~n26274 & ~n55511 ;
  assign n55514 = ~n55512 & n55513 ;
  assign n55515 = n15334 & ~n55505 ;
  assign n55516 = ~n55514 & n55515 ;
  assign n55517 = ~n55509 & ~n55516 ;
  assign n55518 = ~n15364 & ~n55517 ;
  assign n55519 = ~n55502 & ~n55518 ;
  assign n55520 = n8355 & ~n55519 ;
  assign n55492 = \P1_P1_rEIP_reg[11]/NET0131  & ~n53883 ;
  assign n55521 = \P1_P1_PhyAddrPointer_reg[11]/NET0131  & n8361 ;
  assign n55522 = ~n8357 & ~n55521 ;
  assign n55523 = ~n55492 & n55522 ;
  assign n55524 = ~n55520 & n55523 ;
  assign n55525 = ~n55501 & n55524 ;
  assign n55528 = ~n36710 & ~n36733 ;
  assign n55529 = ~n52047 & ~n55528 ;
  assign n55531 = n43598 & n55529 ;
  assign n55530 = ~n43598 & ~n55529 ;
  assign n55532 = ~\P1_P1_DataWidth_reg[1]/NET0131  & ~n55530 ;
  assign n55533 = ~n55531 & n55532 ;
  assign n55527 = \P1_P1_DataWidth_reg[1]/NET0131  & ~\P1_P1_rEIP_reg[12]/NET0131  ;
  assign n55534 = n8282 & ~n55527 ;
  assign n55535 = ~n55533 & n55534 ;
  assign n55536 = \P1_P1_rEIP_reg[12]/NET0131  & ~n50559 ;
  assign n55538 = \P1_P1_rEIP_reg[12]/NET0131  & n51675 ;
  assign n55539 = ~\P1_P1_rEIP_reg[12]/NET0131  & ~n51675 ;
  assign n55540 = ~n55538 & ~n55539 ;
  assign n55541 = n26275 & ~n55540 ;
  assign n55537 = ~\P1_P1_EBX_reg[12]/NET0131  & ~n26275 ;
  assign n55542 = n24502 & ~n55537 ;
  assign n55543 = ~n55541 & n55542 ;
  assign n55545 = \P1_P1_EBX_reg[31]/NET0131  & ~n51696 ;
  assign n55547 = \P1_P1_EBX_reg[12]/NET0131  & ~n55545 ;
  assign n55546 = ~\P1_P1_EBX_reg[12]/NET0131  & n55545 ;
  assign n55548 = ~n26274 & ~n55546 ;
  assign n55549 = ~n55547 & n55548 ;
  assign n55544 = n26274 & ~n55540 ;
  assign n55550 = n15334 & ~n55544 ;
  assign n55551 = ~n55549 & n55550 ;
  assign n55552 = ~n55543 & ~n55551 ;
  assign n55553 = ~n15364 & ~n55552 ;
  assign n55554 = ~n55536 & ~n55553 ;
  assign n55555 = n8355 & ~n55554 ;
  assign n55526 = \P1_P1_rEIP_reg[12]/NET0131  & ~n53883 ;
  assign n55556 = \P1_P1_PhyAddrPointer_reg[12]/NET0131  & n8361 ;
  assign n55557 = ~n8357 & ~n55556 ;
  assign n55558 = ~n55526 & n55557 ;
  assign n55559 = ~n55555 & n55558 ;
  assign n55560 = ~n55535 & n55559 ;
  assign n55563 = ~\P1_P1_PhyAddrPointer_reg[0]/NET0131  & n39557 ;
  assign n55564 = ~n36733 & ~n55563 ;
  assign n55566 = n43616 & ~n55564 ;
  assign n55565 = ~n43616 & n55564 ;
  assign n55567 = ~\P1_P1_DataWidth_reg[1]/NET0131  & ~n55565 ;
  assign n55568 = ~n55566 & n55567 ;
  assign n55562 = \P1_P1_DataWidth_reg[1]/NET0131  & ~\P1_P1_rEIP_reg[13]/NET0131  ;
  assign n55569 = n8282 & ~n55562 ;
  assign n55570 = ~n55568 & n55569 ;
  assign n55571 = \P1_P1_rEIP_reg[13]/NET0131  & ~n50559 ;
  assign n55573 = ~\P1_P1_rEIP_reg[13]/NET0131  & ~n55538 ;
  assign n55574 = ~n51676 & ~n55573 ;
  assign n55575 = n26275 & ~n55574 ;
  assign n55572 = ~\P1_P1_EBX_reg[13]/NET0131  & ~n26275 ;
  assign n55576 = n24502 & ~n55572 ;
  assign n55577 = ~n55575 & n55576 ;
  assign n55579 = \P1_P1_EBX_reg[31]/NET0131  & ~n51697 ;
  assign n55580 = ~\P1_P1_EBX_reg[13]/NET0131  & ~n55579 ;
  assign n55581 = \P1_P1_EBX_reg[13]/NET0131  & n55579 ;
  assign n55582 = ~n55580 & ~n55581 ;
  assign n55583 = ~n26274 & ~n55582 ;
  assign n55578 = n26274 & ~n55574 ;
  assign n55584 = n15334 & ~n55578 ;
  assign n55585 = ~n55583 & n55584 ;
  assign n55586 = ~n55577 & ~n55585 ;
  assign n55587 = ~n15364 & ~n55586 ;
  assign n55588 = ~n55571 & ~n55587 ;
  assign n55589 = n8355 & ~n55588 ;
  assign n55561 = \P1_P1_rEIP_reg[13]/NET0131  & ~n53883 ;
  assign n55590 = \P1_P1_PhyAddrPointer_reg[13]/NET0131  & n8361 ;
  assign n55591 = ~n8357 & ~n55590 ;
  assign n55592 = ~n55561 & n55591 ;
  assign n55593 = ~n55589 & n55592 ;
  assign n55594 = ~n55570 & n55593 ;
  assign n55597 = \P1_P1_PhyAddrPointer_reg[13]/NET0131  & n55563 ;
  assign n55598 = ~n36733 & ~n55597 ;
  assign n55600 = n41679 & ~n55598 ;
  assign n55599 = ~n41679 & n55598 ;
  assign n55601 = ~\P1_P1_DataWidth_reg[1]/NET0131  & ~n55599 ;
  assign n55602 = ~n55600 & n55601 ;
  assign n55596 = \P1_P1_DataWidth_reg[1]/NET0131  & ~\P1_P1_rEIP_reg[14]/NET0131  ;
  assign n55603 = n8282 & ~n55596 ;
  assign n55604 = ~n55602 & n55603 ;
  assign n55613 = \P1_P1_EBX_reg[31]/NET0131  & ~n51698 ;
  assign n55615 = \P1_P1_EBX_reg[14]/NET0131  & ~n55613 ;
  assign n55614 = ~\P1_P1_EBX_reg[14]/NET0131  & n55613 ;
  assign n55616 = ~n26274 & ~n55614 ;
  assign n55617 = ~n55615 & n55616 ;
  assign n55607 = ~\P1_P1_rEIP_reg[14]/NET0131  & ~n51676 ;
  assign n55608 = ~n51677 & ~n55607 ;
  assign n55609 = n26274 & ~n55608 ;
  assign n55618 = n24504 & ~n55609 ;
  assign n55619 = ~n55617 & n55618 ;
  assign n55605 = \P1_P1_rEIP_reg[14]/NET0131  & ~n50559 ;
  assign n55610 = ~n26158 & n55609 ;
  assign n55606 = ~\P1_P1_EBX_reg[14]/NET0131  & ~n26275 ;
  assign n55611 = n24503 & ~n55606 ;
  assign n55612 = ~n55610 & n55611 ;
  assign n55620 = ~n55605 & ~n55612 ;
  assign n55621 = ~n55619 & n55620 ;
  assign n55622 = n8355 & ~n55621 ;
  assign n55595 = \P1_P1_rEIP_reg[14]/NET0131  & ~n53883 ;
  assign n55623 = \P1_P1_PhyAddrPointer_reg[14]/NET0131  & n8361 ;
  assign n55624 = ~n8357 & ~n55623 ;
  assign n55625 = ~n55595 & n55624 ;
  assign n55626 = ~n55622 & n55625 ;
  assign n55627 = ~n55604 & n55626 ;
  assign n55630 = n36714 & n52046 ;
  assign n55631 = ~n36733 & ~n55630 ;
  assign n55633 = ~n43647 & n55631 ;
  assign n55632 = n43647 & ~n55631 ;
  assign n55634 = ~\P1_P1_DataWidth_reg[1]/NET0131  & ~n55632 ;
  assign n55635 = ~n55633 & n55634 ;
  assign n55629 = \P1_P1_DataWidth_reg[1]/NET0131  & ~\P1_P1_rEIP_reg[16]/NET0131  ;
  assign n55636 = n8282 & ~n55629 ;
  assign n55637 = ~n55635 & n55636 ;
  assign n55638 = \P1_P1_rEIP_reg[16]/NET0131  & ~n50559 ;
  assign n55640 = ~\P1_P1_rEIP_reg[16]/NET0131  & ~n51678 ;
  assign n55641 = ~n51679 & ~n55640 ;
  assign n55642 = n26274 & ~n55641 ;
  assign n55643 = ~n26158 & n55642 ;
  assign n55639 = ~\P1_P1_EBX_reg[16]/NET0131  & ~n26275 ;
  assign n55644 = n24502 & ~n55639 ;
  assign n55645 = ~n55643 & n55644 ;
  assign n55646 = \P1_P1_EBX_reg[31]/NET0131  & ~n51700 ;
  assign n55648 = ~\P1_P1_EBX_reg[16]/NET0131  & n55646 ;
  assign n55647 = \P1_P1_EBX_reg[16]/NET0131  & ~n55646 ;
  assign n55649 = ~n26274 & ~n55647 ;
  assign n55650 = ~n55648 & n55649 ;
  assign n55651 = n15334 & ~n55642 ;
  assign n55652 = ~n55650 & n55651 ;
  assign n55653 = ~n55645 & ~n55652 ;
  assign n55654 = ~n15364 & ~n55653 ;
  assign n55655 = ~n55638 & ~n55654 ;
  assign n55656 = n8355 & ~n55655 ;
  assign n55628 = \P1_P1_rEIP_reg[16]/NET0131  & ~n53883 ;
  assign n55657 = \P1_P1_PhyAddrPointer_reg[16]/NET0131  & n8361 ;
  assign n55658 = ~n8357 & ~n55657 ;
  assign n55659 = ~n55628 & n55658 ;
  assign n55660 = ~n55656 & n55659 ;
  assign n55661 = ~n55637 & n55660 ;
  assign n55664 = ~\P1_P1_PhyAddrPointer_reg[18]/NET0131  & ~n36733 ;
  assign n55665 = ~n51763 & ~n55664 ;
  assign n55667 = ~n41716 & ~n55665 ;
  assign n55666 = n41716 & n55665 ;
  assign n55668 = ~\P1_P1_DataWidth_reg[1]/NET0131  & ~n55666 ;
  assign n55669 = ~n55667 & n55668 ;
  assign n55663 = \P1_P1_DataWidth_reg[1]/NET0131  & ~\P1_P1_rEIP_reg[19]/NET0131  ;
  assign n55670 = n8282 & ~n55663 ;
  assign n55671 = ~n55669 & n55670 ;
  assign n55672 = \P1_P1_rEIP_reg[19]/NET0131  & ~n50559 ;
  assign n55674 = ~\P1_P1_rEIP_reg[19]/NET0131  & ~n53962 ;
  assign n55675 = ~n51680 & ~n55674 ;
  assign n55676 = n26274 & ~n55675 ;
  assign n55677 = ~n26158 & n55676 ;
  assign n55673 = ~\P1_P1_EBX_reg[19]/NET0131  & ~n26275 ;
  assign n55678 = n24502 & ~n55673 ;
  assign n55679 = ~n55677 & n55678 ;
  assign n55680 = \P1_P1_EBX_reg[31]/NET0131  & ~n51703 ;
  assign n55682 = ~\P1_P1_EBX_reg[19]/NET0131  & n55680 ;
  assign n55681 = \P1_P1_EBX_reg[19]/NET0131  & ~n55680 ;
  assign n55683 = ~n26274 & ~n55681 ;
  assign n55684 = ~n55682 & n55683 ;
  assign n55685 = n15334 & ~n55676 ;
  assign n55686 = ~n55684 & n55685 ;
  assign n55687 = ~n55679 & ~n55686 ;
  assign n55688 = ~n15364 & ~n55687 ;
  assign n55689 = ~n55672 & ~n55688 ;
  assign n55690 = n8355 & ~n55689 ;
  assign n55662 = \P1_P1_rEIP_reg[19]/NET0131  & ~n53883 ;
  assign n55691 = \P1_P1_PhyAddrPointer_reg[19]/NET0131  & n8361 ;
  assign n55692 = ~n8357 & ~n55691 ;
  assign n55693 = ~n55662 & n55692 ;
  assign n55694 = ~n55690 & n55693 ;
  assign n55695 = ~n55671 & n55694 ;
  assign n55698 = \P1_P1_PhyAddrPointer_reg[7]/NET0131  & n54080 ;
  assign n55699 = ~n36733 & ~n55698 ;
  assign n55701 = n43740 & ~n55699 ;
  assign n55700 = ~n43740 & n55699 ;
  assign n55702 = ~\P1_P1_DataWidth_reg[1]/NET0131  & ~n55700 ;
  assign n55703 = ~n55701 & n55702 ;
  assign n55697 = \P1_P1_DataWidth_reg[1]/NET0131  & ~\P1_P1_rEIP_reg[8]/NET0131  ;
  assign n55704 = n8282 & ~n55697 ;
  assign n55705 = ~n55703 & n55704 ;
  assign n55706 = \P1_P1_rEIP_reg[8]/NET0131  & ~n50559 ;
  assign n55707 = ~\P1_P1_rEIP_reg[8]/NET0131  & ~n51671 ;
  assign n55708 = ~n51672 & ~n55707 ;
  assign n55709 = n26274 & ~n55708 ;
  assign n55710 = ~n26158 & n55709 ;
  assign n55711 = ~\P1_P1_EBX_reg[8]/NET0131  & ~n26275 ;
  assign n55712 = ~n55710 & ~n55711 ;
  assign n55713 = n24502 & n55712 ;
  assign n55714 = \P1_P1_EBX_reg[31]/NET0131  & ~n51692 ;
  assign n55716 = ~\P1_P1_EBX_reg[8]/NET0131  & n55714 ;
  assign n55715 = \P1_P1_EBX_reg[8]/NET0131  & ~n55714 ;
  assign n55717 = ~n26274 & ~n55715 ;
  assign n55718 = ~n55716 & n55717 ;
  assign n55719 = n15334 & ~n55709 ;
  assign n55720 = ~n55718 & n55719 ;
  assign n55721 = ~n55713 & ~n55720 ;
  assign n55722 = ~n15364 & ~n55721 ;
  assign n55723 = ~n55706 & ~n55722 ;
  assign n55724 = n8355 & ~n55723 ;
  assign n55696 = \P1_P1_rEIP_reg[8]/NET0131  & ~n53883 ;
  assign n55725 = \P1_P1_PhyAddrPointer_reg[8]/NET0131  & n8361 ;
  assign n55726 = ~n8357 & ~n55725 ;
  assign n55727 = ~n55696 & n55726 ;
  assign n55728 = ~n55724 & n55727 ;
  assign n55729 = ~n55705 & n55728 ;
  assign n55732 = ~\P1_P1_PhyAddrPointer_reg[0]/NET0131  & n41666 ;
  assign n55733 = ~n36733 & ~n55732 ;
  assign n55735 = n45036 & ~n55733 ;
  assign n55734 = ~n45036 & n55733 ;
  assign n55736 = ~\P1_P1_DataWidth_reg[1]/NET0131  & ~n55734 ;
  assign n55737 = ~n55735 & n55736 ;
  assign n55731 = \P1_P1_DataWidth_reg[1]/NET0131  & ~\P1_P1_rEIP_reg[9]/NET0131  ;
  assign n55738 = n8282 & ~n55731 ;
  assign n55739 = ~n55737 & n55738 ;
  assign n55740 = \P1_P1_rEIP_reg[9]/NET0131  & ~n50559 ;
  assign n55741 = ~\P1_P1_rEIP_reg[9]/NET0131  & ~n51672 ;
  assign n55742 = ~n51673 & ~n55741 ;
  assign n55743 = n26274 & ~n55742 ;
  assign n55744 = ~n26158 & n55743 ;
  assign n55745 = ~\P1_P1_EBX_reg[9]/NET0131  & ~n26275 ;
  assign n55746 = n24502 & ~n55745 ;
  assign n55747 = ~n55744 & n55746 ;
  assign n55748 = \P1_P1_EBX_reg[31]/NET0131  & ~n51693 ;
  assign n55750 = ~\P1_P1_EBX_reg[9]/NET0131  & n55748 ;
  assign n55749 = \P1_P1_EBX_reg[9]/NET0131  & ~n55748 ;
  assign n55751 = ~n26274 & ~n55749 ;
  assign n55752 = ~n55750 & n55751 ;
  assign n55753 = n15334 & ~n55743 ;
  assign n55754 = ~n55752 & n55753 ;
  assign n55755 = ~n55747 & ~n55754 ;
  assign n55756 = ~n15364 & ~n55755 ;
  assign n55757 = ~n55740 & ~n55756 ;
  assign n55758 = n8355 & ~n55757 ;
  assign n55730 = \P1_P1_rEIP_reg[9]/NET0131  & ~n53883 ;
  assign n55759 = \P1_P1_PhyAddrPointer_reg[9]/NET0131  & n8361 ;
  assign n55760 = ~n8357 & ~n55759 ;
  assign n55761 = ~n55730 & n55760 ;
  assign n55762 = ~n55758 & n55761 ;
  assign n55763 = ~n55739 & n55762 ;
  assign n55766 = ~\P2_P2_PhyAddrPointer_reg[0]/NET0131  & n41815 ;
  assign n55767 = n36792 & ~n55766 ;
  assign n55769 = n45060 & ~n55767 ;
  assign n55768 = ~n45060 & n55767 ;
  assign n55770 = ~\P2_P2_DataWidth_reg[1]/NET0131  & ~n55768 ;
  assign n55771 = ~n55769 & n55770 ;
  assign n55765 = \P2_P2_DataWidth_reg[1]/NET0131  & ~\P2_P2_rEIP_reg[10]/NET0131  ;
  assign n55772 = n26794 & ~n55765 ;
  assign n55773 = ~n55771 & n55772 ;
  assign n55774 = \P2_P2_rEIP_reg[10]/NET0131  & ~n50640 ;
  assign n55776 = \P2_P2_rEIP_reg[9]/NET0131  & n52099 ;
  assign n55777 = \P2_P2_rEIP_reg[10]/NET0131  & n55776 ;
  assign n55778 = ~\P2_P2_rEIP_reg[10]/NET0131  & ~n55776 ;
  assign n55779 = ~n55777 & ~n55778 ;
  assign n55780 = n50649 & ~n55779 ;
  assign n55781 = ~n26650 & n55780 ;
  assign n55775 = ~\P2_P2_EBX_reg[10]/NET0131  & ~n50642 ;
  assign n55782 = n26643 & ~n55775 ;
  assign n55783 = ~n55781 & n55782 ;
  assign n55784 = \P2_P2_EBX_reg[31]/NET0131  & ~n52121 ;
  assign n55786 = ~\P2_P2_EBX_reg[10]/NET0131  & n55784 ;
  assign n55785 = \P2_P2_EBX_reg[10]/NET0131  & ~n55784 ;
  assign n55787 = ~n50649 & ~n55785 ;
  assign n55788 = ~n55786 & n55787 ;
  assign n55789 = n26633 & ~n55780 ;
  assign n55790 = ~n55788 & n55789 ;
  assign n55791 = ~n55783 & ~n55790 ;
  assign n55792 = ~n26640 & ~n55791 ;
  assign n55793 = ~n55774 & ~n55792 ;
  assign n55794 = n26792 & ~n55793 ;
  assign n55764 = \P2_P2_rEIP_reg[10]/NET0131  & ~n54099 ;
  assign n55795 = \P2_P2_PhyAddrPointer_reg[10]/NET0131  & n27637 ;
  assign n55796 = ~n28046 & ~n55795 ;
  assign n55797 = ~n55764 & n55796 ;
  assign n55798 = ~n55794 & n55797 ;
  assign n55799 = ~n55773 & n55798 ;
  assign n55802 = n36768 & n52485 ;
  assign n55803 = n36792 & ~n55802 ;
  assign n55805 = n41819 & ~n55803 ;
  assign n55804 = ~n41819 & n55803 ;
  assign n55806 = ~\P2_P2_DataWidth_reg[1]/NET0131  & ~n55804 ;
  assign n55807 = ~n55805 & n55806 ;
  assign n55801 = \P2_P2_DataWidth_reg[1]/NET0131  & ~\P2_P2_rEIP_reg[11]/NET0131  ;
  assign n55808 = n26794 & ~n55801 ;
  assign n55809 = ~n55807 & n55808 ;
  assign n55810 = \P2_P2_rEIP_reg[11]/NET0131  & ~n50640 ;
  assign n55812 = ~\P2_P2_rEIP_reg[11]/NET0131  & ~n55777 ;
  assign n55813 = n52105 & n55776 ;
  assign n55814 = ~n55812 & ~n55813 ;
  assign n55815 = n50649 & ~n55814 ;
  assign n55816 = ~n26650 & n55815 ;
  assign n55811 = ~\P2_P2_EBX_reg[11]/NET0131  & ~n50642 ;
  assign n55817 = n26643 & ~n55811 ;
  assign n55818 = ~n55816 & n55817 ;
  assign n55819 = \P2_P2_EBX_reg[31]/NET0131  & ~n52122 ;
  assign n55821 = \P2_P2_EBX_reg[11]/NET0131  & ~n55819 ;
  assign n55820 = ~\P2_P2_EBX_reg[11]/NET0131  & n55819 ;
  assign n55822 = ~n50649 & ~n55820 ;
  assign n55823 = ~n55821 & n55822 ;
  assign n55824 = n26633 & ~n55815 ;
  assign n55825 = ~n55823 & n55824 ;
  assign n55826 = ~n55818 & ~n55825 ;
  assign n55827 = ~n26640 & ~n55826 ;
  assign n55828 = ~n55810 & ~n55827 ;
  assign n55829 = n26792 & ~n55828 ;
  assign n55800 = \P2_P2_rEIP_reg[11]/NET0131  & ~n54099 ;
  assign n55830 = \P2_P2_PhyAddrPointer_reg[11]/NET0131  & n27637 ;
  assign n55831 = ~n28046 & ~n55830 ;
  assign n55832 = ~n55800 & n55831 ;
  assign n55833 = ~n55829 & n55832 ;
  assign n55834 = ~n55809 & n55833 ;
  assign n55837 = ~\P2_P2_PhyAddrPointer_reg[0]/NET0131  & n41818 ;
  assign n55838 = n36792 & ~n55837 ;
  assign n55840 = n43758 & ~n55838 ;
  assign n55839 = ~n43758 & n55838 ;
  assign n55841 = ~\P2_P2_DataWidth_reg[1]/NET0131  & ~n55839 ;
  assign n55842 = ~n55840 & n55841 ;
  assign n55836 = \P2_P2_DataWidth_reg[1]/NET0131  & ~\P2_P2_rEIP_reg[12]/NET0131  ;
  assign n55843 = n26794 & ~n55836 ;
  assign n55844 = ~n55842 & n55843 ;
  assign n55845 = \P2_P2_rEIP_reg[12]/NET0131  & ~n50640 ;
  assign n55847 = \P2_P2_rEIP_reg[12]/NET0131  & n55813 ;
  assign n55848 = ~\P2_P2_rEIP_reg[12]/NET0131  & ~n55813 ;
  assign n55849 = ~n55847 & ~n55848 ;
  assign n55850 = n50649 & ~n55849 ;
  assign n55851 = ~n26650 & n55850 ;
  assign n55846 = ~\P2_P2_EBX_reg[12]/NET0131  & ~n50642 ;
  assign n55852 = n26643 & ~n55846 ;
  assign n55853 = ~n55851 & n55852 ;
  assign n55854 = \P2_P2_EBX_reg[31]/NET0131  & ~n52123 ;
  assign n55856 = \P2_P2_EBX_reg[12]/NET0131  & ~n55854 ;
  assign n55855 = ~\P2_P2_EBX_reg[12]/NET0131  & n55854 ;
  assign n55857 = ~n50649 & ~n55855 ;
  assign n55858 = ~n55856 & n55857 ;
  assign n55859 = n26633 & ~n55850 ;
  assign n55860 = ~n55858 & n55859 ;
  assign n55861 = ~n55853 & ~n55860 ;
  assign n55862 = ~n26640 & ~n55861 ;
  assign n55863 = ~n55845 & ~n55862 ;
  assign n55864 = n26792 & ~n55863 ;
  assign n55835 = \P2_P2_rEIP_reg[12]/NET0131  & ~n54099 ;
  assign n55865 = \P2_P2_PhyAddrPointer_reg[12]/NET0131  & n27637 ;
  assign n55866 = ~n28046 & ~n55865 ;
  assign n55867 = ~n55835 & n55866 ;
  assign n55868 = ~n55864 & n55867 ;
  assign n55869 = ~n55844 & n55868 ;
  assign n55872 = n36770 & n52152 ;
  assign n55873 = n36792 & ~n55872 ;
  assign n55875 = n43766 & ~n55873 ;
  assign n55874 = ~n43766 & n55873 ;
  assign n55876 = ~\P2_P2_DataWidth_reg[1]/NET0131  & ~n55874 ;
  assign n55877 = ~n55875 & n55876 ;
  assign n55871 = \P2_P2_DataWidth_reg[1]/NET0131  & ~\P2_P2_rEIP_reg[13]/NET0131  ;
  assign n55878 = n26794 & ~n55871 ;
  assign n55879 = ~n55877 & n55878 ;
  assign n55880 = \P2_P2_rEIP_reg[13]/NET0131  & ~n50640 ;
  assign n55882 = ~\P2_P2_rEIP_reg[13]/NET0131  & ~n55847 ;
  assign n55883 = \P2_P2_rEIP_reg[13]/NET0131  & n55847 ;
  assign n55884 = ~n55882 & ~n55883 ;
  assign n55885 = n50649 & ~n55884 ;
  assign n55886 = ~n26650 & n55885 ;
  assign n55881 = ~\P2_P2_EBX_reg[13]/NET0131  & ~n50642 ;
  assign n55887 = n26643 & ~n55881 ;
  assign n55888 = ~n55886 & n55887 ;
  assign n55889 = \P2_P2_EBX_reg[31]/NET0131  & ~n52124 ;
  assign n55891 = \P2_P2_EBX_reg[13]/NET0131  & ~n55889 ;
  assign n55890 = ~\P2_P2_EBX_reg[13]/NET0131  & n55889 ;
  assign n55892 = ~n50649 & ~n55890 ;
  assign n55893 = ~n55891 & n55892 ;
  assign n55894 = n26633 & ~n55885 ;
  assign n55895 = ~n55893 & n55894 ;
  assign n55896 = ~n55888 & ~n55895 ;
  assign n55897 = ~n26640 & ~n55896 ;
  assign n55898 = ~n55880 & ~n55897 ;
  assign n55899 = n26792 & ~n55898 ;
  assign n55870 = \P2_P2_rEIP_reg[13]/NET0131  & ~n54099 ;
  assign n55900 = \P2_P2_PhyAddrPointer_reg[13]/NET0131  & n27637 ;
  assign n55901 = ~n28046 & ~n55900 ;
  assign n55902 = ~n55870 & n55901 ;
  assign n55903 = ~n55899 & n55902 ;
  assign n55904 = ~n55879 & n55903 ;
  assign n55907 = n36792 & ~n52084 ;
  assign n55909 = n41827 & ~n55907 ;
  assign n55908 = ~n41827 & n55907 ;
  assign n55910 = ~\P2_P2_DataWidth_reg[1]/NET0131  & ~n55908 ;
  assign n55911 = ~n55909 & n55910 ;
  assign n55906 = \P2_P2_DataWidth_reg[1]/NET0131  & ~\P2_P2_rEIP_reg[14]/NET0131  ;
  assign n55912 = n26794 & ~n55906 ;
  assign n55913 = ~n55911 & n55912 ;
  assign n55914 = \P2_P2_rEIP_reg[14]/NET0131  & ~n50640 ;
  assign n55915 = \P2_P2_EBX_reg[14]/NET0131  & ~n50642 ;
  assign n55916 = ~\P2_P2_rEIP_reg[14]/NET0131  & ~n55883 ;
  assign n55917 = n50649 & ~n54111 ;
  assign n55918 = ~n55916 & n55917 ;
  assign n55919 = ~n26650 & n55918 ;
  assign n55920 = ~n55915 & ~n55919 ;
  assign n55921 = n26643 & ~n55920 ;
  assign n55922 = \P2_P2_EBX_reg[31]/NET0131  & ~n52125 ;
  assign n55924 = ~\P2_P2_EBX_reg[14]/NET0131  & ~n55922 ;
  assign n55923 = \P2_P2_EBX_reg[14]/NET0131  & n55922 ;
  assign n55925 = ~n50649 & ~n55923 ;
  assign n55926 = ~n55924 & n55925 ;
  assign n55927 = ~n55918 & ~n55926 ;
  assign n55928 = n26633 & ~n55927 ;
  assign n55929 = ~n55921 & ~n55928 ;
  assign n55930 = ~n26640 & ~n55929 ;
  assign n55931 = ~n55914 & ~n55930 ;
  assign n55932 = n26792 & ~n55931 ;
  assign n55905 = \P2_P2_rEIP_reg[14]/NET0131  & ~n54099 ;
  assign n55933 = \P2_P2_PhyAddrPointer_reg[14]/NET0131  & n27637 ;
  assign n55934 = ~n28046 & ~n55933 ;
  assign n55935 = ~n55905 & n55934 ;
  assign n55936 = ~n55932 & n55935 ;
  assign n55937 = ~n55913 & n55936 ;
  assign n55940 = ~\P2_P2_PhyAddrPointer_reg[0]/NET0131  & n39651 ;
  assign n55941 = n36792 & ~n55940 ;
  assign n55943 = n43796 & ~n55941 ;
  assign n55942 = ~n43796 & n55941 ;
  assign n55944 = ~\P2_P2_DataWidth_reg[1]/NET0131  & ~n55942 ;
  assign n55945 = ~n55943 & n55944 ;
  assign n55939 = \P2_P2_DataWidth_reg[1]/NET0131  & ~\P2_P2_rEIP_reg[16]/NET0131  ;
  assign n55946 = n26794 & ~n55939 ;
  assign n55947 = ~n55945 & n55946 ;
  assign n55948 = \P2_P2_rEIP_reg[16]/NET0131  & ~n50640 ;
  assign n55950 = ~\P2_P2_rEIP_reg[16]/NET0131  & ~n54112 ;
  assign n55951 = ~n54146 & ~n55950 ;
  assign n55952 = n50642 & ~n55951 ;
  assign n55949 = ~\P2_P2_EBX_reg[16]/NET0131  & ~n50642 ;
  assign n55953 = n26643 & ~n55949 ;
  assign n55954 = ~n55952 & n55953 ;
  assign n55956 = \P2_P2_EBX_reg[31]/NET0131  & ~n52127 ;
  assign n55958 = \P2_P2_EBX_reg[16]/NET0131  & ~n55956 ;
  assign n55957 = ~\P2_P2_EBX_reg[16]/NET0131  & n55956 ;
  assign n55959 = ~n50649 & ~n55957 ;
  assign n55960 = ~n55958 & n55959 ;
  assign n55955 = n50649 & ~n55951 ;
  assign n55961 = n26633 & ~n55955 ;
  assign n55962 = ~n55960 & n55961 ;
  assign n55963 = ~n55954 & ~n55962 ;
  assign n55964 = ~n26640 & ~n55963 ;
  assign n55965 = ~n55948 & ~n55964 ;
  assign n55966 = n26792 & ~n55965 ;
  assign n55938 = \P2_P2_rEIP_reg[16]/NET0131  & ~n54099 ;
  assign n55967 = \P2_P2_PhyAddrPointer_reg[16]/NET0131  & n27637 ;
  assign n55968 = ~n28046 & ~n55967 ;
  assign n55969 = ~n55938 & n55968 ;
  assign n55970 = ~n55966 & n55969 ;
  assign n55971 = ~n55947 & n55970 ;
  assign n55974 = n36776 & n52085 ;
  assign n55975 = n36792 & ~n55974 ;
  assign n55977 = n41861 & ~n55975 ;
  assign n55976 = ~n41861 & n55975 ;
  assign n55978 = ~\P2_P2_DataWidth_reg[1]/NET0131  & ~n55976 ;
  assign n55979 = ~n55977 & n55978 ;
  assign n55973 = \P2_P2_DataWidth_reg[1]/NET0131  & ~\P2_P2_rEIP_reg[19]/NET0131  ;
  assign n55980 = n26794 & ~n55973 ;
  assign n55981 = ~n55979 & n55980 ;
  assign n55982 = \P2_P2_rEIP_reg[19]/NET0131  & ~n50640 ;
  assign n55984 = ~\P2_P2_rEIP_reg[19]/NET0131  & ~n54183 ;
  assign n55985 = ~n52110 & ~n55984 ;
  assign n55986 = n50642 & ~n55985 ;
  assign n55983 = ~\P2_P2_EBX_reg[19]/NET0131  & ~n50642 ;
  assign n55987 = n26643 & ~n55983 ;
  assign n55988 = ~n55986 & n55987 ;
  assign n55990 = \P2_P2_EBX_reg[31]/NET0131  & ~n52130 ;
  assign n55992 = ~\P2_P2_EBX_reg[19]/NET0131  & n55990 ;
  assign n55991 = \P2_P2_EBX_reg[19]/NET0131  & ~n55990 ;
  assign n55993 = ~n50649 & ~n55991 ;
  assign n55994 = ~n55992 & n55993 ;
  assign n55989 = n50649 & ~n55985 ;
  assign n55995 = n26633 & ~n55989 ;
  assign n55996 = ~n55994 & n55995 ;
  assign n55997 = ~n55988 & ~n55996 ;
  assign n55998 = ~n26640 & ~n55997 ;
  assign n55999 = ~n55982 & ~n55998 ;
  assign n56000 = n26792 & ~n55999 ;
  assign n55972 = \P2_P2_rEIP_reg[19]/NET0131  & ~n54099 ;
  assign n56001 = \P2_P2_PhyAddrPointer_reg[19]/NET0131  & n27637 ;
  assign n56002 = ~n28046 & ~n56001 ;
  assign n56003 = ~n55972 & n56002 ;
  assign n56004 = ~n56000 & n56003 ;
  assign n56005 = ~n55981 & n56004 ;
  assign n56008 = ~\P2_P2_PhyAddrPointer_reg[0]/NET0131  & n41813 ;
  assign n56009 = n36792 & ~n56008 ;
  assign n56011 = n43884 & ~n56009 ;
  assign n56010 = ~n43884 & n56009 ;
  assign n56012 = ~\P2_P2_DataWidth_reg[1]/NET0131  & ~n56010 ;
  assign n56013 = ~n56011 & n56012 ;
  assign n56007 = \P2_P2_DataWidth_reg[1]/NET0131  & ~\P2_P2_rEIP_reg[8]/NET0131  ;
  assign n56014 = n26794 & ~n56007 ;
  assign n56015 = ~n56013 & n56014 ;
  assign n56016 = \P2_P2_rEIP_reg[8]/NET0131  & ~n50640 ;
  assign n56017 = ~\P2_P2_EBX_reg[8]/NET0131  & ~n50642 ;
  assign n56018 = ~\P2_P2_rEIP_reg[8]/NET0131  & ~n52098 ;
  assign n56019 = ~n52099 & ~n56018 ;
  assign n56020 = n50642 & ~n56019 ;
  assign n56021 = ~n56017 & ~n56020 ;
  assign n56022 = n26643 & n56021 ;
  assign n56023 = n50649 & ~n56019 ;
  assign n56024 = \P2_P2_EBX_reg[31]/NET0131  & ~n52119 ;
  assign n56026 = ~\P2_P2_EBX_reg[8]/NET0131  & n56024 ;
  assign n56025 = \P2_P2_EBX_reg[8]/NET0131  & ~n56024 ;
  assign n56027 = ~n50649 & ~n56025 ;
  assign n56028 = ~n56026 & n56027 ;
  assign n56029 = ~n56023 & ~n56028 ;
  assign n56030 = n26633 & n56029 ;
  assign n56031 = ~n56022 & ~n56030 ;
  assign n56032 = ~n26640 & ~n56031 ;
  assign n56033 = ~n56016 & ~n56032 ;
  assign n56034 = n26792 & ~n56033 ;
  assign n56006 = \P2_P2_rEIP_reg[8]/NET0131  & ~n54099 ;
  assign n56035 = \P2_P2_PhyAddrPointer_reg[8]/NET0131  & n27637 ;
  assign n56036 = ~n28046 & ~n56035 ;
  assign n56037 = ~n56006 & n56036 ;
  assign n56038 = ~n56034 & n56037 ;
  assign n56039 = ~n56015 & n56038 ;
  assign n56042 = n36766 & n52152 ;
  assign n56043 = n36792 & ~n56042 ;
  assign n56045 = n45103 & ~n56043 ;
  assign n56044 = ~n45103 & n56043 ;
  assign n56046 = ~\P2_P2_DataWidth_reg[1]/NET0131  & ~n56044 ;
  assign n56047 = ~n56045 & n56046 ;
  assign n56041 = \P2_P2_DataWidth_reg[1]/NET0131  & ~\P2_P2_rEIP_reg[9]/NET0131  ;
  assign n56048 = n26794 & ~n56041 ;
  assign n56049 = ~n56047 & n56048 ;
  assign n56050 = \P2_P2_rEIP_reg[9]/NET0131  & ~n50640 ;
  assign n56052 = ~\P2_P2_rEIP_reg[9]/NET0131  & ~n52099 ;
  assign n56053 = ~n55776 & ~n56052 ;
  assign n56054 = n50649 & ~n56053 ;
  assign n56055 = ~n26650 & n56054 ;
  assign n56051 = ~\P2_P2_EBX_reg[9]/NET0131  & ~n50642 ;
  assign n56056 = n26643 & ~n56051 ;
  assign n56057 = ~n56055 & n56056 ;
  assign n56058 = \P2_P2_EBX_reg[31]/NET0131  & ~n52120 ;
  assign n56060 = \P2_P2_EBX_reg[9]/NET0131  & ~n56058 ;
  assign n56059 = ~\P2_P2_EBX_reg[9]/NET0131  & n56058 ;
  assign n56061 = ~n50649 & ~n56059 ;
  assign n56062 = ~n56060 & n56061 ;
  assign n56063 = n26633 & ~n56054 ;
  assign n56064 = ~n56062 & n56063 ;
  assign n56065 = ~n56057 & ~n56064 ;
  assign n56066 = ~n26640 & ~n56065 ;
  assign n56067 = ~n56050 & ~n56066 ;
  assign n56068 = n26792 & ~n56067 ;
  assign n56040 = \P2_P2_rEIP_reg[9]/NET0131  & ~n54099 ;
  assign n56069 = \P2_P2_PhyAddrPointer_reg[9]/NET0131  & n27637 ;
  assign n56070 = ~n28046 & ~n56069 ;
  assign n56071 = ~n56040 & n56070 ;
  assign n56072 = ~n56068 & n56071 ;
  assign n56073 = ~n56049 & n56072 ;
  assign n56076 = \P2_P3_PhyAddrPointer_reg[0]/NET0131  & ~n36863 ;
  assign n56077 = ~n36863 & ~n39839 ;
  assign n56078 = ~n56076 & ~n56077 ;
  assign n56080 = ~n45179 & ~n56078 ;
  assign n56079 = n45179 & n56078 ;
  assign n56081 = ~\P2_P3_DataWidth_reg[1]/NET0131  & ~n56079 ;
  assign n56082 = ~n56080 & n56081 ;
  assign n56075 = \P2_P3_DataWidth_reg[1]/NET0131  & ~\P2_P3_rEIP_reg[10]/NET0131  ;
  assign n56083 = n27315 & ~n56075 ;
  assign n56084 = ~n56082 & n56083 ;
  assign n56085 = \P2_P3_rEIP_reg[10]/NET0131  & ~n27277 ;
  assign n56087 = ~\P2_P3_rEIP_reg[10]/NET0131  & ~n52554 ;
  assign n56088 = ~n52555 & ~n56087 ;
  assign n56089 = n50735 & ~n56088 ;
  assign n56086 = ~\P2_P3_EBX_reg[10]/NET0131  & ~n50735 ;
  assign n56090 = n27121 & ~n56086 ;
  assign n56091 = ~n56089 & n56090 ;
  assign n56093 = \P2_P3_EBX_reg[31]/NET0131  & ~n52530 ;
  assign n56095 = ~\P2_P3_EBX_reg[10]/NET0131  & n56093 ;
  assign n56094 = \P2_P3_EBX_reg[10]/NET0131  & ~n56093 ;
  assign n56096 = ~n27302 & ~n56094 ;
  assign n56097 = ~n56095 & n56096 ;
  assign n56092 = n27302 & ~n56088 ;
  assign n56098 = n27122 & ~n56092 ;
  assign n56099 = ~n56097 & n56098 ;
  assign n56100 = ~n56091 & ~n56099 ;
  assign n56101 = ~n27177 & ~n56100 ;
  assign n56102 = ~n56085 & ~n56101 ;
  assign n56103 = n27308 & ~n56102 ;
  assign n56074 = \P2_P3_rEIP_reg[10]/NET0131  & ~n54653 ;
  assign n56104 = \P2_P3_PhyAddrPointer_reg[10]/NET0131  & n27651 ;
  assign n56105 = ~n32864 & ~n56104 ;
  assign n56106 = ~n56074 & n56105 ;
  assign n56107 = ~n56103 & n56106 ;
  assign n56108 = ~n56084 & n56107 ;
  assign n56111 = ~n36863 & ~n39840 ;
  assign n56112 = ~n56076 & ~n56111 ;
  assign n56114 = ~n42073 & ~n56112 ;
  assign n56113 = n42073 & n56112 ;
  assign n56115 = ~\P2_P3_DataWidth_reg[1]/NET0131  & ~n56113 ;
  assign n56116 = ~n56114 & n56115 ;
  assign n56110 = \P2_P3_DataWidth_reg[1]/NET0131  & ~\P2_P3_rEIP_reg[11]/NET0131  ;
  assign n56117 = n27315 & ~n56110 ;
  assign n56118 = ~n56116 & n56117 ;
  assign n56119 = \P2_P3_rEIP_reg[11]/NET0131  & ~n27277 ;
  assign n56120 = ~\P2_P3_rEIP_reg[11]/NET0131  & ~n52555 ;
  assign n56121 = ~n52556 & ~n56120 ;
  assign n56122 = n27302 & ~n56121 ;
  assign n56123 = ~n27148 & n56122 ;
  assign n56124 = ~\P2_P3_EBX_reg[11]/NET0131  & ~n50735 ;
  assign n56125 = n27121 & ~n56124 ;
  assign n56126 = ~n56123 & n56125 ;
  assign n56127 = \P2_P3_EBX_reg[31]/NET0131  & ~n52531 ;
  assign n56129 = \P2_P3_EBX_reg[11]/NET0131  & ~n56127 ;
  assign n56128 = ~\P2_P3_EBX_reg[11]/NET0131  & n56127 ;
  assign n56130 = ~n27302 & ~n56128 ;
  assign n56131 = ~n56129 & n56130 ;
  assign n56132 = n27122 & ~n56122 ;
  assign n56133 = ~n56131 & n56132 ;
  assign n56134 = ~n56126 & ~n56133 ;
  assign n56135 = ~n27177 & ~n56134 ;
  assign n56136 = ~n56119 & ~n56135 ;
  assign n56137 = n27308 & ~n56136 ;
  assign n56109 = \P2_P3_rEIP_reg[11]/NET0131  & ~n54653 ;
  assign n56138 = \P2_P3_PhyAddrPointer_reg[11]/NET0131  & n27651 ;
  assign n56139 = ~n32864 & ~n56138 ;
  assign n56140 = ~n56109 & n56139 ;
  assign n56141 = ~n56137 & n56140 ;
  assign n56142 = ~n56118 & n56141 ;
  assign n56145 = ~n36863 & ~n39841 ;
  assign n56146 = ~n56076 & ~n56145 ;
  assign n56148 = ~n44034 & ~n56146 ;
  assign n56147 = n44034 & n56146 ;
  assign n56149 = ~\P2_P3_DataWidth_reg[1]/NET0131  & ~n56147 ;
  assign n56150 = ~n56148 & n56149 ;
  assign n56144 = \P2_P3_DataWidth_reg[1]/NET0131  & ~\P2_P3_rEIP_reg[12]/NET0131  ;
  assign n56151 = n27315 & ~n56144 ;
  assign n56152 = ~n56150 & n56151 ;
  assign n56161 = \P2_P3_EBX_reg[31]/NET0131  & ~n52532 ;
  assign n56163 = \P2_P3_EBX_reg[12]/NET0131  & ~n56161 ;
  assign n56162 = ~\P2_P3_EBX_reg[12]/NET0131  & n56161 ;
  assign n56164 = ~n27302 & ~n56162 ;
  assign n56165 = ~n56163 & n56164 ;
  assign n56155 = ~\P2_P3_rEIP_reg[12]/NET0131  & ~n52556 ;
  assign n56156 = ~n52557 & ~n56155 ;
  assign n56157 = n27302 & ~n56156 ;
  assign n56166 = n46587 & ~n56157 ;
  assign n56167 = ~n56165 & n56166 ;
  assign n56153 = \P2_P3_rEIP_reg[12]/NET0131  & ~n27277 ;
  assign n56158 = ~n27148 & n56157 ;
  assign n56154 = ~\P2_P3_EBX_reg[12]/NET0131  & ~n50735 ;
  assign n56159 = n47747 & ~n56154 ;
  assign n56160 = ~n56158 & n56159 ;
  assign n56168 = ~n56153 & ~n56160 ;
  assign n56169 = ~n56167 & n56168 ;
  assign n56170 = n27308 & ~n56169 ;
  assign n56143 = \P2_P3_rEIP_reg[12]/NET0131  & ~n54653 ;
  assign n56171 = \P2_P3_PhyAddrPointer_reg[12]/NET0131  & n27651 ;
  assign n56172 = ~n32864 & ~n56171 ;
  assign n56173 = ~n56143 & n56172 ;
  assign n56174 = ~n56170 & n56173 ;
  assign n56175 = ~n56152 & n56174 ;
  assign n56179 = n44056 & ~n54743 ;
  assign n56178 = ~n44056 & n54743 ;
  assign n56180 = ~\P2_P3_DataWidth_reg[1]/NET0131  & ~n56178 ;
  assign n56181 = ~n56179 & n56180 ;
  assign n56177 = \P2_P3_DataWidth_reg[1]/NET0131  & ~\P2_P3_rEIP_reg[13]/NET0131  ;
  assign n56182 = n27315 & ~n56177 ;
  assign n56183 = ~n56181 & n56182 ;
  assign n56184 = \P2_P3_rEIP_reg[13]/NET0131  & ~n27277 ;
  assign n56186 = ~\P2_P3_rEIP_reg[13]/NET0131  & ~n52557 ;
  assign n56187 = ~n52558 & ~n56186 ;
  assign n56188 = n27302 & ~n56187 ;
  assign n56189 = ~n27148 & n56188 ;
  assign n56185 = ~\P2_P3_EBX_reg[13]/NET0131  & ~n50735 ;
  assign n56190 = n27121 & ~n56185 ;
  assign n56191 = ~n56189 & n56190 ;
  assign n56192 = \P2_P3_EBX_reg[31]/NET0131  & ~n52533 ;
  assign n56194 = \P2_P3_EBX_reg[13]/NET0131  & ~n56192 ;
  assign n56193 = ~\P2_P3_EBX_reg[13]/NET0131  & n56192 ;
  assign n56195 = ~n27302 & ~n56193 ;
  assign n56196 = ~n56194 & n56195 ;
  assign n56197 = n27122 & ~n56188 ;
  assign n56198 = ~n56196 & n56197 ;
  assign n56199 = ~n56191 & ~n56198 ;
  assign n56200 = ~n27177 & ~n56199 ;
  assign n56201 = ~n56184 & ~n56200 ;
  assign n56202 = n27308 & ~n56201 ;
  assign n56176 = \P2_P3_rEIP_reg[13]/NET0131  & ~n54653 ;
  assign n56203 = \P2_P3_PhyAddrPointer_reg[13]/NET0131  & n27651 ;
  assign n56204 = ~n32864 & ~n56203 ;
  assign n56205 = ~n56176 & n56204 ;
  assign n56206 = ~n56202 & n56205 ;
  assign n56207 = ~n56183 & n56206 ;
  assign n56210 = \P2_P3_PhyAddrPointer_reg[13]/NET0131  & n52576 ;
  assign n56211 = ~n36863 & ~n56210 ;
  assign n56213 = n42086 & ~n56211 ;
  assign n56212 = ~n42086 & n56211 ;
  assign n56214 = ~\P2_P3_DataWidth_reg[1]/NET0131  & ~n56212 ;
  assign n56215 = ~n56213 & n56214 ;
  assign n56209 = \P2_P3_DataWidth_reg[1]/NET0131  & ~\P2_P3_rEIP_reg[14]/NET0131  ;
  assign n56216 = n27315 & ~n56209 ;
  assign n56217 = ~n56215 & n56216 ;
  assign n56218 = \P2_P3_rEIP_reg[14]/NET0131  & ~n27277 ;
  assign n56220 = ~\P2_P3_rEIP_reg[14]/NET0131  & ~n52558 ;
  assign n56221 = ~n52559 & ~n56220 ;
  assign n56222 = n50735 & ~n56221 ;
  assign n56219 = ~\P2_P3_EBX_reg[14]/NET0131  & ~n50735 ;
  assign n56223 = n27121 & ~n56219 ;
  assign n56224 = ~n56222 & n56223 ;
  assign n56226 = \P2_P3_EBX_reg[31]/NET0131  & ~n52534 ;
  assign n56227 = ~\P2_P3_EBX_reg[14]/NET0131  & ~n56226 ;
  assign n56228 = \P2_P3_EBX_reg[14]/NET0131  & n56226 ;
  assign n56229 = ~n56227 & ~n56228 ;
  assign n56230 = ~n27302 & ~n56229 ;
  assign n56225 = n27302 & ~n56221 ;
  assign n56231 = n27122 & ~n56225 ;
  assign n56232 = ~n56230 & n56231 ;
  assign n56233 = ~n56224 & ~n56232 ;
  assign n56234 = ~n27177 & ~n56233 ;
  assign n56235 = ~n56218 & ~n56234 ;
  assign n56236 = n27308 & ~n56235 ;
  assign n56208 = \P2_P3_rEIP_reg[14]/NET0131  & ~n54653 ;
  assign n56237 = \P2_P3_PhyAddrPointer_reg[14]/NET0131  & n27651 ;
  assign n56238 = ~n32864 & ~n56237 ;
  assign n56239 = ~n56208 & n56238 ;
  assign n56240 = ~n56236 & n56239 ;
  assign n56241 = ~n56217 & n56240 ;
  assign n56244 = ~\P2_P3_PhyAddrPointer_reg[15]/NET0131  & ~n36863 ;
  assign n56245 = ~n54658 & ~n56244 ;
  assign n56247 = ~n44070 & ~n56245 ;
  assign n56246 = n44070 & n56245 ;
  assign n56248 = ~\P2_P3_DataWidth_reg[1]/NET0131  & ~n56246 ;
  assign n56249 = ~n56247 & n56248 ;
  assign n56243 = \P2_P3_DataWidth_reg[1]/NET0131  & ~\P2_P3_rEIP_reg[16]/NET0131  ;
  assign n56250 = n27315 & ~n56243 ;
  assign n56251 = ~n56249 & n56250 ;
  assign n56255 = \P2_P3_EBX_reg[31]/NET0131  & ~n52536 ;
  assign n56257 = \P2_P3_EBX_reg[16]/NET0131  & ~n56255 ;
  assign n56256 = ~\P2_P3_EBX_reg[16]/NET0131  & n56255 ;
  assign n56258 = ~n27302 & ~n56256 ;
  assign n56259 = ~n56257 & n56258 ;
  assign n56252 = ~\P2_P3_rEIP_reg[16]/NET0131  & ~n52560 ;
  assign n56253 = ~n52561 & ~n56252 ;
  assign n56254 = n27302 & ~n56253 ;
  assign n56260 = n46587 & ~n56254 ;
  assign n56261 = ~n56259 & n56260 ;
  assign n56262 = \P2_P3_rEIP_reg[16]/NET0131  & ~n27277 ;
  assign n56264 = ~n27148 & n56254 ;
  assign n56263 = ~\P2_P3_EBX_reg[16]/NET0131  & ~n50735 ;
  assign n56265 = n47747 & ~n56263 ;
  assign n56266 = ~n56264 & n56265 ;
  assign n56267 = ~n56262 & ~n56266 ;
  assign n56268 = ~n56261 & n56267 ;
  assign n56269 = n27308 & ~n56268 ;
  assign n56242 = \P2_P3_rEIP_reg[16]/NET0131  & ~n54653 ;
  assign n56270 = \P2_P3_PhyAddrPointer_reg[16]/NET0131  & n27651 ;
  assign n56271 = ~n32864 & ~n56270 ;
  assign n56272 = ~n56242 & n56271 ;
  assign n56273 = ~n56269 & n56272 ;
  assign n56274 = ~n56251 & n56273 ;
  assign n56296 = ~n36863 & ~n52577 ;
  assign n56298 = n42116 & ~n56296 ;
  assign n56297 = ~n42116 & n56296 ;
  assign n56299 = ~\P2_P3_DataWidth_reg[1]/NET0131  & ~n56297 ;
  assign n56300 = ~n56298 & n56299 ;
  assign n56295 = \P2_P3_DataWidth_reg[1]/NET0131  & ~\P2_P3_rEIP_reg[19]/NET0131  ;
  assign n56301 = n27315 & ~n56295 ;
  assign n56302 = ~n56300 & n56301 ;
  assign n56276 = \P2_P3_rEIP_reg[19]/NET0131  & ~n27277 ;
  assign n56278 = ~\P2_P3_rEIP_reg[19]/NET0131  & ~n52563 ;
  assign n56279 = ~n52564 & ~n56278 ;
  assign n56280 = n50735 & ~n56279 ;
  assign n56277 = ~\P2_P3_EBX_reg[19]/NET0131  & ~n50735 ;
  assign n56281 = n27121 & ~n56277 ;
  assign n56282 = ~n56280 & n56281 ;
  assign n56284 = \P2_P3_EBX_reg[31]/NET0131  & ~n52539 ;
  assign n56286 = ~\P2_P3_EBX_reg[19]/NET0131  & n56284 ;
  assign n56285 = \P2_P3_EBX_reg[19]/NET0131  & ~n56284 ;
  assign n56287 = ~n27302 & ~n56285 ;
  assign n56288 = ~n56286 & n56287 ;
  assign n56283 = n27302 & ~n56279 ;
  assign n56289 = n27122 & ~n56283 ;
  assign n56290 = ~n56288 & n56289 ;
  assign n56291 = ~n56282 & ~n56290 ;
  assign n56292 = ~n27177 & ~n56291 ;
  assign n56293 = ~n56276 & ~n56292 ;
  assign n56294 = n27308 & ~n56293 ;
  assign n56275 = \P2_P3_rEIP_reg[19]/NET0131  & ~n54653 ;
  assign n56303 = \P2_P3_PhyAddrPointer_reg[19]/NET0131  & n27651 ;
  assign n56304 = ~n32864 & ~n56303 ;
  assign n56305 = ~n56275 & n56304 ;
  assign n56306 = ~n56294 & n56305 ;
  assign n56307 = ~n56302 & n56306 ;
  assign n56310 = \P2_P3_PhyAddrPointer_reg[7]/NET0131  & n54825 ;
  assign n56311 = ~n36863 & ~n56310 ;
  assign n56313 = ~n44159 & n56311 ;
  assign n56312 = n44159 & ~n56311 ;
  assign n56314 = ~\P2_P3_DataWidth_reg[1]/NET0131  & ~n56312 ;
  assign n56315 = ~n56313 & n56314 ;
  assign n56309 = \P2_P3_DataWidth_reg[1]/NET0131  & ~\P2_P3_rEIP_reg[8]/NET0131  ;
  assign n56316 = n27315 & ~n56309 ;
  assign n56317 = ~n56315 & n56316 ;
  assign n56318 = \P2_P3_rEIP_reg[8]/NET0131  & ~n27277 ;
  assign n56319 = ~\P2_P3_rEIP_reg[8]/NET0131  & ~n52552 ;
  assign n56320 = ~n52553 & ~n56319 ;
  assign n56321 = n27302 & ~n56320 ;
  assign n56322 = ~n27148 & n56321 ;
  assign n56323 = ~\P2_P3_EBX_reg[8]/NET0131  & ~n50735 ;
  assign n56324 = ~n56322 & ~n56323 ;
  assign n56325 = n47747 & n56324 ;
  assign n56326 = \P2_P3_EBX_reg[31]/NET0131  & ~n52528 ;
  assign n56328 = ~\P2_P3_EBX_reg[8]/NET0131  & n56326 ;
  assign n56327 = \P2_P3_EBX_reg[8]/NET0131  & ~n56326 ;
  assign n56329 = ~n27302 & ~n56327 ;
  assign n56330 = ~n56328 & n56329 ;
  assign n56331 = ~n56321 & ~n56330 ;
  assign n56332 = n46587 & n56331 ;
  assign n56333 = ~n56325 & ~n56332 ;
  assign n56334 = ~n56318 & n56333 ;
  assign n56335 = n27308 & ~n56334 ;
  assign n56308 = \P2_P3_rEIP_reg[8]/NET0131  & ~n54653 ;
  assign n56336 = \P2_P3_PhyAddrPointer_reg[8]/NET0131  & n27651 ;
  assign n56337 = ~n32864 & ~n56336 ;
  assign n56338 = ~n56308 & n56337 ;
  assign n56339 = ~n56335 & n56338 ;
  assign n56340 = ~n56317 & n56339 ;
  assign n56343 = n36840 & n50708 ;
  assign n56344 = ~n36863 & ~n56343 ;
  assign n56346 = ~n45237 & n56344 ;
  assign n56345 = n45237 & ~n56344 ;
  assign n56347 = ~\P2_P3_DataWidth_reg[1]/NET0131  & ~n56345 ;
  assign n56348 = ~n56346 & n56347 ;
  assign n56342 = \P2_P3_DataWidth_reg[1]/NET0131  & ~\P2_P3_rEIP_reg[9]/NET0131  ;
  assign n56349 = n27315 & ~n56342 ;
  assign n56350 = ~n56348 & n56349 ;
  assign n56351 = \P2_P3_rEIP_reg[9]/NET0131  & ~n27277 ;
  assign n56352 = ~\P2_P3_rEIP_reg[9]/NET0131  & ~n52553 ;
  assign n56353 = ~n52554 & ~n56352 ;
  assign n56354 = n27302 & ~n56353 ;
  assign n56355 = ~n27148 & n56354 ;
  assign n56356 = ~\P2_P3_EBX_reg[9]/NET0131  & ~n50735 ;
  assign n56357 = ~n56355 & ~n56356 ;
  assign n56358 = n47747 & n56357 ;
  assign n56359 = \P2_P3_EBX_reg[31]/NET0131  & ~n52529 ;
  assign n56361 = ~\P2_P3_EBX_reg[9]/NET0131  & n56359 ;
  assign n56360 = \P2_P3_EBX_reg[9]/NET0131  & ~n56359 ;
  assign n56362 = ~n27302 & ~n56360 ;
  assign n56363 = ~n56361 & n56362 ;
  assign n56364 = ~n56354 & ~n56363 ;
  assign n56365 = n46587 & n56364 ;
  assign n56366 = ~n56358 & ~n56365 ;
  assign n56367 = ~n56351 & n56366 ;
  assign n56368 = n27308 & ~n56367 ;
  assign n56341 = \P2_P3_rEIP_reg[9]/NET0131  & ~n54653 ;
  assign n56369 = \P2_P3_PhyAddrPointer_reg[9]/NET0131  & n27651 ;
  assign n56370 = ~n32864 & ~n56369 ;
  assign n56371 = ~n56341 & n56370 ;
  assign n56372 = ~n56368 & n56371 ;
  assign n56373 = ~n56350 & n56372 ;
  assign n56377 = \P2_P3_PhyAddrPointer_reg[1]/NET0131  & n56076 ;
  assign n56376 = ~\P2_P3_PhyAddrPointer_reg[1]/NET0131  & ~n56076 ;
  assign n56378 = ~\P2_P3_DataWidth_reg[1]/NET0131  & ~n56376 ;
  assign n56379 = ~n56377 & n56378 ;
  assign n56375 = \P2_P3_DataWidth_reg[1]/NET0131  & ~\P2_P3_rEIP_reg[1]/NET0131  ;
  assign n56380 = n27315 & ~n56375 ;
  assign n56381 = ~n56379 & n56380 ;
  assign n56383 = ~\P2_P3_EBX_reg[1]/NET0131  & ~n50735 ;
  assign n56384 = n47747 & ~n56383 ;
  assign n56386 = \P2_P3_EBX_reg[1]/NET0131  & ~\P2_P3_EBX_reg[31]/NET0131  ;
  assign n56387 = ~n46618 & n52846 ;
  assign n56388 = ~n56386 & ~n56387 ;
  assign n56389 = ~n27302 & n56388 ;
  assign n56390 = n46587 & ~n56389 ;
  assign n56391 = ~n56384 & ~n56390 ;
  assign n56392 = \P2_P3_rEIP_reg[1]/NET0131  & n27302 ;
  assign n56393 = ~n56391 & ~n56392 ;
  assign n56395 = \P2_P3_rEIP_reg[1]/NET0131  & ~n27277 ;
  assign n56385 = n27148 & n56384 ;
  assign n56394 = n27221 & n54634 ;
  assign n56396 = ~n56385 & ~n56394 ;
  assign n56397 = ~n56395 & n56396 ;
  assign n56398 = ~n56393 & n56397 ;
  assign n56399 = n27308 & ~n56398 ;
  assign n56374 = \P2_P3_PhyAddrPointer_reg[1]/NET0131  & n27651 ;
  assign n56382 = \P2_P3_rEIP_reg[1]/NET0131  & ~n50703 ;
  assign n56400 = ~n56374 & ~n56382 ;
  assign n56401 = ~n56399 & n56400 ;
  assign n56402 = ~n56381 & n56401 ;
  assign n56403 = ~n26104 & n50414 ;
  assign n56404 = \P2_P1_rEIP_reg[0]/NET0131  & ~n56403 ;
  assign n56405 = ~\P2_P1_InstQueueRd_Addr_reg[0]/NET0131  & n21067 ;
  assign n56406 = \P2_P1_EBX_reg[0]/NET0131  & ~n26103 ;
  assign n56407 = n24898 & n56406 ;
  assign n56408 = ~n56405 & ~n56407 ;
  assign n56409 = ~n21081 & ~n56408 ;
  assign n56410 = \P2_P1_rEIP_reg[0]/NET0131  & n50422 ;
  assign n56411 = \P2_P1_EBX_reg[0]/NET0131  & ~n50422 ;
  assign n56412 = ~n21081 & n56411 ;
  assign n56413 = ~n56410 & ~n56412 ;
  assign n56414 = n21062 & ~n56413 ;
  assign n56415 = ~n56409 & ~n56414 ;
  assign n56416 = ~n56404 & n56415 ;
  assign n56417 = n11623 & ~n56416 ;
  assign n56418 = ~n11625 & ~n26108 ;
  assign n56419 = \P2_P1_PhyAddrPointer_reg[0]/NET0131  & ~n56418 ;
  assign n56420 = ~n27681 & n50411 ;
  assign n56421 = \P2_P1_rEIP_reg[0]/NET0131  & ~n56420 ;
  assign n56422 = ~n56419 & ~n56421 ;
  assign n56423 = ~n56417 & n56422 ;
  assign n56433 = n25769 & n25914 ;
  assign n56434 = n48371 & ~n56433 ;
  assign n56435 = \P1_P2_rEIP_reg[0]/NET0131  & ~n56434 ;
  assign n56428 = ~\P1_P2_InstQueueRd_Addr_reg[0]/NET0131  & n25761 ;
  assign n56429 = \P1_P2_EBX_reg[0]/NET0131  & ~n48443 ;
  assign n56430 = n25757 & n56429 ;
  assign n56431 = ~n56428 & ~n56430 ;
  assign n56432 = ~n25770 & ~n56431 ;
  assign n56436 = \P1_P2_rEIP_reg[0]/NET0131  & n48373 ;
  assign n56437 = \P1_P2_EBX_reg[0]/NET0131  & ~n48373 ;
  assign n56438 = ~n25770 & n56437 ;
  assign n56439 = ~n56436 & ~n56438 ;
  assign n56440 = n25776 & ~n56439 ;
  assign n56441 = ~n56432 & ~n56440 ;
  assign n56442 = ~n56435 & n56441 ;
  assign n56443 = n25918 & ~n56442 ;
  assign n56424 = ~n25929 & ~n27675 ;
  assign n56425 = \P1_P2_PhyAddrPointer_reg[0]/NET0131  & ~n56424 ;
  assign n56426 = ~n25933 & n48452 ;
  assign n56427 = \P1_P2_rEIP_reg[0]/NET0131  & ~n56426 ;
  assign n56444 = ~n56425 & ~n56427 ;
  assign n56445 = ~n56443 & n56444 ;
  assign n56452 = ~\P2_P1_EBX_reg[29]/NET0131  & n51117 ;
  assign n56453 = \P2_P1_EBX_reg[31]/NET0131  & ~n56452 ;
  assign n56455 = ~\P2_P1_EBX_reg[30]/NET0131  & n56453 ;
  assign n56454 = \P2_P1_EBX_reg[30]/NET0131  & ~n56453 ;
  assign n56456 = ~n50422 & ~n56454 ;
  assign n56457 = ~n56455 & n56456 ;
  assign n56448 = ~\P2_P1_rEIP_reg[30]/NET0131  & ~n51114 ;
  assign n56449 = \P2_P1_rEIP_reg[30]/NET0131  & n51114 ;
  assign n56450 = ~n56448 & ~n56449 ;
  assign n56451 = n50422 & ~n56450 ;
  assign n56458 = n24901 & ~n56451 ;
  assign n56459 = ~n56457 & n56458 ;
  assign n56447 = \P2_P1_rEIP_reg[30]/NET0131  & ~n50414 ;
  assign n56461 = n26103 & ~n56450 ;
  assign n56460 = ~\P2_P1_EBX_reg[30]/NET0131  & ~n26103 ;
  assign n56462 = n24899 & ~n56460 ;
  assign n56463 = ~n56461 & n56462 ;
  assign n56464 = ~n56447 & ~n56463 ;
  assign n56465 = ~n56459 & n56464 ;
  assign n56466 = n11623 & ~n56465 ;
  assign n56469 = ~n39540 & n51134 ;
  assign n56470 = n36672 & ~n56469 ;
  assign n56472 = n37942 & ~n56470 ;
  assign n56471 = ~n37942 & n56470 ;
  assign n56473 = ~\P2_P1_DataWidth_reg[1]/NET0131  & ~n56471 ;
  assign n56474 = ~n56472 & n56473 ;
  assign n56468 = \P2_P1_DataWidth_reg[1]/NET0131  & ~\P2_P1_rEIP_reg[30]/NET0131  ;
  assign n56475 = n11609 & ~n56468 ;
  assign n56476 = ~n56474 & n56475 ;
  assign n56446 = \P2_P1_PhyAddrPointer_reg[30]/NET0131  & n11625 ;
  assign n56467 = \P2_P1_rEIP_reg[30]/NET0131  & ~n50411 ;
  assign n56477 = ~n56446 & ~n56467 ;
  assign n56478 = ~n56476 & n56477 ;
  assign n56479 = ~n56466 & n56478 ;
  assign n56482 = ~\P2_P1_rEIP_reg[31]/NET0131  & ~n56449 ;
  assign n56483 = \P2_P1_rEIP_reg[31]/NET0131  & n56449 ;
  assign n56484 = ~n56482 & ~n56483 ;
  assign n56485 = n50422 & n56484 ;
  assign n56486 = ~\P2_P1_EBX_reg[30]/NET0131  & \P2_P1_EBX_reg[31]/NET0131  ;
  assign n56487 = ~n50422 & n56486 ;
  assign n56488 = n56452 & n56487 ;
  assign n56489 = ~n56485 & ~n56488 ;
  assign n56490 = n24901 & ~n56489 ;
  assign n56481 = \P2_P1_rEIP_reg[31]/NET0131  & ~n50414 ;
  assign n56492 = n26103 & ~n56484 ;
  assign n56491 = ~\P2_P1_EBX_reg[31]/NET0131  & ~n26103 ;
  assign n56493 = n24899 & ~n56491 ;
  assign n56494 = ~n56492 & n56493 ;
  assign n56495 = ~n56481 & ~n56494 ;
  assign n56496 = ~n56490 & n56495 ;
  assign n56497 = n11623 & ~n56496 ;
  assign n56498 = \P2_P1_DataWidth_reg[1]/NET0131  & \P2_P1_rEIP_reg[31]/NET0131  ;
  assign n56499 = ~\P2_P1_DataWidth_reg[1]/NET0131  & ~n37942 ;
  assign n56500 = n56469 & n56499 ;
  assign n56501 = n36672 & n56500 ;
  assign n56502 = ~n56498 & ~n56501 ;
  assign n56503 = n11609 & ~n56502 ;
  assign n56480 = \P2_P1_PhyAddrPointer_reg[31]/NET0131  & n11625 ;
  assign n56504 = \P2_P1_rEIP_reg[31]/NET0131  & ~n50411 ;
  assign n56505 = ~n56480 & ~n56504 ;
  assign n56506 = ~n56503 & n56505 ;
  assign n56507 = ~n56497 & n56506 ;
  assign n56512 = \P1_P1_rEIP_reg[0]/NET0131  & ~n50559 ;
  assign n56518 = ~\P1_P1_EBX_reg[0]/NET0131  & n26158 ;
  assign n56514 = \P1_P1_EBX_reg[0]/NET0131  & ~n26274 ;
  assign n56515 = \P1_P1_rEIP_reg[0]/NET0131  & n26274 ;
  assign n56516 = ~n56514 & ~n56515 ;
  assign n56519 = ~n26158 & n56516 ;
  assign n56520 = ~n56518 & ~n56519 ;
  assign n56521 = n24502 & n56520 ;
  assign n56513 = ~\P1_P1_InstQueueRd_Addr_reg[0]/NET0131  & n15382 ;
  assign n56517 = n15334 & ~n56516 ;
  assign n56522 = ~n56513 & ~n56517 ;
  assign n56523 = ~n56521 & n56522 ;
  assign n56524 = ~n15364 & ~n56523 ;
  assign n56525 = ~n56512 & ~n56524 ;
  assign n56526 = n8355 & ~n56525 ;
  assign n56508 = ~n8361 & ~n26280 ;
  assign n56509 = \P1_P1_PhyAddrPointer_reg[0]/NET0131  & ~n56508 ;
  assign n56510 = ~n27791 & n50583 ;
  assign n56511 = \P1_P1_rEIP_reg[0]/NET0131  & ~n56510 ;
  assign n56527 = ~n56509 & ~n56511 ;
  assign n56528 = ~n56526 & n56527 ;
  assign n56531 = \P1_P1_PhyAddrPointer_reg[31]/NET0131  & ~n36729 ;
  assign n56532 = ~n51894 & ~n56531 ;
  assign n56534 = n37960 & n56532 ;
  assign n56533 = ~n37960 & ~n56532 ;
  assign n56535 = ~\P1_P1_DataWidth_reg[1]/NET0131  & ~n56533 ;
  assign n56536 = ~n56534 & n56535 ;
  assign n56530 = \P1_P1_DataWidth_reg[1]/NET0131  & ~\P1_P1_rEIP_reg[30]/NET0131  ;
  assign n56537 = n8282 & ~n56530 ;
  assign n56538 = ~n56536 & n56537 ;
  assign n56548 = ~\P1_P1_EBX_reg[29]/NET0131  & n52025 ;
  assign n56549 = \P1_P1_EBX_reg[31]/NET0131  & ~n56548 ;
  assign n56551 = ~\P1_P1_EBX_reg[30]/NET0131  & n56549 ;
  assign n56550 = \P1_P1_EBX_reg[30]/NET0131  & ~n56549 ;
  assign n56552 = ~n26274 & ~n56550 ;
  assign n56553 = ~n56551 & n56552 ;
  assign n56541 = \P1_P1_rEIP_reg[30]/NET0131  & n52022 ;
  assign n56542 = ~\P1_P1_rEIP_reg[30]/NET0131  & ~n52022 ;
  assign n56543 = ~n56541 & ~n56542 ;
  assign n56544 = n26274 & ~n56543 ;
  assign n56554 = n24504 & ~n56544 ;
  assign n56555 = ~n56553 & n56554 ;
  assign n56539 = \P1_P1_rEIP_reg[30]/NET0131  & ~n50559 ;
  assign n56545 = ~n26158 & n56544 ;
  assign n56540 = ~\P1_P1_EBX_reg[30]/NET0131  & ~n26275 ;
  assign n56546 = n24503 & ~n56540 ;
  assign n56547 = ~n56545 & n56546 ;
  assign n56556 = ~n56539 & ~n56547 ;
  assign n56557 = ~n56555 & n56556 ;
  assign n56558 = n8355 & ~n56557 ;
  assign n56529 = \P1_P1_PhyAddrPointer_reg[30]/NET0131  & n8361 ;
  assign n56559 = \P1_P1_rEIP_reg[30]/NET0131  & ~n50583 ;
  assign n56560 = ~n56529 & ~n56559 ;
  assign n56561 = ~n56558 & n56560 ;
  assign n56562 = ~n56538 & n56561 ;
  assign n56565 = \P1_P1_rEIP_reg[31]/NET0131  & ~n56541 ;
  assign n56566 = ~\P1_P1_rEIP_reg[31]/NET0131  & n56541 ;
  assign n56567 = ~n56565 & ~n56566 ;
  assign n56568 = n26275 & n56567 ;
  assign n56564 = ~\P1_P1_EBX_reg[31]/NET0131  & ~n26275 ;
  assign n56569 = n24502 & ~n56564 ;
  assign n56570 = ~n56568 & n56569 ;
  assign n56571 = n50559 & ~n56570 ;
  assign n56572 = \P1_P1_rEIP_reg[31]/NET0131  & ~n56571 ;
  assign n56573 = n26274 & ~n56567 ;
  assign n56574 = ~\P1_P1_EBX_reg[30]/NET0131  & \P1_P1_EBX_reg[31]/NET0131  ;
  assign n56575 = ~n26274 & n56574 ;
  assign n56576 = n56548 & n56575 ;
  assign n56577 = ~n56573 & ~n56576 ;
  assign n56578 = n15334 & ~n56577 ;
  assign n56579 = ~n56570 & ~n56578 ;
  assign n56580 = ~n15364 & ~n56579 ;
  assign n56581 = ~n56572 & ~n56580 ;
  assign n56582 = n8355 & ~n56581 ;
  assign n56583 = \P1_P1_DataWidth_reg[1]/NET0131  & \P1_P1_rEIP_reg[31]/NET0131  ;
  assign n56584 = ~\P1_P1_DataWidth_reg[1]/NET0131  & n51893 ;
  assign n56585 = n36732 & n56584 ;
  assign n56586 = ~n56583 & ~n56585 ;
  assign n56587 = n8282 & ~n56586 ;
  assign n56563 = \P1_P1_PhyAddrPointer_reg[31]/NET0131  & n8361 ;
  assign n56588 = \P1_P1_rEIP_reg[31]/NET0131  & ~n50583 ;
  assign n56589 = ~n56563 & ~n56588 ;
  assign n56590 = ~n56587 & n56589 ;
  assign n56591 = ~n56582 & n56590 ;
  assign n56596 = ~n26788 & n50640 ;
  assign n56597 = \P2_P2_rEIP_reg[0]/NET0131  & ~n56596 ;
  assign n56599 = ~\P2_P2_EBX_reg[0]/NET0131  & ~n50649 ;
  assign n56600 = ~\P2_P2_rEIP_reg[0]/NET0131  & n50649 ;
  assign n56601 = ~n56599 & ~n56600 ;
  assign n56602 = n47684 & n56601 ;
  assign n56598 = ~\P2_P2_InstQueueRd_Addr_reg[0]/NET0131  & n50638 ;
  assign n56603 = \P2_P2_EBX_reg[0]/NET0131  & ~n50642 ;
  assign n56604 = n26786 & n56603 ;
  assign n56605 = ~n56598 & ~n56604 ;
  assign n56606 = ~n56602 & n56605 ;
  assign n56607 = ~n56597 & n56606 ;
  assign n56608 = n26792 & ~n56607 ;
  assign n56592 = ~n26795 & ~n27637 ;
  assign n56593 = \P2_P2_PhyAddrPointer_reg[0]/NET0131  & ~n56592 ;
  assign n56594 = ~n26800 & n50636 ;
  assign n56595 = \P2_P2_rEIP_reg[0]/NET0131  & ~n56594 ;
  assign n56609 = ~n56593 & ~n56595 ;
  assign n56610 = ~n56608 & n56609 ;
  assign n56621 = ~\P2_P2_EBX_reg[29]/NET0131  & n52456 ;
  assign n56622 = \P2_P2_EBX_reg[31]/NET0131  & ~n56621 ;
  assign n56624 = ~\P2_P2_EBX_reg[30]/NET0131  & n56622 ;
  assign n56623 = \P2_P2_EBX_reg[30]/NET0131  & ~n56622 ;
  assign n56625 = ~n50649 & ~n56623 ;
  assign n56626 = ~n56624 & n56625 ;
  assign n56614 = \P2_P2_rEIP_reg[30]/NET0131  & n52446 ;
  assign n56615 = ~\P2_P2_rEIP_reg[30]/NET0131  & ~n52446 ;
  assign n56616 = ~n56614 & ~n56615 ;
  assign n56617 = n50649 & ~n56616 ;
  assign n56627 = n47684 & ~n56617 ;
  assign n56628 = ~n56626 & n56627 ;
  assign n56612 = \P2_P2_rEIP_reg[30]/NET0131  & ~n50640 ;
  assign n56618 = ~n26650 & n56617 ;
  assign n56613 = ~\P2_P2_EBX_reg[30]/NET0131  & ~n50642 ;
  assign n56619 = n26786 & ~n56613 ;
  assign n56620 = ~n56618 & n56619 ;
  assign n56629 = ~n56612 & ~n56620 ;
  assign n56630 = ~n56628 & n56629 ;
  assign n56631 = n26792 & ~n56630 ;
  assign n56635 = ~n39742 & n52333 ;
  assign n56636 = n52470 & n56635 ;
  assign n56638 = \P2_P2_PhyAddrPointer_reg[31]/NET0131  & ~n56636 ;
  assign n56639 = n37977 & ~n56638 ;
  assign n56634 = n36792 & ~n37977 ;
  assign n56637 = n56634 & ~n56636 ;
  assign n56640 = ~\P2_P2_DataWidth_reg[1]/NET0131  & ~n56637 ;
  assign n56641 = ~n56639 & n56640 ;
  assign n56633 = \P2_P2_DataWidth_reg[1]/NET0131  & ~\P2_P2_rEIP_reg[30]/NET0131  ;
  assign n56642 = n26794 & ~n56633 ;
  assign n56643 = ~n56641 & n56642 ;
  assign n56611 = \P2_P2_PhyAddrPointer_reg[30]/NET0131  & n27637 ;
  assign n56632 = \P2_P2_rEIP_reg[30]/NET0131  & ~n50636 ;
  assign n56644 = ~n56611 & ~n56632 ;
  assign n56645 = ~n56643 & n56644 ;
  assign n56646 = ~n56631 & n56645 ;
  assign n56648 = \P2_P2_DataWidth_reg[1]/NET0131  & \P2_P2_rEIP_reg[31]/NET0131  ;
  assign n56649 = ~\P2_P2_DataWidth_reg[1]/NET0131  & n56634 ;
  assign n56650 = n56636 & n56649 ;
  assign n56651 = ~n56648 & ~n56650 ;
  assign n56652 = n26794 & ~n56651 ;
  assign n56654 = ~\P2_P2_rEIP_reg[31]/NET0131  & ~n56614 ;
  assign n56655 = \P2_P2_rEIP_reg[31]/NET0131  & n56614 ;
  assign n56656 = ~n56654 & ~n56655 ;
  assign n56657 = n50649 & n56656 ;
  assign n56658 = ~\P2_P2_EBX_reg[30]/NET0131  & \P2_P2_EBX_reg[31]/NET0131  ;
  assign n56659 = ~n50649 & n56658 ;
  assign n56660 = n56621 & n56659 ;
  assign n56661 = ~n56657 & ~n56660 ;
  assign n56662 = n47684 & ~n56661 ;
  assign n56653 = \P2_P2_rEIP_reg[31]/NET0131  & ~n50640 ;
  assign n56664 = n50642 & ~n56656 ;
  assign n56663 = ~\P2_P2_EBX_reg[31]/NET0131  & ~n50642 ;
  assign n56665 = n26786 & ~n56663 ;
  assign n56666 = ~n56664 & n56665 ;
  assign n56667 = ~n56653 & ~n56666 ;
  assign n56668 = ~n56662 & n56667 ;
  assign n56669 = n26792 & ~n56668 ;
  assign n56647 = \P2_P2_PhyAddrPointer_reg[31]/NET0131  & n27637 ;
  assign n56670 = \P2_P2_rEIP_reg[31]/NET0131  & ~n50636 ;
  assign n56671 = ~n56647 & ~n56670 ;
  assign n56672 = ~n56669 & n56671 ;
  assign n56673 = ~n56652 & n56672 ;
  assign n56675 = ~n27303 & ~n46587 ;
  assign n56676 = n27302 & ~n56675 ;
  assign n56677 = n27277 & ~n56676 ;
  assign n56678 = \P2_P3_rEIP_reg[0]/NET0131  & ~n56677 ;
  assign n56674 = ~\P2_P3_InstQueueRd_Addr_reg[0]/NET0131  & n54634 ;
  assign n56679 = ~n27302 & n46587 ;
  assign n56680 = n47747 & ~n50735 ;
  assign n56681 = ~n56679 & ~n56680 ;
  assign n56682 = \P2_P3_EBX_reg[0]/NET0131  & ~n56681 ;
  assign n56683 = ~n56674 & ~n56682 ;
  assign n56684 = ~n56678 & n56683 ;
  assign n56685 = n27308 & ~n56684 ;
  assign n56686 = ~n27316 & ~n27651 ;
  assign n56687 = \P2_P3_PhyAddrPointer_reg[0]/NET0131  & ~n56686 ;
  assign n56688 = ~n27325 & n50703 ;
  assign n56689 = \P2_P3_rEIP_reg[0]/NET0131  & ~n56688 ;
  assign n56690 = ~n56687 & ~n56689 ;
  assign n56691 = ~n56685 & n56690 ;
  assign n56703 = \P2_P3_rEIP_reg[25]/NET0131  & ~n27277 ;
  assign n56704 = ~\P2_P3_EBX_reg[25]/NET0131  & ~n50735 ;
  assign n56705 = n47747 & ~n56704 ;
  assign n56706 = \P2_P3_EBX_reg[31]/NET0131  & ~n52729 ;
  assign n56708 = ~\P2_P3_EBX_reg[25]/NET0131  & n56706 ;
  assign n56707 = \P2_P3_EBX_reg[25]/NET0131  & ~n56706 ;
  assign n56709 = ~n27302 & ~n56707 ;
  assign n56710 = ~n56708 & n56709 ;
  assign n56711 = n46587 & ~n56710 ;
  assign n56712 = ~n56705 & ~n56711 ;
  assign n56713 = ~\P2_P3_rEIP_reg[25]/NET0131  & ~n52697 ;
  assign n56714 = ~n52736 & ~n56713 ;
  assign n56715 = n27148 & n56705 ;
  assign n56716 = n27302 & ~n56715 ;
  assign n56717 = ~n56714 & n56716 ;
  assign n56718 = ~n56712 & ~n56717 ;
  assign n56719 = ~n56703 & ~n56718 ;
  assign n56720 = n27308 & ~n56719 ;
  assign n56694 = ~n36853 & ~n36863 ;
  assign n56695 = ~n52648 & ~n56694 ;
  assign n56697 = ~n44150 & ~n56695 ;
  assign n56696 = n44150 & n56695 ;
  assign n56698 = ~\P2_P3_DataWidth_reg[1]/NET0131  & ~n56696 ;
  assign n56699 = ~n56697 & n56698 ;
  assign n56693 = \P2_P3_DataWidth_reg[1]/NET0131  & ~\P2_P3_rEIP_reg[25]/NET0131  ;
  assign n56700 = n27315 & ~n56693 ;
  assign n56701 = ~n56699 & n56700 ;
  assign n56692 = \P2_P3_PhyAddrPointer_reg[25]/NET0131  & n27651 ;
  assign n56702 = \P2_P3_rEIP_reg[25]/NET0131  & ~n50703 ;
  assign n56721 = ~n56692 & ~n56702 ;
  assign n56722 = ~n56701 & n56721 ;
  assign n56723 = ~n56720 & n56722 ;
  assign n56741 = ~\P2_P3_EBX_reg[28]/NET0131  & n52803 ;
  assign n56742 = \P2_P3_EBX_reg[31]/NET0131  & ~n56741 ;
  assign n56744 = ~\P2_P3_EBX_reg[29]/NET0131  & n56742 ;
  assign n56743 = \P2_P3_EBX_reg[29]/NET0131  & ~n56742 ;
  assign n56745 = ~n27302 & ~n56743 ;
  assign n56746 = ~n56744 & n56745 ;
  assign n56727 = ~\P2_P3_rEIP_reg[29]/NET0131  & ~n52800 ;
  assign n56728 = \P2_P3_rEIP_reg[29]/NET0131  & n52800 ;
  assign n56729 = ~n56727 & ~n56728 ;
  assign n56730 = n27302 & ~n56729 ;
  assign n56747 = n46587 & ~n56730 ;
  assign n56748 = ~n56746 & n56747 ;
  assign n56726 = ~\P2_P3_EBX_reg[29]/NET0131  & ~n27302 ;
  assign n56731 = n27178 & ~n56726 ;
  assign n56732 = ~n56730 & n56731 ;
  assign n56725 = \P2_P3_rEIP_reg[29]/NET0131  & n27177 ;
  assign n56733 = \P2_P3_EBX_reg[29]/NET0131  & n27148 ;
  assign n56734 = ~n27177 & n56733 ;
  assign n56735 = ~n56725 & ~n56734 ;
  assign n56736 = ~n56732 & n56735 ;
  assign n56737 = n27121 & ~n56736 ;
  assign n56738 = n27121 & ~n27124 ;
  assign n56739 = \P2_P3_rEIP_reg[29]/NET0131  & ~n56738 ;
  assign n56740 = ~n27277 & n56739 ;
  assign n56749 = ~n56737 & ~n56740 ;
  assign n56750 = ~n56748 & n56749 ;
  assign n56751 = n27308 & ~n56750 ;
  assign n56754 = ~n39910 & n52821 ;
  assign n56755 = ~n36863 & ~n56754 ;
  assign n56757 = n39928 & ~n56755 ;
  assign n56756 = ~n39928 & n56755 ;
  assign n56758 = ~\P2_P3_DataWidth_reg[1]/NET0131  & ~n56756 ;
  assign n56759 = ~n56757 & n56758 ;
  assign n56753 = \P2_P3_DataWidth_reg[1]/NET0131  & ~\P2_P3_rEIP_reg[29]/NET0131  ;
  assign n56760 = n27315 & ~n56753 ;
  assign n56761 = ~n56759 & n56760 ;
  assign n56724 = \P2_P3_PhyAddrPointer_reg[29]/NET0131  & n27651 ;
  assign n56752 = \P2_P3_rEIP_reg[29]/NET0131  & ~n50703 ;
  assign n56762 = ~n56724 & ~n56752 ;
  assign n56763 = ~n56761 & n56762 ;
  assign n56764 = ~n56751 & n56763 ;
  assign n56775 = ~\P2_P3_EBX_reg[29]/NET0131  & n56741 ;
  assign n56776 = \P2_P3_EBX_reg[31]/NET0131  & ~n56775 ;
  assign n56777 = ~\P2_P3_EBX_reg[30]/NET0131  & ~n56776 ;
  assign n56778 = \P2_P3_EBX_reg[30]/NET0131  & n56776 ;
  assign n56779 = ~n56777 & ~n56778 ;
  assign n56780 = ~n27302 & ~n56779 ;
  assign n56768 = \P2_P3_rEIP_reg[30]/NET0131  & n56728 ;
  assign n56769 = ~\P2_P3_rEIP_reg[30]/NET0131  & ~n56728 ;
  assign n56770 = ~n56768 & ~n56769 ;
  assign n56774 = n27302 & ~n56770 ;
  assign n56781 = n46587 & ~n56774 ;
  assign n56782 = ~n56780 & n56781 ;
  assign n56766 = \P2_P3_rEIP_reg[30]/NET0131  & ~n27277 ;
  assign n56771 = n50735 & ~n56770 ;
  assign n56767 = ~\P2_P3_EBX_reg[30]/NET0131  & ~n50735 ;
  assign n56772 = n47747 & ~n56767 ;
  assign n56773 = ~n56771 & n56772 ;
  assign n56783 = ~n56766 & ~n56773 ;
  assign n56784 = ~n56782 & n56783 ;
  assign n56785 = n27308 & ~n56784 ;
  assign n56788 = ~n39928 & n56754 ;
  assign n56789 = ~n36863 & ~n56788 ;
  assign n56791 = n38018 & ~n56789 ;
  assign n56790 = ~n38018 & n56789 ;
  assign n56792 = ~\P2_P3_DataWidth_reg[1]/NET0131  & ~n56790 ;
  assign n56793 = ~n56791 & n56792 ;
  assign n56787 = \P2_P3_DataWidth_reg[1]/NET0131  & ~\P2_P3_rEIP_reg[30]/NET0131  ;
  assign n56794 = n27315 & ~n56787 ;
  assign n56795 = ~n56793 & n56794 ;
  assign n56765 = \P2_P3_PhyAddrPointer_reg[30]/NET0131  & n27651 ;
  assign n56786 = \P2_P3_rEIP_reg[30]/NET0131  & ~n50703 ;
  assign n56796 = ~n56765 & ~n56786 ;
  assign n56797 = ~n56795 & n56796 ;
  assign n56798 = ~n56785 & n56797 ;
  assign n56804 = n56676 & ~n56768 ;
  assign n56805 = n27277 & ~n56804 ;
  assign n56806 = \P2_P3_rEIP_reg[31]/NET0131  & ~n56805 ;
  assign n56800 = ~\P2_P3_EBX_reg[30]/NET0131  & n56679 ;
  assign n56801 = n56775 & n56800 ;
  assign n56802 = ~n56680 & ~n56801 ;
  assign n56803 = \P2_P3_EBX_reg[31]/NET0131  & ~n56802 ;
  assign n56807 = ~\P2_P3_rEIP_reg[31]/NET0131  & n56676 ;
  assign n56808 = n56768 & n56807 ;
  assign n56809 = ~n56803 & ~n56808 ;
  assign n56810 = ~n56806 & n56809 ;
  assign n56811 = n27308 & ~n56810 ;
  assign n56812 = \P2_P3_DataWidth_reg[1]/NET0131  & \P2_P3_rEIP_reg[31]/NET0131  ;
  assign n56813 = ~\P2_P3_DataWidth_reg[1]/NET0131  & ~n38018 ;
  assign n56814 = n56788 & n56813 ;
  assign n56815 = ~n36863 & n56814 ;
  assign n56816 = ~n56812 & ~n56815 ;
  assign n56817 = n27315 & ~n56816 ;
  assign n56799 = \P2_P3_PhyAddrPointer_reg[31]/NET0131  & n27651 ;
  assign n56818 = \P2_P3_rEIP_reg[31]/NET0131  & ~n50703 ;
  assign n56819 = ~n56799 & ~n56818 ;
  assign n56820 = ~n56817 & n56819 ;
  assign n56821 = ~n56811 & n56820 ;
  assign n56823 = ~n26158 & n28731 ;
  assign n56824 = \P1_P1_Datao_reg[27]/NET0131  & ~n26162 ;
  assign n56825 = ~n56823 & ~n56824 ;
  assign n56826 = n8355 & ~n56825 ;
  assign n56822 = \P1_P1_uWord_reg[11]/NET0131  & n27790 ;
  assign n56827 = \P1_P1_Datao_reg[27]/NET0131  & ~n48479 ;
  assign n56828 = ~n56822 & ~n56827 ;
  assign n56829 = ~n56826 & n56828 ;
  assign n56831 = \P2_P2_Datao_reg[27]/NET0131  & ~n26699 ;
  assign n56832 = ~\P2_P2_EAX_reg[27]/NET0131  & ~n47670 ;
  assign n56833 = n26786 & ~n47671 ;
  assign n56834 = ~n56832 & n56833 ;
  assign n56835 = ~n26650 & n56834 ;
  assign n56836 = ~n56831 & ~n56835 ;
  assign n56837 = n26792 & ~n56836 ;
  assign n56830 = \P2_P2_uWord_reg[11]/NET0131  & n48491 ;
  assign n56838 = \P2_P2_Datao_reg[27]/NET0131  & ~n48508 ;
  assign n56839 = ~n56830 & ~n56838 ;
  assign n56840 = ~n56837 & n56839 ;
  assign n56849 = ~n27223 & n27308 ;
  assign n56850 = n48540 & ~n56849 ;
  assign n56851 = \P2_P3_Datao_reg[27]/NET0131  & ~n56850 ;
  assign n56841 = ~n27148 & n27308 ;
  assign n56842 = \P2_P3_EAX_reg[25]/NET0131  & n48531 ;
  assign n56843 = \P2_P3_EAX_reg[26]/NET0131  & n56842 ;
  assign n56845 = \P2_P3_EAX_reg[27]/NET0131  & n56843 ;
  assign n56844 = ~\P2_P3_EAX_reg[27]/NET0131  & ~n56843 ;
  assign n56846 = n47747 & ~n56844 ;
  assign n56847 = ~n56845 & n56846 ;
  assign n56848 = n56841 & n56847 ;
  assign n56852 = \P2_P3_uWord_reg[11]/NET0131  & n48523 ;
  assign n56853 = ~n56848 & ~n56852 ;
  assign n56854 = ~n56851 & n56853 ;
  assign n56856 = ~\P1_P2_EAX_reg[27]/NET0131  & ~n47557 ;
  assign n56857 = ~n47558 & ~n56856 ;
  assign n56858 = ~n25768 & ~n56857 ;
  assign n56859 = n47570 & ~n56858 ;
  assign n56860 = n48554 & ~n56859 ;
  assign n56861 = \P1_P2_Datao_reg[27]/NET0131  & ~n56860 ;
  assign n56862 = n47570 & n56857 ;
  assign n56863 = ~n25768 & n56862 ;
  assign n56864 = ~n56861 & ~n56863 ;
  assign n56865 = n25918 & ~n56864 ;
  assign n56855 = \P1_P2_uWord_reg[11]/NET0131  & n25922 ;
  assign n56866 = \P1_P2_Datao_reg[27]/NET0131  & ~n48566 ;
  assign n56867 = ~n56855 & ~n56866 ;
  assign n56868 = ~n56865 & n56867 ;
  assign n56870 = ~n25958 & ~n29514 ;
  assign n56871 = n24899 & ~n56870 ;
  assign n56872 = n48584 & ~n56871 ;
  assign n56873 = \P2_P1_Datao_reg[27]/NET0131  & ~n56872 ;
  assign n56874 = n26006 & n29515 ;
  assign n56875 = ~n56873 & ~n56874 ;
  assign n56876 = n11623 & ~n56875 ;
  assign n56869 = \P2_P1_uWord_reg[11]/NET0131  & n48581 ;
  assign n56877 = \P2_P1_Datao_reg[27]/NET0131  & ~n48594 ;
  assign n56878 = ~n56869 & ~n56877 ;
  assign n56879 = ~n56876 & n56878 ;
  assign n56882 = ~\P2_P1_EBX_reg[25]/NET0131  & ~n46253 ;
  assign n56883 = n25981 & ~n46254 ;
  assign n56884 = ~n56882 & n56883 ;
  assign n56880 = \P2_P1_EBX_reg[25]/NET0131  & n46227 ;
  assign n56881 = n23782 & n46225 ;
  assign n56885 = ~n56880 & ~n56881 ;
  assign n56886 = ~n56884 & n56885 ;
  assign n56887 = n11623 & ~n56886 ;
  assign n56888 = \P2_P1_EBX_reg[25]/NET0131  & ~n21100 ;
  assign n56889 = ~n56887 & ~n56888 ;
  assign n56890 = ~n25783 & n25918 ;
  assign n56891 = \P1_P2_More_reg/NET0131  & ~n43212 ;
  assign n56892 = ~n56890 & ~n56891 ;
  assign n56893 = n11623 & ~n26062 ;
  assign n56894 = \P2_P1_More_reg/NET0131  & ~n21100 ;
  assign n56895 = ~n56893 & ~n56894 ;
  assign n56896 = ~n25700 & n47570 ;
  assign n56897 = ~n53116 & ~n56896 ;
  assign n56898 = n25918 & n56897 ;
  assign n56899 = n47529 & ~n56898 ;
  assign n56900 = \P1_P2_lWord_reg[0]/NET0131  & ~n56899 ;
  assign n56901 = \P1_P2_EAX_reg[0]/NET0131  & n47570 ;
  assign n56902 = ~n46749 & n53116 ;
  assign n56903 = ~n56901 & ~n56902 ;
  assign n56904 = n25918 & ~n56903 ;
  assign n56905 = ~n56900 & ~n56904 ;
  assign n56906 = \P1_P2_lWord_reg[10]/NET0131  & ~n53114 ;
  assign n56907 = \P1_P2_EAX_reg[10]/NET0131  & n47570 ;
  assign n56908 = n25776 & n47733 ;
  assign n56909 = ~n56907 & ~n56908 ;
  assign n56910 = n25918 & ~n56909 ;
  assign n56911 = ~n56906 & ~n56910 ;
  assign n56912 = \P1_P2_lWord_reg[11]/NET0131  & ~n53114 ;
  assign n56913 = \P1_P2_EAX_reg[11]/NET0131  & n47570 ;
  assign n56914 = n25776 & n44817 ;
  assign n56915 = ~n56913 & ~n56914 ;
  assign n56916 = n25918 & ~n56915 ;
  assign n56917 = ~n56912 & ~n56916 ;
  assign n56918 = \P1_P2_lWord_reg[12]/NET0131  & ~n53114 ;
  assign n56919 = \P1_P2_EAX_reg[12]/NET0131  & n47570 ;
  assign n56920 = n25776 & n49531 ;
  assign n56921 = ~n56919 & ~n56920 ;
  assign n56922 = n25918 & ~n56921 ;
  assign n56923 = ~n56918 & ~n56922 ;
  assign n56924 = \P1_P2_lWord_reg[13]/NET0131  & ~n53114 ;
  assign n56925 = \P1_P2_EAX_reg[13]/NET0131  & n47570 ;
  assign n56926 = n25776 & n48347 ;
  assign n56927 = ~n56925 & ~n56926 ;
  assign n56928 = n25918 & ~n56927 ;
  assign n56929 = ~n56924 & ~n56928 ;
  assign n56930 = \P1_P2_lWord_reg[14]/NET0131  & ~n53114 ;
  assign n56931 = \P1_P2_EAX_reg[14]/NET0131  & n47570 ;
  assign n56932 = n25776 & n46685 ;
  assign n56933 = ~n56931 & ~n56932 ;
  assign n56934 = n25918 & ~n56933 ;
  assign n56935 = ~n56930 & ~n56934 ;
  assign n56936 = \P1_P2_lWord_reg[15]/NET0131  & ~n53114 ;
  assign n56937 = n25776 & n48288 ;
  assign n56938 = \P1_P2_EAX_reg[15]/NET0131  & n25757 ;
  assign n56939 = ~n56937 & ~n56938 ;
  assign n56940 = ~n25770 & n25918 ;
  assign n56941 = ~n56939 & n56940 ;
  assign n56942 = ~n56936 & ~n56941 ;
  assign n56943 = \P1_P2_lWord_reg[1]/NET0131  & ~n56899 ;
  assign n56944 = \P1_P2_EAX_reg[1]/NET0131  & n47570 ;
  assign n56945 = ~n40746 & n53116 ;
  assign n56946 = ~n56944 & ~n56945 ;
  assign n56947 = n25918 & ~n56946 ;
  assign n56948 = ~n56943 & ~n56947 ;
  assign n56949 = \P1_P2_lWord_reg[2]/NET0131  & ~n56899 ;
  assign n56950 = \P1_P2_EAX_reg[2]/NET0131  & n47570 ;
  assign n56951 = n25776 & ~n35963 ;
  assign n56952 = n25773 & n56951 ;
  assign n56953 = ~n56950 & ~n56952 ;
  assign n56954 = n25918 & ~n56953 ;
  assign n56955 = ~n56949 & ~n56954 ;
  assign n56956 = \P1_P2_lWord_reg[3]/NET0131  & ~n56899 ;
  assign n56957 = \P1_P2_EAX_reg[3]/NET0131  & n47570 ;
  assign n56958 = n25776 & ~n29832 ;
  assign n56959 = n25773 & n56958 ;
  assign n56960 = ~n56957 & ~n56959 ;
  assign n56961 = n25918 & ~n56960 ;
  assign n56962 = ~n56956 & ~n56961 ;
  assign n56963 = \P1_P2_lWord_reg[4]/NET0131  & ~n53114 ;
  assign n56964 = \P1_P2_EAX_reg[4]/NET0131  & n47570 ;
  assign n56965 = ~n53117 & ~n56964 ;
  assign n56966 = n25918 & ~n56965 ;
  assign n56967 = ~n56963 & ~n56966 ;
  assign n56968 = \P1_P2_lWord_reg[5]/NET0131  & ~n56899 ;
  assign n56969 = ~n29860 & n53116 ;
  assign n56970 = \P1_P2_EAX_reg[5]/NET0131  & n47570 ;
  assign n56971 = ~n56969 & ~n56970 ;
  assign n56972 = n25918 & ~n56971 ;
  assign n56973 = ~n56968 & ~n56972 ;
  assign n56974 = \P1_P2_lWord_reg[6]/NET0131  & ~n56899 ;
  assign n56975 = \P1_P2_EAX_reg[6]/NET0131  & n47570 ;
  assign n56976 = ~n34449 & n53116 ;
  assign n56977 = ~n56975 & ~n56976 ;
  assign n56978 = n25918 & ~n56977 ;
  assign n56979 = ~n56974 & ~n56978 ;
  assign n56980 = \P1_P2_lWord_reg[7]/NET0131  & ~n56899 ;
  assign n56981 = \P1_P2_EAX_reg[7]/NET0131  & n47570 ;
  assign n56982 = n25776 & ~n28931 ;
  assign n56983 = n25773 & n56982 ;
  assign n56984 = ~n56981 & ~n56983 ;
  assign n56985 = n25918 & ~n56984 ;
  assign n56986 = ~n56980 & ~n56985 ;
  assign n56987 = \P1_P2_lWord_reg[8]/NET0131  & ~n53114 ;
  assign n56988 = \P1_P2_EAX_reg[8]/NET0131  & n25757 ;
  assign n56989 = ~n48661 & ~n56988 ;
  assign n56990 = n56940 & ~n56989 ;
  assign n56991 = ~n56987 & ~n56990 ;
  assign n56992 = \P1_P2_lWord_reg[9]/NET0131  & ~n53114 ;
  assign n56993 = \P1_P2_EAX_reg[9]/NET0131  & n47570 ;
  assign n56994 = ~n49721 & n53116 ;
  assign n56995 = ~n56993 & ~n56994 ;
  assign n56996 = n25918 & ~n56995 ;
  assign n56997 = ~n56992 & ~n56996 ;
  assign n56998 = n8355 & ~n26259 ;
  assign n56999 = \P1_P1_More_reg/NET0131  & ~n15326 ;
  assign n57000 = ~n56998 & ~n56999 ;
  assign n57001 = \P2_P1_uWord_reg[3]/NET0131  & ~n25156 ;
  assign n57002 = ~\P2_P1_EAX_reg[19]/NET0131  & ~n27390 ;
  assign n57003 = ~n27391 & ~n57002 ;
  assign n57004 = n24899 & n57003 ;
  assign n57005 = ~n47523 & ~n57004 ;
  assign n57006 = n11623 & ~n57005 ;
  assign n57007 = ~n57001 & ~n57006 ;
  assign n57008 = \P1_P2_uWord_reg[11]/NET0131  & ~n47529 ;
  assign n57009 = \P1_P2_uWord_reg[11]/NET0131  & ~n47572 ;
  assign n57010 = ~n56914 & ~n57009 ;
  assign n57011 = ~n56862 & n57010 ;
  assign n57012 = n25918 & ~n57011 ;
  assign n57013 = ~n57008 & ~n57012 ;
  assign n57014 = \P2_P2_EAX_reg[16]/NET0131  & ~n44508 ;
  assign n57047 = ~n44736 & ~n48181 ;
  assign n57048 = \P2_P2_EAX_reg[16]/NET0131  & ~n57047 ;
  assign n57056 = ~\P2_P2_EAX_reg[16]/NET0131  & n44732 ;
  assign n57057 = n44719 & n57056 ;
  assign n57049 = \P2_P2_EAX_reg[16]/NET0131  & ~n26641 ;
  assign n57053 = n26641 & ~n46792 ;
  assign n57054 = ~n57049 & ~n57053 ;
  assign n57055 = n26638 & ~n57054 ;
  assign n57026 = \P2_P2_InstQueue_reg[1][0]/NET0131  & n26330 ;
  assign n57024 = \P2_P2_InstQueue_reg[2][0]/NET0131  & n26325 ;
  assign n57015 = \P2_P2_InstQueue_reg[9][0]/NET0131  & n26300 ;
  assign n57016 = \P2_P2_InstQueue_reg[14][0]/NET0131  & n26310 ;
  assign n57031 = ~n57015 & ~n57016 ;
  assign n57041 = ~n57024 & n57031 ;
  assign n57042 = ~n57026 & n57041 ;
  assign n57027 = \P2_P2_InstQueue_reg[8][0]/NET0131  & n26318 ;
  assign n57028 = \P2_P2_InstQueue_reg[11][0]/NET0131  & n26334 ;
  assign n57036 = ~n57027 & ~n57028 ;
  assign n57029 = \P2_P2_InstQueue_reg[15][0]/NET0131  & n26313 ;
  assign n57030 = \P2_P2_InstQueue_reg[7][0]/NET0131  & n26307 ;
  assign n57037 = ~n57029 & ~n57030 ;
  assign n57038 = n57036 & n57037 ;
  assign n57021 = \P2_P2_InstQueue_reg[4][0]/NET0131  & n26338 ;
  assign n57022 = \P2_P2_InstQueue_reg[12][0]/NET0131  & n26304 ;
  assign n57034 = ~n57021 & ~n57022 ;
  assign n57023 = \P2_P2_InstQueue_reg[3][0]/NET0131  & n26322 ;
  assign n57025 = \P2_P2_InstQueue_reg[10][0]/NET0131  & n26327 ;
  assign n57035 = ~n57023 & ~n57025 ;
  assign n57039 = n57034 & n57035 ;
  assign n57017 = \P2_P2_InstQueue_reg[0][0]/NET0131  & n26336 ;
  assign n57018 = \P2_P2_InstQueue_reg[6][0]/NET0131  & n26332 ;
  assign n57032 = ~n57017 & ~n57018 ;
  assign n57019 = \P2_P2_InstQueue_reg[5][0]/NET0131  & n26316 ;
  assign n57020 = \P2_P2_InstQueue_reg[13][0]/NET0131  & n26320 ;
  assign n57033 = ~n57019 & ~n57020 ;
  assign n57040 = n57032 & n57033 ;
  assign n57043 = n57039 & n57040 ;
  assign n57044 = n57038 & n57043 ;
  assign n57045 = n57042 & n57044 ;
  assign n57046 = n44510 & ~n57045 ;
  assign n57050 = n26641 & ~n46777 ;
  assign n57051 = ~n57049 & ~n57050 ;
  assign n57052 = n26633 & ~n57051 ;
  assign n57058 = ~n57046 & ~n57052 ;
  assign n57059 = ~n57055 & n57058 ;
  assign n57060 = ~n57057 & n57059 ;
  assign n57061 = ~n57048 & n57060 ;
  assign n57062 = n26792 & ~n57061 ;
  assign n57063 = ~n57014 & ~n57062 ;
  assign n57064 = \P2_P2_EAX_reg[17]/NET0131  & ~n44508 ;
  assign n57065 = ~n44721 & n44732 ;
  assign n57067 = ~n44736 & ~n57065 ;
  assign n57068 = \P2_P2_EAX_reg[17]/NET0131  & ~n57067 ;
  assign n57066 = n44720 & n57065 ;
  assign n57101 = \P2_P2_EAX_reg[17]/NET0131  & ~n26641 ;
  assign n57105 = ~n53130 & ~n57101 ;
  assign n57106 = n26633 & ~n57105 ;
  assign n57080 = \P2_P2_InstQueue_reg[1][1]/NET0131  & n26330 ;
  assign n57078 = \P2_P2_InstQueue_reg[2][1]/NET0131  & n26325 ;
  assign n57069 = \P2_P2_InstQueue_reg[9][1]/NET0131  & n26300 ;
  assign n57070 = \P2_P2_InstQueue_reg[13][1]/NET0131  & n26320 ;
  assign n57085 = ~n57069 & ~n57070 ;
  assign n57095 = ~n57078 & n57085 ;
  assign n57096 = ~n57080 & n57095 ;
  assign n57081 = \P2_P2_InstQueue_reg[4][1]/NET0131  & n26338 ;
  assign n57082 = \P2_P2_InstQueue_reg[7][1]/NET0131  & n26307 ;
  assign n57090 = ~n57081 & ~n57082 ;
  assign n57083 = \P2_P2_InstQueue_reg[12][1]/NET0131  & n26304 ;
  assign n57084 = \P2_P2_InstQueue_reg[11][1]/NET0131  & n26334 ;
  assign n57091 = ~n57083 & ~n57084 ;
  assign n57092 = n57090 & n57091 ;
  assign n57075 = \P2_P2_InstQueue_reg[15][1]/NET0131  & n26313 ;
  assign n57076 = \P2_P2_InstQueue_reg[5][1]/NET0131  & n26316 ;
  assign n57088 = ~n57075 & ~n57076 ;
  assign n57077 = \P2_P2_InstQueue_reg[14][1]/NET0131  & n26310 ;
  assign n57079 = \P2_P2_InstQueue_reg[10][1]/NET0131  & n26327 ;
  assign n57089 = ~n57077 & ~n57079 ;
  assign n57093 = n57088 & n57089 ;
  assign n57071 = \P2_P2_InstQueue_reg[8][1]/NET0131  & n26318 ;
  assign n57072 = \P2_P2_InstQueue_reg[0][1]/NET0131  & n26336 ;
  assign n57086 = ~n57071 & ~n57072 ;
  assign n57073 = \P2_P2_InstQueue_reg[6][1]/NET0131  & n26332 ;
  assign n57074 = \P2_P2_InstQueue_reg[3][1]/NET0131  & n26322 ;
  assign n57087 = ~n57073 & ~n57074 ;
  assign n57094 = n57086 & n57087 ;
  assign n57097 = n57093 & n57094 ;
  assign n57098 = n57092 & n57097 ;
  assign n57099 = n57096 & n57098 ;
  assign n57100 = n44510 & ~n57099 ;
  assign n57102 = n26641 & ~n40789 ;
  assign n57103 = ~n57101 & ~n57102 ;
  assign n57104 = n26638 & ~n57103 ;
  assign n57107 = ~n57100 & ~n57104 ;
  assign n57108 = ~n57106 & n57107 ;
  assign n57109 = ~n57066 & n57108 ;
  assign n57110 = ~n57068 & n57109 ;
  assign n57111 = n26792 & ~n57110 ;
  assign n57112 = ~n57064 & ~n57111 ;
  assign n57113 = \P2_P2_EAX_reg[18]/NET0131  & ~n44508 ;
  assign n57146 = n46402 & ~n57065 ;
  assign n57147 = \P2_P2_EAX_reg[18]/NET0131  & ~n57146 ;
  assign n57152 = ~\P2_P2_EAX_reg[18]/NET0131  & n44732 ;
  assign n57153 = n44721 & n57152 ;
  assign n57125 = \P2_P2_InstQueue_reg[1][2]/NET0131  & n26330 ;
  assign n57123 = \P2_P2_InstQueue_reg[2][2]/NET0131  & n26325 ;
  assign n57114 = \P2_P2_InstQueue_reg[9][2]/NET0131  & n26300 ;
  assign n57115 = \P2_P2_InstQueue_reg[3][2]/NET0131  & n26322 ;
  assign n57130 = ~n57114 & ~n57115 ;
  assign n57140 = ~n57123 & n57130 ;
  assign n57141 = ~n57125 & n57140 ;
  assign n57126 = \P2_P2_InstQueue_reg[4][2]/NET0131  & n26338 ;
  assign n57127 = \P2_P2_InstQueue_reg[7][2]/NET0131  & n26307 ;
  assign n57135 = ~n57126 & ~n57127 ;
  assign n57128 = \P2_P2_InstQueue_reg[0][2]/NET0131  & n26336 ;
  assign n57129 = \P2_P2_InstQueue_reg[12][2]/NET0131  & n26304 ;
  assign n57136 = ~n57128 & ~n57129 ;
  assign n57137 = n57135 & n57136 ;
  assign n57120 = \P2_P2_InstQueue_reg[11][2]/NET0131  & n26334 ;
  assign n57121 = \P2_P2_InstQueue_reg[6][2]/NET0131  & n26332 ;
  assign n57133 = ~n57120 & ~n57121 ;
  assign n57122 = \P2_P2_InstQueue_reg[5][2]/NET0131  & n26316 ;
  assign n57124 = \P2_P2_InstQueue_reg[10][2]/NET0131  & n26327 ;
  assign n57134 = ~n57122 & ~n57124 ;
  assign n57138 = n57133 & n57134 ;
  assign n57116 = \P2_P2_InstQueue_reg[13][2]/NET0131  & n26320 ;
  assign n57117 = \P2_P2_InstQueue_reg[14][2]/NET0131  & n26310 ;
  assign n57131 = ~n57116 & ~n57117 ;
  assign n57118 = \P2_P2_InstQueue_reg[8][2]/NET0131  & n26318 ;
  assign n57119 = \P2_P2_InstQueue_reg[15][2]/NET0131  & n26313 ;
  assign n57132 = ~n57118 & ~n57119 ;
  assign n57139 = n57131 & n57132 ;
  assign n57142 = n57138 & n57139 ;
  assign n57143 = n57137 & n57142 ;
  assign n57144 = n57141 & n57143 ;
  assign n57145 = n44510 & ~n57144 ;
  assign n57148 = n26638 & ~n36006 ;
  assign n57149 = n26633 & ~n35991 ;
  assign n57150 = ~n57148 & ~n57149 ;
  assign n57151 = n26641 & ~n57150 ;
  assign n57154 = ~n57145 & ~n57151 ;
  assign n57155 = ~n57153 & n57154 ;
  assign n57156 = ~n57147 & n57155 ;
  assign n57157 = n26792 & ~n57156 ;
  assign n57158 = ~n57113 & ~n57157 ;
  assign n57159 = \P2_P2_EAX_reg[19]/NET0131  & ~n44508 ;
  assign n57161 = ~\P2_P2_EAX_reg[19]/NET0131  & ~n44722 ;
  assign n57162 = ~n44723 & n44732 ;
  assign n57163 = ~n57161 & n57162 ;
  assign n57160 = \P2_P2_EAX_reg[19]/NET0131  & ~n46402 ;
  assign n57164 = n26638 & ~n29903 ;
  assign n57165 = n26633 & ~n29888 ;
  assign n57166 = ~n57164 & ~n57165 ;
  assign n57167 = n26641 & ~n57166 ;
  assign n57179 = \P2_P2_InstQueue_reg[1][3]/NET0131  & n26330 ;
  assign n57177 = \P2_P2_InstQueue_reg[2][3]/NET0131  & n26325 ;
  assign n57168 = \P2_P2_InstQueue_reg[9][3]/NET0131  & n26300 ;
  assign n57169 = \P2_P2_InstQueue_reg[0][3]/NET0131  & n26336 ;
  assign n57184 = ~n57168 & ~n57169 ;
  assign n57194 = ~n57177 & n57184 ;
  assign n57195 = ~n57179 & n57194 ;
  assign n57180 = \P2_P2_InstQueue_reg[12][3]/NET0131  & n26304 ;
  assign n57181 = \P2_P2_InstQueue_reg[14][3]/NET0131  & n26310 ;
  assign n57189 = ~n57180 & ~n57181 ;
  assign n57182 = \P2_P2_InstQueue_reg[3][3]/NET0131  & n26322 ;
  assign n57183 = \P2_P2_InstQueue_reg[6][3]/NET0131  & n26332 ;
  assign n57190 = ~n57182 & ~n57183 ;
  assign n57191 = n57189 & n57190 ;
  assign n57174 = \P2_P2_InstQueue_reg[8][3]/NET0131  & n26318 ;
  assign n57175 = \P2_P2_InstQueue_reg[15][3]/NET0131  & n26313 ;
  assign n57187 = ~n57174 & ~n57175 ;
  assign n57176 = \P2_P2_InstQueue_reg[4][3]/NET0131  & n26338 ;
  assign n57178 = \P2_P2_InstQueue_reg[10][3]/NET0131  & n26327 ;
  assign n57188 = ~n57176 & ~n57178 ;
  assign n57192 = n57187 & n57188 ;
  assign n57170 = \P2_P2_InstQueue_reg[13][3]/NET0131  & n26320 ;
  assign n57171 = \P2_P2_InstQueue_reg[11][3]/NET0131  & n26334 ;
  assign n57185 = ~n57170 & ~n57171 ;
  assign n57172 = \P2_P2_InstQueue_reg[5][3]/NET0131  & n26316 ;
  assign n57173 = \P2_P2_InstQueue_reg[7][3]/NET0131  & n26307 ;
  assign n57186 = ~n57172 & ~n57173 ;
  assign n57193 = n57185 & n57186 ;
  assign n57196 = n57192 & n57193 ;
  assign n57197 = n57191 & n57196 ;
  assign n57198 = n57195 & n57197 ;
  assign n57199 = n44510 & ~n57198 ;
  assign n57200 = ~n57167 & ~n57199 ;
  assign n57201 = ~n57160 & n57200 ;
  assign n57202 = ~n57163 & n57201 ;
  assign n57203 = n26792 & ~n57202 ;
  assign n57204 = ~n57159 & ~n57203 ;
  assign n57206 = ~\P2_P2_EAX_reg[20]/NET0131  & ~n44723 ;
  assign n57207 = ~n44724 & n44732 ;
  assign n57208 = ~n57206 & n57207 ;
  assign n57205 = \P2_P2_EAX_reg[20]/NET0131  & ~n46402 ;
  assign n57209 = n26633 & ~n28016 ;
  assign n57210 = n26638 & ~n28037 ;
  assign n57211 = ~n57209 & ~n57210 ;
  assign n57212 = n26641 & ~n57211 ;
  assign n57224 = \P2_P2_InstQueue_reg[1][4]/NET0131  & n26330 ;
  assign n57222 = \P2_P2_InstQueue_reg[2][4]/NET0131  & n26325 ;
  assign n57213 = \P2_P2_InstQueue_reg[9][4]/NET0131  & n26300 ;
  assign n57214 = \P2_P2_InstQueue_reg[0][4]/NET0131  & n26336 ;
  assign n57229 = ~n57213 & ~n57214 ;
  assign n57239 = ~n57222 & n57229 ;
  assign n57240 = ~n57224 & n57239 ;
  assign n57225 = \P2_P2_InstQueue_reg[5][4]/NET0131  & n26316 ;
  assign n57226 = \P2_P2_InstQueue_reg[3][4]/NET0131  & n26322 ;
  assign n57234 = ~n57225 & ~n57226 ;
  assign n57227 = \P2_P2_InstQueue_reg[4][4]/NET0131  & n26338 ;
  assign n57228 = \P2_P2_InstQueue_reg[12][4]/NET0131  & n26304 ;
  assign n57235 = ~n57227 & ~n57228 ;
  assign n57236 = n57234 & n57235 ;
  assign n57219 = \P2_P2_InstQueue_reg[6][4]/NET0131  & n26332 ;
  assign n57220 = \P2_P2_InstQueue_reg[13][4]/NET0131  & n26320 ;
  assign n57232 = ~n57219 & ~n57220 ;
  assign n57221 = \P2_P2_InstQueue_reg[11][4]/NET0131  & n26334 ;
  assign n57223 = \P2_P2_InstQueue_reg[10][4]/NET0131  & n26327 ;
  assign n57233 = ~n57221 & ~n57223 ;
  assign n57237 = n57232 & n57233 ;
  assign n57215 = \P2_P2_InstQueue_reg[7][4]/NET0131  & n26307 ;
  assign n57216 = \P2_P2_InstQueue_reg[14][4]/NET0131  & n26310 ;
  assign n57230 = ~n57215 & ~n57216 ;
  assign n57217 = \P2_P2_InstQueue_reg[8][4]/NET0131  & n26318 ;
  assign n57218 = \P2_P2_InstQueue_reg[15][4]/NET0131  & n26313 ;
  assign n57231 = ~n57217 & ~n57218 ;
  assign n57238 = n57230 & n57231 ;
  assign n57241 = n57237 & n57238 ;
  assign n57242 = n57236 & n57241 ;
  assign n57243 = n57240 & n57242 ;
  assign n57244 = n44510 & ~n57243 ;
  assign n57245 = ~n57212 & ~n57244 ;
  assign n57246 = ~n57205 & n57245 ;
  assign n57247 = ~n57208 & n57246 ;
  assign n57248 = n26792 & ~n57247 ;
  assign n57249 = \P2_P2_EAX_reg[20]/NET0131  & ~n44508 ;
  assign n57250 = ~n57248 & ~n57249 ;
  assign n57251 = \P2_P2_EAX_reg[21]/NET0131  & ~n44508 ;
  assign n57253 = ~\P2_P2_EAX_reg[21]/NET0131  & ~n44724 ;
  assign n57254 = ~n44725 & n44732 ;
  assign n57255 = ~n57253 & n57254 ;
  assign n57252 = \P2_P2_EAX_reg[21]/NET0131  & ~n46402 ;
  assign n57256 = n26638 & ~n39038 ;
  assign n57257 = n26633 & ~n39023 ;
  assign n57258 = ~n57256 & ~n57257 ;
  assign n57259 = n26641 & ~n57258 ;
  assign n57271 = \P2_P2_InstQueue_reg[1][5]/NET0131  & n26330 ;
  assign n57269 = \P2_P2_InstQueue_reg[2][5]/NET0131  & n26325 ;
  assign n57260 = \P2_P2_InstQueue_reg[9][5]/NET0131  & n26300 ;
  assign n57261 = \P2_P2_InstQueue_reg[13][5]/NET0131  & n26320 ;
  assign n57276 = ~n57260 & ~n57261 ;
  assign n57286 = ~n57269 & n57276 ;
  assign n57287 = ~n57271 & n57286 ;
  assign n57272 = \P2_P2_InstQueue_reg[7][5]/NET0131  & n26307 ;
  assign n57273 = \P2_P2_InstQueue_reg[12][5]/NET0131  & n26304 ;
  assign n57281 = ~n57272 & ~n57273 ;
  assign n57274 = \P2_P2_InstQueue_reg[5][5]/NET0131  & n26316 ;
  assign n57275 = \P2_P2_InstQueue_reg[6][5]/NET0131  & n26332 ;
  assign n57282 = ~n57274 & ~n57275 ;
  assign n57283 = n57281 & n57282 ;
  assign n57266 = \P2_P2_InstQueue_reg[15][5]/NET0131  & n26313 ;
  assign n57267 = \P2_P2_InstQueue_reg[11][5]/NET0131  & n26334 ;
  assign n57279 = ~n57266 & ~n57267 ;
  assign n57268 = \P2_P2_InstQueue_reg[4][5]/NET0131  & n26338 ;
  assign n57270 = \P2_P2_InstQueue_reg[10][5]/NET0131  & n26327 ;
  assign n57280 = ~n57268 & ~n57270 ;
  assign n57284 = n57279 & n57280 ;
  assign n57262 = \P2_P2_InstQueue_reg[3][5]/NET0131  & n26322 ;
  assign n57263 = \P2_P2_InstQueue_reg[0][5]/NET0131  & n26336 ;
  assign n57277 = ~n57262 & ~n57263 ;
  assign n57264 = \P2_P2_InstQueue_reg[14][5]/NET0131  & n26310 ;
  assign n57265 = \P2_P2_InstQueue_reg[8][5]/NET0131  & n26318 ;
  assign n57278 = ~n57264 & ~n57265 ;
  assign n57285 = n57277 & n57278 ;
  assign n57288 = n57284 & n57285 ;
  assign n57289 = n57283 & n57288 ;
  assign n57290 = n57287 & n57289 ;
  assign n57291 = n44510 & ~n57290 ;
  assign n57292 = ~n57259 & ~n57291 ;
  assign n57293 = ~n57252 & n57292 ;
  assign n57294 = ~n57255 & n57293 ;
  assign n57295 = n26792 & ~n57294 ;
  assign n57296 = ~n57251 & ~n57295 ;
  assign n57297 = \P2_P2_EAX_reg[22]/NET0131  & ~n44508 ;
  assign n57299 = ~\P2_P2_EAX_reg[22]/NET0131  & ~n44725 ;
  assign n57300 = ~n44726 & n44732 ;
  assign n57301 = ~n57299 & n57300 ;
  assign n57298 = \P2_P2_EAX_reg[22]/NET0131  & ~n46402 ;
  assign n57302 = n26638 & ~n34492 ;
  assign n57303 = n26633 & ~n34477 ;
  assign n57304 = ~n57302 & ~n57303 ;
  assign n57305 = n26641 & ~n57304 ;
  assign n57317 = \P2_P2_InstQueue_reg[1][6]/NET0131  & n26330 ;
  assign n57315 = \P2_P2_InstQueue_reg[2][6]/NET0131  & n26325 ;
  assign n57306 = \P2_P2_InstQueue_reg[9][6]/NET0131  & n26300 ;
  assign n57307 = \P2_P2_InstQueue_reg[15][6]/NET0131  & n26313 ;
  assign n57322 = ~n57306 & ~n57307 ;
  assign n57332 = ~n57315 & n57322 ;
  assign n57333 = ~n57317 & n57332 ;
  assign n57318 = \P2_P2_InstQueue_reg[12][6]/NET0131  & n26304 ;
  assign n57319 = \P2_P2_InstQueue_reg[14][6]/NET0131  & n26310 ;
  assign n57327 = ~n57318 & ~n57319 ;
  assign n57320 = \P2_P2_InstQueue_reg[11][6]/NET0131  & n26334 ;
  assign n57321 = \P2_P2_InstQueue_reg[6][6]/NET0131  & n26332 ;
  assign n57328 = ~n57320 & ~n57321 ;
  assign n57329 = n57327 & n57328 ;
  assign n57312 = \P2_P2_InstQueue_reg[3][6]/NET0131  & n26322 ;
  assign n57313 = \P2_P2_InstQueue_reg[7][6]/NET0131  & n26307 ;
  assign n57325 = ~n57312 & ~n57313 ;
  assign n57314 = \P2_P2_InstQueue_reg[0][6]/NET0131  & n26336 ;
  assign n57316 = \P2_P2_InstQueue_reg[10][6]/NET0131  & n26327 ;
  assign n57326 = ~n57314 & ~n57316 ;
  assign n57330 = n57325 & n57326 ;
  assign n57308 = \P2_P2_InstQueue_reg[5][6]/NET0131  & n26316 ;
  assign n57309 = \P2_P2_InstQueue_reg[8][6]/NET0131  & n26318 ;
  assign n57323 = ~n57308 & ~n57309 ;
  assign n57310 = \P2_P2_InstQueue_reg[13][6]/NET0131  & n26320 ;
  assign n57311 = \P2_P2_InstQueue_reg[4][6]/NET0131  & n26338 ;
  assign n57324 = ~n57310 & ~n57311 ;
  assign n57331 = n57323 & n57324 ;
  assign n57334 = n57330 & n57331 ;
  assign n57335 = n57329 & n57334 ;
  assign n57336 = n57333 & n57335 ;
  assign n57337 = n44510 & ~n57336 ;
  assign n57338 = ~n57305 & ~n57337 ;
  assign n57339 = ~n57298 & n57338 ;
  assign n57340 = ~n57301 & n57339 ;
  assign n57341 = n26792 & ~n57340 ;
  assign n57342 = ~n57297 & ~n57341 ;
  assign n57347 = ~\P2_P2_EAX_reg[23]/NET0131  & ~n44726 ;
  assign n57348 = ~n44727 & n44732 ;
  assign n57349 = ~n57347 & n57348 ;
  assign n57350 = \P2_P2_EAX_reg[23]/NET0131  & n44736 ;
  assign n57351 = \P2_P2_EAX_reg[23]/NET0131  & ~n26641 ;
  assign n57354 = n26641 & ~n28963 ;
  assign n57355 = ~n57351 & ~n57354 ;
  assign n57356 = n26638 & ~n57355 ;
  assign n57343 = n44541 & n44572 ;
  assign n57344 = n26611 & ~n44573 ;
  assign n57345 = ~n57343 & n57344 ;
  assign n57346 = n26582 & n57345 ;
  assign n57352 = ~n48889 & ~n57351 ;
  assign n57353 = n26633 & ~n57352 ;
  assign n57357 = ~n57346 & ~n57353 ;
  assign n57358 = ~n57356 & n57357 ;
  assign n57359 = ~n57350 & n57358 ;
  assign n57360 = ~n57349 & n57359 ;
  assign n57361 = n26792 & ~n57360 ;
  assign n57362 = \P2_P2_EAX_reg[23]/NET0131  & ~n44508 ;
  assign n57363 = ~n57361 & ~n57362 ;
  assign n57364 = \P2_P2_EAX_reg[24]/NET0131  & ~n44508 ;
  assign n57368 = ~n44736 & ~n57348 ;
  assign n57369 = \P2_P2_EAX_reg[24]/NET0131  & ~n57368 ;
  assign n57376 = ~\P2_P2_EAX_reg[24]/NET0131  & n44732 ;
  assign n57377 = n44727 & n57376 ;
  assign n57370 = \P2_P2_EAX_reg[24]/NET0131  & ~n26641 ;
  assign n57374 = ~n48902 & ~n57370 ;
  assign n57375 = n26633 & ~n57374 ;
  assign n57365 = ~n44573 & n44604 ;
  assign n57366 = ~n44605 & ~n57365 ;
  assign n57367 = n44510 & n57366 ;
  assign n57371 = n26641 & ~n46788 ;
  assign n57372 = ~n57370 & ~n57371 ;
  assign n57373 = n26638 & ~n57372 ;
  assign n57378 = ~n57367 & ~n57373 ;
  assign n57379 = ~n57375 & n57378 ;
  assign n57380 = ~n57377 & n57379 ;
  assign n57381 = ~n57369 & n57380 ;
  assign n57382 = n26792 & ~n57381 ;
  assign n57383 = ~n57364 & ~n57382 ;
  assign n57384 = \P2_P2_EAX_reg[28]/NET0131  & ~n44508 ;
  assign n57387 = \P2_P2_EAX_reg[28]/NET0131  & ~n44737 ;
  assign n57385 = ~\P2_P2_EAX_reg[28]/NET0131  & n44732 ;
  assign n57386 = n44731 & n57385 ;
  assign n57391 = ~n44702 & n46318 ;
  assign n57392 = ~n46319 & ~n57391 ;
  assign n57393 = n44510 & n57392 ;
  assign n57388 = \P2_P2_EAX_reg[28]/NET0131  & ~n26641 ;
  assign n57389 = ~n48789 & ~n57388 ;
  assign n57390 = n26633 & ~n57389 ;
  assign n57394 = n26641 & ~n28030 ;
  assign n57395 = ~n57388 & ~n57394 ;
  assign n57396 = n26638 & ~n57395 ;
  assign n57397 = ~n57390 & ~n57396 ;
  assign n57398 = ~n57393 & n57397 ;
  assign n57399 = ~n57386 & n57398 ;
  assign n57400 = ~n57387 & n57399 ;
  assign n57401 = n26792 & ~n57400 ;
  assign n57402 = ~n57384 & ~n57401 ;
  assign n57405 = ~\P2_P2_EBX_reg[25]/NET0131  & ~n46443 ;
  assign n57406 = n26662 & ~n46444 ;
  assign n57407 = ~n57405 & n57406 ;
  assign n57403 = \P2_P2_EBX_reg[25]/NET0131  & n46417 ;
  assign n57404 = n46416 & n53144 ;
  assign n57408 = ~n57403 & ~n57404 ;
  assign n57409 = ~n57407 & n57408 ;
  assign n57410 = n26792 & ~n57409 ;
  assign n57411 = \P2_P2_EBX_reg[25]/NET0131  & ~n44508 ;
  assign n57412 = ~n57410 & ~n57411 ;
  assign n57415 = ~\P1_P3_EBX_reg[25]/NET0131  & ~n46505 ;
  assign n57416 = n9108 & ~n46506 ;
  assign n57417 = ~n57415 & n57416 ;
  assign n57413 = \P1_P3_EBX_reg[25]/NET0131  & n46480 ;
  assign n57414 = n22358 & n46479 ;
  assign n57418 = ~n57413 & ~n57414 ;
  assign n57419 = ~n57417 & n57418 ;
  assign n57420 = n9241 & ~n57419 ;
  assign n57421 = \P1_P3_EBX_reg[25]/NET0131  & ~n16968 ;
  assign n57422 = ~n57420 & ~n57421 ;
  assign n57423 = ~n26658 & n26792 ;
  assign n57424 = \P2_P2_More_reg/NET0131  & ~n44508 ;
  assign n57425 = ~n57423 & ~n57424 ;
  assign n57428 = ~\P1_P1_EBX_reg[25]/NET0131  & ~n46560 ;
  assign n57429 = n26146 & ~n46561 ;
  assign n57430 = ~n57428 & n57429 ;
  assign n57426 = n23944 & n46535 ;
  assign n57427 = \P1_P1_EBX_reg[25]/NET0131  & ~n46533 ;
  assign n57431 = ~n57426 & ~n57427 ;
  assign n57432 = ~n57430 & n57431 ;
  assign n57433 = n8355 & ~n57432 ;
  assign n57434 = \P1_P1_EBX_reg[25]/NET0131  & ~n15326 ;
  assign n57435 = ~n57433 & ~n57434 ;
  assign n57436 = n26792 & ~n47686 ;
  assign n57437 = n47642 & ~n57436 ;
  assign n57438 = \P2_P2_lWord_reg[0]/NET0131  & ~n57437 ;
  assign n57439 = n26633 & n57050 ;
  assign n57440 = \P2_P2_EAX_reg[0]/NET0131  & n26786 ;
  assign n57441 = ~n57439 & ~n57440 ;
  assign n57442 = n26792 & ~n57441 ;
  assign n57443 = ~n57438 & ~n57442 ;
  assign n57444 = \P2_P2_lWord_reg[10]/NET0131  & ~n57437 ;
  assign n57445 = ~n47590 & n47676 ;
  assign n57446 = \P2_P2_EAX_reg[10]/NET0131  & n26643 ;
  assign n57447 = ~n57445 & ~n57446 ;
  assign n57448 = ~n26640 & n26792 ;
  assign n57449 = ~n57447 & n57448 ;
  assign n57450 = ~n57444 & ~n57449 ;
  assign n57451 = \P2_P2_lWord_reg[11]/NET0131  & ~n47642 ;
  assign n57452 = ~n26633 & ~n26786 ;
  assign n57453 = ~n32741 & ~n47683 ;
  assign n57454 = ~n57452 & n57453 ;
  assign n57455 = \P2_P2_lWord_reg[11]/NET0131  & ~n57454 ;
  assign n57456 = n26633 & n44744 ;
  assign n57457 = \P2_P2_EAX_reg[11]/NET0131  & n26786 ;
  assign n57458 = ~n57456 & ~n57457 ;
  assign n57459 = ~n57455 & n57458 ;
  assign n57460 = n26792 & ~n57459 ;
  assign n57461 = ~n57451 & ~n57460 ;
  assign n57462 = \P2_P2_lWord_reg[12]/NET0131  & ~n57437 ;
  assign n57463 = \P2_P2_EAX_reg[12]/NET0131  & n26643 ;
  assign n57464 = ~n47680 & ~n57463 ;
  assign n57465 = n57448 & ~n57464 ;
  assign n57466 = ~n57462 & ~n57465 ;
  assign n57467 = \P2_P2_lWord_reg[13]/NET0131  & ~n57437 ;
  assign n57468 = \P2_P2_EAX_reg[13]/NET0131  & n26643 ;
  assign n57469 = n47676 & ~n48208 ;
  assign n57470 = ~n57468 & ~n57469 ;
  assign n57471 = n57448 & ~n57470 ;
  assign n57472 = ~n57467 & ~n57471 ;
  assign n57473 = \P2_P2_lWord_reg[14]/NET0131  & ~n57437 ;
  assign n57474 = \P2_P2_EAX_reg[14]/NET0131  & n26643 ;
  assign n57475 = ~n46283 & n47676 ;
  assign n57476 = ~n57474 & ~n57475 ;
  assign n57477 = n57448 & ~n57476 ;
  assign n57478 = ~n57473 & ~n57477 ;
  assign n57479 = \P1_P1_uWord_reg[3]/NET0131  & ~n24515 ;
  assign n57481 = \P1_P1_uWord_reg[3]/NET0131  & n25363 ;
  assign n57482 = ~n24648 & ~n57481 ;
  assign n57483 = n15334 & ~n57482 ;
  assign n57480 = \P1_P1_uWord_reg[3]/NET0131  & n24505 ;
  assign n57484 = ~\P1_P1_EAX_reg[19]/NET0131  & ~n25350 ;
  assign n57485 = ~n25351 & ~n57484 ;
  assign n57486 = n24503 & n57485 ;
  assign n57487 = ~n57480 & ~n57486 ;
  assign n57488 = ~n57483 & n57487 ;
  assign n57489 = n8355 & ~n57488 ;
  assign n57490 = ~n57479 & ~n57489 ;
  assign n57491 = \P2_P2_lWord_reg[15]/NET0131  & ~n57437 ;
  assign n57492 = n47676 & ~n48189 ;
  assign n57493 = \P2_P2_EAX_reg[15]/NET0131  & n26643 ;
  assign n57494 = ~n57492 & ~n57493 ;
  assign n57495 = n57448 & ~n57494 ;
  assign n57496 = ~n57491 & ~n57495 ;
  assign n57497 = \P2_P2_EAX_reg[1]/NET0131  & n26643 ;
  assign n57498 = ~n40774 & n47676 ;
  assign n57499 = ~n57497 & ~n57498 ;
  assign n57500 = ~n26640 & ~n57499 ;
  assign n57501 = \P2_P2_lWord_reg[1]/NET0131  & ~n47686 ;
  assign n57502 = ~n57500 & ~n57501 ;
  assign n57503 = n26792 & ~n57502 ;
  assign n57504 = \P2_P2_lWord_reg[1]/NET0131  & ~n47642 ;
  assign n57505 = ~n57503 & ~n57504 ;
  assign n57506 = \P2_P2_EAX_reg[2]/NET0131  & n26643 ;
  assign n57507 = ~n26286 & n57149 ;
  assign n57508 = ~n57506 & ~n57507 ;
  assign n57509 = ~n26640 & ~n57508 ;
  assign n57510 = \P2_P2_lWord_reg[2]/NET0131  & ~n47686 ;
  assign n57511 = ~n57509 & ~n57510 ;
  assign n57512 = n26792 & ~n57511 ;
  assign n57513 = \P2_P2_lWord_reg[2]/NET0131  & ~n47642 ;
  assign n57514 = ~n57512 & ~n57513 ;
  assign n57515 = \P2_P2_EAX_reg[3]/NET0131  & n26643 ;
  assign n57516 = ~n29888 & n47676 ;
  assign n57517 = ~n57515 & ~n57516 ;
  assign n57518 = ~n26640 & ~n57517 ;
  assign n57519 = \P2_P2_lWord_reg[3]/NET0131  & ~n47686 ;
  assign n57520 = ~n57518 & ~n57519 ;
  assign n57521 = n26792 & ~n57520 ;
  assign n57522 = \P2_P2_lWord_reg[3]/NET0131  & ~n47642 ;
  assign n57523 = ~n57521 & ~n57522 ;
  assign n57524 = \P2_P2_EAX_reg[4]/NET0131  & n26643 ;
  assign n57525 = ~n28016 & n47676 ;
  assign n57526 = ~n57524 & ~n57525 ;
  assign n57527 = ~n26640 & ~n57526 ;
  assign n57528 = \P2_P2_lWord_reg[4]/NET0131  & ~n47686 ;
  assign n57529 = ~n57527 & ~n57528 ;
  assign n57530 = n26792 & ~n57529 ;
  assign n57531 = \P2_P2_lWord_reg[4]/NET0131  & ~n47642 ;
  assign n57532 = ~n57530 & ~n57531 ;
  assign n57533 = \P2_P2_EAX_reg[5]/NET0131  & n26643 ;
  assign n57534 = ~n39023 & n47676 ;
  assign n57535 = ~n57533 & ~n57534 ;
  assign n57536 = ~n26640 & ~n57535 ;
  assign n57537 = \P2_P2_lWord_reg[5]/NET0131  & ~n47686 ;
  assign n57538 = ~n57536 & ~n57537 ;
  assign n57539 = n26792 & ~n57538 ;
  assign n57540 = \P2_P2_lWord_reg[5]/NET0131  & ~n47642 ;
  assign n57541 = ~n57539 & ~n57540 ;
  assign n57542 = \P2_P2_EAX_reg[6]/NET0131  & n26643 ;
  assign n57543 = ~n34477 & n47676 ;
  assign n57544 = ~n57542 & ~n57543 ;
  assign n57545 = ~n26640 & ~n57544 ;
  assign n57546 = \P2_P2_lWord_reg[6]/NET0131  & ~n47686 ;
  assign n57547 = ~n57545 & ~n57546 ;
  assign n57548 = n26792 & ~n57547 ;
  assign n57549 = \P2_P2_lWord_reg[6]/NET0131  & ~n47642 ;
  assign n57550 = ~n57548 & ~n57549 ;
  assign n57551 = \P2_P2_EAX_reg[7]/NET0131  & n26643 ;
  assign n57552 = ~n28951 & n47676 ;
  assign n57553 = ~n57551 & ~n57552 ;
  assign n57554 = ~n26640 & ~n57553 ;
  assign n57555 = \P2_P2_lWord_reg[7]/NET0131  & ~n47686 ;
  assign n57556 = ~n57554 & ~n57555 ;
  assign n57557 = n26792 & ~n57556 ;
  assign n57558 = \P2_P2_lWord_reg[7]/NET0131  & ~n47642 ;
  assign n57559 = ~n57557 & ~n57558 ;
  assign n57560 = \P2_P2_lWord_reg[8]/NET0131  & ~n57437 ;
  assign n57561 = \P2_P2_EAX_reg[8]/NET0131  & n26643 ;
  assign n57562 = ~n49031 & ~n57561 ;
  assign n57563 = n57448 & ~n57562 ;
  assign n57564 = ~n57560 & ~n57563 ;
  assign n57565 = \P2_P2_lWord_reg[9]/NET0131  & ~n57437 ;
  assign n57566 = \P2_P2_EAX_reg[9]/NET0131  & n26643 ;
  assign n57567 = n47676 & ~n48946 ;
  assign n57568 = ~n57566 & ~n57567 ;
  assign n57569 = n57448 & ~n57568 ;
  assign n57570 = ~n57565 & ~n57569 ;
  assign n57571 = \P2_P2_uWord_reg[11]/NET0131  & ~n47642 ;
  assign n57572 = \P2_P2_uWord_reg[11]/NET0131  & ~n47686 ;
  assign n57573 = ~n57456 & ~n57572 ;
  assign n57574 = ~n56834 & n57573 ;
  assign n57575 = n26792 & ~n57574 ;
  assign n57576 = ~n57571 & ~n57575 ;
  assign n57609 = ~\P2_P3_EAX_reg[16]/NET0131  & ~n42847 ;
  assign n57610 = n42539 & ~n42848 ;
  assign n57611 = ~n57609 & n57610 ;
  assign n57612 = \P2_P3_EAX_reg[16]/NET0131  & n42542 ;
  assign n57613 = \P2_P3_EAX_reg[16]/NET0131  & ~n27227 ;
  assign n57617 = ~n53248 & ~n57613 ;
  assign n57618 = n27122 & ~n57617 ;
  assign n57586 = \P2_P3_InstQueue_reg[10][0]/NET0131  & n26839 ;
  assign n57577 = \P2_P3_InstQueue_reg[4][0]/NET0131  & n26831 ;
  assign n57578 = \P2_P3_InstQueue_reg[3][0]/NET0131  & n26812 ;
  assign n57593 = ~n57577 & ~n57578 ;
  assign n57602 = ~n57586 & n57593 ;
  assign n57587 = \P2_P3_InstQueue_reg[2][0]/NET0131  & n26837 ;
  assign n57590 = \P2_P3_InstQueue_reg[1][0]/NET0131  & n26845 ;
  assign n57603 = ~n57587 & ~n57590 ;
  assign n57604 = n57602 & n57603 ;
  assign n57592 = \P2_P3_InstQueue_reg[6][0]/NET0131  & n26847 ;
  assign n57589 = \P2_P3_InstQueue_reg[11][0]/NET0131  & n26827 ;
  assign n57591 = \P2_P3_InstQueue_reg[8][0]/NET0131  & n26822 ;
  assign n57598 = ~n57589 & ~n57591 ;
  assign n57599 = ~n57592 & n57598 ;
  assign n57583 = \P2_P3_InstQueue_reg[5][0]/NET0131  & n26843 ;
  assign n57584 = \P2_P3_InstQueue_reg[12][0]/NET0131  & n26833 ;
  assign n57596 = ~n57583 & ~n57584 ;
  assign n57585 = \P2_P3_InstQueue_reg[15][0]/NET0131  & n26829 ;
  assign n57588 = \P2_P3_InstQueue_reg[9][0]/NET0131  & n26841 ;
  assign n57597 = ~n57585 & ~n57588 ;
  assign n57600 = n57596 & n57597 ;
  assign n57579 = \P2_P3_InstQueue_reg[14][0]/NET0131  & n26849 ;
  assign n57580 = \P2_P3_InstQueue_reg[7][0]/NET0131  & n26815 ;
  assign n57594 = ~n57579 & ~n57580 ;
  assign n57581 = \P2_P3_InstQueue_reg[0][0]/NET0131  & n26825 ;
  assign n57582 = \P2_P3_InstQueue_reg[13][0]/NET0131  & n26819 ;
  assign n57595 = ~n57581 & ~n57582 ;
  assign n57601 = n57594 & n57595 ;
  assign n57605 = n57600 & n57601 ;
  assign n57606 = n57599 & n57605 ;
  assign n57607 = n57604 & n57606 ;
  assign n57608 = n42538 & ~n57607 ;
  assign n57614 = \P2_buf2_reg[16]/NET0131  & n27227 ;
  assign n57615 = ~n57613 & ~n57614 ;
  assign n57616 = n27186 & ~n57615 ;
  assign n57619 = ~n57608 & ~n57616 ;
  assign n57620 = ~n57618 & n57619 ;
  assign n57621 = ~n57612 & n57620 ;
  assign n57622 = ~n57611 & n57621 ;
  assign n57623 = n27308 & ~n57622 ;
  assign n57624 = \P2_P3_EAX_reg[16]/NET0131  & ~n42872 ;
  assign n57625 = ~n57623 & ~n57624 ;
  assign n57626 = \P2_P3_EAX_reg[17]/NET0131  & ~n42872 ;
  assign n57659 = ~n42542 & ~n57610 ;
  assign n57660 = \P2_P3_EAX_reg[17]/NET0131  & ~n57659 ;
  assign n57668 = ~\P2_P3_EAX_reg[17]/NET0131  & n42539 ;
  assign n57669 = n42848 & n57668 ;
  assign n57662 = \P2_P3_EAX_reg[17]/NET0131  & ~n27227 ;
  assign n57665 = \P2_buf2_reg[17]/NET0131  & n27227 ;
  assign n57666 = ~n57662 & ~n57665 ;
  assign n57667 = n27186 & ~n57666 ;
  assign n57635 = \P2_P3_InstQueue_reg[1][1]/NET0131  & n26845 ;
  assign n57627 = \P2_P3_InstQueue_reg[4][1]/NET0131  & n26831 ;
  assign n57628 = \P2_P3_InstQueue_reg[8][1]/NET0131  & n26822 ;
  assign n57643 = ~n57627 & ~n57628 ;
  assign n57652 = ~n57635 & n57643 ;
  assign n57637 = \P2_P3_InstQueue_reg[2][1]/NET0131  & n26837 ;
  assign n57638 = \P2_P3_InstQueue_reg[10][1]/NET0131  & n26839 ;
  assign n57653 = ~n57637 & ~n57638 ;
  assign n57654 = n57652 & n57653 ;
  assign n57642 = \P2_P3_InstQueue_reg[0][1]/NET0131  & n26825 ;
  assign n57640 = \P2_P3_InstQueue_reg[14][1]/NET0131  & n26849 ;
  assign n57641 = \P2_P3_InstQueue_reg[6][1]/NET0131  & n26847 ;
  assign n57648 = ~n57640 & ~n57641 ;
  assign n57649 = ~n57642 & n57648 ;
  assign n57633 = \P2_P3_InstQueue_reg[3][1]/NET0131  & n26812 ;
  assign n57634 = \P2_P3_InstQueue_reg[7][1]/NET0131  & n26815 ;
  assign n57646 = ~n57633 & ~n57634 ;
  assign n57636 = \P2_P3_InstQueue_reg[9][1]/NET0131  & n26841 ;
  assign n57639 = \P2_P3_InstQueue_reg[13][1]/NET0131  & n26819 ;
  assign n57647 = ~n57636 & ~n57639 ;
  assign n57650 = n57646 & n57647 ;
  assign n57629 = \P2_P3_InstQueue_reg[5][1]/NET0131  & n26843 ;
  assign n57630 = \P2_P3_InstQueue_reg[12][1]/NET0131  & n26833 ;
  assign n57644 = ~n57629 & ~n57630 ;
  assign n57631 = \P2_P3_InstQueue_reg[11][1]/NET0131  & n26827 ;
  assign n57632 = \P2_P3_InstQueue_reg[15][1]/NET0131  & n26829 ;
  assign n57645 = ~n57631 & ~n57632 ;
  assign n57651 = n57644 & n57645 ;
  assign n57655 = n57650 & n57651 ;
  assign n57656 = n57649 & n57655 ;
  assign n57657 = n57654 & n57656 ;
  assign n57658 = n42538 & ~n57657 ;
  assign n57661 = \P2_buf2_reg[1]/NET0131  & n27227 ;
  assign n57663 = ~n57661 & ~n57662 ;
  assign n57664 = n27122 & ~n57663 ;
  assign n57670 = ~n57658 & ~n57664 ;
  assign n57671 = ~n57667 & n57670 ;
  assign n57672 = ~n57669 & n57671 ;
  assign n57673 = ~n57660 & n57672 ;
  assign n57674 = n27308 & ~n57673 ;
  assign n57675 = ~n57626 & ~n57674 ;
  assign n57677 = ~\P2_P3_EAX_reg[18]/NET0131  & ~n42849 ;
  assign n57678 = n42539 & ~n42850 ;
  assign n57679 = ~n57677 & n57678 ;
  assign n57676 = \P2_P3_EAX_reg[18]/NET0131  & ~n42543 ;
  assign n57680 = \P2_buf2_reg[2]/NET0131  & n27122 ;
  assign n57681 = \P2_buf2_reg[18]/NET0131  & n27186 ;
  assign n57682 = ~n57680 & ~n57681 ;
  assign n57683 = n27227 & ~n57682 ;
  assign n57692 = \P2_P3_InstQueue_reg[1][2]/NET0131  & n26845 ;
  assign n57684 = \P2_P3_InstQueue_reg[0][2]/NET0131  & n26825 ;
  assign n57685 = \P2_P3_InstQueue_reg[3][2]/NET0131  & n26812 ;
  assign n57700 = ~n57684 & ~n57685 ;
  assign n57709 = ~n57692 & n57700 ;
  assign n57694 = \P2_P3_InstQueue_reg[10][2]/NET0131  & n26839 ;
  assign n57695 = \P2_P3_InstQueue_reg[2][2]/NET0131  & n26837 ;
  assign n57710 = ~n57694 & ~n57695 ;
  assign n57711 = n57709 & n57710 ;
  assign n57699 = \P2_P3_InstQueue_reg[14][2]/NET0131  & n26849 ;
  assign n57697 = \P2_P3_InstQueue_reg[6][2]/NET0131  & n26847 ;
  assign n57698 = \P2_P3_InstQueue_reg[5][2]/NET0131  & n26843 ;
  assign n57705 = ~n57697 & ~n57698 ;
  assign n57706 = ~n57699 & n57705 ;
  assign n57690 = \P2_P3_InstQueue_reg[11][2]/NET0131  & n26827 ;
  assign n57691 = \P2_P3_InstQueue_reg[8][2]/NET0131  & n26822 ;
  assign n57703 = ~n57690 & ~n57691 ;
  assign n57693 = \P2_P3_InstQueue_reg[9][2]/NET0131  & n26841 ;
  assign n57696 = \P2_P3_InstQueue_reg[13][2]/NET0131  & n26819 ;
  assign n57704 = ~n57693 & ~n57696 ;
  assign n57707 = n57703 & n57704 ;
  assign n57686 = \P2_P3_InstQueue_reg[7][2]/NET0131  & n26815 ;
  assign n57687 = \P2_P3_InstQueue_reg[4][2]/NET0131  & n26831 ;
  assign n57701 = ~n57686 & ~n57687 ;
  assign n57688 = \P2_P3_InstQueue_reg[15][2]/NET0131  & n26829 ;
  assign n57689 = \P2_P3_InstQueue_reg[12][2]/NET0131  & n26833 ;
  assign n57702 = ~n57688 & ~n57689 ;
  assign n57708 = n57701 & n57702 ;
  assign n57712 = n57707 & n57708 ;
  assign n57713 = n57706 & n57712 ;
  assign n57714 = n57711 & n57713 ;
  assign n57715 = n42538 & ~n57714 ;
  assign n57716 = ~n57683 & ~n57715 ;
  assign n57717 = ~n57676 & n57716 ;
  assign n57718 = ~n57679 & n57717 ;
  assign n57719 = n27308 & ~n57718 ;
  assign n57720 = \P2_P3_EAX_reg[18]/NET0131  & ~n42872 ;
  assign n57721 = ~n57719 & ~n57720 ;
  assign n57722 = \P2_P3_EAX_reg[19]/NET0131  & ~n42872 ;
  assign n57755 = n42543 & ~n57678 ;
  assign n57756 = \P2_P3_EAX_reg[19]/NET0131  & ~n57755 ;
  assign n57761 = ~\P2_P3_EAX_reg[19]/NET0131  & n42539 ;
  assign n57762 = n42850 & n57761 ;
  assign n57731 = \P2_P3_InstQueue_reg[1][3]/NET0131  & n26845 ;
  assign n57723 = \P2_P3_InstQueue_reg[4][3]/NET0131  & n26831 ;
  assign n57724 = \P2_P3_InstQueue_reg[13][3]/NET0131  & n26819 ;
  assign n57739 = ~n57723 & ~n57724 ;
  assign n57748 = ~n57731 & n57739 ;
  assign n57733 = \P2_P3_InstQueue_reg[2][3]/NET0131  & n26837 ;
  assign n57734 = \P2_P3_InstQueue_reg[10][3]/NET0131  & n26839 ;
  assign n57749 = ~n57733 & ~n57734 ;
  assign n57750 = n57748 & n57749 ;
  assign n57738 = \P2_P3_InstQueue_reg[15][3]/NET0131  & n26829 ;
  assign n57736 = \P2_P3_InstQueue_reg[11][3]/NET0131  & n26827 ;
  assign n57737 = \P2_P3_InstQueue_reg[6][3]/NET0131  & n26847 ;
  assign n57744 = ~n57736 & ~n57737 ;
  assign n57745 = ~n57738 & n57744 ;
  assign n57729 = \P2_P3_InstQueue_reg[3][3]/NET0131  & n26812 ;
  assign n57730 = \P2_P3_InstQueue_reg[8][3]/NET0131  & n26822 ;
  assign n57742 = ~n57729 & ~n57730 ;
  assign n57732 = \P2_P3_InstQueue_reg[9][3]/NET0131  & n26841 ;
  assign n57735 = \P2_P3_InstQueue_reg[14][3]/NET0131  & n26849 ;
  assign n57743 = ~n57732 & ~n57735 ;
  assign n57746 = n57742 & n57743 ;
  assign n57725 = \P2_P3_InstQueue_reg[5][3]/NET0131  & n26843 ;
  assign n57726 = \P2_P3_InstQueue_reg[0][3]/NET0131  & n26825 ;
  assign n57740 = ~n57725 & ~n57726 ;
  assign n57727 = \P2_P3_InstQueue_reg[7][3]/NET0131  & n26815 ;
  assign n57728 = \P2_P3_InstQueue_reg[12][3]/NET0131  & n26833 ;
  assign n57741 = ~n57727 & ~n57728 ;
  assign n57747 = n57740 & n57741 ;
  assign n57751 = n57746 & n57747 ;
  assign n57752 = n57745 & n57751 ;
  assign n57753 = n57750 & n57752 ;
  assign n57754 = n42538 & ~n57753 ;
  assign n57757 = \P2_buf2_reg[3]/NET0131  & n27122 ;
  assign n57758 = \P2_buf2_reg[19]/NET0131  & n27186 ;
  assign n57759 = ~n57757 & ~n57758 ;
  assign n57760 = n27227 & ~n57759 ;
  assign n57763 = ~n57754 & ~n57760 ;
  assign n57764 = ~n57762 & n57763 ;
  assign n57765 = ~n57756 & n57764 ;
  assign n57766 = n27308 & ~n57765 ;
  assign n57767 = ~n57722 & ~n57766 ;
  assign n57768 = \P2_P3_EAX_reg[20]/NET0131  & ~n42872 ;
  assign n57801 = n42539 & ~n46591 ;
  assign n57802 = ~n42542 & ~n57801 ;
  assign n57803 = \P2_P3_EAX_reg[20]/NET0131  & ~n57802 ;
  assign n57810 = ~\P2_P3_EAX_reg[20]/NET0131  & n42539 ;
  assign n57811 = n46591 & n57810 ;
  assign n57804 = \P2_P3_EAX_reg[20]/NET0131  & ~n27227 ;
  assign n57808 = ~n53434 & ~n57804 ;
  assign n57809 = n27122 & ~n57808 ;
  assign n57778 = \P2_P3_InstQueue_reg[2][4]/NET0131  & n26837 ;
  assign n57769 = \P2_P3_InstQueue_reg[6][4]/NET0131  & n26847 ;
  assign n57770 = \P2_P3_InstQueue_reg[5][4]/NET0131  & n26843 ;
  assign n57785 = ~n57769 & ~n57770 ;
  assign n57794 = ~n57778 & n57785 ;
  assign n57779 = \P2_P3_InstQueue_reg[10][4]/NET0131  & n26839 ;
  assign n57782 = \P2_P3_InstQueue_reg[1][4]/NET0131  & n26845 ;
  assign n57795 = ~n57779 & ~n57782 ;
  assign n57796 = n57794 & n57795 ;
  assign n57784 = \P2_P3_InstQueue_reg[15][4]/NET0131  & n26829 ;
  assign n57781 = \P2_P3_InstQueue_reg[11][4]/NET0131  & n26827 ;
  assign n57783 = \P2_P3_InstQueue_reg[0][4]/NET0131  & n26825 ;
  assign n57790 = ~n57781 & ~n57783 ;
  assign n57791 = ~n57784 & n57790 ;
  assign n57775 = \P2_P3_InstQueue_reg[4][4]/NET0131  & n26831 ;
  assign n57776 = \P2_P3_InstQueue_reg[14][4]/NET0131  & n26849 ;
  assign n57788 = ~n57775 & ~n57776 ;
  assign n57777 = \P2_P3_InstQueue_reg[3][4]/NET0131  & n26812 ;
  assign n57780 = \P2_P3_InstQueue_reg[9][4]/NET0131  & n26841 ;
  assign n57789 = ~n57777 & ~n57780 ;
  assign n57792 = n57788 & n57789 ;
  assign n57771 = \P2_P3_InstQueue_reg[12][4]/NET0131  & n26833 ;
  assign n57772 = \P2_P3_InstQueue_reg[8][4]/NET0131  & n26822 ;
  assign n57786 = ~n57771 & ~n57772 ;
  assign n57773 = \P2_P3_InstQueue_reg[13][4]/NET0131  & n26819 ;
  assign n57774 = \P2_P3_InstQueue_reg[7][4]/NET0131  & n26815 ;
  assign n57787 = ~n57773 & ~n57774 ;
  assign n57793 = n57786 & n57787 ;
  assign n57797 = n57792 & n57793 ;
  assign n57798 = n57791 & n57797 ;
  assign n57799 = n57796 & n57798 ;
  assign n57800 = n42538 & ~n57799 ;
  assign n57805 = \P2_buf2_reg[20]/NET0131  & n27227 ;
  assign n57806 = ~n57804 & ~n57805 ;
  assign n57807 = n27186 & ~n57806 ;
  assign n57812 = ~n57800 & ~n57807 ;
  assign n57813 = ~n57809 & n57812 ;
  assign n57814 = ~n57811 & n57813 ;
  assign n57815 = ~n57803 & n57814 ;
  assign n57816 = n27308 & ~n57815 ;
  assign n57817 = ~n57768 & ~n57816 ;
  assign n57818 = \P2_P3_EAX_reg[21]/NET0131  & ~n42872 ;
  assign n57820 = \P2_P3_EAX_reg[20]/NET0131  & n46591 ;
  assign n57822 = \P2_P3_EAX_reg[21]/NET0131  & n57820 ;
  assign n57821 = ~\P2_P3_EAX_reg[21]/NET0131  & ~n57820 ;
  assign n57823 = n42539 & ~n57821 ;
  assign n57824 = ~n57822 & n57823 ;
  assign n57825 = \P2_P3_EAX_reg[21]/NET0131  & ~n42543 ;
  assign n57858 = \P2_buf2_reg[21]/NET0131  & n46606 ;
  assign n57819 = n46587 & n53314 ;
  assign n57834 = \P2_P3_InstQueue_reg[1][5]/NET0131  & n26845 ;
  assign n57826 = \P2_P3_InstQueue_reg[3][5]/NET0131  & n26812 ;
  assign n57827 = \P2_P3_InstQueue_reg[15][5]/NET0131  & n26829 ;
  assign n57842 = ~n57826 & ~n57827 ;
  assign n57851 = ~n57834 & n57842 ;
  assign n57836 = \P2_P3_InstQueue_reg[2][5]/NET0131  & n26837 ;
  assign n57837 = \P2_P3_InstQueue_reg[10][5]/NET0131  & n26839 ;
  assign n57852 = ~n57836 & ~n57837 ;
  assign n57853 = n57851 & n57852 ;
  assign n57841 = \P2_P3_InstQueue_reg[4][5]/NET0131  & n26831 ;
  assign n57839 = \P2_P3_InstQueue_reg[6][5]/NET0131  & n26847 ;
  assign n57840 = \P2_P3_InstQueue_reg[14][5]/NET0131  & n26849 ;
  assign n57847 = ~n57839 & ~n57840 ;
  assign n57848 = ~n57841 & n57847 ;
  assign n57832 = \P2_P3_InstQueue_reg[13][5]/NET0131  & n26819 ;
  assign n57833 = \P2_P3_InstQueue_reg[0][5]/NET0131  & n26825 ;
  assign n57845 = ~n57832 & ~n57833 ;
  assign n57835 = \P2_P3_InstQueue_reg[9][5]/NET0131  & n26841 ;
  assign n57838 = \P2_P3_InstQueue_reg[11][5]/NET0131  & n26827 ;
  assign n57846 = ~n57835 & ~n57838 ;
  assign n57849 = n57845 & n57846 ;
  assign n57828 = \P2_P3_InstQueue_reg[12][5]/NET0131  & n26833 ;
  assign n57829 = \P2_P3_InstQueue_reg[8][5]/NET0131  & n26822 ;
  assign n57843 = ~n57828 & ~n57829 ;
  assign n57830 = \P2_P3_InstQueue_reg[7][5]/NET0131  & n26815 ;
  assign n57831 = \P2_P3_InstQueue_reg[5][5]/NET0131  & n26843 ;
  assign n57844 = ~n57830 & ~n57831 ;
  assign n57850 = n57843 & n57844 ;
  assign n57854 = n57849 & n57850 ;
  assign n57855 = n57848 & n57854 ;
  assign n57856 = n57853 & n57855 ;
  assign n57857 = n42538 & ~n57856 ;
  assign n57859 = ~n57819 & ~n57857 ;
  assign n57860 = ~n57858 & n57859 ;
  assign n57861 = ~n57825 & n57860 ;
  assign n57862 = ~n57824 & n57861 ;
  assign n57863 = n27308 & ~n57862 ;
  assign n57864 = ~n57818 & ~n57863 ;
  assign n57865 = \P2_P3_EAX_reg[22]/NET0131  & ~n42872 ;
  assign n57867 = \P2_P3_EAX_reg[22]/NET0131  & n57822 ;
  assign n57868 = n42539 & ~n57867 ;
  assign n57869 = ~\P2_P3_EAX_reg[22]/NET0131  & ~n57822 ;
  assign n57870 = n57868 & ~n57869 ;
  assign n57871 = ~n42542 & ~n45740 ;
  assign n57872 = \P2_P3_EAX_reg[22]/NET0131  & ~n57871 ;
  assign n57884 = \P2_P3_InstQueue_reg[1][6]/NET0131  & n26845 ;
  assign n57876 = \P2_P3_InstQueue_reg[5][6]/NET0131  & n26843 ;
  assign n57877 = \P2_P3_InstQueue_reg[3][6]/NET0131  & n26812 ;
  assign n57892 = ~n57876 & ~n57877 ;
  assign n57901 = ~n57884 & n57892 ;
  assign n57886 = \P2_P3_InstQueue_reg[10][6]/NET0131  & n26839 ;
  assign n57887 = \P2_P3_InstQueue_reg[2][6]/NET0131  & n26837 ;
  assign n57902 = ~n57886 & ~n57887 ;
  assign n57903 = n57901 & n57902 ;
  assign n57891 = \P2_P3_InstQueue_reg[7][6]/NET0131  & n26815 ;
  assign n57889 = \P2_P3_InstQueue_reg[8][6]/NET0131  & n26822 ;
  assign n57890 = \P2_P3_InstQueue_reg[11][6]/NET0131  & n26827 ;
  assign n57897 = ~n57889 & ~n57890 ;
  assign n57898 = ~n57891 & n57897 ;
  assign n57882 = \P2_P3_InstQueue_reg[4][6]/NET0131  & n26831 ;
  assign n57883 = \P2_P3_InstQueue_reg[14][6]/NET0131  & n26849 ;
  assign n57895 = ~n57882 & ~n57883 ;
  assign n57885 = \P2_P3_InstQueue_reg[9][6]/NET0131  & n26841 ;
  assign n57888 = \P2_P3_InstQueue_reg[15][6]/NET0131  & n26829 ;
  assign n57896 = ~n57885 & ~n57888 ;
  assign n57899 = n57895 & n57896 ;
  assign n57878 = \P2_P3_InstQueue_reg[0][6]/NET0131  & n26825 ;
  assign n57879 = \P2_P3_InstQueue_reg[6][6]/NET0131  & n26847 ;
  assign n57893 = ~n57878 & ~n57879 ;
  assign n57880 = \P2_P3_InstQueue_reg[12][6]/NET0131  & n26833 ;
  assign n57881 = \P2_P3_InstQueue_reg[13][6]/NET0131  & n26819 ;
  assign n57894 = ~n57880 & ~n57881 ;
  assign n57900 = n57893 & n57894 ;
  assign n57904 = n57899 & n57900 ;
  assign n57905 = n57898 & n57904 ;
  assign n57906 = n57903 & n57905 ;
  assign n57907 = n42538 & ~n57906 ;
  assign n57866 = \P2_buf2_reg[22]/NET0131  & n46606 ;
  assign n57873 = \P2_P3_EAX_reg[22]/NET0131  & ~n27227 ;
  assign n57874 = ~n53333 & ~n57873 ;
  assign n57875 = n27122 & ~n57874 ;
  assign n57908 = ~n57866 & ~n57875 ;
  assign n57909 = ~n57907 & n57908 ;
  assign n57910 = ~n57872 & n57909 ;
  assign n57911 = ~n57870 & n57910 ;
  assign n57912 = n27308 & ~n57911 ;
  assign n57913 = ~n57865 & ~n57912 ;
  assign n57914 = \P2_P3_EAX_reg[23]/NET0131  & ~n42872 ;
  assign n57918 = n42543 & ~n57868 ;
  assign n57919 = \P2_P3_EAX_reg[23]/NET0131  & ~n57918 ;
  assign n57924 = ~\P2_P3_EAX_reg[23]/NET0131  & n42539 ;
  assign n57925 = n57867 & n57924 ;
  assign n57915 = n42575 & n42606 ;
  assign n57916 = ~n42607 & ~n57915 ;
  assign n57917 = n42538 & n57916 ;
  assign n57920 = \P2_buf2_reg[7]/NET0131  & n27122 ;
  assign n57921 = \P2_buf2_reg[23]/NET0131  & n27186 ;
  assign n57922 = ~n57920 & ~n57921 ;
  assign n57923 = n27227 & ~n57922 ;
  assign n57926 = ~n57917 & ~n57923 ;
  assign n57927 = ~n57925 & n57926 ;
  assign n57928 = ~n57919 & n57927 ;
  assign n57929 = n27308 & ~n57928 ;
  assign n57930 = ~n57914 & ~n57929 ;
  assign n57931 = \P2_P3_EAX_reg[24]/NET0131  & ~n42872 ;
  assign n57935 = \P2_P3_EAX_reg[23]/NET0131  & n57867 ;
  assign n57936 = n42539 & ~n57935 ;
  assign n57937 = n42543 & ~n57936 ;
  assign n57938 = \P2_P3_EAX_reg[24]/NET0131  & ~n57937 ;
  assign n57942 = ~\P2_P3_EAX_reg[24]/NET0131  & n42539 ;
  assign n57943 = n57935 & n57942 ;
  assign n57932 = ~n42607 & n42638 ;
  assign n57933 = ~n42639 & ~n57932 ;
  assign n57934 = n42538 & n57933 ;
  assign n57939 = \P2_buf2_reg[24]/NET0131  & n27186 ;
  assign n57940 = ~n49640 & ~n57939 ;
  assign n57941 = n27227 & ~n57940 ;
  assign n57944 = ~n57934 & ~n57941 ;
  assign n57945 = ~n57943 & n57944 ;
  assign n57946 = ~n57938 & n57945 ;
  assign n57947 = n27308 & ~n57946 ;
  assign n57948 = ~n57931 & ~n57947 ;
  assign n57949 = \P2_P3_EAX_reg[28]/NET0131  & ~n42872 ;
  assign n57951 = ~\P2_P3_EAX_reg[28]/NET0131  & ~n46595 ;
  assign n57952 = n42539 & ~n46596 ;
  assign n57953 = ~n57951 & n57952 ;
  assign n57954 = \P2_P3_EAX_reg[28]/NET0131  & ~n48259 ;
  assign n57955 = ~n42735 & n42766 ;
  assign n57956 = ~n42767 & ~n57955 ;
  assign n57957 = n42538 & n57956 ;
  assign n57950 = n46587 & n47755 ;
  assign n57959 = ~\P2_buf2_reg[28]/NET0131  & n27227 ;
  assign n57958 = ~\P2_P3_EAX_reg[28]/NET0131  & ~n27227 ;
  assign n57960 = n27186 & ~n57958 ;
  assign n57961 = ~n57959 & n57960 ;
  assign n57962 = ~n57950 & ~n57961 ;
  assign n57963 = ~n57957 & n57962 ;
  assign n57964 = ~n57954 & n57963 ;
  assign n57965 = ~n57953 & n57964 ;
  assign n57966 = n27308 & ~n57965 ;
  assign n57967 = ~n57949 & ~n57966 ;
  assign n57970 = ~\P2_P3_EBX_reg[25]/NET0131  & ~n46641 ;
  assign n57971 = n27133 & ~n46642 ;
  assign n57972 = ~n57970 & n57971 ;
  assign n57968 = \P2_P3_EBX_reg[25]/NET0131  & n46615 ;
  assign n57969 = n46614 & n53275 ;
  assign n57973 = ~n57968 & ~n57969 ;
  assign n57974 = ~n57972 & n57973 ;
  assign n57975 = n27308 & ~n57974 ;
  assign n57976 = \P2_P3_EBX_reg[25]/NET0131  & ~n42872 ;
  assign n57977 = ~n57975 & ~n57976 ;
  assign n57978 = \P1_P2_EAX_reg[16]/NET0131  & ~n43212 ;
  assign n58011 = \P1_P2_EAX_reg[16]/NET0131  & ~n43168 ;
  assign n58012 = ~\P1_P2_EAX_reg[16]/NET0131  & ~n43185 ;
  assign n58013 = n43164 & ~n43186 ;
  assign n58014 = ~n58012 & n58013 ;
  assign n58015 = n25773 & n46761 ;
  assign n58016 = ~\P1_P2_EAX_reg[16]/NET0131  & ~n25773 ;
  assign n58017 = ~n58015 & ~n58016 ;
  assign n58018 = n25774 & n58017 ;
  assign n57990 = \P1_P2_InstQueue_reg[9][0]/NET0131  & n25453 ;
  assign n57983 = \P1_P2_InstQueue_reg[10][0]/NET0131  & n25435 ;
  assign n57979 = \P1_P2_InstQueue_reg[4][0]/NET0131  & n25428 ;
  assign n57980 = \P1_P2_InstQueue_reg[12][0]/NET0131  & n25457 ;
  assign n57995 = ~n57979 & ~n57980 ;
  assign n58005 = ~n57983 & n57995 ;
  assign n58006 = ~n57990 & n58005 ;
  assign n57991 = \P1_P2_InstQueue_reg[11][0]/NET0131  & n25455 ;
  assign n57992 = \P1_P2_InstQueue_reg[5][0]/NET0131  & n25444 ;
  assign n58000 = ~n57991 & ~n57992 ;
  assign n57993 = \P1_P2_InstQueue_reg[0][0]/NET0131  & n25442 ;
  assign n57994 = \P1_P2_InstQueue_reg[3][0]/NET0131  & n25425 ;
  assign n58001 = ~n57993 & ~n57994 ;
  assign n58002 = n58000 & n58001 ;
  assign n57986 = \P1_P2_InstQueue_reg[15][0]/NET0131  & n25422 ;
  assign n57987 = \P1_P2_InstQueue_reg[14][0]/NET0131  & n25459 ;
  assign n57998 = ~n57986 & ~n57987 ;
  assign n57988 = \P1_P2_InstQueue_reg[2][0]/NET0131  & n25446 ;
  assign n57989 = \P1_P2_InstQueue_reg[8][0]/NET0131  & n25449 ;
  assign n57999 = ~n57988 & ~n57989 ;
  assign n58003 = n57998 & n57999 ;
  assign n57981 = \P1_P2_InstQueue_reg[7][0]/NET0131  & n25461 ;
  assign n57982 = \P1_P2_InstQueue_reg[1][0]/NET0131  & n25431 ;
  assign n57996 = ~n57981 & ~n57982 ;
  assign n57984 = \P1_P2_InstQueue_reg[13][0]/NET0131  & n25440 ;
  assign n57985 = \P1_P2_InstQueue_reg[6][0]/NET0131  & n25437 ;
  assign n57997 = ~n57984 & ~n57985 ;
  assign n58004 = n57996 & n57997 ;
  assign n58007 = n58003 & n58004 ;
  assign n58008 = n58002 & n58007 ;
  assign n58009 = n58006 & n58008 ;
  assign n58010 = n42875 & ~n58009 ;
  assign n58019 = ~n56902 & ~n58010 ;
  assign n58020 = ~n58018 & n58019 ;
  assign n58021 = ~n58014 & n58020 ;
  assign n58022 = ~n58011 & n58021 ;
  assign n58023 = n25918 & ~n58022 ;
  assign n58024 = ~n57978 & ~n58023 ;
  assign n58025 = \P1_P2_EAX_reg[17]/NET0131  & ~n43212 ;
  assign n58058 = ~n25775 & ~n43167 ;
  assign n58059 = ~n58013 & n58058 ;
  assign n58060 = \P1_P2_EAX_reg[17]/NET0131  & ~n58059 ;
  assign n58065 = ~\P1_P2_EAX_reg[17]/NET0131  & n43164 ;
  assign n58066 = n43186 & n58065 ;
  assign n58064 = n34212 & ~n40758 ;
  assign n58037 = \P1_P2_InstQueue_reg[9][1]/NET0131  & n25453 ;
  assign n58030 = \P1_P2_InstQueue_reg[10][1]/NET0131  & n25435 ;
  assign n58026 = \P1_P2_InstQueue_reg[5][1]/NET0131  & n25444 ;
  assign n58027 = \P1_P2_InstQueue_reg[8][1]/NET0131  & n25449 ;
  assign n58042 = ~n58026 & ~n58027 ;
  assign n58052 = ~n58030 & n58042 ;
  assign n58053 = ~n58037 & n58052 ;
  assign n58038 = \P1_P2_InstQueue_reg[4][1]/NET0131  & n25428 ;
  assign n58039 = \P1_P2_InstQueue_reg[11][1]/NET0131  & n25455 ;
  assign n58047 = ~n58038 & ~n58039 ;
  assign n58040 = \P1_P2_InstQueue_reg[6][1]/NET0131  & n25437 ;
  assign n58041 = \P1_P2_InstQueue_reg[13][1]/NET0131  & n25440 ;
  assign n58048 = ~n58040 & ~n58041 ;
  assign n58049 = n58047 & n58048 ;
  assign n58033 = \P1_P2_InstQueue_reg[3][1]/NET0131  & n25425 ;
  assign n58034 = \P1_P2_InstQueue_reg[15][1]/NET0131  & n25422 ;
  assign n58045 = ~n58033 & ~n58034 ;
  assign n58035 = \P1_P2_InstQueue_reg[2][1]/NET0131  & n25446 ;
  assign n58036 = \P1_P2_InstQueue_reg[12][1]/NET0131  & n25457 ;
  assign n58046 = ~n58035 & ~n58036 ;
  assign n58050 = n58045 & n58046 ;
  assign n58028 = \P1_P2_InstQueue_reg[0][1]/NET0131  & n25442 ;
  assign n58029 = \P1_P2_InstQueue_reg[1][1]/NET0131  & n25431 ;
  assign n58043 = ~n58028 & ~n58029 ;
  assign n58031 = \P1_P2_InstQueue_reg[7][1]/NET0131  & n25461 ;
  assign n58032 = \P1_P2_InstQueue_reg[14][1]/NET0131  & n25459 ;
  assign n58044 = ~n58031 & ~n58032 ;
  assign n58051 = n58043 & n58044 ;
  assign n58054 = n58050 & n58051 ;
  assign n58055 = n58049 & n58054 ;
  assign n58056 = n58053 & n58055 ;
  assign n58057 = n42875 & ~n58056 ;
  assign n58061 = \P1_P2_EAX_reg[17]/NET0131  & ~n25773 ;
  assign n58062 = ~n53356 & ~n58061 ;
  assign n58063 = n25776 & ~n58062 ;
  assign n58067 = ~n58057 & ~n58063 ;
  assign n58068 = ~n58064 & n58067 ;
  assign n58069 = ~n58066 & n58068 ;
  assign n58070 = ~n58060 & n58069 ;
  assign n58071 = n25918 & ~n58070 ;
  assign n58072 = ~n58025 & ~n58071 ;
  assign n58074 = ~\P1_P2_EAX_reg[18]/NET0131  & ~n43187 ;
  assign n58075 = n43164 & ~n43188 ;
  assign n58076 = ~n58074 & n58075 ;
  assign n58073 = \P1_P2_EAX_reg[18]/NET0131  & ~n43169 ;
  assign n58077 = n25774 & ~n35975 ;
  assign n58078 = ~n56951 & ~n58077 ;
  assign n58079 = n25773 & ~n58078 ;
  assign n58091 = \P1_P2_InstQueue_reg[9][2]/NET0131  & n25453 ;
  assign n58084 = \P1_P2_InstQueue_reg[10][2]/NET0131  & n25435 ;
  assign n58080 = \P1_P2_InstQueue_reg[15][2]/NET0131  & n25422 ;
  assign n58081 = \P1_P2_InstQueue_reg[3][2]/NET0131  & n25425 ;
  assign n58096 = ~n58080 & ~n58081 ;
  assign n58106 = ~n58084 & n58096 ;
  assign n58107 = ~n58091 & n58106 ;
  assign n58092 = \P1_P2_InstQueue_reg[8][2]/NET0131  & n25449 ;
  assign n58093 = \P1_P2_InstQueue_reg[7][2]/NET0131  & n25461 ;
  assign n58101 = ~n58092 & ~n58093 ;
  assign n58094 = \P1_P2_InstQueue_reg[12][2]/NET0131  & n25457 ;
  assign n58095 = \P1_P2_InstQueue_reg[5][2]/NET0131  & n25444 ;
  assign n58102 = ~n58094 & ~n58095 ;
  assign n58103 = n58101 & n58102 ;
  assign n58087 = \P1_P2_InstQueue_reg[14][2]/NET0131  & n25459 ;
  assign n58088 = \P1_P2_InstQueue_reg[0][2]/NET0131  & n25442 ;
  assign n58099 = ~n58087 & ~n58088 ;
  assign n58089 = \P1_P2_InstQueue_reg[2][2]/NET0131  & n25446 ;
  assign n58090 = \P1_P2_InstQueue_reg[13][2]/NET0131  & n25440 ;
  assign n58100 = ~n58089 & ~n58090 ;
  assign n58104 = n58099 & n58100 ;
  assign n58082 = \P1_P2_InstQueue_reg[4][2]/NET0131  & n25428 ;
  assign n58083 = \P1_P2_InstQueue_reg[1][2]/NET0131  & n25431 ;
  assign n58097 = ~n58082 & ~n58083 ;
  assign n58085 = \P1_P2_InstQueue_reg[6][2]/NET0131  & n25437 ;
  assign n58086 = \P1_P2_InstQueue_reg[11][2]/NET0131  & n25455 ;
  assign n58098 = ~n58085 & ~n58086 ;
  assign n58105 = n58097 & n58098 ;
  assign n58108 = n58104 & n58105 ;
  assign n58109 = n58103 & n58108 ;
  assign n58110 = n58107 & n58109 ;
  assign n58111 = n42875 & ~n58110 ;
  assign n58112 = ~n58079 & ~n58111 ;
  assign n58113 = ~n58073 & n58112 ;
  assign n58114 = ~n58076 & n58113 ;
  assign n58115 = n25918 & ~n58114 ;
  assign n58116 = \P1_P2_EAX_reg[18]/NET0131  & ~n43212 ;
  assign n58117 = ~n58115 & ~n58116 ;
  assign n58118 = \P1_P2_EAX_reg[19]/NET0131  & ~n43212 ;
  assign n58151 = n43169 & ~n58075 ;
  assign n58152 = \P1_P2_EAX_reg[19]/NET0131  & ~n58151 ;
  assign n58156 = ~\P1_P2_EAX_reg[19]/NET0131  & n43164 ;
  assign n58157 = n43188 & n58156 ;
  assign n58130 = \P1_P2_InstQueue_reg[9][3]/NET0131  & n25453 ;
  assign n58123 = \P1_P2_InstQueue_reg[10][3]/NET0131  & n25435 ;
  assign n58119 = \P1_P2_InstQueue_reg[7][3]/NET0131  & n25461 ;
  assign n58120 = \P1_P2_InstQueue_reg[11][3]/NET0131  & n25455 ;
  assign n58135 = ~n58119 & ~n58120 ;
  assign n58145 = ~n58123 & n58135 ;
  assign n58146 = ~n58130 & n58145 ;
  assign n58131 = \P1_P2_InstQueue_reg[12][3]/NET0131  & n25457 ;
  assign n58132 = \P1_P2_InstQueue_reg[13][3]/NET0131  & n25440 ;
  assign n58140 = ~n58131 & ~n58132 ;
  assign n58133 = \P1_P2_InstQueue_reg[6][3]/NET0131  & n25437 ;
  assign n58134 = \P1_P2_InstQueue_reg[3][3]/NET0131  & n25425 ;
  assign n58141 = ~n58133 & ~n58134 ;
  assign n58142 = n58140 & n58141 ;
  assign n58126 = \P1_P2_InstQueue_reg[15][3]/NET0131  & n25422 ;
  assign n58127 = \P1_P2_InstQueue_reg[8][3]/NET0131  & n25449 ;
  assign n58138 = ~n58126 & ~n58127 ;
  assign n58128 = \P1_P2_InstQueue_reg[2][3]/NET0131  & n25446 ;
  assign n58129 = \P1_P2_InstQueue_reg[4][3]/NET0131  & n25428 ;
  assign n58139 = ~n58128 & ~n58129 ;
  assign n58143 = n58138 & n58139 ;
  assign n58121 = \P1_P2_InstQueue_reg[0][3]/NET0131  & n25442 ;
  assign n58122 = \P1_P2_InstQueue_reg[1][3]/NET0131  & n25431 ;
  assign n58136 = ~n58121 & ~n58122 ;
  assign n58124 = \P1_P2_InstQueue_reg[14][3]/NET0131  & n25459 ;
  assign n58125 = \P1_P2_InstQueue_reg[5][3]/NET0131  & n25444 ;
  assign n58137 = ~n58124 & ~n58125 ;
  assign n58144 = n58136 & n58137 ;
  assign n58147 = n58143 & n58144 ;
  assign n58148 = n58142 & n58147 ;
  assign n58149 = n58146 & n58148 ;
  assign n58150 = n42875 & ~n58149 ;
  assign n58153 = n25774 & ~n29844 ;
  assign n58154 = ~n56958 & ~n58153 ;
  assign n58155 = n25773 & ~n58154 ;
  assign n58158 = ~n58150 & ~n58155 ;
  assign n58159 = ~n58157 & n58158 ;
  assign n58160 = ~n58152 & n58159 ;
  assign n58161 = n25918 & ~n58160 ;
  assign n58162 = ~n58118 & ~n58161 ;
  assign n58164 = ~\P1_P2_EAX_reg[20]/NET0131  & ~n43189 ;
  assign n58165 = n43164 & ~n43190 ;
  assign n58166 = ~n58164 & n58165 ;
  assign n58163 = \P1_P2_EAX_reg[20]/NET0131  & ~n43169 ;
  assign n58167 = n25776 & ~n27937 ;
  assign n58168 = n25774 & ~n27955 ;
  assign n58169 = ~n58167 & ~n58168 ;
  assign n58170 = n25773 & ~n58169 ;
  assign n58182 = \P1_P2_InstQueue_reg[9][4]/NET0131  & n25453 ;
  assign n58175 = \P1_P2_InstQueue_reg[10][4]/NET0131  & n25435 ;
  assign n58171 = \P1_P2_InstQueue_reg[7][4]/NET0131  & n25461 ;
  assign n58172 = \P1_P2_InstQueue_reg[11][4]/NET0131  & n25455 ;
  assign n58187 = ~n58171 & ~n58172 ;
  assign n58197 = ~n58175 & n58187 ;
  assign n58198 = ~n58182 & n58197 ;
  assign n58183 = \P1_P2_InstQueue_reg[12][4]/NET0131  & n25457 ;
  assign n58184 = \P1_P2_InstQueue_reg[15][4]/NET0131  & n25422 ;
  assign n58192 = ~n58183 & ~n58184 ;
  assign n58185 = \P1_P2_InstQueue_reg[6][4]/NET0131  & n25437 ;
  assign n58186 = \P1_P2_InstQueue_reg[3][4]/NET0131  & n25425 ;
  assign n58193 = ~n58185 & ~n58186 ;
  assign n58194 = n58192 & n58193 ;
  assign n58178 = \P1_P2_InstQueue_reg[13][4]/NET0131  & n25440 ;
  assign n58179 = \P1_P2_InstQueue_reg[8][4]/NET0131  & n25449 ;
  assign n58190 = ~n58178 & ~n58179 ;
  assign n58180 = \P1_P2_InstQueue_reg[2][4]/NET0131  & n25446 ;
  assign n58181 = \P1_P2_InstQueue_reg[4][4]/NET0131  & n25428 ;
  assign n58191 = ~n58180 & ~n58181 ;
  assign n58195 = n58190 & n58191 ;
  assign n58173 = \P1_P2_InstQueue_reg[0][4]/NET0131  & n25442 ;
  assign n58174 = \P1_P2_InstQueue_reg[1][4]/NET0131  & n25431 ;
  assign n58188 = ~n58173 & ~n58174 ;
  assign n58176 = \P1_P2_InstQueue_reg[14][4]/NET0131  & n25459 ;
  assign n58177 = \P1_P2_InstQueue_reg[5][4]/NET0131  & n25444 ;
  assign n58189 = ~n58176 & ~n58177 ;
  assign n58196 = n58188 & n58189 ;
  assign n58199 = n58195 & n58196 ;
  assign n58200 = n58194 & n58199 ;
  assign n58201 = n58198 & n58200 ;
  assign n58202 = n42875 & ~n58201 ;
  assign n58203 = ~n58170 & ~n58202 ;
  assign n58204 = ~n58163 & n58203 ;
  assign n58205 = ~n58166 & n58204 ;
  assign n58206 = n25918 & ~n58205 ;
  assign n58207 = \P1_P2_EAX_reg[20]/NET0131  & ~n43212 ;
  assign n58208 = ~n58206 & ~n58207 ;
  assign n58209 = \P1_P2_EAX_reg[21]/NET0131  & ~n43212 ;
  assign n58211 = ~\P1_P2_EAX_reg[21]/NET0131  & ~n43190 ;
  assign n58212 = n43164 & ~n43191 ;
  assign n58213 = ~n58211 & n58212 ;
  assign n58210 = \P1_P2_EAX_reg[21]/NET0131  & ~n43169 ;
  assign n58246 = ~n29872 & n34212 ;
  assign n58225 = \P1_P2_InstQueue_reg[9][5]/NET0131  & n25453 ;
  assign n58218 = \P1_P2_InstQueue_reg[10][5]/NET0131  & n25435 ;
  assign n58214 = \P1_P2_InstQueue_reg[12][5]/NET0131  & n25457 ;
  assign n58215 = \P1_P2_InstQueue_reg[8][5]/NET0131  & n25449 ;
  assign n58230 = ~n58214 & ~n58215 ;
  assign n58240 = ~n58218 & n58230 ;
  assign n58241 = ~n58225 & n58240 ;
  assign n58226 = \P1_P2_InstQueue_reg[15][5]/NET0131  & n25422 ;
  assign n58227 = \P1_P2_InstQueue_reg[5][5]/NET0131  & n25444 ;
  assign n58235 = ~n58226 & ~n58227 ;
  assign n58228 = \P1_P2_InstQueue_reg[0][5]/NET0131  & n25442 ;
  assign n58229 = \P1_P2_InstQueue_reg[3][5]/NET0131  & n25425 ;
  assign n58236 = ~n58228 & ~n58229 ;
  assign n58237 = n58235 & n58236 ;
  assign n58221 = \P1_P2_InstQueue_reg[14][5]/NET0131  & n25459 ;
  assign n58222 = \P1_P2_InstQueue_reg[13][5]/NET0131  & n25440 ;
  assign n58233 = ~n58221 & ~n58222 ;
  assign n58223 = \P1_P2_InstQueue_reg[2][5]/NET0131  & n25446 ;
  assign n58224 = \P1_P2_InstQueue_reg[4][5]/NET0131  & n25428 ;
  assign n58234 = ~n58223 & ~n58224 ;
  assign n58238 = n58233 & n58234 ;
  assign n58216 = \P1_P2_InstQueue_reg[11][5]/NET0131  & n25455 ;
  assign n58217 = \P1_P2_InstQueue_reg[1][5]/NET0131  & n25431 ;
  assign n58231 = ~n58216 & ~n58217 ;
  assign n58219 = \P1_P2_InstQueue_reg[6][5]/NET0131  & n25437 ;
  assign n58220 = \P1_P2_InstQueue_reg[7][5]/NET0131  & n25461 ;
  assign n58232 = ~n58219 & ~n58220 ;
  assign n58239 = n58231 & n58232 ;
  assign n58242 = n58238 & n58239 ;
  assign n58243 = n58237 & n58242 ;
  assign n58244 = n58241 & n58243 ;
  assign n58245 = n42875 & ~n58244 ;
  assign n58247 = ~n56969 & ~n58245 ;
  assign n58248 = ~n58246 & n58247 ;
  assign n58249 = ~n58210 & n58248 ;
  assign n58250 = ~n58213 & n58249 ;
  assign n58251 = n25918 & ~n58250 ;
  assign n58252 = ~n58209 & ~n58251 ;
  assign n58254 = ~\P1_P2_EAX_reg[22]/NET0131  & ~n43191 ;
  assign n58255 = n43164 & ~n43192 ;
  assign n58256 = ~n58254 & n58255 ;
  assign n58253 = \P1_P2_EAX_reg[22]/NET0131  & ~n43169 ;
  assign n58289 = n34212 & ~n34461 ;
  assign n58268 = \P1_P2_InstQueue_reg[9][6]/NET0131  & n25453 ;
  assign n58261 = \P1_P2_InstQueue_reg[10][6]/NET0131  & n25435 ;
  assign n58257 = \P1_P2_InstQueue_reg[12][6]/NET0131  & n25457 ;
  assign n58258 = \P1_P2_InstQueue_reg[6][6]/NET0131  & n25437 ;
  assign n58273 = ~n58257 & ~n58258 ;
  assign n58283 = ~n58261 & n58273 ;
  assign n58284 = ~n58268 & n58283 ;
  assign n58269 = \P1_P2_InstQueue_reg[3][6]/NET0131  & n25425 ;
  assign n58270 = \P1_P2_InstQueue_reg[5][6]/NET0131  & n25444 ;
  assign n58278 = ~n58269 & ~n58270 ;
  assign n58271 = \P1_P2_InstQueue_reg[4][6]/NET0131  & n25428 ;
  assign n58272 = \P1_P2_InstQueue_reg[7][6]/NET0131  & n25461 ;
  assign n58279 = ~n58271 & ~n58272 ;
  assign n58280 = n58278 & n58279 ;
  assign n58264 = \P1_P2_InstQueue_reg[13][6]/NET0131  & n25440 ;
  assign n58265 = \P1_P2_InstQueue_reg[8][6]/NET0131  & n25449 ;
  assign n58276 = ~n58264 & ~n58265 ;
  assign n58266 = \P1_P2_InstQueue_reg[2][6]/NET0131  & n25446 ;
  assign n58267 = \P1_P2_InstQueue_reg[0][6]/NET0131  & n25442 ;
  assign n58277 = ~n58266 & ~n58267 ;
  assign n58281 = n58276 & n58277 ;
  assign n58259 = \P1_P2_InstQueue_reg[15][6]/NET0131  & n25422 ;
  assign n58260 = \P1_P2_InstQueue_reg[1][6]/NET0131  & n25431 ;
  assign n58274 = ~n58259 & ~n58260 ;
  assign n58262 = \P1_P2_InstQueue_reg[14][6]/NET0131  & n25459 ;
  assign n58263 = \P1_P2_InstQueue_reg[11][6]/NET0131  & n25455 ;
  assign n58275 = ~n58262 & ~n58263 ;
  assign n58282 = n58274 & n58275 ;
  assign n58285 = n58281 & n58282 ;
  assign n58286 = n58280 & n58285 ;
  assign n58287 = n58284 & n58286 ;
  assign n58288 = n42875 & ~n58287 ;
  assign n58290 = ~n56976 & ~n58288 ;
  assign n58291 = ~n58289 & n58290 ;
  assign n58292 = ~n58253 & n58291 ;
  assign n58293 = ~n58256 & n58292 ;
  assign n58294 = n25918 & ~n58293 ;
  assign n58295 = \P1_P2_EAX_reg[22]/NET0131  & ~n43212 ;
  assign n58296 = ~n58294 & ~n58295 ;
  assign n58297 = \P1_P2_EAX_reg[23]/NET0131  & ~n43212 ;
  assign n58299 = ~\P1_P2_EAX_reg[23]/NET0131  & ~n43192 ;
  assign n58300 = n43164 & ~n43193 ;
  assign n58301 = ~n58299 & n58300 ;
  assign n58298 = \P1_P2_EAX_reg[23]/NET0131  & ~n43169 ;
  assign n58302 = n25774 & ~n28939 ;
  assign n58303 = ~n56982 & ~n58302 ;
  assign n58304 = n25773 & ~n58303 ;
  assign n58305 = n42906 & n42937 ;
  assign n58306 = ~n42938 & ~n58305 ;
  assign n58307 = n42875 & n58306 ;
  assign n58308 = ~n58304 & ~n58307 ;
  assign n58309 = ~n58298 & n58308 ;
  assign n58310 = ~n58301 & n58309 ;
  assign n58311 = n25918 & ~n58310 ;
  assign n58312 = ~n58297 & ~n58311 ;
  assign n58313 = ~n27297 & n27308 ;
  assign n58314 = \P2_P3_More_reg/NET0131  & ~n42872 ;
  assign n58315 = ~n58313 & ~n58314 ;
  assign n58317 = ~\P1_P2_EAX_reg[24]/NET0131  & ~n43193 ;
  assign n58318 = n43164 & ~n43194 ;
  assign n58319 = ~n58317 & n58318 ;
  assign n58316 = \P1_P2_EAX_reg[24]/NET0131  & ~n43169 ;
  assign n58320 = n25774 & ~n46757 ;
  assign n58321 = ~n48660 & ~n58320 ;
  assign n58322 = n25773 & ~n58321 ;
  assign n58323 = ~n42938 & n42969 ;
  assign n58324 = ~n42970 & ~n58323 ;
  assign n58325 = n42875 & n58324 ;
  assign n58326 = ~n58322 & ~n58325 ;
  assign n58327 = ~n58316 & n58326 ;
  assign n58328 = ~n58319 & n58327 ;
  assign n58329 = n25918 & ~n58328 ;
  assign n58330 = \P1_P2_EAX_reg[24]/NET0131  & ~n43212 ;
  assign n58331 = ~n58329 & ~n58330 ;
  assign n58332 = \P1_P2_EAX_reg[28]/NET0131  & ~n43212 ;
  assign n58333 = ~n43167 & ~n44811 ;
  assign n58334 = \P1_P2_EAX_reg[28]/NET0131  & ~n58333 ;
  assign n58344 = ~\P1_P2_EAX_reg[28]/NET0131  & n43164 ;
  assign n58345 = n43197 & n58344 ;
  assign n58338 = ~n43066 & n43097 ;
  assign n58339 = ~n43098 & ~n58338 ;
  assign n58340 = n42875 & n58339 ;
  assign n58335 = \P1_P2_EAX_reg[28]/NET0131  & ~n25773 ;
  assign n58336 = ~n49531 & ~n58335 ;
  assign n58337 = n25776 & ~n58336 ;
  assign n58341 = n25773 & ~n27948 ;
  assign n58342 = ~n58335 & ~n58341 ;
  assign n58343 = n25774 & ~n58342 ;
  assign n58346 = ~n58337 & ~n58343 ;
  assign n58347 = ~n58340 & n58346 ;
  assign n58348 = ~n58345 & n58347 ;
  assign n58349 = ~n58334 & n58348 ;
  assign n58350 = n25918 & ~n58349 ;
  assign n58351 = ~n58332 & ~n58350 ;
  assign n58352 = \P2_P3_uWord_reg[11]/NET0131  & ~n47752 ;
  assign n58353 = n27122 & n44800 ;
  assign n58354 = ~n56847 & ~n58353 ;
  assign n58355 = n27308 & ~n58354 ;
  assign n58356 = ~n58352 & ~n58355 ;
  assign n58359 = ~\P1_P2_EBX_reg[25]/NET0131  & ~n46721 ;
  assign n58360 = n25803 & ~n46722 ;
  assign n58361 = ~n58359 & n58360 ;
  assign n58357 = \P1_P2_EBX_reg[25]/NET0131  & n46695 ;
  assign n58358 = n46694 & n53373 ;
  assign n58362 = ~n58357 & ~n58358 ;
  assign n58363 = ~n58361 & n58362 ;
  assign n58364 = n25918 & ~n58363 ;
  assign n58365 = \P1_P2_EBX_reg[25]/NET0131  & ~n43212 ;
  assign n58366 = ~n58364 & ~n58365 ;
  assign n58370 = n25918 & ~n39340 ;
  assign n58371 = ~n27607 & n43211 ;
  assign n58372 = ~n58370 & n58371 ;
  assign n58373 = \P1_P2_PhyAddrPointer_reg[0]/NET0131  & ~n58372 ;
  assign n58367 = n25701 & n45964 ;
  assign n58368 = ~n45967 & ~n58367 ;
  assign n58369 = n25918 & ~n58368 ;
  assign n58374 = ~n45955 & ~n58369 ;
  assign n58375 = ~n58373 & n58374 ;
  assign n58379 = n11612 & n36678 ;
  assign n58380 = n11622 & ~n58379 ;
  assign n58381 = n11611 & ~n11615 ;
  assign n58382 = ~n11624 & ~n58381 ;
  assign n58383 = ~n58380 & n58382 ;
  assign n58384 = \P2_P1_PhyAddrPointer_reg[0]/NET0131  & ~n58383 ;
  assign n58376 = n25945 & n45259 ;
  assign n58377 = ~n45257 & ~n58376 ;
  assign n58378 = n11623 & ~n58377 ;
  assign n58385 = ~n45253 & ~n58378 ;
  assign n58386 = ~n58384 & n58385 ;
  assign n58390 = n8355 & ~n41658 ;
  assign n58391 = n15323 & ~n26113 ;
  assign n58392 = n48477 & n58391 ;
  assign n58393 = ~n58390 & n58392 ;
  assign n58394 = \P1_P1_PhyAddrPointer_reg[0]/NET0131  & ~n58393 ;
  assign n58387 = n26126 & n45677 ;
  assign n58388 = ~n45684 & ~n58387 ;
  assign n58389 = n8355 & ~n58388 ;
  assign n58395 = ~n45672 & ~n58389 ;
  assign n58396 = ~n58394 & n58395 ;
  assign n58400 = n26792 & ~n41873 ;
  assign n58401 = ~n26794 & n45043 ;
  assign n58402 = n54098 & n58401 ;
  assign n58403 = ~n58400 & n58402 ;
  assign n58404 = \P2_P2_PhyAddrPointer_reg[0]/NET0131  & ~n58403 ;
  assign n58397 = n26621 & n45474 ;
  assign n58398 = ~n45482 & ~n58397 ;
  assign n58399 = n26792 & ~n58398 ;
  assign n58405 = ~n45470 & ~n58399 ;
  assign n58406 = ~n58404 & n58405 ;
  assign n58409 = n8955 & n49732 ;
  assign n58408 = ~\P1_P3_InstQueue_reg[0][3]/NET0131  & ~n49732 ;
  assign n58410 = n10046 & ~n58408 ;
  assign n58411 = ~n58409 & n58410 ;
  assign n58407 = \P1_P3_InstQueue_reg[0][3]/NET0131  & ~n49750 ;
  assign n58412 = \P1_buf2_reg[27]/NET0131  & n49739 ;
  assign n58413 = \P1_buf2_reg[19]/NET0131  & ~n49739 ;
  assign n58414 = n49742 & n58413 ;
  assign n58415 = ~n58412 & ~n58414 ;
  assign n58416 = n11698 & ~n58415 ;
  assign n58417 = \P1_buf2_reg[3]/NET0131  & n49760 ;
  assign n58418 = ~n58416 & ~n58417 ;
  assign n58419 = ~n58407 & n58418 ;
  assign n58420 = ~n58411 & n58419 ;
  assign n58423 = n8828 & n49732 ;
  assign n58422 = ~\P1_P3_InstQueue_reg[0][6]/NET0131  & ~n49732 ;
  assign n58424 = n10046 & ~n58422 ;
  assign n58425 = ~n58423 & n58424 ;
  assign n58421 = \P1_P3_InstQueue_reg[0][6]/NET0131  & ~n49750 ;
  assign n58426 = \P1_buf2_reg[30]/NET0131  & n49739 ;
  assign n58427 = \P1_buf2_reg[22]/NET0131  & ~n49739 ;
  assign n58428 = n49742 & n58427 ;
  assign n58429 = ~n58426 & ~n58428 ;
  assign n58430 = n11698 & ~n58429 ;
  assign n58431 = \P1_buf2_reg[6]/NET0131  & n49760 ;
  assign n58432 = ~n58430 & ~n58431 ;
  assign n58433 = ~n58421 & n58432 ;
  assign n58434 = ~n58425 & n58433 ;
  assign n58437 = n8955 & n49766 ;
  assign n58436 = ~\P1_P3_InstQueue_reg[10][3]/NET0131  & ~n49766 ;
  assign n58438 = n10046 & ~n58436 ;
  assign n58439 = ~n58437 & n58438 ;
  assign n58435 = \P1_P3_InstQueue_reg[10][3]/NET0131  & ~n49776 ;
  assign n58440 = \P1_buf2_reg[27]/NET0131  & n49770 ;
  assign n58441 = \P1_buf2_reg[19]/NET0131  & n49771 ;
  assign n58442 = ~n58440 & ~n58441 ;
  assign n58443 = n11698 & ~n58442 ;
  assign n58444 = \P1_buf2_reg[3]/NET0131  & n49786 ;
  assign n58445 = ~n58443 & ~n58444 ;
  assign n58446 = ~n58435 & n58445 ;
  assign n58447 = ~n58439 & n58446 ;
  assign n58450 = n8828 & n49766 ;
  assign n58449 = ~\P1_P3_InstQueue_reg[10][6]/NET0131  & ~n49766 ;
  assign n58451 = n10046 & ~n58449 ;
  assign n58452 = ~n58450 & n58451 ;
  assign n58448 = \P1_P3_InstQueue_reg[10][6]/NET0131  & ~n49776 ;
  assign n58453 = \P1_buf2_reg[30]/NET0131  & n49770 ;
  assign n58454 = \P1_buf2_reg[22]/NET0131  & n49771 ;
  assign n58455 = ~n58453 & ~n58454 ;
  assign n58456 = n11698 & ~n58455 ;
  assign n58457 = \P1_buf2_reg[6]/NET0131  & n49786 ;
  assign n58458 = ~n58456 & ~n58457 ;
  assign n58459 = ~n58448 & n58458 ;
  assign n58460 = ~n58452 & n58459 ;
  assign n58463 = n8955 & n49792 ;
  assign n58462 = ~\P1_P3_InstQueue_reg[11][3]/NET0131  & ~n49792 ;
  assign n58464 = n10046 & ~n58462 ;
  assign n58465 = ~n58463 & n58464 ;
  assign n58461 = \P1_P3_InstQueue_reg[11][3]/NET0131  & ~n49798 ;
  assign n58466 = \P1_buf2_reg[27]/NET0131  & n49771 ;
  assign n58467 = \P1_buf2_reg[19]/NET0131  & n49768 ;
  assign n58468 = ~n58466 & ~n58467 ;
  assign n58469 = n11698 & ~n58468 ;
  assign n58470 = \P1_buf2_reg[3]/NET0131  & n49808 ;
  assign n58471 = ~n58469 & ~n58470 ;
  assign n58472 = ~n58461 & n58471 ;
  assign n58473 = ~n58465 & n58472 ;
  assign n58476 = n8828 & n49792 ;
  assign n58475 = ~\P1_P3_InstQueue_reg[11][6]/NET0131  & ~n49792 ;
  assign n58477 = n10046 & ~n58475 ;
  assign n58478 = ~n58476 & n58477 ;
  assign n58474 = \P1_P3_InstQueue_reg[11][6]/NET0131  & ~n49798 ;
  assign n58479 = \P1_buf2_reg[30]/NET0131  & n49771 ;
  assign n58480 = \P1_buf2_reg[22]/NET0131  & n49768 ;
  assign n58481 = ~n58479 & ~n58480 ;
  assign n58482 = n11698 & ~n58481 ;
  assign n58483 = \P1_buf2_reg[6]/NET0131  & n49808 ;
  assign n58484 = ~n58482 & ~n58483 ;
  assign n58485 = ~n58474 & n58484 ;
  assign n58486 = ~n58478 & n58485 ;
  assign n58489 = n8955 & n49814 ;
  assign n58488 = ~\P1_P3_InstQueue_reg[12][3]/NET0131  & ~n49814 ;
  assign n58490 = n10046 & ~n58488 ;
  assign n58491 = ~n58489 & n58490 ;
  assign n58487 = \P1_P3_InstQueue_reg[12][3]/NET0131  & ~n49819 ;
  assign n58492 = \P1_buf2_reg[27]/NET0131  & n49768 ;
  assign n58493 = \P1_buf2_reg[19]/NET0131  & n49766 ;
  assign n58494 = ~n58492 & ~n58493 ;
  assign n58495 = n11698 & ~n58494 ;
  assign n58496 = \P1_buf2_reg[3]/NET0131  & n49829 ;
  assign n58497 = ~n58495 & ~n58496 ;
  assign n58498 = ~n58487 & n58497 ;
  assign n58499 = ~n58491 & n58498 ;
  assign n58502 = n8828 & n49814 ;
  assign n58501 = ~\P1_P3_InstQueue_reg[12][6]/NET0131  & ~n49814 ;
  assign n58503 = n10046 & ~n58501 ;
  assign n58504 = ~n58502 & n58503 ;
  assign n58500 = \P1_P3_InstQueue_reg[12][6]/NET0131  & ~n49819 ;
  assign n58505 = \P1_buf2_reg[30]/NET0131  & n49768 ;
  assign n58506 = \P1_buf2_reg[22]/NET0131  & n49766 ;
  assign n58507 = ~n58505 & ~n58506 ;
  assign n58508 = n11698 & ~n58507 ;
  assign n58509 = \P1_buf2_reg[6]/NET0131  & n49829 ;
  assign n58510 = ~n58508 & ~n58509 ;
  assign n58511 = ~n58500 & n58510 ;
  assign n58512 = ~n58504 & n58511 ;
  assign n58515 = n8955 & n49739 ;
  assign n58514 = ~\P1_P3_InstQueue_reg[13][3]/NET0131  & ~n49739 ;
  assign n58516 = n10046 & ~n58514 ;
  assign n58517 = ~n58515 & n58516 ;
  assign n58513 = \P1_P3_InstQueue_reg[13][3]/NET0131  & ~n49838 ;
  assign n58518 = \P1_buf2_reg[27]/NET0131  & n49766 ;
  assign n58519 = \P1_buf2_reg[19]/NET0131  & ~n49766 ;
  assign n58520 = n49792 & n58519 ;
  assign n58521 = ~n58518 & ~n58520 ;
  assign n58522 = n11698 & ~n58521 ;
  assign n58523 = \P1_buf2_reg[3]/NET0131  & n49848 ;
  assign n58524 = ~n58522 & ~n58523 ;
  assign n58525 = ~n58513 & n58524 ;
  assign n58526 = ~n58517 & n58525 ;
  assign n58529 = n8828 & n49739 ;
  assign n58528 = ~\P1_P3_InstQueue_reg[13][6]/NET0131  & ~n49739 ;
  assign n58530 = n10046 & ~n58528 ;
  assign n58531 = ~n58529 & n58530 ;
  assign n58527 = \P1_P3_InstQueue_reg[13][6]/NET0131  & ~n49838 ;
  assign n58532 = \P1_buf2_reg[30]/NET0131  & n49766 ;
  assign n58533 = \P1_buf2_reg[22]/NET0131  & ~n49766 ;
  assign n58534 = n49792 & n58533 ;
  assign n58535 = ~n58532 & ~n58534 ;
  assign n58536 = n11698 & ~n58535 ;
  assign n58537 = \P1_buf2_reg[6]/NET0131  & n49848 ;
  assign n58538 = ~n58536 & ~n58537 ;
  assign n58539 = ~n58527 & n58538 ;
  assign n58540 = ~n58531 & n58539 ;
  assign n58543 = n8955 & n49742 ;
  assign n58542 = ~\P1_P3_InstQueue_reg[14][3]/NET0131  & ~n49742 ;
  assign n58544 = n10046 & ~n58542 ;
  assign n58545 = ~n58543 & n58544 ;
  assign n58541 = \P1_P3_InstQueue_reg[14][3]/NET0131  & ~n49856 ;
  assign n58546 = \P1_buf2_reg[27]/NET0131  & n49792 ;
  assign n58547 = \P1_buf2_reg[19]/NET0131  & ~n49792 ;
  assign n58548 = n49814 & n58547 ;
  assign n58549 = ~n58546 & ~n58548 ;
  assign n58550 = n11698 & ~n58549 ;
  assign n58551 = \P1_buf2_reg[3]/NET0131  & n49866 ;
  assign n58552 = ~n58550 & ~n58551 ;
  assign n58553 = ~n58541 & n58552 ;
  assign n58554 = ~n58545 & n58553 ;
  assign n58557 = n8828 & n49742 ;
  assign n58556 = ~\P1_P3_InstQueue_reg[14][6]/NET0131  & ~n49742 ;
  assign n58558 = n10046 & ~n58556 ;
  assign n58559 = ~n58557 & n58558 ;
  assign n58555 = \P1_P3_InstQueue_reg[14][6]/NET0131  & ~n49856 ;
  assign n58560 = \P1_buf2_reg[30]/NET0131  & n49792 ;
  assign n58561 = \P1_buf2_reg[22]/NET0131  & ~n49792 ;
  assign n58562 = n49814 & n58561 ;
  assign n58563 = ~n58560 & ~n58562 ;
  assign n58564 = n11698 & ~n58563 ;
  assign n58565 = \P1_buf2_reg[6]/NET0131  & n49866 ;
  assign n58566 = ~n58564 & ~n58565 ;
  assign n58567 = ~n58555 & n58566 ;
  assign n58568 = ~n58559 & n58567 ;
  assign n58571 = n8955 & n49735 ;
  assign n58570 = ~\P1_P3_InstQueue_reg[15][3]/NET0131  & ~n49735 ;
  assign n58572 = n10046 & ~n58570 ;
  assign n58573 = ~n58571 & n58572 ;
  assign n58569 = \P1_P3_InstQueue_reg[15][3]/NET0131  & ~n49875 ;
  assign n58574 = \P1_buf2_reg[27]/NET0131  & n49814 ;
  assign n58575 = \P1_buf2_reg[19]/NET0131  & n49739 ;
  assign n58576 = ~n58574 & ~n58575 ;
  assign n58577 = n11698 & ~n58576 ;
  assign n58578 = \P1_buf2_reg[3]/NET0131  & n49885 ;
  assign n58579 = ~n58577 & ~n58578 ;
  assign n58580 = ~n58569 & n58579 ;
  assign n58581 = ~n58573 & n58580 ;
  assign n58584 = n8828 & n49735 ;
  assign n58583 = ~\P1_P3_InstQueue_reg[15][6]/NET0131  & ~n49735 ;
  assign n58585 = n10046 & ~n58583 ;
  assign n58586 = ~n58584 & n58585 ;
  assign n58582 = \P1_P3_InstQueue_reg[15][6]/NET0131  & ~n49875 ;
  assign n58587 = \P1_buf2_reg[30]/NET0131  & n49814 ;
  assign n58588 = \P1_buf2_reg[22]/NET0131  & n49739 ;
  assign n58589 = ~n58587 & ~n58588 ;
  assign n58590 = n11698 & ~n58589 ;
  assign n58591 = \P1_buf2_reg[6]/NET0131  & n49885 ;
  assign n58592 = ~n58590 & ~n58591 ;
  assign n58593 = ~n58582 & n58592 ;
  assign n58594 = ~n58586 & n58593 ;
  assign n58597 = n8955 & n49890 ;
  assign n58596 = ~\P1_P3_InstQueue_reg[1][3]/NET0131  & ~n49890 ;
  assign n58598 = n10046 & ~n58596 ;
  assign n58599 = ~n58597 & n58598 ;
  assign n58595 = \P1_P3_InstQueue_reg[1][3]/NET0131  & ~n49895 ;
  assign n58600 = \P1_buf2_reg[27]/NET0131  & n49742 ;
  assign n58601 = \P1_buf2_reg[19]/NET0131  & n49735 ;
  assign n58602 = ~n58600 & ~n58601 ;
  assign n58603 = n11698 & ~n58602 ;
  assign n58604 = \P1_buf2_reg[3]/NET0131  & n49905 ;
  assign n58605 = ~n58603 & ~n58604 ;
  assign n58606 = ~n58595 & n58605 ;
  assign n58607 = ~n58599 & n58606 ;
  assign n58610 = n8828 & n49890 ;
  assign n58609 = ~\P1_P3_InstQueue_reg[1][6]/NET0131  & ~n49890 ;
  assign n58611 = n10046 & ~n58609 ;
  assign n58612 = ~n58610 & n58611 ;
  assign n58608 = \P1_P3_InstQueue_reg[1][6]/NET0131  & ~n49895 ;
  assign n58613 = \P1_buf2_reg[30]/NET0131  & n49742 ;
  assign n58614 = \P1_buf2_reg[22]/NET0131  & n49735 ;
  assign n58615 = ~n58613 & ~n58614 ;
  assign n58616 = n11698 & ~n58615 ;
  assign n58617 = \P1_buf2_reg[6]/NET0131  & n49905 ;
  assign n58618 = ~n58616 & ~n58617 ;
  assign n58619 = ~n58608 & n58618 ;
  assign n58620 = ~n58612 & n58619 ;
  assign n58623 = n8955 & n49910 ;
  assign n58622 = ~\P1_P3_InstQueue_reg[2][3]/NET0131  & ~n49910 ;
  assign n58624 = n10046 & ~n58622 ;
  assign n58625 = ~n58623 & n58624 ;
  assign n58621 = \P1_P3_InstQueue_reg[2][3]/NET0131  & ~n49915 ;
  assign n58626 = \P1_buf2_reg[27]/NET0131  & n49735 ;
  assign n58627 = \P1_buf2_reg[19]/NET0131  & n49732 ;
  assign n58628 = ~n58626 & ~n58627 ;
  assign n58629 = n11698 & ~n58628 ;
  assign n58630 = \P1_buf2_reg[3]/NET0131  & n49925 ;
  assign n58631 = ~n58629 & ~n58630 ;
  assign n58632 = ~n58621 & n58631 ;
  assign n58633 = ~n58625 & n58632 ;
  assign n58636 = n8828 & n49910 ;
  assign n58635 = ~\P1_P3_InstQueue_reg[2][6]/NET0131  & ~n49910 ;
  assign n58637 = n10046 & ~n58635 ;
  assign n58638 = ~n58636 & n58637 ;
  assign n58634 = \P1_P3_InstQueue_reg[2][6]/NET0131  & ~n49915 ;
  assign n58639 = \P1_buf2_reg[30]/NET0131  & n49735 ;
  assign n58640 = \P1_buf2_reg[22]/NET0131  & n49732 ;
  assign n58641 = ~n58639 & ~n58640 ;
  assign n58642 = n11698 & ~n58641 ;
  assign n58643 = \P1_buf2_reg[6]/NET0131  & n49925 ;
  assign n58644 = ~n58642 & ~n58643 ;
  assign n58645 = ~n58634 & n58644 ;
  assign n58646 = ~n58638 & n58645 ;
  assign n58649 = n8955 & n49930 ;
  assign n58648 = ~\P1_P3_InstQueue_reg[3][3]/NET0131  & ~n49930 ;
  assign n58650 = n10046 & ~n58648 ;
  assign n58651 = ~n58649 & n58650 ;
  assign n58647 = \P1_P3_InstQueue_reg[3][3]/NET0131  & ~n49935 ;
  assign n58652 = \P1_buf2_reg[27]/NET0131  & n49732 ;
  assign n58653 = \P1_buf2_reg[19]/NET0131  & ~n49732 ;
  assign n58654 = n49890 & n58653 ;
  assign n58655 = ~n58652 & ~n58654 ;
  assign n58656 = n11698 & ~n58655 ;
  assign n58657 = \P1_buf2_reg[3]/NET0131  & n49945 ;
  assign n58658 = ~n58656 & ~n58657 ;
  assign n58659 = ~n58647 & n58658 ;
  assign n58660 = ~n58651 & n58659 ;
  assign n58663 = n8828 & n49930 ;
  assign n58662 = ~\P1_P3_InstQueue_reg[3][6]/NET0131  & ~n49930 ;
  assign n58664 = n10046 & ~n58662 ;
  assign n58665 = ~n58663 & n58664 ;
  assign n58661 = \P1_P3_InstQueue_reg[3][6]/NET0131  & ~n49935 ;
  assign n58666 = \P1_buf2_reg[30]/NET0131  & n49732 ;
  assign n58667 = \P1_buf2_reg[22]/NET0131  & ~n49732 ;
  assign n58668 = n49890 & n58667 ;
  assign n58669 = ~n58666 & ~n58668 ;
  assign n58670 = n11698 & ~n58669 ;
  assign n58671 = \P1_buf2_reg[6]/NET0131  & n49945 ;
  assign n58672 = ~n58670 & ~n58671 ;
  assign n58673 = ~n58661 & n58672 ;
  assign n58674 = ~n58665 & n58673 ;
  assign n58677 = n8955 & n49950 ;
  assign n58676 = ~\P1_P3_InstQueue_reg[4][3]/NET0131  & ~n49950 ;
  assign n58678 = n10046 & ~n58676 ;
  assign n58679 = ~n58677 & n58678 ;
  assign n58675 = \P1_P3_InstQueue_reg[4][3]/NET0131  & ~n49955 ;
  assign n58680 = \P1_buf2_reg[27]/NET0131  & n49890 ;
  assign n58681 = \P1_buf2_reg[19]/NET0131  & ~n49890 ;
  assign n58682 = n49910 & n58681 ;
  assign n58683 = ~n58680 & ~n58682 ;
  assign n58684 = n11698 & ~n58683 ;
  assign n58685 = \P1_buf2_reg[3]/NET0131  & n49965 ;
  assign n58686 = ~n58684 & ~n58685 ;
  assign n58687 = ~n58675 & n58686 ;
  assign n58688 = ~n58679 & n58687 ;
  assign n58691 = n8828 & n49950 ;
  assign n58690 = ~\P1_P3_InstQueue_reg[4][6]/NET0131  & ~n49950 ;
  assign n58692 = n10046 & ~n58690 ;
  assign n58693 = ~n58691 & n58692 ;
  assign n58689 = \P1_P3_InstQueue_reg[4][6]/NET0131  & ~n49955 ;
  assign n58694 = \P1_buf2_reg[30]/NET0131  & n49890 ;
  assign n58695 = \P1_buf2_reg[22]/NET0131  & ~n49890 ;
  assign n58696 = n49910 & n58695 ;
  assign n58697 = ~n58694 & ~n58696 ;
  assign n58698 = n11698 & ~n58697 ;
  assign n58699 = \P1_buf2_reg[6]/NET0131  & n49965 ;
  assign n58700 = ~n58698 & ~n58699 ;
  assign n58701 = ~n58689 & n58700 ;
  assign n58702 = ~n58693 & n58701 ;
  assign n58705 = n8955 & n49970 ;
  assign n58704 = ~\P1_P3_InstQueue_reg[5][3]/NET0131  & ~n49970 ;
  assign n58706 = n10046 & ~n58704 ;
  assign n58707 = ~n58705 & n58706 ;
  assign n58703 = \P1_P3_InstQueue_reg[5][3]/NET0131  & ~n49975 ;
  assign n58708 = \P1_buf2_reg[27]/NET0131  & n49910 ;
  assign n58709 = \P1_buf2_reg[19]/NET0131  & ~n49910 ;
  assign n58710 = n49930 & n58709 ;
  assign n58711 = ~n58708 & ~n58710 ;
  assign n58712 = n11698 & ~n58711 ;
  assign n58713 = \P1_buf2_reg[3]/NET0131  & n49985 ;
  assign n58714 = ~n58712 & ~n58713 ;
  assign n58715 = ~n58703 & n58714 ;
  assign n58716 = ~n58707 & n58715 ;
  assign n58719 = n8828 & n49970 ;
  assign n58718 = ~\P1_P3_InstQueue_reg[5][6]/NET0131  & ~n49970 ;
  assign n58720 = n10046 & ~n58718 ;
  assign n58721 = ~n58719 & n58720 ;
  assign n58717 = \P1_P3_InstQueue_reg[5][6]/NET0131  & ~n49975 ;
  assign n58722 = \P1_buf2_reg[30]/NET0131  & n49910 ;
  assign n58723 = \P1_buf2_reg[22]/NET0131  & ~n49910 ;
  assign n58724 = n49930 & n58723 ;
  assign n58725 = ~n58722 & ~n58724 ;
  assign n58726 = n11698 & ~n58725 ;
  assign n58727 = \P1_buf2_reg[6]/NET0131  & n49985 ;
  assign n58728 = ~n58726 & ~n58727 ;
  assign n58729 = ~n58717 & n58728 ;
  assign n58730 = ~n58721 & n58729 ;
  assign n58733 = n8955 & n49990 ;
  assign n58732 = ~\P1_P3_InstQueue_reg[6][3]/NET0131  & ~n49990 ;
  assign n58734 = n10046 & ~n58732 ;
  assign n58735 = ~n58733 & n58734 ;
  assign n58731 = \P1_P3_InstQueue_reg[6][3]/NET0131  & ~n49995 ;
  assign n58736 = \P1_buf2_reg[27]/NET0131  & n49930 ;
  assign n58737 = \P1_buf2_reg[19]/NET0131  & ~n49930 ;
  assign n58738 = n49950 & n58737 ;
  assign n58739 = ~n58736 & ~n58738 ;
  assign n58740 = n11698 & ~n58739 ;
  assign n58741 = \P1_buf2_reg[3]/NET0131  & n50005 ;
  assign n58742 = ~n58740 & ~n58741 ;
  assign n58743 = ~n58731 & n58742 ;
  assign n58744 = ~n58735 & n58743 ;
  assign n58747 = n27054 & n50021 ;
  assign n58746 = ~\P2_P3_InstQueue_reg[0][3]/NET0131  & ~n50021 ;
  assign n58748 = n27788 & ~n58746 ;
  assign n58749 = ~n58747 & n58748 ;
  assign n58745 = \P2_P3_InstQueue_reg[0][3]/NET0131  & ~n50030 ;
  assign n58750 = \P2_buf2_reg[27]/NET0131  & n50012 ;
  assign n58751 = \P2_buf2_reg[19]/NET0131  & n50015 ;
  assign n58752 = ~n58750 & ~n58751 ;
  assign n58753 = n27325 & ~n58752 ;
  assign n58754 = \P2_buf2_reg[3]/NET0131  & n50040 ;
  assign n58755 = ~n58753 & ~n58754 ;
  assign n58756 = ~n58745 & n58755 ;
  assign n58757 = ~n58749 & n58756 ;
  assign n58760 = n8828 & n49990 ;
  assign n58759 = ~\P1_P3_InstQueue_reg[6][6]/NET0131  & ~n49990 ;
  assign n58761 = n10046 & ~n58759 ;
  assign n58762 = ~n58760 & n58761 ;
  assign n58758 = \P1_P3_InstQueue_reg[6][6]/NET0131  & ~n49995 ;
  assign n58763 = \P1_buf2_reg[30]/NET0131  & n49930 ;
  assign n58764 = \P1_buf2_reg[22]/NET0131  & ~n49930 ;
  assign n58765 = n49950 & n58764 ;
  assign n58766 = ~n58763 & ~n58765 ;
  assign n58767 = n11698 & ~n58766 ;
  assign n58768 = \P1_buf2_reg[6]/NET0131  & n50005 ;
  assign n58769 = ~n58767 & ~n58768 ;
  assign n58770 = ~n58758 & n58769 ;
  assign n58771 = ~n58762 & n58770 ;
  assign n58774 = n26927 & n50021 ;
  assign n58773 = ~\P2_P3_InstQueue_reg[0][6]/NET0131  & ~n50021 ;
  assign n58775 = n27788 & ~n58773 ;
  assign n58776 = ~n58774 & n58775 ;
  assign n58772 = \P2_P3_InstQueue_reg[0][6]/NET0131  & ~n50030 ;
  assign n58777 = \P2_buf2_reg[30]/NET0131  & n50012 ;
  assign n58778 = \P2_buf2_reg[22]/NET0131  & n50015 ;
  assign n58779 = ~n58777 & ~n58778 ;
  assign n58780 = n27325 & ~n58779 ;
  assign n58781 = \P2_buf2_reg[6]/NET0131  & n50040 ;
  assign n58782 = ~n58780 & ~n58781 ;
  assign n58783 = ~n58772 & n58782 ;
  assign n58784 = ~n58776 & n58783 ;
  assign n58787 = n27054 & n50051 ;
  assign n58786 = ~\P2_P3_InstQueue_reg[10][3]/NET0131  & ~n50051 ;
  assign n58788 = n27788 & ~n58786 ;
  assign n58789 = ~n58787 & n58788 ;
  assign n58785 = \P2_P3_InstQueue_reg[10][3]/NET0131  & ~n50056 ;
  assign n58790 = \P2_buf2_reg[19]/NET0131  & n50045 ;
  assign n58791 = \P2_buf2_reg[27]/NET0131  & n50046 ;
  assign n58792 = ~n58790 & ~n58791 ;
  assign n58793 = n27325 & ~n58792 ;
  assign n58794 = \P2_buf2_reg[3]/NET0131  & n50066 ;
  assign n58795 = ~n58793 & ~n58794 ;
  assign n58796 = ~n58785 & n58795 ;
  assign n58797 = ~n58789 & n58796 ;
  assign n58800 = n26927 & n50051 ;
  assign n58799 = ~\P2_P3_InstQueue_reg[10][6]/NET0131  & ~n50051 ;
  assign n58801 = n27788 & ~n58799 ;
  assign n58802 = ~n58800 & n58801 ;
  assign n58798 = \P2_P3_InstQueue_reg[10][6]/NET0131  & ~n50056 ;
  assign n58803 = \P2_buf2_reg[22]/NET0131  & n50045 ;
  assign n58804 = \P2_buf2_reg[30]/NET0131  & n50046 ;
  assign n58805 = ~n58803 & ~n58804 ;
  assign n58806 = n27325 & ~n58805 ;
  assign n58807 = \P2_buf2_reg[6]/NET0131  & n50066 ;
  assign n58808 = ~n58806 & ~n58807 ;
  assign n58809 = ~n58798 & n58808 ;
  assign n58810 = ~n58802 & n58809 ;
  assign n58813 = n8955 & n49770 ;
  assign n58812 = ~\P1_P3_InstQueue_reg[7][3]/NET0131  & ~n49770 ;
  assign n58814 = n10046 & ~n58812 ;
  assign n58815 = ~n58813 & n58814 ;
  assign n58811 = \P1_P3_InstQueue_reg[7][3]/NET0131  & ~n50075 ;
  assign n58816 = \P1_buf2_reg[27]/NET0131  & n49950 ;
  assign n58817 = \P1_buf2_reg[19]/NET0131  & ~n49950 ;
  assign n58818 = n49970 & n58817 ;
  assign n58819 = ~n58816 & ~n58818 ;
  assign n58820 = n11698 & ~n58819 ;
  assign n58821 = \P1_buf2_reg[3]/NET0131  & n50085 ;
  assign n58822 = ~n58820 & ~n58821 ;
  assign n58823 = ~n58811 & n58822 ;
  assign n58824 = ~n58815 & n58823 ;
  assign n58827 = n27054 & n50094 ;
  assign n58826 = ~\P2_P3_InstQueue_reg[11][3]/NET0131  & ~n50094 ;
  assign n58828 = n27788 & ~n58826 ;
  assign n58829 = ~n58827 & n58828 ;
  assign n58825 = \P2_P3_InstQueue_reg[11][3]/NET0131  & ~n50097 ;
  assign n58830 = \P2_buf2_reg[27]/NET0131  & n50045 ;
  assign n58831 = \P2_buf2_reg[19]/NET0131  & n50053 ;
  assign n58832 = ~n58830 & ~n58831 ;
  assign n58833 = n27325 & ~n58832 ;
  assign n58834 = \P2_buf2_reg[3]/NET0131  & n50107 ;
  assign n58835 = ~n58833 & ~n58834 ;
  assign n58836 = ~n58825 & n58835 ;
  assign n58837 = ~n58829 & n58836 ;
  assign n58840 = n8828 & n49770 ;
  assign n58839 = ~\P1_P3_InstQueue_reg[7][6]/NET0131  & ~n49770 ;
  assign n58841 = n10046 & ~n58839 ;
  assign n58842 = ~n58840 & n58841 ;
  assign n58838 = \P1_P3_InstQueue_reg[7][6]/NET0131  & ~n50075 ;
  assign n58843 = \P1_buf2_reg[30]/NET0131  & n49950 ;
  assign n58844 = \P1_buf2_reg[22]/NET0131  & ~n49950 ;
  assign n58845 = n49970 & n58844 ;
  assign n58846 = ~n58843 & ~n58845 ;
  assign n58847 = n11698 & ~n58846 ;
  assign n58848 = \P1_buf2_reg[6]/NET0131  & n50085 ;
  assign n58849 = ~n58847 & ~n58848 ;
  assign n58850 = ~n58838 & n58849 ;
  assign n58851 = ~n58842 & n58850 ;
  assign n58854 = n26927 & n50094 ;
  assign n58853 = ~\P2_P3_InstQueue_reg[11][6]/NET0131  & ~n50094 ;
  assign n58855 = n27788 & ~n58853 ;
  assign n58856 = ~n58854 & n58855 ;
  assign n58852 = \P2_P3_InstQueue_reg[11][6]/NET0131  & ~n50097 ;
  assign n58857 = \P2_buf2_reg[30]/NET0131  & n50045 ;
  assign n58858 = \P2_buf2_reg[22]/NET0131  & n50053 ;
  assign n58859 = ~n58857 & ~n58858 ;
  assign n58860 = n27325 & ~n58859 ;
  assign n58861 = \P2_buf2_reg[6]/NET0131  & n50107 ;
  assign n58862 = ~n58860 & ~n58861 ;
  assign n58863 = ~n58852 & n58862 ;
  assign n58864 = ~n58856 & n58863 ;
  assign n58867 = n27054 & n50115 ;
  assign n58866 = ~\P2_P3_InstQueue_reg[12][3]/NET0131  & ~n50115 ;
  assign n58868 = n27788 & ~n58866 ;
  assign n58869 = ~n58867 & n58868 ;
  assign n58865 = \P2_P3_InstQueue_reg[12][3]/NET0131  & ~n50118 ;
  assign n58870 = \P2_buf2_reg[27]/NET0131  & n50053 ;
  assign n58871 = \P2_buf2_reg[19]/NET0131  & n50051 ;
  assign n58872 = ~n58870 & ~n58871 ;
  assign n58873 = n27325 & ~n58872 ;
  assign n58874 = \P2_buf2_reg[3]/NET0131  & n50128 ;
  assign n58875 = ~n58873 & ~n58874 ;
  assign n58876 = ~n58865 & n58875 ;
  assign n58877 = ~n58869 & n58876 ;
  assign n58880 = n26927 & n50115 ;
  assign n58879 = ~\P2_P3_InstQueue_reg[12][6]/NET0131  & ~n50115 ;
  assign n58881 = n27788 & ~n58879 ;
  assign n58882 = ~n58880 & n58881 ;
  assign n58878 = \P2_P3_InstQueue_reg[12][6]/NET0131  & ~n50118 ;
  assign n58883 = \P2_buf2_reg[30]/NET0131  & n50053 ;
  assign n58884 = \P2_buf2_reg[22]/NET0131  & n50051 ;
  assign n58885 = ~n58883 & ~n58884 ;
  assign n58886 = n27325 & ~n58885 ;
  assign n58887 = \P2_buf2_reg[6]/NET0131  & n50128 ;
  assign n58888 = ~n58886 & ~n58887 ;
  assign n58889 = ~n58878 & n58888 ;
  assign n58890 = ~n58882 & n58889 ;
  assign n58893 = n8955 & n49771 ;
  assign n58892 = ~\P1_P3_InstQueue_reg[8][3]/NET0131  & ~n49771 ;
  assign n58894 = n10046 & ~n58892 ;
  assign n58895 = ~n58893 & n58894 ;
  assign n58891 = \P1_P3_InstQueue_reg[8][3]/NET0131  & ~n50136 ;
  assign n58896 = \P1_buf2_reg[27]/NET0131  & n49970 ;
  assign n58897 = \P1_buf2_reg[19]/NET0131  & ~n49970 ;
  assign n58898 = n49990 & n58897 ;
  assign n58899 = ~n58896 & ~n58898 ;
  assign n58900 = n11698 & ~n58899 ;
  assign n58901 = \P1_buf2_reg[3]/NET0131  & n50146 ;
  assign n58902 = ~n58900 & ~n58901 ;
  assign n58903 = ~n58891 & n58902 ;
  assign n58904 = ~n58895 & n58903 ;
  assign n58907 = n27054 & n50012 ;
  assign n58906 = ~\P2_P3_InstQueue_reg[13][3]/NET0131  & ~n50012 ;
  assign n58908 = n27788 & ~n58906 ;
  assign n58909 = ~n58907 & n58908 ;
  assign n58905 = \P2_P3_InstQueue_reg[13][3]/NET0131  & ~n50155 ;
  assign n58910 = \P2_buf2_reg[27]/NET0131  & n50051 ;
  assign n58911 = \P2_buf2_reg[19]/NET0131  & n50094 ;
  assign n58912 = ~n58910 & ~n58911 ;
  assign n58913 = n27325 & ~n58912 ;
  assign n58914 = \P2_buf2_reg[3]/NET0131  & n50165 ;
  assign n58915 = ~n58913 & ~n58914 ;
  assign n58916 = ~n58905 & n58915 ;
  assign n58917 = ~n58909 & n58916 ;
  assign n58920 = n8828 & n49771 ;
  assign n58919 = ~\P1_P3_InstQueue_reg[8][6]/NET0131  & ~n49771 ;
  assign n58921 = n10046 & ~n58919 ;
  assign n58922 = ~n58920 & n58921 ;
  assign n58918 = \P1_P3_InstQueue_reg[8][6]/NET0131  & ~n50136 ;
  assign n58923 = \P1_buf2_reg[30]/NET0131  & n49970 ;
  assign n58924 = \P1_buf2_reg[22]/NET0131  & ~n49970 ;
  assign n58925 = n49990 & n58924 ;
  assign n58926 = ~n58923 & ~n58925 ;
  assign n58927 = n11698 & ~n58926 ;
  assign n58928 = \P1_buf2_reg[6]/NET0131  & n50146 ;
  assign n58929 = ~n58927 & ~n58928 ;
  assign n58930 = ~n58918 & n58929 ;
  assign n58931 = ~n58922 & n58930 ;
  assign n58934 = n26927 & n50012 ;
  assign n58933 = ~\P2_P3_InstQueue_reg[13][6]/NET0131  & ~n50012 ;
  assign n58935 = n27788 & ~n58933 ;
  assign n58936 = ~n58934 & n58935 ;
  assign n58932 = \P2_P3_InstQueue_reg[13][6]/NET0131  & ~n50155 ;
  assign n58937 = \P2_buf2_reg[30]/NET0131  & n50051 ;
  assign n58938 = \P2_buf2_reg[22]/NET0131  & n50094 ;
  assign n58939 = ~n58937 & ~n58938 ;
  assign n58940 = n27325 & ~n58939 ;
  assign n58941 = \P2_buf2_reg[6]/NET0131  & n50165 ;
  assign n58942 = ~n58940 & ~n58941 ;
  assign n58943 = ~n58932 & n58942 ;
  assign n58944 = ~n58936 & n58943 ;
  assign n58947 = n27054 & n50015 ;
  assign n58946 = ~\P2_P3_InstQueue_reg[14][3]/NET0131  & ~n50015 ;
  assign n58948 = n27788 & ~n58946 ;
  assign n58949 = ~n58947 & n58948 ;
  assign n58945 = \P2_P3_InstQueue_reg[14][3]/NET0131  & ~n50173 ;
  assign n58950 = \P2_buf2_reg[27]/NET0131  & n50094 ;
  assign n58951 = \P2_buf2_reg[19]/NET0131  & n50115 ;
  assign n58952 = ~n58950 & ~n58951 ;
  assign n58953 = n27325 & ~n58952 ;
  assign n58954 = \P2_buf2_reg[3]/NET0131  & n50183 ;
  assign n58955 = ~n58953 & ~n58954 ;
  assign n58956 = ~n58945 & n58955 ;
  assign n58957 = ~n58949 & n58956 ;
  assign n58960 = n26927 & n50015 ;
  assign n58959 = ~\P2_P3_InstQueue_reg[14][6]/NET0131  & ~n50015 ;
  assign n58961 = n27788 & ~n58959 ;
  assign n58962 = ~n58960 & n58961 ;
  assign n58958 = \P2_P3_InstQueue_reg[14][6]/NET0131  & ~n50173 ;
  assign n58963 = \P2_buf2_reg[30]/NET0131  & n50094 ;
  assign n58964 = \P2_buf2_reg[22]/NET0131  & n50115 ;
  assign n58965 = ~n58963 & ~n58964 ;
  assign n58966 = n27325 & ~n58965 ;
  assign n58967 = \P2_buf2_reg[6]/NET0131  & n50183 ;
  assign n58968 = ~n58966 & ~n58967 ;
  assign n58969 = ~n58958 & n58968 ;
  assign n58970 = ~n58962 & n58969 ;
  assign n58973 = n8955 & n49768 ;
  assign n58972 = ~\P1_P3_InstQueue_reg[9][3]/NET0131  & ~n49768 ;
  assign n58974 = n10046 & ~n58972 ;
  assign n58975 = ~n58973 & n58974 ;
  assign n58971 = \P1_P3_InstQueue_reg[9][3]/NET0131  & ~n50191 ;
  assign n58976 = \P1_buf2_reg[27]/NET0131  & n49990 ;
  assign n58977 = \P1_buf2_reg[19]/NET0131  & n49770 ;
  assign n58978 = ~n58976 & ~n58977 ;
  assign n58979 = n11698 & ~n58978 ;
  assign n58980 = \P1_buf2_reg[3]/NET0131  & n50201 ;
  assign n58981 = ~n58979 & ~n58980 ;
  assign n58982 = ~n58971 & n58981 ;
  assign n58983 = ~n58975 & n58982 ;
  assign n58986 = n27054 & n50024 ;
  assign n58985 = ~\P2_P3_InstQueue_reg[15][3]/NET0131  & ~n50024 ;
  assign n58987 = n27788 & ~n58985 ;
  assign n58988 = ~n58986 & n58987 ;
  assign n58984 = \P2_P3_InstQueue_reg[15][3]/NET0131  & ~n50210 ;
  assign n58989 = \P2_buf2_reg[27]/NET0131  & n50115 ;
  assign n58990 = \P2_buf2_reg[19]/NET0131  & n50012 ;
  assign n58991 = ~n58989 & ~n58990 ;
  assign n58992 = n27325 & ~n58991 ;
  assign n58993 = \P2_buf2_reg[3]/NET0131  & n50220 ;
  assign n58994 = ~n58992 & ~n58993 ;
  assign n58995 = ~n58984 & n58994 ;
  assign n58996 = ~n58988 & n58995 ;
  assign n58999 = n8828 & n49768 ;
  assign n58998 = ~\P1_P3_InstQueue_reg[9][6]/NET0131  & ~n49768 ;
  assign n59000 = n10046 & ~n58998 ;
  assign n59001 = ~n58999 & n59000 ;
  assign n58997 = \P1_P3_InstQueue_reg[9][6]/NET0131  & ~n50191 ;
  assign n59002 = \P1_buf2_reg[30]/NET0131  & n49990 ;
  assign n59003 = \P1_buf2_reg[22]/NET0131  & n49770 ;
  assign n59004 = ~n59002 & ~n59003 ;
  assign n59005 = n11698 & ~n59004 ;
  assign n59006 = \P1_buf2_reg[6]/NET0131  & n50201 ;
  assign n59007 = ~n59005 & ~n59006 ;
  assign n59008 = ~n58997 & n59007 ;
  assign n59009 = ~n59001 & n59008 ;
  assign n59012 = n26927 & n50024 ;
  assign n59011 = ~\P2_P3_InstQueue_reg[15][6]/NET0131  & ~n50024 ;
  assign n59013 = n27788 & ~n59011 ;
  assign n59014 = ~n59012 & n59013 ;
  assign n59010 = \P2_P3_InstQueue_reg[15][6]/NET0131  & ~n50210 ;
  assign n59015 = \P2_buf2_reg[30]/NET0131  & n50115 ;
  assign n59016 = \P2_buf2_reg[22]/NET0131  & n50012 ;
  assign n59017 = ~n59015 & ~n59016 ;
  assign n59018 = n27325 & ~n59017 ;
  assign n59019 = \P2_buf2_reg[6]/NET0131  & n50220 ;
  assign n59020 = ~n59018 & ~n59019 ;
  assign n59021 = ~n59010 & n59020 ;
  assign n59022 = ~n59014 & n59021 ;
  assign n59025 = n27054 & n50227 ;
  assign n59024 = ~\P2_P3_InstQueue_reg[1][3]/NET0131  & ~n50227 ;
  assign n59026 = n27788 & ~n59024 ;
  assign n59027 = ~n59025 & n59026 ;
  assign n59023 = \P2_P3_InstQueue_reg[1][3]/NET0131  & ~n50230 ;
  assign n59028 = \P2_buf2_reg[27]/NET0131  & n50015 ;
  assign n59029 = \P2_buf2_reg[19]/NET0131  & n50024 ;
  assign n59030 = ~n59028 & ~n59029 ;
  assign n59031 = n27325 & ~n59030 ;
  assign n59032 = \P2_buf2_reg[3]/NET0131  & n50240 ;
  assign n59033 = ~n59031 & ~n59032 ;
  assign n59034 = ~n59023 & n59033 ;
  assign n59035 = ~n59027 & n59034 ;
  assign n59039 = n9241 & ~n37992 ;
  assign n59040 = ~n9245 & ~n10031 ;
  assign n59041 = n17458 & n59040 ;
  assign n59042 = ~n59039 & n59041 ;
  assign n59043 = \P1_P3_PhyAddrPointer_reg[0]/NET0131  & ~n59042 ;
  assign n59036 = n9064 & n45654 ;
  assign n59037 = ~n45661 & ~n59036 ;
  assign n59038 = n9241 & ~n59037 ;
  assign n59044 = ~n45650 & ~n59038 ;
  assign n59045 = ~n59043 & n59044 ;
  assign n59048 = n26927 & n50227 ;
  assign n59047 = ~\P2_P3_InstQueue_reg[1][6]/NET0131  & ~n50227 ;
  assign n59049 = n27788 & ~n59047 ;
  assign n59050 = ~n59048 & n59049 ;
  assign n59046 = \P2_P3_InstQueue_reg[1][6]/NET0131  & ~n50230 ;
  assign n59051 = \P2_buf2_reg[30]/NET0131  & n50015 ;
  assign n59052 = \P2_buf2_reg[22]/NET0131  & n50024 ;
  assign n59053 = ~n59051 & ~n59052 ;
  assign n59054 = n27325 & ~n59053 ;
  assign n59055 = \P2_buf2_reg[6]/NET0131  & n50240 ;
  assign n59056 = ~n59054 & ~n59055 ;
  assign n59057 = ~n59046 & n59056 ;
  assign n59058 = ~n59050 & n59057 ;
  assign n59061 = n27054 & n50247 ;
  assign n59060 = ~\P2_P3_InstQueue_reg[2][3]/NET0131  & ~n50247 ;
  assign n59062 = n27788 & ~n59060 ;
  assign n59063 = ~n59061 & n59062 ;
  assign n59059 = \P2_P3_InstQueue_reg[2][3]/NET0131  & ~n50250 ;
  assign n59064 = \P2_buf2_reg[19]/NET0131  & n50021 ;
  assign n59065 = \P2_buf2_reg[27]/NET0131  & n50024 ;
  assign n59066 = ~n59064 & ~n59065 ;
  assign n59067 = n27325 & ~n59066 ;
  assign n59068 = \P2_buf2_reg[3]/NET0131  & n50260 ;
  assign n59069 = ~n59067 & ~n59068 ;
  assign n59070 = ~n59059 & n59069 ;
  assign n59071 = ~n59063 & n59070 ;
  assign n59074 = n26927 & n50247 ;
  assign n59073 = ~\P2_P3_InstQueue_reg[2][6]/NET0131  & ~n50247 ;
  assign n59075 = n27788 & ~n59073 ;
  assign n59076 = ~n59074 & n59075 ;
  assign n59072 = \P2_P3_InstQueue_reg[2][6]/NET0131  & ~n50250 ;
  assign n59077 = \P2_buf2_reg[22]/NET0131  & n50021 ;
  assign n59078 = \P2_buf2_reg[30]/NET0131  & n50024 ;
  assign n59079 = ~n59077 & ~n59078 ;
  assign n59080 = n27325 & ~n59079 ;
  assign n59081 = \P2_buf2_reg[6]/NET0131  & n50260 ;
  assign n59082 = ~n59080 & ~n59081 ;
  assign n59083 = ~n59072 & n59082 ;
  assign n59084 = ~n59076 & n59083 ;
  assign n59087 = n27054 & n50267 ;
  assign n59086 = ~\P2_P3_InstQueue_reg[3][3]/NET0131  & ~n50267 ;
  assign n59088 = n27788 & ~n59086 ;
  assign n59089 = ~n59087 & n59088 ;
  assign n59085 = \P2_P3_InstQueue_reg[3][3]/NET0131  & ~n50270 ;
  assign n59090 = \P2_buf2_reg[27]/NET0131  & n50021 ;
  assign n59091 = \P2_buf2_reg[19]/NET0131  & n50227 ;
  assign n59092 = ~n59090 & ~n59091 ;
  assign n59093 = n27325 & ~n59092 ;
  assign n59094 = \P2_buf2_reg[3]/NET0131  & n50280 ;
  assign n59095 = ~n59093 & ~n59094 ;
  assign n59096 = ~n59085 & n59095 ;
  assign n59097 = ~n59089 & n59096 ;
  assign n59100 = n26927 & n50267 ;
  assign n59099 = ~\P2_P3_InstQueue_reg[3][6]/NET0131  & ~n50267 ;
  assign n59101 = n27788 & ~n59099 ;
  assign n59102 = ~n59100 & n59101 ;
  assign n59098 = \P2_P3_InstQueue_reg[3][6]/NET0131  & ~n50270 ;
  assign n59103 = \P2_buf2_reg[30]/NET0131  & n50021 ;
  assign n59104 = \P2_buf2_reg[22]/NET0131  & n50227 ;
  assign n59105 = ~n59103 & ~n59104 ;
  assign n59106 = n27325 & ~n59105 ;
  assign n59107 = \P2_buf2_reg[6]/NET0131  & n50280 ;
  assign n59108 = ~n59106 & ~n59107 ;
  assign n59109 = ~n59098 & n59108 ;
  assign n59110 = ~n59102 & n59109 ;
  assign n59113 = n27054 & n50287 ;
  assign n59112 = ~\P2_P3_InstQueue_reg[4][3]/NET0131  & ~n50287 ;
  assign n59114 = n27788 & ~n59112 ;
  assign n59115 = ~n59113 & n59114 ;
  assign n59111 = \P2_P3_InstQueue_reg[4][3]/NET0131  & ~n50290 ;
  assign n59116 = \P2_buf2_reg[27]/NET0131  & n50227 ;
  assign n59117 = \P2_buf2_reg[19]/NET0131  & n50247 ;
  assign n59118 = ~n59116 & ~n59117 ;
  assign n59119 = n27325 & ~n59118 ;
  assign n59120 = \P2_buf2_reg[3]/NET0131  & n50300 ;
  assign n59121 = ~n59119 & ~n59120 ;
  assign n59122 = ~n59111 & n59121 ;
  assign n59123 = ~n59115 & n59122 ;
  assign n59126 = n26927 & n50287 ;
  assign n59125 = ~\P2_P3_InstQueue_reg[4][6]/NET0131  & ~n50287 ;
  assign n59127 = n27788 & ~n59125 ;
  assign n59128 = ~n59126 & n59127 ;
  assign n59124 = \P2_P3_InstQueue_reg[4][6]/NET0131  & ~n50290 ;
  assign n59129 = \P2_buf2_reg[30]/NET0131  & n50227 ;
  assign n59130 = \P2_buf2_reg[22]/NET0131  & n50247 ;
  assign n59131 = ~n59129 & ~n59130 ;
  assign n59132 = n27325 & ~n59131 ;
  assign n59133 = \P2_buf2_reg[6]/NET0131  & n50300 ;
  assign n59134 = ~n59132 & ~n59133 ;
  assign n59135 = ~n59124 & n59134 ;
  assign n59136 = ~n59128 & n59135 ;
  assign n59139 = n27054 & n50307 ;
  assign n59138 = ~\P2_P3_InstQueue_reg[5][3]/NET0131  & ~n50307 ;
  assign n59140 = n27788 & ~n59138 ;
  assign n59141 = ~n59139 & n59140 ;
  assign n59137 = \P2_P3_InstQueue_reg[5][3]/NET0131  & ~n50310 ;
  assign n59142 = \P2_buf2_reg[27]/NET0131  & n50247 ;
  assign n59143 = \P2_buf2_reg[19]/NET0131  & n50267 ;
  assign n59144 = ~n59142 & ~n59143 ;
  assign n59145 = n27325 & ~n59144 ;
  assign n59146 = \P2_buf2_reg[3]/NET0131  & n50320 ;
  assign n59147 = ~n59145 & ~n59146 ;
  assign n59148 = ~n59137 & n59147 ;
  assign n59149 = ~n59141 & n59148 ;
  assign n59152 = n26927 & n50307 ;
  assign n59151 = ~\P2_P3_InstQueue_reg[5][6]/NET0131  & ~n50307 ;
  assign n59153 = n27788 & ~n59151 ;
  assign n59154 = ~n59152 & n59153 ;
  assign n59150 = \P2_P3_InstQueue_reg[5][6]/NET0131  & ~n50310 ;
  assign n59155 = \P2_buf2_reg[30]/NET0131  & n50247 ;
  assign n59156 = \P2_buf2_reg[22]/NET0131  & n50267 ;
  assign n59157 = ~n59155 & ~n59156 ;
  assign n59158 = n27325 & ~n59157 ;
  assign n59159 = \P2_buf2_reg[6]/NET0131  & n50320 ;
  assign n59160 = ~n59158 & ~n59159 ;
  assign n59161 = ~n59150 & n59160 ;
  assign n59162 = ~n59154 & n59161 ;
  assign n59165 = n27054 & n50327 ;
  assign n59164 = ~\P2_P3_InstQueue_reg[6][3]/NET0131  & ~n50327 ;
  assign n59166 = n27788 & ~n59164 ;
  assign n59167 = ~n59165 & n59166 ;
  assign n59163 = \P2_P3_InstQueue_reg[6][3]/NET0131  & ~n50330 ;
  assign n59168 = \P2_buf2_reg[27]/NET0131  & n50267 ;
  assign n59169 = \P2_buf2_reg[19]/NET0131  & n50287 ;
  assign n59170 = ~n59168 & ~n59169 ;
  assign n59171 = n27325 & ~n59170 ;
  assign n59172 = \P2_buf2_reg[3]/NET0131  & n50340 ;
  assign n59173 = ~n59171 & ~n59172 ;
  assign n59174 = ~n59163 & n59173 ;
  assign n59175 = ~n59167 & n59174 ;
  assign n59178 = n26927 & n50327 ;
  assign n59177 = ~\P2_P3_InstQueue_reg[6][6]/NET0131  & ~n50327 ;
  assign n59179 = n27788 & ~n59177 ;
  assign n59180 = ~n59178 & n59179 ;
  assign n59176 = \P2_P3_InstQueue_reg[6][6]/NET0131  & ~n50330 ;
  assign n59181 = \P2_buf2_reg[30]/NET0131  & n50267 ;
  assign n59182 = \P2_buf2_reg[22]/NET0131  & n50287 ;
  assign n59183 = ~n59181 & ~n59182 ;
  assign n59184 = n27325 & ~n59183 ;
  assign n59185 = \P2_buf2_reg[6]/NET0131  & n50340 ;
  assign n59186 = ~n59184 & ~n59185 ;
  assign n59187 = ~n59176 & n59186 ;
  assign n59188 = ~n59180 & n59187 ;
  assign n59191 = n27054 & n50046 ;
  assign n59190 = ~\P2_P3_InstQueue_reg[7][3]/NET0131  & ~n50046 ;
  assign n59192 = n27788 & ~n59190 ;
  assign n59193 = ~n59191 & n59192 ;
  assign n59189 = \P2_P3_InstQueue_reg[7][3]/NET0131  & ~n50349 ;
  assign n59194 = \P2_buf2_reg[27]/NET0131  & n50287 ;
  assign n59195 = \P2_buf2_reg[19]/NET0131  & n50307 ;
  assign n59196 = ~n59194 & ~n59195 ;
  assign n59197 = n27325 & ~n59196 ;
  assign n59198 = \P2_buf2_reg[3]/NET0131  & n50359 ;
  assign n59199 = ~n59197 & ~n59198 ;
  assign n59200 = ~n59189 & n59199 ;
  assign n59201 = ~n59193 & n59200 ;
  assign n59204 = n26927 & n50046 ;
  assign n59203 = ~\P2_P3_InstQueue_reg[7][6]/NET0131  & ~n50046 ;
  assign n59205 = n27788 & ~n59203 ;
  assign n59206 = ~n59204 & n59205 ;
  assign n59202 = \P2_P3_InstQueue_reg[7][6]/NET0131  & ~n50349 ;
  assign n59207 = \P2_buf2_reg[30]/NET0131  & n50287 ;
  assign n59208 = \P2_buf2_reg[22]/NET0131  & n50307 ;
  assign n59209 = ~n59207 & ~n59208 ;
  assign n59210 = n27325 & ~n59209 ;
  assign n59211 = \P2_buf2_reg[6]/NET0131  & n50359 ;
  assign n59212 = ~n59210 & ~n59211 ;
  assign n59213 = ~n59202 & n59212 ;
  assign n59214 = ~n59206 & n59213 ;
  assign n59217 = n27054 & n50045 ;
  assign n59216 = ~\P2_P3_InstQueue_reg[8][3]/NET0131  & ~n50045 ;
  assign n59218 = n27788 & ~n59216 ;
  assign n59219 = ~n59217 & n59218 ;
  assign n59215 = \P2_P3_InstQueue_reg[8][3]/NET0131  & ~n50367 ;
  assign n59220 = \P2_buf2_reg[27]/NET0131  & n50307 ;
  assign n59221 = \P2_buf2_reg[19]/NET0131  & n50327 ;
  assign n59222 = ~n59220 & ~n59221 ;
  assign n59223 = n27325 & ~n59222 ;
  assign n59224 = \P2_buf2_reg[3]/NET0131  & n50377 ;
  assign n59225 = ~n59223 & ~n59224 ;
  assign n59226 = ~n59215 & n59225 ;
  assign n59227 = ~n59219 & n59226 ;
  assign n59230 = n26927 & n50045 ;
  assign n59229 = ~\P2_P3_InstQueue_reg[8][6]/NET0131  & ~n50045 ;
  assign n59231 = n27788 & ~n59229 ;
  assign n59232 = ~n59230 & n59231 ;
  assign n59228 = \P2_P3_InstQueue_reg[8][6]/NET0131  & ~n50367 ;
  assign n59233 = \P2_buf2_reg[30]/NET0131  & n50307 ;
  assign n59234 = \P2_buf2_reg[22]/NET0131  & n50327 ;
  assign n59235 = ~n59233 & ~n59234 ;
  assign n59236 = n27325 & ~n59235 ;
  assign n59237 = \P2_buf2_reg[6]/NET0131  & n50377 ;
  assign n59238 = ~n59236 & ~n59237 ;
  assign n59239 = ~n59228 & n59238 ;
  assign n59240 = ~n59232 & n59239 ;
  assign n59243 = n27054 & n50053 ;
  assign n59242 = ~\P2_P3_InstQueue_reg[9][3]/NET0131  & ~n50053 ;
  assign n59244 = n27788 & ~n59242 ;
  assign n59245 = ~n59243 & n59244 ;
  assign n59241 = \P2_P3_InstQueue_reg[9][3]/NET0131  & ~n50385 ;
  assign n59246 = \P2_buf2_reg[27]/NET0131  & n50327 ;
  assign n59247 = \P2_buf2_reg[19]/NET0131  & n50046 ;
  assign n59248 = ~n59246 & ~n59247 ;
  assign n59249 = n27325 & ~n59248 ;
  assign n59250 = \P2_buf2_reg[3]/NET0131  & n50395 ;
  assign n59251 = ~n59249 & ~n59250 ;
  assign n59252 = ~n59241 & n59251 ;
  assign n59253 = ~n59245 & n59252 ;
  assign n59256 = n26927 & n50053 ;
  assign n59255 = ~\P2_P3_InstQueue_reg[9][6]/NET0131  & ~n50053 ;
  assign n59257 = n27788 & ~n59255 ;
  assign n59258 = ~n59256 & n59257 ;
  assign n59254 = \P2_P3_InstQueue_reg[9][6]/NET0131  & ~n50385 ;
  assign n59259 = \P2_buf2_reg[30]/NET0131  & n50327 ;
  assign n59260 = \P2_buf2_reg[22]/NET0131  & n50046 ;
  assign n59261 = ~n59259 & ~n59260 ;
  assign n59262 = n27325 & ~n59261 ;
  assign n59263 = \P2_buf2_reg[6]/NET0131  & n50395 ;
  assign n59264 = ~n59262 & ~n59263 ;
  assign n59265 = ~n59254 & n59264 ;
  assign n59266 = ~n59258 & n59265 ;
  assign n59270 = n27308 & ~n39857 ;
  assign n59271 = ~n27315 & n27319 ;
  assign n59272 = n42870 & n59271 ;
  assign n59273 = ~n59270 & n59272 ;
  assign n59274 = \P2_P3_PhyAddrPointer_reg[0]/NET0131  & ~n59273 ;
  assign n59267 = n27284 & ~n45699 ;
  assign n59268 = ~n45703 & ~n59267 ;
  assign n59269 = n27308 & ~n59268 ;
  assign n59275 = ~n45695 & ~n59269 ;
  assign n59276 = ~n59274 & n59275 ;
  assign n59279 = n36644 & n50476 ;
  assign n59280 = n36672 & ~n59279 ;
  assign n59282 = ~n47880 & n59280 ;
  assign n59281 = n47880 & ~n59280 ;
  assign n59283 = ~\P2_P1_DataWidth_reg[1]/NET0131  & ~n59281 ;
  assign n59284 = ~n59282 & n59283 ;
  assign n59278 = \P2_P1_DataWidth_reg[1]/NET0131  & ~\P2_P1_rEIP_reg[5]/NET0131  ;
  assign n59285 = n11609 & ~n59278 ;
  assign n59286 = ~n59284 & n59285 ;
  assign n59287 = \P2_P1_rEIP_reg[5]/NET0131  & ~n50414 ;
  assign n59288 = ~\P2_P1_rEIP_reg[5]/NET0131  & ~n50766 ;
  assign n59289 = ~n50767 & ~n59288 ;
  assign n59290 = n50422 & ~n59289 ;
  assign n59291 = ~n25958 & n59290 ;
  assign n59292 = ~\P2_P1_EBX_reg[5]/NET0131  & ~n26103 ;
  assign n59293 = ~n59291 & ~n59292 ;
  assign n59294 = n24898 & n59293 ;
  assign n59295 = \P2_P1_EBX_reg[31]/NET0131  & ~n50790 ;
  assign n59297 = \P2_P1_EBX_reg[5]/NET0131  & ~n59295 ;
  assign n59296 = ~\P2_P1_EBX_reg[5]/NET0131  & n59295 ;
  assign n59298 = ~n50422 & ~n59296 ;
  assign n59299 = ~n59297 & n59298 ;
  assign n59300 = ~n59290 & ~n59299 ;
  assign n59301 = n21062 & n59300 ;
  assign n59302 = ~n59294 & ~n59301 ;
  assign n59303 = ~n21081 & ~n59302 ;
  assign n59304 = ~n59287 & ~n59303 ;
  assign n59305 = n11623 & ~n59304 ;
  assign n59277 = \P2_P1_rEIP_reg[5]/NET0131  & ~n53464 ;
  assign n59306 = \P2_P1_PhyAddrPointer_reg[5]/NET0131  & n11625 ;
  assign n59307 = ~n11616 & ~n59306 ;
  assign n59308 = ~n59277 & n59307 ;
  assign n59309 = ~n59305 & n59308 ;
  assign n59310 = ~n59286 & n59309 ;
  assign n59313 = ~n36628 & ~n53810 ;
  assign n59315 = ~n47806 & n59313 ;
  assign n59314 = n47806 & ~n59313 ;
  assign n59316 = ~\P1_P2_DataWidth_reg[1]/NET0131  & ~n59314 ;
  assign n59317 = ~n59315 & n59316 ;
  assign n59312 = \P1_P2_DataWidth_reg[1]/NET0131  & ~\P1_P2_rEIP_reg[5]/NET0131  ;
  assign n59318 = n25928 & ~n59312 ;
  assign n59319 = ~n59317 & n59318 ;
  assign n59320 = \P1_P2_rEIP_reg[5]/NET0131  & ~n48371 ;
  assign n59321 = \P1_P2_EBX_reg[31]/NET0131  & ~n48410 ;
  assign n59323 = \P1_P2_EBX_reg[5]/NET0131  & n59321 ;
  assign n59322 = ~\P1_P2_EBX_reg[5]/NET0131  & ~n59321 ;
  assign n59324 = ~n48373 & ~n59322 ;
  assign n59325 = ~n59323 & n59324 ;
  assign n59326 = ~\P1_P2_rEIP_reg[5]/NET0131  & ~n48382 ;
  assign n59327 = ~\P1_P2_DataWidth_reg[1]/NET0131  & ~n48383 ;
  assign n59328 = ~n59326 & n59327 ;
  assign n59329 = ~n25415 & n59328 ;
  assign n59330 = ~n59325 & ~n59329 ;
  assign n59331 = n25776 & ~n59330 ;
  assign n59332 = \P1_P2_EBX_reg[5]/NET0131  & ~n48443 ;
  assign n59333 = n25769 & n59328 ;
  assign n59334 = ~n59332 & ~n59333 ;
  assign n59335 = n25757 & ~n59334 ;
  assign n59336 = ~n59331 & ~n59335 ;
  assign n59337 = ~n25770 & ~n59336 ;
  assign n59338 = ~n59320 & ~n59337 ;
  assign n59339 = n25918 & ~n59338 ;
  assign n59311 = \P1_P2_rEIP_reg[5]/NET0131  & ~n53566 ;
  assign n59340 = \P1_P2_PhyAddrPointer_reg[5]/NET0131  & n27675 ;
  assign n59341 = ~n27967 & ~n59340 ;
  assign n59342 = ~n59311 & n59341 ;
  assign n59343 = ~n59339 & n59342 ;
  assign n59344 = ~n59319 & n59343 ;
  assign n59347 = n36703 & n52046 ;
  assign n59348 = ~n36733 & ~n59347 ;
  assign n59350 = n47940 & ~n59348 ;
  assign n59349 = ~n47940 & n59348 ;
  assign n59351 = ~\P1_P1_DataWidth_reg[1]/NET0131  & ~n59349 ;
  assign n59352 = ~n59350 & n59351 ;
  assign n59346 = \P1_P1_DataWidth_reg[1]/NET0131  & ~\P1_P1_rEIP_reg[5]/NET0131  ;
  assign n59353 = n8282 & ~n59346 ;
  assign n59354 = ~n59352 & n59353 ;
  assign n59355 = \P1_P1_rEIP_reg[5]/NET0131  & ~n50559 ;
  assign n59356 = ~\P1_P1_rEIP_reg[5]/NET0131  & ~n51668 ;
  assign n59357 = ~n51669 & ~n59356 ;
  assign n59358 = n26275 & ~n59357 ;
  assign n59359 = ~\P1_P1_EBX_reg[5]/NET0131  & ~n26275 ;
  assign n59360 = ~n59358 & ~n59359 ;
  assign n59361 = n24502 & n59360 ;
  assign n59362 = n26274 & ~n59357 ;
  assign n59363 = \P1_P1_EBX_reg[31]/NET0131  & ~n51689 ;
  assign n59365 = \P1_P1_EBX_reg[5]/NET0131  & ~n59363 ;
  assign n59364 = ~\P1_P1_EBX_reg[5]/NET0131  & n59363 ;
  assign n59366 = ~n26274 & ~n59364 ;
  assign n59367 = ~n59365 & n59366 ;
  assign n59368 = ~n59362 & ~n59367 ;
  assign n59369 = n15334 & n59368 ;
  assign n59370 = ~n59361 & ~n59369 ;
  assign n59371 = ~n15364 & ~n59370 ;
  assign n59372 = ~n59355 & ~n59371 ;
  assign n59373 = n8355 & ~n59372 ;
  assign n59345 = \P1_P1_rEIP_reg[5]/NET0131  & ~n53883 ;
  assign n59374 = \P1_P1_PhyAddrPointer_reg[5]/NET0131  & n8361 ;
  assign n59375 = ~n8357 & ~n59374 ;
  assign n59376 = ~n59345 & n59375 ;
  assign n59377 = ~n59373 & n59376 ;
  assign n59378 = ~n59354 & n59377 ;
  assign n59381 = n36762 & n52485 ;
  assign n59382 = n36792 & ~n59381 ;
  assign n59384 = n47983 & ~n59382 ;
  assign n59383 = ~n47983 & n59382 ;
  assign n59385 = ~\P2_P2_DataWidth_reg[1]/NET0131  & ~n59383 ;
  assign n59386 = ~n59384 & n59385 ;
  assign n59380 = \P2_P2_DataWidth_reg[1]/NET0131  & ~\P2_P2_rEIP_reg[5]/NET0131  ;
  assign n59387 = n26794 & ~n59380 ;
  assign n59388 = ~n59386 & n59387 ;
  assign n59389 = \P2_P2_rEIP_reg[5]/NET0131  & ~n50640 ;
  assign n59390 = ~\P2_P2_rEIP_reg[5]/NET0131  & ~n52095 ;
  assign n59391 = ~n52096 & ~n59390 ;
  assign n59392 = n50649 & ~n59391 ;
  assign n59393 = ~n26650 & n59392 ;
  assign n59394 = ~\P2_P2_EBX_reg[5]/NET0131  & ~n50642 ;
  assign n59395 = ~n59393 & ~n59394 ;
  assign n59396 = n26786 & n59395 ;
  assign n59397 = \P2_P2_EBX_reg[31]/NET0131  & ~n52116 ;
  assign n59399 = \P2_P2_EBX_reg[5]/NET0131  & ~n59397 ;
  assign n59398 = ~\P2_P2_EBX_reg[5]/NET0131  & n59397 ;
  assign n59400 = ~n50649 & ~n59398 ;
  assign n59401 = ~n59399 & n59400 ;
  assign n59402 = ~n59392 & ~n59401 ;
  assign n59403 = n47684 & n59402 ;
  assign n59404 = ~n59396 & ~n59403 ;
  assign n59405 = ~n59389 & n59404 ;
  assign n59406 = n26792 & ~n59405 ;
  assign n59379 = \P2_P2_rEIP_reg[5]/NET0131  & ~n54099 ;
  assign n59407 = \P2_P2_PhyAddrPointer_reg[5]/NET0131  & n27637 ;
  assign n59408 = ~n28046 & ~n59407 ;
  assign n59409 = ~n59379 & n59408 ;
  assign n59410 = ~n59406 & n59409 ;
  assign n59411 = ~n59388 & n59410 ;
  assign n59414 = n36836 & n50708 ;
  assign n59415 = ~n36863 & ~n59414 ;
  assign n59417 = ~n48107 & n59415 ;
  assign n59416 = n48107 & ~n59415 ;
  assign n59418 = ~\P2_P3_DataWidth_reg[1]/NET0131  & ~n59416 ;
  assign n59419 = ~n59417 & n59418 ;
  assign n59413 = \P2_P3_DataWidth_reg[1]/NET0131  & ~\P2_P3_rEIP_reg[5]/NET0131  ;
  assign n59420 = n27315 & ~n59413 ;
  assign n59421 = ~n59419 & n59420 ;
  assign n59429 = ~\P2_P3_rEIP_reg[5]/NET0131  & ~n52549 ;
  assign n59430 = ~n52550 & ~n59429 ;
  assign n59431 = n56676 & n59430 ;
  assign n59424 = \P2_P3_EBX_reg[31]/NET0131  & ~n52525 ;
  assign n59425 = ~\P2_P3_EBX_reg[5]/NET0131  & ~n59424 ;
  assign n59426 = \P2_P3_EBX_reg[5]/NET0131  & n59424 ;
  assign n59427 = ~n59425 & ~n59426 ;
  assign n59428 = n56679 & n59427 ;
  assign n59422 = \P2_P3_rEIP_reg[5]/NET0131  & ~n27277 ;
  assign n59423 = \P2_P3_EBX_reg[5]/NET0131  & n56680 ;
  assign n59432 = ~n59422 & ~n59423 ;
  assign n59433 = ~n59428 & n59432 ;
  assign n59434 = ~n59431 & n59433 ;
  assign n59435 = n27308 & ~n59434 ;
  assign n59412 = \P2_P3_rEIP_reg[5]/NET0131  & ~n54653 ;
  assign n59436 = \P2_P3_PhyAddrPointer_reg[5]/NET0131  & n27651 ;
  assign n59437 = ~n32864 & ~n59436 ;
  assign n59438 = ~n59412 & n59437 ;
  assign n59439 = ~n59435 & n59438 ;
  assign n59440 = ~n59421 & n59439 ;
  assign n59442 = \P1_P2_PhyAddrPointer_reg[1]/NET0131  & ~n39340 ;
  assign n59443 = n46153 & ~n59442 ;
  assign n59444 = n25918 & ~n59443 ;
  assign n59445 = ~n25933 & n39352 ;
  assign n59446 = \P1_P2_PhyAddrPointer_reg[1]/NET0131  & ~n59445 ;
  assign n59441 = ~\P1_P2_PhyAddrPointer_reg[1]/NET0131  & n36630 ;
  assign n59447 = ~n46126 & ~n59441 ;
  assign n59448 = ~n59446 & n59447 ;
  assign n59449 = ~n59444 & n59448 ;
  assign n59450 = \P2_P1_PhyAddrPointer_reg[1]/NET0131  & ~n36678 ;
  assign n59451 = n45290 & ~n59450 ;
  assign n59452 = n11623 & ~n59451 ;
  assign n59453 = ~\P2_P1_PhyAddrPointer_reg[1]/NET0131  & ~n36674 ;
  assign n59454 = \P2_P1_PhyAddrPointer_reg[1]/NET0131  & ~n11624 ;
  assign n59455 = n50409 & n59454 ;
  assign n59456 = ~n27681 & n59455 ;
  assign n59457 = ~n59453 & ~n59456 ;
  assign n59458 = ~n45272 & ~n59457 ;
  assign n59459 = ~n59452 & n59458 ;
  assign n59460 = \P1_P1_PhyAddrPointer_reg[1]/NET0131  & ~n41658 ;
  assign n59461 = n45898 & ~n59460 ;
  assign n59462 = n8355 & ~n59461 ;
  assign n59463 = ~\P1_P1_PhyAddrPointer_reg[1]/NET0131  & n36701 ;
  assign n59464 = \P1_P1_PhyAddrPointer_reg[1]/NET0131  & ~n8349 ;
  assign n59465 = n50581 & n59464 ;
  assign n59466 = ~n27791 & n59465 ;
  assign n59467 = ~n59463 & ~n59466 ;
  assign n59468 = ~n45878 & ~n59467 ;
  assign n59469 = ~n59462 & n59468 ;
  assign n59471 = \P2_P2_PhyAddrPointer_reg[1]/NET0131  & ~n41873 ;
  assign n59472 = n45522 & ~n59471 ;
  assign n59473 = n26792 & ~n59472 ;
  assign n59474 = ~n26800 & n36758 ;
  assign n59475 = \P2_P2_PhyAddrPointer_reg[1]/NET0131  & ~n59474 ;
  assign n59470 = ~\P2_P2_PhyAddrPointer_reg[1]/NET0131  & ~n36760 ;
  assign n59476 = ~n45489 & ~n59470 ;
  assign n59477 = ~n59475 & n59476 ;
  assign n59478 = ~n59473 & n59477 ;
  assign n59480 = \P1_P3_PhyAddrPointer_reg[1]/NET0131  & ~n37992 ;
  assign n59481 = n18430 & ~n59480 ;
  assign n59482 = n9241 & ~n59481 ;
  assign n59483 = ~n11698 & n36816 ;
  assign n59484 = \P1_P3_PhyAddrPointer_reg[1]/NET0131  & ~n59483 ;
  assign n59479 = ~\P1_P3_PhyAddrPointer_reg[1]/NET0131  & ~n36810 ;
  assign n59485 = ~n18339 & ~n59479 ;
  assign n59486 = ~n59484 & n59485 ;
  assign n59487 = ~n59482 & n59486 ;
  assign n59490 = \P2_P3_PhyAddrPointer_reg[1]/NET0131  & ~n39857 ;
  assign n59489 = n27284 & ~n45727 ;
  assign n59491 = ~n45738 & ~n59489 ;
  assign n59492 = ~n59490 & n59491 ;
  assign n59493 = n27308 & ~n59492 ;
  assign n59494 = ~n27325 & n36873 ;
  assign n59495 = \P2_P3_PhyAddrPointer_reg[1]/NET0131  & ~n59494 ;
  assign n59488 = ~\P2_P3_PhyAddrPointer_reg[1]/NET0131  & ~n36831 ;
  assign n59496 = ~n45713 & ~n59488 ;
  assign n59497 = ~n59495 & n59496 ;
  assign n59498 = ~n59493 & n59497 ;
  assign n59500 = ~n26158 & ~n57485 ;
  assign n59501 = n24503 & ~n59500 ;
  assign n59502 = n53011 & ~n59501 ;
  assign n59503 = \P1_P1_Datao_reg[19]/NET0131  & ~n59502 ;
  assign n59504 = ~n26158 & n57486 ;
  assign n59505 = ~n59503 & ~n59504 ;
  assign n59506 = n8355 & ~n59505 ;
  assign n59499 = \P1_P1_uWord_reg[3]/NET0131  & n27790 ;
  assign n59507 = \P1_P1_Datao_reg[19]/NET0131  & ~n48479 ;
  assign n59508 = ~n59499 & ~n59507 ;
  assign n59509 = ~n59506 & n59508 ;
  assign n59511 = ~n26158 & ~n40738 ;
  assign n59512 = n24503 & ~n59511 ;
  assign n59513 = n53011 & ~n59512 ;
  assign n59514 = \P1_P1_Datao_reg[23]/NET0131  & ~n59513 ;
  assign n59515 = ~n26158 & n40739 ;
  assign n59516 = ~n59514 & ~n59515 ;
  assign n59517 = n8355 & ~n59516 ;
  assign n59510 = \P1_P1_uWord_reg[7]/NET0131  & n27790 ;
  assign n59518 = \P1_P1_Datao_reg[23]/NET0131  & ~n48479 ;
  assign n59519 = ~n59510 & ~n59518 ;
  assign n59520 = ~n59517 & n59519 ;
  assign n59522 = ~n26699 & n26792 ;
  assign n59523 = n48508 & ~n59522 ;
  assign n59524 = \P2_P2_Datao_reg[19]/NET0131  & ~n59523 ;
  assign n59521 = \P2_P2_uWord_reg[3]/NET0131  & n48491 ;
  assign n59525 = ~\P2_P2_EAX_reg[19]/NET0131  & ~n47662 ;
  assign n59526 = ~n47663 & ~n59525 ;
  assign n59527 = n26643 & n59526 ;
  assign n59528 = n26692 & n26792 ;
  assign n59529 = n59527 & n59528 ;
  assign n59530 = ~n59521 & ~n59529 ;
  assign n59531 = ~n59524 & n59530 ;
  assign n59533 = \P2_P2_Datao_reg[23]/NET0131  & ~n26699 ;
  assign n59534 = ~\P2_P2_EAX_reg[23]/NET0131  & ~n47666 ;
  assign n59535 = n26643 & ~n47667 ;
  assign n59536 = ~n59534 & n59535 ;
  assign n59537 = n26692 & n59536 ;
  assign n59538 = ~n59533 & ~n59537 ;
  assign n59539 = n26792 & ~n59538 ;
  assign n59532 = \P2_P2_uWord_reg[7]/NET0131  & n48491 ;
  assign n59540 = \P2_P2_Datao_reg[23]/NET0131  & ~n48508 ;
  assign n59541 = ~n59532 & ~n59540 ;
  assign n59542 = ~n59539 & n59541 ;
  assign n59544 = \P2_P3_Datao_reg[19]/NET0131  & ~n56850 ;
  assign n59543 = \P2_P3_uWord_reg[3]/NET0131  & n48523 ;
  assign n59545 = ~\P2_P3_EAX_reg[19]/NET0131  & ~n47775 ;
  assign n59546 = ~n47776 & ~n59545 ;
  assign n59547 = n47747 & n59546 ;
  assign n59548 = n56841 & n59547 ;
  assign n59549 = ~n59543 & ~n59548 ;
  assign n59550 = ~n59544 & n59549 ;
  assign n59552 = \P2_P3_Datao_reg[23]/NET0131  & ~n27223 ;
  assign n59553 = ~\P2_P3_EAX_reg[23]/NET0131  & ~n48528 ;
  assign n59554 = n27121 & ~n48529 ;
  assign n59555 = ~n59553 & n59554 ;
  assign n59556 = n27178 & n59555 ;
  assign n59557 = ~n59552 & ~n59556 ;
  assign n59558 = n27308 & ~n59557 ;
  assign n59551 = \P2_P3_uWord_reg[7]/NET0131  & n48523 ;
  assign n59559 = \P2_P3_Datao_reg[23]/NET0131  & ~n48540 ;
  assign n59560 = ~n59551 & ~n59559 ;
  assign n59561 = ~n59558 & n59560 ;
  assign n59563 = ~\P1_P2_EAX_reg[19]/NET0131  & ~n47549 ;
  assign n59564 = ~n47550 & ~n59563 ;
  assign n59565 = n47570 & n59564 ;
  assign n59566 = ~n25768 & n59565 ;
  assign n59567 = \P1_P2_Datao_reg[19]/NET0131  & ~n25847 ;
  assign n59568 = ~n59566 & ~n59567 ;
  assign n59569 = n25918 & ~n59568 ;
  assign n59562 = \P1_P2_uWord_reg[3]/NET0131  & n25922 ;
  assign n59570 = \P1_P2_Datao_reg[19]/NET0131  & ~n48566 ;
  assign n59571 = ~n59562 & ~n59570 ;
  assign n59572 = ~n59569 & n59571 ;
  assign n59574 = \P1_P2_Datao_reg[23]/NET0131  & ~n25847 ;
  assign n59575 = ~\P1_P2_EAX_reg[23]/NET0131  & ~n47553 ;
  assign n59576 = ~n47554 & n47570 ;
  assign n59577 = ~n59575 & n59576 ;
  assign n59578 = ~n25768 & n59577 ;
  assign n59579 = ~n59574 & ~n59578 ;
  assign n59580 = n25918 & ~n59579 ;
  assign n59573 = \P1_P2_uWord_reg[7]/NET0131  & n25922 ;
  assign n59581 = \P1_P2_Datao_reg[23]/NET0131  & ~n48566 ;
  assign n59582 = ~n59573 & ~n59581 ;
  assign n59583 = ~n59580 & n59582 ;
  assign n59585 = ~n25958 & ~n57003 ;
  assign n59586 = n24899 & ~n59585 ;
  assign n59587 = n48584 & ~n59586 ;
  assign n59588 = \P2_P1_Datao_reg[19]/NET0131  & ~n59587 ;
  assign n59589 = ~n25958 & n57004 ;
  assign n59590 = ~n59588 & ~n59589 ;
  assign n59591 = n11623 & ~n59590 ;
  assign n59584 = \P2_P1_uWord_reg[3]/NET0131  & n48581 ;
  assign n59592 = \P2_P1_Datao_reg[19]/NET0131  & ~n48594 ;
  assign n59593 = ~n59584 & ~n59592 ;
  assign n59594 = ~n59591 & n59593 ;
  assign n59596 = ~n25958 & ~n40723 ;
  assign n59597 = n24899 & ~n59596 ;
  assign n59598 = n48584 & ~n59597 ;
  assign n59599 = \P2_P1_Datao_reg[23]/NET0131  & ~n59598 ;
  assign n59600 = n26006 & n40724 ;
  assign n59601 = ~n59599 & ~n59600 ;
  assign n59602 = n11623 & ~n59601 ;
  assign n59595 = \P2_P1_uWord_reg[7]/NET0131  & n48581 ;
  assign n59603 = \P2_P1_Datao_reg[23]/NET0131  & ~n48594 ;
  assign n59604 = ~n59595 & ~n59603 ;
  assign n59605 = ~n59602 & n59604 ;
  assign n59608 = ~\P1_P2_EBX_reg[18]/NET0131  & ~n46714 ;
  assign n59609 = n25803 & ~n46715 ;
  assign n59610 = ~n59608 & n59609 ;
  assign n59606 = \P1_P2_EBX_reg[18]/NET0131  & n46695 ;
  assign n59607 = n46694 & ~n58110 ;
  assign n59611 = ~n59606 & ~n59607 ;
  assign n59612 = ~n59610 & n59611 ;
  assign n59613 = n25918 & ~n59612 ;
  assign n59614 = \P1_P2_EBX_reg[18]/NET0131  & ~n43212 ;
  assign n59615 = ~n59613 & ~n59614 ;
  assign n59617 = \P2_P1_EBX_reg[10]/NET0131  & n46227 ;
  assign n59616 = ~n27470 & n46225 ;
  assign n59618 = ~\P2_P1_EBX_reg[10]/NET0131  & ~n46238 ;
  assign n59619 = ~n46239 & ~n59618 ;
  assign n59620 = n25981 & n59619 ;
  assign n59621 = ~n59616 & ~n59620 ;
  assign n59622 = ~n59617 & n59621 ;
  assign n59623 = n11623 & ~n59622 ;
  assign n59624 = \P2_P1_EBX_reg[10]/NET0131  & ~n21100 ;
  assign n59625 = ~n59623 & ~n59624 ;
  assign n59627 = \P2_P1_EBX_reg[11]/NET0131  & n46227 ;
  assign n59626 = ~n25405 & n46225 ;
  assign n59628 = ~\P2_P1_EBX_reg[11]/NET0131  & ~n46239 ;
  assign n59629 = n25981 & ~n46240 ;
  assign n59630 = ~n59628 & n59629 ;
  assign n59631 = ~n59626 & ~n59630 ;
  assign n59632 = ~n59627 & n59631 ;
  assign n59633 = n11623 & ~n59632 ;
  assign n59634 = \P2_P1_EBX_reg[11]/NET0131  & ~n21100 ;
  assign n59635 = ~n59633 & ~n59634 ;
  assign n59636 = \P2_P1_EBX_reg[12]/NET0131  & ~n21100 ;
  assign n59638 = ~n46227 & ~n59629 ;
  assign n59639 = \P2_P1_EBX_reg[12]/NET0131  & ~n59638 ;
  assign n59637 = ~n25208 & n46225 ;
  assign n59640 = ~\P2_P1_EBX_reg[12]/NET0131  & n25981 ;
  assign n59641 = n46240 & n59640 ;
  assign n59642 = ~n59637 & ~n59641 ;
  assign n59643 = ~n59639 & n59642 ;
  assign n59644 = n11623 & ~n59643 ;
  assign n59645 = ~n59636 & ~n59644 ;
  assign n59648 = ~\P2_P1_EBX_reg[13]/NET0131  & ~n46241 ;
  assign n59649 = n25981 & ~n46242 ;
  assign n59650 = ~n59648 & n59649 ;
  assign n59646 = \P2_P1_EBX_reg[13]/NET0131  & n46227 ;
  assign n59647 = ~n25096 & n46225 ;
  assign n59651 = ~n59646 & ~n59647 ;
  assign n59652 = ~n59650 & n59651 ;
  assign n59653 = n11623 & ~n59652 ;
  assign n59654 = \P2_P1_EBX_reg[13]/NET0131  & ~n21100 ;
  assign n59655 = ~n59653 & ~n59654 ;
  assign n59658 = ~\P2_P1_EBX_reg[14]/NET0131  & ~n46242 ;
  assign n59659 = n25981 & ~n46243 ;
  assign n59660 = ~n59658 & n59659 ;
  assign n59656 = ~n24745 & n46225 ;
  assign n59657 = \P2_P1_EBX_reg[14]/NET0131  & n46227 ;
  assign n59661 = ~n59656 & ~n59657 ;
  assign n59662 = ~n59660 & n59661 ;
  assign n59663 = n11623 & ~n59662 ;
  assign n59664 = \P2_P1_EBX_reg[14]/NET0131  & ~n21100 ;
  assign n59665 = ~n59663 & ~n59664 ;
  assign n59668 = ~\P2_P1_EBX_reg[15]/NET0131  & ~n46243 ;
  assign n59669 = n25981 & ~n46244 ;
  assign n59670 = ~n59668 & n59669 ;
  assign n59666 = ~n24789 & n46225 ;
  assign n59667 = \P2_P1_EBX_reg[15]/NET0131  & n46227 ;
  assign n59671 = ~n59666 & ~n59667 ;
  assign n59672 = ~n59670 & n59671 ;
  assign n59673 = n11623 & ~n59672 ;
  assign n59674 = \P2_P1_EBX_reg[15]/NET0131  & ~n21100 ;
  assign n59675 = ~n59673 & ~n59674 ;
  assign n59678 = ~\P2_P1_EBX_reg[16]/NET0131  & ~n46244 ;
  assign n59679 = n25981 & ~n46245 ;
  assign n59680 = ~n59678 & n59679 ;
  assign n59676 = ~n25248 & n46225 ;
  assign n59677 = \P2_P1_EBX_reg[16]/NET0131  & n46227 ;
  assign n59681 = ~n59676 & ~n59677 ;
  assign n59682 = ~n59680 & n59681 ;
  assign n59683 = n11623 & ~n59682 ;
  assign n59684 = \P2_P1_EBX_reg[16]/NET0131  & ~n21100 ;
  assign n59685 = ~n59683 & ~n59684 ;
  assign n59688 = ~\P2_P1_EBX_reg[17]/NET0131  & ~n46245 ;
  assign n59689 = n25981 & ~n46246 ;
  assign n59690 = ~n59688 & n59689 ;
  assign n59686 = \P2_P1_EBX_reg[17]/NET0131  & n46227 ;
  assign n59687 = ~n25134 & n46225 ;
  assign n59691 = ~n59686 & ~n59687 ;
  assign n59692 = ~n59690 & n59691 ;
  assign n59693 = n11623 & ~n59692 ;
  assign n59694 = \P2_P1_EBX_reg[17]/NET0131  & ~n21100 ;
  assign n59695 = ~n59693 & ~n59694 ;
  assign n59698 = ~\P2_P1_EBX_reg[18]/NET0131  & ~n46246 ;
  assign n59699 = n25981 & ~n46247 ;
  assign n59700 = ~n59698 & n59699 ;
  assign n59696 = \P2_P1_EBX_reg[18]/NET0131  & n46227 ;
  assign n59697 = ~n24828 & n46225 ;
  assign n59701 = ~n59696 & ~n59697 ;
  assign n59702 = ~n59700 & n59701 ;
  assign n59703 = n11623 & ~n59702 ;
  assign n59704 = \P2_P1_EBX_reg[18]/NET0131  & ~n21100 ;
  assign n59705 = ~n59703 & ~n59704 ;
  assign n59708 = ~\P2_P1_EBX_reg[19]/NET0131  & ~n46247 ;
  assign n59709 = n25981 & ~n46248 ;
  assign n59710 = ~n59708 & n59709 ;
  assign n59706 = \P2_P1_EBX_reg[19]/NET0131  & n46227 ;
  assign n59707 = ~n24480 & n46225 ;
  assign n59711 = ~n59706 & ~n59707 ;
  assign n59712 = ~n59710 & n59711 ;
  assign n59713 = n11623 & ~n59712 ;
  assign n59714 = \P2_P1_EBX_reg[19]/NET0131  & ~n21100 ;
  assign n59715 = ~n59713 & ~n59714 ;
  assign n59718 = ~\P2_P1_EBX_reg[20]/NET0131  & ~n46248 ;
  assign n59719 = n25981 & ~n46249 ;
  assign n59720 = ~n59718 & n59719 ;
  assign n59716 = \P2_P1_EBX_reg[20]/NET0131  & n46227 ;
  assign n59717 = ~n24878 & n46225 ;
  assign n59721 = ~n59716 & ~n59717 ;
  assign n59722 = ~n59720 & n59721 ;
  assign n59723 = n11623 & ~n59722 ;
  assign n59724 = \P2_P1_EBX_reg[20]/NET0131  & ~n21100 ;
  assign n59725 = ~n59723 & ~n59724 ;
  assign n59728 = ~\P2_P1_EBX_reg[21]/NET0131  & ~n46249 ;
  assign n59729 = n25981 & ~n46250 ;
  assign n59730 = ~n59728 & n59729 ;
  assign n59726 = \P2_P1_EBX_reg[21]/NET0131  & n46227 ;
  assign n59727 = ~n24240 & n46225 ;
  assign n59731 = ~n59726 & ~n59727 ;
  assign n59732 = ~n59730 & n59731 ;
  assign n59733 = n11623 & ~n59732 ;
  assign n59734 = \P2_P1_EBX_reg[21]/NET0131  & ~n21100 ;
  assign n59735 = ~n59733 & ~n59734 ;
  assign n59738 = ~\P2_P1_EBX_reg[22]/NET0131  & ~n46250 ;
  assign n59739 = n25981 & ~n46251 ;
  assign n59740 = ~n59738 & n59739 ;
  assign n59736 = \P2_P1_EBX_reg[22]/NET0131  & n46227 ;
  assign n59737 = ~n24290 & n46225 ;
  assign n59741 = ~n59736 & ~n59737 ;
  assign n59742 = ~n59740 & n59741 ;
  assign n59743 = n11623 & ~n59742 ;
  assign n59744 = \P2_P1_EBX_reg[22]/NET0131  & ~n21100 ;
  assign n59745 = ~n59743 & ~n59744 ;
  assign n59748 = ~\P2_P1_EBX_reg[23]/NET0131  & ~n46251 ;
  assign n59749 = n25981 & ~n46252 ;
  assign n59750 = ~n59748 & n59749 ;
  assign n59746 = n24104 & n46225 ;
  assign n59747 = \P2_P1_EBX_reg[23]/NET0131  & n46227 ;
  assign n59751 = ~n59746 & ~n59747 ;
  assign n59752 = ~n59750 & n59751 ;
  assign n59753 = n11623 & ~n59752 ;
  assign n59754 = \P2_P1_EBX_reg[23]/NET0131  & ~n21100 ;
  assign n59755 = ~n59753 & ~n59754 ;
  assign n59758 = ~\P2_P1_EBX_reg[24]/NET0131  & ~n46252 ;
  assign n59759 = n25981 & ~n46253 ;
  assign n59760 = ~n59758 & n59759 ;
  assign n59756 = n23728 & n46225 ;
  assign n59757 = \P2_P1_EBX_reg[24]/NET0131  & n46227 ;
  assign n59761 = ~n59756 & ~n59757 ;
  assign n59762 = ~n59760 & n59761 ;
  assign n59763 = n11623 & ~n59762 ;
  assign n59764 = \P2_P1_EBX_reg[24]/NET0131  & ~n21100 ;
  assign n59765 = ~n59763 & ~n59764 ;
  assign n59768 = ~\P2_P1_EBX_reg[28]/NET0131  & ~n46257 ;
  assign n59769 = n25981 & ~n46267 ;
  assign n59770 = ~n59768 & n59769 ;
  assign n59766 = \P2_P1_EBX_reg[28]/NET0131  & n46227 ;
  assign n59767 = n22795 & n46225 ;
  assign n59771 = ~n59766 & ~n59767 ;
  assign n59772 = ~n59770 & n59771 ;
  assign n59773 = n11623 & ~n59772 ;
  assign n59774 = \P2_P1_EBX_reg[28]/NET0131  & ~n21100 ;
  assign n59775 = ~n59773 & ~n59774 ;
  assign n59777 = \P2_P1_EBX_reg[8]/NET0131  & n46227 ;
  assign n59776 = ~n27716 & n46225 ;
  assign n59778 = ~\P2_P1_EBX_reg[8]/NET0131  & ~n46236 ;
  assign n59779 = ~n46237 & ~n59778 ;
  assign n59780 = n25981 & n59779 ;
  assign n59781 = ~n59776 & ~n59780 ;
  assign n59782 = ~n59777 & n59781 ;
  assign n59783 = n11623 & ~n59782 ;
  assign n59784 = \P2_P1_EBX_reg[8]/NET0131  & ~n21100 ;
  assign n59785 = ~n59783 & ~n59784 ;
  assign n59787 = \P2_P1_EBX_reg[9]/NET0131  & n46227 ;
  assign n59786 = ~n27524 & n46225 ;
  assign n59788 = ~\P2_P1_EBX_reg[9]/NET0131  & ~n46237 ;
  assign n59789 = ~n46238 & ~n59788 ;
  assign n59790 = n25981 & n59789 ;
  assign n59791 = ~n59786 & ~n59790 ;
  assign n59792 = ~n59787 & n59791 ;
  assign n59793 = n11623 & ~n59792 ;
  assign n59794 = \P2_P1_EBX_reg[9]/NET0131  & ~n21100 ;
  assign n59795 = ~n59793 & ~n59794 ;
  assign n59796 = n11623 & ~n25966 ;
  assign n59797 = \P2_P1_Flush_reg/NET0131  & ~n21100 ;
  assign n59798 = ~n59796 & ~n59797 ;
  assign n59799 = ~n25883 & n25918 ;
  assign n59800 = \P1_P2_Flush_reg/NET0131  & ~n43212 ;
  assign n59801 = ~n59799 & ~n59800 ;
  assign n59802 = \P2_P1_uWord_reg[0]/NET0131  & ~n25156 ;
  assign n59803 = ~\P2_P1_EAX_reg[16]/NET0131  & ~n27387 ;
  assign n59804 = ~n27388 & ~n59803 ;
  assign n59805 = n24899 & n59804 ;
  assign n59806 = n21062 & n25254 ;
  assign n59807 = ~n59805 & ~n59806 ;
  assign n59808 = n11623 & ~n59807 ;
  assign n59809 = ~n59802 & ~n59808 ;
  assign n59810 = \P2_P1_uWord_reg[1]/NET0131  & ~n24913 ;
  assign n59814 = \P2_P1_uWord_reg[1]/NET0131  & ~n25154 ;
  assign n59811 = ~\P2_P1_EAX_reg[17]/NET0131  & ~n27388 ;
  assign n59812 = ~n27389 & ~n59811 ;
  assign n59813 = n24899 & n59812 ;
  assign n59815 = n21062 & n25140 ;
  assign n59816 = ~n59813 & ~n59815 ;
  assign n59817 = ~n59814 & n59816 ;
  assign n59818 = n11623 & ~n59817 ;
  assign n59819 = ~n59810 & ~n59818 ;
  assign n59820 = \P2_P1_uWord_reg[2]/NET0131  & ~n25156 ;
  assign n59821 = ~\P2_P1_EAX_reg[18]/NET0131  & ~n27389 ;
  assign n59822 = ~n27390 & ~n59821 ;
  assign n59823 = n24899 & n59822 ;
  assign n59824 = ~n53109 & ~n59823 ;
  assign n59825 = n11623 & ~n59824 ;
  assign n59826 = ~n59820 & ~n59825 ;
  assign n59827 = \P1_P2_uWord_reg[0]/NET0131  & ~n47529 ;
  assign n59828 = \P1_P2_uWord_reg[0]/NET0131  & ~n47572 ;
  assign n59829 = ~\P1_P2_EAX_reg[16]/NET0131  & ~n47546 ;
  assign n59830 = ~n47547 & ~n59829 ;
  assign n59831 = n47570 & n59830 ;
  assign n59832 = ~n56902 & ~n59831 ;
  assign n59833 = ~n59828 & n59832 ;
  assign n59834 = n25918 & ~n59833 ;
  assign n59835 = ~n59827 & ~n59834 ;
  assign n59836 = \P1_P2_uWord_reg[10]/NET0131  & ~n53114 ;
  assign n59837 = n25776 & n47732 ;
  assign n59838 = ~\P1_P2_EAX_reg[26]/NET0131  & ~n47556 ;
  assign n59839 = n25757 & ~n47557 ;
  assign n59840 = ~n59838 & n59839 ;
  assign n59841 = ~n59837 & ~n59840 ;
  assign n59842 = n56940 & ~n59841 ;
  assign n59843 = ~n59836 & ~n59842 ;
  assign n59844 = \P1_P2_uWord_reg[13]/NET0131  & ~n47529 ;
  assign n59846 = ~\P1_P2_EAX_reg[29]/NET0131  & ~n47560 ;
  assign n59845 = \P1_P2_EAX_reg[29]/NET0131  & n47560 ;
  assign n59847 = n47570 & ~n59845 ;
  assign n59848 = ~n59846 & n59847 ;
  assign n59849 = \P1_P2_uWord_reg[13]/NET0131  & n56897 ;
  assign n59850 = ~n56926 & ~n59849 ;
  assign n59851 = ~n59848 & n59850 ;
  assign n59852 = n25918 & ~n59851 ;
  assign n59853 = ~n59844 & ~n59852 ;
  assign n59854 = \P1_P2_uWord_reg[14]/NET0131  & ~n47529 ;
  assign n59855 = n25776 & n46684 ;
  assign n59856 = \P1_P2_EAX_reg[30]/NET0131  & ~n59845 ;
  assign n59857 = ~\P1_P2_EAX_reg[30]/NET0131  & n59845 ;
  assign n59858 = ~n59856 & ~n59857 ;
  assign n59859 = n25757 & ~n59858 ;
  assign n59860 = ~n59855 & ~n59859 ;
  assign n59861 = ~n25770 & ~n59860 ;
  assign n59862 = \P1_P2_uWord_reg[14]/NET0131  & ~n47572 ;
  assign n59863 = ~n59861 & ~n59862 ;
  assign n59864 = n25918 & ~n59863 ;
  assign n59865 = ~n59854 & ~n59864 ;
  assign n59866 = \P1_P2_uWord_reg[1]/NET0131  & ~n47529 ;
  assign n59870 = \P1_P2_uWord_reg[1]/NET0131  & ~n47572 ;
  assign n59867 = ~\P1_P2_EAX_reg[17]/NET0131  & ~n47547 ;
  assign n59868 = ~n47548 & ~n59867 ;
  assign n59869 = n47570 & n59868 ;
  assign n59871 = ~n56945 & ~n59869 ;
  assign n59872 = ~n59870 & n59871 ;
  assign n59873 = n25918 & ~n59872 ;
  assign n59874 = ~n59866 & ~n59873 ;
  assign n59875 = \P1_P2_uWord_reg[2]/NET0131  & ~n47529 ;
  assign n59879 = \P1_P2_uWord_reg[2]/NET0131  & n47571 ;
  assign n59876 = ~\P1_P2_EAX_reg[18]/NET0131  & ~n47548 ;
  assign n59877 = ~n47549 & ~n59876 ;
  assign n59878 = n47570 & n59877 ;
  assign n59880 = \P1_P2_uWord_reg[2]/NET0131  & n25415 ;
  assign n59881 = ~n53383 & ~n59880 ;
  assign n59882 = n25776 & ~n59881 ;
  assign n59883 = ~n59878 & ~n59882 ;
  assign n59884 = ~n59879 & n59883 ;
  assign n59885 = n25918 & ~n59884 ;
  assign n59886 = ~n59875 & ~n59885 ;
  assign n59887 = \P1_P2_uWord_reg[3]/NET0131  & ~n47529 ;
  assign n59888 = \P1_P2_uWord_reg[3]/NET0131  & n47571 ;
  assign n59889 = \P1_P2_uWord_reg[3]/NET0131  & n25415 ;
  assign n59890 = ~n53394 & ~n59889 ;
  assign n59891 = n25776 & ~n59890 ;
  assign n59892 = ~n59565 & ~n59891 ;
  assign n59893 = ~n59888 & n59892 ;
  assign n59894 = n25918 & ~n59893 ;
  assign n59895 = ~n59887 & ~n59894 ;
  assign n59896 = \P1_P2_uWord_reg[5]/NET0131  & ~n53114 ;
  assign n59897 = ~\P1_P2_EAX_reg[21]/NET0131  & ~n47551 ;
  assign n59898 = ~n47552 & ~n59897 ;
  assign n59899 = n47570 & n59898 ;
  assign n59900 = ~n56969 & ~n59899 ;
  assign n59901 = n25918 & ~n59900 ;
  assign n59902 = ~n59896 & ~n59901 ;
  assign n59903 = \P1_P2_uWord_reg[6]/NET0131  & ~n47529 ;
  assign n59904 = \P1_P2_uWord_reg[6]/NET0131  & ~n47572 ;
  assign n59905 = ~\P1_P2_EAX_reg[22]/NET0131  & ~n47552 ;
  assign n59906 = ~n47553 & ~n59905 ;
  assign n59907 = n47570 & n59906 ;
  assign n59908 = ~n56976 & ~n59907 ;
  assign n59909 = ~n59904 & n59908 ;
  assign n59910 = n25918 & ~n59909 ;
  assign n59911 = ~n59903 & ~n59910 ;
  assign n59912 = \P1_P2_uWord_reg[7]/NET0131  & ~n47529 ;
  assign n59913 = \P1_P2_uWord_reg[7]/NET0131  & ~n47572 ;
  assign n59914 = ~n56983 & ~n59577 ;
  assign n59915 = ~n59913 & n59914 ;
  assign n59916 = n25918 & ~n59915 ;
  assign n59917 = ~n59912 & ~n59916 ;
  assign n59918 = \P1_P2_uWord_reg[9]/NET0131  & ~n47529 ;
  assign n59920 = ~\P1_P2_EAX_reg[25]/NET0131  & ~n47555 ;
  assign n59921 = ~n47556 & ~n59920 ;
  assign n59922 = n47570 & n59921 ;
  assign n59919 = \P1_P2_uWord_reg[9]/NET0131  & ~n47572 ;
  assign n59923 = ~n56994 & ~n59919 ;
  assign n59924 = ~n59922 & n59923 ;
  assign n59925 = n25918 & ~n59924 ;
  assign n59926 = ~n59918 & ~n59925 ;
  assign n59928 = \P2_P2_EBX_reg[10]/NET0131  & n46417 ;
  assign n59927 = n46416 & ~n48701 ;
  assign n59929 = ~\P2_P2_EBX_reg[10]/NET0131  & ~n46428 ;
  assign n59930 = ~n46429 & ~n59929 ;
  assign n59931 = n26662 & n59930 ;
  assign n59932 = ~n59927 & ~n59931 ;
  assign n59933 = ~n59928 & n59932 ;
  assign n59934 = n26792 & ~n59933 ;
  assign n59935 = \P2_P2_EBX_reg[10]/NET0131  & ~n44508 ;
  assign n59936 = ~n59934 & ~n59935 ;
  assign n59938 = \P2_P2_EBX_reg[11]/NET0131  & n46417 ;
  assign n59937 = n46416 & ~n48742 ;
  assign n59939 = ~\P2_P2_EBX_reg[11]/NET0131  & ~n46429 ;
  assign n59940 = n26662 & ~n46430 ;
  assign n59941 = ~n59939 & n59940 ;
  assign n59942 = ~n59937 & ~n59941 ;
  assign n59943 = ~n59938 & n59942 ;
  assign n59944 = n26792 & ~n59943 ;
  assign n59945 = \P2_P2_EBX_reg[11]/NET0131  & ~n44508 ;
  assign n59946 = ~n59944 & ~n59945 ;
  assign n59947 = \P2_P2_EBX_reg[12]/NET0131  & ~n44508 ;
  assign n59949 = ~n46417 & ~n59940 ;
  assign n59950 = \P2_P2_EBX_reg[12]/NET0131  & ~n59949 ;
  assign n59948 = n46416 & ~n48787 ;
  assign n59951 = ~\P2_P2_EBX_reg[12]/NET0131  & n46430 ;
  assign n59952 = n26662 & n59951 ;
  assign n59953 = ~n59948 & ~n59952 ;
  assign n59954 = ~n59950 & n59953 ;
  assign n59955 = n26792 & ~n59954 ;
  assign n59956 = ~n59947 & ~n59955 ;
  assign n59959 = ~\P2_P2_EBX_reg[13]/NET0131  & ~n46431 ;
  assign n59960 = n26662 & ~n46432 ;
  assign n59961 = ~n59959 & n59960 ;
  assign n59957 = \P2_P2_EBX_reg[13]/NET0131  & n46417 ;
  assign n59958 = n46416 & ~n48832 ;
  assign n59962 = ~n59957 & ~n59958 ;
  assign n59963 = ~n59961 & n59962 ;
  assign n59964 = n26792 & ~n59963 ;
  assign n59965 = \P2_P2_EBX_reg[13]/NET0131  & ~n44508 ;
  assign n59966 = ~n59964 & ~n59965 ;
  assign n59969 = ~\P2_P2_EBX_reg[14]/NET0131  & ~n46432 ;
  assign n59970 = n26662 & ~n46433 ;
  assign n59971 = ~n59969 & n59970 ;
  assign n59967 = n46416 & ~n48877 ;
  assign n59968 = \P2_P2_EBX_reg[14]/NET0131  & n46417 ;
  assign n59972 = ~n59967 & ~n59968 ;
  assign n59973 = ~n59971 & n59972 ;
  assign n59974 = n26792 & ~n59973 ;
  assign n59975 = \P2_P2_EBX_reg[14]/NET0131  & ~n44508 ;
  assign n59976 = ~n59974 & ~n59975 ;
  assign n59979 = ~\P2_P2_EBX_reg[15]/NET0131  & ~n46433 ;
  assign n59980 = n26662 & ~n46434 ;
  assign n59981 = ~n59979 & n59980 ;
  assign n59977 = n46416 & ~n48178 ;
  assign n59978 = \P2_P2_EBX_reg[15]/NET0131  & n46417 ;
  assign n59982 = ~n59977 & ~n59978 ;
  assign n59983 = ~n59981 & n59982 ;
  assign n59984 = n26792 & ~n59983 ;
  assign n59985 = \P2_P2_EBX_reg[15]/NET0131  & ~n44508 ;
  assign n59986 = ~n59984 & ~n59985 ;
  assign n59989 = ~\P2_P2_EBX_reg[16]/NET0131  & ~n46434 ;
  assign n59990 = n26662 & ~n46435 ;
  assign n59991 = ~n59989 & n59990 ;
  assign n59987 = n46416 & ~n57045 ;
  assign n59988 = \P2_P2_EBX_reg[16]/NET0131  & n46417 ;
  assign n59992 = ~n59987 & ~n59988 ;
  assign n59993 = ~n59991 & n59992 ;
  assign n59994 = n26792 & ~n59993 ;
  assign n59995 = \P2_P2_EBX_reg[16]/NET0131  & ~n44508 ;
  assign n59996 = ~n59994 & ~n59995 ;
  assign n59999 = ~\P2_P2_EBX_reg[17]/NET0131  & ~n46435 ;
  assign n60000 = n26662 & ~n46436 ;
  assign n60001 = ~n59999 & n60000 ;
  assign n59997 = \P2_P2_EBX_reg[17]/NET0131  & n46417 ;
  assign n59998 = n46416 & ~n57099 ;
  assign n60002 = ~n59997 & ~n59998 ;
  assign n60003 = ~n60001 & n60002 ;
  assign n60004 = n26792 & ~n60003 ;
  assign n60005 = \P2_P2_EBX_reg[17]/NET0131  & ~n44508 ;
  assign n60006 = ~n60004 & ~n60005 ;
  assign n60009 = ~\P2_P2_EBX_reg[18]/NET0131  & ~n46436 ;
  assign n60010 = n26662 & ~n46437 ;
  assign n60011 = ~n60009 & n60010 ;
  assign n60007 = \P2_P2_EBX_reg[18]/NET0131  & n46417 ;
  assign n60008 = n46416 & ~n57144 ;
  assign n60012 = ~n60007 & ~n60008 ;
  assign n60013 = ~n60011 & n60012 ;
  assign n60014 = n26792 & ~n60013 ;
  assign n60015 = \P2_P2_EBX_reg[18]/NET0131  & ~n44508 ;
  assign n60016 = ~n60014 & ~n60015 ;
  assign n60019 = ~\P2_P2_EBX_reg[19]/NET0131  & ~n46437 ;
  assign n60020 = n26662 & ~n46438 ;
  assign n60021 = ~n60019 & n60020 ;
  assign n60017 = \P2_P2_EBX_reg[19]/NET0131  & n46417 ;
  assign n60018 = n46416 & ~n57198 ;
  assign n60022 = ~n60017 & ~n60018 ;
  assign n60023 = ~n60021 & n60022 ;
  assign n60024 = n26792 & ~n60023 ;
  assign n60025 = \P2_P2_EBX_reg[19]/NET0131  & ~n44508 ;
  assign n60026 = ~n60024 & ~n60025 ;
  assign n60029 = ~\P2_P2_EBX_reg[20]/NET0131  & ~n46438 ;
  assign n60030 = n26662 & ~n46439 ;
  assign n60031 = ~n60029 & n60030 ;
  assign n60027 = n46416 & ~n57243 ;
  assign n60028 = \P2_P2_EBX_reg[20]/NET0131  & n46417 ;
  assign n60032 = ~n60027 & ~n60028 ;
  assign n60033 = ~n60031 & n60032 ;
  assign n60034 = n26792 & ~n60033 ;
  assign n60035 = \P2_P2_EBX_reg[20]/NET0131  & ~n44508 ;
  assign n60036 = ~n60034 & ~n60035 ;
  assign n60039 = ~\P2_P2_EBX_reg[21]/NET0131  & ~n46439 ;
  assign n60040 = n26662 & ~n46440 ;
  assign n60041 = ~n60039 & n60040 ;
  assign n60037 = \P2_P2_EBX_reg[21]/NET0131  & n46417 ;
  assign n60038 = n46416 & ~n57290 ;
  assign n60042 = ~n60037 & ~n60038 ;
  assign n60043 = ~n60041 & n60042 ;
  assign n60044 = n26792 & ~n60043 ;
  assign n60045 = \P2_P2_EBX_reg[21]/NET0131  & ~n44508 ;
  assign n60046 = ~n60044 & ~n60045 ;
  assign n60049 = ~\P2_P2_EBX_reg[22]/NET0131  & ~n46440 ;
  assign n60050 = n26662 & ~n46441 ;
  assign n60051 = ~n60049 & n60050 ;
  assign n60047 = \P2_P2_EBX_reg[22]/NET0131  & n46417 ;
  assign n60048 = n46416 & ~n57336 ;
  assign n60052 = ~n60047 & ~n60048 ;
  assign n60053 = ~n60051 & n60052 ;
  assign n60054 = n26792 & ~n60053 ;
  assign n60055 = \P2_P2_EBX_reg[22]/NET0131  & ~n44508 ;
  assign n60056 = ~n60054 & ~n60055 ;
  assign n60059 = ~\P2_P2_EBX_reg[23]/NET0131  & ~n46441 ;
  assign n60060 = n26662 & ~n46442 ;
  assign n60061 = ~n60059 & n60060 ;
  assign n60057 = n26578 & n57345 ;
  assign n60058 = \P2_P2_EBX_reg[23]/NET0131  & n46417 ;
  assign n60062 = ~n60057 & ~n60058 ;
  assign n60063 = ~n60061 & n60062 ;
  assign n60064 = n26792 & ~n60063 ;
  assign n60065 = \P2_P2_EBX_reg[23]/NET0131  & ~n44508 ;
  assign n60066 = ~n60064 & ~n60065 ;
  assign n60067 = \P2_P2_EBX_reg[24]/NET0131  & ~n44508 ;
  assign n60070 = ~\P2_P2_EBX_reg[24]/NET0131  & ~n46442 ;
  assign n60071 = n26662 & ~n46443 ;
  assign n60072 = ~n60070 & n60071 ;
  assign n60068 = \P2_P2_EBX_reg[24]/NET0131  & n46417 ;
  assign n60069 = n46416 & n57366 ;
  assign n60073 = ~n60068 & ~n60069 ;
  assign n60074 = ~n60072 & n60073 ;
  assign n60075 = n26792 & ~n60074 ;
  assign n60076 = ~n60067 & ~n60075 ;
  assign n60079 = ~\P2_P2_EBX_reg[28]/NET0131  & ~n46447 ;
  assign n60080 = n26662 & ~n46458 ;
  assign n60081 = ~n60079 & n60080 ;
  assign n60077 = \P2_P2_EBX_reg[28]/NET0131  & n46417 ;
  assign n60078 = n46416 & n57392 ;
  assign n60082 = ~n60077 & ~n60078 ;
  assign n60083 = ~n60081 & n60082 ;
  assign n60084 = n26792 & ~n60083 ;
  assign n60085 = \P2_P2_EBX_reg[28]/NET0131  & ~n44508 ;
  assign n60086 = ~n60084 & ~n60085 ;
  assign n60088 = \P2_P2_EBX_reg[8]/NET0131  & n46417 ;
  assign n60087 = n46416 & ~n48934 ;
  assign n60089 = ~\P2_P2_EBX_reg[8]/NET0131  & ~n46426 ;
  assign n60090 = ~n46427 & ~n60089 ;
  assign n60091 = n26662 & n60090 ;
  assign n60092 = ~n60087 & ~n60091 ;
  assign n60093 = ~n60088 & n60092 ;
  assign n60094 = n26792 & ~n60093 ;
  assign n60095 = \P2_P2_EBX_reg[8]/NET0131  & ~n44508 ;
  assign n60096 = ~n60094 & ~n60095 ;
  assign n60098 = \P2_P2_EBX_reg[9]/NET0131  & n46417 ;
  assign n60097 = n46416 & ~n48979 ;
  assign n60099 = ~\P2_P2_EBX_reg[9]/NET0131  & ~n46427 ;
  assign n60100 = ~n46428 & ~n60099 ;
  assign n60101 = n26662 & n60100 ;
  assign n60102 = ~n60097 & ~n60101 ;
  assign n60103 = ~n60098 & n60102 ;
  assign n60104 = n26792 & ~n60103 ;
  assign n60105 = \P2_P2_EBX_reg[9]/NET0131  & ~n44508 ;
  assign n60106 = ~n60104 & ~n60105 ;
  assign n60107 = ~n26751 & n26792 ;
  assign n60108 = \P2_P2_Flush_reg/NET0131  & ~n44508 ;
  assign n60109 = ~n60107 & ~n60108 ;
  assign n60111 = \P1_P3_EBX_reg[10]/NET0131  & n46480 ;
  assign n60110 = ~n17156 & n46479 ;
  assign n60112 = ~\P1_P3_EBX_reg[10]/NET0131  & ~n46490 ;
  assign n60113 = ~n46491 & ~n60112 ;
  assign n60114 = n9108 & n60113 ;
  assign n60115 = ~n60110 & ~n60114 ;
  assign n60116 = ~n60111 & n60115 ;
  assign n60117 = n9241 & ~n60116 ;
  assign n60118 = \P1_P3_EBX_reg[10]/NET0131  & ~n16968 ;
  assign n60119 = ~n60117 & ~n60118 ;
  assign n60121 = \P1_P3_EBX_reg[11]/NET0131  & n46480 ;
  assign n60120 = ~n17021 & n46479 ;
  assign n60122 = ~\P1_P3_EBX_reg[11]/NET0131  & ~n46491 ;
  assign n60123 = n9108 & ~n46492 ;
  assign n60124 = ~n60122 & n60123 ;
  assign n60125 = ~n60120 & ~n60124 ;
  assign n60126 = ~n60121 & n60125 ;
  assign n60127 = n9241 & ~n60126 ;
  assign n60128 = \P1_P3_EBX_reg[11]/NET0131  & ~n16968 ;
  assign n60129 = ~n60127 & ~n60128 ;
  assign n60131 = \P1_P1_EBX_reg[10]/NET0131  & ~n46533 ;
  assign n60130 = ~n27364 & n46535 ;
  assign n60132 = ~\P1_P1_EBX_reg[10]/NET0131  & ~n46545 ;
  assign n60133 = ~n46546 & ~n60132 ;
  assign n60134 = n26146 & n60133 ;
  assign n60135 = ~n60130 & ~n60134 ;
  assign n60136 = ~n60131 & n60135 ;
  assign n60137 = n8355 & ~n60136 ;
  assign n60138 = \P1_P1_EBX_reg[10]/NET0131  & ~n15326 ;
  assign n60139 = ~n60137 & ~n60138 ;
  assign n60142 = ~\P1_P3_EBX_reg[12]/NET0131  & ~n46492 ;
  assign n60143 = n9108 & ~n46493 ;
  assign n60144 = ~n60142 & n60143 ;
  assign n60140 = \P1_P3_EBX_reg[12]/NET0131  & n46480 ;
  assign n60141 = ~n17070 & n46479 ;
  assign n60145 = ~n60140 & ~n60141 ;
  assign n60146 = ~n60144 & n60145 ;
  assign n60147 = n9241 & ~n60146 ;
  assign n60148 = \P1_P3_EBX_reg[12]/NET0131  & ~n16968 ;
  assign n60149 = ~n60147 & ~n60148 ;
  assign n60152 = ~\P1_P3_EBX_reg[13]/NET0131  & ~n46493 ;
  assign n60153 = n9108 & ~n46494 ;
  assign n60154 = ~n60152 & n60153 ;
  assign n60150 = ~n17113 & n46479 ;
  assign n60151 = \P1_P3_EBX_reg[13]/NET0131  & n46480 ;
  assign n60155 = ~n60150 & ~n60151 ;
  assign n60156 = ~n60154 & n60155 ;
  assign n60157 = n9241 & ~n60156 ;
  assign n60158 = \P1_P3_EBX_reg[13]/NET0131  & ~n16968 ;
  assign n60159 = ~n60157 & ~n60158 ;
  assign n60162 = ~\P1_P3_EBX_reg[14]/NET0131  & ~n46494 ;
  assign n60163 = n9108 & ~n46495 ;
  assign n60164 = ~n60162 & n60163 ;
  assign n60160 = ~n17201 & n46479 ;
  assign n60161 = \P1_P3_EBX_reg[14]/NET0131  & n46480 ;
  assign n60165 = ~n60160 & ~n60161 ;
  assign n60166 = ~n60164 & n60165 ;
  assign n60167 = n9241 & ~n60166 ;
  assign n60168 = \P1_P3_EBX_reg[14]/NET0131  & ~n16968 ;
  assign n60169 = ~n60167 & ~n60168 ;
  assign n60172 = ~\P1_P3_EBX_reg[15]/NET0131  & ~n46495 ;
  assign n60173 = n9108 & ~n46496 ;
  assign n60174 = ~n60172 & n60173 ;
  assign n60170 = ~n17242 & n46479 ;
  assign n60171 = \P1_P3_EBX_reg[15]/NET0131  & n46480 ;
  assign n60175 = ~n60170 & ~n60171 ;
  assign n60176 = ~n60174 & n60175 ;
  assign n60177 = n9241 & ~n60176 ;
  assign n60178 = \P1_P3_EBX_reg[15]/NET0131  & ~n16968 ;
  assign n60179 = ~n60177 & ~n60178 ;
  assign n60182 = ~\P1_P3_EBX_reg[16]/NET0131  & ~n46496 ;
  assign n60183 = n9108 & ~n46497 ;
  assign n60184 = ~n60182 & n60183 ;
  assign n60180 = ~n18789 & n46479 ;
  assign n60181 = \P1_P3_EBX_reg[16]/NET0131  & n46480 ;
  assign n60185 = ~n60180 & ~n60181 ;
  assign n60186 = ~n60184 & n60185 ;
  assign n60187 = n9241 & ~n60186 ;
  assign n60188 = \P1_P3_EBX_reg[16]/NET0131  & ~n16968 ;
  assign n60189 = ~n60187 & ~n60188 ;
  assign n60192 = ~\P1_P3_EBX_reg[17]/NET0131  & ~n46497 ;
  assign n60193 = n9108 & ~n46498 ;
  assign n60194 = ~n60192 & n60193 ;
  assign n60190 = \P1_P3_EBX_reg[17]/NET0131  & n46480 ;
  assign n60191 = ~n21146 & n46479 ;
  assign n60195 = ~n60190 & ~n60191 ;
  assign n60196 = ~n60194 & n60195 ;
  assign n60197 = n9241 & ~n60196 ;
  assign n60198 = \P1_P3_EBX_reg[17]/NET0131  & ~n16968 ;
  assign n60199 = ~n60197 & ~n60198 ;
  assign n60201 = \P1_P1_EBX_reg[11]/NET0131  & ~n46533 ;
  assign n60200 = ~n25323 & n46535 ;
  assign n60202 = ~\P1_P1_EBX_reg[11]/NET0131  & ~n46546 ;
  assign n60203 = n26146 & ~n46547 ;
  assign n60204 = ~n60202 & n60203 ;
  assign n60205 = ~n60200 & ~n60204 ;
  assign n60206 = ~n60201 & n60205 ;
  assign n60207 = n8355 & ~n60206 ;
  assign n60208 = \P1_P1_EBX_reg[11]/NET0131  & ~n15326 ;
  assign n60209 = ~n60207 & ~n60208 ;
  assign n60212 = ~\P1_P3_EBX_reg[18]/NET0131  & ~n46498 ;
  assign n60213 = n9108 & ~n46499 ;
  assign n60214 = ~n60212 & n60213 ;
  assign n60210 = \P1_P3_EBX_reg[18]/NET0131  & n46480 ;
  assign n60211 = ~n18849 & n46479 ;
  assign n60215 = ~n60210 & ~n60211 ;
  assign n60216 = ~n60214 & n60215 ;
  assign n60217 = n9241 & ~n60216 ;
  assign n60218 = \P1_P3_EBX_reg[18]/NET0131  & ~n16968 ;
  assign n60219 = ~n60217 & ~n60218 ;
  assign n60222 = ~\P1_P3_EBX_reg[19]/NET0131  & ~n46499 ;
  assign n60223 = n9108 & ~n46500 ;
  assign n60224 = ~n60222 & n60223 ;
  assign n60220 = \P1_P3_EBX_reg[19]/NET0131  & n46480 ;
  assign n60221 = ~n21200 & n46479 ;
  assign n60225 = ~n60220 & ~n60221 ;
  assign n60226 = ~n60224 & n60225 ;
  assign n60227 = n9241 & ~n60226 ;
  assign n60228 = \P1_P3_EBX_reg[19]/NET0131  & ~n16968 ;
  assign n60229 = ~n60227 & ~n60228 ;
  assign n60232 = ~\P1_P3_EBX_reg[20]/NET0131  & ~n46500 ;
  assign n60233 = n9108 & ~n46501 ;
  assign n60234 = ~n60232 & n60233 ;
  assign n60230 = ~n21243 & n46479 ;
  assign n60231 = \P1_P3_EBX_reg[20]/NET0131  & n46480 ;
  assign n60235 = ~n60230 & ~n60231 ;
  assign n60236 = ~n60234 & n60235 ;
  assign n60237 = n9241 & ~n60236 ;
  assign n60238 = \P1_P3_EBX_reg[20]/NET0131  & ~n16968 ;
  assign n60239 = ~n60237 & ~n60238 ;
  assign n60241 = \P1_P1_EBX_reg[12]/NET0131  & ~n46533 ;
  assign n60240 = ~n24958 & n46535 ;
  assign n60242 = ~\P1_P1_EBX_reg[12]/NET0131  & ~n46547 ;
  assign n60243 = n26146 & ~n46548 ;
  assign n60244 = ~n60242 & n60243 ;
  assign n60245 = ~n60240 & ~n60244 ;
  assign n60246 = ~n60241 & n60245 ;
  assign n60247 = n8355 & ~n60246 ;
  assign n60248 = \P1_P1_EBX_reg[12]/NET0131  & ~n15326 ;
  assign n60249 = ~n60247 & ~n60248 ;
  assign n60252 = ~\P1_P3_EBX_reg[21]/NET0131  & ~n46501 ;
  assign n60253 = n9108 & ~n46502 ;
  assign n60254 = ~n60252 & n60253 ;
  assign n60250 = \P1_P3_EBX_reg[21]/NET0131  & n46480 ;
  assign n60251 = ~n21295 & n46479 ;
  assign n60255 = ~n60250 & ~n60251 ;
  assign n60256 = ~n60254 & n60255 ;
  assign n60257 = n9241 & ~n60256 ;
  assign n60258 = \P1_P3_EBX_reg[21]/NET0131  & ~n16968 ;
  assign n60259 = ~n60257 & ~n60258 ;
  assign n60262 = ~\P1_P3_EBX_reg[22]/NET0131  & ~n46502 ;
  assign n60263 = n9108 & ~n46503 ;
  assign n60264 = ~n60262 & n60263 ;
  assign n60260 = \P1_P3_EBX_reg[22]/NET0131  & n46480 ;
  assign n60261 = ~n21343 & n46479 ;
  assign n60265 = ~n60260 & ~n60261 ;
  assign n60266 = ~n60264 & n60265 ;
  assign n60267 = n9241 & ~n60266 ;
  assign n60268 = \P1_P3_EBX_reg[22]/NET0131  & ~n16968 ;
  assign n60269 = ~n60267 & ~n60268 ;
  assign n60272 = ~\P1_P3_EBX_reg[23]/NET0131  & ~n46503 ;
  assign n60273 = n9108 & ~n46504 ;
  assign n60274 = ~n60272 & n60273 ;
  assign n60270 = \P1_P3_EBX_reg[23]/NET0131  & n46480 ;
  assign n60271 = n21415 & n46479 ;
  assign n60275 = ~n60270 & ~n60271 ;
  assign n60276 = ~n60274 & n60275 ;
  assign n60277 = n9241 & ~n60276 ;
  assign n60278 = \P1_P3_EBX_reg[23]/NET0131  & ~n16968 ;
  assign n60279 = ~n60277 & ~n60278 ;
  assign n60280 = \P1_P3_EBX_reg[24]/NET0131  & ~n16968 ;
  assign n60283 = ~\P1_P3_EBX_reg[24]/NET0131  & ~n46504 ;
  assign n60284 = n9108 & ~n46505 ;
  assign n60285 = ~n60283 & n60284 ;
  assign n60281 = \P1_P3_EBX_reg[24]/NET0131  & n46480 ;
  assign n60282 = n21467 & n46479 ;
  assign n60286 = ~n60281 & ~n60282 ;
  assign n60287 = ~n60285 & n60286 ;
  assign n60288 = n9241 & ~n60287 ;
  assign n60289 = ~n60280 & ~n60288 ;
  assign n60292 = ~\P1_P1_EBX_reg[13]/NET0131  & ~n46548 ;
  assign n60293 = n26146 & ~n46549 ;
  assign n60294 = ~n60292 & n60293 ;
  assign n60290 = \P1_P1_EBX_reg[13]/NET0131  & ~n46533 ;
  assign n60291 = ~n24551 & n46535 ;
  assign n60295 = ~n60290 & ~n60291 ;
  assign n60296 = ~n60294 & n60295 ;
  assign n60297 = n8355 & ~n60296 ;
  assign n60298 = \P1_P1_EBX_reg[13]/NET0131  & ~n15326 ;
  assign n60299 = ~n60297 & ~n60298 ;
  assign n60302 = ~\P1_P3_EBX_reg[28]/NET0131  & ~n46509 ;
  assign n60303 = n9108 & ~n46520 ;
  assign n60304 = ~n60302 & n60303 ;
  assign n60300 = \P1_P3_EBX_reg[28]/NET0131  & n46480 ;
  assign n60301 = n21940 & n46479 ;
  assign n60305 = ~n60300 & ~n60301 ;
  assign n60306 = ~n60304 & n60305 ;
  assign n60307 = n9241 & ~n60306 ;
  assign n60308 = \P1_P3_EBX_reg[28]/NET0131  & ~n16968 ;
  assign n60309 = ~n60307 & ~n60308 ;
  assign n60312 = ~\P1_P1_EBX_reg[14]/NET0131  & ~n46549 ;
  assign n60313 = n26146 & ~n46550 ;
  assign n60314 = ~n60312 & n60313 ;
  assign n60310 = ~n24339 & n46535 ;
  assign n60311 = \P1_P1_EBX_reg[14]/NET0131  & ~n46533 ;
  assign n60315 = ~n60310 & ~n60311 ;
  assign n60316 = ~n60314 & n60315 ;
  assign n60317 = n8355 & ~n60316 ;
  assign n60318 = \P1_P1_EBX_reg[14]/NET0131  & ~n15326 ;
  assign n60319 = ~n60317 & ~n60318 ;
  assign n60322 = ~\P1_P1_EBX_reg[15]/NET0131  & ~n46550 ;
  assign n60323 = n26146 & ~n46551 ;
  assign n60324 = ~n60322 & n60323 ;
  assign n60320 = ~n24392 & n46535 ;
  assign n60321 = \P1_P1_EBX_reg[15]/NET0131  & ~n46533 ;
  assign n60325 = ~n60320 & ~n60321 ;
  assign n60326 = ~n60324 & n60325 ;
  assign n60327 = n8355 & ~n60326 ;
  assign n60328 = \P1_P1_EBX_reg[15]/NET0131  & ~n15326 ;
  assign n60329 = ~n60327 & ~n60328 ;
  assign n60332 = ~\P1_P1_EBX_reg[16]/NET0131  & ~n46551 ;
  assign n60333 = n26146 & ~n46552 ;
  assign n60334 = ~n60332 & n60333 ;
  assign n60330 = ~n25005 & n46535 ;
  assign n60331 = \P1_P1_EBX_reg[16]/NET0131  & ~n46533 ;
  assign n60335 = ~n60330 & ~n60331 ;
  assign n60336 = ~n60334 & n60335 ;
  assign n60337 = n8355 & ~n60336 ;
  assign n60338 = \P1_P1_EBX_reg[16]/NET0131  & ~n15326 ;
  assign n60339 = ~n60337 & ~n60338 ;
  assign n60341 = \P1_P3_EBX_reg[8]/NET0131  & n46480 ;
  assign n60340 = ~n17326 & n46479 ;
  assign n60342 = ~\P1_P3_EBX_reg[8]/NET0131  & ~n46488 ;
  assign n60343 = ~n46489 & ~n60342 ;
  assign n60344 = n9108 & n60343 ;
  assign n60345 = ~n60340 & ~n60344 ;
  assign n60346 = ~n60341 & n60345 ;
  assign n60347 = n9241 & ~n60346 ;
  assign n60348 = \P1_P3_EBX_reg[8]/NET0131  & ~n16968 ;
  assign n60349 = ~n60347 & ~n60348 ;
  assign n60351 = \P1_P3_EBX_reg[9]/NET0131  & n46480 ;
  assign n60350 = ~n17368 & n46479 ;
  assign n60352 = ~\P1_P3_EBX_reg[9]/NET0131  & ~n46489 ;
  assign n60353 = ~n46490 & ~n60352 ;
  assign n60354 = n9108 & n60353 ;
  assign n60355 = ~n60350 & ~n60354 ;
  assign n60356 = ~n60351 & n60355 ;
  assign n60357 = n9241 & ~n60356 ;
  assign n60358 = \P1_P3_EBX_reg[9]/NET0131  & ~n16968 ;
  assign n60359 = ~n60357 & ~n60358 ;
  assign n60362 = ~\P1_P1_EBX_reg[17]/NET0131  & ~n46552 ;
  assign n60363 = n26146 & ~n46553 ;
  assign n60364 = ~n60362 & n60363 ;
  assign n60360 = \P1_P1_EBX_reg[17]/NET0131  & ~n46533 ;
  assign n60361 = ~n25048 & n46535 ;
  assign n60365 = ~n60360 & ~n60361 ;
  assign n60366 = ~n60364 & n60365 ;
  assign n60367 = n8355 & ~n60366 ;
  assign n60368 = \P1_P1_EBX_reg[17]/NET0131  & ~n15326 ;
  assign n60369 = ~n60367 & ~n60368 ;
  assign n60372 = ~\P1_P1_EBX_reg[18]/NET0131  & ~n46553 ;
  assign n60373 = n26146 & ~n46554 ;
  assign n60374 = ~n60372 & n60373 ;
  assign n60370 = ~n24599 & n46535 ;
  assign n60371 = \P1_P1_EBX_reg[18]/NET0131  & ~n46533 ;
  assign n60375 = ~n60370 & ~n60371 ;
  assign n60376 = ~n60374 & n60375 ;
  assign n60377 = n8355 & ~n60376 ;
  assign n60378 = \P1_P1_EBX_reg[18]/NET0131  & ~n15326 ;
  assign n60379 = ~n60377 & ~n60378 ;
  assign n60382 = ~\P1_P1_EBX_reg[19]/NET0131  & ~n46554 ;
  assign n60383 = n26146 & ~n46555 ;
  assign n60384 = ~n60382 & n60383 ;
  assign n60380 = \P1_P1_EBX_reg[19]/NET0131  & ~n46533 ;
  assign n60381 = ~n24638 & n46535 ;
  assign n60385 = ~n60380 & ~n60381 ;
  assign n60386 = ~n60384 & n60385 ;
  assign n60387 = n8355 & ~n60386 ;
  assign n60388 = \P1_P1_EBX_reg[19]/NET0131  & ~n15326 ;
  assign n60389 = ~n60387 & ~n60388 ;
  assign n60392 = ~\P1_P1_EBX_reg[20]/NET0131  & ~n46555 ;
  assign n60393 = n26146 & ~n46556 ;
  assign n60394 = ~n60392 & n60393 ;
  assign n60390 = ~n24689 & n46535 ;
  assign n60391 = \P1_P1_EBX_reg[20]/NET0131  & ~n46533 ;
  assign n60395 = ~n60390 & ~n60391 ;
  assign n60396 = ~n60394 & n60395 ;
  assign n60397 = n8355 & ~n60396 ;
  assign n60398 = \P1_P1_EBX_reg[20]/NET0131  & ~n15326 ;
  assign n60399 = ~n60397 & ~n60398 ;
  assign n60402 = ~\P1_P1_EBX_reg[21]/NET0131  & ~n46556 ;
  assign n60403 = n26146 & ~n46557 ;
  assign n60404 = ~n60402 & n60403 ;
  assign n60400 = ~n24430 & n46535 ;
  assign n60401 = \P1_P1_EBX_reg[21]/NET0131  & ~n46533 ;
  assign n60405 = ~n60400 & ~n60401 ;
  assign n60406 = ~n60404 & n60405 ;
  assign n60407 = n8355 & ~n60406 ;
  assign n60408 = \P1_P1_EBX_reg[21]/NET0131  & ~n15326 ;
  assign n60409 = ~n60407 & ~n60408 ;
  assign n60412 = ~\P1_P1_EBX_reg[22]/NET0131  & ~n46557 ;
  assign n60413 = n26146 & ~n46558 ;
  assign n60414 = ~n60412 & n60413 ;
  assign n60410 = \P1_P1_EBX_reg[22]/NET0131  & ~n46533 ;
  assign n60411 = ~n24200 & n46535 ;
  assign n60415 = ~n60410 & ~n60411 ;
  assign n60416 = ~n60414 & n60415 ;
  assign n60417 = n8355 & ~n60416 ;
  assign n60418 = \P1_P1_EBX_reg[22]/NET0131  & ~n15326 ;
  assign n60419 = ~n60417 & ~n60418 ;
  assign n60422 = ~\P1_P1_EBX_reg[23]/NET0131  & ~n46558 ;
  assign n60423 = n26146 & ~n46559 ;
  assign n60424 = ~n60422 & n60423 ;
  assign n60420 = n24138 & n26122 ;
  assign n60421 = \P1_P1_EBX_reg[23]/NET0131  & ~n46533 ;
  assign n60425 = ~n60420 & ~n60421 ;
  assign n60426 = ~n60424 & n60425 ;
  assign n60427 = n8355 & ~n60426 ;
  assign n60428 = \P1_P1_EBX_reg[23]/NET0131  & ~n15326 ;
  assign n60429 = ~n60427 & ~n60428 ;
  assign n60430 = n15334 & n25363 ;
  assign n60431 = ~n24505 & ~n60430 ;
  assign n60432 = n8355 & ~n60431 ;
  assign n60433 = n24515 & ~n60432 ;
  assign n60434 = \P1_P1_uWord_reg[0]/NET0131  & ~n60433 ;
  assign n60435 = ~n7924 & n23946 ;
  assign n60436 = ~\P1_P1_EAX_reg[16]/NET0131  & ~n25347 ;
  assign n60437 = ~n25348 & ~n60436 ;
  assign n60438 = n24502 & n60437 ;
  assign n60439 = ~n60435 & ~n60438 ;
  assign n60440 = n8355 & ~n15364 ;
  assign n60441 = ~n60439 & n60440 ;
  assign n60442 = ~n60434 & ~n60441 ;
  assign n60447 = ~\P1_P1_EBX_reg[24]/NET0131  & ~n46559 ;
  assign n60448 = n26146 & ~n46560 ;
  assign n60449 = ~n60447 & n60448 ;
  assign n60443 = \P1_P1_EBX_reg[24]/NET0131  & n46531 ;
  assign n60444 = \P1_P1_EBX_reg[24]/NET0131  & ~n15428 ;
  assign n60445 = ~n23920 & ~n60444 ;
  assign n60446 = n26122 & ~n60445 ;
  assign n60450 = ~n60443 & ~n60446 ;
  assign n60451 = ~n60449 & n60450 ;
  assign n60452 = n8355 & ~n60451 ;
  assign n60453 = \P1_P1_EBX_reg[24]/NET0131  & ~n15326 ;
  assign n60454 = ~n60452 & ~n60453 ;
  assign n60455 = \P1_P1_uWord_reg[1]/NET0131  & ~n24515 ;
  assign n60459 = \P1_P1_uWord_reg[1]/NET0131  & ~n60431 ;
  assign n60456 = ~\P1_P1_EAX_reg[17]/NET0131  & ~n25348 ;
  assign n60457 = ~n25349 & ~n60456 ;
  assign n60458 = n24503 & n60457 ;
  assign n60460 = ~n25051 & ~n60458 ;
  assign n60461 = ~n60459 & n60460 ;
  assign n60462 = n8355 & ~n60461 ;
  assign n60463 = ~n60455 & ~n60462 ;
  assign n60464 = \P1_P1_uWord_reg[2]/NET0131  & ~n60433 ;
  assign n60465 = ~\P1_P1_EAX_reg[18]/NET0131  & ~n25349 ;
  assign n60466 = ~n25350 & ~n60465 ;
  assign n60467 = n24503 & n60466 ;
  assign n60468 = ~n24601 & ~n60467 ;
  assign n60469 = n8355 & ~n60468 ;
  assign n60470 = ~n60464 & ~n60469 ;
  assign n60473 = ~\P1_P1_EBX_reg[28]/NET0131  & ~n46564 ;
  assign n60474 = n26146 & ~n46575 ;
  assign n60475 = ~n60473 & n60474 ;
  assign n60471 = \P1_P1_EBX_reg[28]/NET0131  & ~n46533 ;
  assign n60472 = n22817 & n46535 ;
  assign n60476 = ~n60471 & ~n60472 ;
  assign n60477 = ~n60475 & n60476 ;
  assign n60478 = n8355 & ~n60477 ;
  assign n60479 = \P1_P1_EBX_reg[28]/NET0131  & ~n15326 ;
  assign n60480 = ~n60478 & ~n60479 ;
  assign n60482 = \P1_P1_EBX_reg[8]/NET0131  & ~n46533 ;
  assign n60481 = ~n27778 & n46535 ;
  assign n60483 = ~\P1_P1_EBX_reg[8]/NET0131  & ~n46543 ;
  assign n60484 = ~n46544 & ~n60483 ;
  assign n60485 = n26146 & n60484 ;
  assign n60486 = ~n60481 & ~n60485 ;
  assign n60487 = ~n60482 & n60486 ;
  assign n60488 = n8355 & ~n60487 ;
  assign n60489 = \P1_P1_EBX_reg[8]/NET0131  & ~n15326 ;
  assign n60490 = ~n60488 & ~n60489 ;
  assign n60491 = \P2_P2_uWord_reg[0]/NET0131  & ~n47642 ;
  assign n60498 = \P2_P2_uWord_reg[0]/NET0131  & n47685 ;
  assign n60492 = ~\P2_P2_EAX_reg[16]/NET0131  & ~n47659 ;
  assign n60493 = ~n47660 & ~n60492 ;
  assign n60494 = n26786 & n60493 ;
  assign n60495 = \P2_P2_uWord_reg[0]/NET0131  & n26286 ;
  assign n60496 = ~n57050 & ~n60495 ;
  assign n60497 = n26633 & ~n60496 ;
  assign n60499 = ~n60494 & ~n60497 ;
  assign n60500 = ~n60498 & n60499 ;
  assign n60501 = n26792 & ~n60500 ;
  assign n60502 = ~n60491 & ~n60501 ;
  assign n60503 = \P2_P2_uWord_reg[10]/NET0131  & ~n47642 ;
  assign n60504 = ~\P2_P2_EAX_reg[26]/NET0131  & ~n47669 ;
  assign n60505 = ~n47670 & ~n60504 ;
  assign n60506 = n26643 & n60505 ;
  assign n60507 = ~n57445 & ~n60506 ;
  assign n60508 = ~n26640 & ~n60507 ;
  assign n60509 = \P2_P2_uWord_reg[10]/NET0131  & ~n47686 ;
  assign n60510 = ~n60508 & ~n60509 ;
  assign n60511 = n26792 & ~n60510 ;
  assign n60512 = ~n60503 & ~n60511 ;
  assign n60514 = \P1_P1_EBX_reg[9]/NET0131  & ~n46533 ;
  assign n60513 = ~n27584 & n46535 ;
  assign n60515 = ~\P1_P1_EBX_reg[9]/NET0131  & ~n46544 ;
  assign n60516 = ~n46545 & ~n60515 ;
  assign n60517 = n26146 & n60516 ;
  assign n60518 = ~n60513 & ~n60517 ;
  assign n60519 = ~n60514 & n60518 ;
  assign n60520 = n8355 & ~n60519 ;
  assign n60521 = \P1_P1_EBX_reg[9]/NET0131  & ~n15326 ;
  assign n60522 = ~n60520 & ~n60521 ;
  assign n60523 = \P2_P2_uWord_reg[13]/NET0131  & ~n57437 ;
  assign n60525 = ~\P2_P2_EAX_reg[29]/NET0131  & ~n47673 ;
  assign n60524 = \P2_P2_EAX_reg[29]/NET0131  & n47673 ;
  assign n60526 = n26643 & ~n60524 ;
  assign n60527 = ~n60525 & n60526 ;
  assign n60528 = ~n57469 & ~n60527 ;
  assign n60529 = n57448 & ~n60528 ;
  assign n60530 = ~n60523 & ~n60529 ;
  assign n60531 = \P2_P2_uWord_reg[14]/NET0131  & ~n57437 ;
  assign n60533 = \P2_P2_EAX_reg[30]/NET0131  & n60524 ;
  assign n60532 = ~\P2_P2_EAX_reg[30]/NET0131  & ~n60524 ;
  assign n60534 = n26643 & ~n60532 ;
  assign n60535 = ~n60533 & n60534 ;
  assign n60536 = ~n57475 & ~n60535 ;
  assign n60537 = n57448 & ~n60536 ;
  assign n60538 = ~n60531 & ~n60537 ;
  assign n60539 = \P2_P2_uWord_reg[1]/NET0131  & ~n47642 ;
  assign n60546 = \P2_P2_uWord_reg[1]/NET0131  & n47685 ;
  assign n60540 = ~\P2_P2_EAX_reg[17]/NET0131  & ~n47660 ;
  assign n60541 = ~n47661 & ~n60540 ;
  assign n60542 = n26786 & n60541 ;
  assign n60543 = \P2_P2_uWord_reg[1]/NET0131  & n26286 ;
  assign n60544 = ~n53130 & ~n60543 ;
  assign n60545 = n26633 & ~n60544 ;
  assign n60547 = ~n60542 & ~n60545 ;
  assign n60548 = ~n60546 & n60547 ;
  assign n60549 = n26792 & ~n60548 ;
  assign n60550 = ~n60539 & ~n60549 ;
  assign n60551 = ~\P2_P2_EAX_reg[18]/NET0131  & ~n47661 ;
  assign n60552 = ~n47662 & ~n60551 ;
  assign n60553 = n26643 & n60552 ;
  assign n60554 = ~n57507 & ~n60553 ;
  assign n60555 = ~n26640 & ~n60554 ;
  assign n60556 = \P2_P2_uWord_reg[2]/NET0131  & ~n47686 ;
  assign n60557 = ~n60555 & ~n60556 ;
  assign n60558 = n26792 & ~n60557 ;
  assign n60559 = \P2_P2_uWord_reg[2]/NET0131  & ~n47642 ;
  assign n60560 = ~n60558 & ~n60559 ;
  assign n60561 = ~n57516 & ~n59527 ;
  assign n60562 = ~n26640 & ~n60561 ;
  assign n60563 = \P2_P2_uWord_reg[3]/NET0131  & ~n47686 ;
  assign n60564 = ~n60562 & ~n60563 ;
  assign n60565 = n26792 & ~n60564 ;
  assign n60566 = \P2_P2_uWord_reg[3]/NET0131  & ~n47642 ;
  assign n60567 = ~n60565 & ~n60566 ;
  assign n60568 = \P2_P2_uWord_reg[5]/NET0131  & ~n47642 ;
  assign n60575 = \P2_P2_uWord_reg[5]/NET0131  & n47685 ;
  assign n60569 = ~\P2_P2_EAX_reg[21]/NET0131  & ~n47664 ;
  assign n60570 = ~n47665 & ~n60569 ;
  assign n60571 = n26786 & n60570 ;
  assign n60572 = \P2_P2_uWord_reg[5]/NET0131  & n26286 ;
  assign n60573 = ~n53198 & ~n60572 ;
  assign n60574 = n26633 & ~n60573 ;
  assign n60576 = ~n60571 & ~n60574 ;
  assign n60577 = ~n60575 & n60576 ;
  assign n60578 = n26792 & ~n60577 ;
  assign n60579 = ~n60568 & ~n60578 ;
  assign n60580 = n8355 & ~n26270 ;
  assign n60581 = \P1_P1_Flush_reg/NET0131  & ~n15326 ;
  assign n60582 = ~n60580 & ~n60581 ;
  assign n60583 = \P2_P2_uWord_reg[6]/NET0131  & ~n47642 ;
  assign n60590 = \P2_P2_uWord_reg[6]/NET0131  & n47685 ;
  assign n60584 = ~\P2_P2_EAX_reg[22]/NET0131  & ~n47665 ;
  assign n60585 = n26786 & ~n47666 ;
  assign n60586 = ~n60584 & n60585 ;
  assign n60587 = \P2_P2_uWord_reg[6]/NET0131  & n26286 ;
  assign n60588 = ~n53212 & ~n60587 ;
  assign n60589 = n26633 & ~n60588 ;
  assign n60591 = ~n60586 & ~n60589 ;
  assign n60592 = ~n60590 & n60591 ;
  assign n60593 = n26792 & ~n60592 ;
  assign n60594 = ~n60583 & ~n60593 ;
  assign n60595 = \P2_P2_uWord_reg[7]/NET0131  & ~n57437 ;
  assign n60596 = ~n57552 & ~n59536 ;
  assign n60597 = n57448 & ~n60596 ;
  assign n60598 = ~n60595 & ~n60597 ;
  assign n60599 = \P2_P2_uWord_reg[9]/NET0131  & ~n57437 ;
  assign n60600 = ~\P2_P2_EAX_reg[25]/NET0131  & ~n47668 ;
  assign n60601 = ~n47669 & ~n60600 ;
  assign n60602 = n26643 & n60601 ;
  assign n60603 = ~n57567 & ~n60602 ;
  assign n60604 = n57448 & ~n60603 ;
  assign n60605 = ~n60599 & ~n60604 ;
  assign n60607 = \P2_P3_EBX_reg[10]/NET0131  & n46615 ;
  assign n60606 = n46614 & ~n49074 ;
  assign n60608 = ~\P2_P3_EBX_reg[10]/NET0131  & ~n46626 ;
  assign n60609 = ~n46627 & ~n60608 ;
  assign n60610 = n27133 & n60609 ;
  assign n60611 = ~n60606 & ~n60610 ;
  assign n60612 = ~n60607 & n60611 ;
  assign n60613 = n27308 & ~n60612 ;
  assign n60614 = \P2_P3_EBX_reg[10]/NET0131  & ~n42872 ;
  assign n60615 = ~n60613 & ~n60614 ;
  assign n60617 = \P2_P3_EBX_reg[11]/NET0131  & n46615 ;
  assign n60616 = n46614 & ~n49116 ;
  assign n60618 = ~\P2_P3_EBX_reg[11]/NET0131  & ~n46627 ;
  assign n60619 = n27133 & ~n46628 ;
  assign n60620 = ~n60618 & n60619 ;
  assign n60621 = ~n60616 & ~n60620 ;
  assign n60622 = ~n60617 & n60621 ;
  assign n60623 = n27308 & ~n60622 ;
  assign n60624 = \P2_P3_EBX_reg[11]/NET0131  & ~n42872 ;
  assign n60625 = ~n60623 & ~n60624 ;
  assign n60626 = \P2_P3_EBX_reg[12]/NET0131  & ~n42872 ;
  assign n60628 = ~n46615 & ~n60619 ;
  assign n60629 = \P2_P3_EBX_reg[12]/NET0131  & ~n60628 ;
  assign n60627 = n46614 & ~n49162 ;
  assign n60630 = ~\P2_P3_EBX_reg[12]/NET0131  & n46628 ;
  assign n60631 = n27133 & n60630 ;
  assign n60632 = ~n60627 & ~n60631 ;
  assign n60633 = ~n60629 & n60632 ;
  assign n60634 = n27308 & ~n60633 ;
  assign n60635 = ~n60626 & ~n60634 ;
  assign n60638 = ~\P2_P3_EBX_reg[13]/NET0131  & ~n46629 ;
  assign n60639 = n27133 & ~n46630 ;
  assign n60640 = ~n60638 & n60639 ;
  assign n60636 = \P2_P3_EBX_reg[13]/NET0131  & n46615 ;
  assign n60637 = n46614 & ~n49204 ;
  assign n60641 = ~n60636 & ~n60637 ;
  assign n60642 = ~n60640 & n60641 ;
  assign n60643 = n27308 & ~n60642 ;
  assign n60644 = \P2_P3_EBX_reg[13]/NET0131  & ~n42872 ;
  assign n60645 = ~n60643 & ~n60644 ;
  assign n60648 = ~\P2_P3_EBX_reg[14]/NET0131  & ~n46630 ;
  assign n60649 = n27133 & ~n46631 ;
  assign n60650 = ~n60648 & n60649 ;
  assign n60646 = n46614 & ~n49250 ;
  assign n60647 = \P2_P3_EBX_reg[14]/NET0131  & n46615 ;
  assign n60651 = ~n60646 & ~n60647 ;
  assign n60652 = ~n60650 & n60651 ;
  assign n60653 = n27308 & ~n60652 ;
  assign n60654 = \P2_P3_EBX_reg[14]/NET0131  & ~n42872 ;
  assign n60655 = ~n60653 & ~n60654 ;
  assign n60658 = ~\P2_P3_EBX_reg[15]/NET0131  & ~n46631 ;
  assign n60659 = n27133 & ~n46632 ;
  assign n60660 = ~n60658 & n60659 ;
  assign n60656 = \P2_P3_EBX_reg[15]/NET0131  & n46615 ;
  assign n60657 = n46614 & ~n49295 ;
  assign n60661 = ~n60656 & ~n60657 ;
  assign n60662 = ~n60660 & n60661 ;
  assign n60663 = n27308 & ~n60662 ;
  assign n60664 = \P2_P3_EBX_reg[15]/NET0131  & ~n42872 ;
  assign n60665 = ~n60663 & ~n60664 ;
  assign n60668 = ~\P2_P3_EBX_reg[16]/NET0131  & ~n46632 ;
  assign n60669 = n27133 & ~n46633 ;
  assign n60670 = ~n60668 & n60669 ;
  assign n60666 = n46614 & ~n57607 ;
  assign n60667 = \P2_P3_EBX_reg[16]/NET0131  & n46615 ;
  assign n60671 = ~n60666 & ~n60667 ;
  assign n60672 = ~n60670 & n60671 ;
  assign n60673 = n27308 & ~n60672 ;
  assign n60674 = \P2_P3_EBX_reg[16]/NET0131  & ~n42872 ;
  assign n60675 = ~n60673 & ~n60674 ;
  assign n60678 = ~\P2_P3_EBX_reg[17]/NET0131  & ~n46633 ;
  assign n60679 = n27133 & ~n46634 ;
  assign n60680 = ~n60678 & n60679 ;
  assign n60676 = \P2_P3_EBX_reg[17]/NET0131  & n46615 ;
  assign n60677 = n46614 & ~n57657 ;
  assign n60681 = ~n60676 & ~n60677 ;
  assign n60682 = ~n60680 & n60681 ;
  assign n60683 = n27308 & ~n60682 ;
  assign n60684 = \P2_P3_EBX_reg[17]/NET0131  & ~n42872 ;
  assign n60685 = ~n60683 & ~n60684 ;
  assign n60688 = ~\P2_P3_EBX_reg[18]/NET0131  & ~n46634 ;
  assign n60689 = n27133 & ~n46635 ;
  assign n60690 = ~n60688 & n60689 ;
  assign n60686 = \P2_P3_EBX_reg[18]/NET0131  & n46615 ;
  assign n60687 = n46614 & ~n57714 ;
  assign n60691 = ~n60686 & ~n60687 ;
  assign n60692 = ~n60690 & n60691 ;
  assign n60693 = n27308 & ~n60692 ;
  assign n60694 = \P2_P3_EBX_reg[18]/NET0131  & ~n42872 ;
  assign n60695 = ~n60693 & ~n60694 ;
  assign n60698 = ~\P2_P3_EBX_reg[19]/NET0131  & ~n46635 ;
  assign n60699 = n27133 & ~n46636 ;
  assign n60700 = ~n60698 & n60699 ;
  assign n60696 = n46614 & ~n57753 ;
  assign n60697 = \P2_P3_EBX_reg[19]/NET0131  & n46615 ;
  assign n60701 = ~n60696 & ~n60697 ;
  assign n60702 = ~n60700 & n60701 ;
  assign n60703 = n27308 & ~n60702 ;
  assign n60704 = \P2_P3_EBX_reg[19]/NET0131  & ~n42872 ;
  assign n60705 = ~n60703 & ~n60704 ;
  assign n60708 = ~\P2_P3_EBX_reg[20]/NET0131  & ~n46636 ;
  assign n60709 = n27133 & ~n46637 ;
  assign n60710 = ~n60708 & n60709 ;
  assign n60706 = n46614 & ~n57799 ;
  assign n60707 = \P2_P3_EBX_reg[20]/NET0131  & n46615 ;
  assign n60711 = ~n60706 & ~n60707 ;
  assign n60712 = ~n60710 & n60711 ;
  assign n60713 = n27308 & ~n60712 ;
  assign n60714 = \P2_P3_EBX_reg[20]/NET0131  & ~n42872 ;
  assign n60715 = ~n60713 & ~n60714 ;
  assign n60718 = ~\P2_P3_EBX_reg[21]/NET0131  & ~n46637 ;
  assign n60719 = n27133 & ~n46638 ;
  assign n60720 = ~n60718 & n60719 ;
  assign n60716 = \P2_P3_EBX_reg[21]/NET0131  & n46615 ;
  assign n60717 = n46614 & ~n57856 ;
  assign n60721 = ~n60716 & ~n60717 ;
  assign n60722 = ~n60720 & n60721 ;
  assign n60723 = n27308 & ~n60722 ;
  assign n60724 = \P2_P3_EBX_reg[21]/NET0131  & ~n42872 ;
  assign n60725 = ~n60723 & ~n60724 ;
  assign n60728 = ~\P2_P3_EBX_reg[22]/NET0131  & ~n46638 ;
  assign n60729 = n27133 & ~n46639 ;
  assign n60730 = ~n60728 & n60729 ;
  assign n60726 = \P2_P3_EBX_reg[22]/NET0131  & n46615 ;
  assign n60727 = n46614 & ~n57906 ;
  assign n60731 = ~n60726 & ~n60727 ;
  assign n60732 = ~n60730 & n60731 ;
  assign n60733 = n27308 & ~n60732 ;
  assign n60734 = \P2_P3_EBX_reg[22]/NET0131  & ~n42872 ;
  assign n60735 = ~n60733 & ~n60734 ;
  assign n60736 = \P2_P3_EBX_reg[23]/NET0131  & ~n42872 ;
  assign n60739 = ~\P2_P3_EBX_reg[23]/NET0131  & ~n46639 ;
  assign n60740 = n27133 & ~n46640 ;
  assign n60741 = ~n60739 & n60740 ;
  assign n60737 = \P2_P3_EBX_reg[23]/NET0131  & n46615 ;
  assign n60738 = n46614 & n57916 ;
  assign n60742 = ~n60737 & ~n60738 ;
  assign n60743 = ~n60741 & n60742 ;
  assign n60744 = n27308 & ~n60743 ;
  assign n60745 = ~n60736 & ~n60744 ;
  assign n60748 = ~\P2_P3_EBX_reg[24]/NET0131  & ~n46640 ;
  assign n60749 = n27133 & ~n46641 ;
  assign n60750 = ~n60748 & n60749 ;
  assign n60746 = \P2_P3_EBX_reg[24]/NET0131  & n46615 ;
  assign n60747 = n46614 & n57933 ;
  assign n60751 = ~n60746 & ~n60747 ;
  assign n60752 = ~n60750 & n60751 ;
  assign n60753 = n27308 & ~n60752 ;
  assign n60754 = \P2_P3_EBX_reg[24]/NET0131  & ~n42872 ;
  assign n60755 = ~n60753 & ~n60754 ;
  assign n60758 = ~\P2_P3_EBX_reg[28]/NET0131  & ~n46645 ;
  assign n60759 = n27133 & ~n46655 ;
  assign n60760 = ~n60758 & n60759 ;
  assign n60756 = \P2_P3_EBX_reg[28]/NET0131  & n46615 ;
  assign n60757 = n46614 & n57956 ;
  assign n60761 = ~n60756 & ~n60757 ;
  assign n60762 = ~n60760 & n60761 ;
  assign n60763 = n27308 & ~n60762 ;
  assign n60764 = \P2_P3_EBX_reg[28]/NET0131  & ~n42872 ;
  assign n60765 = ~n60763 & ~n60764 ;
  assign n60767 = \P2_P3_EBX_reg[8]/NET0131  & n46615 ;
  assign n60766 = n46614 & ~n49347 ;
  assign n60768 = ~\P2_P3_EBX_reg[8]/NET0131  & ~n46624 ;
  assign n60769 = ~n46625 & ~n60768 ;
  assign n60770 = n27133 & n60769 ;
  assign n60771 = ~n60766 & ~n60770 ;
  assign n60772 = ~n60767 & n60771 ;
  assign n60773 = n27308 & ~n60772 ;
  assign n60774 = \P2_P3_EBX_reg[8]/NET0131  & ~n42872 ;
  assign n60775 = ~n60773 & ~n60774 ;
  assign n60777 = \P2_P3_EBX_reg[9]/NET0131  & n46615 ;
  assign n60776 = n46614 & ~n49389 ;
  assign n60778 = ~\P2_P3_EBX_reg[9]/NET0131  & ~n46625 ;
  assign n60779 = ~n46626 & ~n60778 ;
  assign n60780 = n27133 & n60779 ;
  assign n60781 = ~n60776 & ~n60780 ;
  assign n60782 = ~n60777 & n60781 ;
  assign n60783 = n27308 & ~n60782 ;
  assign n60784 = \P2_P3_EBX_reg[9]/NET0131  & ~n42872 ;
  assign n60785 = ~n60783 & ~n60784 ;
  assign n60786 = ~n27286 & n27308 ;
  assign n60787 = \P2_P3_Flush_reg/NET0131  & ~n42872 ;
  assign n60788 = ~n60786 & ~n60787 ;
  assign n60789 = \P2_P3_uWord_reg[0]/NET0131  & ~n47752 ;
  assign n60790 = ~\P2_P3_EAX_reg[16]/NET0131  & ~n47772 ;
  assign n60791 = ~n47773 & ~n60790 ;
  assign n60792 = n47747 & n60791 ;
  assign n60793 = n27122 & n53248 ;
  assign n60794 = ~n60792 & ~n60793 ;
  assign n60795 = n27308 & ~n60794 ;
  assign n60796 = ~n60789 & ~n60795 ;
  assign n60797 = \P2_P3_uWord_reg[10]/NET0131  & ~n47752 ;
  assign n60798 = ~n27192 & n47696 ;
  assign n60799 = \P2_P3_EAX_reg[26]/NET0131  & n47777 ;
  assign n60800 = ~\P2_P3_EAX_reg[26]/NET0131  & ~n47777 ;
  assign n60801 = ~n60799 & ~n60800 ;
  assign n60802 = n27121 & n60801 ;
  assign n60803 = ~n60798 & ~n60802 ;
  assign n60804 = n47754 & ~n60803 ;
  assign n60805 = ~n60797 & ~n60804 ;
  assign n60806 = \P2_P3_uWord_reg[13]/NET0131  & ~n47746 ;
  assign n60808 = \P2_P3_EAX_reg[28]/NET0131  & n56845 ;
  assign n60810 = \P2_P3_EAX_reg[29]/NET0131  & n60808 ;
  assign n60809 = ~\P2_P3_EAX_reg[29]/NET0131  & ~n60808 ;
  assign n60811 = n47747 & ~n60809 ;
  assign n60812 = ~n60810 & n60811 ;
  assign n60807 = \P2_P3_uWord_reg[13]/NET0131  & ~n47750 ;
  assign n60813 = ~n48264 & ~n60807 ;
  assign n60814 = ~n60812 & n60813 ;
  assign n60815 = n27308 & ~n60814 ;
  assign n60816 = ~n60806 & ~n60815 ;
  assign n60817 = \P2_P3_uWord_reg[14]/NET0131  & ~n47752 ;
  assign n60818 = n27122 & n46588 ;
  assign n60819 = \P2_P3_EAX_reg[29]/NET0131  & n47779 ;
  assign n60820 = \P2_P3_EAX_reg[30]/NET0131  & n60819 ;
  assign n60821 = ~\P2_P3_EAX_reg[30]/NET0131  & ~n60819 ;
  assign n60822 = ~n60820 & ~n60821 ;
  assign n60823 = n27121 & n60822 ;
  assign n60824 = ~n60818 & ~n60823 ;
  assign n60825 = n47754 & ~n60824 ;
  assign n60826 = ~n60817 & ~n60825 ;
  assign n60827 = \P2_P3_uWord_reg[1]/NET0131  & ~n47752 ;
  assign n60828 = ~\P2_P3_EAX_reg[17]/NET0131  & ~n47773 ;
  assign n60829 = ~n47774 & ~n60828 ;
  assign n60830 = n47747 & n60829 ;
  assign n60831 = n27122 & n57661 ;
  assign n60832 = ~n60830 & ~n60831 ;
  assign n60833 = n27308 & ~n60832 ;
  assign n60834 = ~n60827 & ~n60833 ;
  assign n60835 = \P2_P3_uWord_reg[2]/NET0131  & ~n47746 ;
  assign n60840 = \P2_P3_uWord_reg[2]/NET0131  & n47748 ;
  assign n60836 = \P2_buf2_reg[2]/NET0131  & n27227 ;
  assign n60837 = \P2_P3_uWord_reg[2]/NET0131  & n27192 ;
  assign n60838 = ~n60836 & ~n60837 ;
  assign n60839 = n27122 & ~n60838 ;
  assign n60841 = ~\P2_P3_EAX_reg[18]/NET0131  & ~n47774 ;
  assign n60842 = ~n47775 & ~n60841 ;
  assign n60843 = n47747 & n60842 ;
  assign n60844 = ~n60839 & ~n60843 ;
  assign n60845 = ~n60840 & n60844 ;
  assign n60846 = n27308 & ~n60845 ;
  assign n60847 = ~n60835 & ~n60846 ;
  assign n60848 = \P2_P3_uWord_reg[3]/NET0131  & ~n47746 ;
  assign n60853 = \P2_P3_uWord_reg[3]/NET0131  & n47748 ;
  assign n60849 = \P2_buf2_reg[3]/NET0131  & n27227 ;
  assign n60850 = \P2_P3_uWord_reg[3]/NET0131  & n27192 ;
  assign n60851 = ~n60849 & ~n60850 ;
  assign n60852 = n27122 & ~n60851 ;
  assign n60854 = ~n59547 & ~n60852 ;
  assign n60855 = ~n60853 & n60854 ;
  assign n60856 = n27308 & ~n60855 ;
  assign n60857 = ~n60848 & ~n60856 ;
  assign n60858 = \P2_P3_uWord_reg[5]/NET0131  & ~n47752 ;
  assign n60859 = n27122 & n53314 ;
  assign n60860 = ~\P2_P3_EAX_reg[21]/NET0131  & ~n48526 ;
  assign n60861 = ~n48527 & ~n60860 ;
  assign n60862 = n27121 & n60861 ;
  assign n60863 = ~n60859 & ~n60862 ;
  assign n60864 = n47754 & ~n60863 ;
  assign n60865 = ~n60858 & ~n60864 ;
  assign n60866 = \P2_P3_uWord_reg[6]/NET0131  & ~n47752 ;
  assign n60867 = \P2_buf2_reg[6]/NET0131  & ~n27192 ;
  assign n60868 = n27122 & n60867 ;
  assign n60869 = ~\P2_P3_EAX_reg[22]/NET0131  & ~n48527 ;
  assign n60870 = n27121 & ~n48528 ;
  assign n60871 = ~n60869 & n60870 ;
  assign n60872 = ~n60868 & ~n60871 ;
  assign n60873 = n47754 & ~n60872 ;
  assign n60874 = ~n60866 & ~n60873 ;
  assign n60875 = \P2_P3_uWord_reg[7]/NET0131  & ~n47752 ;
  assign n60876 = ~n27192 & n57920 ;
  assign n60877 = ~n59555 & ~n60876 ;
  assign n60878 = n47754 & ~n60877 ;
  assign n60879 = ~n60875 & ~n60878 ;
  assign n60880 = \P2_P3_uWord_reg[9]/NET0131  & ~n47746 ;
  assign n60885 = \P2_P3_uWord_reg[9]/NET0131  & n47748 ;
  assign n60881 = \P2_buf2_reg[9]/NET0131  & n27227 ;
  assign n60882 = \P2_P3_uWord_reg[9]/NET0131  & n27192 ;
  assign n60883 = ~n60881 & ~n60882 ;
  assign n60884 = n27122 & ~n60883 ;
  assign n60886 = ~\P2_P3_EAX_reg[25]/NET0131  & ~n48531 ;
  assign n60887 = ~n56842 & ~n60886 ;
  assign n60888 = n47747 & n60887 ;
  assign n60889 = ~n60884 & ~n60888 ;
  assign n60890 = ~n60885 & n60889 ;
  assign n60891 = n27308 & ~n60890 ;
  assign n60892 = ~n60880 & ~n60891 ;
  assign n60894 = \P1_P2_EBX_reg[10]/NET0131  & n46695 ;
  assign n60893 = n46694 & ~n49443 ;
  assign n60895 = ~\P1_P2_EBX_reg[10]/NET0131  & ~n46706 ;
  assign n60896 = ~n46707 & ~n60895 ;
  assign n60897 = n25803 & n60896 ;
  assign n60898 = ~n60893 & ~n60897 ;
  assign n60899 = ~n60894 & n60898 ;
  assign n60900 = n25918 & ~n60899 ;
  assign n60901 = \P1_P2_EBX_reg[10]/NET0131  & ~n43212 ;
  assign n60902 = ~n60900 & ~n60901 ;
  assign n60904 = \P1_P2_EBX_reg[11]/NET0131  & n46695 ;
  assign n60903 = n46694 & ~n49484 ;
  assign n60905 = ~\P1_P2_EBX_reg[11]/NET0131  & ~n46707 ;
  assign n60906 = ~n46708 & ~n60905 ;
  assign n60907 = n25803 & n60906 ;
  assign n60908 = ~n60903 & ~n60907 ;
  assign n60909 = ~n60904 & n60908 ;
  assign n60910 = n25918 & ~n60909 ;
  assign n60911 = \P1_P2_EBX_reg[11]/NET0131  & ~n43212 ;
  assign n60912 = ~n60910 & ~n60911 ;
  assign n60914 = \P1_P2_EBX_reg[12]/NET0131  & n46695 ;
  assign n60913 = n46694 & ~n49528 ;
  assign n60915 = ~\P1_P2_EBX_reg[12]/NET0131  & ~n46708 ;
  assign n60916 = n25803 & ~n46709 ;
  assign n60917 = ~n60915 & n60916 ;
  assign n60918 = ~n60913 & ~n60917 ;
  assign n60919 = ~n60914 & n60918 ;
  assign n60920 = n25918 & ~n60919 ;
  assign n60921 = \P1_P2_EBX_reg[12]/NET0131  & ~n43212 ;
  assign n60922 = ~n60920 & ~n60921 ;
  assign n60923 = \P1_P2_EBX_reg[13]/NET0131  & ~n43212 ;
  assign n60925 = ~n46695 & ~n60916 ;
  assign n60926 = \P1_P2_EBX_reg[13]/NET0131  & ~n60925 ;
  assign n60924 = n46694 & ~n49573 ;
  assign n60927 = ~\P1_P2_EBX_reg[13]/NET0131  & n25803 ;
  assign n60928 = n46709 & n60927 ;
  assign n60929 = ~n60924 & ~n60928 ;
  assign n60930 = ~n60926 & n60929 ;
  assign n60931 = n25918 & ~n60930 ;
  assign n60932 = ~n60923 & ~n60931 ;
  assign n60935 = ~\P1_P2_EBX_reg[14]/NET0131  & ~n46710 ;
  assign n60936 = n25803 & ~n46711 ;
  assign n60937 = ~n60935 & n60936 ;
  assign n60933 = n46694 & ~n49616 ;
  assign n60934 = \P1_P2_EBX_reg[14]/NET0131  & n46695 ;
  assign n60938 = ~n60933 & ~n60934 ;
  assign n60939 = ~n60937 & n60938 ;
  assign n60940 = n25918 & ~n60939 ;
  assign n60941 = \P1_P2_EBX_reg[14]/NET0131  & ~n43212 ;
  assign n60942 = ~n60940 & ~n60941 ;
  assign n60945 = ~\P1_P2_EBX_reg[15]/NET0131  & ~n46711 ;
  assign n60946 = n25803 & ~n46712 ;
  assign n60947 = ~n60945 & n60946 ;
  assign n60943 = n46694 & ~n48324 ;
  assign n60944 = \P1_P2_EBX_reg[15]/NET0131  & n46695 ;
  assign n60948 = ~n60943 & ~n60944 ;
  assign n60949 = ~n60947 & n60948 ;
  assign n60950 = n25918 & ~n60949 ;
  assign n60951 = \P1_P2_EBX_reg[15]/NET0131  & ~n43212 ;
  assign n60952 = ~n60950 & ~n60951 ;
  assign n60955 = ~\P1_P2_EBX_reg[16]/NET0131  & ~n46712 ;
  assign n60956 = n25803 & ~n46713 ;
  assign n60957 = ~n60955 & n60956 ;
  assign n60953 = n46694 & ~n58009 ;
  assign n60954 = \P1_P2_EBX_reg[16]/NET0131  & n46695 ;
  assign n60958 = ~n60953 & ~n60954 ;
  assign n60959 = ~n60957 & n60958 ;
  assign n60960 = n25918 & ~n60959 ;
  assign n60961 = \P1_P2_EBX_reg[16]/NET0131  & ~n43212 ;
  assign n60962 = ~n60960 & ~n60961 ;
  assign n60965 = ~\P1_P2_EBX_reg[17]/NET0131  & ~n46713 ;
  assign n60966 = n25803 & ~n46714 ;
  assign n60967 = ~n60965 & n60966 ;
  assign n60963 = \P1_P2_EBX_reg[17]/NET0131  & n46695 ;
  assign n60964 = n46694 & ~n58056 ;
  assign n60968 = ~n60963 & ~n60964 ;
  assign n60969 = ~n60967 & n60968 ;
  assign n60970 = n25918 & ~n60969 ;
  assign n60971 = \P1_P2_EBX_reg[17]/NET0131  & ~n43212 ;
  assign n60972 = ~n60970 & ~n60971 ;
  assign n60975 = ~\P1_P2_EBX_reg[19]/NET0131  & ~n46715 ;
  assign n60976 = n25803 & ~n46716 ;
  assign n60977 = ~n60975 & n60976 ;
  assign n60973 = \P1_P2_EBX_reg[19]/NET0131  & n46695 ;
  assign n60974 = n46694 & ~n58149 ;
  assign n60978 = ~n60973 & ~n60974 ;
  assign n60979 = ~n60977 & n60978 ;
  assign n60980 = n25918 & ~n60979 ;
  assign n60981 = \P1_P2_EBX_reg[19]/NET0131  & ~n43212 ;
  assign n60982 = ~n60980 & ~n60981 ;
  assign n60985 = ~\P1_P2_EBX_reg[20]/NET0131  & ~n46716 ;
  assign n60986 = n25803 & ~n46717 ;
  assign n60987 = ~n60985 & n60986 ;
  assign n60983 = n46694 & ~n58201 ;
  assign n60984 = \P1_P2_EBX_reg[20]/NET0131  & n46695 ;
  assign n60988 = ~n60983 & ~n60984 ;
  assign n60989 = ~n60987 & n60988 ;
  assign n60990 = n25918 & ~n60989 ;
  assign n60991 = \P1_P2_EBX_reg[20]/NET0131  & ~n43212 ;
  assign n60992 = ~n60990 & ~n60991 ;
  assign n60995 = ~\P1_P2_EBX_reg[21]/NET0131  & ~n46717 ;
  assign n60996 = n25803 & ~n46718 ;
  assign n60997 = ~n60995 & n60996 ;
  assign n60993 = \P1_P2_EBX_reg[21]/NET0131  & n46695 ;
  assign n60994 = n46694 & ~n58244 ;
  assign n60998 = ~n60993 & ~n60994 ;
  assign n60999 = ~n60997 & n60998 ;
  assign n61000 = n25918 & ~n60999 ;
  assign n61001 = \P1_P2_EBX_reg[21]/NET0131  & ~n43212 ;
  assign n61002 = ~n61000 & ~n61001 ;
  assign n61005 = ~\P1_P2_EBX_reg[22]/NET0131  & ~n46718 ;
  assign n61006 = n25803 & ~n46719 ;
  assign n61007 = ~n61005 & n61006 ;
  assign n61003 = \P1_P2_EBX_reg[22]/NET0131  & n46695 ;
  assign n61004 = n46694 & ~n58287 ;
  assign n61008 = ~n61003 & ~n61004 ;
  assign n61009 = ~n61007 & n61008 ;
  assign n61010 = n25918 & ~n61009 ;
  assign n61011 = \P1_P2_EBX_reg[22]/NET0131  & ~n43212 ;
  assign n61012 = ~n61010 & ~n61011 ;
  assign n61013 = \P1_P2_EBX_reg[23]/NET0131  & ~n43212 ;
  assign n61016 = ~\P1_P2_EBX_reg[23]/NET0131  & ~n46719 ;
  assign n61017 = n25803 & ~n46720 ;
  assign n61018 = ~n61016 & n61017 ;
  assign n61014 = n46694 & n58306 ;
  assign n61015 = \P1_P2_EBX_reg[23]/NET0131  & n46695 ;
  assign n61019 = ~n61014 & ~n61015 ;
  assign n61020 = ~n61018 & n61019 ;
  assign n61021 = n25918 & ~n61020 ;
  assign n61022 = ~n61013 & ~n61021 ;
  assign n61025 = ~\P1_P2_EBX_reg[24]/NET0131  & ~n46720 ;
  assign n61026 = n25803 & ~n46721 ;
  assign n61027 = ~n61025 & n61026 ;
  assign n61023 = n46694 & n58324 ;
  assign n61024 = \P1_P2_EBX_reg[24]/NET0131  & n46695 ;
  assign n61028 = ~n61023 & ~n61024 ;
  assign n61029 = ~n61027 & n61028 ;
  assign n61030 = n25918 & ~n61029 ;
  assign n61031 = \P1_P2_EBX_reg[24]/NET0131  & ~n43212 ;
  assign n61032 = ~n61030 & ~n61031 ;
  assign n61035 = ~\P1_P2_EBX_reg[28]/NET0131  & ~n46724 ;
  assign n61036 = n25803 & ~n46736 ;
  assign n61037 = ~n61035 & n61036 ;
  assign n61033 = \P1_P2_EBX_reg[28]/NET0131  & n46695 ;
  assign n61034 = n46694 & n58339 ;
  assign n61038 = ~n61033 & ~n61034 ;
  assign n61039 = ~n61037 & n61038 ;
  assign n61040 = n25918 & ~n61039 ;
  assign n61041 = \P1_P2_EBX_reg[28]/NET0131  & ~n43212 ;
  assign n61042 = ~n61040 & ~n61041 ;
  assign n61044 = \P1_P2_EBX_reg[8]/NET0131  & n46695 ;
  assign n61043 = n46694 & ~n49676 ;
  assign n61045 = ~\P1_P2_EBX_reg[8]/NET0131  & ~n46704 ;
  assign n61046 = ~n46705 & ~n61045 ;
  assign n61047 = n25803 & n61046 ;
  assign n61048 = ~n61043 & ~n61047 ;
  assign n61049 = ~n61044 & n61048 ;
  assign n61050 = n25918 & ~n61049 ;
  assign n61051 = \P1_P2_EBX_reg[8]/NET0131  & ~n43212 ;
  assign n61052 = ~n61050 & ~n61051 ;
  assign n61054 = \P1_P2_EBX_reg[9]/NET0131  & n46695 ;
  assign n61053 = n46694 & ~n49717 ;
  assign n61055 = ~\P1_P2_EBX_reg[9]/NET0131  & ~n46705 ;
  assign n61056 = ~n46706 & ~n61055 ;
  assign n61057 = n25803 & n61056 ;
  assign n61058 = ~n61053 & ~n61057 ;
  assign n61059 = ~n61054 & n61058 ;
  assign n61060 = n25918 & ~n61059 ;
  assign n61061 = \P1_P2_EBX_reg[9]/NET0131  & ~n43212 ;
  assign n61062 = ~n61060 & ~n61061 ;
  assign n61064 = \P1_P1_Datao_reg[30]/NET0131  & ~n26162 ;
  assign n61065 = n25362 & ~n26158 ;
  assign n61066 = ~n61064 & ~n61065 ;
  assign n61067 = n8355 & ~n61066 ;
  assign n61063 = \P1_P1_uWord_reg[14]/NET0131  & n27790 ;
  assign n61068 = \P1_P1_Datao_reg[30]/NET0131  & ~n48479 ;
  assign n61069 = ~n61063 & ~n61068 ;
  assign n61070 = ~n61067 & n61069 ;
  assign n61073 = \P2_P2_CodeFetch_reg/NET0131  & n26792 ;
  assign n61074 = ~n26697 & n61073 ;
  assign n61075 = ~n26698 & n61074 ;
  assign n61071 = ~n27614 & ~n48507 ;
  assign n61072 = \P2_P2_CodeFetch_reg/NET0131  & ~n61071 ;
  assign n61076 = ~n26292 & ~n61072 ;
  assign n61077 = ~n61075 & n61076 ;
  assign n61079 = \P2_P2_Datao_reg[30]/NET0131  & ~n26699 ;
  assign n61080 = n26692 & n60535 ;
  assign n61081 = ~n61079 & ~n61080 ;
  assign n61082 = n26792 & ~n61081 ;
  assign n61078 = \P2_P2_uWord_reg[14]/NET0131  & n48491 ;
  assign n61083 = \P2_P2_Datao_reg[30]/NET0131  & ~n48508 ;
  assign n61084 = ~n61078 & ~n61083 ;
  assign n61085 = ~n61082 & n61084 ;
  assign n61086 = ~n9195 & n9241 ;
  assign n61087 = n22872 & ~n61086 ;
  assign n61088 = \P1_P3_CodeFetch_reg/NET0131  & ~n61087 ;
  assign n61089 = ~n9247 & ~n61088 ;
  assign n61091 = n9162 & n22895 ;
  assign n61092 = \P1_P3_Datao_reg[30]/NET0131  & ~n9165 ;
  assign n61093 = ~n61091 & ~n61092 ;
  assign n61094 = n9241 & ~n61093 ;
  assign n61095 = ~n9245 & ~n10037 ;
  assign n61096 = n16493 & n61095 ;
  assign n61097 = \P1_P3_Datao_reg[30]/NET0131  & ~n61096 ;
  assign n61090 = \P1_P3_uWord_reg[14]/NET0131  & n43256 ;
  assign n61098 = \P1_P3_Datao_reg[30]/NET0131  & ~n8731 ;
  assign n61099 = n10029 & n61098 ;
  assign n61100 = ~n61090 & ~n61099 ;
  assign n61101 = ~n61097 & n61100 ;
  assign n61102 = ~n61094 & n61101 ;
  assign n61105 = \P2_P3_CodeFetch_reg/NET0131  & n27308 ;
  assign n61106 = ~n27256 & n61105 ;
  assign n61107 = ~n54647 & n61106 ;
  assign n61103 = ~n27649 & n32869 ;
  assign n61104 = \P2_P3_CodeFetch_reg/NET0131  & ~n61103 ;
  assign n61108 = ~n27311 & ~n61104 ;
  assign n61109 = ~n61107 & n61108 ;
  assign n61112 = \P1_P2_CodeFetch_reg/NET0131  & n25918 ;
  assign n61113 = ~n48371 & n61112 ;
  assign n61110 = ~n27606 & n31486 ;
  assign n61111 = \P1_P2_CodeFetch_reg/NET0131  & ~n61110 ;
  assign n61114 = ~n25418 & ~n61111 ;
  assign n61115 = ~n61113 & n61114 ;
  assign n61117 = \P2_P3_Datao_reg[30]/NET0131  & ~n27223 ;
  assign n61118 = n27303 & n60822 ;
  assign n61119 = ~n61117 & ~n61118 ;
  assign n61120 = n27308 & ~n61119 ;
  assign n61116 = \P2_P3_uWord_reg[14]/NET0131  & n48523 ;
  assign n61121 = \P2_P3_Datao_reg[30]/NET0131  & ~n48540 ;
  assign n61122 = ~n61116 & ~n61121 ;
  assign n61123 = ~n61120 & n61122 ;
  assign n61126 = \P1_P1_CodeFetch_reg/NET0131  & n8355 ;
  assign n61127 = ~n50559 & n61126 ;
  assign n61124 = ~n8348 & n34163 ;
  assign n61125 = \P1_P1_CodeFetch_reg/NET0131  & ~n61124 ;
  assign n61128 = ~n8359 & ~n61125 ;
  assign n61129 = ~n61127 & n61128 ;
  assign n61131 = ~n25768 & n59858 ;
  assign n61132 = n47570 & ~n61131 ;
  assign n61133 = n48554 & ~n61132 ;
  assign n61134 = \P1_P2_Datao_reg[30]/NET0131  & ~n61133 ;
  assign n61135 = n25841 & n59859 ;
  assign n61136 = ~n61134 & ~n61135 ;
  assign n61137 = n25918 & ~n61136 ;
  assign n61130 = \P1_P2_uWord_reg[14]/NET0131  & n25922 ;
  assign n61138 = \P1_P2_Datao_reg[30]/NET0131  & ~n48566 ;
  assign n61139 = ~n61130 & ~n61138 ;
  assign n61140 = ~n61137 & n61139 ;
  assign n61141 = \P2_P3_lWord_reg[0]/NET0131  & ~n47752 ;
  assign n61142 = \P2_P3_EAX_reg[0]/NET0131  & n47747 ;
  assign n61143 = ~n60793 & ~n61142 ;
  assign n61144 = n27308 & ~n61143 ;
  assign n61145 = ~n61141 & ~n61144 ;
  assign n61146 = \P2_P3_lWord_reg[10]/NET0131  & n47748 ;
  assign n61147 = \P2_buf2_reg[10]/NET0131  & n27227 ;
  assign n61148 = \P2_P3_lWord_reg[10]/NET0131  & n27192 ;
  assign n61149 = ~n61147 & ~n61148 ;
  assign n61150 = n27122 & ~n61149 ;
  assign n61151 = \P2_P3_EAX_reg[10]/NET0131  & n47747 ;
  assign n61152 = ~n61150 & ~n61151 ;
  assign n61153 = ~n61146 & n61152 ;
  assign n61154 = n27308 & ~n61153 ;
  assign n61155 = \P2_P3_lWord_reg[10]/NET0131  & ~n47746 ;
  assign n61156 = ~n61154 & ~n61155 ;
  assign n61157 = \P2_P3_lWord_reg[11]/NET0131  & ~n47752 ;
  assign n61158 = \P2_P3_EAX_reg[11]/NET0131  & n47747 ;
  assign n61159 = ~n58353 & ~n61158 ;
  assign n61160 = n27308 & ~n61159 ;
  assign n61161 = ~n61157 & ~n61160 ;
  assign n61162 = \P2_P3_lWord_reg[12]/NET0131  & n47748 ;
  assign n61163 = \P2_P3_lWord_reg[12]/NET0131  & n27192 ;
  assign n61164 = \P2_buf2_reg[12]/NET0131  & n27227 ;
  assign n61165 = ~n61163 & ~n61164 ;
  assign n61166 = n27122 & ~n61165 ;
  assign n61167 = \P2_P3_EAX_reg[12]/NET0131  & n47747 ;
  assign n61168 = ~n61166 & ~n61167 ;
  assign n61169 = ~n61162 & n61168 ;
  assign n61170 = n27308 & ~n61169 ;
  assign n61171 = \P2_P3_lWord_reg[12]/NET0131  & ~n47746 ;
  assign n61172 = ~n61170 & ~n61171 ;
  assign n61173 = \P2_P3_lWord_reg[13]/NET0131  & n47748 ;
  assign n61174 = \P2_P3_lWord_reg[13]/NET0131  & n27192 ;
  assign n61175 = ~n49206 & ~n61174 ;
  assign n61176 = n27122 & ~n61175 ;
  assign n61177 = \P2_P3_EAX_reg[13]/NET0131  & n47747 ;
  assign n61178 = ~n61176 & ~n61177 ;
  assign n61179 = ~n61173 & n61178 ;
  assign n61180 = n27308 & ~n61179 ;
  assign n61181 = \P2_P3_lWord_reg[13]/NET0131  & ~n47746 ;
  assign n61182 = ~n61180 & ~n61181 ;
  assign n61183 = \P2_P3_lWord_reg[14]/NET0131  & n47748 ;
  assign n61184 = \P2_P3_lWord_reg[14]/NET0131  & n27192 ;
  assign n61185 = ~n49253 & ~n61184 ;
  assign n61186 = n27122 & ~n61185 ;
  assign n61187 = \P2_P3_EAX_reg[14]/NET0131  & n47747 ;
  assign n61188 = ~n61186 & ~n61187 ;
  assign n61189 = ~n61183 & n61188 ;
  assign n61190 = n27308 & ~n61189 ;
  assign n61191 = \P2_P3_lWord_reg[14]/NET0131  & ~n47746 ;
  assign n61192 = ~n61190 & ~n61191 ;
  assign n61193 = \P2_P3_lWord_reg[15]/NET0131  & n47748 ;
  assign n61194 = \P2_P3_lWord_reg[15]/NET0131  & n27192 ;
  assign n61195 = ~n49298 & ~n61194 ;
  assign n61196 = n27122 & ~n61195 ;
  assign n61197 = \P2_P3_EAX_reg[15]/NET0131  & n47747 ;
  assign n61198 = ~n61196 & ~n61197 ;
  assign n61199 = ~n61193 & n61198 ;
  assign n61200 = n27308 & ~n61199 ;
  assign n61201 = \P2_P3_lWord_reg[15]/NET0131  & ~n47746 ;
  assign n61202 = ~n61200 & ~n61201 ;
  assign n61203 = \P2_P3_lWord_reg[1]/NET0131  & ~n47752 ;
  assign n61204 = \P2_P3_EAX_reg[1]/NET0131  & n47747 ;
  assign n61205 = ~n60831 & ~n61204 ;
  assign n61206 = n27308 & ~n61205 ;
  assign n61207 = ~n61203 & ~n61206 ;
  assign n61208 = \P2_P3_lWord_reg[2]/NET0131  & n47748 ;
  assign n61209 = \P2_P3_lWord_reg[2]/NET0131  & n27192 ;
  assign n61210 = ~n60836 & ~n61209 ;
  assign n61211 = n27122 & ~n61210 ;
  assign n61212 = \P2_P3_EAX_reg[2]/NET0131  & n47747 ;
  assign n61213 = ~n61211 & ~n61212 ;
  assign n61214 = ~n61208 & n61213 ;
  assign n61215 = n27308 & ~n61214 ;
  assign n61216 = \P2_P3_lWord_reg[2]/NET0131  & ~n47746 ;
  assign n61217 = ~n61215 & ~n61216 ;
  assign n61218 = \P2_P3_lWord_reg[3]/NET0131  & n47748 ;
  assign n61219 = \P2_P3_lWord_reg[3]/NET0131  & n27192 ;
  assign n61220 = ~n60849 & ~n61219 ;
  assign n61221 = n27122 & ~n61220 ;
  assign n61222 = \P2_P3_EAX_reg[3]/NET0131  & n47747 ;
  assign n61223 = ~n61221 & ~n61222 ;
  assign n61224 = ~n61218 & n61223 ;
  assign n61225 = n27308 & ~n61224 ;
  assign n61226 = \P2_P3_lWord_reg[3]/NET0131  & ~n47746 ;
  assign n61227 = ~n61225 & ~n61226 ;
  assign n61228 = \P2_P3_lWord_reg[4]/NET0131  & ~n47752 ;
  assign n61229 = \P2_P3_EAX_reg[4]/NET0131  & n47747 ;
  assign n61230 = ~n53435 & ~n61229 ;
  assign n61231 = n27308 & ~n61230 ;
  assign n61232 = ~n61228 & ~n61231 ;
  assign n61233 = \P2_P3_lWord_reg[5]/NET0131  & n47748 ;
  assign n61234 = \P2_P3_lWord_reg[5]/NET0131  & n27192 ;
  assign n61235 = \P2_buf2_reg[5]/NET0131  & n27227 ;
  assign n61236 = ~n61234 & ~n61235 ;
  assign n61237 = n27122 & ~n61236 ;
  assign n61238 = \P2_P3_EAX_reg[5]/NET0131  & n47747 ;
  assign n61239 = ~n61237 & ~n61238 ;
  assign n61240 = ~n61233 & n61239 ;
  assign n61241 = n27308 & ~n61240 ;
  assign n61242 = \P2_P3_lWord_reg[5]/NET0131  & ~n47746 ;
  assign n61243 = ~n61241 & ~n61242 ;
  assign n61244 = \P2_P3_lWord_reg[6]/NET0131  & ~n47752 ;
  assign n61245 = \P2_P3_EAX_reg[6]/NET0131  & n47747 ;
  assign n61246 = n46587 & n60867 ;
  assign n61247 = ~n61245 & ~n61246 ;
  assign n61248 = n27308 & ~n61247 ;
  assign n61249 = ~n61244 & ~n61248 ;
  assign n61250 = \P2_P3_lWord_reg[7]/NET0131  & n47748 ;
  assign n61251 = \P2_buf2_reg[7]/NET0131  & n27227 ;
  assign n61252 = \P2_P3_lWord_reg[7]/NET0131  & n27192 ;
  assign n61253 = ~n61251 & ~n61252 ;
  assign n61254 = n27122 & ~n61253 ;
  assign n61255 = \P2_P3_EAX_reg[7]/NET0131  & n47747 ;
  assign n61256 = ~n61254 & ~n61255 ;
  assign n61257 = ~n61250 & n61256 ;
  assign n61258 = n27308 & ~n61257 ;
  assign n61259 = \P2_P3_lWord_reg[7]/NET0131  & ~n47746 ;
  assign n61260 = ~n61258 & ~n61259 ;
  assign n61261 = \P2_P3_lWord_reg[8]/NET0131  & n47748 ;
  assign n61262 = \P2_buf2_reg[8]/NET0131  & n27227 ;
  assign n61263 = \P2_P3_lWord_reg[8]/NET0131  & n27192 ;
  assign n61264 = ~n61262 & ~n61263 ;
  assign n61265 = n27122 & ~n61264 ;
  assign n61266 = \P2_P3_EAX_reg[8]/NET0131  & n47747 ;
  assign n61267 = ~n61265 & ~n61266 ;
  assign n61268 = ~n61261 & n61267 ;
  assign n61269 = n27308 & ~n61268 ;
  assign n61270 = \P2_P3_lWord_reg[8]/NET0131  & ~n47746 ;
  assign n61271 = ~n61269 & ~n61270 ;
  assign n61272 = \P2_P3_lWord_reg[9]/NET0131  & n47748 ;
  assign n61273 = \P2_P3_lWord_reg[9]/NET0131  & n27192 ;
  assign n61274 = ~n60881 & ~n61273 ;
  assign n61275 = n27122 & ~n61274 ;
  assign n61276 = \P2_P3_EAX_reg[9]/NET0131  & n47747 ;
  assign n61277 = ~n61275 & ~n61276 ;
  assign n61278 = ~n61272 & n61277 ;
  assign n61279 = n27308 & ~n61278 ;
  assign n61280 = \P2_P3_lWord_reg[9]/NET0131  & ~n47746 ;
  assign n61281 = ~n61279 & ~n61280 ;
  assign n61284 = \P2_P1_CodeFetch_reg/NET0131  & n11623 ;
  assign n61285 = ~n50414 & n61284 ;
  assign n61282 = ~n11615 & n32171 ;
  assign n61283 = \P2_P1_CodeFetch_reg/NET0131  & ~n61282 ;
  assign n61286 = ~n11618 & ~n61283 ;
  assign n61287 = ~n61285 & n61286 ;
  assign n61289 = \P2_P1_Datao_reg[30]/NET0131  & ~n26030 ;
  assign n61290 = n26006 & n27405 ;
  assign n61291 = ~n61289 & ~n61290 ;
  assign n61292 = n11623 & ~n61291 ;
  assign n61288 = \P2_P1_uWord_reg[14]/NET0131  & n48581 ;
  assign n61293 = \P2_P1_Datao_reg[30]/NET0131  & ~n48594 ;
  assign n61294 = ~n61288 & ~n61293 ;
  assign n61295 = ~n61292 & n61294 ;
  assign n61297 = \P1_P2_EBX_reg[5]/NET0131  & n46695 ;
  assign n61296 = \P1_P2_InstQueue_reg[0][5]/NET0131  & n46694 ;
  assign n61298 = ~\P1_P2_EBX_reg[5]/NET0131  & ~n46701 ;
  assign n61299 = n25803 & ~n46702 ;
  assign n61300 = ~n61298 & n61299 ;
  assign n61301 = ~n61296 & ~n61300 ;
  assign n61302 = ~n61297 & n61301 ;
  assign n61303 = n25918 & ~n61302 ;
  assign n61304 = \P1_P2_EBX_reg[5]/NET0131  & ~n43212 ;
  assign n61305 = ~n61303 & ~n61304 ;
  assign n61306 = n11623 & n46227 ;
  assign n61307 = n21100 & ~n61306 ;
  assign n61308 = \P2_P1_EBX_reg[0]/NET0131  & ~n61307 ;
  assign n61309 = ~\P2_P1_EBX_reg[0]/NET0131  & n25981 ;
  assign n61310 = \P2_P1_InstQueue_reg[0][0]/NET0131  & n46225 ;
  assign n61311 = ~n61309 & ~n61310 ;
  assign n61312 = n11623 & ~n61311 ;
  assign n61313 = ~n61308 & ~n61312 ;
  assign n61315 = \P2_P1_EBX_reg[1]/NET0131  & n48137 ;
  assign n61314 = n25981 & n50424 ;
  assign n61316 = ~\P2_P1_EBX_reg[1]/NET0131  & ~n20720 ;
  assign n61317 = ~\P2_P1_InstQueue_reg[0][1]/NET0131  & n20720 ;
  assign n61318 = ~n61316 & ~n61317 ;
  assign n61319 = n25986 & n61318 ;
  assign n61320 = ~n61314 & ~n61319 ;
  assign n61321 = ~n61315 & n61320 ;
  assign n61322 = n11623 & ~n61321 ;
  assign n61323 = \P2_P1_EBX_reg[1]/NET0131  & ~n21100 ;
  assign n61324 = ~n61322 & ~n61323 ;
  assign n61325 = \P2_P1_EBX_reg[2]/NET0131  & ~n21100 ;
  assign n61327 = n25981 & ~n46230 ;
  assign n61328 = ~n46227 & ~n61327 ;
  assign n61329 = \P2_P1_EBX_reg[2]/NET0131  & ~n61328 ;
  assign n61326 = \P2_P1_InstQueue_reg[0][2]/NET0131  & n46225 ;
  assign n61330 = ~\P2_P1_EBX_reg[2]/NET0131  & n46230 ;
  assign n61331 = n25981 & n61330 ;
  assign n61332 = ~n61326 & ~n61331 ;
  assign n61333 = ~n61329 & n61332 ;
  assign n61334 = n11623 & ~n61333 ;
  assign n61335 = ~n61325 & ~n61334 ;
  assign n61340 = \P2_P1_EBX_reg[3]/NET0131  & n48137 ;
  assign n61336 = ~\P2_P1_EBX_reg[3]/NET0131  & ~n20720 ;
  assign n61337 = ~\P2_P1_InstQueue_reg[0][3]/NET0131  & n20720 ;
  assign n61338 = ~n61336 & ~n61337 ;
  assign n61339 = n25986 & n61338 ;
  assign n61341 = ~\P2_P1_EBX_reg[3]/NET0131  & ~n46231 ;
  assign n61342 = n25981 & ~n46232 ;
  assign n61343 = ~n61341 & n61342 ;
  assign n61344 = ~n61339 & ~n61343 ;
  assign n61345 = ~n61340 & n61344 ;
  assign n61346 = n11623 & ~n61345 ;
  assign n61347 = \P2_P1_EBX_reg[3]/NET0131  & ~n21100 ;
  assign n61348 = ~n61346 & ~n61347 ;
  assign n61349 = \P2_P1_EBX_reg[4]/NET0131  & ~n21100 ;
  assign n61351 = ~n46227 & ~n61342 ;
  assign n61352 = \P2_P1_EBX_reg[4]/NET0131  & ~n61351 ;
  assign n61350 = \P2_P1_InstQueue_reg[0][4]/NET0131  & n46225 ;
  assign n61353 = ~\P2_P1_EBX_reg[4]/NET0131  & n46232 ;
  assign n61354 = n25981 & n61353 ;
  assign n61355 = ~n61350 & ~n61354 ;
  assign n61356 = ~n61352 & n61355 ;
  assign n61357 = n11623 & ~n61356 ;
  assign n61358 = ~n61349 & ~n61357 ;
  assign n61363 = \P2_P1_EBX_reg[5]/NET0131  & n48137 ;
  assign n61359 = ~\P2_P1_EBX_reg[5]/NET0131  & ~n20720 ;
  assign n61360 = ~\P2_P1_InstQueue_reg[0][5]/NET0131  & n20720 ;
  assign n61361 = ~n61359 & ~n61360 ;
  assign n61362 = n25986 & n61361 ;
  assign n61364 = ~\P2_P1_EBX_reg[5]/NET0131  & ~n46233 ;
  assign n61365 = n25981 & ~n46234 ;
  assign n61366 = ~n61364 & n61365 ;
  assign n61367 = ~n61362 & ~n61366 ;
  assign n61368 = ~n61363 & n61367 ;
  assign n61369 = n11623 & ~n61368 ;
  assign n61370 = \P2_P1_EBX_reg[5]/NET0131  & ~n21100 ;
  assign n61371 = ~n61369 & ~n61370 ;
  assign n61372 = \P2_P1_EBX_reg[6]/NET0131  & ~n21100 ;
  assign n61374 = ~n46227 & ~n61365 ;
  assign n61375 = \P2_P1_EBX_reg[6]/NET0131  & ~n61374 ;
  assign n61373 = \P2_P1_InstQueue_reg[0][6]/NET0131  & n46225 ;
  assign n61376 = ~\P2_P1_EBX_reg[6]/NET0131  & n46234 ;
  assign n61377 = n25981 & n61376 ;
  assign n61378 = ~n61373 & ~n61377 ;
  assign n61379 = ~n61375 & n61378 ;
  assign n61380 = n11623 & ~n61379 ;
  assign n61381 = ~n61372 & ~n61380 ;
  assign n61385 = \P2_P1_EBX_reg[7]/NET0131  & n48137 ;
  assign n61382 = ~\P2_P1_EBX_reg[7]/NET0131  & ~n46235 ;
  assign n61383 = ~n46236 & ~n61382 ;
  assign n61384 = n25981 & n61383 ;
  assign n61386 = ~\P2_P1_EBX_reg[7]/NET0131  & ~n20720 ;
  assign n61387 = ~\P2_P1_InstQueue_reg[0][7]/NET0131  & n20720 ;
  assign n61388 = ~n61386 & ~n61387 ;
  assign n61389 = n25986 & n61388 ;
  assign n61390 = ~n61384 & ~n61389 ;
  assign n61391 = ~n61385 & n61390 ;
  assign n61392 = n11623 & ~n61391 ;
  assign n61393 = \P2_P1_EBX_reg[7]/NET0131  & ~n21100 ;
  assign n61394 = ~n61392 & ~n61393 ;
  assign n61395 = \P2_P1_lWord_reg[0]/NET0131  & ~n34408 ;
  assign n61396 = \P2_P1_EAX_reg[0]/NET0131  & n24899 ;
  assign n61397 = ~n59806 & ~n61396 ;
  assign n61398 = n11623 & ~n61397 ;
  assign n61399 = ~n61395 & ~n61398 ;
  assign n61400 = \P2_P1_lWord_reg[1]/NET0131  & ~n34408 ;
  assign n61401 = \P2_P1_EAX_reg[1]/NET0131  & n24899 ;
  assign n61402 = ~n59815 & ~n61401 ;
  assign n61403 = n11623 & ~n61402 ;
  assign n61404 = ~n61400 & ~n61403 ;
  assign n61405 = n26792 & n46417 ;
  assign n61406 = n44508 & ~n61405 ;
  assign n61407 = \P2_P2_EBX_reg[0]/NET0131  & ~n61406 ;
  assign n61408 = ~\P2_P2_EBX_reg[0]/NET0131  & n26662 ;
  assign n61409 = \P2_P2_InstQueue_reg[0][0]/NET0131  & n46416 ;
  assign n61410 = ~n61408 & ~n61409 ;
  assign n61411 = n26792 & ~n61410 ;
  assign n61412 = ~n61407 & ~n61411 ;
  assign n61413 = \P1_P1_EAX_reg[0]/NET0131  & n24502 ;
  assign n61414 = ~n60435 & ~n61413 ;
  assign n61415 = ~n15364 & ~n61414 ;
  assign n61416 = \P1_P1_lWord_reg[0]/NET0131  & ~n24506 ;
  assign n61417 = ~n61415 & ~n61416 ;
  assign n61418 = n8355 & ~n61417 ;
  assign n61419 = \P1_P1_lWord_reg[0]/NET0131  & ~n24515 ;
  assign n61420 = ~n61418 & ~n61419 ;
  assign n61422 = ~n26578 & ~n26662 ;
  assign n61423 = \P2_P2_EBX_reg[1]/NET0131  & n61422 ;
  assign n61421 = n26662 & n50651 ;
  assign n61424 = ~\P2_P2_EBX_reg[1]/NET0131  & ~n26611 ;
  assign n61425 = ~\P2_P2_InstQueue_reg[0][1]/NET0131  & n26611 ;
  assign n61426 = ~n61424 & ~n61425 ;
  assign n61427 = n26578 & n61426 ;
  assign n61428 = ~n61421 & ~n61427 ;
  assign n61429 = ~n61423 & n61428 ;
  assign n61430 = n26792 & ~n61429 ;
  assign n61431 = \P2_P2_EBX_reg[1]/NET0131  & ~n44508 ;
  assign n61432 = ~n61430 & ~n61431 ;
  assign n61433 = \P2_P2_EBX_reg[2]/NET0131  & ~n44508 ;
  assign n61437 = ~n26662 & n46416 ;
  assign n61435 = n26662 & n46420 ;
  assign n61438 = \P2_P2_EBX_reg[2]/NET0131  & ~n61435 ;
  assign n61439 = ~n61437 & n61438 ;
  assign n61434 = \P2_P2_InstQueue_reg[0][2]/NET0131  & n46416 ;
  assign n61436 = ~\P2_P2_EBX_reg[2]/NET0131  & n61435 ;
  assign n61440 = ~n61434 & ~n61436 ;
  assign n61441 = ~n61439 & n61440 ;
  assign n61442 = n26792 & ~n61441 ;
  assign n61443 = ~n61433 & ~n61442 ;
  assign n61448 = ~n26578 & n26662 ;
  assign n61449 = ~n46416 & ~n61448 ;
  assign n61450 = \P2_P2_EBX_reg[3]/NET0131  & n61449 ;
  assign n61444 = \P2_P2_InstQueue_reg[0][3]/NET0131  & n46416 ;
  assign n61445 = ~\P2_P2_EBX_reg[3]/NET0131  & ~n46421 ;
  assign n61446 = ~n46422 & ~n61445 ;
  assign n61447 = n26662 & n61446 ;
  assign n61451 = ~n61444 & ~n61447 ;
  assign n61452 = ~n61450 & n61451 ;
  assign n61453 = n26792 & ~n61452 ;
  assign n61454 = \P2_P2_EBX_reg[3]/NET0131  & ~n44508 ;
  assign n61455 = ~n61453 & ~n61454 ;
  assign n61456 = \P2_P2_EBX_reg[4]/NET0131  & ~n44508 ;
  assign n61458 = n26662 & n46422 ;
  assign n61460 = \P2_P2_EBX_reg[4]/NET0131  & ~n61458 ;
  assign n61461 = ~n61437 & n61460 ;
  assign n61457 = \P2_P2_InstQueue_reg[0][4]/NET0131  & n46416 ;
  assign n61459 = ~\P2_P2_EBX_reg[4]/NET0131  & n61458 ;
  assign n61462 = ~n61457 & ~n61459 ;
  assign n61463 = ~n61461 & n61462 ;
  assign n61464 = n26792 & ~n61463 ;
  assign n61465 = ~n61456 & ~n61464 ;
  assign n61470 = \P2_P2_EBX_reg[5]/NET0131  & n61449 ;
  assign n61466 = \P2_P2_InstQueue_reg[0][5]/NET0131  & n46416 ;
  assign n61467 = ~\P2_P2_EBX_reg[5]/NET0131  & ~n46423 ;
  assign n61468 = ~n46424 & ~n61467 ;
  assign n61469 = n26662 & n61468 ;
  assign n61471 = ~n61466 & ~n61469 ;
  assign n61472 = ~n61470 & n61471 ;
  assign n61473 = n26792 & ~n61472 ;
  assign n61474 = \P2_P2_EBX_reg[5]/NET0131  & ~n44508 ;
  assign n61475 = ~n61473 & ~n61474 ;
  assign n61476 = \P2_P2_EBX_reg[6]/NET0131  & ~n44508 ;
  assign n61478 = n26662 & n46424 ;
  assign n61480 = \P2_P2_EBX_reg[6]/NET0131  & ~n61478 ;
  assign n61481 = ~n61437 & n61480 ;
  assign n61477 = \P2_P2_InstQueue_reg[0][6]/NET0131  & n46416 ;
  assign n61479 = ~\P2_P2_EBX_reg[6]/NET0131  & n61478 ;
  assign n61482 = ~n61477 & ~n61479 ;
  assign n61483 = ~n61481 & n61482 ;
  assign n61484 = n26792 & ~n61483 ;
  assign n61485 = ~n61476 & ~n61484 ;
  assign n61489 = \P2_P2_EBX_reg[7]/NET0131  & n61422 ;
  assign n61486 = ~\P2_P2_EBX_reg[7]/NET0131  & ~n46425 ;
  assign n61487 = ~n46426 & ~n61486 ;
  assign n61488 = n26662 & n61487 ;
  assign n61490 = ~\P2_P2_EBX_reg[7]/NET0131  & ~n26611 ;
  assign n61491 = ~\P2_P2_InstQueue_reg[0][7]/NET0131  & n26611 ;
  assign n61492 = ~n61490 & ~n61491 ;
  assign n61493 = n26578 & n61492 ;
  assign n61494 = ~n61488 & ~n61493 ;
  assign n61495 = ~n61489 & n61494 ;
  assign n61496 = n26792 & ~n61495 ;
  assign n61497 = \P2_P2_EBX_reg[7]/NET0131  & ~n44508 ;
  assign n61498 = ~n61496 & ~n61497 ;
  assign n61499 = \P1_P1_EAX_reg[1]/NET0131  & n24502 ;
  assign n61500 = ~n25050 & ~n61499 ;
  assign n61501 = ~n15364 & ~n61500 ;
  assign n61502 = \P1_P1_lWord_reg[1]/NET0131  & ~n24506 ;
  assign n61503 = ~n61501 & ~n61502 ;
  assign n61504 = n8355 & ~n61503 ;
  assign n61505 = \P1_P1_lWord_reg[1]/NET0131  & ~n24515 ;
  assign n61506 = ~n61504 & ~n61505 ;
  assign n61508 = \P1_P2_EBX_reg[1]/NET0131  & n48360 ;
  assign n61507 = n25803 & n50457 ;
  assign n61509 = ~\P1_P2_EBX_reg[1]/NET0131  & ~n25747 ;
  assign n61510 = ~\P1_P2_InstQueue_reg[0][1]/NET0131  & n25747 ;
  assign n61511 = ~n61509 & ~n61510 ;
  assign n61512 = n25738 & n61511 ;
  assign n61513 = ~n61507 & ~n61512 ;
  assign n61514 = ~n61508 & n61513 ;
  assign n61515 = n25918 & ~n61514 ;
  assign n61516 = \P1_P2_EBX_reg[1]/NET0131  & ~n43212 ;
  assign n61517 = ~n61515 & ~n61516 ;
  assign n61518 = n8355 & ~n46533 ;
  assign n61519 = n15326 & ~n61518 ;
  assign n61520 = \P1_P1_EBX_reg[0]/NET0131  & ~n61519 ;
  assign n61521 = \P1_P1_InstQueue_reg[0][0]/NET0131  & n46535 ;
  assign n61522 = ~\P1_P1_EBX_reg[0]/NET0131  & n26146 ;
  assign n61523 = ~n61521 & ~n61522 ;
  assign n61524 = n8355 & ~n61523 ;
  assign n61525 = ~n61520 & ~n61524 ;
  assign n61526 = n9241 & n46480 ;
  assign n61527 = n16968 & ~n61526 ;
  assign n61528 = \P1_P3_EBX_reg[0]/NET0131  & ~n61527 ;
  assign n61529 = ~\P1_P3_EBX_reg[0]/NET0131  & n9108 ;
  assign n61530 = \P1_P3_InstQueue_reg[0][0]/NET0131  & n46479 ;
  assign n61531 = ~n61529 & ~n61530 ;
  assign n61532 = n9241 & ~n61531 ;
  assign n61533 = ~n61528 & ~n61532 ;
  assign n61540 = \P1_P3_EBX_reg[1]/NET0131  & ~n9057 ;
  assign n61541 = ~n9108 & n61540 ;
  assign n61534 = ~\P1_P3_EBX_reg[1]/NET0131  & ~n9049 ;
  assign n61535 = ~\P1_P3_InstQueue_reg[0][1]/NET0131  & n9049 ;
  assign n61536 = ~n61534 & ~n61535 ;
  assign n61537 = n9057 & n61536 ;
  assign n61538 = ~n16501 & ~n19132 ;
  assign n61539 = n9108 & n61538 ;
  assign n61542 = ~n61537 & ~n61539 ;
  assign n61543 = ~n61541 & n61542 ;
  assign n61544 = n9241 & ~n61543 ;
  assign n61545 = \P1_P3_EBX_reg[1]/NET0131  & ~n16968 ;
  assign n61546 = ~n61544 & ~n61545 ;
  assign n61548 = \P1_P3_EBX_reg[2]/NET0131  & n46480 ;
  assign n61547 = \P1_P3_InstQueue_reg[0][2]/NET0131  & n46479 ;
  assign n61549 = ~\P1_P3_EBX_reg[2]/NET0131  & ~n19132 ;
  assign n61550 = ~n46483 & ~n61549 ;
  assign n61551 = n9108 & n61550 ;
  assign n61552 = ~n61547 & ~n61551 ;
  assign n61553 = ~n61548 & n61552 ;
  assign n61554 = n9241 & ~n61553 ;
  assign n61555 = \P1_P3_EBX_reg[2]/NET0131  & ~n16968 ;
  assign n61556 = ~n61554 & ~n61555 ;
  assign n61558 = \P1_P3_EBX_reg[3]/NET0131  & n46480 ;
  assign n61557 = \P1_P3_InstQueue_reg[0][3]/NET0131  & n46479 ;
  assign n61559 = ~\P1_P3_EBX_reg[3]/NET0131  & ~n46483 ;
  assign n61560 = ~n46484 & ~n61559 ;
  assign n61561 = n9108 & n61560 ;
  assign n61562 = ~n61557 & ~n61561 ;
  assign n61563 = ~n61558 & n61562 ;
  assign n61564 = n9241 & ~n61563 ;
  assign n61565 = \P1_P3_EBX_reg[3]/NET0131  & ~n16968 ;
  assign n61566 = ~n61564 & ~n61565 ;
  assign n61568 = \P1_P3_EBX_reg[5]/NET0131  & n46480 ;
  assign n61567 = \P1_P3_InstQueue_reg[0][5]/NET0131  & n46479 ;
  assign n61569 = ~\P1_P3_EBX_reg[5]/NET0131  & ~n46485 ;
  assign n61570 = ~n46486 & ~n61569 ;
  assign n61571 = n9108 & n61570 ;
  assign n61572 = ~n61567 & ~n61571 ;
  assign n61573 = ~n61568 & n61572 ;
  assign n61574 = n9241 & ~n61573 ;
  assign n61575 = \P1_P3_EBX_reg[5]/NET0131  & ~n16968 ;
  assign n61576 = ~n61574 & ~n61575 ;
  assign n61578 = \P1_P3_EBX_reg[4]/NET0131  & n46480 ;
  assign n61577 = \P1_P3_InstQueue_reg[0][4]/NET0131  & n46479 ;
  assign n61579 = ~\P1_P3_EBX_reg[4]/NET0131  & ~n46484 ;
  assign n61580 = ~n46485 & ~n61579 ;
  assign n61581 = n9108 & n61580 ;
  assign n61582 = ~n61577 & ~n61581 ;
  assign n61583 = ~n61578 & n61582 ;
  assign n61584 = n9241 & ~n61583 ;
  assign n61585 = \P1_P3_EBX_reg[4]/NET0131  & ~n16968 ;
  assign n61586 = ~n61584 & ~n61585 ;
  assign n61588 = \P1_P3_EBX_reg[6]/NET0131  & n46480 ;
  assign n61587 = \P1_P3_InstQueue_reg[0][6]/NET0131  & n46479 ;
  assign n61589 = ~\P1_P3_EBX_reg[6]/NET0131  & ~n46486 ;
  assign n61590 = ~n46487 & ~n61589 ;
  assign n61591 = n9108 & n61590 ;
  assign n61592 = ~n61587 & ~n61591 ;
  assign n61593 = ~n61588 & n61592 ;
  assign n61594 = n9241 & ~n61593 ;
  assign n61595 = \P1_P3_EBX_reg[6]/NET0131  & ~n16968 ;
  assign n61596 = ~n61594 & ~n61595 ;
  assign n61598 = \P1_P3_EBX_reg[7]/NET0131  & n46480 ;
  assign n61597 = \P1_P3_InstQueue_reg[0][7]/NET0131  & n46479 ;
  assign n61599 = ~\P1_P3_EBX_reg[7]/NET0131  & ~n46487 ;
  assign n61600 = ~n46488 & ~n61599 ;
  assign n61601 = n9108 & n61600 ;
  assign n61602 = ~n61597 & ~n61601 ;
  assign n61603 = ~n61598 & n61602 ;
  assign n61604 = n9241 & ~n61603 ;
  assign n61605 = \P1_P3_EBX_reg[7]/NET0131  & ~n16968 ;
  assign n61606 = ~n61604 & ~n61605 ;
  assign n61608 = \P1_P1_EBX_reg[1]/NET0131  & n46531 ;
  assign n61607 = n26146 & n50563 ;
  assign n61609 = ~\P1_P1_EBX_reg[1]/NET0131  & ~n15428 ;
  assign n61610 = ~\P1_P1_InstQueue_reg[0][1]/NET0131  & n15428 ;
  assign n61611 = ~n61609 & ~n61610 ;
  assign n61612 = n26122 & n61611 ;
  assign n61613 = ~n61607 & ~n61612 ;
  assign n61614 = ~n61608 & n61613 ;
  assign n61615 = n8355 & ~n61614 ;
  assign n61616 = \P1_P1_EBX_reg[1]/NET0131  & ~n15326 ;
  assign n61617 = ~n61615 & ~n61616 ;
  assign n61618 = \P1_P1_EBX_reg[2]/NET0131  & ~n15326 ;
  assign n61620 = n26146 & ~n46537 ;
  assign n61621 = n46533 & ~n61620 ;
  assign n61622 = \P1_P1_EBX_reg[2]/NET0131  & ~n61621 ;
  assign n61619 = \P1_P1_InstQueue_reg[0][2]/NET0131  & n46535 ;
  assign n61623 = ~\P1_P1_EBX_reg[2]/NET0131  & n46537 ;
  assign n61624 = n26146 & n61623 ;
  assign n61625 = ~n61619 & ~n61624 ;
  assign n61626 = ~n61622 & n61625 ;
  assign n61627 = n8355 & ~n61626 ;
  assign n61628 = ~n61618 & ~n61627 ;
  assign n61633 = \P1_P1_EBX_reg[3]/NET0131  & n46531 ;
  assign n61629 = ~\P1_P1_EBX_reg[3]/NET0131  & ~n15428 ;
  assign n61630 = ~\P1_P1_InstQueue_reg[0][3]/NET0131  & n15428 ;
  assign n61631 = ~n61629 & ~n61630 ;
  assign n61632 = n26122 & n61631 ;
  assign n61634 = ~\P1_P1_EBX_reg[3]/NET0131  & ~n46538 ;
  assign n61635 = n26146 & ~n46539 ;
  assign n61636 = ~n61634 & n61635 ;
  assign n61637 = ~n61632 & ~n61636 ;
  assign n61638 = ~n61633 & n61637 ;
  assign n61639 = n8355 & ~n61638 ;
  assign n61640 = \P1_P1_EBX_reg[3]/NET0131  & ~n15326 ;
  assign n61641 = ~n61639 & ~n61640 ;
  assign n61642 = \P1_P1_EBX_reg[4]/NET0131  & ~n15326 ;
  assign n61644 = n46533 & ~n61635 ;
  assign n61645 = \P1_P1_EBX_reg[4]/NET0131  & ~n61644 ;
  assign n61643 = \P1_P1_InstQueue_reg[0][4]/NET0131  & n46535 ;
  assign n61646 = ~\P1_P1_EBX_reg[4]/NET0131  & n46539 ;
  assign n61647 = n26146 & n61646 ;
  assign n61648 = ~n61643 & ~n61647 ;
  assign n61649 = ~n61645 & n61648 ;
  assign n61650 = n8355 & ~n61649 ;
  assign n61651 = ~n61642 & ~n61650 ;
  assign n61656 = \P1_P1_EBX_reg[5]/NET0131  & n46531 ;
  assign n61652 = ~\P1_P1_EBX_reg[5]/NET0131  & ~n15428 ;
  assign n61653 = ~\P1_P1_InstQueue_reg[0][5]/NET0131  & n15428 ;
  assign n61654 = ~n61652 & ~n61653 ;
  assign n61655 = n26122 & n61654 ;
  assign n61657 = ~\P1_P1_EBX_reg[5]/NET0131  & ~n46540 ;
  assign n61658 = n26146 & ~n46541 ;
  assign n61659 = ~n61657 & n61658 ;
  assign n61660 = ~n61655 & ~n61659 ;
  assign n61661 = ~n61656 & n61660 ;
  assign n61662 = n8355 & ~n61661 ;
  assign n61663 = \P1_P1_EBX_reg[5]/NET0131  & ~n15326 ;
  assign n61664 = ~n61662 & ~n61663 ;
  assign n61665 = \P1_P1_EBX_reg[6]/NET0131  & ~n15326 ;
  assign n61667 = n46533 & ~n61658 ;
  assign n61668 = \P1_P1_EBX_reg[6]/NET0131  & ~n61667 ;
  assign n61666 = \P1_P1_InstQueue_reg[0][6]/NET0131  & n46535 ;
  assign n61669 = ~\P1_P1_EBX_reg[6]/NET0131  & n46541 ;
  assign n61670 = n26146 & n61669 ;
  assign n61671 = ~n61666 & ~n61670 ;
  assign n61672 = ~n61668 & n61671 ;
  assign n61673 = n8355 & ~n61672 ;
  assign n61674 = ~n61665 & ~n61673 ;
  assign n61678 = \P1_P1_EBX_reg[7]/NET0131  & n46531 ;
  assign n61675 = ~\P1_P1_EBX_reg[7]/NET0131  & ~n46542 ;
  assign n61676 = ~n46543 & ~n61675 ;
  assign n61677 = n26146 & n61676 ;
  assign n61679 = ~\P1_P1_EBX_reg[7]/NET0131  & ~n15428 ;
  assign n61680 = ~\P1_P1_InstQueue_reg[0][7]/NET0131  & n15428 ;
  assign n61681 = ~n61679 & ~n61680 ;
  assign n61682 = n26122 & n61681 ;
  assign n61683 = ~n61677 & ~n61682 ;
  assign n61684 = ~n61678 & n61683 ;
  assign n61685 = n8355 & ~n61684 ;
  assign n61686 = \P1_P1_EBX_reg[7]/NET0131  & ~n15326 ;
  assign n61687 = ~n61685 & ~n61686 ;
  assign n61689 = \P1_P2_EBX_reg[3]/NET0131  & n46695 ;
  assign n61688 = \P1_P2_InstQueue_reg[0][3]/NET0131  & n46694 ;
  assign n61690 = ~\P1_P2_EBX_reg[3]/NET0131  & ~n46699 ;
  assign n61691 = n25803 & ~n46700 ;
  assign n61692 = ~n61690 & n61691 ;
  assign n61693 = ~n61688 & ~n61692 ;
  assign n61694 = ~n61689 & n61693 ;
  assign n61695 = n25918 & ~n61694 ;
  assign n61696 = \P1_P2_EBX_reg[3]/NET0131  & ~n43212 ;
  assign n61697 = ~n61695 & ~n61696 ;
  assign n61698 = n27308 & n46615 ;
  assign n61699 = n42872 & ~n61698 ;
  assign n61700 = \P2_P3_EBX_reg[0]/NET0131  & ~n61699 ;
  assign n61701 = ~\P2_P3_EBX_reg[0]/NET0131  & n27133 ;
  assign n61702 = \P2_P3_InstQueue_reg[0][0]/NET0131  & n46614 ;
  assign n61703 = ~n61701 & ~n61702 ;
  assign n61704 = n27308 & ~n61703 ;
  assign n61705 = ~n61700 & ~n61704 ;
  assign n61712 = \P2_P3_EBX_reg[1]/NET0131  & ~n27108 ;
  assign n61713 = ~n27133 & n61712 ;
  assign n61706 = ~\P2_P3_EBX_reg[1]/NET0131  & ~n27206 ;
  assign n61707 = ~\P2_P3_InstQueue_reg[0][1]/NET0131  & n27206 ;
  assign n61708 = ~n61706 & ~n61707 ;
  assign n61709 = n27108 & n61708 ;
  assign n61710 = ~n46618 & ~n50720 ;
  assign n61711 = n27133 & n61710 ;
  assign n61714 = ~n61709 & ~n61711 ;
  assign n61715 = ~n61713 & n61714 ;
  assign n61716 = n27308 & ~n61715 ;
  assign n61717 = \P2_P3_EBX_reg[1]/NET0131  & ~n42872 ;
  assign n61718 = ~n61716 & ~n61717 ;
  assign n61720 = \P2_P3_EBX_reg[2]/NET0131  & n46615 ;
  assign n61719 = \P2_P3_InstQueue_reg[0][2]/NET0131  & n46614 ;
  assign n61721 = ~\P2_P3_EBX_reg[2]/NET0131  & ~n46618 ;
  assign n61722 = n27133 & ~n46619 ;
  assign n61723 = ~n61721 & n61722 ;
  assign n61724 = ~n61719 & ~n61723 ;
  assign n61725 = ~n61720 & n61724 ;
  assign n61726 = n27308 & ~n61725 ;
  assign n61727 = \P2_P3_EBX_reg[2]/NET0131  & ~n42872 ;
  assign n61728 = ~n61726 & ~n61727 ;
  assign n61729 = \P2_P3_EBX_reg[3]/NET0131  & ~n42872 ;
  assign n61731 = ~n46615 & ~n61722 ;
  assign n61732 = \P2_P3_EBX_reg[3]/NET0131  & ~n61731 ;
  assign n61730 = \P2_P3_InstQueue_reg[0][3]/NET0131  & n46614 ;
  assign n61733 = ~\P2_P3_EBX_reg[3]/NET0131  & n46619 ;
  assign n61734 = n27133 & n61733 ;
  assign n61735 = ~n61730 & ~n61734 ;
  assign n61736 = ~n61732 & n61735 ;
  assign n61737 = n27308 & ~n61736 ;
  assign n61738 = ~n61729 & ~n61737 ;
  assign n61740 = \P2_P3_EBX_reg[4]/NET0131  & n46615 ;
  assign n61739 = \P2_P3_InstQueue_reg[0][4]/NET0131  & n46614 ;
  assign n61741 = ~\P2_P3_EBX_reg[4]/NET0131  & ~n46620 ;
  assign n61742 = n27133 & ~n46621 ;
  assign n61743 = ~n61741 & n61742 ;
  assign n61744 = ~n61739 & ~n61743 ;
  assign n61745 = ~n61740 & n61744 ;
  assign n61746 = n27308 & ~n61745 ;
  assign n61747 = \P2_P3_EBX_reg[4]/NET0131  & ~n42872 ;
  assign n61748 = ~n61746 & ~n61747 ;
  assign n61749 = \P2_P3_EBX_reg[5]/NET0131  & ~n42872 ;
  assign n61751 = ~n46615 & ~n61742 ;
  assign n61752 = \P2_P3_EBX_reg[5]/NET0131  & ~n61751 ;
  assign n61750 = \P2_P3_InstQueue_reg[0][5]/NET0131  & n46614 ;
  assign n61753 = ~\P2_P3_EBX_reg[5]/NET0131  & n46621 ;
  assign n61754 = n27133 & n61753 ;
  assign n61755 = ~n61750 & ~n61754 ;
  assign n61756 = ~n61752 & n61755 ;
  assign n61757 = n27308 & ~n61756 ;
  assign n61758 = ~n61749 & ~n61757 ;
  assign n61760 = \P2_P3_EBX_reg[6]/NET0131  & n46615 ;
  assign n61759 = \P2_P3_InstQueue_reg[0][6]/NET0131  & n46614 ;
  assign n61761 = ~\P2_P3_EBX_reg[6]/NET0131  & ~n46622 ;
  assign n61762 = n27133 & ~n46623 ;
  assign n61763 = ~n61761 & n61762 ;
  assign n61764 = ~n61759 & ~n61763 ;
  assign n61765 = ~n61760 & n61764 ;
  assign n61766 = n27308 & ~n61765 ;
  assign n61767 = \P2_P3_EBX_reg[6]/NET0131  & ~n42872 ;
  assign n61768 = ~n61766 & ~n61767 ;
  assign n61769 = \P2_P3_EBX_reg[7]/NET0131  & ~n42872 ;
  assign n61771 = ~n46615 & ~n61762 ;
  assign n61772 = \P2_P3_EBX_reg[7]/NET0131  & ~n61771 ;
  assign n61770 = \P2_P3_InstQueue_reg[0][7]/NET0131  & n46614 ;
  assign n61773 = ~\P2_P3_EBX_reg[7]/NET0131  & n46623 ;
  assign n61774 = n27133 & n61773 ;
  assign n61775 = ~n61770 & ~n61774 ;
  assign n61776 = ~n61772 & n61775 ;
  assign n61777 = n27308 & ~n61776 ;
  assign n61778 = ~n61769 & ~n61777 ;
  assign n61779 = n25918 & n46695 ;
  assign n61780 = n43212 & ~n61779 ;
  assign n61781 = \P1_P2_EBX_reg[0]/NET0131  & ~n61780 ;
  assign n61782 = ~\P1_P2_EBX_reg[0]/NET0131  & n25803 ;
  assign n61783 = \P1_P2_InstQueue_reg[0][0]/NET0131  & n46694 ;
  assign n61784 = ~n61782 & ~n61783 ;
  assign n61785 = n25918 & ~n61784 ;
  assign n61786 = ~n61781 & ~n61785 ;
  assign n61788 = \P1_P2_EBX_reg[2]/NET0131  & n46695 ;
  assign n61787 = \P1_P2_InstQueue_reg[0][2]/NET0131  & n46694 ;
  assign n61789 = ~\P1_P2_EBX_reg[2]/NET0131  & ~n46698 ;
  assign n61790 = ~n46699 & ~n61789 ;
  assign n61791 = n25803 & n61790 ;
  assign n61792 = ~n61787 & ~n61791 ;
  assign n61793 = ~n61788 & n61792 ;
  assign n61794 = n25918 & ~n61793 ;
  assign n61795 = \P1_P2_EBX_reg[2]/NET0131  & ~n43212 ;
  assign n61796 = ~n61794 & ~n61795 ;
  assign n61797 = \P1_P2_EBX_reg[4]/NET0131  & ~n43212 ;
  assign n61799 = ~n46695 & ~n61691 ;
  assign n61800 = \P1_P2_EBX_reg[4]/NET0131  & ~n61799 ;
  assign n61798 = \P1_P2_InstQueue_reg[0][4]/NET0131  & n46694 ;
  assign n61801 = ~\P1_P2_EBX_reg[4]/NET0131  & n46700 ;
  assign n61802 = n25803 & n61801 ;
  assign n61803 = ~n61798 & ~n61802 ;
  assign n61804 = ~n61800 & n61803 ;
  assign n61805 = n25918 & ~n61804 ;
  assign n61806 = ~n61797 & ~n61805 ;
  assign n61807 = \P1_P2_EBX_reg[6]/NET0131  & ~n43212 ;
  assign n61809 = ~n46695 & ~n61299 ;
  assign n61810 = \P1_P2_EBX_reg[6]/NET0131  & ~n61809 ;
  assign n61808 = \P1_P2_InstQueue_reg[0][6]/NET0131  & n46694 ;
  assign n61811 = ~\P1_P2_EBX_reg[6]/NET0131  & n46702 ;
  assign n61812 = n25803 & n61811 ;
  assign n61813 = ~n61808 & ~n61812 ;
  assign n61814 = ~n61810 & n61813 ;
  assign n61815 = n25918 & ~n61814 ;
  assign n61816 = ~n61807 & ~n61815 ;
  assign n61820 = \P1_P2_EBX_reg[7]/NET0131  & n48360 ;
  assign n61817 = ~\P1_P2_EBX_reg[7]/NET0131  & ~n46703 ;
  assign n61818 = ~n46704 & ~n61817 ;
  assign n61819 = n25803 & n61818 ;
  assign n61821 = ~\P1_P2_EBX_reg[7]/NET0131  & ~n25747 ;
  assign n61822 = ~\P1_P2_InstQueue_reg[0][7]/NET0131  & n25747 ;
  assign n61823 = ~n61821 & ~n61822 ;
  assign n61824 = n25738 & n61823 ;
  assign n61825 = ~n61819 & ~n61824 ;
  assign n61826 = ~n61820 & n61825 ;
  assign n61827 = n25918 & ~n61826 ;
  assign n61828 = \P1_P2_EBX_reg[7]/NET0131  & ~n43212 ;
  assign n61829 = ~n61827 & ~n61828 ;
  assign n61831 = \P1_P1_Datao_reg[16]/NET0131  & ~n26162 ;
  assign n61832 = n26175 & n60438 ;
  assign n61833 = ~n61831 & ~n61832 ;
  assign n61834 = n8355 & ~n61833 ;
  assign n61830 = \P1_P1_uWord_reg[0]/NET0131  & n27790 ;
  assign n61835 = \P1_P1_Datao_reg[16]/NET0131  & ~n48479 ;
  assign n61836 = ~n61830 & ~n61835 ;
  assign n61837 = ~n61834 & n61836 ;
  assign n61839 = ~n26158 & n60467 ;
  assign n61840 = \P1_P1_Datao_reg[18]/NET0131  & ~n26162 ;
  assign n61841 = ~n61839 & ~n61840 ;
  assign n61842 = n8355 & ~n61841 ;
  assign n61838 = \P1_P1_uWord_reg[2]/NET0131  & n27790 ;
  assign n61843 = \P1_P1_Datao_reg[18]/NET0131  & ~n48479 ;
  assign n61844 = ~n61838 & ~n61843 ;
  assign n61845 = ~n61842 & n61844 ;
  assign n61847 = n8355 & ~n26162 ;
  assign n61848 = n48479 & ~n61847 ;
  assign n61849 = \P1_P1_Datao_reg[21]/NET0131  & ~n61848 ;
  assign n61846 = \P1_P1_uWord_reg[5]/NET0131  & n27790 ;
  assign n61850 = n8355 & ~n26158 ;
  assign n61851 = n44768 & n61850 ;
  assign n61852 = ~n61846 & ~n61851 ;
  assign n61853 = ~n61849 & n61852 ;
  assign n61855 = ~n26158 & n44780 ;
  assign n61856 = \P1_P1_Datao_reg[22]/NET0131  & ~n26162 ;
  assign n61857 = ~n61855 & ~n61856 ;
  assign n61858 = n8355 & ~n61857 ;
  assign n61854 = \P1_P1_uWord_reg[6]/NET0131  & n27790 ;
  assign n61859 = \P1_P1_Datao_reg[22]/NET0131  & ~n48479 ;
  assign n61860 = ~n61854 & ~n61859 ;
  assign n61861 = ~n61858 & n61860 ;
  assign n61863 = ~n26158 & ~n34441 ;
  assign n61864 = n24503 & ~n61863 ;
  assign n61865 = n53011 & ~n61864 ;
  assign n61866 = \P1_P1_Datao_reg[25]/NET0131  & ~n61865 ;
  assign n61867 = ~n26158 & n34442 ;
  assign n61868 = ~n61866 & ~n61867 ;
  assign n61869 = n8355 & ~n61868 ;
  assign n61862 = \P1_P1_uWord_reg[9]/NET0131  & n27790 ;
  assign n61870 = \P1_P1_Datao_reg[25]/NET0131  & ~n48479 ;
  assign n61871 = ~n61862 & ~n61870 ;
  assign n61872 = ~n61869 & n61871 ;
  assign n61874 = \P1_P1_Datao_reg[26]/NET0131  & ~n26162 ;
  assign n61875 = ~n26158 & n34181 ;
  assign n61876 = ~n61874 & ~n61875 ;
  assign n61877 = n8355 & ~n61876 ;
  assign n61873 = \P1_P1_uWord_reg[10]/NET0131  & n27790 ;
  assign n61878 = \P1_P1_Datao_reg[26]/NET0131  & ~n48479 ;
  assign n61879 = ~n61873 & ~n61878 ;
  assign n61880 = ~n61877 & n61879 ;
  assign n61882 = ~n26158 & ~n27431 ;
  assign n61883 = n24503 & ~n61882 ;
  assign n61884 = n53011 & ~n61883 ;
  assign n61885 = \P1_P1_Datao_reg[29]/NET0131  & ~n61884 ;
  assign n61886 = ~n26158 & n27432 ;
  assign n61887 = ~n61885 & ~n61886 ;
  assign n61888 = n8355 & ~n61887 ;
  assign n61881 = \P1_P1_uWord_reg[13]/NET0131  & n27790 ;
  assign n61889 = \P1_P1_Datao_reg[29]/NET0131  & ~n48479 ;
  assign n61890 = ~n61881 & ~n61889 ;
  assign n61891 = ~n61888 & n61890 ;
  assign n61893 = ~n26158 & n60458 ;
  assign n61894 = \P1_P1_Datao_reg[17]/NET0131  & ~n26162 ;
  assign n61895 = ~n61893 & ~n61894 ;
  assign n61896 = n8355 & ~n61895 ;
  assign n61892 = \P1_P1_uWord_reg[1]/NET0131  & n27790 ;
  assign n61897 = \P1_P1_Datao_reg[17]/NET0131  & ~n48479 ;
  assign n61898 = ~n61892 & ~n61897 ;
  assign n61899 = ~n61896 & n61898 ;
  assign n61901 = \P2_P2_Datao_reg[16]/NET0131  & ~n26699 ;
  assign n61902 = ~n26650 & n60494 ;
  assign n61903 = ~n61901 & ~n61902 ;
  assign n61904 = n26792 & ~n61903 ;
  assign n61900 = \P2_P2_uWord_reg[0]/NET0131  & n48491 ;
  assign n61905 = \P2_P2_Datao_reg[16]/NET0131  & ~n48508 ;
  assign n61906 = ~n61900 & ~n61905 ;
  assign n61907 = ~n61904 & n61906 ;
  assign n61909 = ~n26650 & n60542 ;
  assign n61910 = \P2_P2_Datao_reg[17]/NET0131  & ~n26699 ;
  assign n61911 = ~n61909 & ~n61910 ;
  assign n61912 = n26792 & ~n61911 ;
  assign n61908 = \P2_P2_uWord_reg[1]/NET0131  & n48491 ;
  assign n61913 = \P2_P2_Datao_reg[17]/NET0131  & ~n48508 ;
  assign n61914 = ~n61908 & ~n61913 ;
  assign n61915 = ~n61912 & n61914 ;
  assign n61917 = ~n26650 & ~n60552 ;
  assign n61918 = n26786 & ~n61917 ;
  assign n61919 = n48494 & ~n61918 ;
  assign n61920 = \P2_P2_Datao_reg[18]/NET0131  & ~n61919 ;
  assign n61921 = n26692 & n60553 ;
  assign n61922 = ~n61920 & ~n61921 ;
  assign n61923 = n26792 & ~n61922 ;
  assign n61916 = \P2_P2_uWord_reg[2]/NET0131  & n48491 ;
  assign n61924 = \P2_P2_Datao_reg[18]/NET0131  & ~n48508 ;
  assign n61925 = ~n61916 & ~n61924 ;
  assign n61926 = ~n61923 & n61925 ;
  assign n61928 = \P2_P2_Datao_reg[21]/NET0131  & ~n26699 ;
  assign n61929 = ~n26650 & n60571 ;
  assign n61930 = ~n61928 & ~n61929 ;
  assign n61931 = n26792 & ~n61930 ;
  assign n61927 = \P2_P2_uWord_reg[5]/NET0131  & n48491 ;
  assign n61932 = \P2_P2_Datao_reg[21]/NET0131  & ~n48508 ;
  assign n61933 = ~n61927 & ~n61932 ;
  assign n61934 = ~n61931 & n61933 ;
  assign n61936 = \P2_P2_Datao_reg[22]/NET0131  & ~n26699 ;
  assign n61937 = ~n26650 & n60586 ;
  assign n61938 = ~n61936 & ~n61937 ;
  assign n61939 = n26792 & ~n61938 ;
  assign n61935 = \P2_P2_uWord_reg[6]/NET0131  & n48491 ;
  assign n61940 = \P2_P2_Datao_reg[22]/NET0131  & ~n48508 ;
  assign n61941 = ~n61935 & ~n61940 ;
  assign n61942 = ~n61939 & n61941 ;
  assign n61944 = ~n26650 & ~n60601 ;
  assign n61945 = n26786 & ~n61944 ;
  assign n61946 = n48494 & ~n61945 ;
  assign n61947 = \P2_P2_Datao_reg[25]/NET0131  & ~n61946 ;
  assign n61948 = n26692 & n60602 ;
  assign n61949 = ~n61947 & ~n61948 ;
  assign n61950 = n26792 & ~n61949 ;
  assign n61943 = \P2_P2_uWord_reg[9]/NET0131  & n48491 ;
  assign n61951 = \P2_P2_Datao_reg[25]/NET0131  & ~n48508 ;
  assign n61952 = ~n61943 & ~n61951 ;
  assign n61953 = ~n61950 & n61952 ;
  assign n61955 = ~n26650 & ~n60505 ;
  assign n61956 = n26786 & ~n61955 ;
  assign n61957 = n48494 & ~n61956 ;
  assign n61958 = \P2_P2_Datao_reg[26]/NET0131  & ~n61957 ;
  assign n61959 = n26692 & n60506 ;
  assign n61960 = ~n61958 & ~n61959 ;
  assign n61961 = n26792 & ~n61960 ;
  assign n61954 = \P2_P2_uWord_reg[10]/NET0131  & n48491 ;
  assign n61962 = \P2_P2_Datao_reg[26]/NET0131  & ~n48508 ;
  assign n61963 = ~n61954 & ~n61962 ;
  assign n61964 = ~n61961 & n61963 ;
  assign n61966 = \P2_P2_Datao_reg[29]/NET0131  & ~n26699 ;
  assign n61967 = n26692 & n60527 ;
  assign n61968 = ~n61966 & ~n61967 ;
  assign n61969 = n26792 & ~n61968 ;
  assign n61965 = \P2_P2_uWord_reg[13]/NET0131  & n48491 ;
  assign n61970 = \P2_P2_Datao_reg[29]/NET0131  & ~n48508 ;
  assign n61971 = ~n61965 & ~n61970 ;
  assign n61972 = ~n61969 & n61971 ;
  assign n61974 = \P2_P3_Datao_reg[16]/NET0131  & ~n27223 ;
  assign n61975 = ~n27148 & n60792 ;
  assign n61976 = ~n61974 & ~n61975 ;
  assign n61977 = n27308 & ~n61976 ;
  assign n61973 = \P2_P3_uWord_reg[0]/NET0131  & n48523 ;
  assign n61978 = \P2_P3_Datao_reg[16]/NET0131  & ~n48540 ;
  assign n61979 = ~n61973 & ~n61978 ;
  assign n61980 = ~n61977 & n61979 ;
  assign n61982 = \P2_P3_Datao_reg[17]/NET0131  & ~n27223 ;
  assign n61983 = ~n27148 & n60830 ;
  assign n61984 = ~n61982 & ~n61983 ;
  assign n61985 = n27308 & ~n61984 ;
  assign n61981 = \P2_P3_uWord_reg[1]/NET0131  & n48523 ;
  assign n61986 = \P2_P3_Datao_reg[17]/NET0131  & ~n48540 ;
  assign n61987 = ~n61981 & ~n61986 ;
  assign n61988 = ~n61985 & n61987 ;
  assign n61990 = \P2_P3_Datao_reg[18]/NET0131  & ~n27223 ;
  assign n61991 = ~n27148 & n60843 ;
  assign n61992 = ~n61990 & ~n61991 ;
  assign n61993 = n27308 & ~n61992 ;
  assign n61989 = \P2_P3_uWord_reg[2]/NET0131  & n48523 ;
  assign n61994 = \P2_P3_Datao_reg[18]/NET0131  & ~n48540 ;
  assign n61995 = ~n61989 & ~n61994 ;
  assign n61996 = ~n61993 & n61995 ;
  assign n61998 = \P2_P3_Datao_reg[21]/NET0131  & ~n27223 ;
  assign n61999 = n27303 & n60861 ;
  assign n62000 = ~n61998 & ~n61999 ;
  assign n62001 = n27308 & ~n62000 ;
  assign n61997 = \P2_P3_uWord_reg[5]/NET0131  & n48523 ;
  assign n62002 = \P2_P3_Datao_reg[21]/NET0131  & ~n48540 ;
  assign n62003 = ~n61997 & ~n62002 ;
  assign n62004 = ~n62001 & n62003 ;
  assign n62006 = \P2_P3_Datao_reg[22]/NET0131  & ~n56850 ;
  assign n62005 = \P2_P3_uWord_reg[6]/NET0131  & n48523 ;
  assign n62007 = ~n27177 & n56841 ;
  assign n62008 = n60871 & n62007 ;
  assign n62009 = ~n62005 & ~n62008 ;
  assign n62010 = ~n62006 & n62009 ;
  assign n62012 = \P2_P3_Datao_reg[25]/NET0131  & ~n56850 ;
  assign n62011 = \P2_P3_uWord_reg[9]/NET0131  & n48523 ;
  assign n62013 = n56841 & n60888 ;
  assign n62014 = ~n62011 & ~n62013 ;
  assign n62015 = ~n62012 & n62014 ;
  assign n62017 = \P2_P3_Datao_reg[26]/NET0131  & ~n27223 ;
  assign n62018 = n27303 & n60801 ;
  assign n62019 = ~n62017 & ~n62018 ;
  assign n62020 = n27308 & ~n62019 ;
  assign n62016 = \P2_P3_uWord_reg[10]/NET0131  & n48523 ;
  assign n62021 = \P2_P3_Datao_reg[26]/NET0131  & ~n48540 ;
  assign n62022 = ~n62016 & ~n62021 ;
  assign n62023 = ~n62020 & n62022 ;
  assign n62025 = \P2_P3_Datao_reg[29]/NET0131  & ~n27223 ;
  assign n62026 = ~n27148 & n60812 ;
  assign n62027 = ~n62025 & ~n62026 ;
  assign n62028 = n27308 & ~n62027 ;
  assign n62024 = \P2_P3_uWord_reg[13]/NET0131  & n48523 ;
  assign n62029 = \P2_P3_Datao_reg[29]/NET0131  & ~n48540 ;
  assign n62030 = ~n62024 & ~n62029 ;
  assign n62031 = ~n62028 & n62030 ;
  assign n62033 = ~n25768 & ~n59830 ;
  assign n62034 = n47570 & ~n62033 ;
  assign n62035 = n48554 & ~n62034 ;
  assign n62036 = \P1_P2_Datao_reg[16]/NET0131  & ~n62035 ;
  assign n62037 = ~n25768 & n59831 ;
  assign n62038 = ~n62036 & ~n62037 ;
  assign n62039 = n25918 & ~n62038 ;
  assign n62032 = \P1_P2_uWord_reg[0]/NET0131  & n25922 ;
  assign n62040 = \P1_P2_Datao_reg[16]/NET0131  & ~n48566 ;
  assign n62041 = ~n62032 & ~n62040 ;
  assign n62042 = ~n62039 & n62041 ;
  assign n62044 = ~n25768 & n59869 ;
  assign n62045 = \P1_P2_Datao_reg[17]/NET0131  & ~n25847 ;
  assign n62046 = ~n62044 & ~n62045 ;
  assign n62047 = n25918 & ~n62046 ;
  assign n62043 = \P1_P2_uWord_reg[1]/NET0131  & n25922 ;
  assign n62048 = \P1_P2_Datao_reg[17]/NET0131  & ~n48566 ;
  assign n62049 = ~n62043 & ~n62048 ;
  assign n62050 = ~n62047 & n62049 ;
  assign n62052 = ~n25768 & n59878 ;
  assign n62053 = \P1_P2_Datao_reg[18]/NET0131  & ~n25847 ;
  assign n62054 = ~n62052 & ~n62053 ;
  assign n62055 = n25918 & ~n62054 ;
  assign n62051 = \P1_P2_uWord_reg[2]/NET0131  & n25922 ;
  assign n62056 = \P1_P2_Datao_reg[18]/NET0131  & ~n48566 ;
  assign n62057 = ~n62051 & ~n62056 ;
  assign n62058 = ~n62055 & n62057 ;
  assign n62060 = ~n25768 & n59899 ;
  assign n62061 = \P1_P2_Datao_reg[21]/NET0131  & ~n25847 ;
  assign n62062 = ~n62060 & ~n62061 ;
  assign n62063 = n25918 & ~n62062 ;
  assign n62059 = \P1_P2_uWord_reg[5]/NET0131  & n25922 ;
  assign n62064 = \P1_P2_Datao_reg[21]/NET0131  & ~n48566 ;
  assign n62065 = ~n62059 & ~n62064 ;
  assign n62066 = ~n62063 & n62065 ;
  assign n62068 = ~n25768 & ~n59906 ;
  assign n62069 = n47570 & ~n62068 ;
  assign n62070 = n48554 & ~n62069 ;
  assign n62071 = \P1_P2_Datao_reg[22]/NET0131  & ~n62070 ;
  assign n62072 = ~n25768 & n59907 ;
  assign n62073 = ~n62071 & ~n62072 ;
  assign n62074 = n25918 & ~n62073 ;
  assign n62067 = \P1_P2_uWord_reg[6]/NET0131  & n25922 ;
  assign n62075 = \P1_P2_Datao_reg[22]/NET0131  & ~n48566 ;
  assign n62076 = ~n62067 & ~n62075 ;
  assign n62077 = ~n62074 & n62076 ;
  assign n62079 = ~n25768 & ~n59921 ;
  assign n62080 = n47570 & ~n62079 ;
  assign n62081 = n48554 & ~n62080 ;
  assign n62082 = \P1_P2_Datao_reg[25]/NET0131  & ~n62081 ;
  assign n62083 = ~n25768 & n59922 ;
  assign n62084 = ~n62082 & ~n62083 ;
  assign n62085 = n25918 & ~n62084 ;
  assign n62078 = \P1_P2_uWord_reg[9]/NET0131  & n25922 ;
  assign n62086 = \P1_P2_Datao_reg[25]/NET0131  & ~n48566 ;
  assign n62087 = ~n62078 & ~n62086 ;
  assign n62088 = ~n62085 & n62087 ;
  assign n62093 = n25841 & n25918 ;
  assign n62094 = n59840 & n62093 ;
  assign n62089 = ~n25847 & n25918 ;
  assign n62090 = n48566 & ~n62089 ;
  assign n62091 = \P1_P2_Datao_reg[26]/NET0131  & ~n62090 ;
  assign n62092 = \P1_P2_uWord_reg[10]/NET0131  & n25922 ;
  assign n62095 = ~n62091 & ~n62092 ;
  assign n62096 = ~n62094 & n62095 ;
  assign n62098 = ~n25768 & n59848 ;
  assign n62099 = \P1_P2_Datao_reg[29]/NET0131  & ~n25847 ;
  assign n62100 = ~n62098 & ~n62099 ;
  assign n62101 = n25918 & ~n62100 ;
  assign n62097 = \P1_P2_uWord_reg[13]/NET0131  & n25922 ;
  assign n62102 = \P1_P2_Datao_reg[29]/NET0131  & ~n48566 ;
  assign n62103 = ~n62097 & ~n62102 ;
  assign n62104 = ~n62101 & n62103 ;
  assign n62106 = ~n25958 & ~n44492 ;
  assign n62107 = n24899 & ~n62106 ;
  assign n62108 = n48584 & ~n62107 ;
  assign n62109 = \P2_P1_Datao_reg[21]/NET0131  & ~n62108 ;
  assign n62110 = ~n25958 & n44493 ;
  assign n62111 = ~n62109 & ~n62110 ;
  assign n62112 = n11623 & ~n62111 ;
  assign n62105 = \P2_P1_uWord_reg[5]/NET0131  & n48581 ;
  assign n62113 = \P2_P1_Datao_reg[21]/NET0131  & ~n48594 ;
  assign n62114 = ~n62105 & ~n62113 ;
  assign n62115 = ~n62112 & n62114 ;
  assign n62117 = ~n25958 & ~n59804 ;
  assign n62118 = n24899 & ~n62117 ;
  assign n62119 = n48584 & ~n62118 ;
  assign n62120 = \P2_P1_Datao_reg[16]/NET0131  & ~n62119 ;
  assign n62121 = ~n25958 & n59805 ;
  assign n62122 = ~n62120 & ~n62121 ;
  assign n62123 = n11623 & ~n62122 ;
  assign n62116 = \P2_P1_uWord_reg[0]/NET0131  & n48581 ;
  assign n62124 = \P2_P1_Datao_reg[16]/NET0131  & ~n48594 ;
  assign n62125 = ~n62116 & ~n62124 ;
  assign n62126 = ~n62123 & n62125 ;
  assign n62128 = ~n25958 & ~n59812 ;
  assign n62129 = n24899 & ~n62128 ;
  assign n62130 = n48584 & ~n62129 ;
  assign n62131 = \P2_P1_Datao_reg[17]/NET0131  & ~n62130 ;
  assign n62132 = ~n25958 & n59813 ;
  assign n62133 = ~n62131 & ~n62132 ;
  assign n62134 = n11623 & ~n62133 ;
  assign n62127 = \P2_P1_uWord_reg[1]/NET0131  & n48581 ;
  assign n62135 = \P2_P1_Datao_reg[17]/NET0131  & ~n48594 ;
  assign n62136 = ~n62127 & ~n62135 ;
  assign n62137 = ~n62134 & n62136 ;
  assign n62139 = ~n25958 & ~n59822 ;
  assign n62140 = n24899 & ~n62139 ;
  assign n62141 = n48584 & ~n62140 ;
  assign n62142 = \P2_P1_Datao_reg[18]/NET0131  & ~n62141 ;
  assign n62143 = ~n25958 & n59823 ;
  assign n62144 = ~n62142 & ~n62143 ;
  assign n62145 = n11623 & ~n62144 ;
  assign n62138 = \P2_P1_uWord_reg[2]/NET0131  & n48581 ;
  assign n62146 = \P2_P1_Datao_reg[18]/NET0131  & ~n48594 ;
  assign n62147 = ~n62138 & ~n62146 ;
  assign n62148 = ~n62145 & n62147 ;
  assign n62150 = ~n25958 & ~n44501 ;
  assign n62151 = n24899 & ~n62150 ;
  assign n62152 = n48584 & ~n62151 ;
  assign n62153 = \P2_P1_Datao_reg[22]/NET0131  & ~n62152 ;
  assign n62154 = ~n25958 & n44502 ;
  assign n62155 = ~n62153 & ~n62154 ;
  assign n62156 = n11623 & ~n62155 ;
  assign n62149 = \P2_P1_uWord_reg[6]/NET0131  & n48581 ;
  assign n62157 = \P2_P1_Datao_reg[22]/NET0131  & ~n48594 ;
  assign n62158 = ~n62149 & ~n62157 ;
  assign n62159 = ~n62156 & n62158 ;
  assign n62161 = ~n25958 & n34419 ;
  assign n62162 = \P2_P1_Datao_reg[25]/NET0131  & ~n26030 ;
  assign n62163 = ~n62161 & ~n62162 ;
  assign n62164 = n11623 & ~n62163 ;
  assign n62160 = \P2_P1_uWord_reg[9]/NET0131  & n48581 ;
  assign n62165 = \P2_P1_Datao_reg[25]/NET0131  & ~n48594 ;
  assign n62166 = ~n62160 & ~n62165 ;
  assign n62167 = ~n62164 & n62166 ;
  assign n62169 = ~n25958 & ~n34171 ;
  assign n62170 = n24899 & ~n62169 ;
  assign n62171 = n48584 & ~n62170 ;
  assign n62172 = \P2_P1_Datao_reg[26]/NET0131  & ~n62171 ;
  assign n62173 = n26006 & n34172 ;
  assign n62174 = ~n62172 & ~n62173 ;
  assign n62175 = n11623 & ~n62174 ;
  assign n62168 = \P2_P1_uWord_reg[10]/NET0131  & n48581 ;
  assign n62176 = \P2_P1_Datao_reg[26]/NET0131  & ~n48594 ;
  assign n62177 = ~n62168 & ~n62176 ;
  assign n62178 = ~n62175 & n62177 ;
  assign n62180 = \P2_P1_Datao_reg[29]/NET0131  & ~n26030 ;
  assign n62181 = n26006 & n27544 ;
  assign n62182 = ~n62180 & ~n62181 ;
  assign n62183 = n11623 & ~n62182 ;
  assign n62179 = \P2_P1_uWord_reg[13]/NET0131  & n48581 ;
  assign n62184 = \P2_P1_Datao_reg[29]/NET0131  & ~n48594 ;
  assign n62185 = ~n62179 & ~n62184 ;
  assign n62186 = ~n62183 & n62185 ;
  assign n62187 = ~\P2_P1_Flush_reg/NET0131  & n27486 ;
  assign n62188 = n11626 & ~n48581 ;
  assign n62189 = ~n62187 & n62188 ;
  assign n62190 = n52907 & n62189 ;
  assign n62191 = \P2_P1_InstQueueWr_Addr_reg[2]/NET0131  & ~n62190 ;
  assign n62192 = ~n11597 & ~n36673 ;
  assign n62193 = \P2_P1_InstQueueWr_Addr_reg[2]/NET0131  & ~n62192 ;
  assign n62194 = ~n12341 & ~n62193 ;
  assign n62195 = ~n11692 & ~n62194 ;
  assign n62196 = n11597 & ~n12341 ;
  assign n62197 = ~\P2_P1_InstQueueWr_Addr_reg[2]/NET0131  & ~n11594 ;
  assign n62198 = ~n27681 & n62197 ;
  assign n62199 = ~n62196 & n62198 ;
  assign n62200 = ~n11872 & ~n62199 ;
  assign n62201 = ~n62195 & n62200 ;
  assign n62202 = ~n62191 & ~n62201 ;
  assign n62203 = ~\P2_P2_Flush_reg/NET0131  & n27642 ;
  assign n62204 = ~n26792 & ~n27637 ;
  assign n62205 = ~n48491 & n62204 ;
  assign n62206 = ~n62203 & n62205 ;
  assign n62207 = n52964 & n62206 ;
  assign n62208 = \P2_P2_InstQueueWr_Addr_reg[2]/NET0131  & ~n62207 ;
  assign n62209 = \P2_P2_DataWidth_reg[1]/NET0131  & \P2_P2_InstQueueWr_Addr_reg[2]/NET0131  ;
  assign n62210 = ~n27977 & n62209 ;
  assign n62211 = ~n28400 & ~n28948 ;
  assign n62212 = ~n62210 & n62211 ;
  assign n62213 = ~n27613 & ~n62212 ;
  assign n62214 = n27981 & ~n28948 ;
  assign n62215 = ~\P2_P2_InstQueueWr_Addr_reg[2]/NET0131  & ~n27978 ;
  assign n62216 = ~n26800 & n62215 ;
  assign n62217 = ~n62214 & n62216 ;
  assign n62218 = ~n28386 & ~n62217 ;
  assign n62219 = ~n62213 & n62218 ;
  assign n62220 = ~n62208 & ~n62219 ;
  assign n62223 = n8987 & n49732 ;
  assign n62222 = ~\P1_P3_InstQueue_reg[0][2]/NET0131  & ~n49732 ;
  assign n62224 = n10046 & ~n62222 ;
  assign n62225 = ~n62223 & n62224 ;
  assign n62221 = \P1_P3_InstQueue_reg[0][2]/NET0131  & ~n49750 ;
  assign n62226 = \P1_buf2_reg[26]/NET0131  & n49739 ;
  assign n62227 = \P1_buf2_reg[18]/NET0131  & ~n49739 ;
  assign n62228 = n49742 & n62227 ;
  assign n62229 = ~n62226 & ~n62228 ;
  assign n62230 = n11698 & ~n62229 ;
  assign n62231 = \P1_buf2_reg[2]/NET0131  & n49760 ;
  assign n62232 = ~n62230 & ~n62231 ;
  assign n62233 = ~n62221 & n62232 ;
  assign n62234 = ~n62225 & n62233 ;
  assign n62237 = n8987 & n49766 ;
  assign n62236 = ~\P1_P3_InstQueue_reg[10][2]/NET0131  & ~n49766 ;
  assign n62238 = n10046 & ~n62236 ;
  assign n62239 = ~n62237 & n62238 ;
  assign n62235 = \P1_P3_InstQueue_reg[10][2]/NET0131  & ~n49776 ;
  assign n62240 = \P1_buf2_reg[26]/NET0131  & n49770 ;
  assign n62241 = \P1_buf2_reg[18]/NET0131  & n49771 ;
  assign n62242 = ~n62240 & ~n62241 ;
  assign n62243 = n11698 & ~n62242 ;
  assign n62244 = \P1_buf2_reg[2]/NET0131  & n49786 ;
  assign n62245 = ~n62243 & ~n62244 ;
  assign n62246 = ~n62235 & n62245 ;
  assign n62247 = ~n62239 & n62246 ;
  assign n62250 = n8987 & n49792 ;
  assign n62249 = ~\P1_P3_InstQueue_reg[11][2]/NET0131  & ~n49792 ;
  assign n62251 = n10046 & ~n62249 ;
  assign n62252 = ~n62250 & n62251 ;
  assign n62248 = \P1_P3_InstQueue_reg[11][2]/NET0131  & ~n49798 ;
  assign n62253 = \P1_buf2_reg[26]/NET0131  & n49771 ;
  assign n62254 = \P1_buf2_reg[18]/NET0131  & n49768 ;
  assign n62255 = ~n62253 & ~n62254 ;
  assign n62256 = n11698 & ~n62255 ;
  assign n62257 = \P1_buf2_reg[2]/NET0131  & n49808 ;
  assign n62258 = ~n62256 & ~n62257 ;
  assign n62259 = ~n62248 & n62258 ;
  assign n62260 = ~n62252 & n62259 ;
  assign n62263 = n8987 & n49814 ;
  assign n62262 = ~\P1_P3_InstQueue_reg[12][2]/NET0131  & ~n49814 ;
  assign n62264 = n10046 & ~n62262 ;
  assign n62265 = ~n62263 & n62264 ;
  assign n62261 = \P1_P3_InstQueue_reg[12][2]/NET0131  & ~n49819 ;
  assign n62266 = \P1_buf2_reg[26]/NET0131  & n49768 ;
  assign n62267 = \P1_buf2_reg[18]/NET0131  & n49766 ;
  assign n62268 = ~n62266 & ~n62267 ;
  assign n62269 = n11698 & ~n62268 ;
  assign n62270 = \P1_buf2_reg[2]/NET0131  & n49829 ;
  assign n62271 = ~n62269 & ~n62270 ;
  assign n62272 = ~n62261 & n62271 ;
  assign n62273 = ~n62265 & n62272 ;
  assign n62276 = n8987 & n49739 ;
  assign n62275 = ~\P1_P3_InstQueue_reg[13][2]/NET0131  & ~n49739 ;
  assign n62277 = n10046 & ~n62275 ;
  assign n62278 = ~n62276 & n62277 ;
  assign n62274 = \P1_P3_InstQueue_reg[13][2]/NET0131  & ~n49838 ;
  assign n62279 = \P1_buf2_reg[26]/NET0131  & n49766 ;
  assign n62280 = \P1_buf2_reg[18]/NET0131  & ~n49766 ;
  assign n62281 = n49792 & n62280 ;
  assign n62282 = ~n62279 & ~n62281 ;
  assign n62283 = n11698 & ~n62282 ;
  assign n62284 = \P1_buf2_reg[2]/NET0131  & n49848 ;
  assign n62285 = ~n62283 & ~n62284 ;
  assign n62286 = ~n62274 & n62285 ;
  assign n62287 = ~n62278 & n62286 ;
  assign n62290 = n8987 & n49742 ;
  assign n62289 = ~\P1_P3_InstQueue_reg[14][2]/NET0131  & ~n49742 ;
  assign n62291 = n10046 & ~n62289 ;
  assign n62292 = ~n62290 & n62291 ;
  assign n62288 = \P1_P3_InstQueue_reg[14][2]/NET0131  & ~n49856 ;
  assign n62293 = \P1_buf2_reg[26]/NET0131  & n49792 ;
  assign n62294 = \P1_buf2_reg[18]/NET0131  & ~n49792 ;
  assign n62295 = n49814 & n62294 ;
  assign n62296 = ~n62293 & ~n62295 ;
  assign n62297 = n11698 & ~n62296 ;
  assign n62298 = \P1_buf2_reg[2]/NET0131  & n49866 ;
  assign n62299 = ~n62297 & ~n62298 ;
  assign n62300 = ~n62288 & n62299 ;
  assign n62301 = ~n62292 & n62300 ;
  assign n62304 = n8987 & n49735 ;
  assign n62303 = ~\P1_P3_InstQueue_reg[15][2]/NET0131  & ~n49735 ;
  assign n62305 = n10046 & ~n62303 ;
  assign n62306 = ~n62304 & n62305 ;
  assign n62302 = \P1_P3_InstQueue_reg[15][2]/NET0131  & ~n49875 ;
  assign n62307 = \P1_buf2_reg[26]/NET0131  & n49814 ;
  assign n62308 = \P1_buf2_reg[18]/NET0131  & n49739 ;
  assign n62309 = ~n62307 & ~n62308 ;
  assign n62310 = n11698 & ~n62309 ;
  assign n62311 = \P1_buf2_reg[2]/NET0131  & n49885 ;
  assign n62312 = ~n62310 & ~n62311 ;
  assign n62313 = ~n62302 & n62312 ;
  assign n62314 = ~n62306 & n62313 ;
  assign n62317 = n8987 & n49890 ;
  assign n62316 = ~\P1_P3_InstQueue_reg[1][2]/NET0131  & ~n49890 ;
  assign n62318 = n10046 & ~n62316 ;
  assign n62319 = ~n62317 & n62318 ;
  assign n62315 = \P1_P3_InstQueue_reg[1][2]/NET0131  & ~n49895 ;
  assign n62320 = \P1_buf2_reg[26]/NET0131  & n49742 ;
  assign n62321 = \P1_buf2_reg[18]/NET0131  & n49735 ;
  assign n62322 = ~n62320 & ~n62321 ;
  assign n62323 = n11698 & ~n62322 ;
  assign n62324 = \P1_buf2_reg[2]/NET0131  & n49905 ;
  assign n62325 = ~n62323 & ~n62324 ;
  assign n62326 = ~n62315 & n62325 ;
  assign n62327 = ~n62319 & n62326 ;
  assign n62330 = n8987 & n49910 ;
  assign n62329 = ~\P1_P3_InstQueue_reg[2][2]/NET0131  & ~n49910 ;
  assign n62331 = n10046 & ~n62329 ;
  assign n62332 = ~n62330 & n62331 ;
  assign n62328 = \P1_P3_InstQueue_reg[2][2]/NET0131  & ~n49915 ;
  assign n62333 = \P1_buf2_reg[26]/NET0131  & n49735 ;
  assign n62334 = \P1_buf2_reg[18]/NET0131  & n49732 ;
  assign n62335 = ~n62333 & ~n62334 ;
  assign n62336 = n11698 & ~n62335 ;
  assign n62337 = \P1_buf2_reg[2]/NET0131  & n49925 ;
  assign n62338 = ~n62336 & ~n62337 ;
  assign n62339 = ~n62328 & n62338 ;
  assign n62340 = ~n62332 & n62339 ;
  assign n62343 = n8987 & n49930 ;
  assign n62342 = ~\P1_P3_InstQueue_reg[3][2]/NET0131  & ~n49930 ;
  assign n62344 = n10046 & ~n62342 ;
  assign n62345 = ~n62343 & n62344 ;
  assign n62341 = \P1_P3_InstQueue_reg[3][2]/NET0131  & ~n49935 ;
  assign n62346 = \P1_buf2_reg[26]/NET0131  & n49732 ;
  assign n62347 = \P1_buf2_reg[18]/NET0131  & ~n49732 ;
  assign n62348 = n49890 & n62347 ;
  assign n62349 = ~n62346 & ~n62348 ;
  assign n62350 = n11698 & ~n62349 ;
  assign n62351 = \P1_buf2_reg[2]/NET0131  & n49945 ;
  assign n62352 = ~n62350 & ~n62351 ;
  assign n62353 = ~n62341 & n62352 ;
  assign n62354 = ~n62345 & n62353 ;
  assign n62357 = n8987 & n49950 ;
  assign n62356 = ~\P1_P3_InstQueue_reg[4][2]/NET0131  & ~n49950 ;
  assign n62358 = n10046 & ~n62356 ;
  assign n62359 = ~n62357 & n62358 ;
  assign n62355 = \P1_P3_InstQueue_reg[4][2]/NET0131  & ~n49955 ;
  assign n62360 = \P1_buf2_reg[26]/NET0131  & n49890 ;
  assign n62361 = \P1_buf2_reg[18]/NET0131  & ~n49890 ;
  assign n62362 = n49910 & n62361 ;
  assign n62363 = ~n62360 & ~n62362 ;
  assign n62364 = n11698 & ~n62363 ;
  assign n62365 = \P1_buf2_reg[2]/NET0131  & n49965 ;
  assign n62366 = ~n62364 & ~n62365 ;
  assign n62367 = ~n62355 & n62366 ;
  assign n62368 = ~n62359 & n62367 ;
  assign n62371 = n8987 & n49970 ;
  assign n62370 = ~\P1_P3_InstQueue_reg[5][2]/NET0131  & ~n49970 ;
  assign n62372 = n10046 & ~n62370 ;
  assign n62373 = ~n62371 & n62372 ;
  assign n62369 = \P1_P3_InstQueue_reg[5][2]/NET0131  & ~n49975 ;
  assign n62374 = \P1_buf2_reg[26]/NET0131  & n49910 ;
  assign n62375 = \P1_buf2_reg[18]/NET0131  & ~n49910 ;
  assign n62376 = n49930 & n62375 ;
  assign n62377 = ~n62374 & ~n62376 ;
  assign n62378 = n11698 & ~n62377 ;
  assign n62379 = \P1_buf2_reg[2]/NET0131  & n49985 ;
  assign n62380 = ~n62378 & ~n62379 ;
  assign n62381 = ~n62369 & n62380 ;
  assign n62382 = ~n62373 & n62381 ;
  assign n62385 = n8987 & n49990 ;
  assign n62384 = ~\P1_P3_InstQueue_reg[6][2]/NET0131  & ~n49990 ;
  assign n62386 = n10046 & ~n62384 ;
  assign n62387 = ~n62385 & n62386 ;
  assign n62383 = \P1_P3_InstQueue_reg[6][2]/NET0131  & ~n49995 ;
  assign n62388 = \P1_buf2_reg[26]/NET0131  & n49930 ;
  assign n62389 = \P1_buf2_reg[18]/NET0131  & ~n49930 ;
  assign n62390 = n49950 & n62389 ;
  assign n62391 = ~n62388 & ~n62390 ;
  assign n62392 = n11698 & ~n62391 ;
  assign n62393 = \P1_buf2_reg[2]/NET0131  & n50005 ;
  assign n62394 = ~n62392 & ~n62393 ;
  assign n62395 = ~n62383 & n62394 ;
  assign n62396 = ~n62387 & n62395 ;
  assign n62399 = n26959 & n50021 ;
  assign n62398 = ~\P2_P3_InstQueue_reg[0][2]/NET0131  & ~n50021 ;
  assign n62400 = n27788 & ~n62398 ;
  assign n62401 = ~n62399 & n62400 ;
  assign n62397 = \P2_P3_InstQueue_reg[0][2]/NET0131  & ~n50030 ;
  assign n62402 = \P2_buf2_reg[26]/NET0131  & n50012 ;
  assign n62403 = \P2_buf2_reg[18]/NET0131  & n50015 ;
  assign n62404 = ~n62402 & ~n62403 ;
  assign n62405 = n27325 & ~n62404 ;
  assign n62406 = \P2_buf2_reg[2]/NET0131  & n50040 ;
  assign n62407 = ~n62405 & ~n62406 ;
  assign n62408 = ~n62397 & n62407 ;
  assign n62409 = ~n62401 & n62408 ;
  assign n62412 = n26959 & n50051 ;
  assign n62411 = ~\P2_P3_InstQueue_reg[10][2]/NET0131  & ~n50051 ;
  assign n62413 = n27788 & ~n62411 ;
  assign n62414 = ~n62412 & n62413 ;
  assign n62410 = \P2_P3_InstQueue_reg[10][2]/NET0131  & ~n50056 ;
  assign n62415 = \P2_buf2_reg[18]/NET0131  & n50045 ;
  assign n62416 = \P2_buf2_reg[26]/NET0131  & n50046 ;
  assign n62417 = ~n62415 & ~n62416 ;
  assign n62418 = n27325 & ~n62417 ;
  assign n62419 = \P2_buf2_reg[2]/NET0131  & n50066 ;
  assign n62420 = ~n62418 & ~n62419 ;
  assign n62421 = ~n62410 & n62420 ;
  assign n62422 = ~n62414 & n62421 ;
  assign n62425 = n8987 & n49770 ;
  assign n62424 = ~\P1_P3_InstQueue_reg[7][2]/NET0131  & ~n49770 ;
  assign n62426 = n10046 & ~n62424 ;
  assign n62427 = ~n62425 & n62426 ;
  assign n62423 = \P1_P3_InstQueue_reg[7][2]/NET0131  & ~n50075 ;
  assign n62428 = \P1_buf2_reg[26]/NET0131  & n49950 ;
  assign n62429 = \P1_buf2_reg[18]/NET0131  & ~n49950 ;
  assign n62430 = n49970 & n62429 ;
  assign n62431 = ~n62428 & ~n62430 ;
  assign n62432 = n11698 & ~n62431 ;
  assign n62433 = \P1_buf2_reg[2]/NET0131  & n50085 ;
  assign n62434 = ~n62432 & ~n62433 ;
  assign n62435 = ~n62423 & n62434 ;
  assign n62436 = ~n62427 & n62435 ;
  assign n62439 = n26959 & n50094 ;
  assign n62438 = ~\P2_P3_InstQueue_reg[11][2]/NET0131  & ~n50094 ;
  assign n62440 = n27788 & ~n62438 ;
  assign n62441 = ~n62439 & n62440 ;
  assign n62437 = \P2_P3_InstQueue_reg[11][2]/NET0131  & ~n50097 ;
  assign n62442 = \P2_buf2_reg[26]/NET0131  & n50045 ;
  assign n62443 = \P2_buf2_reg[18]/NET0131  & n50053 ;
  assign n62444 = ~n62442 & ~n62443 ;
  assign n62445 = n27325 & ~n62444 ;
  assign n62446 = \P2_buf2_reg[2]/NET0131  & n50107 ;
  assign n62447 = ~n62445 & ~n62446 ;
  assign n62448 = ~n62437 & n62447 ;
  assign n62449 = ~n62441 & n62448 ;
  assign n62452 = n26959 & n50115 ;
  assign n62451 = ~\P2_P3_InstQueue_reg[12][2]/NET0131  & ~n50115 ;
  assign n62453 = n27788 & ~n62451 ;
  assign n62454 = ~n62452 & n62453 ;
  assign n62450 = \P2_P3_InstQueue_reg[12][2]/NET0131  & ~n50118 ;
  assign n62455 = \P2_buf2_reg[26]/NET0131  & n50053 ;
  assign n62456 = \P2_buf2_reg[18]/NET0131  & n50051 ;
  assign n62457 = ~n62455 & ~n62456 ;
  assign n62458 = n27325 & ~n62457 ;
  assign n62459 = \P2_buf2_reg[2]/NET0131  & n50128 ;
  assign n62460 = ~n62458 & ~n62459 ;
  assign n62461 = ~n62450 & n62460 ;
  assign n62462 = ~n62454 & n62461 ;
  assign n62465 = n8987 & n49771 ;
  assign n62464 = ~\P1_P3_InstQueue_reg[8][2]/NET0131  & ~n49771 ;
  assign n62466 = n10046 & ~n62464 ;
  assign n62467 = ~n62465 & n62466 ;
  assign n62463 = \P1_P3_InstQueue_reg[8][2]/NET0131  & ~n50136 ;
  assign n62468 = \P1_buf2_reg[26]/NET0131  & n49970 ;
  assign n62469 = \P1_buf2_reg[18]/NET0131  & ~n49970 ;
  assign n62470 = n49990 & n62469 ;
  assign n62471 = ~n62468 & ~n62470 ;
  assign n62472 = n11698 & ~n62471 ;
  assign n62473 = \P1_buf2_reg[2]/NET0131  & n50146 ;
  assign n62474 = ~n62472 & ~n62473 ;
  assign n62475 = ~n62463 & n62474 ;
  assign n62476 = ~n62467 & n62475 ;
  assign n62479 = n26959 & n50012 ;
  assign n62478 = ~\P2_P3_InstQueue_reg[13][2]/NET0131  & ~n50012 ;
  assign n62480 = n27788 & ~n62478 ;
  assign n62481 = ~n62479 & n62480 ;
  assign n62477 = \P2_P3_InstQueue_reg[13][2]/NET0131  & ~n50155 ;
  assign n62482 = \P2_buf2_reg[26]/NET0131  & n50051 ;
  assign n62483 = \P2_buf2_reg[18]/NET0131  & n50094 ;
  assign n62484 = ~n62482 & ~n62483 ;
  assign n62485 = n27325 & ~n62484 ;
  assign n62486 = \P2_buf2_reg[2]/NET0131  & n50165 ;
  assign n62487 = ~n62485 & ~n62486 ;
  assign n62488 = ~n62477 & n62487 ;
  assign n62489 = ~n62481 & n62488 ;
  assign n62492 = n26959 & n50015 ;
  assign n62491 = ~\P2_P3_InstQueue_reg[14][2]/NET0131  & ~n50015 ;
  assign n62493 = n27788 & ~n62491 ;
  assign n62494 = ~n62492 & n62493 ;
  assign n62490 = \P2_P3_InstQueue_reg[14][2]/NET0131  & ~n50173 ;
  assign n62495 = \P2_buf2_reg[26]/NET0131  & n50094 ;
  assign n62496 = \P2_buf2_reg[18]/NET0131  & n50115 ;
  assign n62497 = ~n62495 & ~n62496 ;
  assign n62498 = n27325 & ~n62497 ;
  assign n62499 = \P2_buf2_reg[2]/NET0131  & n50183 ;
  assign n62500 = ~n62498 & ~n62499 ;
  assign n62501 = ~n62490 & n62500 ;
  assign n62502 = ~n62494 & n62501 ;
  assign n62505 = n8987 & n49768 ;
  assign n62504 = ~\P1_P3_InstQueue_reg[9][2]/NET0131  & ~n49768 ;
  assign n62506 = n10046 & ~n62504 ;
  assign n62507 = ~n62505 & n62506 ;
  assign n62503 = \P1_P3_InstQueue_reg[9][2]/NET0131  & ~n50191 ;
  assign n62508 = \P1_buf2_reg[26]/NET0131  & n49990 ;
  assign n62509 = \P1_buf2_reg[18]/NET0131  & n49770 ;
  assign n62510 = ~n62508 & ~n62509 ;
  assign n62511 = n11698 & ~n62510 ;
  assign n62512 = \P1_buf2_reg[2]/NET0131  & n50201 ;
  assign n62513 = ~n62511 & ~n62512 ;
  assign n62514 = ~n62503 & n62513 ;
  assign n62515 = ~n62507 & n62514 ;
  assign n62518 = n26959 & n50024 ;
  assign n62517 = ~\P2_P3_InstQueue_reg[15][2]/NET0131  & ~n50024 ;
  assign n62519 = n27788 & ~n62517 ;
  assign n62520 = ~n62518 & n62519 ;
  assign n62516 = \P2_P3_InstQueue_reg[15][2]/NET0131  & ~n50210 ;
  assign n62521 = \P2_buf2_reg[26]/NET0131  & n50115 ;
  assign n62522 = \P2_buf2_reg[18]/NET0131  & n50012 ;
  assign n62523 = ~n62521 & ~n62522 ;
  assign n62524 = n27325 & ~n62523 ;
  assign n62525 = \P2_buf2_reg[2]/NET0131  & n50220 ;
  assign n62526 = ~n62524 & ~n62525 ;
  assign n62527 = ~n62516 & n62526 ;
  assign n62528 = ~n62520 & n62527 ;
  assign n62531 = n26959 & n50227 ;
  assign n62530 = ~\P2_P3_InstQueue_reg[1][2]/NET0131  & ~n50227 ;
  assign n62532 = n27788 & ~n62530 ;
  assign n62533 = ~n62531 & n62532 ;
  assign n62529 = \P2_P3_InstQueue_reg[1][2]/NET0131  & ~n50230 ;
  assign n62534 = \P2_buf2_reg[26]/NET0131  & n50015 ;
  assign n62535 = \P2_buf2_reg[18]/NET0131  & n50024 ;
  assign n62536 = ~n62534 & ~n62535 ;
  assign n62537 = n27325 & ~n62536 ;
  assign n62538 = \P2_buf2_reg[2]/NET0131  & n50240 ;
  assign n62539 = ~n62537 & ~n62538 ;
  assign n62540 = ~n62529 & n62539 ;
  assign n62541 = ~n62533 & n62540 ;
  assign n62544 = n26959 & n50247 ;
  assign n62543 = ~\P2_P3_InstQueue_reg[2][2]/NET0131  & ~n50247 ;
  assign n62545 = n27788 & ~n62543 ;
  assign n62546 = ~n62544 & n62545 ;
  assign n62542 = \P2_P3_InstQueue_reg[2][2]/NET0131  & ~n50250 ;
  assign n62547 = \P2_buf2_reg[18]/NET0131  & n50021 ;
  assign n62548 = \P2_buf2_reg[26]/NET0131  & n50024 ;
  assign n62549 = ~n62547 & ~n62548 ;
  assign n62550 = n27325 & ~n62549 ;
  assign n62551 = \P2_buf2_reg[2]/NET0131  & n50260 ;
  assign n62552 = ~n62550 & ~n62551 ;
  assign n62553 = ~n62542 & n62552 ;
  assign n62554 = ~n62546 & n62553 ;
  assign n62557 = n26959 & n50267 ;
  assign n62556 = ~\P2_P3_InstQueue_reg[3][2]/NET0131  & ~n50267 ;
  assign n62558 = n27788 & ~n62556 ;
  assign n62559 = ~n62557 & n62558 ;
  assign n62555 = \P2_P3_InstQueue_reg[3][2]/NET0131  & ~n50270 ;
  assign n62560 = \P2_buf2_reg[26]/NET0131  & n50021 ;
  assign n62561 = \P2_buf2_reg[18]/NET0131  & n50227 ;
  assign n62562 = ~n62560 & ~n62561 ;
  assign n62563 = n27325 & ~n62562 ;
  assign n62564 = \P2_buf2_reg[2]/NET0131  & n50280 ;
  assign n62565 = ~n62563 & ~n62564 ;
  assign n62566 = ~n62555 & n62565 ;
  assign n62567 = ~n62559 & n62566 ;
  assign n62570 = n26959 & n50287 ;
  assign n62569 = ~\P2_P3_InstQueue_reg[4][2]/NET0131  & ~n50287 ;
  assign n62571 = n27788 & ~n62569 ;
  assign n62572 = ~n62570 & n62571 ;
  assign n62568 = \P2_P3_InstQueue_reg[4][2]/NET0131  & ~n50290 ;
  assign n62573 = \P2_buf2_reg[26]/NET0131  & n50227 ;
  assign n62574 = \P2_buf2_reg[18]/NET0131  & n50247 ;
  assign n62575 = ~n62573 & ~n62574 ;
  assign n62576 = n27325 & ~n62575 ;
  assign n62577 = \P2_buf2_reg[2]/NET0131  & n50300 ;
  assign n62578 = ~n62576 & ~n62577 ;
  assign n62579 = ~n62568 & n62578 ;
  assign n62580 = ~n62572 & n62579 ;
  assign n62583 = n26959 & n50307 ;
  assign n62582 = ~\P2_P3_InstQueue_reg[5][2]/NET0131  & ~n50307 ;
  assign n62584 = n27788 & ~n62582 ;
  assign n62585 = ~n62583 & n62584 ;
  assign n62581 = \P2_P3_InstQueue_reg[5][2]/NET0131  & ~n50310 ;
  assign n62586 = \P2_buf2_reg[26]/NET0131  & n50247 ;
  assign n62587 = \P2_buf2_reg[18]/NET0131  & n50267 ;
  assign n62588 = ~n62586 & ~n62587 ;
  assign n62589 = n27325 & ~n62588 ;
  assign n62590 = \P2_buf2_reg[2]/NET0131  & n50320 ;
  assign n62591 = ~n62589 & ~n62590 ;
  assign n62592 = ~n62581 & n62591 ;
  assign n62593 = ~n62585 & n62592 ;
  assign n62596 = n26959 & n50327 ;
  assign n62595 = ~\P2_P3_InstQueue_reg[6][2]/NET0131  & ~n50327 ;
  assign n62597 = n27788 & ~n62595 ;
  assign n62598 = ~n62596 & n62597 ;
  assign n62594 = \P2_P3_InstQueue_reg[6][2]/NET0131  & ~n50330 ;
  assign n62599 = \P2_buf2_reg[26]/NET0131  & n50267 ;
  assign n62600 = \P2_buf2_reg[18]/NET0131  & n50287 ;
  assign n62601 = ~n62599 & ~n62600 ;
  assign n62602 = n27325 & ~n62601 ;
  assign n62603 = \P2_buf2_reg[2]/NET0131  & n50340 ;
  assign n62604 = ~n62602 & ~n62603 ;
  assign n62605 = ~n62594 & n62604 ;
  assign n62606 = ~n62598 & n62605 ;
  assign n62609 = n26959 & n50046 ;
  assign n62608 = ~\P2_P3_InstQueue_reg[7][2]/NET0131  & ~n50046 ;
  assign n62610 = n27788 & ~n62608 ;
  assign n62611 = ~n62609 & n62610 ;
  assign n62607 = \P2_P3_InstQueue_reg[7][2]/NET0131  & ~n50349 ;
  assign n62612 = \P2_buf2_reg[26]/NET0131  & n50287 ;
  assign n62613 = \P2_buf2_reg[18]/NET0131  & n50307 ;
  assign n62614 = ~n62612 & ~n62613 ;
  assign n62615 = n27325 & ~n62614 ;
  assign n62616 = \P2_buf2_reg[2]/NET0131  & n50359 ;
  assign n62617 = ~n62615 & ~n62616 ;
  assign n62618 = ~n62607 & n62617 ;
  assign n62619 = ~n62611 & n62618 ;
  assign n62622 = n26959 & n50045 ;
  assign n62621 = ~\P2_P3_InstQueue_reg[8][2]/NET0131  & ~n50045 ;
  assign n62623 = n27788 & ~n62621 ;
  assign n62624 = ~n62622 & n62623 ;
  assign n62620 = \P2_P3_InstQueue_reg[8][2]/NET0131  & ~n50367 ;
  assign n62625 = \P2_buf2_reg[26]/NET0131  & n50307 ;
  assign n62626 = \P2_buf2_reg[18]/NET0131  & n50327 ;
  assign n62627 = ~n62625 & ~n62626 ;
  assign n62628 = n27325 & ~n62627 ;
  assign n62629 = \P2_buf2_reg[2]/NET0131  & n50377 ;
  assign n62630 = ~n62628 & ~n62629 ;
  assign n62631 = ~n62620 & n62630 ;
  assign n62632 = ~n62624 & n62631 ;
  assign n62635 = n26959 & n50053 ;
  assign n62634 = ~\P2_P3_InstQueue_reg[9][2]/NET0131  & ~n50053 ;
  assign n62636 = n27788 & ~n62634 ;
  assign n62637 = ~n62635 & n62636 ;
  assign n62633 = \P2_P3_InstQueue_reg[9][2]/NET0131  & ~n50385 ;
  assign n62638 = \P2_buf2_reg[26]/NET0131  & n50327 ;
  assign n62639 = \P2_buf2_reg[18]/NET0131  & n50046 ;
  assign n62640 = ~n62638 & ~n62639 ;
  assign n62641 = n27325 & ~n62640 ;
  assign n62642 = \P2_buf2_reg[2]/NET0131  & n50395 ;
  assign n62643 = ~n62641 & ~n62642 ;
  assign n62644 = ~n62633 & n62643 ;
  assign n62645 = ~n62637 & n62644 ;
  assign n62649 = ~\P1_P1_EAX_reg[13]/NET0131  & n26162 ;
  assign n62648 = ~\P1_P1_Datao_reg[13]/NET0131  & ~n26162 ;
  assign n62650 = n8355 & ~n62648 ;
  assign n62651 = ~n62649 & n62650 ;
  assign n62646 = \P1_P1_lWord_reg[13]/NET0131  & n27790 ;
  assign n62647 = \P1_P1_Datao_reg[13]/NET0131  & ~n48479 ;
  assign n62652 = ~n62646 & ~n62647 ;
  assign n62653 = ~n62651 & n62652 ;
  assign n62657 = ~\P1_P1_EAX_reg[14]/NET0131  & n26162 ;
  assign n62656 = ~\P1_P1_Datao_reg[14]/NET0131  & ~n26162 ;
  assign n62658 = n8355 & ~n62656 ;
  assign n62659 = ~n62657 & n62658 ;
  assign n62654 = \P1_P1_lWord_reg[14]/NET0131  & n27790 ;
  assign n62655 = \P1_P1_Datao_reg[14]/NET0131  & ~n48479 ;
  assign n62660 = ~n62654 & ~n62655 ;
  assign n62661 = ~n62659 & n62660 ;
  assign n62665 = ~\P1_P1_EAX_reg[1]/NET0131  & n26162 ;
  assign n62664 = ~\P1_P1_Datao_reg[1]/NET0131  & ~n26162 ;
  assign n62666 = n8355 & ~n62664 ;
  assign n62667 = ~n62665 & n62666 ;
  assign n62662 = \P1_P1_lWord_reg[1]/NET0131  & n27790 ;
  assign n62663 = \P1_P1_Datao_reg[1]/NET0131  & ~n48479 ;
  assign n62668 = ~n62662 & ~n62663 ;
  assign n62669 = ~n62667 & n62668 ;
  assign n62673 = ~\P1_P1_EAX_reg[2]/NET0131  & n26162 ;
  assign n62672 = ~\P1_P1_Datao_reg[2]/NET0131  & ~n26162 ;
  assign n62674 = n8355 & ~n62672 ;
  assign n62675 = ~n62673 & n62674 ;
  assign n62670 = \P1_P1_lWord_reg[2]/NET0131  & n27790 ;
  assign n62671 = \P1_P1_Datao_reg[2]/NET0131  & ~n48479 ;
  assign n62676 = ~n62670 & ~n62671 ;
  assign n62677 = ~n62675 & n62676 ;
  assign n62681 = ~\P1_P1_EAX_reg[3]/NET0131  & n26162 ;
  assign n62680 = ~\P1_P1_Datao_reg[3]/NET0131  & ~n26162 ;
  assign n62682 = n8355 & ~n62680 ;
  assign n62683 = ~n62681 & n62682 ;
  assign n62678 = \P1_P1_lWord_reg[3]/NET0131  & n27790 ;
  assign n62679 = \P1_P1_Datao_reg[3]/NET0131  & ~n48479 ;
  assign n62684 = ~n62678 & ~n62679 ;
  assign n62685 = ~n62683 & n62684 ;
  assign n62689 = ~\P1_P1_EAX_reg[4]/NET0131  & n26162 ;
  assign n62688 = ~\P1_P1_Datao_reg[4]/NET0131  & ~n26162 ;
  assign n62690 = n8355 & ~n62688 ;
  assign n62691 = ~n62689 & n62690 ;
  assign n62686 = \P1_P1_lWord_reg[4]/NET0131  & n27790 ;
  assign n62687 = \P1_P1_Datao_reg[4]/NET0131  & ~n48479 ;
  assign n62692 = ~n62686 & ~n62687 ;
  assign n62693 = ~n62691 & n62692 ;
  assign n62697 = ~\P1_P1_EAX_reg[5]/NET0131  & n26162 ;
  assign n62696 = ~\P1_P1_Datao_reg[5]/NET0131  & ~n26162 ;
  assign n62698 = n8355 & ~n62696 ;
  assign n62699 = ~n62697 & n62698 ;
  assign n62694 = \P1_P1_lWord_reg[5]/NET0131  & n27790 ;
  assign n62695 = \P1_P1_Datao_reg[5]/NET0131  & ~n48479 ;
  assign n62700 = ~n62694 & ~n62695 ;
  assign n62701 = ~n62699 & n62700 ;
  assign n62705 = ~\P1_P1_EAX_reg[6]/NET0131  & n26162 ;
  assign n62704 = ~\P1_P1_Datao_reg[6]/NET0131  & ~n26162 ;
  assign n62706 = n8355 & ~n62704 ;
  assign n62707 = ~n62705 & n62706 ;
  assign n62702 = \P1_P1_lWord_reg[6]/NET0131  & n27790 ;
  assign n62703 = \P1_P1_Datao_reg[6]/NET0131  & ~n48479 ;
  assign n62708 = ~n62702 & ~n62703 ;
  assign n62709 = ~n62707 & n62708 ;
  assign n62713 = ~\P1_P1_EAX_reg[7]/NET0131  & n26162 ;
  assign n62712 = ~\P1_P1_Datao_reg[7]/NET0131  & ~n26162 ;
  assign n62714 = n8355 & ~n62712 ;
  assign n62715 = ~n62713 & n62714 ;
  assign n62710 = \P1_P1_lWord_reg[7]/NET0131  & n27790 ;
  assign n62711 = \P1_P1_Datao_reg[7]/NET0131  & ~n48479 ;
  assign n62716 = ~n62710 & ~n62711 ;
  assign n62717 = ~n62715 & n62716 ;
  assign n62721 = ~\P1_P1_EAX_reg[8]/NET0131  & n26162 ;
  assign n62720 = ~\P1_P1_Datao_reg[8]/NET0131  & ~n26162 ;
  assign n62722 = n8355 & ~n62720 ;
  assign n62723 = ~n62721 & n62722 ;
  assign n62718 = \P1_P1_lWord_reg[8]/NET0131  & n27790 ;
  assign n62719 = \P1_P1_Datao_reg[8]/NET0131  & ~n48479 ;
  assign n62724 = ~n62718 & ~n62719 ;
  assign n62725 = ~n62723 & n62724 ;
  assign n62729 = ~\P1_P1_EAX_reg[9]/NET0131  & n26162 ;
  assign n62728 = ~\P1_P1_Datao_reg[9]/NET0131  & ~n26162 ;
  assign n62730 = n8355 & ~n62728 ;
  assign n62731 = ~n62729 & n62730 ;
  assign n62726 = \P1_P1_lWord_reg[9]/NET0131  & n27790 ;
  assign n62727 = \P1_P1_Datao_reg[9]/NET0131  & ~n48479 ;
  assign n62732 = ~n62726 & ~n62727 ;
  assign n62733 = ~n62731 & n62732 ;
  assign n62737 = ~\P2_P2_EAX_reg[0]/NET0131  & n26699 ;
  assign n62736 = ~\P2_P2_Datao_reg[0]/NET0131  & ~n26699 ;
  assign n62738 = n26792 & ~n62736 ;
  assign n62739 = ~n62737 & n62738 ;
  assign n62734 = \P2_P2_lWord_reg[0]/NET0131  & n48491 ;
  assign n62735 = \P2_P2_Datao_reg[0]/NET0131  & ~n48508 ;
  assign n62740 = ~n62734 & ~n62735 ;
  assign n62741 = ~n62739 & n62740 ;
  assign n62745 = ~\P2_P2_EAX_reg[10]/NET0131  & n26699 ;
  assign n62744 = ~\P2_P2_Datao_reg[10]/NET0131  & ~n26699 ;
  assign n62746 = n26792 & ~n62744 ;
  assign n62747 = ~n62745 & n62746 ;
  assign n62742 = \P2_P2_lWord_reg[10]/NET0131  & n48491 ;
  assign n62743 = \P2_P2_Datao_reg[10]/NET0131  & ~n48508 ;
  assign n62748 = ~n62742 & ~n62743 ;
  assign n62749 = ~n62747 & n62748 ;
  assign n62753 = ~\P2_P2_EAX_reg[11]/NET0131  & n26699 ;
  assign n62752 = ~\P2_P2_Datao_reg[11]/NET0131  & ~n26699 ;
  assign n62754 = n26792 & ~n62752 ;
  assign n62755 = ~n62753 & n62754 ;
  assign n62750 = \P2_P2_lWord_reg[11]/NET0131  & n48491 ;
  assign n62751 = \P2_P2_Datao_reg[11]/NET0131  & ~n48508 ;
  assign n62756 = ~n62750 & ~n62751 ;
  assign n62757 = ~n62755 & n62756 ;
  assign n62761 = ~\P2_P2_EAX_reg[12]/NET0131  & n26699 ;
  assign n62760 = ~\P2_P2_Datao_reg[12]/NET0131  & ~n26699 ;
  assign n62762 = n26792 & ~n62760 ;
  assign n62763 = ~n62761 & n62762 ;
  assign n62758 = \P2_P2_lWord_reg[12]/NET0131  & n48491 ;
  assign n62759 = \P2_P2_Datao_reg[12]/NET0131  & ~n48508 ;
  assign n62764 = ~n62758 & ~n62759 ;
  assign n62765 = ~n62763 & n62764 ;
  assign n62769 = ~\P2_P2_EAX_reg[13]/NET0131  & n26699 ;
  assign n62768 = ~\P2_P2_Datao_reg[13]/NET0131  & ~n26699 ;
  assign n62770 = n26792 & ~n62768 ;
  assign n62771 = ~n62769 & n62770 ;
  assign n62766 = \P2_P2_lWord_reg[13]/NET0131  & n48491 ;
  assign n62767 = \P2_P2_Datao_reg[13]/NET0131  & ~n48508 ;
  assign n62772 = ~n62766 & ~n62767 ;
  assign n62773 = ~n62771 & n62772 ;
  assign n62777 = ~\P2_P2_EAX_reg[14]/NET0131  & n26699 ;
  assign n62776 = ~\P2_P2_Datao_reg[14]/NET0131  & ~n26699 ;
  assign n62778 = n26792 & ~n62776 ;
  assign n62779 = ~n62777 & n62778 ;
  assign n62774 = \P2_P2_lWord_reg[14]/NET0131  & n48491 ;
  assign n62775 = \P2_P2_Datao_reg[14]/NET0131  & ~n48508 ;
  assign n62780 = ~n62774 & ~n62775 ;
  assign n62781 = ~n62779 & n62780 ;
  assign n62785 = ~\P2_P2_EAX_reg[15]/NET0131  & n26699 ;
  assign n62784 = ~\P2_P2_Datao_reg[15]/NET0131  & ~n26699 ;
  assign n62786 = n26792 & ~n62784 ;
  assign n62787 = ~n62785 & n62786 ;
  assign n62782 = \P2_P2_lWord_reg[15]/NET0131  & n48491 ;
  assign n62783 = \P2_P2_Datao_reg[15]/NET0131  & ~n48508 ;
  assign n62788 = ~n62782 & ~n62783 ;
  assign n62789 = ~n62787 & n62788 ;
  assign n62793 = ~\P2_P2_EAX_reg[1]/NET0131  & n26699 ;
  assign n62792 = ~\P2_P2_Datao_reg[1]/NET0131  & ~n26699 ;
  assign n62794 = n26792 & ~n62792 ;
  assign n62795 = ~n62793 & n62794 ;
  assign n62790 = \P2_P2_lWord_reg[1]/NET0131  & n48491 ;
  assign n62791 = \P2_P2_Datao_reg[1]/NET0131  & ~n48508 ;
  assign n62796 = ~n62790 & ~n62791 ;
  assign n62797 = ~n62795 & n62796 ;
  assign n62801 = ~\P2_P2_EAX_reg[2]/NET0131  & n26699 ;
  assign n62800 = ~\P2_P2_Datao_reg[2]/NET0131  & ~n26699 ;
  assign n62802 = n26792 & ~n62800 ;
  assign n62803 = ~n62801 & n62802 ;
  assign n62798 = \P2_P2_lWord_reg[2]/NET0131  & n48491 ;
  assign n62799 = \P2_P2_Datao_reg[2]/NET0131  & ~n48508 ;
  assign n62804 = ~n62798 & ~n62799 ;
  assign n62805 = ~n62803 & n62804 ;
  assign n62809 = ~\P2_P2_EAX_reg[3]/NET0131  & n26699 ;
  assign n62808 = ~\P2_P2_Datao_reg[3]/NET0131  & ~n26699 ;
  assign n62810 = n26792 & ~n62808 ;
  assign n62811 = ~n62809 & n62810 ;
  assign n62806 = \P2_P2_lWord_reg[3]/NET0131  & n48491 ;
  assign n62807 = \P2_P2_Datao_reg[3]/NET0131  & ~n48508 ;
  assign n62812 = ~n62806 & ~n62807 ;
  assign n62813 = ~n62811 & n62812 ;
  assign n62817 = ~\P2_P2_EAX_reg[4]/NET0131  & n26699 ;
  assign n62816 = ~\P2_P2_Datao_reg[4]/NET0131  & ~n26699 ;
  assign n62818 = n26792 & ~n62816 ;
  assign n62819 = ~n62817 & n62818 ;
  assign n62814 = \P2_P2_lWord_reg[4]/NET0131  & n48491 ;
  assign n62815 = \P2_P2_Datao_reg[4]/NET0131  & ~n48508 ;
  assign n62820 = ~n62814 & ~n62815 ;
  assign n62821 = ~n62819 & n62820 ;
  assign n62825 = ~\P2_P2_EAX_reg[5]/NET0131  & n26699 ;
  assign n62824 = ~\P2_P2_Datao_reg[5]/NET0131  & ~n26699 ;
  assign n62826 = n26792 & ~n62824 ;
  assign n62827 = ~n62825 & n62826 ;
  assign n62822 = \P2_P2_lWord_reg[5]/NET0131  & n48491 ;
  assign n62823 = \P2_P2_Datao_reg[5]/NET0131  & ~n48508 ;
  assign n62828 = ~n62822 & ~n62823 ;
  assign n62829 = ~n62827 & n62828 ;
  assign n62833 = ~\P2_P2_EAX_reg[6]/NET0131  & n26699 ;
  assign n62832 = ~\P2_P2_Datao_reg[6]/NET0131  & ~n26699 ;
  assign n62834 = n26792 & ~n62832 ;
  assign n62835 = ~n62833 & n62834 ;
  assign n62830 = \P2_P2_lWord_reg[6]/NET0131  & n48491 ;
  assign n62831 = \P2_P2_Datao_reg[6]/NET0131  & ~n48508 ;
  assign n62836 = ~n62830 & ~n62831 ;
  assign n62837 = ~n62835 & n62836 ;
  assign n62841 = ~\P2_P2_EAX_reg[7]/NET0131  & n26699 ;
  assign n62840 = ~\P2_P2_Datao_reg[7]/NET0131  & ~n26699 ;
  assign n62842 = n26792 & ~n62840 ;
  assign n62843 = ~n62841 & n62842 ;
  assign n62838 = \P2_P2_lWord_reg[7]/NET0131  & n48491 ;
  assign n62839 = \P2_P2_Datao_reg[7]/NET0131  & ~n48508 ;
  assign n62844 = ~n62838 & ~n62839 ;
  assign n62845 = ~n62843 & n62844 ;
  assign n62849 = ~\P2_P2_EAX_reg[8]/NET0131  & n26699 ;
  assign n62848 = ~\P2_P2_Datao_reg[8]/NET0131  & ~n26699 ;
  assign n62850 = n26792 & ~n62848 ;
  assign n62851 = ~n62849 & n62850 ;
  assign n62846 = \P2_P2_lWord_reg[8]/NET0131  & n48491 ;
  assign n62847 = \P2_P2_Datao_reg[8]/NET0131  & ~n48508 ;
  assign n62852 = ~n62846 & ~n62847 ;
  assign n62853 = ~n62851 & n62852 ;
  assign n62857 = ~\P2_P2_EAX_reg[9]/NET0131  & n26699 ;
  assign n62856 = ~\P2_P2_Datao_reg[9]/NET0131  & ~n26699 ;
  assign n62858 = n26792 & ~n62856 ;
  assign n62859 = ~n62857 & n62858 ;
  assign n62854 = \P2_P2_lWord_reg[9]/NET0131  & n48491 ;
  assign n62855 = \P2_P2_Datao_reg[9]/NET0131  & ~n48508 ;
  assign n62860 = ~n62854 & ~n62855 ;
  assign n62861 = ~n62859 & n62860 ;
  assign n62865 = ~\P2_P3_EAX_reg[0]/NET0131  & n27223 ;
  assign n62864 = ~\P2_P3_Datao_reg[0]/NET0131  & ~n27223 ;
  assign n62866 = n27308 & ~n62864 ;
  assign n62867 = ~n62865 & n62866 ;
  assign n62862 = \P2_P3_lWord_reg[0]/NET0131  & n48523 ;
  assign n62863 = \P2_P3_Datao_reg[0]/NET0131  & ~n48540 ;
  assign n62868 = ~n62862 & ~n62863 ;
  assign n62869 = ~n62867 & n62868 ;
  assign n62873 = ~\P2_P3_EAX_reg[10]/NET0131  & n27223 ;
  assign n62872 = ~\P2_P3_Datao_reg[10]/NET0131  & ~n27223 ;
  assign n62874 = n27308 & ~n62872 ;
  assign n62875 = ~n62873 & n62874 ;
  assign n62870 = \P2_P3_lWord_reg[10]/NET0131  & n48523 ;
  assign n62871 = \P2_P3_Datao_reg[10]/NET0131  & ~n48540 ;
  assign n62876 = ~n62870 & ~n62871 ;
  assign n62877 = ~n62875 & n62876 ;
  assign n62881 = ~\P2_P3_EAX_reg[11]/NET0131  & n27223 ;
  assign n62880 = ~\P2_P3_Datao_reg[11]/NET0131  & ~n27223 ;
  assign n62882 = n27308 & ~n62880 ;
  assign n62883 = ~n62881 & n62882 ;
  assign n62878 = \P2_P3_lWord_reg[11]/NET0131  & n48523 ;
  assign n62879 = \P2_P3_Datao_reg[11]/NET0131  & ~n48540 ;
  assign n62884 = ~n62878 & ~n62879 ;
  assign n62885 = ~n62883 & n62884 ;
  assign n62889 = ~\P2_P3_EAX_reg[12]/NET0131  & n27223 ;
  assign n62888 = ~\P2_P3_Datao_reg[12]/NET0131  & ~n27223 ;
  assign n62890 = n27308 & ~n62888 ;
  assign n62891 = ~n62889 & n62890 ;
  assign n62886 = \P2_P3_lWord_reg[12]/NET0131  & n48523 ;
  assign n62887 = \P2_P3_Datao_reg[12]/NET0131  & ~n48540 ;
  assign n62892 = ~n62886 & ~n62887 ;
  assign n62893 = ~n62891 & n62892 ;
  assign n62897 = ~\P2_P3_EAX_reg[13]/NET0131  & n27223 ;
  assign n62896 = ~\P2_P3_Datao_reg[13]/NET0131  & ~n27223 ;
  assign n62898 = n27308 & ~n62896 ;
  assign n62899 = ~n62897 & n62898 ;
  assign n62894 = \P2_P3_lWord_reg[13]/NET0131  & n48523 ;
  assign n62895 = \P2_P3_Datao_reg[13]/NET0131  & ~n48540 ;
  assign n62900 = ~n62894 & ~n62895 ;
  assign n62901 = ~n62899 & n62900 ;
  assign n62905 = ~\P2_P3_EAX_reg[14]/NET0131  & n27223 ;
  assign n62904 = ~\P2_P3_Datao_reg[14]/NET0131  & ~n27223 ;
  assign n62906 = n27308 & ~n62904 ;
  assign n62907 = ~n62905 & n62906 ;
  assign n62902 = \P2_P3_lWord_reg[14]/NET0131  & n48523 ;
  assign n62903 = \P2_P3_Datao_reg[14]/NET0131  & ~n48540 ;
  assign n62908 = ~n62902 & ~n62903 ;
  assign n62909 = ~n62907 & n62908 ;
  assign n62913 = ~\P2_P3_EAX_reg[15]/NET0131  & n27223 ;
  assign n62912 = ~\P2_P3_Datao_reg[15]/NET0131  & ~n27223 ;
  assign n62914 = n27308 & ~n62912 ;
  assign n62915 = ~n62913 & n62914 ;
  assign n62910 = \P2_P3_lWord_reg[15]/NET0131  & n48523 ;
  assign n62911 = \P2_P3_Datao_reg[15]/NET0131  & ~n48540 ;
  assign n62916 = ~n62910 & ~n62911 ;
  assign n62917 = ~n62915 & n62916 ;
  assign n62921 = ~\P2_P3_EAX_reg[1]/NET0131  & n27223 ;
  assign n62920 = ~\P2_P3_Datao_reg[1]/NET0131  & ~n27223 ;
  assign n62922 = n27308 & ~n62920 ;
  assign n62923 = ~n62921 & n62922 ;
  assign n62918 = \P2_P3_lWord_reg[1]/NET0131  & n48523 ;
  assign n62919 = \P2_P3_Datao_reg[1]/NET0131  & ~n48540 ;
  assign n62924 = ~n62918 & ~n62919 ;
  assign n62925 = ~n62923 & n62924 ;
  assign n62929 = ~\P2_P3_EAX_reg[2]/NET0131  & n27223 ;
  assign n62928 = ~\P2_P3_Datao_reg[2]/NET0131  & ~n27223 ;
  assign n62930 = n27308 & ~n62928 ;
  assign n62931 = ~n62929 & n62930 ;
  assign n62926 = \P2_P3_lWord_reg[2]/NET0131  & n48523 ;
  assign n62927 = \P2_P3_Datao_reg[2]/NET0131  & ~n48540 ;
  assign n62932 = ~n62926 & ~n62927 ;
  assign n62933 = ~n62931 & n62932 ;
  assign n62937 = ~\P2_P3_EAX_reg[3]/NET0131  & n27223 ;
  assign n62936 = ~\P2_P3_Datao_reg[3]/NET0131  & ~n27223 ;
  assign n62938 = n27308 & ~n62936 ;
  assign n62939 = ~n62937 & n62938 ;
  assign n62934 = \P2_P3_lWord_reg[3]/NET0131  & n48523 ;
  assign n62935 = \P2_P3_Datao_reg[3]/NET0131  & ~n48540 ;
  assign n62940 = ~n62934 & ~n62935 ;
  assign n62941 = ~n62939 & n62940 ;
  assign n62945 = ~\P2_P3_EAX_reg[4]/NET0131  & n27223 ;
  assign n62944 = ~\P2_P3_Datao_reg[4]/NET0131  & ~n27223 ;
  assign n62946 = n27308 & ~n62944 ;
  assign n62947 = ~n62945 & n62946 ;
  assign n62942 = \P2_P3_lWord_reg[4]/NET0131  & n48523 ;
  assign n62943 = \P2_P3_Datao_reg[4]/NET0131  & ~n48540 ;
  assign n62948 = ~n62942 & ~n62943 ;
  assign n62949 = ~n62947 & n62948 ;
  assign n62953 = ~\P2_P3_EAX_reg[5]/NET0131  & n27223 ;
  assign n62952 = ~\P2_P3_Datao_reg[5]/NET0131  & ~n27223 ;
  assign n62954 = n27308 & ~n62952 ;
  assign n62955 = ~n62953 & n62954 ;
  assign n62950 = \P2_P3_lWord_reg[5]/NET0131  & n48523 ;
  assign n62951 = \P2_P3_Datao_reg[5]/NET0131  & ~n48540 ;
  assign n62956 = ~n62950 & ~n62951 ;
  assign n62957 = ~n62955 & n62956 ;
  assign n62961 = ~\P2_P3_EAX_reg[6]/NET0131  & n27223 ;
  assign n62960 = ~\P2_P3_Datao_reg[6]/NET0131  & ~n27223 ;
  assign n62962 = n27308 & ~n62960 ;
  assign n62963 = ~n62961 & n62962 ;
  assign n62958 = \P2_P3_lWord_reg[6]/NET0131  & n48523 ;
  assign n62959 = \P2_P3_Datao_reg[6]/NET0131  & ~n48540 ;
  assign n62964 = ~n62958 & ~n62959 ;
  assign n62965 = ~n62963 & n62964 ;
  assign n62969 = ~\P2_P3_EAX_reg[7]/NET0131  & n27223 ;
  assign n62968 = ~\P2_P3_Datao_reg[7]/NET0131  & ~n27223 ;
  assign n62970 = n27308 & ~n62968 ;
  assign n62971 = ~n62969 & n62970 ;
  assign n62966 = \P2_P3_lWord_reg[7]/NET0131  & n48523 ;
  assign n62967 = \P2_P3_Datao_reg[7]/NET0131  & ~n48540 ;
  assign n62972 = ~n62966 & ~n62967 ;
  assign n62973 = ~n62971 & n62972 ;
  assign n62977 = ~\P2_P3_EAX_reg[8]/NET0131  & n27223 ;
  assign n62976 = ~\P2_P3_Datao_reg[8]/NET0131  & ~n27223 ;
  assign n62978 = n27308 & ~n62976 ;
  assign n62979 = ~n62977 & n62978 ;
  assign n62974 = \P2_P3_lWord_reg[8]/NET0131  & n48523 ;
  assign n62975 = \P2_P3_Datao_reg[8]/NET0131  & ~n48540 ;
  assign n62980 = ~n62974 & ~n62975 ;
  assign n62981 = ~n62979 & n62980 ;
  assign n62985 = ~\P2_P3_EAX_reg[9]/NET0131  & n27223 ;
  assign n62984 = ~\P2_P3_Datao_reg[9]/NET0131  & ~n27223 ;
  assign n62986 = n27308 & ~n62984 ;
  assign n62987 = ~n62985 & n62986 ;
  assign n62982 = \P2_P3_lWord_reg[9]/NET0131  & n48523 ;
  assign n62983 = \P2_P3_Datao_reg[9]/NET0131  & ~n48540 ;
  assign n62988 = ~n62982 & ~n62983 ;
  assign n62989 = ~n62987 & n62988 ;
  assign n62993 = ~\P1_P2_EAX_reg[0]/NET0131  & n25847 ;
  assign n62992 = ~\P1_P2_Datao_reg[0]/NET0131  & ~n25847 ;
  assign n62994 = n25918 & ~n62992 ;
  assign n62995 = ~n62993 & n62994 ;
  assign n62990 = \P1_P2_lWord_reg[0]/NET0131  & n25922 ;
  assign n62991 = \P1_P2_Datao_reg[0]/NET0131  & ~n48566 ;
  assign n62996 = ~n62990 & ~n62991 ;
  assign n62997 = ~n62995 & n62996 ;
  assign n63001 = ~\P1_P2_EAX_reg[10]/NET0131  & n25847 ;
  assign n63000 = ~\P1_P2_Datao_reg[10]/NET0131  & ~n25847 ;
  assign n63002 = n25918 & ~n63000 ;
  assign n63003 = ~n63001 & n63002 ;
  assign n62998 = \P1_P2_lWord_reg[10]/NET0131  & n25922 ;
  assign n62999 = \P1_P2_Datao_reg[10]/NET0131  & ~n48566 ;
  assign n63004 = ~n62998 & ~n62999 ;
  assign n63005 = ~n63003 & n63004 ;
  assign n63009 = ~\P1_P2_EAX_reg[11]/NET0131  & n25847 ;
  assign n63008 = ~\P1_P2_Datao_reg[11]/NET0131  & ~n25847 ;
  assign n63010 = n25918 & ~n63008 ;
  assign n63011 = ~n63009 & n63010 ;
  assign n63006 = \P1_P2_lWord_reg[11]/NET0131  & n25922 ;
  assign n63007 = \P1_P2_Datao_reg[11]/NET0131  & ~n48566 ;
  assign n63012 = ~n63006 & ~n63007 ;
  assign n63013 = ~n63011 & n63012 ;
  assign n63017 = ~\P1_P2_EAX_reg[12]/NET0131  & n25847 ;
  assign n63016 = ~\P1_P2_Datao_reg[12]/NET0131  & ~n25847 ;
  assign n63018 = n25918 & ~n63016 ;
  assign n63019 = ~n63017 & n63018 ;
  assign n63014 = \P1_P2_lWord_reg[12]/NET0131  & n25922 ;
  assign n63015 = \P1_P2_Datao_reg[12]/NET0131  & ~n48566 ;
  assign n63020 = ~n63014 & ~n63015 ;
  assign n63021 = ~n63019 & n63020 ;
  assign n63025 = ~\P1_P2_EAX_reg[13]/NET0131  & n25847 ;
  assign n63024 = ~\P1_P2_Datao_reg[13]/NET0131  & ~n25847 ;
  assign n63026 = n25918 & ~n63024 ;
  assign n63027 = ~n63025 & n63026 ;
  assign n63022 = \P1_P2_lWord_reg[13]/NET0131  & n25922 ;
  assign n63023 = \P1_P2_Datao_reg[13]/NET0131  & ~n48566 ;
  assign n63028 = ~n63022 & ~n63023 ;
  assign n63029 = ~n63027 & n63028 ;
  assign n63033 = ~\P1_P2_EAX_reg[14]/NET0131  & n25847 ;
  assign n63032 = ~\P1_P2_Datao_reg[14]/NET0131  & ~n25847 ;
  assign n63034 = n25918 & ~n63032 ;
  assign n63035 = ~n63033 & n63034 ;
  assign n63030 = \P1_P2_lWord_reg[14]/NET0131  & n25922 ;
  assign n63031 = \P1_P2_Datao_reg[14]/NET0131  & ~n48566 ;
  assign n63036 = ~n63030 & ~n63031 ;
  assign n63037 = ~n63035 & n63036 ;
  assign n63041 = ~\P1_P2_EAX_reg[15]/NET0131  & n25847 ;
  assign n63040 = ~\P1_P2_Datao_reg[15]/NET0131  & ~n25847 ;
  assign n63042 = n25918 & ~n63040 ;
  assign n63043 = ~n63041 & n63042 ;
  assign n63038 = \P1_P2_lWord_reg[15]/NET0131  & n25922 ;
  assign n63039 = \P1_P2_Datao_reg[15]/NET0131  & ~n48566 ;
  assign n63044 = ~n63038 & ~n63039 ;
  assign n63045 = ~n63043 & n63044 ;
  assign n63049 = ~\P1_P2_EAX_reg[1]/NET0131  & n25847 ;
  assign n63048 = ~\P1_P2_Datao_reg[1]/NET0131  & ~n25847 ;
  assign n63050 = n25918 & ~n63048 ;
  assign n63051 = ~n63049 & n63050 ;
  assign n63046 = \P1_P2_lWord_reg[1]/NET0131  & n25922 ;
  assign n63047 = \P1_P2_Datao_reg[1]/NET0131  & ~n48566 ;
  assign n63052 = ~n63046 & ~n63047 ;
  assign n63053 = ~n63051 & n63052 ;
  assign n63057 = ~\P1_P2_EAX_reg[2]/NET0131  & n25847 ;
  assign n63056 = ~\P1_P2_Datao_reg[2]/NET0131  & ~n25847 ;
  assign n63058 = n25918 & ~n63056 ;
  assign n63059 = ~n63057 & n63058 ;
  assign n63054 = \P1_P2_lWord_reg[2]/NET0131  & n25922 ;
  assign n63055 = \P1_P2_Datao_reg[2]/NET0131  & ~n48566 ;
  assign n63060 = ~n63054 & ~n63055 ;
  assign n63061 = ~n63059 & n63060 ;
  assign n63065 = ~\P1_P2_EAX_reg[3]/NET0131  & n25847 ;
  assign n63064 = ~\P1_P2_Datao_reg[3]/NET0131  & ~n25847 ;
  assign n63066 = n25918 & ~n63064 ;
  assign n63067 = ~n63065 & n63066 ;
  assign n63062 = \P1_P2_lWord_reg[3]/NET0131  & n25922 ;
  assign n63063 = \P1_P2_Datao_reg[3]/NET0131  & ~n48566 ;
  assign n63068 = ~n63062 & ~n63063 ;
  assign n63069 = ~n63067 & n63068 ;
  assign n63073 = ~\P1_P2_EAX_reg[4]/NET0131  & n25847 ;
  assign n63072 = ~\P1_P2_Datao_reg[4]/NET0131  & ~n25847 ;
  assign n63074 = n25918 & ~n63072 ;
  assign n63075 = ~n63073 & n63074 ;
  assign n63070 = \P1_P2_lWord_reg[4]/NET0131  & n25922 ;
  assign n63071 = \P1_P2_Datao_reg[4]/NET0131  & ~n48566 ;
  assign n63076 = ~n63070 & ~n63071 ;
  assign n63077 = ~n63075 & n63076 ;
  assign n63081 = ~\P1_P2_EAX_reg[5]/NET0131  & n25847 ;
  assign n63080 = ~\P1_P2_Datao_reg[5]/NET0131  & ~n25847 ;
  assign n63082 = n25918 & ~n63080 ;
  assign n63083 = ~n63081 & n63082 ;
  assign n63078 = \P1_P2_lWord_reg[5]/NET0131  & n25922 ;
  assign n63079 = \P1_P2_Datao_reg[5]/NET0131  & ~n48566 ;
  assign n63084 = ~n63078 & ~n63079 ;
  assign n63085 = ~n63083 & n63084 ;
  assign n63089 = ~\P1_P2_EAX_reg[6]/NET0131  & n25847 ;
  assign n63088 = ~\P1_P2_Datao_reg[6]/NET0131  & ~n25847 ;
  assign n63090 = n25918 & ~n63088 ;
  assign n63091 = ~n63089 & n63090 ;
  assign n63086 = \P1_P2_lWord_reg[6]/NET0131  & n25922 ;
  assign n63087 = \P1_P2_Datao_reg[6]/NET0131  & ~n48566 ;
  assign n63092 = ~n63086 & ~n63087 ;
  assign n63093 = ~n63091 & n63092 ;
  assign n63097 = ~\P1_P2_EAX_reg[7]/NET0131  & n25847 ;
  assign n63096 = ~\P1_P2_Datao_reg[7]/NET0131  & ~n25847 ;
  assign n63098 = n25918 & ~n63096 ;
  assign n63099 = ~n63097 & n63098 ;
  assign n63094 = \P1_P2_lWord_reg[7]/NET0131  & n25922 ;
  assign n63095 = \P1_P2_Datao_reg[7]/NET0131  & ~n48566 ;
  assign n63100 = ~n63094 & ~n63095 ;
  assign n63101 = ~n63099 & n63100 ;
  assign n63105 = ~\P1_P2_EAX_reg[8]/NET0131  & n25847 ;
  assign n63104 = ~\P1_P2_Datao_reg[8]/NET0131  & ~n25847 ;
  assign n63106 = n25918 & ~n63104 ;
  assign n63107 = ~n63105 & n63106 ;
  assign n63102 = \P1_P2_lWord_reg[8]/NET0131  & n25922 ;
  assign n63103 = \P1_P2_Datao_reg[8]/NET0131  & ~n48566 ;
  assign n63108 = ~n63102 & ~n63103 ;
  assign n63109 = ~n63107 & n63108 ;
  assign n63113 = ~\P1_P2_EAX_reg[9]/NET0131  & n25847 ;
  assign n63112 = ~\P1_P2_Datao_reg[9]/NET0131  & ~n25847 ;
  assign n63114 = n25918 & ~n63112 ;
  assign n63115 = ~n63113 & n63114 ;
  assign n63110 = \P1_P2_lWord_reg[9]/NET0131  & n25922 ;
  assign n63111 = \P1_P2_Datao_reg[9]/NET0131  & ~n48566 ;
  assign n63116 = ~n63110 & ~n63111 ;
  assign n63117 = ~n63115 & n63116 ;
  assign n63121 = ~\P1_P1_EAX_reg[12]/NET0131  & n26162 ;
  assign n63120 = ~\P1_P1_Datao_reg[12]/NET0131  & ~n26162 ;
  assign n63122 = n8355 & ~n63120 ;
  assign n63123 = ~n63121 & n63122 ;
  assign n63118 = \P1_P1_lWord_reg[12]/NET0131  & n27790 ;
  assign n63119 = \P1_P1_Datao_reg[12]/NET0131  & ~n48479 ;
  assign n63124 = ~n63118 & ~n63119 ;
  assign n63125 = ~n63123 & n63124 ;
  assign n63129 = ~\P2_P1_EAX_reg[7]/NET0131  & n26030 ;
  assign n63128 = ~\P2_P1_Datao_reg[7]/NET0131  & ~n26030 ;
  assign n63130 = n11623 & ~n63128 ;
  assign n63131 = ~n63129 & n63130 ;
  assign n63126 = \P2_P1_lWord_reg[7]/NET0131  & n48581 ;
  assign n63127 = \P2_P1_Datao_reg[7]/NET0131  & ~n48594 ;
  assign n63132 = ~n63126 & ~n63127 ;
  assign n63133 = ~n63131 & n63132 ;
  assign n63137 = ~\P1_P1_EAX_reg[15]/NET0131  & n26162 ;
  assign n63136 = ~\P1_P1_Datao_reg[15]/NET0131  & ~n26162 ;
  assign n63138 = n8355 & ~n63136 ;
  assign n63139 = ~n63137 & n63138 ;
  assign n63134 = \P1_P1_lWord_reg[15]/NET0131  & n27790 ;
  assign n63135 = \P1_P1_Datao_reg[15]/NET0131  & ~n48479 ;
  assign n63140 = ~n63134 & ~n63135 ;
  assign n63141 = ~n63139 & n63140 ;
  assign n63145 = ~\P2_P1_EAX_reg[0]/NET0131  & n26030 ;
  assign n63144 = ~\P2_P1_Datao_reg[0]/NET0131  & ~n26030 ;
  assign n63146 = n11623 & ~n63144 ;
  assign n63147 = ~n63145 & n63146 ;
  assign n63142 = \P2_P1_lWord_reg[0]/NET0131  & n48581 ;
  assign n63143 = \P2_P1_Datao_reg[0]/NET0131  & ~n48594 ;
  assign n63148 = ~n63142 & ~n63143 ;
  assign n63149 = ~n63147 & n63148 ;
  assign n63153 = ~\P2_P1_EAX_reg[10]/NET0131  & n26030 ;
  assign n63152 = ~\P2_P1_Datao_reg[10]/NET0131  & ~n26030 ;
  assign n63154 = n11623 & ~n63152 ;
  assign n63155 = ~n63153 & n63154 ;
  assign n63150 = \P2_P1_lWord_reg[10]/NET0131  & n48581 ;
  assign n63151 = \P2_P1_Datao_reg[10]/NET0131  & ~n48594 ;
  assign n63156 = ~n63150 & ~n63151 ;
  assign n63157 = ~n63155 & n63156 ;
  assign n63161 = ~\P2_P1_EAX_reg[11]/NET0131  & n26030 ;
  assign n63160 = ~\P2_P1_Datao_reg[11]/NET0131  & ~n26030 ;
  assign n63162 = n11623 & ~n63160 ;
  assign n63163 = ~n63161 & n63162 ;
  assign n63158 = \P2_P1_lWord_reg[11]/NET0131  & n48581 ;
  assign n63159 = \P2_P1_Datao_reg[11]/NET0131  & ~n48594 ;
  assign n63164 = ~n63158 & ~n63159 ;
  assign n63165 = ~n63163 & n63164 ;
  assign n63169 = ~\P2_P1_EAX_reg[12]/NET0131  & n26030 ;
  assign n63168 = ~\P2_P1_Datao_reg[12]/NET0131  & ~n26030 ;
  assign n63170 = n11623 & ~n63168 ;
  assign n63171 = ~n63169 & n63170 ;
  assign n63166 = \P2_P1_lWord_reg[12]/NET0131  & n48581 ;
  assign n63167 = \P2_P1_Datao_reg[12]/NET0131  & ~n48594 ;
  assign n63172 = ~n63166 & ~n63167 ;
  assign n63173 = ~n63171 & n63172 ;
  assign n63177 = ~\P2_P1_EAX_reg[13]/NET0131  & n26030 ;
  assign n63176 = ~\P2_P1_Datao_reg[13]/NET0131  & ~n26030 ;
  assign n63178 = n11623 & ~n63176 ;
  assign n63179 = ~n63177 & n63178 ;
  assign n63174 = \P2_P1_lWord_reg[13]/NET0131  & n48581 ;
  assign n63175 = \P2_P1_Datao_reg[13]/NET0131  & ~n48594 ;
  assign n63180 = ~n63174 & ~n63175 ;
  assign n63181 = ~n63179 & n63180 ;
  assign n63185 = ~\P2_P1_EAX_reg[14]/NET0131  & n26030 ;
  assign n63184 = ~\P2_P1_Datao_reg[14]/NET0131  & ~n26030 ;
  assign n63186 = n11623 & ~n63184 ;
  assign n63187 = ~n63185 & n63186 ;
  assign n63182 = \P2_P1_lWord_reg[14]/NET0131  & n48581 ;
  assign n63183 = \P2_P1_Datao_reg[14]/NET0131  & ~n48594 ;
  assign n63188 = ~n63182 & ~n63183 ;
  assign n63189 = ~n63187 & n63188 ;
  assign n63193 = ~\P2_P1_EAX_reg[15]/NET0131  & n26030 ;
  assign n63192 = ~\P2_P1_Datao_reg[15]/NET0131  & ~n26030 ;
  assign n63194 = n11623 & ~n63192 ;
  assign n63195 = ~n63193 & n63194 ;
  assign n63190 = \P2_P1_lWord_reg[15]/NET0131  & n48581 ;
  assign n63191 = \P2_P1_Datao_reg[15]/NET0131  & ~n48594 ;
  assign n63196 = ~n63190 & ~n63191 ;
  assign n63197 = ~n63195 & n63196 ;
  assign n63201 = ~\P2_P1_EAX_reg[1]/NET0131  & n26030 ;
  assign n63200 = ~\P2_P1_Datao_reg[1]/NET0131  & ~n26030 ;
  assign n63202 = n11623 & ~n63200 ;
  assign n63203 = ~n63201 & n63202 ;
  assign n63198 = \P2_P1_lWord_reg[1]/NET0131  & n48581 ;
  assign n63199 = \P2_P1_Datao_reg[1]/NET0131  & ~n48594 ;
  assign n63204 = ~n63198 & ~n63199 ;
  assign n63205 = ~n63203 & n63204 ;
  assign n63209 = ~\P2_P1_EAX_reg[2]/NET0131  & n26030 ;
  assign n63208 = ~\P2_P1_Datao_reg[2]/NET0131  & ~n26030 ;
  assign n63210 = n11623 & ~n63208 ;
  assign n63211 = ~n63209 & n63210 ;
  assign n63206 = \P2_P1_lWord_reg[2]/NET0131  & n48581 ;
  assign n63207 = \P2_P1_Datao_reg[2]/NET0131  & ~n48594 ;
  assign n63212 = ~n63206 & ~n63207 ;
  assign n63213 = ~n63211 & n63212 ;
  assign n63217 = ~\P2_P1_EAX_reg[3]/NET0131  & n26030 ;
  assign n63216 = ~\P2_P1_Datao_reg[3]/NET0131  & ~n26030 ;
  assign n63218 = n11623 & ~n63216 ;
  assign n63219 = ~n63217 & n63218 ;
  assign n63214 = \P2_P1_lWord_reg[3]/NET0131  & n48581 ;
  assign n63215 = \P2_P1_Datao_reg[3]/NET0131  & ~n48594 ;
  assign n63220 = ~n63214 & ~n63215 ;
  assign n63221 = ~n63219 & n63220 ;
  assign n63225 = ~\P2_P1_EAX_reg[4]/NET0131  & n26030 ;
  assign n63224 = ~\P2_P1_Datao_reg[4]/NET0131  & ~n26030 ;
  assign n63226 = n11623 & ~n63224 ;
  assign n63227 = ~n63225 & n63226 ;
  assign n63222 = \P2_P1_lWord_reg[4]/NET0131  & n48581 ;
  assign n63223 = \P2_P1_Datao_reg[4]/NET0131  & ~n48594 ;
  assign n63228 = ~n63222 & ~n63223 ;
  assign n63229 = ~n63227 & n63228 ;
  assign n63233 = ~\P2_P1_EAX_reg[5]/NET0131  & n26030 ;
  assign n63232 = ~\P2_P1_Datao_reg[5]/NET0131  & ~n26030 ;
  assign n63234 = n11623 & ~n63232 ;
  assign n63235 = ~n63233 & n63234 ;
  assign n63230 = \P2_P1_lWord_reg[5]/NET0131  & n48581 ;
  assign n63231 = \P2_P1_Datao_reg[5]/NET0131  & ~n48594 ;
  assign n63236 = ~n63230 & ~n63231 ;
  assign n63237 = ~n63235 & n63236 ;
  assign n63241 = ~\P2_P1_EAX_reg[6]/NET0131  & n26030 ;
  assign n63240 = ~\P2_P1_Datao_reg[6]/NET0131  & ~n26030 ;
  assign n63242 = n11623 & ~n63240 ;
  assign n63243 = ~n63241 & n63242 ;
  assign n63238 = \P2_P1_lWord_reg[6]/NET0131  & n48581 ;
  assign n63239 = \P2_P1_Datao_reg[6]/NET0131  & ~n48594 ;
  assign n63244 = ~n63238 & ~n63239 ;
  assign n63245 = ~n63243 & n63244 ;
  assign n63249 = ~\P2_P1_EAX_reg[8]/NET0131  & n26030 ;
  assign n63248 = ~\P2_P1_Datao_reg[8]/NET0131  & ~n26030 ;
  assign n63250 = n11623 & ~n63248 ;
  assign n63251 = ~n63249 & n63250 ;
  assign n63246 = \P2_P1_lWord_reg[8]/NET0131  & n48581 ;
  assign n63247 = \P2_P1_Datao_reg[8]/NET0131  & ~n48594 ;
  assign n63252 = ~n63246 & ~n63247 ;
  assign n63253 = ~n63251 & n63252 ;
  assign n63257 = ~\P2_P1_EAX_reg[9]/NET0131  & n26030 ;
  assign n63256 = ~\P2_P1_Datao_reg[9]/NET0131  & ~n26030 ;
  assign n63258 = n11623 & ~n63256 ;
  assign n63259 = ~n63257 & n63258 ;
  assign n63254 = \P2_P1_lWord_reg[9]/NET0131  & n48581 ;
  assign n63255 = \P2_P1_Datao_reg[9]/NET0131  & ~n48594 ;
  assign n63260 = ~n63254 & ~n63255 ;
  assign n63261 = ~n63259 & n63260 ;
  assign n63265 = ~\P1_P1_EAX_reg[10]/NET0131  & n26162 ;
  assign n63264 = ~\P1_P1_Datao_reg[10]/NET0131  & ~n26162 ;
  assign n63266 = n8355 & ~n63264 ;
  assign n63267 = ~n63265 & n63266 ;
  assign n63262 = \P1_P1_lWord_reg[10]/NET0131  & n27790 ;
  assign n63263 = \P1_P1_Datao_reg[10]/NET0131  & ~n48479 ;
  assign n63268 = ~n63262 & ~n63263 ;
  assign n63269 = ~n63267 & n63268 ;
  assign n63273 = ~\P1_P1_EAX_reg[0]/NET0131  & n26162 ;
  assign n63272 = ~\P1_P1_Datao_reg[0]/NET0131  & ~n26162 ;
  assign n63274 = n8355 & ~n63272 ;
  assign n63275 = ~n63273 & n63274 ;
  assign n63270 = \P1_P1_lWord_reg[0]/NET0131  & n27790 ;
  assign n63271 = \P1_P1_Datao_reg[0]/NET0131  & ~n48479 ;
  assign n63276 = ~n63270 & ~n63271 ;
  assign n63277 = ~n63275 & n63276 ;
  assign n63281 = ~\P1_P1_EAX_reg[11]/NET0131  & n26162 ;
  assign n63280 = ~\P1_P1_Datao_reg[11]/NET0131  & ~n26162 ;
  assign n63282 = n8355 & ~n63280 ;
  assign n63283 = ~n63281 & n63282 ;
  assign n63278 = \P1_P1_lWord_reg[11]/NET0131  & n27790 ;
  assign n63279 = \P1_P1_Datao_reg[11]/NET0131  & ~n48479 ;
  assign n63284 = ~n63278 & ~n63279 ;
  assign n63285 = ~n63283 & n63284 ;
  assign n63290 = ~n11919 & n27681 ;
  assign n63293 = ~n11861 & n63290 ;
  assign n63294 = ~n36674 & ~n63293 ;
  assign n63286 = ~\P2_P1_InstQueueWr_Addr_reg[3]/NET0131  & ~n11872 ;
  assign n63287 = ~n11873 & ~n63286 ;
  assign n63295 = ~n11864 & ~n63287 ;
  assign n63296 = ~n11865 & ~n63295 ;
  assign n63297 = ~n63294 & n63296 ;
  assign n63289 = \P2_P1_InstQueueWr_Addr_reg[3]/NET0131  & ~n62190 ;
  assign n63288 = n11692 & n63287 ;
  assign n63291 = ~n11918 & ~n12131 ;
  assign n63292 = n63290 & ~n63291 ;
  assign n63298 = ~n63288 & ~n63292 ;
  assign n63299 = ~n63289 & n63298 ;
  assign n63300 = ~n63297 & n63299 ;
  assign n63305 = n26800 & ~n28438 ;
  assign n63308 = ~n28397 & n63305 ;
  assign n63309 = n36760 & ~n63308 ;
  assign n63301 = ~\P2_P2_InstQueueWr_Addr_reg[3]/NET0131  & ~n28386 ;
  assign n63302 = ~n28387 & ~n63301 ;
  assign n63310 = ~n28400 & ~n63302 ;
  assign n63311 = ~n28401 & ~n63310 ;
  assign n63312 = ~n63309 & n63311 ;
  assign n63304 = \P2_P2_InstQueueWr_Addr_reg[3]/NET0131  & ~n62207 ;
  assign n63303 = n27613 & n63302 ;
  assign n63306 = ~n28437 & ~n28610 ;
  assign n63307 = n63305 & ~n63306 ;
  assign n63313 = ~n63303 & ~n63307 ;
  assign n63314 = ~n63304 & n63313 ;
  assign n63315 = ~n63312 & n63314 ;
  assign n63316 = \P2_P1_InstQueueWr_Addr_reg[1]/NET0131  & ~n62189 ;
  assign n63317 = ~\P2_P1_InstQueueWr_Addr_reg[0]/NET0131  & n11692 ;
  assign n63318 = \P2_P1_InstQueueWr_Addr_reg[1]/NET0131  & n52907 ;
  assign n63319 = ~n27681 & n63318 ;
  assign n63320 = ~n63317 & n63319 ;
  assign n63321 = \P2_P1_InstQueueWr_Addr_reg[0]/NET0131  & n11692 ;
  assign n63322 = ~\P2_P1_InstQueueWr_Addr_reg[1]/NET0131  & ~n63321 ;
  assign n63323 = ~n36674 & n63322 ;
  assign n63324 = ~n63320 & ~n63323 ;
  assign n63325 = ~n63316 & ~n63324 ;
  assign n63326 = \P2_P2_InstQueueWr_Addr_reg[1]/NET0131  & ~n62206 ;
  assign n63327 = ~\P2_P2_InstQueueWr_Addr_reg[0]/NET0131  & n27613 ;
  assign n63328 = \P2_P2_InstQueueWr_Addr_reg[1]/NET0131  & n52964 ;
  assign n63329 = ~n26800 & n63328 ;
  assign n63330 = ~n63327 & n63329 ;
  assign n63331 = \P2_P2_InstQueueWr_Addr_reg[0]/NET0131  & n27613 ;
  assign n63332 = ~\P2_P2_InstQueueWr_Addr_reg[1]/NET0131  & ~n63331 ;
  assign n63333 = n36760 & n63332 ;
  assign n63334 = ~n63330 & ~n63333 ;
  assign n63335 = ~n63326 & ~n63334 ;
  assign n63338 = ~n11623 & n43231 ;
  assign n63339 = \P2_P1_InstQueueWr_Addr_reg[0]/NET0131  & ~n63338 ;
  assign n63336 = ~\P2_P1_Flush_reg/NET0131  & ~\P2_P1_InstQueueWr_Addr_reg[0]/NET0131  ;
  assign n63337 = n27486 & ~n63336 ;
  assign n63340 = ~n63317 & ~n63337 ;
  assign n63341 = ~n63339 & n63340 ;
  assign n63344 = ~n27977 & n45045 ;
  assign n63345 = n62205 & n63344 ;
  assign n63346 = \P2_P2_InstQueueWr_Addr_reg[0]/NET0131  & ~n63345 ;
  assign n63342 = ~\P2_P2_Flush_reg/NET0131  & ~\P2_P2_InstQueueWr_Addr_reg[0]/NET0131  ;
  assign n63343 = n27642 & ~n63342 ;
  assign n63347 = ~n63327 & ~n63343 ;
  assign n63348 = ~n63346 & n63347 ;
  assign n63350 = ~\P2_P2_rEIP_reg[0]/NET0131  & ~\P2_P2_rEIP_reg[1]/NET0131  ;
  assign n63351 = \P2_P2_rEIP_reg[31]/NET0131  & ~n63350 ;
  assign n63352 = \P2_P2_rEIP_reg[2]/NET0131  & n63351 ;
  assign n63353 = \P2_P2_rEIP_reg[3]/NET0131  & n63352 ;
  assign n63354 = \P2_P2_rEIP_reg[4]/NET0131  & n63353 ;
  assign n63355 = \P2_P2_rEIP_reg[5]/NET0131  & n63354 ;
  assign n63356 = \P2_P2_rEIP_reg[6]/NET0131  & n63355 ;
  assign n63357 = \P2_P2_rEIP_reg[7]/NET0131  & n63356 ;
  assign n63358 = \P2_P2_rEIP_reg[8]/NET0131  & n63357 ;
  assign n63359 = n52307 & n63358 ;
  assign n63360 = \P2_P2_rEIP_reg[26]/NET0131  & n63359 ;
  assign n63361 = \P2_P2_rEIP_reg[27]/NET0131  & n63360 ;
  assign n63362 = \P2_P2_rEIP_reg[28]/NET0131  & n63361 ;
  assign n63363 = \P2_P2_rEIP_reg[29]/NET0131  & n63362 ;
  assign n63365 = \P2_P2_rEIP_reg[30]/NET0131  & n63363 ;
  assign n63364 = ~\P2_P2_rEIP_reg[30]/NET0131  & ~n63363 ;
  assign n63366 = n26647 & ~n63364 ;
  assign n63367 = ~n63365 & n63366 ;
  assign n63349 = \P2_P2_Address_reg[28]/NET0131  & ~n26646 ;
  assign n63368 = \P2_P2_rEIP_reg[0]/NET0131  & \P2_P2_rEIP_reg[31]/NET0131  ;
  assign n63369 = n52343 & n63368 ;
  assign n63370 = \P2_P2_rEIP_reg[27]/NET0131  & n63369 ;
  assign n63371 = \P2_P2_rEIP_reg[28]/NET0131  & n63370 ;
  assign n63374 = \P2_P2_rEIP_reg[29]/NET0131  & n63371 ;
  assign n63372 = ~\P2_P2_rEIP_reg[29]/NET0131  & ~n63371 ;
  assign n63373 = \P2_P2_State_reg[2]/NET0131  & n26646 ;
  assign n63375 = ~n63372 & n63373 ;
  assign n63376 = ~n63374 & n63375 ;
  assign n63377 = ~n63349 & ~n63376 ;
  assign n63378 = ~n63367 & n63377 ;
  assign n63380 = ~\P1_P1_rEIP_reg[0]/NET0131  & ~\P1_P1_rEIP_reg[1]/NET0131  ;
  assign n63381 = \P1_P1_rEIP_reg[31]/NET0131  & ~n63380 ;
  assign n63382 = \P1_P1_rEIP_reg[2]/NET0131  & n63381 ;
  assign n63383 = \P1_P1_rEIP_reg[3]/NET0131  & n63382 ;
  assign n63384 = \P1_P1_rEIP_reg[4]/NET0131  & n63383 ;
  assign n63385 = \P1_P1_rEIP_reg[5]/NET0131  & n63384 ;
  assign n63386 = \P1_P1_rEIP_reg[6]/NET0131  & n63385 ;
  assign n63387 = \P1_P1_rEIP_reg[7]/NET0131  & n63386 ;
  assign n63388 = \P1_P1_rEIP_reg[8]/NET0131  & n63387 ;
  assign n63389 = \P1_P1_rEIP_reg[9]/NET0131  & n63388 ;
  assign n63390 = \P1_P1_rEIP_reg[10]/NET0131  & n63389 ;
  assign n63391 = \P1_P1_rEIP_reg[11]/NET0131  & n63390 ;
  assign n63392 = n51667 & n63391 ;
  assign n63393 = \P1_P1_rEIP_reg[14]/NET0131  & n63392 ;
  assign n63394 = n51845 & n63393 ;
  assign n63395 = n51950 & n63394 ;
  assign n63396 = n52021 & n63395 ;
  assign n63398 = \P1_P1_rEIP_reg[30]/NET0131  & n63396 ;
  assign n63397 = ~\P1_P1_rEIP_reg[30]/NET0131  & ~n63396 ;
  assign n63399 = n26155 & ~n63397 ;
  assign n63400 = ~n63398 & n63399 ;
  assign n63379 = \P1_P1_Address_reg[28]/NET0131  & ~n26154 ;
  assign n63402 = \P1_P1_rEIP_reg[0]/NET0131  & \P1_P1_rEIP_reg[31]/NET0131  ;
  assign n63411 = n51847 & n63402 ;
  assign n63412 = \P1_P1_rEIP_reg[25]/NET0131  & n63411 ;
  assign n63413 = \P1_P1_rEIP_reg[26]/NET0131  & n63412 ;
  assign n63414 = n52021 & n63413 ;
  assign n63401 = \P1_P1_State_reg[2]/NET0131  & n26154 ;
  assign n63403 = n51674 & n63402 ;
  assign n63404 = \P1_P1_rEIP_reg[11]/NET0131  & n63403 ;
  assign n63405 = n51667 & n63404 ;
  assign n63406 = \P1_P1_rEIP_reg[14]/NET0131  & n63405 ;
  assign n63407 = n51845 & n63406 ;
  assign n63408 = n51951 & n63407 ;
  assign n63409 = \P1_P1_rEIP_reg[28]/NET0131  & n63408 ;
  assign n63410 = ~\P1_P1_rEIP_reg[29]/NET0131  & ~n63409 ;
  assign n63415 = n63401 & ~n63410 ;
  assign n63416 = ~n63414 & n63415 ;
  assign n63417 = ~n63379 & ~n63416 ;
  assign n63418 = ~n63400 & n63417 ;
  assign n63427 = ~\P1_P2_rEIP_reg[0]/NET0131  & ~\P1_P2_rEIP_reg[1]/NET0131  ;
  assign n63428 = \P1_P2_rEIP_reg[31]/NET0131  & ~n63427 ;
  assign n63429 = \P1_P2_rEIP_reg[2]/NET0131  & n63428 ;
  assign n63430 = \P1_P2_rEIP_reg[3]/NET0131  & n63429 ;
  assign n63431 = \P1_P2_rEIP_reg[4]/NET0131  & n63430 ;
  assign n63432 = \P1_P2_rEIP_reg[5]/NET0131  & n63431 ;
  assign n63433 = \P1_P2_rEIP_reg[6]/NET0131  & n63432 ;
  assign n63434 = \P1_P2_rEIP_reg[7]/NET0131  & n63433 ;
  assign n63435 = \P1_P2_rEIP_reg[8]/NET0131  & n63434 ;
  assign n63436 = n48395 & n63435 ;
  assign n63437 = n48377 & n63436 ;
  assign n63438 = \P1_P2_rEIP_reg[21]/NET0131  & n63437 ;
  assign n63439 = \P1_P2_rEIP_reg[22]/NET0131  & n63438 ;
  assign n63440 = n48375 & n63439 ;
  assign n63441 = \P1_P2_rEIP_reg[26]/NET0131  & n63440 ;
  assign n63442 = \P1_P2_rEIP_reg[27]/NET0131  & n63441 ;
  assign n63443 = n48400 & n63442 ;
  assign n63445 = \P1_P2_rEIP_reg[30]/NET0131  & n63443 ;
  assign n63444 = ~\P1_P2_rEIP_reg[30]/NET0131  & ~n63443 ;
  assign n63446 = n25765 & ~n63444 ;
  assign n63447 = ~n63445 & n63446 ;
  assign n63419 = \P1_P2_Address_reg[28]/NET0131  & ~n25764 ;
  assign n63421 = \P1_P2_rEIP_reg[0]/NET0131  & \P1_P2_rEIP_reg[31]/NET0131  ;
  assign n63422 = n51560 & n63421 ;
  assign n63424 = \P1_P2_rEIP_reg[29]/NET0131  & n63422 ;
  assign n63420 = \P1_P2_State_reg[2]/NET0131  & n25764 ;
  assign n63423 = ~\P1_P2_rEIP_reg[29]/NET0131  & ~n63422 ;
  assign n63425 = n63420 & ~n63423 ;
  assign n63426 = ~n63424 & n63425 ;
  assign n63448 = ~n63419 & ~n63426 ;
  assign n63449 = ~n63447 & n63448 ;
  assign n63475 = \P2_P1_rEIP_reg[0]/NET0131  & \P2_P1_rEIP_reg[31]/NET0131  ;
  assign n63476 = n51010 & n63475 ;
  assign n63477 = \P2_P1_rEIP_reg[26]/NET0131  & n63476 ;
  assign n63478 = n51080 & n63477 ;
  assign n63481 = \P2_P1_rEIP_reg[29]/NET0131  & n63478 ;
  assign n63479 = ~\P2_P1_rEIP_reg[29]/NET0131  & ~n63478 ;
  assign n63480 = \P2_P1_State_reg[2]/NET0131  & n25954 ;
  assign n63482 = ~n63479 & n63480 ;
  assign n63483 = ~n63481 & n63482 ;
  assign n63450 = \P2_P1_Address_reg[28]/NET0131  & ~n25954 ;
  assign n63451 = ~\P2_P1_rEIP_reg[0]/NET0131  & ~\P2_P1_rEIP_reg[1]/NET0131  ;
  assign n63452 = \P2_P1_rEIP_reg[31]/NET0131  & ~n63451 ;
  assign n63453 = \P2_P1_rEIP_reg[2]/NET0131  & n63452 ;
  assign n63454 = \P2_P1_rEIP_reg[3]/NET0131  & n63453 ;
  assign n63455 = \P2_P1_rEIP_reg[4]/NET0131  & n63454 ;
  assign n63456 = \P2_P1_rEIP_reg[5]/NET0131  & n63455 ;
  assign n63457 = \P2_P1_rEIP_reg[6]/NET0131  & n63456 ;
  assign n63458 = \P2_P1_rEIP_reg[7]/NET0131  & n63457 ;
  assign n63459 = \P2_P1_rEIP_reg[8]/NET0131  & n63458 ;
  assign n63460 = \P2_P1_rEIP_reg[9]/NET0131  & n63459 ;
  assign n63461 = n50772 & n63460 ;
  assign n63462 = n50966 & n63461 ;
  assign n63463 = n50764 & n63462 ;
  assign n63464 = n50781 & n63463 ;
  assign n63465 = n50965 & n63464 ;
  assign n63466 = n51009 & n63465 ;
  assign n63467 = \P2_P1_rEIP_reg[26]/NET0131  & n63466 ;
  assign n63468 = \P2_P1_rEIP_reg[27]/NET0131  & n63467 ;
  assign n63469 = \P2_P1_rEIP_reg[28]/NET0131  & n63468 ;
  assign n63470 = \P2_P1_rEIP_reg[29]/NET0131  & n63469 ;
  assign n63472 = \P2_P1_rEIP_reg[30]/NET0131  & n63470 ;
  assign n63471 = ~\P2_P1_rEIP_reg[30]/NET0131  & ~n63470 ;
  assign n63473 = n25955 & ~n63471 ;
  assign n63474 = ~n63472 & n63473 ;
  assign n63484 = ~n63450 & ~n63474 ;
  assign n63485 = ~n63483 & n63484 ;
  assign n63486 = ~\P1_P1_Flush_reg/NET0131  & n27623 ;
  assign n63487 = ~n8355 & ~n8361 ;
  assign n63488 = ~n27790 & n63487 ;
  assign n63489 = ~n63486 & n63488 ;
  assign n63490 = n52935 & n63489 ;
  assign n63491 = \P1_P1_InstQueueWr_Addr_reg[2]/NET0131  & ~n63490 ;
  assign n63493 = \P1_P1_DataWidth_reg[1]/NET0131  & \P1_P1_InstQueueWr_Addr_reg[2]/NET0131  ;
  assign n63494 = ~n8287 & n63493 ;
  assign n63492 = ~n8282 & ~n8287 ;
  assign n63495 = ~n8371 & ~n63492 ;
  assign n63496 = ~n63494 & n63495 ;
  assign n63497 = ~n8350 & ~n63496 ;
  assign n63498 = n8143 & ~n63492 ;
  assign n63499 = ~\P1_P1_InstQueueWr_Addr_reg[2]/NET0131  & ~n8140 ;
  assign n63500 = ~n27791 & n63499 ;
  assign n63501 = ~n63498 & n63500 ;
  assign n63502 = ~n8377 & ~n63501 ;
  assign n63503 = ~n63497 & n63502 ;
  assign n63504 = ~n63491 & ~n63503 ;
  assign n63505 = ~\P1_P2_Flush_reg/NET0131  & n27673 ;
  assign n63506 = ~n25918 & ~n25922 ;
  assign n63507 = ~n27675 & n63506 ;
  assign n63508 = ~n63505 & n63507 ;
  assign n63509 = n52882 & n63508 ;
  assign n63510 = \P1_P2_InstQueueWr_Addr_reg[2]/NET0131  & ~n63509 ;
  assign n63511 = ~n27902 & ~n36629 ;
  assign n63512 = \P1_P2_InstQueueWr_Addr_reg[2]/NET0131  & ~n63511 ;
  assign n63513 = ~n28928 & ~n63512 ;
  assign n63514 = ~n27608 & ~n63513 ;
  assign n63515 = n27902 & ~n28928 ;
  assign n63516 = ~\P1_P2_InstQueueWr_Addr_reg[2]/NET0131  & ~n27899 ;
  assign n63517 = ~n25933 & n63516 ;
  assign n63518 = ~n63515 & n63517 ;
  assign n63519 = ~n28056 & ~n63518 ;
  assign n63520 = ~n63514 & n63519 ;
  assign n63521 = ~n63510 & ~n63520 ;
  assign n63522 = ~\P1_P3_Flush_reg/NET0131  & n10041 ;
  assign n63523 = ~n9241 & n43257 ;
  assign n63524 = ~n63522 & n63523 ;
  assign n63525 = ~n21771 & n63524 ;
  assign n63526 = \P1_P3_InstQueueWr_Addr_reg[2]/NET0131  & ~n63525 ;
  assign n63528 = \P1_P3_DataWidth_reg[1]/NET0131  & \P1_P3_InstQueueWr_Addr_reg[2]/NET0131  ;
  assign n63529 = ~n16492 & n63528 ;
  assign n63527 = ~n9245 & ~n16492 ;
  assign n63530 = ~n49741 & ~n63527 ;
  assign n63531 = ~n63529 & n63530 ;
  assign n63532 = ~n10046 & ~n63531 ;
  assign n63533 = n49740 & ~n63527 ;
  assign n63534 = ~\P1_P3_InstQueueWr_Addr_reg[2]/NET0131  & ~n49733 ;
  assign n63535 = ~n11698 & n63534 ;
  assign n63536 = ~n63533 & n63535 ;
  assign n63537 = ~n49734 & ~n63536 ;
  assign n63538 = ~n63532 & n63537 ;
  assign n63539 = ~n63526 & ~n63538 ;
  assign n63542 = n8860 & n49732 ;
  assign n63541 = ~\P1_P3_InstQueue_reg[0][5]/NET0131  & ~n49732 ;
  assign n63543 = n10046 & ~n63541 ;
  assign n63544 = ~n63542 & n63543 ;
  assign n63540 = \P1_P3_InstQueue_reg[0][5]/NET0131  & ~n49750 ;
  assign n63545 = \P1_buf2_reg[29]/NET0131  & n49739 ;
  assign n63546 = \P1_buf2_reg[21]/NET0131  & ~n49739 ;
  assign n63547 = n49742 & n63546 ;
  assign n63548 = ~n63545 & ~n63547 ;
  assign n63549 = n11698 & ~n63548 ;
  assign n63550 = \P1_buf2_reg[5]/NET0131  & n49760 ;
  assign n63551 = ~n63549 & ~n63550 ;
  assign n63552 = ~n63540 & n63551 ;
  assign n63553 = ~n63544 & n63552 ;
  assign n63556 = n8860 & n49766 ;
  assign n63555 = ~\P1_P3_InstQueue_reg[10][5]/NET0131  & ~n49766 ;
  assign n63557 = n10046 & ~n63555 ;
  assign n63558 = ~n63556 & n63557 ;
  assign n63554 = \P1_P3_InstQueue_reg[10][5]/NET0131  & ~n49776 ;
  assign n63559 = \P1_buf2_reg[29]/NET0131  & n49770 ;
  assign n63560 = \P1_buf2_reg[21]/NET0131  & n49771 ;
  assign n63561 = ~n63559 & ~n63560 ;
  assign n63562 = n11698 & ~n63561 ;
  assign n63563 = \P1_buf2_reg[5]/NET0131  & n49786 ;
  assign n63564 = ~n63562 & ~n63563 ;
  assign n63565 = ~n63554 & n63564 ;
  assign n63566 = ~n63558 & n63565 ;
  assign n63569 = n8860 & n49792 ;
  assign n63568 = ~\P1_P3_InstQueue_reg[11][5]/NET0131  & ~n49792 ;
  assign n63570 = n10046 & ~n63568 ;
  assign n63571 = ~n63569 & n63570 ;
  assign n63567 = \P1_P3_InstQueue_reg[11][5]/NET0131  & ~n49798 ;
  assign n63572 = \P1_buf2_reg[29]/NET0131  & n49771 ;
  assign n63573 = \P1_buf2_reg[21]/NET0131  & n49768 ;
  assign n63574 = ~n63572 & ~n63573 ;
  assign n63575 = n11698 & ~n63574 ;
  assign n63576 = \P1_buf2_reg[5]/NET0131  & n49808 ;
  assign n63577 = ~n63575 & ~n63576 ;
  assign n63578 = ~n63567 & n63577 ;
  assign n63579 = ~n63571 & n63578 ;
  assign n63582 = n8860 & n49814 ;
  assign n63581 = ~\P1_P3_InstQueue_reg[12][5]/NET0131  & ~n49814 ;
  assign n63583 = n10046 & ~n63581 ;
  assign n63584 = ~n63582 & n63583 ;
  assign n63580 = \P1_P3_InstQueue_reg[12][5]/NET0131  & ~n49819 ;
  assign n63585 = \P1_buf2_reg[29]/NET0131  & n49768 ;
  assign n63586 = \P1_buf2_reg[21]/NET0131  & n49766 ;
  assign n63587 = ~n63585 & ~n63586 ;
  assign n63588 = n11698 & ~n63587 ;
  assign n63589 = \P1_buf2_reg[5]/NET0131  & n49829 ;
  assign n63590 = ~n63588 & ~n63589 ;
  assign n63591 = ~n63580 & n63590 ;
  assign n63592 = ~n63584 & n63591 ;
  assign n63595 = n8860 & n49739 ;
  assign n63594 = ~\P1_P3_InstQueue_reg[13][5]/NET0131  & ~n49739 ;
  assign n63596 = n10046 & ~n63594 ;
  assign n63597 = ~n63595 & n63596 ;
  assign n63593 = \P1_P3_InstQueue_reg[13][5]/NET0131  & ~n49838 ;
  assign n63598 = \P1_buf2_reg[29]/NET0131  & n49766 ;
  assign n63599 = \P1_buf2_reg[21]/NET0131  & ~n49766 ;
  assign n63600 = n49792 & n63599 ;
  assign n63601 = ~n63598 & ~n63600 ;
  assign n63602 = n11698 & ~n63601 ;
  assign n63603 = \P1_buf2_reg[5]/NET0131  & n49848 ;
  assign n63604 = ~n63602 & ~n63603 ;
  assign n63605 = ~n63593 & n63604 ;
  assign n63606 = ~n63597 & n63605 ;
  assign n63609 = n8860 & n49742 ;
  assign n63608 = ~\P1_P3_InstQueue_reg[14][5]/NET0131  & ~n49742 ;
  assign n63610 = n10046 & ~n63608 ;
  assign n63611 = ~n63609 & n63610 ;
  assign n63607 = \P1_P3_InstQueue_reg[14][5]/NET0131  & ~n49856 ;
  assign n63612 = \P1_buf2_reg[29]/NET0131  & n49792 ;
  assign n63613 = \P1_buf2_reg[21]/NET0131  & ~n49792 ;
  assign n63614 = n49814 & n63613 ;
  assign n63615 = ~n63612 & ~n63614 ;
  assign n63616 = n11698 & ~n63615 ;
  assign n63617 = \P1_buf2_reg[5]/NET0131  & n49866 ;
  assign n63618 = ~n63616 & ~n63617 ;
  assign n63619 = ~n63607 & n63618 ;
  assign n63620 = ~n63611 & n63619 ;
  assign n63623 = n8860 & n49735 ;
  assign n63622 = ~\P1_P3_InstQueue_reg[15][5]/NET0131  & ~n49735 ;
  assign n63624 = n10046 & ~n63622 ;
  assign n63625 = ~n63623 & n63624 ;
  assign n63621 = \P1_P3_InstQueue_reg[15][5]/NET0131  & ~n49875 ;
  assign n63626 = \P1_buf2_reg[29]/NET0131  & n49814 ;
  assign n63627 = \P1_buf2_reg[21]/NET0131  & n49739 ;
  assign n63628 = ~n63626 & ~n63627 ;
  assign n63629 = n11698 & ~n63628 ;
  assign n63630 = \P1_buf2_reg[5]/NET0131  & n49885 ;
  assign n63631 = ~n63629 & ~n63630 ;
  assign n63632 = ~n63621 & n63631 ;
  assign n63633 = ~n63625 & n63632 ;
  assign n63636 = n8860 & n49890 ;
  assign n63635 = ~\P1_P3_InstQueue_reg[1][5]/NET0131  & ~n49890 ;
  assign n63637 = n10046 & ~n63635 ;
  assign n63638 = ~n63636 & n63637 ;
  assign n63634 = \P1_P3_InstQueue_reg[1][5]/NET0131  & ~n49895 ;
  assign n63639 = \P1_buf2_reg[29]/NET0131  & n49742 ;
  assign n63640 = \P1_buf2_reg[21]/NET0131  & n49735 ;
  assign n63641 = ~n63639 & ~n63640 ;
  assign n63642 = n11698 & ~n63641 ;
  assign n63643 = \P1_buf2_reg[5]/NET0131  & n49905 ;
  assign n63644 = ~n63642 & ~n63643 ;
  assign n63645 = ~n63634 & n63644 ;
  assign n63646 = ~n63638 & n63645 ;
  assign n63649 = n8860 & n49910 ;
  assign n63648 = ~\P1_P3_InstQueue_reg[2][5]/NET0131  & ~n49910 ;
  assign n63650 = n10046 & ~n63648 ;
  assign n63651 = ~n63649 & n63650 ;
  assign n63647 = \P1_P3_InstQueue_reg[2][5]/NET0131  & ~n49915 ;
  assign n63652 = \P1_buf2_reg[29]/NET0131  & n49735 ;
  assign n63653 = \P1_buf2_reg[21]/NET0131  & n49732 ;
  assign n63654 = ~n63652 & ~n63653 ;
  assign n63655 = n11698 & ~n63654 ;
  assign n63656 = \P1_buf2_reg[5]/NET0131  & n49925 ;
  assign n63657 = ~n63655 & ~n63656 ;
  assign n63658 = ~n63647 & n63657 ;
  assign n63659 = ~n63651 & n63658 ;
  assign n63662 = n8860 & n49930 ;
  assign n63661 = ~\P1_P3_InstQueue_reg[3][5]/NET0131  & ~n49930 ;
  assign n63663 = n10046 & ~n63661 ;
  assign n63664 = ~n63662 & n63663 ;
  assign n63660 = \P1_P3_InstQueue_reg[3][5]/NET0131  & ~n49935 ;
  assign n63665 = \P1_buf2_reg[29]/NET0131  & n49732 ;
  assign n63666 = \P1_buf2_reg[21]/NET0131  & ~n49732 ;
  assign n63667 = n49890 & n63666 ;
  assign n63668 = ~n63665 & ~n63667 ;
  assign n63669 = n11698 & ~n63668 ;
  assign n63670 = \P1_buf2_reg[5]/NET0131  & n49945 ;
  assign n63671 = ~n63669 & ~n63670 ;
  assign n63672 = ~n63660 & n63671 ;
  assign n63673 = ~n63664 & n63672 ;
  assign n63676 = n8860 & n49950 ;
  assign n63675 = ~\P1_P3_InstQueue_reg[4][5]/NET0131  & ~n49950 ;
  assign n63677 = n10046 & ~n63675 ;
  assign n63678 = ~n63676 & n63677 ;
  assign n63674 = \P1_P3_InstQueue_reg[4][5]/NET0131  & ~n49955 ;
  assign n63679 = \P1_buf2_reg[29]/NET0131  & n49890 ;
  assign n63680 = \P1_buf2_reg[21]/NET0131  & ~n49890 ;
  assign n63681 = n49910 & n63680 ;
  assign n63682 = ~n63679 & ~n63681 ;
  assign n63683 = n11698 & ~n63682 ;
  assign n63684 = \P1_buf2_reg[5]/NET0131  & n49965 ;
  assign n63685 = ~n63683 & ~n63684 ;
  assign n63686 = ~n63674 & n63685 ;
  assign n63687 = ~n63678 & n63686 ;
  assign n63690 = n8860 & n49970 ;
  assign n63689 = ~\P1_P3_InstQueue_reg[5][5]/NET0131  & ~n49970 ;
  assign n63691 = n10046 & ~n63689 ;
  assign n63692 = ~n63690 & n63691 ;
  assign n63688 = \P1_P3_InstQueue_reg[5][5]/NET0131  & ~n49975 ;
  assign n63693 = \P1_buf2_reg[29]/NET0131  & n49910 ;
  assign n63694 = \P1_buf2_reg[21]/NET0131  & ~n49910 ;
  assign n63695 = n49930 & n63694 ;
  assign n63696 = ~n63693 & ~n63695 ;
  assign n63697 = n11698 & ~n63696 ;
  assign n63698 = \P1_buf2_reg[5]/NET0131  & n49985 ;
  assign n63699 = ~n63697 & ~n63698 ;
  assign n63700 = ~n63688 & n63699 ;
  assign n63701 = ~n63692 & n63700 ;
  assign n63702 = ~\P2_P3_Flush_reg/NET0131  & n27661 ;
  assign n63703 = ~n27308 & ~n27651 ;
  assign n63704 = ~n48523 & n63703 ;
  assign n63705 = ~n63702 & n63704 ;
  assign n63706 = n52996 & n63705 ;
  assign n63707 = \P2_P3_InstQueueWr_Addr_reg[2]/NET0131  & ~n63706 ;
  assign n63708 = ~n27315 & ~n32867 ;
  assign n63714 = n50013 & ~n63708 ;
  assign n63715 = ~\P2_P3_InstQueueWr_Addr_reg[2]/NET0131  & ~n50022 ;
  assign n63716 = ~n27325 & n63715 ;
  assign n63717 = ~n63714 & n63716 ;
  assign n63709 = \P2_P3_DataWidth_reg[1]/NET0131  & \P2_P3_InstQueueWr_Addr_reg[2]/NET0131  ;
  assign n63710 = ~n32867 & n63709 ;
  assign n63711 = ~n50014 & ~n63710 ;
  assign n63712 = ~n63708 & n63711 ;
  assign n63713 = ~n27788 & ~n63712 ;
  assign n63718 = ~n50023 & ~n63713 ;
  assign n63719 = ~n63717 & n63718 ;
  assign n63720 = ~n63707 & ~n63719 ;
  assign n63723 = n8860 & n49990 ;
  assign n63722 = ~\P1_P3_InstQueue_reg[6][5]/NET0131  & ~n49990 ;
  assign n63724 = n10046 & ~n63722 ;
  assign n63725 = ~n63723 & n63724 ;
  assign n63721 = \P1_P3_InstQueue_reg[6][5]/NET0131  & ~n49995 ;
  assign n63726 = \P1_buf2_reg[29]/NET0131  & n49930 ;
  assign n63727 = \P1_buf2_reg[21]/NET0131  & ~n49930 ;
  assign n63728 = n49950 & n63727 ;
  assign n63729 = ~n63726 & ~n63728 ;
  assign n63730 = n11698 & ~n63729 ;
  assign n63731 = \P1_buf2_reg[5]/NET0131  & n50005 ;
  assign n63732 = ~n63730 & ~n63731 ;
  assign n63733 = ~n63721 & n63732 ;
  assign n63734 = ~n63725 & n63733 ;
  assign n63737 = n26865 & n50021 ;
  assign n63736 = ~\P2_P3_InstQueue_reg[0][5]/NET0131  & ~n50021 ;
  assign n63738 = n27788 & ~n63736 ;
  assign n63739 = ~n63737 & n63738 ;
  assign n63735 = \P2_P3_InstQueue_reg[0][5]/NET0131  & ~n50030 ;
  assign n63740 = \P2_buf2_reg[29]/NET0131  & n50012 ;
  assign n63741 = \P2_buf2_reg[21]/NET0131  & n50015 ;
  assign n63742 = ~n63740 & ~n63741 ;
  assign n63743 = n27325 & ~n63742 ;
  assign n63744 = \P2_buf2_reg[5]/NET0131  & n50040 ;
  assign n63745 = ~n63743 & ~n63744 ;
  assign n63746 = ~n63735 & n63745 ;
  assign n63747 = ~n63739 & n63746 ;
  assign n63750 = n26865 & n50051 ;
  assign n63749 = ~\P2_P3_InstQueue_reg[10][5]/NET0131  & ~n50051 ;
  assign n63751 = n27788 & ~n63749 ;
  assign n63752 = ~n63750 & n63751 ;
  assign n63748 = \P2_P3_InstQueue_reg[10][5]/NET0131  & ~n50056 ;
  assign n63753 = \P2_buf2_reg[21]/NET0131  & n50045 ;
  assign n63754 = \P2_buf2_reg[29]/NET0131  & n50046 ;
  assign n63755 = ~n63753 & ~n63754 ;
  assign n63756 = n27325 & ~n63755 ;
  assign n63757 = \P2_buf2_reg[5]/NET0131  & n50066 ;
  assign n63758 = ~n63756 & ~n63757 ;
  assign n63759 = ~n63748 & n63758 ;
  assign n63760 = ~n63752 & n63759 ;
  assign n63763 = n8860 & n49770 ;
  assign n63762 = ~\P1_P3_InstQueue_reg[7][5]/NET0131  & ~n49770 ;
  assign n63764 = n10046 & ~n63762 ;
  assign n63765 = ~n63763 & n63764 ;
  assign n63761 = \P1_P3_InstQueue_reg[7][5]/NET0131  & ~n50075 ;
  assign n63766 = \P1_buf2_reg[29]/NET0131  & n49950 ;
  assign n63767 = \P1_buf2_reg[21]/NET0131  & ~n49950 ;
  assign n63768 = n49970 & n63767 ;
  assign n63769 = ~n63766 & ~n63768 ;
  assign n63770 = n11698 & ~n63769 ;
  assign n63771 = \P1_buf2_reg[5]/NET0131  & n50085 ;
  assign n63772 = ~n63770 & ~n63771 ;
  assign n63773 = ~n63761 & n63772 ;
  assign n63774 = ~n63765 & n63773 ;
  assign n63777 = n26865 & n50094 ;
  assign n63776 = ~\P2_P3_InstQueue_reg[11][5]/NET0131  & ~n50094 ;
  assign n63778 = n27788 & ~n63776 ;
  assign n63779 = ~n63777 & n63778 ;
  assign n63775 = \P2_P3_InstQueue_reg[11][5]/NET0131  & ~n50097 ;
  assign n63780 = \P2_buf2_reg[29]/NET0131  & n50045 ;
  assign n63781 = \P2_buf2_reg[21]/NET0131  & n50053 ;
  assign n63782 = ~n63780 & ~n63781 ;
  assign n63783 = n27325 & ~n63782 ;
  assign n63784 = \P2_buf2_reg[5]/NET0131  & n50107 ;
  assign n63785 = ~n63783 & ~n63784 ;
  assign n63786 = ~n63775 & n63785 ;
  assign n63787 = ~n63779 & n63786 ;
  assign n63790 = n26865 & n50115 ;
  assign n63789 = ~\P2_P3_InstQueue_reg[12][5]/NET0131  & ~n50115 ;
  assign n63791 = n27788 & ~n63789 ;
  assign n63792 = ~n63790 & n63791 ;
  assign n63788 = \P2_P3_InstQueue_reg[12][5]/NET0131  & ~n50118 ;
  assign n63793 = \P2_buf2_reg[29]/NET0131  & n50053 ;
  assign n63794 = \P2_buf2_reg[21]/NET0131  & n50051 ;
  assign n63795 = ~n63793 & ~n63794 ;
  assign n63796 = n27325 & ~n63795 ;
  assign n63797 = \P2_buf2_reg[5]/NET0131  & n50128 ;
  assign n63798 = ~n63796 & ~n63797 ;
  assign n63799 = ~n63788 & n63798 ;
  assign n63800 = ~n63792 & n63799 ;
  assign n63803 = n8860 & n49771 ;
  assign n63802 = ~\P1_P3_InstQueue_reg[8][5]/NET0131  & ~n49771 ;
  assign n63804 = n10046 & ~n63802 ;
  assign n63805 = ~n63803 & n63804 ;
  assign n63801 = \P1_P3_InstQueue_reg[8][5]/NET0131  & ~n50136 ;
  assign n63806 = \P1_buf2_reg[29]/NET0131  & n49970 ;
  assign n63807 = \P1_buf2_reg[21]/NET0131  & ~n49970 ;
  assign n63808 = n49990 & n63807 ;
  assign n63809 = ~n63806 & ~n63808 ;
  assign n63810 = n11698 & ~n63809 ;
  assign n63811 = \P1_buf2_reg[5]/NET0131  & n50146 ;
  assign n63812 = ~n63810 & ~n63811 ;
  assign n63813 = ~n63801 & n63812 ;
  assign n63814 = ~n63805 & n63813 ;
  assign n63817 = n26865 & n50012 ;
  assign n63816 = ~\P2_P3_InstQueue_reg[13][5]/NET0131  & ~n50012 ;
  assign n63818 = n27788 & ~n63816 ;
  assign n63819 = ~n63817 & n63818 ;
  assign n63815 = \P2_P3_InstQueue_reg[13][5]/NET0131  & ~n50155 ;
  assign n63820 = \P2_buf2_reg[29]/NET0131  & n50051 ;
  assign n63821 = \P2_buf2_reg[21]/NET0131  & n50094 ;
  assign n63822 = ~n63820 & ~n63821 ;
  assign n63823 = n27325 & ~n63822 ;
  assign n63824 = \P2_buf2_reg[5]/NET0131  & n50165 ;
  assign n63825 = ~n63823 & ~n63824 ;
  assign n63826 = ~n63815 & n63825 ;
  assign n63827 = ~n63819 & n63826 ;
  assign n63830 = n26865 & n50015 ;
  assign n63829 = ~\P2_P3_InstQueue_reg[14][5]/NET0131  & ~n50015 ;
  assign n63831 = n27788 & ~n63829 ;
  assign n63832 = ~n63830 & n63831 ;
  assign n63828 = \P2_P3_InstQueue_reg[14][5]/NET0131  & ~n50173 ;
  assign n63833 = \P2_buf2_reg[29]/NET0131  & n50094 ;
  assign n63834 = \P2_buf2_reg[21]/NET0131  & n50115 ;
  assign n63835 = ~n63833 & ~n63834 ;
  assign n63836 = n27325 & ~n63835 ;
  assign n63837 = \P2_buf2_reg[5]/NET0131  & n50183 ;
  assign n63838 = ~n63836 & ~n63837 ;
  assign n63839 = ~n63828 & n63838 ;
  assign n63840 = ~n63832 & n63839 ;
  assign n63843 = n8860 & n49768 ;
  assign n63842 = ~\P1_P3_InstQueue_reg[9][5]/NET0131  & ~n49768 ;
  assign n63844 = n10046 & ~n63842 ;
  assign n63845 = ~n63843 & n63844 ;
  assign n63841 = \P1_P3_InstQueue_reg[9][5]/NET0131  & ~n50191 ;
  assign n63846 = \P1_buf2_reg[29]/NET0131  & n49990 ;
  assign n63847 = \P1_buf2_reg[21]/NET0131  & n49770 ;
  assign n63848 = ~n63846 & ~n63847 ;
  assign n63849 = n11698 & ~n63848 ;
  assign n63850 = \P1_buf2_reg[5]/NET0131  & n50201 ;
  assign n63851 = ~n63849 & ~n63850 ;
  assign n63852 = ~n63841 & n63851 ;
  assign n63853 = ~n63845 & n63852 ;
  assign n63856 = n26865 & n50024 ;
  assign n63855 = ~\P2_P3_InstQueue_reg[15][5]/NET0131  & ~n50024 ;
  assign n63857 = n27788 & ~n63855 ;
  assign n63858 = ~n63856 & n63857 ;
  assign n63854 = \P2_P3_InstQueue_reg[15][5]/NET0131  & ~n50210 ;
  assign n63859 = \P2_buf2_reg[29]/NET0131  & n50115 ;
  assign n63860 = \P2_buf2_reg[21]/NET0131  & n50012 ;
  assign n63861 = ~n63859 & ~n63860 ;
  assign n63862 = n27325 & ~n63861 ;
  assign n63863 = \P2_buf2_reg[5]/NET0131  & n50220 ;
  assign n63864 = ~n63862 & ~n63863 ;
  assign n63865 = ~n63854 & n63864 ;
  assign n63866 = ~n63858 & n63865 ;
  assign n63869 = n26865 & n50227 ;
  assign n63868 = ~\P2_P3_InstQueue_reg[1][5]/NET0131  & ~n50227 ;
  assign n63870 = n27788 & ~n63868 ;
  assign n63871 = ~n63869 & n63870 ;
  assign n63867 = \P2_P3_InstQueue_reg[1][5]/NET0131  & ~n50230 ;
  assign n63872 = \P2_buf2_reg[29]/NET0131  & n50015 ;
  assign n63873 = \P2_buf2_reg[21]/NET0131  & n50024 ;
  assign n63874 = ~n63872 & ~n63873 ;
  assign n63875 = n27325 & ~n63874 ;
  assign n63876 = \P2_buf2_reg[5]/NET0131  & n50240 ;
  assign n63877 = ~n63875 & ~n63876 ;
  assign n63878 = ~n63867 & n63877 ;
  assign n63879 = ~n63871 & n63878 ;
  assign n63882 = n26865 & n50247 ;
  assign n63881 = ~\P2_P3_InstQueue_reg[2][5]/NET0131  & ~n50247 ;
  assign n63883 = n27788 & ~n63881 ;
  assign n63884 = ~n63882 & n63883 ;
  assign n63880 = \P2_P3_InstQueue_reg[2][5]/NET0131  & ~n50250 ;
  assign n63885 = \P2_buf2_reg[21]/NET0131  & n50021 ;
  assign n63886 = \P2_buf2_reg[29]/NET0131  & n50024 ;
  assign n63887 = ~n63885 & ~n63886 ;
  assign n63888 = n27325 & ~n63887 ;
  assign n63889 = \P2_buf2_reg[5]/NET0131  & n50260 ;
  assign n63890 = ~n63888 & ~n63889 ;
  assign n63891 = ~n63880 & n63890 ;
  assign n63892 = ~n63884 & n63891 ;
  assign n63895 = n26865 & n50267 ;
  assign n63894 = ~\P2_P3_InstQueue_reg[3][5]/NET0131  & ~n50267 ;
  assign n63896 = n27788 & ~n63894 ;
  assign n63897 = ~n63895 & n63896 ;
  assign n63893 = \P2_P3_InstQueue_reg[3][5]/NET0131  & ~n50270 ;
  assign n63898 = \P2_buf2_reg[29]/NET0131  & n50021 ;
  assign n63899 = \P2_buf2_reg[21]/NET0131  & n50227 ;
  assign n63900 = ~n63898 & ~n63899 ;
  assign n63901 = n27325 & ~n63900 ;
  assign n63902 = \P2_buf2_reg[5]/NET0131  & n50280 ;
  assign n63903 = ~n63901 & ~n63902 ;
  assign n63904 = ~n63893 & n63903 ;
  assign n63905 = ~n63897 & n63904 ;
  assign n63908 = n26865 & n50287 ;
  assign n63907 = ~\P2_P3_InstQueue_reg[4][5]/NET0131  & ~n50287 ;
  assign n63909 = n27788 & ~n63907 ;
  assign n63910 = ~n63908 & n63909 ;
  assign n63906 = \P2_P3_InstQueue_reg[4][5]/NET0131  & ~n50290 ;
  assign n63911 = \P2_buf2_reg[29]/NET0131  & n50227 ;
  assign n63912 = \P2_buf2_reg[21]/NET0131  & n50247 ;
  assign n63913 = ~n63911 & ~n63912 ;
  assign n63914 = n27325 & ~n63913 ;
  assign n63915 = \P2_buf2_reg[5]/NET0131  & n50300 ;
  assign n63916 = ~n63914 & ~n63915 ;
  assign n63917 = ~n63906 & n63916 ;
  assign n63918 = ~n63910 & n63917 ;
  assign n63921 = n26865 & n50307 ;
  assign n63920 = ~\P2_P3_InstQueue_reg[5][5]/NET0131  & ~n50307 ;
  assign n63922 = n27788 & ~n63920 ;
  assign n63923 = ~n63921 & n63922 ;
  assign n63919 = \P2_P3_InstQueue_reg[5][5]/NET0131  & ~n50310 ;
  assign n63924 = \P2_buf2_reg[29]/NET0131  & n50247 ;
  assign n63925 = \P2_buf2_reg[21]/NET0131  & n50267 ;
  assign n63926 = ~n63924 & ~n63925 ;
  assign n63927 = n27325 & ~n63926 ;
  assign n63928 = \P2_buf2_reg[5]/NET0131  & n50320 ;
  assign n63929 = ~n63927 & ~n63928 ;
  assign n63930 = ~n63919 & n63929 ;
  assign n63931 = ~n63923 & n63930 ;
  assign n63934 = n26865 & n50327 ;
  assign n63933 = ~\P2_P3_InstQueue_reg[6][5]/NET0131  & ~n50327 ;
  assign n63935 = n27788 & ~n63933 ;
  assign n63936 = ~n63934 & n63935 ;
  assign n63932 = \P2_P3_InstQueue_reg[6][5]/NET0131  & ~n50330 ;
  assign n63937 = \P2_buf2_reg[29]/NET0131  & n50267 ;
  assign n63938 = \P2_buf2_reg[21]/NET0131  & n50287 ;
  assign n63939 = ~n63937 & ~n63938 ;
  assign n63940 = n27325 & ~n63939 ;
  assign n63941 = \P2_buf2_reg[5]/NET0131  & n50340 ;
  assign n63942 = ~n63940 & ~n63941 ;
  assign n63943 = ~n63932 & n63942 ;
  assign n63944 = ~n63936 & n63943 ;
  assign n63947 = n26865 & n50046 ;
  assign n63946 = ~\P2_P3_InstQueue_reg[7][5]/NET0131  & ~n50046 ;
  assign n63948 = n27788 & ~n63946 ;
  assign n63949 = ~n63947 & n63948 ;
  assign n63945 = \P2_P3_InstQueue_reg[7][5]/NET0131  & ~n50349 ;
  assign n63950 = \P2_buf2_reg[29]/NET0131  & n50287 ;
  assign n63951 = \P2_buf2_reg[21]/NET0131  & n50307 ;
  assign n63952 = ~n63950 & ~n63951 ;
  assign n63953 = n27325 & ~n63952 ;
  assign n63954 = \P2_buf2_reg[5]/NET0131  & n50359 ;
  assign n63955 = ~n63953 & ~n63954 ;
  assign n63956 = ~n63945 & n63955 ;
  assign n63957 = ~n63949 & n63956 ;
  assign n63960 = n26865 & n50045 ;
  assign n63959 = ~\P2_P3_InstQueue_reg[8][5]/NET0131  & ~n50045 ;
  assign n63961 = n27788 & ~n63959 ;
  assign n63962 = ~n63960 & n63961 ;
  assign n63958 = \P2_P3_InstQueue_reg[8][5]/NET0131  & ~n50367 ;
  assign n63963 = \P2_buf2_reg[29]/NET0131  & n50307 ;
  assign n63964 = \P2_buf2_reg[21]/NET0131  & n50327 ;
  assign n63965 = ~n63963 & ~n63964 ;
  assign n63966 = n27325 & ~n63965 ;
  assign n63967 = \P2_buf2_reg[5]/NET0131  & n50377 ;
  assign n63968 = ~n63966 & ~n63967 ;
  assign n63969 = ~n63958 & n63968 ;
  assign n63970 = ~n63962 & n63969 ;
  assign n63973 = n26865 & n50053 ;
  assign n63972 = ~\P2_P3_InstQueue_reg[9][5]/NET0131  & ~n50053 ;
  assign n63974 = n27788 & ~n63972 ;
  assign n63975 = ~n63973 & n63974 ;
  assign n63971 = \P2_P3_InstQueue_reg[9][5]/NET0131  & ~n50385 ;
  assign n63976 = \P2_buf2_reg[29]/NET0131  & n50327 ;
  assign n63977 = \P2_buf2_reg[21]/NET0131  & n50046 ;
  assign n63978 = ~n63976 & ~n63977 ;
  assign n63979 = n27325 & ~n63978 ;
  assign n63980 = \P2_buf2_reg[5]/NET0131  & n50395 ;
  assign n63981 = ~n63979 & ~n63980 ;
  assign n63982 = ~n63971 & n63981 ;
  assign n63983 = ~n63975 & n63982 ;
  assign n63985 = n52097 & n63368 ;
  assign n63986 = \P2_P2_rEIP_reg[7]/NET0131  & n63985 ;
  assign n63987 = \P2_P2_rEIP_reg[8]/NET0131  & n63986 ;
  assign n63988 = \P2_P2_rEIP_reg[9]/NET0131  & n63987 ;
  assign n63989 = n52105 & n63988 ;
  assign n63990 = n52104 & n63989 ;
  assign n63991 = \P2_P2_rEIP_reg[14]/NET0131  & n63990 ;
  assign n63992 = \P2_P2_rEIP_reg[15]/NET0131  & n63991 ;
  assign n63993 = \P2_P2_rEIP_reg[16]/NET0131  & n63992 ;
  assign n63994 = ~\P2_P2_rEIP_reg[17]/NET0131  & ~n63993 ;
  assign n63995 = n54148 & n63368 ;
  assign n63996 = n63373 & ~n63995 ;
  assign n63997 = ~n63994 & n63996 ;
  assign n63984 = \P2_P2_Address_reg[16]/NET0131  & ~n26646 ;
  assign n63998 = n52108 & n63358 ;
  assign n63999 = n52101 & n63998 ;
  assign n64001 = \P2_P2_rEIP_reg[18]/NET0131  & n63999 ;
  assign n64000 = ~\P2_P2_rEIP_reg[18]/NET0131  & ~n63999 ;
  assign n64002 = n26647 & ~n64000 ;
  assign n64003 = ~n64001 & n64002 ;
  assign n64004 = ~n63984 & ~n64003 ;
  assign n64005 = ~n63997 & n64004 ;
  assign n64007 = \P1_P1_rEIP_reg[15]/NET0131  & n63393 ;
  assign n64008 = \P1_P1_rEIP_reg[16]/NET0131  & n64007 ;
  assign n64009 = \P1_P1_rEIP_reg[17]/NET0131  & n64008 ;
  assign n64010 = ~\P1_P1_rEIP_reg[18]/NET0131  & ~n64009 ;
  assign n64011 = n51665 & n64008 ;
  assign n64012 = n26155 & ~n64011 ;
  assign n64013 = ~n64010 & n64012 ;
  assign n64006 = \P1_P1_Address_reg[16]/NET0131  & ~n26154 ;
  assign n64014 = n51679 & n63402 ;
  assign n64016 = ~\P1_P1_rEIP_reg[17]/NET0131  & ~n64014 ;
  assign n64015 = \P1_P1_rEIP_reg[17]/NET0131  & n64014 ;
  assign n64017 = n63401 & ~n64015 ;
  assign n64018 = ~n64016 & n64017 ;
  assign n64019 = ~n64006 & ~n64018 ;
  assign n64020 = ~n64013 & n64019 ;
  assign n64022 = \P1_P2_rEIP_reg[11]/NET0131  & n48391 ;
  assign n64023 = n54902 & n63421 ;
  assign n64024 = n64022 & n64023 ;
  assign n64025 = \P1_P2_rEIP_reg[15]/NET0131  & n64024 ;
  assign n64026 = \P1_P2_rEIP_reg[16]/NET0131  & n64025 ;
  assign n64028 = \P1_P2_rEIP_reg[17]/NET0131  & n64026 ;
  assign n64027 = ~\P1_P2_rEIP_reg[17]/NET0131  & ~n64026 ;
  assign n64029 = n63420 & ~n64027 ;
  assign n64030 = ~n64028 & n64029 ;
  assign n64021 = \P1_P2_Address_reg[16]/NET0131  & ~n25764 ;
  assign n64031 = \P1_P2_rEIP_reg[9]/NET0131  & n63435 ;
  assign n64032 = n48392 & n64031 ;
  assign n64033 = n51198 & n64032 ;
  assign n64034 = n48387 & n64033 ;
  assign n64035 = ~\P1_P2_rEIP_reg[18]/NET0131  & ~n64034 ;
  assign n64036 = n25765 & ~n63436 ;
  assign n64037 = ~n64035 & n64036 ;
  assign n64038 = ~n64021 & ~n64037 ;
  assign n64039 = ~n64030 & n64038 ;
  assign n64042 = \P2_P1_rEIP_reg[18]/NET0131  & n63463 ;
  assign n64041 = ~\P2_P1_rEIP_reg[18]/NET0131  & ~n63463 ;
  assign n64043 = n25955 & ~n64041 ;
  assign n64044 = ~n64042 & n64043 ;
  assign n64040 = \P2_P1_Address_reg[16]/NET0131  & ~n25954 ;
  assign n64053 = n50776 & n63475 ;
  assign n64045 = n50768 & n63475 ;
  assign n64046 = \P2_P1_rEIP_reg[7]/NET0131  & n64045 ;
  assign n64047 = \P2_P1_rEIP_reg[8]/NET0131  & n64046 ;
  assign n64048 = \P2_P1_rEIP_reg[9]/NET0131  & n64047 ;
  assign n64049 = n50772 & n64048 ;
  assign n64050 = n50966 & n64049 ;
  assign n64051 = n50763 & n64050 ;
  assign n64052 = ~\P2_P1_rEIP_reg[17]/NET0131  & ~n64051 ;
  assign n64054 = n63480 & ~n64052 ;
  assign n64055 = ~n64053 & n64054 ;
  assign n64056 = ~n64040 & ~n64055 ;
  assign n64057 = ~n64044 & n64056 ;
  assign n64059 = ~\P1_P3_rEIP_reg[0]/NET0131  & ~\P1_P3_rEIP_reg[1]/NET0131  ;
  assign n64060 = \P1_P3_rEIP_reg[31]/NET0131  & ~n64059 ;
  assign n64061 = \P1_P3_rEIP_reg[2]/NET0131  & n64060 ;
  assign n64062 = \P1_P3_rEIP_reg[3]/NET0131  & n64061 ;
  assign n64063 = \P1_P3_rEIP_reg[4]/NET0131  & n64062 ;
  assign n64064 = \P1_P3_rEIP_reg[5]/NET0131  & n64063 ;
  assign n64065 = \P1_P3_rEIP_reg[6]/NET0131  & n64064 ;
  assign n64066 = \P1_P3_rEIP_reg[7]/NET0131  & n64065 ;
  assign n64067 = \P1_P3_rEIP_reg[8]/NET0131  & n64066 ;
  assign n64068 = \P1_P3_rEIP_reg[9]/NET0131  & n64067 ;
  assign n64069 = \P1_P3_rEIP_reg[10]/NET0131  & n64068 ;
  assign n64070 = \P1_P3_rEIP_reg[11]/NET0131  & n64069 ;
  assign n64071 = \P1_P3_rEIP_reg[12]/NET0131  & n64070 ;
  assign n64072 = \P1_P3_rEIP_reg[13]/NET0131  & n64071 ;
  assign n64073 = \P1_P3_rEIP_reg[14]/NET0131  & n64072 ;
  assign n64074 = \P1_P3_rEIP_reg[15]/NET0131  & n64073 ;
  assign n64075 = \P1_P3_rEIP_reg[16]/NET0131  & n64074 ;
  assign n64076 = \P1_P3_rEIP_reg[17]/NET0131  & n64075 ;
  assign n64078 = \P1_P3_rEIP_reg[18]/NET0131  & n64076 ;
  assign n64077 = ~\P1_P3_rEIP_reg[18]/NET0131  & ~n64076 ;
  assign n64079 = n9092 & ~n64077 ;
  assign n64080 = ~n64078 & n64079 ;
  assign n64058 = \P1_P3_Address_reg[16]/NET0131  & ~n9091 ;
  assign n64081 = \P1_P3_rEIP_reg[0]/NET0131  & \P1_P3_rEIP_reg[31]/NET0131  ;
  assign n64082 = n16578 & n64081 ;
  assign n64083 = \P1_P3_rEIP_reg[13]/NET0131  & n64082 ;
  assign n64084 = \P1_P3_rEIP_reg[14]/NET0131  & n64083 ;
  assign n64085 = \P1_P3_rEIP_reg[15]/NET0131  & n64084 ;
  assign n64086 = \P1_P3_rEIP_reg[16]/NET0131  & n64085 ;
  assign n64088 = ~\P1_P3_rEIP_reg[17]/NET0131  & ~n64086 ;
  assign n64087 = \P1_P3_rEIP_reg[17]/NET0131  & n64086 ;
  assign n64089 = n22115 & ~n64087 ;
  assign n64090 = ~n64088 & n64089 ;
  assign n64091 = ~n64058 & ~n64090 ;
  assign n64092 = ~n64080 & n64091 ;
  assign n64101 = ~\P2_P3_rEIP_reg[0]/NET0131  & ~\P2_P3_rEIP_reg[1]/NET0131  ;
  assign n64102 = \P2_P3_rEIP_reg[31]/NET0131  & ~n64101 ;
  assign n64103 = \P2_P3_rEIP_reg[2]/NET0131  & n64102 ;
  assign n64104 = \P2_P3_rEIP_reg[3]/NET0131  & n64103 ;
  assign n64105 = \P2_P3_rEIP_reg[4]/NET0131  & n64104 ;
  assign n64106 = \P2_P3_rEIP_reg[5]/NET0131  & n64105 ;
  assign n64107 = \P2_P3_rEIP_reg[6]/NET0131  & n64106 ;
  assign n64108 = \P2_P3_rEIP_reg[7]/NET0131  & n64107 ;
  assign n64109 = \P2_P3_rEIP_reg[8]/NET0131  & n64108 ;
  assign n64110 = \P2_P3_rEIP_reg[9]/NET0131  & n64109 ;
  assign n64111 = \P2_P3_rEIP_reg[10]/NET0131  & n64110 ;
  assign n64112 = \P2_P3_rEIP_reg[11]/NET0131  & n64111 ;
  assign n64113 = \P2_P3_rEIP_reg[12]/NET0131  & n64112 ;
  assign n64114 = \P2_P3_rEIP_reg[13]/NET0131  & n64113 ;
  assign n64115 = \P2_P3_rEIP_reg[14]/NET0131  & n64114 ;
  assign n64116 = \P2_P3_rEIP_reg[15]/NET0131  & n64115 ;
  assign n64117 = \P2_P3_rEIP_reg[16]/NET0131  & n64116 ;
  assign n64118 = \P2_P3_rEIP_reg[17]/NET0131  & n64117 ;
  assign n64120 = ~\P2_P3_rEIP_reg[18]/NET0131  & ~n64118 ;
  assign n64119 = \P2_P3_rEIP_reg[18]/NET0131  & n64118 ;
  assign n64121 = n27145 & ~n64119 ;
  assign n64122 = ~n64120 & n64121 ;
  assign n64093 = \P2_P3_Address_reg[16]/NET0131  & ~n27144 ;
  assign n64095 = \P2_P3_rEIP_reg[0]/NET0131  & \P2_P3_rEIP_reg[31]/NET0131  ;
  assign n64097 = n52561 & n64095 ;
  assign n64098 = ~\P2_P3_rEIP_reg[17]/NET0131  & ~n64097 ;
  assign n64094 = \P2_P3_State_reg[2]/NET0131  & n27144 ;
  assign n64096 = n52562 & n64095 ;
  assign n64099 = n64094 & ~n64096 ;
  assign n64100 = ~n64098 & n64099 ;
  assign n64123 = ~n64093 & ~n64100 ;
  assign n64124 = ~n64122 & n64123 ;
  assign n64125 = ~\P1_P2_InstQueueWr_Addr_reg[3]/NET0131  & ~n28056 ;
  assign n64126 = ~n28057 & ~n64125 ;
  assign n64128 = ~n28067 & n64126 ;
  assign n64129 = ~n28302 & ~n64128 ;
  assign n64130 = ~n28064 & ~n64129 ;
  assign n64131 = ~n28107 & ~n28280 ;
  assign n64132 = ~n64130 & n64131 ;
  assign n64133 = n25933 & ~n28108 ;
  assign n64134 = ~n64132 & n64133 ;
  assign n64135 = \P1_P2_InstQueueWr_Addr_reg[3]/NET0131  & ~n63509 ;
  assign n64127 = n27608 & n64126 ;
  assign n64136 = n36630 & ~n64129 ;
  assign n64137 = ~n64127 & ~n64136 ;
  assign n64138 = ~n64135 & n64137 ;
  assign n64139 = ~n64134 & n64138 ;
  assign n64140 = ~\P1_P1_InstQueueWr_Addr_reg[3]/NET0131  & ~n8377 ;
  assign n64141 = ~n8378 & ~n64140 ;
  assign n64143 = ~n8371 & n64141 ;
  assign n64144 = ~n8640 & ~n64143 ;
  assign n64145 = ~n8374 & ~n64144 ;
  assign n64146 = ~n8426 & ~n8616 ;
  assign n64147 = ~n64145 & n64146 ;
  assign n64148 = ~n8427 & n27791 ;
  assign n64149 = ~n64147 & n64148 ;
  assign n64150 = \P1_P1_InstQueueWr_Addr_reg[3]/NET0131  & ~n63490 ;
  assign n64142 = n8350 & n64141 ;
  assign n64151 = ~n36701 & ~n64144 ;
  assign n64152 = ~n64142 & ~n64151 ;
  assign n64153 = ~n64150 & n64152 ;
  assign n64154 = ~n64149 & n64153 ;
  assign n64159 = n11698 & ~n49814 ;
  assign n64162 = ~n49738 & n64159 ;
  assign n64163 = n36810 & ~n64162 ;
  assign n64155 = \P1_P3_InstQueueWr_Addr_reg[3]/NET0131  & ~n49734 ;
  assign n64156 = ~n49770 & ~n64155 ;
  assign n64164 = ~n49741 & n64156 ;
  assign n64165 = ~n49742 & ~n64164 ;
  assign n64166 = ~n64163 & n64165 ;
  assign n64158 = \P1_P3_InstQueueWr_Addr_reg[3]/NET0131  & ~n63525 ;
  assign n64157 = n10046 & ~n64156 ;
  assign n64160 = ~n49813 & ~n49970 ;
  assign n64161 = n64159 & ~n64160 ;
  assign n64167 = ~n64157 & ~n64161 ;
  assign n64168 = ~n64158 & n64167 ;
  assign n64169 = ~n64166 & n64168 ;
  assign n64170 = ~\P2_P3_InstQueueWr_Addr_reg[3]/NET0131  & ~n50023 ;
  assign n64171 = ~n50024 & ~n64170 ;
  assign n64172 = ~n50014 & n64171 ;
  assign n64173 = ~n50327 & ~n64172 ;
  assign n64175 = ~n50011 & ~n64173 ;
  assign n64176 = ~n50114 & ~n50307 ;
  assign n64177 = ~n64175 & n64176 ;
  assign n64178 = n27325 & ~n50115 ;
  assign n64179 = ~n64177 & n64178 ;
  assign n64180 = \P2_P3_InstQueueWr_Addr_reg[3]/NET0131  & ~n63706 ;
  assign n64174 = ~n36831 & ~n64173 ;
  assign n64181 = n27788 & n64171 ;
  assign n64182 = ~n64174 & ~n64181 ;
  assign n64183 = ~n64180 & n64182 ;
  assign n64184 = ~n64179 & n64183 ;
  assign n64185 = \P1_P1_InstQueueWr_Addr_reg[1]/NET0131  & ~n63489 ;
  assign n64186 = ~\P1_P1_InstQueueWr_Addr_reg[0]/NET0131  & n8350 ;
  assign n64187 = \P1_P1_InstQueueWr_Addr_reg[1]/NET0131  & n52935 ;
  assign n64188 = ~n27791 & n64187 ;
  assign n64189 = ~n64186 & n64188 ;
  assign n64190 = \P1_P1_InstQueueWr_Addr_reg[0]/NET0131  & n8350 ;
  assign n64191 = ~\P1_P1_InstQueueWr_Addr_reg[1]/NET0131  & ~n64190 ;
  assign n64192 = n36701 & n64191 ;
  assign n64193 = ~n64189 & ~n64192 ;
  assign n64194 = ~n64185 & ~n64193 ;
  assign n64195 = \P1_P2_InstQueueWr_Addr_reg[1]/NET0131  & ~n63508 ;
  assign n64196 = ~\P1_P2_InstQueueWr_Addr_reg[0]/NET0131  & n27608 ;
  assign n64197 = \P1_P2_InstQueueWr_Addr_reg[1]/NET0131  & n52882 ;
  assign n64198 = ~n25933 & n64197 ;
  assign n64199 = ~n64196 & n64198 ;
  assign n64200 = \P1_P2_InstQueueWr_Addr_reg[0]/NET0131  & n27608 ;
  assign n64201 = ~\P1_P2_InstQueueWr_Addr_reg[1]/NET0131  & ~n64200 ;
  assign n64202 = ~n36630 & n64201 ;
  assign n64203 = ~n64199 & ~n64202 ;
  assign n64204 = ~n64195 & ~n64203 ;
  assign n64205 = \P1_P3_InstQueueWr_Addr_reg[1]/NET0131  & ~n63524 ;
  assign n64206 = ~\P1_P3_InstQueueWr_Addr_reg[0]/NET0131  & n10046 ;
  assign n64207 = \P1_P3_InstQueueWr_Addr_reg[1]/NET0131  & ~n21771 ;
  assign n64208 = ~n11698 & n64207 ;
  assign n64209 = ~n64206 & n64208 ;
  assign n64210 = \P1_P3_InstQueueWr_Addr_reg[0]/NET0131  & n10046 ;
  assign n64211 = ~\P1_P3_InstQueueWr_Addr_reg[1]/NET0131  & ~n64210 ;
  assign n64212 = n36810 & n64211 ;
  assign n64213 = ~n64209 & ~n64212 ;
  assign n64214 = ~n64205 & ~n64213 ;
  assign n64215 = \P2_P3_InstQueueWr_Addr_reg[1]/NET0131  & ~n63705 ;
  assign n64216 = ~\P2_P3_InstQueueWr_Addr_reg[0]/NET0131  & n27788 ;
  assign n64217 = \P2_P3_InstQueueWr_Addr_reg[1]/NET0131  & n52996 ;
  assign n64218 = ~n27325 & n64217 ;
  assign n64219 = ~n64216 & n64218 ;
  assign n64220 = \P2_P3_InstQueueWr_Addr_reg[0]/NET0131  & n27788 ;
  assign n64221 = ~\P2_P3_InstQueueWr_Addr_reg[1]/NET0131  & ~n64220 ;
  assign n64222 = n36831 & n64221 ;
  assign n64223 = ~n64219 & ~n64222 ;
  assign n64224 = ~n64215 & ~n64223 ;
  assign n64227 = ~n27308 & n43272 ;
  assign n64228 = \P2_P3_InstQueueWr_Addr_reg[0]/NET0131  & ~n64227 ;
  assign n64225 = ~\P2_P3_Flush_reg/NET0131  & ~\P2_P3_InstQueueWr_Addr_reg[0]/NET0131  ;
  assign n64226 = n27661 & ~n64225 ;
  assign n64229 = ~n64216 & ~n64226 ;
  assign n64230 = ~n64228 & n64229 ;
  assign n64233 = ~n25918 & n43218 ;
  assign n64234 = \P1_P2_InstQueueWr_Addr_reg[0]/NET0131  & ~n64233 ;
  assign n64231 = ~\P1_P2_Flush_reg/NET0131  & ~\P1_P2_InstQueueWr_Addr_reg[0]/NET0131  ;
  assign n64232 = n27673 & ~n64231 ;
  assign n64235 = ~n64196 & ~n64232 ;
  assign n64236 = ~n64234 & n64235 ;
  assign n64239 = n26990 & n50012 ;
  assign n64238 = ~\P2_P3_InstQueue_reg[13][1]/NET0131  & ~n50012 ;
  assign n64240 = n27788 & ~n64238 ;
  assign n64241 = ~n64239 & n64240 ;
  assign n64237 = \P2_P3_InstQueue_reg[13][1]/NET0131  & ~n50155 ;
  assign n64242 = \P2_buf2_reg[25]/NET0131  & n50051 ;
  assign n64243 = \P2_buf2_reg[17]/NET0131  & n50094 ;
  assign n64244 = ~n64242 & ~n64243 ;
  assign n64245 = n27325 & ~n64244 ;
  assign n64246 = \P2_buf2_reg[1]/NET0131  & n50165 ;
  assign n64247 = ~n64245 & ~n64246 ;
  assign n64248 = ~n64237 & n64247 ;
  assign n64249 = ~n64241 & n64248 ;
  assign n64252 = n9018 & n49735 ;
  assign n64251 = ~\P1_P3_InstQueue_reg[15][1]/NET0131  & ~n49735 ;
  assign n64253 = n10046 & ~n64251 ;
  assign n64254 = ~n64252 & n64253 ;
  assign n64250 = \P1_P3_InstQueue_reg[15][1]/NET0131  & ~n49875 ;
  assign n64255 = \P1_buf2_reg[25]/NET0131  & n49814 ;
  assign n64256 = \P1_buf2_reg[17]/NET0131  & n49739 ;
  assign n64257 = ~n64255 & ~n64256 ;
  assign n64258 = n11698 & ~n64257 ;
  assign n64259 = \P1_buf2_reg[1]/NET0131  & n49885 ;
  assign n64260 = ~n64258 & ~n64259 ;
  assign n64261 = ~n64250 & n64260 ;
  assign n64262 = ~n64254 & n64261 ;
  assign n64265 = ~n9241 & n43259 ;
  assign n64266 = \P1_P3_InstQueueWr_Addr_reg[0]/NET0131  & ~n64265 ;
  assign n64263 = ~\P1_P3_Flush_reg/NET0131  & ~\P1_P3_InstQueueWr_Addr_reg[0]/NET0131  ;
  assign n64264 = n10041 & ~n64263 ;
  assign n64267 = ~n64206 & ~n64264 ;
  assign n64268 = ~n64266 & n64267 ;
  assign n64271 = n9018 & n49732 ;
  assign n64270 = ~\P1_P3_InstQueue_reg[0][1]/NET0131  & ~n49732 ;
  assign n64272 = n10046 & ~n64270 ;
  assign n64273 = ~n64271 & n64272 ;
  assign n64269 = \P1_P3_InstQueue_reg[0][1]/NET0131  & ~n49750 ;
  assign n64274 = \P1_buf2_reg[25]/NET0131  & n49739 ;
  assign n64275 = \P1_buf2_reg[17]/NET0131  & ~n49739 ;
  assign n64276 = n49742 & n64275 ;
  assign n64277 = ~n64274 & ~n64276 ;
  assign n64278 = n11698 & ~n64277 ;
  assign n64279 = \P1_buf2_reg[1]/NET0131  & n49760 ;
  assign n64280 = ~n64278 & ~n64279 ;
  assign n64281 = ~n64269 & n64280 ;
  assign n64282 = ~n64273 & n64281 ;
  assign n64285 = n9018 & n49766 ;
  assign n64284 = ~\P1_P3_InstQueue_reg[10][1]/NET0131  & ~n49766 ;
  assign n64286 = n10046 & ~n64284 ;
  assign n64287 = ~n64285 & n64286 ;
  assign n64283 = \P1_P3_InstQueue_reg[10][1]/NET0131  & ~n49776 ;
  assign n64288 = \P1_buf2_reg[25]/NET0131  & n49770 ;
  assign n64289 = \P1_buf2_reg[17]/NET0131  & n49771 ;
  assign n64290 = ~n64288 & ~n64289 ;
  assign n64291 = n11698 & ~n64290 ;
  assign n64292 = \P1_buf2_reg[1]/NET0131  & n49786 ;
  assign n64293 = ~n64291 & ~n64292 ;
  assign n64294 = ~n64283 & n64293 ;
  assign n64295 = ~n64287 & n64294 ;
  assign n64298 = n8924 & n49792 ;
  assign n64297 = ~\P1_P3_InstQueue_reg[11][0]/NET0131  & ~n49792 ;
  assign n64299 = n10046 & ~n64297 ;
  assign n64300 = ~n64298 & n64299 ;
  assign n64296 = \P1_P3_InstQueue_reg[11][0]/NET0131  & ~n49798 ;
  assign n64301 = \P1_buf2_reg[24]/NET0131  & n49771 ;
  assign n64302 = \P1_buf2_reg[16]/NET0131  & n49768 ;
  assign n64303 = ~n64301 & ~n64302 ;
  assign n64304 = n11698 & ~n64303 ;
  assign n64305 = \P1_buf2_reg[0]/NET0131  & n49808 ;
  assign n64306 = ~n64304 & ~n64305 ;
  assign n64307 = ~n64296 & n64306 ;
  assign n64308 = ~n64300 & n64307 ;
  assign n64311 = n9018 & n49792 ;
  assign n64310 = ~\P1_P3_InstQueue_reg[11][1]/NET0131  & ~n49792 ;
  assign n64312 = n10046 & ~n64310 ;
  assign n64313 = ~n64311 & n64312 ;
  assign n64309 = \P1_P3_InstQueue_reg[11][1]/NET0131  & ~n49798 ;
  assign n64314 = \P1_buf2_reg[25]/NET0131  & n49771 ;
  assign n64315 = \P1_buf2_reg[17]/NET0131  & n49768 ;
  assign n64316 = ~n64314 & ~n64315 ;
  assign n64317 = n11698 & ~n64316 ;
  assign n64318 = \P1_buf2_reg[1]/NET0131  & n49808 ;
  assign n64319 = ~n64317 & ~n64318 ;
  assign n64320 = ~n64309 & n64319 ;
  assign n64321 = ~n64313 & n64320 ;
  assign n64324 = n9018 & n49814 ;
  assign n64323 = ~\P1_P3_InstQueue_reg[12][1]/NET0131  & ~n49814 ;
  assign n64325 = n10046 & ~n64323 ;
  assign n64326 = ~n64324 & n64325 ;
  assign n64322 = \P1_P3_InstQueue_reg[12][1]/NET0131  & ~n49819 ;
  assign n64327 = \P1_buf2_reg[25]/NET0131  & n49768 ;
  assign n64328 = \P1_buf2_reg[17]/NET0131  & n49766 ;
  assign n64329 = ~n64327 & ~n64328 ;
  assign n64330 = n11698 & ~n64329 ;
  assign n64331 = \P1_buf2_reg[1]/NET0131  & n49829 ;
  assign n64332 = ~n64330 & ~n64331 ;
  assign n64333 = ~n64322 & n64332 ;
  assign n64334 = ~n64326 & n64333 ;
  assign n64337 = n9018 & n49739 ;
  assign n64336 = ~\P1_P3_InstQueue_reg[13][1]/NET0131  & ~n49739 ;
  assign n64338 = n10046 & ~n64336 ;
  assign n64339 = ~n64337 & n64338 ;
  assign n64335 = \P1_P3_InstQueue_reg[13][1]/NET0131  & ~n49838 ;
  assign n64340 = \P1_buf2_reg[25]/NET0131  & n49766 ;
  assign n64341 = \P1_buf2_reg[17]/NET0131  & ~n49766 ;
  assign n64342 = n49792 & n64341 ;
  assign n64343 = ~n64340 & ~n64342 ;
  assign n64344 = n11698 & ~n64343 ;
  assign n64345 = \P1_buf2_reg[1]/NET0131  & n49848 ;
  assign n64346 = ~n64344 & ~n64345 ;
  assign n64347 = ~n64335 & n64346 ;
  assign n64348 = ~n64339 & n64347 ;
  assign n64351 = n9018 & n49742 ;
  assign n64350 = ~\P1_P3_InstQueue_reg[14][1]/NET0131  & ~n49742 ;
  assign n64352 = n10046 & ~n64350 ;
  assign n64353 = ~n64351 & n64352 ;
  assign n64349 = \P1_P3_InstQueue_reg[14][1]/NET0131  & ~n49856 ;
  assign n64354 = \P1_buf2_reg[25]/NET0131  & n49792 ;
  assign n64355 = \P1_buf2_reg[17]/NET0131  & ~n49792 ;
  assign n64356 = n49814 & n64355 ;
  assign n64357 = ~n64354 & ~n64356 ;
  assign n64358 = n11698 & ~n64357 ;
  assign n64359 = \P1_buf2_reg[1]/NET0131  & n49866 ;
  assign n64360 = ~n64358 & ~n64359 ;
  assign n64361 = ~n64349 & n64360 ;
  assign n64362 = ~n64353 & n64361 ;
  assign n64365 = n9018 & n49890 ;
  assign n64364 = ~\P1_P3_InstQueue_reg[1][1]/NET0131  & ~n49890 ;
  assign n64366 = n10046 & ~n64364 ;
  assign n64367 = ~n64365 & n64366 ;
  assign n64363 = \P1_P3_InstQueue_reg[1][1]/NET0131  & ~n49895 ;
  assign n64368 = \P1_buf2_reg[25]/NET0131  & n49742 ;
  assign n64369 = \P1_buf2_reg[17]/NET0131  & n49735 ;
  assign n64370 = ~n64368 & ~n64369 ;
  assign n64371 = n11698 & ~n64370 ;
  assign n64372 = \P1_buf2_reg[1]/NET0131  & n49905 ;
  assign n64373 = ~n64371 & ~n64372 ;
  assign n64374 = ~n64363 & n64373 ;
  assign n64375 = ~n64367 & n64374 ;
  assign n64378 = n9018 & n49910 ;
  assign n64377 = ~\P1_P3_InstQueue_reg[2][1]/NET0131  & ~n49910 ;
  assign n64379 = n10046 & ~n64377 ;
  assign n64380 = ~n64378 & n64379 ;
  assign n64376 = \P1_P3_InstQueue_reg[2][1]/NET0131  & ~n49915 ;
  assign n64381 = \P1_buf2_reg[25]/NET0131  & n49735 ;
  assign n64382 = \P1_buf2_reg[17]/NET0131  & n49732 ;
  assign n64383 = ~n64381 & ~n64382 ;
  assign n64384 = n11698 & ~n64383 ;
  assign n64385 = \P1_buf2_reg[1]/NET0131  & n49925 ;
  assign n64386 = ~n64384 & ~n64385 ;
  assign n64387 = ~n64376 & n64386 ;
  assign n64388 = ~n64380 & n64387 ;
  assign n64391 = n8924 & n49930 ;
  assign n64390 = ~\P1_P3_InstQueue_reg[3][0]/NET0131  & ~n49930 ;
  assign n64392 = n10046 & ~n64390 ;
  assign n64393 = ~n64391 & n64392 ;
  assign n64389 = \P1_P3_InstQueue_reg[3][0]/NET0131  & ~n49935 ;
  assign n64394 = \P1_buf2_reg[24]/NET0131  & n49732 ;
  assign n64395 = \P1_buf2_reg[16]/NET0131  & ~n49732 ;
  assign n64396 = n49890 & n64395 ;
  assign n64397 = ~n64394 & ~n64396 ;
  assign n64398 = n11698 & ~n64397 ;
  assign n64399 = \P1_buf2_reg[0]/NET0131  & n49945 ;
  assign n64400 = ~n64398 & ~n64399 ;
  assign n64401 = ~n64389 & n64400 ;
  assign n64402 = ~n64393 & n64401 ;
  assign n64405 = n9018 & n49930 ;
  assign n64404 = ~\P1_P3_InstQueue_reg[3][1]/NET0131  & ~n49930 ;
  assign n64406 = n10046 & ~n64404 ;
  assign n64407 = ~n64405 & n64406 ;
  assign n64403 = \P1_P3_InstQueue_reg[3][1]/NET0131  & ~n49935 ;
  assign n64408 = \P1_buf2_reg[25]/NET0131  & n49732 ;
  assign n64409 = \P1_buf2_reg[17]/NET0131  & ~n49732 ;
  assign n64410 = n49890 & n64409 ;
  assign n64411 = ~n64408 & ~n64410 ;
  assign n64412 = n11698 & ~n64411 ;
  assign n64413 = \P1_buf2_reg[1]/NET0131  & n49945 ;
  assign n64414 = ~n64412 & ~n64413 ;
  assign n64415 = ~n64403 & n64414 ;
  assign n64416 = ~n64407 & n64415 ;
  assign n64419 = n9018 & n49950 ;
  assign n64418 = ~\P1_P3_InstQueue_reg[4][1]/NET0131  & ~n49950 ;
  assign n64420 = n10046 & ~n64418 ;
  assign n64421 = ~n64419 & n64420 ;
  assign n64417 = \P1_P3_InstQueue_reg[4][1]/NET0131  & ~n49955 ;
  assign n64422 = \P1_buf2_reg[25]/NET0131  & n49890 ;
  assign n64423 = \P1_buf2_reg[17]/NET0131  & ~n49890 ;
  assign n64424 = n49910 & n64423 ;
  assign n64425 = ~n64422 & ~n64424 ;
  assign n64426 = n11698 & ~n64425 ;
  assign n64427 = \P1_buf2_reg[1]/NET0131  & n49965 ;
  assign n64428 = ~n64426 & ~n64427 ;
  assign n64429 = ~n64417 & n64428 ;
  assign n64430 = ~n64421 & n64429 ;
  assign n64433 = n9018 & n49970 ;
  assign n64432 = ~\P1_P3_InstQueue_reg[5][1]/NET0131  & ~n49970 ;
  assign n64434 = n10046 & ~n64432 ;
  assign n64435 = ~n64433 & n64434 ;
  assign n64431 = \P1_P3_InstQueue_reg[5][1]/NET0131  & ~n49975 ;
  assign n64436 = \P1_buf2_reg[25]/NET0131  & n49910 ;
  assign n64437 = \P1_buf2_reg[17]/NET0131  & ~n49910 ;
  assign n64438 = n49930 & n64437 ;
  assign n64439 = ~n64436 & ~n64438 ;
  assign n64440 = n11698 & ~n64439 ;
  assign n64441 = \P1_buf2_reg[1]/NET0131  & n49985 ;
  assign n64442 = ~n64440 & ~n64441 ;
  assign n64443 = ~n64431 & n64442 ;
  assign n64444 = ~n64435 & n64443 ;
  assign n64447 = n9018 & n49990 ;
  assign n64446 = ~\P1_P3_InstQueue_reg[6][1]/NET0131  & ~n49990 ;
  assign n64448 = n10046 & ~n64446 ;
  assign n64449 = ~n64447 & n64448 ;
  assign n64445 = \P1_P3_InstQueue_reg[6][1]/NET0131  & ~n49995 ;
  assign n64450 = \P1_buf2_reg[25]/NET0131  & n49930 ;
  assign n64451 = \P1_buf2_reg[17]/NET0131  & ~n49930 ;
  assign n64452 = n49950 & n64451 ;
  assign n64453 = ~n64450 & ~n64452 ;
  assign n64454 = n11698 & ~n64453 ;
  assign n64455 = \P1_buf2_reg[1]/NET0131  & n50005 ;
  assign n64456 = ~n64454 & ~n64455 ;
  assign n64457 = ~n64445 & n64456 ;
  assign n64458 = ~n64449 & n64457 ;
  assign n64461 = n26990 & n50021 ;
  assign n64460 = ~\P2_P3_InstQueue_reg[0][1]/NET0131  & ~n50021 ;
  assign n64462 = n27788 & ~n64460 ;
  assign n64463 = ~n64461 & n64462 ;
  assign n64459 = \P2_P3_InstQueue_reg[0][1]/NET0131  & ~n50030 ;
  assign n64464 = \P2_buf2_reg[25]/NET0131  & n50012 ;
  assign n64465 = \P2_buf2_reg[17]/NET0131  & n50015 ;
  assign n64466 = ~n64464 & ~n64465 ;
  assign n64467 = n27325 & ~n64466 ;
  assign n64468 = \P2_buf2_reg[1]/NET0131  & n50040 ;
  assign n64469 = ~n64467 & ~n64468 ;
  assign n64470 = ~n64459 & n64469 ;
  assign n64471 = ~n64463 & n64470 ;
  assign n64474 = n8924 & n49770 ;
  assign n64473 = ~\P1_P3_InstQueue_reg[7][0]/NET0131  & ~n49770 ;
  assign n64475 = n10046 & ~n64473 ;
  assign n64476 = ~n64474 & n64475 ;
  assign n64472 = \P1_P3_InstQueue_reg[7][0]/NET0131  & ~n50075 ;
  assign n64477 = \P1_buf2_reg[24]/NET0131  & n49950 ;
  assign n64478 = \P1_buf2_reg[16]/NET0131  & ~n49950 ;
  assign n64479 = n49970 & n64478 ;
  assign n64480 = ~n64477 & ~n64479 ;
  assign n64481 = n11698 & ~n64480 ;
  assign n64482 = \P1_buf2_reg[0]/NET0131  & n50085 ;
  assign n64483 = ~n64481 & ~n64482 ;
  assign n64484 = ~n64472 & n64483 ;
  assign n64485 = ~n64476 & n64484 ;
  assign n64488 = n26990 & n50051 ;
  assign n64487 = ~\P2_P3_InstQueue_reg[10][1]/NET0131  & ~n50051 ;
  assign n64489 = n27788 & ~n64487 ;
  assign n64490 = ~n64488 & n64489 ;
  assign n64486 = \P2_P3_InstQueue_reg[10][1]/NET0131  & ~n50056 ;
  assign n64491 = \P2_buf2_reg[17]/NET0131  & n50045 ;
  assign n64492 = \P2_buf2_reg[25]/NET0131  & n50046 ;
  assign n64493 = ~n64491 & ~n64492 ;
  assign n64494 = n27325 & ~n64493 ;
  assign n64495 = \P2_buf2_reg[1]/NET0131  & n50066 ;
  assign n64496 = ~n64494 & ~n64495 ;
  assign n64497 = ~n64486 & n64496 ;
  assign n64498 = ~n64490 & n64497 ;
  assign n64501 = n9018 & n49770 ;
  assign n64500 = ~\P1_P3_InstQueue_reg[7][1]/NET0131  & ~n49770 ;
  assign n64502 = n10046 & ~n64500 ;
  assign n64503 = ~n64501 & n64502 ;
  assign n64499 = \P1_P3_InstQueue_reg[7][1]/NET0131  & ~n50075 ;
  assign n64504 = \P1_buf2_reg[25]/NET0131  & n49950 ;
  assign n64505 = \P1_buf2_reg[17]/NET0131  & ~n49950 ;
  assign n64506 = n49970 & n64505 ;
  assign n64507 = ~n64504 & ~n64506 ;
  assign n64508 = n11698 & ~n64507 ;
  assign n64509 = \P1_buf2_reg[1]/NET0131  & n50085 ;
  assign n64510 = ~n64508 & ~n64509 ;
  assign n64511 = ~n64499 & n64510 ;
  assign n64512 = ~n64503 & n64511 ;
  assign n64515 = n27022 & n50094 ;
  assign n64514 = ~\P2_P3_InstQueue_reg[11][0]/NET0131  & ~n50094 ;
  assign n64516 = n27788 & ~n64514 ;
  assign n64517 = ~n64515 & n64516 ;
  assign n64513 = \P2_P3_InstQueue_reg[11][0]/NET0131  & ~n50097 ;
  assign n64518 = \P2_buf2_reg[24]/NET0131  & n50045 ;
  assign n64519 = \P2_buf2_reg[16]/NET0131  & n50053 ;
  assign n64520 = ~n64518 & ~n64519 ;
  assign n64521 = n27325 & ~n64520 ;
  assign n64522 = \P2_buf2_reg[0]/NET0131  & n50107 ;
  assign n64523 = ~n64521 & ~n64522 ;
  assign n64524 = ~n64513 & n64523 ;
  assign n64525 = ~n64517 & n64524 ;
  assign n64528 = n26990 & n50094 ;
  assign n64527 = ~\P2_P3_InstQueue_reg[11][1]/NET0131  & ~n50094 ;
  assign n64529 = n27788 & ~n64527 ;
  assign n64530 = ~n64528 & n64529 ;
  assign n64526 = \P2_P3_InstQueue_reg[11][1]/NET0131  & ~n50097 ;
  assign n64531 = \P2_buf2_reg[25]/NET0131  & n50045 ;
  assign n64532 = \P2_buf2_reg[17]/NET0131  & n50053 ;
  assign n64533 = ~n64531 & ~n64532 ;
  assign n64534 = n27325 & ~n64533 ;
  assign n64535 = \P2_buf2_reg[1]/NET0131  & n50107 ;
  assign n64536 = ~n64534 & ~n64535 ;
  assign n64537 = ~n64526 & n64536 ;
  assign n64538 = ~n64530 & n64537 ;
  assign n64541 = n26990 & n50115 ;
  assign n64540 = ~\P2_P3_InstQueue_reg[12][1]/NET0131  & ~n50115 ;
  assign n64542 = n27788 & ~n64540 ;
  assign n64543 = ~n64541 & n64542 ;
  assign n64539 = \P2_P3_InstQueue_reg[12][1]/NET0131  & ~n50118 ;
  assign n64544 = \P2_buf2_reg[25]/NET0131  & n50053 ;
  assign n64545 = \P2_buf2_reg[17]/NET0131  & n50051 ;
  assign n64546 = ~n64544 & ~n64545 ;
  assign n64547 = n27325 & ~n64546 ;
  assign n64548 = \P2_buf2_reg[1]/NET0131  & n50128 ;
  assign n64549 = ~n64547 & ~n64548 ;
  assign n64550 = ~n64539 & n64549 ;
  assign n64551 = ~n64543 & n64550 ;
  assign n64554 = n9018 & n49771 ;
  assign n64553 = ~\P1_P3_InstQueue_reg[8][1]/NET0131  & ~n49771 ;
  assign n64555 = n10046 & ~n64553 ;
  assign n64556 = ~n64554 & n64555 ;
  assign n64552 = \P1_P3_InstQueue_reg[8][1]/NET0131  & ~n50136 ;
  assign n64557 = \P1_buf2_reg[25]/NET0131  & n49970 ;
  assign n64558 = \P1_buf2_reg[17]/NET0131  & ~n49970 ;
  assign n64559 = n49990 & n64558 ;
  assign n64560 = ~n64557 & ~n64559 ;
  assign n64561 = n11698 & ~n64560 ;
  assign n64562 = \P1_buf2_reg[1]/NET0131  & n50146 ;
  assign n64563 = ~n64561 & ~n64562 ;
  assign n64564 = ~n64552 & n64563 ;
  assign n64565 = ~n64556 & n64564 ;
  assign n64568 = n26990 & n50015 ;
  assign n64567 = ~\P2_P3_InstQueue_reg[14][1]/NET0131  & ~n50015 ;
  assign n64569 = n27788 & ~n64567 ;
  assign n64570 = ~n64568 & n64569 ;
  assign n64566 = \P2_P3_InstQueue_reg[14][1]/NET0131  & ~n50173 ;
  assign n64571 = \P2_buf2_reg[25]/NET0131  & n50094 ;
  assign n64572 = \P2_buf2_reg[17]/NET0131  & n50115 ;
  assign n64573 = ~n64571 & ~n64572 ;
  assign n64574 = n27325 & ~n64573 ;
  assign n64575 = \P2_buf2_reg[1]/NET0131  & n50183 ;
  assign n64576 = ~n64574 & ~n64575 ;
  assign n64577 = ~n64566 & n64576 ;
  assign n64578 = ~n64570 & n64577 ;
  assign n64581 = n9018 & n49768 ;
  assign n64580 = ~\P1_P3_InstQueue_reg[9][1]/NET0131  & ~n49768 ;
  assign n64582 = n10046 & ~n64580 ;
  assign n64583 = ~n64581 & n64582 ;
  assign n64579 = \P1_P3_InstQueue_reg[9][1]/NET0131  & ~n50191 ;
  assign n64584 = \P1_buf2_reg[25]/NET0131  & n49990 ;
  assign n64585 = \P1_buf2_reg[17]/NET0131  & n49770 ;
  assign n64586 = ~n64584 & ~n64585 ;
  assign n64587 = n11698 & ~n64586 ;
  assign n64588 = \P1_buf2_reg[1]/NET0131  & n50201 ;
  assign n64589 = ~n64587 & ~n64588 ;
  assign n64590 = ~n64579 & n64589 ;
  assign n64591 = ~n64583 & n64590 ;
  assign n64594 = n26990 & n50024 ;
  assign n64593 = ~\P2_P3_InstQueue_reg[15][1]/NET0131  & ~n50024 ;
  assign n64595 = n27788 & ~n64593 ;
  assign n64596 = ~n64594 & n64595 ;
  assign n64592 = \P2_P3_InstQueue_reg[15][1]/NET0131  & ~n50210 ;
  assign n64597 = \P2_buf2_reg[25]/NET0131  & n50115 ;
  assign n64598 = \P2_buf2_reg[17]/NET0131  & n50012 ;
  assign n64599 = ~n64597 & ~n64598 ;
  assign n64600 = n27325 & ~n64599 ;
  assign n64601 = \P2_buf2_reg[1]/NET0131  & n50220 ;
  assign n64602 = ~n64600 & ~n64601 ;
  assign n64603 = ~n64592 & n64602 ;
  assign n64604 = ~n64596 & n64603 ;
  assign n64607 = n26990 & n50227 ;
  assign n64606 = ~\P2_P3_InstQueue_reg[1][1]/NET0131  & ~n50227 ;
  assign n64608 = n27788 & ~n64606 ;
  assign n64609 = ~n64607 & n64608 ;
  assign n64605 = \P2_P3_InstQueue_reg[1][1]/NET0131  & ~n50230 ;
  assign n64610 = \P2_buf2_reg[25]/NET0131  & n50015 ;
  assign n64611 = \P2_buf2_reg[17]/NET0131  & n50024 ;
  assign n64612 = ~n64610 & ~n64611 ;
  assign n64613 = n27325 & ~n64612 ;
  assign n64614 = \P2_buf2_reg[1]/NET0131  & n50240 ;
  assign n64615 = ~n64613 & ~n64614 ;
  assign n64616 = ~n64605 & n64615 ;
  assign n64617 = ~n64609 & n64616 ;
  assign n64620 = n26990 & n50247 ;
  assign n64619 = ~\P2_P3_InstQueue_reg[2][1]/NET0131  & ~n50247 ;
  assign n64621 = n27788 & ~n64619 ;
  assign n64622 = ~n64620 & n64621 ;
  assign n64618 = \P2_P3_InstQueue_reg[2][1]/NET0131  & ~n50250 ;
  assign n64623 = \P2_buf2_reg[17]/NET0131  & n50021 ;
  assign n64624 = \P2_buf2_reg[25]/NET0131  & n50024 ;
  assign n64625 = ~n64623 & ~n64624 ;
  assign n64626 = n27325 & ~n64625 ;
  assign n64627 = \P2_buf2_reg[1]/NET0131  & n50260 ;
  assign n64628 = ~n64626 & ~n64627 ;
  assign n64629 = ~n64618 & n64628 ;
  assign n64630 = ~n64622 & n64629 ;
  assign n64633 = n27022 & n50267 ;
  assign n64632 = ~\P2_P3_InstQueue_reg[3][0]/NET0131  & ~n50267 ;
  assign n64634 = n27788 & ~n64632 ;
  assign n64635 = ~n64633 & n64634 ;
  assign n64631 = \P2_P3_InstQueue_reg[3][0]/NET0131  & ~n50270 ;
  assign n64636 = \P2_buf2_reg[24]/NET0131  & n50021 ;
  assign n64637 = \P2_buf2_reg[16]/NET0131  & n50227 ;
  assign n64638 = ~n64636 & ~n64637 ;
  assign n64639 = n27325 & ~n64638 ;
  assign n64640 = \P2_buf2_reg[0]/NET0131  & n50280 ;
  assign n64641 = ~n64639 & ~n64640 ;
  assign n64642 = ~n64631 & n64641 ;
  assign n64643 = ~n64635 & n64642 ;
  assign n64646 = n26990 & n50267 ;
  assign n64645 = ~\P2_P3_InstQueue_reg[3][1]/NET0131  & ~n50267 ;
  assign n64647 = n27788 & ~n64645 ;
  assign n64648 = ~n64646 & n64647 ;
  assign n64644 = \P2_P3_InstQueue_reg[3][1]/NET0131  & ~n50270 ;
  assign n64649 = \P2_buf2_reg[25]/NET0131  & n50021 ;
  assign n64650 = \P2_buf2_reg[17]/NET0131  & n50227 ;
  assign n64651 = ~n64649 & ~n64650 ;
  assign n64652 = n27325 & ~n64651 ;
  assign n64653 = \P2_buf2_reg[1]/NET0131  & n50280 ;
  assign n64654 = ~n64652 & ~n64653 ;
  assign n64655 = ~n64644 & n64654 ;
  assign n64656 = ~n64648 & n64655 ;
  assign n64659 = n26990 & n50287 ;
  assign n64658 = ~\P2_P3_InstQueue_reg[4][1]/NET0131  & ~n50287 ;
  assign n64660 = n27788 & ~n64658 ;
  assign n64661 = ~n64659 & n64660 ;
  assign n64657 = \P2_P3_InstQueue_reg[4][1]/NET0131  & ~n50290 ;
  assign n64662 = \P2_buf2_reg[25]/NET0131  & n50227 ;
  assign n64663 = \P2_buf2_reg[17]/NET0131  & n50247 ;
  assign n64664 = ~n64662 & ~n64663 ;
  assign n64665 = n27325 & ~n64664 ;
  assign n64666 = \P2_buf2_reg[1]/NET0131  & n50300 ;
  assign n64667 = ~n64665 & ~n64666 ;
  assign n64668 = ~n64657 & n64667 ;
  assign n64669 = ~n64661 & n64668 ;
  assign n64672 = n26990 & n50307 ;
  assign n64671 = ~\P2_P3_InstQueue_reg[5][1]/NET0131  & ~n50307 ;
  assign n64673 = n27788 & ~n64671 ;
  assign n64674 = ~n64672 & n64673 ;
  assign n64670 = \P2_P3_InstQueue_reg[5][1]/NET0131  & ~n50310 ;
  assign n64675 = \P2_buf2_reg[25]/NET0131  & n50247 ;
  assign n64676 = \P2_buf2_reg[17]/NET0131  & n50267 ;
  assign n64677 = ~n64675 & ~n64676 ;
  assign n64678 = n27325 & ~n64677 ;
  assign n64679 = \P2_buf2_reg[1]/NET0131  & n50320 ;
  assign n64680 = ~n64678 & ~n64679 ;
  assign n64681 = ~n64670 & n64680 ;
  assign n64682 = ~n64674 & n64681 ;
  assign n64685 = n26990 & n50327 ;
  assign n64684 = ~\P2_P3_InstQueue_reg[6][1]/NET0131  & ~n50327 ;
  assign n64686 = n27788 & ~n64684 ;
  assign n64687 = ~n64685 & n64686 ;
  assign n64683 = \P2_P3_InstQueue_reg[6][1]/NET0131  & ~n50330 ;
  assign n64688 = \P2_buf2_reg[25]/NET0131  & n50267 ;
  assign n64689 = \P2_buf2_reg[17]/NET0131  & n50287 ;
  assign n64690 = ~n64688 & ~n64689 ;
  assign n64691 = n27325 & ~n64690 ;
  assign n64692 = \P2_buf2_reg[1]/NET0131  & n50340 ;
  assign n64693 = ~n64691 & ~n64692 ;
  assign n64694 = ~n64683 & n64693 ;
  assign n64695 = ~n64687 & n64694 ;
  assign n64698 = n27022 & n50046 ;
  assign n64697 = ~\P2_P3_InstQueue_reg[7][0]/NET0131  & ~n50046 ;
  assign n64699 = n27788 & ~n64697 ;
  assign n64700 = ~n64698 & n64699 ;
  assign n64696 = \P2_P3_InstQueue_reg[7][0]/NET0131  & ~n50349 ;
  assign n64701 = \P2_buf2_reg[24]/NET0131  & n50287 ;
  assign n64702 = \P2_buf2_reg[16]/NET0131  & n50307 ;
  assign n64703 = ~n64701 & ~n64702 ;
  assign n64704 = n27325 & ~n64703 ;
  assign n64705 = \P2_buf2_reg[0]/NET0131  & n50359 ;
  assign n64706 = ~n64704 & ~n64705 ;
  assign n64707 = ~n64696 & n64706 ;
  assign n64708 = ~n64700 & n64707 ;
  assign n64711 = n26990 & n50046 ;
  assign n64710 = ~\P2_P3_InstQueue_reg[7][1]/NET0131  & ~n50046 ;
  assign n64712 = n27788 & ~n64710 ;
  assign n64713 = ~n64711 & n64712 ;
  assign n64709 = \P2_P3_InstQueue_reg[7][1]/NET0131  & ~n50349 ;
  assign n64714 = \P2_buf2_reg[25]/NET0131  & n50287 ;
  assign n64715 = \P2_buf2_reg[17]/NET0131  & n50307 ;
  assign n64716 = ~n64714 & ~n64715 ;
  assign n64717 = n27325 & ~n64716 ;
  assign n64718 = \P2_buf2_reg[1]/NET0131  & n50359 ;
  assign n64719 = ~n64717 & ~n64718 ;
  assign n64720 = ~n64709 & n64719 ;
  assign n64721 = ~n64713 & n64720 ;
  assign n64724 = n26990 & n50045 ;
  assign n64723 = ~\P2_P3_InstQueue_reg[8][1]/NET0131  & ~n50045 ;
  assign n64725 = n27788 & ~n64723 ;
  assign n64726 = ~n64724 & n64725 ;
  assign n64722 = \P2_P3_InstQueue_reg[8][1]/NET0131  & ~n50367 ;
  assign n64727 = \P2_buf2_reg[25]/NET0131  & n50307 ;
  assign n64728 = \P2_buf2_reg[17]/NET0131  & n50327 ;
  assign n64729 = ~n64727 & ~n64728 ;
  assign n64730 = n27325 & ~n64729 ;
  assign n64731 = \P2_buf2_reg[1]/NET0131  & n50377 ;
  assign n64732 = ~n64730 & ~n64731 ;
  assign n64733 = ~n64722 & n64732 ;
  assign n64734 = ~n64726 & n64733 ;
  assign n64737 = n26990 & n50053 ;
  assign n64736 = ~\P2_P3_InstQueue_reg[9][1]/NET0131  & ~n50053 ;
  assign n64738 = n27788 & ~n64736 ;
  assign n64739 = ~n64737 & n64738 ;
  assign n64735 = \P2_P3_InstQueue_reg[9][1]/NET0131  & ~n50385 ;
  assign n64740 = \P2_buf2_reg[25]/NET0131  & n50327 ;
  assign n64741 = \P2_buf2_reg[17]/NET0131  & n50046 ;
  assign n64742 = ~n64740 & ~n64741 ;
  assign n64743 = n27325 & ~n64742 ;
  assign n64744 = \P2_buf2_reg[1]/NET0131  & n50395 ;
  assign n64745 = ~n64743 & ~n64744 ;
  assign n64746 = ~n64735 & n64745 ;
  assign n64747 = ~n64739 & n64746 ;
  assign n64750 = ~n8355 & n43284 ;
  assign n64751 = \P1_P1_InstQueueWr_Addr_reg[0]/NET0131  & ~n64750 ;
  assign n64748 = ~\P1_P1_Flush_reg/NET0131  & ~\P1_P1_InstQueueWr_Addr_reg[0]/NET0131  ;
  assign n64749 = n27623 & ~n64748 ;
  assign n64752 = ~n64186 & ~n64749 ;
  assign n64753 = ~n64751 & n64752 ;
  assign n64759 = ~\P2_P1_rEIP_reg[26]/NET0131  & ~n63466 ;
  assign n64760 = n25955 & ~n63467 ;
  assign n64761 = ~n64759 & n64760 ;
  assign n64754 = \P2_P1_Address_reg[24]/NET0131  & ~n25954 ;
  assign n64756 = ~\P2_P1_rEIP_reg[25]/NET0131  & ~n64047 ;
  assign n64755 = n50975 & n64047 ;
  assign n64757 = n63480 & ~n64755 ;
  assign n64758 = ~n64756 & n64757 ;
  assign n64762 = ~n64754 & ~n64758 ;
  assign n64763 = ~n64761 & n64762 ;
  assign n64770 = ~\P2_P2_rEIP_reg[26]/NET0131  & ~n63359 ;
  assign n64771 = n26647 & ~n63360 ;
  assign n64772 = ~n64770 & n64771 ;
  assign n64764 = \P2_P2_Address_reg[24]/NET0131  & ~n26646 ;
  assign n64765 = n52306 & n63987 ;
  assign n64767 = \P2_P2_rEIP_reg[25]/NET0131  & n64765 ;
  assign n64766 = ~\P2_P2_rEIP_reg[25]/NET0131  & ~n64765 ;
  assign n64768 = n63373 & ~n64766 ;
  assign n64769 = ~n64767 & n64768 ;
  assign n64773 = ~n64764 & ~n64769 ;
  assign n64774 = ~n64772 & n64773 ;
  assign n64776 = \P1_P1_rEIP_reg[24]/NET0131  & n63394 ;
  assign n64777 = \P1_P1_rEIP_reg[25]/NET0131  & n64776 ;
  assign n64778 = ~\P1_P1_rEIP_reg[26]/NET0131  & ~n64777 ;
  assign n64779 = n26155 & ~n63395 ;
  assign n64780 = ~n64778 & n64779 ;
  assign n64775 = \P1_P1_Address_reg[24]/NET0131  & ~n26154 ;
  assign n64781 = ~\P1_P1_rEIP_reg[25]/NET0131  & ~n63411 ;
  assign n64782 = n63401 & ~n63412 ;
  assign n64783 = ~n64781 & n64782 ;
  assign n64784 = ~n64775 & ~n64783 ;
  assign n64785 = ~n64780 & n64784 ;
  assign n64792 = ~\P1_P2_rEIP_reg[26]/NET0131  & ~n63440 ;
  assign n64793 = n25765 & ~n63441 ;
  assign n64794 = ~n64792 & n64793 ;
  assign n64786 = \P1_P2_Address_reg[24]/NET0131  & ~n25764 ;
  assign n64787 = n48386 & n63421 ;
  assign n64789 = ~n51408 & n64787 ;
  assign n64788 = ~\P1_P2_rEIP_reg[25]/NET0131  & ~n64787 ;
  assign n64790 = n63420 & ~n64788 ;
  assign n64791 = ~n64789 & n64790 ;
  assign n64795 = ~n64786 & ~n64791 ;
  assign n64796 = ~n64794 & n64795 ;
  assign n64798 = n50765 & n63461 ;
  assign n64799 = ~\P2_P1_rEIP_reg[14]/NET0131  & ~n64798 ;
  assign n64800 = n25955 & ~n63462 ;
  assign n64801 = ~n64799 & n64800 ;
  assign n64797 = \P2_P1_Address_reg[12]/NET0131  & ~n25954 ;
  assign n64802 = \P2_P1_rEIP_reg[12]/NET0131  & n64049 ;
  assign n64803 = ~\P2_P1_rEIP_reg[13]/NET0131  & ~n64802 ;
  assign n64804 = n50765 & n64049 ;
  assign n64805 = n63480 & ~n64804 ;
  assign n64806 = ~n64803 & n64805 ;
  assign n64807 = ~n64797 & ~n64806 ;
  assign n64808 = ~n64801 & n64807 ;
  assign n64814 = ~\P1_P1_rEIP_reg[14]/NET0131  & ~n63392 ;
  assign n64815 = n26155 & ~n63393 ;
  assign n64816 = ~n64814 & n64815 ;
  assign n64809 = \P1_P1_Address_reg[12]/NET0131  & ~n26154 ;
  assign n64810 = \P1_P1_rEIP_reg[12]/NET0131  & n63404 ;
  assign n64811 = ~\P1_P1_rEIP_reg[13]/NET0131  & ~n64810 ;
  assign n64812 = n63401 & ~n63405 ;
  assign n64813 = ~n64811 & n64812 ;
  assign n64817 = ~n64809 & ~n64813 ;
  assign n64818 = ~n64816 & n64817 ;
  assign n64820 = \P2_P2_rEIP_reg[9]/NET0131  & n63358 ;
  assign n64821 = n52105 & n64820 ;
  assign n64822 = n52104 & n64821 ;
  assign n64823 = ~\P2_P2_rEIP_reg[14]/NET0131  & ~n64822 ;
  assign n64824 = n26647 & ~n63998 ;
  assign n64825 = ~n64823 & n64824 ;
  assign n64819 = \P2_P2_Address_reg[12]/NET0131  & ~n26646 ;
  assign n64826 = \P2_P2_rEIP_reg[12]/NET0131  & n63989 ;
  assign n64827 = ~\P2_P2_rEIP_reg[13]/NET0131  & ~n64826 ;
  assign n64828 = n63373 & ~n63990 ;
  assign n64829 = ~n64827 & n64828 ;
  assign n64830 = ~n64819 & ~n64829 ;
  assign n64831 = ~n64825 & n64830 ;
  assign n64833 = ~\P1_P3_rEIP_reg[14]/NET0131  & ~n64072 ;
  assign n64834 = n9092 & ~n64073 ;
  assign n64835 = ~n64833 & n64834 ;
  assign n64832 = \P1_P3_Address_reg[12]/NET0131  & ~n9091 ;
  assign n64836 = ~\P1_P3_rEIP_reg[13]/NET0131  & ~n64082 ;
  assign n64837 = n22115 & ~n64083 ;
  assign n64838 = ~n64836 & n64837 ;
  assign n64839 = ~n64832 & ~n64838 ;
  assign n64840 = ~n64835 & n64839 ;
  assign n64842 = n48390 & n64032 ;
  assign n64843 = ~\P1_P2_rEIP_reg[14]/NET0131  & ~n64842 ;
  assign n64844 = \P1_P2_rEIP_reg[10]/NET0131  & n64031 ;
  assign n64845 = n64022 & n64844 ;
  assign n64846 = n25765 & ~n64845 ;
  assign n64847 = ~n64843 & n64846 ;
  assign n64841 = \P1_P2_Address_reg[12]/NET0131  & ~n25764 ;
  assign n64848 = n48393 & n64787 ;
  assign n64849 = \P1_P2_rEIP_reg[12]/NET0131  & n64848 ;
  assign n64851 = \P1_P2_rEIP_reg[13]/NET0131  & n64849 ;
  assign n64850 = ~\P1_P2_rEIP_reg[13]/NET0131  & ~n64849 ;
  assign n64852 = n63420 & ~n64850 ;
  assign n64853 = ~n64851 & n64852 ;
  assign n64854 = ~n64841 & ~n64853 ;
  assign n64855 = ~n64847 & n64854 ;
  assign n64857 = ~\P2_P3_rEIP_reg[14]/NET0131  & ~n64114 ;
  assign n64858 = n27145 & ~n64115 ;
  assign n64859 = ~n64857 & n64858 ;
  assign n64856 = \P2_P3_Address_reg[12]/NET0131  & ~n27144 ;
  assign n64860 = n52557 & n64095 ;
  assign n64862 = ~\P2_P3_rEIP_reg[13]/NET0131  & ~n64860 ;
  assign n64861 = \P2_P3_rEIP_reg[13]/NET0131  & n64860 ;
  assign n64863 = n64094 & ~n64861 ;
  assign n64864 = ~n64862 & n64863 ;
  assign n64865 = ~n64856 & ~n64864 ;
  assign n64866 = ~n64859 & n64865 ;
  assign n64869 = n27022 & n50327 ;
  assign n64868 = ~\P2_P3_InstQueue_reg[6][0]/NET0131  & ~n50327 ;
  assign n64870 = n27788 & ~n64868 ;
  assign n64871 = ~n64869 & n64870 ;
  assign n64867 = \P2_P3_InstQueue_reg[6][0]/NET0131  & ~n50330 ;
  assign n64872 = \P2_buf2_reg[24]/NET0131  & n50267 ;
  assign n64873 = \P2_buf2_reg[16]/NET0131  & n50287 ;
  assign n64874 = ~n64872 & ~n64873 ;
  assign n64875 = n27325 & ~n64874 ;
  assign n64876 = \P2_buf2_reg[0]/NET0131  & n50340 ;
  assign n64877 = ~n64875 & ~n64876 ;
  assign n64878 = ~n64867 & n64877 ;
  assign n64879 = ~n64871 & n64878 ;
  assign n64882 = n8924 & n49732 ;
  assign n64881 = ~\P1_P3_InstQueue_reg[0][0]/NET0131  & ~n49732 ;
  assign n64883 = n10046 & ~n64881 ;
  assign n64884 = ~n64882 & n64883 ;
  assign n64880 = \P1_P3_InstQueue_reg[0][0]/NET0131  & ~n49750 ;
  assign n64885 = \P1_buf2_reg[24]/NET0131  & n49739 ;
  assign n64886 = \P1_buf2_reg[16]/NET0131  & ~n49739 ;
  assign n64887 = n49742 & n64886 ;
  assign n64888 = ~n64885 & ~n64887 ;
  assign n64889 = n11698 & ~n64888 ;
  assign n64890 = \P1_buf2_reg[0]/NET0131  & n49760 ;
  assign n64891 = ~n64889 & ~n64890 ;
  assign n64892 = ~n64880 & n64891 ;
  assign n64893 = ~n64884 & n64892 ;
  assign n64896 = n8924 & n49766 ;
  assign n64895 = ~\P1_P3_InstQueue_reg[10][0]/NET0131  & ~n49766 ;
  assign n64897 = n10046 & ~n64895 ;
  assign n64898 = ~n64896 & n64897 ;
  assign n64894 = \P1_P3_InstQueue_reg[10][0]/NET0131  & ~n49776 ;
  assign n64899 = \P1_buf2_reg[24]/NET0131  & n49770 ;
  assign n64900 = \P1_buf2_reg[16]/NET0131  & n49771 ;
  assign n64901 = ~n64899 & ~n64900 ;
  assign n64902 = n11698 & ~n64901 ;
  assign n64903 = \P1_buf2_reg[0]/NET0131  & n49786 ;
  assign n64904 = ~n64902 & ~n64903 ;
  assign n64905 = ~n64894 & n64904 ;
  assign n64906 = ~n64898 & n64905 ;
  assign n64909 = n8924 & n49814 ;
  assign n64908 = ~\P1_P3_InstQueue_reg[12][0]/NET0131  & ~n49814 ;
  assign n64910 = n10046 & ~n64908 ;
  assign n64911 = ~n64909 & n64910 ;
  assign n64907 = \P1_P3_InstQueue_reg[12][0]/NET0131  & ~n49819 ;
  assign n64912 = \P1_buf2_reg[24]/NET0131  & n49768 ;
  assign n64913 = \P1_buf2_reg[16]/NET0131  & n49766 ;
  assign n64914 = ~n64912 & ~n64913 ;
  assign n64915 = n11698 & ~n64914 ;
  assign n64916 = \P1_buf2_reg[0]/NET0131  & n49829 ;
  assign n64917 = ~n64915 & ~n64916 ;
  assign n64918 = ~n64907 & n64917 ;
  assign n64919 = ~n64911 & n64918 ;
  assign n64922 = n8924 & n49739 ;
  assign n64921 = ~\P1_P3_InstQueue_reg[13][0]/NET0131  & ~n49739 ;
  assign n64923 = n10046 & ~n64921 ;
  assign n64924 = ~n64922 & n64923 ;
  assign n64920 = \P1_P3_InstQueue_reg[13][0]/NET0131  & ~n49838 ;
  assign n64925 = \P1_buf2_reg[24]/NET0131  & n49766 ;
  assign n64926 = \P1_buf2_reg[16]/NET0131  & ~n49766 ;
  assign n64927 = n49792 & n64926 ;
  assign n64928 = ~n64925 & ~n64927 ;
  assign n64929 = n11698 & ~n64928 ;
  assign n64930 = \P1_buf2_reg[0]/NET0131  & n49848 ;
  assign n64931 = ~n64929 & ~n64930 ;
  assign n64932 = ~n64920 & n64931 ;
  assign n64933 = ~n64924 & n64932 ;
  assign n64936 = n8924 & n49742 ;
  assign n64935 = ~\P1_P3_InstQueue_reg[14][0]/NET0131  & ~n49742 ;
  assign n64937 = n10046 & ~n64935 ;
  assign n64938 = ~n64936 & n64937 ;
  assign n64934 = \P1_P3_InstQueue_reg[14][0]/NET0131  & ~n49856 ;
  assign n64939 = \P1_buf2_reg[24]/NET0131  & n49792 ;
  assign n64940 = \P1_buf2_reg[16]/NET0131  & ~n49792 ;
  assign n64941 = n49814 & n64940 ;
  assign n64942 = ~n64939 & ~n64941 ;
  assign n64943 = n11698 & ~n64942 ;
  assign n64944 = \P1_buf2_reg[0]/NET0131  & n49866 ;
  assign n64945 = ~n64943 & ~n64944 ;
  assign n64946 = ~n64934 & n64945 ;
  assign n64947 = ~n64938 & n64946 ;
  assign n64950 = n8924 & n49735 ;
  assign n64949 = ~\P1_P3_InstQueue_reg[15][0]/NET0131  & ~n49735 ;
  assign n64951 = n10046 & ~n64949 ;
  assign n64952 = ~n64950 & n64951 ;
  assign n64948 = \P1_P3_InstQueue_reg[15][0]/NET0131  & ~n49875 ;
  assign n64953 = \P1_buf2_reg[24]/NET0131  & n49814 ;
  assign n64954 = \P1_buf2_reg[16]/NET0131  & n49739 ;
  assign n64955 = ~n64953 & ~n64954 ;
  assign n64956 = n11698 & ~n64955 ;
  assign n64957 = \P1_buf2_reg[0]/NET0131  & n49885 ;
  assign n64958 = ~n64956 & ~n64957 ;
  assign n64959 = ~n64948 & n64958 ;
  assign n64960 = ~n64952 & n64959 ;
  assign n64963 = n8924 & n49890 ;
  assign n64962 = ~\P1_P3_InstQueue_reg[1][0]/NET0131  & ~n49890 ;
  assign n64964 = n10046 & ~n64962 ;
  assign n64965 = ~n64963 & n64964 ;
  assign n64961 = \P1_P3_InstQueue_reg[1][0]/NET0131  & ~n49895 ;
  assign n64966 = \P1_buf2_reg[24]/NET0131  & n49742 ;
  assign n64967 = \P1_buf2_reg[16]/NET0131  & n49735 ;
  assign n64968 = ~n64966 & ~n64967 ;
  assign n64969 = n11698 & ~n64968 ;
  assign n64970 = \P1_buf2_reg[0]/NET0131  & n49905 ;
  assign n64971 = ~n64969 & ~n64970 ;
  assign n64972 = ~n64961 & n64971 ;
  assign n64973 = ~n64965 & n64972 ;
  assign n64976 = n8924 & n49910 ;
  assign n64975 = ~\P1_P3_InstQueue_reg[2][0]/NET0131  & ~n49910 ;
  assign n64977 = n10046 & ~n64975 ;
  assign n64978 = ~n64976 & n64977 ;
  assign n64974 = \P1_P3_InstQueue_reg[2][0]/NET0131  & ~n49915 ;
  assign n64979 = \P1_buf2_reg[24]/NET0131  & n49735 ;
  assign n64980 = \P1_buf2_reg[16]/NET0131  & n49732 ;
  assign n64981 = ~n64979 & ~n64980 ;
  assign n64982 = n11698 & ~n64981 ;
  assign n64983 = \P1_buf2_reg[0]/NET0131  & n49925 ;
  assign n64984 = ~n64982 & ~n64983 ;
  assign n64985 = ~n64974 & n64984 ;
  assign n64986 = ~n64978 & n64985 ;
  assign n64989 = n8924 & n49950 ;
  assign n64988 = ~\P1_P3_InstQueue_reg[4][0]/NET0131  & ~n49950 ;
  assign n64990 = n10046 & ~n64988 ;
  assign n64991 = ~n64989 & n64990 ;
  assign n64987 = \P1_P3_InstQueue_reg[4][0]/NET0131  & ~n49955 ;
  assign n64992 = \P1_buf2_reg[24]/NET0131  & n49890 ;
  assign n64993 = \P1_buf2_reg[16]/NET0131  & ~n49890 ;
  assign n64994 = n49910 & n64993 ;
  assign n64995 = ~n64992 & ~n64994 ;
  assign n64996 = n11698 & ~n64995 ;
  assign n64997 = \P1_buf2_reg[0]/NET0131  & n49965 ;
  assign n64998 = ~n64996 & ~n64997 ;
  assign n64999 = ~n64987 & n64998 ;
  assign n65000 = ~n64991 & n64999 ;
  assign n65003 = n8924 & n49970 ;
  assign n65002 = ~\P1_P3_InstQueue_reg[5][0]/NET0131  & ~n49970 ;
  assign n65004 = n10046 & ~n65002 ;
  assign n65005 = ~n65003 & n65004 ;
  assign n65001 = \P1_P3_InstQueue_reg[5][0]/NET0131  & ~n49975 ;
  assign n65006 = \P1_buf2_reg[24]/NET0131  & n49910 ;
  assign n65007 = \P1_buf2_reg[16]/NET0131  & ~n49910 ;
  assign n65008 = n49930 & n65007 ;
  assign n65009 = ~n65006 & ~n65008 ;
  assign n65010 = n11698 & ~n65009 ;
  assign n65011 = \P1_buf2_reg[0]/NET0131  & n49985 ;
  assign n65012 = ~n65010 & ~n65011 ;
  assign n65013 = ~n65001 & n65012 ;
  assign n65014 = ~n65005 & n65013 ;
  assign n65017 = n8924 & n49990 ;
  assign n65016 = ~\P1_P3_InstQueue_reg[6][0]/NET0131  & ~n49990 ;
  assign n65018 = n10046 & ~n65016 ;
  assign n65019 = ~n65017 & n65018 ;
  assign n65015 = \P1_P3_InstQueue_reg[6][0]/NET0131  & ~n49995 ;
  assign n65020 = \P1_buf2_reg[24]/NET0131  & n49930 ;
  assign n65021 = \P1_buf2_reg[16]/NET0131  & ~n49930 ;
  assign n65022 = n49950 & n65021 ;
  assign n65023 = ~n65020 & ~n65022 ;
  assign n65024 = n11698 & ~n65023 ;
  assign n65025 = \P1_buf2_reg[0]/NET0131  & n50005 ;
  assign n65026 = ~n65024 & ~n65025 ;
  assign n65027 = ~n65015 & n65026 ;
  assign n65028 = ~n65019 & n65027 ;
  assign n65031 = n27022 & n50021 ;
  assign n65030 = ~\P2_P3_InstQueue_reg[0][0]/NET0131  & ~n50021 ;
  assign n65032 = n27788 & ~n65030 ;
  assign n65033 = ~n65031 & n65032 ;
  assign n65029 = \P2_P3_InstQueue_reg[0][0]/NET0131  & ~n50030 ;
  assign n65034 = \P2_buf2_reg[24]/NET0131  & n50012 ;
  assign n65035 = \P2_buf2_reg[16]/NET0131  & n50015 ;
  assign n65036 = ~n65034 & ~n65035 ;
  assign n65037 = n27325 & ~n65036 ;
  assign n65038 = \P2_buf2_reg[0]/NET0131  & n50040 ;
  assign n65039 = ~n65037 & ~n65038 ;
  assign n65040 = ~n65029 & n65039 ;
  assign n65041 = ~n65033 & n65040 ;
  assign n65044 = n27022 & n50051 ;
  assign n65043 = ~\P2_P3_InstQueue_reg[10][0]/NET0131  & ~n50051 ;
  assign n65045 = n27788 & ~n65043 ;
  assign n65046 = ~n65044 & n65045 ;
  assign n65042 = \P2_P3_InstQueue_reg[10][0]/NET0131  & ~n50056 ;
  assign n65047 = \P2_buf2_reg[16]/NET0131  & n50045 ;
  assign n65048 = \P2_buf2_reg[24]/NET0131  & n50046 ;
  assign n65049 = ~n65047 & ~n65048 ;
  assign n65050 = n27325 & ~n65049 ;
  assign n65051 = \P2_buf2_reg[0]/NET0131  & n50066 ;
  assign n65052 = ~n65050 & ~n65051 ;
  assign n65053 = ~n65042 & n65052 ;
  assign n65054 = ~n65046 & n65053 ;
  assign n65057 = n27022 & n50115 ;
  assign n65056 = ~\P2_P3_InstQueue_reg[12][0]/NET0131  & ~n50115 ;
  assign n65058 = n27788 & ~n65056 ;
  assign n65059 = ~n65057 & n65058 ;
  assign n65055 = \P2_P3_InstQueue_reg[12][0]/NET0131  & ~n50118 ;
  assign n65060 = \P2_buf2_reg[24]/NET0131  & n50053 ;
  assign n65061 = \P2_buf2_reg[16]/NET0131  & n50051 ;
  assign n65062 = ~n65060 & ~n65061 ;
  assign n65063 = n27325 & ~n65062 ;
  assign n65064 = \P2_buf2_reg[0]/NET0131  & n50128 ;
  assign n65065 = ~n65063 & ~n65064 ;
  assign n65066 = ~n65055 & n65065 ;
  assign n65067 = ~n65059 & n65066 ;
  assign n65070 = n8924 & n49771 ;
  assign n65069 = ~\P1_P3_InstQueue_reg[8][0]/NET0131  & ~n49771 ;
  assign n65071 = n10046 & ~n65069 ;
  assign n65072 = ~n65070 & n65071 ;
  assign n65068 = \P1_P3_InstQueue_reg[8][0]/NET0131  & ~n50136 ;
  assign n65073 = \P1_buf2_reg[24]/NET0131  & n49970 ;
  assign n65074 = \P1_buf2_reg[16]/NET0131  & ~n49970 ;
  assign n65075 = n49990 & n65074 ;
  assign n65076 = ~n65073 & ~n65075 ;
  assign n65077 = n11698 & ~n65076 ;
  assign n65078 = \P1_buf2_reg[0]/NET0131  & n50146 ;
  assign n65079 = ~n65077 & ~n65078 ;
  assign n65080 = ~n65068 & n65079 ;
  assign n65081 = ~n65072 & n65080 ;
  assign n65084 = n27022 & n50012 ;
  assign n65083 = ~\P2_P3_InstQueue_reg[13][0]/NET0131  & ~n50012 ;
  assign n65085 = n27788 & ~n65083 ;
  assign n65086 = ~n65084 & n65085 ;
  assign n65082 = \P2_P3_InstQueue_reg[13][0]/NET0131  & ~n50155 ;
  assign n65087 = \P2_buf2_reg[24]/NET0131  & n50051 ;
  assign n65088 = \P2_buf2_reg[16]/NET0131  & n50094 ;
  assign n65089 = ~n65087 & ~n65088 ;
  assign n65090 = n27325 & ~n65089 ;
  assign n65091 = \P2_buf2_reg[0]/NET0131  & n50165 ;
  assign n65092 = ~n65090 & ~n65091 ;
  assign n65093 = ~n65082 & n65092 ;
  assign n65094 = ~n65086 & n65093 ;
  assign n65097 = n27022 & n50015 ;
  assign n65096 = ~\P2_P3_InstQueue_reg[14][0]/NET0131  & ~n50015 ;
  assign n65098 = n27788 & ~n65096 ;
  assign n65099 = ~n65097 & n65098 ;
  assign n65095 = \P2_P3_InstQueue_reg[14][0]/NET0131  & ~n50173 ;
  assign n65100 = \P2_buf2_reg[24]/NET0131  & n50094 ;
  assign n65101 = \P2_buf2_reg[16]/NET0131  & n50115 ;
  assign n65102 = ~n65100 & ~n65101 ;
  assign n65103 = n27325 & ~n65102 ;
  assign n65104 = \P2_buf2_reg[0]/NET0131  & n50183 ;
  assign n65105 = ~n65103 & ~n65104 ;
  assign n65106 = ~n65095 & n65105 ;
  assign n65107 = ~n65099 & n65106 ;
  assign n65110 = n8924 & n49768 ;
  assign n65109 = ~\P1_P3_InstQueue_reg[9][0]/NET0131  & ~n49768 ;
  assign n65111 = n10046 & ~n65109 ;
  assign n65112 = ~n65110 & n65111 ;
  assign n65108 = \P1_P3_InstQueue_reg[9][0]/NET0131  & ~n50191 ;
  assign n65113 = \P1_buf2_reg[24]/NET0131  & n49990 ;
  assign n65114 = \P1_buf2_reg[16]/NET0131  & n49770 ;
  assign n65115 = ~n65113 & ~n65114 ;
  assign n65116 = n11698 & ~n65115 ;
  assign n65117 = \P1_buf2_reg[0]/NET0131  & n50201 ;
  assign n65118 = ~n65116 & ~n65117 ;
  assign n65119 = ~n65108 & n65118 ;
  assign n65120 = ~n65112 & n65119 ;
  assign n65123 = n27022 & n50024 ;
  assign n65122 = ~\P2_P3_InstQueue_reg[15][0]/NET0131  & ~n50024 ;
  assign n65124 = n27788 & ~n65122 ;
  assign n65125 = ~n65123 & n65124 ;
  assign n65121 = \P2_P3_InstQueue_reg[15][0]/NET0131  & ~n50210 ;
  assign n65126 = \P2_buf2_reg[24]/NET0131  & n50115 ;
  assign n65127 = \P2_buf2_reg[16]/NET0131  & n50012 ;
  assign n65128 = ~n65126 & ~n65127 ;
  assign n65129 = n27325 & ~n65128 ;
  assign n65130 = \P2_buf2_reg[0]/NET0131  & n50220 ;
  assign n65131 = ~n65129 & ~n65130 ;
  assign n65132 = ~n65121 & n65131 ;
  assign n65133 = ~n65125 & n65132 ;
  assign n65136 = n27022 & n50227 ;
  assign n65135 = ~\P2_P3_InstQueue_reg[1][0]/NET0131  & ~n50227 ;
  assign n65137 = n27788 & ~n65135 ;
  assign n65138 = ~n65136 & n65137 ;
  assign n65134 = \P2_P3_InstQueue_reg[1][0]/NET0131  & ~n50230 ;
  assign n65139 = \P2_buf2_reg[24]/NET0131  & n50015 ;
  assign n65140 = \P2_buf2_reg[16]/NET0131  & n50024 ;
  assign n65141 = ~n65139 & ~n65140 ;
  assign n65142 = n27325 & ~n65141 ;
  assign n65143 = \P2_buf2_reg[0]/NET0131  & n50240 ;
  assign n65144 = ~n65142 & ~n65143 ;
  assign n65145 = ~n65134 & n65144 ;
  assign n65146 = ~n65138 & n65145 ;
  assign n65149 = n27022 & n50287 ;
  assign n65148 = ~\P2_P3_InstQueue_reg[4][0]/NET0131  & ~n50287 ;
  assign n65150 = n27788 & ~n65148 ;
  assign n65151 = ~n65149 & n65150 ;
  assign n65147 = \P2_P3_InstQueue_reg[4][0]/NET0131  & ~n50290 ;
  assign n65152 = \P2_buf2_reg[24]/NET0131  & n50227 ;
  assign n65153 = \P2_buf2_reg[16]/NET0131  & n50247 ;
  assign n65154 = ~n65152 & ~n65153 ;
  assign n65155 = n27325 & ~n65154 ;
  assign n65156 = \P2_buf2_reg[0]/NET0131  & n50300 ;
  assign n65157 = ~n65155 & ~n65156 ;
  assign n65158 = ~n65147 & n65157 ;
  assign n65159 = ~n65151 & n65158 ;
  assign n65162 = n27022 & n50307 ;
  assign n65161 = ~\P2_P3_InstQueue_reg[5][0]/NET0131  & ~n50307 ;
  assign n65163 = n27788 & ~n65161 ;
  assign n65164 = ~n65162 & n65163 ;
  assign n65160 = \P2_P3_InstQueue_reg[5][0]/NET0131  & ~n50310 ;
  assign n65165 = \P2_buf2_reg[24]/NET0131  & n50247 ;
  assign n65166 = \P2_buf2_reg[16]/NET0131  & n50267 ;
  assign n65167 = ~n65165 & ~n65166 ;
  assign n65168 = n27325 & ~n65167 ;
  assign n65169 = \P2_buf2_reg[0]/NET0131  & n50320 ;
  assign n65170 = ~n65168 & ~n65169 ;
  assign n65171 = ~n65160 & n65170 ;
  assign n65172 = ~n65164 & n65171 ;
  assign n65175 = n27022 & n50045 ;
  assign n65174 = ~\P2_P3_InstQueue_reg[8][0]/NET0131  & ~n50045 ;
  assign n65176 = n27788 & ~n65174 ;
  assign n65177 = ~n65175 & n65176 ;
  assign n65173 = \P2_P3_InstQueue_reg[8][0]/NET0131  & ~n50367 ;
  assign n65178 = \P2_buf2_reg[24]/NET0131  & n50307 ;
  assign n65179 = \P2_buf2_reg[16]/NET0131  & n50327 ;
  assign n65180 = ~n65178 & ~n65179 ;
  assign n65181 = n27325 & ~n65180 ;
  assign n65182 = \P2_buf2_reg[0]/NET0131  & n50377 ;
  assign n65183 = ~n65181 & ~n65182 ;
  assign n65184 = ~n65173 & n65183 ;
  assign n65185 = ~n65177 & n65184 ;
  assign n65188 = n27022 & n50053 ;
  assign n65187 = ~\P2_P3_InstQueue_reg[9][0]/NET0131  & ~n50053 ;
  assign n65189 = n27788 & ~n65187 ;
  assign n65190 = ~n65188 & n65189 ;
  assign n65186 = \P2_P3_InstQueue_reg[9][0]/NET0131  & ~n50385 ;
  assign n65191 = \P2_buf2_reg[24]/NET0131  & n50327 ;
  assign n65192 = \P2_buf2_reg[16]/NET0131  & n50046 ;
  assign n65193 = ~n65191 & ~n65192 ;
  assign n65194 = n27325 & ~n65193 ;
  assign n65195 = \P2_buf2_reg[0]/NET0131  & n50395 ;
  assign n65196 = ~n65194 & ~n65195 ;
  assign n65197 = ~n65186 & n65196 ;
  assign n65198 = ~n65190 & n65197 ;
  assign n65201 = n27022 & n50247 ;
  assign n65200 = ~\P2_P3_InstQueue_reg[2][0]/NET0131  & ~n50247 ;
  assign n65202 = n27788 & ~n65200 ;
  assign n65203 = ~n65201 & n65202 ;
  assign n65199 = \P2_P3_InstQueue_reg[2][0]/NET0131  & ~n50250 ;
  assign n65204 = \P2_buf2_reg[16]/NET0131  & n50021 ;
  assign n65205 = \P2_buf2_reg[24]/NET0131  & n50024 ;
  assign n65206 = ~n65204 & ~n65205 ;
  assign n65207 = n27325 & ~n65206 ;
  assign n65208 = \P2_buf2_reg[0]/NET0131  & n50260 ;
  assign n65209 = ~n65207 & ~n65208 ;
  assign n65210 = ~n65199 & n65209 ;
  assign n65211 = ~n65203 & n65210 ;
  assign n65217 = \P2_P1_rEIP_reg[21]/NET0131  & n63464 ;
  assign n65219 = \P2_P1_rEIP_reg[22]/NET0131  & n65217 ;
  assign n65218 = ~\P2_P1_rEIP_reg[22]/NET0131  & ~n65217 ;
  assign n65220 = n25955 & ~n65218 ;
  assign n65221 = ~n65219 & n65220 ;
  assign n65212 = \P2_P1_Address_reg[20]/NET0131  & ~n25954 ;
  assign n65214 = ~n50836 & n63475 ;
  assign n65213 = ~\P2_P1_rEIP_reg[21]/NET0131  & ~n63475 ;
  assign n65215 = n63480 & ~n65213 ;
  assign n65216 = ~n65214 & n65215 ;
  assign n65222 = ~n65212 & ~n65216 ;
  assign n65223 = ~n65221 & n65222 ;
  assign n65225 = n52103 & n63991 ;
  assign n65226 = \P2_P2_rEIP_reg[20]/NET0131  & n65225 ;
  assign n65228 = \P2_P2_rEIP_reg[21]/NET0131  & n65226 ;
  assign n65227 = ~\P2_P2_rEIP_reg[21]/NET0131  & ~n65226 ;
  assign n65229 = n63373 & ~n65227 ;
  assign n65230 = ~n65228 & n65229 ;
  assign n65224 = \P2_P2_Address_reg[20]/NET0131  & ~n26646 ;
  assign n65231 = n52305 & n63358 ;
  assign n65233 = ~\P2_P2_rEIP_reg[22]/NET0131  & ~n65231 ;
  assign n65232 = \P2_P2_rEIP_reg[22]/NET0131  & n65231 ;
  assign n65234 = n26647 & ~n65232 ;
  assign n65235 = ~n65233 & n65234 ;
  assign n65236 = ~n65224 & ~n65235 ;
  assign n65237 = ~n65230 & n65236 ;
  assign n65244 = n51682 & n63402 ;
  assign n65245 = ~\P1_P1_rEIP_reg[21]/NET0131  & ~n65244 ;
  assign n65246 = n51737 & n63402 ;
  assign n65247 = n63401 & ~n65246 ;
  assign n65248 = ~n65245 & n65247 ;
  assign n65238 = \P1_P1_Address_reg[20]/NET0131  & ~n26154 ;
  assign n65239 = n51736 & n63393 ;
  assign n65240 = ~\P1_P1_rEIP_reg[22]/NET0131  & ~n65239 ;
  assign n65241 = n51844 & n63393 ;
  assign n65242 = n26155 & ~n65241 ;
  assign n65243 = ~n65240 & n65242 ;
  assign n65249 = ~n65238 & ~n65243 ;
  assign n65250 = ~n65248 & n65249 ;
  assign n65254 = n51238 & n64028 ;
  assign n65255 = ~\P1_P2_rEIP_reg[21]/NET0131  & ~n65254 ;
  assign n65252 = n48389 & n64024 ;
  assign n65253 = n48378 & n65252 ;
  assign n65256 = n63420 & ~n65253 ;
  assign n65257 = ~n65255 & n65256 ;
  assign n65251 = \P1_P2_Address_reg[20]/NET0131  & ~n25764 ;
  assign n65258 = ~\P1_P2_rEIP_reg[22]/NET0131  & ~n63438 ;
  assign n65259 = n25765 & ~n63439 ;
  assign n65260 = ~n65258 & n65259 ;
  assign n65261 = ~n65251 & ~n65260 ;
  assign n65262 = ~n65257 & n65261 ;
  assign n65265 = ~\P2_P2_rEIP_reg[10]/NET0131  & ~n64820 ;
  assign n65264 = \P2_P2_rEIP_reg[10]/NET0131  & n64820 ;
  assign n65266 = n26647 & ~n65264 ;
  assign n65267 = ~n65265 & n65266 ;
  assign n65263 = \P2_P2_Address_reg[8]/NET0131  & ~n26646 ;
  assign n65268 = ~\P2_P2_rEIP_reg[9]/NET0131  & ~n63987 ;
  assign n65269 = n63373 & ~n63988 ;
  assign n65270 = ~n65268 & n65269 ;
  assign n65271 = ~n65263 & ~n65270 ;
  assign n65272 = ~n65267 & n65271 ;
  assign n65278 = ~\P1_P3_rEIP_reg[10]/NET0131  & ~n64068 ;
  assign n65279 = n9092 & ~n64069 ;
  assign n65280 = ~n65278 & n65279 ;
  assign n65273 = \P1_P3_Address_reg[8]/NET0131  & ~n9091 ;
  assign n65275 = ~n17916 & n64081 ;
  assign n65274 = ~\P1_P3_rEIP_reg[9]/NET0131  & ~n64081 ;
  assign n65276 = n22115 & ~n65274 ;
  assign n65277 = ~n65275 & n65276 ;
  assign n65281 = ~n65273 & ~n65277 ;
  assign n65282 = ~n65280 & n65281 ;
  assign n65284 = ~\P1_P1_rEIP_reg[10]/NET0131  & ~n63389 ;
  assign n65285 = n26155 & ~n63390 ;
  assign n65286 = ~n65284 & n65285 ;
  assign n65283 = \P1_P1_Address_reg[8]/NET0131  & ~n26154 ;
  assign n65287 = n51670 & n63402 ;
  assign n65288 = \P1_P1_rEIP_reg[7]/NET0131  & n65287 ;
  assign n65289 = \P1_P1_rEIP_reg[8]/NET0131  & n65288 ;
  assign n65291 = ~\P1_P1_rEIP_reg[9]/NET0131  & ~n65289 ;
  assign n65290 = \P1_P1_rEIP_reg[9]/NET0131  & n65289 ;
  assign n65292 = n63401 & ~n65290 ;
  assign n65293 = ~n65291 & n65292 ;
  assign n65294 = ~n65283 & ~n65293 ;
  assign n65295 = ~n65286 & n65294 ;
  assign n65297 = ~\P2_P3_rEIP_reg[10]/NET0131  & ~n64110 ;
  assign n65298 = n27145 & ~n64111 ;
  assign n65299 = ~n65297 & n65298 ;
  assign n65296 = \P2_P3_Address_reg[8]/NET0131  & ~n27144 ;
  assign n65300 = n52551 & n64095 ;
  assign n65301 = \P2_P3_rEIP_reg[7]/NET0131  & n65300 ;
  assign n65302 = \P2_P3_rEIP_reg[8]/NET0131  & n65301 ;
  assign n65304 = ~\P2_P3_rEIP_reg[9]/NET0131  & ~n65302 ;
  assign n65303 = \P2_P3_rEIP_reg[9]/NET0131  & n65302 ;
  assign n65305 = n64094 & ~n65303 ;
  assign n65306 = ~n65304 & n65305 ;
  assign n65307 = ~n65296 & ~n65306 ;
  assign n65308 = ~n65299 & n65307 ;
  assign n65310 = ~\P1_P2_rEIP_reg[10]/NET0131  & ~n64031 ;
  assign n65311 = n25765 & ~n64844 ;
  assign n65312 = ~n65310 & n65311 ;
  assign n65309 = \P1_P2_Address_reg[8]/NET0131  & ~n25764 ;
  assign n65314 = n51239 & n63421 ;
  assign n65313 = ~\P1_P2_rEIP_reg[9]/NET0131  & ~n64787 ;
  assign n65315 = n63420 & ~n65313 ;
  assign n65316 = ~n65314 & n65315 ;
  assign n65317 = ~n65309 & ~n65316 ;
  assign n65318 = ~n65312 & n65317 ;
  assign n65321 = ~\P2_P1_rEIP_reg[10]/NET0131  & ~n63460 ;
  assign n65320 = \P2_P1_rEIP_reg[10]/NET0131  & n63460 ;
  assign n65322 = n25955 & ~n65320 ;
  assign n65323 = ~n65321 & n65322 ;
  assign n65319 = \P2_P1_Address_reg[8]/NET0131  & ~n25954 ;
  assign n65324 = ~\P2_P1_rEIP_reg[9]/NET0131  & ~n64047 ;
  assign n65325 = n63480 & ~n64048 ;
  assign n65326 = ~n65324 & n65325 ;
  assign n65327 = ~n65319 & ~n65326 ;
  assign n65328 = ~n65323 & n65327 ;
  assign n65329 = \P3_rd_reg/NET0131  & \P4_IR_reg[28]/NET0131  ;
  assign n65330 = \P2_P3_Datao_reg[28]/NET0131  & ~\P3_rd_reg/NET0131  ;
  assign n65331 = ~n65329 & ~n65330 ;
  assign n65333 = ~\P2_P2_rEIP_reg[6]/NET0131  & ~n63355 ;
  assign n65334 = n26647 & ~n63356 ;
  assign n65335 = ~n65333 & n65334 ;
  assign n65332 = \P2_P2_Address_reg[4]/NET0131  & ~n26646 ;
  assign n65336 = \P2_P2_rEIP_reg[1]/NET0131  & n63368 ;
  assign n65337 = \P2_P2_rEIP_reg[2]/NET0131  & n65336 ;
  assign n65338 = \P2_P2_rEIP_reg[3]/NET0131  & n65337 ;
  assign n65339 = \P2_P2_rEIP_reg[4]/NET0131  & n65338 ;
  assign n65341 = ~\P2_P2_rEIP_reg[5]/NET0131  & ~n65339 ;
  assign n65340 = \P2_P2_rEIP_reg[5]/NET0131  & n65339 ;
  assign n65342 = n63373 & ~n65340 ;
  assign n65343 = ~n65341 & n65342 ;
  assign n65344 = ~n65332 & ~n65343 ;
  assign n65345 = ~n65335 & n65344 ;
  assign n65355 = ~\P1_P3_rEIP_reg[6]/NET0131  & ~n64064 ;
  assign n65356 = n9092 & ~n64065 ;
  assign n65357 = ~n65355 & n65356 ;
  assign n65346 = \P1_P3_Address_reg[4]/NET0131  & ~n9091 ;
  assign n65347 = \P1_P3_rEIP_reg[1]/NET0131  & n64081 ;
  assign n65348 = \P1_P3_rEIP_reg[2]/NET0131  & n65347 ;
  assign n65349 = \P1_P3_rEIP_reg[3]/NET0131  & n65348 ;
  assign n65350 = \P1_P3_rEIP_reg[4]/NET0131  & n65349 ;
  assign n65352 = \P1_P3_rEIP_reg[5]/NET0131  & n65350 ;
  assign n65351 = ~\P1_P3_rEIP_reg[5]/NET0131  & ~n65350 ;
  assign n65353 = n22115 & ~n65351 ;
  assign n65354 = ~n65352 & n65353 ;
  assign n65358 = ~n65346 & ~n65354 ;
  assign n65359 = ~n65357 & n65358 ;
  assign n65361 = ~\P1_P1_rEIP_reg[6]/NET0131  & ~n63385 ;
  assign n65362 = n26155 & ~n63386 ;
  assign n65363 = ~n65361 & n65362 ;
  assign n65360 = \P1_P1_Address_reg[4]/NET0131  & ~n26154 ;
  assign n65364 = \P1_P1_rEIP_reg[1]/NET0131  & n63402 ;
  assign n65365 = \P1_P1_rEIP_reg[2]/NET0131  & n65364 ;
  assign n65366 = \P1_P1_rEIP_reg[3]/NET0131  & n65365 ;
  assign n65367 = \P1_P1_rEIP_reg[4]/NET0131  & n65366 ;
  assign n65369 = ~\P1_P1_rEIP_reg[5]/NET0131  & ~n65367 ;
  assign n65368 = \P1_P1_rEIP_reg[5]/NET0131  & n65367 ;
  assign n65370 = n63401 & ~n65368 ;
  assign n65371 = ~n65369 & n65370 ;
  assign n65372 = ~n65360 & ~n65371 ;
  assign n65373 = ~n65363 & n65372 ;
  assign n65375 = ~\P2_P3_rEIP_reg[6]/NET0131  & ~n64106 ;
  assign n65376 = n27145 & ~n64107 ;
  assign n65377 = ~n65375 & n65376 ;
  assign n65374 = \P2_P3_Address_reg[4]/NET0131  & ~n27144 ;
  assign n65378 = \P2_P3_rEIP_reg[1]/NET0131  & n64095 ;
  assign n65379 = \P2_P3_rEIP_reg[2]/NET0131  & n65378 ;
  assign n65380 = \P2_P3_rEIP_reg[3]/NET0131  & n65379 ;
  assign n65381 = \P2_P3_rEIP_reg[4]/NET0131  & n65380 ;
  assign n65383 = ~\P2_P3_rEIP_reg[5]/NET0131  & ~n65381 ;
  assign n65382 = \P2_P3_rEIP_reg[5]/NET0131  & n65381 ;
  assign n65384 = n64094 & ~n65382 ;
  assign n65385 = ~n65383 & n65384 ;
  assign n65386 = ~n65374 & ~n65385 ;
  assign n65387 = ~n65377 & n65386 ;
  assign n65389 = ~\P1_P2_rEIP_reg[6]/NET0131  & ~n63432 ;
  assign n65390 = n25765 & ~n63433 ;
  assign n65391 = ~n65389 & n65390 ;
  assign n65388 = \P1_P2_Address_reg[4]/NET0131  & ~n25764 ;
  assign n65392 = \P1_P2_rEIP_reg[1]/NET0131  & n63421 ;
  assign n65393 = \P1_P2_rEIP_reg[2]/NET0131  & n65392 ;
  assign n65394 = \P1_P2_rEIP_reg[3]/NET0131  & n65393 ;
  assign n65395 = \P1_P2_rEIP_reg[4]/NET0131  & n65394 ;
  assign n65396 = ~\P1_P2_rEIP_reg[5]/NET0131  & ~n65395 ;
  assign n65397 = n48383 & n63421 ;
  assign n65398 = n63420 & ~n65397 ;
  assign n65399 = ~n65396 & n65398 ;
  assign n65400 = ~n65388 & ~n65399 ;
  assign n65401 = ~n65391 & n65400 ;
  assign n65403 = ~\P2_P1_rEIP_reg[6]/NET0131  & ~n63456 ;
  assign n65404 = n25955 & ~n63457 ;
  assign n65405 = ~n65403 & n65404 ;
  assign n65402 = \P2_P1_Address_reg[4]/NET0131  & ~n25954 ;
  assign n65406 = \P2_P1_rEIP_reg[1]/NET0131  & n63475 ;
  assign n65407 = \P2_P1_rEIP_reg[2]/NET0131  & n65406 ;
  assign n65408 = \P2_P1_rEIP_reg[3]/NET0131  & n65407 ;
  assign n65409 = \P2_P1_rEIP_reg[4]/NET0131  & n65408 ;
  assign n65411 = ~\P2_P1_rEIP_reg[5]/NET0131  & ~n65409 ;
  assign n65410 = \P2_P1_rEIP_reg[5]/NET0131  & n65409 ;
  assign n65412 = n63480 & ~n65410 ;
  assign n65413 = ~n65411 & n65412 ;
  assign n65414 = ~n65402 & ~n65413 ;
  assign n65415 = ~n65405 & n65414 ;
  assign n65417 = ~\P1_P3_rEIP_reg[17]/NET0131  & ~n64075 ;
  assign n65418 = n9092 & ~n64076 ;
  assign n65419 = ~n65417 & n65418 ;
  assign n65416 = \P1_P3_Address_reg[15]/NET0131  & ~n9091 ;
  assign n65420 = ~\P1_P3_rEIP_reg[16]/NET0131  & ~n64085 ;
  assign n65421 = n22115 & ~n64086 ;
  assign n65422 = ~n65420 & n65421 ;
  assign n65423 = ~n65416 & ~n65422 ;
  assign n65424 = ~n65419 & n65423 ;
  assign n65426 = ~\P2_P3_rEIP_reg[17]/NET0131  & ~n64117 ;
  assign n65427 = n27145 & ~n64118 ;
  assign n65428 = ~n65426 & n65427 ;
  assign n65425 = \P2_P3_Address_reg[15]/NET0131  & ~n27144 ;
  assign n65429 = n52560 & n64095 ;
  assign n65430 = ~\P2_P3_rEIP_reg[16]/NET0131  & ~n65429 ;
  assign n65431 = n64094 & ~n64097 ;
  assign n65432 = ~n65430 & n65431 ;
  assign n65433 = ~n65425 & ~n65432 ;
  assign n65434 = ~n65428 & n65433 ;
  assign n65436 = ~\P2_P2_rEIP_reg[16]/NET0131  & ~n63992 ;
  assign n65437 = n63373 & ~n63993 ;
  assign n65438 = ~n65436 & n65437 ;
  assign n65435 = \P2_P2_Address_reg[15]/NET0131  & ~n26646 ;
  assign n65439 = \P2_P2_rEIP_reg[15]/NET0131  & n63998 ;
  assign n65440 = \P2_P2_rEIP_reg[16]/NET0131  & n65439 ;
  assign n65441 = ~\P2_P2_rEIP_reg[17]/NET0131  & ~n65440 ;
  assign n65442 = n26647 & ~n63999 ;
  assign n65443 = ~n65441 & n65442 ;
  assign n65444 = ~n65435 & ~n65443 ;
  assign n65445 = ~n65438 & n65444 ;
  assign n65447 = ~\P2_P2_rEIP_reg[29]/NET0131  & ~n63362 ;
  assign n65448 = n26647 & ~n63363 ;
  assign n65449 = ~n65447 & n65448 ;
  assign n65446 = \P2_P2_Address_reg[27]/NET0131  & ~n26646 ;
  assign n65450 = ~\P2_P2_rEIP_reg[28]/NET0131  & ~n63370 ;
  assign n65451 = ~n63371 & n63373 ;
  assign n65452 = ~n65450 & n65451 ;
  assign n65453 = ~n65446 & ~n65452 ;
  assign n65454 = ~n65449 & n65453 ;
  assign n65456 = ~\P1_P1_rEIP_reg[17]/NET0131  & ~n64008 ;
  assign n65457 = n26155 & ~n64009 ;
  assign n65458 = ~n65456 & n65457 ;
  assign n65455 = \P1_P1_Address_reg[15]/NET0131  & ~n26154 ;
  assign n65459 = \P1_P1_rEIP_reg[15]/NET0131  & n63406 ;
  assign n65460 = ~\P1_P1_rEIP_reg[16]/NET0131  & ~n65459 ;
  assign n65461 = n63401 & ~n64014 ;
  assign n65462 = ~n65460 & n65461 ;
  assign n65463 = ~n65455 & ~n65462 ;
  assign n65464 = ~n65458 & n65463 ;
  assign n65467 = ~n51988 & n63402 ;
  assign n65466 = ~\P1_P1_rEIP_reg[28]/NET0131  & ~n63402 ;
  assign n65468 = n63401 & ~n65466 ;
  assign n65469 = ~n65467 & n65468 ;
  assign n65465 = \P1_P1_Address_reg[27]/NET0131  & ~n26154 ;
  assign n65470 = n52020 & n63395 ;
  assign n65471 = ~\P1_P1_rEIP_reg[29]/NET0131  & ~n65470 ;
  assign n65472 = n26155 & ~n63396 ;
  assign n65473 = ~n65471 & n65472 ;
  assign n65474 = ~n65465 & ~n65473 ;
  assign n65475 = ~n65469 & n65474 ;
  assign n65480 = \P1_P2_rEIP_reg[16]/NET0131  & n64033 ;
  assign n65481 = ~\P1_P2_rEIP_reg[17]/NET0131  & ~n65480 ;
  assign n65482 = n25765 & ~n64034 ;
  assign n65483 = ~n65481 & n65482 ;
  assign n65476 = \P1_P2_Address_reg[15]/NET0131  & ~n25764 ;
  assign n65477 = ~\P1_P2_rEIP_reg[16]/NET0131  & ~n64025 ;
  assign n65478 = n63420 & ~n64026 ;
  assign n65479 = ~n65477 & n65478 ;
  assign n65484 = ~n65476 & ~n65479 ;
  assign n65485 = ~n65483 & n65484 ;
  assign n65492 = \P1_P2_rEIP_reg[28]/NET0131  & n63442 ;
  assign n65493 = ~\P1_P2_rEIP_reg[29]/NET0131  & ~n65492 ;
  assign n65494 = n25765 & ~n63443 ;
  assign n65495 = ~n65493 & n65494 ;
  assign n65486 = \P1_P2_Address_reg[27]/NET0131  & ~n25764 ;
  assign n65489 = n51521 & n63421 ;
  assign n65487 = n51519 & n63421 ;
  assign n65488 = ~\P1_P2_rEIP_reg[28]/NET0131  & ~n65487 ;
  assign n65490 = n63420 & ~n65488 ;
  assign n65491 = ~n65489 & n65490 ;
  assign n65496 = ~n65486 & ~n65491 ;
  assign n65497 = ~n65495 & n65496 ;
  assign n65499 = \P2_P1_rEIP_reg[15]/NET0131  & n63462 ;
  assign n65500 = \P2_P1_rEIP_reg[16]/NET0131  & n65499 ;
  assign n65501 = ~\P2_P1_rEIP_reg[17]/NET0131  & ~n65500 ;
  assign n65502 = n25955 & ~n63463 ;
  assign n65503 = ~n65501 & n65502 ;
  assign n65498 = \P2_P1_Address_reg[15]/NET0131  & ~n25954 ;
  assign n65504 = \P2_P1_rEIP_reg[15]/NET0131  & n64050 ;
  assign n65505 = ~\P2_P1_rEIP_reg[16]/NET0131  & ~n65504 ;
  assign n65506 = n63480 & ~n64051 ;
  assign n65507 = ~n65505 & n65506 ;
  assign n65508 = ~n65498 & ~n65507 ;
  assign n65509 = ~n65503 & n65508 ;
  assign n65514 = \P2_P1_rEIP_reg[27]/NET0131  & n63477 ;
  assign n65515 = ~\P2_P1_rEIP_reg[28]/NET0131  & ~n65514 ;
  assign n65516 = ~n63478 & n63480 ;
  assign n65517 = ~n65515 & n65516 ;
  assign n65510 = \P2_P1_Address_reg[27]/NET0131  & ~n25954 ;
  assign n65511 = ~\P2_P1_rEIP_reg[29]/NET0131  & ~n63469 ;
  assign n65512 = n25955 & ~n63470 ;
  assign n65513 = ~n65511 & n65512 ;
  assign n65518 = ~n65510 & ~n65513 ;
  assign n65519 = ~n65517 & n65518 ;
  assign n65520 = \P3_rd_reg/NET0131  & \P4_IR_reg[27]/NET0131  ;
  assign n65521 = \P2_P3_Datao_reg[27]/NET0131  & ~\P3_rd_reg/NET0131  ;
  assign n65522 = ~n65520 & ~n65521 ;
  assign n65528 = n52234 & n63368 ;
  assign n65529 = ~\P2_P2_rEIP_reg[24]/NET0131  & ~n65528 ;
  assign n65530 = n63373 & ~n64765 ;
  assign n65531 = ~n65529 & n65530 ;
  assign n65523 = \P2_P2_Address_reg[23]/NET0131  & ~n26646 ;
  assign n65524 = n52306 & n63358 ;
  assign n65525 = ~\P2_P2_rEIP_reg[25]/NET0131  & ~n65524 ;
  assign n65526 = n26647 & ~n63359 ;
  assign n65527 = ~n65525 & n65526 ;
  assign n65532 = ~n65523 & ~n65527 ;
  assign n65533 = ~n65531 & n65532 ;
  assign n65538 = ~\P1_P1_rEIP_reg[25]/NET0131  & ~n64776 ;
  assign n65539 = n26155 & ~n64777 ;
  assign n65540 = ~n65538 & n65539 ;
  assign n65534 = \P1_P1_Address_reg[23]/NET0131  & ~n26154 ;
  assign n65535 = ~\P1_P1_rEIP_reg[24]/NET0131  & ~n63407 ;
  assign n65536 = n63401 & ~n63411 ;
  assign n65537 = ~n65535 & n65536 ;
  assign n65541 = ~n65534 & ~n65537 ;
  assign n65542 = ~n65540 & n65541 ;
  assign n65550 = ~n51408 & n63435 ;
  assign n65549 = ~\P1_P2_rEIP_reg[25]/NET0131  & ~n63435 ;
  assign n65551 = n25765 & ~n65549 ;
  assign n65552 = ~n65550 & n65551 ;
  assign n65543 = \P1_P2_Address_reg[23]/NET0131  & ~n25764 ;
  assign n65544 = n48385 & n63421 ;
  assign n65546 = n51352 & n65544 ;
  assign n65545 = ~\P1_P2_rEIP_reg[24]/NET0131  & ~n65544 ;
  assign n65547 = n63420 & ~n65545 ;
  assign n65548 = ~n65546 & n65547 ;
  assign n65553 = ~n65543 & ~n65548 ;
  assign n65554 = ~n65552 & n65553 ;
  assign n65557 = ~n50931 & n63475 ;
  assign n65556 = ~\P2_P1_rEIP_reg[24]/NET0131  & ~n63475 ;
  assign n65558 = n63480 & ~n65556 ;
  assign n65559 = ~n65557 & n65558 ;
  assign n65555 = \P2_P1_Address_reg[23]/NET0131  & ~n25954 ;
  assign n65560 = n50972 & n63459 ;
  assign n65561 = ~\P2_P1_rEIP_reg[25]/NET0131  & ~n65560 ;
  assign n65562 = n25955 & ~n65561 ;
  assign n65563 = ~n63466 & n65562 ;
  assign n65564 = ~n65555 & ~n65563 ;
  assign n65565 = ~n65559 & n65564 ;
  assign n65567 = \P2_P1_rEIP_reg[12]/NET0131  & n63461 ;
  assign n65568 = ~\P2_P1_rEIP_reg[13]/NET0131  & ~n65567 ;
  assign n65569 = n25955 & ~n64798 ;
  assign n65570 = ~n65568 & n65569 ;
  assign n65566 = \P2_P1_Address_reg[11]/NET0131  & ~n25954 ;
  assign n65571 = ~\P2_P1_rEIP_reg[12]/NET0131  & ~n64049 ;
  assign n65572 = n63480 & ~n64802 ;
  assign n65573 = ~n65571 & n65572 ;
  assign n65574 = ~n65566 & ~n65573 ;
  assign n65575 = ~n65570 & n65574 ;
  assign n65577 = \P1_P1_rEIP_reg[12]/NET0131  & n63391 ;
  assign n65578 = ~\P1_P1_rEIP_reg[13]/NET0131  & ~n65577 ;
  assign n65579 = n26155 & ~n63392 ;
  assign n65580 = ~n65578 & n65579 ;
  assign n65576 = \P1_P1_Address_reg[11]/NET0131  & ~n26154 ;
  assign n65581 = ~\P1_P1_rEIP_reg[12]/NET0131  & ~n63404 ;
  assign n65582 = n63401 & ~n64810 ;
  assign n65583 = ~n65581 & n65582 ;
  assign n65584 = ~n65576 & ~n65583 ;
  assign n65585 = ~n65580 & n65584 ;
  assign n65587 = \P2_P2_rEIP_reg[12]/NET0131  & n64821 ;
  assign n65588 = ~\P2_P2_rEIP_reg[13]/NET0131  & ~n65587 ;
  assign n65589 = n26647 & ~n64822 ;
  assign n65590 = ~n65588 & n65589 ;
  assign n65586 = \P2_P2_Address_reg[11]/NET0131  & ~n26646 ;
  assign n65591 = ~\P2_P2_rEIP_reg[12]/NET0131  & ~n63989 ;
  assign n65592 = n63373 & ~n64826 ;
  assign n65593 = ~n65591 & n65592 ;
  assign n65594 = ~n65586 & ~n65593 ;
  assign n65595 = ~n65590 & n65594 ;
  assign n65597 = ~\P1_P3_rEIP_reg[13]/NET0131  & ~n64071 ;
  assign n65598 = n9092 & ~n64072 ;
  assign n65599 = ~n65597 & n65598 ;
  assign n65596 = \P1_P3_Address_reg[11]/NET0131  & ~n9091 ;
  assign n65600 = n16577 & n64081 ;
  assign n65601 = ~\P1_P3_rEIP_reg[12]/NET0131  & ~n65600 ;
  assign n65602 = n22115 & ~n64082 ;
  assign n65603 = ~n65601 & n65602 ;
  assign n65604 = ~n65596 & ~n65603 ;
  assign n65605 = ~n65599 & n65604 ;
  assign n65607 = \P1_P2_rEIP_reg[12]/NET0131  & n64032 ;
  assign n65608 = ~\P1_P2_rEIP_reg[13]/NET0131  & ~n65607 ;
  assign n65609 = n25765 & ~n64842 ;
  assign n65610 = ~n65608 & n65609 ;
  assign n65606 = \P1_P2_Address_reg[11]/NET0131  & ~n25764 ;
  assign n65611 = ~\P1_P2_rEIP_reg[12]/NET0131  & ~n64848 ;
  assign n65612 = n63420 & ~n64849 ;
  assign n65613 = ~n65611 & n65612 ;
  assign n65614 = ~n65606 & ~n65613 ;
  assign n65615 = ~n65610 & n65614 ;
  assign n65621 = ~\P2_P3_rEIP_reg[13]/NET0131  & ~n64113 ;
  assign n65622 = n27145 & ~n64114 ;
  assign n65623 = ~n65621 & n65622 ;
  assign n65616 = \P2_P3_Address_reg[11]/NET0131  & ~n27144 ;
  assign n65618 = ~n56156 & n64095 ;
  assign n65617 = ~\P2_P3_rEIP_reg[12]/NET0131  & ~n64095 ;
  assign n65619 = n64094 & ~n65617 ;
  assign n65620 = ~n65618 & n65619 ;
  assign n65624 = ~n65616 & ~n65620 ;
  assign n65625 = ~n65623 & n65624 ;
  assign n65626 = \P3_rd_reg/NET0131  & \P4_IR_reg[24]/NET0131  ;
  assign n65627 = \P2_P3_Datao_reg[24]/NET0131  & ~\P3_rd_reg/NET0131  ;
  assign n65628 = ~n65626 & ~n65627 ;
  assign n65630 = ~\P2_P2_rEIP_reg[5]/NET0131  & ~n63354 ;
  assign n65631 = n26647 & ~n63355 ;
  assign n65632 = ~n65630 & n65631 ;
  assign n65629 = \P2_P2_Address_reg[3]/NET0131  & ~n26646 ;
  assign n65633 = ~\P2_P2_rEIP_reg[4]/NET0131  & ~n65338 ;
  assign n65634 = n63373 & ~n65339 ;
  assign n65635 = ~n65633 & n65634 ;
  assign n65636 = ~n65629 & ~n65635 ;
  assign n65637 = ~n65632 & n65636 ;
  assign n65639 = ~\P1_P3_rEIP_reg[5]/NET0131  & ~n64063 ;
  assign n65640 = n9092 & ~n64064 ;
  assign n65641 = ~n65639 & n65640 ;
  assign n65638 = \P1_P3_Address_reg[3]/NET0131  & ~n9091 ;
  assign n65642 = ~\P1_P3_rEIP_reg[4]/NET0131  & ~n65349 ;
  assign n65643 = n22115 & ~n65350 ;
  assign n65644 = ~n65642 & n65643 ;
  assign n65645 = ~n65638 & ~n65644 ;
  assign n65646 = ~n65641 & n65645 ;
  assign n65648 = ~\P1_P1_rEIP_reg[5]/NET0131  & ~n63384 ;
  assign n65649 = n26155 & ~n63385 ;
  assign n65650 = ~n65648 & n65649 ;
  assign n65647 = \P1_P1_Address_reg[3]/NET0131  & ~n26154 ;
  assign n65651 = ~\P1_P1_rEIP_reg[4]/NET0131  & ~n65366 ;
  assign n65652 = n63401 & ~n65367 ;
  assign n65653 = ~n65651 & n65652 ;
  assign n65654 = ~n65647 & ~n65653 ;
  assign n65655 = ~n65650 & n65654 ;
  assign n65657 = ~\P1_P2_rEIP_reg[5]/NET0131  & ~n63431 ;
  assign n65658 = n25765 & ~n63432 ;
  assign n65659 = ~n65657 & n65658 ;
  assign n65656 = \P1_P2_Address_reg[3]/NET0131  & ~n25764 ;
  assign n65660 = ~\P1_P2_rEIP_reg[4]/NET0131  & ~n65394 ;
  assign n65661 = n63420 & ~n65395 ;
  assign n65662 = ~n65660 & n65661 ;
  assign n65663 = ~n65656 & ~n65662 ;
  assign n65664 = ~n65659 & n65663 ;
  assign n65666 = ~\P2_P3_rEIP_reg[5]/NET0131  & ~n64105 ;
  assign n65667 = n27145 & ~n64106 ;
  assign n65668 = ~n65666 & n65667 ;
  assign n65665 = \P2_P3_Address_reg[3]/NET0131  & ~n27144 ;
  assign n65669 = ~\P2_P3_rEIP_reg[4]/NET0131  & ~n65380 ;
  assign n65670 = n64094 & ~n65381 ;
  assign n65671 = ~n65669 & n65670 ;
  assign n65672 = ~n65665 & ~n65671 ;
  assign n65673 = ~n65668 & n65672 ;
  assign n65675 = ~\P2_P1_rEIP_reg[5]/NET0131  & ~n63455 ;
  assign n65676 = n25955 & ~n63456 ;
  assign n65677 = ~n65675 & n65676 ;
  assign n65674 = \P2_P1_Address_reg[3]/NET0131  & ~n25954 ;
  assign n65678 = ~\P2_P1_rEIP_reg[4]/NET0131  & ~n65408 ;
  assign n65679 = n63480 & ~n65409 ;
  assign n65680 = ~n65678 & n65679 ;
  assign n65681 = ~n65674 & ~n65680 ;
  assign n65682 = ~n65677 & n65681 ;
  assign n65684 = ~\P2_P2_rEIP_reg[20]/NET0131  & ~n65225 ;
  assign n65685 = n63373 & ~n65226 ;
  assign n65686 = ~n65684 & n65685 ;
  assign n65683 = \P2_P2_Address_reg[19]/NET0131  & ~n26646 ;
  assign n65687 = n52103 & n63998 ;
  assign n65688 = \P2_P2_rEIP_reg[20]/NET0131  & n65687 ;
  assign n65689 = ~\P2_P2_rEIP_reg[21]/NET0131  & ~n65688 ;
  assign n65690 = n26647 & ~n65231 ;
  assign n65691 = ~n65689 & n65690 ;
  assign n65692 = ~n65683 & ~n65691 ;
  assign n65693 = ~n65686 & n65692 ;
  assign n65699 = n51666 & n64008 ;
  assign n65700 = \P1_P1_rEIP_reg[20]/NET0131  & n65699 ;
  assign n65701 = ~\P1_P1_rEIP_reg[21]/NET0131  & ~n65700 ;
  assign n65702 = n26155 & ~n65239 ;
  assign n65703 = ~n65701 & n65702 ;
  assign n65694 = \P1_P1_Address_reg[19]/NET0131  & ~n26154 ;
  assign n65695 = n51666 & n64014 ;
  assign n65696 = ~\P1_P1_rEIP_reg[20]/NET0131  & ~n65695 ;
  assign n65697 = n63401 & ~n65244 ;
  assign n65698 = ~n65696 & n65697 ;
  assign n65704 = ~n65694 & ~n65698 ;
  assign n65705 = ~n65703 & n65704 ;
  assign n65707 = n51203 & n63421 ;
  assign n65708 = \P1_P2_rEIP_reg[20]/NET0131  & ~n65707 ;
  assign n65709 = \P1_P2_rEIP_reg[19]/NET0131  & ~\P1_P2_rEIP_reg[20]/NET0131  ;
  assign n65710 = n65252 & n65709 ;
  assign n65711 = ~n65708 & ~n65710 ;
  assign n65712 = n63420 & ~n65711 ;
  assign n65706 = \P1_P2_Address_reg[19]/NET0131  & ~n25764 ;
  assign n65713 = ~\P1_P2_rEIP_reg[21]/NET0131  & ~n63437 ;
  assign n65714 = n25765 & ~n63438 ;
  assign n65715 = ~n65713 & n65714 ;
  assign n65716 = ~n65706 & ~n65715 ;
  assign n65717 = ~n65712 & n65716 ;
  assign n65724 = ~\P2_P1_rEIP_reg[21]/NET0131  & ~n63464 ;
  assign n65725 = n25955 & ~n65217 ;
  assign n65726 = ~n65724 & n65725 ;
  assign n65718 = \P2_P1_Address_reg[19]/NET0131  & ~n25954 ;
  assign n65719 = n50780 & n64053 ;
  assign n65721 = \P2_P1_rEIP_reg[20]/NET0131  & n65719 ;
  assign n65720 = ~\P2_P1_rEIP_reg[20]/NET0131  & ~n65719 ;
  assign n65722 = n63480 & ~n65720 ;
  assign n65723 = ~n65721 & n65722 ;
  assign n65727 = ~n65718 & ~n65723 ;
  assign n65728 = ~n65726 & n65727 ;
  assign n65730 = ~\P2_P1_rEIP_reg[9]/NET0131  & ~n63459 ;
  assign n65731 = n25955 & ~n63460 ;
  assign n65732 = ~n65730 & n65731 ;
  assign n65729 = \P2_P1_Address_reg[7]/NET0131  & ~n25954 ;
  assign n65733 = ~\P2_P1_rEIP_reg[8]/NET0131  & ~n64046 ;
  assign n65734 = n63480 & ~n64047 ;
  assign n65735 = ~n65733 & n65734 ;
  assign n65736 = ~n65729 & ~n65735 ;
  assign n65737 = ~n65732 & n65736 ;
  assign n65739 = ~\P2_P2_rEIP_reg[9]/NET0131  & ~n63358 ;
  assign n65740 = n26647 & ~n64820 ;
  assign n65741 = ~n65739 & n65740 ;
  assign n65738 = \P2_P2_Address_reg[7]/NET0131  & ~n26646 ;
  assign n65742 = ~\P2_P2_rEIP_reg[8]/NET0131  & ~n63986 ;
  assign n65743 = n63373 & ~n63987 ;
  assign n65744 = ~n65742 & n65743 ;
  assign n65745 = ~n65738 & ~n65744 ;
  assign n65746 = ~n65741 & n65745 ;
  assign n65752 = ~\P1_P3_rEIP_reg[9]/NET0131  & ~n64067 ;
  assign n65753 = n9092 & ~n64068 ;
  assign n65754 = ~n65752 & n65753 ;
  assign n65747 = \P1_P3_Address_reg[7]/NET0131  & ~n9091 ;
  assign n65749 = ~n17948 & n64081 ;
  assign n65748 = ~\P1_P3_rEIP_reg[8]/NET0131  & ~n64081 ;
  assign n65750 = n22115 & ~n65748 ;
  assign n65751 = ~n65749 & n65750 ;
  assign n65755 = ~n65747 & ~n65751 ;
  assign n65756 = ~n65754 & n65755 ;
  assign n65758 = ~\P1_P1_rEIP_reg[9]/NET0131  & ~n63388 ;
  assign n65759 = n26155 & ~n63389 ;
  assign n65760 = ~n65758 & n65759 ;
  assign n65757 = \P1_P1_Address_reg[7]/NET0131  & ~n26154 ;
  assign n65761 = ~\P1_P1_rEIP_reg[8]/NET0131  & ~n65288 ;
  assign n65762 = n63401 & ~n65289 ;
  assign n65763 = ~n65761 & n65762 ;
  assign n65764 = ~n65757 & ~n65763 ;
  assign n65765 = ~n65760 & n65764 ;
  assign n65767 = ~\P2_P3_rEIP_reg[9]/NET0131  & ~n64109 ;
  assign n65768 = n27145 & ~n64110 ;
  assign n65769 = ~n65767 & n65768 ;
  assign n65766 = \P2_P3_Address_reg[7]/NET0131  & ~n27144 ;
  assign n65770 = ~\P2_P3_rEIP_reg[8]/NET0131  & ~n65301 ;
  assign n65771 = n64094 & ~n65302 ;
  assign n65772 = ~n65770 & n65771 ;
  assign n65773 = ~n65766 & ~n65772 ;
  assign n65774 = ~n65769 & n65773 ;
  assign n65776 = ~\P1_P2_rEIP_reg[9]/NET0131  & ~n63435 ;
  assign n65777 = n25765 & ~n64031 ;
  assign n65778 = ~n65776 & n65777 ;
  assign n65775 = \P1_P2_Address_reg[7]/NET0131  & ~n25764 ;
  assign n65779 = ~\P1_P2_rEIP_reg[8]/NET0131  & ~n65544 ;
  assign n65780 = n63420 & ~n64787 ;
  assign n65781 = ~n65779 & n65780 ;
  assign n65782 = ~n65775 & ~n65781 ;
  assign n65783 = ~n65778 & n65782 ;
  assign n65786 = ~\P1_P1_BE_n_reg[3]/NET0131  & ~\P1_P1_D_C_n_reg/NET0131  ;
  assign n65787 = \P1_P1_M_IO_n_reg/NET0131  & \P1_P1_W_R_n_reg/NET0131  ;
  assign n65788 = n65786 & n65787 ;
  assign n65784 = ~\P1_P1_ADS_n_reg/NET0131  & ~\P1_P1_BE_n_reg[0]/NET0131  ;
  assign n65785 = ~\P1_P1_BE_n_reg[1]/NET0131  & ~\P1_P1_BE_n_reg[2]/NET0131  ;
  assign n65789 = n65784 & n65785 ;
  assign n65790 = n65788 & n65789 ;
  assign n65791 = n7653 & n65790 ;
  assign n65794 = ~\P1_P2_BE_n_reg[3]/NET0131  & ~\P1_P2_D_C_n_reg/NET0131  ;
  assign n65795 = \P1_P2_M_IO_n_reg/NET0131  & \P1_P2_W_R_n_reg/NET0131  ;
  assign n65796 = n65794 & n65795 ;
  assign n65792 = ~\P1_P2_ADS_n_reg/NET0131  & ~\P1_P2_BE_n_reg[0]/NET0131  ;
  assign n65793 = ~\P1_P2_BE_n_reg[1]/NET0131  & ~\P1_P2_BE_n_reg[2]/NET0131  ;
  assign n65797 = n65792 & n65793 ;
  assign n65798 = n65796 & n65797 ;
  assign n65799 = n27934 & n65798 ;
  assign n65800 = \P1_buf1_reg[17]/NET0131  & ~n65799 ;
  assign n65801 = \P1_P2_Datao_reg[17]/NET0131  & n65799 ;
  assign n65802 = ~n65800 & ~n65801 ;
  assign n65803 = ~n65791 & ~n65802 ;
  assign n65804 = \P1_P1_Datao_reg[17]/NET0131  & n65791 ;
  assign n65805 = ~n65803 & ~n65804 ;
  assign n65808 = ~\P2_P1_BE_n_reg[3]/NET0131  & ~\P2_P1_D_C_n_reg/NET0131  ;
  assign n65809 = \P2_P1_M_IO_n_reg/NET0131  & \P2_P1_W_R_n_reg/NET0131  ;
  assign n65810 = n65808 & n65809 ;
  assign n65806 = ~\P2_P1_ADS_n_reg/NET0131  & ~\P2_P1_BE_n_reg[0]/NET0131  ;
  assign n65807 = ~\P2_P1_BE_n_reg[1]/NET0131  & ~\P2_P1_BE_n_reg[2]/NET0131  ;
  assign n65811 = n65806 & n65807 ;
  assign n65812 = n65810 & n65811 ;
  assign n65813 = n10134 & n65812 ;
  assign n65816 = ~\P2_P2_BE_n_reg[3]/NET0131  & ~\P2_P2_D_C_n_reg/NET0131  ;
  assign n65817 = \P2_P2_M_IO_n_reg/NET0131  & \P2_P2_W_R_n_reg/NET0131  ;
  assign n65818 = n65816 & n65817 ;
  assign n65814 = ~\P2_P2_ADS_n_reg/NET0131  & ~\P2_P2_BE_n_reg[0]/NET0131  ;
  assign n65815 = ~\P2_P2_BE_n_reg[1]/NET0131  & ~\P2_P2_BE_n_reg[2]/NET0131  ;
  assign n65819 = n65814 & n65815 ;
  assign n65820 = n65818 & n65819 ;
  assign n65821 = n28013 & n65820 ;
  assign n65822 = \P2_buf1_reg[12]/NET0131  & ~n65821 ;
  assign n65823 = \P2_P2_Datao_reg[12]/NET0131  & n65821 ;
  assign n65824 = ~n65822 & ~n65823 ;
  assign n65825 = ~n65813 & ~n65824 ;
  assign n65826 = \P2_P1_Datao_reg[12]/NET0131  & n65813 ;
  assign n65827 = ~n65825 & ~n65826 ;
  assign n65828 = \P2_buf1_reg[11]/NET0131  & ~n65821 ;
  assign n65829 = \P2_P2_Datao_reg[11]/NET0131  & n65821 ;
  assign n65830 = ~n65828 & ~n65829 ;
  assign n65831 = ~n65813 & ~n65830 ;
  assign n65832 = \P2_P1_Datao_reg[11]/NET0131  & n65813 ;
  assign n65833 = ~n65831 & ~n65832 ;
  assign n65834 = \P2_buf1_reg[14]/NET0131  & ~n65821 ;
  assign n65835 = \P2_P2_Datao_reg[14]/NET0131  & n65821 ;
  assign n65836 = ~n65834 & ~n65835 ;
  assign n65837 = ~n65813 & ~n65836 ;
  assign n65838 = \P2_P1_Datao_reg[14]/NET0131  & n65813 ;
  assign n65839 = ~n65837 & ~n65838 ;
  assign n65840 = \P1_buf1_reg[1]/NET0131  & ~n65799 ;
  assign n65841 = \P1_P2_Datao_reg[1]/NET0131  & n65799 ;
  assign n65842 = ~n65840 & ~n65841 ;
  assign n65843 = ~n65791 & ~n65842 ;
  assign n65844 = \P1_P1_Datao_reg[1]/NET0131  & n65791 ;
  assign n65845 = ~n65843 & ~n65844 ;
  assign n65846 = \P1_buf1_reg[11]/NET0131  & ~n65799 ;
  assign n65847 = \P1_P2_Datao_reg[11]/NET0131  & n65799 ;
  assign n65848 = ~n65846 & ~n65847 ;
  assign n65849 = ~n65791 & ~n65848 ;
  assign n65850 = \P1_P1_Datao_reg[11]/NET0131  & n65791 ;
  assign n65851 = ~n65849 & ~n65850 ;
  assign n65852 = \P2_buf1_reg[9]/NET0131  & ~n65821 ;
  assign n65853 = \P2_P2_Datao_reg[9]/NET0131  & n65821 ;
  assign n65854 = ~n65852 & ~n65853 ;
  assign n65855 = ~n65813 & ~n65854 ;
  assign n65856 = \P2_P1_Datao_reg[9]/NET0131  & n65813 ;
  assign n65857 = ~n65855 & ~n65856 ;
  assign n65858 = \P1_buf1_reg[10]/NET0131  & ~n65799 ;
  assign n65859 = \P1_P2_Datao_reg[10]/NET0131  & n65799 ;
  assign n65860 = ~n65858 & ~n65859 ;
  assign n65861 = ~n65791 & ~n65860 ;
  assign n65862 = \P1_P1_Datao_reg[10]/NET0131  & n65791 ;
  assign n65863 = ~n65861 & ~n65862 ;
  assign n65864 = \P1_buf1_reg[5]/NET0131  & ~n65799 ;
  assign n65865 = \P1_P2_Datao_reg[5]/NET0131  & n65799 ;
  assign n65866 = ~n65864 & ~n65865 ;
  assign n65867 = ~n65791 & ~n65866 ;
  assign n65868 = \P1_P1_Datao_reg[5]/NET0131  & n65791 ;
  assign n65869 = ~n65867 & ~n65868 ;
  assign n65870 = \P2_buf1_reg[5]/NET0131  & ~n65821 ;
  assign n65871 = \P2_P2_Datao_reg[5]/NET0131  & n65821 ;
  assign n65872 = ~n65870 & ~n65871 ;
  assign n65873 = ~n65813 & ~n65872 ;
  assign n65874 = \P2_P1_Datao_reg[5]/NET0131  & n65813 ;
  assign n65875 = ~n65873 & ~n65874 ;
  assign n65876 = \P1_buf1_reg[16]/NET0131  & ~n65799 ;
  assign n65877 = \P1_P2_Datao_reg[16]/NET0131  & n65799 ;
  assign n65878 = ~n65876 & ~n65877 ;
  assign n65879 = ~n65791 & ~n65878 ;
  assign n65880 = \P1_P1_Datao_reg[16]/NET0131  & n65791 ;
  assign n65881 = ~n65879 & ~n65880 ;
  assign n65882 = \P1_buf1_reg[23]/NET0131  & ~n65799 ;
  assign n65883 = \P1_P2_Datao_reg[23]/NET0131  & n65799 ;
  assign n65884 = ~n65882 & ~n65883 ;
  assign n65885 = ~n65791 & ~n65884 ;
  assign n65886 = \P1_P1_Datao_reg[23]/NET0131  & n65791 ;
  assign n65887 = ~n65885 & ~n65886 ;
  assign n65888 = \P2_buf1_reg[0]/NET0131  & ~n65821 ;
  assign n65889 = \P2_P2_Datao_reg[0]/NET0131  & n65821 ;
  assign n65890 = ~n65888 & ~n65889 ;
  assign n65891 = ~n65813 & ~n65890 ;
  assign n65892 = \P2_P1_Datao_reg[0]/NET0131  & n65813 ;
  assign n65893 = ~n65891 & ~n65892 ;
  assign n65894 = \P2_buf1_reg[10]/NET0131  & ~n65821 ;
  assign n65895 = \P2_P2_Datao_reg[10]/NET0131  & n65821 ;
  assign n65896 = ~n65894 & ~n65895 ;
  assign n65897 = ~n65813 & ~n65896 ;
  assign n65898 = \P2_P1_Datao_reg[10]/NET0131  & n65813 ;
  assign n65899 = ~n65897 & ~n65898 ;
  assign n65900 = \P2_buf1_reg[13]/NET0131  & ~n65821 ;
  assign n65901 = \P2_P2_Datao_reg[13]/NET0131  & n65821 ;
  assign n65902 = ~n65900 & ~n65901 ;
  assign n65903 = ~n65813 & ~n65902 ;
  assign n65904 = \P2_P1_Datao_reg[13]/NET0131  & n65813 ;
  assign n65905 = ~n65903 & ~n65904 ;
  assign n65906 = \P2_buf1_reg[15]/NET0131  & ~n65821 ;
  assign n65907 = \P2_P2_Datao_reg[15]/NET0131  & n65821 ;
  assign n65908 = ~n65906 & ~n65907 ;
  assign n65909 = ~n65813 & ~n65908 ;
  assign n65910 = \P2_P1_Datao_reg[15]/NET0131  & n65813 ;
  assign n65911 = ~n65909 & ~n65910 ;
  assign n65912 = \P2_buf1_reg[16]/NET0131  & ~n65821 ;
  assign n65913 = \P2_P2_Datao_reg[16]/NET0131  & n65821 ;
  assign n65914 = ~n65912 & ~n65913 ;
  assign n65915 = ~n65813 & ~n65914 ;
  assign n65916 = \P2_P1_Datao_reg[16]/NET0131  & n65813 ;
  assign n65917 = ~n65915 & ~n65916 ;
  assign n65918 = \P2_buf1_reg[17]/NET0131  & ~n65821 ;
  assign n65919 = \P2_P2_Datao_reg[17]/NET0131  & n65821 ;
  assign n65920 = ~n65918 & ~n65919 ;
  assign n65921 = ~n65813 & ~n65920 ;
  assign n65922 = \P2_P1_Datao_reg[17]/NET0131  & n65813 ;
  assign n65923 = ~n65921 & ~n65922 ;
  assign n65924 = \P2_buf1_reg[18]/NET0131  & ~n65821 ;
  assign n65925 = \P2_P2_Datao_reg[18]/NET0131  & n65821 ;
  assign n65926 = ~n65924 & ~n65925 ;
  assign n65927 = ~n65813 & ~n65926 ;
  assign n65928 = \P2_P1_Datao_reg[18]/NET0131  & n65813 ;
  assign n65929 = ~n65927 & ~n65928 ;
  assign n65930 = \P2_buf1_reg[19]/NET0131  & ~n65821 ;
  assign n65931 = \P2_P2_Datao_reg[19]/NET0131  & n65821 ;
  assign n65932 = ~n65930 & ~n65931 ;
  assign n65933 = ~n65813 & ~n65932 ;
  assign n65934 = \P2_P1_Datao_reg[19]/NET0131  & n65813 ;
  assign n65935 = ~n65933 & ~n65934 ;
  assign n65936 = \P2_buf1_reg[1]/NET0131  & ~n65821 ;
  assign n65937 = \P2_P2_Datao_reg[1]/NET0131  & n65821 ;
  assign n65938 = ~n65936 & ~n65937 ;
  assign n65939 = ~n65813 & ~n65938 ;
  assign n65940 = \P2_P1_Datao_reg[1]/NET0131  & n65813 ;
  assign n65941 = ~n65939 & ~n65940 ;
  assign n65942 = \P2_buf1_reg[20]/NET0131  & ~n65821 ;
  assign n65943 = \P2_P2_Datao_reg[20]/NET0131  & n65821 ;
  assign n65944 = ~n65942 & ~n65943 ;
  assign n65945 = ~n65813 & ~n65944 ;
  assign n65946 = \P2_P1_Datao_reg[20]/NET0131  & n65813 ;
  assign n65947 = ~n65945 & ~n65946 ;
  assign n65948 = \P2_buf1_reg[21]/NET0131  & ~n65821 ;
  assign n65949 = \P2_P2_Datao_reg[21]/NET0131  & n65821 ;
  assign n65950 = ~n65948 & ~n65949 ;
  assign n65951 = ~n65813 & ~n65950 ;
  assign n65952 = \P2_P1_Datao_reg[21]/NET0131  & n65813 ;
  assign n65953 = ~n65951 & ~n65952 ;
  assign n65954 = \P2_buf1_reg[22]/NET0131  & ~n65821 ;
  assign n65955 = \P2_P2_Datao_reg[22]/NET0131  & n65821 ;
  assign n65956 = ~n65954 & ~n65955 ;
  assign n65957 = ~n65813 & ~n65956 ;
  assign n65958 = \P2_P1_Datao_reg[22]/NET0131  & n65813 ;
  assign n65959 = ~n65957 & ~n65958 ;
  assign n65960 = \P2_buf1_reg[23]/NET0131  & ~n65821 ;
  assign n65961 = \P2_P2_Datao_reg[23]/NET0131  & n65821 ;
  assign n65962 = ~n65960 & ~n65961 ;
  assign n65963 = ~n65813 & ~n65962 ;
  assign n65964 = \P2_P1_Datao_reg[23]/NET0131  & n65813 ;
  assign n65965 = ~n65963 & ~n65964 ;
  assign n65966 = \P2_buf1_reg[24]/NET0131  & ~n65821 ;
  assign n65967 = \P2_P2_Datao_reg[24]/NET0131  & n65821 ;
  assign n65968 = ~n65966 & ~n65967 ;
  assign n65969 = ~n65813 & ~n65968 ;
  assign n65970 = \P2_P1_Datao_reg[24]/NET0131  & n65813 ;
  assign n65971 = ~n65969 & ~n65970 ;
  assign n65972 = \P2_buf1_reg[25]/NET0131  & ~n65821 ;
  assign n65973 = \P2_P2_Datao_reg[25]/NET0131  & n65821 ;
  assign n65974 = ~n65972 & ~n65973 ;
  assign n65975 = ~n65813 & ~n65974 ;
  assign n65976 = \P2_P1_Datao_reg[25]/NET0131  & n65813 ;
  assign n65977 = ~n65975 & ~n65976 ;
  assign n65978 = \P2_buf1_reg[26]/NET0131  & ~n65821 ;
  assign n65979 = \P2_P2_Datao_reg[26]/NET0131  & n65821 ;
  assign n65980 = ~n65978 & ~n65979 ;
  assign n65981 = ~n65813 & ~n65980 ;
  assign n65982 = \P2_P1_Datao_reg[26]/NET0131  & n65813 ;
  assign n65983 = ~n65981 & ~n65982 ;
  assign n65984 = \P2_buf1_reg[28]/NET0131  & ~n65821 ;
  assign n65985 = \P2_P2_Datao_reg[28]/NET0131  & n65821 ;
  assign n65986 = ~n65984 & ~n65985 ;
  assign n65987 = ~n65813 & ~n65986 ;
  assign n65988 = \P2_P1_Datao_reg[28]/NET0131  & n65813 ;
  assign n65989 = ~n65987 & ~n65988 ;
  assign n65990 = \P2_buf1_reg[29]/NET0131  & ~n65821 ;
  assign n65991 = \P2_P2_Datao_reg[29]/NET0131  & n65821 ;
  assign n65992 = ~n65990 & ~n65991 ;
  assign n65993 = ~n65813 & ~n65992 ;
  assign n65994 = \P2_P1_Datao_reg[29]/NET0131  & n65813 ;
  assign n65995 = ~n65993 & ~n65994 ;
  assign n65996 = \P2_buf1_reg[2]/NET0131  & ~n65821 ;
  assign n65997 = \P2_P2_Datao_reg[2]/NET0131  & n65821 ;
  assign n65998 = ~n65996 & ~n65997 ;
  assign n65999 = ~n65813 & ~n65998 ;
  assign n66000 = \P2_P1_Datao_reg[2]/NET0131  & n65813 ;
  assign n66001 = ~n65999 & ~n66000 ;
  assign n66002 = \P2_buf1_reg[30]/NET0131  & ~n65821 ;
  assign n66003 = \P2_P2_Datao_reg[30]/NET0131  & n65821 ;
  assign n66004 = ~n66002 & ~n66003 ;
  assign n66005 = ~n65813 & ~n66004 ;
  assign n66006 = \P2_P1_Datao_reg[30]/NET0131  & n65813 ;
  assign n66007 = ~n66005 & ~n66006 ;
  assign n66008 = \P2_buf1_reg[3]/NET0131  & ~n65821 ;
  assign n66009 = \P2_P2_Datao_reg[3]/NET0131  & n65821 ;
  assign n66010 = ~n66008 & ~n66009 ;
  assign n66011 = ~n65813 & ~n66010 ;
  assign n66012 = \P2_P1_Datao_reg[3]/NET0131  & n65813 ;
  assign n66013 = ~n66011 & ~n66012 ;
  assign n66014 = \P2_buf1_reg[4]/NET0131  & ~n65821 ;
  assign n66015 = \P2_P2_Datao_reg[4]/NET0131  & n65821 ;
  assign n66016 = ~n66014 & ~n66015 ;
  assign n66017 = ~n65813 & ~n66016 ;
  assign n66018 = \P2_P1_Datao_reg[4]/NET0131  & n65813 ;
  assign n66019 = ~n66017 & ~n66018 ;
  assign n66020 = \P2_buf1_reg[6]/NET0131  & ~n65821 ;
  assign n66021 = \P2_P2_Datao_reg[6]/NET0131  & n65821 ;
  assign n66022 = ~n66020 & ~n66021 ;
  assign n66023 = ~n65813 & ~n66022 ;
  assign n66024 = \P2_P1_Datao_reg[6]/NET0131  & n65813 ;
  assign n66025 = ~n66023 & ~n66024 ;
  assign n66026 = \P2_buf1_reg[7]/NET0131  & ~n65821 ;
  assign n66027 = \P2_P2_Datao_reg[7]/NET0131  & n65821 ;
  assign n66028 = ~n66026 & ~n66027 ;
  assign n66029 = ~n65813 & ~n66028 ;
  assign n66030 = \P2_P1_Datao_reg[7]/NET0131  & n65813 ;
  assign n66031 = ~n66029 & ~n66030 ;
  assign n66032 = \P2_buf1_reg[8]/NET0131  & ~n65821 ;
  assign n66033 = \P2_P2_Datao_reg[8]/NET0131  & n65821 ;
  assign n66034 = ~n66032 & ~n66033 ;
  assign n66035 = ~n65813 & ~n66034 ;
  assign n66036 = \P2_P1_Datao_reg[8]/NET0131  & n65813 ;
  assign n66037 = ~n66035 & ~n66036 ;
  assign n66038 = \P2_buf1_reg[27]/NET0131  & ~n65821 ;
  assign n66039 = \P2_P2_Datao_reg[27]/NET0131  & n65821 ;
  assign n66040 = ~n66038 & ~n66039 ;
  assign n66041 = ~n65813 & ~n66040 ;
  assign n66042 = \P2_P1_Datao_reg[27]/NET0131  & n65813 ;
  assign n66043 = ~n66041 & ~n66042 ;
  assign n66044 = \P1_buf1_reg[12]/NET0131  & ~n65799 ;
  assign n66045 = \P1_P2_Datao_reg[12]/NET0131  & n65799 ;
  assign n66046 = ~n66044 & ~n66045 ;
  assign n66047 = ~n65791 & ~n66046 ;
  assign n66048 = \P1_P1_Datao_reg[12]/NET0131  & n65791 ;
  assign n66049 = ~n66047 & ~n66048 ;
  assign n66050 = \P1_buf1_reg[13]/NET0131  & ~n65799 ;
  assign n66051 = \P1_P2_Datao_reg[13]/NET0131  & n65799 ;
  assign n66052 = ~n66050 & ~n66051 ;
  assign n66053 = ~n65791 & ~n66052 ;
  assign n66054 = \P1_P1_Datao_reg[13]/NET0131  & n65791 ;
  assign n66055 = ~n66053 & ~n66054 ;
  assign n66056 = \P1_buf1_reg[14]/NET0131  & ~n65799 ;
  assign n66057 = \P1_P2_Datao_reg[14]/NET0131  & n65799 ;
  assign n66058 = ~n66056 & ~n66057 ;
  assign n66059 = ~n65791 & ~n66058 ;
  assign n66060 = \P1_P1_Datao_reg[14]/NET0131  & n65791 ;
  assign n66061 = ~n66059 & ~n66060 ;
  assign n66062 = \P1_buf1_reg[15]/NET0131  & ~n65799 ;
  assign n66063 = \P1_P2_Datao_reg[15]/NET0131  & n65799 ;
  assign n66064 = ~n66062 & ~n66063 ;
  assign n66065 = ~n65791 & ~n66064 ;
  assign n66066 = \P1_P1_Datao_reg[15]/NET0131  & n65791 ;
  assign n66067 = ~n66065 & ~n66066 ;
  assign n66068 = \P1_buf1_reg[18]/NET0131  & ~n65799 ;
  assign n66069 = \P1_P2_Datao_reg[18]/NET0131  & n65799 ;
  assign n66070 = ~n66068 & ~n66069 ;
  assign n66071 = ~n65791 & ~n66070 ;
  assign n66072 = \P1_P1_Datao_reg[18]/NET0131  & n65791 ;
  assign n66073 = ~n66071 & ~n66072 ;
  assign n66074 = \P1_buf1_reg[19]/NET0131  & ~n65799 ;
  assign n66075 = \P1_P2_Datao_reg[19]/NET0131  & n65799 ;
  assign n66076 = ~n66074 & ~n66075 ;
  assign n66077 = ~n65791 & ~n66076 ;
  assign n66078 = \P1_P1_Datao_reg[19]/NET0131  & n65791 ;
  assign n66079 = ~n66077 & ~n66078 ;
  assign n66080 = \P1_buf1_reg[21]/NET0131  & ~n65799 ;
  assign n66081 = \P1_P2_Datao_reg[21]/NET0131  & n65799 ;
  assign n66082 = ~n66080 & ~n66081 ;
  assign n66083 = ~n65791 & ~n66082 ;
  assign n66084 = \P1_P1_Datao_reg[21]/NET0131  & n65791 ;
  assign n66085 = ~n66083 & ~n66084 ;
  assign n66086 = \P1_buf1_reg[22]/NET0131  & ~n65799 ;
  assign n66087 = \P1_P2_Datao_reg[22]/NET0131  & n65799 ;
  assign n66088 = ~n66086 & ~n66087 ;
  assign n66089 = ~n65791 & ~n66088 ;
  assign n66090 = \P1_P1_Datao_reg[22]/NET0131  & n65791 ;
  assign n66091 = ~n66089 & ~n66090 ;
  assign n66092 = \P1_buf1_reg[24]/NET0131  & ~n65799 ;
  assign n66093 = \P1_P2_Datao_reg[24]/NET0131  & n65799 ;
  assign n66094 = ~n66092 & ~n66093 ;
  assign n66095 = ~n65791 & ~n66094 ;
  assign n66096 = \P1_P1_Datao_reg[24]/NET0131  & n65791 ;
  assign n66097 = ~n66095 & ~n66096 ;
  assign n66098 = \P1_buf1_reg[25]/NET0131  & ~n65799 ;
  assign n66099 = \P1_P2_Datao_reg[25]/NET0131  & n65799 ;
  assign n66100 = ~n66098 & ~n66099 ;
  assign n66101 = ~n65791 & ~n66100 ;
  assign n66102 = \P1_P1_Datao_reg[25]/NET0131  & n65791 ;
  assign n66103 = ~n66101 & ~n66102 ;
  assign n66104 = \P1_buf1_reg[29]/NET0131  & ~n65799 ;
  assign n66105 = \P1_P2_Datao_reg[29]/NET0131  & n65799 ;
  assign n66106 = ~n66104 & ~n66105 ;
  assign n66107 = ~n65791 & ~n66106 ;
  assign n66108 = \P1_P1_Datao_reg[29]/NET0131  & n65791 ;
  assign n66109 = ~n66107 & ~n66108 ;
  assign n66110 = \P1_buf1_reg[2]/NET0131  & ~n65799 ;
  assign n66111 = \P1_P2_Datao_reg[2]/NET0131  & n65799 ;
  assign n66112 = ~n66110 & ~n66111 ;
  assign n66113 = ~n65791 & ~n66112 ;
  assign n66114 = \P1_P1_Datao_reg[2]/NET0131  & n65791 ;
  assign n66115 = ~n66113 & ~n66114 ;
  assign n66116 = \P1_buf1_reg[3]/NET0131  & ~n65799 ;
  assign n66117 = \P1_P2_Datao_reg[3]/NET0131  & n65799 ;
  assign n66118 = ~n66116 & ~n66117 ;
  assign n66119 = ~n65791 & ~n66118 ;
  assign n66120 = \P1_P1_Datao_reg[3]/NET0131  & n65791 ;
  assign n66121 = ~n66119 & ~n66120 ;
  assign n66122 = \P1_buf1_reg[6]/NET0131  & ~n65799 ;
  assign n66123 = \P1_P2_Datao_reg[6]/NET0131  & n65799 ;
  assign n66124 = ~n66122 & ~n66123 ;
  assign n66125 = ~n65791 & ~n66124 ;
  assign n66126 = \P1_P1_Datao_reg[6]/NET0131  & n65791 ;
  assign n66127 = ~n66125 & ~n66126 ;
  assign n66128 = \P1_buf1_reg[7]/NET0131  & ~n65799 ;
  assign n66129 = \P1_P2_Datao_reg[7]/NET0131  & n65799 ;
  assign n66130 = ~n66128 & ~n66129 ;
  assign n66131 = ~n65791 & ~n66130 ;
  assign n66132 = \P1_P1_Datao_reg[7]/NET0131  & n65791 ;
  assign n66133 = ~n66131 & ~n66132 ;
  assign n66134 = \P1_buf1_reg[8]/NET0131  & ~n65799 ;
  assign n66135 = \P1_P2_Datao_reg[8]/NET0131  & n65799 ;
  assign n66136 = ~n66134 & ~n66135 ;
  assign n66137 = ~n65791 & ~n66136 ;
  assign n66138 = \P1_P1_Datao_reg[8]/NET0131  & n65791 ;
  assign n66139 = ~n66137 & ~n66138 ;
  assign n66140 = \P1_buf1_reg[9]/NET0131  & ~n65799 ;
  assign n66141 = \P1_P2_Datao_reg[9]/NET0131  & n65799 ;
  assign n66142 = ~n66140 & ~n66141 ;
  assign n66143 = ~n65791 & ~n66142 ;
  assign n66144 = \P1_P1_Datao_reg[9]/NET0131  & n65791 ;
  assign n66145 = ~n66143 & ~n66144 ;
  assign n66146 = \P1_buf1_reg[30]/NET0131  & ~n65799 ;
  assign n66147 = \P1_P2_Datao_reg[30]/NET0131  & n65799 ;
  assign n66148 = ~n66146 & ~n66147 ;
  assign n66149 = ~n65791 & ~n66148 ;
  assign n66150 = \P1_P1_Datao_reg[30]/NET0131  & n65791 ;
  assign n66151 = ~n66149 & ~n66150 ;
  assign n66152 = \P1_buf1_reg[20]/NET0131  & ~n65799 ;
  assign n66153 = \P1_P2_Datao_reg[20]/NET0131  & n65799 ;
  assign n66154 = ~n66152 & ~n66153 ;
  assign n66155 = ~n65791 & ~n66154 ;
  assign n66156 = \P1_P1_Datao_reg[20]/NET0131  & n65791 ;
  assign n66157 = ~n66155 & ~n66156 ;
  assign n66158 = \P1_buf1_reg[0]/NET0131  & ~n65799 ;
  assign n66159 = \P1_P2_Datao_reg[0]/NET0131  & n65799 ;
  assign n66160 = ~n66158 & ~n66159 ;
  assign n66161 = ~n65791 & ~n66160 ;
  assign n66162 = \P1_P1_Datao_reg[0]/NET0131  & n65791 ;
  assign n66163 = ~n66161 & ~n66162 ;
  assign n66164 = \P1_buf1_reg[28]/NET0131  & ~n65799 ;
  assign n66165 = \P1_P2_Datao_reg[28]/NET0131  & n65799 ;
  assign n66166 = ~n66164 & ~n66165 ;
  assign n66167 = ~n65791 & ~n66166 ;
  assign n66168 = \P1_P1_Datao_reg[28]/NET0131  & n65791 ;
  assign n66169 = ~n66167 & ~n66168 ;
  assign n66170 = \P1_buf1_reg[27]/NET0131  & ~n65799 ;
  assign n66171 = \P1_P2_Datao_reg[27]/NET0131  & n65799 ;
  assign n66172 = ~n66170 & ~n66171 ;
  assign n66173 = ~n65791 & ~n66172 ;
  assign n66174 = \P1_P1_Datao_reg[27]/NET0131  & n65791 ;
  assign n66175 = ~n66173 & ~n66174 ;
  assign n66176 = \P1_buf1_reg[4]/NET0131  & ~n65799 ;
  assign n66177 = \P1_P2_Datao_reg[4]/NET0131  & n65799 ;
  assign n66178 = ~n66176 & ~n66177 ;
  assign n66179 = ~n65791 & ~n66178 ;
  assign n66180 = \P1_P1_Datao_reg[4]/NET0131  & n65791 ;
  assign n66181 = ~n66179 & ~n66180 ;
  assign n66182 = \P1_buf1_reg[26]/NET0131  & ~n65799 ;
  assign n66183 = \P1_P2_Datao_reg[26]/NET0131  & n65799 ;
  assign n66184 = ~n66182 & ~n66183 ;
  assign n66185 = ~n65791 & ~n66184 ;
  assign n66186 = \P1_P1_Datao_reg[26]/NET0131  & n65791 ;
  assign n66187 = ~n66185 & ~n66186 ;
  assign n66188 = \P3_rd_reg/NET0131  & \P4_IR_reg[16]/NET0131  ;
  assign n66189 = \P2_P3_Datao_reg[16]/NET0131  & ~\P3_rd_reg/NET0131  ;
  assign n66190 = ~n66188 & ~n66189 ;
  assign n66191 = \P3_rd_reg/NET0131  & \P4_IR_reg[20]/NET0131  ;
  assign n66192 = \P2_P3_Datao_reg[20]/NET0131  & ~\P3_rd_reg/NET0131  ;
  assign n66193 = ~n66191 & ~n66192 ;
  assign n66194 = \P2_P3_Datao_reg[23]/NET0131  & ~\P3_rd_reg/NET0131  ;
  assign n66195 = ~n15744 & ~n66194 ;
  assign n66197 = ~\P2_P2_rEIP_reg[15]/NET0131  & ~n63991 ;
  assign n66198 = n63373 & ~n63992 ;
  assign n66199 = ~n66197 & n66198 ;
  assign n66196 = \P2_P2_Address_reg[14]/NET0131  & ~n26646 ;
  assign n66200 = ~\P2_P2_rEIP_reg[16]/NET0131  & ~n65439 ;
  assign n66201 = n26647 & ~n65440 ;
  assign n66202 = ~n66200 & n66201 ;
  assign n66203 = ~n66196 & ~n66202 ;
  assign n66204 = ~n66199 & n66203 ;
  assign n66206 = ~\P1_P1_rEIP_reg[16]/NET0131  & ~n64007 ;
  assign n66207 = n26155 & ~n64008 ;
  assign n66208 = ~n66206 & n66207 ;
  assign n66205 = \P1_P1_Address_reg[14]/NET0131  & ~n26154 ;
  assign n66209 = ~\P1_P1_rEIP_reg[15]/NET0131  & ~n63406 ;
  assign n66210 = n63401 & ~n65459 ;
  assign n66211 = ~n66209 & n66210 ;
  assign n66212 = ~n66205 & ~n66211 ;
  assign n66213 = ~n66208 & n66212 ;
  assign n66215 = ~\P1_P3_rEIP_reg[16]/NET0131  & ~n64074 ;
  assign n66216 = n9092 & ~n64075 ;
  assign n66217 = ~n66215 & n66216 ;
  assign n66214 = \P1_P3_Address_reg[14]/NET0131  & ~n9091 ;
  assign n66218 = ~\P1_P3_rEIP_reg[15]/NET0131  & ~n64084 ;
  assign n66219 = n22115 & ~n64085 ;
  assign n66220 = ~n66218 & n66219 ;
  assign n66221 = ~n66214 & ~n66220 ;
  assign n66222 = ~n66217 & n66221 ;
  assign n66224 = ~\P1_P2_rEIP_reg[16]/NET0131  & ~n64033 ;
  assign n66225 = n25765 & ~n65480 ;
  assign n66226 = ~n66224 & n66225 ;
  assign n66223 = \P1_P2_Address_reg[14]/NET0131  & ~n25764 ;
  assign n66227 = ~\P1_P2_rEIP_reg[15]/NET0131  & ~n64024 ;
  assign n66228 = n51200 & n65544 ;
  assign n66229 = n63420 & ~n66228 ;
  assign n66230 = ~n66227 & n66229 ;
  assign n66231 = ~n66223 & ~n66230 ;
  assign n66232 = ~n66226 & n66231 ;
  assign n66234 = ~\P2_P3_rEIP_reg[16]/NET0131  & ~n64116 ;
  assign n66235 = n27145 & ~n64117 ;
  assign n66236 = ~n66234 & n66235 ;
  assign n66233 = \P2_P3_Address_reg[14]/NET0131  & ~n27144 ;
  assign n66237 = n52559 & n64095 ;
  assign n66238 = ~\P2_P3_rEIP_reg[15]/NET0131  & ~n66237 ;
  assign n66239 = n64094 & ~n65429 ;
  assign n66240 = ~n66238 & n66239 ;
  assign n66241 = ~n66233 & ~n66240 ;
  assign n66242 = ~n66236 & n66241 ;
  assign n66244 = ~\P2_P1_rEIP_reg[16]/NET0131  & ~n65499 ;
  assign n66245 = n25955 & ~n65500 ;
  assign n66246 = ~n66244 & n66245 ;
  assign n66243 = \P2_P1_Address_reg[14]/NET0131  & ~n25954 ;
  assign n66247 = ~\P2_P1_rEIP_reg[15]/NET0131  & ~n64050 ;
  assign n66248 = n63480 & ~n65504 ;
  assign n66249 = ~n66247 & n66248 ;
  assign n66250 = ~n66243 & ~n66249 ;
  assign n66251 = ~n66246 & n66250 ;
  assign n66253 = ~\P2_P2_rEIP_reg[28]/NET0131  & ~n63361 ;
  assign n66254 = n26647 & ~n63362 ;
  assign n66255 = ~n66253 & n66254 ;
  assign n66252 = \P2_P2_Address_reg[26]/NET0131  & ~n26646 ;
  assign n66256 = ~\P2_P2_rEIP_reg[27]/NET0131  & ~n63369 ;
  assign n66257 = ~n63370 & n63373 ;
  assign n66258 = ~n66256 & n66257 ;
  assign n66259 = ~n66252 & ~n66258 ;
  assign n66260 = ~n66255 & n66259 ;
  assign n66262 = \P1_P1_rEIP_reg[27]/NET0131  & n63395 ;
  assign n66263 = ~\P1_P1_rEIP_reg[28]/NET0131  & ~n66262 ;
  assign n66264 = n26155 & ~n65470 ;
  assign n66265 = ~n66263 & n66264 ;
  assign n66261 = \P1_P1_Address_reg[26]/NET0131  & ~n26154 ;
  assign n66266 = ~\P1_P1_rEIP_reg[27]/NET0131  & ~n63413 ;
  assign n66267 = n63401 & ~n63408 ;
  assign n66268 = ~n66266 & n66267 ;
  assign n66269 = ~n66261 & ~n66268 ;
  assign n66270 = ~n66265 & n66269 ;
  assign n66272 = n51313 & n64033 ;
  assign n66273 = n51516 & n66272 ;
  assign n66275 = \P1_P2_rEIP_reg[28]/NET0131  & n66273 ;
  assign n66274 = ~\P1_P2_rEIP_reg[28]/NET0131  & ~n66273 ;
  assign n66276 = n25765 & ~n66274 ;
  assign n66277 = ~n66275 & n66276 ;
  assign n66271 = \P1_P2_Address_reg[26]/NET0131  & ~n25764 ;
  assign n66278 = n51310 & n63421 ;
  assign n66279 = n48376 & n66278 ;
  assign n66281 = ~\P1_P2_rEIP_reg[27]/NET0131  & ~n66279 ;
  assign n66280 = \P1_P2_rEIP_reg[27]/NET0131  & n66279 ;
  assign n66282 = n63420 & ~n66280 ;
  assign n66283 = ~n66281 & n66282 ;
  assign n66284 = ~n66271 & ~n66283 ;
  assign n66285 = ~n66277 & n66284 ;
  assign n66290 = ~\P2_P1_rEIP_reg[27]/NET0131  & ~n63477 ;
  assign n66291 = n63480 & ~n65514 ;
  assign n66292 = ~n66290 & n66291 ;
  assign n66286 = \P2_P1_Address_reg[26]/NET0131  & ~n25954 ;
  assign n66287 = ~\P2_P1_rEIP_reg[28]/NET0131  & ~n63468 ;
  assign n66288 = n25955 & ~n63469 ;
  assign n66289 = ~n66287 & n66288 ;
  assign n66293 = ~n66286 & ~n66289 ;
  assign n66294 = ~n66292 & n66293 ;
  assign n66300 = \P2_P2_rEIP_reg[22]/NET0131  & n65228 ;
  assign n66301 = ~\P2_P2_rEIP_reg[23]/NET0131  & ~n66300 ;
  assign n66302 = n63373 & ~n65528 ;
  assign n66303 = ~n66301 & n66302 ;
  assign n66295 = \P2_P2_Address_reg[22]/NET0131  & ~n26646 ;
  assign n66296 = \P2_P2_rEIP_reg[23]/NET0131  & n65232 ;
  assign n66297 = ~\P2_P2_rEIP_reg[24]/NET0131  & ~n66296 ;
  assign n66298 = n26647 & ~n65524 ;
  assign n66299 = ~n66297 & n66298 ;
  assign n66304 = ~n66295 & ~n66299 ;
  assign n66305 = ~n66303 & n66304 ;
  assign n66311 = ~\P1_P1_rEIP_reg[24]/NET0131  & ~n63394 ;
  assign n66312 = n26155 & ~n64776 ;
  assign n66313 = ~n66311 & n66312 ;
  assign n66306 = \P1_P1_Address_reg[22]/NET0131  & ~n26154 ;
  assign n66307 = n51774 & n63402 ;
  assign n66308 = ~\P1_P1_rEIP_reg[23]/NET0131  & ~n66307 ;
  assign n66309 = n63401 & ~n63407 ;
  assign n66310 = ~n66308 & n66309 ;
  assign n66314 = ~n66306 & ~n66310 ;
  assign n66315 = ~n66313 & n66314 ;
  assign n66322 = \P1_P2_rEIP_reg[24]/NET0131  & n66272 ;
  assign n66321 = ~\P1_P2_rEIP_reg[24]/NET0131  & ~n66272 ;
  assign n66323 = n25765 & ~n66321 ;
  assign n66324 = ~n66322 & n66323 ;
  assign n66316 = \P1_P2_Address_reg[22]/NET0131  & ~n25764 ;
  assign n66318 = \P1_P2_rEIP_reg[23]/NET0131  & n66278 ;
  assign n66317 = ~\P1_P2_rEIP_reg[23]/NET0131  & ~n66278 ;
  assign n66319 = n63420 & ~n66317 ;
  assign n66320 = ~n66318 & n66319 ;
  assign n66325 = ~n66316 & ~n66320 ;
  assign n66326 = ~n66324 & n66325 ;
  assign n66329 = ~n50896 & n63475 ;
  assign n66328 = ~\P2_P1_rEIP_reg[23]/NET0131  & ~n63475 ;
  assign n66330 = n63480 & ~n66328 ;
  assign n66331 = ~n66329 & n66330 ;
  assign n66327 = \P2_P1_Address_reg[22]/NET0131  & ~n25954 ;
  assign n66332 = ~\P2_P1_rEIP_reg[24]/NET0131  & ~n63465 ;
  assign n66333 = n25955 & ~n65560 ;
  assign n66334 = ~n66332 & n66333 ;
  assign n66335 = ~n66327 & ~n66334 ;
  assign n66336 = ~n66331 & n66335 ;
  assign n66337 = \P3_rd_reg/NET0131  & \P4_IR_reg[12]/NET0131  ;
  assign n66338 = \P2_P3_Datao_reg[12]/NET0131  & ~\P3_rd_reg/NET0131  ;
  assign n66339 = ~n66337 & ~n66338 ;
  assign n66340 = \P3_rd_reg/NET0131  & \P4_IR_reg[15]/NET0131  ;
  assign n66341 = \P2_P3_Datao_reg[15]/NET0131  & ~\P3_rd_reg/NET0131  ;
  assign n66342 = ~n66340 & ~n66341 ;
  assign n66344 = \P2_P3_State_reg[2]/NET0131  & hold_pad ;
  assign n66347 = ~\P2_P3_RequestPending_reg/NET0131  & ~hold_pad ;
  assign n66348 = \P2_P3_State_reg[0]/NET0131  & \P2_P3_State_reg[1]/NET0131  ;
  assign n66349 = ~n66347 & n66348 ;
  assign n66350 = ~n66344 & n66349 ;
  assign n66351 = ~n27192 & ~n66350 ;
  assign n66352 = ~n64094 & ~n66348 ;
  assign n66353 = ~n66351 & ~n66352 ;
  assign n66343 = \P2_P3_State_reg[0]/NET0131  & ~\P2_P3_State_reg[1]/NET0131  ;
  assign n66345 = \P2_P3_RequestPending_reg/NET0131  & ~n66344 ;
  assign n66346 = n66343 & n66345 ;
  assign n66354 = n27148 & ~n66346 ;
  assign n66355 = ~n66353 & n66354 ;
  assign n66359 = ~\P2_P3_State_reg[2]/NET0131  & n66348 ;
  assign n66360 = ~hold_pad & ~n27192 ;
  assign n66361 = \P2_P3_RequestPending_reg/NET0131  & n66360 ;
  assign n66362 = n66359 & ~n66361 ;
  assign n66356 = \P2_P3_State_reg[2]/NET0131  & n66348 ;
  assign n66357 = ~n66343 & ~n66356 ;
  assign n66358 = ~n66345 & ~n66357 ;
  assign n66363 = ~n27145 & ~n27146 ;
  assign n66364 = ~hold_pad & ~na_pad ;
  assign n66365 = \P2_P3_RequestPending_reg/NET0131  & \P2_P3_State_reg[2]/NET0131  ;
  assign n66366 = n66364 & n66365 ;
  assign n66367 = ~n66363 & ~n66366 ;
  assign n66368 = ~n66358 & ~n66367 ;
  assign n66369 = ~n66362 & n66368 ;
  assign n66371 = ~\P1_P1_rEIP_reg[12]/NET0131  & ~n63391 ;
  assign n66372 = n26155 & ~n65577 ;
  assign n66373 = ~n66371 & n66372 ;
  assign n66370 = \P1_P1_Address_reg[10]/NET0131  & ~n26154 ;
  assign n66374 = ~\P1_P1_rEIP_reg[11]/NET0131  & ~n63403 ;
  assign n66375 = n63401 & ~n63404 ;
  assign n66376 = ~n66374 & n66375 ;
  assign n66377 = ~n66370 & ~n66376 ;
  assign n66378 = ~n66373 & n66377 ;
  assign n66380 = ~\P2_P2_rEIP_reg[12]/NET0131  & ~n64821 ;
  assign n66381 = n26647 & ~n65587 ;
  assign n66382 = ~n66380 & n66381 ;
  assign n66379 = \P2_P2_Address_reg[10]/NET0131  & ~n26646 ;
  assign n66383 = n55777 & n63368 ;
  assign n66384 = ~\P2_P2_rEIP_reg[11]/NET0131  & ~n66383 ;
  assign n66385 = n63373 & ~n63989 ;
  assign n66386 = ~n66384 & n66385 ;
  assign n66387 = ~n66379 & ~n66386 ;
  assign n66388 = ~n66382 & n66387 ;
  assign n66394 = ~\P1_P3_rEIP_reg[12]/NET0131  & ~n64070 ;
  assign n66395 = n9092 & ~n64071 ;
  assign n66396 = ~n66394 & n66395 ;
  assign n66389 = \P1_P3_Address_reg[10]/NET0131  & ~n9091 ;
  assign n66391 = ~n17698 & n64081 ;
  assign n66390 = ~\P1_P3_rEIP_reg[11]/NET0131  & ~n64081 ;
  assign n66392 = n22115 & ~n66390 ;
  assign n66393 = ~n66391 & n66392 ;
  assign n66397 = ~n66389 & ~n66393 ;
  assign n66398 = ~n66396 & n66397 ;
  assign n66400 = ~\P1_P2_rEIP_reg[12]/NET0131  & ~n64032 ;
  assign n66401 = n25765 & ~n65607 ;
  assign n66402 = ~n66400 & n66401 ;
  assign n66399 = \P1_P2_Address_reg[10]/NET0131  & ~n25764 ;
  assign n66403 = ~\P1_P2_rEIP_reg[11]/NET0131  & ~n64023 ;
  assign n66404 = n63420 & ~n64848 ;
  assign n66405 = ~n66403 & n66404 ;
  assign n66406 = ~n66399 & ~n66405 ;
  assign n66407 = ~n66402 & n66406 ;
  assign n66413 = ~\P2_P3_rEIP_reg[12]/NET0131  & ~n64112 ;
  assign n66414 = n27145 & ~n64113 ;
  assign n66415 = ~n66413 & n66414 ;
  assign n66408 = \P2_P3_Address_reg[10]/NET0131  & ~n27144 ;
  assign n66410 = ~n56121 & n64095 ;
  assign n66409 = ~\P2_P3_rEIP_reg[11]/NET0131  & ~n64095 ;
  assign n66411 = n64094 & ~n66409 ;
  assign n66412 = ~n66410 & n66411 ;
  assign n66416 = ~n66408 & ~n66412 ;
  assign n66417 = ~n66415 & n66416 ;
  assign n66419 = ~\P2_P1_rEIP_reg[12]/NET0131  & ~n63461 ;
  assign n66420 = n25955 & ~n65567 ;
  assign n66421 = ~n66419 & n66420 ;
  assign n66418 = \P2_P1_Address_reg[10]/NET0131  & ~n25954 ;
  assign n66422 = n54867 & n63475 ;
  assign n66423 = ~\P2_P1_rEIP_reg[11]/NET0131  & ~n66422 ;
  assign n66424 = n63480 & ~n64049 ;
  assign n66425 = ~n66423 & n66424 ;
  assign n66426 = ~n66418 & ~n66425 ;
  assign n66427 = ~n66421 & n66426 ;
  assign n66428 = \P3_rd_reg/NET0131  & \P4_IR_reg[11]/NET0131  ;
  assign n66429 = \P2_P3_Datao_reg[11]/NET0131  & ~\P3_rd_reg/NET0131  ;
  assign n66430 = ~n66428 & ~n66429 ;
  assign n66431 = \P3_rd_reg/NET0131  & \P4_IR_reg[19]/NET0131  ;
  assign n66432 = \P2_P3_Datao_reg[19]/NET0131  & ~\P3_rd_reg/NET0131  ;
  assign n66433 = ~n66431 & ~n66432 ;
  assign n66434 = \P3_rd_reg/NET0131  & \P4_IR_reg[8]/NET0131  ;
  assign n66435 = \P2_P3_Datao_reg[8]/NET0131  & ~\P3_rd_reg/NET0131  ;
  assign n66436 = ~n66434 & ~n66435 ;
  assign n66437 = ~n65791 & n65799 ;
  assign n66438 = ~n65813 & n65821 ;
  assign n66440 = ~\P2_P2_rEIP_reg[4]/NET0131  & ~n63353 ;
  assign n66441 = n26647 & ~n63354 ;
  assign n66442 = ~n66440 & n66441 ;
  assign n66439 = \P2_P2_Address_reg[2]/NET0131  & ~n26646 ;
  assign n66443 = ~\P2_P2_rEIP_reg[3]/NET0131  & ~n65337 ;
  assign n66444 = n63373 & ~n65338 ;
  assign n66445 = ~n66443 & n66444 ;
  assign n66446 = ~n66439 & ~n66445 ;
  assign n66447 = ~n66442 & n66446 ;
  assign n66449 = ~\P1_P3_rEIP_reg[4]/NET0131  & ~n64062 ;
  assign n66450 = n9092 & ~n64063 ;
  assign n66451 = ~n66449 & n66450 ;
  assign n66448 = \P1_P3_Address_reg[2]/NET0131  & ~n9091 ;
  assign n66452 = ~\P1_P3_rEIP_reg[3]/NET0131  & ~n65348 ;
  assign n66453 = n22115 & ~n65349 ;
  assign n66454 = ~n66452 & n66453 ;
  assign n66455 = ~n66448 & ~n66454 ;
  assign n66456 = ~n66451 & n66455 ;
  assign n66458 = ~\P1_P1_rEIP_reg[4]/NET0131  & ~n63383 ;
  assign n66459 = n26155 & ~n63384 ;
  assign n66460 = ~n66458 & n66459 ;
  assign n66457 = \P1_P1_Address_reg[2]/NET0131  & ~n26154 ;
  assign n66461 = ~\P1_P1_rEIP_reg[3]/NET0131  & ~n65365 ;
  assign n66462 = n63401 & ~n65366 ;
  assign n66463 = ~n66461 & n66462 ;
  assign n66464 = ~n66457 & ~n66463 ;
  assign n66465 = ~n66460 & n66464 ;
  assign n66467 = ~\P1_P2_rEIP_reg[4]/NET0131  & ~n63430 ;
  assign n66468 = n25765 & ~n63431 ;
  assign n66469 = ~n66467 & n66468 ;
  assign n66466 = \P1_P2_Address_reg[2]/NET0131  & ~n25764 ;
  assign n66470 = ~\P1_P2_rEIP_reg[3]/NET0131  & ~n65393 ;
  assign n66471 = n63420 & ~n65394 ;
  assign n66472 = ~n66470 & n66471 ;
  assign n66473 = ~n66466 & ~n66472 ;
  assign n66474 = ~n66469 & n66473 ;
  assign n66476 = ~\P2_P3_rEIP_reg[4]/NET0131  & ~n64104 ;
  assign n66477 = n27145 & ~n64105 ;
  assign n66478 = ~n66476 & n66477 ;
  assign n66475 = \P2_P3_Address_reg[2]/NET0131  & ~n27144 ;
  assign n66479 = ~\P2_P3_rEIP_reg[3]/NET0131  & ~n65379 ;
  assign n66480 = n64094 & ~n65380 ;
  assign n66481 = ~n66479 & n66480 ;
  assign n66482 = ~n66475 & ~n66481 ;
  assign n66483 = ~n66478 & n66482 ;
  assign n66485 = ~\P2_P1_rEIP_reg[4]/NET0131  & ~n63454 ;
  assign n66486 = n25955 & ~n63455 ;
  assign n66487 = ~n66485 & n66486 ;
  assign n66484 = \P2_P1_Address_reg[2]/NET0131  & ~n25954 ;
  assign n66488 = ~\P2_P1_rEIP_reg[3]/NET0131  & ~n65407 ;
  assign n66489 = n63480 & ~n65408 ;
  assign n66490 = ~n66488 & n66489 ;
  assign n66491 = ~n66484 & ~n66490 ;
  assign n66492 = ~n66487 & n66491 ;
  assign n66497 = \P2_P2_rEIP_reg[18]/NET0131  & n63995 ;
  assign n66498 = ~\P2_P2_rEIP_reg[19]/NET0131  & ~n66497 ;
  assign n66499 = n63373 & ~n66498 ;
  assign n66500 = ~n65225 & n66499 ;
  assign n66493 = \P2_P2_Address_reg[18]/NET0131  & ~n26646 ;
  assign n66494 = ~\P2_P2_rEIP_reg[20]/NET0131  & ~n65687 ;
  assign n66495 = n26647 & ~n65688 ;
  assign n66496 = ~n66494 & n66495 ;
  assign n66501 = ~n66493 & ~n66496 ;
  assign n66502 = ~n66500 & n66501 ;
  assign n66508 = ~\P1_P1_rEIP_reg[20]/NET0131  & ~n65699 ;
  assign n66509 = n26155 & ~n65700 ;
  assign n66510 = ~n66508 & n66509 ;
  assign n66503 = \P1_P1_Address_reg[18]/NET0131  & ~n26154 ;
  assign n66504 = n51665 & n64014 ;
  assign n66505 = ~\P1_P1_rEIP_reg[19]/NET0131  & ~n66504 ;
  assign n66506 = n63401 & ~n65695 ;
  assign n66507 = ~n66505 & n66506 ;
  assign n66511 = ~n66503 & ~n66507 ;
  assign n66512 = ~n66510 & n66511 ;
  assign n66517 = n48389 & n64845 ;
  assign n66518 = \P1_P2_rEIP_reg[19]/NET0131  & n66517 ;
  assign n66520 = \P1_P2_rEIP_reg[20]/NET0131  & n66518 ;
  assign n66519 = ~\P1_P2_rEIP_reg[20]/NET0131  & ~n66518 ;
  assign n66521 = n25765 & ~n66519 ;
  assign n66522 = ~n66520 & n66521 ;
  assign n66513 = \P1_P2_Address_reg[18]/NET0131  & ~n25764 ;
  assign n66514 = ~\P1_P2_rEIP_reg[19]/NET0131  & ~n65252 ;
  assign n66515 = n63420 & ~n65707 ;
  assign n66516 = ~n66514 & n66515 ;
  assign n66523 = ~n66513 & ~n66516 ;
  assign n66524 = ~n66522 & n66523 ;
  assign n66526 = \P2_P1_rEIP_reg[19]/NET0131  & n64042 ;
  assign n66527 = ~\P2_P1_rEIP_reg[20]/NET0131  & ~n66526 ;
  assign n66528 = n25955 & ~n63464 ;
  assign n66529 = ~n66527 & n66528 ;
  assign n66525 = \P2_P1_Address_reg[18]/NET0131  & ~n25954 ;
  assign n66530 = n50777 & n63475 ;
  assign n66531 = ~\P2_P1_rEIP_reg[19]/NET0131  & ~n66530 ;
  assign n66532 = n63480 & ~n65719 ;
  assign n66533 = ~n66531 & n66532 ;
  assign n66534 = ~n66525 & ~n66533 ;
  assign n66535 = ~n66529 & n66534 ;
  assign n66542 = \P1_P3_rEIP_reg[19]/NET0131  & n64078 ;
  assign n66544 = \P1_P3_rEIP_reg[20]/NET0131  & n66542 ;
  assign n66543 = ~\P1_P3_rEIP_reg[20]/NET0131  & ~n66542 ;
  assign n66545 = n9092 & ~n66543 ;
  assign n66546 = ~n66544 & n66545 ;
  assign n66536 = \P1_P3_Address_reg[18]/NET0131  & ~n9091 ;
  assign n66539 = n16585 & n64081 ;
  assign n66537 = \P1_P3_rEIP_reg[18]/NET0131  & n64087 ;
  assign n66538 = ~\P1_P3_rEIP_reg[19]/NET0131  & ~n66537 ;
  assign n66540 = n22115 & ~n66538 ;
  assign n66541 = ~n66539 & n66540 ;
  assign n66547 = ~n66536 & ~n66541 ;
  assign n66548 = ~n66546 & n66547 ;
  assign n66554 = \P2_P3_rEIP_reg[19]/NET0131  & n64119 ;
  assign n66556 = \P2_P3_rEIP_reg[20]/NET0131  & n66554 ;
  assign n66555 = ~\P2_P3_rEIP_reg[20]/NET0131  & ~n66554 ;
  assign n66557 = n27145 & ~n66555 ;
  assign n66558 = ~n66556 & n66557 ;
  assign n66549 = \P2_P3_Address_reg[18]/NET0131  & ~n27144 ;
  assign n66551 = ~n56279 & n64095 ;
  assign n66550 = ~\P2_P3_rEIP_reg[19]/NET0131  & ~n64095 ;
  assign n66552 = n64094 & ~n66550 ;
  assign n66553 = ~n66551 & n66552 ;
  assign n66559 = ~n66549 & ~n66553 ;
  assign n66560 = ~n66558 & n66559 ;
  assign n66562 = ~\P2_P1_rEIP_reg[8]/NET0131  & ~n63458 ;
  assign n66563 = n25955 & ~n63459 ;
  assign n66564 = ~n66562 & n66563 ;
  assign n66561 = \P2_P1_Address_reg[6]/NET0131  & ~n25954 ;
  assign n66565 = ~\P2_P1_rEIP_reg[7]/NET0131  & ~n64045 ;
  assign n66566 = n63480 & ~n64046 ;
  assign n66567 = ~n66565 & n66566 ;
  assign n66568 = ~n66561 & ~n66567 ;
  assign n66569 = ~n66564 & n66568 ;
  assign n66571 = ~\P2_P2_rEIP_reg[8]/NET0131  & ~n63357 ;
  assign n66572 = n26647 & ~n63358 ;
  assign n66573 = ~n66571 & n66572 ;
  assign n66570 = \P2_P2_Address_reg[6]/NET0131  & ~n26646 ;
  assign n66574 = ~\P2_P2_rEIP_reg[7]/NET0131  & ~n63985 ;
  assign n66575 = n63373 & ~n63986 ;
  assign n66576 = ~n66574 & n66575 ;
  assign n66577 = ~n66570 & ~n66576 ;
  assign n66578 = ~n66573 & n66577 ;
  assign n66580 = ~\P1_P1_rEIP_reg[8]/NET0131  & ~n63387 ;
  assign n66581 = n26155 & ~n63388 ;
  assign n66582 = ~n66580 & n66581 ;
  assign n66579 = \P1_P1_Address_reg[6]/NET0131  & ~n26154 ;
  assign n66583 = ~\P1_P1_rEIP_reg[7]/NET0131  & ~n65287 ;
  assign n66584 = n63401 & ~n65288 ;
  assign n66585 = ~n66583 & n66584 ;
  assign n66586 = ~n66579 & ~n66585 ;
  assign n66587 = ~n66582 & n66586 ;
  assign n66589 = ~\P2_P3_rEIP_reg[8]/NET0131  & ~n64108 ;
  assign n66590 = n27145 & ~n64109 ;
  assign n66591 = ~n66589 & n66590 ;
  assign n66588 = \P2_P3_Address_reg[6]/NET0131  & ~n27144 ;
  assign n66592 = ~\P2_P3_rEIP_reg[7]/NET0131  & ~n65300 ;
  assign n66593 = n64094 & ~n65301 ;
  assign n66594 = ~n66592 & n66593 ;
  assign n66595 = ~n66588 & ~n66594 ;
  assign n66596 = ~n66591 & n66595 ;
  assign n66598 = ~\P1_P2_rEIP_reg[8]/NET0131  & ~n63434 ;
  assign n66599 = n25765 & ~n63435 ;
  assign n66600 = ~n66598 & n66599 ;
  assign n66597 = \P1_P2_Address_reg[6]/NET0131  & ~n25764 ;
  assign n66601 = n48384 & n63421 ;
  assign n66602 = ~\P1_P2_rEIP_reg[7]/NET0131  & ~n66601 ;
  assign n66603 = n63420 & ~n65544 ;
  assign n66604 = ~n66602 & n66603 ;
  assign n66605 = ~n66597 & ~n66604 ;
  assign n66606 = ~n66600 & n66605 ;
  assign n66612 = ~\P1_P3_rEIP_reg[8]/NET0131  & ~n64066 ;
  assign n66613 = n9092 & ~n64067 ;
  assign n66614 = ~n66612 & n66613 ;
  assign n66607 = \P1_P3_Address_reg[6]/NET0131  & ~n9091 ;
  assign n66609 = ~n17619 & n64081 ;
  assign n66608 = ~\P1_P3_rEIP_reg[7]/NET0131  & ~n64081 ;
  assign n66610 = n22115 & ~n66608 ;
  assign n66611 = ~n66609 & n66610 ;
  assign n66615 = ~n66607 & ~n66611 ;
  assign n66616 = ~n66614 & n66615 ;
  assign n66617 = \P3_rd_reg/NET0131  & \P4_IR_reg[30]/NET0131  ;
  assign n66618 = \P2_P3_Datao_reg[30]/NET0131  & ~\P3_rd_reg/NET0131  ;
  assign n66619 = ~n66617 & ~n66618 ;
  assign n66620 = \P3_rd_reg/NET0131  & \P4_IR_reg[4]/NET0131  ;
  assign n66621 = \P2_P3_Datao_reg[4]/NET0131  & ~\P3_rd_reg/NET0131  ;
  assign n66622 = ~n66620 & ~n66621 ;
  assign n66623 = \P3_rd_reg/NET0131  & \P4_IR_reg[7]/NET0131  ;
  assign n66624 = \P2_P3_Datao_reg[7]/NET0131  & ~\P3_rd_reg/NET0131  ;
  assign n66625 = ~n66623 & ~n66624 ;
  assign n66626 = ~\P2_P2_Address_reg[29]/NET0131  & n65820 ;
  assign n66629 = ~\P2_P3_BE_n_reg[3]/NET0131  & ~\P2_P3_D_C_n_reg/NET0131  ;
  assign n66630 = \P2_P3_M_IO_n_reg/NET0131  & ~\P2_P3_W_R_n_reg/NET0131  ;
  assign n66631 = n66629 & n66630 ;
  assign n66627 = ~\P2_P3_ADS_n_reg/NET0131  & ~\P2_P3_BE_n_reg[0]/NET0131  ;
  assign n66628 = ~\P2_P3_BE_n_reg[1]/NET0131  & ~\P2_P3_BE_n_reg[2]/NET0131  ;
  assign n66632 = n66627 & n66628 ;
  assign n66633 = n66631 & n66632 ;
  assign n66634 = ~n66626 & n66633 ;
  assign n66635 = ~\P1_P2_Address_reg[29]/NET0131  & n65798 ;
  assign n66638 = ~\P1_P3_BE_n_reg[3]/NET0131  & ~\P1_P3_D_C_n_reg/NET0131  ;
  assign n66639 = \P1_P3_M_IO_n_reg/NET0131  & ~\P1_P3_W_R_n_reg/NET0131  ;
  assign n66640 = n66638 & n66639 ;
  assign n66636 = ~\P1_P3_ADS_n_reg/NET0131  & ~\P1_P3_BE_n_reg[0]/NET0131  ;
  assign n66637 = ~\P1_P3_BE_n_reg[1]/NET0131  & ~\P1_P3_BE_n_reg[2]/NET0131  ;
  assign n66641 = n66636 & n66637 ;
  assign n66642 = n66640 & n66641 ;
  assign n66643 = ~n66635 & n66642 ;
  assign n66644 = ~\P2_P3_State_reg[2]/NET0131  & n66349 ;
  assign n66645 = n27192 & n66644 ;
  assign n66646 = ~n27147 & ~n66645 ;
  assign n66647 = ~na_pad & ~n66646 ;
  assign n66651 = n66356 & ~n66360 ;
  assign n66648 = \P2_P3_RequestPending_reg/NET0131  & ~\P2_P3_State_reg[2]/NET0131  ;
  assign n66649 = hold_pad & n66343 ;
  assign n66650 = ~n66648 & n66649 ;
  assign n66652 = ~n64094 & ~n66650 ;
  assign n66653 = ~n66651 & n66652 ;
  assign n66654 = ~n66647 & n66653 ;
  assign n66659 = ~\P2_P1_rEIP_reg[26]/NET0131  & ~n63476 ;
  assign n66660 = ~n63477 & n63480 ;
  assign n66661 = ~n66659 & n66660 ;
  assign n66655 = \P2_P1_Address_reg[25]/NET0131  & ~n25954 ;
  assign n66656 = ~\P2_P1_rEIP_reg[27]/NET0131  & ~n63467 ;
  assign n66657 = n25955 & ~n63468 ;
  assign n66658 = ~n66656 & n66657 ;
  assign n66662 = ~n66655 & ~n66658 ;
  assign n66663 = ~n66661 & n66662 ;
  assign n66665 = ~\P2_P2_rEIP_reg[27]/NET0131  & ~n63360 ;
  assign n66666 = n26647 & ~n63361 ;
  assign n66667 = ~n66665 & n66666 ;
  assign n66664 = \P2_P2_Address_reg[25]/NET0131  & ~n26646 ;
  assign n66668 = ~\P2_P2_rEIP_reg[26]/NET0131  & ~n64767 ;
  assign n66669 = ~n63369 & n63373 ;
  assign n66670 = ~n66668 & n66669 ;
  assign n66671 = ~n66664 & ~n66670 ;
  assign n66672 = ~n66667 & n66671 ;
  assign n66674 = ~\P1_P1_rEIP_reg[27]/NET0131  & ~n63395 ;
  assign n66675 = n26155 & ~n66262 ;
  assign n66676 = ~n66674 & n66675 ;
  assign n66673 = \P1_P1_Address_reg[25]/NET0131  & ~n26154 ;
  assign n66677 = ~\P1_P1_rEIP_reg[26]/NET0131  & ~n63412 ;
  assign n66678 = n63401 & ~n63413 ;
  assign n66679 = ~n66677 & n66678 ;
  assign n66680 = ~n66673 & ~n66679 ;
  assign n66681 = ~n66676 & n66680 ;
  assign n66689 = n48379 & n66517 ;
  assign n66690 = n48376 & n66689 ;
  assign n66692 = \P1_P2_rEIP_reg[27]/NET0131  & n66690 ;
  assign n66691 = ~\P1_P2_rEIP_reg[27]/NET0131  & ~n66690 ;
  assign n66693 = n25765 & ~n66691 ;
  assign n66694 = ~n66692 & n66693 ;
  assign n66682 = \P1_P2_Address_reg[25]/NET0131  & ~n25764 ;
  assign n66683 = n48379 & n65252 ;
  assign n66685 = n48375 & n66683 ;
  assign n66686 = ~\P1_P2_rEIP_reg[26]/NET0131  & ~n66685 ;
  assign n66684 = n48376 & n66683 ;
  assign n66687 = n63420 & ~n66684 ;
  assign n66688 = ~n66686 & n66687 ;
  assign n66695 = ~n66682 & ~n66688 ;
  assign n66696 = ~n66694 & n66695 ;
  assign n66703 = \P2_P2_rEIP_reg[31]/NET0131  & n63365 ;
  assign n66702 = ~\P2_P2_rEIP_reg[31]/NET0131  & ~n63365 ;
  assign n66704 = n26647 & ~n66702 ;
  assign n66705 = ~n66703 & n66704 ;
  assign n66697 = \P2_P2_Address_reg[29]/NET0131  & ~n26646 ;
  assign n66699 = \P2_P2_rEIP_reg[0]/NET0131  & n56655 ;
  assign n66698 = ~\P2_P2_rEIP_reg[30]/NET0131  & ~n63374 ;
  assign n66700 = n63373 & ~n66698 ;
  assign n66701 = ~n66699 & n66700 ;
  assign n66706 = ~n66697 & ~n66701 ;
  assign n66707 = ~n66705 & n66706 ;
  assign n66714 = \P1_P1_rEIP_reg[31]/NET0131  & n63398 ;
  assign n66713 = ~\P1_P1_rEIP_reg[31]/NET0131  & ~n63398 ;
  assign n66715 = n26155 & ~n66713 ;
  assign n66716 = ~n66714 & n66715 ;
  assign n66708 = \P1_P1_Address_reg[29]/NET0131  & ~n26154 ;
  assign n66710 = \P1_P1_rEIP_reg[30]/NET0131  & n63414 ;
  assign n66709 = ~\P1_P1_rEIP_reg[30]/NET0131  & ~n63414 ;
  assign n66711 = n63401 & ~n66709 ;
  assign n66712 = ~n66710 & n66711 ;
  assign n66717 = ~n66708 & ~n66712 ;
  assign n66718 = ~n66716 & n66717 ;
  assign n66720 = n48403 & n66692 ;
  assign n66722 = \P1_P2_rEIP_reg[31]/NET0131  & n66720 ;
  assign n66721 = ~\P1_P2_rEIP_reg[31]/NET0131  & ~n66720 ;
  assign n66723 = n25765 & ~n66721 ;
  assign n66724 = ~n66722 & n66723 ;
  assign n66719 = \P1_P2_Address_reg[29]/NET0131  & ~n25764 ;
  assign n66726 = ~n48405 & n63421 ;
  assign n66725 = ~\P1_P2_rEIP_reg[30]/NET0131  & ~n63421 ;
  assign n66727 = n63420 & ~n66725 ;
  assign n66728 = ~n66726 & n66727 ;
  assign n66729 = ~n66719 & ~n66728 ;
  assign n66730 = ~n66724 & n66729 ;
  assign n66737 = \P2_P1_rEIP_reg[31]/NET0131  & n63472 ;
  assign n66736 = ~\P2_P1_rEIP_reg[31]/NET0131  & ~n63472 ;
  assign n66738 = n25955 & ~n66736 ;
  assign n66739 = ~n66737 & n66738 ;
  assign n66731 = \P2_P1_Address_reg[29]/NET0131  & ~n25954 ;
  assign n66733 = \P2_P1_rEIP_reg[0]/NET0131  & n56483 ;
  assign n66732 = ~\P2_P1_rEIP_reg[30]/NET0131  & ~n63481 ;
  assign n66734 = n63480 & ~n66732 ;
  assign n66735 = ~n66733 & n66734 ;
  assign n66740 = ~n66731 & ~n66735 ;
  assign n66741 = ~n66739 & n66740 ;
  assign n66744 = \P1_P2_State_reg[1]/NET0131  & hold_pad ;
  assign n66745 = ~\P1_P2_RequestPending_reg/NET0131  & ~n66744 ;
  assign n66746 = ~\P1_P2_State_reg[2]/NET0131  & ~n66745 ;
  assign n66742 = \P1_P2_State_reg[1]/NET0131  & n25415 ;
  assign n66747 = \P1_P2_RequestPending_reg/NET0131  & ~hold_pad ;
  assign n66748 = ~n66742 & ~n66747 ;
  assign n66749 = ~n66746 & n66748 ;
  assign n66750 = \P1_P2_State_reg[0]/NET0131  & ~n66749 ;
  assign n66743 = \P1_P2_State_reg[2]/NET0131  & n66742 ;
  assign n66751 = n25768 & ~n66743 ;
  assign n66752 = ~n66750 & n66751 ;
  assign n66755 = \P2_P1_State_reg[1]/NET0131  & hold_pad ;
  assign n66756 = ~\P2_P1_RequestPending_reg/NET0131  & ~n66755 ;
  assign n66757 = ~\P2_P1_State_reg[2]/NET0131  & ~n66756 ;
  assign n66753 = \P2_P1_State_reg[1]/NET0131  & n21073 ;
  assign n66758 = \P2_P1_RequestPending_reg/NET0131  & ~hold_pad ;
  assign n66759 = ~n66753 & ~n66758 ;
  assign n66760 = ~n66757 & n66759 ;
  assign n66761 = \P2_P1_State_reg[0]/NET0131  & ~n66760 ;
  assign n66754 = \P2_P1_State_reg[2]/NET0131  & n66753 ;
  assign n66762 = n25958 & ~n66754 ;
  assign n66763 = ~n66761 & n66762 ;
  assign n66766 = \P1_P1_State_reg[1]/NET0131  & hold_pad ;
  assign n66767 = ~\P1_P1_RequestPending_reg/NET0131  & ~n66766 ;
  assign n66768 = ~\P1_P1_State_reg[2]/NET0131  & ~n66767 ;
  assign n66764 = \P1_P1_State_reg[1]/NET0131  & n15335 ;
  assign n66769 = \P1_P1_RequestPending_reg/NET0131  & ~hold_pad ;
  assign n66770 = ~n66764 & ~n66769 ;
  assign n66771 = ~n66768 & n66770 ;
  assign n66772 = \P1_P1_State_reg[0]/NET0131  & ~n66771 ;
  assign n66765 = \P1_P1_State_reg[2]/NET0131  & n66764 ;
  assign n66773 = n26158 & ~n66765 ;
  assign n66774 = ~n66772 & n66773 ;
  assign n66779 = ~hold_pad & ~n26286 ;
  assign n66780 = \P2_P2_State_reg[0]/NET0131  & ~n66779 ;
  assign n66781 = ~\P2_P2_State_reg[2]/NET0131  & ~n66780 ;
  assign n66778 = \P2_P2_State_reg[2]/NET0131  & ~n26286 ;
  assign n66782 = \P2_P2_State_reg[1]/NET0131  & ~n66778 ;
  assign n66783 = ~n66781 & n66782 ;
  assign n66775 = \P2_P2_State_reg[2]/NET0131  & hold_pad ;
  assign n66776 = \P2_P2_RequestPending_reg/NET0131  & ~n66775 ;
  assign n66777 = \P2_P2_State_reg[0]/NET0131  & n66776 ;
  assign n66784 = n26650 & ~n66777 ;
  assign n66785 = ~n66783 & n66784 ;
  assign n66786 = ~\P1_P2_RequestPending_reg/NET0131  & ~\P1_P2_State_reg[1]/NET0131  ;
  assign n66787 = ~\P1_P2_State_reg[2]/NET0131  & ~n66786 ;
  assign n66788 = \P1_P2_State_reg[0]/NET0131  & ~n66787 ;
  assign n66789 = ~n66747 & n66788 ;
  assign n66790 = ~n25415 & n66747 ;
  assign n66791 = \P1_P2_State_reg[1]/NET0131  & ~n66790 ;
  assign n66792 = \P1_P2_State_reg[0]/NET0131  & ~n66791 ;
  assign n66793 = \P1_P2_RequestPending_reg/NET0131  & n66364 ;
  assign n66794 = ~\P1_P2_State_reg[1]/NET0131  & ~n66793 ;
  assign n66795 = \P1_P2_State_reg[2]/NET0131  & ~n66794 ;
  assign n66796 = ~n66792 & ~n66795 ;
  assign n66797 = ~n66789 & ~n66796 ;
  assign n66798 = ~\P2_P1_RequestPending_reg/NET0131  & ~\P2_P1_State_reg[1]/NET0131  ;
  assign n66799 = ~\P2_P1_State_reg[2]/NET0131  & ~n66798 ;
  assign n66800 = \P2_P1_State_reg[0]/NET0131  & ~n66799 ;
  assign n66801 = ~n66758 & n66800 ;
  assign n66802 = ~n21073 & n66758 ;
  assign n66803 = \P2_P1_State_reg[1]/NET0131  & ~n66802 ;
  assign n66804 = \P2_P1_State_reg[0]/NET0131  & ~n66803 ;
  assign n66805 = \P2_P1_RequestPending_reg/NET0131  & n66364 ;
  assign n66806 = ~\P2_P1_State_reg[1]/NET0131  & ~n66805 ;
  assign n66807 = \P2_P1_State_reg[2]/NET0131  & ~n66806 ;
  assign n66808 = ~n66804 & ~n66807 ;
  assign n66809 = ~n66801 & ~n66808 ;
  assign n66811 = ~n15335 & n66769 ;
  assign n66812 = \P1_P1_State_reg[1]/NET0131  & ~n66811 ;
  assign n66813 = \P1_P1_State_reg[0]/NET0131  & ~n66812 ;
  assign n66814 = ~\P1_P1_State_reg[2]/NET0131  & ~n66813 ;
  assign n66810 = na_pad & n26157 ;
  assign n66817 = ~\P1_P1_RequestPending_reg/NET0131  & ~\P1_P1_State_reg[1]/NET0131  ;
  assign n66818 = ~\P1_P1_State_reg[2]/NET0131  & ~n66817 ;
  assign n66815 = ~\P1_P1_State_reg[1]/NET0131  & \P1_P1_State_reg[2]/NET0131  ;
  assign n66816 = ~\P1_P1_State_reg[0]/NET0131  & ~n66815 ;
  assign n66819 = ~n66769 & ~n66816 ;
  assign n66820 = ~n66818 & n66819 ;
  assign n66821 = ~n66810 & ~n66820 ;
  assign n66822 = ~n66814 & n66821 ;
  assign n66831 = ~n26647 & ~n26648 ;
  assign n66832 = \P2_P2_RequestPending_reg/NET0131  & \P2_P2_State_reg[2]/NET0131  ;
  assign n66833 = n66364 & n66832 ;
  assign n66834 = ~n66831 & ~n66833 ;
  assign n66823 = \P2_P2_State_reg[0]/NET0131  & \P2_P2_State_reg[1]/NET0131  ;
  assign n66824 = \P2_P2_State_reg[2]/NET0131  & n66823 ;
  assign n66825 = \P2_P2_State_reg[0]/NET0131  & ~\P2_P2_State_reg[1]/NET0131  ;
  assign n66826 = ~n66824 & ~n66825 ;
  assign n66827 = ~n66776 & ~n66826 ;
  assign n66828 = ~\P2_P2_State_reg[2]/NET0131  & n66823 ;
  assign n66829 = \P2_P2_RequestPending_reg/NET0131  & n66779 ;
  assign n66830 = n66828 & ~n66829 ;
  assign n66835 = ~n66827 & ~n66830 ;
  assign n66836 = ~n66834 & n66835 ;
  assign n66838 = ~\P2_P1_rEIP_reg[15]/NET0131  & ~n63462 ;
  assign n66839 = n25955 & ~n65499 ;
  assign n66840 = ~n66838 & n66839 ;
  assign n66837 = \P2_P1_Address_reg[13]/NET0131  & ~n25954 ;
  assign n66841 = ~\P2_P1_rEIP_reg[14]/NET0131  & ~n64804 ;
  assign n66842 = n63480 & ~n64050 ;
  assign n66843 = ~n66841 & n66842 ;
  assign n66844 = ~n66837 & ~n66843 ;
  assign n66845 = ~n66840 & n66844 ;
  assign n66847 = ~\P1_P1_rEIP_reg[15]/NET0131  & ~n63393 ;
  assign n66848 = n26155 & ~n64007 ;
  assign n66849 = ~n66847 & n66848 ;
  assign n66846 = \P1_P1_Address_reg[13]/NET0131  & ~n26154 ;
  assign n66850 = ~\P1_P1_rEIP_reg[14]/NET0131  & ~n63405 ;
  assign n66851 = n63401 & ~n63406 ;
  assign n66852 = ~n66850 & n66851 ;
  assign n66853 = ~n66846 & ~n66852 ;
  assign n66854 = ~n66849 & n66853 ;
  assign n66856 = ~\P2_P2_rEIP_reg[14]/NET0131  & ~n63990 ;
  assign n66857 = n63373 & ~n63991 ;
  assign n66858 = ~n66856 & n66857 ;
  assign n66855 = \P2_P2_Address_reg[13]/NET0131  & ~n26646 ;
  assign n66859 = ~\P2_P2_rEIP_reg[15]/NET0131  & ~n63998 ;
  assign n66860 = n26647 & ~n65439 ;
  assign n66861 = ~n66859 & n66860 ;
  assign n66862 = ~n66855 & ~n66861 ;
  assign n66863 = ~n66858 & n66862 ;
  assign n66865 = ~\P1_P3_rEIP_reg[15]/NET0131  & ~n64073 ;
  assign n66866 = n9092 & ~n64074 ;
  assign n66867 = ~n66865 & n66866 ;
  assign n66864 = \P1_P3_Address_reg[13]/NET0131  & ~n9091 ;
  assign n66868 = ~\P1_P3_rEIP_reg[14]/NET0131  & ~n64083 ;
  assign n66869 = n22115 & ~n64084 ;
  assign n66870 = ~n66868 & n66869 ;
  assign n66871 = ~n66864 & ~n66870 ;
  assign n66872 = ~n66867 & n66871 ;
  assign n66877 = ~\P1_P2_rEIP_reg[15]/NET0131  & ~n64845 ;
  assign n66878 = n25765 & ~n64033 ;
  assign n66879 = ~n66877 & n66878 ;
  assign n66873 = \P1_P2_Address_reg[13]/NET0131  & ~n25764 ;
  assign n66874 = ~\P1_P2_rEIP_reg[14]/NET0131  & ~n64851 ;
  assign n66875 = n63420 & ~n64024 ;
  assign n66876 = ~n66874 & n66875 ;
  assign n66880 = ~n66873 & ~n66876 ;
  assign n66881 = ~n66879 & n66880 ;
  assign n66883 = ~\P2_P3_rEIP_reg[15]/NET0131  & ~n64115 ;
  assign n66884 = n27145 & ~n64116 ;
  assign n66885 = ~n66883 & n66884 ;
  assign n66882 = \P2_P3_Address_reg[13]/NET0131  & ~n27144 ;
  assign n66886 = ~\P2_P3_rEIP_reg[14]/NET0131  & ~n64861 ;
  assign n66887 = n64094 & ~n66237 ;
  assign n66888 = ~n66886 & n66887 ;
  assign n66889 = ~n66882 & ~n66888 ;
  assign n66890 = ~n66885 & n66889 ;
  assign n66892 = ~\P2_P2_rEIP_reg[11]/NET0131  & ~n65264 ;
  assign n66893 = n26647 & ~n64821 ;
  assign n66894 = ~n66892 & n66893 ;
  assign n66891 = \P2_P2_Address_reg[9]/NET0131  & ~n26646 ;
  assign n66895 = ~\P2_P2_rEIP_reg[10]/NET0131  & ~n63988 ;
  assign n66896 = n63373 & ~n66383 ;
  assign n66897 = ~n66895 & n66896 ;
  assign n66898 = ~n66891 & ~n66897 ;
  assign n66899 = ~n66894 & n66898 ;
  assign n66905 = ~\P1_P3_rEIP_reg[11]/NET0131  & ~n64069 ;
  assign n66906 = n9092 & ~n64070 ;
  assign n66907 = ~n66905 & n66906 ;
  assign n66900 = \P1_P3_Address_reg[9]/NET0131  & ~n9091 ;
  assign n66902 = ~n17643 & n64081 ;
  assign n66901 = ~\P1_P3_rEIP_reg[10]/NET0131  & ~n64081 ;
  assign n66903 = n22115 & ~n66901 ;
  assign n66904 = ~n66902 & n66903 ;
  assign n66908 = ~n66900 & ~n66904 ;
  assign n66909 = ~n66907 & n66908 ;
  assign n66911 = ~\P1_P1_rEIP_reg[11]/NET0131  & ~n63390 ;
  assign n66912 = n26155 & ~n63391 ;
  assign n66913 = ~n66911 & n66912 ;
  assign n66910 = \P1_P1_Address_reg[9]/NET0131  & ~n26154 ;
  assign n66914 = ~\P1_P1_rEIP_reg[10]/NET0131  & ~n65290 ;
  assign n66915 = n63401 & ~n63403 ;
  assign n66916 = ~n66914 & n66915 ;
  assign n66917 = ~n66910 & ~n66916 ;
  assign n66918 = ~n66913 & n66917 ;
  assign n66924 = ~\P2_P3_rEIP_reg[11]/NET0131  & ~n64111 ;
  assign n66925 = n27145 & ~n64112 ;
  assign n66926 = ~n66924 & n66925 ;
  assign n66919 = \P2_P3_Address_reg[9]/NET0131  & ~n27144 ;
  assign n66921 = \P2_P3_rEIP_reg[10]/NET0131  & n65303 ;
  assign n66920 = ~\P2_P3_rEIP_reg[10]/NET0131  & ~n65303 ;
  assign n66922 = n64094 & ~n66920 ;
  assign n66923 = ~n66921 & n66922 ;
  assign n66927 = ~n66919 & ~n66923 ;
  assign n66928 = ~n66926 & n66927 ;
  assign n66933 = ~\P1_P2_rEIP_reg[11]/NET0131  & ~n64844 ;
  assign n66934 = n25765 & ~n64032 ;
  assign n66935 = ~n66933 & n66934 ;
  assign n66929 = \P1_P2_Address_reg[9]/NET0131  & ~n25764 ;
  assign n66930 = ~\P1_P2_rEIP_reg[10]/NET0131  & ~n65314 ;
  assign n66931 = n63420 & ~n64023 ;
  assign n66932 = ~n66930 & n66931 ;
  assign n66936 = ~n66929 & ~n66932 ;
  assign n66937 = ~n66935 & n66936 ;
  assign n66939 = ~\P2_P1_rEIP_reg[11]/NET0131  & ~n65320 ;
  assign n66940 = n25955 & ~n63461 ;
  assign n66941 = ~n66939 & n66940 ;
  assign n66938 = \P2_P1_Address_reg[9]/NET0131  & ~n25954 ;
  assign n66942 = ~\P2_P1_rEIP_reg[10]/NET0131  & ~n64048 ;
  assign n66943 = n63480 & ~n66422 ;
  assign n66944 = ~n66942 & n66943 ;
  assign n66945 = ~n66938 & ~n66944 ;
  assign n66946 = ~n66941 & n66945 ;
  assign n66952 = ~\P2_P1_rEIP_reg[23]/NET0131  & ~n65219 ;
  assign n66953 = n25955 & ~n63465 ;
  assign n66954 = ~n66952 & n66953 ;
  assign n66947 = \P2_P1_Address_reg[21]/NET0131  & ~n25954 ;
  assign n66949 = ~n50871 & n63475 ;
  assign n66948 = ~\P2_P1_rEIP_reg[22]/NET0131  & ~n63475 ;
  assign n66950 = n63480 & ~n66948 ;
  assign n66951 = ~n66949 & n66950 ;
  assign n66955 = ~n66947 & ~n66951 ;
  assign n66956 = ~n66954 & n66955 ;
  assign n66958 = ~\P2_P2_rEIP_reg[22]/NET0131  & ~n65228 ;
  assign n66959 = n63373 & ~n66300 ;
  assign n66960 = ~n66958 & n66959 ;
  assign n66957 = \P2_P2_Address_reg[21]/NET0131  & ~n26646 ;
  assign n66961 = ~\P2_P2_rEIP_reg[23]/NET0131  & ~n65232 ;
  assign n66962 = n26647 & ~n66296 ;
  assign n66963 = ~n66961 & n66962 ;
  assign n66964 = ~n66957 & ~n66963 ;
  assign n66965 = ~n66960 & n66964 ;
  assign n66971 = ~\P1_P2_rEIP_reg[23]/NET0131  & ~n66689 ;
  assign n66972 = n25765 & ~n66272 ;
  assign n66973 = ~n66971 & n66972 ;
  assign n66966 = \P1_P2_Address_reg[21]/NET0131  & ~n25764 ;
  assign n66967 = n51237 & n63421 ;
  assign n66968 = ~\P1_P2_rEIP_reg[22]/NET0131  & ~n66967 ;
  assign n66969 = n63420 & ~n66968 ;
  assign n66970 = ~n66683 & n66969 ;
  assign n66974 = ~n66966 & ~n66970 ;
  assign n66975 = ~n66973 & n66974 ;
  assign n66980 = ~\P1_P1_rEIP_reg[22]/NET0131  & ~n65246 ;
  assign n66981 = n63401 & ~n66307 ;
  assign n66982 = ~n66980 & n66981 ;
  assign n66976 = \P1_P1_Address_reg[21]/NET0131  & ~n26154 ;
  assign n66977 = ~\P1_P1_rEIP_reg[23]/NET0131  & ~n65241 ;
  assign n66978 = n26155 & ~n63394 ;
  assign n66979 = ~n66977 & n66978 ;
  assign n66983 = ~n66976 & ~n66979 ;
  assign n66984 = ~n66982 & n66983 ;
  assign n66985 = \P3_rd_reg/NET0131  & \P4_IR_reg[3]/NET0131  ;
  assign n66986 = \P2_P3_Datao_reg[3]/NET0131  & ~\P3_rd_reg/NET0131  ;
  assign n66987 = ~n66985 & ~n66986 ;
  assign n66988 = \P3_rd_reg/NET0131  & \P4_IR_reg[26]/NET0131  ;
  assign n66989 = \P2_P3_Datao_reg[26]/NET0131  & ~\P3_rd_reg/NET0131  ;
  assign n66990 = ~n66988 & ~n66989 ;
  assign n66996 = \P1_P2_State_reg[0]/NET0131  & \P1_P2_State_reg[1]/NET0131  ;
  assign n66997 = ~\P1_P2_State_reg[2]/NET0131  & n66996 ;
  assign n66998 = ~\P1_P2_RequestPending_reg/NET0131  & ~hold_pad ;
  assign n66999 = ~na_pad & n25415 ;
  assign n67000 = ~n66998 & n66999 ;
  assign n67001 = n66997 & n67000 ;
  assign n66991 = hold_pad & n66788 ;
  assign n66992 = ~\P1_P2_State_reg[1]/NET0131  & na_pad ;
  assign n66993 = ~\P1_P2_State_reg[0]/NET0131  & ~n66992 ;
  assign n66994 = ~n66742 & ~n66993 ;
  assign n66995 = \P1_P2_State_reg[2]/NET0131  & ~n66994 ;
  assign n67002 = ~n66991 & ~n66995 ;
  assign n67003 = ~n67001 & n67002 ;
  assign n67009 = \P2_P1_State_reg[0]/NET0131  & \P2_P1_State_reg[1]/NET0131  ;
  assign n67010 = ~\P2_P1_State_reg[2]/NET0131  & n67009 ;
  assign n67011 = ~\P2_P1_RequestPending_reg/NET0131  & ~hold_pad ;
  assign n67012 = ~na_pad & n21073 ;
  assign n67013 = ~n67011 & n67012 ;
  assign n67014 = n67010 & n67013 ;
  assign n67004 = hold_pad & n66800 ;
  assign n67005 = ~\P2_P1_State_reg[1]/NET0131  & na_pad ;
  assign n67006 = ~\P2_P1_State_reg[0]/NET0131  & ~n67005 ;
  assign n67007 = ~n66753 & ~n67006 ;
  assign n67008 = \P2_P1_State_reg[2]/NET0131  & ~n67007 ;
  assign n67015 = ~n67004 & ~n67008 ;
  assign n67016 = ~n67014 & n67015 ;
  assign n67017 = ~\P2_P2_RequestPending_reg/NET0131  & ~hold_pad ;
  assign n67018 = n26286 & ~n67017 ;
  assign n67019 = n66828 & n67018 ;
  assign n67020 = ~n26649 & ~n67019 ;
  assign n67021 = ~na_pad & ~n67020 ;
  assign n67025 = ~n66779 & n66824 ;
  assign n67022 = \P2_P2_RequestPending_reg/NET0131  & ~\P2_P2_State_reg[2]/NET0131  ;
  assign n67023 = hold_pad & n66825 ;
  assign n67024 = ~n67022 & n67023 ;
  assign n67026 = ~n63373 & ~n67024 ;
  assign n67027 = ~n67025 & n67026 ;
  assign n67028 = ~n67021 & n67027 ;
  assign n67035 = \P1_P1_State_reg[0]/NET0131  & \P1_P1_State_reg[1]/NET0131  ;
  assign n67036 = ~\P1_P1_State_reg[2]/NET0131  & n67035 ;
  assign n67037 = ~\P1_P1_RequestPending_reg/NET0131  & ~hold_pad ;
  assign n67038 = ~na_pad & n15335 ;
  assign n67039 = ~n67037 & n67038 ;
  assign n67040 = n67036 & n67039 ;
  assign n67029 = ~\P1_P1_State_reg[1]/NET0131  & na_pad ;
  assign n67030 = ~\P1_P1_State_reg[0]/NET0131  & ~n67029 ;
  assign n67031 = ~n66764 & ~n67030 ;
  assign n67032 = \P1_P1_State_reg[2]/NET0131  & ~n67031 ;
  assign n67033 = \P1_P1_State_reg[0]/NET0131  & hold_pad ;
  assign n67034 = ~n66818 & n67033 ;
  assign n67041 = ~n67032 & ~n67034 ;
  assign n67042 = ~n67040 & n67041 ;
  assign n67044 = ~\P2_P1_DataWidth_reg[0]/NET0131  & ~\P2_P1_DataWidth_reg[1]/NET0131  ;
  assign n67045 = \P2_P1_DataWidth_reg[0]/NET0131  & \P2_P1_DataWidth_reg[1]/NET0131  ;
  assign n67046 = \P2_P1_rEIP_reg[1]/NET0131  & ~n67045 ;
  assign n67047 = ~n67044 & ~n67046 ;
  assign n67048 = \P2_P1_rEIP_reg[0]/NET0131  & ~n67047 ;
  assign n67043 = ~\P2_P1_rEIP_reg[0]/NET0131  & n50417 ;
  assign n67049 = \P2_P1_ByteEnable_reg[2]/NET0131  & n67045 ;
  assign n67050 = ~n67043 & ~n67049 ;
  assign n67051 = ~n67048 & n67050 ;
  assign n67052 = \P2_P3_DataWidth_reg[0]/NET0131  & \P2_P3_DataWidth_reg[1]/NET0131  ;
  assign n67053 = \P2_P3_ByteEnable_reg[2]/NET0131  & n67052 ;
  assign n67054 = ~\P2_P3_DataWidth_reg[1]/NET0131  & \P2_P3_rEIP_reg[1]/NET0131  ;
  assign n67055 = \P2_P3_DataWidth_reg[0]/NET0131  & ~n67054 ;
  assign n67056 = \P2_P3_rEIP_reg[0]/NET0131  & ~n67055 ;
  assign n67057 = ~n64101 & ~n67056 ;
  assign n67058 = ~n56375 & ~n67057 ;
  assign n67059 = ~n67053 & ~n67058 ;
  assign n67061 = ~\P2_P2_DataWidth_reg[0]/NET0131  & ~\P2_P2_DataWidth_reg[1]/NET0131  ;
  assign n67062 = \P2_P2_DataWidth_reg[0]/NET0131  & \P2_P2_DataWidth_reg[1]/NET0131  ;
  assign n67063 = \P2_P2_rEIP_reg[1]/NET0131  & ~n67062 ;
  assign n67064 = ~n67061 & ~n67063 ;
  assign n67065 = \P2_P2_rEIP_reg[0]/NET0131  & ~n67064 ;
  assign n67060 = ~\P2_P2_rEIP_reg[0]/NET0131  & n50644 ;
  assign n67066 = \P2_P2_ByteEnable_reg[2]/NET0131  & n67062 ;
  assign n67067 = ~n67060 & ~n67066 ;
  assign n67068 = ~n67065 & n67067 ;
  assign n67072 = \P1_P3_DataWidth_reg[0]/NET0131  & \P1_P3_DataWidth_reg[1]/NET0131  ;
  assign n67074 = \P1_P3_rEIP_reg[1]/NET0131  & ~n67072 ;
  assign n67075 = ~\P1_P3_DataWidth_reg[0]/NET0131  & ~\P1_P3_DataWidth_reg[1]/NET0131  ;
  assign n67076 = \P1_P3_rEIP_reg[0]/NET0131  & ~n67075 ;
  assign n67077 = n67074 & n67076 ;
  assign n67069 = ~\P1_P3_DataWidth_reg[0]/NET0131  & \P1_P3_rEIP_reg[0]/NET0131  ;
  assign n67070 = ~n64059 & ~n67069 ;
  assign n67071 = ~\P1_P3_DataWidth_reg[1]/NET0131  & ~n67070 ;
  assign n67073 = \P1_P3_ByteEnable_reg[2]/NET0131  & n67072 ;
  assign n67078 = ~n67071 & ~n67073 ;
  assign n67079 = ~n67077 & n67078 ;
  assign n67081 = ~\P1_P2_DataWidth_reg[0]/NET0131  & ~\P1_P2_DataWidth_reg[1]/NET0131  ;
  assign n67082 = \P1_P2_DataWidth_reg[0]/NET0131  & \P1_P2_DataWidth_reg[1]/NET0131  ;
  assign n67083 = \P1_P2_rEIP_reg[1]/NET0131  & ~n67082 ;
  assign n67084 = ~n67081 & ~n67083 ;
  assign n67085 = \P1_P2_rEIP_reg[0]/NET0131  & ~n67084 ;
  assign n67080 = ~\P1_P2_rEIP_reg[0]/NET0131  & n50452 ;
  assign n67086 = \P1_P2_ByteEnable_reg[2]/NET0131  & n67082 ;
  assign n67087 = ~n67080 & ~n67086 ;
  assign n67088 = ~n67085 & n67087 ;
  assign n67089 = \P1_P1_DataWidth_reg[0]/NET0131  & \P1_P1_DataWidth_reg[1]/NET0131  ;
  assign n67091 = \P1_P1_rEIP_reg[1]/NET0131  & ~n67089 ;
  assign n67092 = \P1_P1_rEIP_reg[0]/NET0131  & n67091 ;
  assign n67090 = \P1_P1_ByteEnable_reg[2]/NET0131  & n67089 ;
  assign n67093 = \P1_P1_DataWidth_reg[0]/NET0131  & \P1_P1_rEIP_reg[0]/NET0131  ;
  assign n67094 = n50568 & ~n67093 ;
  assign n67095 = ~n67090 & ~n67094 ;
  assign n67096 = ~n67092 & n67095 ;
  assign n67099 = ~\P2_P3_DataWidth_reg[0]/NET0131  & ~\P2_P3_DataWidth_reg[1]/NET0131  ;
  assign n67100 = ~\P2_P3_rEIP_reg[0]/NET0131  & n67099 ;
  assign n67097 = \P2_P3_ByteEnable_reg[1]/NET0131  & n67052 ;
  assign n67098 = \P2_P3_rEIP_reg[1]/NET0131  & ~n67052 ;
  assign n67101 = ~n67097 & ~n67098 ;
  assign n67102 = ~n67100 & n67101 ;
  assign n67104 = ~\P1_P2_DataWidth_reg[0]/NET0131  & ~\P1_P2_rEIP_reg[0]/NET0131  ;
  assign n67105 = ~\P1_P2_DataWidth_reg[1]/NET0131  & n67104 ;
  assign n67103 = \P1_P2_ByteEnable_reg[1]/NET0131  & n67082 ;
  assign n67106 = ~n67083 & ~n67103 ;
  assign n67107 = ~n67105 & n67106 ;
  assign n67109 = ~\P2_P1_DataWidth_reg[0]/NET0131  & ~\P2_P1_rEIP_reg[0]/NET0131  ;
  assign n67110 = ~\P2_P1_DataWidth_reg[1]/NET0131  & n67109 ;
  assign n67108 = \P2_P1_ByteEnable_reg[1]/NET0131  & n67045 ;
  assign n67111 = ~n67046 & ~n67108 ;
  assign n67112 = ~n67110 & n67111 ;
  assign n67114 = \P1_P3_ByteEnable_reg[1]/NET0131  & n67072 ;
  assign n67113 = ~\P1_P3_rEIP_reg[0]/NET0131  & n67075 ;
  assign n67115 = ~n67074 & ~n67113 ;
  assign n67116 = ~n67114 & n67115 ;
  assign n67118 = ~\P1_P1_DataWidth_reg[0]/NET0131  & ~\P1_P1_rEIP_reg[0]/NET0131  ;
  assign n67119 = ~\P1_P1_DataWidth_reg[1]/NET0131  & n67118 ;
  assign n67117 = \P1_P1_ByteEnable_reg[1]/NET0131  & n67089 ;
  assign n67120 = ~n67091 & ~n67117 ;
  assign n67121 = ~n67119 & n67120 ;
  assign n67123 = ~\P2_P2_DataWidth_reg[0]/NET0131  & ~\P2_P2_rEIP_reg[0]/NET0131  ;
  assign n67124 = ~\P2_P2_DataWidth_reg[1]/NET0131  & n67123 ;
  assign n67122 = \P2_P2_ByteEnable_reg[1]/NET0131  & n67062 ;
  assign n67125 = ~n67063 & ~n67122 ;
  assign n67126 = ~n67124 & n67125 ;
  assign n67128 = ~\P1_P3_rEIP_reg[19]/NET0131  & ~n64078 ;
  assign n67129 = n9092 & ~n66542 ;
  assign n67130 = ~n67128 & n67129 ;
  assign n67127 = \P1_P3_Address_reg[17]/NET0131  & ~n9091 ;
  assign n67131 = ~\P1_P3_rEIP_reg[18]/NET0131  & ~n64087 ;
  assign n67132 = n22115 & ~n66537 ;
  assign n67133 = ~n67131 & n67132 ;
  assign n67134 = ~n67127 & ~n67133 ;
  assign n67135 = ~n67130 & n67134 ;
  assign n67141 = ~\P2_P3_rEIP_reg[19]/NET0131  & ~n64119 ;
  assign n67142 = n27145 & ~n66554 ;
  assign n67143 = ~n67141 & n67142 ;
  assign n67136 = \P2_P3_Address_reg[17]/NET0131  & ~n27144 ;
  assign n67138 = ~n54726 & n64095 ;
  assign n67137 = ~\P2_P3_rEIP_reg[18]/NET0131  & ~n64095 ;
  assign n67139 = n64094 & ~n67137 ;
  assign n67140 = ~n67138 & n67139 ;
  assign n67144 = ~n67136 & ~n67140 ;
  assign n67145 = ~n67143 & n67144 ;
  assign n67147 = ~\P2_P1_rEIP_reg[3]/NET0131  & ~n63453 ;
  assign n67148 = n25955 & ~n63454 ;
  assign n67149 = ~n67147 & n67148 ;
  assign n67146 = \P2_P1_Address_reg[1]/NET0131  & ~n25954 ;
  assign n67150 = ~\P2_P1_rEIP_reg[2]/NET0131  & ~n65406 ;
  assign n67151 = n63480 & ~n65407 ;
  assign n67152 = ~n67150 & n67151 ;
  assign n67153 = ~n67146 & ~n67152 ;
  assign n67154 = ~n67149 & n67153 ;
  assign n67156 = ~\P1_P1_rEIP_reg[3]/NET0131  & ~n63382 ;
  assign n67157 = n26155 & ~n63383 ;
  assign n67158 = ~n67156 & n67157 ;
  assign n67155 = \P1_P1_Address_reg[1]/NET0131  & ~n26154 ;
  assign n67159 = ~\P1_P1_rEIP_reg[2]/NET0131  & ~n65364 ;
  assign n67160 = n63401 & ~n65365 ;
  assign n67161 = ~n67159 & n67160 ;
  assign n67162 = ~n67155 & ~n67161 ;
  assign n67163 = ~n67158 & n67162 ;
  assign n67165 = ~\P2_P2_rEIP_reg[3]/NET0131  & ~n63352 ;
  assign n67166 = n26647 & ~n63353 ;
  assign n67167 = ~n67165 & n67166 ;
  assign n67164 = \P2_P2_Address_reg[1]/NET0131  & ~n26646 ;
  assign n67168 = ~\P2_P2_rEIP_reg[2]/NET0131  & ~n65336 ;
  assign n67169 = n63373 & ~n65337 ;
  assign n67170 = ~n67168 & n67169 ;
  assign n67171 = ~n67164 & ~n67170 ;
  assign n67172 = ~n67167 & n67171 ;
  assign n67174 = ~\P1_P3_rEIP_reg[3]/NET0131  & ~n64061 ;
  assign n67175 = n9092 & ~n64062 ;
  assign n67176 = ~n67174 & n67175 ;
  assign n67173 = \P1_P3_Address_reg[1]/NET0131  & ~n9091 ;
  assign n67177 = ~\P1_P3_rEIP_reg[2]/NET0131  & ~n65347 ;
  assign n67178 = n22115 & ~n65348 ;
  assign n67179 = ~n67177 & n67178 ;
  assign n67180 = ~n67173 & ~n67179 ;
  assign n67181 = ~n67176 & n67180 ;
  assign n67183 = ~\P2_P3_rEIP_reg[3]/NET0131  & ~n64103 ;
  assign n67184 = n27145 & ~n64104 ;
  assign n67185 = ~n67183 & n67184 ;
  assign n67182 = \P2_P3_Address_reg[1]/NET0131  & ~n27144 ;
  assign n67186 = ~\P2_P3_rEIP_reg[2]/NET0131  & ~n65378 ;
  assign n67187 = n64094 & ~n65379 ;
  assign n67188 = ~n67186 & n67187 ;
  assign n67189 = ~n67182 & ~n67188 ;
  assign n67190 = ~n67185 & n67189 ;
  assign n67192 = ~\P1_P2_rEIP_reg[3]/NET0131  & ~n63429 ;
  assign n67193 = n25765 & ~n63430 ;
  assign n67194 = ~n67192 & n67193 ;
  assign n67191 = \P1_P2_Address_reg[1]/NET0131  & ~n25764 ;
  assign n67195 = ~\P1_P2_rEIP_reg[2]/NET0131  & ~n65392 ;
  assign n67196 = n63420 & ~n65393 ;
  assign n67197 = ~n67195 & n67196 ;
  assign n67198 = ~n67191 & ~n67197 ;
  assign n67199 = ~n67194 & n67198 ;
  assign n67201 = ~\P2_P1_rEIP_reg[19]/NET0131  & ~n64042 ;
  assign n67202 = n25955 & ~n66526 ;
  assign n67203 = ~n67201 & n67202 ;
  assign n67200 = \P2_P1_Address_reg[17]/NET0131  & ~n25954 ;
  assign n67204 = ~\P2_P1_rEIP_reg[18]/NET0131  & ~n64053 ;
  assign n67205 = n63480 & ~n66530 ;
  assign n67206 = ~n67204 & n67205 ;
  assign n67207 = ~n67200 & ~n67206 ;
  assign n67208 = ~n67203 & n67207 ;
  assign n67213 = ~\P2_P2_rEIP_reg[19]/NET0131  & ~n64001 ;
  assign n67214 = n26647 & ~n65687 ;
  assign n67215 = ~n67213 & n67214 ;
  assign n67209 = \P2_P2_Address_reg[17]/NET0131  & ~n26646 ;
  assign n67210 = ~\P2_P2_rEIP_reg[18]/NET0131  & ~n63995 ;
  assign n67211 = n63373 & ~n66497 ;
  assign n67212 = ~n67210 & n67211 ;
  assign n67216 = ~n67209 & ~n67212 ;
  assign n67217 = ~n67215 & n67216 ;
  assign n67222 = ~\P1_P1_rEIP_reg[19]/NET0131  & ~n64011 ;
  assign n67223 = n26155 & ~n65699 ;
  assign n67224 = ~n67222 & n67223 ;
  assign n67218 = \P1_P1_Address_reg[17]/NET0131  & ~n26154 ;
  assign n67219 = ~\P1_P1_rEIP_reg[18]/NET0131  & ~n64015 ;
  assign n67220 = n63401 & ~n66504 ;
  assign n67221 = ~n67219 & n67220 ;
  assign n67225 = ~n67218 & ~n67221 ;
  assign n67226 = ~n67224 & n67225 ;
  assign n67231 = ~\P1_P2_rEIP_reg[18]/NET0131  & ~n64028 ;
  assign n67232 = n63420 & ~n65252 ;
  assign n67233 = ~n67231 & n67232 ;
  assign n67227 = \P1_P2_Address_reg[17]/NET0131  & ~n25764 ;
  assign n67228 = ~\P1_P2_rEIP_reg[19]/NET0131  & ~n66517 ;
  assign n67229 = n25765 & ~n66518 ;
  assign n67230 = ~n67228 & n67229 ;
  assign n67234 = ~n67227 & ~n67230 ;
  assign n67235 = ~n67233 & n67234 ;
  assign n67237 = ~\P2_P2_rEIP_reg[7]/NET0131  & ~n63356 ;
  assign n67238 = n26647 & ~n63357 ;
  assign n67239 = ~n67237 & n67238 ;
  assign n67236 = \P2_P2_Address_reg[5]/NET0131  & ~n26646 ;
  assign n67240 = ~\P2_P2_rEIP_reg[6]/NET0131  & ~n65340 ;
  assign n67241 = n63373 & ~n63985 ;
  assign n67242 = ~n67240 & n67241 ;
  assign n67243 = ~n67236 & ~n67242 ;
  assign n67244 = ~n67239 & n67243 ;
  assign n67250 = ~\P1_P3_rEIP_reg[7]/NET0131  & ~n64065 ;
  assign n67251 = n9092 & ~n64066 ;
  assign n67252 = ~n67250 & n67251 ;
  assign n67245 = \P1_P3_Address_reg[5]/NET0131  & ~n9091 ;
  assign n67247 = ~n17583 & n64081 ;
  assign n67246 = ~\P1_P3_rEIP_reg[6]/NET0131  & ~n64081 ;
  assign n67248 = n22115 & ~n67246 ;
  assign n67249 = ~n67247 & n67248 ;
  assign n67253 = ~n67245 & ~n67249 ;
  assign n67254 = ~n67252 & n67253 ;
  assign n67256 = ~\P1_P1_rEIP_reg[7]/NET0131  & ~n63386 ;
  assign n67257 = n26155 & ~n63387 ;
  assign n67258 = ~n67256 & n67257 ;
  assign n67255 = \P1_P1_Address_reg[5]/NET0131  & ~n26154 ;
  assign n67259 = ~\P1_P1_rEIP_reg[6]/NET0131  & ~n65368 ;
  assign n67260 = n63401 & ~n65287 ;
  assign n67261 = ~n67259 & n67260 ;
  assign n67262 = ~n67255 & ~n67261 ;
  assign n67263 = ~n67258 & n67262 ;
  assign n67265 = ~\P2_P3_rEIP_reg[7]/NET0131  & ~n64107 ;
  assign n67266 = n27145 & ~n64108 ;
  assign n67267 = ~n67265 & n67266 ;
  assign n67264 = \P2_P3_Address_reg[5]/NET0131  & ~n27144 ;
  assign n67268 = ~\P2_P3_rEIP_reg[6]/NET0131  & ~n65382 ;
  assign n67269 = n64094 & ~n65300 ;
  assign n67270 = ~n67268 & n67269 ;
  assign n67271 = ~n67264 & ~n67270 ;
  assign n67272 = ~n67267 & n67271 ;
  assign n67274 = ~\P1_P2_rEIP_reg[7]/NET0131  & ~n63433 ;
  assign n67275 = n25765 & ~n63434 ;
  assign n67276 = ~n67274 & n67275 ;
  assign n67273 = \P1_P2_Address_reg[5]/NET0131  & ~n25764 ;
  assign n67277 = ~\P1_P2_rEIP_reg[6]/NET0131  & ~n65397 ;
  assign n67278 = n63420 & ~n66601 ;
  assign n67279 = ~n67277 & n67278 ;
  assign n67280 = ~n67273 & ~n67279 ;
  assign n67281 = ~n67276 & n67280 ;
  assign n67283 = ~\P2_P1_rEIP_reg[7]/NET0131  & ~n63457 ;
  assign n67284 = n25955 & ~n63458 ;
  assign n67285 = ~n67283 & n67284 ;
  assign n67282 = \P2_P1_Address_reg[5]/NET0131  & ~n25954 ;
  assign n67286 = ~\P2_P1_rEIP_reg[6]/NET0131  & ~n65410 ;
  assign n67287 = n63480 & ~n64045 ;
  assign n67288 = ~n67286 & n67287 ;
  assign n67289 = ~n67282 & ~n67288 ;
  assign n67290 = ~n67285 & n67289 ;
  assign n67291 = \P3_rd_reg/NET0131  & \P4_IR_reg[29]/NET0131  ;
  assign n67292 = \P2_P3_Datao_reg[29]/NET0131  & ~\P3_rd_reg/NET0131  ;
  assign n67293 = ~n67291 & ~n67292 ;
  assign n67294 = \P3_rd_reg/NET0131  & \P4_IR_reg[18]/NET0131  ;
  assign n67295 = \P2_P3_Datao_reg[18]/NET0131  & ~\P3_rd_reg/NET0131  ;
  assign n67296 = ~n67294 & ~n67295 ;
  assign n67297 = \P3_rd_reg/NET0131  & \P4_IR_reg[14]/NET0131  ;
  assign n67298 = \P2_P3_Datao_reg[14]/NET0131  & ~\P3_rd_reg/NET0131  ;
  assign n67299 = ~n67297 & ~n67298 ;
  assign n67300 = \P3_rd_reg/NET0131  & \P4_IR_reg[22]/NET0131  ;
  assign n67301 = \P2_P3_Datao_reg[22]/NET0131  & ~\P3_rd_reg/NET0131  ;
  assign n67302 = ~n67300 & ~n67301 ;
  assign n67303 = \P2_P1_ByteEnable_reg[3]/NET0131  & n67045 ;
  assign n67304 = \P2_P1_rEIP_reg[1]/NET0131  & ~n67109 ;
  assign n67305 = ~\P2_P1_DataWidth_reg[1]/NET0131  & ~n67304 ;
  assign n67306 = ~n67303 & ~n67305 ;
  assign n67307 = \P2_P2_ByteEnable_reg[3]/NET0131  & n67062 ;
  assign n67308 = \P2_P2_rEIP_reg[1]/NET0131  & ~n67123 ;
  assign n67309 = ~\P2_P2_DataWidth_reg[1]/NET0131  & ~n67308 ;
  assign n67310 = ~n67307 & ~n67309 ;
  assign n67311 = \P1_P3_ByteEnable_reg[3]/NET0131  & n67072 ;
  assign n67312 = \P1_P3_rEIP_reg[1]/NET0131  & ~n67113 ;
  assign n67313 = ~\P1_P3_DataWidth_reg[1]/NET0131  & ~n67312 ;
  assign n67314 = ~n67311 & ~n67313 ;
  assign n67315 = \P1_P2_ByteEnable_reg[3]/NET0131  & n67082 ;
  assign n67316 = \P1_P2_rEIP_reg[1]/NET0131  & ~n67104 ;
  assign n67317 = ~\P1_P2_DataWidth_reg[1]/NET0131  & ~n67316 ;
  assign n67318 = ~n67315 & ~n67317 ;
  assign n67319 = \P2_P3_ByteEnable_reg[3]/NET0131  & n67052 ;
  assign n67320 = \P2_P3_rEIP_reg[1]/NET0131  & ~n67100 ;
  assign n67321 = ~\P2_P3_DataWidth_reg[1]/NET0131  & ~n67320 ;
  assign n67322 = ~n67319 & ~n67321 ;
  assign n67323 = \P1_P1_ByteEnable_reg[3]/NET0131  & n67089 ;
  assign n67324 = \P1_P1_rEIP_reg[1]/NET0131  & ~n67118 ;
  assign n67325 = ~\P1_P1_DataWidth_reg[1]/NET0131  & ~n67324 ;
  assign n67326 = ~n67323 & ~n67325 ;
  assign n67327 = \P3_rd_reg/NET0131  & \P4_IR_reg[25]/NET0131  ;
  assign n67328 = \P2_P3_Datao_reg[25]/NET0131  & ~\P3_rd_reg/NET0131  ;
  assign n67329 = ~n67327 & ~n67328 ;
  assign n67330 = \P3_rd_reg/NET0131  & \P4_IR_reg[10]/NET0131  ;
  assign n67331 = \P2_P3_Datao_reg[10]/NET0131  & ~\P3_rd_reg/NET0131  ;
  assign n67332 = ~n67330 & ~n67331 ;
  assign n67333 = \P3_rd_reg/NET0131  & \P4_IR_reg[6]/NET0131  ;
  assign n67334 = \P2_P3_Datao_reg[6]/NET0131  & ~\P3_rd_reg/NET0131  ;
  assign n67335 = ~n67333 & ~n67334 ;
  assign n67336 = \P3_rd_reg/NET0131  & \P4_IR_reg[2]/NET0131  ;
  assign n67337 = \P2_P3_Datao_reg[2]/NET0131  & ~\P3_rd_reg/NET0131  ;
  assign n67338 = ~n67336 & ~n67337 ;
  assign n67339 = \P3_rd_reg/NET0131  & \P4_IR_reg[17]/NET0131  ;
  assign n67340 = \P2_P3_Datao_reg[17]/NET0131  & ~\P3_rd_reg/NET0131  ;
  assign n67341 = ~n67339 & ~n67340 ;
  assign n67342 = \P3_rd_reg/NET0131  & \P4_IR_reg[21]/NET0131  ;
  assign n67343 = \P2_P3_Datao_reg[21]/NET0131  & ~\P3_rd_reg/NET0131  ;
  assign n67344 = ~n67342 & ~n67343 ;
  assign n67346 = ~\P2_P1_rEIP_reg[2]/NET0131  & ~n63452 ;
  assign n67347 = n25955 & ~n63453 ;
  assign n67348 = ~n67346 & n67347 ;
  assign n67345 = \P2_P1_Address_reg[0]/NET0131  & ~n25954 ;
  assign n67349 = ~\P2_P1_rEIP_reg[1]/NET0131  & ~n63475 ;
  assign n67350 = n63480 & ~n65406 ;
  assign n67351 = ~n67349 & n67350 ;
  assign n67352 = ~n67345 & ~n67351 ;
  assign n67353 = ~n67348 & n67352 ;
  assign n67355 = ~\P1_P2_rEIP_reg[2]/NET0131  & ~n63428 ;
  assign n67356 = n25765 & ~n63429 ;
  assign n67357 = ~n67355 & n67356 ;
  assign n67354 = \P1_P2_Address_reg[0]/NET0131  & ~n25764 ;
  assign n67358 = ~\P1_P2_rEIP_reg[1]/NET0131  & ~n63421 ;
  assign n67359 = n63420 & ~n65392 ;
  assign n67360 = ~n67358 & n67359 ;
  assign n67361 = ~n67354 & ~n67360 ;
  assign n67362 = ~n67357 & n67361 ;
  assign n67364 = ~\P1_P1_rEIP_reg[2]/NET0131  & ~n63381 ;
  assign n67365 = n26155 & ~n63382 ;
  assign n67366 = ~n67364 & n67365 ;
  assign n67363 = \P1_P1_Address_reg[0]/NET0131  & ~n26154 ;
  assign n67367 = ~\P1_P1_rEIP_reg[1]/NET0131  & ~n63402 ;
  assign n67368 = n63401 & ~n65364 ;
  assign n67369 = ~n67367 & n67368 ;
  assign n67370 = ~n67363 & ~n67369 ;
  assign n67371 = ~n67366 & n67370 ;
  assign n67373 = ~\P1_P3_rEIP_reg[2]/NET0131  & ~n64060 ;
  assign n67374 = n9092 & ~n64061 ;
  assign n67375 = ~n67373 & n67374 ;
  assign n67372 = \P1_P3_Address_reg[0]/NET0131  & ~n9091 ;
  assign n67376 = ~\P1_P3_rEIP_reg[1]/NET0131  & ~n64081 ;
  assign n67377 = n22115 & ~n65347 ;
  assign n67378 = ~n67376 & n67377 ;
  assign n67379 = ~n67372 & ~n67378 ;
  assign n67380 = ~n67375 & n67379 ;
  assign n67382 = ~\P2_P2_rEIP_reg[2]/NET0131  & ~n63351 ;
  assign n67383 = n26647 & ~n63352 ;
  assign n67384 = ~n67382 & n67383 ;
  assign n67381 = \P2_P2_Address_reg[0]/NET0131  & ~n26646 ;
  assign n67385 = ~\P2_P2_rEIP_reg[1]/NET0131  & ~n63368 ;
  assign n67386 = n63373 & ~n65336 ;
  assign n67387 = ~n67385 & n67386 ;
  assign n67388 = ~n67381 & ~n67387 ;
  assign n67389 = ~n67384 & n67388 ;
  assign n67391 = ~\P2_P3_rEIP_reg[2]/NET0131  & ~n64102 ;
  assign n67392 = n27145 & ~n64103 ;
  assign n67393 = ~n67391 & n67392 ;
  assign n67390 = \P2_P3_Address_reg[0]/NET0131  & ~n27144 ;
  assign n67394 = ~\P2_P3_rEIP_reg[1]/NET0131  & ~n64095 ;
  assign n67395 = n64094 & ~n65378 ;
  assign n67396 = ~n67394 & n67395 ;
  assign n67397 = ~n67390 & ~n67396 ;
  assign n67398 = ~n67393 & n67397 ;
  assign n67399 = \P3_rd_reg/NET0131  & \P4_IR_reg[13]/NET0131  ;
  assign n67400 = \P2_P3_Datao_reg[13]/NET0131  & ~\P3_rd_reg/NET0131  ;
  assign n67401 = ~n67399 & ~n67400 ;
  assign n67402 = \P3_rd_reg/NET0131  & \P4_IR_reg[5]/NET0131  ;
  assign n67403 = \P2_P3_Datao_reg[5]/NET0131  & ~\P3_rd_reg/NET0131  ;
  assign n67404 = ~n67402 & ~n67403 ;
  assign n67405 = \P3_rd_reg/NET0131  & \P4_IR_reg[9]/NET0131  ;
  assign n67406 = \P2_P3_Datao_reg[9]/NET0131  & ~\P3_rd_reg/NET0131  ;
  assign n67407 = ~n67405 & ~n67406 ;
  assign n67408 = ~n26156 & ~n67036 ;
  assign n67409 = ~\P1_P1_DataWidth_reg[1]/NET0131  & n67408 ;
  assign n67410 = ~n26157 & ~n67036 ;
  assign n67411 = ~bs_pad & ~n67410 ;
  assign n67412 = ~n67409 & ~n67411 ;
  assign n67415 = ~n26646 & n66826 ;
  assign n67416 = \P2_P2_DataWidth_reg[1]/NET0131  & ~n67415 ;
  assign n67413 = ~n26649 & ~n66828 ;
  assign n67414 = bs_pad & ~n67413 ;
  assign n67417 = ~\P2_P2_State_reg[2]/NET0131  & n26648 ;
  assign n67418 = ~n67414 & ~n67417 ;
  assign n67419 = ~n67416 & n67418 ;
  assign n67420 = ~n9093 & ~n23019 ;
  assign n67421 = ~\P1_P3_DataWidth_reg[1]/NET0131  & n67420 ;
  assign n67422 = ~n9094 & ~n23019 ;
  assign n67423 = ~bs_pad & ~n67422 ;
  assign n67424 = ~n67421 & ~n67423 ;
  assign n67425 = ~n25766 & ~n66997 ;
  assign n67426 = ~\P1_P2_DataWidth_reg[1]/NET0131  & n67425 ;
  assign n67427 = ~n25767 & ~n66997 ;
  assign n67428 = ~bs_pad & ~n67427 ;
  assign n67429 = ~n67426 & ~n67428 ;
  assign n67430 = ~n27146 & ~n66359 ;
  assign n67431 = ~\P2_P3_DataWidth_reg[1]/NET0131  & n67430 ;
  assign n67432 = ~n27147 & ~n66359 ;
  assign n67433 = ~bs_pad & ~n67432 ;
  assign n67434 = ~n67431 & ~n67433 ;
  assign n67435 = ~n25956 & ~n67010 ;
  assign n67436 = ~\P2_P1_DataWidth_reg[1]/NET0131  & n67435 ;
  assign n67437 = ~n25957 & ~n67010 ;
  assign n67438 = ~bs_pad & ~n67437 ;
  assign n67439 = ~n67436 & ~n67438 ;
  assign n67440 = \P2_P1_DataWidth_reg[0]/NET0131  & n67435 ;
  assign n67441 = ~n67438 & ~n67440 ;
  assign n67442 = \P2_P1_BE_n_reg[1]/NET0131  & ~n25954 ;
  assign n67443 = \P2_P1_ByteEnable_reg[1]/NET0131  & n25954 ;
  assign n67444 = ~n67442 & ~n67443 ;
  assign n67445 = \P2_P1_ADS_n_reg/NET0131  & \P2_P1_State_reg[0]/NET0131  ;
  assign n67446 = n67435 & ~n67445 ;
  assign n67447 = \P1_P2_DataWidth_reg[0]/NET0131  & n67425 ;
  assign n67448 = ~n67428 & ~n67447 ;
  assign n67449 = \P1_P1_DataWidth_reg[0]/NET0131  & n67408 ;
  assign n67450 = ~n67411 & ~n67449 ;
  assign n67451 = \P2_P2_W_R_n_reg/NET0131  & ~n26646 ;
  assign n67452 = ~\P2_P2_ReadRequest_reg/NET0131  & n26646 ;
  assign n67453 = ~n67451 & ~n67452 ;
  assign n67454 = \P1_P3_DataWidth_reg[0]/NET0131  & n67420 ;
  assign n67455 = ~n67423 & ~n67454 ;
  assign n67456 = \P1_P2_M_IO_n_reg/NET0131  & ~n25764 ;
  assign n67457 = \P1_P2_MemoryFetch_reg/NET0131  & n25764 ;
  assign n67458 = ~n67456 & ~n67457 ;
  assign n67459 = \P2_P3_ADS_n_reg/NET0131  & \P2_P3_State_reg[0]/NET0131  ;
  assign n67460 = n67430 & ~n67459 ;
  assign n67461 = \P1_P1_ADS_n_reg/NET0131  & \P1_P1_State_reg[0]/NET0131  ;
  assign n67462 = n67408 & ~n67461 ;
  assign n67463 = \P2_P3_BE_n_reg[2]/NET0131  & ~n27144 ;
  assign n67464 = \P2_P3_ByteEnable_reg[2]/NET0131  & n27144 ;
  assign n67465 = ~n67463 & ~n67464 ;
  assign n67466 = \P2_P1_M_IO_n_reg/NET0131  & ~n25954 ;
  assign n67467 = \P2_P1_MemoryFetch_reg/NET0131  & n25954 ;
  assign n67468 = ~n67466 & ~n67467 ;
  assign n67469 = \P2_P3_BE_n_reg[1]/NET0131  & ~n27144 ;
  assign n67470 = \P2_P3_ByteEnable_reg[1]/NET0131  & n27144 ;
  assign n67471 = ~n67469 & ~n67470 ;
  assign n67472 = \P1_P2_W_R_n_reg/NET0131  & ~n25764 ;
  assign n67473 = ~\P1_P2_ReadRequest_reg/NET0131  & n25764 ;
  assign n67474 = ~n67472 & ~n67473 ;
  assign n67475 = \P2_P3_BE_n_reg[0]/NET0131  & ~n27144 ;
  assign n67476 = \P2_P3_ByteEnable_reg[0]/NET0131  & n27144 ;
  assign n67477 = ~n67475 & ~n67476 ;
  assign n67478 = \P2_P1_BE_n_reg[3]/NET0131  & ~n25954 ;
  assign n67479 = \P2_P1_ByteEnable_reg[3]/NET0131  & n25954 ;
  assign n67480 = ~n67478 & ~n67479 ;
  assign n67481 = \P1_P1_M_IO_n_reg/NET0131  & ~n26154 ;
  assign n67482 = \P1_P1_MemoryFetch_reg/NET0131  & n26154 ;
  assign n67483 = ~n67481 & ~n67482 ;
  assign n67484 = \P2_P2_BE_n_reg[0]/NET0131  & ~n26646 ;
  assign n67485 = \P2_P2_ByteEnable_reg[0]/NET0131  & n26646 ;
  assign n67486 = ~n67484 & ~n67485 ;
  assign n67487 = \P2_P2_BE_n_reg[1]/NET0131  & ~n26646 ;
  assign n67488 = \P2_P2_ByteEnable_reg[1]/NET0131  & n26646 ;
  assign n67489 = ~n67487 & ~n67488 ;
  assign n67490 = \P2_P2_BE_n_reg[2]/NET0131  & ~n26646 ;
  assign n67491 = \P2_P2_ByteEnable_reg[2]/NET0131  & n26646 ;
  assign n67492 = ~n67490 & ~n67491 ;
  assign n67493 = \P2_P2_BE_n_reg[3]/NET0131  & ~n26646 ;
  assign n67494 = \P2_P2_ByteEnable_reg[3]/NET0131  & n26646 ;
  assign n67495 = ~n67493 & ~n67494 ;
  assign n67496 = ~bs_pad & ~n67413 ;
  assign n67497 = \P2_P2_DataWidth_reg[0]/NET0131  & ~n67415 ;
  assign n67498 = ~n67496 & ~n67497 ;
  assign n67499 = \P1_P3_ADS_n_reg/NET0131  & \P1_P3_State_reg[0]/NET0131  ;
  assign n67500 = n67420 & ~n67499 ;
  assign n67501 = \P1_P3_BE_n_reg[0]/NET0131  & ~n9091 ;
  assign n67502 = \P1_P3_ByteEnable_reg[0]/NET0131  & n9091 ;
  assign n67503 = ~n67501 & ~n67502 ;
  assign n67504 = \P1_P3_BE_n_reg[1]/NET0131  & ~n9091 ;
  assign n67505 = \P1_P3_ByteEnable_reg[1]/NET0131  & n9091 ;
  assign n67506 = ~n67504 & ~n67505 ;
  assign n67507 = \P2_P3_DataWidth_reg[0]/NET0131  & n67430 ;
  assign n67508 = ~n67433 & ~n67507 ;
  assign n67509 = \P1_P1_W_R_n_reg/NET0131  & ~n26154 ;
  assign n67510 = ~\P1_P1_ReadRequest_reg/NET0131  & n26154 ;
  assign n67511 = ~n67509 & ~n67510 ;
  assign n67512 = \P2_P1_BE_n_reg[2]/NET0131  & ~n25954 ;
  assign n67513 = \P2_P1_ByteEnable_reg[2]/NET0131  & n25954 ;
  assign n67514 = ~n67512 & ~n67513 ;
  assign n67515 = \P1_P3_BE_n_reg[3]/NET0131  & ~n9091 ;
  assign n67516 = \P1_P3_ByteEnable_reg[3]/NET0131  & n9091 ;
  assign n67517 = ~n67515 & ~n67516 ;
  assign n67518 = \P1_P2_ADS_n_reg/NET0131  & \P1_P2_State_reg[0]/NET0131  ;
  assign n67519 = n67425 & ~n67518 ;
  assign n67520 = \P1_P1_BE_n_reg[0]/NET0131  & ~n26154 ;
  assign n67521 = \P1_P1_ByteEnable_reg[0]/NET0131  & n26154 ;
  assign n67522 = ~n67520 & ~n67521 ;
  assign n67523 = \P1_P1_BE_n_reg[3]/NET0131  & ~n26154 ;
  assign n67524 = \P1_P1_ByteEnable_reg[3]/NET0131  & n26154 ;
  assign n67525 = ~n67523 & ~n67524 ;
  assign n67526 = \P2_P3_BE_n_reg[3]/NET0131  & ~n27144 ;
  assign n67527 = \P2_P3_ByteEnable_reg[3]/NET0131  & n27144 ;
  assign n67528 = ~n67526 & ~n67527 ;
  assign n67529 = \P1_P2_BE_n_reg[0]/NET0131  & ~n25764 ;
  assign n67530 = \P1_P2_ByteEnable_reg[0]/NET0131  & n25764 ;
  assign n67531 = ~n67529 & ~n67530 ;
  assign n67532 = \P1_P2_BE_n_reg[1]/NET0131  & ~n25764 ;
  assign n67533 = \P1_P2_ByteEnable_reg[1]/NET0131  & n25764 ;
  assign n67534 = ~n67532 & ~n67533 ;
  assign n67535 = \P1_P2_BE_n_reg[2]/NET0131  & ~n25764 ;
  assign n67536 = \P1_P2_ByteEnable_reg[2]/NET0131  & n25764 ;
  assign n67537 = ~n67535 & ~n67536 ;
  assign n67538 = \P1_P2_BE_n_reg[3]/NET0131  & ~n25764 ;
  assign n67539 = \P1_P2_ByteEnable_reg[3]/NET0131  & n25764 ;
  assign n67540 = ~n67538 & ~n67539 ;
  assign n67541 = \P2_P2_M_IO_n_reg/NET0131  & ~n26646 ;
  assign n67542 = \P2_P2_MemoryFetch_reg/NET0131  & n26646 ;
  assign n67543 = ~n67541 & ~n67542 ;
  assign n67544 = \P1_P1_BE_n_reg[1]/NET0131  & ~n26154 ;
  assign n67545 = \P1_P1_ByteEnable_reg[1]/NET0131  & n26154 ;
  assign n67546 = ~n67544 & ~n67545 ;
  assign n67547 = \P2_P2_ADS_n_reg/NET0131  & \P2_P2_State_reg[0]/NET0131  ;
  assign n67548 = ~n26648 & ~n67547 ;
  assign n67549 = ~n66828 & n67548 ;
  assign n67550 = \P2_P1_W_R_n_reg/NET0131  & ~n25954 ;
  assign n67551 = ~\P2_P1_ReadRequest_reg/NET0131  & n25954 ;
  assign n67552 = ~n67550 & ~n67551 ;
  assign n67553 = \P2_P3_M_IO_n_reg/NET0131  & ~n27144 ;
  assign n67554 = \P2_P3_MemoryFetch_reg/NET0131  & n27144 ;
  assign n67555 = ~n67553 & ~n67554 ;
  assign n67556 = \P2_P3_W_R_n_reg/NET0131  & ~n27144 ;
  assign n67557 = ~\P2_P3_ReadRequest_reg/NET0131  & n27144 ;
  assign n67558 = ~n67556 & ~n67557 ;
  assign n67559 = \P1_P3_M_IO_n_reg/NET0131  & ~n9091 ;
  assign n67560 = \P1_P3_MemoryFetch_reg/NET0131  & n9091 ;
  assign n67561 = ~n67559 & ~n67560 ;
  assign n67562 = \P2_P1_BE_n_reg[0]/NET0131  & ~n25954 ;
  assign n67563 = \P2_P1_ByteEnable_reg[0]/NET0131  & n25954 ;
  assign n67564 = ~n67562 & ~n67563 ;
  assign n67565 = \P1_P1_BE_n_reg[2]/NET0131  & ~n26154 ;
  assign n67566 = \P1_P1_ByteEnable_reg[2]/NET0131  & n26154 ;
  assign n67567 = ~n67565 & ~n67566 ;
  assign n67568 = \P1_P3_BE_n_reg[2]/NET0131  & ~n9091 ;
  assign n67569 = \P1_P3_ByteEnable_reg[2]/NET0131  & n9091 ;
  assign n67570 = ~n67568 & ~n67569 ;
  assign n67571 = \P1_P3_W_R_n_reg/NET0131  & ~n9091 ;
  assign n67572 = ~\P1_P3_ReadRequest_reg/NET0131  & n9091 ;
  assign n67573 = ~n67571 & ~n67572 ;
  assign n67575 = n66826 & n67413 ;
  assign n67576 = \P2_P2_D_C_n_reg/NET0131  & ~n67575 ;
  assign n67574 = ~\P2_P2_CodeFetch_reg/NET0131  & n26646 ;
  assign n67577 = ~n67417 & ~n67574 ;
  assign n67578 = ~n67576 & n67577 ;
  assign n67579 = ~\P2_P1_State_reg[1]/NET0131  & \P2_P1_State_reg[2]/NET0131  ;
  assign n67580 = ~\P2_P1_State_reg[0]/NET0131  & ~n67579 ;
  assign n67581 = ~\P2_P1_D_C_n_reg/NET0131  & ~n67580 ;
  assign n67582 = \P2_P1_CodeFetch_reg/NET0131  & n25954 ;
  assign n67583 = ~n67581 & ~n67582 ;
  assign n67584 = ~\P1_P1_D_C_n_reg/NET0131  & ~n66816 ;
  assign n67585 = \P1_P1_CodeFetch_reg/NET0131  & n26154 ;
  assign n67586 = ~n67584 & ~n67585 ;
  assign n67587 = ~\P1_P3_State_reg[1]/NET0131  & \P1_P3_State_reg[2]/NET0131  ;
  assign n67588 = ~\P1_P3_State_reg[0]/NET0131  & ~n67587 ;
  assign n67589 = ~\P1_P3_D_C_n_reg/NET0131  & ~n67588 ;
  assign n67590 = \P1_P3_CodeFetch_reg/NET0131  & n9091 ;
  assign n67591 = ~n67589 & ~n67590 ;
  assign n67592 = ~\P1_P2_State_reg[1]/NET0131  & \P1_P2_State_reg[2]/NET0131  ;
  assign n67593 = ~\P1_P2_State_reg[0]/NET0131  & ~n67592 ;
  assign n67594 = ~\P1_P2_D_C_n_reg/NET0131  & ~n67593 ;
  assign n67595 = \P1_P2_CodeFetch_reg/NET0131  & n25764 ;
  assign n67596 = ~n67594 & ~n67595 ;
  assign n67598 = n66357 & n67432 ;
  assign n67599 = \P2_P3_D_C_n_reg/NET0131  & ~n67598 ;
  assign n67597 = ~\P2_P3_CodeFetch_reg/NET0131  & n27144 ;
  assign n67600 = ~\P2_P3_State_reg[2]/NET0131  & n27146 ;
  assign n67601 = ~n67597 & ~n67600 ;
  assign n67602 = ~n67599 & n67601 ;
  assign n67603 = \P3_rd_reg/NET0131  & \P4_IR_reg[1]/NET0131  ;
  assign n67604 = \P2_P3_Datao_reg[1]/NET0131  & ~\P3_rd_reg/NET0131  ;
  assign n67605 = ~n67603 & ~n67604 ;
  assign n67606 = \P4_reg2_reg[28]/NET0131  & ~n20673 ;
  assign n67613 = n18747 & n23843 ;
  assign n67614 = ~n67606 & ~n67613 ;
  assign n67615 = n18483 & ~n67614 ;
  assign n67608 = ~n18740 & n20673 ;
  assign n67607 = ~n22000 & n67606 ;
  assign n67609 = n15790 & n16426 ;
  assign n67610 = ~n67607 & ~n67609 ;
  assign n67611 = ~n67608 & n67610 ;
  assign n67612 = n18666 & ~n67611 ;
  assign n67616 = ~n20681 & n22172 ;
  assign n67617 = \P4_reg2_reg[28]/NET0131  & ~n67616 ;
  assign n67618 = ~n67612 & ~n67617 ;
  assign n67619 = ~n67615 & n67618 ;
  assign n67630 = n11599 & ~n12820 ;
  assign n67625 = n11383 & ~n11920 ;
  assign n67621 = \P2_P1_InstQueue_reg[12][6]/NET0131  & ~n11919 ;
  assign n67626 = ~n11596 & n67621 ;
  assign n67627 = ~n67625 & ~n67626 ;
  assign n67631 = ~n11599 & n67627 ;
  assign n67632 = ~n67630 & ~n67631 ;
  assign n67633 = ~n11577 & ~n67632 ;
  assign n67629 = n11577 & ~n12817 ;
  assign n67634 = n27681 & ~n67629 ;
  assign n67635 = ~n67633 & n67634 ;
  assign n67622 = n11919 & ~n12807 ;
  assign n67623 = ~n67621 & ~n67622 ;
  assign n67624 = n11692 & ~n67623 ;
  assign n67620 = \P2_P1_InstQueue_reg[12][6]/NET0131  & ~n11630 ;
  assign n67628 = n36674 & ~n67627 ;
  assign n67636 = ~n67620 & ~n67628 ;
  assign n67637 = ~n67624 & n67636 ;
  assign n67638 = ~n67635 & n67637 ;
  assign n67649 = n11596 & ~n14576 ;
  assign n67644 = n11378 & ~n11961 ;
  assign n67640 = \P2_P1_InstQueue_reg[13][5]/NET0131  & ~n11862 ;
  assign n67645 = ~n11919 & n67640 ;
  assign n67646 = ~n67644 & ~n67645 ;
  assign n67650 = ~n11596 & n67646 ;
  assign n67651 = ~n67649 & ~n67650 ;
  assign n67652 = ~n11599 & ~n67651 ;
  assign n67648 = n11599 & ~n14573 ;
  assign n67653 = n27681 & ~n67648 ;
  assign n67654 = ~n67652 & n67653 ;
  assign n67641 = n11862 & ~n14612 ;
  assign n67642 = ~n67640 & ~n67641 ;
  assign n67643 = n11692 & ~n67642 ;
  assign n67639 = \P2_P1_InstQueue_reg[13][5]/NET0131  & ~n11630 ;
  assign n67647 = n36674 & ~n67646 ;
  assign n67655 = ~n67639 & ~n67647 ;
  assign n67656 = ~n67643 & n67655 ;
  assign n67657 = ~n67654 & n67656 ;
  assign n67668 = n11873 & ~n14576 ;
  assign n67663 = n11378 & ~n12024 ;
  assign n67659 = \P2_P1_InstQueue_reg[1][5]/NET0131  & ~n12023 ;
  assign n67664 = ~n11871 & n67659 ;
  assign n67665 = ~n67663 & ~n67664 ;
  assign n67669 = ~n11873 & n67665 ;
  assign n67670 = ~n67668 & ~n67669 ;
  assign n67671 = ~n11865 & ~n67670 ;
  assign n67667 = n11865 & ~n14573 ;
  assign n67672 = n27681 & ~n67667 ;
  assign n67673 = ~n67671 & n67672 ;
  assign n67660 = n12023 & ~n14612 ;
  assign n67661 = ~n67659 & ~n67660 ;
  assign n67662 = n11692 & ~n67661 ;
  assign n67658 = \P2_P1_InstQueue_reg[1][5]/NET0131  & ~n11630 ;
  assign n67666 = n36674 & ~n67665 ;
  assign n67674 = ~n67658 & ~n67666 ;
  assign n67675 = ~n67662 & n67674 ;
  assign n67676 = ~n67673 & n67675 ;
  assign n67687 = n11865 & ~n14576 ;
  assign n67682 = n11378 & ~n11874 ;
  assign n67678 = \P2_P1_InstQueue_reg[0][5]/NET0131  & ~n11871 ;
  assign n67683 = ~n11873 & n67678 ;
  assign n67684 = ~n67682 & ~n67683 ;
  assign n67688 = ~n11865 & n67684 ;
  assign n67689 = ~n67687 & ~n67688 ;
  assign n67690 = ~n11862 & ~n67689 ;
  assign n67686 = n11862 & ~n14573 ;
  assign n67691 = n27681 & ~n67686 ;
  assign n67692 = ~n67690 & n67691 ;
  assign n67679 = n11871 & ~n14612 ;
  assign n67680 = ~n67678 & ~n67679 ;
  assign n67681 = n11692 & ~n67680 ;
  assign n67677 = \P2_P1_InstQueue_reg[0][5]/NET0131  & ~n11630 ;
  assign n67685 = n36674 & ~n67684 ;
  assign n67693 = ~n67677 & ~n67685 ;
  assign n67694 = ~n67681 & n67693 ;
  assign n67695 = ~n67692 & n67694 ;
  assign n67706 = n11871 & ~n14576 ;
  assign n67701 = n11378 & ~n12066 ;
  assign n67697 = \P2_P1_InstQueue_reg[2][5]/NET0131  & ~n12065 ;
  assign n67702 = ~n12023 & n67697 ;
  assign n67703 = ~n67701 & ~n67702 ;
  assign n67707 = ~n11871 & n67703 ;
  assign n67708 = ~n67706 & ~n67707 ;
  assign n67709 = ~n11873 & ~n67708 ;
  assign n67705 = n11873 & ~n14573 ;
  assign n67710 = n27681 & ~n67705 ;
  assign n67711 = ~n67709 & n67710 ;
  assign n67698 = n12065 & ~n14612 ;
  assign n67699 = ~n67697 & ~n67698 ;
  assign n67700 = n11692 & ~n67699 ;
  assign n67696 = \P2_P1_InstQueue_reg[2][5]/NET0131  & ~n11630 ;
  assign n67704 = n36674 & ~n67703 ;
  assign n67712 = ~n67696 & ~n67704 ;
  assign n67713 = ~n67700 & n67712 ;
  assign n67714 = ~n67711 & n67713 ;
  assign n67725 = n12109 & ~n14576 ;
  assign n67720 = n11378 & ~n12174 ;
  assign n67716 = \P2_P1_InstQueue_reg[6][5]/NET0131  & ~n12173 ;
  assign n67721 = ~n12131 & n67716 ;
  assign n67722 = ~n67720 & ~n67721 ;
  assign n67726 = ~n12109 & n67722 ;
  assign n67727 = ~n67725 & ~n67726 ;
  assign n67728 = ~n12087 & ~n67727 ;
  assign n67724 = n12087 & ~n14573 ;
  assign n67729 = n27681 & ~n67724 ;
  assign n67730 = ~n67728 & n67729 ;
  assign n67717 = n12173 & ~n14612 ;
  assign n67718 = ~n67716 & ~n67717 ;
  assign n67719 = n11692 & ~n67718 ;
  assign n67715 = \P2_P1_InstQueue_reg[6][5]/NET0131  & ~n11630 ;
  assign n67723 = n36674 & ~n67722 ;
  assign n67731 = ~n67715 & ~n67723 ;
  assign n67732 = ~n67719 & n67731 ;
  assign n67733 = ~n67730 & n67732 ;
  assign n67744 = n11599 & ~n14576 ;
  assign n67739 = n11378 & ~n11920 ;
  assign n67735 = \P2_P1_InstQueue_reg[12][5]/NET0131  & ~n11919 ;
  assign n67740 = ~n11596 & n67735 ;
  assign n67741 = ~n67739 & ~n67740 ;
  assign n67745 = ~n11599 & n67741 ;
  assign n67746 = ~n67744 & ~n67745 ;
  assign n67747 = ~n11577 & ~n67746 ;
  assign n67743 = n11577 & ~n14573 ;
  assign n67748 = n27681 & ~n67743 ;
  assign n67749 = ~n67747 & n67748 ;
  assign n67736 = n11919 & ~n14612 ;
  assign n67737 = ~n67735 & ~n67736 ;
  assign n67738 = n11692 & ~n67737 ;
  assign n67734 = \P2_P1_InstQueue_reg[12][5]/NET0131  & ~n11630 ;
  assign n67742 = n36674 & ~n67741 ;
  assign n67750 = ~n67734 & ~n67742 ;
  assign n67751 = ~n67738 & n67750 ;
  assign n67752 = ~n67749 & n67751 ;
  assign n67763 = n11862 & ~n14576 ;
  assign n67758 = n11378 & ~n12002 ;
  assign n67754 = \P2_P1_InstQueue_reg[15][5]/NET0131  & ~n11873 ;
  assign n67759 = ~n11865 & n67754 ;
  assign n67760 = ~n67758 & ~n67759 ;
  assign n67764 = ~n11862 & n67760 ;
  assign n67765 = ~n67763 & ~n67764 ;
  assign n67766 = ~n11919 & ~n67765 ;
  assign n67762 = n11919 & ~n14573 ;
  assign n67767 = n27681 & ~n67762 ;
  assign n67768 = ~n67766 & n67767 ;
  assign n67755 = n11873 & ~n14612 ;
  assign n67756 = ~n67754 & ~n67755 ;
  assign n67757 = n11692 & ~n67756 ;
  assign n67753 = \P2_P1_InstQueue_reg[15][5]/NET0131  & ~n11630 ;
  assign n67761 = n36674 & ~n67760 ;
  assign n67769 = ~n67753 & ~n67761 ;
  assign n67770 = ~n67757 & n67769 ;
  assign n67771 = ~n67768 & n67770 ;
  assign n67782 = n12173 & ~n14576 ;
  assign n67777 = n11378 & ~n11895 ;
  assign n67773 = \P2_P1_InstQueue_reg[8][5]/NET0131  & ~n10105 ;
  assign n67778 = ~n11891 & n67773 ;
  assign n67779 = ~n67777 & ~n67778 ;
  assign n67783 = ~n12173 & n67779 ;
  assign n67784 = ~n67782 & ~n67783 ;
  assign n67785 = ~n12131 & ~n67784 ;
  assign n67781 = n12131 & ~n14573 ;
  assign n67786 = n27681 & ~n67781 ;
  assign n67787 = ~n67785 & n67786 ;
  assign n67774 = n10105 & ~n14612 ;
  assign n67775 = ~n67773 & ~n67774 ;
  assign n67776 = n11692 & ~n67775 ;
  assign n67772 = \P2_P1_InstQueue_reg[8][5]/NET0131  & ~n11630 ;
  assign n67780 = n36674 & ~n67779 ;
  assign n67788 = ~n67772 & ~n67780 ;
  assign n67789 = ~n67776 & n67788 ;
  assign n67790 = ~n67787 & n67789 ;
  assign n67801 = n12131 & ~n14576 ;
  assign n67796 = n11378 & ~n12195 ;
  assign n67792 = \P2_P1_InstQueue_reg[7][5]/NET0131  & ~n11891 ;
  assign n67797 = ~n12173 & n67792 ;
  assign n67798 = ~n67796 & ~n67797 ;
  assign n67802 = ~n12131 & n67798 ;
  assign n67803 = ~n67801 & ~n67802 ;
  assign n67804 = ~n12109 & ~n67803 ;
  assign n67800 = n12109 & ~n14573 ;
  assign n67805 = n27681 & ~n67800 ;
  assign n67806 = ~n67804 & n67805 ;
  assign n67793 = n11891 & ~n14612 ;
  assign n67794 = ~n67792 & ~n67793 ;
  assign n67795 = n11692 & ~n67794 ;
  assign n67791 = \P2_P1_InstQueue_reg[7][5]/NET0131  & ~n11630 ;
  assign n67799 = n36674 & ~n67798 ;
  assign n67807 = ~n67791 & ~n67799 ;
  assign n67808 = ~n67795 & n67807 ;
  assign n67809 = ~n67806 & n67808 ;
  assign \P3_state_reg[0]/NET0131_syn_2  = ~\P3_rd_reg/NET0131  ;
  assign \_al_n1  = ~1'b0 ;
  assign \aux[0]_pad  = n2835 ;
  assign \aux[1]_pad  = ~n2849 ;
  assign \aux[2]_pad  = n2869 ;
  assign \dout[0]_pad  = n2873 ;
  assign \dout[10]_pad  = n3355 ;
  assign \dout[11]_pad  = ~n3450 ;
  assign \dout[12]_pad  = ~n3548 ;
  assign \dout[13]_pad  = ~n3658 ;
  assign \dout[14]_pad  = n3770 ;
  assign \dout[15]_pad  = ~n3892 ;
  assign \dout[16]_pad  = n4018 ;
  assign \dout[17]_pad  = ~n4156 ;
  assign \dout[18]_pad  = n4290 ;
  assign \dout[19]_pad  = 1'b0 ;
  assign \dout[1]_pad  = ~n4294 ;
  assign \dout[2]_pad  = n4296 ;
  assign \dout[3]_pad  = ~n4300 ;
  assign \dout[4]_pad  = ~n4304 ;
  assign \dout[5]_pad  = ~n4308 ;
  assign \dout[6]_pad  = ~n4312 ;
  assign \dout[7]_pad  = ~n4316 ;
  assign \dout[8]_pad  = n4320 ;
  assign \dout[9]_pad  = n4324 ;
  assign \g326201/_0_  = ~n8370 ;
  assign \g326202/_0_  = ~n8400 ;
  assign \g326203/_0_  = ~n8424 ;
  assign \g326204/_0_  = ~n8449 ;
  assign \g326205/_0_  = ~n8472 ;
  assign \g326206/_0_  = ~n8495 ;
  assign \g326207/_0_  = ~n8518 ;
  assign \g326208/_0_  = ~n8542 ;
  assign \g326209/_0_  = ~n8566 ;
  assign \g326210/_0_  = ~n8590 ;
  assign \g326211/_0_  = ~n8614 ;
  assign \g326212/_0_  = ~n8638 ;
  assign \g326213/_0_  = ~n8662 ;
  assign \g326214/_0_  = ~n8685 ;
  assign \g326215/_0_  = ~n8707 ;
  assign \g326216/_0_  = ~n8730 ;
  assign \g326251/_0_  = ~n9251 ;
  assign \g326255/_0_  = ~n9310 ;
  assign \g326256/_0_  = ~n9369 ;
  assign \g326271/_0_  = ~n9391 ;
  assign \g326272/_0_  = ~n9413 ;
  assign \g326273/_0_  = ~n9433 ;
  assign \g326274/_0_  = ~n9454 ;
  assign \g326275/_0_  = ~n9476 ;
  assign \g326276/_0_  = ~n9498 ;
  assign \g326277/_0_  = ~n9520 ;
  assign \g326278/_0_  = ~n9542 ;
  assign \g326279/_0_  = ~n9564 ;
  assign \g326280/_0_  = ~n9586 ;
  assign \g326281/_0_  = ~n9608 ;
  assign \g326282/_0_  = ~n9630 ;
  assign \g326283/_0_  = ~n9652 ;
  assign \g326284/_0_  = ~n9674 ;
  assign \g326285/_0_  = ~n9696 ;
  assign \g326286/_0_  = ~n9718 ;
  assign \g326287/_0_  = ~n9740 ;
  assign \g326288/_0_  = ~n9762 ;
  assign \g326289/_0_  = ~n9784 ;
  assign \g326290/_0_  = ~n9806 ;
  assign \g326291/_0_  = ~n9828 ;
  assign \g326292/_0_  = ~n9850 ;
  assign \g326293/_0_  = ~n9872 ;
  assign \g326294/_0_  = ~n9894 ;
  assign \g326295/_0_  = ~n9916 ;
  assign \g326296/_0_  = ~n9938 ;
  assign \g326297/_0_  = ~n9960 ;
  assign \g326298/_0_  = ~n9982 ;
  assign \g326299/_0_  = ~n10004 ;
  assign \g326300/_0_  = ~n10026 ;
  assign \g326301/_0_  = ~n10045 ;
  assign \g326335/_0_  = ~n10047 ;
  assign \g326369/_0_  = ~n10102 ;
  assign \g326370/_0_  = ~n11696 ;
  assign \g326371/_0_  = ~n11701 ;
  assign \g326372/_0_  = ~n11721 ;
  assign \g326373/_0_  = ~n11740 ;
  assign \g326374/_0_  = ~n11760 ;
  assign \g326375/_0_  = ~n11780 ;
  assign \g326376/_0_  = ~n11800 ;
  assign \g326377/_0_  = ~n11820 ;
  assign \g326378/_0_  = ~n11840 ;
  assign \g326379/_0_  = ~n11860 ;
  assign \g326380/_0_  = ~n11889 ;
  assign \g326381/_0_  = ~n11912 ;
  assign \g326382/_0_  = ~n11935 ;
  assign \g326383/_0_  = ~n11955 ;
  assign \g326384/_0_  = ~n11976 ;
  assign \g326385/_0_  = ~n11996 ;
  assign \g326386/_0_  = ~n12017 ;
  assign \g326387/_0_  = ~n12039 ;
  assign \g326388/_0_  = ~n12059 ;
  assign \g326389/_0_  = ~n12081 ;
  assign \g326390/_0_  = ~n12103 ;
  assign \g326391/_0_  = ~n12125 ;
  assign \g326392/_0_  = ~n12147 ;
  assign \g326393/_0_  = ~n12167 ;
  assign \g326394/_0_  = ~n12189 ;
  assign \g326395/_0_  = ~n12210 ;
  assign \g326396/_0_  = ~n12230 ;
  assign \g326397/_0_  = ~n12250 ;
  assign \g326398/_0_  = ~n12270 ;
  assign \g326399/_0_  = ~n12290 ;
  assign \g326400/_0_  = ~n12310 ;
  assign \g326401/_0_  = ~n12330 ;
  assign \g326423/_0_  = ~n12386 ;
  assign \g326438/_0_  = ~n12405 ;
  assign \g326439/_0_  = ~n12424 ;
  assign \g326440/_0_  = ~n12443 ;
  assign \g326441/_0_  = ~n12462 ;
  assign \g326442/_0_  = ~n12481 ;
  assign \g326443/_0_  = ~n12500 ;
  assign \g326444/_0_  = ~n12519 ;
  assign \g326445/_0_  = ~n12538 ;
  assign \g326446/_0_  = ~n12557 ;
  assign \g326447/_0_  = ~n12576 ;
  assign \g326448/_0_  = ~n12595 ;
  assign \g326449/_0_  = ~n12614 ;
  assign \g326450/_0_  = ~n12633 ;
  assign \g326451/_0_  = ~n12652 ;
  assign \g326452/_0_  = ~n12671 ;
  assign \g326561/_0_  = ~n12725 ;
  assign \g326571/_0_  = ~n12774 ;
  assign \g326572/_0_  = ~n12828 ;
  assign \g326597/_0_  = ~n12847 ;
  assign \g326598/_0_  = ~n12866 ;
  assign \g326599/_0_  = ~n12885 ;
  assign \g326600/_0_  = ~n12904 ;
  assign \g326601/_0_  = ~n12923 ;
  assign \g326602/_0_  = ~n12942 ;
  assign \g326603/_0_  = ~n12961 ;
  assign \g326604/_0_  = ~n12975 ;
  assign \g326605/_0_  = ~n12994 ;
  assign \g326606/_0_  = ~n13013 ;
  assign \g326607/_0_  = ~n13027 ;
  assign \g326608/_0_  = ~n13046 ;
  assign \g326609/_0_  = ~n13060 ;
  assign \g326611/_0_  = ~n13079 ;
  assign \g326612/_0_  = ~n13093 ;
  assign \g326613/_0_  = ~n13112 ;
  assign \g326614/_0_  = ~n13126 ;
  assign \g326615/_0_  = ~n13145 ;
  assign \g326616/_0_  = ~n13159 ;
  assign \g326617/_0_  = ~n13178 ;
  assign \g326618/_0_  = ~n13192 ;
  assign \g326619/_0_  = ~n13211 ;
  assign \g326620/_0_  = ~n13230 ;
  assign \g326621/_0_  = ~n13244 ;
  assign \g326622/_0_  = ~n13263 ;
  assign \g326623/_0_  = ~n13277 ;
  assign \g326624/_0_  = ~n13296 ;
  assign \g326625/_0_  = ~n13310 ;
  assign \g326626/_0_  = ~n13329 ;
  assign \g326627/_0_  = ~n13343 ;
  assign \g326628/_0_  = ~n13362 ;
  assign \g326629/_0_  = ~n13381 ;
  assign \g326630/_0_  = ~n13395 ;
  assign \g326631/_0_  = ~n13414 ;
  assign \g326632/_0_  = ~n13428 ;
  assign \g326633/_0_  = ~n13447 ;
  assign \g326634/_0_  = ~n13461 ;
  assign \g326635/_0_  = ~n13480 ;
  assign \g326636/_0_  = ~n13494 ;
  assign \g326637/_0_  = ~n13513 ;
  assign \g326638/_0_  = ~n13532 ;
  assign \g326639/_0_  = ~n13551 ;
  assign \g326640/_0_  = ~n13570 ;
  assign \g326641/_0_  = ~n13589 ;
  assign \g326798/_0_  = ~n13646 ;
  assign \g326821/_0_  = ~n13668 ;
  assign \g326822/_0_  = ~n13687 ;
  assign \g326823/_0_  = ~n13709 ;
  assign \g326824/_0_  = ~n13731 ;
  assign \g326825/_0_  = ~n13753 ;
  assign \g326826/_0_  = ~n13775 ;
  assign \g326827/_0_  = ~n13797 ;
  assign \g326828/_0_  = ~n13819 ;
  assign \g326829/_0_  = ~n13841 ;
  assign \g326830/_0_  = ~n13863 ;
  assign \g326831/_0_  = ~n13885 ;
  assign \g326832/_0_  = ~n13907 ;
  assign \g326833/_0_  = ~n13929 ;
  assign \g326834/_0_  = ~n13951 ;
  assign \g326835/_0_  = ~n13973 ;
  assign \g326868/_0_  = ~n14027 ;
  assign \g326887/_0_  = ~n14076 ;
  assign \g326926/_0_  = ~n14095 ;
  assign \g326927/_0_  = ~n14114 ;
  assign \g326928/_0_  = ~n14133 ;
  assign \g326929/_0_  = ~n14152 ;
  assign \g326930/_0_  = ~n14171 ;
  assign \g326931/_0_  = ~n14190 ;
  assign \g326932/_0_  = ~n14209 ;
  assign \g326933/_0_  = ~n14228 ;
  assign \g326934/_0_  = ~n14242 ;
  assign \g326935/_0_  = ~n14256 ;
  assign \g326936/_0_  = ~n14275 ;
  assign \g326937/_0_  = ~n14289 ;
  assign \g326938/_0_  = ~n14303 ;
  assign \g326939/_0_  = ~n14317 ;
  assign \g326940/_0_  = ~n14331 ;
  assign \g326941/_0_  = ~n14345 ;
  assign \g326942/_0_  = ~n14364 ;
  assign \g326943/_0_  = ~n14378 ;
  assign \g326944/_0_  = ~n14392 ;
  assign \g326945/_0_  = ~n14406 ;
  assign \g326946/_0_  = ~n14420 ;
  assign \g326947/_0_  = ~n14439 ;
  assign \g326948/_0_  = ~n14453 ;
  assign \g326949/_0_  = ~n14467 ;
  assign \g326950/_0_  = ~n14481 ;
  assign \g326951/_0_  = ~n14495 ;
  assign \g326952/_0_  = ~n14514 ;
  assign \g326953/_0_  = ~n14533 ;
  assign \g326954/_0_  = ~n14552 ;
  assign \g326955/_0_  = ~n14571 ;
  assign \g327192/_0_  = ~n14620 ;
  assign \g327234/_0_  = ~n14634 ;
  assign \g327237/_0_  = ~n14648 ;
  assign \g327241/_0_  = ~n14662 ;
  assign \g327242/_0_  = ~n14676 ;
  assign \g327243/_0_  = ~n14690 ;
  assign \g327247/_0_  = ~n14704 ;
  assign \g327290/_0_  = ~n14758 ;
  assign \g327311/_0_  = ~n14807 ;
  assign \g327369/_0_  = ~n14826 ;
  assign \g327370/_0_  = ~n14845 ;
  assign \g327371/_0_  = ~n14864 ;
  assign \g327373/_0_  = ~n14883 ;
  assign \g327375/_0_  = ~n14902 ;
  assign \g327377/_0_  = ~n14921 ;
  assign \g327379/_0_  = ~n14940 ;
  assign \g327380/_0_  = ~n14959 ;
  assign \g327381/_0_  = ~n14973 ;
  assign \g327382/_0_  = ~n14987 ;
  assign \g327383/_0_  = ~n15006 ;
  assign \g327384/_0_  = ~n15020 ;
  assign \g327385/_0_  = ~n15034 ;
  assign \g327386/_0_  = ~n15048 ;
  assign \g327387/_0_  = ~n15062 ;
  assign \g327388/_0_  = ~n15081 ;
  assign \g327389/_0_  = ~n15095 ;
  assign \g327390/_0_  = ~n15109 ;
  assign \g327391/_0_  = ~n15123 ;
  assign \g327392/_0_  = ~n15137 ;
  assign \g327393/_0_  = ~n15156 ;
  assign \g327394/_0_  = ~n15170 ;
  assign \g327395/_0_  = ~n15184 ;
  assign \g327396/_0_  = ~n15198 ;
  assign \g327397/_0_  = ~n15212 ;
  assign \g327398/_0_  = ~n15231 ;
  assign \g327399/_0_  = ~n15245 ;
  assign \g327400/_0_  = ~n15264 ;
  assign \g327401/_0_  = ~n15283 ;
  assign \g327402/_0_  = ~n15302 ;
  assign \g327601/_0_  = ~n15321 ;
  assign \g327602/_0_  = ~n15732 ;
  assign \g327698/_0_  = ~n16445 ;
  assign \g327781/_0_  = ~n16528 ;
  assign \g327798/_0_  = ~n16625 ;
  assign \g327799/_0_  = ~n16663 ;
  assign \g327800/_0_  = ~n16704 ;
  assign \g327801/_0_  = ~n16742 ;
  assign \g327802/_0_  = ~n16788 ;
  assign \g327803/_0_  = ~n16831 ;
  assign \g327804/_0_  = ~n16872 ;
  assign \g327805/_0_  = ~n16909 ;
  assign \g327806/_0_  = ~n16947 ;
  assign \g327807/_0_  = ~n16956 ;
  assign \g327826/_0_  = ~n16965 ;
  assign \g327828/_0_  = ~n17029 ;
  assign \g327829/_0_  = ~n17075 ;
  assign \g327830/_0_  = ~n17121 ;
  assign \g327831/_0_  = ~n17163 ;
  assign \g327832/_0_  = ~n17208 ;
  assign \g327833/_0_  = ~n17250 ;
  assign \g327834/_0_  = ~n17292 ;
  assign \g327835/_0_  = ~n17334 ;
  assign \g327836/_0_  = ~n17376 ;
  assign \g327970/_0_  = ~n17425 ;
  assign \g328019/_0_  = ~n17463 ;
  assign \g328020/_0_  = ~n17496 ;
  assign \g328021/_0_  = ~n17529 ;
  assign \g328022/_0_  = ~n17565 ;
  assign \g328023/_0_  = ~n17602 ;
  assign \g328024/_0_  = ~n17638 ;
  assign \g328027/_0_  = ~n17678 ;
  assign \g328028/_0_  = ~n17715 ;
  assign \g328029/_0_  = ~n17750 ;
  assign \g328030/_0_  = ~n17788 ;
  assign \g328031/_0_  = ~n17826 ;
  assign \g328032/_0_  = ~n17860 ;
  assign \g328033/_0_  = ~n17896 ;
  assign \g328034/_0_  = ~n17933 ;
  assign \g328035/_0_  = ~n17968 ;
  assign \g328046/_0_  = ~n17982 ;
  assign \g328048/_0_  = ~n17996 ;
  assign \g328049/_0_  = ~n18010 ;
  assign \g328052/_0_  = ~n18024 ;
  assign \g328054/_0_  = ~n18038 ;
  assign \g328056/_0_  = ~n18052 ;
  assign \g328058/_0_  = ~n18066 ;
  assign \g328059/_0_  = ~n18080 ;
  assign \g328060/_0_  = ~n18094 ;
  assign \g328061/_0_  = ~n18108 ;
  assign \g328062/_0_  = ~n18122 ;
  assign \g328063/_0_  = ~n18136 ;
  assign \g328064/_0_  = ~n18150 ;
  assign \g328065/_0_  = ~n18164 ;
  assign \g328066/_0_  = ~n18178 ;
  assign \g328067/_0_  = ~n18197 ;
  assign \g328068/_0_  = ~n18232 ;
  assign \g328069/_0_  = ~n18273 ;
  assign \g328070/_0_  = ~n18309 ;
  assign \g328071/_0_  = ~n18338 ;
  assign \g328120/_0_  = ~n18448 ;
  assign \g328152/_0_  = ~n18681 ;
  assign \g328153/_0_  = ~n18751 ;
  assign \g328154/_0_  = ~n18799 ;
  assign \g328155/_0_  = ~n18810 ;
  assign \g328156/_0_  = ~n18859 ;
  assign \g328157/_0_  = ~n18900 ;
  assign \g328158/_0_  = ~n18941 ;
  assign \g328159/_0_  = ~n18982 ;
  assign \g328160/_0_  = ~n19025 ;
  assign \g328161/_0_  = ~n19071 ;
  assign \g328257/_0_  = ~n19121 ;
  assign \g328280/_0_  = ~n19151 ;
  assign \g328302/_0_  = ~n19169 ;
  assign \g328303/_0_  = ~n19189 ;
  assign \g328332/_0_  = ~n19386 ;
  assign \g328333/_0_  = ~n19428 ;
  assign \g328334/_0_  = ~n19477 ;
  assign \g328335/_0_  = ~n19525 ;
  assign \g328336/_0_  = ~n19566 ;
  assign \g328337/_0_  = ~n19607 ;
  assign \g328338/_0_  = ~n19664 ;
  assign \g328339/_0_  = ~n19705 ;
  assign \g328340/_0_  = ~n19755 ;
  assign \g328341/_0_  = ~n19801 ;
  assign \g328342/_0_  = ~n19844 ;
  assign \g328343/_0_  = ~n19897 ;
  assign \g328344/_0_  = ~n19947 ;
  assign \g328345/_0_  = ~n19993 ;
  assign \g328346/_0_  = ~n20038 ;
  assign \g328347/_0_  = ~n20081 ;
  assign \g328348/_0_  = ~n20129 ;
  assign \g328349/_0_  = ~n20177 ;
  assign \g328350/_0_  = ~n20219 ;
  assign \g328351/_0_  = ~n20263 ;
  assign \g328352/_0_  = ~n20297 ;
  assign \g328353/_0_  = ~n20336 ;
  assign \g328354/_0_  = ~n20383 ;
  assign \g328355/_0_  = ~n20429 ;
  assign \g328356/_0_  = ~n20465 ;
  assign \g328357/_0_  = ~n20499 ;
  assign \g328358/_0_  = ~n20546 ;
  assign \g328359/_0_  = ~n20586 ;
  assign \g328360/_0_  = ~n20616 ;
  assign \g328361/_0_  = ~n20660 ;
  assign \g328372/_0_  = ~n20667 ;
  assign \g328373/_0_  = ~n20670 ;
  assign \g328374/_0_  = ~n20692 ;
  assign \g328375/_0_  = ~n21102 ;
  assign \g328376/_0_  = ~n21110 ;
  assign \g328377/_0_  = ~n21159 ;
  assign \g328378/_0_  = ~n21207 ;
  assign \g328379/_0_  = ~n21253 ;
  assign \g328380/_0_  = ~n21301 ;
  assign \g328381/_0_  = ~n21349 ;
  assign \g328382/_0_  = ~n21432 ;
  assign \g328383/_0_  = ~n21490 ;
  assign \g328384/_0_  = ~n21678 ;
  assign \g328385/_0_  = ~n21730 ;
  assign \g328569/_0_  = ~n21765 ;
  assign \g328587/_0_  = ~n21781 ;
  assign \g328658/_0_  = ~n21849 ;
  assign \g328662/_3_  = ~n21858 ;
  assign \g328664/_3_  = ~n21861 ;
  assign \g328666/_3_  = ~n21914 ;
  assign \g328669/_3_  = ~n21930 ;
  assign \g328670/_0_  = ~n21950 ;
  assign \g328671/_0_  = ~n21965 ;
  assign \g328672/_0_  = ~n21968 ;
  assign \g328674/_0_  = ~n21971 ;
  assign \g328809/_0_  = ~n22007 ;
  assign \g328810/_0_  = ~n22039 ;
  assign \g328811/_0_  = ~n22072 ;
  assign \g328812/_0_  = ~n22104 ;
  assign \g328856/_0_  = ~n22114 ;
  assign \g328887/_0_  = n22125 ;
  assign \g328931/_0_  = ~n22170 ;
  assign \g328945/_0_  = ~n22186 ;
  assign \g328960/_0_  = ~n22217 ;
  assign \g328991/_0_  = ~n22253 ;
  assign \g328992/_0_  = ~n22276 ;
  assign \g329022/_3_  = ~n22279 ;
  assign \g329024/_3_  = ~n22287 ;
  assign \g329025/_0_  = ~n22295 ;
  assign \g329026/_0_  = ~n22300 ;
  assign \g329027/_0_  = ~n22305 ;
  assign \g329029/_3_  = ~n22332 ;
  assign \g329030/_0_  = ~n22355 ;
  assign \g329032/_0_  = ~n22376 ;
  assign \g329033/_0_  = ~n22395 ;
  assign \g329034/_0_  = ~n22414 ;
  assign \g329182/_0_  = ~n22449 ;
  assign \g329228/_0_  = ~n22482 ;
  assign \g329281/_0_  = ~n22519 ;
  assign \g329301/_0_  = ~n22550 ;
  assign \g329302/_0_  = ~n22559 ;
  assign \g329322/_2_  = ~n22572 ;
  assign \g329324/_3_  = ~n22603 ;
  assign \g329334/_3_  = ~n22606 ;
  assign \g329336/_3_  = ~n22609 ;
  assign \g329338/_3_  = ~n22612 ;
  assign \g329340/_2_  = ~n22631 ;
  assign \g329342/_3_  = ~n22634 ;
  assign \g329343/_0_  = ~n22639 ;
  assign \g329345/_3_  = ~n22653 ;
  assign \g329347/_3_  = ~n22656 ;
  assign \g329349/_3_  = ~n22659 ;
  assign \g329351/_3_  = ~n22662 ;
  assign \g329353/_3_  = ~n22665 ;
  assign \g329355/_3_  = ~n22668 ;
  assign \g329357/_3_  = ~n22671 ;
  assign \g329359/_3_  = ~n22679 ;
  assign \g329360/_0_  = ~n22682 ;
  assign \g329362/_3_  = ~n22692 ;
  assign \g329364/_3_  = ~n22696 ;
  assign \g329366/_3_  = ~n22701 ;
  assign \g329368/_3_  = ~n22717 ;
  assign \g329370/_3_  = ~n22728 ;
  assign \g329372/_3_  = ~n22744 ;
  assign \g329374/_3_  = ~n22760 ;
  assign \g329376/_3_  = ~n22776 ;
  assign \g329378/_3_  = ~n22792 ;
  assign \g329379/_0_  = ~n22814 ;
  assign \g329380/_0_  = ~n22847 ;
  assign \g329381/_0_  = ~n22871 ;
  assign \g329388/_0_  = ~n22904 ;
  assign \g329516/_0_  = ~n22948 ;
  assign \g329517/_0_  = ~n22980 ;
  assign \g329518/_0_  = ~n23013 ;
  assign \g329587/_0_  = ~n23028 ;
  assign \g329605/_0_  = ~n23060 ;
  assign \g329687/_0_  = ~n23100 ;
  assign \g329703/_0_  = ~n23109 ;
  assign \g329709/_3_  = ~n23129 ;
  assign \g329716/_3_  = ~n23137 ;
  assign \g329718/_3_  = ~n23140 ;
  assign \g329720/_3_  = ~n23143 ;
  assign \g329722/_3_  = ~n23151 ;
  assign \g329724/_3_  = ~n23157 ;
  assign \g329725/_0_  = ~n23179 ;
  assign \g329727/_0_  = ~n23203 ;
  assign \g329805/_0_  = ~n23234 ;
  assign \g329807/_0_  = ~n23269 ;
  assign \g329809/_0_  = n23303 ;
  assign \g329810/_0_  = ~n23332 ;
  assign \g329811/_0_  = ~n23364 ;
  assign \g329812/_0_  = ~n23399 ;
  assign \g330065/_3_  = ~n23407 ;
  assign \g330067/_3_  = ~n23430 ;
  assign \g330069/_3_  = ~n23435 ;
  assign \g330071/_3_  = ~n23444 ;
  assign \g330073/_3_  = ~n23447 ;
  assign \g330075/_3_  = ~n23450 ;
  assign \g330077/_3_  = ~n23458 ;
  assign \g330079/_3_  = n23473 ;
  assign \g330081/_3_  = ~n23476 ;
  assign \g330083/_3_  = ~n23479 ;
  assign \g330085/_3_  = ~n23482 ;
  assign \g330087/_3_  = ~n23485 ;
  assign \g330089/_3_  = ~n23507 ;
  assign \g330091/_3_  = ~n23527 ;
  assign \g330093/_3_  = n23540 ;
  assign \g330095/_3_  = ~n23556 ;
  assign \g330097/_3_  = ~n23562 ;
  assign \g330099/_0_  = ~n23587 ;
  assign \g330188/_0_  = ~n23618 ;
  assign \g330337/_0_  = ~n23656 ;
  assign \g330388/_3_  = ~n23676 ;
  assign \g330418/_3_  = ~n23683 ;
  assign \g330420/_3_  = ~n23703 ;
  assign \g330422/_3_  = ~n23711 ;
  assign \g330424/_3_  = ~n23714 ;
  assign \g330426/_3_  = ~n23717 ;
  assign \g330428/_3_  = ~n23725 ;
  assign \g330429/_0_  = ~n23748 ;
  assign \g330431/_3_  = ~n23759 ;
  assign \g330433/_3_  = ~n23776 ;
  assign \g330435/_3_  = ~n23779 ;
  assign \g330436/_0_  = ~n23800 ;
  assign \g330438/_3_  = ~n23803 ;
  assign \g330440/_3_  = ~n23819 ;
  assign \g330441/_0_  = ~n23840 ;
  assign \g330443/_3_  = ~n23853 ;
  assign \g330444/_0_  = ~n23872 ;
  assign \g330446/_3_  = ~n23888 ;
  assign \g330448/_3_  = ~n23904 ;
  assign \g330450/_3_  = ~n23917 ;
  assign \g330451/_0_  = ~n23941 ;
  assign \g330452/_0_  = ~n23962 ;
  assign \g330453/_0_  = ~n23986 ;
  assign \g330535/_0_  = ~n24006 ;
  assign \g330762/_3_  = ~n24009 ;
  assign \g330764/_3_  = ~n24012 ;
  assign \g330766/_3_  = ~n24015 ;
  assign \g330768/_3_  = ~n24037 ;
  assign \g330770/_3_  = ~n24040 ;
  assign \g330772/_3_  = ~n24061 ;
  assign \g330774/_3_  = ~n24077 ;
  assign \g330776/_3_  = ~n24093 ;
  assign \g331141/_3_  = ~n24101 ;
  assign \g331142/_0_  = ~n24122 ;
  assign \g331144/_3_  = ~n24125 ;
  assign \g331145/_0_  = ~n24146 ;
  assign \g331147/_3_  = ~n24157 ;
  assign \g331484/_0_  = ~n24208 ;
  assign \g331485/_0_  = ~n24259 ;
  assign \g331486/_0_  = ~n24307 ;
  assign \g331497/_0_  = ~n24355 ;
  assign \g331498/_0_  = ~n24399 ;
  assign \g331502/_0_  = ~n24449 ;
  assign \g332061/_0_  = ~n24499 ;
  assign \g332062/_0_  = ~n24517 ;
  assign \g332063/_0_  = ~n24558 ;
  assign \g332064/_0_  = ~n24607 ;
  assign \g332065/_0_  = ~n24657 ;
  assign \g332066/_0_  = ~n24706 ;
  assign \g332070/_0_  = ~n24753 ;
  assign \g332071/_0_  = ~n24797 ;
  assign \g332672/_0_  = ~n24847 ;
  assign \g332673/_0_  = ~n24896 ;
  assign \g332678/_0_  = ~n24915 ;
  assign \g332679/_0_  = ~n24922 ;
  assign \g332680/_0_  = ~n24966 ;
  assign \g332681/_0_  = ~n25014 ;
  assign \g332682/_0_  = ~n25061 ;
  assign \g332700/_0_  = ~n25102 ;
  assign \g333449/_0_  = ~n25153 ;
  assign \g333453/_0_  = ~n25163 ;
  assign \g333454/_0_  = ~n25171 ;
  assign \g333462/_0_  = ~n25217 ;
  assign \g333463/_0_  = ~n25266 ;
  assign \g334369/_0_  = ~n25271 ;
  assign \g334370/_0_  = ~n25281 ;
  assign \g335243/_0_  = ~n25287 ;
  assign \g335244/_0_  = ~n25330 ;
  assign \g335965/_0_  = ~n25371 ;
  assign \g335969/_0_  = ~n25414 ;
  assign \g336538/_0_  = ~n25932 ;
  assign \g336539/_0_  = ~n25939 ;
  assign \g336540/_0_  = ~n26112 ;
  assign \g336546/_0_  = ~n26284 ;
  assign \g336551/_0_  = ~n26799 ;
  assign \g336552/_0_  = ~n26805 ;
  assign \g336557/_0_  = ~n27324 ;
  assign \g336558/_0_  = ~n27330 ;
  assign \g336654/_0_  = ~n27371 ;
  assign \g336655/_0_  = ~n27412 ;
  assign \g336656/_0_  = ~n27418 ;
  assign \g336657/_0_  = ~n27436 ;
  assign \g336660/_0_  = ~n27479 ;
  assign \g336850/_0_  = ~n27492 ;
  assign \g337247/_0_  = ~n27533 ;
  assign \g337248/_0_  = ~n27539 ;
  assign \g337249/_0_  = ~n27549 ;
  assign \g337250/_0_  = ~n27592 ;
  assign \g337251/_0_  = ~n27605 ;
  assign \g337629/_0_  = ~n27610 ;
  assign \g337635/_0_  = ~n27611 ;
  assign \g337637/_0_  = ~n27616 ;
  assign \g337879/_0_  = ~\P3_rd_reg/NET0131  ;
  assign \g337905/_0_  = ~n27629 ;
  assign \g337906/_0_  = ~n27646 ;
  assign \g337907/_0_  = ~n27665 ;
  assign \g337916/_0_  = ~n27679 ;
  assign \g337917/_0_  = ~n27684 ;
  assign \g337946/_0_  = ~n27725 ;
  assign \g337947/_0_  = ~n27730 ;
  assign \g337948/_0_  = ~n27740 ;
  assign \g337949/_0_  = ~n27745 ;
  assign \g337950/_0_  = ~n27786 ;
  assign \g338030/_0_  = ~n27787 ;
  assign \g338034/_0_  = ~n27789 ;
  assign \g338388/_0_  = ~n27795 ;
  assign \g338442/_0_  = ~n27846 ;
  assign \g338443/_0_  = ~n27886 ;
  assign \g338513/_0_  = ~n27892 ;
  assign \g338514/_0_  = ~n27897 ;
  assign \g338750/_0_  = ~n27976 ;
  assign \g338759/_0_  = ~n28054 ;
  assign \g338800/_0_  = ~n28083 ;
  assign \g338801/_0_  = ~n28106 ;
  assign \g338802/_0_  = ~n28129 ;
  assign \g338803/_0_  = ~n28150 ;
  assign \g338804/_0_  = ~n28170 ;
  assign \g338805/_0_  = ~n28191 ;
  assign \g338806/_0_  = ~n28213 ;
  assign \g338807/_0_  = ~n28235 ;
  assign \g338808/_0_  = ~n28257 ;
  assign \g338809/_0_  = ~n28279 ;
  assign \g338810/_0_  = ~n28301 ;
  assign \g338811/_0_  = ~n28323 ;
  assign \g338812/_0_  = ~n28344 ;
  assign \g338813/_0_  = ~n28364 ;
  assign \g338814/_0_  = ~n28384 ;
  assign \g338815/_0_  = ~n28413 ;
  assign \g338816/_0_  = ~n28436 ;
  assign \g338817/_0_  = ~n28459 ;
  assign \g338818/_0_  = ~n28480 ;
  assign \g338819/_0_  = ~n28500 ;
  assign \g338820/_0_  = ~n28521 ;
  assign \g338821/_0_  = ~n28543 ;
  assign \g338822/_0_  = ~n28565 ;
  assign \g338823/_0_  = ~n28587 ;
  assign \g338824/_0_  = ~n28609 ;
  assign \g338825/_0_  = ~n28631 ;
  assign \g338826/_0_  = ~n28653 ;
  assign \g338827/_0_  = ~n28674 ;
  assign \g338828/_0_  = ~n28694 ;
  assign \g338829/_0_  = ~n28714 ;
  assign \g338869/_0_  = ~n18658 ;
  assign \g338886/_0_  = ~n28721 ;
  assign \g338887/_0_  = ~n28727 ;
  assign \g338888/_0_  = ~n28739 ;
  assign \g339020/_0_  = ~n28817 ;
  assign \g339021/_0_  = ~n28855 ;
  assign \g339022/_0_  = ~n28877 ;
  assign \g339023/_0_  = ~n28899 ;
  assign \g339024/_0_  = ~n28921 ;
  assign \g339045/_0_  = ~n28945 ;
  assign \g339060/_0_  = ~n28969 ;
  assign \g339125/_0_  = ~n28991 ;
  assign \g339142/_0_  = ~n29007 ;
  assign \g339143/_0_  = ~n29023 ;
  assign \g339144/_0_  = ~n29039 ;
  assign \g339145/_0_  = ~n29055 ;
  assign \g339146/_0_  = ~n29071 ;
  assign \g339147/_0_  = ~n29087 ;
  assign \g339148/_0_  = ~n29103 ;
  assign \g339149/_0_  = ~n29119 ;
  assign \g339150/_0_  = ~n29135 ;
  assign \g339151/_0_  = ~n29151 ;
  assign \g339152/_0_  = ~n29167 ;
  assign \g339153/_0_  = ~n29183 ;
  assign \g339154/_0_  = ~n29199 ;
  assign \g339155/_0_  = ~n29215 ;
  assign \g339156/_0_  = ~n29231 ;
  assign \g339157/_0_  = ~n29247 ;
  assign \g339158/_0_  = ~n29263 ;
  assign \g339159/_0_  = ~n29279 ;
  assign \g339160/_0_  = ~n29295 ;
  assign \g339161/_0_  = ~n29311 ;
  assign \g339162/_0_  = ~n29327 ;
  assign \g339163/_0_  = ~n29343 ;
  assign \g339164/_0_  = ~n29359 ;
  assign \g339165/_0_  = ~n29375 ;
  assign \g339166/_0_  = ~n29391 ;
  assign \g339167/_0_  = ~n29407 ;
  assign \g339168/_0_  = ~n29423 ;
  assign \g339169/_0_  = ~n29439 ;
  assign \g339170/_0_  = ~n29455 ;
  assign \g339171/_0_  = ~n29471 ;
  assign \g339254/_0_  = ~n29512 ;
  assign \g339255/_0_  = ~n29522 ;
  assign \g339257/_0_  = ~n29567 ;
  assign \g339458/_0_  = ~n29589 ;
  assign \g339459/_0_  = ~n29619 ;
  assign \g339460/_0_  = ~n29649 ;
  assign \g339461/_0_  = ~n29679 ;
  assign \g339462/_0_  = ~n29709 ;
  assign \g339463/_0_  = ~n29739 ;
  assign \g339464/_0_  = ~n29761 ;
  assign \g339466/_0_  = ~n29783 ;
  assign \g339469/_0_  = ~n29805 ;
  assign \g339470/_0_  = ~n29827 ;
  assign \g339472/_0_  = ~n29829 ;
  assign \g339504/_0_  = ~n29857 ;
  assign \g339505/_0_  = ~n29885 ;
  assign \g339535/_0_  = ~n29913 ;
  assign \g339601/_0_  = ~n29922 ;
  assign \g339614/_0_  = ~n29941 ;
  assign \g339615/_0_  = ~n29960 ;
  assign \g339616/_0_  = ~n29979 ;
  assign \g339617/_0_  = ~n29998 ;
  assign \g339618/_0_  = ~n30017 ;
  assign \g339619/_0_  = ~n30036 ;
  assign \g339620/_0_  = ~n30055 ;
  assign \g339621/_0_  = ~n30074 ;
  assign \g339622/_0_  = ~n30093 ;
  assign \g339623/_0_  = ~n30112 ;
  assign \g339624/_0_  = ~n30131 ;
  assign \g339625/_0_  = ~n30150 ;
  assign \g339626/_0_  = ~n30169 ;
  assign \g339627/_0_  = ~n30188 ;
  assign \g339628/_0_  = ~n30207 ;
  assign \g339629/_0_  = ~n30226 ;
  assign \g339630/_0_  = ~n30245 ;
  assign \g339631/_0_  = ~n30264 ;
  assign \g339632/_0_  = ~n30283 ;
  assign \g339633/_0_  = ~n30302 ;
  assign \g339634/_0_  = ~n30321 ;
  assign \g339635/_0_  = ~n30340 ;
  assign \g339636/_0_  = ~n30359 ;
  assign \g339637/_0_  = ~n30378 ;
  assign \g339638/_0_  = ~n30397 ;
  assign \g339639/_0_  = ~n30416 ;
  assign \g339640/_0_  = ~n30435 ;
  assign \g339641/_0_  = ~n30454 ;
  assign \g339642/_0_  = ~n30473 ;
  assign \g339643/_0_  = ~n30492 ;
  assign \g339644/_0_  = ~n30511 ;
  assign \g339645/_0_  = ~n30530 ;
  assign \g339646/_0_  = ~n30549 ;
  assign \g339647/_0_  = ~n30568 ;
  assign \g339648/_0_  = ~n30587 ;
  assign \g339649/_0_  = ~n30606 ;
  assign \g339650/_0_  = ~n30625 ;
  assign \g339651/_0_  = ~n30644 ;
  assign \g339652/_0_  = ~n30663 ;
  assign \g339653/_0_  = ~n30682 ;
  assign \g339654/_0_  = ~n30701 ;
  assign \g339655/_0_  = ~n30720 ;
  assign \g339656/_0_  = ~n30739 ;
  assign \g339657/_0_  = ~n30758 ;
  assign \g339658/_0_  = ~n30777 ;
  assign \g339718/_0_  = ~n31491 ;
  assign \g339719/_0_  = ~n32176 ;
  assign \g339720/_0_  = ~n32863 ;
  assign \g339721/_0_  = ~n33513 ;
  assign \g339723/_0_  = ~n34167 ;
  assign \g339725/_0_  = ~n34177 ;
  assign \g339727/_0_  = ~n34189 ;
  assign \g340058/_0_  = ~n18663 ;
  assign \g340102/_0_  = ~n34226 ;
  assign \g340103/_0_  = ~n34260 ;
  assign \g340104/_0_  = ~n34312 ;
  assign \g340106/_0_  = ~n34371 ;
  assign \g340109/_0_  = ~n34404 ;
  assign \g340244/_0_  = ~n34414 ;
  assign \g340245/_0_  = ~n34423 ;
  assign \g340246/_0_  = ~n34433 ;
  assign \g340247/_0_  = ~n34446 ;
  assign \g340464/_0_  = ~n34474 ;
  assign \g340505/_0_  = ~n34502 ;
  assign \g340612/_0_  = ~n34521 ;
  assign \g340613/_0_  = ~n34540 ;
  assign \g340614/_0_  = ~n34559 ;
  assign \g340615/_0_  = ~n34578 ;
  assign \g340616/_0_  = ~n34597 ;
  assign \g340617/_0_  = ~n34616 ;
  assign \g340618/_0_  = ~n34635 ;
  assign \g340619/_0_  = ~n34654 ;
  assign \g340620/_0_  = ~n34673 ;
  assign \g340621/_0_  = ~n34692 ;
  assign \g340622/_0_  = ~n34711 ;
  assign \g340623/_0_  = ~n34730 ;
  assign \g340624/_0_  = ~n34749 ;
  assign \g340625/_0_  = ~n34768 ;
  assign \g340626/_0_  = ~n34787 ;
  assign \g340630/_0_  = ~n34806 ;
  assign \g340631/_0_  = ~n34825 ;
  assign \g340632/_0_  = ~n34844 ;
  assign \g340633/_0_  = ~n34863 ;
  assign \g340634/_0_  = ~n34882 ;
  assign \g340635/_0_  = ~n34901 ;
  assign \g340636/_0_  = ~n34920 ;
  assign \g340637/_0_  = ~n34939 ;
  assign \g340638/_0_  = ~n34958 ;
  assign \g340640/_0_  = ~n34977 ;
  assign \g340641/_0_  = ~n34996 ;
  assign \g340642/_0_  = ~n35015 ;
  assign \g340643/_0_  = ~n35034 ;
  assign \g340644/_0_  = ~n35053 ;
  assign \g340645/_0_  = ~n35072 ;
  assign \g340701/_0_  = ~n35105 ;
  assign \g340702/_0_  = ~n35142 ;
  assign \g340703/_0_  = ~n35198 ;
  assign \g340704/_0_  = ~n35248 ;
  assign \g340714/_0_  = ~n35279 ;
  assign \g340716/_0_  = ~n35310 ;
  assign \g340717/_0_  = ~n35345 ;
  assign \g340718/_0_  = ~n35399 ;
  assign \g340728/_0_  = ~n35435 ;
  assign \g340729/_0_  = ~n35478 ;
  assign \g340730/_0_  = ~n35511 ;
  assign \g340731/_0_  = ~n35544 ;
  assign \g340747/_0_  = ~n35598 ;
  assign \g340748/_0_  = ~n35635 ;
  assign \g340749/_0_  = ~n35684 ;
  assign \g340750/_0_  = ~n35716 ;
  assign \g340751/_0_  = ~n35758 ;
  assign \g340752/_0_  = ~n35797 ;
  assign \g340753/_0_  = ~n35856 ;
  assign \g340754/_0_  = ~n35889 ;
  assign \g340792/_0_  = ~n35899 ;
  assign \g340793/_0_  = ~n35909 ;
  assign \g340794/_0_  = ~n35920 ;
  assign \g340795/_0_  = ~n35934 ;
  assign \g340796/_0_  = ~n35948 ;
  assign \g340797/_0_  = ~n35960 ;
  assign \g340988/_0_  = ~n35988 ;
  assign \g341033/_0_  = ~n36016 ;
  assign \g341191/_0_  = ~n36035 ;
  assign \g341192/_0_  = ~n36054 ;
  assign \g341193/_0_  = ~n36073 ;
  assign \g341194/_0_  = ~n36092 ;
  assign \g341195/_0_  = ~n36111 ;
  assign \g341196/_0_  = ~n36130 ;
  assign \g341197/_0_  = ~n36149 ;
  assign \g341198/_0_  = ~n36168 ;
  assign \g341199/_0_  = ~n36187 ;
  assign \g341200/_0_  = ~n36206 ;
  assign \g341201/_0_  = ~n36225 ;
  assign \g341202/_0_  = ~n36244 ;
  assign \g341203/_0_  = ~n36263 ;
  assign \g341205/_0_  = ~n36282 ;
  assign \g341206/_0_  = ~n36301 ;
  assign \g341207/_0_  = ~n36320 ;
  assign \g341208/_0_  = ~n36339 ;
  assign \g341209/_0_  = ~n36358 ;
  assign \g341210/_0_  = ~n36377 ;
  assign \g341211/_0_  = ~n36396 ;
  assign \g341212/_0_  = ~n36415 ;
  assign \g341213/_0_  = ~n36434 ;
  assign \g341214/_0_  = ~n36453 ;
  assign \g341215/_0_  = ~n36472 ;
  assign \g341216/_0_  = ~n36491 ;
  assign \g341217/_0_  = ~n36510 ;
  assign \g341218/_0_  = ~n36529 ;
  assign \g341219/_0_  = ~n36548 ;
  assign \g341220/_0_  = ~n36567 ;
  assign \g341221/_0_  = ~n36586 ;
  assign \g341241/_0_  = ~n36639 ;
  assign \g341242/_0_  = ~n36692 ;
  assign \g341245/_0_  = ~n36748 ;
  assign \g341248/_0_  = ~n36801 ;
  assign \g341250/_0_  = ~n36821 ;
  assign \g341251/_0_  = ~n36878 ;
  assign \g341339/_0_  = ~n36916 ;
  assign \g341347/_0_  = ~n36954 ;
  assign \g341349/_0_  = ~n36993 ;
  assign \g341350/_0_  = ~n37024 ;
  assign \g341352/_0_  = ~n37052 ;
  assign \g341353/_0_  = ~n37082 ;
  assign \g341354/_0_  = ~n37113 ;
  assign \g341365/_0_  = ~n37142 ;
  assign \g341366/_0_  = ~n37181 ;
  assign \g341367/_0_  = ~n37219 ;
  assign \g341368/_0_  = ~n37253 ;
  assign \g341369/_0_  = ~n37284 ;
  assign \g341370/_0_  = ~n37316 ;
  assign \g341373/_0_  = ~n37346 ;
  assign \g341388/_0_  = ~n37375 ;
  assign \g341389/_0_  = ~n37419 ;
  assign \g341390/_0_  = ~n37450 ;
  assign \g341391/_0_  = ~n37484 ;
  assign \g341392/_0_  = ~n37512 ;
  assign \g341393/_0_  = ~n37544 ;
  assign \g341394/_0_  = ~n37572 ;
  assign \g341395/_0_  = ~n37616 ;
  assign \g341396/_0_  = ~n37646 ;
  assign \g341397/_0_  = ~n37677 ;
  assign \g341398/_0_  = ~n37705 ;
  assign \g341400/_0_  = ~n37734 ;
  assign \g341401/_0_  = ~n37770 ;
  assign \g341419/_0_  = ~n37807 ;
  assign \g341435/_0_  = ~n37846 ;
  assign \g341436/_0_  = ~n37877 ;
  assign \g341455/_0_  = ~n37883 ;
  assign \g341456/_0_  = ~n37889 ;
  assign \g341457/_0_  = ~n37898 ;
  assign \g341458/_0_  = ~n37907 ;
  assign \g342136/_0_  = ~n37929 ;
  assign \g342137/_0_  = ~n37948 ;
  assign \g342141/_0_  = ~n37966 ;
  assign \g342145/_0_  = ~n37990 ;
  assign \g342148/_0_  = ~n38006 ;
  assign \g342149/_0_  = ~n38024 ;
  assign \g342308/_0_  = ~n38052 ;
  assign \g342318/_0_  = ~n38085 ;
  assign \g342322/_0_  = ~n38115 ;
  assign \g342323/_0_  = ~n38146 ;
  assign \g342327/_0_  = ~n38175 ;
  assign \g342331/_0_  = ~n38203 ;
  assign \g342333/_0_  = ~n38231 ;
  assign \g342354/_0_  = ~n38268 ;
  assign \g342355/_0_  = ~n38309 ;
  assign \g342356/_0_  = ~n38342 ;
  assign \g342357/_0_  = ~n38377 ;
  assign \g342358/_0_  = ~n38412 ;
  assign \g342359/_0_  = ~n38442 ;
  assign \g342383/_0_  = ~n38484 ;
  assign \g342384/_0_  = ~n38518 ;
  assign \g342385/_0_  = ~n38551 ;
  assign \g342386/_0_  = ~n38584 ;
  assign \g342387/_0_  = ~n38615 ;
  assign \g342388/_0_  = ~n38648 ;
  assign \g342389/_0_  = ~n38678 ;
  assign \g342390/_0_  = ~n38721 ;
  assign \g342391/_0_  = ~n38749 ;
  assign \g342392/_0_  = ~n38783 ;
  assign \g342393/_0_  = ~n38816 ;
  assign \g342394/_0_  = ~n38846 ;
  assign \g342397/_0_  = ~n38887 ;
  assign \g342398/_0_  = ~n38922 ;
  assign \g342399/_0_  = ~n38960 ;
  assign \g342400/_0_  = ~n38991 ;
  assign \g342401/_0_  = ~n39019 ;
  assign \g342454/u3_syn_4  = n39020 ;
  assign \g342800/_0_  = ~n39048 ;
  assign \g343406/_0_  = ~n39067 ;
  assign \g343407/_0_  = ~n39086 ;
  assign \g343408/_0_  = ~n39105 ;
  assign \g343409/_0_  = ~n39124 ;
  assign \g343410/_0_  = ~n39143 ;
  assign \g343411/_0_  = ~n39162 ;
  assign \g343412/_0_  = ~n39181 ;
  assign \g343413/_0_  = ~n39200 ;
  assign \g343414/_0_  = ~n39219 ;
  assign \g343415/_0_  = ~n39238 ;
  assign \g343416/_0_  = ~n39257 ;
  assign \g343417/_0_  = ~n39276 ;
  assign \g343418/_0_  = ~n39295 ;
  assign \g343419/_0_  = ~n39314 ;
  assign \g343420/_0_  = ~n39333 ;
  assign \g343431/_0_  = ~n39357 ;
  assign \g343432/_0_  = ~n39381 ;
  assign \g343433/_0_  = ~n39404 ;
  assign \g343434/_0_  = ~n39424 ;
  assign \g343435/_0_  = ~n39443 ;
  assign \g343436/_0_  = ~n39466 ;
  assign \g343437/_0_  = ~n39489 ;
  assign \g343439/_0_  = ~n39509 ;
  assign \g343440/_0_  = ~n39528 ;
  assign \g343441/_0_  = ~n39546 ;
  assign \g343443/_0_  = ~n39568 ;
  assign \g343444/_0_  = ~n39591 ;
  assign \g343445/_0_  = ~n39610 ;
  assign \g343446/_0_  = ~n39628 ;
  assign \g343447/_0_  = ~n39646 ;
  assign \g343452/_0_  = ~n39671 ;
  assign \g343453/_0_  = ~n39691 ;
  assign \g343454/_0_  = ~n39712 ;
  assign \g343455/_0_  = ~n39730 ;
  assign \g343456/_0_  = ~n39748 ;
  assign \g343458/_0_  = ~n39762 ;
  assign \g343459/_0_  = ~n39779 ;
  assign \g343460/_0_  = ~n39796 ;
  assign \g343461/_0_  = ~n39812 ;
  assign \g343462/_0_  = ~n39828 ;
  assign \g343463/_0_  = ~n39855 ;
  assign \g343464/_0_  = ~n39881 ;
  assign \g343465/_0_  = ~n39900 ;
  assign \g343466/_0_  = ~n39916 ;
  assign \g343467/_0_  = ~n39934 ;
  assign \g343512/_0_  = ~n39962 ;
  assign \g343514/_0_  = ~n39996 ;
  assign \g343515/_0_  = ~n40024 ;
  assign \g343517/_0_  = ~n40052 ;
  assign \g343524/_0_  = ~n40083 ;
  assign \g343531/_0_  = ~n40111 ;
  assign \g343533/_0_  = ~n40139 ;
  assign \g343534/_0_  = ~n40173 ;
  assign \g343535/_0_  = ~n40201 ;
  assign \g343536/_0_  = ~n40238 ;
  assign \g343537/_0_  = ~n40275 ;
  assign \g343555/_0_  = ~n40306 ;
  assign \g343556/_0_  = ~n40338 ;
  assign \g343557/_0_  = ~n40367 ;
  assign \g343558/_0_  = ~n40395 ;
  assign \g343559/_0_  = ~n40427 ;
  assign \g343560/_0_  = ~n40455 ;
  assign \g343561/_0_  = ~n40489 ;
  assign \g343563/_0_  = ~n40517 ;
  assign \g343564/_0_  = ~n40555 ;
  assign \g343566/_0_  = ~n40593 ;
  assign \g343567/_0_  = ~n40628 ;
  assign \g343568/_0_  = ~n40658 ;
  assign \g343569/_0_  = ~n40689 ;
  assign \g343570/_0_  = ~n40721 ;
  assign \g343699/_0_  = ~n40731 ;
  assign \g343703/_0_  = ~n40743 ;
  assign \g343944/_0_  = ~n40771 ;
  assign \g343992/_0_  = ~n40799 ;
  assign \g344429/_0_  = ~n40818 ;
  assign \g344430/_0_  = ~n40837 ;
  assign \g344431/_0_  = ~n40856 ;
  assign \g344432/_0_  = ~n40875 ;
  assign \g344433/_0_  = ~n40894 ;
  assign \g344434/_0_  = ~n40913 ;
  assign \g344435/_0_  = ~n40932 ;
  assign \g344437/_0_  = ~n40951 ;
  assign \g344438/_0_  = ~n40970 ;
  assign \g344439/_0_  = ~n40989 ;
  assign \g344440/_0_  = ~n41008 ;
  assign \g344441/_0_  = ~n41027 ;
  assign \g344442/_0_  = ~n41046 ;
  assign \g344443/_0_  = ~n41065 ;
  assign \g344444/_0_  = ~n41084 ;
  assign \g344447/_0_  = ~n41103 ;
  assign \g344448/_0_  = ~n41122 ;
  assign \g344449/_0_  = ~n41141 ;
  assign \g344450/_0_  = ~n41160 ;
  assign \g344451/_0_  = ~n41179 ;
  assign \g344452/_0_  = ~n41198 ;
  assign \g344453/_0_  = ~n41217 ;
  assign \g344454/_0_  = ~n41236 ;
  assign \g344455/_0_  = ~n41255 ;
  assign \g344456/_0_  = ~n41274 ;
  assign \g344457/_0_  = ~n41293 ;
  assign \g344458/_0_  = ~n41312 ;
  assign \g344459/_0_  = ~n41331 ;
  assign \g344460/_0_  = ~n41350 ;
  assign \g344461/_0_  = ~n41369 ;
  assign \g344495/_0_  = ~n41392 ;
  assign \g344496/_0_  = ~n41412 ;
  assign \g344497/_0_  = ~n41433 ;
  assign \g344498/_0_  = ~n41449 ;
  assign \g344499/_0_  = ~n41465 ;
  assign \g344500/_0_  = ~n41482 ;
  assign \g344501/_0_  = ~n41500 ;
  assign \g344502/_0_  = ~n41519 ;
  assign \g344503/_0_  = ~n41539 ;
  assign \g344504/_0_  = ~n41565 ;
  assign \g344505/_0_  = ~n41584 ;
  assign \g344506/_0_  = ~n41603 ;
  assign \g344507/_0_  = ~n41622 ;
  assign \g344508/_0_  = ~n41656 ;
  assign \g344511/_0_  = ~n41677 ;
  assign \g344512/_0_  = ~n41698 ;
  assign \g344513/_0_  = ~n41722 ;
  assign \g344514/_0_  = ~n41742 ;
  assign \g344515/_0_  = ~n41761 ;
  assign \g344516/_0_  = ~n41782 ;
  assign \g344517/_0_  = ~n41802 ;
  assign \g344523/_0_  = ~n41825 ;
  assign \g344524/_0_  = ~n41846 ;
  assign \g344525/_0_  = ~n41867 ;
  assign \g344526/_0_  = ~n41887 ;
  assign \g344527/_0_  = ~n41906 ;
  assign \g344528/_0_  = ~n41923 ;
  assign \g344529/_0_  = ~n41941 ;
  assign \g344536/_0_  = ~n41957 ;
  assign \g344537/_0_  = ~n41976 ;
  assign \g344538/_0_  = ~n41992 ;
  assign \g344539/_0_  = ~n42011 ;
  assign \g344540/_0_  = ~n42030 ;
  assign \g344541/_0_  = ~n42046 ;
  assign \g344542/_0_  = ~n42061 ;
  assign \g344543/_0_  = ~n42079 ;
  assign \g344545/_0_  = ~n42098 ;
  assign \g344546/_0_  = ~n42122 ;
  assign \g344547/_0_  = ~n42139 ;
  assign \g344548/_0_  = ~n42158 ;
  assign \g344549/_0_  = ~n42178 ;
  assign \g344550/_0_  = ~n42199 ;
  assign \g344711/_0_  = ~n42226 ;
  assign \g344712/_0_  = ~n42258 ;
  assign \g344729/_0_  = ~n42292 ;
  assign \g344737/_0_  = ~n42319 ;
  assign \g344738/_0_  = ~n42351 ;
  assign \g344783/_0_  = ~n42378 ;
  assign \g344784/_0_  = ~n42414 ;
  assign \g344786/_0_  = ~n42441 ;
  assign \g344791/_0_  = ~n42481 ;
  assign \g344792/_0_  = ~n42513 ;
  assign \g344816/_0_  = ~n42523 ;
  assign \g344819/_0_  = ~n42537 ;
  assign \g344823/_0_  = ~n42874 ;
  assign \g344825/_0_  = ~n43214 ;
  assign \g345116/_0_  = ~n43226 ;
  assign \g345129/_0_  = ~n43239 ;
  assign \g345149/_0_  = ~n43252 ;
  assign \g345161/_0_  = ~n43266 ;
  assign \g345170/_0_  = ~n43280 ;
  assign \g345237/_0_  = ~n43292 ;
  assign \g345313/_0_  = ~n43311 ;
  assign \g345314/_0_  = ~n43329 ;
  assign \g345316/_0_  = ~n43349 ;
  assign \g345317/_0_  = ~n43366 ;
  assign \g345318/_0_  = ~n43384 ;
  assign \g345319/_0_  = ~n43403 ;
  assign \g345320/_0_  = ~n43421 ;
  assign \g345321/_0_  = ~n43442 ;
  assign \g345322/_0_  = ~n43463 ;
  assign \g345323/_0_  = ~n43481 ;
  assign \g345324/_0_  = ~n43499 ;
  assign \g345325/_0_  = ~n43516 ;
  assign \g345326/_0_  = ~n43540 ;
  assign \g345327/_0_  = ~n43558 ;
  assign \g345328/_0_  = ~n43576 ;
  assign \g345329/_0_  = ~n43596 ;
  assign \g345333/_0_  = ~n43614 ;
  assign \g345334/_0_  = ~n43635 ;
  assign \g345335/_0_  = ~n43653 ;
  assign \g345336/_0_  = ~n43671 ;
  assign \g345337/_0_  = ~n43689 ;
  assign \g345338/_0_  = ~n43707 ;
  assign \g345339/_0_  = ~n43724 ;
  assign \g345340/_0_  = ~n43746 ;
  assign \g345349/_0_  = ~n43764 ;
  assign \g345350/_0_  = ~n43785 ;
  assign \g345351/_0_  = ~n43802 ;
  assign \g345352/_0_  = ~n43820 ;
  assign \g345353/_0_  = ~n43838 ;
  assign \g345354/_0_  = ~n43856 ;
  assign \g345355/_0_  = ~n43874 ;
  assign \g345356/_0_  = ~n43890 ;
  assign \g345365/_0_  = ~n43909 ;
  assign \g345366/_0_  = ~n43926 ;
  assign \g345367/_0_  = ~n43945 ;
  assign \g345368/_0_  = ~n43961 ;
  assign \g345369/_0_  = ~n43977 ;
  assign \g345370/_0_  = ~n43991 ;
  assign \g345371/_0_  = ~n44007 ;
  assign \g345373/_0_  = ~n44023 ;
  assign \g345374/_0_  = ~n44046 ;
  assign \g345377/_0_  = ~n44063 ;
  assign \g345378/_0_  = ~n44082 ;
  assign \g345379/_0_  = ~n44102 ;
  assign \g345380/_0_  = ~n44120 ;
  assign \g345381/_0_  = ~n44137 ;
  assign \g345382/_0_  = ~n44155 ;
  assign \g345383/_0_  = ~n44177 ;
  assign \g345488/_0_  = ~n44206 ;
  assign \g345491/_0_  = ~n44233 ;
  assign \g345524/_0_  = ~n44260 ;
  assign \g345525/_0_  = ~n44287 ;
  assign \g345545/_0_  = ~n44314 ;
  assign \g345546/_0_  = ~n44348 ;
  assign \g345574/_0_  = ~n44384 ;
  assign \g345575/_0_  = ~n44411 ;
  assign \g345638/_0_  = ~n44445 ;
  assign \g345639/_0_  = ~n44479 ;
  assign \g345690/_0_  = ~n44485 ;
  assign \g345691/_0_  = ~n44497 ;
  assign \g345692/_0_  = ~n44506 ;
  assign \g345694/_0_  = ~n44755 ;
  assign \g345695/_0_  = ~n44764 ;
  assign \g345698/_0_  = ~n44776 ;
  assign \g345699/_0_  = ~n44788 ;
  assign \g345701/_0_  = ~n44809 ;
  assign \g345703/_0_  = ~n44833 ;
  assign \g346299/_0_  = ~n16244 ;
  assign \g346326/_0_  = ~n15782 ;
  assign \g346364/_0_  = ~n16302 ;
  assign \g346707/_0_  = ~n44845 ;
  assign \g346711/_0_  = ~n44857 ;
  assign \g346721/_0_  = ~n44878 ;
  assign \g346726/_0_  = ~n44890 ;
  assign \g346729/_0_  = ~n44910 ;
  assign \g346730/_0_  = ~n44929 ;
  assign \g346731/_0_  = ~n44950 ;
  assign \g346733/_0_  = ~n44968 ;
  assign \g346735/_0_  = ~n44986 ;
  assign \g346738/_0_  = ~n45006 ;
  assign \g346740/_0_  = ~n45024 ;
  assign \g346741/_0_  = ~n45042 ;
  assign \g346746/_0_  = ~n45058 ;
  assign \g346748/_0_  = ~n45078 ;
  assign \g346750/_0_  = ~n45101 ;
  assign \g346751/_0_  = ~n45120 ;
  assign \g346758/_0_  = ~n45132 ;
  assign \g346759/_0_  = ~n45151 ;
  assign \g346761/_0_  = ~n45167 ;
  assign \g346762/_0_  = ~n45185 ;
  assign \g346763/_0_  = ~n45204 ;
  assign \g346765/_0_  = ~n45225 ;
  assign \g346766/_0_  = ~n45243 ;
  assign \g346965/_0_  = ~n45252 ;
  assign \g346971/_0_  = ~n45271 ;
  assign \g346981/_0_  = ~n45307 ;
  assign \g346986/_0_  = ~n45349 ;
  assign \g346988/_0_  = ~n45392 ;
  assign \g346989/_0_  = ~n45426 ;
  assign \g346994/_0_  = ~n45435 ;
  assign \g346998/_0_  = ~n45469 ;
  assign \g347015/_0_  = ~n45488 ;
  assign \g347016/_0_  = ~n45532 ;
  assign \g347017/_0_  = ~n45568 ;
  assign \g347018/_0_  = ~n45613 ;
  assign \g347019/_0_  = ~n45640 ;
  assign \g347020/_0_  = ~n45649 ;
  assign \g347043/_0_  = ~n45671 ;
  assign \g347050/_0_  = ~n45694 ;
  assign \g347051/_0_  = ~n45712 ;
  assign \g347052/_0_  = ~n45750 ;
  assign \g347053/_0_  = ~n45789 ;
  assign \g347054/_0_  = ~n45836 ;
  assign \g347055/_0_  = ~n45868 ;
  assign \g347056/_0_  = ~n45877 ;
  assign \g347057/_0_  = ~n45906 ;
  assign \g347058/_0_  = ~n45915 ;
  assign \g347059/_0_  = ~n45954 ;
  assign \g347061/_0_  = ~n45972 ;
  assign \g347062/_0_  = ~n46008 ;
  assign \g347063/_0_  = ~n46046 ;
  assign \g347064/_0_  = ~n46085 ;
  assign \g347065/_0_  = ~n46125 ;
  assign \g347066/_0_  = ~n46164 ;
  assign \g347067/_0_  = ~n46174 ;
  assign \g347068/_0_  = ~n46184 ;
  assign \g347069/_0_  = ~n46194 ;
  assign \g347070/_0_  = ~n46204 ;
  assign \g347071/_0_  = ~n46214 ;
  assign \g347083/_0_  = ~n46224 ;
  assign \g347085/_0_  = ~n46264 ;
  assign \g347087/_0_  = ~n46278 ;
  assign \g347089/_0_  = ~n46401 ;
  assign \g347090/_0_  = ~n46415 ;
  assign \g347091/_0_  = ~n46454 ;
  assign \g347092/_0_  = ~n46468 ;
  assign \g347093/_0_  = ~n46478 ;
  assign \g347096/_0_  = ~n46516 ;
  assign \g347097/_0_  = ~n46530 ;
  assign \g347098/_0_  = ~n46571 ;
  assign \g347099/_0_  = ~n46585 ;
  assign \g347100/_0_  = ~n46613 ;
  assign \g347101/_0_  = ~n46652 ;
  assign \g347102/_0_  = ~n46666 ;
  assign \g347104/_0_  = ~n46693 ;
  assign \g347106/_0_  = ~n46732 ;
  assign \g347108/_0_  = ~n46746 ;
  assign \g347318/_0_  = ~n46774 ;
  assign \g347400/_0_  = ~n46802 ;
  assign \g347449/_0_  = ~n15832 ;
  assign \g347477/_0_  = ~n15949 ;
  assign \g347488/_0_  = ~n16061 ;
  assign \g347531/_0_  = ~n15936 ;
  assign \g347537/_0_  = ~n15922 ;
  assign \g347544/_0_  = ~n15909 ;
  assign \g347546/_0_  = ~n15895 ;
  assign \g347553/_0_  = ~n15844 ;
  assign \g347560/_0_  = ~n15820 ;
  assign \g347569/_0_  = ~n16110 ;
  assign \g347575/_0_  = ~n16095 ;
  assign \g347581/_1_  = ~n16083 ;
  assign \g347587/_0_  = ~n16071 ;
  assign \g347592/_0_  = ~n15976 ;
  assign \g347597/_0_  = ~n15963 ;
  assign \g347603/_0_  = ~n16188 ;
  assign \g347610/_0_  = ~n16175 ;
  assign \g347611/_0_  = ~n16006 ;
  assign \g347616/_0_  = ~n15991 ;
  assign \g347624/_0_  = ~n16035 ;
  assign \g347628/_1_  = ~n16021 ;
  assign \g347632/_0_  = ~n16048 ;
  assign \g347641/_0_  = ~n16131 ;
  assign \g347645/_0_  = ~n16147 ;
  assign \g347653/_0_  = ~n15794 ;
  assign \g347661/_0_  = ~n15872 ;
  assign \g347671/_0_  = ~n15856 ;
  assign \g347678/_0_  = ~n15884 ;
  assign \g347881/_0_  = ~n46821 ;
  assign \g347883/_0_  = ~n46840 ;
  assign \g347885/_0_  = ~n46859 ;
  assign \g347886/_0_  = ~n46878 ;
  assign \g347888/_0_  = ~n46897 ;
  assign \g347889/_0_  = ~n46916 ;
  assign \g347890/_0_  = ~n46935 ;
  assign \g347891/_0_  = ~n46954 ;
  assign \g347892/_0_  = ~n46973 ;
  assign \g347893/_0_  = ~n46992 ;
  assign \g347895/_0_  = ~n47011 ;
  assign \g347896/_0_  = ~n47030 ;
  assign \g347897/_0_  = ~n47049 ;
  assign \g347898/_0_  = ~n47068 ;
  assign \g347899/_0_  = ~n47087 ;
  assign \g347902/_0_  = ~n47106 ;
  assign \g347903/_0_  = ~n47125 ;
  assign \g347904/_0_  = ~n47144 ;
  assign \g347906/_0_  = ~n47163 ;
  assign \g347907/_0_  = ~n47182 ;
  assign \g347908/_0_  = ~n47201 ;
  assign \g347909/_0_  = ~n47220 ;
  assign \g347910/_0_  = ~n47239 ;
  assign \g347911/_0_  = ~n47258 ;
  assign \g347912/_0_  = ~n47277 ;
  assign \g347913/_0_  = ~n47296 ;
  assign \g347914/_0_  = ~n47315 ;
  assign \g347915/_0_  = ~n47334 ;
  assign \g347916/_0_  = ~n47353 ;
  assign \g347917/_0_  = ~n47372 ;
  assign \g347974/_0_  = ~n47393 ;
  assign \g347977/_0_  = ~n47416 ;
  assign \g347983/_0_  = ~n47439 ;
  assign \g347999/_0_  = ~n47460 ;
  assign \g348012/_0_  = ~n47476 ;
  assign \g348015/_0_  = ~n47500 ;
  assign \g348288/_0_  = ~n47510 ;
  assign \g348291/_0_  = ~n47520 ;
  assign \g348292/_0_  = ~n47526 ;
  assign \g348293/_0_  = ~n47576 ;
  assign \g348294/_0_  = ~n47601 ;
  assign \g348295/_0_  = ~n47611 ;
  assign \g348296/_0_  = ~n47620 ;
  assign \g348300/_0_  = ~n47630 ;
  assign \g348301/_0_  = ~n47640 ;
  assign \g348302/_0_  = ~n47690 ;
  assign \g348303/_0_  = ~n47708 ;
  assign \g348304/_0_  = ~n47718 ;
  assign \g348307/_0_  = ~n47744 ;
  assign \g348308/_0_  = ~n47785 ;
  assign \g349018/_0_  = ~n47803 ;
  assign \g349020/_0_  = ~n47825 ;
  assign \g349021/_0_  = ~n47843 ;
  assign \g349025/_0_  = ~n47866 ;
  assign \g349026/_0_  = ~n47885 ;
  assign \g349027/_0_  = ~n47903 ;
  assign \g349035/_0_  = ~n47926 ;
  assign \g349036/_0_  = ~n47945 ;
  assign \g349037/_0_  = ~n47963 ;
  assign \g349049/_0_  = ~n47981 ;
  assign \g349050/_0_  = ~n48002 ;
  assign \g349051/_0_  = ~n48021 ;
  assign \g349070/_0_  = ~n48037 ;
  assign \g349071/_0_  = ~n48054 ;
  assign \g349072/_0_  = ~n48071 ;
  assign \g349076/_0_  = ~n48094 ;
  assign \g349077/_0_  = ~n48113 ;
  assign \g349078/_0_  = ~n48133 ;
  assign \g349326/_0_  = ~n48146 ;
  assign \g349333/_0_  = ~n48197 ;
  assign \g349334/_0_  = ~n48221 ;
  assign \g349335/_0_  = ~n48231 ;
  assign \g349343/_0_  = ~n48241 ;
  assign \g349345/_0_  = ~n48253 ;
  assign \g349349/_0_  = ~n48273 ;
  assign \g349350/_0_  = ~n48283 ;
  assign \g349355/_0_  = ~n48332 ;
  assign \g349357/_0_  = ~n48356 ;
  assign \g349358/_0_  = ~n48369 ;
  assign \g349873/_0_  = ~n48469 ;
  assign \g350037/_0_  = ~n48482 ;
  assign \g350042/_0_  = ~n48490 ;
  assign \g350050/_0_  = ~n48511 ;
  assign \g350051/_0_  = ~n48522 ;
  assign \g350089/_0_  = ~n48543 ;
  assign \g350090/_0_  = ~n48551 ;
  assign \g350093/_0_  = ~n48569 ;
  assign \g350094/_0_  = ~n48580 ;
  assign \g350096/_0_  = ~n48597 ;
  assign \g350097/_0_  = ~n48608 ;
  assign \g350165/_0_  = ~n48618 ;
  assign \g350166/_0_  = ~n48628 ;
  assign \g350168/_0_  = ~n48638 ;
  assign \g350170/_0_  = ~n48645 ;
  assign \g350171/_0_  = ~n48655 ;
  assign \g350172/_0_  = ~n48667 ;
  assign \g350173/_0_  = ~n48710 ;
  assign \g350174/_0_  = ~n48751 ;
  assign \g350175/_0_  = ~n48797 ;
  assign \g350176/_0_  = ~n48841 ;
  assign \g350177/_0_  = ~n48886 ;
  assign \g350178/_0_  = ~n48897 ;
  assign \g350179/_0_  = ~n48942 ;
  assign \g350180/_0_  = ~n48987 ;
  assign \g350181/_0_  = ~n48997 ;
  assign \g350183/_0_  = ~n49007 ;
  assign \g350184/_0_  = ~n49019 ;
  assign \g350185/_0_  = ~n49029 ;
  assign \g350186/_0_  = ~n49037 ;
  assign \g350187/_0_  = ~n49080 ;
  assign \g350188/_0_  = ~n49125 ;
  assign \g350189/_0_  = ~n49168 ;
  assign \g350190/_0_  = ~n49214 ;
  assign \g350191/_0_  = ~n49260 ;
  assign \g350192/_0_  = ~n49305 ;
  assign \g350193/_0_  = ~n49315 ;
  assign \g350194/_0_  = ~n49356 ;
  assign \g350195/_0_  = ~n49397 ;
  assign \g350196/_0_  = ~n49407 ;
  assign \g350197/_0_  = ~n49450 ;
  assign \g350198/_0_  = ~n49492 ;
  assign \g350199/_0_  = ~n49538 ;
  assign \g350200/_0_  = ~n49582 ;
  assign \g350201/_0_  = ~n49625 ;
  assign \g350202/_0_  = ~n49638 ;
  assign \g350203/_0_  = ~n49644 ;
  assign \g350204/_0_  = ~n49685 ;
  assign \g350205/_0_  = ~n49729 ;
  assign \g350654/_0_  = ~n49764 ;
  assign \g350655/_0_  = ~n49790 ;
  assign \g350656/_0_  = ~n49812 ;
  assign \g350658/_0_  = ~n49833 ;
  assign \g350660/_0_  = ~n49852 ;
  assign \g350661/_0_  = ~n49870 ;
  assign \g350662/_0_  = ~n49889 ;
  assign \g350663/_0_  = ~n49909 ;
  assign \g350664/_0_  = ~n49929 ;
  assign \g350665/_0_  = ~n49949 ;
  assign \g350666/_0_  = ~n49969 ;
  assign \g350667/_0_  = ~n49989 ;
  assign \g350668/_0_  = ~n50009 ;
  assign \g350669/_0_  = ~n50044 ;
  assign \g350670/_0_  = ~n50070 ;
  assign \g350671/_0_  = ~n50089 ;
  assign \g350672/_0_  = ~n50111 ;
  assign \g350673/_0_  = ~n50132 ;
  assign \g350674/_0_  = ~n50150 ;
  assign \g350675/_0_  = ~n50169 ;
  assign \g350676/_0_  = ~n50187 ;
  assign \g350677/_0_  = ~n50205 ;
  assign \g350678/_0_  = ~n50224 ;
  assign \g350679/_0_  = ~n50244 ;
  assign \g350680/_0_  = ~n50264 ;
  assign \g350681/_0_  = ~n50284 ;
  assign \g350682/_0_  = ~n50304 ;
  assign \g350683/_0_  = ~n50324 ;
  assign \g350684/_0_  = ~n50344 ;
  assign \g350685/_0_  = ~n50363 ;
  assign \g350686/_0_  = ~n50381 ;
  assign \g350687/_0_  = ~n50399 ;
  assign \g350723/_0_  = ~n50437 ;
  assign \g350724/_0_  = ~n50471 ;
  assign \g350725/_0_  = ~n50513 ;
  assign \g350726/_0_  = ~n50549 ;
  assign \g350727/_0_  = ~n50587 ;
  assign \g350728/_0_  = ~n50625 ;
  assign \g350729/_0_  = ~n50664 ;
  assign \g350730/_0_  = ~n50702 ;
  assign \g350731/_0_  = ~n50748 ;
  assign \g350814/_0_  = ~n50820 ;
  assign \g350815/_0_  = ~n50856 ;
  assign \g350816/_0_  = ~n50891 ;
  assign \g350817/_0_  = ~n50925 ;
  assign \g350818/_0_  = ~n50959 ;
  assign \g350819/_0_  = ~n51005 ;
  assign \g350820/_0_  = ~n51041 ;
  assign \g350821/_0_  = ~n51075 ;
  assign \g350822/_0_  = ~n51110 ;
  assign \g350823/_0_  = ~n51144 ;
  assign \g350824/_0_  = ~n51177 ;
  assign \g350825/_0_  = ~n51226 ;
  assign \g350826/_0_  = ~n51265 ;
  assign \g350827/_0_  = ~n51296 ;
  assign \g350828/_0_  = ~n51336 ;
  assign \g350829/_0_  = ~n51377 ;
  assign \g350830/_0_  = ~n51429 ;
  assign \g350831/_0_  = ~n51463 ;
  assign \g350832/_0_  = ~n51498 ;
  assign \g350833/_0_  = ~n51542 ;
  assign \g350834/_0_  = ~n51583 ;
  assign \g350835/_0_  = ~n51620 ;
  assign \g350836/_0_  = ~n51650 ;
  assign \g350839/_0_  = ~n51719 ;
  assign \g350840/_0_  = ~n51758 ;
  assign \g350842/_0_  = ~n51795 ;
  assign \g350843/_0_  = ~n51830 ;
  assign \g350844/_0_  = ~n51868 ;
  assign \g350845/_0_  = ~n51903 ;
  assign \g350846/_0_  = ~n51937 ;
  assign \g350847/_0_  = ~n51973 ;
  assign \g350848/_0_  = ~n52007 ;
  assign \g350849/_0_  = ~n52043 ;
  assign \g350850/_0_  = ~n52081 ;
  assign \g350852/_0_  = ~n52149 ;
  assign \g350853/_0_  = ~n52186 ;
  assign \g350854/_0_  = ~n52220 ;
  assign \g350856/_0_  = ~n52255 ;
  assign \g350857/_0_  = ~n52292 ;
  assign \g350858/_0_  = ~n52330 ;
  assign \g350859/_0_  = ~n52370 ;
  assign \g350860/_0_  = ~n52407 ;
  assign \g350861/_0_  = ~n52442 ;
  assign \g350862/_0_  = ~n52482 ;
  assign \g350863/_0_  = ~n52519 ;
  assign \g350866/_0_  = ~n52588 ;
  assign \g350867/_0_  = ~n52623 ;
  assign \g350868/_0_  = ~n52657 ;
  assign \g350869/_0_  = ~n52692 ;
  assign \g350870/_0_  = ~n52726 ;
  assign \g350871/_0_  = ~n52763 ;
  assign \g350872/_0_  = ~n52797 ;
  assign \g350873/_0_  = ~n52831 ;
  assign \g350874/_0_  = ~n52864 ;
  assign \g350952/_0_  = ~n52877 ;
  assign \g350959/_0_  = ~n52891 ;
  assign \g350961/_0_  = ~n52903 ;
  assign \g350964/_0_  = ~n52919 ;
  assign \g350974/_0_  = ~n52931 ;
  assign \g350977/_0_  = ~n52946 ;
  assign \g351003/_0_  = ~n52961 ;
  assign \g351005/_0_  = ~n52972 ;
  assign \g351037/_0_  = ~n52984 ;
  assign \g351045/_0_  = ~n52995 ;
  assign \g351048/_0_  = ~n53008 ;
  assign \g351129/_0_  = ~n53021 ;
  assign \g351147/_0_  = ~n53035 ;
  assign \g351169/_0_  = ~n53046 ;
  assign \g351171/_0_  = ~n53060 ;
  assign \g351175/_0_  = ~n53071 ;
  assign \g351195/_0_  = ~n53086 ;
  assign \g351196/_0_  = ~n53099 ;
  assign \g351197/_0_  = ~n53106 ;
  assign \g351198/_0_  = ~n53112 ;
  assign \g351201/_0_  = ~n53120 ;
  assign \g351202/_0_  = ~n53128 ;
  assign \g351203/_0_  = ~n53141 ;
  assign \g351204/_0_  = ~n53159 ;
  assign \g351205/_0_  = ~n53169 ;
  assign \g351206/_0_  = ~n53179 ;
  assign \g351207/_0_  = ~n53190 ;
  assign \g351208/_0_  = ~n53205 ;
  assign \g351209/_0_  = ~n53219 ;
  assign \g351210/_0_  = ~n53228 ;
  assign \g351211/_0_  = ~n53235 ;
  assign \g351214/_0_  = ~n53244 ;
  assign \g351215/_0_  = ~n53253 ;
  assign \g351216/_0_  = ~n53265 ;
  assign \g351217/_0_  = ~n53282 ;
  assign \g351218/_0_  = ~n53292 ;
  assign \g351219/_0_  = ~n53302 ;
  assign \g351220/_0_  = ~n53312 ;
  assign \g351221/_0_  = ~n53325 ;
  assign \g351222/_0_  = ~n53340 ;
  assign \g351223/_0_  = ~n53348 ;
  assign \g351224/_0_  = ~n53363 ;
  assign \g351225/_0_  = ~n53380 ;
  assign \g351226/_0_  = ~n53391 ;
  assign \g351227/_0_  = ~n53402 ;
  assign \g351228/_0_  = ~n53412 ;
  assign \g351229/_0_  = ~n53422 ;
  assign \g351230/_0_  = ~n53432 ;
  assign \g351231/_0_  = ~n53438 ;
  assign \g351671/_0_  = ~n53445 ;
  assign \g351699/_0_  = ~n53451 ;
  assign \g351703/_0_  = ~n53457 ;
  assign \g351704/_0_  = ~n53463 ;
  assign \g351709/_0_  = ~n53497 ;
  assign \g351711/_0_  = ~n53531 ;
  assign \g351712/_0_  = ~n53564 ;
  assign \g351715/_0_  = ~n53603 ;
  assign \g351716/_0_  = ~n53635 ;
  assign \g351717/_0_  = ~n53668 ;
  assign \g351721/_0_  = ~n53701 ;
  assign \g351722/_0_  = ~n53707 ;
  assign \g351723/_0_  = ~n53740 ;
  assign \g351724/_0_  = ~n53773 ;
  assign \g351725/_0_  = ~n53807 ;
  assign \g351726/_0_  = ~n53842 ;
  assign \g351727/_0_  = ~n53876 ;
  assign \g351728/_0_  = ~n53882 ;
  assign \g351739/_0_  = ~n53917 ;
  assign \g351741/_0_  = ~n53950 ;
  assign \g351742/_0_  = ~n53983 ;
  assign \g351750/_0_  = ~n54017 ;
  assign \g351752/_0_  = ~n54051 ;
  assign \g351753/_0_  = ~n54057 ;
  assign \g351756/_0_  = ~n54091 ;
  assign \g351757/_0_  = ~n54097 ;
  assign \g351759/_0_  = ~n54134 ;
  assign \g351760/_0_  = ~n54170 ;
  assign \g351761/_0_  = ~n54205 ;
  assign \g351766/_0_  = ~n54237 ;
  assign \g351767/_0_  = ~n54270 ;
  assign \g351768/_0_  = ~n54303 ;
  assign \g351771/_0_  = ~n54314 ;
  assign \g351772/_0_  = ~n54324 ;
  assign \g351773/_0_  = ~n54334 ;
  assign \g351775/_0_  = ~n54344 ;
  assign \g351776/_0_  = ~n54354 ;
  assign \g351779/_0_  = ~n54364 ;
  assign \g351780/_0_  = ~n54374 ;
  assign \g351782/_0_  = ~n54384 ;
  assign \g351785/_0_  = ~n54394 ;
  assign \g351786/_0_  = ~n54404 ;
  assign \g351788/_0_  = ~n54414 ;
  assign \g351789/_0_  = ~n54424 ;
  assign \g351790/_0_  = ~n54435 ;
  assign \g351791/_0_  = ~n54445 ;
  assign \g351792/_0_  = ~n54455 ;
  assign \g351793/_0_  = ~n54465 ;
  assign \g351794/_0_  = ~n54475 ;
  assign \g351795/_0_  = ~n54485 ;
  assign \g351796/_0_  = ~n54495 ;
  assign \g351797/_0_  = ~n54505 ;
  assign \g351798/_0_  = ~n54515 ;
  assign \g351799/_0_  = ~n54525 ;
  assign \g351800/_0_  = ~n54535 ;
  assign \g351801/_0_  = ~n54542 ;
  assign \g351802/_0_  = ~n54552 ;
  assign \g351803/_0_  = ~n54562 ;
  assign \g351804/_0_  = ~n54572 ;
  assign \g351805/_0_  = ~n54582 ;
  assign \g351806/_0_  = ~n54592 ;
  assign \g351807/_0_  = ~n54602 ;
  assign \g351808/_0_  = ~n54612 ;
  assign \g351809/_0_  = ~n54622 ;
  assign \g351810/_0_  = ~n54632 ;
  assign \g351811/_0_  = ~n54639 ;
  assign \g351812/_0_  = ~n54645 ;
  assign \g351814/_0_  = ~n54652 ;
  assign \g351817/_0_  = ~n54687 ;
  assign \g351818/_0_  = ~n54721 ;
  assign \g351819/_0_  = ~n54756 ;
  assign \g351821/_0_  = ~n54789 ;
  assign \g351822/_0_  = ~n54822 ;
  assign \g351823/_0_  = ~n54855 ;
  assign \g351841/_0_  = ~n54889 ;
  assign \g351842/_0_  = ~n54925 ;
  assign \g351843/_0_  = ~n54959 ;
  assign \g351844/_0_  = ~n54992 ;
  assign \g351845/_0_  = ~n55024 ;
  assign \g351846/_0_  = ~n55057 ;
  assign \g351847/_0_  = ~n55090 ;
  assign \g351848/_0_  = ~n55125 ;
  assign \g351849/_0_  = ~n55158 ;
  assign \g351850/_0_  = ~n55193 ;
  assign \g351851/_0_  = ~n55225 ;
  assign \g351852/_0_  = ~n55257 ;
  assign \g351853/_0_  = ~n55295 ;
  assign \g351854/_0_  = ~n55326 ;
  assign \g351855/_0_  = ~n55359 ;
  assign \g351856/_0_  = ~n55392 ;
  assign \g351857/_0_  = ~n55424 ;
  assign \g351858/_0_  = ~n55457 ;
  assign \g351859/_0_  = ~n55491 ;
  assign \g351860/_0_  = ~n55525 ;
  assign \g351861/_0_  = ~n55560 ;
  assign \g351862/_0_  = ~n55594 ;
  assign \g351863/_0_  = ~n55627 ;
  assign \g351864/_0_  = ~n55661 ;
  assign \g351865/_0_  = ~n55695 ;
  assign \g351866/_0_  = ~n55729 ;
  assign \g351867/_0_  = ~n55763 ;
  assign \g351868/_0_  = ~n55799 ;
  assign \g351869/_0_  = ~n55834 ;
  assign \g351870/_0_  = ~n55869 ;
  assign \g351871/_0_  = ~n55904 ;
  assign \g351872/_0_  = ~n55937 ;
  assign \g351873/_0_  = ~n55971 ;
  assign \g351874/_0_  = ~n56005 ;
  assign \g351875/_0_  = ~n56039 ;
  assign \g351876/_0_  = ~n56073 ;
  assign \g351877/_0_  = ~n56108 ;
  assign \g351878/_0_  = ~n56142 ;
  assign \g351879/_0_  = ~n56175 ;
  assign \g351880/_0_  = ~n56207 ;
  assign \g351881/_0_  = ~n56241 ;
  assign \g351882/_0_  = ~n56274 ;
  assign \g351883/_0_  = ~n56307 ;
  assign \g351884/_0_  = ~n56340 ;
  assign \g351885/_0_  = ~n56373 ;
  assign \g351889/_0_  = ~n56402 ;
  assign \g351920/_0_  = ~n56423 ;
  assign \g351921/_0_  = ~n56445 ;
  assign \g351922/_0_  = ~n56479 ;
  assign \g351923/_0_  = ~n56507 ;
  assign \g351924/_0_  = ~n56528 ;
  assign \g351925/_0_  = ~n56562 ;
  assign \g351926/_0_  = ~n56591 ;
  assign \g351927/_0_  = ~n56610 ;
  assign \g351928/_0_  = ~n56646 ;
  assign \g351929/_0_  = ~n56673 ;
  assign \g351930/_0_  = ~n56691 ;
  assign \g351954/_0_  = ~n56723 ;
  assign \g351955/_0_  = ~n56764 ;
  assign \g351956/_0_  = ~n56798 ;
  assign \g351957/_0_  = ~n56821 ;
  assign \g352167/_0_  = ~n56829 ;
  assign \g352178/_0_  = ~n56840 ;
  assign \g352211/_0_  = ~n56854 ;
  assign \g352215/_0_  = ~n56868 ;
  assign \g352219/_0_  = ~n56879 ;
  assign \g352237/_0_  = ~n56889 ;
  assign \g352238/_0_  = ~n56892 ;
  assign \g352239/_0_  = ~n56895 ;
  assign \g352240/_0_  = ~n56905 ;
  assign \g352241/_0_  = ~n56911 ;
  assign \g352242/_0_  = ~n56917 ;
  assign \g352243/_0_  = ~n56923 ;
  assign \g352244/_0_  = ~n56929 ;
  assign \g352245/_0_  = ~n56935 ;
  assign \g352246/_0_  = ~n56942 ;
  assign \g352247/_0_  = ~n56948 ;
  assign \g352248/_0_  = ~n56955 ;
  assign \g352249/_0_  = ~n56962 ;
  assign \g352250/_0_  = ~n56967 ;
  assign \g352251/_0_  = ~n56973 ;
  assign \g352252/_0_  = ~n56979 ;
  assign \g352253/_0_  = ~n56986 ;
  assign \g352254/_0_  = ~n56991 ;
  assign \g352255/_0_  = ~n56997 ;
  assign \g352256/_0_  = ~n57000 ;
  assign \g352257/_0_  = ~n57007 ;
  assign \g352258/_0_  = ~n57013 ;
  assign \g352259/_0_  = ~n57063 ;
  assign \g352260/_0_  = ~n57112 ;
  assign \g352261/_0_  = ~n57158 ;
  assign \g352262/_0_  = ~n57204 ;
  assign \g352263/_0_  = ~n57250 ;
  assign \g352264/_0_  = ~n57296 ;
  assign \g352265/_0_  = ~n57342 ;
  assign \g352266/_0_  = ~n57363 ;
  assign \g352267/_0_  = ~n57383 ;
  assign \g352268/_0_  = ~n57402 ;
  assign \g352269/_0_  = ~n57412 ;
  assign \g352271/_0_  = ~n57422 ;
  assign \g352272/_0_  = ~n57425 ;
  assign \g352273/_0_  = ~n57435 ;
  assign \g352274/_0_  = ~n57443 ;
  assign \g352275/_0_  = ~n57450 ;
  assign \g352276/_0_  = ~n57461 ;
  assign \g352277/_0_  = ~n57466 ;
  assign \g352278/_0_  = ~n57472 ;
  assign \g352279/_0_  = ~n57478 ;
  assign \g352280/_0_  = ~n57490 ;
  assign \g352281/_0_  = ~n57496 ;
  assign \g352282/_0_  = ~n57505 ;
  assign \g352283/_0_  = ~n57514 ;
  assign \g352284/_0_  = ~n57523 ;
  assign \g352285/_0_  = ~n57532 ;
  assign \g352286/_0_  = ~n57541 ;
  assign \g352287/_0_  = ~n57550 ;
  assign \g352288/_0_  = ~n57559 ;
  assign \g352289/_0_  = ~n57564 ;
  assign \g352290/_0_  = ~n57570 ;
  assign \g352291/_0_  = ~n57576 ;
  assign \g352292/_0_  = ~n57625 ;
  assign \g352293/_0_  = ~n57675 ;
  assign \g352294/_0_  = ~n57721 ;
  assign \g352295/_0_  = ~n57767 ;
  assign \g352296/_0_  = ~n57817 ;
  assign \g352297/_0_  = ~n57864 ;
  assign \g352298/_0_  = ~n57913 ;
  assign \g352299/_0_  = ~n57930 ;
  assign \g352300/_0_  = ~n57948 ;
  assign \g352301/_0_  = ~n57967 ;
  assign \g352302/_0_  = ~n57977 ;
  assign \g352303/_0_  = ~n58024 ;
  assign \g352304/_0_  = ~n58072 ;
  assign \g352305/_0_  = ~n58117 ;
  assign \g352306/_0_  = ~n58162 ;
  assign \g352307/_0_  = ~n58208 ;
  assign \g352308/_0_  = ~n58252 ;
  assign \g352309/_0_  = ~n58296 ;
  assign \g352310/_0_  = ~n58312 ;
  assign \g352311/_0_  = ~n58315 ;
  assign \g352312/_0_  = ~n58331 ;
  assign \g352313/_0_  = ~n58351 ;
  assign \g352314/_0_  = ~n58356 ;
  assign \g352315/_0_  = ~n58366 ;
  assign \g352525/_0_  = ~n58375 ;
  assign \g352527/_0_  = ~n58386 ;
  assign \g352529/_0_  = ~n58396 ;
  assign \g352547/_0_  = ~n58406 ;
  assign \g352553/_0_  = ~n58420 ;
  assign \g352554/_0_  = ~n58434 ;
  assign \g352556/_0_  = ~n58447 ;
  assign \g352558/_0_  = ~n58460 ;
  assign \g352559/_0_  = ~n58473 ;
  assign \g352560/_0_  = ~n58486 ;
  assign \g352561/_0_  = ~n58499 ;
  assign \g352563/_0_  = ~n58512 ;
  assign \g352564/_0_  = ~n58526 ;
  assign \g352565/_0_  = ~n58540 ;
  assign \g352567/_0_  = ~n58554 ;
  assign \g352568/_0_  = ~n58568 ;
  assign \g352569/_0_  = ~n58581 ;
  assign \g352570/_0_  = ~n58594 ;
  assign \g352572/_0_  = ~n58607 ;
  assign \g352574/_0_  = ~n58620 ;
  assign \g352575/_0_  = ~n58633 ;
  assign \g352577/_0_  = ~n58646 ;
  assign \g352579/_0_  = ~n58660 ;
  assign \g352581/_0_  = ~n58674 ;
  assign \g352583/_0_  = ~n58688 ;
  assign \g352584/_0_  = ~n58702 ;
  assign \g352585/_0_  = ~n58716 ;
  assign \g352586/_0_  = ~n58730 ;
  assign \g352587/_0_  = ~n58744 ;
  assign \g352588/_0_  = ~n58757 ;
  assign \g352589/_0_  = ~n58771 ;
  assign \g352590/_0_  = ~n58784 ;
  assign \g352591/_0_  = ~n58797 ;
  assign \g352592/_0_  = ~n58810 ;
  assign \g352593/_0_  = ~n58824 ;
  assign \g352594/_0_  = ~n58837 ;
  assign \g352595/_0_  = ~n58851 ;
  assign \g352596/_0_  = ~n58864 ;
  assign \g352597/_0_  = ~n58877 ;
  assign \g352598/_0_  = ~n58890 ;
  assign \g352599/_0_  = ~n58904 ;
  assign \g352600/_0_  = ~n58917 ;
  assign \g352601/_0_  = ~n58931 ;
  assign \g352602/_0_  = ~n58944 ;
  assign \g352603/_0_  = ~n58957 ;
  assign \g352605/_0_  = ~n58970 ;
  assign \g352606/_0_  = ~n58983 ;
  assign \g352607/_0_  = ~n58996 ;
  assign \g352608/_0_  = ~n59009 ;
  assign \g352609/_0_  = ~n59022 ;
  assign \g352610/_0_  = ~n59035 ;
  assign \g352611/_0_  = ~n59045 ;
  assign \g352612/_0_  = ~n59058 ;
  assign \g352613/_0_  = ~n59071 ;
  assign \g352614/_0_  = ~n59084 ;
  assign \g352615/_0_  = ~n59097 ;
  assign \g352616/_0_  = ~n59110 ;
  assign \g352617/_0_  = ~n59123 ;
  assign \g352618/_0_  = ~n59136 ;
  assign \g352619/_0_  = ~n59149 ;
  assign \g352620/_0_  = ~n59162 ;
  assign \g352621/_0_  = ~n59175 ;
  assign \g352622/_0_  = ~n59188 ;
  assign \g352623/_0_  = ~n59201 ;
  assign \g352624/_0_  = ~n59214 ;
  assign \g352625/_0_  = ~n59227 ;
  assign \g352626/_0_  = ~n59240 ;
  assign \g352627/_0_  = ~n59253 ;
  assign \g352628/_0_  = ~n59266 ;
  assign \g352629/_0_  = ~n59276 ;
  assign \g352662/_0_  = ~n59310 ;
  assign \g352663/_0_  = ~n59344 ;
  assign \g352666/_0_  = ~n59378 ;
  assign \g352667/_0_  = ~n59411 ;
  assign \g352668/_0_  = ~n59440 ;
  assign \g352676/_0_  = ~n59449 ;
  assign \g352677/_0_  = ~n59459 ;
  assign \g352678/_0_  = ~n59469 ;
  assign \g352683/_0_  = ~n59478 ;
  assign \g352684/_0_  = ~n59487 ;
  assign \g352685/_0_  = ~n59498 ;
  assign \g353014/_0_  = ~n59509 ;
  assign \g353016/_0_  = ~n59520 ;
  assign \g353035/_0_  = ~n59531 ;
  assign \g353036/_0_  = ~n59542 ;
  assign \g353065/_0_  = ~n59550 ;
  assign \g353067/_0_  = ~n59561 ;
  assign \g353071/_0_  = ~n59572 ;
  assign \g353073/_0_  = ~n59583 ;
  assign \g353085/_0_  = ~n59594 ;
  assign \g353087/_0_  = ~n59605 ;
  assign \g353116/_0_  = ~n59615 ;
  assign \g353119/_0_  = ~n59625 ;
  assign \g353120/_0_  = ~n59635 ;
  assign \g353121/_0_  = ~n59645 ;
  assign \g353122/_0_  = ~n59655 ;
  assign \g353123/_0_  = ~n59665 ;
  assign \g353124/_0_  = ~n59675 ;
  assign \g353125/_0_  = ~n59685 ;
  assign \g353126/_0_  = ~n59695 ;
  assign \g353127/_0_  = ~n59705 ;
  assign \g353128/_0_  = ~n59715 ;
  assign \g353130/_0_  = ~n59725 ;
  assign \g353131/_0_  = ~n59735 ;
  assign \g353132/_0_  = ~n59745 ;
  assign \g353133/_0_  = ~n59755 ;
  assign \g353134/_0_  = ~n59765 ;
  assign \g353135/_0_  = ~n59775 ;
  assign \g353136/_0_  = ~n59785 ;
  assign \g353137/_0_  = ~n59795 ;
  assign \g353138/_0_  = ~n59798 ;
  assign \g353142/_0_  = ~n59801 ;
  assign \g353148/_0_  = ~n59809 ;
  assign \g353149/_0_  = ~n59819 ;
  assign \g353150/_0_  = ~n59826 ;
  assign \g353151/_0_  = ~n59835 ;
  assign \g353152/_0_  = ~n59843 ;
  assign \g353153/_0_  = ~n59853 ;
  assign \g353154/_0_  = ~n59865 ;
  assign \g353155/_0_  = ~n59874 ;
  assign \g353157/_0_  = ~n59886 ;
  assign \g353158/_0_  = ~n59895 ;
  assign \g353159/_0_  = ~n59902 ;
  assign \g353160/_0_  = ~n59911 ;
  assign \g353161/_0_  = ~n59917 ;
  assign \g353162/_0_  = ~n59926 ;
  assign \g353163/_0_  = ~n59936 ;
  assign \g353164/_0_  = ~n59946 ;
  assign \g353165/_0_  = ~n59956 ;
  assign \g353166/_0_  = ~n59966 ;
  assign \g353167/_0_  = ~n59976 ;
  assign \g353168/_0_  = ~n59986 ;
  assign \g353169/_0_  = ~n59996 ;
  assign \g353170/_0_  = ~n60006 ;
  assign \g353171/_0_  = ~n60016 ;
  assign \g353172/_0_  = ~n60026 ;
  assign \g353173/_0_  = ~n60036 ;
  assign \g353174/_0_  = ~n60046 ;
  assign \g353175/_0_  = ~n60056 ;
  assign \g353176/_0_  = ~n60066 ;
  assign \g353177/_0_  = ~n60076 ;
  assign \g353178/_0_  = ~n60086 ;
  assign \g353179/_0_  = ~n60096 ;
  assign \g353180/_0_  = ~n60106 ;
  assign \g353181/_0_  = ~n60109 ;
  assign \g353184/_0_  = ~n60119 ;
  assign \g353185/_0_  = ~n60129 ;
  assign \g353186/_0_  = ~n60139 ;
  assign \g353187/_0_  = ~n60149 ;
  assign \g353188/_0_  = ~n60159 ;
  assign \g353189/_0_  = ~n60169 ;
  assign \g353190/_0_  = ~n60179 ;
  assign \g353191/_0_  = ~n60189 ;
  assign \g353192/_0_  = ~n60199 ;
  assign \g353193/_0_  = ~n60209 ;
  assign \g353194/_0_  = ~n60219 ;
  assign \g353195/_0_  = ~n60229 ;
  assign \g353196/_0_  = ~n60239 ;
  assign \g353197/_0_  = ~n60249 ;
  assign \g353198/_0_  = ~n60259 ;
  assign \g353199/_0_  = ~n60269 ;
  assign \g353200/_0_  = ~n60279 ;
  assign \g353201/_0_  = ~n60289 ;
  assign \g353202/_0_  = ~n60299 ;
  assign \g353203/_0_  = ~n60309 ;
  assign \g353204/_0_  = ~n60319 ;
  assign \g353205/_0_  = ~n60329 ;
  assign \g353206/_0_  = ~n60339 ;
  assign \g353207/_0_  = ~n60349 ;
  assign \g353208/_0_  = ~n60359 ;
  assign \g353209/_0_  = ~n60369 ;
  assign \g353210/_0_  = ~n60379 ;
  assign \g353211/_0_  = ~n60389 ;
  assign \g353212/_0_  = ~n60399 ;
  assign \g353213/_0_  = ~n60409 ;
  assign \g353214/_0_  = ~n60419 ;
  assign \g353215/_0_  = ~n60429 ;
  assign \g353216/_0_  = ~n60442 ;
  assign \g353217/_0_  = ~n60454 ;
  assign \g353218/_0_  = ~n60463 ;
  assign \g353219/_0_  = ~n60470 ;
  assign \g353220/_0_  = ~n60480 ;
  assign \g353221/_0_  = ~n60490 ;
  assign \g353222/_0_  = ~n60502 ;
  assign \g353223/_0_  = ~n60512 ;
  assign \g353224/_0_  = ~n60522 ;
  assign \g353225/_0_  = ~n60530 ;
  assign \g353226/_0_  = ~n60538 ;
  assign \g353227/_0_  = ~n60550 ;
  assign \g353228/_0_  = ~n60560 ;
  assign \g353229/_0_  = ~n60567 ;
  assign \g353230/_0_  = ~n60579 ;
  assign \g353231/_0_  = ~n60582 ;
  assign \g353232/_0_  = ~n60594 ;
  assign \g353233/_0_  = ~n60598 ;
  assign \g353234/_0_  = ~n60605 ;
  assign \g353235/_0_  = ~n60615 ;
  assign \g353236/_0_  = ~n60625 ;
  assign \g353237/_0_  = ~n60635 ;
  assign \g353238/_0_  = ~n60645 ;
  assign \g353239/_0_  = ~n60655 ;
  assign \g353240/_0_  = ~n60665 ;
  assign \g353241/_0_  = ~n60675 ;
  assign \g353242/_0_  = ~n60685 ;
  assign \g353243/_0_  = ~n60695 ;
  assign \g353244/_0_  = ~n60705 ;
  assign \g353245/_0_  = ~n60715 ;
  assign \g353246/_0_  = ~n60725 ;
  assign \g353247/_0_  = ~n60735 ;
  assign \g353248/_0_  = ~n60745 ;
  assign \g353249/_0_  = ~n60755 ;
  assign \g353250/_0_  = ~n60765 ;
  assign \g353251/_0_  = ~n60775 ;
  assign \g353252/_0_  = ~n60785 ;
  assign \g353253/_0_  = ~n60788 ;
  assign \g353254/_0_  = ~n60796 ;
  assign \g353255/_0_  = ~n60805 ;
  assign \g353256/_0_  = ~n60816 ;
  assign \g353257/_0_  = ~n60826 ;
  assign \g353258/_0_  = ~n60834 ;
  assign \g353259/_0_  = ~n60847 ;
  assign \g353260/_0_  = ~n60857 ;
  assign \g353261/_0_  = ~n60865 ;
  assign \g353262/_0_  = ~n60874 ;
  assign \g353263/_0_  = ~n60879 ;
  assign \g353264/_0_  = ~n60892 ;
  assign \g353265/_0_  = ~n60902 ;
  assign \g353266/_0_  = ~n60912 ;
  assign \g353267/_0_  = ~n60922 ;
  assign \g353268/_0_  = ~n60932 ;
  assign \g353269/_0_  = ~n60942 ;
  assign \g353270/_0_  = ~n60952 ;
  assign \g353271/_0_  = ~n60962 ;
  assign \g353272/_0_  = ~n60972 ;
  assign \g353273/_0_  = ~n60982 ;
  assign \g353274/_0_  = ~n60992 ;
  assign \g353275/_0_  = ~n61002 ;
  assign \g353276/_0_  = ~n61012 ;
  assign \g353277/_0_  = ~n61022 ;
  assign \g353278/_0_  = ~n61032 ;
  assign \g353279/_0_  = ~n61042 ;
  assign \g353280/_0_  = ~n61052 ;
  assign \g353281/_0_  = ~n61062 ;
  assign \g354206/_0_  = ~n61070 ;
  assign \g354214/_0_  = ~n61077 ;
  assign \g354216/_0_  = ~n61085 ;
  assign \g354217/_0_  = ~n61089 ;
  assign \g354222/_0_  = ~n61102 ;
  assign \g354278/_0_  = ~n61109 ;
  assign \g354282/_0_  = ~n61115 ;
  assign \g354284/_0_  = ~n61123 ;
  assign \g354289/_0_  = ~n61129 ;
  assign \g354301/_0_  = ~n61140 ;
  assign \g354330/_0_  = ~n61145 ;
  assign \g354331/_0_  = ~n61156 ;
  assign \g354332/_0_  = ~n61161 ;
  assign \g354333/_0_  = ~n61172 ;
  assign \g354335/_0_  = ~n61182 ;
  assign \g354336/_0_  = ~n61192 ;
  assign \g354337/_0_  = ~n61202 ;
  assign \g354338/_0_  = ~n61207 ;
  assign \g354339/_0_  = ~n61217 ;
  assign \g354340/_0_  = ~n61227 ;
  assign \g354341/_0_  = ~n61232 ;
  assign \g354342/_0_  = ~n61243 ;
  assign \g354343/_0_  = ~n61249 ;
  assign \g354344/_0_  = ~n61260 ;
  assign \g354345/_0_  = ~n61271 ;
  assign \g354346/_0_  = ~n61281 ;
  assign \g354358/_0_  = ~n61287 ;
  assign \g354364/_0_  = ~n61295 ;
  assign \g354442/_0_  = ~n61305 ;
  assign \g354444/_0_  = ~n61313 ;
  assign \g354445/_0_  = ~n61324 ;
  assign \g354447/_0_  = ~n61335 ;
  assign \g354448/_0_  = ~n61348 ;
  assign \g354449/_0_  = ~n61358 ;
  assign \g354450/_0_  = ~n61371 ;
  assign \g354451/_0_  = ~n61381 ;
  assign \g354452/_0_  = ~n61394 ;
  assign \g354455/_0_  = ~n61399 ;
  assign \g354456/_0_  = ~n61404 ;
  assign \g354464/_0_  = ~n61412 ;
  assign \g354465/_0_  = ~n61420 ;
  assign \g354466/_0_  = ~n61432 ;
  assign \g354468/_0_  = ~n61443 ;
  assign \g354469/_0_  = ~n61455 ;
  assign \g354470/_0_  = ~n61465 ;
  assign \g354471/_0_  = ~n61475 ;
  assign \g354472/_0_  = ~n61485 ;
  assign \g354473/_0_  = ~n61498 ;
  assign \g354474/_0_  = ~n61506 ;
  assign \g354477/_0_  = ~n61517 ;
  assign \g354478/_0_  = ~n61525 ;
  assign \g354479/_0_  = ~n61533 ;
  assign \g354480/_0_  = ~n61546 ;
  assign \g354482/_0_  = ~n61556 ;
  assign \g354483/_0_  = ~n61566 ;
  assign \g354484/_0_  = ~n61576 ;
  assign \g354485/_0_  = ~n61586 ;
  assign \g354486/_0_  = ~n61596 ;
  assign \g354487/_0_  = ~n61606 ;
  assign \g354488/_0_  = ~n61617 ;
  assign \g354490/_0_  = ~n61628 ;
  assign \g354491/_0_  = ~n61641 ;
  assign \g354492/_0_  = ~n61651 ;
  assign \g354493/_0_  = ~n61664 ;
  assign \g354494/_0_  = ~n61674 ;
  assign \g354495/_0_  = ~n61687 ;
  assign \g354504/_0_  = ~n61697 ;
  assign \g354505/_0_  = ~n61705 ;
  assign \g354506/_0_  = ~n61718 ;
  assign \g354508/_0_  = ~n61728 ;
  assign \g354509/_0_  = ~n61738 ;
  assign \g354510/_0_  = ~n61748 ;
  assign \g354511/_0_  = ~n61758 ;
  assign \g354512/_0_  = ~n61768 ;
  assign \g354513/_0_  = ~n61778 ;
  assign \g354522/_0_  = ~n61786 ;
  assign \g354524/_0_  = ~n61796 ;
  assign \g354525/_0_  = ~n61806 ;
  assign \g354526/_0_  = ~n61816 ;
  assign \g354527/_0_  = ~n61829 ;
  assign \g354920/_1_  = n18665 ;
  assign \g355460/_0_  = ~n61837 ;
  assign \g355461/_0_  = ~n61845 ;
  assign \g355463/_0_  = ~n61853 ;
  assign \g355464/_0_  = ~n61861 ;
  assign \g355466/_0_  = ~n61872 ;
  assign \g355467/_0_  = ~n61880 ;
  assign \g355470/_0_  = ~n61891 ;
  assign \g355471/_0_  = ~n61899 ;
  assign \g355475/_0_  = ~n61907 ;
  assign \g355476/_0_  = ~n61915 ;
  assign \g355477/_0_  = ~n61926 ;
  assign \g355479/_0_  = ~n61934 ;
  assign \g355480/_0_  = ~n61942 ;
  assign \g355481/_0_  = ~n61953 ;
  assign \g355482/_0_  = ~n61964 ;
  assign \g355483/_0_  = ~n61972 ;
  assign \g355508/_0_  = ~n61980 ;
  assign \g355509/_0_  = ~n61988 ;
  assign \g355510/_0_  = ~n61996 ;
  assign \g355511/_0_  = ~n62004 ;
  assign \g355512/_0_  = ~n62010 ;
  assign \g355513/_0_  = ~n62015 ;
  assign \g355514/_0_  = ~n62023 ;
  assign \g355515/_0_  = ~n62031 ;
  assign \g355520/_0_  = ~n62042 ;
  assign \g355521/_0_  = ~n62050 ;
  assign \g355523/_0_  = ~n62058 ;
  assign \g355525/_0_  = ~n62066 ;
  assign \g355527/_0_  = ~n62077 ;
  assign \g355530/_0_  = ~n62088 ;
  assign \g355532/_0_  = ~n62096 ;
  assign \g355534/_0_  = ~n62104 ;
  assign \g355564/_0_  = ~n62115 ;
  assign \g355565/_0_  = ~n62126 ;
  assign \g355566/_0_  = ~n62137 ;
  assign \g355567/_0_  = ~n62148 ;
  assign \g355568/_0_  = ~n62159 ;
  assign \g355569/_0_  = ~n62167 ;
  assign \g355570/_0_  = ~n62178 ;
  assign \g355571/_0_  = ~n62186 ;
  assign \g355980/_0_  = ~n62202 ;
  assign \g356052/_0_  = ~n62220 ;
  assign \g356106/_0_  = ~n62234 ;
  assign \g356111/_0_  = ~n62247 ;
  assign \g356114/_0_  = ~n62260 ;
  assign \g356117/_0_  = ~n62273 ;
  assign \g356122/_0_  = ~n62287 ;
  assign \g356126/_0_  = ~n62301 ;
  assign \g356129/_0_  = ~n62314 ;
  assign \g356133/_0_  = ~n62327 ;
  assign \g356142/_0_  = ~n62340 ;
  assign \g356148/_0_  = ~n62354 ;
  assign \g356151/_0_  = ~n62368 ;
  assign \g356155/_0_  = ~n62382 ;
  assign \g356160/_0_  = ~n62396 ;
  assign \g356162/_0_  = ~n62409 ;
  assign \g356165/_0_  = ~n62422 ;
  assign \g356167/_0_  = ~n62436 ;
  assign \g356170/_0_  = ~n62449 ;
  assign \g356174/_0_  = ~n62462 ;
  assign \g356176/_0_  = ~n62476 ;
  assign \g356179/_0_  = ~n62489 ;
  assign \g356183/_0_  = ~n62502 ;
  assign \g356185/_0_  = ~n62515 ;
  assign \g356189/_0_  = ~n62528 ;
  assign \g356193/_0_  = ~n62541 ;
  assign \g356196/_0_  = ~n62554 ;
  assign \g356199/_0_  = ~n62567 ;
  assign \g356202/_0_  = ~n62580 ;
  assign \g356205/_0_  = ~n62593 ;
  assign \g356207/_0_  = ~n62606 ;
  assign \g356210/_0_  = ~n62619 ;
  assign \g356213/_0_  = ~n62632 ;
  assign \g356215/_0_  = ~n62645 ;
  assign \g357046/_0_  = ~n62653 ;
  assign \g357047/_0_  = ~n62661 ;
  assign \g357048/_0_  = ~n62669 ;
  assign \g357051/_0_  = ~n62677 ;
  assign \g357052/_0_  = ~n62685 ;
  assign \g357053/_0_  = ~n62693 ;
  assign \g357054/_0_  = ~n62701 ;
  assign \g357055/_0_  = ~n62709 ;
  assign \g357056/_0_  = ~n62717 ;
  assign \g357057/_0_  = ~n62725 ;
  assign \g357058/_0_  = ~n62733 ;
  assign \g357059/_0_  = ~n62741 ;
  assign \g357060/_0_  = ~n62749 ;
  assign \g357061/_0_  = ~n62757 ;
  assign \g357062/_0_  = ~n62765 ;
  assign \g357063/_0_  = ~n62773 ;
  assign \g357064/_0_  = ~n62781 ;
  assign \g357065/_0_  = ~n62789 ;
  assign \g357066/_0_  = ~n62797 ;
  assign \g357067/_0_  = ~n62805 ;
  assign \g357068/_0_  = ~n62813 ;
  assign \g357069/_0_  = ~n62821 ;
  assign \g357070/_0_  = ~n62829 ;
  assign \g357071/_0_  = ~n62837 ;
  assign \g357072/_0_  = ~n62845 ;
  assign \g357073/_0_  = ~n62853 ;
  assign \g357074/_0_  = ~n62861 ;
  assign \g357099/_0_  = ~n62869 ;
  assign \g357100/_0_  = ~n62877 ;
  assign \g357101/_0_  = ~n62885 ;
  assign \g357102/_0_  = ~n62893 ;
  assign \g357103/_0_  = ~n62901 ;
  assign \g357104/_0_  = ~n62909 ;
  assign \g357105/_0_  = ~n62917 ;
  assign \g357106/_0_  = ~n62925 ;
  assign \g357107/_0_  = ~n62933 ;
  assign \g357108/_0_  = ~n62941 ;
  assign \g357109/_0_  = ~n62949 ;
  assign \g357110/_0_  = ~n62957 ;
  assign \g357111/_0_  = ~n62965 ;
  assign \g357112/_0_  = ~n62973 ;
  assign \g357113/_0_  = ~n62981 ;
  assign \g357114/_0_  = ~n62989 ;
  assign \g357116/_0_  = ~n62997 ;
  assign \g357119/_0_  = ~n63005 ;
  assign \g357121/_0_  = ~n63013 ;
  assign \g357122/_0_  = ~n63021 ;
  assign \g357123/_0_  = ~n63029 ;
  assign \g357124/_0_  = ~n63037 ;
  assign \g357125/_0_  = ~n63045 ;
  assign \g357126/_0_  = ~n63053 ;
  assign \g357128/_0_  = ~n63061 ;
  assign \g357129/_0_  = ~n63069 ;
  assign \g357130/_0_  = ~n63077 ;
  assign \g357131/_0_  = ~n63085 ;
  assign \g357132/_0_  = ~n63093 ;
  assign \g357133/_0_  = ~n63101 ;
  assign \g357134/_0_  = ~n63109 ;
  assign \g357135/_0_  = ~n63117 ;
  assign \g357142/_0_  = ~n63125 ;
  assign \g357144/_0_  = ~n63133 ;
  assign \g357145/_0_  = ~n63141 ;
  assign \g357146/_0_  = ~n63149 ;
  assign \g357147/_0_  = ~n63157 ;
  assign \g357148/_0_  = ~n63165 ;
  assign \g357149/_0_  = ~n63173 ;
  assign \g357150/_0_  = ~n63181 ;
  assign \g357151/_0_  = ~n63189 ;
  assign \g357152/_0_  = ~n63197 ;
  assign \g357153/_0_  = ~n63205 ;
  assign \g357154/_0_  = ~n63213 ;
  assign \g357155/_0_  = ~n63221 ;
  assign \g357156/_0_  = ~n63229 ;
  assign \g357157/_0_  = ~n63237 ;
  assign \g357158/_0_  = ~n63245 ;
  assign \g357160/_0_  = ~n63253 ;
  assign \g357161/_0_  = ~n63261 ;
  assign \g357163/_0_  = ~n63269 ;
  assign \g357164/_0_  = ~n63277 ;
  assign \g357165/_0_  = ~n63285 ;
  assign \g357288/_0_  = ~n63300 ;
  assign \g357289/_0_  = ~n63315 ;
  assign \g357413/_0_  = ~n63325 ;
  assign \g357414/_0_  = ~n63335 ;
  assign \g357464/_0_  = ~n63341 ;
  assign \g357510/_0_  = ~n63348 ;
  assign \g357733/_0_  = ~n63378 ;
  assign \g357769/_0_  = ~n63418 ;
  assign \g357781/_0_  = ~n63449 ;
  assign \g357828/_0_  = ~n63485 ;
  assign \g358792/_0_  = ~n63504 ;
  assign \g358802/_0_  = ~n63521 ;
  assign \g359042/_0_  = ~n63539 ;
  assign \g359043/_0_  = ~n63553 ;
  assign \g359045/_0_  = ~n63566 ;
  assign \g359048/_0_  = ~n63579 ;
  assign \g359051/_0_  = ~n63592 ;
  assign \g359053/_0_  = ~n63606 ;
  assign \g359057/_0_  = ~n63620 ;
  assign \g359060/_0_  = ~n63633 ;
  assign \g359064/_0_  = ~n63646 ;
  assign \g359070/_0_  = ~n63659 ;
  assign \g359074/_0_  = ~n63673 ;
  assign \g359077/_0_  = ~n63687 ;
  assign \g359080/_0_  = ~n63701 ;
  assign \g359086/_0_  = ~n63720 ;
  assign \g359087/_0_  = ~n63734 ;
  assign \g359088/_0_  = ~n63747 ;
  assign \g359090/_0_  = ~n63760 ;
  assign \g359092/_0_  = ~n63774 ;
  assign \g359094/_0_  = ~n63787 ;
  assign \g359096/_0_  = ~n63800 ;
  assign \g359097/_0_  = ~n63814 ;
  assign \g359099/_0_  = ~n63827 ;
  assign \g359101/_0_  = ~n63840 ;
  assign \g359102/_0_  = ~n63853 ;
  assign \g359104/_0_  = ~n63866 ;
  assign \g359106/_0_  = ~n63879 ;
  assign \g359107/_0_  = ~n63892 ;
  assign \g359108/_0_  = ~n63905 ;
  assign \g359110/_0_  = ~n63918 ;
  assign \g359111/_0_  = ~n63931 ;
  assign \g359112/_0_  = ~n63944 ;
  assign \g359113/_0_  = ~n63957 ;
  assign \g359116/_0_  = ~n63970 ;
  assign \g359118/_0_  = ~n63983 ;
  assign \g359572/_0_  = ~n64005 ;
  assign \g359573/_0_  = ~n64020 ;
  assign \g359577/_0_  = ~n64039 ;
  assign \g359585/_0_  = ~n64057 ;
  assign \g359887/_0_  = ~n64092 ;
  assign \g359888/_0_  = ~n64124 ;
  assign \g360077/_0_  = ~n64139 ;
  assign \g360083/_0_  = ~n64154 ;
  assign \g360113/_0_  = ~n64169 ;
  assign \g360124/_0_  = ~n64184 ;
  assign \g360302/_0_  = ~n64194 ;
  assign \g360303/_0_  = ~n64204 ;
  assign \g360304/_0_  = ~n64214 ;
  assign \g360305/_0_  = ~n64224 ;
  assign \g360320/_0_  = ~n64230 ;
  assign \g360325/_0_  = ~n64236 ;
  assign \g360361/_0_  = ~n64249 ;
  assign \g360371/_0_  = ~n64262 ;
  assign \g360440/_0_  = ~n64268 ;
  assign \g360441/_0_  = ~n64282 ;
  assign \g360443/_0_  = ~n64295 ;
  assign \g360445/_0_  = ~n64308 ;
  assign \g360446/_0_  = ~n64321 ;
  assign \g360448/_0_  = ~n64334 ;
  assign \g360450/_0_  = ~n64348 ;
  assign \g360453/_0_  = ~n64362 ;
  assign \g360462/_0_  = ~n64375 ;
  assign \g360469/_0_  = ~n64388 ;
  assign \g360476/_0_  = ~n64402 ;
  assign \g360478/_0_  = ~n64416 ;
  assign \g360480/_0_  = ~n64430 ;
  assign \g360485/_0_  = ~n64444 ;
  assign \g360487/_0_  = ~n64458 ;
  assign \g360489/_0_  = ~n64471 ;
  assign \g360491/_0_  = ~n64485 ;
  assign \g360492/_0_  = ~n64498 ;
  assign \g360494/_0_  = ~n64512 ;
  assign \g360497/_0_  = ~n64525 ;
  assign \g360498/_0_  = ~n64538 ;
  assign \g360504/_0_  = ~n64551 ;
  assign \g360506/_0_  = ~n64565 ;
  assign \g360514/_0_  = ~n64578 ;
  assign \g360516/_0_  = ~n64591 ;
  assign \g360518/_0_  = ~n64604 ;
  assign \g360522/_0_  = ~n64617 ;
  assign \g360524/_0_  = ~n64630 ;
  assign \g360527/_0_  = ~n64643 ;
  assign \g360528/_0_  = ~n64656 ;
  assign \g360530/_0_  = ~n64669 ;
  assign \g360533/_0_  = ~n64682 ;
  assign \g360535/_0_  = ~n64695 ;
  assign \g360538/_0_  = ~n64708 ;
  assign \g360539/_0_  = ~n64721 ;
  assign \g360542/_0_  = ~n64734 ;
  assign \g360546/_0_  = ~n64747 ;
  assign \g360593/_0_  = ~n64753 ;
  assign \g361116/_0_  = ~n64763 ;
  assign \g361128/_0_  = ~n64774 ;
  assign \g361132/_0_  = ~n64785 ;
  assign \g361137/_0_  = ~n64796 ;
  assign \g361616/_0_  = ~n64808 ;
  assign \g361624/_0_  = ~n64818 ;
  assign \g361626/_0_  = ~n64831 ;
  assign \g361627/_0_  = ~n64840 ;
  assign \g361630/_0_  = ~n64855 ;
  assign \g361631/_0_  = ~n64866 ;
  assign \g362129/_0_  = ~n64879 ;
  assign \g362558/_0_  = ~n64893 ;
  assign \g362560/_0_  = ~n64906 ;
  assign \g362564/_0_  = ~n64919 ;
  assign \g362567/_0_  = ~n64933 ;
  assign \g362575/_0_  = ~n64947 ;
  assign \g362586/_0_  = ~n64960 ;
  assign \g362598/_0_  = ~n64973 ;
  assign \g362608/_0_  = ~n64986 ;
  assign \g362627/_0_  = ~n65000 ;
  assign \g362638/_0_  = ~n65014 ;
  assign \g362648/_0_  = ~n65028 ;
  assign \g362650/_0_  = ~n65041 ;
  assign \g362653/_0_  = ~n65054 ;
  assign \g362663/_0_  = ~n65067 ;
  assign \g362664/_0_  = ~n65081 ;
  assign \g362667/_0_  = ~n65094 ;
  assign \g362671/_0_  = ~n65107 ;
  assign \g362673/_0_  = ~n65120 ;
  assign \g362676/_0_  = ~n65133 ;
  assign \g362679/_0_  = ~n65146 ;
  assign \g362686/_0_  = ~n65159 ;
  assign \g362688/_0_  = ~n65172 ;
  assign \g362693/_0_  = ~n65185 ;
  assign \g362697/_0_  = ~n65198 ;
  assign \g362703/_0_  = ~n65211 ;
  assign \g363274/_0_  = ~n65223 ;
  assign \g363290/_0_  = ~n65237 ;
  assign \g363294/_0_  = ~n65250 ;
  assign \g363303/_0_  = ~n65262 ;
  assign \g363608/_0_  = ~n65272 ;
  assign \g363609/_0_  = ~n65282 ;
  assign \g363615/_0_  = ~n65295 ;
  assign \g363616/_0_  = ~n65308 ;
  assign \g363617/_0_  = ~n65318 ;
  assign \g363627/_0_  = ~n65328 ;
  assign \g363818/_3_  = ~n65331 ;
  assign \g365385/_0_  = ~n65345 ;
  assign \g365388/_0_  = ~n65359 ;
  assign \g365391/_0_  = ~n65373 ;
  assign \g365393/_0_  = ~n65387 ;
  assign \g365394/_0_  = ~n65401 ;
  assign \g365398/_0_  = ~n65415 ;
  assign \g365474/_0_  = ~n65424 ;
  assign \g365477/_0_  = ~n65434 ;
  assign \g366167/_0_  = ~n65445 ;
  assign \g366168/_0_  = ~n65454 ;
  assign \g366169/_0_  = ~n65464 ;
  assign \g366170/_0_  = ~n65475 ;
  assign \g366171/_0_  = ~n65485 ;
  assign \g366172/_0_  = ~n65497 ;
  assign \g366173/_0_  = ~n65509 ;
  assign \g366174/_0_  = ~n65519 ;
  assign \g366523/_3_  = ~n65522 ;
  assign \g369170/_0_  = ~n65533 ;
  assign \g369171/_0_  = ~n65542 ;
  assign \g369173/_0_  = ~n65554 ;
  assign \g369177/_0_  = ~n65565 ;
  assign \g369289/_0_  = ~n65575 ;
  assign \g369290/_0_  = ~n65585 ;
  assign \g369291/_0_  = ~n65595 ;
  assign \g369292/_0_  = ~n65605 ;
  assign \g369293/_0_  = ~n65615 ;
  assign \g369294/_0_  = ~n65625 ;
  assign \g369453/_3_  = ~n65628 ;
  assign \g371379/_0_  = ~n65637 ;
  assign \g371381/_0_  = ~n65646 ;
  assign \g371384/_0_  = ~n65655 ;
  assign \g371386/_0_  = ~n65664 ;
  assign \g371387/_0_  = ~n65673 ;
  assign \g371391/_0_  = ~n65682 ;
  assign \g372221/_0_  = ~n65693 ;
  assign \g372222/_0_  = ~n65705 ;
  assign \g372232/_0_  = ~n65717 ;
  assign \g372246/_0_  = ~n65728 ;
  assign \g372249/_0_  = ~n65737 ;
  assign \g372250/_0_  = ~n65746 ;
  assign \g372251/_0_  = ~n65756 ;
  assign \g372252/_0_  = ~n65765 ;
  assign \g372253/_0_  = ~n65774 ;
  assign \g372254/_0_  = ~n65783 ;
  assign \g372454/_3_  = ~n65805 ;
  assign \g372455/_3_  = ~n65827 ;
  assign \g372456/_3_  = ~n65833 ;
  assign \g372457/_3_  = ~n65839 ;
  assign \g372458/_3_  = ~n65845 ;
  assign \g372459/_3_  = ~n65851 ;
  assign \g372460/_3_  = ~n65857 ;
  assign \g372461/_3_  = ~n65863 ;
  assign \g372462/_3_  = ~n65869 ;
  assign \g372463/_3_  = ~n65875 ;
  assign \g372464/_3_  = ~n65881 ;
  assign \g372465/_3_  = ~n65887 ;
  assign \g372466/_3_  = ~n65893 ;
  assign \g372467/_3_  = ~n65899 ;
  assign \g372468/_3_  = ~n65905 ;
  assign \g372469/_3_  = ~n65911 ;
  assign \g372470/_3_  = ~n65917 ;
  assign \g372471/_3_  = ~n65923 ;
  assign \g372472/_3_  = ~n65929 ;
  assign \g372473/_3_  = ~n65935 ;
  assign \g372474/_3_  = ~n65941 ;
  assign \g372475/_3_  = ~n65947 ;
  assign \g372476/_3_  = ~n65953 ;
  assign \g372477/_3_  = ~n65959 ;
  assign \g372478/_3_  = ~n65965 ;
  assign \g372479/_3_  = ~n65971 ;
  assign \g372480/_3_  = ~n65977 ;
  assign \g372481/_3_  = ~n65983 ;
  assign \g372482/_3_  = ~n65989 ;
  assign \g372483/_3_  = ~n65995 ;
  assign \g372484/_3_  = ~n66001 ;
  assign \g372485/_3_  = ~n66007 ;
  assign \g372487/_3_  = ~n66013 ;
  assign \g372488/_3_  = ~n66019 ;
  assign \g372489/_3_  = ~n66025 ;
  assign \g372490/_3_  = ~n66031 ;
  assign \g372491/_3_  = ~n66037 ;
  assign \g372492/_3_  = ~n66043 ;
  assign \g372493/_3_  = ~n66049 ;
  assign \g372494/_3_  = ~n66055 ;
  assign \g372495/_3_  = ~n66061 ;
  assign \g372496/_3_  = ~n66067 ;
  assign \g372497/_3_  = ~n66073 ;
  assign \g372498/_3_  = ~n66079 ;
  assign \g372499/_3_  = ~n66085 ;
  assign \g372500/_3_  = ~n66091 ;
  assign \g372501/_3_  = ~n66097 ;
  assign \g372502/_3_  = ~n66103 ;
  assign \g372503/_3_  = ~n66109 ;
  assign \g372504/_3_  = ~n66115 ;
  assign \g372506/_3_  = ~n66121 ;
  assign \g372507/_3_  = ~n66127 ;
  assign \g372508/_3_  = ~n66133 ;
  assign \g372509/_3_  = ~n66139 ;
  assign \g372510/_3_  = ~n66145 ;
  assign \g372511/_3_  = ~n66151 ;
  assign \g372512/_3_  = ~n66157 ;
  assign \g372513/_3_  = ~n66163 ;
  assign \g372514/_3_  = ~n66169 ;
  assign \g372515/_3_  = ~n66175 ;
  assign \g372516/_3_  = ~n66181 ;
  assign \g372517/_3_  = ~n66187 ;
  assign \g372531/_3_  = ~n66190 ;
  assign \g372532/_3_  = ~n66193 ;
  assign \g372533/_3_  = ~n66195 ;
  assign \g374644/_0_  = ~n66204 ;
  assign \g374645/_0_  = ~n66213 ;
  assign \g374648/_0_  = ~n66222 ;
  assign \g374697/_0_  = ~n66232 ;
  assign \g374701/_0_  = ~n66242 ;
  assign \g374749/_0_  = ~n66251 ;
  assign \g374956/_0_  = ~n66260 ;
  assign \g374961/_0_  = ~n66270 ;
  assign \g374965/_0_  = ~n66285 ;
  assign \g374982/_0_  = ~n66294 ;
  assign \g375071/_0_  = ~n66305 ;
  assign \g375073/_0_  = ~n66315 ;
  assign \g375075/_0_  = ~n66326 ;
  assign \g375078/_0_  = ~n66336 ;
  assign \g375315/_3_  = ~n66339 ;
  assign \g375316/_3_  = ~n66342 ;
  assign \g376101/_0_  = ~n66355 ;
  assign \g376479/_0_  = ~n66369 ;
  assign \g377693/_0_  = ~n66378 ;
  assign \g377694/_0_  = ~n66388 ;
  assign \g377695/_0_  = ~n66398 ;
  assign \g377720/_0_  = ~n66407 ;
  assign \g377721/_0_  = ~n66417 ;
  assign \g377722/_0_  = ~n66427 ;
  assign \g378092/_3_  = ~n66430 ;
  assign \g378093/_3_  = ~n66433 ;
  assign \g378094/_3_  = ~n66436 ;
  assign \g378523/_0_  = ~n66437 ;
  assign \g378524/_0_  = ~n66438 ;
  assign \g382190/_0_  = ~n66447 ;
  assign \g382191/_0_  = ~n66456 ;
  assign \g382192/_0_  = ~n66465 ;
  assign \g382193/_0_  = ~n66474 ;
  assign \g382194/_0_  = ~n66483 ;
  assign \g382195/_0_  = ~n66492 ;
  assign \g382279/_0_  = ~n66502 ;
  assign \g382284/_0_  = ~n66512 ;
  assign \g382292/_0_  = ~n66524 ;
  assign \g382299/_0_  = ~n66535 ;
  assign \g382534/_0_  = ~n66548 ;
  assign \g382535/_0_  = ~n66560 ;
  assign \g382555/_0_  = ~n66569 ;
  assign \g382562/_0_  = ~n66578 ;
  assign \g382563/_0_  = ~n66587 ;
  assign \g382564/_0_  = ~n66596 ;
  assign \g382565/_0_  = ~n66606 ;
  assign \g382571/_0_  = ~n66616 ;
  assign \g382773/_3_  = ~n66619 ;
  assign \g382774/_3_  = ~n66622 ;
  assign \g382775/_3_  = ~n66625 ;
  assign \g383503/_2_  = ~n65813 ;
  assign \g383932/_2_  = ~n65791 ;
  assign \g384194/_0_  = ~n66634 ;
  assign \g384195/_0_  = ~n66643 ;
  assign \g384208/_0_  = ~n66654 ;
  assign \g385644/_0_  = ~n66663 ;
  assign \g385649/_0_  = ~n66672 ;
  assign \g385654/_0_  = ~n66681 ;
  assign \g385672/_0_  = ~n66696 ;
  assign \g385812/_0_  = ~n66707 ;
  assign \g385813/_0_  = ~n66718 ;
  assign \g385816/_0_  = ~n66730 ;
  assign \g385819/_0_  = ~n66741 ;
  assign \g386657/_0_  = ~n66752 ;
  assign \g386660/_0_  = ~n66763 ;
  assign \g386710/_0_  = ~n66774 ;
  assign \g386868/_0_  = ~n66785 ;
  assign \g387282/_0_  = ~n66797 ;
  assign \g387284/_0_  = ~n66809 ;
  assign \g387287/_0_  = ~n66822 ;
  assign \g387292/_0_  = ~n66836 ;
  assign \g387559/_0_  = ~n66845 ;
  assign \g387560/_0_  = ~n66854 ;
  assign \g387561/_0_  = ~n66863 ;
  assign \g387562/_0_  = ~n66872 ;
  assign \g387563/_0_  = ~n66881 ;
  assign \g387564/_0_  = ~n66890 ;
  assign \g387735/_0_  = ~n66899 ;
  assign \g387736/_0_  = ~n66909 ;
  assign \g387738/_0_  = ~n66918 ;
  assign \g387739/_0_  = ~n66928 ;
  assign \g387740/_0_  = ~n66937 ;
  assign \g387743/_0_  = ~n66946 ;
  assign \g387788/_0_  = ~n66956 ;
  assign \g387793/_0_  = ~n66965 ;
  assign \g387796/_0_  = ~n66975 ;
  assign \g387803/_0_  = ~n66984 ;
  assign \g388323/_3_  = ~n66987 ;
  assign \g388332/_3_  = ~n66990 ;
  assign \g388543/_0_  = ~n67003 ;
  assign \g388544/_0_  = ~n67016 ;
  assign \g388545/_0_  = ~n67028 ;
  assign \g388547/_0_  = ~n67042 ;
  assign \g388585/_0_  = ~n67051 ;
  assign \g388694/_0_  = ~n67059 ;
  assign \g388830/_0_  = ~n67068 ;
  assign \g388869/_0_  = ~n67079 ;
  assign \g388998/_0_  = ~n67088 ;
  assign \g389009/_0_  = ~n67096 ;
  assign \g389221/_0_  = ~n67102 ;
  assign \g389225/_0_  = ~n67107 ;
  assign \g389226/_0_  = ~n67112 ;
  assign \g389231/_0_  = ~n67116 ;
  assign \g389234/_0_  = ~n67121 ;
  assign \g389242/_0_  = ~n67126 ;
  assign \g389368/_2_  = ~n66635 ;
  assign \g389368/_2__syn_2  = n66635 ;
  assign \g389369/_2_  = ~n66626 ;
  assign \g389369/_2__syn_2  = n66626 ;
  assign \g389746/_0_  = ~n67135 ;
  assign \g389751/_0_  = ~n67145 ;
  assign \g389774/_0_  = ~n67154 ;
  assign \g389776/_0_  = ~n67163 ;
  assign \g389777/_0_  = ~n67172 ;
  assign \g389779/_0_  = ~n67181 ;
  assign \g389781/_0_  = ~n67190 ;
  assign \g389784/_0_  = ~n67199 ;
  assign \g389787/_0_  = ~n67208 ;
  assign \g389796/_0_  = ~n67217 ;
  assign \g389797/_0_  = ~n67226 ;
  assign \g389801/_0_  = ~n67235 ;
  assign \g390034/_0_  = ~n67244 ;
  assign \g390035/_0_  = ~n67254 ;
  assign \g390037/_0_  = ~n67263 ;
  assign \g390038/_0_  = ~n67272 ;
  assign \g390039/_0_  = ~n67281 ;
  assign \g390043/_0_  = ~n67290 ;
  assign \g390303/_3_  = ~n67293 ;
  assign \g390322/_3_  = ~n67296 ;
  assign \g390323/_3_  = ~n67299 ;
  assign \g390324/_3_  = ~n67302 ;
  assign \g390706/_0_  = ~n67306 ;
  assign \g390876/_0_  = ~n67310 ;
  assign \g390894/_0_  = ~n67314 ;
  assign \g390968/_0_  = ~n67318 ;
  assign \g391050/_0_  = ~n67322 ;
  assign \g391077/_0_  = ~n67326 ;
  assign \g392543/_3_  = ~n67329 ;
  assign \g392565/_3_  = ~n67332 ;
  assign \g392566/_3_  = ~n67335 ;
  assign \g394544/_3_  = ~n67338 ;
  assign \g394545/_3_  = ~n67341 ;
  assign \g394586/_3_  = ~n67344 ;
  assign \g395723/_0_  = ~n67353 ;
  assign \g395757/_0_  = ~n67362 ;
  assign \g395821/_0_  = ~n67371 ;
  assign \g395857/_0_  = ~n67380 ;
  assign \g395858/_0_  = ~n67389 ;
  assign \g395929/_0_  = ~n67398 ;
  assign \g396850/_3_  = ~n67401 ;
  assign \g396876/_3_  = ~n67404 ;
  assign \g396877/_3_  = ~n67407 ;
  assign \g397026/_1_  = ~n67045 ;
  assign \g397035/_1_  = ~n67082 ;
  assign \g397074/_1_  = ~n67062 ;
  assign \g397144/_1_  = ~n67052 ;
  assign \g397344/_1_  = ~n67089 ;
  assign \g397418/_1_  = ~n67072 ;
  assign \g397980/_0_  = n67412 ;
  assign \g398209/_0_  = ~n67419 ;
  assign \g398361/_0_  = n67424 ;
  assign \g398409/_0_  = n67429 ;
  assign \g398458/_0_  = n67434 ;
  assign \g398728/_0_  = n67439 ;
  assign \g401059/_0_  = ~n67441 ;
  assign \g401066/_0_  = ~n67444 ;
  assign \g401091/_0_  = ~n67446 ;
  assign \g401127/_0_  = ~n67448 ;
  assign \g401160/_0_  = ~n67450 ;
  assign \g401368/_0_  = ~n67453 ;
  assign \g401408/_0_  = ~n67455 ;
  assign \g401455/_0_  = ~n67458 ;
  assign \g401485/_0_  = ~n67460 ;
  assign \g401487/_0_  = ~n67462 ;
  assign \g401506/_0_  = ~n67465 ;
  assign \g401515/_0_  = ~n67468 ;
  assign \g401534/_0_  = ~n67471 ;
  assign \g401549/_0_  = ~n67474 ;
  assign \g401554/_0_  = ~n67477 ;
  assign \g401555/_0_  = ~n67480 ;
  assign \g401592/_0_  = ~n67483 ;
  assign \g401616/_0_  = ~n67486 ;
  assign \g401617/_0_  = ~n67489 ;
  assign \g401618/_0_  = ~n67492 ;
  assign \g401619/_0_  = ~n67495 ;
  assign \g401635/_0_  = ~n67498 ;
  assign \g401657/_0_  = ~n67500 ;
  assign \g401671/_0_  = ~n67503 ;
  assign \g401672/_0_  = ~n67506 ;
  assign \g401684/_0_  = ~n67508 ;
  assign \g401704/_0_  = ~n67511 ;
  assign \g401794/_0_  = ~n67514 ;
  assign \g401807/_0_  = ~n67517 ;
  assign \g401919/_0_  = ~n67519 ;
  assign \g401932/_0_  = ~n67522 ;
  assign \g401935/_0_  = ~n67525 ;
  assign \g401951/_0_  = ~n67528 ;
  assign \g401959/_0_  = ~n67531 ;
  assign \g401961/_0_  = ~n67534 ;
  assign \g401962/_0_  = ~n67537 ;
  assign \g401963/_0_  = ~n67540 ;
  assign \g401998/_0_  = ~n67543 ;
  assign \g402049/_0_  = ~n67546 ;
  assign \g402057/_0_  = ~n67549 ;
  assign \g402063/_0_  = ~n67552 ;
  assign \g402165/_0_  = ~n67555 ;
  assign \g402194/_0_  = ~n67558 ;
  assign \g402298/_0_  = ~n67561 ;
  assign \g402302/_0_  = ~n67564 ;
  assign \g402336/_0_  = ~n67567 ;
  assign \g402346/_0_  = ~n67570 ;
  assign \g402398/_0_  = ~n67573 ;
  assign \g402909/_0_  = ~n67578 ;
  assign \g402910/_0_  = n67583 ;
  assign \g402911/_0_  = n67586 ;
  assign \g402912/_0_  = n67591 ;
  assign \g402913/_0_  = n67596 ;
  assign \g402914/_0_  = ~n67602 ;
  assign \g403206/_3_  = ~n67605 ;
  assign \g427842/_1_  = ~n63451 ;
  assign \g427994/_0_  = ~n64059 ;
  assign \g428519/_1_  = ~n63427 ;
  assign \g429040/_1_  = ~n64101 ;
  assign \g429357/_0_  = ~n63380 ;
  assign \g429711/_1_  = ~n63350 ;
  assign \g440733/_0_  = ~n15809 ;
  assign \g440782/_0_  = ~n67619 ;
  assign \g441022/_0_  = ~n67638 ;
  assign \g441242/_0_  = ~n67657 ;
  assign \g441305/_0_  = ~n67676 ;
  assign \g441317/_0_  = ~n67695 ;
  assign \g441329/_0_  = ~n67714 ;
  assign \g441341/_0_  = ~n67733 ;
  assign \g441370/_0_  = ~n67752 ;
  assign \g441382/_0_  = ~n67771 ;
  assign \g441394/_0_  = ~n67790 ;
  assign \g441939/_0_  = ~n67809 ;
endmodule
