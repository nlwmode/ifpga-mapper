module top( \ac97_reset_pad_o__pad  , \dma_ack_i[0]_pad  , \dma_ack_i[1]_pad  , \dma_ack_i[2]_pad  , \dma_ack_i[3]_pad  , \dma_ack_i[4]_pad  , \dma_ack_i[5]_pad  , \dma_ack_i[6]_pad  , \dma_ack_i[7]_pad  , \dma_ack_i[8]_pad  , \dma_req_o[0]_pad  , \dma_req_o[1]_pad  , \dma_req_o[2]_pad  , \dma_req_o[3]_pad  , \dma_req_o[4]_pad  , \dma_req_o[5]_pad  , \dma_req_o[6]_pad  , \dma_req_o[7]_pad  , \dma_req_o[8]_pad  , \in_valid_s_reg[0]/NET0131  , \in_valid_s_reg[1]/NET0131  , \in_valid_s_reg[2]/NET0131  , suspended_o_pad , \u0_slt0_r_reg[0]/P0001  , \u0_slt0_r_reg[10]/P0001  , \u0_slt0_r_reg[11]/P0001  , \u0_slt0_r_reg[12]/P0001  , \u0_slt0_r_reg[13]/P0001  , \u0_slt0_r_reg[14]/P0001  , \u0_slt0_r_reg[1]/P0001  , \u0_slt0_r_reg[2]/P0001  , \u0_slt0_r_reg[3]/P0001  , \u0_slt0_r_reg[4]/P0001  , \u0_slt0_r_reg[5]/P0001  , \u0_slt0_r_reg[6]/P0001  , \u0_slt0_r_reg[7]/P0001  , \u0_slt0_r_reg[8]/P0001  , \u0_slt0_r_reg[9]/P0001  , \u0_slt1_r_reg[0]/P0001  , \u0_slt1_r_reg[10]/P0001  , \u0_slt1_r_reg[11]/P0001  , \u0_slt1_r_reg[12]/P0001  , \u0_slt1_r_reg[13]/P0001  , \u0_slt1_r_reg[14]/P0001  , \u0_slt1_r_reg[15]/P0001  , \u0_slt1_r_reg[16]/P0001  , \u0_slt1_r_reg[17]/P0001  , \u0_slt1_r_reg[18]/P0001  , \u0_slt1_r_reg[19]/P0001  , \u0_slt1_r_reg[1]/P0001  , \u0_slt1_r_reg[2]/P0001  , \u0_slt1_r_reg[3]/P0001  , \u0_slt1_r_reg[4]/P0001  , \u0_slt1_r_reg[5]/P0001  , \u0_slt1_r_reg[6]/P0001  , \u0_slt1_r_reg[7]/P0001  , \u0_slt1_r_reg[8]/P0001  , \u0_slt1_r_reg[9]/P0001  , \u0_slt2_r_reg[0]/P0001  , \u0_slt2_r_reg[10]/P0001  , \u0_slt2_r_reg[11]/P0001  , \u0_slt2_r_reg[12]/P0001  , \u0_slt2_r_reg[13]/P0001  , \u0_slt2_r_reg[14]/P0001  , \u0_slt2_r_reg[15]/P0001  , \u0_slt2_r_reg[16]/P0001  , \u0_slt2_r_reg[17]/P0001  , \u0_slt2_r_reg[18]/P0001  , \u0_slt2_r_reg[19]/P0001  , \u0_slt2_r_reg[1]/P0001  , \u0_slt2_r_reg[2]/P0001  , \u0_slt2_r_reg[3]/P0001  , \u0_slt2_r_reg[4]/P0001  , \u0_slt2_r_reg[5]/P0001  , \u0_slt2_r_reg[6]/P0001  , \u0_slt2_r_reg[7]/P0001  , \u0_slt2_r_reg[8]/P0001  , \u0_slt2_r_reg[9]/P0001  , \u0_slt3_r_reg[0]/P0001  , \u0_slt3_r_reg[10]/P0001  , \u0_slt3_r_reg[11]/P0001  , \u0_slt3_r_reg[12]/P0001  , \u0_slt3_r_reg[13]/P0001  , \u0_slt3_r_reg[14]/P0001  , \u0_slt3_r_reg[15]/P0001  , \u0_slt3_r_reg[16]/P0001  , \u0_slt3_r_reg[17]/P0001  , \u0_slt3_r_reg[18]/P0001  , \u0_slt3_r_reg[19]/P0001  , \u0_slt3_r_reg[1]/P0001  , \u0_slt3_r_reg[2]/P0001  , \u0_slt3_r_reg[3]/P0001  , \u0_slt3_r_reg[4]/P0001  , \u0_slt3_r_reg[5]/P0001  , \u0_slt3_r_reg[6]/P0001  , \u0_slt3_r_reg[7]/P0001  , \u0_slt3_r_reg[8]/P0001  , \u0_slt3_r_reg[9]/P0001  , \u0_slt4_r_reg[0]/P0001  , \u0_slt4_r_reg[10]/P0001  , \u0_slt4_r_reg[11]/P0001  , \u0_slt4_r_reg[12]/P0001  , \u0_slt4_r_reg[13]/P0001  , \u0_slt4_r_reg[14]/P0001  , \u0_slt4_r_reg[15]/P0001  , \u0_slt4_r_reg[16]/P0001  , \u0_slt4_r_reg[17]/P0001  , \u0_slt4_r_reg[18]/P0001  , \u0_slt4_r_reg[19]/P0001  , \u0_slt4_r_reg[1]/P0001  , \u0_slt4_r_reg[2]/P0001  , \u0_slt4_r_reg[3]/P0001  , \u0_slt4_r_reg[4]/P0001  , \u0_slt4_r_reg[5]/P0001  , \u0_slt4_r_reg[6]/P0001  , \u0_slt4_r_reg[7]/P0001  , \u0_slt4_r_reg[8]/P0001  , \u0_slt4_r_reg[9]/P0001  , \u0_slt5_r_reg[0]/P0001  , \u0_slt5_r_reg[10]/P0001  , \u0_slt5_r_reg[11]/P0001  , \u0_slt5_r_reg[12]/P0001  , \u0_slt5_r_reg[13]/P0001  , \u0_slt5_r_reg[14]/P0001  , \u0_slt5_r_reg[15]/P0001  , \u0_slt5_r_reg[16]/P0001  , \u0_slt5_r_reg[17]/P0001  , \u0_slt5_r_reg[18]/P0001  , \u0_slt5_r_reg[19]/P0001  , \u0_slt5_r_reg[1]/P0001  , \u0_slt5_r_reg[2]/P0001  , \u0_slt5_r_reg[3]/P0001  , \u0_slt5_r_reg[4]/P0001  , \u0_slt5_r_reg[5]/P0001  , \u0_slt5_r_reg[6]/P0001  , \u0_slt5_r_reg[7]/P0001  , \u0_slt5_r_reg[8]/P0001  , \u0_slt5_r_reg[9]/P0001  , \u0_slt6_r_reg[0]/P0001  , \u0_slt6_r_reg[10]/P0001  , \u0_slt6_r_reg[11]/P0001  , \u0_slt6_r_reg[12]/P0001  , \u0_slt6_r_reg[13]/P0001  , \u0_slt6_r_reg[14]/P0001  , \u0_slt6_r_reg[15]/P0001  , \u0_slt6_r_reg[16]/P0001  , \u0_slt6_r_reg[17]/P0001  , \u0_slt6_r_reg[18]/P0001  , \u0_slt6_r_reg[19]/P0001  , \u0_slt6_r_reg[1]/P0001  , \u0_slt6_r_reg[2]/P0001  , \u0_slt6_r_reg[3]/P0001  , \u0_slt6_r_reg[4]/P0001  , \u0_slt6_r_reg[5]/P0001  , \u0_slt6_r_reg[6]/P0001  , \u0_slt6_r_reg[7]/P0001  , \u0_slt6_r_reg[8]/P0001  , \u0_slt6_r_reg[9]/P0001  , \u0_slt7_r_reg[0]/P0001  , \u0_slt7_r_reg[10]/P0001  , \u0_slt7_r_reg[11]/P0001  , \u0_slt7_r_reg[12]/P0001  , \u0_slt7_r_reg[13]/P0001  , \u0_slt7_r_reg[14]/P0001  , \u0_slt7_r_reg[15]/P0001  , \u0_slt7_r_reg[16]/P0001  , \u0_slt7_r_reg[17]/P0001  , \u0_slt7_r_reg[18]/P0001  , \u0_slt7_r_reg[19]/P0001  , \u0_slt7_r_reg[1]/P0001  , \u0_slt7_r_reg[2]/P0001  , \u0_slt7_r_reg[3]/P0001  , \u0_slt7_r_reg[4]/P0001  , \u0_slt7_r_reg[5]/P0001  , \u0_slt7_r_reg[6]/P0001  , \u0_slt7_r_reg[7]/P0001  , \u0_slt7_r_reg[8]/P0001  , \u0_slt7_r_reg[9]/P0001  , \u0_slt8_r_reg[0]/P0001  , \u0_slt8_r_reg[10]/P0001  , \u0_slt8_r_reg[11]/P0001  , \u0_slt8_r_reg[12]/P0001  , \u0_slt8_r_reg[13]/P0001  , \u0_slt8_r_reg[14]/P0001  , \u0_slt8_r_reg[15]/P0001  , \u0_slt8_r_reg[16]/P0001  , \u0_slt8_r_reg[17]/P0001  , \u0_slt8_r_reg[18]/P0001  , \u0_slt8_r_reg[19]/P0001  , \u0_slt8_r_reg[1]/P0001  , \u0_slt8_r_reg[2]/P0001  , \u0_slt8_r_reg[3]/P0001  , \u0_slt8_r_reg[4]/P0001  , \u0_slt8_r_reg[5]/P0001  , \u0_slt8_r_reg[6]/P0001  , \u0_slt8_r_reg[7]/P0001  , \u0_slt8_r_reg[8]/P0001  , \u0_slt8_r_reg[9]/P0001  , \u0_slt9_r_reg[0]/P0001  , \u0_slt9_r_reg[10]/P0001  , \u0_slt9_r_reg[11]/P0001  , \u0_slt9_r_reg[12]/P0001  , \u0_slt9_r_reg[13]/P0001  , \u0_slt9_r_reg[14]/P0001  , \u0_slt9_r_reg[15]/P0001  , \u0_slt9_r_reg[16]/P0001  , \u0_slt9_r_reg[17]/P0001  , \u0_slt9_r_reg[18]/P0001  , \u0_slt9_r_reg[19]/P0001  , \u0_slt9_r_reg[1]/P0001  , \u0_slt9_r_reg[2]/P0001  , \u0_slt9_r_reg[3]/P0001  , \u0_slt9_r_reg[4]/P0001  , \u0_slt9_r_reg[5]/P0001  , \u0_slt9_r_reg[6]/P0001  , \u0_slt9_r_reg[7]/P0001  , \u0_slt9_r_reg[8]/P0001  , \u0_slt9_r_reg[9]/P0001  , \u10_din_tmp1_reg[0]/P0001  , \u10_din_tmp1_reg[10]/P0001  , \u10_din_tmp1_reg[11]/P0001  , \u10_din_tmp1_reg[12]/P0001  , \u10_din_tmp1_reg[13]/P0001  , \u10_din_tmp1_reg[14]/P0001  , \u10_din_tmp1_reg[15]/P0001  , \u10_din_tmp1_reg[1]/P0001  , \u10_din_tmp1_reg[2]/P0001  , \u10_din_tmp1_reg[3]/P0001  , \u10_din_tmp1_reg[4]/P0001  , \u10_din_tmp1_reg[5]/P0001  , \u10_din_tmp1_reg[6]/P0001  , \u10_din_tmp1_reg[7]/P0001  , \u10_din_tmp1_reg[8]/P0001  , \u10_din_tmp1_reg[9]/P0001  , \u10_dout_reg[0]/P0001  , \u10_dout_reg[10]/P0001  , \u10_dout_reg[11]/P0001  , \u10_dout_reg[12]/P0001  , \u10_dout_reg[13]/P0001  , \u10_dout_reg[14]/P0001  , \u10_dout_reg[15]/P0001  , \u10_dout_reg[16]/P0001  , \u10_dout_reg[17]/P0001  , \u10_dout_reg[18]/P0001  , \u10_dout_reg[19]/P0001  , \u10_dout_reg[1]/P0001  , \u10_dout_reg[20]/P0001  , \u10_dout_reg[21]/P0001  , \u10_dout_reg[22]/P0001  , \u10_dout_reg[23]/P0001  , \u10_dout_reg[24]/P0001  , \u10_dout_reg[25]/P0001  , \u10_dout_reg[26]/P0001  , \u10_dout_reg[27]/P0001  , \u10_dout_reg[28]/P0001  , \u10_dout_reg[29]/P0001  , \u10_dout_reg[2]/P0001  , \u10_dout_reg[30]/P0001  , \u10_dout_reg[31]/P0001  , \u10_dout_reg[3]/P0001  , \u10_dout_reg[4]/P0001  , \u10_dout_reg[5]/P0001  , \u10_dout_reg[6]/P0001  , \u10_dout_reg[7]/P0001  , \u10_dout_reg[8]/P0001  , \u10_dout_reg[9]/P0001  , \u10_empty_reg/P0001  , \u10_full_reg/NET0131  , \u10_mem_reg[0][0]/P0001  , \u10_mem_reg[0][10]/P0001  , \u10_mem_reg[0][11]/P0001  , \u10_mem_reg[0][12]/P0001  , \u10_mem_reg[0][13]/P0001  , \u10_mem_reg[0][14]/P0001  , \u10_mem_reg[0][15]/P0001  , \u10_mem_reg[0][16]/P0001  , \u10_mem_reg[0][17]/P0001  , \u10_mem_reg[0][18]/P0001  , \u10_mem_reg[0][19]/P0001  , \u10_mem_reg[0][1]/P0001  , \u10_mem_reg[0][20]/P0001  , \u10_mem_reg[0][21]/P0001  , \u10_mem_reg[0][22]/P0001  , \u10_mem_reg[0][23]/P0001  , \u10_mem_reg[0][24]/P0001  , \u10_mem_reg[0][25]/P0001  , \u10_mem_reg[0][26]/P0001  , \u10_mem_reg[0][27]/P0001  , \u10_mem_reg[0][28]/P0001  , \u10_mem_reg[0][29]/P0001  , \u10_mem_reg[0][2]/P0001  , \u10_mem_reg[0][30]/P0001  , \u10_mem_reg[0][31]/P0001  , \u10_mem_reg[0][3]/P0001  , \u10_mem_reg[0][4]/P0001  , \u10_mem_reg[0][5]/P0001  , \u10_mem_reg[0][6]/P0001  , \u10_mem_reg[0][7]/P0001  , \u10_mem_reg[0][8]/P0001  , \u10_mem_reg[0][9]/P0001  , \u10_mem_reg[1][0]/P0001  , \u10_mem_reg[1][10]/P0001  , \u10_mem_reg[1][11]/P0001  , \u10_mem_reg[1][12]/P0001  , \u10_mem_reg[1][13]/P0001  , \u10_mem_reg[1][14]/P0001  , \u10_mem_reg[1][15]/P0001  , \u10_mem_reg[1][16]/P0001  , \u10_mem_reg[1][17]/P0001  , \u10_mem_reg[1][18]/P0001  , \u10_mem_reg[1][19]/P0001  , \u10_mem_reg[1][1]/P0001  , \u10_mem_reg[1][20]/P0001  , \u10_mem_reg[1][21]/P0001  , \u10_mem_reg[1][22]/P0001  , \u10_mem_reg[1][23]/P0001  , \u10_mem_reg[1][24]/P0001  , \u10_mem_reg[1][25]/P0001  , \u10_mem_reg[1][26]/P0001  , \u10_mem_reg[1][27]/P0001  , \u10_mem_reg[1][28]/P0001  , \u10_mem_reg[1][29]/P0001  , \u10_mem_reg[1][2]/P0001  , \u10_mem_reg[1][30]/P0001  , \u10_mem_reg[1][31]/P0001  , \u10_mem_reg[1][3]/P0001  , \u10_mem_reg[1][4]/P0001  , \u10_mem_reg[1][5]/P0001  , \u10_mem_reg[1][6]/P0001  , \u10_mem_reg[1][7]/P0001  , \u10_mem_reg[1][8]/P0001  , \u10_mem_reg[1][9]/P0001  , \u10_mem_reg[2][0]/P0001  , \u10_mem_reg[2][10]/P0001  , \u10_mem_reg[2][11]/P0001  , \u10_mem_reg[2][12]/P0001  , \u10_mem_reg[2][13]/P0001  , \u10_mem_reg[2][14]/P0001  , \u10_mem_reg[2][15]/P0001  , \u10_mem_reg[2][16]/P0001  , \u10_mem_reg[2][17]/P0001  , \u10_mem_reg[2][18]/P0001  , \u10_mem_reg[2][19]/P0001  , \u10_mem_reg[2][1]/P0001  , \u10_mem_reg[2][20]/P0001  , \u10_mem_reg[2][21]/P0001  , \u10_mem_reg[2][22]/P0001  , \u10_mem_reg[2][23]/P0001  , \u10_mem_reg[2][24]/P0001  , \u10_mem_reg[2][25]/P0001  , \u10_mem_reg[2][26]/P0001  , \u10_mem_reg[2][27]/P0001  , \u10_mem_reg[2][28]/P0001  , \u10_mem_reg[2][29]/P0001  , \u10_mem_reg[2][2]/P0001  , \u10_mem_reg[2][30]/P0001  , \u10_mem_reg[2][31]/P0001  , \u10_mem_reg[2][3]/P0001  , \u10_mem_reg[2][4]/P0001  , \u10_mem_reg[2][5]/P0001  , \u10_mem_reg[2][6]/P0001  , \u10_mem_reg[2][7]/P0001  , \u10_mem_reg[2][8]/P0001  , \u10_mem_reg[2][9]/P0001  , \u10_mem_reg[3][0]/P0001  , \u10_mem_reg[3][10]/P0001  , \u10_mem_reg[3][11]/P0001  , \u10_mem_reg[3][12]/P0001  , \u10_mem_reg[3][13]/P0001  , \u10_mem_reg[3][14]/P0001  , \u10_mem_reg[3][15]/P0001  , \u10_mem_reg[3][16]/P0001  , \u10_mem_reg[3][17]/P0001  , \u10_mem_reg[3][18]/P0001  , \u10_mem_reg[3][19]/P0001  , \u10_mem_reg[3][1]/P0001  , \u10_mem_reg[3][20]/P0001  , \u10_mem_reg[3][21]/P0001  , \u10_mem_reg[3][22]/P0001  , \u10_mem_reg[3][23]/P0001  , \u10_mem_reg[3][24]/P0001  , \u10_mem_reg[3][25]/P0001  , \u10_mem_reg[3][26]/P0001  , \u10_mem_reg[3][27]/P0001  , \u10_mem_reg[3][28]/P0001  , \u10_mem_reg[3][29]/P0001  , \u10_mem_reg[3][2]/P0001  , \u10_mem_reg[3][30]/P0001  , \u10_mem_reg[3][31]/P0001  , \u10_mem_reg[3][3]/P0001  , \u10_mem_reg[3][4]/P0001  , \u10_mem_reg[3][5]/P0001  , \u10_mem_reg[3][6]/P0001  , \u10_mem_reg[3][7]/P0001  , \u10_mem_reg[3][8]/P0001  , \u10_mem_reg[3][9]/P0001  , \u10_rp_reg[0]/P0001  , \u10_rp_reg[1]/P0001  , \u10_rp_reg[2]/P0001  , \u10_status_reg[0]/P0001  , \u10_status_reg[1]/P0001  , \u10_wp_reg[0]/NET0131  , \u10_wp_reg[1]/P0001  , \u10_wp_reg[2]/P0001  , \u10_wp_reg[3]/P0001  , \u11_din_tmp1_reg[0]/P0001  , \u11_din_tmp1_reg[10]/P0001  , \u11_din_tmp1_reg[11]/P0001  , \u11_din_tmp1_reg[12]/P0001  , \u11_din_tmp1_reg[13]/P0001  , \u11_din_tmp1_reg[14]/P0001  , \u11_din_tmp1_reg[15]/P0001  , \u11_din_tmp1_reg[1]/P0001  , \u11_din_tmp1_reg[2]/P0001  , \u11_din_tmp1_reg[3]/P0001  , \u11_din_tmp1_reg[4]/P0001  , \u11_din_tmp1_reg[5]/P0001  , \u11_din_tmp1_reg[6]/P0001  , \u11_din_tmp1_reg[7]/P0001  , \u11_din_tmp1_reg[8]/P0001  , \u11_din_tmp1_reg[9]/P0001  , \u11_dout_reg[0]/P0001  , \u11_dout_reg[10]/P0001  , \u11_dout_reg[11]/P0001  , \u11_dout_reg[12]/P0001  , \u11_dout_reg[13]/P0001  , \u11_dout_reg[14]/P0001  , \u11_dout_reg[15]/P0001  , \u11_dout_reg[16]/P0001  , \u11_dout_reg[17]/P0001  , \u11_dout_reg[18]/P0001  , \u11_dout_reg[19]/P0001  , \u11_dout_reg[1]/P0001  , \u11_dout_reg[20]/P0001  , \u11_dout_reg[21]/P0001  , \u11_dout_reg[22]/P0001  , \u11_dout_reg[23]/P0001  , \u11_dout_reg[24]/P0001  , \u11_dout_reg[25]/P0001  , \u11_dout_reg[26]/P0001  , \u11_dout_reg[27]/P0001  , \u11_dout_reg[28]/P0001  , \u11_dout_reg[29]/P0001  , \u11_dout_reg[2]/P0001  , \u11_dout_reg[30]/P0001  , \u11_dout_reg[31]/P0001  , \u11_dout_reg[3]/P0001  , \u11_dout_reg[4]/P0001  , \u11_dout_reg[5]/P0001  , \u11_dout_reg[6]/P0001  , \u11_dout_reg[7]/P0001  , \u11_dout_reg[8]/P0001  , \u11_dout_reg[9]/P0001  , \u11_empty_reg/P0001  , \u11_full_reg/NET0131  , \u11_mem_reg[0][0]/P0001  , \u11_mem_reg[0][10]/P0001  , \u11_mem_reg[0][11]/P0001  , \u11_mem_reg[0][12]/P0001  , \u11_mem_reg[0][13]/P0001  , \u11_mem_reg[0][14]/P0001  , \u11_mem_reg[0][15]/P0001  , \u11_mem_reg[0][16]/P0001  , \u11_mem_reg[0][17]/P0001  , \u11_mem_reg[0][18]/P0001  , \u11_mem_reg[0][19]/P0001  , \u11_mem_reg[0][1]/P0001  , \u11_mem_reg[0][20]/P0001  , \u11_mem_reg[0][21]/P0001  , \u11_mem_reg[0][22]/P0001  , \u11_mem_reg[0][23]/P0001  , \u11_mem_reg[0][24]/P0001  , \u11_mem_reg[0][25]/P0001  , \u11_mem_reg[0][26]/P0001  , \u11_mem_reg[0][27]/P0001  , \u11_mem_reg[0][28]/P0001  , \u11_mem_reg[0][29]/P0001  , \u11_mem_reg[0][2]/P0001  , \u11_mem_reg[0][30]/P0001  , \u11_mem_reg[0][31]/P0001  , \u11_mem_reg[0][3]/P0001  , \u11_mem_reg[0][4]/P0001  , \u11_mem_reg[0][5]/P0001  , \u11_mem_reg[0][6]/P0001  , \u11_mem_reg[0][7]/P0001  , \u11_mem_reg[0][8]/P0001  , \u11_mem_reg[0][9]/P0001  , \u11_mem_reg[1][0]/P0001  , \u11_mem_reg[1][10]/P0001  , \u11_mem_reg[1][11]/P0001  , \u11_mem_reg[1][12]/P0001  , \u11_mem_reg[1][13]/P0001  , \u11_mem_reg[1][14]/P0001  , \u11_mem_reg[1][15]/P0001  , \u11_mem_reg[1][16]/P0001  , \u11_mem_reg[1][17]/P0001  , \u11_mem_reg[1][18]/P0001  , \u11_mem_reg[1][19]/P0001  , \u11_mem_reg[1][1]/P0001  , \u11_mem_reg[1][20]/P0001  , \u11_mem_reg[1][21]/P0001  , \u11_mem_reg[1][22]/P0001  , \u11_mem_reg[1][23]/P0001  , \u11_mem_reg[1][24]/P0001  , \u11_mem_reg[1][25]/P0001  , \u11_mem_reg[1][26]/P0001  , \u11_mem_reg[1][27]/P0001  , \u11_mem_reg[1][28]/P0001  , \u11_mem_reg[1][29]/P0001  , \u11_mem_reg[1][2]/P0001  , \u11_mem_reg[1][30]/P0001  , \u11_mem_reg[1][31]/P0001  , \u11_mem_reg[1][3]/P0001  , \u11_mem_reg[1][4]/P0001  , \u11_mem_reg[1][5]/P0001  , \u11_mem_reg[1][6]/P0001  , \u11_mem_reg[1][7]/P0001  , \u11_mem_reg[1][8]/P0001  , \u11_mem_reg[1][9]/P0001  , \u11_mem_reg[2][0]/P0001  , \u11_mem_reg[2][10]/P0001  , \u11_mem_reg[2][11]/P0001  , \u11_mem_reg[2][12]/P0001  , \u11_mem_reg[2][13]/P0001  , \u11_mem_reg[2][14]/P0001  , \u11_mem_reg[2][15]/P0001  , \u11_mem_reg[2][16]/P0001  , \u11_mem_reg[2][17]/P0001  , \u11_mem_reg[2][18]/P0001  , \u11_mem_reg[2][19]/P0001  , \u11_mem_reg[2][1]/P0001  , \u11_mem_reg[2][20]/P0001  , \u11_mem_reg[2][21]/P0001  , \u11_mem_reg[2][22]/P0001  , \u11_mem_reg[2][23]/P0001  , \u11_mem_reg[2][24]/P0001  , \u11_mem_reg[2][25]/P0001  , \u11_mem_reg[2][26]/P0001  , \u11_mem_reg[2][27]/P0001  , \u11_mem_reg[2][28]/P0001  , \u11_mem_reg[2][29]/P0001  , \u11_mem_reg[2][2]/P0001  , \u11_mem_reg[2][30]/P0001  , \u11_mem_reg[2][31]/P0001  , \u11_mem_reg[2][3]/P0001  , \u11_mem_reg[2][4]/P0001  , \u11_mem_reg[2][5]/P0001  , \u11_mem_reg[2][6]/P0001  , \u11_mem_reg[2][7]/P0001  , \u11_mem_reg[2][8]/P0001  , \u11_mem_reg[2][9]/P0001  , \u11_mem_reg[3][0]/P0001  , \u11_mem_reg[3][10]/P0001  , \u11_mem_reg[3][11]/P0001  , \u11_mem_reg[3][12]/P0001  , \u11_mem_reg[3][13]/P0001  , \u11_mem_reg[3][14]/P0001  , \u11_mem_reg[3][15]/P0001  , \u11_mem_reg[3][16]/P0001  , \u11_mem_reg[3][17]/P0001  , \u11_mem_reg[3][18]/P0001  , \u11_mem_reg[3][19]/P0001  , \u11_mem_reg[3][1]/P0001  , \u11_mem_reg[3][20]/P0001  , \u11_mem_reg[3][21]/P0001  , \u11_mem_reg[3][22]/P0001  , \u11_mem_reg[3][23]/P0001  , \u11_mem_reg[3][24]/P0001  , \u11_mem_reg[3][25]/P0001  , \u11_mem_reg[3][26]/P0001  , \u11_mem_reg[3][27]/P0001  , \u11_mem_reg[3][28]/P0001  , \u11_mem_reg[3][29]/P0001  , \u11_mem_reg[3][2]/P0001  , \u11_mem_reg[3][30]/P0001  , \u11_mem_reg[3][31]/P0001  , \u11_mem_reg[3][3]/P0001  , \u11_mem_reg[3][4]/P0001  , \u11_mem_reg[3][5]/P0001  , \u11_mem_reg[3][6]/P0001  , \u11_mem_reg[3][7]/P0001  , \u11_mem_reg[3][8]/P0001  , \u11_mem_reg[3][9]/P0001  , \u11_rp_reg[0]/P0001  , \u11_rp_reg[1]/P0001  , \u11_rp_reg[2]/P0001  , \u11_status_reg[0]/P0001  , \u11_status_reg[1]/P0001  , \u11_wp_reg[0]/NET0131  , \u11_wp_reg[1]/P0001  , \u11_wp_reg[2]/P0001  , \u11_wp_reg[3]/P0001  , \u12_dout_reg[0]/P0001  , \u12_dout_reg[10]/P0001  , \u12_dout_reg[11]/P0001  , \u12_dout_reg[12]/P0001  , \u12_dout_reg[13]/P0001  , \u12_dout_reg[14]/P0001  , \u12_dout_reg[15]/P0001  , \u12_dout_reg[16]/P0001  , \u12_dout_reg[17]/P0001  , \u12_dout_reg[18]/P0001  , \u12_dout_reg[19]/P0001  , \u12_dout_reg[1]/P0001  , \u12_dout_reg[20]/P0001  , \u12_dout_reg[21]/P0001  , \u12_dout_reg[22]/P0001  , \u12_dout_reg[23]/P0001  , \u12_dout_reg[24]/P0001  , \u12_dout_reg[25]/P0001  , \u12_dout_reg[26]/P0001  , \u12_dout_reg[27]/P0001  , \u12_dout_reg[28]/P0001  , \u12_dout_reg[29]/P0001  , \u12_dout_reg[2]/P0001  , \u12_dout_reg[30]/P0001  , \u12_dout_reg[31]/P0001  , \u12_dout_reg[3]/P0001  , \u12_dout_reg[4]/P0001  , \u12_dout_reg[5]/P0001  , \u12_dout_reg[6]/P0001  , \u12_dout_reg[7]/P0001  , \u12_dout_reg[8]/P0001  , \u12_dout_reg[9]/P0001  , \u12_i3_re_reg/NET0131  , \u12_i4_re_reg/P0001  , \u12_i6_re_reg/NET0131  , \u12_o3_we_reg/P0001  , \u12_o4_we_reg/P0001  , \u12_o6_we_reg/P0001  , \u12_o7_we_reg/P0001  , \u12_o8_we_reg/P0001  , \u12_o9_we_reg/P0001  , \u12_re1_reg/P0001  , \u12_re2_reg/NET0131  , \u12_rf_we_reg/P0001  , \u12_we1_reg/P0001  , \u12_we2_reg/P0001  , \u13_ac97_rst_force_reg/P0001  , \u13_crac_dout_r_reg[0]/P0001  , \u13_crac_dout_r_reg[10]/P0001  , \u13_crac_dout_r_reg[11]/P0001  , \u13_crac_dout_r_reg[12]/P0001  , \u13_crac_dout_r_reg[13]/P0001  , \u13_crac_dout_r_reg[14]/P0001  , \u13_crac_dout_r_reg[15]/P0001  , \u13_crac_dout_r_reg[1]/P0001  , \u13_crac_dout_r_reg[2]/P0001  , \u13_crac_dout_r_reg[3]/P0001  , \u13_crac_dout_r_reg[4]/P0001  , \u13_crac_dout_r_reg[5]/P0001  , \u13_crac_dout_r_reg[6]/P0001  , \u13_crac_dout_r_reg[7]/P0001  , \u13_crac_dout_r_reg[8]/P0001  , \u13_crac_dout_r_reg[9]/P0001  , \u13_crac_r_reg[0]/NET0131  , \u13_crac_r_reg[1]/NET0131  , \u13_crac_r_reg[2]/NET0131  , \u13_crac_r_reg[3]/NET0131  , \u13_crac_r_reg[4]/NET0131  , \u13_crac_r_reg[5]/NET0131  , \u13_crac_r_reg[6]/NET0131  , \u13_crac_r_reg[7]/NET0131  , \u13_icc_r_reg[0]/NET0131  , \u13_icc_r_reg[10]/NET0131  , \u13_icc_r_reg[11]/NET0131  , \u13_icc_r_reg[12]/NET0131  , \u13_icc_r_reg[13]/NET0131  , \u13_icc_r_reg[14]/NET0131  , \u13_icc_r_reg[15]/NET0131  , \u13_icc_r_reg[16]/NET0131  , \u13_icc_r_reg[17]/NET0131  , \u13_icc_r_reg[18]/NET0131  , \u13_icc_r_reg[19]/NET0131  , \u13_icc_r_reg[1]/NET0131  , \u13_icc_r_reg[20]/NET0131  , \u13_icc_r_reg[21]/NET0131  , \u13_icc_r_reg[22]/NET0131  , \u13_icc_r_reg[23]/NET0131  , \u13_icc_r_reg[2]/NET0131  , \u13_icc_r_reg[3]/NET0131  , \u13_icc_r_reg[4]/NET0131  , \u13_icc_r_reg[5]/NET0131  , \u13_icc_r_reg[6]/NET0131  , \u13_icc_r_reg[7]/NET0131  , \u13_icc_r_reg[8]/NET0131  , \u13_icc_r_reg[9]/NET0131  , \u13_intm_r_reg[0]/NET0131  , \u13_intm_r_reg[10]/NET0131  , \u13_intm_r_reg[11]/NET0131  , \u13_intm_r_reg[12]/NET0131  , \u13_intm_r_reg[13]/NET0131  , \u13_intm_r_reg[14]/NET0131  , \u13_intm_r_reg[15]/NET0131  , \u13_intm_r_reg[16]/NET0131  , \u13_intm_r_reg[17]/NET0131  , \u13_intm_r_reg[18]/NET0131  , \u13_intm_r_reg[19]/NET0131  , \u13_intm_r_reg[1]/NET0131  , \u13_intm_r_reg[20]/NET0131  , \u13_intm_r_reg[21]/NET0131  , \u13_intm_r_reg[22]/NET0131  , \u13_intm_r_reg[23]/NET0131  , \u13_intm_r_reg[24]/NET0131  , \u13_intm_r_reg[25]/NET0131  , \u13_intm_r_reg[26]/NET0131  , \u13_intm_r_reg[27]/NET0131  , \u13_intm_r_reg[28]/NET0131  , \u13_intm_r_reg[2]/NET0131  , \u13_intm_r_reg[3]/NET0131  , \u13_intm_r_reg[4]/NET0131  , \u13_intm_r_reg[5]/NET0131  , \u13_intm_r_reg[6]/NET0131  , \u13_intm_r_reg[7]/NET0131  , \u13_intm_r_reg[8]/NET0131  , \u13_intm_r_reg[9]/NET0131  , \u13_ints_r_reg[0]/NET0131  , \u13_ints_r_reg[10]/NET0131  , \u13_ints_r_reg[11]/NET0131  , \u13_ints_r_reg[12]/NET0131  , \u13_ints_r_reg[13]/NET0131  , \u13_ints_r_reg[14]/NET0131  , \u13_ints_r_reg[15]/NET0131  , \u13_ints_r_reg[16]/NET0131  , \u13_ints_r_reg[17]/NET0131  , \u13_ints_r_reg[18]/NET0131  , \u13_ints_r_reg[19]/NET0131  , \u13_ints_r_reg[1]/NET0131  , \u13_ints_r_reg[20]/NET0131  , \u13_ints_r_reg[21]/NET0131  , \u13_ints_r_reg[22]/NET0131  , \u13_ints_r_reg[23]/NET0131  , \u13_ints_r_reg[24]/NET0131  , \u13_ints_r_reg[25]/NET0131  , \u13_ints_r_reg[26]/NET0131  , \u13_ints_r_reg[27]/NET0131  , \u13_ints_r_reg[28]/NET0131  , \u13_ints_r_reg[2]/NET0131  , \u13_ints_r_reg[3]/NET0131  , \u13_ints_r_reg[4]/NET0131  , \u13_ints_r_reg[5]/NET0131  , \u13_ints_r_reg[6]/NET0131  , \u13_ints_r_reg[7]/NET0131  , \u13_ints_r_reg[8]/NET0131  , \u13_ints_r_reg[9]/NET0131  , \u13_occ0_r_reg[0]/NET0131  , \u13_occ0_r_reg[10]/NET0131  , \u13_occ0_r_reg[11]/NET0131  , \u13_occ0_r_reg[12]/NET0131  , \u13_occ0_r_reg[13]/NET0131  , \u13_occ0_r_reg[14]/NET0131  , \u13_occ0_r_reg[15]/NET0131  , \u13_occ0_r_reg[16]/NET0131  , \u13_occ0_r_reg[17]/NET0131  , \u13_occ0_r_reg[18]/NET0131  , \u13_occ0_r_reg[19]/NET0131  , \u13_occ0_r_reg[1]/NET0131  , \u13_occ0_r_reg[20]/NET0131  , \u13_occ0_r_reg[21]/NET0131  , \u13_occ0_r_reg[22]/NET0131  , \u13_occ0_r_reg[23]/NET0131  , \u13_occ0_r_reg[24]/NET0131  , \u13_occ0_r_reg[25]/NET0131  , \u13_occ0_r_reg[26]/NET0131  , \u13_occ0_r_reg[27]/NET0131  , \u13_occ0_r_reg[28]/NET0131  , \u13_occ0_r_reg[29]/NET0131  , \u13_occ0_r_reg[2]/NET0131  , \u13_occ0_r_reg[30]/NET0131  , \u13_occ0_r_reg[31]/NET0131  , \u13_occ0_r_reg[3]/NET0131  , \u13_occ0_r_reg[4]/NET0131  , \u13_occ0_r_reg[5]/NET0131  , \u13_occ0_r_reg[6]/NET0131  , \u13_occ0_r_reg[7]/NET0131  , \u13_occ0_r_reg[8]/NET0131  , \u13_occ0_r_reg[9]/NET0131  , \u13_occ1_r_reg[0]/NET0131  , \u13_occ1_r_reg[10]/NET0131  , \u13_occ1_r_reg[11]/NET0131  , \u13_occ1_r_reg[12]/NET0131  , \u13_occ1_r_reg[13]/NET0131  , \u13_occ1_r_reg[14]/NET0131  , \u13_occ1_r_reg[15]/NET0131  , \u13_occ1_r_reg[1]/NET0131  , \u13_occ1_r_reg[2]/NET0131  , \u13_occ1_r_reg[3]/NET0131  , \u13_occ1_r_reg[4]/NET0131  , \u13_occ1_r_reg[5]/NET0131  , \u13_occ1_r_reg[6]/NET0131  , \u13_occ1_r_reg[7]/NET0131  , \u13_occ1_r_reg[8]/NET0131  , \u13_occ1_r_reg[9]/NET0131  , \u13_resume_req_reg/P0001  , \u14_crac_valid_r_reg/P0001  , \u14_crac_wr_r_reg/P0001  , \u14_u0_en_out_l2_reg/P0001  , \u14_u0_en_out_l_reg/NET0131  , \u14_u0_full_empty_r_reg/P0001  , \u14_u1_en_out_l2_reg/P0001  , \u14_u1_en_out_l_reg/NET0131  , \u14_u1_full_empty_r_reg/P0001  , \u14_u2_en_out_l2_reg/P0001  , \u14_u2_en_out_l_reg/NET0131  , \u14_u2_full_empty_r_reg/P0001  , \u14_u3_en_out_l2_reg/P0001  , \u14_u3_en_out_l_reg/NET0131  , \u14_u3_full_empty_r_reg/P0001  , \u14_u4_en_out_l2_reg/P0001  , \u14_u4_en_out_l_reg/NET0131  , \u14_u4_full_empty_r_reg/P0001  , \u14_u5_en_out_l2_reg/P0001  , \u14_u5_en_out_l_reg/NET0131  , \u14_u5_full_empty_r_reg/P0001  , \u14_u6_en_out_l2_reg/P0001  , \u14_u6_en_out_l_reg/NET0131  , \u14_u6_full_empty_r_reg/P0001  , \u14_u7_en_out_l2_reg/P0001  , \u14_u7_en_out_l_reg/NET0131  , \u14_u7_full_empty_r_reg/P0001  , \u14_u8_en_out_l2_reg/P0001  , \u14_u8_en_out_l_reg/NET0131  , \u14_u8_full_empty_r_reg/P0001  , \u15_crac_din_reg[0]/NET0131  , \u15_crac_din_reg[10]/NET0131  , \u15_crac_din_reg[11]/NET0131  , \u15_crac_din_reg[12]/NET0131  , \u15_crac_din_reg[13]/NET0131  , \u15_crac_din_reg[14]/NET0131  , \u15_crac_din_reg[15]/NET0131  , \u15_crac_din_reg[1]/NET0131  , \u15_crac_din_reg[2]/NET0131  , \u15_crac_din_reg[3]/NET0131  , \u15_crac_din_reg[4]/NET0131  , \u15_crac_din_reg[5]/NET0131  , \u15_crac_din_reg[6]/NET0131  , \u15_crac_din_reg[7]/NET0131  , \u15_crac_din_reg[8]/NET0131  , \u15_crac_din_reg[9]/NET0131  , \u15_crac_rd_done_reg/P0001  , \u15_crac_rd_reg/NET0131  , \u15_crac_we_r_reg/P0001  , \u15_crac_wr_reg/NET0131  , \u15_rdd1_reg/NET0131  , \u15_rdd2_reg/NET0131  , \u15_rdd3_reg/NET0131  , \u15_valid_r_reg/P0001  , \u16_u0_dma_req_r1_reg/P0001  , \u16_u1_dma_req_r1_reg/P0001  , \u16_u2_dma_req_r1_reg/P0001  , \u16_u3_dma_req_r1_reg/P0001  , \u16_u4_dma_req_r1_reg/P0001  , \u16_u5_dma_req_r1_reg/P0001  , \u16_u6_dma_req_r1_reg/P0001  , \u16_u7_dma_req_r1_reg/P0001  , \u16_u8_dma_req_r1_reg/P0001  , \u17_int_set_reg[0]/NET0131  , \u17_int_set_reg[1]/NET0131  , \u17_int_set_reg[2]/NET0131  , \u18_int_set_reg[0]/NET0131  , \u18_int_set_reg[1]/NET0131  , \u18_int_set_reg[2]/NET0131  , \u19_int_set_reg[0]/NET0131  , \u19_int_set_reg[1]/NET0131  , \u19_int_set_reg[2]/NET0131  , \u1_slt0_reg[11]/P0001  , \u1_slt0_reg[12]/P0001  , \u1_slt0_reg[15]/P0001  , \u1_slt0_reg[9]/P0001  , \u1_slt1_reg[10]/P0001  , \u1_slt1_reg[11]/P0001  , \u1_slt1_reg[5]/P0001  , \u1_slt1_reg[6]/P0001  , \u1_slt1_reg[7]/P0001  , \u1_slt1_reg[8]/P0001  , \u1_slt3_reg[0]/P0001  , \u1_slt3_reg[10]/P0001  , \u1_slt3_reg[11]/P0001  , \u1_slt3_reg[12]/P0001  , \u1_slt3_reg[13]/P0001  , \u1_slt3_reg[14]/P0001  , \u1_slt3_reg[15]/P0001  , \u1_slt3_reg[16]/P0001  , \u1_slt3_reg[17]/P0001  , \u1_slt3_reg[18]/P0001  , \u1_slt3_reg[19]/P0001  , \u1_slt3_reg[1]/P0001  , \u1_slt3_reg[2]/P0001  , \u1_slt3_reg[3]/P0001  , \u1_slt3_reg[4]/P0001  , \u1_slt3_reg[5]/P0001  , \u1_slt3_reg[6]/P0001  , \u1_slt3_reg[7]/P0001  , \u1_slt3_reg[8]/P0001  , \u1_slt3_reg[9]/P0001  , \u1_slt4_reg[0]/P0001  , \u1_slt4_reg[10]/P0001  , \u1_slt4_reg[11]/P0001  , \u1_slt4_reg[12]/P0001  , \u1_slt4_reg[13]/P0001  , \u1_slt4_reg[14]/P0001  , \u1_slt4_reg[15]/P0001  , \u1_slt4_reg[16]/P0001  , \u1_slt4_reg[17]/P0001  , \u1_slt4_reg[18]/P0001  , \u1_slt4_reg[19]/P0001  , \u1_slt4_reg[1]/P0001  , \u1_slt4_reg[2]/P0001  , \u1_slt4_reg[3]/P0001  , \u1_slt4_reg[4]/P0001  , \u1_slt4_reg[5]/P0001  , \u1_slt4_reg[6]/P0001  , \u1_slt4_reg[7]/P0001  , \u1_slt4_reg[8]/P0001  , \u1_slt4_reg[9]/P0001  , \u1_slt6_reg[0]/P0001  , \u1_slt6_reg[10]/P0001  , \u1_slt6_reg[11]/P0001  , \u1_slt6_reg[12]/P0001  , \u1_slt6_reg[13]/P0001  , \u1_slt6_reg[14]/P0001  , \u1_slt6_reg[15]/P0001  , \u1_slt6_reg[16]/P0001  , \u1_slt6_reg[17]/P0001  , \u1_slt6_reg[18]/P0001  , \u1_slt6_reg[19]/P0001  , \u1_slt6_reg[1]/P0001  , \u1_slt6_reg[2]/P0001  , \u1_slt6_reg[3]/P0001  , \u1_slt6_reg[4]/P0001  , \u1_slt6_reg[5]/P0001  , \u1_slt6_reg[6]/P0001  , \u1_slt6_reg[7]/P0001  , \u1_slt6_reg[8]/P0001  , \u1_slt6_reg[9]/P0001  , \u1_sr_reg[10]/P0001  , \u1_sr_reg[11]/P0001  , \u1_sr_reg[12]/P0001  , \u1_sr_reg[15]/P0001  , \u1_sr_reg[5]/P0001  , \u1_sr_reg[6]/P0001  , \u1_sr_reg[7]/P0001  , \u1_sr_reg[8]/P0001  , \u1_sr_reg[9]/P0001  , \u20_int_set_reg[0]/NET0131  , \u20_int_set_reg[1]/NET0131  , \u20_int_set_reg[2]/NET0131  , \u21_int_set_reg[0]/NET0131  , \u21_int_set_reg[1]/NET0131  , \u21_int_set_reg[2]/NET0131  , \u22_int_set_reg[0]/NET0131  , \u22_int_set_reg[1]/NET0131  , \u22_int_set_reg[2]/NET0131  , \u23_int_set_reg[0]/NET0131  , \u23_int_set_reg[1]/NET0131  , \u23_int_set_reg[2]/NET0131  , \u24_int_set_reg[0]/NET0131  , \u24_int_set_reg[1]/NET0131  , \u24_int_set_reg[2]/NET0131  , \u25_int_set_reg[0]/NET0131  , \u25_int_set_reg[1]/NET0131  , \u25_int_set_reg[2]/NET0131  , \u26_cnt_reg[0]/NET0131  , \u26_cnt_reg[1]/NET0131  , \u26_cnt_reg[2]/NET0131  , \u26_ps_cnt_reg[0]/NET0131  , \u26_ps_cnt_reg[1]/NET0131  , \u26_ps_cnt_reg[2]/NET0131  , \u26_ps_cnt_reg[3]/NET0131  , \u26_ps_cnt_reg[4]/NET0131  , \u26_ps_cnt_reg[5]/NET0131  , \u2_bit_clk_e_reg/P0001  , \u2_bit_clk_r1_reg/P0001  , \u2_bit_clk_r_reg/P0001  , \u2_cnt_reg[0]/NET0131  , \u2_cnt_reg[1]/NET0131  , \u2_cnt_reg[2]/NET0131  , \u2_cnt_reg[3]/NET0131  , \u2_cnt_reg[4]/NET0131  , \u2_cnt_reg[5]/NET0131  , \u2_cnt_reg[6]/NET0131  , \u2_cnt_reg[7]/NET0131  , \u2_ld_reg/P0001  , \u2_out_le_reg[0]/P0001  , \u2_out_le_reg[1]/P0001  , \u2_res_cnt_reg[0]/P0001  , \u2_res_cnt_reg[1]/P0001  , \u2_res_cnt_reg[2]/P0001  , \u2_res_cnt_reg[3]/P0001  , \u2_sync_beat_reg/P0001  , \u2_sync_resume_reg/NET0131  , \u2_to_cnt_reg[0]/NET0131  , \u2_to_cnt_reg[1]/NET0131  , \u2_to_cnt_reg[2]/NET0131  , \u2_to_cnt_reg[3]/NET0131  , \u2_to_cnt_reg[4]/NET0131  , \u2_to_cnt_reg[5]/NET0131  , \u3_dout_reg[0]/P0001  , \u3_dout_reg[10]/P0001  , \u3_dout_reg[11]/P0001  , \u3_dout_reg[12]/P0001  , \u3_dout_reg[13]/P0001  , \u3_dout_reg[14]/P0001  , \u3_dout_reg[15]/P0001  , \u3_dout_reg[16]/P0001  , \u3_dout_reg[17]/P0001  , \u3_dout_reg[18]/P0001  , \u3_dout_reg[19]/P0001  , \u3_dout_reg[1]/P0001  , \u3_dout_reg[2]/P0001  , \u3_dout_reg[3]/P0001  , \u3_dout_reg[4]/P0001  , \u3_dout_reg[5]/P0001  , \u3_dout_reg[6]/P0001  , \u3_dout_reg[7]/P0001  , \u3_dout_reg[8]/P0001  , \u3_dout_reg[9]/P0001  , \u3_empty_reg/NET0131  , \u3_mem_reg[0][0]/NET0131  , \u3_mem_reg[0][10]/NET0131  , \u3_mem_reg[0][11]/NET0131  , \u3_mem_reg[0][12]/NET0131  , \u3_mem_reg[0][13]/NET0131  , \u3_mem_reg[0][14]/NET0131  , \u3_mem_reg[0][15]/NET0131  , \u3_mem_reg[0][16]/NET0131  , \u3_mem_reg[0][17]/NET0131  , \u3_mem_reg[0][18]/NET0131  , \u3_mem_reg[0][19]/NET0131  , \u3_mem_reg[0][1]/NET0131  , \u3_mem_reg[0][20]/NET0131  , \u3_mem_reg[0][21]/NET0131  , \u3_mem_reg[0][22]/NET0131  , \u3_mem_reg[0][23]/NET0131  , \u3_mem_reg[0][24]/NET0131  , \u3_mem_reg[0][25]/NET0131  , \u3_mem_reg[0][26]/NET0131  , \u3_mem_reg[0][27]/NET0131  , \u3_mem_reg[0][28]/NET0131  , \u3_mem_reg[0][29]/NET0131  , \u3_mem_reg[0][2]/NET0131  , \u3_mem_reg[0][30]/NET0131  , \u3_mem_reg[0][31]/NET0131  , \u3_mem_reg[0][3]/NET0131  , \u3_mem_reg[0][4]/NET0131  , \u3_mem_reg[0][5]/NET0131  , \u3_mem_reg[0][6]/NET0131  , \u3_mem_reg[0][7]/NET0131  , \u3_mem_reg[0][8]/NET0131  , \u3_mem_reg[0][9]/NET0131  , \u3_mem_reg[1][0]/NET0131  , \u3_mem_reg[1][10]/NET0131  , \u3_mem_reg[1][11]/NET0131  , \u3_mem_reg[1][12]/NET0131  , \u3_mem_reg[1][13]/NET0131  , \u3_mem_reg[1][14]/NET0131  , \u3_mem_reg[1][15]/NET0131  , \u3_mem_reg[1][16]/NET0131  , \u3_mem_reg[1][17]/NET0131  , \u3_mem_reg[1][18]/NET0131  , \u3_mem_reg[1][19]/NET0131  , \u3_mem_reg[1][1]/NET0131  , \u3_mem_reg[1][20]/NET0131  , \u3_mem_reg[1][21]/NET0131  , \u3_mem_reg[1][22]/NET0131  , \u3_mem_reg[1][23]/NET0131  , \u3_mem_reg[1][24]/NET0131  , \u3_mem_reg[1][25]/NET0131  , \u3_mem_reg[1][26]/NET0131  , \u3_mem_reg[1][27]/NET0131  , \u3_mem_reg[1][28]/NET0131  , \u3_mem_reg[1][29]/NET0131  , \u3_mem_reg[1][2]/NET0131  , \u3_mem_reg[1][30]/NET0131  , \u3_mem_reg[1][31]/NET0131  , \u3_mem_reg[1][3]/NET0131  , \u3_mem_reg[1][4]/NET0131  , \u3_mem_reg[1][5]/NET0131  , \u3_mem_reg[1][6]/NET0131  , \u3_mem_reg[1][7]/NET0131  , \u3_mem_reg[1][8]/NET0131  , \u3_mem_reg[1][9]/NET0131  , \u3_mem_reg[2][0]/NET0131  , \u3_mem_reg[2][10]/NET0131  , \u3_mem_reg[2][11]/NET0131  , \u3_mem_reg[2][12]/NET0131  , \u3_mem_reg[2][13]/NET0131  , \u3_mem_reg[2][14]/NET0131  , \u3_mem_reg[2][15]/NET0131  , \u3_mem_reg[2][16]/NET0131  , \u3_mem_reg[2][17]/NET0131  , \u3_mem_reg[2][18]/NET0131  , \u3_mem_reg[2][19]/NET0131  , \u3_mem_reg[2][1]/NET0131  , \u3_mem_reg[2][20]/NET0131  , \u3_mem_reg[2][21]/NET0131  , \u3_mem_reg[2][22]/NET0131  , \u3_mem_reg[2][23]/NET0131  , \u3_mem_reg[2][24]/NET0131  , \u3_mem_reg[2][25]/NET0131  , \u3_mem_reg[2][26]/NET0131  , \u3_mem_reg[2][27]/NET0131  , \u3_mem_reg[2][28]/NET0131  , \u3_mem_reg[2][29]/NET0131  , \u3_mem_reg[2][2]/NET0131  , \u3_mem_reg[2][30]/NET0131  , \u3_mem_reg[2][31]/NET0131  , \u3_mem_reg[2][3]/NET0131  , \u3_mem_reg[2][4]/NET0131  , \u3_mem_reg[2][5]/NET0131  , \u3_mem_reg[2][6]/NET0131  , \u3_mem_reg[2][7]/NET0131  , \u3_mem_reg[2][8]/NET0131  , \u3_mem_reg[2][9]/NET0131  , \u3_mem_reg[3][0]/NET0131  , \u3_mem_reg[3][10]/NET0131  , \u3_mem_reg[3][11]/NET0131  , \u3_mem_reg[3][12]/NET0131  , \u3_mem_reg[3][13]/NET0131  , \u3_mem_reg[3][14]/NET0131  , \u3_mem_reg[3][15]/NET0131  , \u3_mem_reg[3][16]/NET0131  , \u3_mem_reg[3][17]/NET0131  , \u3_mem_reg[3][18]/NET0131  , \u3_mem_reg[3][19]/NET0131  , \u3_mem_reg[3][1]/NET0131  , \u3_mem_reg[3][20]/NET0131  , \u3_mem_reg[3][21]/NET0131  , \u3_mem_reg[3][22]/NET0131  , \u3_mem_reg[3][23]/NET0131  , \u3_mem_reg[3][24]/NET0131  , \u3_mem_reg[3][25]/NET0131  , \u3_mem_reg[3][26]/NET0131  , \u3_mem_reg[3][27]/NET0131  , \u3_mem_reg[3][28]/NET0131  , \u3_mem_reg[3][29]/NET0131  , \u3_mem_reg[3][2]/NET0131  , \u3_mem_reg[3][30]/NET0131  , \u3_mem_reg[3][31]/NET0131  , \u3_mem_reg[3][3]/NET0131  , \u3_mem_reg[3][4]/NET0131  , \u3_mem_reg[3][5]/NET0131  , \u3_mem_reg[3][6]/NET0131  , \u3_mem_reg[3][7]/NET0131  , \u3_mem_reg[3][8]/NET0131  , \u3_mem_reg[3][9]/NET0131  , \u3_rp_reg[0]/P0001  , \u3_rp_reg[1]/NET0131  , \u3_rp_reg[2]/NET0131  , \u3_rp_reg[3]/NET0131  , \u3_status_reg[0]/P0001  , \u3_status_reg[1]/P0001  , \u3_wp_reg[0]/P0001  , \u3_wp_reg[1]/NET0131  , \u3_wp_reg[2]/P0001  , \u4_dout_reg[0]/P0001  , \u4_dout_reg[10]/P0001  , \u4_dout_reg[11]/P0001  , \u4_dout_reg[12]/P0001  , \u4_dout_reg[13]/P0001  , \u4_dout_reg[14]/P0001  , \u4_dout_reg[15]/P0001  , \u4_dout_reg[16]/P0001  , \u4_dout_reg[17]/P0001  , \u4_dout_reg[18]/P0001  , \u4_dout_reg[19]/P0001  , \u4_dout_reg[1]/P0001  , \u4_dout_reg[2]/P0001  , \u4_dout_reg[3]/P0001  , \u4_dout_reg[4]/P0001  , \u4_dout_reg[5]/P0001  , \u4_dout_reg[6]/P0001  , \u4_dout_reg[7]/P0001  , \u4_dout_reg[8]/P0001  , \u4_dout_reg[9]/P0001  , \u4_empty_reg/NET0131  , \u4_mem_reg[0][0]/NET0131  , \u4_mem_reg[0][10]/NET0131  , \u4_mem_reg[0][11]/NET0131  , \u4_mem_reg[0][12]/NET0131  , \u4_mem_reg[0][13]/NET0131  , \u4_mem_reg[0][14]/NET0131  , \u4_mem_reg[0][15]/NET0131  , \u4_mem_reg[0][16]/NET0131  , \u4_mem_reg[0][17]/NET0131  , \u4_mem_reg[0][18]/NET0131  , \u4_mem_reg[0][19]/NET0131  , \u4_mem_reg[0][1]/NET0131  , \u4_mem_reg[0][20]/NET0131  , \u4_mem_reg[0][21]/NET0131  , \u4_mem_reg[0][22]/NET0131  , \u4_mem_reg[0][23]/NET0131  , \u4_mem_reg[0][24]/NET0131  , \u4_mem_reg[0][25]/NET0131  , \u4_mem_reg[0][26]/NET0131  , \u4_mem_reg[0][27]/NET0131  , \u4_mem_reg[0][28]/NET0131  , \u4_mem_reg[0][29]/NET0131  , \u4_mem_reg[0][2]/NET0131  , \u4_mem_reg[0][30]/NET0131  , \u4_mem_reg[0][31]/NET0131  , \u4_mem_reg[0][3]/NET0131  , \u4_mem_reg[0][4]/NET0131  , \u4_mem_reg[0][5]/NET0131  , \u4_mem_reg[0][6]/NET0131  , \u4_mem_reg[0][7]/NET0131  , \u4_mem_reg[0][8]/NET0131  , \u4_mem_reg[0][9]/NET0131  , \u4_mem_reg[1][0]/NET0131  , \u4_mem_reg[1][10]/NET0131  , \u4_mem_reg[1][11]/NET0131  , \u4_mem_reg[1][12]/NET0131  , \u4_mem_reg[1][13]/NET0131  , \u4_mem_reg[1][14]/NET0131  , \u4_mem_reg[1][15]/NET0131  , \u4_mem_reg[1][16]/NET0131  , \u4_mem_reg[1][17]/NET0131  , \u4_mem_reg[1][18]/NET0131  , \u4_mem_reg[1][19]/NET0131  , \u4_mem_reg[1][1]/NET0131  , \u4_mem_reg[1][20]/NET0131  , \u4_mem_reg[1][21]/NET0131  , \u4_mem_reg[1][22]/NET0131  , \u4_mem_reg[1][23]/NET0131  , \u4_mem_reg[1][24]/NET0131  , \u4_mem_reg[1][25]/NET0131  , \u4_mem_reg[1][26]/NET0131  , \u4_mem_reg[1][27]/NET0131  , \u4_mem_reg[1][28]/NET0131  , \u4_mem_reg[1][29]/NET0131  , \u4_mem_reg[1][2]/NET0131  , \u4_mem_reg[1][30]/NET0131  , \u4_mem_reg[1][31]/NET0131  , \u4_mem_reg[1][3]/NET0131  , \u4_mem_reg[1][4]/NET0131  , \u4_mem_reg[1][5]/NET0131  , \u4_mem_reg[1][6]/NET0131  , \u4_mem_reg[1][7]/NET0131  , \u4_mem_reg[1][8]/NET0131  , \u4_mem_reg[1][9]/NET0131  , \u4_mem_reg[2][0]/NET0131  , \u4_mem_reg[2][10]/NET0131  , \u4_mem_reg[2][11]/NET0131  , \u4_mem_reg[2][12]/NET0131  , \u4_mem_reg[2][13]/NET0131  , \u4_mem_reg[2][14]/NET0131  , \u4_mem_reg[2][15]/NET0131  , \u4_mem_reg[2][16]/NET0131  , \u4_mem_reg[2][17]/NET0131  , \u4_mem_reg[2][18]/NET0131  , \u4_mem_reg[2][19]/NET0131  , \u4_mem_reg[2][1]/NET0131  , \u4_mem_reg[2][20]/NET0131  , \u4_mem_reg[2][21]/NET0131  , \u4_mem_reg[2][22]/NET0131  , \u4_mem_reg[2][23]/NET0131  , \u4_mem_reg[2][24]/NET0131  , \u4_mem_reg[2][25]/NET0131  , \u4_mem_reg[2][26]/NET0131  , \u4_mem_reg[2][27]/NET0131  , \u4_mem_reg[2][28]/NET0131  , \u4_mem_reg[2][29]/NET0131  , \u4_mem_reg[2][2]/NET0131  , \u4_mem_reg[2][30]/NET0131  , \u4_mem_reg[2][31]/NET0131  , \u4_mem_reg[2][3]/NET0131  , \u4_mem_reg[2][4]/NET0131  , \u4_mem_reg[2][5]/NET0131  , \u4_mem_reg[2][6]/NET0131  , \u4_mem_reg[2][7]/NET0131  , \u4_mem_reg[2][8]/NET0131  , \u4_mem_reg[2][9]/NET0131  , \u4_mem_reg[3][0]/NET0131  , \u4_mem_reg[3][10]/NET0131  , \u4_mem_reg[3][11]/NET0131  , \u4_mem_reg[3][12]/NET0131  , \u4_mem_reg[3][13]/NET0131  , \u4_mem_reg[3][14]/NET0131  , \u4_mem_reg[3][15]/NET0131  , \u4_mem_reg[3][16]/NET0131  , \u4_mem_reg[3][17]/NET0131  , \u4_mem_reg[3][18]/NET0131  , \u4_mem_reg[3][19]/NET0131  , \u4_mem_reg[3][1]/NET0131  , \u4_mem_reg[3][20]/NET0131  , \u4_mem_reg[3][21]/NET0131  , \u4_mem_reg[3][22]/NET0131  , \u4_mem_reg[3][23]/NET0131  , \u4_mem_reg[3][24]/NET0131  , \u4_mem_reg[3][25]/NET0131  , \u4_mem_reg[3][26]/NET0131  , \u4_mem_reg[3][27]/NET0131  , \u4_mem_reg[3][28]/NET0131  , \u4_mem_reg[3][29]/NET0131  , \u4_mem_reg[3][2]/NET0131  , \u4_mem_reg[3][30]/NET0131  , \u4_mem_reg[3][31]/NET0131  , \u4_mem_reg[3][3]/NET0131  , \u4_mem_reg[3][4]/NET0131  , \u4_mem_reg[3][5]/NET0131  , \u4_mem_reg[3][6]/NET0131  , \u4_mem_reg[3][7]/NET0131  , \u4_mem_reg[3][8]/NET0131  , \u4_mem_reg[3][9]/NET0131  , \u4_rp_reg[0]/P0001  , \u4_rp_reg[1]/NET0131  , \u4_rp_reg[2]/NET0131  , \u4_rp_reg[3]/NET0131  , \u4_status_reg[0]/P0001  , \u4_status_reg[1]/P0001  , \u4_wp_reg[0]/P0001  , \u4_wp_reg[1]/NET0131  , \u4_wp_reg[2]/P0001  , \u5_dout_reg[0]/P0001  , \u5_dout_reg[10]/P0001  , \u5_dout_reg[11]/P0001  , \u5_dout_reg[12]/P0001  , \u5_dout_reg[13]/P0001  , \u5_dout_reg[14]/P0001  , \u5_dout_reg[15]/P0001  , \u5_dout_reg[16]/P0001  , \u5_dout_reg[17]/P0001  , \u5_dout_reg[18]/P0001  , \u5_dout_reg[19]/P0001  , \u5_dout_reg[1]/P0001  , \u5_dout_reg[2]/P0001  , \u5_dout_reg[3]/P0001  , \u5_dout_reg[4]/P0001  , \u5_dout_reg[5]/P0001  , \u5_dout_reg[6]/P0001  , \u5_dout_reg[7]/P0001  , \u5_dout_reg[8]/P0001  , \u5_dout_reg[9]/P0001  , \u5_empty_reg/NET0131  , \u5_mem_reg[0][0]/NET0131  , \u5_mem_reg[0][10]/NET0131  , \u5_mem_reg[0][11]/NET0131  , \u5_mem_reg[0][12]/NET0131  , \u5_mem_reg[0][13]/NET0131  , \u5_mem_reg[0][14]/NET0131  , \u5_mem_reg[0][15]/NET0131  , \u5_mem_reg[0][16]/NET0131  , \u5_mem_reg[0][17]/NET0131  , \u5_mem_reg[0][18]/NET0131  , \u5_mem_reg[0][19]/NET0131  , \u5_mem_reg[0][1]/NET0131  , \u5_mem_reg[0][20]/NET0131  , \u5_mem_reg[0][21]/NET0131  , \u5_mem_reg[0][22]/NET0131  , \u5_mem_reg[0][23]/NET0131  , \u5_mem_reg[0][24]/NET0131  , \u5_mem_reg[0][25]/NET0131  , \u5_mem_reg[0][26]/NET0131  , \u5_mem_reg[0][27]/NET0131  , \u5_mem_reg[0][28]/NET0131  , \u5_mem_reg[0][29]/NET0131  , \u5_mem_reg[0][2]/NET0131  , \u5_mem_reg[0][30]/NET0131  , \u5_mem_reg[0][31]/NET0131  , \u5_mem_reg[0][3]/NET0131  , \u5_mem_reg[0][4]/NET0131  , \u5_mem_reg[0][5]/NET0131  , \u5_mem_reg[0][6]/NET0131  , \u5_mem_reg[0][7]/NET0131  , \u5_mem_reg[0][8]/NET0131  , \u5_mem_reg[0][9]/NET0131  , \u5_mem_reg[1][0]/NET0131  , \u5_mem_reg[1][10]/NET0131  , \u5_mem_reg[1][11]/NET0131  , \u5_mem_reg[1][12]/NET0131  , \u5_mem_reg[1][13]/NET0131  , \u5_mem_reg[1][14]/NET0131  , \u5_mem_reg[1][15]/NET0131  , \u5_mem_reg[1][16]/NET0131  , \u5_mem_reg[1][17]/NET0131  , \u5_mem_reg[1][18]/NET0131  , \u5_mem_reg[1][19]/NET0131  , \u5_mem_reg[1][1]/NET0131  , \u5_mem_reg[1][20]/NET0131  , \u5_mem_reg[1][21]/NET0131  , \u5_mem_reg[1][22]/NET0131  , \u5_mem_reg[1][23]/NET0131  , \u5_mem_reg[1][24]/NET0131  , \u5_mem_reg[1][25]/NET0131  , \u5_mem_reg[1][26]/NET0131  , \u5_mem_reg[1][27]/NET0131  , \u5_mem_reg[1][28]/NET0131  , \u5_mem_reg[1][29]/NET0131  , \u5_mem_reg[1][2]/NET0131  , \u5_mem_reg[1][30]/NET0131  , \u5_mem_reg[1][31]/NET0131  , \u5_mem_reg[1][3]/NET0131  , \u5_mem_reg[1][4]/NET0131  , \u5_mem_reg[1][5]/NET0131  , \u5_mem_reg[1][6]/NET0131  , \u5_mem_reg[1][7]/NET0131  , \u5_mem_reg[1][8]/NET0131  , \u5_mem_reg[1][9]/NET0131  , \u5_mem_reg[2][0]/NET0131  , \u5_mem_reg[2][10]/NET0131  , \u5_mem_reg[2][11]/NET0131  , \u5_mem_reg[2][12]/NET0131  , \u5_mem_reg[2][13]/NET0131  , \u5_mem_reg[2][14]/NET0131  , \u5_mem_reg[2][15]/NET0131  , \u5_mem_reg[2][16]/NET0131  , \u5_mem_reg[2][17]/NET0131  , \u5_mem_reg[2][18]/NET0131  , \u5_mem_reg[2][19]/NET0131  , \u5_mem_reg[2][1]/NET0131  , \u5_mem_reg[2][20]/NET0131  , \u5_mem_reg[2][21]/NET0131  , \u5_mem_reg[2][22]/NET0131  , \u5_mem_reg[2][23]/NET0131  , \u5_mem_reg[2][24]/NET0131  , \u5_mem_reg[2][25]/NET0131  , \u5_mem_reg[2][26]/NET0131  , \u5_mem_reg[2][27]/NET0131  , \u5_mem_reg[2][28]/NET0131  , \u5_mem_reg[2][29]/NET0131  , \u5_mem_reg[2][2]/NET0131  , \u5_mem_reg[2][30]/NET0131  , \u5_mem_reg[2][31]/NET0131  , \u5_mem_reg[2][3]/NET0131  , \u5_mem_reg[2][4]/NET0131  , \u5_mem_reg[2][5]/NET0131  , \u5_mem_reg[2][6]/NET0131  , \u5_mem_reg[2][7]/NET0131  , \u5_mem_reg[2][8]/NET0131  , \u5_mem_reg[2][9]/NET0131  , \u5_mem_reg[3][0]/NET0131  , \u5_mem_reg[3][10]/NET0131  , \u5_mem_reg[3][11]/NET0131  , \u5_mem_reg[3][12]/NET0131  , \u5_mem_reg[3][13]/NET0131  , \u5_mem_reg[3][14]/NET0131  , \u5_mem_reg[3][15]/NET0131  , \u5_mem_reg[3][16]/NET0131  , \u5_mem_reg[3][17]/NET0131  , \u5_mem_reg[3][18]/NET0131  , \u5_mem_reg[3][19]/NET0131  , \u5_mem_reg[3][1]/NET0131  , \u5_mem_reg[3][20]/NET0131  , \u5_mem_reg[3][21]/NET0131  , \u5_mem_reg[3][22]/NET0131  , \u5_mem_reg[3][23]/NET0131  , \u5_mem_reg[3][24]/NET0131  , \u5_mem_reg[3][25]/NET0131  , \u5_mem_reg[3][26]/NET0131  , \u5_mem_reg[3][27]/NET0131  , \u5_mem_reg[3][28]/NET0131  , \u5_mem_reg[3][29]/NET0131  , \u5_mem_reg[3][2]/NET0131  , \u5_mem_reg[3][30]/NET0131  , \u5_mem_reg[3][31]/NET0131  , \u5_mem_reg[3][3]/NET0131  , \u5_mem_reg[3][4]/NET0131  , \u5_mem_reg[3][5]/NET0131  , \u5_mem_reg[3][6]/NET0131  , \u5_mem_reg[3][7]/NET0131  , \u5_mem_reg[3][8]/NET0131  , \u5_mem_reg[3][9]/NET0131  , \u5_rp_reg[0]/P0001  , \u5_rp_reg[1]/NET0131  , \u5_rp_reg[2]/NET0131  , \u5_rp_reg[3]/NET0131  , \u5_status_reg[0]/P0001  , \u5_status_reg[1]/P0001  , \u5_wp_reg[0]/P0001  , \u5_wp_reg[1]/NET0131  , \u5_wp_reg[2]/P0001  , \u6_dout_reg[0]/P0001  , \u6_dout_reg[10]/P0001  , \u6_dout_reg[11]/P0001  , \u6_dout_reg[12]/P0001  , \u6_dout_reg[13]/P0001  , \u6_dout_reg[14]/P0001  , \u6_dout_reg[15]/P0001  , \u6_dout_reg[16]/P0001  , \u6_dout_reg[17]/P0001  , \u6_dout_reg[18]/P0001  , \u6_dout_reg[19]/P0001  , \u6_dout_reg[1]/P0001  , \u6_dout_reg[2]/P0001  , \u6_dout_reg[3]/P0001  , \u6_dout_reg[4]/P0001  , \u6_dout_reg[5]/P0001  , \u6_dout_reg[6]/P0001  , \u6_dout_reg[7]/P0001  , \u6_dout_reg[8]/P0001  , \u6_dout_reg[9]/P0001  , \u6_empty_reg/NET0131  , \u6_mem_reg[0][0]/NET0131  , \u6_mem_reg[0][10]/NET0131  , \u6_mem_reg[0][11]/NET0131  , \u6_mem_reg[0][12]/NET0131  , \u6_mem_reg[0][13]/NET0131  , \u6_mem_reg[0][14]/NET0131  , \u6_mem_reg[0][15]/NET0131  , \u6_mem_reg[0][16]/NET0131  , \u6_mem_reg[0][17]/NET0131  , \u6_mem_reg[0][18]/NET0131  , \u6_mem_reg[0][19]/NET0131  , \u6_mem_reg[0][1]/NET0131  , \u6_mem_reg[0][20]/NET0131  , \u6_mem_reg[0][21]/NET0131  , \u6_mem_reg[0][22]/NET0131  , \u6_mem_reg[0][23]/NET0131  , \u6_mem_reg[0][24]/NET0131  , \u6_mem_reg[0][25]/NET0131  , \u6_mem_reg[0][26]/NET0131  , \u6_mem_reg[0][27]/NET0131  , \u6_mem_reg[0][28]/NET0131  , \u6_mem_reg[0][29]/NET0131  , \u6_mem_reg[0][2]/NET0131  , \u6_mem_reg[0][30]/NET0131  , \u6_mem_reg[0][31]/NET0131  , \u6_mem_reg[0][3]/NET0131  , \u6_mem_reg[0][4]/NET0131  , \u6_mem_reg[0][5]/NET0131  , \u6_mem_reg[0][6]/NET0131  , \u6_mem_reg[0][7]/NET0131  , \u6_mem_reg[0][8]/NET0131  , \u6_mem_reg[0][9]/NET0131  , \u6_mem_reg[1][0]/NET0131  , \u6_mem_reg[1][10]/NET0131  , \u6_mem_reg[1][11]/NET0131  , \u6_mem_reg[1][12]/NET0131  , \u6_mem_reg[1][13]/NET0131  , \u6_mem_reg[1][14]/NET0131  , \u6_mem_reg[1][15]/NET0131  , \u6_mem_reg[1][16]/NET0131  , \u6_mem_reg[1][17]/NET0131  , \u6_mem_reg[1][18]/NET0131  , \u6_mem_reg[1][19]/NET0131  , \u6_mem_reg[1][1]/NET0131  , \u6_mem_reg[1][20]/NET0131  , \u6_mem_reg[1][21]/NET0131  , \u6_mem_reg[1][22]/NET0131  , \u6_mem_reg[1][23]/NET0131  , \u6_mem_reg[1][24]/NET0131  , \u6_mem_reg[1][25]/NET0131  , \u6_mem_reg[1][26]/NET0131  , \u6_mem_reg[1][27]/NET0131  , \u6_mem_reg[1][28]/NET0131  , \u6_mem_reg[1][29]/NET0131  , \u6_mem_reg[1][2]/NET0131  , \u6_mem_reg[1][30]/NET0131  , \u6_mem_reg[1][31]/NET0131  , \u6_mem_reg[1][3]/NET0131  , \u6_mem_reg[1][4]/NET0131  , \u6_mem_reg[1][5]/NET0131  , \u6_mem_reg[1][6]/NET0131  , \u6_mem_reg[1][7]/NET0131  , \u6_mem_reg[1][8]/NET0131  , \u6_mem_reg[1][9]/NET0131  , \u6_mem_reg[2][0]/NET0131  , \u6_mem_reg[2][10]/NET0131  , \u6_mem_reg[2][11]/NET0131  , \u6_mem_reg[2][12]/NET0131  , \u6_mem_reg[2][13]/NET0131  , \u6_mem_reg[2][14]/NET0131  , \u6_mem_reg[2][15]/NET0131  , \u6_mem_reg[2][16]/NET0131  , \u6_mem_reg[2][17]/NET0131  , \u6_mem_reg[2][18]/NET0131  , \u6_mem_reg[2][19]/NET0131  , \u6_mem_reg[2][1]/NET0131  , \u6_mem_reg[2][20]/NET0131  , \u6_mem_reg[2][21]/NET0131  , \u6_mem_reg[2][22]/NET0131  , \u6_mem_reg[2][23]/NET0131  , \u6_mem_reg[2][24]/NET0131  , \u6_mem_reg[2][25]/NET0131  , \u6_mem_reg[2][26]/NET0131  , \u6_mem_reg[2][27]/NET0131  , \u6_mem_reg[2][28]/NET0131  , \u6_mem_reg[2][29]/NET0131  , \u6_mem_reg[2][2]/NET0131  , \u6_mem_reg[2][30]/NET0131  , \u6_mem_reg[2][31]/NET0131  , \u6_mem_reg[2][3]/NET0131  , \u6_mem_reg[2][4]/NET0131  , \u6_mem_reg[2][5]/NET0131  , \u6_mem_reg[2][6]/NET0131  , \u6_mem_reg[2][7]/NET0131  , \u6_mem_reg[2][8]/NET0131  , \u6_mem_reg[2][9]/NET0131  , \u6_mem_reg[3][0]/NET0131  , \u6_mem_reg[3][10]/NET0131  , \u6_mem_reg[3][11]/NET0131  , \u6_mem_reg[3][12]/NET0131  , \u6_mem_reg[3][13]/NET0131  , \u6_mem_reg[3][14]/NET0131  , \u6_mem_reg[3][15]/NET0131  , \u6_mem_reg[3][16]/NET0131  , \u6_mem_reg[3][17]/NET0131  , \u6_mem_reg[3][18]/NET0131  , \u6_mem_reg[3][19]/NET0131  , \u6_mem_reg[3][1]/NET0131  , \u6_mem_reg[3][20]/NET0131  , \u6_mem_reg[3][21]/NET0131  , \u6_mem_reg[3][22]/NET0131  , \u6_mem_reg[3][23]/NET0131  , \u6_mem_reg[3][24]/NET0131  , \u6_mem_reg[3][25]/NET0131  , \u6_mem_reg[3][26]/NET0131  , \u6_mem_reg[3][27]/NET0131  , \u6_mem_reg[3][28]/NET0131  , \u6_mem_reg[3][29]/NET0131  , \u6_mem_reg[3][2]/NET0131  , \u6_mem_reg[3][30]/NET0131  , \u6_mem_reg[3][31]/NET0131  , \u6_mem_reg[3][3]/NET0131  , \u6_mem_reg[3][4]/NET0131  , \u6_mem_reg[3][5]/NET0131  , \u6_mem_reg[3][6]/NET0131  , \u6_mem_reg[3][7]/NET0131  , \u6_mem_reg[3][8]/NET0131  , \u6_mem_reg[3][9]/NET0131  , \u6_rp_reg[0]/P0001  , \u6_rp_reg[1]/NET0131  , \u6_rp_reg[2]/NET0131  , \u6_rp_reg[3]/NET0131  , \u6_status_reg[0]/P0001  , \u6_status_reg[1]/P0001  , \u6_wp_reg[0]/P0001  , \u6_wp_reg[1]/NET0131  , \u6_wp_reg[2]/P0001  , \u7_dout_reg[0]/P0001  , \u7_dout_reg[10]/P0001  , \u7_dout_reg[11]/P0001  , \u7_dout_reg[12]/P0001  , \u7_dout_reg[13]/P0001  , \u7_dout_reg[14]/P0001  , \u7_dout_reg[15]/P0001  , \u7_dout_reg[16]/P0001  , \u7_dout_reg[17]/P0001  , \u7_dout_reg[18]/P0001  , \u7_dout_reg[19]/P0001  , \u7_dout_reg[1]/P0001  , \u7_dout_reg[2]/P0001  , \u7_dout_reg[3]/P0001  , \u7_dout_reg[4]/P0001  , \u7_dout_reg[5]/P0001  , \u7_dout_reg[6]/P0001  , \u7_dout_reg[7]/P0001  , \u7_dout_reg[8]/P0001  , \u7_dout_reg[9]/P0001  , \u7_empty_reg/NET0131  , \u7_mem_reg[0][0]/NET0131  , \u7_mem_reg[0][10]/NET0131  , \u7_mem_reg[0][11]/NET0131  , \u7_mem_reg[0][12]/NET0131  , \u7_mem_reg[0][13]/NET0131  , \u7_mem_reg[0][14]/NET0131  , \u7_mem_reg[0][15]/NET0131  , \u7_mem_reg[0][16]/NET0131  , \u7_mem_reg[0][17]/NET0131  , \u7_mem_reg[0][18]/NET0131  , \u7_mem_reg[0][19]/NET0131  , \u7_mem_reg[0][1]/NET0131  , \u7_mem_reg[0][20]/NET0131  , \u7_mem_reg[0][21]/NET0131  , \u7_mem_reg[0][22]/NET0131  , \u7_mem_reg[0][23]/NET0131  , \u7_mem_reg[0][24]/NET0131  , \u7_mem_reg[0][25]/NET0131  , \u7_mem_reg[0][26]/NET0131  , \u7_mem_reg[0][27]/NET0131  , \u7_mem_reg[0][28]/NET0131  , \u7_mem_reg[0][29]/NET0131  , \u7_mem_reg[0][2]/NET0131  , \u7_mem_reg[0][30]/NET0131  , \u7_mem_reg[0][31]/NET0131  , \u7_mem_reg[0][3]/NET0131  , \u7_mem_reg[0][4]/NET0131  , \u7_mem_reg[0][5]/NET0131  , \u7_mem_reg[0][6]/NET0131  , \u7_mem_reg[0][7]/NET0131  , \u7_mem_reg[0][8]/NET0131  , \u7_mem_reg[0][9]/NET0131  , \u7_mem_reg[1][0]/NET0131  , \u7_mem_reg[1][10]/NET0131  , \u7_mem_reg[1][11]/NET0131  , \u7_mem_reg[1][12]/NET0131  , \u7_mem_reg[1][13]/NET0131  , \u7_mem_reg[1][14]/NET0131  , \u7_mem_reg[1][15]/NET0131  , \u7_mem_reg[1][16]/NET0131  , \u7_mem_reg[1][17]/NET0131  , \u7_mem_reg[1][18]/NET0131  , \u7_mem_reg[1][19]/NET0131  , \u7_mem_reg[1][1]/NET0131  , \u7_mem_reg[1][20]/NET0131  , \u7_mem_reg[1][21]/NET0131  , \u7_mem_reg[1][22]/NET0131  , \u7_mem_reg[1][23]/NET0131  , \u7_mem_reg[1][24]/NET0131  , \u7_mem_reg[1][25]/NET0131  , \u7_mem_reg[1][26]/NET0131  , \u7_mem_reg[1][27]/NET0131  , \u7_mem_reg[1][28]/NET0131  , \u7_mem_reg[1][29]/NET0131  , \u7_mem_reg[1][2]/NET0131  , \u7_mem_reg[1][30]/NET0131  , \u7_mem_reg[1][31]/NET0131  , \u7_mem_reg[1][3]/NET0131  , \u7_mem_reg[1][4]/NET0131  , \u7_mem_reg[1][5]/NET0131  , \u7_mem_reg[1][6]/NET0131  , \u7_mem_reg[1][7]/NET0131  , \u7_mem_reg[1][8]/NET0131  , \u7_mem_reg[1][9]/NET0131  , \u7_mem_reg[2][0]/NET0131  , \u7_mem_reg[2][10]/NET0131  , \u7_mem_reg[2][11]/NET0131  , \u7_mem_reg[2][12]/NET0131  , \u7_mem_reg[2][13]/NET0131  , \u7_mem_reg[2][14]/NET0131  , \u7_mem_reg[2][15]/NET0131  , \u7_mem_reg[2][16]/NET0131  , \u7_mem_reg[2][17]/NET0131  , \u7_mem_reg[2][18]/NET0131  , \u7_mem_reg[2][19]/NET0131  , \u7_mem_reg[2][1]/NET0131  , \u7_mem_reg[2][20]/NET0131  , \u7_mem_reg[2][21]/NET0131  , \u7_mem_reg[2][22]/NET0131  , \u7_mem_reg[2][23]/NET0131  , \u7_mem_reg[2][24]/NET0131  , \u7_mem_reg[2][25]/NET0131  , \u7_mem_reg[2][26]/NET0131  , \u7_mem_reg[2][27]/NET0131  , \u7_mem_reg[2][28]/NET0131  , \u7_mem_reg[2][29]/NET0131  , \u7_mem_reg[2][2]/NET0131  , \u7_mem_reg[2][30]/NET0131  , \u7_mem_reg[2][31]/NET0131  , \u7_mem_reg[2][3]/NET0131  , \u7_mem_reg[2][4]/NET0131  , \u7_mem_reg[2][5]/NET0131  , \u7_mem_reg[2][6]/NET0131  , \u7_mem_reg[2][7]/NET0131  , \u7_mem_reg[2][8]/NET0131  , \u7_mem_reg[2][9]/NET0131  , \u7_mem_reg[3][0]/NET0131  , \u7_mem_reg[3][10]/NET0131  , \u7_mem_reg[3][11]/NET0131  , \u7_mem_reg[3][12]/NET0131  , \u7_mem_reg[3][13]/NET0131  , \u7_mem_reg[3][14]/NET0131  , \u7_mem_reg[3][15]/NET0131  , \u7_mem_reg[3][16]/NET0131  , \u7_mem_reg[3][17]/NET0131  , \u7_mem_reg[3][18]/NET0131  , \u7_mem_reg[3][19]/NET0131  , \u7_mem_reg[3][1]/NET0131  , \u7_mem_reg[3][20]/NET0131  , \u7_mem_reg[3][21]/NET0131  , \u7_mem_reg[3][22]/NET0131  , \u7_mem_reg[3][23]/NET0131  , \u7_mem_reg[3][24]/NET0131  , \u7_mem_reg[3][25]/NET0131  , \u7_mem_reg[3][26]/NET0131  , \u7_mem_reg[3][27]/NET0131  , \u7_mem_reg[3][28]/NET0131  , \u7_mem_reg[3][29]/NET0131  , \u7_mem_reg[3][2]/NET0131  , \u7_mem_reg[3][30]/NET0131  , \u7_mem_reg[3][31]/NET0131  , \u7_mem_reg[3][3]/NET0131  , \u7_mem_reg[3][4]/NET0131  , \u7_mem_reg[3][5]/NET0131  , \u7_mem_reg[3][6]/NET0131  , \u7_mem_reg[3][7]/NET0131  , \u7_mem_reg[3][8]/NET0131  , \u7_mem_reg[3][9]/NET0131  , \u7_rp_reg[0]/P0001  , \u7_rp_reg[1]/NET0131  , \u7_rp_reg[2]/NET0131  , \u7_rp_reg[3]/NET0131  , \u7_status_reg[0]/P0001  , \u7_status_reg[1]/P0001  , \u7_wp_reg[0]/P0001  , \u7_wp_reg[1]/NET0131  , \u7_wp_reg[2]/P0001  , \u8_dout_reg[0]/P0001  , \u8_dout_reg[10]/P0001  , \u8_dout_reg[11]/P0001  , \u8_dout_reg[12]/P0001  , \u8_dout_reg[13]/P0001  , \u8_dout_reg[14]/P0001  , \u8_dout_reg[15]/P0001  , \u8_dout_reg[16]/P0001  , \u8_dout_reg[17]/P0001  , \u8_dout_reg[18]/P0001  , \u8_dout_reg[19]/P0001  , \u8_dout_reg[1]/P0001  , \u8_dout_reg[2]/P0001  , \u8_dout_reg[3]/P0001  , \u8_dout_reg[4]/P0001  , \u8_dout_reg[5]/P0001  , \u8_dout_reg[6]/P0001  , \u8_dout_reg[7]/P0001  , \u8_dout_reg[8]/P0001  , \u8_dout_reg[9]/P0001  , \u8_empty_reg/NET0131  , \u8_mem_reg[0][0]/NET0131  , \u8_mem_reg[0][10]/NET0131  , \u8_mem_reg[0][11]/NET0131  , \u8_mem_reg[0][12]/NET0131  , \u8_mem_reg[0][13]/NET0131  , \u8_mem_reg[0][14]/NET0131  , \u8_mem_reg[0][15]/NET0131  , \u8_mem_reg[0][16]/NET0131  , \u8_mem_reg[0][17]/NET0131  , \u8_mem_reg[0][18]/NET0131  , \u8_mem_reg[0][19]/NET0131  , \u8_mem_reg[0][1]/NET0131  , \u8_mem_reg[0][20]/NET0131  , \u8_mem_reg[0][21]/NET0131  , \u8_mem_reg[0][22]/NET0131  , \u8_mem_reg[0][23]/NET0131  , \u8_mem_reg[0][24]/NET0131  , \u8_mem_reg[0][25]/NET0131  , \u8_mem_reg[0][26]/NET0131  , \u8_mem_reg[0][27]/NET0131  , \u8_mem_reg[0][28]/NET0131  , \u8_mem_reg[0][29]/NET0131  , \u8_mem_reg[0][2]/NET0131  , \u8_mem_reg[0][30]/NET0131  , \u8_mem_reg[0][31]/NET0131  , \u8_mem_reg[0][3]/NET0131  , \u8_mem_reg[0][4]/NET0131  , \u8_mem_reg[0][5]/NET0131  , \u8_mem_reg[0][6]/NET0131  , \u8_mem_reg[0][7]/NET0131  , \u8_mem_reg[0][8]/NET0131  , \u8_mem_reg[0][9]/NET0131  , \u8_mem_reg[1][0]/NET0131  , \u8_mem_reg[1][10]/NET0131  , \u8_mem_reg[1][11]/NET0131  , \u8_mem_reg[1][12]/NET0131  , \u8_mem_reg[1][13]/NET0131  , \u8_mem_reg[1][14]/NET0131  , \u8_mem_reg[1][15]/NET0131  , \u8_mem_reg[1][16]/NET0131  , \u8_mem_reg[1][17]/NET0131  , \u8_mem_reg[1][18]/NET0131  , \u8_mem_reg[1][19]/NET0131  , \u8_mem_reg[1][1]/NET0131  , \u8_mem_reg[1][20]/NET0131  , \u8_mem_reg[1][21]/NET0131  , \u8_mem_reg[1][22]/NET0131  , \u8_mem_reg[1][23]/NET0131  , \u8_mem_reg[1][24]/NET0131  , \u8_mem_reg[1][25]/NET0131  , \u8_mem_reg[1][26]/NET0131  , \u8_mem_reg[1][27]/NET0131  , \u8_mem_reg[1][28]/NET0131  , \u8_mem_reg[1][29]/NET0131  , \u8_mem_reg[1][2]/NET0131  , \u8_mem_reg[1][30]/NET0131  , \u8_mem_reg[1][31]/NET0131  , \u8_mem_reg[1][3]/NET0131  , \u8_mem_reg[1][4]/NET0131  , \u8_mem_reg[1][5]/NET0131  , \u8_mem_reg[1][6]/NET0131  , \u8_mem_reg[1][7]/NET0131  , \u8_mem_reg[1][8]/NET0131  , \u8_mem_reg[1][9]/NET0131  , \u8_mem_reg[2][0]/NET0131  , \u8_mem_reg[2][10]/NET0131  , \u8_mem_reg[2][11]/NET0131  , \u8_mem_reg[2][12]/NET0131  , \u8_mem_reg[2][13]/NET0131  , \u8_mem_reg[2][14]/NET0131  , \u8_mem_reg[2][15]/NET0131  , \u8_mem_reg[2][16]/NET0131  , \u8_mem_reg[2][17]/NET0131  , \u8_mem_reg[2][18]/NET0131  , \u8_mem_reg[2][19]/NET0131  , \u8_mem_reg[2][1]/NET0131  , \u8_mem_reg[2][20]/NET0131  , \u8_mem_reg[2][21]/NET0131  , \u8_mem_reg[2][22]/NET0131  , \u8_mem_reg[2][23]/NET0131  , \u8_mem_reg[2][24]/NET0131  , \u8_mem_reg[2][25]/NET0131  , \u8_mem_reg[2][26]/NET0131  , \u8_mem_reg[2][27]/NET0131  , \u8_mem_reg[2][28]/NET0131  , \u8_mem_reg[2][29]/NET0131  , \u8_mem_reg[2][2]/NET0131  , \u8_mem_reg[2][30]/NET0131  , \u8_mem_reg[2][31]/NET0131  , \u8_mem_reg[2][3]/NET0131  , \u8_mem_reg[2][4]/NET0131  , \u8_mem_reg[2][5]/NET0131  , \u8_mem_reg[2][6]/NET0131  , \u8_mem_reg[2][7]/NET0131  , \u8_mem_reg[2][8]/NET0131  , \u8_mem_reg[2][9]/NET0131  , \u8_mem_reg[3][0]/NET0131  , \u8_mem_reg[3][10]/NET0131  , \u8_mem_reg[3][11]/NET0131  , \u8_mem_reg[3][12]/NET0131  , \u8_mem_reg[3][13]/NET0131  , \u8_mem_reg[3][14]/NET0131  , \u8_mem_reg[3][15]/NET0131  , \u8_mem_reg[3][16]/NET0131  , \u8_mem_reg[3][17]/NET0131  , \u8_mem_reg[3][18]/NET0131  , \u8_mem_reg[3][19]/NET0131  , \u8_mem_reg[3][1]/NET0131  , \u8_mem_reg[3][20]/NET0131  , \u8_mem_reg[3][21]/NET0131  , \u8_mem_reg[3][22]/NET0131  , \u8_mem_reg[3][23]/NET0131  , \u8_mem_reg[3][24]/NET0131  , \u8_mem_reg[3][25]/NET0131  , \u8_mem_reg[3][26]/NET0131  , \u8_mem_reg[3][27]/NET0131  , \u8_mem_reg[3][28]/NET0131  , \u8_mem_reg[3][29]/NET0131  , \u8_mem_reg[3][2]/NET0131  , \u8_mem_reg[3][30]/NET0131  , \u8_mem_reg[3][31]/NET0131  , \u8_mem_reg[3][3]/NET0131  , \u8_mem_reg[3][4]/NET0131  , \u8_mem_reg[3][5]/NET0131  , \u8_mem_reg[3][6]/NET0131  , \u8_mem_reg[3][7]/NET0131  , \u8_mem_reg[3][8]/NET0131  , \u8_mem_reg[3][9]/NET0131  , \u8_rp_reg[0]/P0001  , \u8_rp_reg[1]/NET0131  , \u8_rp_reg[2]/NET0131  , \u8_rp_reg[3]/NET0131  , \u8_status_reg[0]/P0001  , \u8_status_reg[1]/P0001  , \u8_wp_reg[0]/P0001  , \u8_wp_reg[1]/NET0131  , \u8_wp_reg[2]/P0001  , \u9_din_tmp1_reg[0]/P0001  , \u9_din_tmp1_reg[10]/P0001  , \u9_din_tmp1_reg[11]/P0001  , \u9_din_tmp1_reg[12]/P0001  , \u9_din_tmp1_reg[13]/P0001  , \u9_din_tmp1_reg[14]/P0001  , \u9_din_tmp1_reg[15]/P0001  , \u9_din_tmp1_reg[1]/P0001  , \u9_din_tmp1_reg[2]/P0001  , \u9_din_tmp1_reg[3]/P0001  , \u9_din_tmp1_reg[4]/P0001  , \u9_din_tmp1_reg[5]/P0001  , \u9_din_tmp1_reg[6]/P0001  , \u9_din_tmp1_reg[7]/P0001  , \u9_din_tmp1_reg[8]/P0001  , \u9_din_tmp1_reg[9]/P0001  , \u9_dout_reg[0]/P0001  , \u9_dout_reg[10]/P0001  , \u9_dout_reg[11]/P0001  , \u9_dout_reg[12]/P0001  , \u9_dout_reg[13]/P0001  , \u9_dout_reg[14]/P0001  , \u9_dout_reg[15]/P0001  , \u9_dout_reg[16]/P0001  , \u9_dout_reg[17]/P0001  , \u9_dout_reg[18]/P0001  , \u9_dout_reg[19]/P0001  , \u9_dout_reg[1]/P0001  , \u9_dout_reg[20]/P0001  , \u9_dout_reg[21]/P0001  , \u9_dout_reg[22]/P0001  , \u9_dout_reg[23]/P0001  , \u9_dout_reg[24]/P0001  , \u9_dout_reg[25]/P0001  , \u9_dout_reg[26]/P0001  , \u9_dout_reg[27]/P0001  , \u9_dout_reg[28]/P0001  , \u9_dout_reg[29]/P0001  , \u9_dout_reg[2]/P0001  , \u9_dout_reg[30]/P0001  , \u9_dout_reg[31]/P0001  , \u9_dout_reg[3]/P0001  , \u9_dout_reg[4]/P0001  , \u9_dout_reg[5]/P0001  , \u9_dout_reg[6]/P0001  , \u9_dout_reg[7]/P0001  , \u9_dout_reg[8]/P0001  , \u9_dout_reg[9]/P0001  , \u9_empty_reg/P0001  , \u9_full_reg/NET0131  , \u9_mem_reg[0][0]/P0001  , \u9_mem_reg[0][10]/P0001  , \u9_mem_reg[0][11]/P0001  , \u9_mem_reg[0][12]/P0001  , \u9_mem_reg[0][13]/P0001  , \u9_mem_reg[0][14]/P0001  , \u9_mem_reg[0][15]/P0001  , \u9_mem_reg[0][16]/P0001  , \u9_mem_reg[0][17]/P0001  , \u9_mem_reg[0][18]/P0001  , \u9_mem_reg[0][19]/P0001  , \u9_mem_reg[0][1]/P0001  , \u9_mem_reg[0][20]/P0001  , \u9_mem_reg[0][21]/P0001  , \u9_mem_reg[0][22]/P0001  , \u9_mem_reg[0][23]/P0001  , \u9_mem_reg[0][24]/P0001  , \u9_mem_reg[0][25]/P0001  , \u9_mem_reg[0][26]/P0001  , \u9_mem_reg[0][27]/P0001  , \u9_mem_reg[0][28]/P0001  , \u9_mem_reg[0][29]/P0001  , \u9_mem_reg[0][2]/P0001  , \u9_mem_reg[0][30]/P0001  , \u9_mem_reg[0][31]/P0001  , \u9_mem_reg[0][3]/P0001  , \u9_mem_reg[0][4]/P0001  , \u9_mem_reg[0][5]/P0001  , \u9_mem_reg[0][6]/P0001  , \u9_mem_reg[0][7]/P0001  , \u9_mem_reg[0][8]/P0001  , \u9_mem_reg[0][9]/P0001  , \u9_mem_reg[1][0]/P0001  , \u9_mem_reg[1][10]/P0001  , \u9_mem_reg[1][11]/P0001  , \u9_mem_reg[1][12]/P0001  , \u9_mem_reg[1][13]/P0001  , \u9_mem_reg[1][14]/P0001  , \u9_mem_reg[1][15]/P0001  , \u9_mem_reg[1][16]/P0001  , \u9_mem_reg[1][17]/P0001  , \u9_mem_reg[1][18]/P0001  , \u9_mem_reg[1][19]/P0001  , \u9_mem_reg[1][1]/P0001  , \u9_mem_reg[1][20]/P0001  , \u9_mem_reg[1][21]/P0001  , \u9_mem_reg[1][22]/P0001  , \u9_mem_reg[1][23]/P0001  , \u9_mem_reg[1][24]/P0001  , \u9_mem_reg[1][25]/P0001  , \u9_mem_reg[1][26]/P0001  , \u9_mem_reg[1][27]/P0001  , \u9_mem_reg[1][28]/P0001  , \u9_mem_reg[1][29]/P0001  , \u9_mem_reg[1][2]/P0001  , \u9_mem_reg[1][30]/P0001  , \u9_mem_reg[1][31]/P0001  , \u9_mem_reg[1][3]/P0001  , \u9_mem_reg[1][4]/P0001  , \u9_mem_reg[1][5]/P0001  , \u9_mem_reg[1][6]/P0001  , \u9_mem_reg[1][7]/P0001  , \u9_mem_reg[1][8]/P0001  , \u9_mem_reg[1][9]/P0001  , \u9_mem_reg[2][0]/P0001  , \u9_mem_reg[2][10]/P0001  , \u9_mem_reg[2][11]/P0001  , \u9_mem_reg[2][12]/P0001  , \u9_mem_reg[2][13]/P0001  , \u9_mem_reg[2][14]/P0001  , \u9_mem_reg[2][15]/P0001  , \u9_mem_reg[2][16]/P0001  , \u9_mem_reg[2][17]/P0001  , \u9_mem_reg[2][18]/P0001  , \u9_mem_reg[2][19]/P0001  , \u9_mem_reg[2][1]/P0001  , \u9_mem_reg[2][20]/P0001  , \u9_mem_reg[2][21]/P0001  , \u9_mem_reg[2][22]/P0001  , \u9_mem_reg[2][23]/P0001  , \u9_mem_reg[2][24]/P0001  , \u9_mem_reg[2][25]/P0001  , \u9_mem_reg[2][26]/P0001  , \u9_mem_reg[2][27]/P0001  , \u9_mem_reg[2][28]/P0001  , \u9_mem_reg[2][29]/P0001  , \u9_mem_reg[2][2]/P0001  , \u9_mem_reg[2][30]/P0001  , \u9_mem_reg[2][31]/P0001  , \u9_mem_reg[2][3]/P0001  , \u9_mem_reg[2][4]/P0001  , \u9_mem_reg[2][5]/P0001  , \u9_mem_reg[2][6]/P0001  , \u9_mem_reg[2][7]/P0001  , \u9_mem_reg[2][8]/P0001  , \u9_mem_reg[2][9]/P0001  , \u9_mem_reg[3][0]/P0001  , \u9_mem_reg[3][10]/P0001  , \u9_mem_reg[3][11]/P0001  , \u9_mem_reg[3][12]/P0001  , \u9_mem_reg[3][13]/P0001  , \u9_mem_reg[3][14]/P0001  , \u9_mem_reg[3][15]/P0001  , \u9_mem_reg[3][16]/P0001  , \u9_mem_reg[3][17]/P0001  , \u9_mem_reg[3][18]/P0001  , \u9_mem_reg[3][19]/P0001  , \u9_mem_reg[3][1]/P0001  , \u9_mem_reg[3][20]/P0001  , \u9_mem_reg[3][21]/P0001  , \u9_mem_reg[3][22]/P0001  , \u9_mem_reg[3][23]/P0001  , \u9_mem_reg[3][24]/P0001  , \u9_mem_reg[3][25]/P0001  , \u9_mem_reg[3][26]/P0001  , \u9_mem_reg[3][27]/P0001  , \u9_mem_reg[3][28]/P0001  , \u9_mem_reg[3][29]/P0001  , \u9_mem_reg[3][2]/P0001  , \u9_mem_reg[3][30]/P0001  , \u9_mem_reg[3][31]/P0001  , \u9_mem_reg[3][3]/P0001  , \u9_mem_reg[3][4]/P0001  , \u9_mem_reg[3][5]/P0001  , \u9_mem_reg[3][6]/P0001  , \u9_mem_reg[3][7]/P0001  , \u9_mem_reg[3][8]/P0001  , \u9_mem_reg[3][9]/P0001  , \u9_rp_reg[0]/P0001  , \u9_rp_reg[1]/P0001  , \u9_rp_reg[2]/P0001  , \u9_status_reg[0]/P0001  , \u9_status_reg[1]/P0001  , \u9_wp_reg[0]/NET0131  , \u9_wp_reg[1]/P0001  , \u9_wp_reg[2]/P0001  , \u9_wp_reg[3]/P0001  , \valid_s_reg/NET0131  , wb_ack_o_pad , \wb_addr_i[29]_pad  , \wb_addr_i[2]_pad  , \wb_addr_i[30]_pad  , \wb_addr_i[31]_pad  , \wb_addr_i[3]_pad  , \wb_addr_i[4]_pad  , \wb_addr_i[5]_pad  , \wb_addr_i[6]_pad  , wb_cyc_i_pad , wb_stb_i_pad , wb_we_i_pad , \_al_n1  , \g16/_0_  , \g23/_0_  , \g29500/_0_  , \g29503/_3_  , \g29505/_3_  , \g29507/_3_  , \g29509/_3_  , \g29511/_0_  , \g29513/_3_  , \g29515/_3_  , \g29517/_3_  , \g29519/_0_  , \g29522/_0_  , \g29524/_0_  , \g29526/_0_  , \g29528/_0_  , \g29530/_0_  , \g29532/_0_  , \g29534/_3_  , \g29536/_3_  , \g29538/_3_  , \g29540/_3_  , \g29542/_3_  , \g29544/_3_  , \g29546/_3_  , \g29548/_3_  , \g29550/_0_  , \g29552/_0_  , \g29554/_0_  , \g29556/_0_  , \g29558/_0_  , \g29560/_0_  , \g29562/_0_  , \g29564/_0_  , \g29566/_0_  , \g29568/_0_  , \g29570/_0_  , \g29572/_0_  , \g29574/_3_  , \g29576/_3_  , \g29578/_3_  , \g29580/_3_  , \g29582/_3_  , \g29584/_3_  , \g29586/_3_  , \g29588/_3_  , \g29590/_3_  , \g29592/_3_  , \g29594/_3_  , \g29596/_3_  , \g29598/_3_  , \g29600/_3_  , \g29602/_3_  , \g29604/_3_  , \g29606/_0_  , \g29608/_0_  , \g29610/_0_  , \g29612/_0_  , \g29614/_3_  , \g29616/_3_  , \g29618/_3_  , \g29620/_3_  , \g29622/_3_  , \g29624/_3_  , \g29626/_3_  , \g29628/_3_  , \g29630/_3_  , \g29632/_3_  , \g29634/_3_  , \g29636/_3_  , \g29638/_3_  , \g29640/_3_  , \g29642/_3_  , \g29644/_3_  , \g29646/_3_  , \g29648/_3_  , \g29650/_3_  , \g29652/_3_  , \g29654/_3_  , \g29656/_3_  , \g29658/_3_  , \g29660/_3_  , \g29662/_3_  , \g29664/_3_  , \g29666/_3_  , \g29668/_3_  , \g29670/_3_  , \g29672/_3_  , \g29674/_3_  , \g29676/_3_  , \g29678/_3_  , \g29680/_3_  , \g29682/_3_  , \g29684/_3_  , \g29686/_3_  , \g29688/_3_  , \g29690/_3_  , \g29692/_3_  , \g29694/_0_  , \g29696/_0_  , \g29698/_0_  , \g29700/_0_  , \g29702/_0_  , \g29704/_0_  , \g29706/_0_  , \g29708/_0_  , \g29710/_0_  , \g29712/_0_  , \g29714/_0_  , \g29716/_0_  , \g29718/_0_  , \g29720/_0_  , \g29722/_0_  , \g29724/_0_  , \g29726/_0_  , \g29728/_0_  , \g29730/_0_  , \g29732/_0_  , \g29734/_3_  , \g29736/_3_  , \g29738/_3_  , \g29740/_3_  , \g29742/_3_  , \g29744/_3_  , \g29746/_3_  , \g29748/_3_  , \g29750/_3_  , \g29752/_3_  , \g29754/_3_  , \g29756/_3_  , \g29758/_3_  , \g29760/_3_  , \g29762/_3_  , \g29764/_3_  , \g29766/_3_  , \g29768/_3_  , \g29770/_3_  , \g29772/_3_  , \g29774/_3_  , \g29776/_3_  , \g29778/_3_  , \g29780/_3_  , \g29782/_3_  , \g29784/_3_  , \g29786/_3_  , \g29788/_3_  , \g29790/_3_  , \g29792/_3_  , \g29794/_3_  , \g29796/_3_  , \g29798/_3_  , \g29800/_3_  , \g29802/_3_  , \g29804/_3_  , \g29806/_3_  , \g29808/_3_  , \g29810/_3_  , \g29812/_3_  , \g29814/_3_  , \g29816/_3_  , \g29818/_3_  , \g29820/_3_  , \g29822/_3_  , \g29824/_3_  , \g29826/_3_  , \g29828/_3_  , \g29830/_3_  , \g29832/_3_  , \g29834/_3_  , \g29836/_3_  , \g29838/_3_  , \g29840/_3_  , \g29842/_3_  , \g29844/_3_  , \g29846/_3_  , \g29848/_3_  , \g29850/_3_  , \g29852/_3_  , \g29854/_3_  , \g29856/_3_  , \g29858/_3_  , \g29860/_3_  , \g29862/_3_  , \g29864/_3_  , \g29866/_3_  , \g29868/_3_  , \g29870/_3_  , \g29872/_3_  , \g29874/_3_  , \g29876/_3_  , \g29878/_3_  , \g29880/_3_  , \g29904/_0_  , \g29905/_0_  , \g29906/_0_  , \g29907/_0_  , \g29908/_0_  , \g29909/_0_  , \g29914/_3_  , \g29952/_0_  , \g29953/_0_  , \g29954/_0_  , \g29955/_0_  , \g29956/_0_  , \g29957/_0_  , \g29975/_0_  , \g29976/_0_  , \g29977/_0_  , \g29978/_0_  , \g29979/_0_  , \g29980/_0_  , \g29989/_3_  , \g30020/_0_  , \g30021/_0_  , \g30045/_0_  , \g30046/_0_  , \g30047/_0_  , \g30048/_0_  , \g30049/_0_  , \g30050/_0_  , \g30051/_0_  , \g30052/_0_  , \g30053/_0_  , \g30054/_0_  , \g30062/_0_  , \g30063/_0_  , \g30064/_0_  , \g30065/_0_  , \g30066/_0_  , \g30067/_0_  , \g30068/_0_  , \g30069/_0_  , \g30070/_0_  , \g30071/_0_  , \g30072/_0_  , \g30073/_0_  , \g30074/_0_  , \g30075/_0_  , \g30136/_3_  , \g30707/_0_  , \g30708/_0_  , \g30711/_0_  , \g30714/_0_  , \g30715/_0_  , \g30720/_0_  , \g30725/_0_  , \g30741/_0_  , \g30742/_0_  , \g30743/_0_  , \g30744/_0_  , \g30745/_0_  , \g30746/_0_  , \g30747/_0_  , \g30748/_0_  , \g30749/_0_  , \g30750/_0_  , \g30751/_0_  , \g30752/_0_  , \g30789/_0_  , \g30790/_0_  , \g30791/_0_  , \g30792/_0_  , \g30793/_0_  , \g30794/_0_  , \g30795/_0_  , \g30796/_0_  , \g30797/_0_  , \g30798/_0_  , \g30799/_0_  , \g30800/_0_  , \g30801/_0_  , \g30802/_0_  , \g30803/_0_  , \g30804/_0_  , \g30805/_0_  , \g30806/_0_  , \g30807/_0_  , \g30808/_0_  , \g30809/_0_  , \g30810/_0_  , \g30811/_0_  , \g30812/_0_  , \g30813/_0_  , \g30814/_0_  , \g30815/_0_  , \g30816/_0_  , \g30817/_0_  , \g30818/_0_  , \g30819/_0_  , \g30820/_0_  , \g30821/_0_  , \g30822/_0_  , \g30823/_0_  , \g30824/_0_  , \g30825/_0_  , \g30826/_0_  , \g30827/_0_  , \g30828/_0_  , \g30829/_0_  , \g30830/_0_  , \g30831/_0_  , \g30832/_0_  , \g30833/_0_  , \g30834/_0_  , \g30835/_0_  , \g30836/_0_  , \g30837/_0_  , \g30838/_0_  , \g30839/_0_  , \g30840/_0_  , \g30841/_0_  , \g30842/_0_  , \g30843/_0_  , \g30844/_0_  , \g30845/_0_  , \g30846/_0_  , \g30847/_0_  , \g30848/_0_  , \g30849/_0_  , \g30850/_0_  , \g30851/_0_  , \g30852/_0_  , \g30853/_0_  , \g30854/_0_  , \g30855/_0_  , \g30856/_0_  , \g30857/_0_  , \g30858/_0_  , \g30859/_0_  , \g30860/_0_  , \g30861/_0_  , \g30862/_0_  , \g30863/_0_  , \g30864/_0_  , \g30865/_0_  , \g30866/_0_  , \g30867/_0_  , \g30868/_0_  , \g30869/_0_  , \g30870/_0_  , \g30871/_0_  , \g30872/_0_  , \g30873/_0_  , \g30874/_0_  , \g30875/_0_  , \g30876/_0_  , \g30877/_0_  , \g30878/_0_  , \g30879/_0_  , \g30880/_0_  , \g30881/_0_  , \g30882/_0_  , \g30883/_0_  , \g30884/_0_  , \g30885/_0_  , \g30886/_0_  , \g30887/_0_  , \g30888/_0_  , \g30889/_0_  , \g30890/_0_  , \g30891/_0_  , \g30892/_0_  , \g30893/_0_  , \g30894/_0_  , \g30895/_0_  , \g30896/_0_  , \g30897/_0_  , \g30898/_0_  , \g30899/_0_  , \g30900/_0_  , \g30901/_0_  , \g30902/_0_  , \g30906/_0_  , \g30907/_0_  , \g30908/_0_  , \g30909/_0_  , \g30910/_0_  , \g30911/_0_  , \g30918/_0_  , \g30919/_0_  , \g30920/_0_  , \g30921/_0_  , \g30922/_0_  , \g30923/_0_  , \g30924/_0_  , \g30925/_0_  , \g30926/_0_  , \g30946/_0_  , \g30947/_0_  , \g30948/_0_  , \g30949/_0_  , \g30950/_0_  , \g30951/_0_  , \g30952/_0_  , \g30953/_0_  , \g30954/_0_  , \g30955/_0_  , \g30956/_0_  , \g30957/_0_  , \g30958/_0_  , \g30959/_0_  , \g30960/_0_  , \g30961/_0_  , \g30962/_0_  , \g30963/_0_  , \g30964/_0_  , \g30965/_0_  , \g30966/_0_  , \g30967/_0_  , \g30968/_0_  , \g30969/_0_  , \g30970/_0_  , \g30971/_0_  , \g30972/_0_  , \g30973/_0_  , \g30974/_0_  , \g30975/_0_  , \g30976/_0_  , \g30977/_0_  , \g30978/_0_  , \g30979/_0_  , \g30980/_0_  , \g30981/_0_  , \g30982/_0_  , \g30983/_0_  , \g30984/_0_  , \g30985/_0_  , \g30986/_0_  , \g30987/_0_  , \g30988/_0_  , \g30989/_0_  , \g30990/_0_  , \g30991/_0_  , \g30992/_0_  , \g30993/_0_  , \g30994/_0_  , \g30995/_0_  , \g30996/_0_  , \g30997/_0_  , \g30998/_0_  , \g30999/_0_  , \g31000/_0_  , \g31001/_0_  , \g31002/_0_  , \g31003/_0_  , \g31004/_0_  , \g31005/_0_  , \g31006/_0_  , \g31007/_0_  , \g31008/_0_  , \g31009/_0_  , \g31010/_0_  , \g31011/_0_  , \g31012/_0_  , \g31013/_0_  , \g31014/_0_  , \g31015/_0_  , \g31016/_0_  , \g31017/_0_  , \g31018/_0_  , \g31019/_0_  , \g31020/_0_  , \g31021/_0_  , \g31022/_0_  , \g31023/_0_  , \g31024/_0_  , \g31025/_0_  , \g31026/_0_  , \g31027/_0_  , \g31028/_0_  , \g31029/_0_  , \g31030/_0_  , \g31031/_0_  , \g31032/_0_  , \g31033/_0_  , \g31034/_0_  , \g31035/_0_  , \g31036/_0_  , \g31037/_0_  , \g31038/_0_  , \g31039/_0_  , \g31040/_0_  , \g31041/_0_  , \g31042/_0_  , \g31043/_0_  , \g31044/_0_  , \g31045/_0_  , \g31046/_0_  , \g31047/_0_  , \g31048/_0_  , \g31049/_0_  , \g31050/_0_  , \g31051/_0_  , \g31052/_0_  , \g31053/_0_  , \g31054/_0_  , \g31055/_0_  , \g31056/_0_  , \g31057/_0_  , \g31058/_0_  , \g31059/_0_  , \g31060/_0_  , \g31061/_0_  , \g31062/_0_  , \g31063/_0_  , \g31064/_0_  , \g31065/_0_  , \g31066/_0_  , \g31067/_0_  , \g31068/_0_  , \g31069/_0_  , \g31070/_0_  , \g31071/_0_  , \g31072/_0_  , \g31073/_0_  , \g31074/_0_  , \g31075/_0_  , \g31076/_0_  , \g31077/_0_  , \g31084/u3_syn_4  , \g31085/u3_syn_4  , \g31096/u3_syn_4  , \g31115/u3_syn_4  , \g31136/u3_syn_4  , \g31158/u3_syn_4  , \g31176/u3_syn_4  , \g31193/u3_syn_4  , \g31195/u3_syn_4  , \g31247/u3_syn_4  , \g31280/u3_syn_4  , \g31285/u3_syn_4  , \g31568/_0_  , \g31631/_0_  , \g31672/_0_  , \g31731/_0_  , \g31732/_0_  , \g31742/_2_  , \g31744/_2_  , \g31746/_2_  , \g31748/_2_  , \g31751/_2_  , \g31754/_2_  , \g31756/_2_  , \g31758/_2_  , \g31760/_2_  , \g31761/_0_  , \g31789/_0_  , \g31807/_3_  , \g31825/_3_  , \g32607/_0_  , \g32608/_0_  , \g32609/_0_  , \g32610/_0_  , \g32611/_0_  , \g32612/_0_  , \g32613/_0_  , \g32614/_0_  , \g32615/_0_  , \g32616/_0_  , \g32617/_0_  , \g32618/_0_  , \g32645/_0__syn_2  , \g32687/_0__syn_2  , \g32749/_0__syn_2  , \g32757/_0_  , \g32758/_0_  , \g32759/_0_  , \g32760/_0_  , \g32761/_0_  , \g32762/_0_  , \g32763/_0_  , \g32764/_0_  , \g32765/_0_  , \g32769/_0_  , \g32835/_1_  , \g32839/_0_  , \g32844/_0_  , \g32901/_1_  , \g32902/_0_  , \g32963/_1_  , \g32972/_0_  , \g32977/_0_  , \g32979/_0_  , \g32980/_0_  , \g32981/_0_  , \g32982/_0_  , \g32983/_0_  , \g32987/_0_  , \g33018/_0_  , \g33019/_0_  , \g33088/_0_  , \g33261/_0_  , \g33264/_0_  , \g33275/_0_  , \g33276/_0_  , \g33277/_0_  , \g33371/_0_  , \g33382/_0_  , \g33401/_0_  , \g33402/_0_  , \g33403/_0_  , \g33404/_0_  , \g33405/_0_  , \g33406/_0_  , \g33407/_0_  , \g33408/_0_  , \g33409/_0_  , \g33410/_0_  , \g33411/_0_  , \g33412/_0_  , \g33413/_0_  , \g33414/_0_  , \g33415/_0_  , \g33416/_0_  , \g33417/_0_  , \g33418/_0_  , \g33419/_0_  , \g33420/_0_  , \g33421/_0_  , \g33422/_0_  , \g33423/_0_  , \g33424/_0_  , \g33425/_0_  , \g33426/_0_  , \g33427/_0_  , \g33428/_0_  , \g33429/_0_  , \g33430/_0_  , \g33431/_0_  , \g33432/_0_  , \g33433/_0_  , \g33434/_0_  , \g33435/_0_  , \g33436/_0_  , \g33437/_0_  , \g33438/_0_  , \g33439/_0_  , \g33440/_0_  , \g33441/_0_  , \g33442/_0_  , \g33443/_0_  , \g33444/_0_  , \g33445/_0_  , \g33446/_0_  , \g33447/_0_  , \g33448/_0_  , \g33449/_0_  , \g33450/_0_  , \g33451/_0_  , \g33452/_0_  , \g33453/_0_  , \g33454/_0_  , \g33455/_0_  , \g33456/_0_  , \g33457/_0_  , \g33458/_0_  , \g33459/_0_  , \g33460/_0_  , \g33461/_0_  , \g33462/_0_  , \g33463/_0_  , \g33464/_0_  , \g33465/_0_  , \g33466/_0_  , \g33467/_0_  , \g33468/_0_  , \g33469/_0_  , \g33470/_0_  , \g33471/_0_  , \g33472/_0_  , \g33473/_0_  , \g33474/_0_  , \g33475/_0_  , \g33476/_0_  , \g33477/_0_  , \g33478/_0_  , \g33479/_0_  , \g33480/_0_  , \g33481/_0_  , \g33482/_0_  , \g33483/_0_  , \g33484/_0_  , \g33485/_0_  , \g33486/_0_  , \g33487/_0_  , \g33488/_0_  , \g33489/_0_  , \g33490/_0_  , \g33491/_0_  , \g33492/_0_  , \g33493/_0_  , \g33494/_0_  , \g33495/_0_  , \g33496/_0_  , \g33497/_0_  , \g33498/_0_  , \g33499/_0_  , \g33500/_0_  , \g33501/_0_  , \g33502/_0_  , \g33503/_0_  , \g33504/_0_  , \g33505/_0_  , \g33506/_0_  , \g33507/_0_  , \g33508/_0_  , \g33509/_0_  , \g33510/_0_  , \g33511/_0_  , \g33512/_0_  , \g33513/_0_  , \g33514/_0_  , \g33515/_0_  , \g33516/_0_  , \g33517/_0_  , \g33518/_0_  , \g33519/_0_  , \g33520/_0_  , \g33521/_0_  , \g33522/_0_  , \g33523/_0_  , \g33524/_0_  , \g33525/_0_  , \g33526/_0_  , \g33527/_0_  , \g33528/_0_  , \g33529/_0_  , \g33530/_0_  , \g33531/_0_  , \g33532/_0_  , \g33533/_0_  , \g33534/_0_  , \g33535/_0_  , \g33536/_0_  , \g33537/_0_  , \g33538/_0_  , \g33539/_0_  , \g33540/_0_  , \g33541/_0_  , \g33542/_0_  , \g33543/_0_  , \g33544/_0_  , \g33545/_0_  , \g33546/_0_  , \g33547/_0_  , \g33548/_0_  , \g33549/_0_  , \g33550/_0_  , \g33551/_0_  , \g33552/_0_  , \g33553/_0_  , \g33554/_0_  , \g33555/_0_  , \g33556/_0_  , \g33557/_0_  , \g33558/_0_  , \g33559/_0_  , \g33560/_0_  , \g33561/_0_  , \g33562/_0_  , \g33563/_0_  , \g33564/_0_  , \g33565/_0_  , \g33566/_0_  , \g33567/_0_  , \g33568/_0_  , \g33569/_0_  , \g33570/_0_  , \g33571/_0_  , \g33572/_0_  , \g33573/_0_  , \g33574/_0_  , \g33575/_0_  , \g33576/_0_  , \g33577/_0_  , \g33578/_0_  , \g33579/_0_  , \g33580/_0_  , \g33581/_0_  , \g33582/_0_  , \g33583/_0_  , \g33584/_0_  , \g33585/_0_  , \g33586/_0_  , \g33587/_0_  , \g33588/_0_  , \g33589/_0_  , \g33590/_0_  , \g33591/_0_  , \g33592/_0_  , \g33593/_0_  , \g33594/_0_  , \g33595/_0_  , \g33596/_0_  , \g33597/_0_  , \g33598/_0_  , \g33599/_0_  , \g33600/_0_  , \g33601/_0_  , \g33602/_0_  , \g33603/_0_  , \g33604/_0_  , \g33605/_0_  , \g33606/_0_  , \g33607/_0_  , \g33608/_0_  , \g33609/_0_  , \g33610/_0_  , \g33611/_0_  , \g33612/_0_  , \g33613/_0_  , \g33614/_0_  , \g33615/_0_  , \g33616/_0_  , \g33617/_0_  , \g33618/_0_  , \g33619/_0_  , \g33620/_0_  , \g33621/_0_  , \g33622/_0_  , \g33623/_0_  , \g33624/_0_  , \g33625/_0_  , \g33626/_0_  , \g33627/_0_  , \g33628/_0_  , \g33629/_0_  , \g33630/_0_  , \g33631/_0_  , \g33632/_0_  , \g33633/_0_  , \g33634/_0_  , \g33635/_0_  , \g33636/_0_  , \g33637/_0_  , \g33638/_0_  , \g33639/_0_  , \g33640/_0_  , \g33641/_0_  , \g33642/_0_  , \g33643/_0_  , \g33644/_0_  , \g33645/_0_  , \g33646/_0_  , \g33647/_0_  , \g33648/_0_  , \g33649/_0_  , \g33650/_0_  , \g33651/_0_  , \g33652/_0_  , \g33653/_0_  , \g33654/_0_  , \g33655/_0_  , \g33656/_0_  , \g33657/_0_  , \g33658/_0_  , \g33659/_0_  , \g33660/_0_  , \g33661/_0_  , \g33662/_0_  , \g33663/_0_  , \g33664/_0_  , \g33665/_0_  , \g33666/_0_  , \g33667/_0_  , \g33668/_0_  , \g33669/_0_  , \g33670/_0_  , \g33671/_0_  , \g33672/_0_  , \g33673/_0_  , \g33674/_0_  , \g33675/_0_  , \g33676/_0_  , \g33677/_0_  , \g33678/_0_  , \g33679/_0_  , \g33680/_0_  , \g33681/_0_  , \g33682/_0_  , \g33683/_0_  , \g33684/_0_  , \g33685/_0_  , \g33686/_0_  , \g33687/_0_  , \g33688/_0_  , \g33689/_0_  , \g33690/_0_  , \g33691/_0_  , \g33692/_0_  , \g33693/_0_  , \g33694/_0_  , \g33695/_0_  , \g33696/_0_  , \g33697/_0_  , \g33698/_0_  , \g33699/_0_  , \g33700/_0_  , \g33701/_0_  , \g33702/_0_  , \g33703/_0_  , \g33704/_0_  , \g33705/_0_  , \g33706/_0_  , \g33707/_0_  , \g33708/_0_  , \g33709/_0_  , \g33710/_0_  , \g33711/_0_  , \g33712/_0_  , \g33713/_0_  , \g33714/_0_  , \g33715/_0_  , \g33716/_0_  , \g33717/_0_  , \g33718/_0_  , \g33719/_0_  , \g33720/_0_  , \g33721/_0_  , \g33722/_0_  , \g33723/_0_  , \g33724/_0_  , \g33725/_0_  , \g33726/_0_  , \g33727/_0_  , \g33728/_0_  , \g33729/_0_  , \g33730/_0_  , \g33731/_0_  , \g33732/_0_  , \g33733/_0_  , \g33734/_0_  , \g33735/_0_  , \g33736/_0_  , \g33737/_0_  , \g33738/_0_  , \g33739/_0_  , \g33740/_0_  , \g33741/_0_  , \g33742/_0_  , \g33743/_0_  , \g33744/_0_  , \g33745/_0_  , \g33746/_0_  , \g33747/_0_  , \g33748/_0_  , \g33749/_0_  , \g33750/_0_  , \g33751/_0_  , \g33752/_0_  , \g33753/_0_  , \g33754/_0_  , \g33755/_0_  , \g33756/_0_  , \g33757/_0_  , \g33758/_0_  , \g33759/_0_  , \g33760/_0_  , \g33761/_0_  , \g33762/_0_  , \g33763/_0_  , \g33764/_0_  , \g33765/_0_  , \g33766/_0_  , \g33767/_0_  , \g33768/_0_  , \g33769/_0_  , \g33770/_0_  , \g33771/_0_  , \g33772/_0_  , \g33773/_0_  , \g33774/_0_  , \g33775/_0_  , \g33776/_0_  , \g33777/_0_  , \g33778/_0_  , \g33779/_0_  , \g33780/_0_  , \g33781/_0_  , \g33782/_0_  , \g33783/_0_  , \g33784/_0_  , \g33785/_0_  , \g33786/_0_  , \g33787/_0_  , \g33788/_0_  , \g33789/_0_  , \g33790/_0_  , \g33791/_0_  , \g33792/_0_  , \g33793/_0_  , \g33794/_0_  , \g33795/_0_  , \g33796/_0_  , \g33797/_0_  , \g33798/_0_  , \g33799/_0_  , \g33800/_0_  , \g33801/_0_  , \g33802/_0_  , \g33803/_0_  , \g33804/_0_  , \g33805/_0_  , \g33806/_0_  , \g33807/_0_  , \g33808/_0_  , \g33809/_0_  , \g33810/_0_  , \g33811/_0_  , \g33812/_0_  , \g33813/_0_  , \g33814/_0_  , \g33815/_0_  , \g33816/_0_  , \g33817/_0_  , \g33818/_0_  , \g33819/_0_  , \g33820/_0_  , \g33821/_0_  , \g33822/_0_  , \g33823/_0_  , \g33824/_0_  , \g33825/_0_  , \g33826/_0_  , \g33827/_0_  , \g33828/_0_  , \g33829/_0_  , \g33830/_0_  , \g33831/_0_  , \g33832/_0_  , \g33833/_0_  , \g33834/_0_  , \g33835/_0_  , \g33836/_0_  , \g33837/_0_  , \g33838/_0_  , \g33839/_0_  , \g33840/_0_  , \g33841/_0_  , \g33842/_0_  , \g33843/_0_  , \g33844/_0_  , \g33845/_0_  , \g33846/_0_  , \g33847/_0_  , \g33848/_0_  , \g33849/_0_  , \g33850/_0_  , \g33851/_0_  , \g33852/_0_  , \g33853/_0_  , \g33854/_0_  , \g33855/_0_  , \g33856/_0_  , \g33857/_0_  , \g33858/_0_  , \g33859/_0_  , \g33860/_0_  , \g33861/_0_  , \g33862/_0_  , \g33863/_0_  , \g33864/_0_  , \g33865/_0_  , \g33866/_0_  , \g33867/_0_  , \g33868/_0_  , \g33869/_0_  , \g33870/_0_  , \g33871/_0_  , \g33872/_0_  , \g33873/_0_  , \g33874/_0_  , \g33875/_0_  , \g33876/_0_  , \g33877/_0_  , \g33878/_0_  , \g33879/_0_  , \g33880/_0_  , \g33881/_0_  , \g33882/_0_  , \g33883/_0_  , \g33884/_0_  , \g33885/_0_  , \g33886/_0_  , \g33887/_0_  , \g33888/_0_  , \g33889/_0_  , \g33890/_0_  , \g33891/_0_  , \g33892/_0_  , \g33893/_0_  , \g33894/_0_  , \g33895/_0_  , \g33896/_0_  , \g33897/_0_  , \g33898/_0_  , \g33899/_0_  , \g33900/_0_  , \g33901/_0_  , \g33902/_0_  , \g33903/_0_  , \g33904/_0_  , \g33905/_0_  , \g33906/_0_  , \g33907/_0_  , \g33908/_0_  , \g33909/_0_  , \g33910/_0_  , \g33911/_0_  , \g33912/_0_  , \g33913/_0_  , \g33914/_0_  , \g33915/_0_  , \g33916/_0_  , \g33917/_0_  , \g33918/_0_  , \g33919/_0_  , \g33920/_0_  , \g33921/_0_  , \g33922/_0_  , \g33923/_0_  , \g33924/_0_  , \g33925/_0_  , \g33926/_0_  , \g33927/_0_  , \g33928/_0_  , \g33929/_0_  , \g33930/_0_  , \g33931/_0_  , \g33932/_0_  , \g33933/_0_  , \g33934/_0_  , \g33935/_0_  , \g33936/_0_  , \g33937/_0_  , \g33938/_0_  , \g33939/_0_  , \g33940/_0_  , \g33941/_0_  , \g33942/_0_  , \g33943/_0_  , \g33944/_0_  , \g33945/_0_  , \g33946/_0_  , \g33947/_0_  , \g33948/_0_  , \g33949/_0_  , \g33950/_0_  , \g33951/_0_  , \g33952/_0_  , \g33953/_0_  , \g33954/_0_  , \g33955/_0_  , \g33956/_0_  , \g33957/_0_  , \g33958/_0_  , \g33959/_0_  , \g33960/_0_  , \g33961/_0_  , \g33962/_0_  , \g33963/_0_  , \g33964/_0_  , \g33965/_0_  , \g33966/_0_  , \g33967/_0_  , \g33968/_0_  , \g33969/_0_  , \g33970/_0_  , \g33971/_0_  , \g33972/_0_  , \g33973/_0_  , \g33974/_0_  , \g33975/_0_  , \g33976/_0_  , \g33977/u3_syn_4  , \g33981/u3_syn_4  , \g34014/u3_syn_4  , \g34047/u3_syn_4  , \g34084/u3_syn_4  , \g34123/u3_syn_4  , \g34306/_0_  , \g34316/_0_  , \g34324/_0_  , \g34326/_0_  , \g34328/_0_  , \g34331/_0_  , \g34333/_0_  , \g34344/_0_  , \g34347/_0_  , \g34351/_0_  , \g34361/_0_  , \g34368/_0_  , \g34377/_0_  , \g34385/_0_  , \g34393/_0_  , \g34414/_1_  , \g34451/_1_  , \g34476/_1_  , \g34487/_0_  , \g34490/_1_  , \g34715/_0_  , \g34878/_0_  , \g34882/_0_  , \g34883/_0_  , \g34893/_0_  , \g34896/_0_  , \g34898/_0_  , \g34899/_0_  , \g34916/_3_  , \g35264/_0_  , \g35265/_0_  , \g35266/_0_  , \g35267/_0_  , \g35268/_0_  , \g35269/_0_  , \g35270/_0_  , \g35271/_0_  , \g35272/_0_  , \g35273/_0_  , \g35274/_0_  , \g35275/_0_  , \g35276/_0_  , \g35277/_0_  , \g35278/_0_  , \g35279/_0_  , \g35283/_0_  , \g35287/_0_  , \g35294/_0_  , \g35300/_0_  , \g35304/_0_  , \g35308/_0_  , \g35312/_0_  , \g35316/_0_  , \g35318/_0_  , \g35326/_0_  , \g35334/_0_  , \g35336/_0_  , \g35337/_0_  , \g35338/_0_  , \g35357/_0_  , \g35358/_0_  , \g35359/_0_  , \g35419/_0_  , \g35438/_0_  , \g35439/_0_  , \g35440/_0_  , \g35441/_0_  , \g35442/_0_  , \g35444/_0_  , \g35445/_0_  , \g35446/_0_  , \g35447/_0_  , \g35448/_0_  , \g35449/_0_  , \g35450/_0_  , \g35451/_0_  , \g35452/_0_  , \g35463/_0_  , \g35464/_0_  , \g35466/_0_  , \g35485/_2_  , \g35495/_0_  , \g35496/_0_  , \g35499/_0_  , \g35500/_0_  , \g35501/_0_  , \g35502/_0_  , \g35563/_0_  , \g35633/_0_  , \g35717/_0_  , \g35718/_0_  , \g35719/_0_  , \g35809/_0_  , \g35810/_0_  , \g35811/_0_  , \g35812/_0_  , \g35813/_0_  , \g35814/_0_  , \g35815/_0_  , \g35816/_0_  , \g35817/_0_  , \g35818/_0_  , \g35819/_0_  , \g35820/_0_  , \g35821/_0_  , \g35822/_0_  , \g35823/_0_  , \g35824/_0_  , \g35825/_0_  , \g35826/_0_  , \g35827/_0_  , \g35830/_0_  , \g35833/_0_  , \g35835/_0_  , \g35836/_0_  , \g35837/_0_  , \g35839/_0_  , \g35840/_0_  , \g35841/_0_  , \g35843/_0_  , \g35844/_0_  , \g35845/_0_  , \g35853/_0_  , \g35854/_0_  , \g35855/_0_  , \g35856/_0_  , \g36306/_0_  , \g36414/_0_  , \g36415/_0_  , \g36449/_0_  , \g36550/_0_  , \g36551/_0_  , \g36553/_0_  , \g36560/_0_  , \g36562/_3_  , \g36563/_0_  , \g36612/_0_  , \g36614/_2_  , \g36695/_0_  , \g36784/_0_  , \g36785/_0_  , \g36786/_0_  , \g36787/_0_  , \g36788/_0_  , \g36789/_0_  , \g36790/_0_  , \g36791/_0_  , \g36792/_0_  , \g36793/_0_  , \g36794/_0_  , \g36796/_0_  , \g36797/_0_  , \g36798/_0_  , \g36799/_0_  , \g36800/_0_  , \g36801/_0_  , \g36802/_0_  , \g36803/_0_  , \g36804/_0_  , \g36805/_0_  , \g36806/_0_  , \g36807/_0_  , \g36808/_0_  , \g36809/_0_  , \g36810/_0_  , \g36811/_0_  , \g36813/_0_  , \g36814/_0_  , \g36815/_0_  , \g36820/_0_  , \g36825/_0_  , \g36832/_0_  , \g36846/_0_  , \g36855/_0_  , \g36857/_0_  , \g36859/_0_  , \g36860/_0_  , \g36861/_0_  , \g36862/_0_  , \g36863/_0_  , \g36864/_0_  , \g36867/_0_  , \g36870/_0_  , \g36871/_0_  , \g36877/_0_  , \g36879/_0_  , \g36892/_0_  , \g36893/_0_  , \g36901/_0_  , \g36909/_0_  , \g36914/_0_  , \g36919/_0_  , \g36922/_0_  , \g36923/_0_  , \g36927/_0_  , \g36930/_0_  , \g36931/_0_  , \g36933/_0_  , \g36934/_0_  , \g36935/_0_  , \g36936/_0_  , \g36937/_0_  , \g36938/_0_  , \g36939/_0_  , \g36940/_0_  , \g36941/_0_  , \g36943/_0_  , \g36944/_0_  , \g36945/_0_  , \g36946/_0_  , \g36947/_0_  , \g36948/_0_  , \g36949/_0_  , \g36950/_0_  , \g36951/_0_  , \g36952/_0_  , \g36953/_0_  , \g36954/_0_  , \g36957/_0_  , \g36958/_0_  , \g36959/_0_  , \g36960/_0_  , \g36961/_0_  , \g36962/_0_  , \g36963/_0_  , \g36970/_0_  , \g36977/_0_  , \g36986/_0_  , \g36991/_0_  , \g36994/_0_  , \g37015/_0_  , \g37057/_0_  , \g37073/_0_  , \g37128/_0_  , \g37129/_0_  , \g37138/_0_  , \g37139/_0_  , \g37140/_0_  , \g37141/_0_  , \g37142/_0_  , \g37143/_0_  , \g37144/_0_  , \g37145/_0_  , \g37146/_0_  , \g37147/_0_  , \g37148/_0_  , \g37149/_0_  , \g37150/_0_  , \g37151/_0_  , \g37152/_0_  , \g37153/_0_  , \g37154/_0_  , \g37155/_0_  , \g37156/_0_  , \g37157/_0_  , \g37158/_0_  , \g37159/_0_  , \g37160/_0_  , \g37161/_0_  , \g37162/_0_  , \g37163/_0_  , \g37164/_0_  , \g37165/_0_  , \g37166/_0_  , \g37167/_0_  , \g37168/_0_  , \g37169/_0_  , \g37170/_0_  , \g37171/_0_  , \g37172/_0_  , \g37173/_0_  , \g37174/_0_  , \g37175/_0_  , \g37176/_0_  , \g37177/_0_  , \g37178/_0_  , \g37179/_0_  , \g37180/_0_  , \g37181/_0_  , \g37182/_0_  , \g37183/_0_  , \g37184/_0_  , \g37185/_0_  , \g37187/_0_  , \g37188/_0_  , \g37190/_0_  , \g37191/_0_  , \g37192/_0_  , \g37193/_0_  , \g37194/_0_  , \g37372/_3_  , \g37377/_0_  , \g37378/_0_  , \g37379/_0_  , \g37380/_0_  , \g37381/_0_  , \g37382/_0_  , \g37383/_0_  , \g37384/_0_  , \g37385/_0_  , \g37386/_0_  , \g37387/_0_  , \g37388/_0_  , \g37389/_0_  , \g37390/_0_  , \g37391/_0_  , \g37392/_0_  , \g37393/_0_  , \g37394/_0_  , \g37395/_0_  , \g37396/_0_  , \g37397/_0_  , \g37398/_0_  , \g37399/_0_  , \g37400/_0_  , \g37401/_0_  , \g37402/_0_  , \g37403/_0_  , \g37404/_0_  , \g37405/_0_  , \g37406/_0_  , \g37407/_0_  , \g37408/_0_  , \g37409/_0_  , \g37410/_0_  , \g37411/_0_  , \g37412/_0_  , \g37413/_0_  , \g37576/_3_  , \g37590/_2_  , \g40278/_0_  , \g40379/_0_  , \g40389/_2_  , \g40390/_2_  , \g40391/_0_  , \g40393/_2_  , \g40395/_0_  , \g40397/_0_  , \g40400/_0_  , \g40402/_0_  , \g45458/_0_  , \g45675/_0_  , \g45677/_0_  , \g45678/_0_  , \g45682/_0_  , sync_pad_o_pad , \u14_u0_full_empty_r_reg/P0001_reg_syn_3  , \u14_u1_full_empty_r_reg/P0001_reg_syn_3  , \u14_u2_full_empty_r_reg/P0001_reg_syn_3  , \u14_u3_full_empty_r_reg/P0001_reg_syn_3  , \u14_u4_full_empty_r_reg/P0001_reg_syn_3  , \u14_u5_full_empty_r_reg/P0001_reg_syn_3  , \u14_u6_full_empty_r_reg/P0001_reg_syn_3  , \u14_u7_full_empty_r_reg/P0001_reg_syn_3  , \u14_u8_full_empty_r_reg/P0001_reg_syn_3  , \u1_slt0_reg[11]/P0001_reg_syn_3  , \u1_slt0_reg[12]/P0001_reg_syn_3  , \u1_slt0_reg[15]/P0001_reg_syn_3  , \u1_slt0_reg[9]/P0001_reg_syn_3  , \u1_slt1_reg[10]/P0001_reg_syn_3  , \u1_slt1_reg[11]/P0001_reg_syn_3  , \u1_slt1_reg[5]/P0001_reg_syn_3  , \u1_slt1_reg[6]/P0001_reg_syn_3  , \u1_slt1_reg[7]/P0001_reg_syn_3  , \u1_slt1_reg[8]/P0001_reg_syn_3  , wb_err_o_pad );
  input \ac97_reset_pad_o__pad  ;
  input \dma_ack_i[0]_pad  ;
  input \dma_ack_i[1]_pad  ;
  input \dma_ack_i[2]_pad  ;
  input \dma_ack_i[3]_pad  ;
  input \dma_ack_i[4]_pad  ;
  input \dma_ack_i[5]_pad  ;
  input \dma_ack_i[6]_pad  ;
  input \dma_ack_i[7]_pad  ;
  input \dma_ack_i[8]_pad  ;
  input \dma_req_o[0]_pad  ;
  input \dma_req_o[1]_pad  ;
  input \dma_req_o[2]_pad  ;
  input \dma_req_o[3]_pad  ;
  input \dma_req_o[4]_pad  ;
  input \dma_req_o[5]_pad  ;
  input \dma_req_o[6]_pad  ;
  input \dma_req_o[7]_pad  ;
  input \dma_req_o[8]_pad  ;
  input \in_valid_s_reg[0]/NET0131  ;
  input \in_valid_s_reg[1]/NET0131  ;
  input \in_valid_s_reg[2]/NET0131  ;
  input suspended_o_pad ;
  input \u0_slt0_r_reg[0]/P0001  ;
  input \u0_slt0_r_reg[10]/P0001  ;
  input \u0_slt0_r_reg[11]/P0001  ;
  input \u0_slt0_r_reg[12]/P0001  ;
  input \u0_slt0_r_reg[13]/P0001  ;
  input \u0_slt0_r_reg[14]/P0001  ;
  input \u0_slt0_r_reg[1]/P0001  ;
  input \u0_slt0_r_reg[2]/P0001  ;
  input \u0_slt0_r_reg[3]/P0001  ;
  input \u0_slt0_r_reg[4]/P0001  ;
  input \u0_slt0_r_reg[5]/P0001  ;
  input \u0_slt0_r_reg[6]/P0001  ;
  input \u0_slt0_r_reg[7]/P0001  ;
  input \u0_slt0_r_reg[8]/P0001  ;
  input \u0_slt0_r_reg[9]/P0001  ;
  input \u0_slt1_r_reg[0]/P0001  ;
  input \u0_slt1_r_reg[10]/P0001  ;
  input \u0_slt1_r_reg[11]/P0001  ;
  input \u0_slt1_r_reg[12]/P0001  ;
  input \u0_slt1_r_reg[13]/P0001  ;
  input \u0_slt1_r_reg[14]/P0001  ;
  input \u0_slt1_r_reg[15]/P0001  ;
  input \u0_slt1_r_reg[16]/P0001  ;
  input \u0_slt1_r_reg[17]/P0001  ;
  input \u0_slt1_r_reg[18]/P0001  ;
  input \u0_slt1_r_reg[19]/P0001  ;
  input \u0_slt1_r_reg[1]/P0001  ;
  input \u0_slt1_r_reg[2]/P0001  ;
  input \u0_slt1_r_reg[3]/P0001  ;
  input \u0_slt1_r_reg[4]/P0001  ;
  input \u0_slt1_r_reg[5]/P0001  ;
  input \u0_slt1_r_reg[6]/P0001  ;
  input \u0_slt1_r_reg[7]/P0001  ;
  input \u0_slt1_r_reg[8]/P0001  ;
  input \u0_slt1_r_reg[9]/P0001  ;
  input \u0_slt2_r_reg[0]/P0001  ;
  input \u0_slt2_r_reg[10]/P0001  ;
  input \u0_slt2_r_reg[11]/P0001  ;
  input \u0_slt2_r_reg[12]/P0001  ;
  input \u0_slt2_r_reg[13]/P0001  ;
  input \u0_slt2_r_reg[14]/P0001  ;
  input \u0_slt2_r_reg[15]/P0001  ;
  input \u0_slt2_r_reg[16]/P0001  ;
  input \u0_slt2_r_reg[17]/P0001  ;
  input \u0_slt2_r_reg[18]/P0001  ;
  input \u0_slt2_r_reg[19]/P0001  ;
  input \u0_slt2_r_reg[1]/P0001  ;
  input \u0_slt2_r_reg[2]/P0001  ;
  input \u0_slt2_r_reg[3]/P0001  ;
  input \u0_slt2_r_reg[4]/P0001  ;
  input \u0_slt2_r_reg[5]/P0001  ;
  input \u0_slt2_r_reg[6]/P0001  ;
  input \u0_slt2_r_reg[7]/P0001  ;
  input \u0_slt2_r_reg[8]/P0001  ;
  input \u0_slt2_r_reg[9]/P0001  ;
  input \u0_slt3_r_reg[0]/P0001  ;
  input \u0_slt3_r_reg[10]/P0001  ;
  input \u0_slt3_r_reg[11]/P0001  ;
  input \u0_slt3_r_reg[12]/P0001  ;
  input \u0_slt3_r_reg[13]/P0001  ;
  input \u0_slt3_r_reg[14]/P0001  ;
  input \u0_slt3_r_reg[15]/P0001  ;
  input \u0_slt3_r_reg[16]/P0001  ;
  input \u0_slt3_r_reg[17]/P0001  ;
  input \u0_slt3_r_reg[18]/P0001  ;
  input \u0_slt3_r_reg[19]/P0001  ;
  input \u0_slt3_r_reg[1]/P0001  ;
  input \u0_slt3_r_reg[2]/P0001  ;
  input \u0_slt3_r_reg[3]/P0001  ;
  input \u0_slt3_r_reg[4]/P0001  ;
  input \u0_slt3_r_reg[5]/P0001  ;
  input \u0_slt3_r_reg[6]/P0001  ;
  input \u0_slt3_r_reg[7]/P0001  ;
  input \u0_slt3_r_reg[8]/P0001  ;
  input \u0_slt3_r_reg[9]/P0001  ;
  input \u0_slt4_r_reg[0]/P0001  ;
  input \u0_slt4_r_reg[10]/P0001  ;
  input \u0_slt4_r_reg[11]/P0001  ;
  input \u0_slt4_r_reg[12]/P0001  ;
  input \u0_slt4_r_reg[13]/P0001  ;
  input \u0_slt4_r_reg[14]/P0001  ;
  input \u0_slt4_r_reg[15]/P0001  ;
  input \u0_slt4_r_reg[16]/P0001  ;
  input \u0_slt4_r_reg[17]/P0001  ;
  input \u0_slt4_r_reg[18]/P0001  ;
  input \u0_slt4_r_reg[19]/P0001  ;
  input \u0_slt4_r_reg[1]/P0001  ;
  input \u0_slt4_r_reg[2]/P0001  ;
  input \u0_slt4_r_reg[3]/P0001  ;
  input \u0_slt4_r_reg[4]/P0001  ;
  input \u0_slt4_r_reg[5]/P0001  ;
  input \u0_slt4_r_reg[6]/P0001  ;
  input \u0_slt4_r_reg[7]/P0001  ;
  input \u0_slt4_r_reg[8]/P0001  ;
  input \u0_slt4_r_reg[9]/P0001  ;
  input \u0_slt5_r_reg[0]/P0001  ;
  input \u0_slt5_r_reg[10]/P0001  ;
  input \u0_slt5_r_reg[11]/P0001  ;
  input \u0_slt5_r_reg[12]/P0001  ;
  input \u0_slt5_r_reg[13]/P0001  ;
  input \u0_slt5_r_reg[14]/P0001  ;
  input \u0_slt5_r_reg[15]/P0001  ;
  input \u0_slt5_r_reg[16]/P0001  ;
  input \u0_slt5_r_reg[17]/P0001  ;
  input \u0_slt5_r_reg[18]/P0001  ;
  input \u0_slt5_r_reg[19]/P0001  ;
  input \u0_slt5_r_reg[1]/P0001  ;
  input \u0_slt5_r_reg[2]/P0001  ;
  input \u0_slt5_r_reg[3]/P0001  ;
  input \u0_slt5_r_reg[4]/P0001  ;
  input \u0_slt5_r_reg[5]/P0001  ;
  input \u0_slt5_r_reg[6]/P0001  ;
  input \u0_slt5_r_reg[7]/P0001  ;
  input \u0_slt5_r_reg[8]/P0001  ;
  input \u0_slt5_r_reg[9]/P0001  ;
  input \u0_slt6_r_reg[0]/P0001  ;
  input \u0_slt6_r_reg[10]/P0001  ;
  input \u0_slt6_r_reg[11]/P0001  ;
  input \u0_slt6_r_reg[12]/P0001  ;
  input \u0_slt6_r_reg[13]/P0001  ;
  input \u0_slt6_r_reg[14]/P0001  ;
  input \u0_slt6_r_reg[15]/P0001  ;
  input \u0_slt6_r_reg[16]/P0001  ;
  input \u0_slt6_r_reg[17]/P0001  ;
  input \u0_slt6_r_reg[18]/P0001  ;
  input \u0_slt6_r_reg[19]/P0001  ;
  input \u0_slt6_r_reg[1]/P0001  ;
  input \u0_slt6_r_reg[2]/P0001  ;
  input \u0_slt6_r_reg[3]/P0001  ;
  input \u0_slt6_r_reg[4]/P0001  ;
  input \u0_slt6_r_reg[5]/P0001  ;
  input \u0_slt6_r_reg[6]/P0001  ;
  input \u0_slt6_r_reg[7]/P0001  ;
  input \u0_slt6_r_reg[8]/P0001  ;
  input \u0_slt6_r_reg[9]/P0001  ;
  input \u0_slt7_r_reg[0]/P0001  ;
  input \u0_slt7_r_reg[10]/P0001  ;
  input \u0_slt7_r_reg[11]/P0001  ;
  input \u0_slt7_r_reg[12]/P0001  ;
  input \u0_slt7_r_reg[13]/P0001  ;
  input \u0_slt7_r_reg[14]/P0001  ;
  input \u0_slt7_r_reg[15]/P0001  ;
  input \u0_slt7_r_reg[16]/P0001  ;
  input \u0_slt7_r_reg[17]/P0001  ;
  input \u0_slt7_r_reg[18]/P0001  ;
  input \u0_slt7_r_reg[19]/P0001  ;
  input \u0_slt7_r_reg[1]/P0001  ;
  input \u0_slt7_r_reg[2]/P0001  ;
  input \u0_slt7_r_reg[3]/P0001  ;
  input \u0_slt7_r_reg[4]/P0001  ;
  input \u0_slt7_r_reg[5]/P0001  ;
  input \u0_slt7_r_reg[6]/P0001  ;
  input \u0_slt7_r_reg[7]/P0001  ;
  input \u0_slt7_r_reg[8]/P0001  ;
  input \u0_slt7_r_reg[9]/P0001  ;
  input \u0_slt8_r_reg[0]/P0001  ;
  input \u0_slt8_r_reg[10]/P0001  ;
  input \u0_slt8_r_reg[11]/P0001  ;
  input \u0_slt8_r_reg[12]/P0001  ;
  input \u0_slt8_r_reg[13]/P0001  ;
  input \u0_slt8_r_reg[14]/P0001  ;
  input \u0_slt8_r_reg[15]/P0001  ;
  input \u0_slt8_r_reg[16]/P0001  ;
  input \u0_slt8_r_reg[17]/P0001  ;
  input \u0_slt8_r_reg[18]/P0001  ;
  input \u0_slt8_r_reg[19]/P0001  ;
  input \u0_slt8_r_reg[1]/P0001  ;
  input \u0_slt8_r_reg[2]/P0001  ;
  input \u0_slt8_r_reg[3]/P0001  ;
  input \u0_slt8_r_reg[4]/P0001  ;
  input \u0_slt8_r_reg[5]/P0001  ;
  input \u0_slt8_r_reg[6]/P0001  ;
  input \u0_slt8_r_reg[7]/P0001  ;
  input \u0_slt8_r_reg[8]/P0001  ;
  input \u0_slt8_r_reg[9]/P0001  ;
  input \u0_slt9_r_reg[0]/P0001  ;
  input \u0_slt9_r_reg[10]/P0001  ;
  input \u0_slt9_r_reg[11]/P0001  ;
  input \u0_slt9_r_reg[12]/P0001  ;
  input \u0_slt9_r_reg[13]/P0001  ;
  input \u0_slt9_r_reg[14]/P0001  ;
  input \u0_slt9_r_reg[15]/P0001  ;
  input \u0_slt9_r_reg[16]/P0001  ;
  input \u0_slt9_r_reg[17]/P0001  ;
  input \u0_slt9_r_reg[18]/P0001  ;
  input \u0_slt9_r_reg[19]/P0001  ;
  input \u0_slt9_r_reg[1]/P0001  ;
  input \u0_slt9_r_reg[2]/P0001  ;
  input \u0_slt9_r_reg[3]/P0001  ;
  input \u0_slt9_r_reg[4]/P0001  ;
  input \u0_slt9_r_reg[5]/P0001  ;
  input \u0_slt9_r_reg[6]/P0001  ;
  input \u0_slt9_r_reg[7]/P0001  ;
  input \u0_slt9_r_reg[8]/P0001  ;
  input \u0_slt9_r_reg[9]/P0001  ;
  input \u10_din_tmp1_reg[0]/P0001  ;
  input \u10_din_tmp1_reg[10]/P0001  ;
  input \u10_din_tmp1_reg[11]/P0001  ;
  input \u10_din_tmp1_reg[12]/P0001  ;
  input \u10_din_tmp1_reg[13]/P0001  ;
  input \u10_din_tmp1_reg[14]/P0001  ;
  input \u10_din_tmp1_reg[15]/P0001  ;
  input \u10_din_tmp1_reg[1]/P0001  ;
  input \u10_din_tmp1_reg[2]/P0001  ;
  input \u10_din_tmp1_reg[3]/P0001  ;
  input \u10_din_tmp1_reg[4]/P0001  ;
  input \u10_din_tmp1_reg[5]/P0001  ;
  input \u10_din_tmp1_reg[6]/P0001  ;
  input \u10_din_tmp1_reg[7]/P0001  ;
  input \u10_din_tmp1_reg[8]/P0001  ;
  input \u10_din_tmp1_reg[9]/P0001  ;
  input \u10_dout_reg[0]/P0001  ;
  input \u10_dout_reg[10]/P0001  ;
  input \u10_dout_reg[11]/P0001  ;
  input \u10_dout_reg[12]/P0001  ;
  input \u10_dout_reg[13]/P0001  ;
  input \u10_dout_reg[14]/P0001  ;
  input \u10_dout_reg[15]/P0001  ;
  input \u10_dout_reg[16]/P0001  ;
  input \u10_dout_reg[17]/P0001  ;
  input \u10_dout_reg[18]/P0001  ;
  input \u10_dout_reg[19]/P0001  ;
  input \u10_dout_reg[1]/P0001  ;
  input \u10_dout_reg[20]/P0001  ;
  input \u10_dout_reg[21]/P0001  ;
  input \u10_dout_reg[22]/P0001  ;
  input \u10_dout_reg[23]/P0001  ;
  input \u10_dout_reg[24]/P0001  ;
  input \u10_dout_reg[25]/P0001  ;
  input \u10_dout_reg[26]/P0001  ;
  input \u10_dout_reg[27]/P0001  ;
  input \u10_dout_reg[28]/P0001  ;
  input \u10_dout_reg[29]/P0001  ;
  input \u10_dout_reg[2]/P0001  ;
  input \u10_dout_reg[30]/P0001  ;
  input \u10_dout_reg[31]/P0001  ;
  input \u10_dout_reg[3]/P0001  ;
  input \u10_dout_reg[4]/P0001  ;
  input \u10_dout_reg[5]/P0001  ;
  input \u10_dout_reg[6]/P0001  ;
  input \u10_dout_reg[7]/P0001  ;
  input \u10_dout_reg[8]/P0001  ;
  input \u10_dout_reg[9]/P0001  ;
  input \u10_empty_reg/P0001  ;
  input \u10_full_reg/NET0131  ;
  input \u10_mem_reg[0][0]/P0001  ;
  input \u10_mem_reg[0][10]/P0001  ;
  input \u10_mem_reg[0][11]/P0001  ;
  input \u10_mem_reg[0][12]/P0001  ;
  input \u10_mem_reg[0][13]/P0001  ;
  input \u10_mem_reg[0][14]/P0001  ;
  input \u10_mem_reg[0][15]/P0001  ;
  input \u10_mem_reg[0][16]/P0001  ;
  input \u10_mem_reg[0][17]/P0001  ;
  input \u10_mem_reg[0][18]/P0001  ;
  input \u10_mem_reg[0][19]/P0001  ;
  input \u10_mem_reg[0][1]/P0001  ;
  input \u10_mem_reg[0][20]/P0001  ;
  input \u10_mem_reg[0][21]/P0001  ;
  input \u10_mem_reg[0][22]/P0001  ;
  input \u10_mem_reg[0][23]/P0001  ;
  input \u10_mem_reg[0][24]/P0001  ;
  input \u10_mem_reg[0][25]/P0001  ;
  input \u10_mem_reg[0][26]/P0001  ;
  input \u10_mem_reg[0][27]/P0001  ;
  input \u10_mem_reg[0][28]/P0001  ;
  input \u10_mem_reg[0][29]/P0001  ;
  input \u10_mem_reg[0][2]/P0001  ;
  input \u10_mem_reg[0][30]/P0001  ;
  input \u10_mem_reg[0][31]/P0001  ;
  input \u10_mem_reg[0][3]/P0001  ;
  input \u10_mem_reg[0][4]/P0001  ;
  input \u10_mem_reg[0][5]/P0001  ;
  input \u10_mem_reg[0][6]/P0001  ;
  input \u10_mem_reg[0][7]/P0001  ;
  input \u10_mem_reg[0][8]/P0001  ;
  input \u10_mem_reg[0][9]/P0001  ;
  input \u10_mem_reg[1][0]/P0001  ;
  input \u10_mem_reg[1][10]/P0001  ;
  input \u10_mem_reg[1][11]/P0001  ;
  input \u10_mem_reg[1][12]/P0001  ;
  input \u10_mem_reg[1][13]/P0001  ;
  input \u10_mem_reg[1][14]/P0001  ;
  input \u10_mem_reg[1][15]/P0001  ;
  input \u10_mem_reg[1][16]/P0001  ;
  input \u10_mem_reg[1][17]/P0001  ;
  input \u10_mem_reg[1][18]/P0001  ;
  input \u10_mem_reg[1][19]/P0001  ;
  input \u10_mem_reg[1][1]/P0001  ;
  input \u10_mem_reg[1][20]/P0001  ;
  input \u10_mem_reg[1][21]/P0001  ;
  input \u10_mem_reg[1][22]/P0001  ;
  input \u10_mem_reg[1][23]/P0001  ;
  input \u10_mem_reg[1][24]/P0001  ;
  input \u10_mem_reg[1][25]/P0001  ;
  input \u10_mem_reg[1][26]/P0001  ;
  input \u10_mem_reg[1][27]/P0001  ;
  input \u10_mem_reg[1][28]/P0001  ;
  input \u10_mem_reg[1][29]/P0001  ;
  input \u10_mem_reg[1][2]/P0001  ;
  input \u10_mem_reg[1][30]/P0001  ;
  input \u10_mem_reg[1][31]/P0001  ;
  input \u10_mem_reg[1][3]/P0001  ;
  input \u10_mem_reg[1][4]/P0001  ;
  input \u10_mem_reg[1][5]/P0001  ;
  input \u10_mem_reg[1][6]/P0001  ;
  input \u10_mem_reg[1][7]/P0001  ;
  input \u10_mem_reg[1][8]/P0001  ;
  input \u10_mem_reg[1][9]/P0001  ;
  input \u10_mem_reg[2][0]/P0001  ;
  input \u10_mem_reg[2][10]/P0001  ;
  input \u10_mem_reg[2][11]/P0001  ;
  input \u10_mem_reg[2][12]/P0001  ;
  input \u10_mem_reg[2][13]/P0001  ;
  input \u10_mem_reg[2][14]/P0001  ;
  input \u10_mem_reg[2][15]/P0001  ;
  input \u10_mem_reg[2][16]/P0001  ;
  input \u10_mem_reg[2][17]/P0001  ;
  input \u10_mem_reg[2][18]/P0001  ;
  input \u10_mem_reg[2][19]/P0001  ;
  input \u10_mem_reg[2][1]/P0001  ;
  input \u10_mem_reg[2][20]/P0001  ;
  input \u10_mem_reg[2][21]/P0001  ;
  input \u10_mem_reg[2][22]/P0001  ;
  input \u10_mem_reg[2][23]/P0001  ;
  input \u10_mem_reg[2][24]/P0001  ;
  input \u10_mem_reg[2][25]/P0001  ;
  input \u10_mem_reg[2][26]/P0001  ;
  input \u10_mem_reg[2][27]/P0001  ;
  input \u10_mem_reg[2][28]/P0001  ;
  input \u10_mem_reg[2][29]/P0001  ;
  input \u10_mem_reg[2][2]/P0001  ;
  input \u10_mem_reg[2][30]/P0001  ;
  input \u10_mem_reg[2][31]/P0001  ;
  input \u10_mem_reg[2][3]/P0001  ;
  input \u10_mem_reg[2][4]/P0001  ;
  input \u10_mem_reg[2][5]/P0001  ;
  input \u10_mem_reg[2][6]/P0001  ;
  input \u10_mem_reg[2][7]/P0001  ;
  input \u10_mem_reg[2][8]/P0001  ;
  input \u10_mem_reg[2][9]/P0001  ;
  input \u10_mem_reg[3][0]/P0001  ;
  input \u10_mem_reg[3][10]/P0001  ;
  input \u10_mem_reg[3][11]/P0001  ;
  input \u10_mem_reg[3][12]/P0001  ;
  input \u10_mem_reg[3][13]/P0001  ;
  input \u10_mem_reg[3][14]/P0001  ;
  input \u10_mem_reg[3][15]/P0001  ;
  input \u10_mem_reg[3][16]/P0001  ;
  input \u10_mem_reg[3][17]/P0001  ;
  input \u10_mem_reg[3][18]/P0001  ;
  input \u10_mem_reg[3][19]/P0001  ;
  input \u10_mem_reg[3][1]/P0001  ;
  input \u10_mem_reg[3][20]/P0001  ;
  input \u10_mem_reg[3][21]/P0001  ;
  input \u10_mem_reg[3][22]/P0001  ;
  input \u10_mem_reg[3][23]/P0001  ;
  input \u10_mem_reg[3][24]/P0001  ;
  input \u10_mem_reg[3][25]/P0001  ;
  input \u10_mem_reg[3][26]/P0001  ;
  input \u10_mem_reg[3][27]/P0001  ;
  input \u10_mem_reg[3][28]/P0001  ;
  input \u10_mem_reg[3][29]/P0001  ;
  input \u10_mem_reg[3][2]/P0001  ;
  input \u10_mem_reg[3][30]/P0001  ;
  input \u10_mem_reg[3][31]/P0001  ;
  input \u10_mem_reg[3][3]/P0001  ;
  input \u10_mem_reg[3][4]/P0001  ;
  input \u10_mem_reg[3][5]/P0001  ;
  input \u10_mem_reg[3][6]/P0001  ;
  input \u10_mem_reg[3][7]/P0001  ;
  input \u10_mem_reg[3][8]/P0001  ;
  input \u10_mem_reg[3][9]/P0001  ;
  input \u10_rp_reg[0]/P0001  ;
  input \u10_rp_reg[1]/P0001  ;
  input \u10_rp_reg[2]/P0001  ;
  input \u10_status_reg[0]/P0001  ;
  input \u10_status_reg[1]/P0001  ;
  input \u10_wp_reg[0]/NET0131  ;
  input \u10_wp_reg[1]/P0001  ;
  input \u10_wp_reg[2]/P0001  ;
  input \u10_wp_reg[3]/P0001  ;
  input \u11_din_tmp1_reg[0]/P0001  ;
  input \u11_din_tmp1_reg[10]/P0001  ;
  input \u11_din_tmp1_reg[11]/P0001  ;
  input \u11_din_tmp1_reg[12]/P0001  ;
  input \u11_din_tmp1_reg[13]/P0001  ;
  input \u11_din_tmp1_reg[14]/P0001  ;
  input \u11_din_tmp1_reg[15]/P0001  ;
  input \u11_din_tmp1_reg[1]/P0001  ;
  input \u11_din_tmp1_reg[2]/P0001  ;
  input \u11_din_tmp1_reg[3]/P0001  ;
  input \u11_din_tmp1_reg[4]/P0001  ;
  input \u11_din_tmp1_reg[5]/P0001  ;
  input \u11_din_tmp1_reg[6]/P0001  ;
  input \u11_din_tmp1_reg[7]/P0001  ;
  input \u11_din_tmp1_reg[8]/P0001  ;
  input \u11_din_tmp1_reg[9]/P0001  ;
  input \u11_dout_reg[0]/P0001  ;
  input \u11_dout_reg[10]/P0001  ;
  input \u11_dout_reg[11]/P0001  ;
  input \u11_dout_reg[12]/P0001  ;
  input \u11_dout_reg[13]/P0001  ;
  input \u11_dout_reg[14]/P0001  ;
  input \u11_dout_reg[15]/P0001  ;
  input \u11_dout_reg[16]/P0001  ;
  input \u11_dout_reg[17]/P0001  ;
  input \u11_dout_reg[18]/P0001  ;
  input \u11_dout_reg[19]/P0001  ;
  input \u11_dout_reg[1]/P0001  ;
  input \u11_dout_reg[20]/P0001  ;
  input \u11_dout_reg[21]/P0001  ;
  input \u11_dout_reg[22]/P0001  ;
  input \u11_dout_reg[23]/P0001  ;
  input \u11_dout_reg[24]/P0001  ;
  input \u11_dout_reg[25]/P0001  ;
  input \u11_dout_reg[26]/P0001  ;
  input \u11_dout_reg[27]/P0001  ;
  input \u11_dout_reg[28]/P0001  ;
  input \u11_dout_reg[29]/P0001  ;
  input \u11_dout_reg[2]/P0001  ;
  input \u11_dout_reg[30]/P0001  ;
  input \u11_dout_reg[31]/P0001  ;
  input \u11_dout_reg[3]/P0001  ;
  input \u11_dout_reg[4]/P0001  ;
  input \u11_dout_reg[5]/P0001  ;
  input \u11_dout_reg[6]/P0001  ;
  input \u11_dout_reg[7]/P0001  ;
  input \u11_dout_reg[8]/P0001  ;
  input \u11_dout_reg[9]/P0001  ;
  input \u11_empty_reg/P0001  ;
  input \u11_full_reg/NET0131  ;
  input \u11_mem_reg[0][0]/P0001  ;
  input \u11_mem_reg[0][10]/P0001  ;
  input \u11_mem_reg[0][11]/P0001  ;
  input \u11_mem_reg[0][12]/P0001  ;
  input \u11_mem_reg[0][13]/P0001  ;
  input \u11_mem_reg[0][14]/P0001  ;
  input \u11_mem_reg[0][15]/P0001  ;
  input \u11_mem_reg[0][16]/P0001  ;
  input \u11_mem_reg[0][17]/P0001  ;
  input \u11_mem_reg[0][18]/P0001  ;
  input \u11_mem_reg[0][19]/P0001  ;
  input \u11_mem_reg[0][1]/P0001  ;
  input \u11_mem_reg[0][20]/P0001  ;
  input \u11_mem_reg[0][21]/P0001  ;
  input \u11_mem_reg[0][22]/P0001  ;
  input \u11_mem_reg[0][23]/P0001  ;
  input \u11_mem_reg[0][24]/P0001  ;
  input \u11_mem_reg[0][25]/P0001  ;
  input \u11_mem_reg[0][26]/P0001  ;
  input \u11_mem_reg[0][27]/P0001  ;
  input \u11_mem_reg[0][28]/P0001  ;
  input \u11_mem_reg[0][29]/P0001  ;
  input \u11_mem_reg[0][2]/P0001  ;
  input \u11_mem_reg[0][30]/P0001  ;
  input \u11_mem_reg[0][31]/P0001  ;
  input \u11_mem_reg[0][3]/P0001  ;
  input \u11_mem_reg[0][4]/P0001  ;
  input \u11_mem_reg[0][5]/P0001  ;
  input \u11_mem_reg[0][6]/P0001  ;
  input \u11_mem_reg[0][7]/P0001  ;
  input \u11_mem_reg[0][8]/P0001  ;
  input \u11_mem_reg[0][9]/P0001  ;
  input \u11_mem_reg[1][0]/P0001  ;
  input \u11_mem_reg[1][10]/P0001  ;
  input \u11_mem_reg[1][11]/P0001  ;
  input \u11_mem_reg[1][12]/P0001  ;
  input \u11_mem_reg[1][13]/P0001  ;
  input \u11_mem_reg[1][14]/P0001  ;
  input \u11_mem_reg[1][15]/P0001  ;
  input \u11_mem_reg[1][16]/P0001  ;
  input \u11_mem_reg[1][17]/P0001  ;
  input \u11_mem_reg[1][18]/P0001  ;
  input \u11_mem_reg[1][19]/P0001  ;
  input \u11_mem_reg[1][1]/P0001  ;
  input \u11_mem_reg[1][20]/P0001  ;
  input \u11_mem_reg[1][21]/P0001  ;
  input \u11_mem_reg[1][22]/P0001  ;
  input \u11_mem_reg[1][23]/P0001  ;
  input \u11_mem_reg[1][24]/P0001  ;
  input \u11_mem_reg[1][25]/P0001  ;
  input \u11_mem_reg[1][26]/P0001  ;
  input \u11_mem_reg[1][27]/P0001  ;
  input \u11_mem_reg[1][28]/P0001  ;
  input \u11_mem_reg[1][29]/P0001  ;
  input \u11_mem_reg[1][2]/P0001  ;
  input \u11_mem_reg[1][30]/P0001  ;
  input \u11_mem_reg[1][31]/P0001  ;
  input \u11_mem_reg[1][3]/P0001  ;
  input \u11_mem_reg[1][4]/P0001  ;
  input \u11_mem_reg[1][5]/P0001  ;
  input \u11_mem_reg[1][6]/P0001  ;
  input \u11_mem_reg[1][7]/P0001  ;
  input \u11_mem_reg[1][8]/P0001  ;
  input \u11_mem_reg[1][9]/P0001  ;
  input \u11_mem_reg[2][0]/P0001  ;
  input \u11_mem_reg[2][10]/P0001  ;
  input \u11_mem_reg[2][11]/P0001  ;
  input \u11_mem_reg[2][12]/P0001  ;
  input \u11_mem_reg[2][13]/P0001  ;
  input \u11_mem_reg[2][14]/P0001  ;
  input \u11_mem_reg[2][15]/P0001  ;
  input \u11_mem_reg[2][16]/P0001  ;
  input \u11_mem_reg[2][17]/P0001  ;
  input \u11_mem_reg[2][18]/P0001  ;
  input \u11_mem_reg[2][19]/P0001  ;
  input \u11_mem_reg[2][1]/P0001  ;
  input \u11_mem_reg[2][20]/P0001  ;
  input \u11_mem_reg[2][21]/P0001  ;
  input \u11_mem_reg[2][22]/P0001  ;
  input \u11_mem_reg[2][23]/P0001  ;
  input \u11_mem_reg[2][24]/P0001  ;
  input \u11_mem_reg[2][25]/P0001  ;
  input \u11_mem_reg[2][26]/P0001  ;
  input \u11_mem_reg[2][27]/P0001  ;
  input \u11_mem_reg[2][28]/P0001  ;
  input \u11_mem_reg[2][29]/P0001  ;
  input \u11_mem_reg[2][2]/P0001  ;
  input \u11_mem_reg[2][30]/P0001  ;
  input \u11_mem_reg[2][31]/P0001  ;
  input \u11_mem_reg[2][3]/P0001  ;
  input \u11_mem_reg[2][4]/P0001  ;
  input \u11_mem_reg[2][5]/P0001  ;
  input \u11_mem_reg[2][6]/P0001  ;
  input \u11_mem_reg[2][7]/P0001  ;
  input \u11_mem_reg[2][8]/P0001  ;
  input \u11_mem_reg[2][9]/P0001  ;
  input \u11_mem_reg[3][0]/P0001  ;
  input \u11_mem_reg[3][10]/P0001  ;
  input \u11_mem_reg[3][11]/P0001  ;
  input \u11_mem_reg[3][12]/P0001  ;
  input \u11_mem_reg[3][13]/P0001  ;
  input \u11_mem_reg[3][14]/P0001  ;
  input \u11_mem_reg[3][15]/P0001  ;
  input \u11_mem_reg[3][16]/P0001  ;
  input \u11_mem_reg[3][17]/P0001  ;
  input \u11_mem_reg[3][18]/P0001  ;
  input \u11_mem_reg[3][19]/P0001  ;
  input \u11_mem_reg[3][1]/P0001  ;
  input \u11_mem_reg[3][20]/P0001  ;
  input \u11_mem_reg[3][21]/P0001  ;
  input \u11_mem_reg[3][22]/P0001  ;
  input \u11_mem_reg[3][23]/P0001  ;
  input \u11_mem_reg[3][24]/P0001  ;
  input \u11_mem_reg[3][25]/P0001  ;
  input \u11_mem_reg[3][26]/P0001  ;
  input \u11_mem_reg[3][27]/P0001  ;
  input \u11_mem_reg[3][28]/P0001  ;
  input \u11_mem_reg[3][29]/P0001  ;
  input \u11_mem_reg[3][2]/P0001  ;
  input \u11_mem_reg[3][30]/P0001  ;
  input \u11_mem_reg[3][31]/P0001  ;
  input \u11_mem_reg[3][3]/P0001  ;
  input \u11_mem_reg[3][4]/P0001  ;
  input \u11_mem_reg[3][5]/P0001  ;
  input \u11_mem_reg[3][6]/P0001  ;
  input \u11_mem_reg[3][7]/P0001  ;
  input \u11_mem_reg[3][8]/P0001  ;
  input \u11_mem_reg[3][9]/P0001  ;
  input \u11_rp_reg[0]/P0001  ;
  input \u11_rp_reg[1]/P0001  ;
  input \u11_rp_reg[2]/P0001  ;
  input \u11_status_reg[0]/P0001  ;
  input \u11_status_reg[1]/P0001  ;
  input \u11_wp_reg[0]/NET0131  ;
  input \u11_wp_reg[1]/P0001  ;
  input \u11_wp_reg[2]/P0001  ;
  input \u11_wp_reg[3]/P0001  ;
  input \u12_dout_reg[0]/P0001  ;
  input \u12_dout_reg[10]/P0001  ;
  input \u12_dout_reg[11]/P0001  ;
  input \u12_dout_reg[12]/P0001  ;
  input \u12_dout_reg[13]/P0001  ;
  input \u12_dout_reg[14]/P0001  ;
  input \u12_dout_reg[15]/P0001  ;
  input \u12_dout_reg[16]/P0001  ;
  input \u12_dout_reg[17]/P0001  ;
  input \u12_dout_reg[18]/P0001  ;
  input \u12_dout_reg[19]/P0001  ;
  input \u12_dout_reg[1]/P0001  ;
  input \u12_dout_reg[20]/P0001  ;
  input \u12_dout_reg[21]/P0001  ;
  input \u12_dout_reg[22]/P0001  ;
  input \u12_dout_reg[23]/P0001  ;
  input \u12_dout_reg[24]/P0001  ;
  input \u12_dout_reg[25]/P0001  ;
  input \u12_dout_reg[26]/P0001  ;
  input \u12_dout_reg[27]/P0001  ;
  input \u12_dout_reg[28]/P0001  ;
  input \u12_dout_reg[29]/P0001  ;
  input \u12_dout_reg[2]/P0001  ;
  input \u12_dout_reg[30]/P0001  ;
  input \u12_dout_reg[31]/P0001  ;
  input \u12_dout_reg[3]/P0001  ;
  input \u12_dout_reg[4]/P0001  ;
  input \u12_dout_reg[5]/P0001  ;
  input \u12_dout_reg[6]/P0001  ;
  input \u12_dout_reg[7]/P0001  ;
  input \u12_dout_reg[8]/P0001  ;
  input \u12_dout_reg[9]/P0001  ;
  input \u12_i3_re_reg/NET0131  ;
  input \u12_i4_re_reg/P0001  ;
  input \u12_i6_re_reg/NET0131  ;
  input \u12_o3_we_reg/P0001  ;
  input \u12_o4_we_reg/P0001  ;
  input \u12_o6_we_reg/P0001  ;
  input \u12_o7_we_reg/P0001  ;
  input \u12_o8_we_reg/P0001  ;
  input \u12_o9_we_reg/P0001  ;
  input \u12_re1_reg/P0001  ;
  input \u12_re2_reg/NET0131  ;
  input \u12_rf_we_reg/P0001  ;
  input \u12_we1_reg/P0001  ;
  input \u12_we2_reg/P0001  ;
  input \u13_ac97_rst_force_reg/P0001  ;
  input \u13_crac_dout_r_reg[0]/P0001  ;
  input \u13_crac_dout_r_reg[10]/P0001  ;
  input \u13_crac_dout_r_reg[11]/P0001  ;
  input \u13_crac_dout_r_reg[12]/P0001  ;
  input \u13_crac_dout_r_reg[13]/P0001  ;
  input \u13_crac_dout_r_reg[14]/P0001  ;
  input \u13_crac_dout_r_reg[15]/P0001  ;
  input \u13_crac_dout_r_reg[1]/P0001  ;
  input \u13_crac_dout_r_reg[2]/P0001  ;
  input \u13_crac_dout_r_reg[3]/P0001  ;
  input \u13_crac_dout_r_reg[4]/P0001  ;
  input \u13_crac_dout_r_reg[5]/P0001  ;
  input \u13_crac_dout_r_reg[6]/P0001  ;
  input \u13_crac_dout_r_reg[7]/P0001  ;
  input \u13_crac_dout_r_reg[8]/P0001  ;
  input \u13_crac_dout_r_reg[9]/P0001  ;
  input \u13_crac_r_reg[0]/NET0131  ;
  input \u13_crac_r_reg[1]/NET0131  ;
  input \u13_crac_r_reg[2]/NET0131  ;
  input \u13_crac_r_reg[3]/NET0131  ;
  input \u13_crac_r_reg[4]/NET0131  ;
  input \u13_crac_r_reg[5]/NET0131  ;
  input \u13_crac_r_reg[6]/NET0131  ;
  input \u13_crac_r_reg[7]/NET0131  ;
  input \u13_icc_r_reg[0]/NET0131  ;
  input \u13_icc_r_reg[10]/NET0131  ;
  input \u13_icc_r_reg[11]/NET0131  ;
  input \u13_icc_r_reg[12]/NET0131  ;
  input \u13_icc_r_reg[13]/NET0131  ;
  input \u13_icc_r_reg[14]/NET0131  ;
  input \u13_icc_r_reg[15]/NET0131  ;
  input \u13_icc_r_reg[16]/NET0131  ;
  input \u13_icc_r_reg[17]/NET0131  ;
  input \u13_icc_r_reg[18]/NET0131  ;
  input \u13_icc_r_reg[19]/NET0131  ;
  input \u13_icc_r_reg[1]/NET0131  ;
  input \u13_icc_r_reg[20]/NET0131  ;
  input \u13_icc_r_reg[21]/NET0131  ;
  input \u13_icc_r_reg[22]/NET0131  ;
  input \u13_icc_r_reg[23]/NET0131  ;
  input \u13_icc_r_reg[2]/NET0131  ;
  input \u13_icc_r_reg[3]/NET0131  ;
  input \u13_icc_r_reg[4]/NET0131  ;
  input \u13_icc_r_reg[5]/NET0131  ;
  input \u13_icc_r_reg[6]/NET0131  ;
  input \u13_icc_r_reg[7]/NET0131  ;
  input \u13_icc_r_reg[8]/NET0131  ;
  input \u13_icc_r_reg[9]/NET0131  ;
  input \u13_intm_r_reg[0]/NET0131  ;
  input \u13_intm_r_reg[10]/NET0131  ;
  input \u13_intm_r_reg[11]/NET0131  ;
  input \u13_intm_r_reg[12]/NET0131  ;
  input \u13_intm_r_reg[13]/NET0131  ;
  input \u13_intm_r_reg[14]/NET0131  ;
  input \u13_intm_r_reg[15]/NET0131  ;
  input \u13_intm_r_reg[16]/NET0131  ;
  input \u13_intm_r_reg[17]/NET0131  ;
  input \u13_intm_r_reg[18]/NET0131  ;
  input \u13_intm_r_reg[19]/NET0131  ;
  input \u13_intm_r_reg[1]/NET0131  ;
  input \u13_intm_r_reg[20]/NET0131  ;
  input \u13_intm_r_reg[21]/NET0131  ;
  input \u13_intm_r_reg[22]/NET0131  ;
  input \u13_intm_r_reg[23]/NET0131  ;
  input \u13_intm_r_reg[24]/NET0131  ;
  input \u13_intm_r_reg[25]/NET0131  ;
  input \u13_intm_r_reg[26]/NET0131  ;
  input \u13_intm_r_reg[27]/NET0131  ;
  input \u13_intm_r_reg[28]/NET0131  ;
  input \u13_intm_r_reg[2]/NET0131  ;
  input \u13_intm_r_reg[3]/NET0131  ;
  input \u13_intm_r_reg[4]/NET0131  ;
  input \u13_intm_r_reg[5]/NET0131  ;
  input \u13_intm_r_reg[6]/NET0131  ;
  input \u13_intm_r_reg[7]/NET0131  ;
  input \u13_intm_r_reg[8]/NET0131  ;
  input \u13_intm_r_reg[9]/NET0131  ;
  input \u13_ints_r_reg[0]/NET0131  ;
  input \u13_ints_r_reg[10]/NET0131  ;
  input \u13_ints_r_reg[11]/NET0131  ;
  input \u13_ints_r_reg[12]/NET0131  ;
  input \u13_ints_r_reg[13]/NET0131  ;
  input \u13_ints_r_reg[14]/NET0131  ;
  input \u13_ints_r_reg[15]/NET0131  ;
  input \u13_ints_r_reg[16]/NET0131  ;
  input \u13_ints_r_reg[17]/NET0131  ;
  input \u13_ints_r_reg[18]/NET0131  ;
  input \u13_ints_r_reg[19]/NET0131  ;
  input \u13_ints_r_reg[1]/NET0131  ;
  input \u13_ints_r_reg[20]/NET0131  ;
  input \u13_ints_r_reg[21]/NET0131  ;
  input \u13_ints_r_reg[22]/NET0131  ;
  input \u13_ints_r_reg[23]/NET0131  ;
  input \u13_ints_r_reg[24]/NET0131  ;
  input \u13_ints_r_reg[25]/NET0131  ;
  input \u13_ints_r_reg[26]/NET0131  ;
  input \u13_ints_r_reg[27]/NET0131  ;
  input \u13_ints_r_reg[28]/NET0131  ;
  input \u13_ints_r_reg[2]/NET0131  ;
  input \u13_ints_r_reg[3]/NET0131  ;
  input \u13_ints_r_reg[4]/NET0131  ;
  input \u13_ints_r_reg[5]/NET0131  ;
  input \u13_ints_r_reg[6]/NET0131  ;
  input \u13_ints_r_reg[7]/NET0131  ;
  input \u13_ints_r_reg[8]/NET0131  ;
  input \u13_ints_r_reg[9]/NET0131  ;
  input \u13_occ0_r_reg[0]/NET0131  ;
  input \u13_occ0_r_reg[10]/NET0131  ;
  input \u13_occ0_r_reg[11]/NET0131  ;
  input \u13_occ0_r_reg[12]/NET0131  ;
  input \u13_occ0_r_reg[13]/NET0131  ;
  input \u13_occ0_r_reg[14]/NET0131  ;
  input \u13_occ0_r_reg[15]/NET0131  ;
  input \u13_occ0_r_reg[16]/NET0131  ;
  input \u13_occ0_r_reg[17]/NET0131  ;
  input \u13_occ0_r_reg[18]/NET0131  ;
  input \u13_occ0_r_reg[19]/NET0131  ;
  input \u13_occ0_r_reg[1]/NET0131  ;
  input \u13_occ0_r_reg[20]/NET0131  ;
  input \u13_occ0_r_reg[21]/NET0131  ;
  input \u13_occ0_r_reg[22]/NET0131  ;
  input \u13_occ0_r_reg[23]/NET0131  ;
  input \u13_occ0_r_reg[24]/NET0131  ;
  input \u13_occ0_r_reg[25]/NET0131  ;
  input \u13_occ0_r_reg[26]/NET0131  ;
  input \u13_occ0_r_reg[27]/NET0131  ;
  input \u13_occ0_r_reg[28]/NET0131  ;
  input \u13_occ0_r_reg[29]/NET0131  ;
  input \u13_occ0_r_reg[2]/NET0131  ;
  input \u13_occ0_r_reg[30]/NET0131  ;
  input \u13_occ0_r_reg[31]/NET0131  ;
  input \u13_occ0_r_reg[3]/NET0131  ;
  input \u13_occ0_r_reg[4]/NET0131  ;
  input \u13_occ0_r_reg[5]/NET0131  ;
  input \u13_occ0_r_reg[6]/NET0131  ;
  input \u13_occ0_r_reg[7]/NET0131  ;
  input \u13_occ0_r_reg[8]/NET0131  ;
  input \u13_occ0_r_reg[9]/NET0131  ;
  input \u13_occ1_r_reg[0]/NET0131  ;
  input \u13_occ1_r_reg[10]/NET0131  ;
  input \u13_occ1_r_reg[11]/NET0131  ;
  input \u13_occ1_r_reg[12]/NET0131  ;
  input \u13_occ1_r_reg[13]/NET0131  ;
  input \u13_occ1_r_reg[14]/NET0131  ;
  input \u13_occ1_r_reg[15]/NET0131  ;
  input \u13_occ1_r_reg[1]/NET0131  ;
  input \u13_occ1_r_reg[2]/NET0131  ;
  input \u13_occ1_r_reg[3]/NET0131  ;
  input \u13_occ1_r_reg[4]/NET0131  ;
  input \u13_occ1_r_reg[5]/NET0131  ;
  input \u13_occ1_r_reg[6]/NET0131  ;
  input \u13_occ1_r_reg[7]/NET0131  ;
  input \u13_occ1_r_reg[8]/NET0131  ;
  input \u13_occ1_r_reg[9]/NET0131  ;
  input \u13_resume_req_reg/P0001  ;
  input \u14_crac_valid_r_reg/P0001  ;
  input \u14_crac_wr_r_reg/P0001  ;
  input \u14_u0_en_out_l2_reg/P0001  ;
  input \u14_u0_en_out_l_reg/NET0131  ;
  input \u14_u0_full_empty_r_reg/P0001  ;
  input \u14_u1_en_out_l2_reg/P0001  ;
  input \u14_u1_en_out_l_reg/NET0131  ;
  input \u14_u1_full_empty_r_reg/P0001  ;
  input \u14_u2_en_out_l2_reg/P0001  ;
  input \u14_u2_en_out_l_reg/NET0131  ;
  input \u14_u2_full_empty_r_reg/P0001  ;
  input \u14_u3_en_out_l2_reg/P0001  ;
  input \u14_u3_en_out_l_reg/NET0131  ;
  input \u14_u3_full_empty_r_reg/P0001  ;
  input \u14_u4_en_out_l2_reg/P0001  ;
  input \u14_u4_en_out_l_reg/NET0131  ;
  input \u14_u4_full_empty_r_reg/P0001  ;
  input \u14_u5_en_out_l2_reg/P0001  ;
  input \u14_u5_en_out_l_reg/NET0131  ;
  input \u14_u5_full_empty_r_reg/P0001  ;
  input \u14_u6_en_out_l2_reg/P0001  ;
  input \u14_u6_en_out_l_reg/NET0131  ;
  input \u14_u6_full_empty_r_reg/P0001  ;
  input \u14_u7_en_out_l2_reg/P0001  ;
  input \u14_u7_en_out_l_reg/NET0131  ;
  input \u14_u7_full_empty_r_reg/P0001  ;
  input \u14_u8_en_out_l2_reg/P0001  ;
  input \u14_u8_en_out_l_reg/NET0131  ;
  input \u14_u8_full_empty_r_reg/P0001  ;
  input \u15_crac_din_reg[0]/NET0131  ;
  input \u15_crac_din_reg[10]/NET0131  ;
  input \u15_crac_din_reg[11]/NET0131  ;
  input \u15_crac_din_reg[12]/NET0131  ;
  input \u15_crac_din_reg[13]/NET0131  ;
  input \u15_crac_din_reg[14]/NET0131  ;
  input \u15_crac_din_reg[15]/NET0131  ;
  input \u15_crac_din_reg[1]/NET0131  ;
  input \u15_crac_din_reg[2]/NET0131  ;
  input \u15_crac_din_reg[3]/NET0131  ;
  input \u15_crac_din_reg[4]/NET0131  ;
  input \u15_crac_din_reg[5]/NET0131  ;
  input \u15_crac_din_reg[6]/NET0131  ;
  input \u15_crac_din_reg[7]/NET0131  ;
  input \u15_crac_din_reg[8]/NET0131  ;
  input \u15_crac_din_reg[9]/NET0131  ;
  input \u15_crac_rd_done_reg/P0001  ;
  input \u15_crac_rd_reg/NET0131  ;
  input \u15_crac_we_r_reg/P0001  ;
  input \u15_crac_wr_reg/NET0131  ;
  input \u15_rdd1_reg/NET0131  ;
  input \u15_rdd2_reg/NET0131  ;
  input \u15_rdd3_reg/NET0131  ;
  input \u15_valid_r_reg/P0001  ;
  input \u16_u0_dma_req_r1_reg/P0001  ;
  input \u16_u1_dma_req_r1_reg/P0001  ;
  input \u16_u2_dma_req_r1_reg/P0001  ;
  input \u16_u3_dma_req_r1_reg/P0001  ;
  input \u16_u4_dma_req_r1_reg/P0001  ;
  input \u16_u5_dma_req_r1_reg/P0001  ;
  input \u16_u6_dma_req_r1_reg/P0001  ;
  input \u16_u7_dma_req_r1_reg/P0001  ;
  input \u16_u8_dma_req_r1_reg/P0001  ;
  input \u17_int_set_reg[0]/NET0131  ;
  input \u17_int_set_reg[1]/NET0131  ;
  input \u17_int_set_reg[2]/NET0131  ;
  input \u18_int_set_reg[0]/NET0131  ;
  input \u18_int_set_reg[1]/NET0131  ;
  input \u18_int_set_reg[2]/NET0131  ;
  input \u19_int_set_reg[0]/NET0131  ;
  input \u19_int_set_reg[1]/NET0131  ;
  input \u19_int_set_reg[2]/NET0131  ;
  input \u1_slt0_reg[11]/P0001  ;
  input \u1_slt0_reg[12]/P0001  ;
  input \u1_slt0_reg[15]/P0001  ;
  input \u1_slt0_reg[9]/P0001  ;
  input \u1_slt1_reg[10]/P0001  ;
  input \u1_slt1_reg[11]/P0001  ;
  input \u1_slt1_reg[5]/P0001  ;
  input \u1_slt1_reg[6]/P0001  ;
  input \u1_slt1_reg[7]/P0001  ;
  input \u1_slt1_reg[8]/P0001  ;
  input \u1_slt3_reg[0]/P0001  ;
  input \u1_slt3_reg[10]/P0001  ;
  input \u1_slt3_reg[11]/P0001  ;
  input \u1_slt3_reg[12]/P0001  ;
  input \u1_slt3_reg[13]/P0001  ;
  input \u1_slt3_reg[14]/P0001  ;
  input \u1_slt3_reg[15]/P0001  ;
  input \u1_slt3_reg[16]/P0001  ;
  input \u1_slt3_reg[17]/P0001  ;
  input \u1_slt3_reg[18]/P0001  ;
  input \u1_slt3_reg[19]/P0001  ;
  input \u1_slt3_reg[1]/P0001  ;
  input \u1_slt3_reg[2]/P0001  ;
  input \u1_slt3_reg[3]/P0001  ;
  input \u1_slt3_reg[4]/P0001  ;
  input \u1_slt3_reg[5]/P0001  ;
  input \u1_slt3_reg[6]/P0001  ;
  input \u1_slt3_reg[7]/P0001  ;
  input \u1_slt3_reg[8]/P0001  ;
  input \u1_slt3_reg[9]/P0001  ;
  input \u1_slt4_reg[0]/P0001  ;
  input \u1_slt4_reg[10]/P0001  ;
  input \u1_slt4_reg[11]/P0001  ;
  input \u1_slt4_reg[12]/P0001  ;
  input \u1_slt4_reg[13]/P0001  ;
  input \u1_slt4_reg[14]/P0001  ;
  input \u1_slt4_reg[15]/P0001  ;
  input \u1_slt4_reg[16]/P0001  ;
  input \u1_slt4_reg[17]/P0001  ;
  input \u1_slt4_reg[18]/P0001  ;
  input \u1_slt4_reg[19]/P0001  ;
  input \u1_slt4_reg[1]/P0001  ;
  input \u1_slt4_reg[2]/P0001  ;
  input \u1_slt4_reg[3]/P0001  ;
  input \u1_slt4_reg[4]/P0001  ;
  input \u1_slt4_reg[5]/P0001  ;
  input \u1_slt4_reg[6]/P0001  ;
  input \u1_slt4_reg[7]/P0001  ;
  input \u1_slt4_reg[8]/P0001  ;
  input \u1_slt4_reg[9]/P0001  ;
  input \u1_slt6_reg[0]/P0001  ;
  input \u1_slt6_reg[10]/P0001  ;
  input \u1_slt6_reg[11]/P0001  ;
  input \u1_slt6_reg[12]/P0001  ;
  input \u1_slt6_reg[13]/P0001  ;
  input \u1_slt6_reg[14]/P0001  ;
  input \u1_slt6_reg[15]/P0001  ;
  input \u1_slt6_reg[16]/P0001  ;
  input \u1_slt6_reg[17]/P0001  ;
  input \u1_slt6_reg[18]/P0001  ;
  input \u1_slt6_reg[19]/P0001  ;
  input \u1_slt6_reg[1]/P0001  ;
  input \u1_slt6_reg[2]/P0001  ;
  input \u1_slt6_reg[3]/P0001  ;
  input \u1_slt6_reg[4]/P0001  ;
  input \u1_slt6_reg[5]/P0001  ;
  input \u1_slt6_reg[6]/P0001  ;
  input \u1_slt6_reg[7]/P0001  ;
  input \u1_slt6_reg[8]/P0001  ;
  input \u1_slt6_reg[9]/P0001  ;
  input \u1_sr_reg[10]/P0001  ;
  input \u1_sr_reg[11]/P0001  ;
  input \u1_sr_reg[12]/P0001  ;
  input \u1_sr_reg[15]/P0001  ;
  input \u1_sr_reg[5]/P0001  ;
  input \u1_sr_reg[6]/P0001  ;
  input \u1_sr_reg[7]/P0001  ;
  input \u1_sr_reg[8]/P0001  ;
  input \u1_sr_reg[9]/P0001  ;
  input \u20_int_set_reg[0]/NET0131  ;
  input \u20_int_set_reg[1]/NET0131  ;
  input \u20_int_set_reg[2]/NET0131  ;
  input \u21_int_set_reg[0]/NET0131  ;
  input \u21_int_set_reg[1]/NET0131  ;
  input \u21_int_set_reg[2]/NET0131  ;
  input \u22_int_set_reg[0]/NET0131  ;
  input \u22_int_set_reg[1]/NET0131  ;
  input \u22_int_set_reg[2]/NET0131  ;
  input \u23_int_set_reg[0]/NET0131  ;
  input \u23_int_set_reg[1]/NET0131  ;
  input \u23_int_set_reg[2]/NET0131  ;
  input \u24_int_set_reg[0]/NET0131  ;
  input \u24_int_set_reg[1]/NET0131  ;
  input \u24_int_set_reg[2]/NET0131  ;
  input \u25_int_set_reg[0]/NET0131  ;
  input \u25_int_set_reg[1]/NET0131  ;
  input \u25_int_set_reg[2]/NET0131  ;
  input \u26_cnt_reg[0]/NET0131  ;
  input \u26_cnt_reg[1]/NET0131  ;
  input \u26_cnt_reg[2]/NET0131  ;
  input \u26_ps_cnt_reg[0]/NET0131  ;
  input \u26_ps_cnt_reg[1]/NET0131  ;
  input \u26_ps_cnt_reg[2]/NET0131  ;
  input \u26_ps_cnt_reg[3]/NET0131  ;
  input \u26_ps_cnt_reg[4]/NET0131  ;
  input \u26_ps_cnt_reg[5]/NET0131  ;
  input \u2_bit_clk_e_reg/P0001  ;
  input \u2_bit_clk_r1_reg/P0001  ;
  input \u2_bit_clk_r_reg/P0001  ;
  input \u2_cnt_reg[0]/NET0131  ;
  input \u2_cnt_reg[1]/NET0131  ;
  input \u2_cnt_reg[2]/NET0131  ;
  input \u2_cnt_reg[3]/NET0131  ;
  input \u2_cnt_reg[4]/NET0131  ;
  input \u2_cnt_reg[5]/NET0131  ;
  input \u2_cnt_reg[6]/NET0131  ;
  input \u2_cnt_reg[7]/NET0131  ;
  input \u2_ld_reg/P0001  ;
  input \u2_out_le_reg[0]/P0001  ;
  input \u2_out_le_reg[1]/P0001  ;
  input \u2_res_cnt_reg[0]/P0001  ;
  input \u2_res_cnt_reg[1]/P0001  ;
  input \u2_res_cnt_reg[2]/P0001  ;
  input \u2_res_cnt_reg[3]/P0001  ;
  input \u2_sync_beat_reg/P0001  ;
  input \u2_sync_resume_reg/NET0131  ;
  input \u2_to_cnt_reg[0]/NET0131  ;
  input \u2_to_cnt_reg[1]/NET0131  ;
  input \u2_to_cnt_reg[2]/NET0131  ;
  input \u2_to_cnt_reg[3]/NET0131  ;
  input \u2_to_cnt_reg[4]/NET0131  ;
  input \u2_to_cnt_reg[5]/NET0131  ;
  input \u3_dout_reg[0]/P0001  ;
  input \u3_dout_reg[10]/P0001  ;
  input \u3_dout_reg[11]/P0001  ;
  input \u3_dout_reg[12]/P0001  ;
  input \u3_dout_reg[13]/P0001  ;
  input \u3_dout_reg[14]/P0001  ;
  input \u3_dout_reg[15]/P0001  ;
  input \u3_dout_reg[16]/P0001  ;
  input \u3_dout_reg[17]/P0001  ;
  input \u3_dout_reg[18]/P0001  ;
  input \u3_dout_reg[19]/P0001  ;
  input \u3_dout_reg[1]/P0001  ;
  input \u3_dout_reg[2]/P0001  ;
  input \u3_dout_reg[3]/P0001  ;
  input \u3_dout_reg[4]/P0001  ;
  input \u3_dout_reg[5]/P0001  ;
  input \u3_dout_reg[6]/P0001  ;
  input \u3_dout_reg[7]/P0001  ;
  input \u3_dout_reg[8]/P0001  ;
  input \u3_dout_reg[9]/P0001  ;
  input \u3_empty_reg/NET0131  ;
  input \u3_mem_reg[0][0]/NET0131  ;
  input \u3_mem_reg[0][10]/NET0131  ;
  input \u3_mem_reg[0][11]/NET0131  ;
  input \u3_mem_reg[0][12]/NET0131  ;
  input \u3_mem_reg[0][13]/NET0131  ;
  input \u3_mem_reg[0][14]/NET0131  ;
  input \u3_mem_reg[0][15]/NET0131  ;
  input \u3_mem_reg[0][16]/NET0131  ;
  input \u3_mem_reg[0][17]/NET0131  ;
  input \u3_mem_reg[0][18]/NET0131  ;
  input \u3_mem_reg[0][19]/NET0131  ;
  input \u3_mem_reg[0][1]/NET0131  ;
  input \u3_mem_reg[0][20]/NET0131  ;
  input \u3_mem_reg[0][21]/NET0131  ;
  input \u3_mem_reg[0][22]/NET0131  ;
  input \u3_mem_reg[0][23]/NET0131  ;
  input \u3_mem_reg[0][24]/NET0131  ;
  input \u3_mem_reg[0][25]/NET0131  ;
  input \u3_mem_reg[0][26]/NET0131  ;
  input \u3_mem_reg[0][27]/NET0131  ;
  input \u3_mem_reg[0][28]/NET0131  ;
  input \u3_mem_reg[0][29]/NET0131  ;
  input \u3_mem_reg[0][2]/NET0131  ;
  input \u3_mem_reg[0][30]/NET0131  ;
  input \u3_mem_reg[0][31]/NET0131  ;
  input \u3_mem_reg[0][3]/NET0131  ;
  input \u3_mem_reg[0][4]/NET0131  ;
  input \u3_mem_reg[0][5]/NET0131  ;
  input \u3_mem_reg[0][6]/NET0131  ;
  input \u3_mem_reg[0][7]/NET0131  ;
  input \u3_mem_reg[0][8]/NET0131  ;
  input \u3_mem_reg[0][9]/NET0131  ;
  input \u3_mem_reg[1][0]/NET0131  ;
  input \u3_mem_reg[1][10]/NET0131  ;
  input \u3_mem_reg[1][11]/NET0131  ;
  input \u3_mem_reg[1][12]/NET0131  ;
  input \u3_mem_reg[1][13]/NET0131  ;
  input \u3_mem_reg[1][14]/NET0131  ;
  input \u3_mem_reg[1][15]/NET0131  ;
  input \u3_mem_reg[1][16]/NET0131  ;
  input \u3_mem_reg[1][17]/NET0131  ;
  input \u3_mem_reg[1][18]/NET0131  ;
  input \u3_mem_reg[1][19]/NET0131  ;
  input \u3_mem_reg[1][1]/NET0131  ;
  input \u3_mem_reg[1][20]/NET0131  ;
  input \u3_mem_reg[1][21]/NET0131  ;
  input \u3_mem_reg[1][22]/NET0131  ;
  input \u3_mem_reg[1][23]/NET0131  ;
  input \u3_mem_reg[1][24]/NET0131  ;
  input \u3_mem_reg[1][25]/NET0131  ;
  input \u3_mem_reg[1][26]/NET0131  ;
  input \u3_mem_reg[1][27]/NET0131  ;
  input \u3_mem_reg[1][28]/NET0131  ;
  input \u3_mem_reg[1][29]/NET0131  ;
  input \u3_mem_reg[1][2]/NET0131  ;
  input \u3_mem_reg[1][30]/NET0131  ;
  input \u3_mem_reg[1][31]/NET0131  ;
  input \u3_mem_reg[1][3]/NET0131  ;
  input \u3_mem_reg[1][4]/NET0131  ;
  input \u3_mem_reg[1][5]/NET0131  ;
  input \u3_mem_reg[1][6]/NET0131  ;
  input \u3_mem_reg[1][7]/NET0131  ;
  input \u3_mem_reg[1][8]/NET0131  ;
  input \u3_mem_reg[1][9]/NET0131  ;
  input \u3_mem_reg[2][0]/NET0131  ;
  input \u3_mem_reg[2][10]/NET0131  ;
  input \u3_mem_reg[2][11]/NET0131  ;
  input \u3_mem_reg[2][12]/NET0131  ;
  input \u3_mem_reg[2][13]/NET0131  ;
  input \u3_mem_reg[2][14]/NET0131  ;
  input \u3_mem_reg[2][15]/NET0131  ;
  input \u3_mem_reg[2][16]/NET0131  ;
  input \u3_mem_reg[2][17]/NET0131  ;
  input \u3_mem_reg[2][18]/NET0131  ;
  input \u3_mem_reg[2][19]/NET0131  ;
  input \u3_mem_reg[2][1]/NET0131  ;
  input \u3_mem_reg[2][20]/NET0131  ;
  input \u3_mem_reg[2][21]/NET0131  ;
  input \u3_mem_reg[2][22]/NET0131  ;
  input \u3_mem_reg[2][23]/NET0131  ;
  input \u3_mem_reg[2][24]/NET0131  ;
  input \u3_mem_reg[2][25]/NET0131  ;
  input \u3_mem_reg[2][26]/NET0131  ;
  input \u3_mem_reg[2][27]/NET0131  ;
  input \u3_mem_reg[2][28]/NET0131  ;
  input \u3_mem_reg[2][29]/NET0131  ;
  input \u3_mem_reg[2][2]/NET0131  ;
  input \u3_mem_reg[2][30]/NET0131  ;
  input \u3_mem_reg[2][31]/NET0131  ;
  input \u3_mem_reg[2][3]/NET0131  ;
  input \u3_mem_reg[2][4]/NET0131  ;
  input \u3_mem_reg[2][5]/NET0131  ;
  input \u3_mem_reg[2][6]/NET0131  ;
  input \u3_mem_reg[2][7]/NET0131  ;
  input \u3_mem_reg[2][8]/NET0131  ;
  input \u3_mem_reg[2][9]/NET0131  ;
  input \u3_mem_reg[3][0]/NET0131  ;
  input \u3_mem_reg[3][10]/NET0131  ;
  input \u3_mem_reg[3][11]/NET0131  ;
  input \u3_mem_reg[3][12]/NET0131  ;
  input \u3_mem_reg[3][13]/NET0131  ;
  input \u3_mem_reg[3][14]/NET0131  ;
  input \u3_mem_reg[3][15]/NET0131  ;
  input \u3_mem_reg[3][16]/NET0131  ;
  input \u3_mem_reg[3][17]/NET0131  ;
  input \u3_mem_reg[3][18]/NET0131  ;
  input \u3_mem_reg[3][19]/NET0131  ;
  input \u3_mem_reg[3][1]/NET0131  ;
  input \u3_mem_reg[3][20]/NET0131  ;
  input \u3_mem_reg[3][21]/NET0131  ;
  input \u3_mem_reg[3][22]/NET0131  ;
  input \u3_mem_reg[3][23]/NET0131  ;
  input \u3_mem_reg[3][24]/NET0131  ;
  input \u3_mem_reg[3][25]/NET0131  ;
  input \u3_mem_reg[3][26]/NET0131  ;
  input \u3_mem_reg[3][27]/NET0131  ;
  input \u3_mem_reg[3][28]/NET0131  ;
  input \u3_mem_reg[3][29]/NET0131  ;
  input \u3_mem_reg[3][2]/NET0131  ;
  input \u3_mem_reg[3][30]/NET0131  ;
  input \u3_mem_reg[3][31]/NET0131  ;
  input \u3_mem_reg[3][3]/NET0131  ;
  input \u3_mem_reg[3][4]/NET0131  ;
  input \u3_mem_reg[3][5]/NET0131  ;
  input \u3_mem_reg[3][6]/NET0131  ;
  input \u3_mem_reg[3][7]/NET0131  ;
  input \u3_mem_reg[3][8]/NET0131  ;
  input \u3_mem_reg[3][9]/NET0131  ;
  input \u3_rp_reg[0]/P0001  ;
  input \u3_rp_reg[1]/NET0131  ;
  input \u3_rp_reg[2]/NET0131  ;
  input \u3_rp_reg[3]/NET0131  ;
  input \u3_status_reg[0]/P0001  ;
  input \u3_status_reg[1]/P0001  ;
  input \u3_wp_reg[0]/P0001  ;
  input \u3_wp_reg[1]/NET0131  ;
  input \u3_wp_reg[2]/P0001  ;
  input \u4_dout_reg[0]/P0001  ;
  input \u4_dout_reg[10]/P0001  ;
  input \u4_dout_reg[11]/P0001  ;
  input \u4_dout_reg[12]/P0001  ;
  input \u4_dout_reg[13]/P0001  ;
  input \u4_dout_reg[14]/P0001  ;
  input \u4_dout_reg[15]/P0001  ;
  input \u4_dout_reg[16]/P0001  ;
  input \u4_dout_reg[17]/P0001  ;
  input \u4_dout_reg[18]/P0001  ;
  input \u4_dout_reg[19]/P0001  ;
  input \u4_dout_reg[1]/P0001  ;
  input \u4_dout_reg[2]/P0001  ;
  input \u4_dout_reg[3]/P0001  ;
  input \u4_dout_reg[4]/P0001  ;
  input \u4_dout_reg[5]/P0001  ;
  input \u4_dout_reg[6]/P0001  ;
  input \u4_dout_reg[7]/P0001  ;
  input \u4_dout_reg[8]/P0001  ;
  input \u4_dout_reg[9]/P0001  ;
  input \u4_empty_reg/NET0131  ;
  input \u4_mem_reg[0][0]/NET0131  ;
  input \u4_mem_reg[0][10]/NET0131  ;
  input \u4_mem_reg[0][11]/NET0131  ;
  input \u4_mem_reg[0][12]/NET0131  ;
  input \u4_mem_reg[0][13]/NET0131  ;
  input \u4_mem_reg[0][14]/NET0131  ;
  input \u4_mem_reg[0][15]/NET0131  ;
  input \u4_mem_reg[0][16]/NET0131  ;
  input \u4_mem_reg[0][17]/NET0131  ;
  input \u4_mem_reg[0][18]/NET0131  ;
  input \u4_mem_reg[0][19]/NET0131  ;
  input \u4_mem_reg[0][1]/NET0131  ;
  input \u4_mem_reg[0][20]/NET0131  ;
  input \u4_mem_reg[0][21]/NET0131  ;
  input \u4_mem_reg[0][22]/NET0131  ;
  input \u4_mem_reg[0][23]/NET0131  ;
  input \u4_mem_reg[0][24]/NET0131  ;
  input \u4_mem_reg[0][25]/NET0131  ;
  input \u4_mem_reg[0][26]/NET0131  ;
  input \u4_mem_reg[0][27]/NET0131  ;
  input \u4_mem_reg[0][28]/NET0131  ;
  input \u4_mem_reg[0][29]/NET0131  ;
  input \u4_mem_reg[0][2]/NET0131  ;
  input \u4_mem_reg[0][30]/NET0131  ;
  input \u4_mem_reg[0][31]/NET0131  ;
  input \u4_mem_reg[0][3]/NET0131  ;
  input \u4_mem_reg[0][4]/NET0131  ;
  input \u4_mem_reg[0][5]/NET0131  ;
  input \u4_mem_reg[0][6]/NET0131  ;
  input \u4_mem_reg[0][7]/NET0131  ;
  input \u4_mem_reg[0][8]/NET0131  ;
  input \u4_mem_reg[0][9]/NET0131  ;
  input \u4_mem_reg[1][0]/NET0131  ;
  input \u4_mem_reg[1][10]/NET0131  ;
  input \u4_mem_reg[1][11]/NET0131  ;
  input \u4_mem_reg[1][12]/NET0131  ;
  input \u4_mem_reg[1][13]/NET0131  ;
  input \u4_mem_reg[1][14]/NET0131  ;
  input \u4_mem_reg[1][15]/NET0131  ;
  input \u4_mem_reg[1][16]/NET0131  ;
  input \u4_mem_reg[1][17]/NET0131  ;
  input \u4_mem_reg[1][18]/NET0131  ;
  input \u4_mem_reg[1][19]/NET0131  ;
  input \u4_mem_reg[1][1]/NET0131  ;
  input \u4_mem_reg[1][20]/NET0131  ;
  input \u4_mem_reg[1][21]/NET0131  ;
  input \u4_mem_reg[1][22]/NET0131  ;
  input \u4_mem_reg[1][23]/NET0131  ;
  input \u4_mem_reg[1][24]/NET0131  ;
  input \u4_mem_reg[1][25]/NET0131  ;
  input \u4_mem_reg[1][26]/NET0131  ;
  input \u4_mem_reg[1][27]/NET0131  ;
  input \u4_mem_reg[1][28]/NET0131  ;
  input \u4_mem_reg[1][29]/NET0131  ;
  input \u4_mem_reg[1][2]/NET0131  ;
  input \u4_mem_reg[1][30]/NET0131  ;
  input \u4_mem_reg[1][31]/NET0131  ;
  input \u4_mem_reg[1][3]/NET0131  ;
  input \u4_mem_reg[1][4]/NET0131  ;
  input \u4_mem_reg[1][5]/NET0131  ;
  input \u4_mem_reg[1][6]/NET0131  ;
  input \u4_mem_reg[1][7]/NET0131  ;
  input \u4_mem_reg[1][8]/NET0131  ;
  input \u4_mem_reg[1][9]/NET0131  ;
  input \u4_mem_reg[2][0]/NET0131  ;
  input \u4_mem_reg[2][10]/NET0131  ;
  input \u4_mem_reg[2][11]/NET0131  ;
  input \u4_mem_reg[2][12]/NET0131  ;
  input \u4_mem_reg[2][13]/NET0131  ;
  input \u4_mem_reg[2][14]/NET0131  ;
  input \u4_mem_reg[2][15]/NET0131  ;
  input \u4_mem_reg[2][16]/NET0131  ;
  input \u4_mem_reg[2][17]/NET0131  ;
  input \u4_mem_reg[2][18]/NET0131  ;
  input \u4_mem_reg[2][19]/NET0131  ;
  input \u4_mem_reg[2][1]/NET0131  ;
  input \u4_mem_reg[2][20]/NET0131  ;
  input \u4_mem_reg[2][21]/NET0131  ;
  input \u4_mem_reg[2][22]/NET0131  ;
  input \u4_mem_reg[2][23]/NET0131  ;
  input \u4_mem_reg[2][24]/NET0131  ;
  input \u4_mem_reg[2][25]/NET0131  ;
  input \u4_mem_reg[2][26]/NET0131  ;
  input \u4_mem_reg[2][27]/NET0131  ;
  input \u4_mem_reg[2][28]/NET0131  ;
  input \u4_mem_reg[2][29]/NET0131  ;
  input \u4_mem_reg[2][2]/NET0131  ;
  input \u4_mem_reg[2][30]/NET0131  ;
  input \u4_mem_reg[2][31]/NET0131  ;
  input \u4_mem_reg[2][3]/NET0131  ;
  input \u4_mem_reg[2][4]/NET0131  ;
  input \u4_mem_reg[2][5]/NET0131  ;
  input \u4_mem_reg[2][6]/NET0131  ;
  input \u4_mem_reg[2][7]/NET0131  ;
  input \u4_mem_reg[2][8]/NET0131  ;
  input \u4_mem_reg[2][9]/NET0131  ;
  input \u4_mem_reg[3][0]/NET0131  ;
  input \u4_mem_reg[3][10]/NET0131  ;
  input \u4_mem_reg[3][11]/NET0131  ;
  input \u4_mem_reg[3][12]/NET0131  ;
  input \u4_mem_reg[3][13]/NET0131  ;
  input \u4_mem_reg[3][14]/NET0131  ;
  input \u4_mem_reg[3][15]/NET0131  ;
  input \u4_mem_reg[3][16]/NET0131  ;
  input \u4_mem_reg[3][17]/NET0131  ;
  input \u4_mem_reg[3][18]/NET0131  ;
  input \u4_mem_reg[3][19]/NET0131  ;
  input \u4_mem_reg[3][1]/NET0131  ;
  input \u4_mem_reg[3][20]/NET0131  ;
  input \u4_mem_reg[3][21]/NET0131  ;
  input \u4_mem_reg[3][22]/NET0131  ;
  input \u4_mem_reg[3][23]/NET0131  ;
  input \u4_mem_reg[3][24]/NET0131  ;
  input \u4_mem_reg[3][25]/NET0131  ;
  input \u4_mem_reg[3][26]/NET0131  ;
  input \u4_mem_reg[3][27]/NET0131  ;
  input \u4_mem_reg[3][28]/NET0131  ;
  input \u4_mem_reg[3][29]/NET0131  ;
  input \u4_mem_reg[3][2]/NET0131  ;
  input \u4_mem_reg[3][30]/NET0131  ;
  input \u4_mem_reg[3][31]/NET0131  ;
  input \u4_mem_reg[3][3]/NET0131  ;
  input \u4_mem_reg[3][4]/NET0131  ;
  input \u4_mem_reg[3][5]/NET0131  ;
  input \u4_mem_reg[3][6]/NET0131  ;
  input \u4_mem_reg[3][7]/NET0131  ;
  input \u4_mem_reg[3][8]/NET0131  ;
  input \u4_mem_reg[3][9]/NET0131  ;
  input \u4_rp_reg[0]/P0001  ;
  input \u4_rp_reg[1]/NET0131  ;
  input \u4_rp_reg[2]/NET0131  ;
  input \u4_rp_reg[3]/NET0131  ;
  input \u4_status_reg[0]/P0001  ;
  input \u4_status_reg[1]/P0001  ;
  input \u4_wp_reg[0]/P0001  ;
  input \u4_wp_reg[1]/NET0131  ;
  input \u4_wp_reg[2]/P0001  ;
  input \u5_dout_reg[0]/P0001  ;
  input \u5_dout_reg[10]/P0001  ;
  input \u5_dout_reg[11]/P0001  ;
  input \u5_dout_reg[12]/P0001  ;
  input \u5_dout_reg[13]/P0001  ;
  input \u5_dout_reg[14]/P0001  ;
  input \u5_dout_reg[15]/P0001  ;
  input \u5_dout_reg[16]/P0001  ;
  input \u5_dout_reg[17]/P0001  ;
  input \u5_dout_reg[18]/P0001  ;
  input \u5_dout_reg[19]/P0001  ;
  input \u5_dout_reg[1]/P0001  ;
  input \u5_dout_reg[2]/P0001  ;
  input \u5_dout_reg[3]/P0001  ;
  input \u5_dout_reg[4]/P0001  ;
  input \u5_dout_reg[5]/P0001  ;
  input \u5_dout_reg[6]/P0001  ;
  input \u5_dout_reg[7]/P0001  ;
  input \u5_dout_reg[8]/P0001  ;
  input \u5_dout_reg[9]/P0001  ;
  input \u5_empty_reg/NET0131  ;
  input \u5_mem_reg[0][0]/NET0131  ;
  input \u5_mem_reg[0][10]/NET0131  ;
  input \u5_mem_reg[0][11]/NET0131  ;
  input \u5_mem_reg[0][12]/NET0131  ;
  input \u5_mem_reg[0][13]/NET0131  ;
  input \u5_mem_reg[0][14]/NET0131  ;
  input \u5_mem_reg[0][15]/NET0131  ;
  input \u5_mem_reg[0][16]/NET0131  ;
  input \u5_mem_reg[0][17]/NET0131  ;
  input \u5_mem_reg[0][18]/NET0131  ;
  input \u5_mem_reg[0][19]/NET0131  ;
  input \u5_mem_reg[0][1]/NET0131  ;
  input \u5_mem_reg[0][20]/NET0131  ;
  input \u5_mem_reg[0][21]/NET0131  ;
  input \u5_mem_reg[0][22]/NET0131  ;
  input \u5_mem_reg[0][23]/NET0131  ;
  input \u5_mem_reg[0][24]/NET0131  ;
  input \u5_mem_reg[0][25]/NET0131  ;
  input \u5_mem_reg[0][26]/NET0131  ;
  input \u5_mem_reg[0][27]/NET0131  ;
  input \u5_mem_reg[0][28]/NET0131  ;
  input \u5_mem_reg[0][29]/NET0131  ;
  input \u5_mem_reg[0][2]/NET0131  ;
  input \u5_mem_reg[0][30]/NET0131  ;
  input \u5_mem_reg[0][31]/NET0131  ;
  input \u5_mem_reg[0][3]/NET0131  ;
  input \u5_mem_reg[0][4]/NET0131  ;
  input \u5_mem_reg[0][5]/NET0131  ;
  input \u5_mem_reg[0][6]/NET0131  ;
  input \u5_mem_reg[0][7]/NET0131  ;
  input \u5_mem_reg[0][8]/NET0131  ;
  input \u5_mem_reg[0][9]/NET0131  ;
  input \u5_mem_reg[1][0]/NET0131  ;
  input \u5_mem_reg[1][10]/NET0131  ;
  input \u5_mem_reg[1][11]/NET0131  ;
  input \u5_mem_reg[1][12]/NET0131  ;
  input \u5_mem_reg[1][13]/NET0131  ;
  input \u5_mem_reg[1][14]/NET0131  ;
  input \u5_mem_reg[1][15]/NET0131  ;
  input \u5_mem_reg[1][16]/NET0131  ;
  input \u5_mem_reg[1][17]/NET0131  ;
  input \u5_mem_reg[1][18]/NET0131  ;
  input \u5_mem_reg[1][19]/NET0131  ;
  input \u5_mem_reg[1][1]/NET0131  ;
  input \u5_mem_reg[1][20]/NET0131  ;
  input \u5_mem_reg[1][21]/NET0131  ;
  input \u5_mem_reg[1][22]/NET0131  ;
  input \u5_mem_reg[1][23]/NET0131  ;
  input \u5_mem_reg[1][24]/NET0131  ;
  input \u5_mem_reg[1][25]/NET0131  ;
  input \u5_mem_reg[1][26]/NET0131  ;
  input \u5_mem_reg[1][27]/NET0131  ;
  input \u5_mem_reg[1][28]/NET0131  ;
  input \u5_mem_reg[1][29]/NET0131  ;
  input \u5_mem_reg[1][2]/NET0131  ;
  input \u5_mem_reg[1][30]/NET0131  ;
  input \u5_mem_reg[1][31]/NET0131  ;
  input \u5_mem_reg[1][3]/NET0131  ;
  input \u5_mem_reg[1][4]/NET0131  ;
  input \u5_mem_reg[1][5]/NET0131  ;
  input \u5_mem_reg[1][6]/NET0131  ;
  input \u5_mem_reg[1][7]/NET0131  ;
  input \u5_mem_reg[1][8]/NET0131  ;
  input \u5_mem_reg[1][9]/NET0131  ;
  input \u5_mem_reg[2][0]/NET0131  ;
  input \u5_mem_reg[2][10]/NET0131  ;
  input \u5_mem_reg[2][11]/NET0131  ;
  input \u5_mem_reg[2][12]/NET0131  ;
  input \u5_mem_reg[2][13]/NET0131  ;
  input \u5_mem_reg[2][14]/NET0131  ;
  input \u5_mem_reg[2][15]/NET0131  ;
  input \u5_mem_reg[2][16]/NET0131  ;
  input \u5_mem_reg[2][17]/NET0131  ;
  input \u5_mem_reg[2][18]/NET0131  ;
  input \u5_mem_reg[2][19]/NET0131  ;
  input \u5_mem_reg[2][1]/NET0131  ;
  input \u5_mem_reg[2][20]/NET0131  ;
  input \u5_mem_reg[2][21]/NET0131  ;
  input \u5_mem_reg[2][22]/NET0131  ;
  input \u5_mem_reg[2][23]/NET0131  ;
  input \u5_mem_reg[2][24]/NET0131  ;
  input \u5_mem_reg[2][25]/NET0131  ;
  input \u5_mem_reg[2][26]/NET0131  ;
  input \u5_mem_reg[2][27]/NET0131  ;
  input \u5_mem_reg[2][28]/NET0131  ;
  input \u5_mem_reg[2][29]/NET0131  ;
  input \u5_mem_reg[2][2]/NET0131  ;
  input \u5_mem_reg[2][30]/NET0131  ;
  input \u5_mem_reg[2][31]/NET0131  ;
  input \u5_mem_reg[2][3]/NET0131  ;
  input \u5_mem_reg[2][4]/NET0131  ;
  input \u5_mem_reg[2][5]/NET0131  ;
  input \u5_mem_reg[2][6]/NET0131  ;
  input \u5_mem_reg[2][7]/NET0131  ;
  input \u5_mem_reg[2][8]/NET0131  ;
  input \u5_mem_reg[2][9]/NET0131  ;
  input \u5_mem_reg[3][0]/NET0131  ;
  input \u5_mem_reg[3][10]/NET0131  ;
  input \u5_mem_reg[3][11]/NET0131  ;
  input \u5_mem_reg[3][12]/NET0131  ;
  input \u5_mem_reg[3][13]/NET0131  ;
  input \u5_mem_reg[3][14]/NET0131  ;
  input \u5_mem_reg[3][15]/NET0131  ;
  input \u5_mem_reg[3][16]/NET0131  ;
  input \u5_mem_reg[3][17]/NET0131  ;
  input \u5_mem_reg[3][18]/NET0131  ;
  input \u5_mem_reg[3][19]/NET0131  ;
  input \u5_mem_reg[3][1]/NET0131  ;
  input \u5_mem_reg[3][20]/NET0131  ;
  input \u5_mem_reg[3][21]/NET0131  ;
  input \u5_mem_reg[3][22]/NET0131  ;
  input \u5_mem_reg[3][23]/NET0131  ;
  input \u5_mem_reg[3][24]/NET0131  ;
  input \u5_mem_reg[3][25]/NET0131  ;
  input \u5_mem_reg[3][26]/NET0131  ;
  input \u5_mem_reg[3][27]/NET0131  ;
  input \u5_mem_reg[3][28]/NET0131  ;
  input \u5_mem_reg[3][29]/NET0131  ;
  input \u5_mem_reg[3][2]/NET0131  ;
  input \u5_mem_reg[3][30]/NET0131  ;
  input \u5_mem_reg[3][31]/NET0131  ;
  input \u5_mem_reg[3][3]/NET0131  ;
  input \u5_mem_reg[3][4]/NET0131  ;
  input \u5_mem_reg[3][5]/NET0131  ;
  input \u5_mem_reg[3][6]/NET0131  ;
  input \u5_mem_reg[3][7]/NET0131  ;
  input \u5_mem_reg[3][8]/NET0131  ;
  input \u5_mem_reg[3][9]/NET0131  ;
  input \u5_rp_reg[0]/P0001  ;
  input \u5_rp_reg[1]/NET0131  ;
  input \u5_rp_reg[2]/NET0131  ;
  input \u5_rp_reg[3]/NET0131  ;
  input \u5_status_reg[0]/P0001  ;
  input \u5_status_reg[1]/P0001  ;
  input \u5_wp_reg[0]/P0001  ;
  input \u5_wp_reg[1]/NET0131  ;
  input \u5_wp_reg[2]/P0001  ;
  input \u6_dout_reg[0]/P0001  ;
  input \u6_dout_reg[10]/P0001  ;
  input \u6_dout_reg[11]/P0001  ;
  input \u6_dout_reg[12]/P0001  ;
  input \u6_dout_reg[13]/P0001  ;
  input \u6_dout_reg[14]/P0001  ;
  input \u6_dout_reg[15]/P0001  ;
  input \u6_dout_reg[16]/P0001  ;
  input \u6_dout_reg[17]/P0001  ;
  input \u6_dout_reg[18]/P0001  ;
  input \u6_dout_reg[19]/P0001  ;
  input \u6_dout_reg[1]/P0001  ;
  input \u6_dout_reg[2]/P0001  ;
  input \u6_dout_reg[3]/P0001  ;
  input \u6_dout_reg[4]/P0001  ;
  input \u6_dout_reg[5]/P0001  ;
  input \u6_dout_reg[6]/P0001  ;
  input \u6_dout_reg[7]/P0001  ;
  input \u6_dout_reg[8]/P0001  ;
  input \u6_dout_reg[9]/P0001  ;
  input \u6_empty_reg/NET0131  ;
  input \u6_mem_reg[0][0]/NET0131  ;
  input \u6_mem_reg[0][10]/NET0131  ;
  input \u6_mem_reg[0][11]/NET0131  ;
  input \u6_mem_reg[0][12]/NET0131  ;
  input \u6_mem_reg[0][13]/NET0131  ;
  input \u6_mem_reg[0][14]/NET0131  ;
  input \u6_mem_reg[0][15]/NET0131  ;
  input \u6_mem_reg[0][16]/NET0131  ;
  input \u6_mem_reg[0][17]/NET0131  ;
  input \u6_mem_reg[0][18]/NET0131  ;
  input \u6_mem_reg[0][19]/NET0131  ;
  input \u6_mem_reg[0][1]/NET0131  ;
  input \u6_mem_reg[0][20]/NET0131  ;
  input \u6_mem_reg[0][21]/NET0131  ;
  input \u6_mem_reg[0][22]/NET0131  ;
  input \u6_mem_reg[0][23]/NET0131  ;
  input \u6_mem_reg[0][24]/NET0131  ;
  input \u6_mem_reg[0][25]/NET0131  ;
  input \u6_mem_reg[0][26]/NET0131  ;
  input \u6_mem_reg[0][27]/NET0131  ;
  input \u6_mem_reg[0][28]/NET0131  ;
  input \u6_mem_reg[0][29]/NET0131  ;
  input \u6_mem_reg[0][2]/NET0131  ;
  input \u6_mem_reg[0][30]/NET0131  ;
  input \u6_mem_reg[0][31]/NET0131  ;
  input \u6_mem_reg[0][3]/NET0131  ;
  input \u6_mem_reg[0][4]/NET0131  ;
  input \u6_mem_reg[0][5]/NET0131  ;
  input \u6_mem_reg[0][6]/NET0131  ;
  input \u6_mem_reg[0][7]/NET0131  ;
  input \u6_mem_reg[0][8]/NET0131  ;
  input \u6_mem_reg[0][9]/NET0131  ;
  input \u6_mem_reg[1][0]/NET0131  ;
  input \u6_mem_reg[1][10]/NET0131  ;
  input \u6_mem_reg[1][11]/NET0131  ;
  input \u6_mem_reg[1][12]/NET0131  ;
  input \u6_mem_reg[1][13]/NET0131  ;
  input \u6_mem_reg[1][14]/NET0131  ;
  input \u6_mem_reg[1][15]/NET0131  ;
  input \u6_mem_reg[1][16]/NET0131  ;
  input \u6_mem_reg[1][17]/NET0131  ;
  input \u6_mem_reg[1][18]/NET0131  ;
  input \u6_mem_reg[1][19]/NET0131  ;
  input \u6_mem_reg[1][1]/NET0131  ;
  input \u6_mem_reg[1][20]/NET0131  ;
  input \u6_mem_reg[1][21]/NET0131  ;
  input \u6_mem_reg[1][22]/NET0131  ;
  input \u6_mem_reg[1][23]/NET0131  ;
  input \u6_mem_reg[1][24]/NET0131  ;
  input \u6_mem_reg[1][25]/NET0131  ;
  input \u6_mem_reg[1][26]/NET0131  ;
  input \u6_mem_reg[1][27]/NET0131  ;
  input \u6_mem_reg[1][28]/NET0131  ;
  input \u6_mem_reg[1][29]/NET0131  ;
  input \u6_mem_reg[1][2]/NET0131  ;
  input \u6_mem_reg[1][30]/NET0131  ;
  input \u6_mem_reg[1][31]/NET0131  ;
  input \u6_mem_reg[1][3]/NET0131  ;
  input \u6_mem_reg[1][4]/NET0131  ;
  input \u6_mem_reg[1][5]/NET0131  ;
  input \u6_mem_reg[1][6]/NET0131  ;
  input \u6_mem_reg[1][7]/NET0131  ;
  input \u6_mem_reg[1][8]/NET0131  ;
  input \u6_mem_reg[1][9]/NET0131  ;
  input \u6_mem_reg[2][0]/NET0131  ;
  input \u6_mem_reg[2][10]/NET0131  ;
  input \u6_mem_reg[2][11]/NET0131  ;
  input \u6_mem_reg[2][12]/NET0131  ;
  input \u6_mem_reg[2][13]/NET0131  ;
  input \u6_mem_reg[2][14]/NET0131  ;
  input \u6_mem_reg[2][15]/NET0131  ;
  input \u6_mem_reg[2][16]/NET0131  ;
  input \u6_mem_reg[2][17]/NET0131  ;
  input \u6_mem_reg[2][18]/NET0131  ;
  input \u6_mem_reg[2][19]/NET0131  ;
  input \u6_mem_reg[2][1]/NET0131  ;
  input \u6_mem_reg[2][20]/NET0131  ;
  input \u6_mem_reg[2][21]/NET0131  ;
  input \u6_mem_reg[2][22]/NET0131  ;
  input \u6_mem_reg[2][23]/NET0131  ;
  input \u6_mem_reg[2][24]/NET0131  ;
  input \u6_mem_reg[2][25]/NET0131  ;
  input \u6_mem_reg[2][26]/NET0131  ;
  input \u6_mem_reg[2][27]/NET0131  ;
  input \u6_mem_reg[2][28]/NET0131  ;
  input \u6_mem_reg[2][29]/NET0131  ;
  input \u6_mem_reg[2][2]/NET0131  ;
  input \u6_mem_reg[2][30]/NET0131  ;
  input \u6_mem_reg[2][31]/NET0131  ;
  input \u6_mem_reg[2][3]/NET0131  ;
  input \u6_mem_reg[2][4]/NET0131  ;
  input \u6_mem_reg[2][5]/NET0131  ;
  input \u6_mem_reg[2][6]/NET0131  ;
  input \u6_mem_reg[2][7]/NET0131  ;
  input \u6_mem_reg[2][8]/NET0131  ;
  input \u6_mem_reg[2][9]/NET0131  ;
  input \u6_mem_reg[3][0]/NET0131  ;
  input \u6_mem_reg[3][10]/NET0131  ;
  input \u6_mem_reg[3][11]/NET0131  ;
  input \u6_mem_reg[3][12]/NET0131  ;
  input \u6_mem_reg[3][13]/NET0131  ;
  input \u6_mem_reg[3][14]/NET0131  ;
  input \u6_mem_reg[3][15]/NET0131  ;
  input \u6_mem_reg[3][16]/NET0131  ;
  input \u6_mem_reg[3][17]/NET0131  ;
  input \u6_mem_reg[3][18]/NET0131  ;
  input \u6_mem_reg[3][19]/NET0131  ;
  input \u6_mem_reg[3][1]/NET0131  ;
  input \u6_mem_reg[3][20]/NET0131  ;
  input \u6_mem_reg[3][21]/NET0131  ;
  input \u6_mem_reg[3][22]/NET0131  ;
  input \u6_mem_reg[3][23]/NET0131  ;
  input \u6_mem_reg[3][24]/NET0131  ;
  input \u6_mem_reg[3][25]/NET0131  ;
  input \u6_mem_reg[3][26]/NET0131  ;
  input \u6_mem_reg[3][27]/NET0131  ;
  input \u6_mem_reg[3][28]/NET0131  ;
  input \u6_mem_reg[3][29]/NET0131  ;
  input \u6_mem_reg[3][2]/NET0131  ;
  input \u6_mem_reg[3][30]/NET0131  ;
  input \u6_mem_reg[3][31]/NET0131  ;
  input \u6_mem_reg[3][3]/NET0131  ;
  input \u6_mem_reg[3][4]/NET0131  ;
  input \u6_mem_reg[3][5]/NET0131  ;
  input \u6_mem_reg[3][6]/NET0131  ;
  input \u6_mem_reg[3][7]/NET0131  ;
  input \u6_mem_reg[3][8]/NET0131  ;
  input \u6_mem_reg[3][9]/NET0131  ;
  input \u6_rp_reg[0]/P0001  ;
  input \u6_rp_reg[1]/NET0131  ;
  input \u6_rp_reg[2]/NET0131  ;
  input \u6_rp_reg[3]/NET0131  ;
  input \u6_status_reg[0]/P0001  ;
  input \u6_status_reg[1]/P0001  ;
  input \u6_wp_reg[0]/P0001  ;
  input \u6_wp_reg[1]/NET0131  ;
  input \u6_wp_reg[2]/P0001  ;
  input \u7_dout_reg[0]/P0001  ;
  input \u7_dout_reg[10]/P0001  ;
  input \u7_dout_reg[11]/P0001  ;
  input \u7_dout_reg[12]/P0001  ;
  input \u7_dout_reg[13]/P0001  ;
  input \u7_dout_reg[14]/P0001  ;
  input \u7_dout_reg[15]/P0001  ;
  input \u7_dout_reg[16]/P0001  ;
  input \u7_dout_reg[17]/P0001  ;
  input \u7_dout_reg[18]/P0001  ;
  input \u7_dout_reg[19]/P0001  ;
  input \u7_dout_reg[1]/P0001  ;
  input \u7_dout_reg[2]/P0001  ;
  input \u7_dout_reg[3]/P0001  ;
  input \u7_dout_reg[4]/P0001  ;
  input \u7_dout_reg[5]/P0001  ;
  input \u7_dout_reg[6]/P0001  ;
  input \u7_dout_reg[7]/P0001  ;
  input \u7_dout_reg[8]/P0001  ;
  input \u7_dout_reg[9]/P0001  ;
  input \u7_empty_reg/NET0131  ;
  input \u7_mem_reg[0][0]/NET0131  ;
  input \u7_mem_reg[0][10]/NET0131  ;
  input \u7_mem_reg[0][11]/NET0131  ;
  input \u7_mem_reg[0][12]/NET0131  ;
  input \u7_mem_reg[0][13]/NET0131  ;
  input \u7_mem_reg[0][14]/NET0131  ;
  input \u7_mem_reg[0][15]/NET0131  ;
  input \u7_mem_reg[0][16]/NET0131  ;
  input \u7_mem_reg[0][17]/NET0131  ;
  input \u7_mem_reg[0][18]/NET0131  ;
  input \u7_mem_reg[0][19]/NET0131  ;
  input \u7_mem_reg[0][1]/NET0131  ;
  input \u7_mem_reg[0][20]/NET0131  ;
  input \u7_mem_reg[0][21]/NET0131  ;
  input \u7_mem_reg[0][22]/NET0131  ;
  input \u7_mem_reg[0][23]/NET0131  ;
  input \u7_mem_reg[0][24]/NET0131  ;
  input \u7_mem_reg[0][25]/NET0131  ;
  input \u7_mem_reg[0][26]/NET0131  ;
  input \u7_mem_reg[0][27]/NET0131  ;
  input \u7_mem_reg[0][28]/NET0131  ;
  input \u7_mem_reg[0][29]/NET0131  ;
  input \u7_mem_reg[0][2]/NET0131  ;
  input \u7_mem_reg[0][30]/NET0131  ;
  input \u7_mem_reg[0][31]/NET0131  ;
  input \u7_mem_reg[0][3]/NET0131  ;
  input \u7_mem_reg[0][4]/NET0131  ;
  input \u7_mem_reg[0][5]/NET0131  ;
  input \u7_mem_reg[0][6]/NET0131  ;
  input \u7_mem_reg[0][7]/NET0131  ;
  input \u7_mem_reg[0][8]/NET0131  ;
  input \u7_mem_reg[0][9]/NET0131  ;
  input \u7_mem_reg[1][0]/NET0131  ;
  input \u7_mem_reg[1][10]/NET0131  ;
  input \u7_mem_reg[1][11]/NET0131  ;
  input \u7_mem_reg[1][12]/NET0131  ;
  input \u7_mem_reg[1][13]/NET0131  ;
  input \u7_mem_reg[1][14]/NET0131  ;
  input \u7_mem_reg[1][15]/NET0131  ;
  input \u7_mem_reg[1][16]/NET0131  ;
  input \u7_mem_reg[1][17]/NET0131  ;
  input \u7_mem_reg[1][18]/NET0131  ;
  input \u7_mem_reg[1][19]/NET0131  ;
  input \u7_mem_reg[1][1]/NET0131  ;
  input \u7_mem_reg[1][20]/NET0131  ;
  input \u7_mem_reg[1][21]/NET0131  ;
  input \u7_mem_reg[1][22]/NET0131  ;
  input \u7_mem_reg[1][23]/NET0131  ;
  input \u7_mem_reg[1][24]/NET0131  ;
  input \u7_mem_reg[1][25]/NET0131  ;
  input \u7_mem_reg[1][26]/NET0131  ;
  input \u7_mem_reg[1][27]/NET0131  ;
  input \u7_mem_reg[1][28]/NET0131  ;
  input \u7_mem_reg[1][29]/NET0131  ;
  input \u7_mem_reg[1][2]/NET0131  ;
  input \u7_mem_reg[1][30]/NET0131  ;
  input \u7_mem_reg[1][31]/NET0131  ;
  input \u7_mem_reg[1][3]/NET0131  ;
  input \u7_mem_reg[1][4]/NET0131  ;
  input \u7_mem_reg[1][5]/NET0131  ;
  input \u7_mem_reg[1][6]/NET0131  ;
  input \u7_mem_reg[1][7]/NET0131  ;
  input \u7_mem_reg[1][8]/NET0131  ;
  input \u7_mem_reg[1][9]/NET0131  ;
  input \u7_mem_reg[2][0]/NET0131  ;
  input \u7_mem_reg[2][10]/NET0131  ;
  input \u7_mem_reg[2][11]/NET0131  ;
  input \u7_mem_reg[2][12]/NET0131  ;
  input \u7_mem_reg[2][13]/NET0131  ;
  input \u7_mem_reg[2][14]/NET0131  ;
  input \u7_mem_reg[2][15]/NET0131  ;
  input \u7_mem_reg[2][16]/NET0131  ;
  input \u7_mem_reg[2][17]/NET0131  ;
  input \u7_mem_reg[2][18]/NET0131  ;
  input \u7_mem_reg[2][19]/NET0131  ;
  input \u7_mem_reg[2][1]/NET0131  ;
  input \u7_mem_reg[2][20]/NET0131  ;
  input \u7_mem_reg[2][21]/NET0131  ;
  input \u7_mem_reg[2][22]/NET0131  ;
  input \u7_mem_reg[2][23]/NET0131  ;
  input \u7_mem_reg[2][24]/NET0131  ;
  input \u7_mem_reg[2][25]/NET0131  ;
  input \u7_mem_reg[2][26]/NET0131  ;
  input \u7_mem_reg[2][27]/NET0131  ;
  input \u7_mem_reg[2][28]/NET0131  ;
  input \u7_mem_reg[2][29]/NET0131  ;
  input \u7_mem_reg[2][2]/NET0131  ;
  input \u7_mem_reg[2][30]/NET0131  ;
  input \u7_mem_reg[2][31]/NET0131  ;
  input \u7_mem_reg[2][3]/NET0131  ;
  input \u7_mem_reg[2][4]/NET0131  ;
  input \u7_mem_reg[2][5]/NET0131  ;
  input \u7_mem_reg[2][6]/NET0131  ;
  input \u7_mem_reg[2][7]/NET0131  ;
  input \u7_mem_reg[2][8]/NET0131  ;
  input \u7_mem_reg[2][9]/NET0131  ;
  input \u7_mem_reg[3][0]/NET0131  ;
  input \u7_mem_reg[3][10]/NET0131  ;
  input \u7_mem_reg[3][11]/NET0131  ;
  input \u7_mem_reg[3][12]/NET0131  ;
  input \u7_mem_reg[3][13]/NET0131  ;
  input \u7_mem_reg[3][14]/NET0131  ;
  input \u7_mem_reg[3][15]/NET0131  ;
  input \u7_mem_reg[3][16]/NET0131  ;
  input \u7_mem_reg[3][17]/NET0131  ;
  input \u7_mem_reg[3][18]/NET0131  ;
  input \u7_mem_reg[3][19]/NET0131  ;
  input \u7_mem_reg[3][1]/NET0131  ;
  input \u7_mem_reg[3][20]/NET0131  ;
  input \u7_mem_reg[3][21]/NET0131  ;
  input \u7_mem_reg[3][22]/NET0131  ;
  input \u7_mem_reg[3][23]/NET0131  ;
  input \u7_mem_reg[3][24]/NET0131  ;
  input \u7_mem_reg[3][25]/NET0131  ;
  input \u7_mem_reg[3][26]/NET0131  ;
  input \u7_mem_reg[3][27]/NET0131  ;
  input \u7_mem_reg[3][28]/NET0131  ;
  input \u7_mem_reg[3][29]/NET0131  ;
  input \u7_mem_reg[3][2]/NET0131  ;
  input \u7_mem_reg[3][30]/NET0131  ;
  input \u7_mem_reg[3][31]/NET0131  ;
  input \u7_mem_reg[3][3]/NET0131  ;
  input \u7_mem_reg[3][4]/NET0131  ;
  input \u7_mem_reg[3][5]/NET0131  ;
  input \u7_mem_reg[3][6]/NET0131  ;
  input \u7_mem_reg[3][7]/NET0131  ;
  input \u7_mem_reg[3][8]/NET0131  ;
  input \u7_mem_reg[3][9]/NET0131  ;
  input \u7_rp_reg[0]/P0001  ;
  input \u7_rp_reg[1]/NET0131  ;
  input \u7_rp_reg[2]/NET0131  ;
  input \u7_rp_reg[3]/NET0131  ;
  input \u7_status_reg[0]/P0001  ;
  input \u7_status_reg[1]/P0001  ;
  input \u7_wp_reg[0]/P0001  ;
  input \u7_wp_reg[1]/NET0131  ;
  input \u7_wp_reg[2]/P0001  ;
  input \u8_dout_reg[0]/P0001  ;
  input \u8_dout_reg[10]/P0001  ;
  input \u8_dout_reg[11]/P0001  ;
  input \u8_dout_reg[12]/P0001  ;
  input \u8_dout_reg[13]/P0001  ;
  input \u8_dout_reg[14]/P0001  ;
  input \u8_dout_reg[15]/P0001  ;
  input \u8_dout_reg[16]/P0001  ;
  input \u8_dout_reg[17]/P0001  ;
  input \u8_dout_reg[18]/P0001  ;
  input \u8_dout_reg[19]/P0001  ;
  input \u8_dout_reg[1]/P0001  ;
  input \u8_dout_reg[2]/P0001  ;
  input \u8_dout_reg[3]/P0001  ;
  input \u8_dout_reg[4]/P0001  ;
  input \u8_dout_reg[5]/P0001  ;
  input \u8_dout_reg[6]/P0001  ;
  input \u8_dout_reg[7]/P0001  ;
  input \u8_dout_reg[8]/P0001  ;
  input \u8_dout_reg[9]/P0001  ;
  input \u8_empty_reg/NET0131  ;
  input \u8_mem_reg[0][0]/NET0131  ;
  input \u8_mem_reg[0][10]/NET0131  ;
  input \u8_mem_reg[0][11]/NET0131  ;
  input \u8_mem_reg[0][12]/NET0131  ;
  input \u8_mem_reg[0][13]/NET0131  ;
  input \u8_mem_reg[0][14]/NET0131  ;
  input \u8_mem_reg[0][15]/NET0131  ;
  input \u8_mem_reg[0][16]/NET0131  ;
  input \u8_mem_reg[0][17]/NET0131  ;
  input \u8_mem_reg[0][18]/NET0131  ;
  input \u8_mem_reg[0][19]/NET0131  ;
  input \u8_mem_reg[0][1]/NET0131  ;
  input \u8_mem_reg[0][20]/NET0131  ;
  input \u8_mem_reg[0][21]/NET0131  ;
  input \u8_mem_reg[0][22]/NET0131  ;
  input \u8_mem_reg[0][23]/NET0131  ;
  input \u8_mem_reg[0][24]/NET0131  ;
  input \u8_mem_reg[0][25]/NET0131  ;
  input \u8_mem_reg[0][26]/NET0131  ;
  input \u8_mem_reg[0][27]/NET0131  ;
  input \u8_mem_reg[0][28]/NET0131  ;
  input \u8_mem_reg[0][29]/NET0131  ;
  input \u8_mem_reg[0][2]/NET0131  ;
  input \u8_mem_reg[0][30]/NET0131  ;
  input \u8_mem_reg[0][31]/NET0131  ;
  input \u8_mem_reg[0][3]/NET0131  ;
  input \u8_mem_reg[0][4]/NET0131  ;
  input \u8_mem_reg[0][5]/NET0131  ;
  input \u8_mem_reg[0][6]/NET0131  ;
  input \u8_mem_reg[0][7]/NET0131  ;
  input \u8_mem_reg[0][8]/NET0131  ;
  input \u8_mem_reg[0][9]/NET0131  ;
  input \u8_mem_reg[1][0]/NET0131  ;
  input \u8_mem_reg[1][10]/NET0131  ;
  input \u8_mem_reg[1][11]/NET0131  ;
  input \u8_mem_reg[1][12]/NET0131  ;
  input \u8_mem_reg[1][13]/NET0131  ;
  input \u8_mem_reg[1][14]/NET0131  ;
  input \u8_mem_reg[1][15]/NET0131  ;
  input \u8_mem_reg[1][16]/NET0131  ;
  input \u8_mem_reg[1][17]/NET0131  ;
  input \u8_mem_reg[1][18]/NET0131  ;
  input \u8_mem_reg[1][19]/NET0131  ;
  input \u8_mem_reg[1][1]/NET0131  ;
  input \u8_mem_reg[1][20]/NET0131  ;
  input \u8_mem_reg[1][21]/NET0131  ;
  input \u8_mem_reg[1][22]/NET0131  ;
  input \u8_mem_reg[1][23]/NET0131  ;
  input \u8_mem_reg[1][24]/NET0131  ;
  input \u8_mem_reg[1][25]/NET0131  ;
  input \u8_mem_reg[1][26]/NET0131  ;
  input \u8_mem_reg[1][27]/NET0131  ;
  input \u8_mem_reg[1][28]/NET0131  ;
  input \u8_mem_reg[1][29]/NET0131  ;
  input \u8_mem_reg[1][2]/NET0131  ;
  input \u8_mem_reg[1][30]/NET0131  ;
  input \u8_mem_reg[1][31]/NET0131  ;
  input \u8_mem_reg[1][3]/NET0131  ;
  input \u8_mem_reg[1][4]/NET0131  ;
  input \u8_mem_reg[1][5]/NET0131  ;
  input \u8_mem_reg[1][6]/NET0131  ;
  input \u8_mem_reg[1][7]/NET0131  ;
  input \u8_mem_reg[1][8]/NET0131  ;
  input \u8_mem_reg[1][9]/NET0131  ;
  input \u8_mem_reg[2][0]/NET0131  ;
  input \u8_mem_reg[2][10]/NET0131  ;
  input \u8_mem_reg[2][11]/NET0131  ;
  input \u8_mem_reg[2][12]/NET0131  ;
  input \u8_mem_reg[2][13]/NET0131  ;
  input \u8_mem_reg[2][14]/NET0131  ;
  input \u8_mem_reg[2][15]/NET0131  ;
  input \u8_mem_reg[2][16]/NET0131  ;
  input \u8_mem_reg[2][17]/NET0131  ;
  input \u8_mem_reg[2][18]/NET0131  ;
  input \u8_mem_reg[2][19]/NET0131  ;
  input \u8_mem_reg[2][1]/NET0131  ;
  input \u8_mem_reg[2][20]/NET0131  ;
  input \u8_mem_reg[2][21]/NET0131  ;
  input \u8_mem_reg[2][22]/NET0131  ;
  input \u8_mem_reg[2][23]/NET0131  ;
  input \u8_mem_reg[2][24]/NET0131  ;
  input \u8_mem_reg[2][25]/NET0131  ;
  input \u8_mem_reg[2][26]/NET0131  ;
  input \u8_mem_reg[2][27]/NET0131  ;
  input \u8_mem_reg[2][28]/NET0131  ;
  input \u8_mem_reg[2][29]/NET0131  ;
  input \u8_mem_reg[2][2]/NET0131  ;
  input \u8_mem_reg[2][30]/NET0131  ;
  input \u8_mem_reg[2][31]/NET0131  ;
  input \u8_mem_reg[2][3]/NET0131  ;
  input \u8_mem_reg[2][4]/NET0131  ;
  input \u8_mem_reg[2][5]/NET0131  ;
  input \u8_mem_reg[2][6]/NET0131  ;
  input \u8_mem_reg[2][7]/NET0131  ;
  input \u8_mem_reg[2][8]/NET0131  ;
  input \u8_mem_reg[2][9]/NET0131  ;
  input \u8_mem_reg[3][0]/NET0131  ;
  input \u8_mem_reg[3][10]/NET0131  ;
  input \u8_mem_reg[3][11]/NET0131  ;
  input \u8_mem_reg[3][12]/NET0131  ;
  input \u8_mem_reg[3][13]/NET0131  ;
  input \u8_mem_reg[3][14]/NET0131  ;
  input \u8_mem_reg[3][15]/NET0131  ;
  input \u8_mem_reg[3][16]/NET0131  ;
  input \u8_mem_reg[3][17]/NET0131  ;
  input \u8_mem_reg[3][18]/NET0131  ;
  input \u8_mem_reg[3][19]/NET0131  ;
  input \u8_mem_reg[3][1]/NET0131  ;
  input \u8_mem_reg[3][20]/NET0131  ;
  input \u8_mem_reg[3][21]/NET0131  ;
  input \u8_mem_reg[3][22]/NET0131  ;
  input \u8_mem_reg[3][23]/NET0131  ;
  input \u8_mem_reg[3][24]/NET0131  ;
  input \u8_mem_reg[3][25]/NET0131  ;
  input \u8_mem_reg[3][26]/NET0131  ;
  input \u8_mem_reg[3][27]/NET0131  ;
  input \u8_mem_reg[3][28]/NET0131  ;
  input \u8_mem_reg[3][29]/NET0131  ;
  input \u8_mem_reg[3][2]/NET0131  ;
  input \u8_mem_reg[3][30]/NET0131  ;
  input \u8_mem_reg[3][31]/NET0131  ;
  input \u8_mem_reg[3][3]/NET0131  ;
  input \u8_mem_reg[3][4]/NET0131  ;
  input \u8_mem_reg[3][5]/NET0131  ;
  input \u8_mem_reg[3][6]/NET0131  ;
  input \u8_mem_reg[3][7]/NET0131  ;
  input \u8_mem_reg[3][8]/NET0131  ;
  input \u8_mem_reg[3][9]/NET0131  ;
  input \u8_rp_reg[0]/P0001  ;
  input \u8_rp_reg[1]/NET0131  ;
  input \u8_rp_reg[2]/NET0131  ;
  input \u8_rp_reg[3]/NET0131  ;
  input \u8_status_reg[0]/P0001  ;
  input \u8_status_reg[1]/P0001  ;
  input \u8_wp_reg[0]/P0001  ;
  input \u8_wp_reg[1]/NET0131  ;
  input \u8_wp_reg[2]/P0001  ;
  input \u9_din_tmp1_reg[0]/P0001  ;
  input \u9_din_tmp1_reg[10]/P0001  ;
  input \u9_din_tmp1_reg[11]/P0001  ;
  input \u9_din_tmp1_reg[12]/P0001  ;
  input \u9_din_tmp1_reg[13]/P0001  ;
  input \u9_din_tmp1_reg[14]/P0001  ;
  input \u9_din_tmp1_reg[15]/P0001  ;
  input \u9_din_tmp1_reg[1]/P0001  ;
  input \u9_din_tmp1_reg[2]/P0001  ;
  input \u9_din_tmp1_reg[3]/P0001  ;
  input \u9_din_tmp1_reg[4]/P0001  ;
  input \u9_din_tmp1_reg[5]/P0001  ;
  input \u9_din_tmp1_reg[6]/P0001  ;
  input \u9_din_tmp1_reg[7]/P0001  ;
  input \u9_din_tmp1_reg[8]/P0001  ;
  input \u9_din_tmp1_reg[9]/P0001  ;
  input \u9_dout_reg[0]/P0001  ;
  input \u9_dout_reg[10]/P0001  ;
  input \u9_dout_reg[11]/P0001  ;
  input \u9_dout_reg[12]/P0001  ;
  input \u9_dout_reg[13]/P0001  ;
  input \u9_dout_reg[14]/P0001  ;
  input \u9_dout_reg[15]/P0001  ;
  input \u9_dout_reg[16]/P0001  ;
  input \u9_dout_reg[17]/P0001  ;
  input \u9_dout_reg[18]/P0001  ;
  input \u9_dout_reg[19]/P0001  ;
  input \u9_dout_reg[1]/P0001  ;
  input \u9_dout_reg[20]/P0001  ;
  input \u9_dout_reg[21]/P0001  ;
  input \u9_dout_reg[22]/P0001  ;
  input \u9_dout_reg[23]/P0001  ;
  input \u9_dout_reg[24]/P0001  ;
  input \u9_dout_reg[25]/P0001  ;
  input \u9_dout_reg[26]/P0001  ;
  input \u9_dout_reg[27]/P0001  ;
  input \u9_dout_reg[28]/P0001  ;
  input \u9_dout_reg[29]/P0001  ;
  input \u9_dout_reg[2]/P0001  ;
  input \u9_dout_reg[30]/P0001  ;
  input \u9_dout_reg[31]/P0001  ;
  input \u9_dout_reg[3]/P0001  ;
  input \u9_dout_reg[4]/P0001  ;
  input \u9_dout_reg[5]/P0001  ;
  input \u9_dout_reg[6]/P0001  ;
  input \u9_dout_reg[7]/P0001  ;
  input \u9_dout_reg[8]/P0001  ;
  input \u9_dout_reg[9]/P0001  ;
  input \u9_empty_reg/P0001  ;
  input \u9_full_reg/NET0131  ;
  input \u9_mem_reg[0][0]/P0001  ;
  input \u9_mem_reg[0][10]/P0001  ;
  input \u9_mem_reg[0][11]/P0001  ;
  input \u9_mem_reg[0][12]/P0001  ;
  input \u9_mem_reg[0][13]/P0001  ;
  input \u9_mem_reg[0][14]/P0001  ;
  input \u9_mem_reg[0][15]/P0001  ;
  input \u9_mem_reg[0][16]/P0001  ;
  input \u9_mem_reg[0][17]/P0001  ;
  input \u9_mem_reg[0][18]/P0001  ;
  input \u9_mem_reg[0][19]/P0001  ;
  input \u9_mem_reg[0][1]/P0001  ;
  input \u9_mem_reg[0][20]/P0001  ;
  input \u9_mem_reg[0][21]/P0001  ;
  input \u9_mem_reg[0][22]/P0001  ;
  input \u9_mem_reg[0][23]/P0001  ;
  input \u9_mem_reg[0][24]/P0001  ;
  input \u9_mem_reg[0][25]/P0001  ;
  input \u9_mem_reg[0][26]/P0001  ;
  input \u9_mem_reg[0][27]/P0001  ;
  input \u9_mem_reg[0][28]/P0001  ;
  input \u9_mem_reg[0][29]/P0001  ;
  input \u9_mem_reg[0][2]/P0001  ;
  input \u9_mem_reg[0][30]/P0001  ;
  input \u9_mem_reg[0][31]/P0001  ;
  input \u9_mem_reg[0][3]/P0001  ;
  input \u9_mem_reg[0][4]/P0001  ;
  input \u9_mem_reg[0][5]/P0001  ;
  input \u9_mem_reg[0][6]/P0001  ;
  input \u9_mem_reg[0][7]/P0001  ;
  input \u9_mem_reg[0][8]/P0001  ;
  input \u9_mem_reg[0][9]/P0001  ;
  input \u9_mem_reg[1][0]/P0001  ;
  input \u9_mem_reg[1][10]/P0001  ;
  input \u9_mem_reg[1][11]/P0001  ;
  input \u9_mem_reg[1][12]/P0001  ;
  input \u9_mem_reg[1][13]/P0001  ;
  input \u9_mem_reg[1][14]/P0001  ;
  input \u9_mem_reg[1][15]/P0001  ;
  input \u9_mem_reg[1][16]/P0001  ;
  input \u9_mem_reg[1][17]/P0001  ;
  input \u9_mem_reg[1][18]/P0001  ;
  input \u9_mem_reg[1][19]/P0001  ;
  input \u9_mem_reg[1][1]/P0001  ;
  input \u9_mem_reg[1][20]/P0001  ;
  input \u9_mem_reg[1][21]/P0001  ;
  input \u9_mem_reg[1][22]/P0001  ;
  input \u9_mem_reg[1][23]/P0001  ;
  input \u9_mem_reg[1][24]/P0001  ;
  input \u9_mem_reg[1][25]/P0001  ;
  input \u9_mem_reg[1][26]/P0001  ;
  input \u9_mem_reg[1][27]/P0001  ;
  input \u9_mem_reg[1][28]/P0001  ;
  input \u9_mem_reg[1][29]/P0001  ;
  input \u9_mem_reg[1][2]/P0001  ;
  input \u9_mem_reg[1][30]/P0001  ;
  input \u9_mem_reg[1][31]/P0001  ;
  input \u9_mem_reg[1][3]/P0001  ;
  input \u9_mem_reg[1][4]/P0001  ;
  input \u9_mem_reg[1][5]/P0001  ;
  input \u9_mem_reg[1][6]/P0001  ;
  input \u9_mem_reg[1][7]/P0001  ;
  input \u9_mem_reg[1][8]/P0001  ;
  input \u9_mem_reg[1][9]/P0001  ;
  input \u9_mem_reg[2][0]/P0001  ;
  input \u9_mem_reg[2][10]/P0001  ;
  input \u9_mem_reg[2][11]/P0001  ;
  input \u9_mem_reg[2][12]/P0001  ;
  input \u9_mem_reg[2][13]/P0001  ;
  input \u9_mem_reg[2][14]/P0001  ;
  input \u9_mem_reg[2][15]/P0001  ;
  input \u9_mem_reg[2][16]/P0001  ;
  input \u9_mem_reg[2][17]/P0001  ;
  input \u9_mem_reg[2][18]/P0001  ;
  input \u9_mem_reg[2][19]/P0001  ;
  input \u9_mem_reg[2][1]/P0001  ;
  input \u9_mem_reg[2][20]/P0001  ;
  input \u9_mem_reg[2][21]/P0001  ;
  input \u9_mem_reg[2][22]/P0001  ;
  input \u9_mem_reg[2][23]/P0001  ;
  input \u9_mem_reg[2][24]/P0001  ;
  input \u9_mem_reg[2][25]/P0001  ;
  input \u9_mem_reg[2][26]/P0001  ;
  input \u9_mem_reg[2][27]/P0001  ;
  input \u9_mem_reg[2][28]/P0001  ;
  input \u9_mem_reg[2][29]/P0001  ;
  input \u9_mem_reg[2][2]/P0001  ;
  input \u9_mem_reg[2][30]/P0001  ;
  input \u9_mem_reg[2][31]/P0001  ;
  input \u9_mem_reg[2][3]/P0001  ;
  input \u9_mem_reg[2][4]/P0001  ;
  input \u9_mem_reg[2][5]/P0001  ;
  input \u9_mem_reg[2][6]/P0001  ;
  input \u9_mem_reg[2][7]/P0001  ;
  input \u9_mem_reg[2][8]/P0001  ;
  input \u9_mem_reg[2][9]/P0001  ;
  input \u9_mem_reg[3][0]/P0001  ;
  input \u9_mem_reg[3][10]/P0001  ;
  input \u9_mem_reg[3][11]/P0001  ;
  input \u9_mem_reg[3][12]/P0001  ;
  input \u9_mem_reg[3][13]/P0001  ;
  input \u9_mem_reg[3][14]/P0001  ;
  input \u9_mem_reg[3][15]/P0001  ;
  input \u9_mem_reg[3][16]/P0001  ;
  input \u9_mem_reg[3][17]/P0001  ;
  input \u9_mem_reg[3][18]/P0001  ;
  input \u9_mem_reg[3][19]/P0001  ;
  input \u9_mem_reg[3][1]/P0001  ;
  input \u9_mem_reg[3][20]/P0001  ;
  input \u9_mem_reg[3][21]/P0001  ;
  input \u9_mem_reg[3][22]/P0001  ;
  input \u9_mem_reg[3][23]/P0001  ;
  input \u9_mem_reg[3][24]/P0001  ;
  input \u9_mem_reg[3][25]/P0001  ;
  input \u9_mem_reg[3][26]/P0001  ;
  input \u9_mem_reg[3][27]/P0001  ;
  input \u9_mem_reg[3][28]/P0001  ;
  input \u9_mem_reg[3][29]/P0001  ;
  input \u9_mem_reg[3][2]/P0001  ;
  input \u9_mem_reg[3][30]/P0001  ;
  input \u9_mem_reg[3][31]/P0001  ;
  input \u9_mem_reg[3][3]/P0001  ;
  input \u9_mem_reg[3][4]/P0001  ;
  input \u9_mem_reg[3][5]/P0001  ;
  input \u9_mem_reg[3][6]/P0001  ;
  input \u9_mem_reg[3][7]/P0001  ;
  input \u9_mem_reg[3][8]/P0001  ;
  input \u9_mem_reg[3][9]/P0001  ;
  input \u9_rp_reg[0]/P0001  ;
  input \u9_rp_reg[1]/P0001  ;
  input \u9_rp_reg[2]/P0001  ;
  input \u9_status_reg[0]/P0001  ;
  input \u9_status_reg[1]/P0001  ;
  input \u9_wp_reg[0]/NET0131  ;
  input \u9_wp_reg[1]/P0001  ;
  input \u9_wp_reg[2]/P0001  ;
  input \u9_wp_reg[3]/P0001  ;
  input \valid_s_reg/NET0131  ;
  input wb_ack_o_pad ;
  input \wb_addr_i[29]_pad  ;
  input \wb_addr_i[2]_pad  ;
  input \wb_addr_i[30]_pad  ;
  input \wb_addr_i[31]_pad  ;
  input \wb_addr_i[3]_pad  ;
  input \wb_addr_i[4]_pad  ;
  input \wb_addr_i[5]_pad  ;
  input \wb_addr_i[6]_pad  ;
  input wb_cyc_i_pad ;
  input wb_stb_i_pad ;
  input wb_we_i_pad ;
  output \_al_n1  ;
  output \g16/_0_  ;
  output \g23/_0_  ;
  output \g29500/_0_  ;
  output \g29503/_3_  ;
  output \g29505/_3_  ;
  output \g29507/_3_  ;
  output \g29509/_3_  ;
  output \g29511/_0_  ;
  output \g29513/_3_  ;
  output \g29515/_3_  ;
  output \g29517/_3_  ;
  output \g29519/_0_  ;
  output \g29522/_0_  ;
  output \g29524/_0_  ;
  output \g29526/_0_  ;
  output \g29528/_0_  ;
  output \g29530/_0_  ;
  output \g29532/_0_  ;
  output \g29534/_3_  ;
  output \g29536/_3_  ;
  output \g29538/_3_  ;
  output \g29540/_3_  ;
  output \g29542/_3_  ;
  output \g29544/_3_  ;
  output \g29546/_3_  ;
  output \g29548/_3_  ;
  output \g29550/_0_  ;
  output \g29552/_0_  ;
  output \g29554/_0_  ;
  output \g29556/_0_  ;
  output \g29558/_0_  ;
  output \g29560/_0_  ;
  output \g29562/_0_  ;
  output \g29564/_0_  ;
  output \g29566/_0_  ;
  output \g29568/_0_  ;
  output \g29570/_0_  ;
  output \g29572/_0_  ;
  output \g29574/_3_  ;
  output \g29576/_3_  ;
  output \g29578/_3_  ;
  output \g29580/_3_  ;
  output \g29582/_3_  ;
  output \g29584/_3_  ;
  output \g29586/_3_  ;
  output \g29588/_3_  ;
  output \g29590/_3_  ;
  output \g29592/_3_  ;
  output \g29594/_3_  ;
  output \g29596/_3_  ;
  output \g29598/_3_  ;
  output \g29600/_3_  ;
  output \g29602/_3_  ;
  output \g29604/_3_  ;
  output \g29606/_0_  ;
  output \g29608/_0_  ;
  output \g29610/_0_  ;
  output \g29612/_0_  ;
  output \g29614/_3_  ;
  output \g29616/_3_  ;
  output \g29618/_3_  ;
  output \g29620/_3_  ;
  output \g29622/_3_  ;
  output \g29624/_3_  ;
  output \g29626/_3_  ;
  output \g29628/_3_  ;
  output \g29630/_3_  ;
  output \g29632/_3_  ;
  output \g29634/_3_  ;
  output \g29636/_3_  ;
  output \g29638/_3_  ;
  output \g29640/_3_  ;
  output \g29642/_3_  ;
  output \g29644/_3_  ;
  output \g29646/_3_  ;
  output \g29648/_3_  ;
  output \g29650/_3_  ;
  output \g29652/_3_  ;
  output \g29654/_3_  ;
  output \g29656/_3_  ;
  output \g29658/_3_  ;
  output \g29660/_3_  ;
  output \g29662/_3_  ;
  output \g29664/_3_  ;
  output \g29666/_3_  ;
  output \g29668/_3_  ;
  output \g29670/_3_  ;
  output \g29672/_3_  ;
  output \g29674/_3_  ;
  output \g29676/_3_  ;
  output \g29678/_3_  ;
  output \g29680/_3_  ;
  output \g29682/_3_  ;
  output \g29684/_3_  ;
  output \g29686/_3_  ;
  output \g29688/_3_  ;
  output \g29690/_3_  ;
  output \g29692/_3_  ;
  output \g29694/_0_  ;
  output \g29696/_0_  ;
  output \g29698/_0_  ;
  output \g29700/_0_  ;
  output \g29702/_0_  ;
  output \g29704/_0_  ;
  output \g29706/_0_  ;
  output \g29708/_0_  ;
  output \g29710/_0_  ;
  output \g29712/_0_  ;
  output \g29714/_0_  ;
  output \g29716/_0_  ;
  output \g29718/_0_  ;
  output \g29720/_0_  ;
  output \g29722/_0_  ;
  output \g29724/_0_  ;
  output \g29726/_0_  ;
  output \g29728/_0_  ;
  output \g29730/_0_  ;
  output \g29732/_0_  ;
  output \g29734/_3_  ;
  output \g29736/_3_  ;
  output \g29738/_3_  ;
  output \g29740/_3_  ;
  output \g29742/_3_  ;
  output \g29744/_3_  ;
  output \g29746/_3_  ;
  output \g29748/_3_  ;
  output \g29750/_3_  ;
  output \g29752/_3_  ;
  output \g29754/_3_  ;
  output \g29756/_3_  ;
  output \g29758/_3_  ;
  output \g29760/_3_  ;
  output \g29762/_3_  ;
  output \g29764/_3_  ;
  output \g29766/_3_  ;
  output \g29768/_3_  ;
  output \g29770/_3_  ;
  output \g29772/_3_  ;
  output \g29774/_3_  ;
  output \g29776/_3_  ;
  output \g29778/_3_  ;
  output \g29780/_3_  ;
  output \g29782/_3_  ;
  output \g29784/_3_  ;
  output \g29786/_3_  ;
  output \g29788/_3_  ;
  output \g29790/_3_  ;
  output \g29792/_3_  ;
  output \g29794/_3_  ;
  output \g29796/_3_  ;
  output \g29798/_3_  ;
  output \g29800/_3_  ;
  output \g29802/_3_  ;
  output \g29804/_3_  ;
  output \g29806/_3_  ;
  output \g29808/_3_  ;
  output \g29810/_3_  ;
  output \g29812/_3_  ;
  output \g29814/_3_  ;
  output \g29816/_3_  ;
  output \g29818/_3_  ;
  output \g29820/_3_  ;
  output \g29822/_3_  ;
  output \g29824/_3_  ;
  output \g29826/_3_  ;
  output \g29828/_3_  ;
  output \g29830/_3_  ;
  output \g29832/_3_  ;
  output \g29834/_3_  ;
  output \g29836/_3_  ;
  output \g29838/_3_  ;
  output \g29840/_3_  ;
  output \g29842/_3_  ;
  output \g29844/_3_  ;
  output \g29846/_3_  ;
  output \g29848/_3_  ;
  output \g29850/_3_  ;
  output \g29852/_3_  ;
  output \g29854/_3_  ;
  output \g29856/_3_  ;
  output \g29858/_3_  ;
  output \g29860/_3_  ;
  output \g29862/_3_  ;
  output \g29864/_3_  ;
  output \g29866/_3_  ;
  output \g29868/_3_  ;
  output \g29870/_3_  ;
  output \g29872/_3_  ;
  output \g29874/_3_  ;
  output \g29876/_3_  ;
  output \g29878/_3_  ;
  output \g29880/_3_  ;
  output \g29904/_0_  ;
  output \g29905/_0_  ;
  output \g29906/_0_  ;
  output \g29907/_0_  ;
  output \g29908/_0_  ;
  output \g29909/_0_  ;
  output \g29914/_3_  ;
  output \g29952/_0_  ;
  output \g29953/_0_  ;
  output \g29954/_0_  ;
  output \g29955/_0_  ;
  output \g29956/_0_  ;
  output \g29957/_0_  ;
  output \g29975/_0_  ;
  output \g29976/_0_  ;
  output \g29977/_0_  ;
  output \g29978/_0_  ;
  output \g29979/_0_  ;
  output \g29980/_0_  ;
  output \g29989/_3_  ;
  output \g30020/_0_  ;
  output \g30021/_0_  ;
  output \g30045/_0_  ;
  output \g30046/_0_  ;
  output \g30047/_0_  ;
  output \g30048/_0_  ;
  output \g30049/_0_  ;
  output \g30050/_0_  ;
  output \g30051/_0_  ;
  output \g30052/_0_  ;
  output \g30053/_0_  ;
  output \g30054/_0_  ;
  output \g30062/_0_  ;
  output \g30063/_0_  ;
  output \g30064/_0_  ;
  output \g30065/_0_  ;
  output \g30066/_0_  ;
  output \g30067/_0_  ;
  output \g30068/_0_  ;
  output \g30069/_0_  ;
  output \g30070/_0_  ;
  output \g30071/_0_  ;
  output \g30072/_0_  ;
  output \g30073/_0_  ;
  output \g30074/_0_  ;
  output \g30075/_0_  ;
  output \g30136/_3_  ;
  output \g30707/_0_  ;
  output \g30708/_0_  ;
  output \g30711/_0_  ;
  output \g30714/_0_  ;
  output \g30715/_0_  ;
  output \g30720/_0_  ;
  output \g30725/_0_  ;
  output \g30741/_0_  ;
  output \g30742/_0_  ;
  output \g30743/_0_  ;
  output \g30744/_0_  ;
  output \g30745/_0_  ;
  output \g30746/_0_  ;
  output \g30747/_0_  ;
  output \g30748/_0_  ;
  output \g30749/_0_  ;
  output \g30750/_0_  ;
  output \g30751/_0_  ;
  output \g30752/_0_  ;
  output \g30789/_0_  ;
  output \g30790/_0_  ;
  output \g30791/_0_  ;
  output \g30792/_0_  ;
  output \g30793/_0_  ;
  output \g30794/_0_  ;
  output \g30795/_0_  ;
  output \g30796/_0_  ;
  output \g30797/_0_  ;
  output \g30798/_0_  ;
  output \g30799/_0_  ;
  output \g30800/_0_  ;
  output \g30801/_0_  ;
  output \g30802/_0_  ;
  output \g30803/_0_  ;
  output \g30804/_0_  ;
  output \g30805/_0_  ;
  output \g30806/_0_  ;
  output \g30807/_0_  ;
  output \g30808/_0_  ;
  output \g30809/_0_  ;
  output \g30810/_0_  ;
  output \g30811/_0_  ;
  output \g30812/_0_  ;
  output \g30813/_0_  ;
  output \g30814/_0_  ;
  output \g30815/_0_  ;
  output \g30816/_0_  ;
  output \g30817/_0_  ;
  output \g30818/_0_  ;
  output \g30819/_0_  ;
  output \g30820/_0_  ;
  output \g30821/_0_  ;
  output \g30822/_0_  ;
  output \g30823/_0_  ;
  output \g30824/_0_  ;
  output \g30825/_0_  ;
  output \g30826/_0_  ;
  output \g30827/_0_  ;
  output \g30828/_0_  ;
  output \g30829/_0_  ;
  output \g30830/_0_  ;
  output \g30831/_0_  ;
  output \g30832/_0_  ;
  output \g30833/_0_  ;
  output \g30834/_0_  ;
  output \g30835/_0_  ;
  output \g30836/_0_  ;
  output \g30837/_0_  ;
  output \g30838/_0_  ;
  output \g30839/_0_  ;
  output \g30840/_0_  ;
  output \g30841/_0_  ;
  output \g30842/_0_  ;
  output \g30843/_0_  ;
  output \g30844/_0_  ;
  output \g30845/_0_  ;
  output \g30846/_0_  ;
  output \g30847/_0_  ;
  output \g30848/_0_  ;
  output \g30849/_0_  ;
  output \g30850/_0_  ;
  output \g30851/_0_  ;
  output \g30852/_0_  ;
  output \g30853/_0_  ;
  output \g30854/_0_  ;
  output \g30855/_0_  ;
  output \g30856/_0_  ;
  output \g30857/_0_  ;
  output \g30858/_0_  ;
  output \g30859/_0_  ;
  output \g30860/_0_  ;
  output \g30861/_0_  ;
  output \g30862/_0_  ;
  output \g30863/_0_  ;
  output \g30864/_0_  ;
  output \g30865/_0_  ;
  output \g30866/_0_  ;
  output \g30867/_0_  ;
  output \g30868/_0_  ;
  output \g30869/_0_  ;
  output \g30870/_0_  ;
  output \g30871/_0_  ;
  output \g30872/_0_  ;
  output \g30873/_0_  ;
  output \g30874/_0_  ;
  output \g30875/_0_  ;
  output \g30876/_0_  ;
  output \g30877/_0_  ;
  output \g30878/_0_  ;
  output \g30879/_0_  ;
  output \g30880/_0_  ;
  output \g30881/_0_  ;
  output \g30882/_0_  ;
  output \g30883/_0_  ;
  output \g30884/_0_  ;
  output \g30885/_0_  ;
  output \g30886/_0_  ;
  output \g30887/_0_  ;
  output \g30888/_0_  ;
  output \g30889/_0_  ;
  output \g30890/_0_  ;
  output \g30891/_0_  ;
  output \g30892/_0_  ;
  output \g30893/_0_  ;
  output \g30894/_0_  ;
  output \g30895/_0_  ;
  output \g30896/_0_  ;
  output \g30897/_0_  ;
  output \g30898/_0_  ;
  output \g30899/_0_  ;
  output \g30900/_0_  ;
  output \g30901/_0_  ;
  output \g30902/_0_  ;
  output \g30906/_0_  ;
  output \g30907/_0_  ;
  output \g30908/_0_  ;
  output \g30909/_0_  ;
  output \g30910/_0_  ;
  output \g30911/_0_  ;
  output \g30918/_0_  ;
  output \g30919/_0_  ;
  output \g30920/_0_  ;
  output \g30921/_0_  ;
  output \g30922/_0_  ;
  output \g30923/_0_  ;
  output \g30924/_0_  ;
  output \g30925/_0_  ;
  output \g30926/_0_  ;
  output \g30946/_0_  ;
  output \g30947/_0_  ;
  output \g30948/_0_  ;
  output \g30949/_0_  ;
  output \g30950/_0_  ;
  output \g30951/_0_  ;
  output \g30952/_0_  ;
  output \g30953/_0_  ;
  output \g30954/_0_  ;
  output \g30955/_0_  ;
  output \g30956/_0_  ;
  output \g30957/_0_  ;
  output \g30958/_0_  ;
  output \g30959/_0_  ;
  output \g30960/_0_  ;
  output \g30961/_0_  ;
  output \g30962/_0_  ;
  output \g30963/_0_  ;
  output \g30964/_0_  ;
  output \g30965/_0_  ;
  output \g30966/_0_  ;
  output \g30967/_0_  ;
  output \g30968/_0_  ;
  output \g30969/_0_  ;
  output \g30970/_0_  ;
  output \g30971/_0_  ;
  output \g30972/_0_  ;
  output \g30973/_0_  ;
  output \g30974/_0_  ;
  output \g30975/_0_  ;
  output \g30976/_0_  ;
  output \g30977/_0_  ;
  output \g30978/_0_  ;
  output \g30979/_0_  ;
  output \g30980/_0_  ;
  output \g30981/_0_  ;
  output \g30982/_0_  ;
  output \g30983/_0_  ;
  output \g30984/_0_  ;
  output \g30985/_0_  ;
  output \g30986/_0_  ;
  output \g30987/_0_  ;
  output \g30988/_0_  ;
  output \g30989/_0_  ;
  output \g30990/_0_  ;
  output \g30991/_0_  ;
  output \g30992/_0_  ;
  output \g30993/_0_  ;
  output \g30994/_0_  ;
  output \g30995/_0_  ;
  output \g30996/_0_  ;
  output \g30997/_0_  ;
  output \g30998/_0_  ;
  output \g30999/_0_  ;
  output \g31000/_0_  ;
  output \g31001/_0_  ;
  output \g31002/_0_  ;
  output \g31003/_0_  ;
  output \g31004/_0_  ;
  output \g31005/_0_  ;
  output \g31006/_0_  ;
  output \g31007/_0_  ;
  output \g31008/_0_  ;
  output \g31009/_0_  ;
  output \g31010/_0_  ;
  output \g31011/_0_  ;
  output \g31012/_0_  ;
  output \g31013/_0_  ;
  output \g31014/_0_  ;
  output \g31015/_0_  ;
  output \g31016/_0_  ;
  output \g31017/_0_  ;
  output \g31018/_0_  ;
  output \g31019/_0_  ;
  output \g31020/_0_  ;
  output \g31021/_0_  ;
  output \g31022/_0_  ;
  output \g31023/_0_  ;
  output \g31024/_0_  ;
  output \g31025/_0_  ;
  output \g31026/_0_  ;
  output \g31027/_0_  ;
  output \g31028/_0_  ;
  output \g31029/_0_  ;
  output \g31030/_0_  ;
  output \g31031/_0_  ;
  output \g31032/_0_  ;
  output \g31033/_0_  ;
  output \g31034/_0_  ;
  output \g31035/_0_  ;
  output \g31036/_0_  ;
  output \g31037/_0_  ;
  output \g31038/_0_  ;
  output \g31039/_0_  ;
  output \g31040/_0_  ;
  output \g31041/_0_  ;
  output \g31042/_0_  ;
  output \g31043/_0_  ;
  output \g31044/_0_  ;
  output \g31045/_0_  ;
  output \g31046/_0_  ;
  output \g31047/_0_  ;
  output \g31048/_0_  ;
  output \g31049/_0_  ;
  output \g31050/_0_  ;
  output \g31051/_0_  ;
  output \g31052/_0_  ;
  output \g31053/_0_  ;
  output \g31054/_0_  ;
  output \g31055/_0_  ;
  output \g31056/_0_  ;
  output \g31057/_0_  ;
  output \g31058/_0_  ;
  output \g31059/_0_  ;
  output \g31060/_0_  ;
  output \g31061/_0_  ;
  output \g31062/_0_  ;
  output \g31063/_0_  ;
  output \g31064/_0_  ;
  output \g31065/_0_  ;
  output \g31066/_0_  ;
  output \g31067/_0_  ;
  output \g31068/_0_  ;
  output \g31069/_0_  ;
  output \g31070/_0_  ;
  output \g31071/_0_  ;
  output \g31072/_0_  ;
  output \g31073/_0_  ;
  output \g31074/_0_  ;
  output \g31075/_0_  ;
  output \g31076/_0_  ;
  output \g31077/_0_  ;
  output \g31084/u3_syn_4  ;
  output \g31085/u3_syn_4  ;
  output \g31096/u3_syn_4  ;
  output \g31115/u3_syn_4  ;
  output \g31136/u3_syn_4  ;
  output \g31158/u3_syn_4  ;
  output \g31176/u3_syn_4  ;
  output \g31193/u3_syn_4  ;
  output \g31195/u3_syn_4  ;
  output \g31247/u3_syn_4  ;
  output \g31280/u3_syn_4  ;
  output \g31285/u3_syn_4  ;
  output \g31568/_0_  ;
  output \g31631/_0_  ;
  output \g31672/_0_  ;
  output \g31731/_0_  ;
  output \g31732/_0_  ;
  output \g31742/_2_  ;
  output \g31744/_2_  ;
  output \g31746/_2_  ;
  output \g31748/_2_  ;
  output \g31751/_2_  ;
  output \g31754/_2_  ;
  output \g31756/_2_  ;
  output \g31758/_2_  ;
  output \g31760/_2_  ;
  output \g31761/_0_  ;
  output \g31789/_0_  ;
  output \g31807/_3_  ;
  output \g31825/_3_  ;
  output \g32607/_0_  ;
  output \g32608/_0_  ;
  output \g32609/_0_  ;
  output \g32610/_0_  ;
  output \g32611/_0_  ;
  output \g32612/_0_  ;
  output \g32613/_0_  ;
  output \g32614/_0_  ;
  output \g32615/_0_  ;
  output \g32616/_0_  ;
  output \g32617/_0_  ;
  output \g32618/_0_  ;
  output \g32645/_0__syn_2  ;
  output \g32687/_0__syn_2  ;
  output \g32749/_0__syn_2  ;
  output \g32757/_0_  ;
  output \g32758/_0_  ;
  output \g32759/_0_  ;
  output \g32760/_0_  ;
  output \g32761/_0_  ;
  output \g32762/_0_  ;
  output \g32763/_0_  ;
  output \g32764/_0_  ;
  output \g32765/_0_  ;
  output \g32769/_0_  ;
  output \g32835/_1_  ;
  output \g32839/_0_  ;
  output \g32844/_0_  ;
  output \g32901/_1_  ;
  output \g32902/_0_  ;
  output \g32963/_1_  ;
  output \g32972/_0_  ;
  output \g32977/_0_  ;
  output \g32979/_0_  ;
  output \g32980/_0_  ;
  output \g32981/_0_  ;
  output \g32982/_0_  ;
  output \g32983/_0_  ;
  output \g32987/_0_  ;
  output \g33018/_0_  ;
  output \g33019/_0_  ;
  output \g33088/_0_  ;
  output \g33261/_0_  ;
  output \g33264/_0_  ;
  output \g33275/_0_  ;
  output \g33276/_0_  ;
  output \g33277/_0_  ;
  output \g33371/_0_  ;
  output \g33382/_0_  ;
  output \g33401/_0_  ;
  output \g33402/_0_  ;
  output \g33403/_0_  ;
  output \g33404/_0_  ;
  output \g33405/_0_  ;
  output \g33406/_0_  ;
  output \g33407/_0_  ;
  output \g33408/_0_  ;
  output \g33409/_0_  ;
  output \g33410/_0_  ;
  output \g33411/_0_  ;
  output \g33412/_0_  ;
  output \g33413/_0_  ;
  output \g33414/_0_  ;
  output \g33415/_0_  ;
  output \g33416/_0_  ;
  output \g33417/_0_  ;
  output \g33418/_0_  ;
  output \g33419/_0_  ;
  output \g33420/_0_  ;
  output \g33421/_0_  ;
  output \g33422/_0_  ;
  output \g33423/_0_  ;
  output \g33424/_0_  ;
  output \g33425/_0_  ;
  output \g33426/_0_  ;
  output \g33427/_0_  ;
  output \g33428/_0_  ;
  output \g33429/_0_  ;
  output \g33430/_0_  ;
  output \g33431/_0_  ;
  output \g33432/_0_  ;
  output \g33433/_0_  ;
  output \g33434/_0_  ;
  output \g33435/_0_  ;
  output \g33436/_0_  ;
  output \g33437/_0_  ;
  output \g33438/_0_  ;
  output \g33439/_0_  ;
  output \g33440/_0_  ;
  output \g33441/_0_  ;
  output \g33442/_0_  ;
  output \g33443/_0_  ;
  output \g33444/_0_  ;
  output \g33445/_0_  ;
  output \g33446/_0_  ;
  output \g33447/_0_  ;
  output \g33448/_0_  ;
  output \g33449/_0_  ;
  output \g33450/_0_  ;
  output \g33451/_0_  ;
  output \g33452/_0_  ;
  output \g33453/_0_  ;
  output \g33454/_0_  ;
  output \g33455/_0_  ;
  output \g33456/_0_  ;
  output \g33457/_0_  ;
  output \g33458/_0_  ;
  output \g33459/_0_  ;
  output \g33460/_0_  ;
  output \g33461/_0_  ;
  output \g33462/_0_  ;
  output \g33463/_0_  ;
  output \g33464/_0_  ;
  output \g33465/_0_  ;
  output \g33466/_0_  ;
  output \g33467/_0_  ;
  output \g33468/_0_  ;
  output \g33469/_0_  ;
  output \g33470/_0_  ;
  output \g33471/_0_  ;
  output \g33472/_0_  ;
  output \g33473/_0_  ;
  output \g33474/_0_  ;
  output \g33475/_0_  ;
  output \g33476/_0_  ;
  output \g33477/_0_  ;
  output \g33478/_0_  ;
  output \g33479/_0_  ;
  output \g33480/_0_  ;
  output \g33481/_0_  ;
  output \g33482/_0_  ;
  output \g33483/_0_  ;
  output \g33484/_0_  ;
  output \g33485/_0_  ;
  output \g33486/_0_  ;
  output \g33487/_0_  ;
  output \g33488/_0_  ;
  output \g33489/_0_  ;
  output \g33490/_0_  ;
  output \g33491/_0_  ;
  output \g33492/_0_  ;
  output \g33493/_0_  ;
  output \g33494/_0_  ;
  output \g33495/_0_  ;
  output \g33496/_0_  ;
  output \g33497/_0_  ;
  output \g33498/_0_  ;
  output \g33499/_0_  ;
  output \g33500/_0_  ;
  output \g33501/_0_  ;
  output \g33502/_0_  ;
  output \g33503/_0_  ;
  output \g33504/_0_  ;
  output \g33505/_0_  ;
  output \g33506/_0_  ;
  output \g33507/_0_  ;
  output \g33508/_0_  ;
  output \g33509/_0_  ;
  output \g33510/_0_  ;
  output \g33511/_0_  ;
  output \g33512/_0_  ;
  output \g33513/_0_  ;
  output \g33514/_0_  ;
  output \g33515/_0_  ;
  output \g33516/_0_  ;
  output \g33517/_0_  ;
  output \g33518/_0_  ;
  output \g33519/_0_  ;
  output \g33520/_0_  ;
  output \g33521/_0_  ;
  output \g33522/_0_  ;
  output \g33523/_0_  ;
  output \g33524/_0_  ;
  output \g33525/_0_  ;
  output \g33526/_0_  ;
  output \g33527/_0_  ;
  output \g33528/_0_  ;
  output \g33529/_0_  ;
  output \g33530/_0_  ;
  output \g33531/_0_  ;
  output \g33532/_0_  ;
  output \g33533/_0_  ;
  output \g33534/_0_  ;
  output \g33535/_0_  ;
  output \g33536/_0_  ;
  output \g33537/_0_  ;
  output \g33538/_0_  ;
  output \g33539/_0_  ;
  output \g33540/_0_  ;
  output \g33541/_0_  ;
  output \g33542/_0_  ;
  output \g33543/_0_  ;
  output \g33544/_0_  ;
  output \g33545/_0_  ;
  output \g33546/_0_  ;
  output \g33547/_0_  ;
  output \g33548/_0_  ;
  output \g33549/_0_  ;
  output \g33550/_0_  ;
  output \g33551/_0_  ;
  output \g33552/_0_  ;
  output \g33553/_0_  ;
  output \g33554/_0_  ;
  output \g33555/_0_  ;
  output \g33556/_0_  ;
  output \g33557/_0_  ;
  output \g33558/_0_  ;
  output \g33559/_0_  ;
  output \g33560/_0_  ;
  output \g33561/_0_  ;
  output \g33562/_0_  ;
  output \g33563/_0_  ;
  output \g33564/_0_  ;
  output \g33565/_0_  ;
  output \g33566/_0_  ;
  output \g33567/_0_  ;
  output \g33568/_0_  ;
  output \g33569/_0_  ;
  output \g33570/_0_  ;
  output \g33571/_0_  ;
  output \g33572/_0_  ;
  output \g33573/_0_  ;
  output \g33574/_0_  ;
  output \g33575/_0_  ;
  output \g33576/_0_  ;
  output \g33577/_0_  ;
  output \g33578/_0_  ;
  output \g33579/_0_  ;
  output \g33580/_0_  ;
  output \g33581/_0_  ;
  output \g33582/_0_  ;
  output \g33583/_0_  ;
  output \g33584/_0_  ;
  output \g33585/_0_  ;
  output \g33586/_0_  ;
  output \g33587/_0_  ;
  output \g33588/_0_  ;
  output \g33589/_0_  ;
  output \g33590/_0_  ;
  output \g33591/_0_  ;
  output \g33592/_0_  ;
  output \g33593/_0_  ;
  output \g33594/_0_  ;
  output \g33595/_0_  ;
  output \g33596/_0_  ;
  output \g33597/_0_  ;
  output \g33598/_0_  ;
  output \g33599/_0_  ;
  output \g33600/_0_  ;
  output \g33601/_0_  ;
  output \g33602/_0_  ;
  output \g33603/_0_  ;
  output \g33604/_0_  ;
  output \g33605/_0_  ;
  output \g33606/_0_  ;
  output \g33607/_0_  ;
  output \g33608/_0_  ;
  output \g33609/_0_  ;
  output \g33610/_0_  ;
  output \g33611/_0_  ;
  output \g33612/_0_  ;
  output \g33613/_0_  ;
  output \g33614/_0_  ;
  output \g33615/_0_  ;
  output \g33616/_0_  ;
  output \g33617/_0_  ;
  output \g33618/_0_  ;
  output \g33619/_0_  ;
  output \g33620/_0_  ;
  output \g33621/_0_  ;
  output \g33622/_0_  ;
  output \g33623/_0_  ;
  output \g33624/_0_  ;
  output \g33625/_0_  ;
  output \g33626/_0_  ;
  output \g33627/_0_  ;
  output \g33628/_0_  ;
  output \g33629/_0_  ;
  output \g33630/_0_  ;
  output \g33631/_0_  ;
  output \g33632/_0_  ;
  output \g33633/_0_  ;
  output \g33634/_0_  ;
  output \g33635/_0_  ;
  output \g33636/_0_  ;
  output \g33637/_0_  ;
  output \g33638/_0_  ;
  output \g33639/_0_  ;
  output \g33640/_0_  ;
  output \g33641/_0_  ;
  output \g33642/_0_  ;
  output \g33643/_0_  ;
  output \g33644/_0_  ;
  output \g33645/_0_  ;
  output \g33646/_0_  ;
  output \g33647/_0_  ;
  output \g33648/_0_  ;
  output \g33649/_0_  ;
  output \g33650/_0_  ;
  output \g33651/_0_  ;
  output \g33652/_0_  ;
  output \g33653/_0_  ;
  output \g33654/_0_  ;
  output \g33655/_0_  ;
  output \g33656/_0_  ;
  output \g33657/_0_  ;
  output \g33658/_0_  ;
  output \g33659/_0_  ;
  output \g33660/_0_  ;
  output \g33661/_0_  ;
  output \g33662/_0_  ;
  output \g33663/_0_  ;
  output \g33664/_0_  ;
  output \g33665/_0_  ;
  output \g33666/_0_  ;
  output \g33667/_0_  ;
  output \g33668/_0_  ;
  output \g33669/_0_  ;
  output \g33670/_0_  ;
  output \g33671/_0_  ;
  output \g33672/_0_  ;
  output \g33673/_0_  ;
  output \g33674/_0_  ;
  output \g33675/_0_  ;
  output \g33676/_0_  ;
  output \g33677/_0_  ;
  output \g33678/_0_  ;
  output \g33679/_0_  ;
  output \g33680/_0_  ;
  output \g33681/_0_  ;
  output \g33682/_0_  ;
  output \g33683/_0_  ;
  output \g33684/_0_  ;
  output \g33685/_0_  ;
  output \g33686/_0_  ;
  output \g33687/_0_  ;
  output \g33688/_0_  ;
  output \g33689/_0_  ;
  output \g33690/_0_  ;
  output \g33691/_0_  ;
  output \g33692/_0_  ;
  output \g33693/_0_  ;
  output \g33694/_0_  ;
  output \g33695/_0_  ;
  output \g33696/_0_  ;
  output \g33697/_0_  ;
  output \g33698/_0_  ;
  output \g33699/_0_  ;
  output \g33700/_0_  ;
  output \g33701/_0_  ;
  output \g33702/_0_  ;
  output \g33703/_0_  ;
  output \g33704/_0_  ;
  output \g33705/_0_  ;
  output \g33706/_0_  ;
  output \g33707/_0_  ;
  output \g33708/_0_  ;
  output \g33709/_0_  ;
  output \g33710/_0_  ;
  output \g33711/_0_  ;
  output \g33712/_0_  ;
  output \g33713/_0_  ;
  output \g33714/_0_  ;
  output \g33715/_0_  ;
  output \g33716/_0_  ;
  output \g33717/_0_  ;
  output \g33718/_0_  ;
  output \g33719/_0_  ;
  output \g33720/_0_  ;
  output \g33721/_0_  ;
  output \g33722/_0_  ;
  output \g33723/_0_  ;
  output \g33724/_0_  ;
  output \g33725/_0_  ;
  output \g33726/_0_  ;
  output \g33727/_0_  ;
  output \g33728/_0_  ;
  output \g33729/_0_  ;
  output \g33730/_0_  ;
  output \g33731/_0_  ;
  output \g33732/_0_  ;
  output \g33733/_0_  ;
  output \g33734/_0_  ;
  output \g33735/_0_  ;
  output \g33736/_0_  ;
  output \g33737/_0_  ;
  output \g33738/_0_  ;
  output \g33739/_0_  ;
  output \g33740/_0_  ;
  output \g33741/_0_  ;
  output \g33742/_0_  ;
  output \g33743/_0_  ;
  output \g33744/_0_  ;
  output \g33745/_0_  ;
  output \g33746/_0_  ;
  output \g33747/_0_  ;
  output \g33748/_0_  ;
  output \g33749/_0_  ;
  output \g33750/_0_  ;
  output \g33751/_0_  ;
  output \g33752/_0_  ;
  output \g33753/_0_  ;
  output \g33754/_0_  ;
  output \g33755/_0_  ;
  output \g33756/_0_  ;
  output \g33757/_0_  ;
  output \g33758/_0_  ;
  output \g33759/_0_  ;
  output \g33760/_0_  ;
  output \g33761/_0_  ;
  output \g33762/_0_  ;
  output \g33763/_0_  ;
  output \g33764/_0_  ;
  output \g33765/_0_  ;
  output \g33766/_0_  ;
  output \g33767/_0_  ;
  output \g33768/_0_  ;
  output \g33769/_0_  ;
  output \g33770/_0_  ;
  output \g33771/_0_  ;
  output \g33772/_0_  ;
  output \g33773/_0_  ;
  output \g33774/_0_  ;
  output \g33775/_0_  ;
  output \g33776/_0_  ;
  output \g33777/_0_  ;
  output \g33778/_0_  ;
  output \g33779/_0_  ;
  output \g33780/_0_  ;
  output \g33781/_0_  ;
  output \g33782/_0_  ;
  output \g33783/_0_  ;
  output \g33784/_0_  ;
  output \g33785/_0_  ;
  output \g33786/_0_  ;
  output \g33787/_0_  ;
  output \g33788/_0_  ;
  output \g33789/_0_  ;
  output \g33790/_0_  ;
  output \g33791/_0_  ;
  output \g33792/_0_  ;
  output \g33793/_0_  ;
  output \g33794/_0_  ;
  output \g33795/_0_  ;
  output \g33796/_0_  ;
  output \g33797/_0_  ;
  output \g33798/_0_  ;
  output \g33799/_0_  ;
  output \g33800/_0_  ;
  output \g33801/_0_  ;
  output \g33802/_0_  ;
  output \g33803/_0_  ;
  output \g33804/_0_  ;
  output \g33805/_0_  ;
  output \g33806/_0_  ;
  output \g33807/_0_  ;
  output \g33808/_0_  ;
  output \g33809/_0_  ;
  output \g33810/_0_  ;
  output \g33811/_0_  ;
  output \g33812/_0_  ;
  output \g33813/_0_  ;
  output \g33814/_0_  ;
  output \g33815/_0_  ;
  output \g33816/_0_  ;
  output \g33817/_0_  ;
  output \g33818/_0_  ;
  output \g33819/_0_  ;
  output \g33820/_0_  ;
  output \g33821/_0_  ;
  output \g33822/_0_  ;
  output \g33823/_0_  ;
  output \g33824/_0_  ;
  output \g33825/_0_  ;
  output \g33826/_0_  ;
  output \g33827/_0_  ;
  output \g33828/_0_  ;
  output \g33829/_0_  ;
  output \g33830/_0_  ;
  output \g33831/_0_  ;
  output \g33832/_0_  ;
  output \g33833/_0_  ;
  output \g33834/_0_  ;
  output \g33835/_0_  ;
  output \g33836/_0_  ;
  output \g33837/_0_  ;
  output \g33838/_0_  ;
  output \g33839/_0_  ;
  output \g33840/_0_  ;
  output \g33841/_0_  ;
  output \g33842/_0_  ;
  output \g33843/_0_  ;
  output \g33844/_0_  ;
  output \g33845/_0_  ;
  output \g33846/_0_  ;
  output \g33847/_0_  ;
  output \g33848/_0_  ;
  output \g33849/_0_  ;
  output \g33850/_0_  ;
  output \g33851/_0_  ;
  output \g33852/_0_  ;
  output \g33853/_0_  ;
  output \g33854/_0_  ;
  output \g33855/_0_  ;
  output \g33856/_0_  ;
  output \g33857/_0_  ;
  output \g33858/_0_  ;
  output \g33859/_0_  ;
  output \g33860/_0_  ;
  output \g33861/_0_  ;
  output \g33862/_0_  ;
  output \g33863/_0_  ;
  output \g33864/_0_  ;
  output \g33865/_0_  ;
  output \g33866/_0_  ;
  output \g33867/_0_  ;
  output \g33868/_0_  ;
  output \g33869/_0_  ;
  output \g33870/_0_  ;
  output \g33871/_0_  ;
  output \g33872/_0_  ;
  output \g33873/_0_  ;
  output \g33874/_0_  ;
  output \g33875/_0_  ;
  output \g33876/_0_  ;
  output \g33877/_0_  ;
  output \g33878/_0_  ;
  output \g33879/_0_  ;
  output \g33880/_0_  ;
  output \g33881/_0_  ;
  output \g33882/_0_  ;
  output \g33883/_0_  ;
  output \g33884/_0_  ;
  output \g33885/_0_  ;
  output \g33886/_0_  ;
  output \g33887/_0_  ;
  output \g33888/_0_  ;
  output \g33889/_0_  ;
  output \g33890/_0_  ;
  output \g33891/_0_  ;
  output \g33892/_0_  ;
  output \g33893/_0_  ;
  output \g33894/_0_  ;
  output \g33895/_0_  ;
  output \g33896/_0_  ;
  output \g33897/_0_  ;
  output \g33898/_0_  ;
  output \g33899/_0_  ;
  output \g33900/_0_  ;
  output \g33901/_0_  ;
  output \g33902/_0_  ;
  output \g33903/_0_  ;
  output \g33904/_0_  ;
  output \g33905/_0_  ;
  output \g33906/_0_  ;
  output \g33907/_0_  ;
  output \g33908/_0_  ;
  output \g33909/_0_  ;
  output \g33910/_0_  ;
  output \g33911/_0_  ;
  output \g33912/_0_  ;
  output \g33913/_0_  ;
  output \g33914/_0_  ;
  output \g33915/_0_  ;
  output \g33916/_0_  ;
  output \g33917/_0_  ;
  output \g33918/_0_  ;
  output \g33919/_0_  ;
  output \g33920/_0_  ;
  output \g33921/_0_  ;
  output \g33922/_0_  ;
  output \g33923/_0_  ;
  output \g33924/_0_  ;
  output \g33925/_0_  ;
  output \g33926/_0_  ;
  output \g33927/_0_  ;
  output \g33928/_0_  ;
  output \g33929/_0_  ;
  output \g33930/_0_  ;
  output \g33931/_0_  ;
  output \g33932/_0_  ;
  output \g33933/_0_  ;
  output \g33934/_0_  ;
  output \g33935/_0_  ;
  output \g33936/_0_  ;
  output \g33937/_0_  ;
  output \g33938/_0_  ;
  output \g33939/_0_  ;
  output \g33940/_0_  ;
  output \g33941/_0_  ;
  output \g33942/_0_  ;
  output \g33943/_0_  ;
  output \g33944/_0_  ;
  output \g33945/_0_  ;
  output \g33946/_0_  ;
  output \g33947/_0_  ;
  output \g33948/_0_  ;
  output \g33949/_0_  ;
  output \g33950/_0_  ;
  output \g33951/_0_  ;
  output \g33952/_0_  ;
  output \g33953/_0_  ;
  output \g33954/_0_  ;
  output \g33955/_0_  ;
  output \g33956/_0_  ;
  output \g33957/_0_  ;
  output \g33958/_0_  ;
  output \g33959/_0_  ;
  output \g33960/_0_  ;
  output \g33961/_0_  ;
  output \g33962/_0_  ;
  output \g33963/_0_  ;
  output \g33964/_0_  ;
  output \g33965/_0_  ;
  output \g33966/_0_  ;
  output \g33967/_0_  ;
  output \g33968/_0_  ;
  output \g33969/_0_  ;
  output \g33970/_0_  ;
  output \g33971/_0_  ;
  output \g33972/_0_  ;
  output \g33973/_0_  ;
  output \g33974/_0_  ;
  output \g33975/_0_  ;
  output \g33976/_0_  ;
  output \g33977/u3_syn_4  ;
  output \g33981/u3_syn_4  ;
  output \g34014/u3_syn_4  ;
  output \g34047/u3_syn_4  ;
  output \g34084/u3_syn_4  ;
  output \g34123/u3_syn_4  ;
  output \g34306/_0_  ;
  output \g34316/_0_  ;
  output \g34324/_0_  ;
  output \g34326/_0_  ;
  output \g34328/_0_  ;
  output \g34331/_0_  ;
  output \g34333/_0_  ;
  output \g34344/_0_  ;
  output \g34347/_0_  ;
  output \g34351/_0_  ;
  output \g34361/_0_  ;
  output \g34368/_0_  ;
  output \g34377/_0_  ;
  output \g34385/_0_  ;
  output \g34393/_0_  ;
  output \g34414/_1_  ;
  output \g34451/_1_  ;
  output \g34476/_1_  ;
  output \g34487/_0_  ;
  output \g34490/_1_  ;
  output \g34715/_0_  ;
  output \g34878/_0_  ;
  output \g34882/_0_  ;
  output \g34883/_0_  ;
  output \g34893/_0_  ;
  output \g34896/_0_  ;
  output \g34898/_0_  ;
  output \g34899/_0_  ;
  output \g34916/_3_  ;
  output \g35264/_0_  ;
  output \g35265/_0_  ;
  output \g35266/_0_  ;
  output \g35267/_0_  ;
  output \g35268/_0_  ;
  output \g35269/_0_  ;
  output \g35270/_0_  ;
  output \g35271/_0_  ;
  output \g35272/_0_  ;
  output \g35273/_0_  ;
  output \g35274/_0_  ;
  output \g35275/_0_  ;
  output \g35276/_0_  ;
  output \g35277/_0_  ;
  output \g35278/_0_  ;
  output \g35279/_0_  ;
  output \g35283/_0_  ;
  output \g35287/_0_  ;
  output \g35294/_0_  ;
  output \g35300/_0_  ;
  output \g35304/_0_  ;
  output \g35308/_0_  ;
  output \g35312/_0_  ;
  output \g35316/_0_  ;
  output \g35318/_0_  ;
  output \g35326/_0_  ;
  output \g35334/_0_  ;
  output \g35336/_0_  ;
  output \g35337/_0_  ;
  output \g35338/_0_  ;
  output \g35357/_0_  ;
  output \g35358/_0_  ;
  output \g35359/_0_  ;
  output \g35419/_0_  ;
  output \g35438/_0_  ;
  output \g35439/_0_  ;
  output \g35440/_0_  ;
  output \g35441/_0_  ;
  output \g35442/_0_  ;
  output \g35444/_0_  ;
  output \g35445/_0_  ;
  output \g35446/_0_  ;
  output \g35447/_0_  ;
  output \g35448/_0_  ;
  output \g35449/_0_  ;
  output \g35450/_0_  ;
  output \g35451/_0_  ;
  output \g35452/_0_  ;
  output \g35463/_0_  ;
  output \g35464/_0_  ;
  output \g35466/_0_  ;
  output \g35485/_2_  ;
  output \g35495/_0_  ;
  output \g35496/_0_  ;
  output \g35499/_0_  ;
  output \g35500/_0_  ;
  output \g35501/_0_  ;
  output \g35502/_0_  ;
  output \g35563/_0_  ;
  output \g35633/_0_  ;
  output \g35717/_0_  ;
  output \g35718/_0_  ;
  output \g35719/_0_  ;
  output \g35809/_0_  ;
  output \g35810/_0_  ;
  output \g35811/_0_  ;
  output \g35812/_0_  ;
  output \g35813/_0_  ;
  output \g35814/_0_  ;
  output \g35815/_0_  ;
  output \g35816/_0_  ;
  output \g35817/_0_  ;
  output \g35818/_0_  ;
  output \g35819/_0_  ;
  output \g35820/_0_  ;
  output \g35821/_0_  ;
  output \g35822/_0_  ;
  output \g35823/_0_  ;
  output \g35824/_0_  ;
  output \g35825/_0_  ;
  output \g35826/_0_  ;
  output \g35827/_0_  ;
  output \g35830/_0_  ;
  output \g35833/_0_  ;
  output \g35835/_0_  ;
  output \g35836/_0_  ;
  output \g35837/_0_  ;
  output \g35839/_0_  ;
  output \g35840/_0_  ;
  output \g35841/_0_  ;
  output \g35843/_0_  ;
  output \g35844/_0_  ;
  output \g35845/_0_  ;
  output \g35853/_0_  ;
  output \g35854/_0_  ;
  output \g35855/_0_  ;
  output \g35856/_0_  ;
  output \g36306/_0_  ;
  output \g36414/_0_  ;
  output \g36415/_0_  ;
  output \g36449/_0_  ;
  output \g36550/_0_  ;
  output \g36551/_0_  ;
  output \g36553/_0_  ;
  output \g36560/_0_  ;
  output \g36562/_3_  ;
  output \g36563/_0_  ;
  output \g36612/_0_  ;
  output \g36614/_2_  ;
  output \g36695/_0_  ;
  output \g36784/_0_  ;
  output \g36785/_0_  ;
  output \g36786/_0_  ;
  output \g36787/_0_  ;
  output \g36788/_0_  ;
  output \g36789/_0_  ;
  output \g36790/_0_  ;
  output \g36791/_0_  ;
  output \g36792/_0_  ;
  output \g36793/_0_  ;
  output \g36794/_0_  ;
  output \g36796/_0_  ;
  output \g36797/_0_  ;
  output \g36798/_0_  ;
  output \g36799/_0_  ;
  output \g36800/_0_  ;
  output \g36801/_0_  ;
  output \g36802/_0_  ;
  output \g36803/_0_  ;
  output \g36804/_0_  ;
  output \g36805/_0_  ;
  output \g36806/_0_  ;
  output \g36807/_0_  ;
  output \g36808/_0_  ;
  output \g36809/_0_  ;
  output \g36810/_0_  ;
  output \g36811/_0_  ;
  output \g36813/_0_  ;
  output \g36814/_0_  ;
  output \g36815/_0_  ;
  output \g36820/_0_  ;
  output \g36825/_0_  ;
  output \g36832/_0_  ;
  output \g36846/_0_  ;
  output \g36855/_0_  ;
  output \g36857/_0_  ;
  output \g36859/_0_  ;
  output \g36860/_0_  ;
  output \g36861/_0_  ;
  output \g36862/_0_  ;
  output \g36863/_0_  ;
  output \g36864/_0_  ;
  output \g36867/_0_  ;
  output \g36870/_0_  ;
  output \g36871/_0_  ;
  output \g36877/_0_  ;
  output \g36879/_0_  ;
  output \g36892/_0_  ;
  output \g36893/_0_  ;
  output \g36901/_0_  ;
  output \g36909/_0_  ;
  output \g36914/_0_  ;
  output \g36919/_0_  ;
  output \g36922/_0_  ;
  output \g36923/_0_  ;
  output \g36927/_0_  ;
  output \g36930/_0_  ;
  output \g36931/_0_  ;
  output \g36933/_0_  ;
  output \g36934/_0_  ;
  output \g36935/_0_  ;
  output \g36936/_0_  ;
  output \g36937/_0_  ;
  output \g36938/_0_  ;
  output \g36939/_0_  ;
  output \g36940/_0_  ;
  output \g36941/_0_  ;
  output \g36943/_0_  ;
  output \g36944/_0_  ;
  output \g36945/_0_  ;
  output \g36946/_0_  ;
  output \g36947/_0_  ;
  output \g36948/_0_  ;
  output \g36949/_0_  ;
  output \g36950/_0_  ;
  output \g36951/_0_  ;
  output \g36952/_0_  ;
  output \g36953/_0_  ;
  output \g36954/_0_  ;
  output \g36957/_0_  ;
  output \g36958/_0_  ;
  output \g36959/_0_  ;
  output \g36960/_0_  ;
  output \g36961/_0_  ;
  output \g36962/_0_  ;
  output \g36963/_0_  ;
  output \g36970/_0_  ;
  output \g36977/_0_  ;
  output \g36986/_0_  ;
  output \g36991/_0_  ;
  output \g36994/_0_  ;
  output \g37015/_0_  ;
  output \g37057/_0_  ;
  output \g37073/_0_  ;
  output \g37128/_0_  ;
  output \g37129/_0_  ;
  output \g37138/_0_  ;
  output \g37139/_0_  ;
  output \g37140/_0_  ;
  output \g37141/_0_  ;
  output \g37142/_0_  ;
  output \g37143/_0_  ;
  output \g37144/_0_  ;
  output \g37145/_0_  ;
  output \g37146/_0_  ;
  output \g37147/_0_  ;
  output \g37148/_0_  ;
  output \g37149/_0_  ;
  output \g37150/_0_  ;
  output \g37151/_0_  ;
  output \g37152/_0_  ;
  output \g37153/_0_  ;
  output \g37154/_0_  ;
  output \g37155/_0_  ;
  output \g37156/_0_  ;
  output \g37157/_0_  ;
  output \g37158/_0_  ;
  output \g37159/_0_  ;
  output \g37160/_0_  ;
  output \g37161/_0_  ;
  output \g37162/_0_  ;
  output \g37163/_0_  ;
  output \g37164/_0_  ;
  output \g37165/_0_  ;
  output \g37166/_0_  ;
  output \g37167/_0_  ;
  output \g37168/_0_  ;
  output \g37169/_0_  ;
  output \g37170/_0_  ;
  output \g37171/_0_  ;
  output \g37172/_0_  ;
  output \g37173/_0_  ;
  output \g37174/_0_  ;
  output \g37175/_0_  ;
  output \g37176/_0_  ;
  output \g37177/_0_  ;
  output \g37178/_0_  ;
  output \g37179/_0_  ;
  output \g37180/_0_  ;
  output \g37181/_0_  ;
  output \g37182/_0_  ;
  output \g37183/_0_  ;
  output \g37184/_0_  ;
  output \g37185/_0_  ;
  output \g37187/_0_  ;
  output \g37188/_0_  ;
  output \g37190/_0_  ;
  output \g37191/_0_  ;
  output \g37192/_0_  ;
  output \g37193/_0_  ;
  output \g37194/_0_  ;
  output \g37372/_3_  ;
  output \g37377/_0_  ;
  output \g37378/_0_  ;
  output \g37379/_0_  ;
  output \g37380/_0_  ;
  output \g37381/_0_  ;
  output \g37382/_0_  ;
  output \g37383/_0_  ;
  output \g37384/_0_  ;
  output \g37385/_0_  ;
  output \g37386/_0_  ;
  output \g37387/_0_  ;
  output \g37388/_0_  ;
  output \g37389/_0_  ;
  output \g37390/_0_  ;
  output \g37391/_0_  ;
  output \g37392/_0_  ;
  output \g37393/_0_  ;
  output \g37394/_0_  ;
  output \g37395/_0_  ;
  output \g37396/_0_  ;
  output \g37397/_0_  ;
  output \g37398/_0_  ;
  output \g37399/_0_  ;
  output \g37400/_0_  ;
  output \g37401/_0_  ;
  output \g37402/_0_  ;
  output \g37403/_0_  ;
  output \g37404/_0_  ;
  output \g37405/_0_  ;
  output \g37406/_0_  ;
  output \g37407/_0_  ;
  output \g37408/_0_  ;
  output \g37409/_0_  ;
  output \g37410/_0_  ;
  output \g37411/_0_  ;
  output \g37412/_0_  ;
  output \g37413/_0_  ;
  output \g37576/_3_  ;
  output \g37590/_2_  ;
  output \g40278/_0_  ;
  output \g40379/_0_  ;
  output \g40389/_2_  ;
  output \g40390/_2_  ;
  output \g40391/_0_  ;
  output \g40393/_2_  ;
  output \g40395/_0_  ;
  output \g40397/_0_  ;
  output \g40400/_0_  ;
  output \g40402/_0_  ;
  output \g45458/_0_  ;
  output \g45675/_0_  ;
  output \g45677/_0_  ;
  output \g45678/_0_  ;
  output \g45682/_0_  ;
  output sync_pad_o_pad ;
  output \u14_u0_full_empty_r_reg/P0001_reg_syn_3  ;
  output \u14_u1_full_empty_r_reg/P0001_reg_syn_3  ;
  output \u14_u2_full_empty_r_reg/P0001_reg_syn_3  ;
  output \u14_u3_full_empty_r_reg/P0001_reg_syn_3  ;
  output \u14_u4_full_empty_r_reg/P0001_reg_syn_3  ;
  output \u14_u5_full_empty_r_reg/P0001_reg_syn_3  ;
  output \u14_u6_full_empty_r_reg/P0001_reg_syn_3  ;
  output \u14_u7_full_empty_r_reg/P0001_reg_syn_3  ;
  output \u14_u8_full_empty_r_reg/P0001_reg_syn_3  ;
  output \u1_slt0_reg[11]/P0001_reg_syn_3  ;
  output \u1_slt0_reg[12]/P0001_reg_syn_3  ;
  output \u1_slt0_reg[15]/P0001_reg_syn_3  ;
  output \u1_slt0_reg[9]/P0001_reg_syn_3  ;
  output \u1_slt1_reg[10]/P0001_reg_syn_3  ;
  output \u1_slt1_reg[11]/P0001_reg_syn_3  ;
  output \u1_slt1_reg[5]/P0001_reg_syn_3  ;
  output \u1_slt1_reg[6]/P0001_reg_syn_3  ;
  output \u1_slt1_reg[7]/P0001_reg_syn_3  ;
  output \u1_slt1_reg[8]/P0001_reg_syn_3  ;
  output wb_err_o_pad ;
  wire n2146 , n2147 , n2148 , n2149 , n2150 , n2151 , n2152 , n2153 , n2154 , n2155 , n2156 , n2157 , n2158 , n2159 , n2160 , n2161 , n2162 , n2163 , n2164 , n2165 , n2166 , n2167 , n2168 , n2169 , n2170 , n2171 , n2172 , n2173 , n2174 , n2175 , n2176 , n2177 , n2178 , n2179 , n2180 , n2181 , n2182 , n2183 , n2184 , n2185 , n2186 , n2187 , n2188 , n2189 , n2190 , n2191 , n2192 , n2193 , n2194 , n2195 , n2196 , n2197 , n2198 , n2199 , n2200 , n2201 , n2202 , n2203 , n2204 , n2205 , n2206 , n2207 , n2208 , n2209 , n2210 , n2211 , n2212 , n2213 , n2214 , n2215 , n2216 , n2217 , n2218 , n2219 , n2220 , n2221 , n2222 , n2223 , n2224 , n2225 , n2226 , n2227 , n2228 , n2229 , n2230 , n2231 , n2232 , n2233 , n2234 , n2235 , n2236 , n2237 , n2238 , n2239 , n2240 , n2241 , n2242 , n2243 , n2244 , n2245 , n2246 , n2247 , n2248 , n2249 , n2250 , n2251 , n2252 , n2253 , n2254 , n2255 , n2256 , n2257 , n2258 , n2259 , n2260 , n2261 , n2262 , n2263 , n2264 , n2265 , n2266 , n2267 , n2268 , n2269 , n2270 , n2271 , n2272 , n2273 , n2274 , n2275 , n2276 , n2277 , n2278 , n2279 , n2280 , n2281 , n2282 , n2283 , n2284 , n2285 , n2286 , n2287 , n2288 , n2289 , n2290 , n2291 , n2292 , n2293 , n2294 , n2295 , n2296 , n2297 , n2298 , n2299 , n2300 , n2301 , n2302 , n2303 , n2304 , n2305 , n2306 , n2307 , n2308 , n2309 , n2310 , n2311 , n2312 , n2313 , n2314 , n2315 , n2316 , n2317 , n2318 , n2319 , n2320 , n2321 , n2322 , n2323 , n2324 , n2325 , n2326 , n2327 , n2328 , n2329 , n2330 , n2331 , n2332 , n2333 , n2334 , n2335 , n2336 , n2337 , n2338 , n2339 , n2340 , n2341 , n2342 , n2343 , n2344 , n2345 , n2346 , n2347 , n2348 , n2349 , n2350 , n2351 , n2352 , n2353 , n2354 , n2355 , n2356 , n2357 , n2358 , n2359 , n2360 , n2361 , n2362 , n2363 , n2364 , n2365 , n2366 , n2367 , n2368 , n2369 , n2370 , n2371 , n2372 , n2373 , n2374 , n2375 , n2376 , n2377 , n2378 , n2379 , n2380 , n2381 , n2382 , n2383 , n2384 , n2385 , n2386 , n2387 , n2388 , n2389 , n2390 , n2391 , n2392 , n2393 , n2394 , n2395 , n2396 , n2397 , n2398 , n2399 , n2400 , n2401 , n2402 , n2403 , n2404 , n2405 , n2406 , n2407 , n2408 , n2409 , n2410 , n2411 , n2412 , n2413 , n2414 , n2415 , n2416 , n2417 , n2418 , n2419 , n2420 , n2421 , n2422 , n2423 , n2424 , n2425 , n2426 , n2427 , n2428 , n2429 , n2430 , n2431 , n2432 , n2433 , n2434 , n2435 , n2436 , n2437 , n2438 , n2439 , n2440 , n2441 , n2442 , n2443 , n2444 , n2445 , n2446 , n2447 , n2448 , n2449 , n2450 , n2451 , n2452 , n2453 , n2454 , n2455 , n2456 , n2457 , n2458 , n2459 , n2460 , n2461 , n2462 , n2463 , n2464 , n2465 , n2466 , n2467 , n2468 , n2469 , n2470 , n2471 , n2472 , n2473 , n2474 , n2475 , n2476 , n2477 , n2478 , n2479 , n2480 , n2481 , n2482 , n2483 , n2484 , n2485 , n2486 , n2487 , n2488 , n2489 , n2490 , n2491 , n2492 , n2493 , n2494 , n2495 , n2496 , n2497 , n2498 , n2499 , n2500 , n2501 , n2502 , n2503 , n2504 , n2505 , n2506 , n2507 , n2508 , n2509 , n2510 , n2511 , n2512 , n2513 , n2514 , n2515 , n2516 , n2517 , n2518 , n2519 , n2520 , n2521 , n2522 , n2523 , n2524 , n2525 , n2526 , n2527 , n2528 , n2529 , n2530 , n2531 , n2532 , n2533 , n2534 , n2535 , n2536 , n2537 , n2538 , n2539 , n2540 , n2541 , n2542 , n2543 , n2544 , n2545 , n2546 , n2547 , n2548 , n2549 , n2550 , n2551 , n2552 , n2553 , n2554 , n2555 , n2556 , n2557 , n2558 , n2559 , n2560 , n2561 , n2562 , n2563 , n2564 , n2565 , n2566 , n2567 , n2568 , n2569 , n2570 , n2571 , n2572 , n2573 , n2574 , n2575 , n2576 , n2577 , n2578 , n2579 , n2580 , n2581 , n2582 , n2583 , n2584 , n2585 , n2586 , n2587 , n2588 , n2589 , n2590 , n2591 , n2592 , n2593 , n2594 , n2595 , n2596 , n2597 , n2598 , n2599 , n2600 , n2601 , n2602 , n2603 , n2604 , n2605 , n2606 , n2607 , n2608 , n2609 , n2610 , n2611 , n2612 , n2613 , n2614 , n2615 , n2616 , n2617 , n2618 , n2619 , n2620 , n2621 , n2622 , n2623 , n2624 , n2625 , n2626 , n2627 , n2628 , n2629 , n2630 , n2631 , n2632 , n2633 , n2634 , n2635 , n2636 , n2637 , n2638 , n2639 , n2640 , n2641 , n2642 , n2643 , n2644 , n2645 , n2646 , n2647 , n2648 , n2649 , n2650 , n2651 , n2652 , n2653 , n2654 , n2655 , n2656 , n2657 , n2658 , n2659 , n2660 , n2661 , n2662 , n2663 , n2664 , n2665 , n2666 , n2667 , n2668 , n2669 , n2670 , n2671 , n2672 , n2673 , n2674 , n2675 , n2676 , n2677 , n2678 , n2679 , n2680 , n2681 , n2682 , n2683 , n2684 , n2685 , n2686 , n2687 , n2688 , n2689 , n2690 , n2691 , n2692 , n2693 , n2694 , n2695 , n2696 , n2697 , n2698 , n2699 , n2700 , n2701 , n2702 , n2703 , n2704 , n2705 , n2706 , n2707 , n2708 , n2709 , n2710 , n2711 , n2712 , n2713 , n2714 , n2715 , n2716 , n2717 , n2718 , n2719 , n2720 , n2721 , n2722 , n2723 , n2724 , n2725 , n2726 , n2727 , n2728 , n2729 , n2730 , n2731 , n2732 , n2733 , n2734 , n2735 , n2736 , n2737 , n2738 , n2739 , n2740 , n2741 , n2742 , n2743 , n2744 , n2745 , n2746 , n2747 , n2748 , n2749 , n2750 , n2751 , n2752 , n2753 , n2754 , n2755 , n2756 , n2757 , n2758 , n2759 , n2760 , n2761 , n2762 , n2763 , n2764 , n2765 , n2766 , n2767 , n2768 , n2769 , n2770 , n2771 , n2772 , n2773 , n2774 , n2775 , n2776 , n2777 , n2778 , n2779 , n2780 , n2781 , n2782 , n2783 , n2784 , n2785 , n2786 , n2787 , n2788 , n2789 , n2790 , n2791 , n2792 , n2793 , n2794 , n2795 , n2796 , n2797 , n2798 , n2799 , n2800 , n2801 , n2802 , n2803 , n2804 , n2805 , n2806 , n2807 , n2808 , n2809 , n2810 , n2811 , n2812 , n2813 , n2814 , n2815 , n2816 , n2817 , n2818 , n2819 , n2820 , n2821 , n2822 , n2823 , n2824 , n2825 , n2826 , n2827 , n2828 , n2829 , n2830 , n2831 , n2832 , n2833 , n2834 , n2835 , n2836 , n2837 , n2838 , n2839 , n2840 , n2841 , n2842 , n2843 , n2844 , n2845 , n2846 , n2847 , n2848 , n2849 , n2850 , n2851 , n2852 , n2853 , n2854 , n2855 , n2856 , n2857 , n2858 , n2859 , n2860 , n2861 , n2862 , n2863 , n2864 , n2865 , n2866 , n2867 , n2868 , n2869 , n2870 , n2871 , n2872 , n2873 , n2874 , n2875 , n2876 , n2877 , n2878 , n2879 , n2880 , n2881 , n2882 , n2883 , n2884 , n2885 , n2886 , n2887 , n2888 , n2889 , n2890 , n2891 , n2892 , n2893 , n2894 , n2895 , n2896 , n2897 , n2898 , n2899 , n2900 , n2901 , n2902 , n2903 , n2904 , n2905 , n2906 , n2907 , n2908 , n2909 , n2910 , n2911 , n2912 , n2913 , n2914 , n2915 , n2916 , n2917 , n2918 , n2919 , n2920 , n2921 , n2922 , n2923 , n2924 , n2925 , n2926 , n2927 , n2928 , n2929 , n2930 , n2931 , n2932 , n2933 , n2934 , n2935 , n2936 , n2937 , n2938 , n2939 , n2940 , n2941 , n2942 , n2943 , n2944 , n2945 , n2946 , n2947 , n2948 , n2949 , n2950 , n2951 , n2952 , n2953 , n2954 , n2955 , n2956 , n2957 , n2958 , n2959 , n2960 , n2961 , n2962 , n2963 , n2964 , n2965 , n2966 , n2967 , n2968 , n2969 , n2970 , n2971 , n2972 , n2973 , n2974 , n2975 , n2976 , n2977 , n2978 , n2979 , n2980 , n2981 , n2982 , n2983 , n2984 , n2985 , n2986 , n2987 , n2988 , n2989 , n2990 , n2991 , n2992 , n2993 , n2994 , n2995 , n2996 , n2997 , n2998 , n2999 , n3000 , n3001 , n3002 , n3003 , n3004 , n3005 , n3006 , n3007 , n3008 , n3009 , n3010 , n3011 , n3012 , n3013 , n3014 , n3015 , n3016 , n3017 , n3018 , n3019 , n3020 , n3021 , n3022 , n3023 , n3024 , n3025 , n3026 , n3027 , n3028 , n3029 , n3030 , n3031 , n3032 , n3033 , n3034 , n3035 , n3036 , n3037 , n3038 , n3039 , n3040 , n3041 , n3042 , n3043 , n3044 , n3045 , n3046 , n3047 , n3048 , n3049 , n3050 , n3051 , n3052 , n3053 , n3054 , n3055 , n3056 , n3057 , n3058 , n3059 , n3060 , n3061 , n3062 , n3063 , n3064 , n3065 , n3066 , n3067 , n3068 , n3069 , n3070 , n3071 , n3072 , n3073 , n3074 , n3075 , n3076 , n3077 , n3078 , n3079 , n3080 , n3081 , n3082 , n3083 , n3084 , n3085 , n3086 , n3087 , n3088 , n3089 , n3090 , n3091 , n3092 , n3093 , n3094 , n3095 , n3096 , n3097 , n3098 , n3099 , n3100 , n3101 , n3102 , n3103 , n3104 , n3105 , n3106 , n3107 , n3108 , n3109 , n3110 , n3111 , n3112 , n3113 , n3114 , n3115 , n3116 , n3117 , n3118 , n3119 , n3120 , n3121 , n3122 , n3123 , n3124 , n3125 , n3126 , n3127 , n3128 , n3129 , n3130 , n3131 , n3132 , n3133 , n3134 , n3135 , n3136 , n3137 , n3138 , n3139 , n3140 , n3141 , n3142 , n3143 , n3144 , n3145 , n3146 , n3147 , n3148 , n3149 , n3150 , n3151 , n3152 , n3153 , n3154 , n3155 , n3156 , n3157 , n3158 , n3159 , n3160 , n3161 , n3162 , n3163 , n3164 , n3165 , n3166 , n3167 , n3168 , n3169 , n3170 , n3171 , n3172 , n3173 , n3174 , n3175 , n3176 , n3177 , n3178 , n3179 , n3180 , n3181 , n3182 , n3183 , n3184 , n3185 , n3186 , n3187 , n3188 , n3189 , n3190 , n3191 , n3192 , n3193 , n3194 , n3195 , n3196 , n3197 , n3198 , n3199 , n3200 , n3201 , n3202 , n3203 , n3204 , n3205 , n3206 , n3207 , n3208 , n3209 , n3210 , n3211 , n3212 , n3213 , n3214 , n3215 , n3216 , n3217 , n3218 , n3219 , n3220 , n3221 , n3222 , n3223 , n3224 , n3225 , n3226 , n3227 , n3228 , n3229 , n3230 , n3231 , n3232 , n3233 , n3234 , n3235 , n3236 , n3237 , n3238 , n3239 , n3240 , n3241 , n3242 , n3243 , n3244 , n3245 , n3246 , n3247 , n3248 , n3249 , n3250 , n3251 , n3252 , n3253 , n3254 , n3255 , n3256 , n3257 , n3258 , n3259 , n3260 , n3261 , n3262 , n3263 , n3264 , n3265 , n3266 , n3267 , n3268 , n3269 , n3270 , n3271 , n3272 , n3273 , n3274 , n3275 , n3276 , n3277 , n3278 , n3279 , n3280 , n3281 , n3282 , n3283 , n3284 , n3285 , n3286 , n3287 , n3288 , n3289 , n3290 , n3291 , n3292 , n3293 , n3294 , n3295 , n3296 , n3297 , n3298 , n3299 , n3300 , n3301 , n3302 , n3303 , n3304 , n3305 , n3306 , n3307 , n3308 , n3309 , n3310 , n3311 , n3312 , n3313 , n3314 , n3315 , n3316 , n3317 , n3318 , n3319 , n3320 , n3321 , n3322 , n3323 , n3324 , n3325 , n3326 , n3327 , n3328 , n3329 , n3330 , n3331 , n3332 , n3333 , n3334 , n3335 , n3336 , n3337 , n3338 , n3339 , n3340 , n3341 , n3342 , n3343 , n3344 , n3345 , n3346 , n3347 , n3348 , n3349 , n3350 , n3351 , n3352 , n3353 , n3354 , n3355 , n3356 , n3357 , n3358 , n3359 , n3360 , n3361 , n3362 , n3363 , n3364 , n3365 , n3366 , n3367 , n3368 , n3369 , n3370 , n3371 , n3372 , n3373 , n3374 , n3375 , n3376 , n3377 , n3378 , n3379 , n3380 , n3381 , n3382 , n3383 , n3384 , n3385 , n3386 , n3387 , n3388 , n3389 , n3390 , n3391 , n3392 , n3393 , n3394 , n3395 , n3396 , n3397 , n3398 , n3399 , n3400 , n3401 , n3402 , n3403 , n3404 , n3405 , n3406 , n3407 , n3408 , n3409 , n3410 , n3411 , n3412 , n3413 , n3414 , n3415 , n3416 , n3417 , n3418 , n3419 , n3420 , n3421 , n3422 , n3423 , n3424 , n3425 , n3426 , n3427 , n3428 , n3429 , n3430 , n3431 , n3432 , n3433 , n3434 , n3435 , n3436 , n3437 , n3438 , n3439 , n3440 , n3441 , n3442 , n3443 , n3444 , n3445 , n3446 , n3447 , n3448 , n3449 , n3450 , n3451 , n3452 , n3453 , n3454 , n3455 , n3456 , n3457 , n3458 , n3459 , n3460 , n3461 , n3462 , n3463 , n3464 , n3465 , n3466 , n3467 , n3468 , n3469 , n3470 , n3471 , n3472 , n3473 , n3474 , n3475 , n3476 , n3477 , n3478 , n3479 , n3480 , n3481 , n3482 , n3483 , n3484 , n3485 , n3486 , n3487 , n3488 , n3489 , n3490 , n3491 , n3492 , n3493 , n3494 , n3495 , n3496 , n3497 , n3498 , n3499 , n3500 , n3501 , n3502 , n3503 , n3504 , n3505 , n3506 , n3507 , n3508 , n3509 , n3510 , n3511 , n3512 , n3513 , n3514 , n3515 , n3516 , n3517 , n3518 , n3519 , n3520 , n3521 , n3522 , n3523 , n3524 , n3525 , n3526 , n3527 , n3528 , n3529 , n3530 , n3531 , n3532 , n3533 , n3534 , n3535 , n3536 , n3537 , n3538 , n3539 , n3540 , n3541 , n3542 , n3543 , n3544 , n3545 , n3546 , n3547 , n3548 , n3549 , n3550 , n3551 , n3552 , n3553 , n3554 , n3555 , n3556 , n3557 , n3558 , n3559 , n3560 , n3561 , n3562 , n3563 , n3564 , n3565 , n3566 , n3567 , n3568 , n3569 , n3570 , n3571 , n3572 , n3573 , n3574 , n3575 , n3576 , n3577 , n3578 , n3579 , n3580 , n3581 , n3582 , n3583 , n3584 , n3585 , n3586 , n3587 , n3588 , n3589 , n3590 , n3591 , n3592 , n3593 , n3594 , n3595 , n3596 , n3597 , n3598 , n3599 , n3600 , n3601 , n3602 , n3603 , n3604 , n3605 , n3606 , n3607 , n3608 , n3609 , n3610 , n3611 , n3612 , n3613 , n3614 , n3615 , n3616 , n3617 , n3618 , n3619 , n3620 , n3621 , n3622 , n3623 , n3624 , n3625 , n3626 , n3627 , n3628 , n3629 , n3630 , n3631 , n3632 , n3633 , n3634 , n3635 , n3636 , n3637 , n3638 , n3639 , n3640 , n3641 , n3642 , n3643 , n3644 , n3645 , n3646 , n3647 , n3648 , n3649 , n3650 , n3651 , n3652 , n3653 , n3654 , n3655 , n3656 , n3657 , n3658 , n3659 , n3660 , n3661 , n3662 , n3663 , n3664 , n3665 , n3666 , n3667 , n3668 , n3669 , n3670 , n3671 , n3672 , n3673 , n3674 , n3675 , n3676 , n3677 , n3678 , n3679 , n3680 , n3681 , n3682 , n3683 , n3684 , n3685 , n3686 , n3687 , n3688 , n3689 , n3690 , n3691 , n3692 , n3693 , n3694 , n3695 , n3696 , n3697 , n3698 , n3699 , n3700 , n3701 , n3702 , n3703 , n3704 , n3705 , n3706 , n3707 , n3708 , n3709 , n3710 , n3711 , n3712 , n3713 , n3714 , n3715 , n3716 , n3717 , n3718 , n3719 , n3720 , n3721 , n3722 , n3723 , n3724 , n3725 , n3726 , n3727 , n3728 , n3729 , n3730 , n3731 , n3732 , n3733 , n3734 , n3735 , n3736 , n3737 , n3738 , n3739 , n3740 , n3741 , n3742 , n3743 , n3744 , n3745 , n3746 , n3747 , n3748 , n3749 , n3750 , n3751 , n3752 , n3753 , n3754 , n3755 , n3756 , n3757 , n3758 , n3759 , n3760 , n3761 , n3762 , n3763 , n3764 , n3765 , n3766 , n3767 , n3768 , n3769 , n3770 , n3771 , n3772 , n3773 , n3774 , n3775 , n3776 , n3777 , n3778 , n3779 , n3780 , n3781 , n3782 , n3783 , n3784 , n3785 , n3786 , n3787 , n3788 , n3789 , n3790 , n3791 , n3792 , n3793 , n3794 , n3795 , n3796 , n3797 , n3798 , n3799 , n3800 , n3801 , n3802 , n3803 , n3804 , n3805 , n3806 , n3807 , n3808 , n3809 , n3810 , n3811 , n3812 , n3813 , n3814 , n3815 , n3816 , n3817 , n3818 , n3819 , n3820 , n3821 , n3822 , n3823 , n3824 , n3825 , n3826 , n3827 , n3828 , n3829 , n3830 , n3831 , n3832 , n3833 , n3834 , n3835 , n3836 , n3837 , n3838 , n3839 , n3840 , n3841 , n3842 , n3843 , n3844 , n3845 , n3846 , n3847 , n3848 , n3849 , n3850 , n3851 , n3852 , n3853 , n3854 , n3855 , n3856 , n3857 , n3858 , n3859 , n3860 , n3861 , n3862 , n3863 , n3864 , n3865 , n3866 , n3867 , n3868 , n3869 , n3870 , n3871 , n3872 , n3873 , n3874 , n3875 , n3876 , n3877 , n3878 , n3879 , n3880 , n3881 , n3882 , n3883 , n3884 , n3885 , n3886 , n3887 , n3888 , n3889 , n3890 , n3891 , n3892 , n3893 , n3894 , n3895 , n3896 , n3897 , n3898 , n3899 , n3900 , n3901 , n3902 , n3903 , n3904 , n3905 , n3906 , n3907 , n3908 , n3909 , n3910 , n3911 , n3912 , n3913 , n3914 , n3915 , n3916 , n3917 , n3918 , n3919 , n3920 , n3921 , n3922 , n3923 , n3924 , n3925 , n3926 , n3927 , n3928 , n3929 , n3930 , n3931 , n3932 , n3933 , n3934 , n3935 , n3936 , n3937 , n3938 , n3939 , n3940 , n3941 , n3942 , n3943 , n3944 , n3945 , n3946 , n3947 , n3948 , n3949 , n3950 , n3951 , n3952 , n3953 , n3954 , n3955 , n3956 , n3957 , n3958 , n3959 , n3960 , n3961 , n3962 , n3963 , n3964 , n3965 , n3966 , n3967 , n3968 , n3969 , n3970 , n3971 , n3972 , n3973 , n3974 , n3975 , n3976 , n3977 , n3978 , n3979 , n3980 , n3981 , n3982 , n3983 , n3984 , n3985 , n3986 , n3987 , n3988 , n3989 , n3990 , n3991 , n3992 , n3993 , n3994 , n3995 , n3996 , n3997 , n3998 , n3999 , n4000 , n4001 , n4002 , n4003 , n4004 , n4005 , n4006 , n4007 , n4008 , n4009 , n4010 , n4011 , n4012 , n4013 , n4014 , n4015 , n4016 , n4017 , n4018 , n4019 , n4020 , n4021 , n4022 , n4023 , n4024 , n4025 , n4026 , n4027 , n4028 , n4029 , n4030 , n4031 , n4032 , n4033 , n4034 , n4035 , n4036 , n4037 , n4038 , n4039 , n4040 , n4041 , n4042 , n4043 , n4044 , n4045 , n4046 , n4047 , n4048 , n4049 , n4050 , n4051 , n4052 , n4053 , n4054 , n4055 , n4056 , n4057 , n4058 , n4059 , n4060 , n4061 , n4062 , n4063 , n4064 , n4065 , n4066 , n4067 , n4068 , n4069 , n4070 , n4071 , n4072 , n4073 , n4074 , n4075 , n4076 , n4077 , n4078 , n4079 , n4080 , n4081 , n4082 , n4083 , n4084 , n4085 , n4086 , n4087 , n4088 , n4089 , n4090 , n4091 , n4092 , n4093 , n4094 , n4095 , n4096 , n4097 , n4098 , n4099 , n4100 , n4101 , n4102 , n4103 , n4104 , n4105 , n4106 , n4107 , n4108 , n4109 , n4110 , n4111 , n4112 , n4113 , n4114 , n4115 , n4116 , n4117 , n4118 , n4119 , n4120 , n4121 , n4122 , n4123 , n4124 , n4125 , n4126 , n4127 , n4128 , n4129 , n4130 , n4131 , n4132 , n4133 , n4134 , n4135 , n4136 , n4137 , n4138 , n4139 , n4140 , n4141 , n4142 , n4143 , n4144 , n4145 , n4146 , n4147 , n4148 , n4149 , n4150 , n4151 , n4152 , n4153 , n4154 , n4155 , n4156 , n4157 , n4158 , n4159 , n4160 , n4161 , n4162 , n4163 , n4164 , n4165 , n4166 , n4167 , n4168 , n4169 , n4170 , n4171 , n4172 , n4173 , n4174 , n4175 , n4176 , n4177 , n4178 , n4179 , n4180 , n4181 , n4182 , n4183 , n4184 , n4185 , n4186 , n4187 , n4188 , n4189 , n4190 , n4191 , n4192 , n4193 , n4194 , n4195 , n4196 , n4197 , n4198 , n4199 , n4200 , n4201 , n4202 , n4203 , n4204 , n4205 , n4206 , n4207 , n4208 , n4209 , n4210 , n4211 , n4212 , n4213 , n4214 , n4215 , n4216 , n4217 , n4218 , n4219 , n4220 , n4221 , n4222 , n4223 , n4224 , n4225 , n4226 , n4227 , n4228 , n4229 , n4230 , n4231 , n4232 , n4233 , n4234 , n4235 , n4236 , n4237 , n4238 , n4239 , n4240 , n4241 , n4242 , n4243 , n4244 , n4245 , n4246 , n4247 , n4248 , n4249 , n4250 , n4251 , n4252 , n4253 , n4254 , n4255 , n4256 , n4257 , n4258 , n4259 , n4260 , n4261 , n4262 , n4263 , n4264 , n4265 , n4266 , n4267 , n4268 , n4269 , n4270 , n4271 , n4272 , n4273 , n4274 , n4275 , n4276 , n4277 , n4278 , n4279 , n4280 , n4281 , n4282 , n4283 , n4284 , n4285 , n4286 , n4287 , n4288 , n4289 , n4290 , n4291 , n4292 , n4293 , n4294 , n4295 , n4296 , n4297 , n4298 , n4299 , n4300 , n4301 , n4302 , n4303 , n4304 , n4305 , n4306 , n4307 , n4308 , n4309 , n4310 , n4311 , n4312 , n4313 , n4314 , n4315 , n4316 , n4317 , n4318 , n4319 , n4320 , n4321 , n4322 , n4323 , n4324 , n4325 , n4326 , n4327 , n4328 , n4329 , n4330 , n4331 , n4332 , n4333 , n4334 , n4335 , n4336 , n4337 , n4338 , n4339 , n4340 , n4341 , n4342 , n4343 , n4344 , n4345 , n4346 , n4347 , n4348 , n4349 , n4350 , n4351 , n4352 , n4353 , n4354 , n4355 , n4356 , n4357 , n4358 , n4359 , n4360 , n4361 , n4362 , n4363 , n4364 , n4365 , n4366 , n4367 , n4368 , n4369 , n4370 , n4371 , n4372 , n4373 , n4374 , n4375 , n4376 , n4377 , n4378 , n4379 , n4380 , n4381 , n4382 , n4383 , n4384 , n4385 , n4386 , n4387 , n4388 , n4389 , n4390 , n4391 , n4392 , n4393 , n4394 , n4395 , n4396 , n4397 , n4398 , n4399 , n4400 , n4401 , n4402 , n4403 , n4404 , n4405 , n4406 , n4407 , n4408 , n4409 , n4410 , n4411 , n4412 , n4413 , n4414 , n4415 , n4416 , n4417 , n4418 , n4419 , n4420 , n4421 , n4422 , n4423 , n4424 , n4425 , n4426 , n4427 , n4428 , n4429 , n4430 , n4431 , n4432 , n4433 , n4434 , n4435 , n4436 , n4437 , n4438 , n4439 , n4440 , n4441 , n4442 , n4443 , n4444 , n4445 , n4446 , n4447 , n4448 , n4449 , n4450 , n4451 , n4452 , n4453 , n4454 , n4455 , n4456 , n4457 , n4458 , n4459 , n4460 , n4461 , n4462 , n4463 , n4464 , n4465 , n4466 , n4467 , n4468 , n4469 , n4470 , n4471 , n4472 , n4473 , n4474 , n4475 , n4476 , n4477 , n4478 , n4479 , n4480 , n4481 , n4482 , n4483 , n4484 , n4485 , n4486 , n4487 , n4488 , n4489 , n4490 , n4491 , n4492 , n4493 , n4494 , n4495 , n4496 , n4497 , n4498 , n4499 , n4500 , n4501 , n4502 , n4503 , n4504 , n4505 , n4506 , n4507 , n4508 , n4509 , n4510 , n4511 , n4512 , n4513 , n4514 , n4515 , n4516 , n4517 , n4518 , n4519 , n4520 , n4521 , n4522 , n4523 , n4524 , n4525 , n4526 , n4527 , n4528 , n4529 , n4530 , n4531 , n4532 , n4533 , n4534 , n4535 , n4536 , n4537 , n4538 , n4539 , n4540 , n4541 , n4542 , n4543 , n4544 , n4545 , n4546 , n4547 , n4548 , n4549 , n4550 , n4551 , n4552 , n4553 , n4554 , n4555 , n4556 , n4557 , n4558 , n4559 , n4560 , n4561 , n4562 , n4563 , n4564 , n4565 , n4566 , n4567 , n4568 , n4569 , n4570 , n4571 , n4572 , n4573 , n4574 , n4575 , n4576 , n4577 , n4578 , n4579 , n4580 , n4581 , n4582 , n4583 , n4584 , n4585 , n4586 , n4587 , n4588 , n4589 , n4590 , n4591 , n4592 , n4593 , n4594 , n4595 , n4596 , n4597 , n4598 , n4599 , n4600 , n4601 , n4602 , n4603 , n4604 , n4605 , n4606 , n4607 , n4608 , n4609 , n4610 , n4611 , n4612 , n4613 , n4614 , n4615 , n4616 , n4617 , n4618 , n4619 , n4620 , n4621 , n4622 , n4623 , n4624 , n4625 , n4626 , n4627 , n4628 , n4629 , n4630 , n4631 , n4632 , n4633 , n4634 , n4635 , n4636 , n4637 , n4638 , n4639 , n4640 , n4641 , n4642 , n4643 , n4644 , n4645 , n4646 , n4647 , n4648 , n4649 , n4650 , n4651 , n4652 , n4653 , n4654 , n4655 , n4656 , n4657 , n4658 , n4659 , n4660 , n4661 , n4662 , n4663 , n4664 , n4665 , n4666 , n4667 , n4668 , n4669 , n4670 , n4671 , n4672 , n4673 , n4674 , n4675 , n4676 , n4677 , n4678 , n4679 , n4680 , n4681 , n4682 , n4683 , n4684 , n4685 , n4686 , n4687 , n4688 , n4689 , n4690 , n4691 , n4692 , n4693 , n4694 , n4695 , n4696 , n4697 , n4698 , n4699 , n4700 , n4701 , n4702 , n4703 , n4704 , n4705 , n4706 , n4707 , n4708 , n4709 , n4710 , n4711 , n4712 , n4713 , n4714 , n4715 , n4716 , n4717 , n4718 , n4719 , n4720 , n4721 , n4722 , n4723 , n4724 , n4725 , n4726 , n4727 , n4728 , n4729 , n4730 , n4731 , n4732 , n4733 , n4734 , n4735 , n4736 , n4737 , n4738 , n4739 , n4740 , n4741 , n4742 , n4743 , n4744 , n4745 , n4746 , n4747 , n4748 , n4749 , n4750 , n4751 , n4752 , n4753 , n4754 , n4755 , n4756 , n4757 , n4758 , n4759 , n4760 , n4761 , n4762 , n4763 , n4764 , n4765 , n4766 , n4767 , n4768 , n4769 , n4770 , n4771 , n4772 , n4773 , n4774 , n4775 , n4776 , n4777 , n4778 , n4779 , n4780 , n4781 , n4782 , n4783 , n4784 , n4785 , n4786 , n4787 , n4788 , n4789 , n4790 , n4791 , n4792 , n4793 , n4794 , n4795 , n4796 , n4797 , n4798 , n4799 , n4800 , n4801 , n4802 , n4803 , n4804 , n4805 , n4806 , n4807 , n4808 , n4809 , n4810 , n4811 , n4812 , n4813 , n4814 , n4815 , n4816 , n4817 , n4818 , n4819 , n4820 , n4821 , n4822 , n4823 , n4824 , n4825 , n4826 , n4827 , n4828 , n4829 , n4830 , n4831 , n4832 , n4833 , n4834 , n4835 , n4836 , n4837 , n4838 , n4839 , n4840 , n4841 , n4842 , n4843 , n4844 , n4845 , n4846 , n4847 , n4848 , n4849 , n4850 , n4851 , n4852 , n4853 , n4854 , n4855 , n4856 , n4857 , n4858 , n4859 , n4860 , n4861 , n4862 , n4863 , n4864 , n4865 , n4866 , n4867 , n4868 , n4869 , n4870 , n4871 , n4872 , n4873 , n4874 , n4875 , n4876 , n4877 , n4878 , n4879 , n4880 , n4881 , n4882 , n4883 , n4884 , n4885 , n4886 , n4887 , n4888 , n4889 , n4890 , n4891 , n4892 , n4893 , n4894 , n4895 , n4896 , n4897 , n4898 , n4899 , n4900 , n4901 , n4902 , n4903 , n4904 , n4905 , n4906 , n4907 , n4908 , n4909 , n4910 , n4911 , n4912 , n4913 , n4914 , n4915 , n4916 , n4917 , n4918 , n4919 , n4920 , n4921 , n4922 , n4923 , n4924 , n4925 , n4926 , n4927 , n4928 , n4929 , n4930 , n4931 , n4932 , n4933 , n4934 , n4935 , n4936 , n4937 , n4938 , n4939 , n4940 , n4941 , n4942 , n4943 , n4944 , n4945 , n4946 , n4947 , n4948 , n4949 , n4950 , n4951 , n4952 , n4953 , n4954 , n4955 , n4956 , n4957 , n4958 , n4959 , n4960 , n4961 , n4962 , n4963 , n4964 , n4965 , n4966 , n4967 , n4968 , n4969 , n4970 , n4971 , n4972 , n4973 , n4974 , n4975 , n4976 , n4977 , n4978 , n4979 , n4980 , n4981 , n4982 , n4983 , n4984 , n4985 , n4986 , n4987 , n4988 , n4989 , n4990 , n4991 , n4992 , n4993 , n4994 , n4995 , n4996 , n4997 , n4998 , n4999 , n5000 , n5001 , n5002 , n5003 , n5004 , n5005 , n5006 , n5007 , n5008 , n5009 , n5010 , n5011 , n5012 , n5013 , n5014 , n5015 , n5016 , n5017 , n5018 , n5019 , n5020 , n5021 , n5022 , n5023 , n5024 , n5025 , n5026 , n5027 , n5028 , n5029 , n5030 , n5031 , n5032 , n5033 , n5034 , n5035 , n5036 , n5037 , n5038 , n5039 , n5040 , n5041 , n5042 , n5043 , n5044 , n5045 , n5046 , n5047 , n5048 , n5049 , n5050 , n5051 , n5052 , n5053 , n5054 , n5055 , n5056 , n5057 , n5058 , n5059 , n5060 , n5061 , n5062 , n5063 , n5064 , n5065 , n5066 , n5067 , n5068 , n5069 , n5070 , n5071 , n5072 , n5073 , n5074 , n5075 , n5076 , n5077 , n5078 , n5079 , n5080 , n5081 , n5082 , n5083 , n5084 , n5085 , n5086 , n5087 , n5088 , n5089 , n5090 , n5091 , n5092 , n5093 , n5094 , n5095 , n5096 , n5097 , n5098 , n5099 , n5100 , n5101 , n5102 , n5103 , n5104 , n5105 , n5106 , n5107 , n5108 , n5109 , n5110 , n5111 , n5112 , n5113 , n5114 , n5115 , n5116 , n5117 , n5118 , n5119 , n5120 , n5121 , n5122 , n5123 , n5124 , n5125 , n5126 , n5127 , n5128 , n5129 , n5130 , n5131 , n5132 , n5133 , n5134 , n5135 , n5136 , n5137 , n5138 , n5139 , n5140 , n5141 , n5142 , n5143 , n5144 , n5145 , n5146 , n5147 , n5148 , n5149 , n5150 , n5151 , n5152 , n5153 , n5154 , n5155 , n5156 , n5157 , n5158 , n5159 , n5160 , n5161 , n5162 , n5163 , n5164 , n5165 , n5166 , n5167 , n5168 , n5169 , n5170 , n5171 , n5172 , n5173 , n5174 , n5175 , n5176 , n5177 , n5178 , n5179 , n5180 , n5181 , n5182 , n5183 , n5184 , n5185 , n5186 , n5187 , n5188 , n5189 , n5190 , n5191 , n5192 , n5193 , n5194 , n5195 , n5196 , n5197 , n5198 , n5199 , n5200 , n5201 , n5202 , n5203 , n5204 , n5205 , n5206 , n5207 , n5208 , n5209 , n5210 , n5211 , n5212 , n5213 , n5214 , n5215 , n5216 , n5217 , n5218 , n5219 , n5220 , n5221 , n5222 , n5223 , n5224 , n5225 , n5226 , n5227 , n5228 , n5229 , n5230 , n5231 , n5232 , n5233 , n5234 , n5235 , n5236 , n5237 , n5238 , n5239 , n5240 , n5241 , n5242 , n5243 , n5244 , n5245 , n5246 , n5247 , n5248 , n5249 , n5250 , n5251 , n5252 , n5253 , n5254 , n5255 , n5256 , n5257 , n5258 , n5259 , n5260 , n5261 , n5262 , n5263 , n5264 , n5265 , n5266 , n5267 , n5268 , n5269 , n5270 , n5271 , n5272 , n5273 , n5274 , n5275 , n5276 , n5277 , n5278 , n5279 , n5280 , n5281 , n5282 , n5283 , n5284 , n5285 , n5286 , n5287 , n5288 , n5289 , n5290 , n5291 , n5292 , n5293 , n5294 , n5295 , n5296 , n5297 , n5298 , n5299 , n5300 , n5301 , n5302 , n5303 , n5304 , n5305 , n5306 , n5307 , n5308 , n5309 , n5310 , n5311 , n5312 , n5313 , n5314 , n5315 , n5316 , n5317 , n5318 , n5319 , n5320 , n5321 , n5322 , n5323 , n5324 , n5325 , n5326 , n5327 , n5328 , n5329 , n5330 , n5331 , n5332 , n5333 , n5334 , n5335 , n5336 , n5337 , n5338 , n5339 , n5340 , n5341 , n5342 , n5343 , n5344 , n5345 , n5346 , n5347 , n5348 , n5349 , n5350 , n5351 , n5352 , n5353 , n5354 , n5355 , n5356 , n5357 , n5358 , n5359 , n5360 , n5361 , n5362 , n5363 , n5364 , n5365 , n5366 , n5367 , n5368 , n5369 , n5370 , n5371 , n5372 , n5373 , n5374 , n5375 , n5376 , n5377 , n5378 , n5379 , n5380 , n5381 , n5382 , n5383 , n5384 , n5385 , n5386 , n5387 , n5388 , n5389 , n5390 , n5391 , n5392 , n5393 , n5394 , n5395 , n5396 , n5397 , n5398 , n5399 , n5400 , n5401 , n5402 , n5403 , n5404 , n5405 , n5406 , n5407 , n5408 , n5409 , n5410 , n5411 , n5412 , n5413 , n5414 , n5415 , n5416 , n5417 , n5418 , n5419 , n5420 , n5421 , n5422 , n5423 , n5424 , n5425 , n5426 , n5427 , n5428 , n5429 , n5430 , n5431 , n5432 , n5433 , n5434 , n5435 , n5436 , n5437 , n5438 , n5439 , n5440 , n5441 , n5442 , n5443 , n5444 , n5445 , n5446 , n5447 , n5448 , n5449 , n5450 , n5451 , n5452 , n5453 , n5454 , n5455 , n5456 , n5457 , n5458 , n5459 , n5460 , n5461 , n5462 , n5463 , n5464 , n5465 , n5466 , n5467 , n5468 , n5469 , n5470 , n5471 , n5472 , n5473 , n5474 , n5475 , n5476 , n5477 , n5478 , n5479 , n5480 , n5481 , n5482 , n5483 , n5484 , n5485 , n5486 , n5487 , n5488 , n5489 , n5490 , n5491 , n5492 , n5493 , n5494 , n5495 , n5496 , n5497 , n5498 , n5499 , n5500 , n5501 , n5502 , n5503 , n5504 , n5505 , n5506 , n5507 , n5508 , n5509 , n5510 , n5511 , n5512 , n5513 , n5514 , n5515 , n5516 , n5517 , n5518 , n5519 , n5520 , n5521 , n5522 , n5523 , n5524 , n5525 , n5526 , n5527 , n5528 , n5529 , n5530 , n5531 , n5532 , n5533 , n5534 , n5535 , n5536 , n5537 , n5538 , n5539 , n5540 , n5541 , n5542 , n5543 , n5544 , n5545 , n5546 , n5547 , n5548 , n5549 , n5550 , n5551 , n5552 , n5553 , n5554 , n5555 , n5556 , n5557 , n5558 , n5559 , n5560 , n5561 , n5562 , n5563 , n5564 , n5565 , n5566 , n5567 , n5568 , n5569 , n5570 , n5571 , n5572 , n5573 , n5574 , n5575 , n5576 , n5577 , n5578 , n5579 , n5580 , n5581 , n5582 , n5583 , n5584 , n5585 , n5586 , n5587 , n5588 , n5589 , n5590 , n5591 , n5592 , n5593 , n5594 , n5595 , n5596 , n5597 , n5598 , n5599 , n5600 , n5601 , n5602 , n5603 , n5604 , n5605 , n5606 , n5607 , n5608 , n5609 , n5610 , n5611 , n5612 , n5613 , n5614 , n5615 , n5616 , n5617 , n5618 , n5619 , n5620 , n5621 , n5622 , n5623 , n5624 , n5625 , n5626 , n5627 , n5628 , n5629 , n5630 , n5631 , n5632 , n5633 , n5634 , n5635 , n5636 , n5637 , n5638 , n5639 , n5640 , n5641 , n5642 , n5643 , n5644 , n5645 , n5646 , n5647 , n5648 , n5649 , n5650 , n5651 , n5652 , n5653 , n5654 , n5655 , n5656 , n5657 , n5658 , n5659 , n5660 , n5661 , n5662 , n5663 , n5664 , n5665 , n5666 , n5667 , n5668 , n5669 , n5670 , n5671 , n5672 , n5673 , n5674 , n5675 , n5676 , n5677 , n5678 , n5679 , n5680 , n5681 , n5682 , n5683 , n5684 , n5685 , n5686 , n5687 , n5688 , n5689 , n5690 , n5691 , n5692 , n5693 , n5694 , n5695 , n5696 , n5697 , n5698 , n5699 , n5700 , n5701 , n5702 , n5703 , n5704 , n5705 , n5706 , n5707 , n5708 , n5709 , n5710 , n5711 , n5712 , n5713 , n5714 , n5715 , n5716 , n5717 , n5718 , n5719 , n5720 , n5721 , n5722 , n5723 , n5724 , n5725 , n5726 , n5727 , n5728 , n5729 , n5730 , n5731 , n5732 , n5733 , n5734 , n5735 , n5736 , n5737 , n5738 , n5739 , n5740 , n5741 , n5742 , n5743 , n5744 , n5745 , n5746 , n5747 , n5748 , n5749 , n5750 , n5751 , n5752 , n5753 , n5754 , n5755 , n5756 , n5757 , n5758 , n5759 , n5760 , n5761 , n5762 , n5763 , n5764 , n5765 , n5766 , n5767 , n5768 , n5769 , n5770 , n5771 , n5772 , n5773 , n5774 , n5775 , n5776 , n5777 , n5778 , n5779 , n5780 , n5781 , n5782 , n5783 , n5784 , n5785 , n5786 , n5787 , n5788 , n5789 , n5790 , n5791 , n5792 , n5793 , n5794 , n5795 , n5796 , n5797 , n5798 , n5799 , n5800 , n5801 , n5802 , n5803 , n5804 , n5805 , n5806 , n5807 , n5808 , n5809 , n5810 , n5811 , n5812 , n5813 , n5814 , n5815 , n5816 , n5817 , n5818 , n5819 , n5820 , n5821 , n5822 , n5823 , n5824 , n5825 , n5826 , n5827 , n5828 , n5829 , n5830 , n5831 , n5832 , n5833 , n5834 , n5835 , n5836 , n5837 , n5838 , n5839 , n5840 , n5841 , n5842 , n5843 , n5844 , n5845 , n5846 , n5847 , n5848 , n5849 , n5850 , n5851 , n5852 , n5853 , n5854 , n5855 , n5856 , n5857 , n5858 , n5859 , n5860 , n5861 , n5862 , n5863 , n5864 , n5865 , n5866 , n5867 , n5868 , n5869 , n5870 , n5871 , n5872 , n5873 , n5874 , n5875 , n5876 , n5877 , n5878 , n5879 , n5880 , n5881 , n5882 , n5883 , n5884 , n5885 , n5886 , n5887 , n5888 , n5889 , n5890 , n5891 , n5892 , n5893 , n5894 , n5895 , n5896 , n5897 , n5898 , n5899 , n5900 , n5901 , n5902 , n5903 , n5904 , n5905 , n5906 , n5907 , n5908 , n5909 , n5910 , n5911 , n5912 , n5913 , n5914 , n5915 , n5916 , n5917 , n5918 , n5919 , n5920 , n5921 , n5922 , n5923 , n5924 , n5925 , n5926 , n5927 , n5928 , n5929 , n5930 , n5931 , n5932 , n5933 , n5934 , n5935 , n5936 , n5937 , n5938 , n5939 , n5940 , n5941 , n5942 , n5943 , n5944 , n5945 , n5946 , n5947 , n5948 , n5949 , n5950 , n5951 , n5952 , n5953 , n5954 , n5955 , n5956 , n5957 , n5958 , n5959 , n5960 , n5961 , n5962 , n5963 , n5964 , n5965 , n5966 , n5967 , n5968 , n5969 , n5970 , n5971 , n5972 , n5973 , n5974 , n5975 , n5976 , n5977 , n5978 , n5979 , n5980 , n5981 , n5982 , n5983 , n5984 , n5985 , n5986 , n5987 , n5988 , n5989 , n5990 , n5991 , n5992 , n5993 , n5994 , n5995 , n5996 , n5997 , n5998 , n5999 , n6000 , n6001 , n6002 , n6003 , n6004 , n6005 , n6006 , n6007 , n6008 , n6009 , n6010 , n6011 , n6012 , n6013 , n6014 , n6015 , n6016 , n6017 , n6018 , n6019 , n6020 , n6021 , n6022 , n6023 , n6024 , n6025 , n6026 , n6027 , n6028 , n6029 , n6030 , n6031 , n6032 , n6033 , n6034 , n6035 , n6036 , n6037 , n6038 , n6039 , n6040 , n6041 , n6042 , n6043 , n6044 , n6045 , n6046 , n6047 , n6048 , n6049 , n6050 , n6051 , n6052 , n6053 , n6054 , n6055 , n6056 , n6057 , n6058 , n6059 , n6060 , n6061 , n6062 , n6063 , n6064 , n6065 , n6066 , n6067 , n6068 , n6069 , n6070 , n6071 , n6072 , n6073 , n6074 , n6075 , n6076 , n6077 , n6078 , n6079 , n6080 , n6081 , n6082 , n6083 , n6084 , n6085 , n6086 , n6087 , n6088 , n6089 , n6090 , n6091 , n6092 , n6093 , n6094 , n6095 , n6096 , n6097 , n6098 , n6099 , n6100 , n6101 , n6102 , n6103 , n6104 , n6105 , n6106 , n6107 , n6108 , n6109 , n6110 , n6111 , n6112 , n6113 , n6114 , n6115 , n6116 , n6117 , n6118 , n6119 , n6120 , n6121 , n6122 , n6123 , n6124 , n6125 , n6126 , n6127 , n6128 , n6129 , n6130 , n6131 , n6132 , n6133 , n6134 , n6135 , n6136 , n6137 , n6138 , n6139 , n6140 , n6141 , n6142 , n6143 , n6144 , n6145 , n6146 , n6147 , n6148 , n6149 , n6150 , n6151 , n6152 , n6153 , n6154 , n6155 , n6156 , n6157 , n6158 , n6159 , n6160 , n6161 , n6162 , n6163 , n6164 , n6165 , n6166 , n6167 , n6168 , n6169 , n6170 , n6171 , n6172 , n6173 , n6174 , n6175 , n6176 , n6177 , n6178 , n6179 , n6180 , n6181 , n6182 , n6183 , n6184 , n6185 , n6186 , n6187 , n6188 , n6189 , n6190 , n6191 , n6192 , n6193 , n6194 , n6195 , n6196 , n6197 , n6198 , n6199 , n6200 , n6201 , n6202 , n6203 , n6204 , n6205 , n6206 , n6207 , n6208 , n6209 , n6210 , n6211 , n6212 , n6213 , n6214 , n6215 , n6216 , n6217 , n6218 , n6219 , n6220 , n6221 , n6222 , n6223 , n6224 , n6225 , n6226 , n6227 , n6228 , n6229 , n6230 , n6231 , n6232 , n6233 , n6234 , n6235 , n6236 , n6237 , n6238 , n6239 , n6240 , n6241 , n6242 , n6243 , n6244 , n6245 , n6246 , n6247 , n6248 , n6249 , n6250 , n6251 , n6252 , n6253 , n6254 , n6255 , n6256 , n6257 , n6258 , n6259 , n6260 , n6261 , n6262 , n6263 , n6264 , n6265 , n6266 , n6267 , n6268 , n6269 , n6270 , n6271 , n6272 , n6273 , n6274 , n6275 , n6276 , n6277 , n6278 , n6279 , n6280 , n6281 , n6282 , n6283 , n6284 , n6285 , n6286 , n6287 , n6288 , n6289 , n6290 , n6291 , n6292 , n6293 , n6294 , n6295 , n6296 , n6297 , n6298 , n6299 , n6300 , n6301 , n6302 , n6303 , n6304 , n6305 , n6306 , n6307 , n6308 , n6309 , n6310 , n6311 , n6312 , n6313 , n6314 , n6315 , n6316 , n6317 , n6318 , n6319 , n6320 , n6321 , n6322 , n6323 , n6324 , n6325 , n6326 , n6327 , n6328 , n6329 , n6330 , n6331 , n6332 , n6333 , n6334 , n6335 , n6336 , n6337 , n6338 , n6339 , n6340 , n6341 , n6342 , n6343 , n6344 , n6345 , n6346 , n6347 , n6348 , n6349 , n6350 , n6351 , n6352 , n6353 , n6354 , n6355 , n6356 , n6357 , n6358 , n6359 , n6360 , n6361 , n6362 , n6363 , n6364 , n6365 , n6366 , n6367 , n6368 , n6369 , n6370 , n6371 , n6372 , n6373 , n6374 , n6375 , n6376 , n6377 , n6378 , n6379 , n6380 , n6381 , n6382 , n6383 , n6384 , n6385 , n6386 , n6387 , n6388 , n6389 , n6390 , n6391 , n6392 , n6393 , n6394 , n6395 , n6396 , n6397 , n6398 , n6399 , n6400 , n6401 , n6402 , n6403 , n6404 , n6405 , n6406 , n6407 , n6408 , n6409 , n6410 , n6411 , n6412 , n6413 , n6414 , n6415 , n6416 , n6417 , n6418 , n6419 , n6420 , n6421 , n6422 , n6423 , n6424 , n6425 , n6426 , n6427 , n6428 , n6429 , n6430 , n6431 , n6432 , n6433 , n6434 , n6435 , n6436 , n6437 , n6438 , n6439 , n6440 , n6441 , n6442 , n6443 , n6444 , n6445 , n6446 , n6447 , n6448 , n6449 , n6450 , n6451 , n6452 , n6453 , n6454 , n6455 , n6456 , n6457 , n6458 , n6459 , n6460 , n6461 , n6462 , n6463 , n6464 , n6465 , n6466 , n6467 , n6468 , n6469 , n6470 , n6471 , n6472 , n6473 , n6474 , n6475 , n6476 , n6477 , n6478 , n6479 , n6480 , n6481 , n6482 , n6483 , n6484 , n6485 , n6486 , n6487 , n6488 , n6489 , n6490 , n6491 , n6492 , n6493 , n6494 , n6495 , n6496 , n6497 , n6498 , n6499 , n6500 , n6501 , n6502 , n6503 , n6504 , n6505 , n6506 , n6507 , n6508 , n6509 , n6510 , n6511 , n6512 , n6513 , n6514 , n6515 , n6516 , n6517 , n6518 , n6519 , n6520 , n6521 , n6522 , n6523 , n6524 , n6525 , n6526 , n6527 , n6528 , n6529 , n6530 , n6531 , n6532 , n6533 , n6534 , n6535 , n6536 , n6537 , n6538 , n6539 , n6540 , n6541 , n6542 , n6543 , n6544 , n6545 , n6546 , n6547 , n6548 , n6549 , n6550 , n6551 , n6552 , n6553 , n6554 , n6555 , n6556 , n6557 , n6558 , n6559 , n6560 , n6561 , n6562 , n6563 , n6564 , n6565 , n6566 , n6567 , n6568 , n6569 , n6570 , n6571 , n6572 , n6573 , n6574 , n6575 , n6576 , n6577 , n6578 , n6579 , n6580 , n6581 , n6582 , n6583 , n6584 , n6585 , n6586 , n6587 , n6588 , n6589 , n6590 , n6591 , n6592 , n6593 , n6594 , n6595 , n6596 , n6597 , n6598 , n6599 , n6600 , n6601 , n6602 , n6603 , n6604 , n6605 , n6606 , n6607 , n6608 , n6609 , n6610 , n6611 , n6612 , n6613 , n6614 , n6615 , n6616 , n6617 , n6618 , n6619 , n6620 , n6621 , n6622 , n6623 , n6624 , n6625 , n6626 , n6627 , n6628 , n6629 , n6630 , n6631 , n6632 , n6633 , n6634 , n6635 , n6636 , n6637 , n6638 , n6639 , n6640 , n6641 , n6642 , n6643 , n6644 , n6645 , n6646 , n6647 , n6648 , n6649 , n6650 , n6651 , n6652 , n6653 , n6654 , n6655 , n6656 , n6657 , n6658 , n6659 , n6660 , n6661 , n6662 , n6663 , n6664 , n6665 , n6666 , n6667 , n6668 , n6669 , n6670 , n6671 , n6672 , n6673 , n6674 , n6675 , n6676 , n6677 , n6678 , n6679 , n6680 , n6681 , n6682 , n6683 , n6684 , n6685 , n6686 , n6687 , n6688 , n6689 , n6690 , n6691 , n6692 , n6693 , n6694 , n6695 , n6696 , n6697 , n6698 , n6699 , n6700 , n6701 , n6702 , n6703 , n6704 , n6705 , n6706 , n6707 , n6708 , n6709 , n6710 , n6711 , n6712 , n6713 , n6714 , n6715 , n6716 , n6717 , n6718 , n6719 , n6720 , n6721 , n6722 , n6723 , n6724 , n6725 , n6726 , n6727 , n6728 , n6729 , n6730 , n6731 , n6732 , n6733 , n6734 , n6735 , n6736 , n6737 , n6738 , n6739 , n6740 , n6741 , n6742 , n6743 , n6744 , n6745 , n6746 , n6747 , n6748 , n6749 , n6750 , n6751 , n6752 , n6753 , n6754 , n6755 , n6756 , n6757 , n6758 , n6759 , n6760 , n6761 , n6762 , n6763 , n6764 , n6765 , n6766 , n6767 , n6768 , n6769 , n6770 , n6771 , n6772 , n6773 , n6774 , n6775 , n6776 , n6777 , n6778 , n6779 , n6780 , n6781 , n6782 , n6783 , n6784 , n6785 , n6786 , n6787 , n6788 , n6789 , n6790 , n6791 , n6792 , n6793 , n6794 , n6795 , n6796 , n6797 , n6798 , n6799 , n6800 , n6801 , n6802 , n6803 , n6804 , n6805 , n6806 , n6807 , n6808 , n6809 , n6810 , n6811 , n6812 , n6813 , n6814 , n6815 , n6816 , n6817 , n6818 , n6819 , n6820 , n6821 , n6822 , n6823 , n6824 , n6825 , n6826 , n6827 , n6828 , n6829 , n6830 , n6831 , n6832 , n6833 , n6834 , n6835 , n6836 , n6837 , n6838 , n6839 , n6840 , n6841 , n6842 , n6843 , n6844 , n6845 , n6846 , n6847 , n6848 , n6849 , n6850 , n6851 , n6852 , n6853 , n6854 , n6855 , n6856 , n6857 , n6858 , n6859 , n6860 , n6861 , n6862 , n6863 , n6864 , n6865 , n6866 , n6867 , n6868 , n6869 , n6870 , n6871 , n6872 , n6873 , n6874 , n6875 , n6876 , n6877 , n6878 , n6879 , n6880 , n6881 , n6882 , n6883 , n6884 , n6885 , n6886 , n6887 , n6888 , n6889 , n6890 , n6891 , n6892 , n6893 , n6894 , n6895 , n6896 , n6897 , n6898 , n6899 , n6900 , n6901 , n6902 , n6903 , n6904 , n6905 , n6906 , n6907 , n6908 , n6909 , n6910 , n6911 , n6912 , n6913 , n6914 , n6915 , n6916 , n6917 , n6918 , n6919 , n6920 , n6921 , n6922 , n6923 , n6924 , n6925 , n6926 , n6927 , n6928 , n6929 , n6930 , n6931 , n6932 , n6933 , n6934 , n6935 , n6936 , n6937 , n6938 , n6939 , n6940 , n6941 , n6942 , n6943 , n6944 , n6945 , n6946 , n6947 , n6948 , n6949 , n6950 , n6951 , n6952 , n6953 , n6954 , n6955 , n6956 , n6957 , n6958 , n6959 , n6960 , n6961 , n6962 , n6963 , n6964 , n6965 , n6966 , n6967 , n6968 , n6969 , n6970 , n6971 , n6972 , n6973 , n6974 , n6975 , n6976 , n6977 , n6978 , n6979 , n6980 , n6981 , n6982 , n6983 , n6984 , n6985 , n6986 , n6987 , n6988 , n6989 , n6990 , n6991 , n6992 , n6993 , n6994 , n6995 , n6996 , n6997 , n6998 , n6999 , n7000 , n7001 , n7002 , n7003 , n7004 , n7005 , n7006 , n7007 , n7008 , n7009 , n7010 , n7011 , n7012 , n7013 , n7014 , n7015 , n7016 , n7017 , n7018 , n7019 , n7020 , n7021 , n7022 , n7023 , n7024 , n7025 , n7026 , n7027 , n7028 , n7029 , n7030 , n7031 , n7032 , n7033 , n7034 , n7035 , n7036 , n7037 , n7038 , n7039 , n7040 , n7041 , n7042 , n7043 , n7044 , n7045 , n7046 , n7047 , n7048 , n7049 , n7050 , n7051 , n7052 , n7053 , n7054 , n7055 , n7056 , n7057 , n7058 , n7059 , n7060 , n7061 , n7062 , n7063 , n7064 , n7065 , n7066 , n7067 , n7068 , n7069 , n7070 , n7071 , n7072 , n7073 , n7074 , n7075 , n7076 , n7077 , n7078 , n7079 , n7080 , n7081 , n7082 , n7083 , n7084 , n7085 , n7086 , n7087 , n7088 , n7089 , n7090 , n7091 , n7092 , n7093 , n7094 , n7095 , n7096 , n7097 , n7098 , n7099 , n7100 , n7101 , n7102 , n7103 , n7104 , n7105 , n7106 , n7107 , n7108 , n7109 , n7110 , n7111 , n7112 , n7113 , n7114 , n7115 , n7116 , n7117 , n7118 , n7119 , n7120 , n7121 , n7122 , n7123 , n7124 , n7125 , n7126 , n7127 , n7128 , n7129 , n7130 , n7131 , n7132 , n7133 , n7134 , n7135 , n7136 , n7137 , n7138 , n7139 , n7140 , n7141 , n7142 , n7143 , n7144 , n7145 , n7146 , n7147 , n7148 , n7149 , n7150 , n7151 , n7152 , n7153 , n7154 , n7155 , n7156 , n7157 , n7158 , n7159 , n7160 , n7161 , n7162 , n7163 , n7164 , n7165 , n7166 , n7167 , n7168 , n7169 , n7170 , n7171 , n7172 , n7173 , n7174 , n7175 , n7176 , n7177 , n7178 , n7179 , n7180 , n7181 , n7182 , n7183 , n7184 , n7185 , n7186 , n7187 , n7188 , n7189 , n7190 , n7191 , n7192 , n7193 , n7194 , n7195 , n7196 , n7197 , n7198 , n7199 , n7200 , n7201 , n7202 , n7203 , n7204 , n7205 , n7206 , n7207 , n7208 , n7209 , n7210 , n7211 , n7212 , n7213 , n7214 , n7215 , n7216 , n7217 , n7218 , n7219 , n7220 , n7221 , n7222 , n7223 , n7224 , n7225 , n7226 , n7227 , n7228 , n7229 , n7230 , n7231 , n7232 , n7233 , n7234 , n7235 , n7236 , n7237 , n7238 , n7239 , n7240 , n7241 , n7242 , n7243 , n7244 , n7245 , n7246 , n7247 , n7248 , n7249 , n7250 , n7251 , n7252 , n7253 , n7254 , n7255 , n7256 , n7257 , n7258 , n7259 , n7260 , n7261 , n7262 , n7263 , n7264 , n7265 , n7266 , n7267 , n7268 , n7269 , n7270 , n7271 , n7272 , n7273 , n7274 , n7275 , n7276 , n7277 , n7278 , n7279 , n7280 , n7281 , n7282 , n7283 , n7284 , n7285 , n7286 , n7287 , n7288 , n7289 , n7290 , n7291 , n7292 , n7293 , n7294 , n7295 , n7296 , n7297 , n7298 , n7299 , n7300 , n7301 , n7302 , n7303 , n7304 , n7305 , n7306 , n7307 , n7308 , n7309 , n7310 , n7311 , n7312 , n7313 , n7314 , n7315 , n7316 , n7317 , n7318 , n7319 , n7320 , n7321 , n7322 , n7323 , n7324 , n7325 , n7326 , n7327 , n7328 , n7329 , n7330 , n7331 , n7332 , n7333 , n7334 , n7335 , n7336 , n7337 , n7338 , n7339 , n7340 , n7341 , n7342 , n7343 , n7344 , n7345 , n7346 , n7347 , n7348 , n7349 , n7350 , n7351 , n7352 , n7353 , n7354 , n7355 , n7356 , n7357 , n7358 , n7359 , n7360 , n7361 , n7362 , n7363 , n7364 , n7365 , n7366 , n7367 , n7368 , n7369 , n7370 , n7371 , n7372 , n7373 , n7374 , n7375 , n7376 , n7377 , n7378 , n7379 , n7380 , n7381 , n7382 , n7383 , n7384 , n7385 , n7386 , n7387 , n7388 , n7389 , n7390 , n7391 , n7392 , n7393 , n7394 , n7395 , n7396 , n7397 , n7398 , n7399 , n7400 , n7401 , n7402 , n7403 , n7404 , n7405 , n7406 , n7407 , n7408 , n7409 , n7410 , n7411 , n7412 , n7413 , n7414 , n7415 , n7416 , n7417 , n7418 , n7419 , n7420 , n7421 , n7422 , n7423 , n7424 , n7425 , n7426 , n7427 , n7428 , n7429 , n7430 , n7431 , n7432 , n7433 , n7434 , n7435 , n7436 , n7437 , n7438 , n7439 , n7440 , n7441 , n7442 , n7443 , n7444 , n7445 , n7446 , n7447 , n7448 , n7449 , n7450 , n7451 , n7452 , n7453 , n7454 , n7455 , n7456 , n7457 , n7458 , n7459 , n7460 , n7461 , n7462 , n7463 , n7464 , n7465 , n7466 , n7467 , n7468 , n7469 , n7470 , n7471 , n7472 , n7473 , n7474 , n7475 , n7476 , n7477 , n7478 , n7479 , n7480 , n7481 , n7482 , n7483 , n7484 , n7485 , n7486 , n7487 , n7488 , n7489 , n7490 , n7491 , n7492 , n7493 , n7494 , n7495 , n7496 , n7497 , n7498 , n7499 , n7500 , n7501 , n7502 , n7503 , n7504 , n7505 , n7506 , n7507 , n7508 , n7509 , n7510 , n7511 , n7512 , n7513 , n7514 , n7515 , n7516 , n7517 , n7518 , n7519 , n7520 , n7521 , n7522 , n7523 , n7524 , n7525 , n7526 , n7527 , n7528 , n7529 , n7530 , n7531 , n7532 , n7533 , n7534 , n7535 , n7536 , n7537 , n7538 , n7539 , n7540 , n7541 , n7542 , n7543 , n7544 , n7545 , n7546 , n7547 , n7548 , n7549 , n7550 , n7551 , n7552 , n7553 , n7554 , n7555 , n7556 , n7557 , n7558 , n7559 , n7560 , n7561 , n7562 , n7563 , n7564 , n7565 , n7566 , n7567 , n7568 , n7569 , n7570 , n7571 , n7572 , n7573 , n7574 , n7575 , n7576 , n7577 , n7578 , n7579 , n7580 , n7581 , n7582 , n7583 , n7584 , n7585 , n7586 , n7587 , n7588 , n7589 , n7590 , n7591 , n7592 , n7593 , n7594 , n7595 , n7596 , n7597 , n7598 , n7599 , n7600 , n7601 , n7602 , n7603 , n7604 , n7605 , n7606 , n7607 , n7608 , n7609 , n7610 , n7611 , n7612 , n7613 , n7614 , n7615 , n7616 , n7617 , n7618 , n7619 , n7620 , n7621 , n7622 , n7623 , n7624 , n7625 , n7626 , n7627 , n7628 , n7629 , n7630 , n7631 , n7632 , n7633 , n7634 , n7635 , n7636 , n7637 , n7638 , n7639 , n7640 , n7641 , n7642 , n7643 , n7644 , n7645 , n7646 , n7647 , n7648 , n7649 , n7650 , n7651 , n7652 , n7653 , n7654 , n7655 , n7656 , n7657 , n7658 , n7659 , n7660 , n7661 , n7662 , n7663 , n7664 , n7665 , n7666 , n7667 , n7668 , n7669 , n7670 , n7671 , n7672 , n7673 , n7674 , n7675 , n7676 , n7677 , n7678 , n7679 , n7680 , n7681 , n7682 , n7683 , n7684 , n7685 , n7686 , n7687 , n7688 , n7689 , n7690 , n7691 , n7692 , n7693 , n7694 , n7695 , n7696 , n7697 , n7698 , n7699 , n7700 , n7701 , n7702 , n7703 , n7704 , n7705 , n7706 , n7707 , n7708 , n7709 , n7710 , n7711 , n7712 , n7713 , n7714 , n7715 , n7716 , n7717 , n7718 , n7719 , n7720 , n7721 , n7722 , n7723 , n7724 , n7725 , n7726 , n7727 , n7728 , n7729 , n7730 , n7731 , n7732 , n7733 , n7734 , n7735 , n7736 , n7737 , n7738 , n7739 , n7740 , n7741 , n7742 , n7743 , n7744 , n7745 , n7746 , n7747 , n7748 , n7749 , n7750 , n7751 , n7752 , n7753 , n7754 , n7755 , n7756 , n7757 , n7758 , n7759 , n7760 , n7761 , n7762 , n7763 , n7764 , n7765 , n7766 , n7767 , n7768 , n7769 , n7770 , n7771 , n7772 , n7773 , n7774 , n7775 , n7776 , n7777 , n7778 , n7779 , n7780 , n7781 , n7782 , n7783 , n7784 , n7785 , n7786 , n7787 , n7788 , n7789 , n7790 , n7791 , n7792 , n7793 , n7794 , n7795 , n7796 , n7797 , n7798 , n7799 , n7800 , n7801 , n7802 , n7803 , n7804 , n7805 , n7806 , n7807 , n7808 , n7809 , n7810 , n7811 , n7812 , n7813 , n7814 , n7815 , n7816 , n7817 , n7818 , n7819 , n7820 , n7821 , n7822 , n7823 , n7824 , n7825 , n7826 , n7827 , n7828 , n7829 , n7830 , n7831 , n7832 , n7833 , n7834 , n7835 , n7836 , n7837 , n7838 , n7839 , n7840 , n7841 , n7842 , n7843 , n7844 , n7845 , n7846 , n7847 , n7848 , n7849 , n7850 , n7851 , n7852 , n7853 , n7854 , n7855 , n7856 , n7857 , n7858 , n7859 , n7860 , n7861 , n7862 , n7863 , n7864 , n7865 , n7866 , n7867 , n7868 , n7869 , n7870 , n7871 , n7872 , n7873 , n7874 , n7875 , n7876 , n7877 , n7878 , n7879 , n7880 , n7881 , n7882 , n7883 , n7884 , n7885 , n7886 , n7887 , n7888 , n7889 , n7890 , n7891 , n7892 , n7893 , n7894 , n7895 , n7896 , n7897 , n7898 , n7899 , n7900 , n7901 , n7902 , n7903 , n7904 , n7905 , n7906 , n7907 , n7908 , n7909 , n7910 , n7911 , n7912 , n7913 , n7914 , n7915 , n7916 , n7917 , n7918 , n7919 , n7920 , n7921 , n7922 , n7923 , n7924 , n7925 , n7926 , n7927 , n7928 , n7929 , n7930 , n7931 , n7932 , n7933 , n7934 , n7935 , n7936 , n7937 , n7938 , n7939 , n7940 , n7941 , n7942 , n7943 , n7944 , n7945 , n7946 , n7947 , n7948 , n7949 , n7950 , n7951 , n7952 , n7953 , n7954 , n7955 , n7956 , n7957 , n7958 , n7959 , n7960 , n7961 , n7962 , n7963 , n7964 , n7965 , n7966 , n7967 , n7968 , n7969 , n7970 , n7971 , n7972 , n7973 , n7974 , n7975 , n7976 , n7977 , n7978 , n7979 , n7980 , n7981 , n7982 , n7983 , n7984 , n7985 , n7986 , n7987 , n7988 , n7989 , n7990 , n7991 , n7992 , n7993 , n7994 , n7995 , n7996 , n7997 , n7998 , n7999 , n8000 , n8001 , n8002 , n8003 , n8004 , n8005 , n8006 , n8007 , n8008 , n8009 , n8010 , n8011 , n8012 , n8013 , n8014 , n8015 , n8016 , n8017 , n8018 , n8019 , n8020 , n8021 , n8022 , n8023 , n8024 , n8025 , n8026 , n8027 , n8028 , n8029 , n8030 , n8031 , n8032 , n8033 , n8034 , n8035 , n8036 , n8037 , n8038 , n8039 , n8040 , n8041 , n8042 , n8043 , n8044 , n8045 , n8046 , n8047 , n8048 , n8049 , n8050 , n8051 , n8052 , n8053 , n8054 , n8055 , n8056 , n8057 , n8058 , n8059 , n8060 , n8061 , n8062 , n8063 , n8064 , n8065 , n8066 , n8067 , n8068 , n8069 , n8070 , n8071 , n8072 , n8073 , n8074 , n8075 , n8076 , n8077 , n8078 , n8079 , n8080 , n8081 , n8082 , n8083 , n8084 , n8085 , n8086 , n8087 , n8088 , n8089 , n8090 , n8091 , n8092 , n8093 , n8094 , n8095 , n8096 , n8097 , n8098 , n8099 , n8100 , n8101 , n8102 , n8103 , n8104 , n8105 , n8106 , n8107 , n8108 , n8109 , n8110 , n8111 , n8112 , n8113 , n8114 , n8115 , n8116 , n8117 , n8118 , n8119 , n8120 , n8121 , n8122 , n8123 , n8124 , n8125 , n8126 , n8127 , n8128 , n8129 , n8130 , n8131 , n8132 , n8133 , n8134 , n8135 , n8136 , n8137 , n8138 , n8139 , n8140 , n8141 , n8142 , n8143 , n8144 , n8145 , n8146 , n8147 , n8148 , n8149 , n8150 , n8151 , n8152 , n8153 , n8154 , n8155 , n8156 , n8157 , n8158 , n8159 , n8160 , n8161 , n8162 , n8163 , n8164 , n8165 , n8166 , n8167 , n8168 , n8169 , n8170 , n8171 , n8172 , n8173 , n8174 , n8175 , n8176 , n8177 , n8178 , n8179 , n8180 , n8181 , n8182 , n8183 , n8184 , n8185 , n8186 , n8187 , n8188 , n8189 , n8190 , n8191 , n8192 , n8193 , n8194 , n8195 , n8196 , n8197 , n8198 , n8199 , n8200 , n8201 , n8202 , n8203 , n8204 , n8205 , n8206 , n8207 , n8208 , n8209 , n8210 , n8211 , n8212 , n8213 , n8214 , n8215 , n8216 , n8217 , n8218 , n8219 , n8220 , n8221 , n8222 , n8223 , n8224 , n8225 , n8226 , n8227 , n8228 , n8229 , n8230 , n8231 , n8232 , n8233 , n8234 , n8235 , n8236 , n8237 , n8238 , n8239 , n8240 , n8241 , n8242 , n8243 , n8244 , n8245 , n8246 , n8247 , n8248 , n8249 , n8250 , n8251 , n8252 , n8253 , n8254 , n8255 , n8256 , n8257 , n8258 , n8259 , n8260 , n8261 , n8262 , n8263 , n8264 , n8265 , n8266 , n8267 , n8268 , n8269 , n8270 , n8271 , n8272 , n8273 , n8274 , n8275 , n8276 , n8277 , n8278 , n8279 , n8280 , n8281 , n8282 , n8283 , n8284 , n8285 , n8286 , n8287 , n8288 , n8289 , n8290 , n8291 , n8292 , n8293 , n8294 , n8295 , n8296 , n8297 , n8298 , n8299 , n8300 , n8301 , n8302 , n8303 , n8304 , n8305 , n8306 , n8307 , n8308 , n8309 , n8310 , n8311 , n8312 , n8313 , n8314 , n8315 , n8316 , n8317 , n8318 , n8319 , n8320 , n8321 , n8322 , n8323 , n8324 , n8325 , n8326 , n8327 , n8328 , n8329 , n8330 , n8331 , n8332 , n8333 , n8334 , n8335 , n8336 , n8337 , n8338 , n8339 , n8340 , n8341 , n8342 , n8343 , n8344 , n8345 , n8346 , n8347 , n8348 , n8349 , n8350 , n8351 , n8352 , n8353 , n8354 , n8355 , n8356 , n8357 , n8358 , n8359 , n8360 , n8361 , n8362 , n8363 , n8364 , n8365 , n8366 , n8367 , n8368 , n8369 , n8370 , n8371 , n8372 , n8373 , n8374 , n8375 , n8376 , n8377 , n8378 , n8379 , n8380 , n8381 , n8382 , n8383 , n8384 , n8385 , n8386 , n8387 , n8388 , n8389 , n8390 , n8391 , n8392 , n8393 , n8394 , n8395 , n8396 , n8397 , n8398 , n8399 , n8400 , n8401 , n8402 , n8403 , n8404 , n8405 , n8406 , n8407 , n8408 , n8409 , n8410 , n8411 , n8412 , n8413 , n8414 , n8415 , n8416 , n8417 , n8418 , n8419 , n8420 , n8421 , n8422 , n8423 , n8424 , n8425 , n8426 , n8427 , n8428 , n8429 , n8430 , n8431 , n8432 , n8433 , n8434 , n8435 , n8436 , n8437 , n8438 , n8439 , n8440 , n8441 , n8442 , n8443 , n8444 , n8445 , n8446 , n8447 , n8448 , n8449 , n8450 , n8451 , n8452 , n8453 , n8454 , n8455 , n8456 , n8457 , n8458 , n8459 , n8460 , n8461 , n8462 , n8463 , n8464 , n8465 , n8466 , n8467 , n8468 , n8469 , n8470 , n8471 , n8472 , n8473 , n8474 , n8475 , n8476 , n8477 , n8478 , n8479 , n8480 , n8481 , n8482 , n8483 , n8484 , n8485 , n8486 , n8487 , n8488 , n8489 , n8490 , n8491 , n8492 , n8493 , n8494 , n8495 , n8496 , n8497 , n8498 , n8499 , n8500 , n8501 , n8502 , n8503 , n8504 , n8505 , n8506 , n8507 , n8508 , n8509 , n8510 , n8511 , n8512 , n8513 , n8514 , n8515 , n8516 , n8517 , n8518 , n8519 , n8520 , n8521 , n8522 , n8523 , n8524 , n8525 , n8526 , n8527 , n8528 , n8529 , n8530 , n8531 , n8532 , n8533 , n8534 , n8535 , n8536 , n8537 , n8538 , n8539 , n8540 , n8541 , n8542 , n8543 , n8544 , n8545 , n8546 , n8547 , n8548 , n8549 , n8550 , n8551 , n8552 , n8553 , n8554 , n8555 , n8556 , n8557 , n8558 , n8559 , n8560 , n8561 , n8562 , n8563 , n8564 , n8565 , n8566 , n8567 , n8568 , n8569 , n8570 , n8571 , n8572 , n8573 , n8574 , n8575 , n8576 , n8577 , n8578 , n8579 , n8580 , n8581 , n8582 , n8583 , n8584 , n8585 , n8586 , n8587 , n8588 , n8589 , n8590 , n8591 , n8592 , n8593 , n8594 , n8595 , n8596 , n8597 , n8598 , n8599 , n8600 , n8601 , n8602 , n8603 , n8604 , n8605 , n8606 , n8607 , n8608 , n8609 , n8610 , n8611 , n8612 , n8613 , n8614 , n8615 , n8616 , n8617 , n8618 , n8619 , n8620 , n8621 , n8622 , n8623 , n8624 , n8625 , n8626 , n8627 , n8628 , n8629 , n8630 , n8631 , n8632 , n8633 , n8634 , n8635 , n8636 , n8637 , n8638 , n8639 , n8640 , n8641 , n8642 , n8643 , n8644 , n8645 , n8646 , n8647 , n8648 , n8649 , n8650 , n8651 , n8652 , n8653 , n8654 , n8655 , n8656 , n8657 , n8658 , n8659 , n8660 , n8661 , n8662 , n8663 , n8664 , n8665 , n8666 , n8667 , n8668 , n8669 , n8670 , n8671 , n8672 , n8673 , n8674 , n8675 , n8676 , n8677 , n8678 , n8679 , n8680 , n8681 , n8682 , n8683 , n8684 , n8685 , n8686 , n8687 , n8688 , n8689 , n8690 , n8691 , n8692 , n8693 , n8694 , n8695 , n8696 , n8697 , n8698 , n8699 , n8700 , n8701 , n8702 , n8703 , n8704 , n8705 , n8706 , n8707 , n8708 , n8709 , n8710 , n8711 , n8712 , n8713 , n8714 , n8715 , n8716 , n8717 , n8718 , n8719 , n8720 , n8721 , n8722 , n8723 , n8724 , n8725 , n8726 , n8727 , n8728 , n8729 , n8730 , n8731 , n8732 , n8733 , n8734 , n8735 , n8736 , n8737 , n8738 , n8739 , n8740 , n8741 , n8742 , n8743 , n8744 , n8745 , n8746 , n8747 , n8748 , n8749 , n8750 , n8751 , n8752 , n8753 , n8754 , n8755 , n8756 , n8757 , n8758 , n8759 , n8760 , n8761 , n8762 , n8763 , n8764 , n8765 , n8766 , n8767 , n8768 , n8769 , n8770 , n8771 , n8772 , n8773 , n8774 , n8775 , n8776 , n8777 , n8778 , n8779 , n8780 , n8781 , n8782 , n8783 , n8784 , n8785 , n8786 , n8787 , n8788 , n8789 , n8790 , n8791 , n8792 , n8793 , n8794 , n8795 , n8796 , n8797 , n8798 , n8799 , n8800 , n8801 , n8802 , n8803 , n8804 , n8805 , n8806 , n8807 , n8808 , n8809 , n8810 , n8811 , n8812 , n8813 , n8814 , n8815 , n8816 , n8817 , n8818 , n8819 , n8820 , n8821 , n8822 , n8823 , n8824 , n8825 , n8826 , n8827 , n8828 , n8829 , n8830 , n8831 , n8832 , n8833 , n8834 , n8835 , n8836 , n8837 , n8838 , n8839 , n8840 , n8841 , n8842 , n8843 , n8844 , n8845 , n8846 , n8847 , n8848 , n8849 , n8850 , n8851 , n8852 , n8853 , n8854 , n8855 , n8856 , n8857 , n8858 , n8859 , n8860 , n8861 , n8862 , n8863 , n8864 , n8865 , n8866 , n8867 , n8868 , n8869 , n8870 , n8871 , n8872 , n8873 , n8874 , n8875 , n8876 , n8877 , n8878 , n8879 , n8880 , n8881 , n8882 , n8883 , n8884 , n8885 , n8886 , n8887 , n8888 , n8889 , n8890 , n8891 , n8892 , n8893 , n8894 , n8895 , n8896 , n8897 , n8898 , n8899 , n8900 , n8901 , n8902 , n8903 , n8904 , n8905 , n8906 , n8907 , n8908 , n8909 , n8910 , n8911 , n8912 , n8913 , n8914 , n8915 , n8916 , n8917 , n8918 , n8919 , n8920 , n8921 , n8922 , n8923 , n8924 , n8925 , n8926 , n8927 , n8928 , n8929 , n8930 , n8931 , n8932 , n8933 , n8934 , n8935 , n8936 , n8937 , n8938 , n8939 , n8940 , n8941 , n8942 , n8943 , n8944 , n8945 , n8946 , n8947 , n8948 , n8949 , n8950 , n8951 , n8952 , n8953 , n8954 , n8955 , n8956 , n8957 , n8958 , n8959 , n8960 , n8961 , n8962 , n8963 , n8964 , n8965 , n8966 , n8967 , n8968 , n8969 , n8970 , n8971 , n8972 , n8973 , n8974 , n8975 , n8976 , n8977 , n8978 , n8979 , n8980 , n8981 , n8982 , n8983 , n8984 , n8985 , n8986 , n8987 , n8988 , n8989 , n8990 , n8991 , n8992 , n8993 , n8994 , n8995 , n8996 , n8997 , n8998 , n8999 , n9000 , n9001 , n9002 , n9003 , n9004 , n9005 , n9006 , n9007 , n9008 , n9009 , n9010 , n9011 , n9012 , n9013 , n9014 , n9015 , n9016 , n9017 , n9018 , n9019 , n9020 , n9021 , n9022 , n9023 , n9024 , n9025 , n9026 , n9027 , n9028 , n9029 , n9030 , n9031 , n9032 , n9033 , n9034 , n9035 , n9036 , n9037 , n9038 , n9039 , n9040 , n9041 , n9042 , n9043 , n9044 , n9045 , n9046 , n9047 , n9048 , n9049 , n9050 , n9051 , n9052 , n9053 , n9054 , n9055 , n9056 , n9057 , n9058 , n9059 , n9060 , n9061 , n9062 , n9063 , n9064 , n9065 , n9066 , n9067 , n9068 , n9069 , n9070 , n9071 , n9072 , n9073 , n9074 , n9075 , n9076 , n9077 , n9078 , n9079 , n9080 , n9081 , n9082 , n9083 , n9084 , n9085 , n9086 , n9087 , n9088 , n9089 , n9090 , n9091 , n9092 , n9093 , n9094 , n9095 , n9096 , n9097 , n9098 , n9099 , n9100 , n9101 , n9102 , n9103 , n9104 , n9105 , n9106 , n9107 , n9108 , n9109 , n9110 , n9111 , n9112 , n9113 , n9114 , n9115 , n9116 , n9117 , n9118 , n9119 , n9120 , n9121 , n9122 , n9123 , n9124 , n9125 , n9126 , n9127 , n9128 , n9129 , n9130 , n9131 , n9132 , n9133 , n9134 , n9135 , n9136 , n9137 , n9138 , n9139 , n9140 , n9141 , n9142 , n9143 , n9144 , n9145 , n9146 , n9147 , n9148 , n9149 , n9150 , n9151 , n9152 , n9153 , n9154 , n9155 , n9156 , n9157 , n9158 , n9159 , n9160 , n9161 , n9162 , n9163 , n9164 , n9165 , n9166 , n9167 , n9168 , n9169 , n9170 , n9171 , n9172 , n9173 , n9174 , n9175 , n9176 , n9177 , n9178 , n9179 , n9180 , n9181 , n9182 , n9183 , n9184 , n9185 , n9186 , n9187 , n9188 , n9189 , n9190 , n9191 , n9192 , n9193 , n9194 , n9195 , n9196 , n9197 , n9198 , n9199 , n9200 , n9201 , n9202 , n9203 , n9204 , n9205 , n9206 , n9207 , n9208 , n9209 , n9210 , n9211 , n9212 , n9213 , n9214 , n9215 , n9216 , n9217 , n9218 , n9219 , n9220 , n9221 , n9222 , n9223 , n9224 , n9225 , n9226 , n9227 , n9228 , n9229 , n9230 , n9231 , n9232 , n9233 , n9234 , n9235 , n9236 , n9237 , n9238 , n9239 , n9240 , n9241 , n9242 , n9243 , n9244 , n9245 , n9246 , n9247 , n9248 , n9249 , n9250 , n9251 , n9252 , n9253 , n9254 , n9255 , n9256 , n9257 , n9258 , n9259 , n9260 , n9261 , n9262 , n9263 , n9264 , n9265 , n9266 , n9267 , n9268 , n9269 , n9270 , n9271 , n9272 , n9273 , n9274 , n9275 , n9276 , n9277 , n9278 , n9279 , n9280 , n9281 , n9282 , n9283 , n9284 , n9285 , n9286 , n9287 , n9288 , n9289 , n9290 , n9291 , n9292 , n9293 , n9294 , n9295 , n9296 , n9297 , n9298 , n9299 , n9300 , n9301 , n9302 , n9303 , n9304 , n9305 , n9306 , n9307 , n9308 , n9309 , n9310 , n9311 , n9312 , n9313 , n9314 , n9315 , n9316 , n9317 , n9318 , n9319 , n9320 , n9321 , n9322 , n9323 , n9324 , n9325 , n9326 , n9327 , n9328 , n9329 , n9330 , n9331 , n9332 , n9333 , n9334 , n9335 , n9336 , n9337 , n9338 , n9339 , n9340 , n9341 , n9342 , n9343 , n9344 , n9345 , n9346 , n9347 , n9348 , n9349 , n9350 , n9351 , n9352 , n9353 , n9354 , n9355 , n9356 , n9357 , n9358 , n9359 , n9360 , n9361 , n9362 , n9363 , n9364 , n9365 , n9366 , n9367 , n9368 , n9369 , n9370 , n9371 , n9372 , n9373 , n9374 , n9375 , n9376 , n9377 , n9378 , n9379 , n9380 , n9381 , n9382 , n9383 , n9384 , n9385 , n9386 , n9387 , n9388 , n9389 , n9390 , n9391 , n9392 , n9393 , n9394 , n9395 , n9396 , n9397 , n9398 , n9399 , n9400 , n9401 , n9402 , n9403 , n9404 , n9405 , n9406 , n9407 , n9408 , n9409 , n9410 , n9411 , n9412 , n9413 , n9414 , n9415 , n9416 , n9417 , n9418 , n9419 , n9420 , n9421 , n9422 , n9423 , n9424 , n9425 , n9426 , n9427 , n9428 , n9429 , n9430 , n9431 , n9432 , n9433 , n9434 , n9435 , n9436 , n9437 , n9438 , n9439 , n9440 , n9441 , n9442 , n9443 , n9444 , n9445 , n9446 , n9447 , n9448 , n9449 , n9450 , n9451 , n9452 , n9453 , n9454 , n9455 , n9456 , n9457 , n9458 , n9459 , n9460 , n9461 , n9462 , n9463 , n9464 , n9465 , n9466 , n9467 , n9468 , n9469 , n9470 , n9471 , n9472 , n9473 , n9474 , n9475 , n9476 , n9477 , n9478 , n9479 , n9480 , n9481 , n9482 , n9483 , n9484 , n9485 , n9486 , n9487 , n9488 , n9489 , n9490 , n9491 , n9492 , n9493 , n9494 , n9495 , n9496 , n9497 , n9498 , n9499 , n9500 , n9501 , n9502 , n9503 , n9504 , n9505 , n9506 , n9507 , n9508 , n9509 , n9510 , n9511 , n9512 , n9513 , n9514 , n9515 , n9516 , n9517 , n9518 , n9519 , n9520 , n9521 , n9522 , n9523 , n9524 , n9525 , n9526 , n9527 , n9528 , n9529 , n9530 , n9531 , n9532 , n9533 , n9534 , n9535 , n9536 , n9537 , n9538 , n9539 , n9540 , n9541 , n9542 , n9543 , n9544 , n9545 , n9546 , n9547 , n9548 , n9549 , n9550 , n9551 , n9552 , n9553 , n9554 , n9555 , n9556 , n9557 , n9558 , n9559 , n9560 , n9561 , n9562 , n9563 , n9564 , n9565 , n9566 , n9567 , n9568 , n9569 , n9570 , n9571 , n9572 , n9573 , n9574 , n9575 , n9576 , n9577 , n9578 , n9579 , n9580 , n9581 , n9582 , n9583 , n9584 , n9585 , n9586 , n9587 , n9588 , n9589 , n9590 , n9591 , n9592 , n9593 , n9594 , n9595 , n9596 , n9597 , n9598 , n9599 , n9600 , n9601 , n9602 , n9603 , n9604 , n9605 , n9606 , n9607 , n9608 , n9609 , n9610 , n9611 , n9612 , n9613 , n9614 , n9615 , n9616 , n9617 , n9618 , n9619 , n9620 , n9621 , n9622 , n9623 , n9624 , n9625 , n9626 , n9627 , n9628 , n9629 , n9630 , n9631 , n9632 , n9633 , n9634 , n9635 , n9636 , n9637 , n9638 , n9639 , n9640 , n9641 , n9642 , n9643 , n9644 , n9645 , n9646 , n9647 , n9648 , n9649 , n9650 , n9651 , n9652 , n9653 , n9654 , n9655 , n9656 , n9657 , n9658 , n9659 , n9660 , n9661 , n9662 , n9663 , n9664 , n9665 , n9666 , n9667 , n9668 , n9669 , n9670 , n9671 , n9672 , n9673 , n9674 , n9675 , n9676 , n9677 , n9678 , n9679 , n9680 , n9681 , n9682 , n9683 , n9684 , n9685 , n9686 , n9687 , n9688 , n9689 , n9690 , n9691 , n9692 , n9693 , n9694 , n9695 , n9696 , n9697 , n9698 , n9699 , n9700 , n9701 , n9702 , n9703 , n9704 , n9705 , n9706 , n9707 , n9708 , n9709 , n9710 , n9711 , n9712 , n9713 , n9714 , n9715 , n9716 , n9717 , n9718 , n9719 , n9720 , n9721 , n9722 , n9723 , n9724 , n9725 , n9726 , n9727 , n9728 , n9729 , n9730 , n9731 , n9732 , n9733 , n9734 , n9735 , n9736 , n9737 , n9738 , n9739 , n9740 , n9741 , n9742 , n9743 , n9744 , n9745 , n9746 , n9747 , n9748 , n9749 , n9750 , n9751 , n9752 , n9753 , n9754 , n9755 , n9756 , n9757 , n9758 , n9759 , n9760 , n9761 , n9762 , n9763 , n9764 , n9765 , n9766 , n9767 , n9768 , n9769 , n9770 , n9771 , n9772 , n9773 , n9774 , n9775 , n9776 , n9777 , n9778 , n9779 , n9780 , n9781 , n9782 , n9783 , n9784 , n9785 , n9786 , n9787 , n9788 , n9789 , n9790 , n9791 , n9792 , n9793 , n9794 , n9795 , n9796 , n9797 , n9798 , n9799 , n9800 , n9801 , n9802 , n9803 , n9804 , n9805 , n9806 , n9807 , n9808 , n9809 , n9810 , n9811 , n9812 , n9813 , n9814 , n9815 , n9816 , n9817 , n9818 , n9819 , n9820 , n9821 , n9822 , n9823 , n9824 , n9825 , n9826 , n9827 , n9828 , n9829 , n9830 , n9831 , n9832 , n9833 , n9834 , n9835 , n9836 , n9837 , n9838 , n9839 , n9840 , n9841 , n9842 , n9843 , n9844 , n9845 , n9846 , n9847 , n9848 , n9849 , n9850 , n9851 , n9852 , n9853 , n9854 , n9855 , n9856 , n9857 , n9858 , n9859 , n9860 , n9861 , n9862 , n9863 , n9864 , n9865 , n9866 , n9867 , n9868 , n9869 , n9870 , n9871 , n9872 , n9873 , n9874 , n9875 , n9876 , n9877 , n9878 , n9879 , n9880 , n9881 , n9882 , n9883 , n9884 , n9885 , n9886 , n9887 , n9888 , n9889 , n9890 , n9891 , n9892 , n9893 , n9894 , n9895 , n9896 , n9897 , n9898 , n9899 , n9900 , n9901 , n9902 , n9903 , n9904 , n9905 , n9906 , n9907 , n9908 , n9909 , n9910 , n9911 , n9912 , n9913 , n9914 , n9915 , n9916 , n9917 , n9918 , n9919 , n9920 , n9921 , n9922 , n9923 , n9924 , n9925 , n9926 , n9927 , n9928 , n9929 , n9930 , n9931 , n9932 , n9933 , n9934 , n9935 , n9936 , n9937 , n9938 , n9939 , n9940 , n9941 , n9942 , n9943 , n9944 , n9945 , n9946 , n9947 , n9948 , n9949 , n9950 , n9951 , n9952 , n9953 , n9954 , n9955 , n9956 , n9957 , n9958 , n9959 , n9960 , n9961 , n9962 , n9963 , n9964 , n9965 , n9966 , n9967 , n9968 , n9969 , n9970 , n9971 , n9972 , n9973 , n9974 , n9975 , n9976 , n9977 , n9978 , n9979 , n9980 , n9981 , n9982 , n9983 , n9984 , n9985 , n9986 , n9987 , n9988 , n9989 , n9990 , n9991 , n9992 , n9993 , n9994 , n9995 , n9996 , n9997 , n9998 , n9999 , n10000 , n10001 , n10002 , n10003 , n10004 , n10005 , n10006 , n10007 , n10008 , n10009 , n10010 , n10011 , n10012 , n10013 , n10014 , n10015 , n10016 , n10017 , n10018 , n10019 , n10020 , n10021 , n10022 , n10023 , n10024 , n10025 , n10026 , n10027 , n10028 , n10029 , n10030 , n10031 , n10032 , n10033 , n10034 , n10035 , n10036 , n10037 , n10038 , n10039 , n10040 , n10041 , n10042 , n10043 , n10044 , n10045 , n10046 , n10047 , n10048 , n10049 , n10050 , n10051 , n10052 , n10053 , n10054 , n10055 , n10056 , n10057 , n10058 , n10059 , n10060 , n10061 , n10062 , n10063 , n10064 , n10065 , n10066 , n10067 , n10068 , n10069 , n10070 , n10071 , n10072 , n10073 , n10074 , n10075 , n10076 , n10077 , n10078 , n10079 , n10080 , n10081 , n10082 , n10083 , n10084 , n10085 , n10086 , n10087 , n10088 , n10089 , n10090 , n10091 , n10092 , n10093 , n10094 , n10095 , n10096 , n10097 , n10098 , n10099 , n10100 , n10101 , n10102 , n10103 , n10104 , n10105 , n10106 , n10107 , n10108 , n10109 , n10110 , n10111 , n10112 , n10113 , n10114 , n10115 , n10116 , n10117 , n10118 , n10119 , n10120 , n10121 , n10122 , n10123 , n10124 , n10125 , n10126 , n10127 , n10128 , n10129 , n10130 , n10131 , n10132 , n10133 , n10134 , n10135 , n10136 , n10137 , n10138 , n10139 , n10140 , n10141 , n10142 , n10143 , n10144 , n10145 , n10146 , n10147 , n10148 , n10149 , n10150 , n10151 , n10152 , n10153 , n10154 , n10155 , n10156 , n10157 , n10158 , n10159 , n10160 , n10161 , n10162 , n10163 , n10164 , n10165 , n10166 , n10167 , n10168 , n10169 , n10170 , n10171 , n10172 , n10173 , n10174 , n10175 , n10176 , n10177 , n10178 , n10179 , n10180 , n10181 , n10182 , n10183 , n10184 , n10185 , n10186 , n10187 , n10188 , n10189 , n10190 , n10191 , n10192 , n10193 , n10194 , n10195 , n10196 , n10197 , n10198 , n10199 , n10200 , n10201 , n10202 , n10203 , n10204 , n10205 , n10206 , n10207 , n10208 , n10209 , n10210 , n10211 , n10212 , n10213 , n10214 , n10215 , n10216 , n10217 , n10218 , n10219 , n10220 , n10221 , n10222 , n10223 , n10224 , n10225 , n10226 , n10227 , n10228 , n10229 , n10230 , n10231 , n10232 , n10233 , n10234 , n10235 , n10236 , n10237 , n10238 , n10239 , n10240 , n10241 , n10242 , n10243 , n10244 , n10245 , n10246 , n10247 , n10248 , n10249 , n10250 , n10251 ;
  assign n2146 = ~\dma_ack_i[8]_pad  & \dma_req_o[8]_pad  ;
  assign n2147 = \u11_status_reg[1]/P0001  & \u13_icc_r_reg[21]/NET0131  ;
  assign n2148 = ~\u11_status_reg[0]/P0001  & ~\u13_icc_r_reg[20]/NET0131  ;
  assign n2149 = ~n2147 & n2148 ;
  assign n2150 = ~\u11_status_reg[1]/P0001  & ~\u13_icc_r_reg[21]/NET0131  ;
  assign n2151 = ~\u11_full_reg/NET0131  & ~n2150 ;
  assign n2152 = ~n2149 & n2151 ;
  assign n2153 = \u13_icc_r_reg[16]/NET0131  & ~n2152 ;
  assign n2154 = ~\dma_ack_i[8]_pad  & \u13_icc_r_reg[22]/NET0131  ;
  assign n2155 = n2153 & n2154 ;
  assign n2156 = \u16_u8_dma_req_r1_reg/P0001  & n2155 ;
  assign n2157 = ~n2146 & ~n2156 ;
  assign n2158 = \u14_u5_en_out_l_reg/NET0131  & \valid_s_reg/NET0131  ;
  assign n2159 = ~\u14_u5_en_out_l2_reg/P0001  & n2158 ;
  assign n2160 = ~\u13_occ1_r_reg[10]/NET0131  & ~\u13_occ1_r_reg[11]/NET0131  ;
  assign n2161 = ~\u8_rp_reg[0]/P0001  & n2160 ;
  assign n2162 = n2159 & ~n2161 ;
  assign n2163 = \u8_rp_reg[1]/NET0131  & \u8_rp_reg[2]/NET0131  ;
  assign n2164 = n2162 & n2163 ;
  assign n2166 = \u8_rp_reg[3]/NET0131  & n2164 ;
  assign n2165 = ~\u8_rp_reg[3]/NET0131  & ~n2164 ;
  assign n2167 = \u13_occ1_r_reg[8]/NET0131  & ~n2165 ;
  assign n2168 = ~n2166 & n2167 ;
  assign n2169 = ~\u0_slt0_r_reg[14]/P0001  & ~\u2_ld_reg/P0001  ;
  assign n2173 = ~\u14_u3_en_out_l_reg/NET0131  & ~\u14_u4_en_out_l_reg/NET0131  ;
  assign n2174 = ~\u14_u5_en_out_l_reg/NET0131  & n2173 ;
  assign n2170 = ~\u14_crac_wr_r_reg/P0001  & \u2_ld_reg/P0001  ;
  assign n2171 = ~\u14_crac_valid_r_reg/P0001  & ~\u14_u0_en_out_l_reg/NET0131  ;
  assign n2172 = ~\u14_u1_en_out_l_reg/NET0131  & ~\u14_u2_en_out_l_reg/NET0131  ;
  assign n2175 = n2171 & n2172 ;
  assign n2176 = n2170 & n2175 ;
  assign n2177 = n2174 & n2176 ;
  assign n2178 = ~n2169 & ~n2177 ;
  assign n2179 = \u14_crac_valid_r_reg/P0001  & \u2_ld_reg/P0001  ;
  assign n2180 = \u0_slt0_r_reg[13]/P0001  & ~\u2_ld_reg/P0001  ;
  assign n2181 = ~n2179 & ~n2180 ;
  assign n2182 = ~\u0_slt0_r_reg[12]/P0001  & ~\u2_ld_reg/P0001  ;
  assign n2183 = ~n2170 & ~n2182 ;
  assign n2184 = \u0_slt0_r_reg[11]/P0001  & ~\u2_ld_reg/P0001  ;
  assign n2185 = \u14_u0_en_out_l_reg/NET0131  & \u2_ld_reg/P0001  ;
  assign n2186 = ~n2184 & ~n2185 ;
  assign n2187 = \u14_u1_en_out_l_reg/NET0131  & \u2_ld_reg/P0001  ;
  assign n2188 = \u0_slt0_r_reg[10]/P0001  & ~\u2_ld_reg/P0001  ;
  assign n2189 = ~n2187 & ~n2188 ;
  assign n2190 = \u0_slt0_r_reg[9]/P0001  & ~\u2_ld_reg/P0001  ;
  assign n2191 = \u14_u2_en_out_l_reg/NET0131  & \u2_ld_reg/P0001  ;
  assign n2192 = \u0_slt0_r_reg[8]/P0001  & ~\u2_ld_reg/P0001  ;
  assign n2193 = ~n2191 & ~n2192 ;
  assign n2194 = \u14_u3_en_out_l_reg/NET0131  & \u2_ld_reg/P0001  ;
  assign n2195 = \u0_slt0_r_reg[7]/P0001  & ~\u2_ld_reg/P0001  ;
  assign n2196 = ~n2194 & ~n2195 ;
  assign n2197 = \u14_u4_en_out_l_reg/NET0131  & \u2_ld_reg/P0001  ;
  assign n2198 = \u0_slt0_r_reg[6]/P0001  & ~\u2_ld_reg/P0001  ;
  assign n2199 = ~n2197 & ~n2198 ;
  assign n2200 = \u0_slt0_r_reg[5]/P0001  & ~\u2_ld_reg/P0001  ;
  assign n2201 = \u14_u5_en_out_l_reg/NET0131  & \u2_ld_reg/P0001  ;
  assign n2202 = ~n2200 & ~n2201 ;
  assign n2203 = \u0_slt0_r_reg[4]/P0001  & ~\u2_ld_reg/P0001  ;
  assign n2204 = \u0_slt0_r_reg[3]/P0001  & ~\u2_ld_reg/P0001  ;
  assign n2205 = \u0_slt0_r_reg[2]/P0001  & ~\u2_ld_reg/P0001  ;
  assign n2206 = \u0_slt0_r_reg[1]/P0001  & ~\u2_ld_reg/P0001  ;
  assign n2207 = \u0_slt0_r_reg[0]/P0001  & ~\u2_ld_reg/P0001  ;
  assign n2208 = \u0_slt1_r_reg[19]/P0001  & ~\u2_ld_reg/P0001  ;
  assign n2209 = \u13_crac_r_reg[7]/NET0131  & \u2_ld_reg/P0001  ;
  assign n2210 = \u0_slt1_r_reg[18]/P0001  & ~\u2_ld_reg/P0001  ;
  assign n2211 = ~n2209 & ~n2210 ;
  assign n2212 = \u13_crac_r_reg[6]/NET0131  & \u2_ld_reg/P0001  ;
  assign n2213 = \u0_slt1_r_reg[17]/P0001  & ~\u2_ld_reg/P0001  ;
  assign n2214 = ~n2212 & ~n2213 ;
  assign n2215 = \u13_crac_r_reg[5]/NET0131  & \u2_ld_reg/P0001  ;
  assign n2216 = \u0_slt1_r_reg[16]/P0001  & ~\u2_ld_reg/P0001  ;
  assign n2217 = ~n2215 & ~n2216 ;
  assign n2218 = \u13_crac_r_reg[4]/NET0131  & \u2_ld_reg/P0001  ;
  assign n2219 = \u0_slt1_r_reg[15]/P0001  & ~\u2_ld_reg/P0001  ;
  assign n2220 = ~n2218 & ~n2219 ;
  assign n2221 = \u13_crac_r_reg[3]/NET0131  & \u2_ld_reg/P0001  ;
  assign n2222 = \u0_slt1_r_reg[14]/P0001  & ~\u2_ld_reg/P0001  ;
  assign n2223 = ~n2221 & ~n2222 ;
  assign n2224 = \u13_crac_r_reg[2]/NET0131  & \u2_ld_reg/P0001  ;
  assign n2225 = \u0_slt1_r_reg[13]/P0001  & ~\u2_ld_reg/P0001  ;
  assign n2226 = ~n2224 & ~n2225 ;
  assign n2227 = \u13_crac_r_reg[1]/NET0131  & \u2_ld_reg/P0001  ;
  assign n2228 = \u0_slt1_r_reg[12]/P0001  & ~\u2_ld_reg/P0001  ;
  assign n2229 = ~n2227 & ~n2228 ;
  assign n2230 = \u13_crac_r_reg[0]/NET0131  & \u2_ld_reg/P0001  ;
  assign n2231 = \u0_slt1_r_reg[11]/P0001  & ~\u2_ld_reg/P0001  ;
  assign n2232 = ~n2230 & ~n2231 ;
  assign n2233 = \u0_slt1_r_reg[10]/P0001  & ~\u2_ld_reg/P0001  ;
  assign n2234 = \u0_slt1_r_reg[9]/P0001  & ~\u2_ld_reg/P0001  ;
  assign n2235 = \u0_slt1_r_reg[8]/P0001  & ~\u2_ld_reg/P0001  ;
  assign n2236 = \u0_slt1_r_reg[7]/P0001  & ~\u2_ld_reg/P0001  ;
  assign n2237 = \u0_slt1_r_reg[6]/P0001  & ~\u2_ld_reg/P0001  ;
  assign n2238 = \u0_slt1_r_reg[5]/P0001  & ~\u2_ld_reg/P0001  ;
  assign n2239 = \u0_slt1_r_reg[4]/P0001  & ~\u2_ld_reg/P0001  ;
  assign n2240 = \u0_slt1_r_reg[3]/P0001  & ~\u2_ld_reg/P0001  ;
  assign n2241 = \u0_slt1_r_reg[2]/P0001  & ~\u2_ld_reg/P0001  ;
  assign n2242 = \u0_slt1_r_reg[1]/P0001  & ~\u2_ld_reg/P0001  ;
  assign n2243 = \u0_slt1_r_reg[0]/P0001  & ~\u2_ld_reg/P0001  ;
  assign n2244 = \u0_slt2_r_reg[19]/P0001  & ~\u2_ld_reg/P0001  ;
  assign n2245 = \u13_crac_dout_r_reg[15]/P0001  & \u2_ld_reg/P0001  ;
  assign n2246 = \u0_slt2_r_reg[18]/P0001  & ~\u2_ld_reg/P0001  ;
  assign n2247 = ~n2245 & ~n2246 ;
  assign n2248 = \u13_crac_dout_r_reg[14]/P0001  & \u2_ld_reg/P0001  ;
  assign n2249 = \u0_slt2_r_reg[17]/P0001  & ~\u2_ld_reg/P0001  ;
  assign n2250 = ~n2248 & ~n2249 ;
  assign n2251 = \u13_crac_dout_r_reg[13]/P0001  & \u2_ld_reg/P0001  ;
  assign n2252 = \u0_slt2_r_reg[16]/P0001  & ~\u2_ld_reg/P0001  ;
  assign n2253 = ~n2251 & ~n2252 ;
  assign n2254 = \u13_crac_dout_r_reg[12]/P0001  & \u2_ld_reg/P0001  ;
  assign n2255 = \u0_slt2_r_reg[15]/P0001  & ~\u2_ld_reg/P0001  ;
  assign n2256 = ~n2254 & ~n2255 ;
  assign n2257 = \u13_crac_dout_r_reg[11]/P0001  & \u2_ld_reg/P0001  ;
  assign n2258 = \u0_slt2_r_reg[14]/P0001  & ~\u2_ld_reg/P0001  ;
  assign n2259 = ~n2257 & ~n2258 ;
  assign n2260 = \u13_crac_dout_r_reg[10]/P0001  & \u2_ld_reg/P0001  ;
  assign n2261 = \u0_slt2_r_reg[13]/P0001  & ~\u2_ld_reg/P0001  ;
  assign n2262 = ~n2260 & ~n2261 ;
  assign n2263 = \u13_crac_dout_r_reg[9]/P0001  & \u2_ld_reg/P0001  ;
  assign n2264 = \u0_slt2_r_reg[12]/P0001  & ~\u2_ld_reg/P0001  ;
  assign n2265 = ~n2263 & ~n2264 ;
  assign n2266 = \u13_crac_dout_r_reg[8]/P0001  & \u2_ld_reg/P0001  ;
  assign n2267 = \u0_slt2_r_reg[11]/P0001  & ~\u2_ld_reg/P0001  ;
  assign n2268 = ~n2266 & ~n2267 ;
  assign n2269 = \u13_crac_dout_r_reg[7]/P0001  & \u2_ld_reg/P0001  ;
  assign n2270 = \u0_slt2_r_reg[10]/P0001  & ~\u2_ld_reg/P0001  ;
  assign n2271 = ~n2269 & ~n2270 ;
  assign n2272 = \u13_crac_dout_r_reg[6]/P0001  & \u2_ld_reg/P0001  ;
  assign n2273 = \u0_slt2_r_reg[9]/P0001  & ~\u2_ld_reg/P0001  ;
  assign n2274 = ~n2272 & ~n2273 ;
  assign n2275 = \u13_crac_dout_r_reg[5]/P0001  & \u2_ld_reg/P0001  ;
  assign n2276 = \u0_slt2_r_reg[8]/P0001  & ~\u2_ld_reg/P0001  ;
  assign n2277 = ~n2275 & ~n2276 ;
  assign n2278 = \u13_crac_dout_r_reg[4]/P0001  & \u2_ld_reg/P0001  ;
  assign n2279 = \u0_slt2_r_reg[7]/P0001  & ~\u2_ld_reg/P0001  ;
  assign n2280 = ~n2278 & ~n2279 ;
  assign n2281 = \u13_crac_dout_r_reg[3]/P0001  & \u2_ld_reg/P0001  ;
  assign n2282 = \u0_slt2_r_reg[6]/P0001  & ~\u2_ld_reg/P0001  ;
  assign n2283 = ~n2281 & ~n2282 ;
  assign n2284 = \u13_crac_dout_r_reg[2]/P0001  & \u2_ld_reg/P0001  ;
  assign n2285 = \u0_slt2_r_reg[5]/P0001  & ~\u2_ld_reg/P0001  ;
  assign n2286 = ~n2284 & ~n2285 ;
  assign n2287 = \u13_crac_dout_r_reg[1]/P0001  & \u2_ld_reg/P0001  ;
  assign n2288 = \u0_slt2_r_reg[4]/P0001  & ~\u2_ld_reg/P0001  ;
  assign n2289 = ~n2287 & ~n2288 ;
  assign n2290 = \u13_crac_dout_r_reg[0]/P0001  & \u2_ld_reg/P0001  ;
  assign n2291 = \u0_slt2_r_reg[3]/P0001  & ~\u2_ld_reg/P0001  ;
  assign n2292 = ~n2290 & ~n2291 ;
  assign n2293 = \u0_slt2_r_reg[2]/P0001  & ~\u2_ld_reg/P0001  ;
  assign n2294 = \u0_slt2_r_reg[1]/P0001  & ~\u2_ld_reg/P0001  ;
  assign n2295 = \u0_slt2_r_reg[0]/P0001  & ~\u2_ld_reg/P0001  ;
  assign n2296 = \u0_slt3_r_reg[19]/P0001  & ~\u2_ld_reg/P0001  ;
  assign n2297 = \u2_ld_reg/P0001  & \u3_dout_reg[19]/P0001  ;
  assign n2298 = \u0_slt3_r_reg[18]/P0001  & ~\u2_ld_reg/P0001  ;
  assign n2299 = ~n2297 & ~n2298 ;
  assign n2300 = \u2_ld_reg/P0001  & \u3_dout_reg[18]/P0001  ;
  assign n2301 = \u0_slt3_r_reg[17]/P0001  & ~\u2_ld_reg/P0001  ;
  assign n2302 = ~n2300 & ~n2301 ;
  assign n2303 = \u2_ld_reg/P0001  & \u3_dout_reg[17]/P0001  ;
  assign n2304 = \u0_slt3_r_reg[16]/P0001  & ~\u2_ld_reg/P0001  ;
  assign n2305 = ~n2303 & ~n2304 ;
  assign n2306 = \u2_ld_reg/P0001  & \u3_dout_reg[16]/P0001  ;
  assign n2307 = \u0_slt3_r_reg[15]/P0001  & ~\u2_ld_reg/P0001  ;
  assign n2308 = ~n2306 & ~n2307 ;
  assign n2309 = \u2_ld_reg/P0001  & \u3_dout_reg[15]/P0001  ;
  assign n2310 = \u0_slt3_r_reg[14]/P0001  & ~\u2_ld_reg/P0001  ;
  assign n2311 = ~n2309 & ~n2310 ;
  assign n2312 = \u2_ld_reg/P0001  & \u3_dout_reg[14]/P0001  ;
  assign n2313 = \u0_slt3_r_reg[13]/P0001  & ~\u2_ld_reg/P0001  ;
  assign n2314 = ~n2312 & ~n2313 ;
  assign n2315 = \u2_ld_reg/P0001  & \u3_dout_reg[13]/P0001  ;
  assign n2316 = \u0_slt3_r_reg[12]/P0001  & ~\u2_ld_reg/P0001  ;
  assign n2317 = ~n2315 & ~n2316 ;
  assign n2318 = \u2_ld_reg/P0001  & \u3_dout_reg[12]/P0001  ;
  assign n2319 = \u0_slt3_r_reg[11]/P0001  & ~\u2_ld_reg/P0001  ;
  assign n2320 = ~n2318 & ~n2319 ;
  assign n2321 = \u2_ld_reg/P0001  & \u3_dout_reg[11]/P0001  ;
  assign n2322 = \u0_slt3_r_reg[10]/P0001  & ~\u2_ld_reg/P0001  ;
  assign n2323 = ~n2321 & ~n2322 ;
  assign n2324 = \u2_ld_reg/P0001  & \u3_dout_reg[10]/P0001  ;
  assign n2325 = \u0_slt3_r_reg[9]/P0001  & ~\u2_ld_reg/P0001  ;
  assign n2326 = ~n2324 & ~n2325 ;
  assign n2327 = \u2_ld_reg/P0001  & \u3_dout_reg[9]/P0001  ;
  assign n2328 = \u0_slt3_r_reg[8]/P0001  & ~\u2_ld_reg/P0001  ;
  assign n2329 = ~n2327 & ~n2328 ;
  assign n2330 = \u2_ld_reg/P0001  & \u3_dout_reg[8]/P0001  ;
  assign n2331 = \u0_slt3_r_reg[7]/P0001  & ~\u2_ld_reg/P0001  ;
  assign n2332 = ~n2330 & ~n2331 ;
  assign n2333 = \u2_ld_reg/P0001  & \u3_dout_reg[7]/P0001  ;
  assign n2334 = \u0_slt3_r_reg[6]/P0001  & ~\u2_ld_reg/P0001  ;
  assign n2335 = ~n2333 & ~n2334 ;
  assign n2336 = \u2_ld_reg/P0001  & \u3_dout_reg[6]/P0001  ;
  assign n2337 = \u0_slt3_r_reg[5]/P0001  & ~\u2_ld_reg/P0001  ;
  assign n2338 = ~n2336 & ~n2337 ;
  assign n2339 = \u2_ld_reg/P0001  & \u3_dout_reg[5]/P0001  ;
  assign n2340 = \u0_slt3_r_reg[4]/P0001  & ~\u2_ld_reg/P0001  ;
  assign n2341 = ~n2339 & ~n2340 ;
  assign n2342 = \u2_ld_reg/P0001  & \u3_dout_reg[4]/P0001  ;
  assign n2343 = \u0_slt3_r_reg[3]/P0001  & ~\u2_ld_reg/P0001  ;
  assign n2344 = ~n2342 & ~n2343 ;
  assign n2345 = \u2_ld_reg/P0001  & \u3_dout_reg[3]/P0001  ;
  assign n2346 = \u0_slt3_r_reg[2]/P0001  & ~\u2_ld_reg/P0001  ;
  assign n2347 = ~n2345 & ~n2346 ;
  assign n2348 = \u2_ld_reg/P0001  & \u3_dout_reg[2]/P0001  ;
  assign n2349 = \u0_slt3_r_reg[1]/P0001  & ~\u2_ld_reg/P0001  ;
  assign n2350 = ~n2348 & ~n2349 ;
  assign n2351 = \u2_ld_reg/P0001  & \u3_dout_reg[1]/P0001  ;
  assign n2352 = \u0_slt3_r_reg[0]/P0001  & ~\u2_ld_reg/P0001  ;
  assign n2353 = ~n2351 & ~n2352 ;
  assign n2354 = \u2_ld_reg/P0001  & \u3_dout_reg[0]/P0001  ;
  assign n2355 = \u0_slt4_r_reg[19]/P0001  & ~\u2_ld_reg/P0001  ;
  assign n2356 = ~n2354 & ~n2355 ;
  assign n2357 = \u2_ld_reg/P0001  & \u4_dout_reg[19]/P0001  ;
  assign n2358 = \u0_slt4_r_reg[18]/P0001  & ~\u2_ld_reg/P0001  ;
  assign n2359 = ~n2357 & ~n2358 ;
  assign n2360 = \u2_ld_reg/P0001  & \u4_dout_reg[18]/P0001  ;
  assign n2361 = \u0_slt4_r_reg[17]/P0001  & ~\u2_ld_reg/P0001  ;
  assign n2362 = ~n2360 & ~n2361 ;
  assign n2363 = \u2_ld_reg/P0001  & \u4_dout_reg[17]/P0001  ;
  assign n2364 = \u0_slt4_r_reg[16]/P0001  & ~\u2_ld_reg/P0001  ;
  assign n2365 = ~n2363 & ~n2364 ;
  assign n2366 = \u2_ld_reg/P0001  & \u4_dout_reg[16]/P0001  ;
  assign n2367 = \u0_slt4_r_reg[15]/P0001  & ~\u2_ld_reg/P0001  ;
  assign n2368 = ~n2366 & ~n2367 ;
  assign n2369 = \u2_ld_reg/P0001  & \u4_dout_reg[15]/P0001  ;
  assign n2370 = \u0_slt4_r_reg[14]/P0001  & ~\u2_ld_reg/P0001  ;
  assign n2371 = ~n2369 & ~n2370 ;
  assign n2372 = \u2_ld_reg/P0001  & \u4_dout_reg[14]/P0001  ;
  assign n2373 = \u0_slt4_r_reg[13]/P0001  & ~\u2_ld_reg/P0001  ;
  assign n2374 = ~n2372 & ~n2373 ;
  assign n2375 = \u2_ld_reg/P0001  & \u4_dout_reg[13]/P0001  ;
  assign n2376 = \u0_slt4_r_reg[12]/P0001  & ~\u2_ld_reg/P0001  ;
  assign n2377 = ~n2375 & ~n2376 ;
  assign n2378 = \u2_ld_reg/P0001  & \u4_dout_reg[12]/P0001  ;
  assign n2379 = \u0_slt4_r_reg[11]/P0001  & ~\u2_ld_reg/P0001  ;
  assign n2380 = ~n2378 & ~n2379 ;
  assign n2381 = \u2_ld_reg/P0001  & \u4_dout_reg[11]/P0001  ;
  assign n2382 = \u0_slt4_r_reg[10]/P0001  & ~\u2_ld_reg/P0001  ;
  assign n2383 = ~n2381 & ~n2382 ;
  assign n2384 = \u2_ld_reg/P0001  & \u4_dout_reg[10]/P0001  ;
  assign n2385 = \u0_slt4_r_reg[9]/P0001  & ~\u2_ld_reg/P0001  ;
  assign n2386 = ~n2384 & ~n2385 ;
  assign n2387 = \u2_ld_reg/P0001  & \u4_dout_reg[9]/P0001  ;
  assign n2388 = \u0_slt4_r_reg[8]/P0001  & ~\u2_ld_reg/P0001  ;
  assign n2389 = ~n2387 & ~n2388 ;
  assign n2390 = \u2_ld_reg/P0001  & \u4_dout_reg[8]/P0001  ;
  assign n2391 = \u0_slt4_r_reg[7]/P0001  & ~\u2_ld_reg/P0001  ;
  assign n2392 = ~n2390 & ~n2391 ;
  assign n2393 = \u2_ld_reg/P0001  & \u4_dout_reg[7]/P0001  ;
  assign n2394 = \u0_slt4_r_reg[6]/P0001  & ~\u2_ld_reg/P0001  ;
  assign n2395 = ~n2393 & ~n2394 ;
  assign n2396 = \u2_ld_reg/P0001  & \u4_dout_reg[6]/P0001  ;
  assign n2397 = \u0_slt4_r_reg[5]/P0001  & ~\u2_ld_reg/P0001  ;
  assign n2398 = ~n2396 & ~n2397 ;
  assign n2399 = \u2_ld_reg/P0001  & \u4_dout_reg[5]/P0001  ;
  assign n2400 = \u0_slt4_r_reg[4]/P0001  & ~\u2_ld_reg/P0001  ;
  assign n2401 = ~n2399 & ~n2400 ;
  assign n2402 = \u2_ld_reg/P0001  & \u4_dout_reg[4]/P0001  ;
  assign n2403 = \u0_slt4_r_reg[3]/P0001  & ~\u2_ld_reg/P0001  ;
  assign n2404 = ~n2402 & ~n2403 ;
  assign n2405 = \u2_ld_reg/P0001  & \u4_dout_reg[3]/P0001  ;
  assign n2406 = \u0_slt4_r_reg[2]/P0001  & ~\u2_ld_reg/P0001  ;
  assign n2407 = ~n2405 & ~n2406 ;
  assign n2408 = \u2_ld_reg/P0001  & \u4_dout_reg[2]/P0001  ;
  assign n2409 = \u0_slt4_r_reg[1]/P0001  & ~\u2_ld_reg/P0001  ;
  assign n2410 = ~n2408 & ~n2409 ;
  assign n2411 = \u2_ld_reg/P0001  & \u4_dout_reg[1]/P0001  ;
  assign n2412 = \u0_slt4_r_reg[0]/P0001  & ~\u2_ld_reg/P0001  ;
  assign n2413 = ~n2411 & ~n2412 ;
  assign n2414 = \u2_ld_reg/P0001  & \u4_dout_reg[0]/P0001  ;
  assign n2415 = \u0_slt5_r_reg[19]/P0001  & ~\u2_ld_reg/P0001  ;
  assign n2416 = ~n2414 & ~n2415 ;
  assign n2417 = \u0_slt5_r_reg[18]/P0001  & ~\u2_ld_reg/P0001  ;
  assign n2418 = \u0_slt5_r_reg[17]/P0001  & ~\u2_ld_reg/P0001  ;
  assign n2419 = \u0_slt5_r_reg[16]/P0001  & ~\u2_ld_reg/P0001  ;
  assign n2420 = \u0_slt5_r_reg[15]/P0001  & ~\u2_ld_reg/P0001  ;
  assign n2421 = \u0_slt5_r_reg[14]/P0001  & ~\u2_ld_reg/P0001  ;
  assign n2422 = \u0_slt5_r_reg[13]/P0001  & ~\u2_ld_reg/P0001  ;
  assign n2423 = \u0_slt5_r_reg[12]/P0001  & ~\u2_ld_reg/P0001  ;
  assign n2424 = \u0_slt5_r_reg[11]/P0001  & ~\u2_ld_reg/P0001  ;
  assign n2425 = \u0_slt5_r_reg[10]/P0001  & ~\u2_ld_reg/P0001  ;
  assign n2426 = \u0_slt5_r_reg[9]/P0001  & ~\u2_ld_reg/P0001  ;
  assign n2427 = \u0_slt5_r_reg[8]/P0001  & ~\u2_ld_reg/P0001  ;
  assign n2428 = \u0_slt5_r_reg[7]/P0001  & ~\u2_ld_reg/P0001  ;
  assign n2429 = \u0_slt5_r_reg[6]/P0001  & ~\u2_ld_reg/P0001  ;
  assign n2430 = \u0_slt5_r_reg[5]/P0001  & ~\u2_ld_reg/P0001  ;
  assign n2431 = \u0_slt5_r_reg[4]/P0001  & ~\u2_ld_reg/P0001  ;
  assign n2432 = \u0_slt5_r_reg[3]/P0001  & ~\u2_ld_reg/P0001  ;
  assign n2433 = \u0_slt5_r_reg[2]/P0001  & ~\u2_ld_reg/P0001  ;
  assign n2434 = \u0_slt5_r_reg[1]/P0001  & ~\u2_ld_reg/P0001  ;
  assign n2435 = \u0_slt5_r_reg[0]/P0001  & ~\u2_ld_reg/P0001  ;
  assign n2436 = \u0_slt6_r_reg[19]/P0001  & ~\u2_ld_reg/P0001  ;
  assign n2437 = \u2_ld_reg/P0001  & \u5_dout_reg[19]/P0001  ;
  assign n2438 = \u0_slt6_r_reg[18]/P0001  & ~\u2_ld_reg/P0001  ;
  assign n2439 = ~n2437 & ~n2438 ;
  assign n2440 = \u2_ld_reg/P0001  & \u5_dout_reg[18]/P0001  ;
  assign n2441 = \u0_slt6_r_reg[17]/P0001  & ~\u2_ld_reg/P0001  ;
  assign n2442 = ~n2440 & ~n2441 ;
  assign n2443 = \u2_ld_reg/P0001  & \u5_dout_reg[17]/P0001  ;
  assign n2444 = \u0_slt6_r_reg[16]/P0001  & ~\u2_ld_reg/P0001  ;
  assign n2445 = ~n2443 & ~n2444 ;
  assign n2446 = \u2_ld_reg/P0001  & \u5_dout_reg[16]/P0001  ;
  assign n2447 = \u0_slt6_r_reg[15]/P0001  & ~\u2_ld_reg/P0001  ;
  assign n2448 = ~n2446 & ~n2447 ;
  assign n2449 = \u2_ld_reg/P0001  & \u5_dout_reg[15]/P0001  ;
  assign n2450 = \u0_slt6_r_reg[14]/P0001  & ~\u2_ld_reg/P0001  ;
  assign n2451 = ~n2449 & ~n2450 ;
  assign n2452 = \u2_ld_reg/P0001  & \u5_dout_reg[14]/P0001  ;
  assign n2453 = \u0_slt6_r_reg[13]/P0001  & ~\u2_ld_reg/P0001  ;
  assign n2454 = ~n2452 & ~n2453 ;
  assign n2455 = \u2_ld_reg/P0001  & \u5_dout_reg[13]/P0001  ;
  assign n2456 = \u0_slt6_r_reg[12]/P0001  & ~\u2_ld_reg/P0001  ;
  assign n2457 = ~n2455 & ~n2456 ;
  assign n2458 = \u2_ld_reg/P0001  & \u5_dout_reg[12]/P0001  ;
  assign n2459 = \u0_slt6_r_reg[11]/P0001  & ~\u2_ld_reg/P0001  ;
  assign n2460 = ~n2458 & ~n2459 ;
  assign n2461 = \u2_ld_reg/P0001  & \u5_dout_reg[11]/P0001  ;
  assign n2462 = \u0_slt6_r_reg[10]/P0001  & ~\u2_ld_reg/P0001  ;
  assign n2463 = ~n2461 & ~n2462 ;
  assign n2464 = \u2_ld_reg/P0001  & \u5_dout_reg[10]/P0001  ;
  assign n2465 = \u0_slt6_r_reg[9]/P0001  & ~\u2_ld_reg/P0001  ;
  assign n2466 = ~n2464 & ~n2465 ;
  assign n2467 = \u2_ld_reg/P0001  & \u5_dout_reg[9]/P0001  ;
  assign n2468 = \u0_slt6_r_reg[8]/P0001  & ~\u2_ld_reg/P0001  ;
  assign n2469 = ~n2467 & ~n2468 ;
  assign n2470 = \u2_ld_reg/P0001  & \u5_dout_reg[8]/P0001  ;
  assign n2471 = \u0_slt6_r_reg[7]/P0001  & ~\u2_ld_reg/P0001  ;
  assign n2472 = ~n2470 & ~n2471 ;
  assign n2473 = \u2_ld_reg/P0001  & \u5_dout_reg[7]/P0001  ;
  assign n2474 = \u0_slt6_r_reg[6]/P0001  & ~\u2_ld_reg/P0001  ;
  assign n2475 = ~n2473 & ~n2474 ;
  assign n2476 = \u2_ld_reg/P0001  & \u5_dout_reg[6]/P0001  ;
  assign n2477 = \u0_slt6_r_reg[5]/P0001  & ~\u2_ld_reg/P0001  ;
  assign n2478 = ~n2476 & ~n2477 ;
  assign n2479 = \u2_ld_reg/P0001  & \u5_dout_reg[5]/P0001  ;
  assign n2480 = \u0_slt6_r_reg[4]/P0001  & ~\u2_ld_reg/P0001  ;
  assign n2481 = ~n2479 & ~n2480 ;
  assign n2482 = \u2_ld_reg/P0001  & \u5_dout_reg[4]/P0001  ;
  assign n2483 = \u0_slt6_r_reg[3]/P0001  & ~\u2_ld_reg/P0001  ;
  assign n2484 = ~n2482 & ~n2483 ;
  assign n2485 = \u2_ld_reg/P0001  & \u5_dout_reg[3]/P0001  ;
  assign n2486 = \u0_slt6_r_reg[2]/P0001  & ~\u2_ld_reg/P0001  ;
  assign n2487 = ~n2485 & ~n2486 ;
  assign n2488 = \u2_ld_reg/P0001  & \u5_dout_reg[2]/P0001  ;
  assign n2489 = \u0_slt6_r_reg[1]/P0001  & ~\u2_ld_reg/P0001  ;
  assign n2490 = ~n2488 & ~n2489 ;
  assign n2491 = \u2_ld_reg/P0001  & \u5_dout_reg[1]/P0001  ;
  assign n2492 = \u0_slt6_r_reg[0]/P0001  & ~\u2_ld_reg/P0001  ;
  assign n2493 = ~n2491 & ~n2492 ;
  assign n2494 = \u2_ld_reg/P0001  & \u5_dout_reg[0]/P0001  ;
  assign n2495 = \u0_slt7_r_reg[19]/P0001  & ~\u2_ld_reg/P0001  ;
  assign n2496 = ~n2494 & ~n2495 ;
  assign n2497 = \u2_ld_reg/P0001  & \u6_dout_reg[19]/P0001  ;
  assign n2498 = \u0_slt7_r_reg[18]/P0001  & ~\u2_ld_reg/P0001  ;
  assign n2499 = ~n2497 & ~n2498 ;
  assign n2500 = \u2_ld_reg/P0001  & \u6_dout_reg[18]/P0001  ;
  assign n2501 = \u0_slt7_r_reg[17]/P0001  & ~\u2_ld_reg/P0001  ;
  assign n2502 = ~n2500 & ~n2501 ;
  assign n2503 = \u2_ld_reg/P0001  & \u6_dout_reg[17]/P0001  ;
  assign n2504 = \u0_slt7_r_reg[16]/P0001  & ~\u2_ld_reg/P0001  ;
  assign n2505 = ~n2503 & ~n2504 ;
  assign n2506 = \u2_ld_reg/P0001  & \u6_dout_reg[16]/P0001  ;
  assign n2507 = \u0_slt7_r_reg[15]/P0001  & ~\u2_ld_reg/P0001  ;
  assign n2508 = ~n2506 & ~n2507 ;
  assign n2509 = \u2_ld_reg/P0001  & \u6_dout_reg[15]/P0001  ;
  assign n2510 = \u0_slt7_r_reg[14]/P0001  & ~\u2_ld_reg/P0001  ;
  assign n2511 = ~n2509 & ~n2510 ;
  assign n2512 = \u2_ld_reg/P0001  & \u6_dout_reg[14]/P0001  ;
  assign n2513 = \u0_slt7_r_reg[13]/P0001  & ~\u2_ld_reg/P0001  ;
  assign n2514 = ~n2512 & ~n2513 ;
  assign n2515 = \u2_ld_reg/P0001  & \u6_dout_reg[13]/P0001  ;
  assign n2516 = \u0_slt7_r_reg[12]/P0001  & ~\u2_ld_reg/P0001  ;
  assign n2517 = ~n2515 & ~n2516 ;
  assign n2518 = \u2_ld_reg/P0001  & \u6_dout_reg[12]/P0001  ;
  assign n2519 = \u0_slt7_r_reg[11]/P0001  & ~\u2_ld_reg/P0001  ;
  assign n2520 = ~n2518 & ~n2519 ;
  assign n2521 = \u2_ld_reg/P0001  & \u6_dout_reg[11]/P0001  ;
  assign n2522 = \u0_slt7_r_reg[10]/P0001  & ~\u2_ld_reg/P0001  ;
  assign n2523 = ~n2521 & ~n2522 ;
  assign n2524 = \u2_ld_reg/P0001  & \u6_dout_reg[10]/P0001  ;
  assign n2525 = \u0_slt7_r_reg[9]/P0001  & ~\u2_ld_reg/P0001  ;
  assign n2526 = ~n2524 & ~n2525 ;
  assign n2527 = \u2_ld_reg/P0001  & \u6_dout_reg[9]/P0001  ;
  assign n2528 = \u0_slt7_r_reg[8]/P0001  & ~\u2_ld_reg/P0001  ;
  assign n2529 = ~n2527 & ~n2528 ;
  assign n2530 = \u2_ld_reg/P0001  & \u6_dout_reg[8]/P0001  ;
  assign n2531 = \u0_slt7_r_reg[7]/P0001  & ~\u2_ld_reg/P0001  ;
  assign n2532 = ~n2530 & ~n2531 ;
  assign n2533 = \u2_ld_reg/P0001  & \u6_dout_reg[7]/P0001  ;
  assign n2534 = \u0_slt7_r_reg[6]/P0001  & ~\u2_ld_reg/P0001  ;
  assign n2535 = ~n2533 & ~n2534 ;
  assign n2536 = \u2_ld_reg/P0001  & \u6_dout_reg[6]/P0001  ;
  assign n2537 = \u0_slt7_r_reg[5]/P0001  & ~\u2_ld_reg/P0001  ;
  assign n2538 = ~n2536 & ~n2537 ;
  assign n2539 = \u2_ld_reg/P0001  & \u6_dout_reg[5]/P0001  ;
  assign n2540 = \u0_slt7_r_reg[4]/P0001  & ~\u2_ld_reg/P0001  ;
  assign n2541 = ~n2539 & ~n2540 ;
  assign n2542 = \u2_ld_reg/P0001  & \u6_dout_reg[4]/P0001  ;
  assign n2543 = \u0_slt7_r_reg[3]/P0001  & ~\u2_ld_reg/P0001  ;
  assign n2544 = ~n2542 & ~n2543 ;
  assign n2545 = \u2_ld_reg/P0001  & \u6_dout_reg[3]/P0001  ;
  assign n2546 = \u0_slt7_r_reg[2]/P0001  & ~\u2_ld_reg/P0001  ;
  assign n2547 = ~n2545 & ~n2546 ;
  assign n2548 = \u2_ld_reg/P0001  & \u6_dout_reg[2]/P0001  ;
  assign n2549 = \u0_slt7_r_reg[1]/P0001  & ~\u2_ld_reg/P0001  ;
  assign n2550 = ~n2548 & ~n2549 ;
  assign n2551 = \u2_ld_reg/P0001  & \u6_dout_reg[1]/P0001  ;
  assign n2552 = \u0_slt7_r_reg[0]/P0001  & ~\u2_ld_reg/P0001  ;
  assign n2553 = ~n2551 & ~n2552 ;
  assign n2554 = \u2_ld_reg/P0001  & \u6_dout_reg[0]/P0001  ;
  assign n2555 = \u0_slt8_r_reg[19]/P0001  & ~\u2_ld_reg/P0001  ;
  assign n2556 = ~n2554 & ~n2555 ;
  assign n2557 = \u2_ld_reg/P0001  & \u7_dout_reg[19]/P0001  ;
  assign n2558 = \u0_slt8_r_reg[18]/P0001  & ~\u2_ld_reg/P0001  ;
  assign n2559 = ~n2557 & ~n2558 ;
  assign n2560 = \u2_ld_reg/P0001  & \u7_dout_reg[18]/P0001  ;
  assign n2561 = \u0_slt8_r_reg[17]/P0001  & ~\u2_ld_reg/P0001  ;
  assign n2562 = ~n2560 & ~n2561 ;
  assign n2563 = \u2_ld_reg/P0001  & \u7_dout_reg[17]/P0001  ;
  assign n2564 = \u0_slt8_r_reg[16]/P0001  & ~\u2_ld_reg/P0001  ;
  assign n2565 = ~n2563 & ~n2564 ;
  assign n2566 = \u2_ld_reg/P0001  & \u7_dout_reg[16]/P0001  ;
  assign n2567 = \u0_slt8_r_reg[15]/P0001  & ~\u2_ld_reg/P0001  ;
  assign n2568 = ~n2566 & ~n2567 ;
  assign n2569 = \u2_ld_reg/P0001  & \u7_dout_reg[15]/P0001  ;
  assign n2570 = \u0_slt8_r_reg[14]/P0001  & ~\u2_ld_reg/P0001  ;
  assign n2571 = ~n2569 & ~n2570 ;
  assign n2572 = \u2_ld_reg/P0001  & \u7_dout_reg[14]/P0001  ;
  assign n2573 = \u0_slt8_r_reg[13]/P0001  & ~\u2_ld_reg/P0001  ;
  assign n2574 = ~n2572 & ~n2573 ;
  assign n2575 = \u2_ld_reg/P0001  & \u7_dout_reg[13]/P0001  ;
  assign n2576 = \u0_slt8_r_reg[12]/P0001  & ~\u2_ld_reg/P0001  ;
  assign n2577 = ~n2575 & ~n2576 ;
  assign n2578 = \u2_ld_reg/P0001  & \u7_dout_reg[12]/P0001  ;
  assign n2579 = \u0_slt8_r_reg[11]/P0001  & ~\u2_ld_reg/P0001  ;
  assign n2580 = ~n2578 & ~n2579 ;
  assign n2581 = \u2_ld_reg/P0001  & \u7_dout_reg[11]/P0001  ;
  assign n2582 = \u0_slt8_r_reg[10]/P0001  & ~\u2_ld_reg/P0001  ;
  assign n2583 = ~n2581 & ~n2582 ;
  assign n2584 = \u2_ld_reg/P0001  & \u7_dout_reg[10]/P0001  ;
  assign n2585 = \u0_slt8_r_reg[9]/P0001  & ~\u2_ld_reg/P0001  ;
  assign n2586 = ~n2584 & ~n2585 ;
  assign n2587 = \u2_ld_reg/P0001  & \u7_dout_reg[9]/P0001  ;
  assign n2588 = \u0_slt8_r_reg[8]/P0001  & ~\u2_ld_reg/P0001  ;
  assign n2589 = ~n2587 & ~n2588 ;
  assign n2590 = \u2_ld_reg/P0001  & \u7_dout_reg[8]/P0001  ;
  assign n2591 = \u0_slt8_r_reg[7]/P0001  & ~\u2_ld_reg/P0001  ;
  assign n2592 = ~n2590 & ~n2591 ;
  assign n2593 = \u2_ld_reg/P0001  & \u7_dout_reg[7]/P0001  ;
  assign n2594 = \u0_slt8_r_reg[6]/P0001  & ~\u2_ld_reg/P0001  ;
  assign n2595 = ~n2593 & ~n2594 ;
  assign n2596 = \u2_ld_reg/P0001  & \u7_dout_reg[6]/P0001  ;
  assign n2597 = \u0_slt8_r_reg[5]/P0001  & ~\u2_ld_reg/P0001  ;
  assign n2598 = ~n2596 & ~n2597 ;
  assign n2599 = \u2_ld_reg/P0001  & \u7_dout_reg[5]/P0001  ;
  assign n2600 = \u0_slt8_r_reg[4]/P0001  & ~\u2_ld_reg/P0001  ;
  assign n2601 = ~n2599 & ~n2600 ;
  assign n2602 = \u2_ld_reg/P0001  & \u7_dout_reg[4]/P0001  ;
  assign n2603 = \u0_slt8_r_reg[3]/P0001  & ~\u2_ld_reg/P0001  ;
  assign n2604 = ~n2602 & ~n2603 ;
  assign n2605 = \u2_ld_reg/P0001  & \u7_dout_reg[3]/P0001  ;
  assign n2606 = \u0_slt8_r_reg[2]/P0001  & ~\u2_ld_reg/P0001  ;
  assign n2607 = ~n2605 & ~n2606 ;
  assign n2608 = \u2_ld_reg/P0001  & \u7_dout_reg[2]/P0001  ;
  assign n2609 = \u0_slt8_r_reg[1]/P0001  & ~\u2_ld_reg/P0001  ;
  assign n2610 = ~n2608 & ~n2609 ;
  assign n2611 = \u2_ld_reg/P0001  & \u7_dout_reg[1]/P0001  ;
  assign n2612 = \u0_slt8_r_reg[0]/P0001  & ~\u2_ld_reg/P0001  ;
  assign n2613 = ~n2611 & ~n2612 ;
  assign n2614 = \u2_ld_reg/P0001  & \u7_dout_reg[0]/P0001  ;
  assign n2615 = \u0_slt9_r_reg[19]/P0001  & ~\u2_ld_reg/P0001  ;
  assign n2616 = ~n2614 & ~n2615 ;
  assign n2617 = \u2_ld_reg/P0001  & \u8_dout_reg[19]/P0001  ;
  assign n2618 = \u0_slt9_r_reg[18]/P0001  & ~\u2_ld_reg/P0001  ;
  assign n2619 = ~n2617 & ~n2618 ;
  assign n2620 = \u2_ld_reg/P0001  & \u8_dout_reg[18]/P0001  ;
  assign n2621 = \u0_slt9_r_reg[17]/P0001  & ~\u2_ld_reg/P0001  ;
  assign n2622 = ~n2620 & ~n2621 ;
  assign n2623 = \u2_ld_reg/P0001  & \u8_dout_reg[17]/P0001  ;
  assign n2624 = \u0_slt9_r_reg[16]/P0001  & ~\u2_ld_reg/P0001  ;
  assign n2625 = ~n2623 & ~n2624 ;
  assign n2626 = \u2_ld_reg/P0001  & \u8_dout_reg[16]/P0001  ;
  assign n2627 = \u0_slt9_r_reg[15]/P0001  & ~\u2_ld_reg/P0001  ;
  assign n2628 = ~n2626 & ~n2627 ;
  assign n2629 = \u2_ld_reg/P0001  & \u8_dout_reg[15]/P0001  ;
  assign n2630 = \u0_slt9_r_reg[14]/P0001  & ~\u2_ld_reg/P0001  ;
  assign n2631 = ~n2629 & ~n2630 ;
  assign n2632 = \u2_ld_reg/P0001  & \u8_dout_reg[14]/P0001  ;
  assign n2633 = \u0_slt9_r_reg[13]/P0001  & ~\u2_ld_reg/P0001  ;
  assign n2634 = ~n2632 & ~n2633 ;
  assign n2635 = \u2_ld_reg/P0001  & \u8_dout_reg[13]/P0001  ;
  assign n2636 = \u0_slt9_r_reg[12]/P0001  & ~\u2_ld_reg/P0001  ;
  assign n2637 = ~n2635 & ~n2636 ;
  assign n2638 = \u2_ld_reg/P0001  & \u8_dout_reg[12]/P0001  ;
  assign n2639 = \u0_slt9_r_reg[11]/P0001  & ~\u2_ld_reg/P0001  ;
  assign n2640 = ~n2638 & ~n2639 ;
  assign n2641 = \u2_ld_reg/P0001  & \u8_dout_reg[11]/P0001  ;
  assign n2642 = \u0_slt9_r_reg[10]/P0001  & ~\u2_ld_reg/P0001  ;
  assign n2643 = ~n2641 & ~n2642 ;
  assign n2644 = \u2_ld_reg/P0001  & \u8_dout_reg[10]/P0001  ;
  assign n2645 = \u0_slt9_r_reg[9]/P0001  & ~\u2_ld_reg/P0001  ;
  assign n2646 = ~n2644 & ~n2645 ;
  assign n2647 = \u2_ld_reg/P0001  & \u8_dout_reg[9]/P0001  ;
  assign n2648 = \u0_slt9_r_reg[8]/P0001  & ~\u2_ld_reg/P0001  ;
  assign n2649 = ~n2647 & ~n2648 ;
  assign n2650 = \u2_ld_reg/P0001  & \u8_dout_reg[8]/P0001  ;
  assign n2651 = \u0_slt9_r_reg[7]/P0001  & ~\u2_ld_reg/P0001  ;
  assign n2652 = ~n2650 & ~n2651 ;
  assign n2653 = \u2_ld_reg/P0001  & \u8_dout_reg[7]/P0001  ;
  assign n2654 = \u0_slt9_r_reg[6]/P0001  & ~\u2_ld_reg/P0001  ;
  assign n2655 = ~n2653 & ~n2654 ;
  assign n2656 = \u2_ld_reg/P0001  & \u8_dout_reg[6]/P0001  ;
  assign n2657 = \u0_slt9_r_reg[5]/P0001  & ~\u2_ld_reg/P0001  ;
  assign n2658 = ~n2656 & ~n2657 ;
  assign n2659 = ~\dma_ack_i[0]_pad  & \dma_req_o[0]_pad  ;
  assign n2661 = \u13_occ0_r_reg[5]/NET0131  & \u3_status_reg[1]/P0001  ;
  assign n2662 = ~\u13_occ0_r_reg[4]/NET0131  & ~\u3_status_reg[0]/P0001  ;
  assign n2663 = ~n2661 & n2662 ;
  assign n2660 = ~\u13_occ0_r_reg[5]/NET0131  & ~\u3_status_reg[1]/P0001  ;
  assign n2664 = ~\u3_empty_reg/NET0131  & ~n2660 ;
  assign n2665 = ~n2663 & n2664 ;
  assign n2666 = \u13_occ0_r_reg[0]/NET0131  & ~n2665 ;
  assign n2667 = ~\dma_ack_i[0]_pad  & \u13_occ0_r_reg[6]/NET0131  ;
  assign n2668 = n2666 & n2667 ;
  assign n2669 = \u16_u0_dma_req_r1_reg/P0001  & n2668 ;
  assign n2670 = ~n2659 & ~n2669 ;
  assign n2671 = ~\dma_ack_i[1]_pad  & \dma_req_o[1]_pad  ;
  assign n2673 = \u13_occ0_r_reg[13]/NET0131  & \u4_status_reg[1]/P0001  ;
  assign n2674 = ~\u13_occ0_r_reg[12]/NET0131  & ~\u4_status_reg[0]/P0001  ;
  assign n2675 = ~n2673 & n2674 ;
  assign n2672 = ~\u13_occ0_r_reg[13]/NET0131  & ~\u4_status_reg[1]/P0001  ;
  assign n2676 = ~\u4_empty_reg/NET0131  & ~n2672 ;
  assign n2677 = ~n2675 & n2676 ;
  assign n2678 = \u13_occ0_r_reg[8]/NET0131  & ~n2677 ;
  assign n2679 = ~\dma_ack_i[1]_pad  & \u13_occ0_r_reg[14]/NET0131  ;
  assign n2680 = n2678 & n2679 ;
  assign n2681 = \u16_u1_dma_req_r1_reg/P0001  & n2680 ;
  assign n2682 = ~n2671 & ~n2681 ;
  assign n2683 = ~\dma_ack_i[2]_pad  & \dma_req_o[2]_pad  ;
  assign n2685 = \u13_occ0_r_reg[21]/NET0131  & \u5_status_reg[1]/P0001  ;
  assign n2686 = ~\u13_occ0_r_reg[20]/NET0131  & ~\u5_status_reg[0]/P0001  ;
  assign n2687 = ~n2685 & n2686 ;
  assign n2684 = ~\u13_occ0_r_reg[21]/NET0131  & ~\u5_status_reg[1]/P0001  ;
  assign n2688 = ~\u5_empty_reg/NET0131  & ~n2684 ;
  assign n2689 = ~n2687 & n2688 ;
  assign n2690 = \u13_occ0_r_reg[16]/NET0131  & ~n2689 ;
  assign n2691 = ~\dma_ack_i[2]_pad  & \u13_occ0_r_reg[22]/NET0131  ;
  assign n2692 = n2690 & n2691 ;
  assign n2693 = \u16_u2_dma_req_r1_reg/P0001  & n2692 ;
  assign n2694 = ~n2683 & ~n2693 ;
  assign n2695 = ~\dma_ack_i[3]_pad  & \dma_req_o[3]_pad  ;
  assign n2697 = \u13_occ0_r_reg[29]/NET0131  & \u6_status_reg[1]/P0001  ;
  assign n2698 = ~\u13_occ0_r_reg[28]/NET0131  & ~\u6_status_reg[0]/P0001  ;
  assign n2699 = ~n2697 & n2698 ;
  assign n2696 = ~\u13_occ0_r_reg[29]/NET0131  & ~\u6_status_reg[1]/P0001  ;
  assign n2700 = ~\u6_empty_reg/NET0131  & ~n2696 ;
  assign n2701 = ~n2699 & n2700 ;
  assign n2702 = \u13_occ0_r_reg[24]/NET0131  & ~n2701 ;
  assign n2703 = ~\dma_ack_i[3]_pad  & \u13_occ0_r_reg[30]/NET0131  ;
  assign n2704 = n2702 & n2703 ;
  assign n2705 = \u16_u3_dma_req_r1_reg/P0001  & n2704 ;
  assign n2706 = ~n2695 & ~n2705 ;
  assign n2707 = ~\dma_ack_i[4]_pad  & \dma_req_o[4]_pad  ;
  assign n2709 = \u13_occ1_r_reg[5]/NET0131  & \u7_status_reg[1]/P0001  ;
  assign n2710 = ~\u13_occ1_r_reg[4]/NET0131  & ~\u7_status_reg[0]/P0001  ;
  assign n2711 = ~n2709 & n2710 ;
  assign n2708 = ~\u13_occ1_r_reg[5]/NET0131  & ~\u7_status_reg[1]/P0001  ;
  assign n2712 = ~\u7_empty_reg/NET0131  & ~n2708 ;
  assign n2713 = ~n2711 & n2712 ;
  assign n2714 = \u13_occ1_r_reg[0]/NET0131  & ~n2713 ;
  assign n2715 = ~\dma_ack_i[4]_pad  & \u13_occ1_r_reg[6]/NET0131  ;
  assign n2716 = n2714 & n2715 ;
  assign n2717 = \u16_u4_dma_req_r1_reg/P0001  & n2716 ;
  assign n2718 = ~n2707 & ~n2717 ;
  assign n2719 = ~\dma_ack_i[5]_pad  & \dma_req_o[5]_pad  ;
  assign n2721 = \u13_occ1_r_reg[13]/NET0131  & \u8_status_reg[1]/P0001  ;
  assign n2722 = ~\u13_occ1_r_reg[12]/NET0131  & ~\u8_status_reg[0]/P0001  ;
  assign n2723 = ~n2721 & n2722 ;
  assign n2720 = ~\u13_occ1_r_reg[13]/NET0131  & ~\u8_status_reg[1]/P0001  ;
  assign n2724 = ~\u8_empty_reg/NET0131  & ~n2720 ;
  assign n2725 = ~n2723 & n2724 ;
  assign n2726 = \u13_occ1_r_reg[8]/NET0131  & ~n2725 ;
  assign n2727 = ~\dma_ack_i[5]_pad  & \u13_occ1_r_reg[14]/NET0131  ;
  assign n2728 = n2726 & n2727 ;
  assign n2729 = \u16_u5_dma_req_r1_reg/P0001  & n2728 ;
  assign n2730 = ~n2719 & ~n2729 ;
  assign n2731 = \u2_ld_reg/P0001  & \u8_dout_reg[5]/P0001  ;
  assign n2732 = \u0_slt9_r_reg[4]/P0001  & ~\u2_ld_reg/P0001  ;
  assign n2733 = ~n2731 & ~n2732 ;
  assign n2734 = ~\u13_ints_r_reg[11]/NET0131  & ~\u20_int_set_reg[0]/NET0131  ;
  assign n2735 = wb_cyc_i_pad & wb_stb_i_pad ;
  assign n2736 = ~\u12_re2_reg/NET0131  & ~wb_we_i_pad ;
  assign n2737 = n2735 & n2736 ;
  assign n2738 = \u12_re1_reg/P0001  & n2737 ;
  assign n2739 = ~\wb_addr_i[5]_pad  & ~\wb_addr_i[6]_pad  ;
  assign n2740 = ~\wb_addr_i[2]_pad  & \wb_addr_i[3]_pad  ;
  assign n2741 = \wb_addr_i[4]_pad  & n2740 ;
  assign n2742 = n2739 & n2741 ;
  assign n2743 = n2738 & n2742 ;
  assign n2744 = ~n2734 & ~n2743 ;
  assign n2745 = ~\u13_ints_r_reg[14]/NET0131  & ~\u21_int_set_reg[0]/NET0131  ;
  assign n2746 = ~n2743 & ~n2745 ;
  assign n2747 = ~\u13_ints_r_reg[17]/NET0131  & ~\u22_int_set_reg[0]/NET0131  ;
  assign n2748 = ~n2743 & ~n2747 ;
  assign n2749 = ~\u13_ints_r_reg[2]/NET0131  & ~\u17_int_set_reg[0]/NET0131  ;
  assign n2750 = ~n2743 & ~n2749 ;
  assign n2751 = ~\u13_ints_r_reg[5]/NET0131  & ~\u18_int_set_reg[0]/NET0131  ;
  assign n2752 = ~n2743 & ~n2751 ;
  assign n2753 = ~\u13_ints_r_reg[8]/NET0131  & ~\u19_int_set_reg[0]/NET0131  ;
  assign n2754 = ~n2743 & ~n2753 ;
  assign n2755 = \u2_ld_reg/P0001  & \u8_dout_reg[4]/P0001  ;
  assign n2756 = \u0_slt9_r_reg[3]/P0001  & ~\u2_ld_reg/P0001  ;
  assign n2757 = ~n2755 & ~n2756 ;
  assign n2758 = \u14_u1_en_out_l_reg/NET0131  & \valid_s_reg/NET0131  ;
  assign n2759 = ~\u14_u1_en_out_l2_reg/P0001  & n2758 ;
  assign n2760 = ~\u13_occ0_r_reg[10]/NET0131  & ~\u13_occ0_r_reg[11]/NET0131  ;
  assign n2761 = ~\u4_rp_reg[0]/P0001  & n2760 ;
  assign n2762 = n2759 & ~n2761 ;
  assign n2763 = \u4_rp_reg[1]/NET0131  & n2762 ;
  assign n2764 = ~\u4_rp_reg[2]/NET0131  & ~n2763 ;
  assign n2765 = \u4_rp_reg[1]/NET0131  & \u4_rp_reg[2]/NET0131  ;
  assign n2766 = n2762 & n2765 ;
  assign n2767 = \u13_occ0_r_reg[8]/NET0131  & ~n2766 ;
  assign n2768 = ~n2764 & n2767 ;
  assign n2769 = \u14_u2_en_out_l_reg/NET0131  & \valid_s_reg/NET0131  ;
  assign n2770 = ~\u14_u2_en_out_l2_reg/P0001  & n2769 ;
  assign n2771 = ~\u13_occ0_r_reg[18]/NET0131  & ~\u13_occ0_r_reg[19]/NET0131  ;
  assign n2772 = ~\u5_rp_reg[0]/P0001  & n2771 ;
  assign n2773 = n2770 & ~n2772 ;
  assign n2774 = \u5_rp_reg[1]/NET0131  & n2773 ;
  assign n2775 = ~\u5_rp_reg[2]/NET0131  & ~n2774 ;
  assign n2776 = \u5_rp_reg[1]/NET0131  & \u5_rp_reg[2]/NET0131  ;
  assign n2777 = n2773 & n2776 ;
  assign n2778 = \u13_occ0_r_reg[16]/NET0131  & ~n2777 ;
  assign n2779 = ~n2775 & n2778 ;
  assign n2780 = \u8_rp_reg[1]/NET0131  & n2162 ;
  assign n2781 = ~\u8_rp_reg[2]/NET0131  & ~n2780 ;
  assign n2782 = \u13_occ1_r_reg[8]/NET0131  & ~n2164 ;
  assign n2783 = ~n2781 & n2782 ;
  assign n2784 = ~\u13_occ0_r_reg[2]/NET0131  & ~\u13_occ0_r_reg[3]/NET0131  ;
  assign n2785 = ~\u3_rp_reg[0]/P0001  & n2784 ;
  assign n2786 = ~\u14_u0_en_out_l2_reg/P0001  & \u14_u0_en_out_l_reg/NET0131  ;
  assign n2787 = \valid_s_reg/NET0131  & n2786 ;
  assign n2788 = ~n2785 & n2787 ;
  assign n2789 = \u3_rp_reg[1]/NET0131  & n2788 ;
  assign n2791 = \u3_rp_reg[2]/NET0131  & n2789 ;
  assign n2790 = ~\u3_rp_reg[2]/NET0131  & ~n2789 ;
  assign n2792 = \u13_occ0_r_reg[0]/NET0131  & ~n2790 ;
  assign n2793 = ~n2791 & n2792 ;
  assign n2794 = \u14_u3_en_out_l_reg/NET0131  & \valid_s_reg/NET0131  ;
  assign n2795 = ~\u14_u3_en_out_l2_reg/P0001  & n2794 ;
  assign n2796 = ~\u13_occ0_r_reg[26]/NET0131  & ~\u13_occ0_r_reg[27]/NET0131  ;
  assign n2797 = ~\u6_rp_reg[0]/P0001  & n2796 ;
  assign n2798 = n2795 & ~n2797 ;
  assign n2799 = \u6_rp_reg[1]/NET0131  & n2798 ;
  assign n2800 = ~\u6_rp_reg[2]/NET0131  & ~n2799 ;
  assign n2801 = \u6_rp_reg[1]/NET0131  & \u6_rp_reg[2]/NET0131  ;
  assign n2802 = n2798 & n2801 ;
  assign n2803 = \u13_occ0_r_reg[24]/NET0131  & ~n2802 ;
  assign n2804 = ~n2800 & n2803 ;
  assign n2805 = ~\u13_occ1_r_reg[2]/NET0131  & ~\u13_occ1_r_reg[3]/NET0131  ;
  assign n2806 = ~\u7_rp_reg[0]/P0001  & n2805 ;
  assign n2807 = \u14_u4_en_out_l_reg/NET0131  & \valid_s_reg/NET0131  ;
  assign n2808 = ~\u14_u4_en_out_l2_reg/P0001  & n2807 ;
  assign n2809 = ~n2806 & n2808 ;
  assign n2810 = \u7_rp_reg[1]/NET0131  & n2809 ;
  assign n2812 = \u7_rp_reg[2]/NET0131  & n2810 ;
  assign n2811 = ~\u7_rp_reg[2]/NET0131  & ~n2810 ;
  assign n2813 = \u13_occ1_r_reg[0]/NET0131  & ~n2811 ;
  assign n2814 = ~n2812 & n2813 ;
  assign n2816 = \u3_rp_reg[3]/NET0131  & n2791 ;
  assign n2815 = ~\u3_rp_reg[3]/NET0131  & ~n2791 ;
  assign n2817 = \u13_occ0_r_reg[0]/NET0131  & ~n2815 ;
  assign n2818 = ~n2816 & n2817 ;
  assign n2820 = \u4_rp_reg[3]/NET0131  & n2766 ;
  assign n2819 = ~\u4_rp_reg[3]/NET0131  & ~n2766 ;
  assign n2821 = \u13_occ0_r_reg[8]/NET0131  & ~n2819 ;
  assign n2822 = ~n2820 & n2821 ;
  assign n2823 = ~\u13_ints_r_reg[20]/NET0131  & ~\u23_int_set_reg[0]/NET0131  ;
  assign n2824 = ~n2743 & ~n2823 ;
  assign n2825 = ~\u13_ints_r_reg[23]/NET0131  & ~\u24_int_set_reg[0]/NET0131  ;
  assign n2826 = ~n2743 & ~n2825 ;
  assign n2827 = ~\u13_ints_r_reg[26]/NET0131  & ~\u25_int_set_reg[0]/NET0131  ;
  assign n2828 = ~n2743 & ~n2827 ;
  assign n2830 = \u5_rp_reg[3]/NET0131  & n2777 ;
  assign n2829 = ~\u5_rp_reg[3]/NET0131  & ~n2777 ;
  assign n2831 = \u13_occ0_r_reg[16]/NET0131  & ~n2829 ;
  assign n2832 = ~n2830 & n2831 ;
  assign n2834 = \u6_rp_reg[3]/NET0131  & n2802 ;
  assign n2833 = ~\u6_rp_reg[3]/NET0131  & ~n2802 ;
  assign n2835 = \u13_occ0_r_reg[24]/NET0131  & ~n2833 ;
  assign n2836 = ~n2834 & n2835 ;
  assign n2838 = \u7_rp_reg[3]/NET0131  & n2812 ;
  assign n2837 = ~\u7_rp_reg[3]/NET0131  & ~n2812 ;
  assign n2839 = \u13_occ1_r_reg[0]/NET0131  & ~n2837 ;
  assign n2840 = ~n2838 & n2839 ;
  assign n2841 = ~\u8_rp_reg[1]/NET0131  & ~n2162 ;
  assign n2842 = \u13_occ1_r_reg[8]/NET0131  & ~n2780 ;
  assign n2843 = ~n2841 & n2842 ;
  assign n2844 = ~\u3_rp_reg[1]/NET0131  & ~n2788 ;
  assign n2845 = \u13_occ0_r_reg[0]/NET0131  & ~n2789 ;
  assign n2846 = ~n2844 & n2845 ;
  assign n2847 = ~\u4_rp_reg[1]/NET0131  & ~n2762 ;
  assign n2848 = \u13_occ0_r_reg[8]/NET0131  & ~n2763 ;
  assign n2849 = ~n2847 & n2848 ;
  assign n2850 = ~\u5_rp_reg[1]/NET0131  & ~n2773 ;
  assign n2851 = \u13_occ0_r_reg[16]/NET0131  & ~n2774 ;
  assign n2852 = ~n2850 & n2851 ;
  assign n2853 = ~\u6_rp_reg[1]/NET0131  & ~n2798 ;
  assign n2854 = \u13_occ0_r_reg[24]/NET0131  & ~n2799 ;
  assign n2855 = ~n2853 & n2854 ;
  assign n2856 = ~\u7_rp_reg[1]/NET0131  & ~n2809 ;
  assign n2857 = \u13_occ1_r_reg[0]/NET0131  & ~n2810 ;
  assign n2858 = ~n2856 & n2857 ;
  assign n2859 = \u2_ld_reg/P0001  & \u8_dout_reg[3]/P0001  ;
  assign n2860 = \u0_slt9_r_reg[2]/P0001  & ~\u2_ld_reg/P0001  ;
  assign n2861 = ~n2859 & ~n2860 ;
  assign n2862 = suspended_o_pad & \u13_resume_req_reg/P0001  ;
  assign n2863 = ~\u2_sync_resume_reg/NET0131  & ~n2862 ;
  assign n2864 = \u2_res_cnt_reg[0]/P0001  & ~\u2_res_cnt_reg[1]/P0001  ;
  assign n2865 = \u2_res_cnt_reg[2]/P0001  & ~\u2_res_cnt_reg[3]/P0001  ;
  assign n2866 = n2864 & n2865 ;
  assign n2867 = ~n2863 & ~n2866 ;
  assign n2868 = n2159 & n2160 ;
  assign n2870 = \u8_rp_reg[0]/P0001  & n2868 ;
  assign n2869 = ~\u8_rp_reg[0]/P0001  & ~n2868 ;
  assign n2871 = \u13_occ1_r_reg[8]/NET0131  & ~n2869 ;
  assign n2872 = ~n2870 & n2871 ;
  assign n2873 = n2784 & n2787 ;
  assign n2875 = \u3_rp_reg[0]/P0001  & n2873 ;
  assign n2874 = ~\u3_rp_reg[0]/P0001  & ~n2873 ;
  assign n2876 = \u13_occ0_r_reg[0]/NET0131  & ~n2874 ;
  assign n2877 = ~n2875 & n2876 ;
  assign n2878 = n2759 & n2760 ;
  assign n2880 = \u4_rp_reg[0]/P0001  & n2878 ;
  assign n2879 = ~\u4_rp_reg[0]/P0001  & ~n2878 ;
  assign n2881 = \u13_occ0_r_reg[8]/NET0131  & ~n2879 ;
  assign n2882 = ~n2880 & n2881 ;
  assign n2883 = n2770 & n2771 ;
  assign n2885 = \u5_rp_reg[0]/P0001  & n2883 ;
  assign n2884 = ~\u5_rp_reg[0]/P0001  & ~n2883 ;
  assign n2886 = \u13_occ0_r_reg[16]/NET0131  & ~n2884 ;
  assign n2887 = ~n2885 & n2886 ;
  assign n2888 = n2795 & n2796 ;
  assign n2890 = \u6_rp_reg[0]/P0001  & n2888 ;
  assign n2889 = ~\u6_rp_reg[0]/P0001  & ~n2888 ;
  assign n2891 = \u13_occ0_r_reg[24]/NET0131  & ~n2889 ;
  assign n2892 = ~n2890 & n2891 ;
  assign n2893 = n2805 & n2808 ;
  assign n2895 = \u7_rp_reg[0]/P0001  & n2893 ;
  assign n2894 = ~\u7_rp_reg[0]/P0001  & ~n2893 ;
  assign n2896 = \u13_occ1_r_reg[0]/NET0131  & ~n2894 ;
  assign n2897 = ~n2895 & n2896 ;
  assign n2898 = \u13_occ0_r_reg[8]/NET0131  & ~n2759 ;
  assign n2899 = \u4_dout_reg[0]/P0001  & n2898 ;
  assign n2900 = \u4_mem_reg[3][0]/NET0131  & n2765 ;
  assign n2901 = ~\u4_rp_reg[1]/NET0131  & \u4_rp_reg[2]/NET0131  ;
  assign n2902 = \u4_mem_reg[2][0]/NET0131  & n2901 ;
  assign n2907 = ~n2900 & ~n2902 ;
  assign n2903 = \u4_rp_reg[1]/NET0131  & ~\u4_rp_reg[2]/NET0131  ;
  assign n2904 = \u4_mem_reg[1][0]/NET0131  & n2903 ;
  assign n2905 = ~\u4_rp_reg[1]/NET0131  & ~\u4_rp_reg[2]/NET0131  ;
  assign n2906 = \u4_mem_reg[0][0]/NET0131  & n2905 ;
  assign n2908 = ~n2904 & ~n2906 ;
  assign n2909 = n2907 & n2908 ;
  assign n2910 = ~\u13_occ0_r_reg[10]/NET0131  & \u13_occ0_r_reg[11]/NET0131  ;
  assign n2911 = \u13_occ0_r_reg[8]/NET0131  & n2910 ;
  assign n2912 = n2759 & n2911 ;
  assign n2913 = ~n2909 & n2912 ;
  assign n2914 = ~n2899 & ~n2913 ;
  assign n2915 = \u4_dout_reg[1]/P0001  & n2898 ;
  assign n2916 = \u4_mem_reg[3][1]/NET0131  & n2765 ;
  assign n2917 = \u4_mem_reg[2][1]/NET0131  & n2901 ;
  assign n2920 = ~n2916 & ~n2917 ;
  assign n2918 = \u4_mem_reg[1][1]/NET0131  & n2903 ;
  assign n2919 = \u4_mem_reg[0][1]/NET0131  & n2905 ;
  assign n2921 = ~n2918 & ~n2919 ;
  assign n2922 = n2920 & n2921 ;
  assign n2923 = n2912 & ~n2922 ;
  assign n2924 = ~n2915 & ~n2923 ;
  assign n2925 = \u13_occ0_r_reg[16]/NET0131  & ~n2770 ;
  assign n2926 = \u5_dout_reg[0]/P0001  & n2925 ;
  assign n2927 = \u5_mem_reg[3][0]/NET0131  & n2776 ;
  assign n2928 = \u5_rp_reg[1]/NET0131  & ~\u5_rp_reg[2]/NET0131  ;
  assign n2929 = \u5_mem_reg[1][0]/NET0131  & n2928 ;
  assign n2934 = ~n2927 & ~n2929 ;
  assign n2930 = ~\u5_rp_reg[1]/NET0131  & \u5_rp_reg[2]/NET0131  ;
  assign n2931 = \u5_mem_reg[2][0]/NET0131  & n2930 ;
  assign n2932 = ~\u5_rp_reg[1]/NET0131  & ~\u5_rp_reg[2]/NET0131  ;
  assign n2933 = \u5_mem_reg[0][0]/NET0131  & n2932 ;
  assign n2935 = ~n2931 & ~n2933 ;
  assign n2936 = n2934 & n2935 ;
  assign n2937 = ~\u13_occ0_r_reg[18]/NET0131  & \u13_occ0_r_reg[19]/NET0131  ;
  assign n2938 = \u13_occ0_r_reg[16]/NET0131  & n2937 ;
  assign n2939 = n2770 & n2938 ;
  assign n2940 = ~n2936 & n2939 ;
  assign n2941 = ~n2926 & ~n2940 ;
  assign n2942 = \u5_dout_reg[1]/P0001  & n2925 ;
  assign n2943 = \u5_mem_reg[3][1]/NET0131  & n2776 ;
  assign n2944 = \u5_mem_reg[1][1]/NET0131  & n2928 ;
  assign n2947 = ~n2943 & ~n2944 ;
  assign n2945 = \u5_mem_reg[2][1]/NET0131  & n2930 ;
  assign n2946 = \u5_mem_reg[0][1]/NET0131  & n2932 ;
  assign n2948 = ~n2945 & ~n2946 ;
  assign n2949 = n2947 & n2948 ;
  assign n2950 = n2939 & ~n2949 ;
  assign n2951 = ~n2942 & ~n2950 ;
  assign n2952 = \u13_occ0_r_reg[24]/NET0131  & ~n2795 ;
  assign n2953 = \u6_dout_reg[0]/P0001  & n2952 ;
  assign n2954 = \u6_mem_reg[3][0]/NET0131  & n2801 ;
  assign n2955 = ~\u6_rp_reg[1]/NET0131  & \u6_rp_reg[2]/NET0131  ;
  assign n2956 = \u6_mem_reg[2][0]/NET0131  & n2955 ;
  assign n2961 = ~n2954 & ~n2956 ;
  assign n2957 = \u6_rp_reg[1]/NET0131  & ~\u6_rp_reg[2]/NET0131  ;
  assign n2958 = \u6_mem_reg[1][0]/NET0131  & n2957 ;
  assign n2959 = ~\u6_rp_reg[1]/NET0131  & ~\u6_rp_reg[2]/NET0131  ;
  assign n2960 = \u6_mem_reg[0][0]/NET0131  & n2959 ;
  assign n2962 = ~n2958 & ~n2960 ;
  assign n2963 = n2961 & n2962 ;
  assign n2964 = ~\u13_occ0_r_reg[26]/NET0131  & \u13_occ0_r_reg[27]/NET0131  ;
  assign n2965 = \u13_occ0_r_reg[24]/NET0131  & n2964 ;
  assign n2966 = n2795 & n2965 ;
  assign n2967 = ~n2963 & n2966 ;
  assign n2968 = ~n2953 & ~n2967 ;
  assign n2969 = \u6_dout_reg[1]/P0001  & n2952 ;
  assign n2970 = \u6_mem_reg[2][1]/NET0131  & n2955 ;
  assign n2971 = \u6_mem_reg[1][1]/NET0131  & n2957 ;
  assign n2974 = ~n2970 & ~n2971 ;
  assign n2972 = \u6_mem_reg[3][1]/NET0131  & n2801 ;
  assign n2973 = \u6_mem_reg[0][1]/NET0131  & n2959 ;
  assign n2975 = ~n2972 & ~n2973 ;
  assign n2976 = n2974 & n2975 ;
  assign n2977 = n2966 & ~n2976 ;
  assign n2978 = ~n2969 & ~n2977 ;
  assign n2979 = \u13_occ1_r_reg[0]/NET0131  & ~n2808 ;
  assign n2980 = \u7_dout_reg[0]/P0001  & n2979 ;
  assign n2981 = \u7_rp_reg[1]/NET0131  & \u7_rp_reg[2]/NET0131  ;
  assign n2982 = \u7_mem_reg[3][0]/NET0131  & n2981 ;
  assign n2983 = ~\u7_rp_reg[1]/NET0131  & \u7_rp_reg[2]/NET0131  ;
  assign n2984 = \u7_mem_reg[2][0]/NET0131  & n2983 ;
  assign n2989 = ~n2982 & ~n2984 ;
  assign n2985 = \u7_rp_reg[1]/NET0131  & ~\u7_rp_reg[2]/NET0131  ;
  assign n2986 = \u7_mem_reg[1][0]/NET0131  & n2985 ;
  assign n2987 = ~\u7_rp_reg[1]/NET0131  & ~\u7_rp_reg[2]/NET0131  ;
  assign n2988 = \u7_mem_reg[0][0]/NET0131  & n2987 ;
  assign n2990 = ~n2986 & ~n2988 ;
  assign n2991 = n2989 & n2990 ;
  assign n2992 = ~\u13_occ1_r_reg[2]/NET0131  & \u13_occ1_r_reg[3]/NET0131  ;
  assign n2993 = \u13_occ1_r_reg[0]/NET0131  & n2992 ;
  assign n2994 = n2808 & n2993 ;
  assign n2995 = ~n2991 & n2994 ;
  assign n2996 = ~n2980 & ~n2995 ;
  assign n2997 = \u7_dout_reg[1]/P0001  & n2979 ;
  assign n2998 = \u7_mem_reg[3][1]/NET0131  & n2981 ;
  assign n2999 = \u7_mem_reg[2][1]/NET0131  & n2983 ;
  assign n3002 = ~n2998 & ~n2999 ;
  assign n3000 = \u7_mem_reg[1][1]/NET0131  & n2985 ;
  assign n3001 = \u7_mem_reg[0][1]/NET0131  & n2987 ;
  assign n3003 = ~n3000 & ~n3001 ;
  assign n3004 = n3002 & n3003 ;
  assign n3005 = n2994 & ~n3004 ;
  assign n3006 = ~n2997 & ~n3005 ;
  assign n3007 = \u13_occ0_r_reg[0]/NET0131  & ~n2787 ;
  assign n3008 = \u3_dout_reg[0]/P0001  & n3007 ;
  assign n3009 = \u3_rp_reg[1]/NET0131  & \u3_rp_reg[2]/NET0131  ;
  assign n3010 = \u3_mem_reg[3][0]/NET0131  & n3009 ;
  assign n3011 = ~\u3_rp_reg[1]/NET0131  & \u3_rp_reg[2]/NET0131  ;
  assign n3012 = \u3_mem_reg[2][0]/NET0131  & n3011 ;
  assign n3017 = ~n3010 & ~n3012 ;
  assign n3013 = \u3_rp_reg[1]/NET0131  & ~\u3_rp_reg[2]/NET0131  ;
  assign n3014 = \u3_mem_reg[1][0]/NET0131  & n3013 ;
  assign n3015 = ~\u3_rp_reg[1]/NET0131  & ~\u3_rp_reg[2]/NET0131  ;
  assign n3016 = \u3_mem_reg[0][0]/NET0131  & n3015 ;
  assign n3018 = ~n3014 & ~n3016 ;
  assign n3019 = n3017 & n3018 ;
  assign n3020 = ~\u13_occ0_r_reg[2]/NET0131  & \u13_occ0_r_reg[3]/NET0131  ;
  assign n3021 = \u13_occ0_r_reg[0]/NET0131  & n3020 ;
  assign n3022 = n2787 & n3021 ;
  assign n3023 = ~n3019 & n3022 ;
  assign n3024 = ~n3008 & ~n3023 ;
  assign n3025 = \u13_occ1_r_reg[8]/NET0131  & ~n2159 ;
  assign n3026 = \u8_dout_reg[0]/P0001  & n3025 ;
  assign n3027 = \u8_mem_reg[3][0]/NET0131  & n2163 ;
  assign n3028 = ~\u8_rp_reg[1]/NET0131  & \u8_rp_reg[2]/NET0131  ;
  assign n3029 = \u8_mem_reg[2][0]/NET0131  & n3028 ;
  assign n3034 = ~n3027 & ~n3029 ;
  assign n3030 = \u8_rp_reg[1]/NET0131  & ~\u8_rp_reg[2]/NET0131  ;
  assign n3031 = \u8_mem_reg[1][0]/NET0131  & n3030 ;
  assign n3032 = ~\u8_rp_reg[1]/NET0131  & ~\u8_rp_reg[2]/NET0131  ;
  assign n3033 = \u8_mem_reg[0][0]/NET0131  & n3032 ;
  assign n3035 = ~n3031 & ~n3033 ;
  assign n3036 = n3034 & n3035 ;
  assign n3037 = ~\u13_occ1_r_reg[10]/NET0131  & \u13_occ1_r_reg[11]/NET0131  ;
  assign n3038 = \u13_occ1_r_reg[8]/NET0131  & n3037 ;
  assign n3039 = n2159 & n3038 ;
  assign n3040 = ~n3036 & n3039 ;
  assign n3041 = ~n3026 & ~n3040 ;
  assign n3042 = \u3_dout_reg[1]/P0001  & n3007 ;
  assign n3043 = \u3_mem_reg[1][1]/NET0131  & n3013 ;
  assign n3044 = \u3_mem_reg[2][1]/NET0131  & n3011 ;
  assign n3047 = ~n3043 & ~n3044 ;
  assign n3045 = \u3_mem_reg[3][1]/NET0131  & n3009 ;
  assign n3046 = \u3_mem_reg[0][1]/NET0131  & n3015 ;
  assign n3048 = ~n3045 & ~n3046 ;
  assign n3049 = n3047 & n3048 ;
  assign n3050 = n3022 & ~n3049 ;
  assign n3051 = ~n3042 & ~n3050 ;
  assign n3052 = \u8_dout_reg[1]/P0001  & n3025 ;
  assign n3053 = \u8_mem_reg[3][1]/NET0131  & n2163 ;
  assign n3054 = \u8_mem_reg[2][1]/NET0131  & n3028 ;
  assign n3057 = ~n3053 & ~n3054 ;
  assign n3055 = \u8_mem_reg[1][1]/NET0131  & n3030 ;
  assign n3056 = \u8_mem_reg[0][1]/NET0131  & n3032 ;
  assign n3058 = ~n3055 & ~n3056 ;
  assign n3059 = n3057 & n3058 ;
  assign n3060 = n3039 & ~n3059 ;
  assign n3061 = ~n3052 & ~n3060 ;
  assign n3062 = \in_valid_s_reg[2]/NET0131  & \u14_u8_en_out_l_reg/NET0131  ;
  assign n3063 = ~\u14_u8_en_out_l2_reg/P0001  & n3062 ;
  assign n3064 = ~\u13_icc_r_reg[18]/NET0131  & ~\u13_icc_r_reg[19]/NET0131  ;
  assign n3065 = ~\u11_wp_reg[0]/NET0131  & n3064 ;
  assign n3066 = n3063 & ~n3065 ;
  assign n3067 = \u11_wp_reg[1]/P0001  & n3066 ;
  assign n3069 = ~\u11_wp_reg[2]/P0001  & ~n3067 ;
  assign n3068 = \u11_wp_reg[2]/P0001  & n3067 ;
  assign n3070 = \u13_icc_r_reg[16]/NET0131  & ~n3068 ;
  assign n3071 = ~n3069 & n3070 ;
  assign n3081 = \u4_mem_reg[2][22]/NET0131  & n2901 ;
  assign n3085 = \u4_rp_reg[0]/P0001  & ~n3081 ;
  assign n3084 = \u4_mem_reg[0][22]/NET0131  & n2905 ;
  assign n3082 = \u4_mem_reg[3][22]/NET0131  & n2765 ;
  assign n3083 = \u4_mem_reg[1][22]/NET0131  & n2903 ;
  assign n3086 = ~n3082 & ~n3083 ;
  assign n3087 = ~n3084 & n3086 ;
  assign n3088 = n3085 & n3087 ;
  assign n3073 = \u4_mem_reg[3][6]/NET0131  & n2765 ;
  assign n3074 = \u4_mem_reg[2][6]/NET0131  & n2901 ;
  assign n3077 = ~n3073 & ~n3074 ;
  assign n3075 = \u4_mem_reg[0][6]/NET0131  & n2905 ;
  assign n3076 = \u4_mem_reg[1][6]/NET0131  & n2903 ;
  assign n3078 = ~n3075 & ~n3076 ;
  assign n3079 = n3077 & n3078 ;
  assign n3080 = ~\u4_rp_reg[0]/P0001  & n3079 ;
  assign n3089 = n2760 & ~n3080 ;
  assign n3090 = ~n3088 & n3089 ;
  assign n3099 = \u13_occ0_r_reg[10]/NET0131  & ~\u13_occ0_r_reg[11]/NET0131  ;
  assign n3100 = \u4_mem_reg[3][8]/NET0131  & n2765 ;
  assign n3101 = \u4_mem_reg[2][8]/NET0131  & n2901 ;
  assign n3104 = ~n3100 & ~n3101 ;
  assign n3102 = \u4_mem_reg[0][8]/NET0131  & n2905 ;
  assign n3103 = \u4_mem_reg[1][8]/NET0131  & n2903 ;
  assign n3105 = ~n3102 & ~n3103 ;
  assign n3106 = n3104 & n3105 ;
  assign n3107 = n3099 & ~n3106 ;
  assign n3091 = \u4_mem_reg[3][10]/NET0131  & n2765 ;
  assign n3092 = \u4_mem_reg[2][10]/NET0131  & n2901 ;
  assign n3095 = ~n3091 & ~n3092 ;
  assign n3093 = \u4_mem_reg[0][10]/NET0131  & n2905 ;
  assign n3094 = \u4_mem_reg[1][10]/NET0131  & n2903 ;
  assign n3096 = ~n3093 & ~n3094 ;
  assign n3097 = n3095 & n3096 ;
  assign n3098 = n2910 & ~n3097 ;
  assign n3108 = n2759 & ~n3098 ;
  assign n3109 = ~n3107 & n3108 ;
  assign n3110 = ~n3090 & n3109 ;
  assign n3072 = ~\u4_dout_reg[10]/P0001  & ~n2759 ;
  assign n3111 = \u13_occ0_r_reg[8]/NET0131  & ~n3072 ;
  assign n3112 = ~n3110 & n3111 ;
  assign n3122 = \u4_mem_reg[2][23]/NET0131  & n2901 ;
  assign n3126 = \u4_rp_reg[0]/P0001  & ~n3122 ;
  assign n3125 = \u4_mem_reg[0][23]/NET0131  & n2905 ;
  assign n3123 = \u4_mem_reg[3][23]/NET0131  & n2765 ;
  assign n3124 = \u4_mem_reg[1][23]/NET0131  & n2903 ;
  assign n3127 = ~n3123 & ~n3124 ;
  assign n3128 = ~n3125 & n3127 ;
  assign n3129 = n3126 & n3128 ;
  assign n3114 = \u4_mem_reg[1][7]/NET0131  & n2903 ;
  assign n3115 = \u4_mem_reg[2][7]/NET0131  & n2901 ;
  assign n3118 = ~n3114 & ~n3115 ;
  assign n3116 = \u4_mem_reg[3][7]/NET0131  & n2765 ;
  assign n3117 = \u4_mem_reg[0][7]/NET0131  & n2905 ;
  assign n3119 = ~n3116 & ~n3117 ;
  assign n3120 = n3118 & n3119 ;
  assign n3121 = ~\u4_rp_reg[0]/P0001  & n3120 ;
  assign n3130 = n2760 & ~n3121 ;
  assign n3131 = ~n3129 & n3130 ;
  assign n3140 = \u4_mem_reg[1][9]/NET0131  & n2903 ;
  assign n3141 = \u4_mem_reg[3][9]/NET0131  & n2765 ;
  assign n3144 = ~n3140 & ~n3141 ;
  assign n3142 = \u4_mem_reg[2][9]/NET0131  & n2901 ;
  assign n3143 = \u4_mem_reg[0][9]/NET0131  & n2905 ;
  assign n3145 = ~n3142 & ~n3143 ;
  assign n3146 = n3144 & n3145 ;
  assign n3147 = n3099 & ~n3146 ;
  assign n3132 = \u4_mem_reg[3][11]/NET0131  & n2765 ;
  assign n3133 = \u4_mem_reg[1][11]/NET0131  & n2903 ;
  assign n3136 = ~n3132 & ~n3133 ;
  assign n3134 = \u4_mem_reg[2][11]/NET0131  & n2901 ;
  assign n3135 = \u4_mem_reg[0][11]/NET0131  & n2905 ;
  assign n3137 = ~n3134 & ~n3135 ;
  assign n3138 = n3136 & n3137 ;
  assign n3139 = n2910 & ~n3138 ;
  assign n3148 = n2759 & ~n3139 ;
  assign n3149 = ~n3147 & n3148 ;
  assign n3150 = ~n3131 & n3149 ;
  assign n3113 = ~\u4_dout_reg[11]/P0001  & ~n2759 ;
  assign n3151 = \u13_occ0_r_reg[8]/NET0131  & ~n3113 ;
  assign n3152 = ~n3150 & n3151 ;
  assign n3155 = \u4_mem_reg[2][24]/NET0131  & n2901 ;
  assign n3159 = \u4_rp_reg[0]/P0001  & ~n3155 ;
  assign n3158 = \u4_mem_reg[0][24]/NET0131  & n2905 ;
  assign n3156 = \u4_mem_reg[3][24]/NET0131  & n2765 ;
  assign n3157 = \u4_mem_reg[1][24]/NET0131  & n2903 ;
  assign n3160 = ~n3156 & ~n3157 ;
  assign n3161 = ~n3158 & n3160 ;
  assign n3162 = n3159 & n3161 ;
  assign n3154 = ~\u4_rp_reg[0]/P0001  & n3106 ;
  assign n3163 = n2760 & ~n3154 ;
  assign n3164 = ~n3162 & n3163 ;
  assign n3173 = ~n3097 & n3099 ;
  assign n3165 = \u4_mem_reg[3][12]/NET0131  & n2765 ;
  assign n3166 = \u4_mem_reg[2][12]/NET0131  & n2901 ;
  assign n3169 = ~n3165 & ~n3166 ;
  assign n3167 = \u4_mem_reg[0][12]/NET0131  & n2905 ;
  assign n3168 = \u4_mem_reg[1][12]/NET0131  & n2903 ;
  assign n3170 = ~n3167 & ~n3168 ;
  assign n3171 = n3169 & n3170 ;
  assign n3172 = n2910 & ~n3171 ;
  assign n3174 = n2759 & ~n3172 ;
  assign n3175 = ~n3173 & n3174 ;
  assign n3176 = ~n3164 & n3175 ;
  assign n3153 = ~\u4_dout_reg[12]/P0001  & ~n2759 ;
  assign n3177 = \u13_occ0_r_reg[8]/NET0131  & ~n3153 ;
  assign n3178 = ~n3176 & n3177 ;
  assign n3181 = \u4_mem_reg[2][25]/NET0131  & n2901 ;
  assign n3185 = \u4_rp_reg[0]/P0001  & ~n3181 ;
  assign n3184 = \u4_mem_reg[0][25]/NET0131  & n2905 ;
  assign n3182 = \u4_mem_reg[3][25]/NET0131  & n2765 ;
  assign n3183 = \u4_mem_reg[1][25]/NET0131  & n2903 ;
  assign n3186 = ~n3182 & ~n3183 ;
  assign n3187 = ~n3184 & n3186 ;
  assign n3188 = n3185 & n3187 ;
  assign n3180 = ~\u4_rp_reg[0]/P0001  & n3146 ;
  assign n3189 = n2760 & ~n3180 ;
  assign n3190 = ~n3188 & n3189 ;
  assign n3199 = n3099 & ~n3138 ;
  assign n3191 = \u4_mem_reg[1][13]/NET0131  & n2903 ;
  assign n3192 = \u4_mem_reg[3][13]/NET0131  & n2765 ;
  assign n3195 = ~n3191 & ~n3192 ;
  assign n3193 = \u4_mem_reg[2][13]/NET0131  & n2901 ;
  assign n3194 = \u4_mem_reg[0][13]/NET0131  & n2905 ;
  assign n3196 = ~n3193 & ~n3194 ;
  assign n3197 = n3195 & n3196 ;
  assign n3198 = n2910 & ~n3197 ;
  assign n3200 = n2759 & ~n3198 ;
  assign n3201 = ~n3199 & n3200 ;
  assign n3202 = ~n3190 & n3201 ;
  assign n3179 = ~\u4_dout_reg[13]/P0001  & ~n2759 ;
  assign n3203 = \u13_occ0_r_reg[8]/NET0131  & ~n3179 ;
  assign n3204 = ~n3202 & n3203 ;
  assign n3207 = \u4_mem_reg[2][26]/NET0131  & n2901 ;
  assign n3211 = \u4_rp_reg[0]/P0001  & ~n3207 ;
  assign n3210 = \u4_mem_reg[0][26]/NET0131  & n2905 ;
  assign n3208 = \u4_mem_reg[3][26]/NET0131  & n2765 ;
  assign n3209 = \u4_mem_reg[1][26]/NET0131  & n2903 ;
  assign n3212 = ~n3208 & ~n3209 ;
  assign n3213 = ~n3210 & n3212 ;
  assign n3214 = n3211 & n3213 ;
  assign n3206 = ~\u4_rp_reg[0]/P0001  & n3097 ;
  assign n3215 = n2760 & ~n3206 ;
  assign n3216 = ~n3214 & n3215 ;
  assign n3225 = n3099 & ~n3171 ;
  assign n3217 = \u4_mem_reg[1][14]/NET0131  & n2903 ;
  assign n3218 = \u4_mem_reg[2][14]/NET0131  & n2901 ;
  assign n3221 = ~n3217 & ~n3218 ;
  assign n3219 = \u4_mem_reg[0][14]/NET0131  & n2905 ;
  assign n3220 = \u4_mem_reg[3][14]/NET0131  & n2765 ;
  assign n3222 = ~n3219 & ~n3220 ;
  assign n3223 = n3221 & n3222 ;
  assign n3224 = n2910 & ~n3223 ;
  assign n3226 = n2759 & ~n3224 ;
  assign n3227 = ~n3225 & n3226 ;
  assign n3228 = ~n3216 & n3227 ;
  assign n3205 = ~\u4_dout_reg[14]/P0001  & ~n2759 ;
  assign n3229 = \u13_occ0_r_reg[8]/NET0131  & ~n3205 ;
  assign n3230 = ~n3228 & n3229 ;
  assign n3233 = \u4_mem_reg[2][27]/NET0131  & n2901 ;
  assign n3237 = \u4_rp_reg[0]/P0001  & ~n3233 ;
  assign n3236 = \u4_mem_reg[0][27]/NET0131  & n2905 ;
  assign n3234 = \u4_mem_reg[1][27]/NET0131  & n2903 ;
  assign n3235 = \u4_mem_reg[3][27]/NET0131  & n2765 ;
  assign n3238 = ~n3234 & ~n3235 ;
  assign n3239 = ~n3236 & n3238 ;
  assign n3240 = n3237 & n3239 ;
  assign n3232 = ~\u4_rp_reg[0]/P0001  & n3138 ;
  assign n3241 = n2760 & ~n3232 ;
  assign n3242 = ~n3240 & n3241 ;
  assign n3251 = n3099 & ~n3197 ;
  assign n3243 = \u4_mem_reg[2][15]/NET0131  & n2901 ;
  assign n3244 = \u4_mem_reg[0][15]/NET0131  & n2905 ;
  assign n3247 = ~n3243 & ~n3244 ;
  assign n3245 = \u4_mem_reg[1][15]/NET0131  & n2903 ;
  assign n3246 = \u4_mem_reg[3][15]/NET0131  & n2765 ;
  assign n3248 = ~n3245 & ~n3246 ;
  assign n3249 = n3247 & n3248 ;
  assign n3250 = n2910 & ~n3249 ;
  assign n3252 = n2759 & ~n3250 ;
  assign n3253 = ~n3251 & n3252 ;
  assign n3254 = ~n3242 & n3253 ;
  assign n3231 = ~\u4_dout_reg[15]/P0001  & ~n2759 ;
  assign n3255 = \u13_occ0_r_reg[8]/NET0131  & ~n3231 ;
  assign n3256 = ~n3254 & n3255 ;
  assign n3259 = \u4_mem_reg[2][28]/NET0131  & n2901 ;
  assign n3263 = \u4_rp_reg[0]/P0001  & ~n3259 ;
  assign n3262 = \u4_mem_reg[0][28]/NET0131  & n2905 ;
  assign n3260 = \u4_mem_reg[1][28]/NET0131  & n2903 ;
  assign n3261 = \u4_mem_reg[3][28]/NET0131  & n2765 ;
  assign n3264 = ~n3260 & ~n3261 ;
  assign n3265 = ~n3262 & n3264 ;
  assign n3266 = n3263 & n3265 ;
  assign n3258 = ~\u4_rp_reg[0]/P0001  & n3171 ;
  assign n3267 = n2760 & ~n3258 ;
  assign n3268 = ~n3266 & n3267 ;
  assign n3277 = n3099 & ~n3223 ;
  assign n3269 = \u4_mem_reg[3][16]/NET0131  & n2765 ;
  assign n3270 = \u4_mem_reg[2][16]/NET0131  & n2901 ;
  assign n3273 = ~n3269 & ~n3270 ;
  assign n3271 = \u4_mem_reg[0][16]/NET0131  & n2905 ;
  assign n3272 = \u4_mem_reg[1][16]/NET0131  & n2903 ;
  assign n3274 = ~n3271 & ~n3272 ;
  assign n3275 = n3273 & n3274 ;
  assign n3276 = n2910 & ~n3275 ;
  assign n3278 = n2759 & ~n3276 ;
  assign n3279 = ~n3277 & n3278 ;
  assign n3280 = ~n3268 & n3279 ;
  assign n3257 = ~\u4_dout_reg[16]/P0001  & ~n2759 ;
  assign n3281 = \u13_occ0_r_reg[8]/NET0131  & ~n3257 ;
  assign n3282 = ~n3280 & n3281 ;
  assign n3285 = \u4_mem_reg[2][29]/NET0131  & n2901 ;
  assign n3289 = \u4_rp_reg[0]/P0001  & ~n3285 ;
  assign n3288 = \u4_mem_reg[0][29]/NET0131  & n2905 ;
  assign n3286 = \u4_mem_reg[3][29]/NET0131  & n2765 ;
  assign n3287 = \u4_mem_reg[1][29]/NET0131  & n2903 ;
  assign n3290 = ~n3286 & ~n3287 ;
  assign n3291 = ~n3288 & n3290 ;
  assign n3292 = n3289 & n3291 ;
  assign n3284 = ~\u4_rp_reg[0]/P0001  & n3197 ;
  assign n3293 = n2760 & ~n3284 ;
  assign n3294 = ~n3292 & n3293 ;
  assign n3303 = n3099 & ~n3249 ;
  assign n3295 = \u4_mem_reg[3][17]/NET0131  & n2765 ;
  assign n3296 = \u4_mem_reg[2][17]/NET0131  & n2901 ;
  assign n3299 = ~n3295 & ~n3296 ;
  assign n3297 = \u4_mem_reg[1][17]/NET0131  & n2903 ;
  assign n3298 = \u4_mem_reg[0][17]/NET0131  & n2905 ;
  assign n3300 = ~n3297 & ~n3298 ;
  assign n3301 = n3299 & n3300 ;
  assign n3302 = n2910 & ~n3301 ;
  assign n3304 = n2759 & ~n3302 ;
  assign n3305 = ~n3303 & n3304 ;
  assign n3306 = ~n3294 & n3305 ;
  assign n3283 = ~\u4_dout_reg[17]/P0001  & ~n2759 ;
  assign n3307 = \u13_occ0_r_reg[8]/NET0131  & ~n3283 ;
  assign n3308 = ~n3306 & n3307 ;
  assign n3309 = \in_valid_s_reg[0]/NET0131  & \u14_u6_en_out_l_reg/NET0131  ;
  assign n3310 = ~\u14_u6_en_out_l2_reg/P0001  & n3309 ;
  assign n3311 = ~\u13_icc_r_reg[2]/NET0131  & ~\u13_icc_r_reg[3]/NET0131  ;
  assign n3312 = ~\u9_wp_reg[0]/NET0131  & n3311 ;
  assign n3313 = n3310 & ~n3312 ;
  assign n3314 = \u9_wp_reg[1]/P0001  & n3313 ;
  assign n3316 = ~\u9_wp_reg[2]/P0001  & ~n3314 ;
  assign n3315 = \u9_wp_reg[2]/P0001  & n3314 ;
  assign n3317 = \u13_icc_r_reg[0]/NET0131  & ~n3315 ;
  assign n3318 = ~n3316 & n3317 ;
  assign n3321 = \u4_mem_reg[2][30]/NET0131  & n2901 ;
  assign n3325 = \u4_rp_reg[0]/P0001  & ~n3321 ;
  assign n3324 = \u4_mem_reg[0][30]/NET0131  & n2905 ;
  assign n3322 = \u4_mem_reg[3][30]/NET0131  & n2765 ;
  assign n3323 = \u4_mem_reg[1][30]/NET0131  & n2903 ;
  assign n3326 = ~n3322 & ~n3323 ;
  assign n3327 = ~n3324 & n3326 ;
  assign n3328 = n3325 & n3327 ;
  assign n3320 = ~\u4_rp_reg[0]/P0001  & n3223 ;
  assign n3329 = n2760 & ~n3320 ;
  assign n3330 = ~n3328 & n3329 ;
  assign n3339 = n3099 & ~n3275 ;
  assign n3331 = \u4_mem_reg[1][18]/NET0131  & n2903 ;
  assign n3332 = \u4_mem_reg[3][18]/NET0131  & n2765 ;
  assign n3335 = ~n3331 & ~n3332 ;
  assign n3333 = \u4_mem_reg[2][18]/NET0131  & n2901 ;
  assign n3334 = \u4_mem_reg[0][18]/NET0131  & n2905 ;
  assign n3336 = ~n3333 & ~n3334 ;
  assign n3337 = n3335 & n3336 ;
  assign n3338 = n2910 & ~n3337 ;
  assign n3340 = n2759 & ~n3338 ;
  assign n3341 = ~n3339 & n3340 ;
  assign n3342 = ~n3330 & n3341 ;
  assign n3319 = ~\u4_dout_reg[18]/P0001  & ~n2759 ;
  assign n3343 = \u13_occ0_r_reg[8]/NET0131  & ~n3319 ;
  assign n3344 = ~n3342 & n3343 ;
  assign n3347 = \u4_mem_reg[2][31]/NET0131  & n2901 ;
  assign n3351 = \u4_rp_reg[0]/P0001  & ~n3347 ;
  assign n3350 = \u4_mem_reg[0][31]/NET0131  & n2905 ;
  assign n3348 = \u4_mem_reg[3][31]/NET0131  & n2765 ;
  assign n3349 = \u4_mem_reg[1][31]/NET0131  & n2903 ;
  assign n3352 = ~n3348 & ~n3349 ;
  assign n3353 = ~n3350 & n3352 ;
  assign n3354 = n3351 & n3353 ;
  assign n3346 = ~\u4_rp_reg[0]/P0001  & n3249 ;
  assign n3355 = n2760 & ~n3346 ;
  assign n3356 = ~n3354 & n3355 ;
  assign n3365 = n3099 & ~n3301 ;
  assign n3357 = \u4_mem_reg[3][19]/NET0131  & n2765 ;
  assign n3358 = \u4_mem_reg[2][19]/NET0131  & n2901 ;
  assign n3361 = ~n3357 & ~n3358 ;
  assign n3359 = \u4_mem_reg[1][19]/NET0131  & n2903 ;
  assign n3360 = \u4_mem_reg[0][19]/NET0131  & n2905 ;
  assign n3362 = ~n3359 & ~n3360 ;
  assign n3363 = n3361 & n3362 ;
  assign n3364 = n2910 & ~n3363 ;
  assign n3366 = n2759 & ~n3364 ;
  assign n3367 = ~n3365 & n3366 ;
  assign n3368 = ~n3356 & n3367 ;
  assign n3345 = ~\u4_dout_reg[19]/P0001  & ~n2759 ;
  assign n3369 = \u13_occ0_r_reg[8]/NET0131  & ~n3345 ;
  assign n3370 = ~n3368 & n3369 ;
  assign n3373 = \u4_mem_reg[1][2]/NET0131  & n2903 ;
  assign n3374 = \u4_mem_reg[0][2]/NET0131  & n2905 ;
  assign n3377 = ~n3373 & ~n3374 ;
  assign n3375 = \u4_mem_reg[2][2]/NET0131  & n2901 ;
  assign n3376 = \u4_mem_reg[3][2]/NET0131  & n2765 ;
  assign n3378 = ~n3375 & ~n3376 ;
  assign n3379 = n3377 & n3378 ;
  assign n3380 = n2910 & ~n3379 ;
  assign n3372 = ~n2909 & n3099 ;
  assign n3381 = n2759 & ~n3372 ;
  assign n3382 = ~n3380 & n3381 ;
  assign n3371 = ~\u4_dout_reg[2]/P0001  & ~n2759 ;
  assign n3383 = \u13_occ0_r_reg[8]/NET0131  & ~n3371 ;
  assign n3384 = ~n3382 & n3383 ;
  assign n3394 = ~n2922 & n3099 ;
  assign n3386 = \u4_mem_reg[2][3]/NET0131  & n2901 ;
  assign n3387 = \u4_mem_reg[3][3]/NET0131  & n2765 ;
  assign n3390 = ~n3386 & ~n3387 ;
  assign n3388 = \u4_mem_reg[1][3]/NET0131  & n2903 ;
  assign n3389 = \u4_mem_reg[0][3]/NET0131  & n2905 ;
  assign n3391 = ~n3388 & ~n3389 ;
  assign n3392 = n3390 & n3391 ;
  assign n3393 = n2910 & ~n3392 ;
  assign n3395 = n2759 & ~n3393 ;
  assign n3396 = ~n3394 & n3395 ;
  assign n3385 = ~\u4_dout_reg[3]/P0001  & ~n2759 ;
  assign n3397 = \u13_occ0_r_reg[8]/NET0131  & ~n3385 ;
  assign n3398 = ~n3396 & n3397 ;
  assign n3401 = \u4_rp_reg[0]/P0001  & n3275 ;
  assign n3400 = ~\u4_rp_reg[0]/P0001  & n2909 ;
  assign n3402 = n2760 & ~n3400 ;
  assign n3403 = ~n3401 & n3402 ;
  assign n3412 = n3099 & ~n3379 ;
  assign n3404 = \u4_mem_reg[3][4]/NET0131  & n2765 ;
  assign n3405 = \u4_mem_reg[2][4]/NET0131  & n2901 ;
  assign n3408 = ~n3404 & ~n3405 ;
  assign n3406 = \u4_mem_reg[0][4]/NET0131  & n2905 ;
  assign n3407 = \u4_mem_reg[1][4]/NET0131  & n2903 ;
  assign n3409 = ~n3406 & ~n3407 ;
  assign n3410 = n3408 & n3409 ;
  assign n3411 = n2910 & ~n3410 ;
  assign n3413 = n2759 & ~n3411 ;
  assign n3414 = ~n3412 & n3413 ;
  assign n3415 = ~n3403 & n3414 ;
  assign n3399 = ~\u4_dout_reg[4]/P0001  & ~n2759 ;
  assign n3416 = \u13_occ0_r_reg[8]/NET0131  & ~n3399 ;
  assign n3417 = ~n3415 & n3416 ;
  assign n3420 = \u4_rp_reg[0]/P0001  & n3301 ;
  assign n3419 = ~\u4_rp_reg[0]/P0001  & n2922 ;
  assign n3421 = n2760 & ~n3419 ;
  assign n3422 = ~n3420 & n3421 ;
  assign n3431 = n3099 & ~n3392 ;
  assign n3423 = \u4_mem_reg[2][5]/NET0131  & n2901 ;
  assign n3424 = \u4_mem_reg[1][5]/NET0131  & n2903 ;
  assign n3427 = ~n3423 & ~n3424 ;
  assign n3425 = \u4_mem_reg[3][5]/NET0131  & n2765 ;
  assign n3426 = \u4_mem_reg[0][5]/NET0131  & n2905 ;
  assign n3428 = ~n3425 & ~n3426 ;
  assign n3429 = n3427 & n3428 ;
  assign n3430 = n2910 & ~n3429 ;
  assign n3432 = n2759 & ~n3430 ;
  assign n3433 = ~n3431 & n3432 ;
  assign n3434 = ~n3422 & n3433 ;
  assign n3418 = ~\u4_dout_reg[5]/P0001  & ~n2759 ;
  assign n3435 = \u13_occ0_r_reg[8]/NET0131  & ~n3418 ;
  assign n3436 = ~n3434 & n3435 ;
  assign n3439 = \u4_rp_reg[0]/P0001  & n3337 ;
  assign n3438 = ~\u4_rp_reg[0]/P0001  & n3379 ;
  assign n3440 = n2760 & ~n3438 ;
  assign n3441 = ~n3439 & n3440 ;
  assign n3443 = n3099 & ~n3410 ;
  assign n3442 = n2910 & ~n3079 ;
  assign n3444 = n2759 & ~n3442 ;
  assign n3445 = ~n3443 & n3444 ;
  assign n3446 = ~n3441 & n3445 ;
  assign n3437 = ~\u4_dout_reg[6]/P0001  & ~n2759 ;
  assign n3447 = \u13_occ0_r_reg[8]/NET0131  & ~n3437 ;
  assign n3448 = ~n3446 & n3447 ;
  assign n3451 = \u4_rp_reg[0]/P0001  & n3363 ;
  assign n3450 = ~\u4_rp_reg[0]/P0001  & n3392 ;
  assign n3452 = n2760 & ~n3450 ;
  assign n3453 = ~n3451 & n3452 ;
  assign n3455 = n3099 & ~n3429 ;
  assign n3454 = n2910 & ~n3120 ;
  assign n3456 = n2759 & ~n3454 ;
  assign n3457 = ~n3455 & n3456 ;
  assign n3458 = ~n3453 & n3457 ;
  assign n3449 = ~\u4_dout_reg[7]/P0001  & ~n2759 ;
  assign n3459 = \u13_occ0_r_reg[8]/NET0131  & ~n3449 ;
  assign n3460 = ~n3458 & n3459 ;
  assign n3463 = \u4_mem_reg[2][20]/NET0131  & n2901 ;
  assign n3467 = \u4_rp_reg[0]/P0001  & ~n3463 ;
  assign n3466 = \u4_mem_reg[0][20]/NET0131  & n2905 ;
  assign n3464 = \u4_mem_reg[3][20]/NET0131  & n2765 ;
  assign n3465 = \u4_mem_reg[1][20]/NET0131  & n2903 ;
  assign n3468 = ~n3464 & ~n3465 ;
  assign n3469 = ~n3466 & n3468 ;
  assign n3470 = n3467 & n3469 ;
  assign n3462 = ~\u4_rp_reg[0]/P0001  & n3410 ;
  assign n3471 = n2760 & ~n3462 ;
  assign n3472 = ~n3470 & n3471 ;
  assign n3474 = ~n3079 & n3099 ;
  assign n3473 = n2910 & ~n3106 ;
  assign n3475 = n2759 & ~n3473 ;
  assign n3476 = ~n3474 & n3475 ;
  assign n3477 = ~n3472 & n3476 ;
  assign n3461 = ~\u4_dout_reg[8]/P0001  & ~n2759 ;
  assign n3478 = \u13_occ0_r_reg[8]/NET0131  & ~n3461 ;
  assign n3479 = ~n3477 & n3478 ;
  assign n3482 = \u4_mem_reg[2][21]/NET0131  & n2901 ;
  assign n3486 = \u4_rp_reg[0]/P0001  & ~n3482 ;
  assign n3485 = \u4_mem_reg[0][21]/NET0131  & n2905 ;
  assign n3483 = \u4_mem_reg[3][21]/NET0131  & n2765 ;
  assign n3484 = \u4_mem_reg[1][21]/NET0131  & n2903 ;
  assign n3487 = ~n3483 & ~n3484 ;
  assign n3488 = ~n3485 & n3487 ;
  assign n3489 = n3486 & n3488 ;
  assign n3481 = ~\u4_rp_reg[0]/P0001  & n3429 ;
  assign n3490 = n2760 & ~n3481 ;
  assign n3491 = ~n3489 & n3490 ;
  assign n3493 = n3099 & ~n3120 ;
  assign n3492 = n2910 & ~n3146 ;
  assign n3494 = n2759 & ~n3492 ;
  assign n3495 = ~n3493 & n3494 ;
  assign n3496 = ~n3491 & n3495 ;
  assign n3480 = ~\u4_dout_reg[9]/P0001  & ~n2759 ;
  assign n3497 = \u13_occ0_r_reg[8]/NET0131  & ~n3480 ;
  assign n3498 = ~n3496 & n3497 ;
  assign n3499 = \in_valid_s_reg[1]/NET0131  & \u14_u7_en_out_l_reg/NET0131  ;
  assign n3500 = ~\u14_u7_en_out_l2_reg/P0001  & n3499 ;
  assign n3501 = ~\u13_icc_r_reg[10]/NET0131  & ~\u13_icc_r_reg[11]/NET0131  ;
  assign n3502 = ~\u10_wp_reg[0]/NET0131  & n3501 ;
  assign n3503 = n3500 & ~n3502 ;
  assign n3504 = \u10_wp_reg[1]/P0001  & n3503 ;
  assign n3506 = ~\u10_wp_reg[2]/P0001  & ~n3504 ;
  assign n3505 = \u10_wp_reg[2]/P0001  & n3504 ;
  assign n3507 = \u13_icc_r_reg[8]/NET0131  & ~n3505 ;
  assign n3508 = ~n3506 & n3507 ;
  assign n3518 = \u5_mem_reg[2][22]/NET0131  & n2930 ;
  assign n3522 = \u5_rp_reg[0]/P0001  & ~n3518 ;
  assign n3521 = \u5_mem_reg[0][22]/NET0131  & n2932 ;
  assign n3519 = \u5_mem_reg[3][22]/NET0131  & n2776 ;
  assign n3520 = \u5_mem_reg[1][22]/NET0131  & n2928 ;
  assign n3523 = ~n3519 & ~n3520 ;
  assign n3524 = ~n3521 & n3523 ;
  assign n3525 = n3522 & n3524 ;
  assign n3510 = \u5_mem_reg[1][6]/NET0131  & n2928 ;
  assign n3511 = \u5_mem_reg[2][6]/NET0131  & n2930 ;
  assign n3514 = ~n3510 & ~n3511 ;
  assign n3512 = \u5_mem_reg[3][6]/NET0131  & n2776 ;
  assign n3513 = \u5_mem_reg[0][6]/NET0131  & n2932 ;
  assign n3515 = ~n3512 & ~n3513 ;
  assign n3516 = n3514 & n3515 ;
  assign n3517 = ~\u5_rp_reg[0]/P0001  & n3516 ;
  assign n3526 = n2771 & ~n3517 ;
  assign n3527 = ~n3525 & n3526 ;
  assign n3536 = \u13_occ0_r_reg[18]/NET0131  & ~\u13_occ0_r_reg[19]/NET0131  ;
  assign n3537 = \u5_mem_reg[2][8]/NET0131  & n2930 ;
  assign n3538 = \u5_mem_reg[1][8]/NET0131  & n2928 ;
  assign n3541 = ~n3537 & ~n3538 ;
  assign n3539 = \u5_mem_reg[3][8]/NET0131  & n2776 ;
  assign n3540 = \u5_mem_reg[0][8]/NET0131  & n2932 ;
  assign n3542 = ~n3539 & ~n3540 ;
  assign n3543 = n3541 & n3542 ;
  assign n3544 = n3536 & ~n3543 ;
  assign n3528 = \u5_mem_reg[2][10]/NET0131  & n2930 ;
  assign n3529 = \u5_mem_reg[1][10]/NET0131  & n2928 ;
  assign n3532 = ~n3528 & ~n3529 ;
  assign n3530 = \u5_mem_reg[3][10]/NET0131  & n2776 ;
  assign n3531 = \u5_mem_reg[0][10]/NET0131  & n2932 ;
  assign n3533 = ~n3530 & ~n3531 ;
  assign n3534 = n3532 & n3533 ;
  assign n3535 = n2937 & ~n3534 ;
  assign n3545 = n2770 & ~n3535 ;
  assign n3546 = ~n3544 & n3545 ;
  assign n3547 = ~n3527 & n3546 ;
  assign n3509 = ~\u5_dout_reg[10]/P0001  & ~n2770 ;
  assign n3548 = \u13_occ0_r_reg[16]/NET0131  & ~n3509 ;
  assign n3549 = ~n3547 & n3548 ;
  assign n3559 = \u5_mem_reg[2][23]/NET0131  & n2930 ;
  assign n3563 = \u5_rp_reg[0]/P0001  & ~n3559 ;
  assign n3562 = \u5_mem_reg[0][23]/NET0131  & n2932 ;
  assign n3560 = \u5_mem_reg[3][23]/NET0131  & n2776 ;
  assign n3561 = \u5_mem_reg[1][23]/NET0131  & n2928 ;
  assign n3564 = ~n3560 & ~n3561 ;
  assign n3565 = ~n3562 & n3564 ;
  assign n3566 = n3563 & n3565 ;
  assign n3551 = \u5_mem_reg[2][7]/NET0131  & n2930 ;
  assign n3552 = \u5_mem_reg[1][7]/NET0131  & n2928 ;
  assign n3555 = ~n3551 & ~n3552 ;
  assign n3553 = \u5_mem_reg[3][7]/NET0131  & n2776 ;
  assign n3554 = \u5_mem_reg[0][7]/NET0131  & n2932 ;
  assign n3556 = ~n3553 & ~n3554 ;
  assign n3557 = n3555 & n3556 ;
  assign n3558 = ~\u5_rp_reg[0]/P0001  & n3557 ;
  assign n3567 = n2771 & ~n3558 ;
  assign n3568 = ~n3566 & n3567 ;
  assign n3577 = \u5_mem_reg[1][9]/NET0131  & n2928 ;
  assign n3578 = \u5_mem_reg[2][9]/NET0131  & n2930 ;
  assign n3581 = ~n3577 & ~n3578 ;
  assign n3579 = \u5_mem_reg[3][9]/NET0131  & n2776 ;
  assign n3580 = \u5_mem_reg[0][9]/NET0131  & n2932 ;
  assign n3582 = ~n3579 & ~n3580 ;
  assign n3583 = n3581 & n3582 ;
  assign n3584 = n3536 & ~n3583 ;
  assign n3569 = \u5_mem_reg[2][11]/NET0131  & n2930 ;
  assign n3570 = \u5_mem_reg[1][11]/NET0131  & n2928 ;
  assign n3573 = ~n3569 & ~n3570 ;
  assign n3571 = \u5_mem_reg[3][11]/NET0131  & n2776 ;
  assign n3572 = \u5_mem_reg[0][11]/NET0131  & n2932 ;
  assign n3574 = ~n3571 & ~n3572 ;
  assign n3575 = n3573 & n3574 ;
  assign n3576 = n2937 & ~n3575 ;
  assign n3585 = n2770 & ~n3576 ;
  assign n3586 = ~n3584 & n3585 ;
  assign n3587 = ~n3568 & n3586 ;
  assign n3550 = ~\u5_dout_reg[11]/P0001  & ~n2770 ;
  assign n3588 = \u13_occ0_r_reg[16]/NET0131  & ~n3550 ;
  assign n3589 = ~n3587 & n3588 ;
  assign n3592 = \u5_mem_reg[2][24]/NET0131  & n2930 ;
  assign n3596 = \u5_rp_reg[0]/P0001  & ~n3592 ;
  assign n3595 = \u5_mem_reg[0][24]/NET0131  & n2932 ;
  assign n3593 = \u5_mem_reg[3][24]/NET0131  & n2776 ;
  assign n3594 = \u5_mem_reg[1][24]/NET0131  & n2928 ;
  assign n3597 = ~n3593 & ~n3594 ;
  assign n3598 = ~n3595 & n3597 ;
  assign n3599 = n3596 & n3598 ;
  assign n3591 = ~\u5_rp_reg[0]/P0001  & n3543 ;
  assign n3600 = n2771 & ~n3591 ;
  assign n3601 = ~n3599 & n3600 ;
  assign n3610 = ~n3534 & n3536 ;
  assign n3602 = \u5_mem_reg[1][12]/NET0131  & n2928 ;
  assign n3603 = \u5_mem_reg[2][12]/NET0131  & n2930 ;
  assign n3606 = ~n3602 & ~n3603 ;
  assign n3604 = \u5_mem_reg[3][12]/NET0131  & n2776 ;
  assign n3605 = \u5_mem_reg[0][12]/NET0131  & n2932 ;
  assign n3607 = ~n3604 & ~n3605 ;
  assign n3608 = n3606 & n3607 ;
  assign n3609 = n2937 & ~n3608 ;
  assign n3611 = n2770 & ~n3609 ;
  assign n3612 = ~n3610 & n3611 ;
  assign n3613 = ~n3601 & n3612 ;
  assign n3590 = ~\u5_dout_reg[12]/P0001  & ~n2770 ;
  assign n3614 = \u13_occ0_r_reg[16]/NET0131  & ~n3590 ;
  assign n3615 = ~n3613 & n3614 ;
  assign n3618 = \u5_mem_reg[2][25]/NET0131  & n2930 ;
  assign n3622 = \u5_rp_reg[0]/P0001  & ~n3618 ;
  assign n3621 = \u5_mem_reg[0][25]/NET0131  & n2932 ;
  assign n3619 = \u5_mem_reg[3][25]/NET0131  & n2776 ;
  assign n3620 = \u5_mem_reg[1][25]/NET0131  & n2928 ;
  assign n3623 = ~n3619 & ~n3620 ;
  assign n3624 = ~n3621 & n3623 ;
  assign n3625 = n3622 & n3624 ;
  assign n3617 = ~\u5_rp_reg[0]/P0001  & n3583 ;
  assign n3626 = n2771 & ~n3617 ;
  assign n3627 = ~n3625 & n3626 ;
  assign n3636 = n3536 & ~n3575 ;
  assign n3628 = \u5_mem_reg[1][13]/NET0131  & n2928 ;
  assign n3629 = \u5_mem_reg[2][13]/NET0131  & n2930 ;
  assign n3632 = ~n3628 & ~n3629 ;
  assign n3630 = \u5_mem_reg[3][13]/NET0131  & n2776 ;
  assign n3631 = \u5_mem_reg[0][13]/NET0131  & n2932 ;
  assign n3633 = ~n3630 & ~n3631 ;
  assign n3634 = n3632 & n3633 ;
  assign n3635 = n2937 & ~n3634 ;
  assign n3637 = n2770 & ~n3635 ;
  assign n3638 = ~n3636 & n3637 ;
  assign n3639 = ~n3627 & n3638 ;
  assign n3616 = ~\u5_dout_reg[13]/P0001  & ~n2770 ;
  assign n3640 = \u13_occ0_r_reg[16]/NET0131  & ~n3616 ;
  assign n3641 = ~n3639 & n3640 ;
  assign n3644 = \u5_mem_reg[2][26]/NET0131  & n2930 ;
  assign n3648 = \u5_rp_reg[0]/P0001  & ~n3644 ;
  assign n3647 = \u5_mem_reg[0][26]/NET0131  & n2932 ;
  assign n3645 = \u5_mem_reg[3][26]/NET0131  & n2776 ;
  assign n3646 = \u5_mem_reg[1][26]/NET0131  & n2928 ;
  assign n3649 = ~n3645 & ~n3646 ;
  assign n3650 = ~n3647 & n3649 ;
  assign n3651 = n3648 & n3650 ;
  assign n3643 = ~\u5_rp_reg[0]/P0001  & n3534 ;
  assign n3652 = n2771 & ~n3643 ;
  assign n3653 = ~n3651 & n3652 ;
  assign n3662 = n3536 & ~n3608 ;
  assign n3654 = \u5_mem_reg[2][14]/NET0131  & n2930 ;
  assign n3655 = \u5_mem_reg[3][14]/NET0131  & n2776 ;
  assign n3658 = ~n3654 & ~n3655 ;
  assign n3656 = \u5_mem_reg[0][14]/NET0131  & n2932 ;
  assign n3657 = \u5_mem_reg[1][14]/NET0131  & n2928 ;
  assign n3659 = ~n3656 & ~n3657 ;
  assign n3660 = n3658 & n3659 ;
  assign n3661 = n2937 & ~n3660 ;
  assign n3663 = n2770 & ~n3661 ;
  assign n3664 = ~n3662 & n3663 ;
  assign n3665 = ~n3653 & n3664 ;
  assign n3642 = ~\u5_dout_reg[14]/P0001  & ~n2770 ;
  assign n3666 = \u13_occ0_r_reg[16]/NET0131  & ~n3642 ;
  assign n3667 = ~n3665 & n3666 ;
  assign n3670 = \u5_mem_reg[2][27]/NET0131  & n2930 ;
  assign n3674 = \u5_rp_reg[0]/P0001  & ~n3670 ;
  assign n3673 = \u5_mem_reg[0][27]/NET0131  & n2932 ;
  assign n3671 = \u5_mem_reg[3][27]/NET0131  & n2776 ;
  assign n3672 = \u5_mem_reg[1][27]/NET0131  & n2928 ;
  assign n3675 = ~n3671 & ~n3672 ;
  assign n3676 = ~n3673 & n3675 ;
  assign n3677 = n3674 & n3676 ;
  assign n3669 = ~\u5_rp_reg[0]/P0001  & n3575 ;
  assign n3678 = n2771 & ~n3669 ;
  assign n3679 = ~n3677 & n3678 ;
  assign n3688 = n3536 & ~n3634 ;
  assign n3680 = \u5_mem_reg[1][15]/NET0131  & n2928 ;
  assign n3681 = \u5_mem_reg[3][15]/NET0131  & n2776 ;
  assign n3684 = ~n3680 & ~n3681 ;
  assign n3682 = \u5_mem_reg[2][15]/NET0131  & n2930 ;
  assign n3683 = \u5_mem_reg[0][15]/NET0131  & n2932 ;
  assign n3685 = ~n3682 & ~n3683 ;
  assign n3686 = n3684 & n3685 ;
  assign n3687 = n2937 & ~n3686 ;
  assign n3689 = n2770 & ~n3687 ;
  assign n3690 = ~n3688 & n3689 ;
  assign n3691 = ~n3679 & n3690 ;
  assign n3668 = ~\u5_dout_reg[15]/P0001  & ~n2770 ;
  assign n3692 = \u13_occ0_r_reg[16]/NET0131  & ~n3668 ;
  assign n3693 = ~n3691 & n3692 ;
  assign n3696 = \u5_mem_reg[2][28]/NET0131  & n2930 ;
  assign n3700 = \u5_rp_reg[0]/P0001  & ~n3696 ;
  assign n3699 = \u5_mem_reg[0][28]/NET0131  & n2932 ;
  assign n3697 = \u5_mem_reg[3][28]/NET0131  & n2776 ;
  assign n3698 = \u5_mem_reg[1][28]/NET0131  & n2928 ;
  assign n3701 = ~n3697 & ~n3698 ;
  assign n3702 = ~n3699 & n3701 ;
  assign n3703 = n3700 & n3702 ;
  assign n3695 = ~\u5_rp_reg[0]/P0001  & n3608 ;
  assign n3704 = n2771 & ~n3695 ;
  assign n3705 = ~n3703 & n3704 ;
  assign n3714 = n3536 & ~n3660 ;
  assign n3706 = \u5_mem_reg[1][16]/NET0131  & n2928 ;
  assign n3707 = \u5_mem_reg[3][16]/NET0131  & n2776 ;
  assign n3710 = ~n3706 & ~n3707 ;
  assign n3708 = \u5_mem_reg[2][16]/NET0131  & n2930 ;
  assign n3709 = \u5_mem_reg[0][16]/NET0131  & n2932 ;
  assign n3711 = ~n3708 & ~n3709 ;
  assign n3712 = n3710 & n3711 ;
  assign n3713 = n2937 & ~n3712 ;
  assign n3715 = n2770 & ~n3713 ;
  assign n3716 = ~n3714 & n3715 ;
  assign n3717 = ~n3705 & n3716 ;
  assign n3694 = ~\u5_dout_reg[16]/P0001  & ~n2770 ;
  assign n3718 = \u13_occ0_r_reg[16]/NET0131  & ~n3694 ;
  assign n3719 = ~n3717 & n3718 ;
  assign n3722 = \u5_mem_reg[2][29]/NET0131  & n2930 ;
  assign n3726 = \u5_rp_reg[0]/P0001  & ~n3722 ;
  assign n3725 = \u5_mem_reg[0][29]/NET0131  & n2932 ;
  assign n3723 = \u5_mem_reg[3][29]/NET0131  & n2776 ;
  assign n3724 = \u5_mem_reg[1][29]/NET0131  & n2928 ;
  assign n3727 = ~n3723 & ~n3724 ;
  assign n3728 = ~n3725 & n3727 ;
  assign n3729 = n3726 & n3728 ;
  assign n3721 = ~\u5_rp_reg[0]/P0001  & n3634 ;
  assign n3730 = n2771 & ~n3721 ;
  assign n3731 = ~n3729 & n3730 ;
  assign n3740 = n3536 & ~n3686 ;
  assign n3732 = \u5_mem_reg[2][17]/NET0131  & n2930 ;
  assign n3733 = \u5_mem_reg[3][17]/NET0131  & n2776 ;
  assign n3736 = ~n3732 & ~n3733 ;
  assign n3734 = \u5_mem_reg[1][17]/NET0131  & n2928 ;
  assign n3735 = \u5_mem_reg[0][17]/NET0131  & n2932 ;
  assign n3737 = ~n3734 & ~n3735 ;
  assign n3738 = n3736 & n3737 ;
  assign n3739 = n2937 & ~n3738 ;
  assign n3741 = n2770 & ~n3739 ;
  assign n3742 = ~n3740 & n3741 ;
  assign n3743 = ~n3731 & n3742 ;
  assign n3720 = ~\u5_dout_reg[17]/P0001  & ~n2770 ;
  assign n3744 = \u13_occ0_r_reg[16]/NET0131  & ~n3720 ;
  assign n3745 = ~n3743 & n3744 ;
  assign n3748 = \u5_mem_reg[2][30]/NET0131  & n2930 ;
  assign n3752 = \u5_rp_reg[0]/P0001  & ~n3748 ;
  assign n3751 = \u5_mem_reg[0][30]/NET0131  & n2932 ;
  assign n3749 = \u5_mem_reg[3][30]/NET0131  & n2776 ;
  assign n3750 = \u5_mem_reg[1][30]/NET0131  & n2928 ;
  assign n3753 = ~n3749 & ~n3750 ;
  assign n3754 = ~n3751 & n3753 ;
  assign n3755 = n3752 & n3754 ;
  assign n3747 = ~\u5_rp_reg[0]/P0001  & n3660 ;
  assign n3756 = n2771 & ~n3747 ;
  assign n3757 = ~n3755 & n3756 ;
  assign n3766 = n3536 & ~n3712 ;
  assign n3758 = \u5_mem_reg[1][18]/NET0131  & n2928 ;
  assign n3759 = \u5_mem_reg[2][18]/NET0131  & n2930 ;
  assign n3762 = ~n3758 & ~n3759 ;
  assign n3760 = \u5_mem_reg[3][18]/NET0131  & n2776 ;
  assign n3761 = \u5_mem_reg[0][18]/NET0131  & n2932 ;
  assign n3763 = ~n3760 & ~n3761 ;
  assign n3764 = n3762 & n3763 ;
  assign n3765 = n2937 & ~n3764 ;
  assign n3767 = n2770 & ~n3765 ;
  assign n3768 = ~n3766 & n3767 ;
  assign n3769 = ~n3757 & n3768 ;
  assign n3746 = ~\u5_dout_reg[18]/P0001  & ~n2770 ;
  assign n3770 = \u13_occ0_r_reg[16]/NET0131  & ~n3746 ;
  assign n3771 = ~n3769 & n3770 ;
  assign n3774 = \u5_mem_reg[2][31]/NET0131  & n2930 ;
  assign n3778 = \u5_rp_reg[0]/P0001  & ~n3774 ;
  assign n3777 = \u5_mem_reg[0][31]/NET0131  & n2932 ;
  assign n3775 = \u5_mem_reg[3][31]/NET0131  & n2776 ;
  assign n3776 = \u5_mem_reg[1][31]/NET0131  & n2928 ;
  assign n3779 = ~n3775 & ~n3776 ;
  assign n3780 = ~n3777 & n3779 ;
  assign n3781 = n3778 & n3780 ;
  assign n3773 = ~\u5_rp_reg[0]/P0001  & n3686 ;
  assign n3782 = n2771 & ~n3773 ;
  assign n3783 = ~n3781 & n3782 ;
  assign n3792 = n3536 & ~n3738 ;
  assign n3784 = \u5_mem_reg[2][19]/NET0131  & n2930 ;
  assign n3785 = \u5_mem_reg[3][19]/NET0131  & n2776 ;
  assign n3788 = ~n3784 & ~n3785 ;
  assign n3786 = \u5_mem_reg[1][19]/NET0131  & n2928 ;
  assign n3787 = \u5_mem_reg[0][19]/NET0131  & n2932 ;
  assign n3789 = ~n3786 & ~n3787 ;
  assign n3790 = n3788 & n3789 ;
  assign n3791 = n2937 & ~n3790 ;
  assign n3793 = n2770 & ~n3791 ;
  assign n3794 = ~n3792 & n3793 ;
  assign n3795 = ~n3783 & n3794 ;
  assign n3772 = ~\u5_dout_reg[19]/P0001  & ~n2770 ;
  assign n3796 = \u13_occ0_r_reg[16]/NET0131  & ~n3772 ;
  assign n3797 = ~n3795 & n3796 ;
  assign n3800 = \u5_mem_reg[1][2]/NET0131  & n2928 ;
  assign n3801 = \u5_mem_reg[0][2]/NET0131  & n2932 ;
  assign n3804 = ~n3800 & ~n3801 ;
  assign n3802 = \u5_mem_reg[2][2]/NET0131  & n2930 ;
  assign n3803 = \u5_mem_reg[3][2]/NET0131  & n2776 ;
  assign n3805 = ~n3802 & ~n3803 ;
  assign n3806 = n3804 & n3805 ;
  assign n3807 = n2937 & ~n3806 ;
  assign n3799 = ~n2936 & n3536 ;
  assign n3808 = n2770 & ~n3799 ;
  assign n3809 = ~n3807 & n3808 ;
  assign n3798 = ~\u5_dout_reg[2]/P0001  & ~n2770 ;
  assign n3810 = \u13_occ0_r_reg[16]/NET0131  & ~n3798 ;
  assign n3811 = ~n3809 & n3810 ;
  assign n3814 = \u5_mem_reg[3][3]/NET0131  & n2776 ;
  assign n3815 = \u5_mem_reg[2][3]/NET0131  & n2930 ;
  assign n3818 = ~n3814 & ~n3815 ;
  assign n3816 = \u5_mem_reg[1][3]/NET0131  & n2928 ;
  assign n3817 = \u5_mem_reg[0][3]/NET0131  & n2932 ;
  assign n3819 = ~n3816 & ~n3817 ;
  assign n3820 = n3818 & n3819 ;
  assign n3821 = n2937 & ~n3820 ;
  assign n3813 = ~n2949 & n3536 ;
  assign n3822 = n2770 & ~n3813 ;
  assign n3823 = ~n3821 & n3822 ;
  assign n3812 = ~\u5_dout_reg[3]/P0001  & ~n2770 ;
  assign n3824 = \u13_occ0_r_reg[16]/NET0131  & ~n3812 ;
  assign n3825 = ~n3823 & n3824 ;
  assign n3828 = \u5_rp_reg[0]/P0001  & n3712 ;
  assign n3827 = ~\u5_rp_reg[0]/P0001  & n2936 ;
  assign n3829 = n2771 & ~n3827 ;
  assign n3830 = ~n3828 & n3829 ;
  assign n3839 = n3536 & ~n3806 ;
  assign n3831 = \u5_mem_reg[3][4]/NET0131  & n2776 ;
  assign n3832 = \u5_mem_reg[1][4]/NET0131  & n2928 ;
  assign n3835 = ~n3831 & ~n3832 ;
  assign n3833 = \u5_mem_reg[2][4]/NET0131  & n2930 ;
  assign n3834 = \u5_mem_reg[0][4]/NET0131  & n2932 ;
  assign n3836 = ~n3833 & ~n3834 ;
  assign n3837 = n3835 & n3836 ;
  assign n3838 = n2937 & ~n3837 ;
  assign n3840 = n2770 & ~n3838 ;
  assign n3841 = ~n3839 & n3840 ;
  assign n3842 = ~n3830 & n3841 ;
  assign n3826 = ~\u5_dout_reg[4]/P0001  & ~n2770 ;
  assign n3843 = \u13_occ0_r_reg[16]/NET0131  & ~n3826 ;
  assign n3844 = ~n3842 & n3843 ;
  assign n3847 = \u5_rp_reg[0]/P0001  & n3738 ;
  assign n3846 = ~\u5_rp_reg[0]/P0001  & n2949 ;
  assign n3848 = n2771 & ~n3846 ;
  assign n3849 = ~n3847 & n3848 ;
  assign n3858 = n3536 & ~n3820 ;
  assign n3850 = \u5_mem_reg[1][5]/NET0131  & n2928 ;
  assign n3851 = \u5_mem_reg[2][5]/NET0131  & n2930 ;
  assign n3854 = ~n3850 & ~n3851 ;
  assign n3852 = \u5_mem_reg[3][5]/NET0131  & n2776 ;
  assign n3853 = \u5_mem_reg[0][5]/NET0131  & n2932 ;
  assign n3855 = ~n3852 & ~n3853 ;
  assign n3856 = n3854 & n3855 ;
  assign n3857 = n2937 & ~n3856 ;
  assign n3859 = n2770 & ~n3857 ;
  assign n3860 = ~n3858 & n3859 ;
  assign n3861 = ~n3849 & n3860 ;
  assign n3845 = ~\u5_dout_reg[5]/P0001  & ~n2770 ;
  assign n3862 = \u13_occ0_r_reg[16]/NET0131  & ~n3845 ;
  assign n3863 = ~n3861 & n3862 ;
  assign n3866 = \u5_rp_reg[0]/P0001  & n3764 ;
  assign n3865 = ~\u5_rp_reg[0]/P0001  & n3806 ;
  assign n3867 = n2771 & ~n3865 ;
  assign n3868 = ~n3866 & n3867 ;
  assign n3870 = n3536 & ~n3837 ;
  assign n3869 = n2937 & ~n3516 ;
  assign n3871 = n2770 & ~n3869 ;
  assign n3872 = ~n3870 & n3871 ;
  assign n3873 = ~n3868 & n3872 ;
  assign n3864 = ~\u5_dout_reg[6]/P0001  & ~n2770 ;
  assign n3874 = \u13_occ0_r_reg[16]/NET0131  & ~n3864 ;
  assign n3875 = ~n3873 & n3874 ;
  assign n3878 = \u5_rp_reg[0]/P0001  & n3790 ;
  assign n3877 = ~\u5_rp_reg[0]/P0001  & n3820 ;
  assign n3879 = n2771 & ~n3877 ;
  assign n3880 = ~n3878 & n3879 ;
  assign n3882 = n3536 & ~n3856 ;
  assign n3881 = n2937 & ~n3557 ;
  assign n3883 = n2770 & ~n3881 ;
  assign n3884 = ~n3882 & n3883 ;
  assign n3885 = ~n3880 & n3884 ;
  assign n3876 = ~\u5_dout_reg[7]/P0001  & ~n2770 ;
  assign n3886 = \u13_occ0_r_reg[16]/NET0131  & ~n3876 ;
  assign n3887 = ~n3885 & n3886 ;
  assign n3890 = \u5_mem_reg[2][20]/NET0131  & n2930 ;
  assign n3894 = \u5_rp_reg[0]/P0001  & ~n3890 ;
  assign n3893 = \u5_mem_reg[0][20]/NET0131  & n2932 ;
  assign n3891 = \u5_mem_reg[3][20]/NET0131  & n2776 ;
  assign n3892 = \u5_mem_reg[1][20]/NET0131  & n2928 ;
  assign n3895 = ~n3891 & ~n3892 ;
  assign n3896 = ~n3893 & n3895 ;
  assign n3897 = n3894 & n3896 ;
  assign n3889 = ~\u5_rp_reg[0]/P0001  & n3837 ;
  assign n3898 = n2771 & ~n3889 ;
  assign n3899 = ~n3897 & n3898 ;
  assign n3901 = ~n3516 & n3536 ;
  assign n3900 = n2937 & ~n3543 ;
  assign n3902 = n2770 & ~n3900 ;
  assign n3903 = ~n3901 & n3902 ;
  assign n3904 = ~n3899 & n3903 ;
  assign n3888 = ~\u5_dout_reg[8]/P0001  & ~n2770 ;
  assign n3905 = \u13_occ0_r_reg[16]/NET0131  & ~n3888 ;
  assign n3906 = ~n3904 & n3905 ;
  assign n3909 = \u5_mem_reg[2][21]/NET0131  & n2930 ;
  assign n3913 = \u5_rp_reg[0]/P0001  & ~n3909 ;
  assign n3912 = \u5_mem_reg[0][21]/NET0131  & n2932 ;
  assign n3910 = \u5_mem_reg[3][21]/NET0131  & n2776 ;
  assign n3911 = \u5_mem_reg[1][21]/NET0131  & n2928 ;
  assign n3914 = ~n3910 & ~n3911 ;
  assign n3915 = ~n3912 & n3914 ;
  assign n3916 = n3913 & n3915 ;
  assign n3908 = ~\u5_rp_reg[0]/P0001  & n3856 ;
  assign n3917 = n2771 & ~n3908 ;
  assign n3918 = ~n3916 & n3917 ;
  assign n3920 = n3536 & ~n3557 ;
  assign n3919 = n2937 & ~n3583 ;
  assign n3921 = n2770 & ~n3919 ;
  assign n3922 = ~n3920 & n3921 ;
  assign n3923 = ~n3918 & n3922 ;
  assign n3907 = ~\u5_dout_reg[9]/P0001  & ~n2770 ;
  assign n3924 = \u13_occ0_r_reg[16]/NET0131  & ~n3907 ;
  assign n3925 = ~n3923 & n3924 ;
  assign n3935 = \u6_mem_reg[2][22]/NET0131  & n2955 ;
  assign n3939 = \u6_rp_reg[0]/P0001  & ~n3935 ;
  assign n3938 = \u6_mem_reg[0][22]/NET0131  & n2959 ;
  assign n3936 = \u6_mem_reg[1][22]/NET0131  & n2957 ;
  assign n3937 = \u6_mem_reg[3][22]/NET0131  & n2801 ;
  assign n3940 = ~n3936 & ~n3937 ;
  assign n3941 = ~n3938 & n3940 ;
  assign n3942 = n3939 & n3941 ;
  assign n3927 = \u6_mem_reg[3][6]/NET0131  & n2801 ;
  assign n3928 = \u6_mem_reg[2][6]/NET0131  & n2955 ;
  assign n3931 = ~n3927 & ~n3928 ;
  assign n3929 = \u6_mem_reg[0][6]/NET0131  & n2959 ;
  assign n3930 = \u6_mem_reg[1][6]/NET0131  & n2957 ;
  assign n3932 = ~n3929 & ~n3930 ;
  assign n3933 = n3931 & n3932 ;
  assign n3934 = ~\u6_rp_reg[0]/P0001  & n3933 ;
  assign n3943 = n2796 & ~n3934 ;
  assign n3944 = ~n3942 & n3943 ;
  assign n3953 = \u13_occ0_r_reg[26]/NET0131  & ~\u13_occ0_r_reg[27]/NET0131  ;
  assign n3954 = \u6_mem_reg[3][8]/NET0131  & n2801 ;
  assign n3955 = \u6_mem_reg[2][8]/NET0131  & n2955 ;
  assign n3958 = ~n3954 & ~n3955 ;
  assign n3956 = \u6_mem_reg[0][8]/NET0131  & n2959 ;
  assign n3957 = \u6_mem_reg[1][8]/NET0131  & n2957 ;
  assign n3959 = ~n3956 & ~n3957 ;
  assign n3960 = n3958 & n3959 ;
  assign n3961 = n3953 & ~n3960 ;
  assign n3945 = \u6_mem_reg[1][10]/NET0131  & n2957 ;
  assign n3946 = \u6_mem_reg[3][10]/NET0131  & n2801 ;
  assign n3949 = ~n3945 & ~n3946 ;
  assign n3947 = \u6_mem_reg[0][10]/NET0131  & n2959 ;
  assign n3948 = \u6_mem_reg[2][10]/NET0131  & n2955 ;
  assign n3950 = ~n3947 & ~n3948 ;
  assign n3951 = n3949 & n3950 ;
  assign n3952 = n2964 & ~n3951 ;
  assign n3962 = n2795 & ~n3952 ;
  assign n3963 = ~n3961 & n3962 ;
  assign n3964 = ~n3944 & n3963 ;
  assign n3926 = ~\u6_dout_reg[10]/P0001  & ~n2795 ;
  assign n3965 = \u13_occ0_r_reg[24]/NET0131  & ~n3926 ;
  assign n3966 = ~n3964 & n3965 ;
  assign n3976 = \u6_mem_reg[2][23]/NET0131  & n2955 ;
  assign n3980 = \u6_rp_reg[0]/P0001  & ~n3976 ;
  assign n3979 = \u6_mem_reg[0][23]/NET0131  & n2959 ;
  assign n3977 = \u6_mem_reg[1][23]/NET0131  & n2957 ;
  assign n3978 = \u6_mem_reg[3][23]/NET0131  & n2801 ;
  assign n3981 = ~n3977 & ~n3978 ;
  assign n3982 = ~n3979 & n3981 ;
  assign n3983 = n3980 & n3982 ;
  assign n3968 = \u6_mem_reg[3][7]/NET0131  & n2801 ;
  assign n3969 = \u6_mem_reg[2][7]/NET0131  & n2955 ;
  assign n3972 = ~n3968 & ~n3969 ;
  assign n3970 = \u6_mem_reg[0][7]/NET0131  & n2959 ;
  assign n3971 = \u6_mem_reg[1][7]/NET0131  & n2957 ;
  assign n3973 = ~n3970 & ~n3971 ;
  assign n3974 = n3972 & n3973 ;
  assign n3975 = ~\u6_rp_reg[0]/P0001  & n3974 ;
  assign n3984 = n2796 & ~n3975 ;
  assign n3985 = ~n3983 & n3984 ;
  assign n3994 = \u6_mem_reg[3][9]/NET0131  & n2801 ;
  assign n3995 = \u6_mem_reg[1][9]/NET0131  & n2957 ;
  assign n3998 = ~n3994 & ~n3995 ;
  assign n3996 = \u6_mem_reg[2][9]/NET0131  & n2955 ;
  assign n3997 = \u6_mem_reg[0][9]/NET0131  & n2959 ;
  assign n3999 = ~n3996 & ~n3997 ;
  assign n4000 = n3998 & n3999 ;
  assign n4001 = n3953 & ~n4000 ;
  assign n3986 = \u6_mem_reg[3][11]/NET0131  & n2801 ;
  assign n3987 = \u6_mem_reg[2][11]/NET0131  & n2955 ;
  assign n3990 = ~n3986 & ~n3987 ;
  assign n3988 = \u6_mem_reg[0][11]/NET0131  & n2959 ;
  assign n3989 = \u6_mem_reg[1][11]/NET0131  & n2957 ;
  assign n3991 = ~n3988 & ~n3989 ;
  assign n3992 = n3990 & n3991 ;
  assign n3993 = n2964 & ~n3992 ;
  assign n4002 = n2795 & ~n3993 ;
  assign n4003 = ~n4001 & n4002 ;
  assign n4004 = ~n3985 & n4003 ;
  assign n3967 = ~\u6_dout_reg[11]/P0001  & ~n2795 ;
  assign n4005 = \u13_occ0_r_reg[24]/NET0131  & ~n3967 ;
  assign n4006 = ~n4004 & n4005 ;
  assign n4009 = \u6_mem_reg[2][24]/NET0131  & n2955 ;
  assign n4013 = \u6_rp_reg[0]/P0001  & ~n4009 ;
  assign n4012 = \u6_mem_reg[0][24]/NET0131  & n2959 ;
  assign n4010 = \u6_mem_reg[1][24]/NET0131  & n2957 ;
  assign n4011 = \u6_mem_reg[3][24]/NET0131  & n2801 ;
  assign n4014 = ~n4010 & ~n4011 ;
  assign n4015 = ~n4012 & n4014 ;
  assign n4016 = n4013 & n4015 ;
  assign n4008 = ~\u6_rp_reg[0]/P0001  & n3960 ;
  assign n4017 = n2796 & ~n4008 ;
  assign n4018 = ~n4016 & n4017 ;
  assign n4027 = ~n3951 & n3953 ;
  assign n4019 = \u6_mem_reg[3][12]/NET0131  & n2801 ;
  assign n4020 = \u6_mem_reg[1][12]/NET0131  & n2957 ;
  assign n4023 = ~n4019 & ~n4020 ;
  assign n4021 = \u6_mem_reg[0][12]/NET0131  & n2959 ;
  assign n4022 = \u6_mem_reg[2][12]/NET0131  & n2955 ;
  assign n4024 = ~n4021 & ~n4022 ;
  assign n4025 = n4023 & n4024 ;
  assign n4026 = n2964 & ~n4025 ;
  assign n4028 = n2795 & ~n4026 ;
  assign n4029 = ~n4027 & n4028 ;
  assign n4030 = ~n4018 & n4029 ;
  assign n4007 = ~\u6_dout_reg[12]/P0001  & ~n2795 ;
  assign n4031 = \u13_occ0_r_reg[24]/NET0131  & ~n4007 ;
  assign n4032 = ~n4030 & n4031 ;
  assign n4035 = \u6_mem_reg[2][25]/NET0131  & n2955 ;
  assign n4039 = \u6_rp_reg[0]/P0001  & ~n4035 ;
  assign n4038 = \u6_mem_reg[0][25]/NET0131  & n2959 ;
  assign n4036 = \u6_mem_reg[1][25]/NET0131  & n2957 ;
  assign n4037 = \u6_mem_reg[3][25]/NET0131  & n2801 ;
  assign n4040 = ~n4036 & ~n4037 ;
  assign n4041 = ~n4038 & n4040 ;
  assign n4042 = n4039 & n4041 ;
  assign n4034 = ~\u6_rp_reg[0]/P0001  & n4000 ;
  assign n4043 = n2796 & ~n4034 ;
  assign n4044 = ~n4042 & n4043 ;
  assign n4053 = n3953 & ~n3992 ;
  assign n4045 = \u6_mem_reg[3][13]/NET0131  & n2801 ;
  assign n4046 = \u6_mem_reg[2][13]/NET0131  & n2955 ;
  assign n4049 = ~n4045 & ~n4046 ;
  assign n4047 = \u6_mem_reg[0][13]/NET0131  & n2959 ;
  assign n4048 = \u6_mem_reg[1][13]/NET0131  & n2957 ;
  assign n4050 = ~n4047 & ~n4048 ;
  assign n4051 = n4049 & n4050 ;
  assign n4052 = n2964 & ~n4051 ;
  assign n4054 = n2795 & ~n4052 ;
  assign n4055 = ~n4053 & n4054 ;
  assign n4056 = ~n4044 & n4055 ;
  assign n4033 = ~\u6_dout_reg[13]/P0001  & ~n2795 ;
  assign n4057 = \u13_occ0_r_reg[24]/NET0131  & ~n4033 ;
  assign n4058 = ~n4056 & n4057 ;
  assign n4061 = \u6_mem_reg[2][26]/NET0131  & n2955 ;
  assign n4065 = \u6_rp_reg[0]/P0001  & ~n4061 ;
  assign n4064 = \u6_mem_reg[0][26]/NET0131  & n2959 ;
  assign n4062 = \u6_mem_reg[1][26]/NET0131  & n2957 ;
  assign n4063 = \u6_mem_reg[3][26]/NET0131  & n2801 ;
  assign n4066 = ~n4062 & ~n4063 ;
  assign n4067 = ~n4064 & n4066 ;
  assign n4068 = n4065 & n4067 ;
  assign n4060 = ~\u6_rp_reg[0]/P0001  & n3951 ;
  assign n4069 = n2796 & ~n4060 ;
  assign n4070 = ~n4068 & n4069 ;
  assign n4079 = n3953 & ~n4025 ;
  assign n4071 = \u6_mem_reg[1][14]/NET0131  & n2957 ;
  assign n4072 = \u6_mem_reg[0][14]/NET0131  & n2959 ;
  assign n4075 = ~n4071 & ~n4072 ;
  assign n4073 = \u6_mem_reg[3][14]/NET0131  & n2801 ;
  assign n4074 = \u6_mem_reg[2][14]/NET0131  & n2955 ;
  assign n4076 = ~n4073 & ~n4074 ;
  assign n4077 = n4075 & n4076 ;
  assign n4078 = n2964 & ~n4077 ;
  assign n4080 = n2795 & ~n4078 ;
  assign n4081 = ~n4079 & n4080 ;
  assign n4082 = ~n4070 & n4081 ;
  assign n4059 = ~\u6_dout_reg[14]/P0001  & ~n2795 ;
  assign n4083 = \u13_occ0_r_reg[24]/NET0131  & ~n4059 ;
  assign n4084 = ~n4082 & n4083 ;
  assign n4087 = \u6_mem_reg[2][27]/NET0131  & n2955 ;
  assign n4091 = \u6_rp_reg[0]/P0001  & ~n4087 ;
  assign n4090 = \u6_mem_reg[0][27]/NET0131  & n2959 ;
  assign n4088 = \u6_mem_reg[3][27]/NET0131  & n2801 ;
  assign n4089 = \u6_mem_reg[1][27]/NET0131  & n2957 ;
  assign n4092 = ~n4088 & ~n4089 ;
  assign n4093 = ~n4090 & n4092 ;
  assign n4094 = n4091 & n4093 ;
  assign n4086 = ~\u6_rp_reg[0]/P0001  & n3992 ;
  assign n4095 = n2796 & ~n4086 ;
  assign n4096 = ~n4094 & n4095 ;
  assign n4105 = n3953 & ~n4051 ;
  assign n4097 = \u6_mem_reg[3][15]/NET0131  & n2801 ;
  assign n4098 = \u6_mem_reg[2][15]/NET0131  & n2955 ;
  assign n4101 = ~n4097 & ~n4098 ;
  assign n4099 = \u6_mem_reg[0][15]/NET0131  & n2959 ;
  assign n4100 = \u6_mem_reg[1][15]/NET0131  & n2957 ;
  assign n4102 = ~n4099 & ~n4100 ;
  assign n4103 = n4101 & n4102 ;
  assign n4104 = n2964 & ~n4103 ;
  assign n4106 = n2795 & ~n4104 ;
  assign n4107 = ~n4105 & n4106 ;
  assign n4108 = ~n4096 & n4107 ;
  assign n4085 = ~\u6_dout_reg[15]/P0001  & ~n2795 ;
  assign n4109 = \u13_occ0_r_reg[24]/NET0131  & ~n4085 ;
  assign n4110 = ~n4108 & n4109 ;
  assign n4113 = \u6_mem_reg[2][28]/NET0131  & n2955 ;
  assign n4117 = \u6_rp_reg[0]/P0001  & ~n4113 ;
  assign n4116 = \u6_mem_reg[0][28]/NET0131  & n2959 ;
  assign n4114 = \u6_mem_reg[1][28]/NET0131  & n2957 ;
  assign n4115 = \u6_mem_reg[3][28]/NET0131  & n2801 ;
  assign n4118 = ~n4114 & ~n4115 ;
  assign n4119 = ~n4116 & n4118 ;
  assign n4120 = n4117 & n4119 ;
  assign n4112 = ~\u6_rp_reg[0]/P0001  & n4025 ;
  assign n4121 = n2796 & ~n4112 ;
  assign n4122 = ~n4120 & n4121 ;
  assign n4131 = n3953 & ~n4077 ;
  assign n4123 = \u6_mem_reg[1][16]/NET0131  & n2957 ;
  assign n4124 = \u6_mem_reg[0][16]/NET0131  & n2959 ;
  assign n4127 = ~n4123 & ~n4124 ;
  assign n4125 = \u6_mem_reg[2][16]/NET0131  & n2955 ;
  assign n4126 = \u6_mem_reg[3][16]/NET0131  & n2801 ;
  assign n4128 = ~n4125 & ~n4126 ;
  assign n4129 = n4127 & n4128 ;
  assign n4130 = n2964 & ~n4129 ;
  assign n4132 = n2795 & ~n4130 ;
  assign n4133 = ~n4131 & n4132 ;
  assign n4134 = ~n4122 & n4133 ;
  assign n4111 = ~\u6_dout_reg[16]/P0001  & ~n2795 ;
  assign n4135 = \u13_occ0_r_reg[24]/NET0131  & ~n4111 ;
  assign n4136 = ~n4134 & n4135 ;
  assign n4139 = \u6_mem_reg[2][29]/NET0131  & n2955 ;
  assign n4143 = \u6_rp_reg[0]/P0001  & ~n4139 ;
  assign n4142 = \u6_mem_reg[0][29]/NET0131  & n2959 ;
  assign n4140 = \u6_mem_reg[3][29]/NET0131  & n2801 ;
  assign n4141 = \u6_mem_reg[1][29]/NET0131  & n2957 ;
  assign n4144 = ~n4140 & ~n4141 ;
  assign n4145 = ~n4142 & n4144 ;
  assign n4146 = n4143 & n4145 ;
  assign n4138 = ~\u6_rp_reg[0]/P0001  & n4051 ;
  assign n4147 = n2796 & ~n4138 ;
  assign n4148 = ~n4146 & n4147 ;
  assign n4157 = n3953 & ~n4103 ;
  assign n4149 = \u6_mem_reg[3][17]/NET0131  & n2801 ;
  assign n4150 = \u6_mem_reg[1][17]/NET0131  & n2957 ;
  assign n4153 = ~n4149 & ~n4150 ;
  assign n4151 = \u6_mem_reg[2][17]/NET0131  & n2955 ;
  assign n4152 = \u6_mem_reg[0][17]/NET0131  & n2959 ;
  assign n4154 = ~n4151 & ~n4152 ;
  assign n4155 = n4153 & n4154 ;
  assign n4156 = n2964 & ~n4155 ;
  assign n4158 = n2795 & ~n4156 ;
  assign n4159 = ~n4157 & n4158 ;
  assign n4160 = ~n4148 & n4159 ;
  assign n4137 = ~\u6_dout_reg[17]/P0001  & ~n2795 ;
  assign n4161 = \u13_occ0_r_reg[24]/NET0131  & ~n4137 ;
  assign n4162 = ~n4160 & n4161 ;
  assign n4165 = \u6_mem_reg[2][30]/NET0131  & n2955 ;
  assign n4169 = \u6_rp_reg[0]/P0001  & ~n4165 ;
  assign n4168 = \u6_mem_reg[0][30]/NET0131  & n2959 ;
  assign n4166 = \u6_mem_reg[3][30]/NET0131  & n2801 ;
  assign n4167 = \u6_mem_reg[1][30]/NET0131  & n2957 ;
  assign n4170 = ~n4166 & ~n4167 ;
  assign n4171 = ~n4168 & n4170 ;
  assign n4172 = n4169 & n4171 ;
  assign n4164 = ~\u6_rp_reg[0]/P0001  & n4077 ;
  assign n4173 = n2796 & ~n4164 ;
  assign n4174 = ~n4172 & n4173 ;
  assign n4183 = n3953 & ~n4129 ;
  assign n4175 = \u6_mem_reg[1][18]/NET0131  & n2957 ;
  assign n4176 = \u6_mem_reg[3][18]/NET0131  & n2801 ;
  assign n4179 = ~n4175 & ~n4176 ;
  assign n4177 = \u6_mem_reg[2][18]/NET0131  & n2955 ;
  assign n4178 = \u6_mem_reg[0][18]/NET0131  & n2959 ;
  assign n4180 = ~n4177 & ~n4178 ;
  assign n4181 = n4179 & n4180 ;
  assign n4182 = n2964 & ~n4181 ;
  assign n4184 = n2795 & ~n4182 ;
  assign n4185 = ~n4183 & n4184 ;
  assign n4186 = ~n4174 & n4185 ;
  assign n4163 = ~\u6_dout_reg[18]/P0001  & ~n2795 ;
  assign n4187 = \u13_occ0_r_reg[24]/NET0131  & ~n4163 ;
  assign n4188 = ~n4186 & n4187 ;
  assign n4191 = \u6_mem_reg[2][31]/NET0131  & n2955 ;
  assign n4195 = \u6_rp_reg[0]/P0001  & ~n4191 ;
  assign n4194 = \u6_mem_reg[0][31]/NET0131  & n2959 ;
  assign n4192 = \u6_mem_reg[3][31]/NET0131  & n2801 ;
  assign n4193 = \u6_mem_reg[1][31]/NET0131  & n2957 ;
  assign n4196 = ~n4192 & ~n4193 ;
  assign n4197 = ~n4194 & n4196 ;
  assign n4198 = n4195 & n4197 ;
  assign n4190 = ~\u6_rp_reg[0]/P0001  & n4103 ;
  assign n4199 = n2796 & ~n4190 ;
  assign n4200 = ~n4198 & n4199 ;
  assign n4209 = n3953 & ~n4155 ;
  assign n4201 = \u6_mem_reg[2][19]/NET0131  & n2955 ;
  assign n4202 = \u6_mem_reg[3][19]/NET0131  & n2801 ;
  assign n4205 = ~n4201 & ~n4202 ;
  assign n4203 = \u6_mem_reg[1][19]/NET0131  & n2957 ;
  assign n4204 = \u6_mem_reg[0][19]/NET0131  & n2959 ;
  assign n4206 = ~n4203 & ~n4204 ;
  assign n4207 = n4205 & n4206 ;
  assign n4208 = n2964 & ~n4207 ;
  assign n4210 = n2795 & ~n4208 ;
  assign n4211 = ~n4209 & n4210 ;
  assign n4212 = ~n4200 & n4211 ;
  assign n4189 = ~\u6_dout_reg[19]/P0001  & ~n2795 ;
  assign n4213 = \u13_occ0_r_reg[24]/NET0131  & ~n4189 ;
  assign n4214 = ~n4212 & n4213 ;
  assign n4217 = \u6_mem_reg[3][2]/NET0131  & n2801 ;
  assign n4218 = \u6_mem_reg[2][2]/NET0131  & n2955 ;
  assign n4221 = ~n4217 & ~n4218 ;
  assign n4219 = \u6_mem_reg[1][2]/NET0131  & n2957 ;
  assign n4220 = \u6_mem_reg[0][2]/NET0131  & n2959 ;
  assign n4222 = ~n4219 & ~n4220 ;
  assign n4223 = n4221 & n4222 ;
  assign n4224 = n2964 & ~n4223 ;
  assign n4216 = ~n2963 & n3953 ;
  assign n4225 = n2795 & ~n4216 ;
  assign n4226 = ~n4224 & n4225 ;
  assign n4215 = ~\u6_dout_reg[2]/P0001  & ~n2795 ;
  assign n4227 = \u13_occ0_r_reg[24]/NET0131  & ~n4215 ;
  assign n4228 = ~n4226 & n4227 ;
  assign n4231 = \u6_mem_reg[3][3]/NET0131  & n2801 ;
  assign n4232 = \u6_mem_reg[1][3]/NET0131  & n2957 ;
  assign n4235 = ~n4231 & ~n4232 ;
  assign n4233 = \u6_mem_reg[2][3]/NET0131  & n2955 ;
  assign n4234 = \u6_mem_reg[0][3]/NET0131  & n2959 ;
  assign n4236 = ~n4233 & ~n4234 ;
  assign n4237 = n4235 & n4236 ;
  assign n4238 = n2964 & ~n4237 ;
  assign n4230 = ~n2976 & n3953 ;
  assign n4239 = n2795 & ~n4230 ;
  assign n4240 = ~n4238 & n4239 ;
  assign n4229 = ~\u6_dout_reg[3]/P0001  & ~n2795 ;
  assign n4241 = \u13_occ0_r_reg[24]/NET0131  & ~n4229 ;
  assign n4242 = ~n4240 & n4241 ;
  assign n4245 = \u6_rp_reg[0]/P0001  & n4129 ;
  assign n4244 = ~\u6_rp_reg[0]/P0001  & n2963 ;
  assign n4246 = n2796 & ~n4244 ;
  assign n4247 = ~n4245 & n4246 ;
  assign n4256 = n3953 & ~n4223 ;
  assign n4248 = \u6_mem_reg[3][4]/NET0131  & n2801 ;
  assign n4249 = \u6_mem_reg[2][4]/NET0131  & n2955 ;
  assign n4252 = ~n4248 & ~n4249 ;
  assign n4250 = \u6_mem_reg[0][4]/NET0131  & n2959 ;
  assign n4251 = \u6_mem_reg[1][4]/NET0131  & n2957 ;
  assign n4253 = ~n4250 & ~n4251 ;
  assign n4254 = n4252 & n4253 ;
  assign n4255 = n2964 & ~n4254 ;
  assign n4257 = n2795 & ~n4255 ;
  assign n4258 = ~n4256 & n4257 ;
  assign n4259 = ~n4247 & n4258 ;
  assign n4243 = ~\u6_dout_reg[4]/P0001  & ~n2795 ;
  assign n4260 = \u13_occ0_r_reg[24]/NET0131  & ~n4243 ;
  assign n4261 = ~n4259 & n4260 ;
  assign n4264 = \u6_rp_reg[0]/P0001  & n4155 ;
  assign n4263 = ~\u6_rp_reg[0]/P0001  & n2976 ;
  assign n4265 = n2796 & ~n4263 ;
  assign n4266 = ~n4264 & n4265 ;
  assign n4275 = n3953 & ~n4237 ;
  assign n4267 = \u6_mem_reg[3][5]/NET0131  & n2801 ;
  assign n4268 = \u6_mem_reg[2][5]/NET0131  & n2955 ;
  assign n4271 = ~n4267 & ~n4268 ;
  assign n4269 = \u6_mem_reg[0][5]/NET0131  & n2959 ;
  assign n4270 = \u6_mem_reg[1][5]/NET0131  & n2957 ;
  assign n4272 = ~n4269 & ~n4270 ;
  assign n4273 = n4271 & n4272 ;
  assign n4274 = n2964 & ~n4273 ;
  assign n4276 = n2795 & ~n4274 ;
  assign n4277 = ~n4275 & n4276 ;
  assign n4278 = ~n4266 & n4277 ;
  assign n4262 = ~\u6_dout_reg[5]/P0001  & ~n2795 ;
  assign n4279 = \u13_occ0_r_reg[24]/NET0131  & ~n4262 ;
  assign n4280 = ~n4278 & n4279 ;
  assign n4283 = \u6_rp_reg[0]/P0001  & n4181 ;
  assign n4282 = ~\u6_rp_reg[0]/P0001  & n4223 ;
  assign n4284 = n2796 & ~n4282 ;
  assign n4285 = ~n4283 & n4284 ;
  assign n4287 = n3953 & ~n4254 ;
  assign n4286 = n2964 & ~n3933 ;
  assign n4288 = n2795 & ~n4286 ;
  assign n4289 = ~n4287 & n4288 ;
  assign n4290 = ~n4285 & n4289 ;
  assign n4281 = ~\u6_dout_reg[6]/P0001  & ~n2795 ;
  assign n4291 = \u13_occ0_r_reg[24]/NET0131  & ~n4281 ;
  assign n4292 = ~n4290 & n4291 ;
  assign n4295 = \u6_rp_reg[0]/P0001  & n4207 ;
  assign n4294 = ~\u6_rp_reg[0]/P0001  & n4237 ;
  assign n4296 = n2796 & ~n4294 ;
  assign n4297 = ~n4295 & n4296 ;
  assign n4299 = n3953 & ~n4273 ;
  assign n4298 = n2964 & ~n3974 ;
  assign n4300 = n2795 & ~n4298 ;
  assign n4301 = ~n4299 & n4300 ;
  assign n4302 = ~n4297 & n4301 ;
  assign n4293 = ~\u6_dout_reg[7]/P0001  & ~n2795 ;
  assign n4303 = \u13_occ0_r_reg[24]/NET0131  & ~n4293 ;
  assign n4304 = ~n4302 & n4303 ;
  assign n4307 = \u6_mem_reg[2][20]/NET0131  & n2955 ;
  assign n4311 = \u6_rp_reg[0]/P0001  & ~n4307 ;
  assign n4310 = \u6_mem_reg[0][20]/NET0131  & n2959 ;
  assign n4308 = \u6_mem_reg[3][20]/NET0131  & n2801 ;
  assign n4309 = \u6_mem_reg[1][20]/NET0131  & n2957 ;
  assign n4312 = ~n4308 & ~n4309 ;
  assign n4313 = ~n4310 & n4312 ;
  assign n4314 = n4311 & n4313 ;
  assign n4306 = ~\u6_rp_reg[0]/P0001  & n4254 ;
  assign n4315 = n2796 & ~n4306 ;
  assign n4316 = ~n4314 & n4315 ;
  assign n4318 = ~n3933 & n3953 ;
  assign n4317 = n2964 & ~n3960 ;
  assign n4319 = n2795 & ~n4317 ;
  assign n4320 = ~n4318 & n4319 ;
  assign n4321 = ~n4316 & n4320 ;
  assign n4305 = ~\u6_dout_reg[8]/P0001  & ~n2795 ;
  assign n4322 = \u13_occ0_r_reg[24]/NET0131  & ~n4305 ;
  assign n4323 = ~n4321 & n4322 ;
  assign n4326 = \u6_mem_reg[2][21]/NET0131  & n2955 ;
  assign n4330 = \u6_rp_reg[0]/P0001  & ~n4326 ;
  assign n4329 = \u6_mem_reg[0][21]/NET0131  & n2959 ;
  assign n4327 = \u6_mem_reg[1][21]/NET0131  & n2957 ;
  assign n4328 = \u6_mem_reg[3][21]/NET0131  & n2801 ;
  assign n4331 = ~n4327 & ~n4328 ;
  assign n4332 = ~n4329 & n4331 ;
  assign n4333 = n4330 & n4332 ;
  assign n4325 = ~\u6_rp_reg[0]/P0001  & n4273 ;
  assign n4334 = n2796 & ~n4325 ;
  assign n4335 = ~n4333 & n4334 ;
  assign n4337 = n3953 & ~n3974 ;
  assign n4336 = n2964 & ~n4000 ;
  assign n4338 = n2795 & ~n4336 ;
  assign n4339 = ~n4337 & n4338 ;
  assign n4340 = ~n4335 & n4339 ;
  assign n4324 = ~\u6_dout_reg[9]/P0001  & ~n2795 ;
  assign n4341 = \u13_occ0_r_reg[24]/NET0131  & ~n4324 ;
  assign n4342 = ~n4340 & n4341 ;
  assign n4344 = \u7_mem_reg[2][6]/NET0131  & n2983 ;
  assign n4345 = \u7_mem_reg[3][6]/NET0131  & n2981 ;
  assign n4348 = ~n4344 & ~n4345 ;
  assign n4346 = \u7_mem_reg[0][6]/NET0131  & n2987 ;
  assign n4347 = \u7_mem_reg[1][6]/NET0131  & n2985 ;
  assign n4349 = ~n4346 & ~n4347 ;
  assign n4350 = n4348 & n4349 ;
  assign n4351 = n2806 & ~n4350 ;
  assign n4378 = n2808 & ~n4351 ;
  assign n4370 = \u7_mem_reg[3][10]/NET0131  & n2981 ;
  assign n4371 = \u7_mem_reg[2][10]/NET0131  & n2983 ;
  assign n4374 = ~n4370 & ~n4371 ;
  assign n4372 = \u7_mem_reg[1][10]/NET0131  & n2985 ;
  assign n4373 = \u7_mem_reg[0][10]/NET0131  & n2987 ;
  assign n4375 = ~n4372 & ~n4373 ;
  assign n4376 = n4374 & n4375 ;
  assign n4377 = n2992 & ~n4376 ;
  assign n4352 = \u13_occ1_r_reg[2]/NET0131  & ~\u13_occ1_r_reg[3]/NET0131  ;
  assign n4353 = \u7_mem_reg[3][8]/NET0131  & n2981 ;
  assign n4354 = \u7_mem_reg[2][8]/NET0131  & n2983 ;
  assign n4357 = ~n4353 & ~n4354 ;
  assign n4355 = \u7_mem_reg[1][8]/NET0131  & n2985 ;
  assign n4356 = \u7_mem_reg[0][8]/NET0131  & n2987 ;
  assign n4358 = ~n4355 & ~n4356 ;
  assign n4359 = n4357 & n4358 ;
  assign n4360 = n4352 & ~n4359 ;
  assign n4361 = \u7_rp_reg[0]/P0001  & n2805 ;
  assign n4362 = \u7_mem_reg[3][22]/NET0131  & n2981 ;
  assign n4363 = \u7_mem_reg[0][22]/NET0131  & n2987 ;
  assign n4366 = ~n4362 & ~n4363 ;
  assign n4364 = \u7_mem_reg[1][22]/NET0131  & n2985 ;
  assign n4365 = \u7_mem_reg[2][22]/NET0131  & n2983 ;
  assign n4367 = ~n4364 & ~n4365 ;
  assign n4368 = n4366 & n4367 ;
  assign n4369 = n4361 & ~n4368 ;
  assign n4379 = ~n4360 & ~n4369 ;
  assign n4380 = ~n4377 & n4379 ;
  assign n4381 = n4378 & n4380 ;
  assign n4343 = ~\u7_dout_reg[10]/P0001  & ~n2808 ;
  assign n4382 = \u13_occ1_r_reg[0]/NET0131  & ~n4343 ;
  assign n4383 = ~n4381 & n4382 ;
  assign n4385 = \u7_mem_reg[1][11]/NET0131  & n2985 ;
  assign n4386 = \u7_mem_reg[2][11]/NET0131  & n2983 ;
  assign n4389 = ~n4385 & ~n4386 ;
  assign n4387 = \u7_mem_reg[0][11]/NET0131  & n2987 ;
  assign n4388 = \u7_mem_reg[3][11]/NET0131  & n2981 ;
  assign n4390 = ~n4387 & ~n4388 ;
  assign n4391 = n4389 & n4390 ;
  assign n4392 = n2992 & ~n4391 ;
  assign n4417 = n2808 & ~n4392 ;
  assign n4409 = \u7_mem_reg[3][9]/NET0131  & n2981 ;
  assign n4410 = \u7_mem_reg[0][9]/NET0131  & n2987 ;
  assign n4413 = ~n4409 & ~n4410 ;
  assign n4411 = \u7_mem_reg[2][9]/NET0131  & n2983 ;
  assign n4412 = \u7_mem_reg[1][9]/NET0131  & n2985 ;
  assign n4414 = ~n4411 & ~n4412 ;
  assign n4415 = n4413 & n4414 ;
  assign n4416 = n4352 & ~n4415 ;
  assign n4393 = \u7_mem_reg[1][7]/NET0131  & n2985 ;
  assign n4394 = \u7_mem_reg[3][7]/NET0131  & n2981 ;
  assign n4397 = ~n4393 & ~n4394 ;
  assign n4395 = \u7_mem_reg[2][7]/NET0131  & n2983 ;
  assign n4396 = \u7_mem_reg[0][7]/NET0131  & n2987 ;
  assign n4398 = ~n4395 & ~n4396 ;
  assign n4399 = n4397 & n4398 ;
  assign n4400 = n2806 & ~n4399 ;
  assign n4401 = \u7_mem_reg[2][23]/NET0131  & n2983 ;
  assign n4402 = \u7_mem_reg[0][23]/NET0131  & n2987 ;
  assign n4405 = ~n4401 & ~n4402 ;
  assign n4403 = \u7_mem_reg[1][23]/NET0131  & n2985 ;
  assign n4404 = \u7_mem_reg[3][23]/NET0131  & n2981 ;
  assign n4406 = ~n4403 & ~n4404 ;
  assign n4407 = n4405 & n4406 ;
  assign n4408 = n4361 & ~n4407 ;
  assign n4418 = ~n4400 & ~n4408 ;
  assign n4419 = ~n4416 & n4418 ;
  assign n4420 = n4417 & n4419 ;
  assign n4384 = ~\u7_dout_reg[11]/P0001  & ~n2808 ;
  assign n4421 = \u13_occ1_r_reg[0]/NET0131  & ~n4384 ;
  assign n4422 = ~n4420 & n4421 ;
  assign n4424 = \u13_icc_r_reg[5]/NET0131  & \u9_status_reg[1]/P0001  ;
  assign n4425 = ~\u13_icc_r_reg[4]/NET0131  & ~\u9_status_reg[0]/P0001  ;
  assign n4426 = ~n4424 & n4425 ;
  assign n4423 = ~\u13_icc_r_reg[5]/NET0131  & ~\u9_status_reg[1]/P0001  ;
  assign n4427 = ~\u9_full_reg/NET0131  & ~n4423 ;
  assign n4428 = ~n4426 & n4427 ;
  assign n4429 = \u13_icc_r_reg[0]/NET0131  & ~n4428 ;
  assign n4432 = \u7_mem_reg[2][24]/NET0131  & n2983 ;
  assign n4436 = \u7_rp_reg[0]/P0001  & ~n4432 ;
  assign n4435 = \u7_mem_reg[0][24]/NET0131  & n2987 ;
  assign n4433 = \u7_mem_reg[3][24]/NET0131  & n2981 ;
  assign n4434 = \u7_mem_reg[1][24]/NET0131  & n2985 ;
  assign n4437 = ~n4433 & ~n4434 ;
  assign n4438 = ~n4435 & n4437 ;
  assign n4439 = n4436 & n4438 ;
  assign n4431 = ~\u7_rp_reg[0]/P0001  & n4359 ;
  assign n4440 = n2805 & ~n4431 ;
  assign n4441 = ~n4439 & n4440 ;
  assign n4450 = n4352 & ~n4376 ;
  assign n4442 = \u7_mem_reg[3][12]/NET0131  & n2981 ;
  assign n4443 = \u7_mem_reg[2][12]/NET0131  & n2983 ;
  assign n4446 = ~n4442 & ~n4443 ;
  assign n4444 = \u7_mem_reg[1][12]/NET0131  & n2985 ;
  assign n4445 = \u7_mem_reg[0][12]/NET0131  & n2987 ;
  assign n4447 = ~n4444 & ~n4445 ;
  assign n4448 = n4446 & n4447 ;
  assign n4449 = n2992 & ~n4448 ;
  assign n4451 = n2808 & ~n4449 ;
  assign n4452 = ~n4450 & n4451 ;
  assign n4453 = ~n4441 & n4452 ;
  assign n4430 = ~\u7_dout_reg[12]/P0001  & ~n2808 ;
  assign n4454 = \u13_occ1_r_reg[0]/NET0131  & ~n4430 ;
  assign n4455 = ~n4453 & n4454 ;
  assign n4456 = \u10_status_reg[1]/P0001  & \u13_icc_r_reg[13]/NET0131  ;
  assign n4457 = ~\u10_status_reg[0]/P0001  & ~\u13_icc_r_reg[12]/NET0131  ;
  assign n4458 = ~n4456 & n4457 ;
  assign n4459 = ~\u10_status_reg[1]/P0001  & ~\u13_icc_r_reg[13]/NET0131  ;
  assign n4460 = ~\u10_full_reg/NET0131  & ~n4459 ;
  assign n4461 = ~n4458 & n4460 ;
  assign n4462 = \u13_icc_r_reg[8]/NET0131  & ~n4461 ;
  assign n4474 = \u7_mem_reg[2][25]/NET0131  & n2983 ;
  assign n4478 = \u7_rp_reg[0]/P0001  & ~n4474 ;
  assign n4477 = \u7_mem_reg[0][25]/NET0131  & n2987 ;
  assign n4475 = \u7_mem_reg[3][25]/NET0131  & n2981 ;
  assign n4476 = \u7_mem_reg[1][25]/NET0131  & n2985 ;
  assign n4479 = ~n4475 & ~n4476 ;
  assign n4480 = ~n4477 & n4479 ;
  assign n4481 = n4478 & n4480 ;
  assign n4473 = ~\u7_rp_reg[0]/P0001  & n4415 ;
  assign n4482 = n2805 & ~n4473 ;
  assign n4483 = ~n4481 & n4482 ;
  assign n4465 = \u7_mem_reg[3][13]/NET0131  & n2981 ;
  assign n4466 = \u7_mem_reg[2][13]/NET0131  & n2983 ;
  assign n4469 = ~n4465 & ~n4466 ;
  assign n4467 = \u7_mem_reg[1][13]/NET0131  & n2985 ;
  assign n4468 = \u7_mem_reg[0][13]/NET0131  & n2987 ;
  assign n4470 = ~n4467 & ~n4468 ;
  assign n4471 = n4469 & n4470 ;
  assign n4472 = n2992 & ~n4471 ;
  assign n4464 = n4352 & ~n4391 ;
  assign n4484 = n2808 & ~n4464 ;
  assign n4485 = ~n4472 & n4484 ;
  assign n4486 = ~n4483 & n4485 ;
  assign n4463 = ~\u7_dout_reg[13]/P0001  & ~n2808 ;
  assign n4487 = \u13_occ1_r_reg[0]/NET0131  & ~n4463 ;
  assign n4488 = ~n4486 & n4487 ;
  assign n4491 = \u7_mem_reg[2][26]/NET0131  & n2983 ;
  assign n4495 = \u7_rp_reg[0]/P0001  & ~n4491 ;
  assign n4494 = \u7_mem_reg[0][26]/NET0131  & n2987 ;
  assign n4492 = \u7_mem_reg[3][26]/NET0131  & n2981 ;
  assign n4493 = \u7_mem_reg[1][26]/NET0131  & n2985 ;
  assign n4496 = ~n4492 & ~n4493 ;
  assign n4497 = ~n4494 & n4496 ;
  assign n4498 = n4495 & n4497 ;
  assign n4490 = ~\u7_rp_reg[0]/P0001  & n4376 ;
  assign n4499 = n2805 & ~n4490 ;
  assign n4500 = ~n4498 & n4499 ;
  assign n4509 = n4352 & ~n4448 ;
  assign n4501 = \u7_mem_reg[3][14]/NET0131  & n2981 ;
  assign n4502 = \u7_mem_reg[2][14]/NET0131  & n2983 ;
  assign n4505 = ~n4501 & ~n4502 ;
  assign n4503 = \u7_mem_reg[1][14]/NET0131  & n2985 ;
  assign n4504 = \u7_mem_reg[0][14]/NET0131  & n2987 ;
  assign n4506 = ~n4503 & ~n4504 ;
  assign n4507 = n4505 & n4506 ;
  assign n4508 = n2992 & ~n4507 ;
  assign n4510 = n2808 & ~n4508 ;
  assign n4511 = ~n4509 & n4510 ;
  assign n4512 = ~n4500 & n4511 ;
  assign n4489 = ~\u7_dout_reg[14]/P0001  & ~n2808 ;
  assign n4513 = \u13_occ1_r_reg[0]/NET0131  & ~n4489 ;
  assign n4514 = ~n4512 & n4513 ;
  assign n4516 = n2806 & ~n4391 ;
  assign n4534 = n2808 & ~n4516 ;
  assign n4526 = \u7_mem_reg[1][15]/NET0131  & n2985 ;
  assign n4527 = \u7_mem_reg[3][15]/NET0131  & n2981 ;
  assign n4530 = ~n4526 & ~n4527 ;
  assign n4528 = \u7_mem_reg[2][15]/NET0131  & n2983 ;
  assign n4529 = \u7_mem_reg[0][15]/NET0131  & n2987 ;
  assign n4531 = ~n4528 & ~n4529 ;
  assign n4532 = n4530 & n4531 ;
  assign n4533 = n2992 & ~n4532 ;
  assign n4517 = n4352 & ~n4471 ;
  assign n4518 = \u7_mem_reg[1][27]/NET0131  & n2985 ;
  assign n4519 = \u7_mem_reg[0][27]/NET0131  & n2987 ;
  assign n4522 = ~n4518 & ~n4519 ;
  assign n4520 = \u7_mem_reg[2][27]/NET0131  & n2983 ;
  assign n4521 = \u7_mem_reg[3][27]/NET0131  & n2981 ;
  assign n4523 = ~n4520 & ~n4521 ;
  assign n4524 = n4522 & n4523 ;
  assign n4525 = n4361 & ~n4524 ;
  assign n4535 = ~n4517 & ~n4525 ;
  assign n4536 = ~n4533 & n4535 ;
  assign n4537 = n4534 & n4536 ;
  assign n4515 = ~\u7_dout_reg[15]/P0001  & ~n2808 ;
  assign n4538 = \u13_occ1_r_reg[0]/NET0131  & ~n4515 ;
  assign n4539 = ~n4537 & n4538 ;
  assign n4542 = \u7_mem_reg[2][28]/NET0131  & n2983 ;
  assign n4546 = \u7_rp_reg[0]/P0001  & ~n4542 ;
  assign n4545 = \u7_mem_reg[0][28]/NET0131  & n2987 ;
  assign n4543 = \u7_mem_reg[3][28]/NET0131  & n2981 ;
  assign n4544 = \u7_mem_reg[1][28]/NET0131  & n2985 ;
  assign n4547 = ~n4543 & ~n4544 ;
  assign n4548 = ~n4545 & n4547 ;
  assign n4549 = n4546 & n4548 ;
  assign n4541 = ~\u7_rp_reg[0]/P0001  & n4448 ;
  assign n4550 = n2805 & ~n4541 ;
  assign n4551 = ~n4549 & n4550 ;
  assign n4560 = n4352 & ~n4507 ;
  assign n4552 = \u7_mem_reg[3][16]/NET0131  & n2981 ;
  assign n4553 = \u7_mem_reg[2][16]/NET0131  & n2983 ;
  assign n4556 = ~n4552 & ~n4553 ;
  assign n4554 = \u7_mem_reg[1][16]/NET0131  & n2985 ;
  assign n4555 = \u7_mem_reg[0][16]/NET0131  & n2987 ;
  assign n4557 = ~n4554 & ~n4555 ;
  assign n4558 = n4556 & n4557 ;
  assign n4559 = n2992 & ~n4558 ;
  assign n4561 = n2808 & ~n4559 ;
  assign n4562 = ~n4560 & n4561 ;
  assign n4563 = ~n4551 & n4562 ;
  assign n4540 = ~\u7_dout_reg[16]/P0001  & ~n2808 ;
  assign n4564 = \u13_occ1_r_reg[0]/NET0131  & ~n4540 ;
  assign n4565 = ~n4563 & n4564 ;
  assign n4568 = \u7_mem_reg[2][29]/NET0131  & n2983 ;
  assign n4572 = \u7_rp_reg[0]/P0001  & ~n4568 ;
  assign n4571 = \u7_mem_reg[0][29]/NET0131  & n2987 ;
  assign n4569 = \u7_mem_reg[3][29]/NET0131  & n2981 ;
  assign n4570 = \u7_mem_reg[1][29]/NET0131  & n2985 ;
  assign n4573 = ~n4569 & ~n4570 ;
  assign n4574 = ~n4571 & n4573 ;
  assign n4575 = n4572 & n4574 ;
  assign n4567 = ~\u7_rp_reg[0]/P0001  & n4471 ;
  assign n4576 = n2805 & ~n4567 ;
  assign n4577 = ~n4575 & n4576 ;
  assign n4586 = n4352 & ~n4532 ;
  assign n4578 = \u7_mem_reg[1][17]/NET0131  & n2985 ;
  assign n4579 = \u7_mem_reg[3][17]/NET0131  & n2981 ;
  assign n4582 = ~n4578 & ~n4579 ;
  assign n4580 = \u7_mem_reg[2][17]/NET0131  & n2983 ;
  assign n4581 = \u7_mem_reg[0][17]/NET0131  & n2987 ;
  assign n4583 = ~n4580 & ~n4581 ;
  assign n4584 = n4582 & n4583 ;
  assign n4585 = n2992 & ~n4584 ;
  assign n4587 = n2808 & ~n4585 ;
  assign n4588 = ~n4586 & n4587 ;
  assign n4589 = ~n4577 & n4588 ;
  assign n4566 = ~\u7_dout_reg[17]/P0001  & ~n2808 ;
  assign n4590 = \u13_occ1_r_reg[0]/NET0131  & ~n4566 ;
  assign n4591 = ~n4589 & n4590 ;
  assign n4594 = \u7_mem_reg[2][30]/NET0131  & n2983 ;
  assign n4598 = \u7_rp_reg[0]/P0001  & ~n4594 ;
  assign n4597 = \u7_mem_reg[0][30]/NET0131  & n2987 ;
  assign n4595 = \u7_mem_reg[3][30]/NET0131  & n2981 ;
  assign n4596 = \u7_mem_reg[1][30]/NET0131  & n2985 ;
  assign n4599 = ~n4595 & ~n4596 ;
  assign n4600 = ~n4597 & n4599 ;
  assign n4601 = n4598 & n4600 ;
  assign n4593 = ~\u7_rp_reg[0]/P0001  & n4507 ;
  assign n4602 = n2805 & ~n4593 ;
  assign n4603 = ~n4601 & n4602 ;
  assign n4612 = n4352 & ~n4558 ;
  assign n4604 = \u7_mem_reg[2][18]/NET0131  & n2983 ;
  assign n4605 = \u7_mem_reg[1][18]/NET0131  & n2985 ;
  assign n4608 = ~n4604 & ~n4605 ;
  assign n4606 = \u7_mem_reg[3][18]/NET0131  & n2981 ;
  assign n4607 = \u7_mem_reg[0][18]/NET0131  & n2987 ;
  assign n4609 = ~n4606 & ~n4607 ;
  assign n4610 = n4608 & n4609 ;
  assign n4611 = n2992 & ~n4610 ;
  assign n4613 = n2808 & ~n4611 ;
  assign n4614 = ~n4612 & n4613 ;
  assign n4615 = ~n4603 & n4614 ;
  assign n4592 = ~\u7_dout_reg[18]/P0001  & ~n2808 ;
  assign n4616 = \u13_occ1_r_reg[0]/NET0131  & ~n4592 ;
  assign n4617 = ~n4615 & n4616 ;
  assign n4620 = \u7_mem_reg[2][31]/NET0131  & n2983 ;
  assign n4624 = \u7_rp_reg[0]/P0001  & ~n4620 ;
  assign n4623 = \u7_mem_reg[0][31]/NET0131  & n2987 ;
  assign n4621 = \u7_mem_reg[3][31]/NET0131  & n2981 ;
  assign n4622 = \u7_mem_reg[1][31]/NET0131  & n2985 ;
  assign n4625 = ~n4621 & ~n4622 ;
  assign n4626 = ~n4623 & n4625 ;
  assign n4627 = n4624 & n4626 ;
  assign n4619 = ~\u7_rp_reg[0]/P0001  & n4532 ;
  assign n4628 = n2805 & ~n4619 ;
  assign n4629 = ~n4627 & n4628 ;
  assign n4638 = n4352 & ~n4584 ;
  assign n4630 = \u7_mem_reg[3][19]/NET0131  & n2981 ;
  assign n4631 = \u7_mem_reg[0][19]/NET0131  & n2987 ;
  assign n4634 = ~n4630 & ~n4631 ;
  assign n4632 = \u7_mem_reg[1][19]/NET0131  & n2985 ;
  assign n4633 = \u7_mem_reg[2][19]/NET0131  & n2983 ;
  assign n4635 = ~n4632 & ~n4633 ;
  assign n4636 = n4634 & n4635 ;
  assign n4637 = n2992 & ~n4636 ;
  assign n4639 = n2808 & ~n4637 ;
  assign n4640 = ~n4638 & n4639 ;
  assign n4641 = ~n4629 & n4640 ;
  assign n4618 = ~\u7_dout_reg[19]/P0001  & ~n2808 ;
  assign n4642 = \u13_occ1_r_reg[0]/NET0131  & ~n4618 ;
  assign n4643 = ~n4641 & n4642 ;
  assign n4646 = \u7_mem_reg[3][2]/NET0131  & n2981 ;
  assign n4647 = \u7_mem_reg[2][2]/NET0131  & n2983 ;
  assign n4650 = ~n4646 & ~n4647 ;
  assign n4648 = \u7_mem_reg[1][2]/NET0131  & n2985 ;
  assign n4649 = \u7_mem_reg[0][2]/NET0131  & n2987 ;
  assign n4651 = ~n4648 & ~n4649 ;
  assign n4652 = n4650 & n4651 ;
  assign n4653 = n2992 & ~n4652 ;
  assign n4645 = ~n2991 & n4352 ;
  assign n4654 = n2808 & ~n4645 ;
  assign n4655 = ~n4653 & n4654 ;
  assign n4644 = ~\u7_dout_reg[2]/P0001  & ~n2808 ;
  assign n4656 = \u13_occ1_r_reg[0]/NET0131  & ~n4644 ;
  assign n4657 = ~n4655 & n4656 ;
  assign n4667 = ~n3004 & n4352 ;
  assign n4659 = \u7_mem_reg[1][3]/NET0131  & n2985 ;
  assign n4660 = \u7_mem_reg[3][3]/NET0131  & n2981 ;
  assign n4663 = ~n4659 & ~n4660 ;
  assign n4661 = \u7_mem_reg[2][3]/NET0131  & n2983 ;
  assign n4662 = \u7_mem_reg[0][3]/NET0131  & n2987 ;
  assign n4664 = ~n4661 & ~n4662 ;
  assign n4665 = n4663 & n4664 ;
  assign n4666 = n2992 & ~n4665 ;
  assign n4668 = n2808 & ~n4666 ;
  assign n4669 = ~n4667 & n4668 ;
  assign n4658 = ~\u7_dout_reg[3]/P0001  & ~n2808 ;
  assign n4670 = \u13_occ1_r_reg[0]/NET0131  & ~n4658 ;
  assign n4671 = ~n4669 & n4670 ;
  assign n4674 = \u7_rp_reg[0]/P0001  & n4558 ;
  assign n4673 = ~\u7_rp_reg[0]/P0001  & n2991 ;
  assign n4675 = n2805 & ~n4673 ;
  assign n4676 = ~n4674 & n4675 ;
  assign n4685 = n4352 & ~n4652 ;
  assign n4677 = \u7_mem_reg[1][4]/NET0131  & n2985 ;
  assign n4678 = \u7_mem_reg[2][4]/NET0131  & n2983 ;
  assign n4681 = ~n4677 & ~n4678 ;
  assign n4679 = \u7_mem_reg[3][4]/NET0131  & n2981 ;
  assign n4680 = \u7_mem_reg[0][4]/NET0131  & n2987 ;
  assign n4682 = ~n4679 & ~n4680 ;
  assign n4683 = n4681 & n4682 ;
  assign n4684 = n2992 & ~n4683 ;
  assign n4686 = n2808 & ~n4684 ;
  assign n4687 = ~n4685 & n4686 ;
  assign n4688 = ~n4676 & n4687 ;
  assign n4672 = ~\u7_dout_reg[4]/P0001  & ~n2808 ;
  assign n4689 = \u13_occ1_r_reg[0]/NET0131  & ~n4672 ;
  assign n4690 = ~n4688 & n4689 ;
  assign n4693 = \u7_rp_reg[0]/P0001  & n4584 ;
  assign n4692 = ~\u7_rp_reg[0]/P0001  & n3004 ;
  assign n4694 = n2805 & ~n4692 ;
  assign n4695 = ~n4693 & n4694 ;
  assign n4704 = n4352 & ~n4665 ;
  assign n4696 = \u7_mem_reg[3][5]/NET0131  & n2981 ;
  assign n4697 = \u7_mem_reg[0][5]/NET0131  & n2987 ;
  assign n4700 = ~n4696 & ~n4697 ;
  assign n4698 = \u7_mem_reg[2][5]/NET0131  & n2983 ;
  assign n4699 = \u7_mem_reg[1][5]/NET0131  & n2985 ;
  assign n4701 = ~n4698 & ~n4699 ;
  assign n4702 = n4700 & n4701 ;
  assign n4703 = n2992 & ~n4702 ;
  assign n4705 = n2808 & ~n4703 ;
  assign n4706 = ~n4704 & n4705 ;
  assign n4707 = ~n4695 & n4706 ;
  assign n4691 = ~\u7_dout_reg[5]/P0001  & ~n2808 ;
  assign n4708 = \u13_occ1_r_reg[0]/NET0131  & ~n4691 ;
  assign n4709 = ~n4707 & n4708 ;
  assign n4714 = \u7_rp_reg[0]/P0001  & n4610 ;
  assign n4713 = ~\u7_rp_reg[0]/P0001  & n4652 ;
  assign n4715 = n2805 & ~n4713 ;
  assign n4716 = ~n4714 & n4715 ;
  assign n4712 = n4352 & ~n4683 ;
  assign n4711 = n2992 & ~n4350 ;
  assign n4717 = n2808 & ~n4711 ;
  assign n4718 = ~n4712 & n4717 ;
  assign n4719 = ~n4716 & n4718 ;
  assign n4710 = ~\u7_dout_reg[6]/P0001  & ~n2808 ;
  assign n4720 = \u13_occ1_r_reg[0]/NET0131  & ~n4710 ;
  assign n4721 = ~n4719 & n4720 ;
  assign n4726 = \u7_rp_reg[0]/P0001  & n4636 ;
  assign n4725 = ~\u7_rp_reg[0]/P0001  & n4665 ;
  assign n4727 = n2805 & ~n4725 ;
  assign n4728 = ~n4726 & n4727 ;
  assign n4724 = n4352 & ~n4702 ;
  assign n4723 = n2992 & ~n4399 ;
  assign n4729 = n2808 & ~n4723 ;
  assign n4730 = ~n4724 & n4729 ;
  assign n4731 = ~n4728 & n4730 ;
  assign n4722 = ~\u7_dout_reg[7]/P0001  & ~n2808 ;
  assign n4732 = \u13_occ1_r_reg[0]/NET0131  & ~n4722 ;
  assign n4733 = ~n4731 & n4732 ;
  assign n4738 = \u7_mem_reg[2][20]/NET0131  & n2983 ;
  assign n4742 = \u7_rp_reg[0]/P0001  & ~n4738 ;
  assign n4741 = \u7_mem_reg[0][20]/NET0131  & n2987 ;
  assign n4739 = \u7_mem_reg[3][20]/NET0131  & n2981 ;
  assign n4740 = \u7_mem_reg[1][20]/NET0131  & n2985 ;
  assign n4743 = ~n4739 & ~n4740 ;
  assign n4744 = ~n4741 & n4743 ;
  assign n4745 = n4742 & n4744 ;
  assign n4737 = ~\u7_rp_reg[0]/P0001  & n4683 ;
  assign n4746 = n2805 & ~n4737 ;
  assign n4747 = ~n4745 & n4746 ;
  assign n4736 = n2992 & ~n4359 ;
  assign n4735 = ~n4350 & n4352 ;
  assign n4748 = n2808 & ~n4735 ;
  assign n4749 = ~n4736 & n4748 ;
  assign n4750 = ~n4747 & n4749 ;
  assign n4734 = ~\u7_dout_reg[8]/P0001  & ~n2808 ;
  assign n4751 = \u13_occ1_r_reg[0]/NET0131  & ~n4734 ;
  assign n4752 = ~n4750 & n4751 ;
  assign n4757 = \u7_mem_reg[2][21]/NET0131  & n2983 ;
  assign n4761 = \u7_rp_reg[0]/P0001  & ~n4757 ;
  assign n4760 = \u7_mem_reg[0][21]/NET0131  & n2987 ;
  assign n4758 = \u7_mem_reg[3][21]/NET0131  & n2981 ;
  assign n4759 = \u7_mem_reg[1][21]/NET0131  & n2985 ;
  assign n4762 = ~n4758 & ~n4759 ;
  assign n4763 = ~n4760 & n4762 ;
  assign n4764 = n4761 & n4763 ;
  assign n4756 = ~\u7_rp_reg[0]/P0001  & n4702 ;
  assign n4765 = n2805 & ~n4756 ;
  assign n4766 = ~n4764 & n4765 ;
  assign n4755 = n2992 & ~n4415 ;
  assign n4754 = n4352 & ~n4399 ;
  assign n4767 = n2808 & ~n4754 ;
  assign n4768 = ~n4755 & n4767 ;
  assign n4769 = ~n4766 & n4768 ;
  assign n4753 = ~\u7_dout_reg[9]/P0001  & ~n2808 ;
  assign n4770 = \u13_occ1_r_reg[0]/NET0131  & ~n4753 ;
  assign n4771 = ~n4769 & n4770 ;
  assign n4781 = \u3_mem_reg[2][22]/NET0131  & n3011 ;
  assign n4785 = \u3_rp_reg[0]/P0001  & ~n4781 ;
  assign n4784 = \u3_mem_reg[0][22]/NET0131  & n3015 ;
  assign n4782 = \u3_mem_reg[3][22]/NET0131  & n3009 ;
  assign n4783 = \u3_mem_reg[1][22]/NET0131  & n3013 ;
  assign n4786 = ~n4782 & ~n4783 ;
  assign n4787 = ~n4784 & n4786 ;
  assign n4788 = n4785 & n4787 ;
  assign n4773 = \u3_mem_reg[3][6]/NET0131  & n3009 ;
  assign n4774 = \u3_mem_reg[2][6]/NET0131  & n3011 ;
  assign n4777 = ~n4773 & ~n4774 ;
  assign n4775 = \u3_mem_reg[1][6]/NET0131  & n3013 ;
  assign n4776 = \u3_mem_reg[0][6]/NET0131  & n3015 ;
  assign n4778 = ~n4775 & ~n4776 ;
  assign n4779 = n4777 & n4778 ;
  assign n4780 = ~\u3_rp_reg[0]/P0001  & n4779 ;
  assign n4789 = n2784 & ~n4780 ;
  assign n4790 = ~n4788 & n4789 ;
  assign n4799 = \u13_occ0_r_reg[2]/NET0131  & ~\u13_occ0_r_reg[3]/NET0131  ;
  assign n4800 = \u3_mem_reg[3][8]/NET0131  & n3009 ;
  assign n4801 = \u3_mem_reg[2][8]/NET0131  & n3011 ;
  assign n4804 = ~n4800 & ~n4801 ;
  assign n4802 = \u3_mem_reg[1][8]/NET0131  & n3013 ;
  assign n4803 = \u3_mem_reg[0][8]/NET0131  & n3015 ;
  assign n4805 = ~n4802 & ~n4803 ;
  assign n4806 = n4804 & n4805 ;
  assign n4807 = n4799 & ~n4806 ;
  assign n4791 = \u3_mem_reg[3][10]/NET0131  & n3009 ;
  assign n4792 = \u3_mem_reg[2][10]/NET0131  & n3011 ;
  assign n4795 = ~n4791 & ~n4792 ;
  assign n4793 = \u3_mem_reg[0][10]/NET0131  & n3015 ;
  assign n4794 = \u3_mem_reg[1][10]/NET0131  & n3013 ;
  assign n4796 = ~n4793 & ~n4794 ;
  assign n4797 = n4795 & n4796 ;
  assign n4798 = n3020 & ~n4797 ;
  assign n4808 = n2787 & ~n4798 ;
  assign n4809 = ~n4807 & n4808 ;
  assign n4810 = ~n4790 & n4809 ;
  assign n4772 = ~\u3_dout_reg[10]/P0001  & ~n2787 ;
  assign n4811 = \u13_occ0_r_reg[0]/NET0131  & ~n4772 ;
  assign n4812 = ~n4810 & n4811 ;
  assign n4814 = \u3_mem_reg[2][9]/NET0131  & n3011 ;
  assign n4815 = \u3_mem_reg[3][9]/NET0131  & n3009 ;
  assign n4818 = ~n4814 & ~n4815 ;
  assign n4816 = \u3_mem_reg[1][9]/NET0131  & n3013 ;
  assign n4817 = \u3_mem_reg[0][9]/NET0131  & n3015 ;
  assign n4819 = ~n4816 & ~n4817 ;
  assign n4820 = n4818 & n4819 ;
  assign n4821 = n4799 & ~n4820 ;
  assign n4847 = n2787 & ~n4821 ;
  assign n4838 = \u3_rp_reg[0]/P0001  & n2784 ;
  assign n4839 = \u3_mem_reg[2][23]/NET0131  & n3011 ;
  assign n4840 = \u3_mem_reg[0][23]/NET0131  & n3015 ;
  assign n4843 = ~n4839 & ~n4840 ;
  assign n4841 = \u3_mem_reg[3][23]/NET0131  & n3009 ;
  assign n4842 = \u3_mem_reg[1][23]/NET0131  & n3013 ;
  assign n4844 = ~n4841 & ~n4842 ;
  assign n4845 = n4843 & n4844 ;
  assign n4846 = n4838 & ~n4845 ;
  assign n4822 = \u3_mem_reg[3][11]/NET0131  & n3009 ;
  assign n4823 = \u3_mem_reg[2][11]/NET0131  & n3011 ;
  assign n4826 = ~n4822 & ~n4823 ;
  assign n4824 = \u3_mem_reg[0][11]/NET0131  & n3015 ;
  assign n4825 = \u3_mem_reg[1][11]/NET0131  & n3013 ;
  assign n4827 = ~n4824 & ~n4825 ;
  assign n4828 = n4826 & n4827 ;
  assign n4829 = n3020 & ~n4828 ;
  assign n4830 = \u3_mem_reg[2][7]/NET0131  & n3011 ;
  assign n4831 = \u3_mem_reg[0][7]/NET0131  & n3015 ;
  assign n4834 = ~n4830 & ~n4831 ;
  assign n4832 = \u3_mem_reg[3][7]/NET0131  & n3009 ;
  assign n4833 = \u3_mem_reg[1][7]/NET0131  & n3013 ;
  assign n4835 = ~n4832 & ~n4833 ;
  assign n4836 = n4834 & n4835 ;
  assign n4837 = n2785 & ~n4836 ;
  assign n4848 = ~n4829 & ~n4837 ;
  assign n4849 = ~n4846 & n4848 ;
  assign n4850 = n4847 & n4849 ;
  assign n4813 = ~\u3_dout_reg[11]/P0001  & ~n2787 ;
  assign n4851 = \u13_occ0_r_reg[0]/NET0131  & ~n4813 ;
  assign n4852 = ~n4850 & n4851 ;
  assign n4855 = \u3_mem_reg[2][24]/NET0131  & n3011 ;
  assign n4859 = \u3_rp_reg[0]/P0001  & ~n4855 ;
  assign n4858 = \u3_mem_reg[0][24]/NET0131  & n3015 ;
  assign n4856 = \u3_mem_reg[3][24]/NET0131  & n3009 ;
  assign n4857 = \u3_mem_reg[1][24]/NET0131  & n3013 ;
  assign n4860 = ~n4856 & ~n4857 ;
  assign n4861 = ~n4858 & n4860 ;
  assign n4862 = n4859 & n4861 ;
  assign n4854 = ~\u3_rp_reg[0]/P0001  & n4806 ;
  assign n4863 = n2784 & ~n4854 ;
  assign n4864 = ~n4862 & n4863 ;
  assign n4873 = ~n4797 & n4799 ;
  assign n4865 = \u3_mem_reg[2][12]/NET0131  & n3011 ;
  assign n4866 = \u3_mem_reg[3][12]/NET0131  & n3009 ;
  assign n4869 = ~n4865 & ~n4866 ;
  assign n4867 = \u3_mem_reg[1][12]/NET0131  & n3013 ;
  assign n4868 = \u3_mem_reg[0][12]/NET0131  & n3015 ;
  assign n4870 = ~n4867 & ~n4868 ;
  assign n4871 = n4869 & n4870 ;
  assign n4872 = n3020 & ~n4871 ;
  assign n4874 = n2787 & ~n4872 ;
  assign n4875 = ~n4873 & n4874 ;
  assign n4876 = ~n4864 & n4875 ;
  assign n4853 = ~\u3_dout_reg[12]/P0001  & ~n2787 ;
  assign n4877 = \u13_occ0_r_reg[0]/NET0131  & ~n4853 ;
  assign n4878 = ~n4876 & n4877 ;
  assign n4880 = n2785 & ~n4820 ;
  assign n4898 = n2787 & ~n4880 ;
  assign n4897 = n4799 & ~n4828 ;
  assign n4881 = \u3_mem_reg[3][13]/NET0131  & n3009 ;
  assign n4882 = \u3_mem_reg[1][13]/NET0131  & n3013 ;
  assign n4885 = ~n4881 & ~n4882 ;
  assign n4883 = \u3_mem_reg[2][13]/NET0131  & n3011 ;
  assign n4884 = \u3_mem_reg[0][13]/NET0131  & n3015 ;
  assign n4886 = ~n4883 & ~n4884 ;
  assign n4887 = n4885 & n4886 ;
  assign n4888 = n3020 & ~n4887 ;
  assign n4889 = \u3_mem_reg[3][25]/NET0131  & n3009 ;
  assign n4890 = \u3_mem_reg[1][25]/NET0131  & n3013 ;
  assign n4893 = ~n4889 & ~n4890 ;
  assign n4891 = \u3_mem_reg[0][25]/NET0131  & n3015 ;
  assign n4892 = \u3_mem_reg[2][25]/NET0131  & n3011 ;
  assign n4894 = ~n4891 & ~n4892 ;
  assign n4895 = n4893 & n4894 ;
  assign n4896 = n4838 & ~n4895 ;
  assign n4899 = ~n4888 & ~n4896 ;
  assign n4900 = ~n4897 & n4899 ;
  assign n4901 = n4898 & n4900 ;
  assign n4879 = ~\u3_dout_reg[13]/P0001  & ~n2787 ;
  assign n4902 = \u13_occ0_r_reg[0]/NET0131  & ~n4879 ;
  assign n4903 = ~n4901 & n4902 ;
  assign n4906 = \u3_mem_reg[2][26]/NET0131  & n3011 ;
  assign n4910 = \u3_rp_reg[0]/P0001  & ~n4906 ;
  assign n4909 = \u3_mem_reg[0][26]/NET0131  & n3015 ;
  assign n4907 = \u3_mem_reg[3][26]/NET0131  & n3009 ;
  assign n4908 = \u3_mem_reg[1][26]/NET0131  & n3013 ;
  assign n4911 = ~n4907 & ~n4908 ;
  assign n4912 = ~n4909 & n4911 ;
  assign n4913 = n4910 & n4912 ;
  assign n4905 = ~\u3_rp_reg[0]/P0001  & n4797 ;
  assign n4914 = n2784 & ~n4905 ;
  assign n4915 = ~n4913 & n4914 ;
  assign n4924 = n4799 & ~n4871 ;
  assign n4916 = \u3_mem_reg[1][14]/NET0131  & n3013 ;
  assign n4917 = \u3_mem_reg[3][14]/NET0131  & n3009 ;
  assign n4920 = ~n4916 & ~n4917 ;
  assign n4918 = \u3_mem_reg[0][14]/NET0131  & n3015 ;
  assign n4919 = \u3_mem_reg[2][14]/NET0131  & n3011 ;
  assign n4921 = ~n4918 & ~n4919 ;
  assign n4922 = n4920 & n4921 ;
  assign n4923 = n3020 & ~n4922 ;
  assign n4925 = n2787 & ~n4923 ;
  assign n4926 = ~n4924 & n4925 ;
  assign n4927 = ~n4915 & n4926 ;
  assign n4904 = ~\u3_dout_reg[14]/P0001  & ~n2787 ;
  assign n4928 = \u13_occ0_r_reg[0]/NET0131  & ~n4904 ;
  assign n4929 = ~n4927 & n4928 ;
  assign n4941 = \u3_mem_reg[2][27]/NET0131  & n3011 ;
  assign n4945 = \u3_rp_reg[0]/P0001  & ~n4941 ;
  assign n4944 = \u3_mem_reg[0][27]/NET0131  & n3015 ;
  assign n4942 = \u3_mem_reg[3][27]/NET0131  & n3009 ;
  assign n4943 = \u3_mem_reg[1][27]/NET0131  & n3013 ;
  assign n4946 = ~n4942 & ~n4943 ;
  assign n4947 = ~n4944 & n4946 ;
  assign n4948 = n4945 & n4947 ;
  assign n4940 = ~\u3_rp_reg[0]/P0001  & n4828 ;
  assign n4949 = n2784 & ~n4940 ;
  assign n4950 = ~n4948 & n4949 ;
  assign n4932 = \u3_mem_reg[3][15]/NET0131  & n3009 ;
  assign n4933 = \u3_mem_reg[2][15]/NET0131  & n3011 ;
  assign n4936 = ~n4932 & ~n4933 ;
  assign n4934 = \u3_mem_reg[1][15]/NET0131  & n3013 ;
  assign n4935 = \u3_mem_reg[0][15]/NET0131  & n3015 ;
  assign n4937 = ~n4934 & ~n4935 ;
  assign n4938 = n4936 & n4937 ;
  assign n4939 = n3020 & ~n4938 ;
  assign n4931 = n4799 & ~n4887 ;
  assign n4951 = n2787 & ~n4931 ;
  assign n4952 = ~n4939 & n4951 ;
  assign n4953 = ~n4950 & n4952 ;
  assign n4930 = ~\u3_dout_reg[15]/P0001  & ~n2787 ;
  assign n4954 = \u13_occ0_r_reg[0]/NET0131  & ~n4930 ;
  assign n4955 = ~n4953 & n4954 ;
  assign n4958 = \u3_mem_reg[2][28]/NET0131  & n3011 ;
  assign n4962 = \u3_rp_reg[0]/P0001  & ~n4958 ;
  assign n4961 = \u3_mem_reg[0][28]/NET0131  & n3015 ;
  assign n4959 = \u3_mem_reg[3][28]/NET0131  & n3009 ;
  assign n4960 = \u3_mem_reg[1][28]/NET0131  & n3013 ;
  assign n4963 = ~n4959 & ~n4960 ;
  assign n4964 = ~n4961 & n4963 ;
  assign n4965 = n4962 & n4964 ;
  assign n4957 = ~\u3_rp_reg[0]/P0001  & n4871 ;
  assign n4966 = n2784 & ~n4957 ;
  assign n4967 = ~n4965 & n4966 ;
  assign n4976 = n4799 & ~n4922 ;
  assign n4968 = \u3_mem_reg[3][16]/NET0131  & n3009 ;
  assign n4969 = \u3_mem_reg[2][16]/NET0131  & n3011 ;
  assign n4972 = ~n4968 & ~n4969 ;
  assign n4970 = \u3_mem_reg[1][16]/NET0131  & n3013 ;
  assign n4971 = \u3_mem_reg[0][16]/NET0131  & n3015 ;
  assign n4973 = ~n4970 & ~n4971 ;
  assign n4974 = n4972 & n4973 ;
  assign n4975 = n3020 & ~n4974 ;
  assign n4977 = n2787 & ~n4975 ;
  assign n4978 = ~n4976 & n4977 ;
  assign n4979 = ~n4967 & n4978 ;
  assign n4956 = ~\u3_dout_reg[16]/P0001  & ~n2787 ;
  assign n4980 = \u13_occ0_r_reg[0]/NET0131  & ~n4956 ;
  assign n4981 = ~n4979 & n4980 ;
  assign n4983 = n4799 & ~n4938 ;
  assign n5001 = n2787 & ~n4983 ;
  assign n4993 = \u3_mem_reg[1][17]/NET0131  & n3013 ;
  assign n4994 = \u3_mem_reg[3][17]/NET0131  & n3009 ;
  assign n4997 = ~n4993 & ~n4994 ;
  assign n4995 = \u3_mem_reg[2][17]/NET0131  & n3011 ;
  assign n4996 = \u3_mem_reg[0][17]/NET0131  & n3015 ;
  assign n4998 = ~n4995 & ~n4996 ;
  assign n4999 = n4997 & n4998 ;
  assign n5000 = n3020 & ~n4999 ;
  assign n4984 = n2785 & ~n4887 ;
  assign n4985 = \u3_mem_reg[3][29]/NET0131  & n3009 ;
  assign n4986 = \u3_mem_reg[0][29]/NET0131  & n3015 ;
  assign n4989 = ~n4985 & ~n4986 ;
  assign n4987 = \u3_mem_reg[2][29]/NET0131  & n3011 ;
  assign n4988 = \u3_mem_reg[1][29]/NET0131  & n3013 ;
  assign n4990 = ~n4987 & ~n4988 ;
  assign n4991 = n4989 & n4990 ;
  assign n4992 = n4838 & ~n4991 ;
  assign n5002 = ~n4984 & ~n4992 ;
  assign n5003 = ~n5000 & n5002 ;
  assign n5004 = n5001 & n5003 ;
  assign n4982 = ~\u3_dout_reg[17]/P0001  & ~n2787 ;
  assign n5005 = \u13_occ0_r_reg[0]/NET0131  & ~n4982 ;
  assign n5006 = ~n5004 & n5005 ;
  assign n5009 = \u3_mem_reg[2][30]/NET0131  & n3011 ;
  assign n5013 = \u3_rp_reg[0]/P0001  & ~n5009 ;
  assign n5012 = \u3_mem_reg[0][30]/NET0131  & n3015 ;
  assign n5010 = \u3_mem_reg[3][30]/NET0131  & n3009 ;
  assign n5011 = \u3_mem_reg[1][30]/NET0131  & n3013 ;
  assign n5014 = ~n5010 & ~n5011 ;
  assign n5015 = ~n5012 & n5014 ;
  assign n5016 = n5013 & n5015 ;
  assign n5008 = ~\u3_rp_reg[0]/P0001  & n4922 ;
  assign n5017 = n2784 & ~n5008 ;
  assign n5018 = ~n5016 & n5017 ;
  assign n5027 = n4799 & ~n4974 ;
  assign n5019 = \u3_mem_reg[1][18]/NET0131  & n3013 ;
  assign n5020 = \u3_mem_reg[3][18]/NET0131  & n3009 ;
  assign n5023 = ~n5019 & ~n5020 ;
  assign n5021 = \u3_mem_reg[2][18]/NET0131  & n3011 ;
  assign n5022 = \u3_mem_reg[0][18]/NET0131  & n3015 ;
  assign n5024 = ~n5021 & ~n5022 ;
  assign n5025 = n5023 & n5024 ;
  assign n5026 = n3020 & ~n5025 ;
  assign n5028 = n2787 & ~n5026 ;
  assign n5029 = ~n5027 & n5028 ;
  assign n5030 = ~n5018 & n5029 ;
  assign n5007 = ~\u3_dout_reg[18]/P0001  & ~n2787 ;
  assign n5031 = \u13_occ0_r_reg[0]/NET0131  & ~n5007 ;
  assign n5032 = ~n5030 & n5031 ;
  assign n5042 = \u8_mem_reg[2][22]/NET0131  & n3028 ;
  assign n5046 = \u8_rp_reg[0]/P0001  & ~n5042 ;
  assign n5045 = \u8_mem_reg[0][22]/NET0131  & n3032 ;
  assign n5043 = \u8_mem_reg[3][22]/NET0131  & n2163 ;
  assign n5044 = \u8_mem_reg[1][22]/NET0131  & n3030 ;
  assign n5047 = ~n5043 & ~n5044 ;
  assign n5048 = ~n5045 & n5047 ;
  assign n5049 = n5046 & n5048 ;
  assign n5034 = \u8_mem_reg[3][6]/NET0131  & n2163 ;
  assign n5035 = \u8_mem_reg[2][6]/NET0131  & n3028 ;
  assign n5038 = ~n5034 & ~n5035 ;
  assign n5036 = \u8_mem_reg[0][6]/NET0131  & n3032 ;
  assign n5037 = \u8_mem_reg[1][6]/NET0131  & n3030 ;
  assign n5039 = ~n5036 & ~n5037 ;
  assign n5040 = n5038 & n5039 ;
  assign n5041 = ~\u8_rp_reg[0]/P0001  & n5040 ;
  assign n5050 = n2160 & ~n5041 ;
  assign n5051 = ~n5049 & n5050 ;
  assign n5060 = \u13_occ1_r_reg[10]/NET0131  & ~\u13_occ1_r_reg[11]/NET0131  ;
  assign n5061 = \u8_mem_reg[3][8]/NET0131  & n2163 ;
  assign n5062 = \u8_mem_reg[2][8]/NET0131  & n3028 ;
  assign n5065 = ~n5061 & ~n5062 ;
  assign n5063 = \u8_mem_reg[0][8]/NET0131  & n3032 ;
  assign n5064 = \u8_mem_reg[1][8]/NET0131  & n3030 ;
  assign n5066 = ~n5063 & ~n5064 ;
  assign n5067 = n5065 & n5066 ;
  assign n5068 = n5060 & ~n5067 ;
  assign n5052 = \u8_mem_reg[3][10]/NET0131  & n2163 ;
  assign n5053 = \u8_mem_reg[2][10]/NET0131  & n3028 ;
  assign n5056 = ~n5052 & ~n5053 ;
  assign n5054 = \u8_mem_reg[0][10]/NET0131  & n3032 ;
  assign n5055 = \u8_mem_reg[1][10]/NET0131  & n3030 ;
  assign n5057 = ~n5054 & ~n5055 ;
  assign n5058 = n5056 & n5057 ;
  assign n5059 = n3037 & ~n5058 ;
  assign n5069 = n2159 & ~n5059 ;
  assign n5070 = ~n5068 & n5069 ;
  assign n5071 = ~n5051 & n5070 ;
  assign n5033 = ~\u8_dout_reg[10]/P0001  & ~n2159 ;
  assign n5072 = \u13_occ1_r_reg[8]/NET0131  & ~n5033 ;
  assign n5073 = ~n5071 & n5072 ;
  assign n5076 = \u3_mem_reg[2][31]/NET0131  & n3011 ;
  assign n5080 = \u3_rp_reg[0]/P0001  & ~n5076 ;
  assign n5079 = \u3_mem_reg[0][31]/NET0131  & n3015 ;
  assign n5077 = \u3_mem_reg[3][31]/NET0131  & n3009 ;
  assign n5078 = \u3_mem_reg[1][31]/NET0131  & n3013 ;
  assign n5081 = ~n5077 & ~n5078 ;
  assign n5082 = ~n5079 & n5081 ;
  assign n5083 = n5080 & n5082 ;
  assign n5075 = ~\u3_rp_reg[0]/P0001  & n4938 ;
  assign n5084 = n2784 & ~n5075 ;
  assign n5085 = ~n5083 & n5084 ;
  assign n5094 = n4799 & ~n4999 ;
  assign n5086 = \u3_mem_reg[2][19]/NET0131  & n3011 ;
  assign n5087 = \u3_mem_reg[0][19]/NET0131  & n3015 ;
  assign n5090 = ~n5086 & ~n5087 ;
  assign n5088 = \u3_mem_reg[1][19]/NET0131  & n3013 ;
  assign n5089 = \u3_mem_reg[3][19]/NET0131  & n3009 ;
  assign n5091 = ~n5088 & ~n5089 ;
  assign n5092 = n5090 & n5091 ;
  assign n5093 = n3020 & ~n5092 ;
  assign n5095 = n2787 & ~n5093 ;
  assign n5096 = ~n5094 & n5095 ;
  assign n5097 = ~n5085 & n5096 ;
  assign n5074 = ~\u3_dout_reg[19]/P0001  & ~n2787 ;
  assign n5098 = \u13_occ0_r_reg[0]/NET0131  & ~n5074 ;
  assign n5099 = ~n5097 & n5098 ;
  assign n5109 = \u8_mem_reg[2][23]/NET0131  & n3028 ;
  assign n5113 = \u8_rp_reg[0]/P0001  & ~n5109 ;
  assign n5112 = \u8_mem_reg[0][23]/NET0131  & n3032 ;
  assign n5110 = \u8_mem_reg[3][23]/NET0131  & n2163 ;
  assign n5111 = \u8_mem_reg[1][23]/NET0131  & n3030 ;
  assign n5114 = ~n5110 & ~n5111 ;
  assign n5115 = ~n5112 & n5114 ;
  assign n5116 = n5113 & n5115 ;
  assign n5101 = \u8_mem_reg[3][7]/NET0131  & n2163 ;
  assign n5102 = \u8_mem_reg[2][7]/NET0131  & n3028 ;
  assign n5105 = ~n5101 & ~n5102 ;
  assign n5103 = \u8_mem_reg[0][7]/NET0131  & n3032 ;
  assign n5104 = \u8_mem_reg[1][7]/NET0131  & n3030 ;
  assign n5106 = ~n5103 & ~n5104 ;
  assign n5107 = n5105 & n5106 ;
  assign n5108 = ~\u8_rp_reg[0]/P0001  & n5107 ;
  assign n5117 = n2160 & ~n5108 ;
  assign n5118 = ~n5116 & n5117 ;
  assign n5127 = \u8_mem_reg[3][9]/NET0131  & n2163 ;
  assign n5128 = \u8_mem_reg[1][9]/NET0131  & n3030 ;
  assign n5131 = ~n5127 & ~n5128 ;
  assign n5129 = \u8_mem_reg[0][9]/NET0131  & n3032 ;
  assign n5130 = \u8_mem_reg[2][9]/NET0131  & n3028 ;
  assign n5132 = ~n5129 & ~n5130 ;
  assign n5133 = n5131 & n5132 ;
  assign n5134 = n5060 & ~n5133 ;
  assign n5119 = \u8_mem_reg[3][11]/NET0131  & n2163 ;
  assign n5120 = \u8_mem_reg[2][11]/NET0131  & n3028 ;
  assign n5123 = ~n5119 & ~n5120 ;
  assign n5121 = \u8_mem_reg[0][11]/NET0131  & n3032 ;
  assign n5122 = \u8_mem_reg[1][11]/NET0131  & n3030 ;
  assign n5124 = ~n5121 & ~n5122 ;
  assign n5125 = n5123 & n5124 ;
  assign n5126 = n3037 & ~n5125 ;
  assign n5135 = n2159 & ~n5126 ;
  assign n5136 = ~n5134 & n5135 ;
  assign n5137 = ~n5118 & n5136 ;
  assign n5100 = ~\u8_dout_reg[11]/P0001  & ~n2159 ;
  assign n5138 = \u13_occ1_r_reg[8]/NET0131  & ~n5100 ;
  assign n5139 = ~n5137 & n5138 ;
  assign n5142 = \u8_mem_reg[2][24]/NET0131  & n3028 ;
  assign n5146 = \u8_rp_reg[0]/P0001  & ~n5142 ;
  assign n5145 = \u8_mem_reg[0][24]/NET0131  & n3032 ;
  assign n5143 = \u8_mem_reg[3][24]/NET0131  & n2163 ;
  assign n5144 = \u8_mem_reg[1][24]/NET0131  & n3030 ;
  assign n5147 = ~n5143 & ~n5144 ;
  assign n5148 = ~n5145 & n5147 ;
  assign n5149 = n5146 & n5148 ;
  assign n5141 = ~\u8_rp_reg[0]/P0001  & n5067 ;
  assign n5150 = n2160 & ~n5141 ;
  assign n5151 = ~n5149 & n5150 ;
  assign n5160 = ~n5058 & n5060 ;
  assign n5152 = \u8_mem_reg[3][12]/NET0131  & n2163 ;
  assign n5153 = \u8_mem_reg[1][12]/NET0131  & n3030 ;
  assign n5156 = ~n5152 & ~n5153 ;
  assign n5154 = \u8_mem_reg[0][12]/NET0131  & n3032 ;
  assign n5155 = \u8_mem_reg[2][12]/NET0131  & n3028 ;
  assign n5157 = ~n5154 & ~n5155 ;
  assign n5158 = n5156 & n5157 ;
  assign n5159 = n3037 & ~n5158 ;
  assign n5161 = n2159 & ~n5159 ;
  assign n5162 = ~n5160 & n5161 ;
  assign n5163 = ~n5151 & n5162 ;
  assign n5140 = ~\u8_dout_reg[12]/P0001  & ~n2159 ;
  assign n5164 = \u13_occ1_r_reg[8]/NET0131  & ~n5140 ;
  assign n5165 = ~n5163 & n5164 ;
  assign n5168 = \u3_mem_reg[3][2]/NET0131  & n3009 ;
  assign n5169 = \u3_mem_reg[2][2]/NET0131  & n3011 ;
  assign n5172 = ~n5168 & ~n5169 ;
  assign n5170 = \u3_mem_reg[1][2]/NET0131  & n3013 ;
  assign n5171 = \u3_mem_reg[0][2]/NET0131  & n3015 ;
  assign n5173 = ~n5170 & ~n5171 ;
  assign n5174 = n5172 & n5173 ;
  assign n5175 = n3020 & ~n5174 ;
  assign n5167 = ~n3019 & n4799 ;
  assign n5176 = n2787 & ~n5167 ;
  assign n5177 = ~n5175 & n5176 ;
  assign n5166 = ~\u3_dout_reg[2]/P0001  & ~n2787 ;
  assign n5178 = \u13_occ0_r_reg[0]/NET0131  & ~n5166 ;
  assign n5179 = ~n5177 & n5178 ;
  assign n5182 = \u8_mem_reg[2][25]/NET0131  & n3028 ;
  assign n5186 = \u8_rp_reg[0]/P0001  & ~n5182 ;
  assign n5185 = \u8_mem_reg[0][25]/NET0131  & n3032 ;
  assign n5183 = \u8_mem_reg[3][25]/NET0131  & n2163 ;
  assign n5184 = \u8_mem_reg[1][25]/NET0131  & n3030 ;
  assign n5187 = ~n5183 & ~n5184 ;
  assign n5188 = ~n5185 & n5187 ;
  assign n5189 = n5186 & n5188 ;
  assign n5181 = ~\u8_rp_reg[0]/P0001  & n5133 ;
  assign n5190 = n2160 & ~n5181 ;
  assign n5191 = ~n5189 & n5190 ;
  assign n5200 = n5060 & ~n5125 ;
  assign n5192 = \u8_mem_reg[3][13]/NET0131  & n2163 ;
  assign n5193 = \u8_mem_reg[2][13]/NET0131  & n3028 ;
  assign n5196 = ~n5192 & ~n5193 ;
  assign n5194 = \u8_mem_reg[0][13]/NET0131  & n3032 ;
  assign n5195 = \u8_mem_reg[1][13]/NET0131  & n3030 ;
  assign n5197 = ~n5194 & ~n5195 ;
  assign n5198 = n5196 & n5197 ;
  assign n5199 = n3037 & ~n5198 ;
  assign n5201 = n2159 & ~n5199 ;
  assign n5202 = ~n5200 & n5201 ;
  assign n5203 = ~n5191 & n5202 ;
  assign n5180 = ~\u8_dout_reg[13]/P0001  & ~n2159 ;
  assign n5204 = \u13_occ1_r_reg[8]/NET0131  & ~n5180 ;
  assign n5205 = ~n5203 & n5204 ;
  assign n5208 = \u3_mem_reg[1][3]/NET0131  & n3013 ;
  assign n5209 = \u3_mem_reg[3][3]/NET0131  & n3009 ;
  assign n5212 = ~n5208 & ~n5209 ;
  assign n5210 = \u3_mem_reg[2][3]/NET0131  & n3011 ;
  assign n5211 = \u3_mem_reg[0][3]/NET0131  & n3015 ;
  assign n5213 = ~n5210 & ~n5211 ;
  assign n5214 = n5212 & n5213 ;
  assign n5215 = n3020 & ~n5214 ;
  assign n5207 = ~n3049 & n4799 ;
  assign n5216 = n2787 & ~n5207 ;
  assign n5217 = ~n5215 & n5216 ;
  assign n5206 = ~\u3_dout_reg[3]/P0001  & ~n2787 ;
  assign n5218 = \u13_occ0_r_reg[0]/NET0131  & ~n5206 ;
  assign n5219 = ~n5217 & n5218 ;
  assign n5222 = \u8_mem_reg[2][26]/NET0131  & n3028 ;
  assign n5226 = \u8_rp_reg[0]/P0001  & ~n5222 ;
  assign n5225 = \u8_mem_reg[0][26]/NET0131  & n3032 ;
  assign n5223 = \u8_mem_reg[3][26]/NET0131  & n2163 ;
  assign n5224 = \u8_mem_reg[1][26]/NET0131  & n3030 ;
  assign n5227 = ~n5223 & ~n5224 ;
  assign n5228 = ~n5225 & n5227 ;
  assign n5229 = n5226 & n5228 ;
  assign n5221 = ~\u8_rp_reg[0]/P0001  & n5058 ;
  assign n5230 = n2160 & ~n5221 ;
  assign n5231 = ~n5229 & n5230 ;
  assign n5240 = n5060 & ~n5158 ;
  assign n5232 = \u8_mem_reg[3][14]/NET0131  & n2163 ;
  assign n5233 = \u8_mem_reg[2][14]/NET0131  & n3028 ;
  assign n5236 = ~n5232 & ~n5233 ;
  assign n5234 = \u8_mem_reg[0][14]/NET0131  & n3032 ;
  assign n5235 = \u8_mem_reg[1][14]/NET0131  & n3030 ;
  assign n5237 = ~n5234 & ~n5235 ;
  assign n5238 = n5236 & n5237 ;
  assign n5239 = n3037 & ~n5238 ;
  assign n5241 = n2159 & ~n5239 ;
  assign n5242 = ~n5240 & n5241 ;
  assign n5243 = ~n5231 & n5242 ;
  assign n5220 = ~\u8_dout_reg[14]/P0001  & ~n2159 ;
  assign n5244 = \u13_occ1_r_reg[8]/NET0131  & ~n5220 ;
  assign n5245 = ~n5243 & n5244 ;
  assign n5248 = \u3_rp_reg[0]/P0001  & n4974 ;
  assign n5247 = ~\u3_rp_reg[0]/P0001  & n3019 ;
  assign n5249 = n2784 & ~n5247 ;
  assign n5250 = ~n5248 & n5249 ;
  assign n5259 = n4799 & ~n5174 ;
  assign n5251 = \u3_mem_reg[3][4]/NET0131  & n3009 ;
  assign n5252 = \u3_mem_reg[2][4]/NET0131  & n3011 ;
  assign n5255 = ~n5251 & ~n5252 ;
  assign n5253 = \u3_mem_reg[0][4]/NET0131  & n3015 ;
  assign n5254 = \u3_mem_reg[1][4]/NET0131  & n3013 ;
  assign n5256 = ~n5253 & ~n5254 ;
  assign n5257 = n5255 & n5256 ;
  assign n5258 = n3020 & ~n5257 ;
  assign n5260 = n2787 & ~n5258 ;
  assign n5261 = ~n5259 & n5260 ;
  assign n5262 = ~n5250 & n5261 ;
  assign n5246 = ~\u3_dout_reg[4]/P0001  & ~n2787 ;
  assign n5263 = \u13_occ0_r_reg[0]/NET0131  & ~n5246 ;
  assign n5264 = ~n5262 & n5263 ;
  assign n5267 = \u8_mem_reg[2][27]/NET0131  & n3028 ;
  assign n5271 = \u8_rp_reg[0]/P0001  & ~n5267 ;
  assign n5270 = \u8_mem_reg[0][27]/NET0131  & n3032 ;
  assign n5268 = \u8_mem_reg[3][27]/NET0131  & n2163 ;
  assign n5269 = \u8_mem_reg[1][27]/NET0131  & n3030 ;
  assign n5272 = ~n5268 & ~n5269 ;
  assign n5273 = ~n5270 & n5272 ;
  assign n5274 = n5271 & n5273 ;
  assign n5266 = ~\u8_rp_reg[0]/P0001  & n5125 ;
  assign n5275 = n2160 & ~n5266 ;
  assign n5276 = ~n5274 & n5275 ;
  assign n5285 = n5060 & ~n5198 ;
  assign n5277 = \u8_mem_reg[3][15]/NET0131  & n2163 ;
  assign n5278 = \u8_mem_reg[2][15]/NET0131  & n3028 ;
  assign n5281 = ~n5277 & ~n5278 ;
  assign n5279 = \u8_mem_reg[0][15]/NET0131  & n3032 ;
  assign n5280 = \u8_mem_reg[1][15]/NET0131  & n3030 ;
  assign n5282 = ~n5279 & ~n5280 ;
  assign n5283 = n5281 & n5282 ;
  assign n5284 = n3037 & ~n5283 ;
  assign n5286 = n2159 & ~n5284 ;
  assign n5287 = ~n5285 & n5286 ;
  assign n5288 = ~n5276 & n5287 ;
  assign n5265 = ~\u8_dout_reg[15]/P0001  & ~n2159 ;
  assign n5289 = \u13_occ1_r_reg[8]/NET0131  & ~n5265 ;
  assign n5290 = ~n5288 & n5289 ;
  assign n5293 = \u3_rp_reg[0]/P0001  & n4999 ;
  assign n5292 = ~\u3_rp_reg[0]/P0001  & n3049 ;
  assign n5294 = n2784 & ~n5292 ;
  assign n5295 = ~n5293 & n5294 ;
  assign n5304 = n4799 & ~n5214 ;
  assign n5296 = \u3_mem_reg[3][5]/NET0131  & n3009 ;
  assign n5297 = \u3_mem_reg[2][5]/NET0131  & n3011 ;
  assign n5300 = ~n5296 & ~n5297 ;
  assign n5298 = \u3_mem_reg[1][5]/NET0131  & n3013 ;
  assign n5299 = \u3_mem_reg[0][5]/NET0131  & n3015 ;
  assign n5301 = ~n5298 & ~n5299 ;
  assign n5302 = n5300 & n5301 ;
  assign n5303 = n3020 & ~n5302 ;
  assign n5305 = n2787 & ~n5303 ;
  assign n5306 = ~n5304 & n5305 ;
  assign n5307 = ~n5295 & n5306 ;
  assign n5291 = ~\u3_dout_reg[5]/P0001  & ~n2787 ;
  assign n5308 = \u13_occ0_r_reg[0]/NET0131  & ~n5291 ;
  assign n5309 = ~n5307 & n5308 ;
  assign n5312 = \u8_mem_reg[2][28]/NET0131  & n3028 ;
  assign n5316 = \u8_rp_reg[0]/P0001  & ~n5312 ;
  assign n5315 = \u8_mem_reg[0][28]/NET0131  & n3032 ;
  assign n5313 = \u8_mem_reg[3][28]/NET0131  & n2163 ;
  assign n5314 = \u8_mem_reg[1][28]/NET0131  & n3030 ;
  assign n5317 = ~n5313 & ~n5314 ;
  assign n5318 = ~n5315 & n5317 ;
  assign n5319 = n5316 & n5318 ;
  assign n5311 = ~\u8_rp_reg[0]/P0001  & n5158 ;
  assign n5320 = n2160 & ~n5311 ;
  assign n5321 = ~n5319 & n5320 ;
  assign n5330 = n5060 & ~n5238 ;
  assign n5322 = \u8_mem_reg[2][16]/NET0131  & n3028 ;
  assign n5323 = \u8_mem_reg[0][16]/NET0131  & n3032 ;
  assign n5326 = ~n5322 & ~n5323 ;
  assign n5324 = \u8_mem_reg[1][16]/NET0131  & n3030 ;
  assign n5325 = \u8_mem_reg[3][16]/NET0131  & n2163 ;
  assign n5327 = ~n5324 & ~n5325 ;
  assign n5328 = n5326 & n5327 ;
  assign n5329 = n3037 & ~n5328 ;
  assign n5331 = n2159 & ~n5329 ;
  assign n5332 = ~n5330 & n5331 ;
  assign n5333 = ~n5321 & n5332 ;
  assign n5310 = ~\u8_dout_reg[16]/P0001  & ~n2159 ;
  assign n5334 = \u13_occ1_r_reg[8]/NET0131  & ~n5310 ;
  assign n5335 = ~n5333 & n5334 ;
  assign n5338 = \u8_mem_reg[2][29]/NET0131  & n3028 ;
  assign n5342 = \u8_rp_reg[0]/P0001  & ~n5338 ;
  assign n5341 = \u8_mem_reg[0][29]/NET0131  & n3032 ;
  assign n5339 = \u8_mem_reg[3][29]/NET0131  & n2163 ;
  assign n5340 = \u8_mem_reg[1][29]/NET0131  & n3030 ;
  assign n5343 = ~n5339 & ~n5340 ;
  assign n5344 = ~n5341 & n5343 ;
  assign n5345 = n5342 & n5344 ;
  assign n5337 = ~\u8_rp_reg[0]/P0001  & n5198 ;
  assign n5346 = n2160 & ~n5337 ;
  assign n5347 = ~n5345 & n5346 ;
  assign n5356 = n5060 & ~n5283 ;
  assign n5348 = \u8_mem_reg[3][17]/NET0131  & n2163 ;
  assign n5349 = \u8_mem_reg[2][17]/NET0131  & n3028 ;
  assign n5352 = ~n5348 & ~n5349 ;
  assign n5350 = \u8_mem_reg[0][17]/NET0131  & n3032 ;
  assign n5351 = \u8_mem_reg[1][17]/NET0131  & n3030 ;
  assign n5353 = ~n5350 & ~n5351 ;
  assign n5354 = n5352 & n5353 ;
  assign n5355 = n3037 & ~n5354 ;
  assign n5357 = n2159 & ~n5355 ;
  assign n5358 = ~n5356 & n5357 ;
  assign n5359 = ~n5347 & n5358 ;
  assign n5336 = ~\u8_dout_reg[17]/P0001  & ~n2159 ;
  assign n5360 = \u13_occ1_r_reg[8]/NET0131  & ~n5336 ;
  assign n5361 = ~n5359 & n5360 ;
  assign n5364 = \u3_rp_reg[0]/P0001  & n5025 ;
  assign n5363 = ~\u3_rp_reg[0]/P0001  & n5174 ;
  assign n5365 = n2784 & ~n5363 ;
  assign n5366 = ~n5364 & n5365 ;
  assign n5368 = n4799 & ~n5257 ;
  assign n5367 = n3020 & ~n4779 ;
  assign n5369 = n2787 & ~n5367 ;
  assign n5370 = ~n5368 & n5369 ;
  assign n5371 = ~n5366 & n5370 ;
  assign n5362 = ~\u3_dout_reg[6]/P0001  & ~n2787 ;
  assign n5372 = \u13_occ0_r_reg[0]/NET0131  & ~n5362 ;
  assign n5373 = ~n5371 & n5372 ;
  assign n5376 = \u3_rp_reg[0]/P0001  & n5092 ;
  assign n5375 = ~\u3_rp_reg[0]/P0001  & n5214 ;
  assign n5377 = n2784 & ~n5375 ;
  assign n5378 = ~n5376 & n5377 ;
  assign n5380 = n4799 & ~n5302 ;
  assign n5379 = n3020 & ~n4836 ;
  assign n5381 = n2787 & ~n5379 ;
  assign n5382 = ~n5380 & n5381 ;
  assign n5383 = ~n5378 & n5382 ;
  assign n5374 = ~\u3_dout_reg[7]/P0001  & ~n2787 ;
  assign n5384 = \u13_occ0_r_reg[0]/NET0131  & ~n5374 ;
  assign n5385 = ~n5383 & n5384 ;
  assign n5388 = \u8_mem_reg[2][30]/NET0131  & n3028 ;
  assign n5392 = \u8_rp_reg[0]/P0001  & ~n5388 ;
  assign n5391 = \u8_mem_reg[0][30]/NET0131  & n3032 ;
  assign n5389 = \u8_mem_reg[3][30]/NET0131  & n2163 ;
  assign n5390 = \u8_mem_reg[1][30]/NET0131  & n3030 ;
  assign n5393 = ~n5389 & ~n5390 ;
  assign n5394 = ~n5391 & n5393 ;
  assign n5395 = n5392 & n5394 ;
  assign n5387 = ~\u8_rp_reg[0]/P0001  & n5238 ;
  assign n5396 = n2160 & ~n5387 ;
  assign n5397 = ~n5395 & n5396 ;
  assign n5406 = n5060 & ~n5328 ;
  assign n5398 = \u8_mem_reg[2][18]/NET0131  & n3028 ;
  assign n5399 = \u8_mem_reg[3][18]/NET0131  & n2163 ;
  assign n5402 = ~n5398 & ~n5399 ;
  assign n5400 = \u8_mem_reg[1][18]/NET0131  & n3030 ;
  assign n5401 = \u8_mem_reg[0][18]/NET0131  & n3032 ;
  assign n5403 = ~n5400 & ~n5401 ;
  assign n5404 = n5402 & n5403 ;
  assign n5405 = n3037 & ~n5404 ;
  assign n5407 = n2159 & ~n5405 ;
  assign n5408 = ~n5406 & n5407 ;
  assign n5409 = ~n5397 & n5408 ;
  assign n5386 = ~\u8_dout_reg[18]/P0001  & ~n2159 ;
  assign n5410 = \u13_occ1_r_reg[8]/NET0131  & ~n5386 ;
  assign n5411 = ~n5409 & n5410 ;
  assign n5414 = \u3_mem_reg[2][20]/NET0131  & n3011 ;
  assign n5418 = \u3_rp_reg[0]/P0001  & ~n5414 ;
  assign n5417 = \u3_mem_reg[0][20]/NET0131  & n3015 ;
  assign n5415 = \u3_mem_reg[3][20]/NET0131  & n3009 ;
  assign n5416 = \u3_mem_reg[1][20]/NET0131  & n3013 ;
  assign n5419 = ~n5415 & ~n5416 ;
  assign n5420 = ~n5417 & n5419 ;
  assign n5421 = n5418 & n5420 ;
  assign n5413 = ~\u3_rp_reg[0]/P0001  & n5257 ;
  assign n5422 = n2784 & ~n5413 ;
  assign n5423 = ~n5421 & n5422 ;
  assign n5425 = ~n4779 & n4799 ;
  assign n5424 = n3020 & ~n4806 ;
  assign n5426 = n2787 & ~n5424 ;
  assign n5427 = ~n5425 & n5426 ;
  assign n5428 = ~n5423 & n5427 ;
  assign n5412 = ~\u3_dout_reg[8]/P0001  & ~n2787 ;
  assign n5429 = \u13_occ0_r_reg[0]/NET0131  & ~n5412 ;
  assign n5430 = ~n5428 & n5429 ;
  assign n5433 = \u8_mem_reg[2][31]/NET0131  & n3028 ;
  assign n5437 = \u8_rp_reg[0]/P0001  & ~n5433 ;
  assign n5436 = \u8_mem_reg[0][31]/NET0131  & n3032 ;
  assign n5434 = \u8_mem_reg[3][31]/NET0131  & n2163 ;
  assign n5435 = \u8_mem_reg[1][31]/NET0131  & n3030 ;
  assign n5438 = ~n5434 & ~n5435 ;
  assign n5439 = ~n5436 & n5438 ;
  assign n5440 = n5437 & n5439 ;
  assign n5432 = ~\u8_rp_reg[0]/P0001  & n5283 ;
  assign n5441 = n2160 & ~n5432 ;
  assign n5442 = ~n5440 & n5441 ;
  assign n5451 = n5060 & ~n5354 ;
  assign n5443 = \u8_mem_reg[1][19]/NET0131  & n3030 ;
  assign n5444 = \u8_mem_reg[3][19]/NET0131  & n2163 ;
  assign n5447 = ~n5443 & ~n5444 ;
  assign n5445 = \u8_mem_reg[2][19]/NET0131  & n3028 ;
  assign n5446 = \u8_mem_reg[0][19]/NET0131  & n3032 ;
  assign n5448 = ~n5445 & ~n5446 ;
  assign n5449 = n5447 & n5448 ;
  assign n5450 = n3037 & ~n5449 ;
  assign n5452 = n2159 & ~n5450 ;
  assign n5453 = ~n5451 & n5452 ;
  assign n5454 = ~n5442 & n5453 ;
  assign n5431 = ~\u8_dout_reg[19]/P0001  & ~n2159 ;
  assign n5455 = \u13_occ1_r_reg[8]/NET0131  & ~n5431 ;
  assign n5456 = ~n5454 & n5455 ;
  assign n5461 = \u3_mem_reg[2][21]/NET0131  & n3011 ;
  assign n5465 = \u3_rp_reg[0]/P0001  & ~n5461 ;
  assign n5464 = \u3_mem_reg[0][21]/NET0131  & n3015 ;
  assign n5462 = \u3_mem_reg[3][21]/NET0131  & n3009 ;
  assign n5463 = \u3_mem_reg[1][21]/NET0131  & n3013 ;
  assign n5466 = ~n5462 & ~n5463 ;
  assign n5467 = ~n5464 & n5466 ;
  assign n5468 = n5465 & n5467 ;
  assign n5460 = ~\u3_rp_reg[0]/P0001  & n5302 ;
  assign n5469 = n2784 & ~n5460 ;
  assign n5470 = ~n5468 & n5469 ;
  assign n5459 = n4799 & ~n4836 ;
  assign n5458 = n3020 & ~n4820 ;
  assign n5471 = n2787 & ~n5458 ;
  assign n5472 = ~n5459 & n5471 ;
  assign n5473 = ~n5470 & n5472 ;
  assign n5457 = ~\u3_dout_reg[9]/P0001  & ~n2787 ;
  assign n5474 = \u13_occ0_r_reg[0]/NET0131  & ~n5457 ;
  assign n5475 = ~n5473 & n5474 ;
  assign n5478 = \u8_mem_reg[3][2]/NET0131  & n2163 ;
  assign n5479 = \u8_mem_reg[0][2]/NET0131  & n3032 ;
  assign n5482 = ~n5478 & ~n5479 ;
  assign n5480 = \u8_mem_reg[1][2]/NET0131  & n3030 ;
  assign n5481 = \u8_mem_reg[2][2]/NET0131  & n3028 ;
  assign n5483 = ~n5480 & ~n5481 ;
  assign n5484 = n5482 & n5483 ;
  assign n5485 = n3037 & ~n5484 ;
  assign n5477 = ~n3036 & n5060 ;
  assign n5486 = n2159 & ~n5477 ;
  assign n5487 = ~n5485 & n5486 ;
  assign n5476 = ~\u8_dout_reg[2]/P0001  & ~n2159 ;
  assign n5488 = \u13_occ1_r_reg[8]/NET0131  & ~n5476 ;
  assign n5489 = ~n5487 & n5488 ;
  assign n5492 = \u8_mem_reg[3][3]/NET0131  & n2163 ;
  assign n5493 = \u8_mem_reg[0][3]/NET0131  & n3032 ;
  assign n5496 = ~n5492 & ~n5493 ;
  assign n5494 = \u8_mem_reg[2][3]/NET0131  & n3028 ;
  assign n5495 = \u8_mem_reg[1][3]/NET0131  & n3030 ;
  assign n5497 = ~n5494 & ~n5495 ;
  assign n5498 = n5496 & n5497 ;
  assign n5499 = n3037 & ~n5498 ;
  assign n5491 = ~n3059 & n5060 ;
  assign n5500 = n2159 & ~n5491 ;
  assign n5501 = ~n5499 & n5500 ;
  assign n5490 = ~\u8_dout_reg[3]/P0001  & ~n2159 ;
  assign n5502 = \u13_occ1_r_reg[8]/NET0131  & ~n5490 ;
  assign n5503 = ~n5501 & n5502 ;
  assign n5506 = \u8_rp_reg[0]/P0001  & n5328 ;
  assign n5505 = ~\u8_rp_reg[0]/P0001  & n3036 ;
  assign n5507 = n2160 & ~n5505 ;
  assign n5508 = ~n5506 & n5507 ;
  assign n5517 = n5060 & ~n5484 ;
  assign n5509 = \u8_mem_reg[3][4]/NET0131  & n2163 ;
  assign n5510 = \u8_mem_reg[2][4]/NET0131  & n3028 ;
  assign n5513 = ~n5509 & ~n5510 ;
  assign n5511 = \u8_mem_reg[0][4]/NET0131  & n3032 ;
  assign n5512 = \u8_mem_reg[1][4]/NET0131  & n3030 ;
  assign n5514 = ~n5511 & ~n5512 ;
  assign n5515 = n5513 & n5514 ;
  assign n5516 = n3037 & ~n5515 ;
  assign n5518 = n2159 & ~n5516 ;
  assign n5519 = ~n5517 & n5518 ;
  assign n5520 = ~n5508 & n5519 ;
  assign n5504 = ~\u8_dout_reg[4]/P0001  & ~n2159 ;
  assign n5521 = \u13_occ1_r_reg[8]/NET0131  & ~n5504 ;
  assign n5522 = ~n5520 & n5521 ;
  assign n5525 = \u8_rp_reg[0]/P0001  & n5354 ;
  assign n5524 = ~\u8_rp_reg[0]/P0001  & n3059 ;
  assign n5526 = n2160 & ~n5524 ;
  assign n5527 = ~n5525 & n5526 ;
  assign n5536 = n5060 & ~n5498 ;
  assign n5528 = \u8_mem_reg[3][5]/NET0131  & n2163 ;
  assign n5529 = \u8_mem_reg[2][5]/NET0131  & n3028 ;
  assign n5532 = ~n5528 & ~n5529 ;
  assign n5530 = \u8_mem_reg[1][5]/NET0131  & n3030 ;
  assign n5531 = \u8_mem_reg[0][5]/NET0131  & n3032 ;
  assign n5533 = ~n5530 & ~n5531 ;
  assign n5534 = n5532 & n5533 ;
  assign n5535 = n3037 & ~n5534 ;
  assign n5537 = n2159 & ~n5535 ;
  assign n5538 = ~n5536 & n5537 ;
  assign n5539 = ~n5527 & n5538 ;
  assign n5523 = ~\u8_dout_reg[5]/P0001  & ~n2159 ;
  assign n5540 = \u13_occ1_r_reg[8]/NET0131  & ~n5523 ;
  assign n5541 = ~n5539 & n5540 ;
  assign n5544 = \u8_rp_reg[0]/P0001  & n5404 ;
  assign n5543 = ~\u8_rp_reg[0]/P0001  & n5484 ;
  assign n5545 = n2160 & ~n5543 ;
  assign n5546 = ~n5544 & n5545 ;
  assign n5548 = n5060 & ~n5515 ;
  assign n5547 = n3037 & ~n5040 ;
  assign n5549 = n2159 & ~n5547 ;
  assign n5550 = ~n5548 & n5549 ;
  assign n5551 = ~n5546 & n5550 ;
  assign n5542 = ~\u8_dout_reg[6]/P0001  & ~n2159 ;
  assign n5552 = \u13_occ1_r_reg[8]/NET0131  & ~n5542 ;
  assign n5553 = ~n5551 & n5552 ;
  assign n5556 = \u8_rp_reg[0]/P0001  & n5449 ;
  assign n5555 = ~\u8_rp_reg[0]/P0001  & n5498 ;
  assign n5557 = n2160 & ~n5555 ;
  assign n5558 = ~n5556 & n5557 ;
  assign n5560 = n5060 & ~n5534 ;
  assign n5559 = n3037 & ~n5107 ;
  assign n5561 = n2159 & ~n5559 ;
  assign n5562 = ~n5560 & n5561 ;
  assign n5563 = ~n5558 & n5562 ;
  assign n5554 = ~\u8_dout_reg[7]/P0001  & ~n2159 ;
  assign n5564 = \u13_occ1_r_reg[8]/NET0131  & ~n5554 ;
  assign n5565 = ~n5563 & n5564 ;
  assign n5568 = \u8_mem_reg[2][20]/NET0131  & n3028 ;
  assign n5572 = \u8_rp_reg[0]/P0001  & ~n5568 ;
  assign n5571 = \u8_mem_reg[0][20]/NET0131  & n3032 ;
  assign n5569 = \u8_mem_reg[3][20]/NET0131  & n2163 ;
  assign n5570 = \u8_mem_reg[1][20]/NET0131  & n3030 ;
  assign n5573 = ~n5569 & ~n5570 ;
  assign n5574 = ~n5571 & n5573 ;
  assign n5575 = n5572 & n5574 ;
  assign n5567 = ~\u8_rp_reg[0]/P0001  & n5515 ;
  assign n5576 = n2160 & ~n5567 ;
  assign n5577 = ~n5575 & n5576 ;
  assign n5579 = ~n5040 & n5060 ;
  assign n5578 = n3037 & ~n5067 ;
  assign n5580 = n2159 & ~n5578 ;
  assign n5581 = ~n5579 & n5580 ;
  assign n5582 = ~n5577 & n5581 ;
  assign n5566 = ~\u8_dout_reg[8]/P0001  & ~n2159 ;
  assign n5583 = \u13_occ1_r_reg[8]/NET0131  & ~n5566 ;
  assign n5584 = ~n5582 & n5583 ;
  assign n5587 = \u8_mem_reg[2][21]/NET0131  & n3028 ;
  assign n5591 = \u8_rp_reg[0]/P0001  & ~n5587 ;
  assign n5590 = \u8_mem_reg[0][21]/NET0131  & n3032 ;
  assign n5588 = \u8_mem_reg[3][21]/NET0131  & n2163 ;
  assign n5589 = \u8_mem_reg[1][21]/NET0131  & n3030 ;
  assign n5592 = ~n5588 & ~n5589 ;
  assign n5593 = ~n5590 & n5592 ;
  assign n5594 = n5591 & n5593 ;
  assign n5586 = ~\u8_rp_reg[0]/P0001  & n5534 ;
  assign n5595 = n2160 & ~n5586 ;
  assign n5596 = ~n5594 & n5595 ;
  assign n5598 = n5060 & ~n5107 ;
  assign n5597 = n3037 & ~n5133 ;
  assign n5599 = n2159 & ~n5597 ;
  assign n5600 = ~n5598 & n5599 ;
  assign n5601 = ~n5596 & n5600 ;
  assign n5585 = ~\u8_dout_reg[9]/P0001  & ~n2159 ;
  assign n5602 = \u13_occ1_r_reg[8]/NET0131  & ~n5585 ;
  assign n5603 = ~n5601 & n5602 ;
  assign n5604 = ~\u11_wp_reg[1]/P0001  & ~n3066 ;
  assign n5605 = \u13_icc_r_reg[16]/NET0131  & ~n3067 ;
  assign n5606 = ~n5604 & n5605 ;
  assign n5607 = ~\u9_wp_reg[1]/P0001  & ~n3313 ;
  assign n5608 = \u13_icc_r_reg[0]/NET0131  & ~n3314 ;
  assign n5609 = ~n5607 & n5608 ;
  assign n5610 = ~\u10_wp_reg[1]/P0001  & ~n3503 ;
  assign n5611 = \u13_icc_r_reg[8]/NET0131  & ~n3504 ;
  assign n5612 = ~n5610 & n5611 ;
  assign n5614 = \u11_wp_reg[3]/P0001  & n3068 ;
  assign n5613 = ~\u11_wp_reg[3]/P0001  & ~n3068 ;
  assign n5615 = \u13_icc_r_reg[16]/NET0131  & ~n5613 ;
  assign n5616 = ~n5614 & n5615 ;
  assign n5618 = \u9_wp_reg[3]/P0001  & n3315 ;
  assign n5617 = ~\u9_wp_reg[3]/P0001  & ~n3315 ;
  assign n5619 = \u13_icc_r_reg[0]/NET0131  & ~n5617 ;
  assign n5620 = ~n5618 & n5619 ;
  assign n5622 = \u10_wp_reg[3]/P0001  & n3505 ;
  assign n5621 = ~\u10_wp_reg[3]/P0001  & ~n3505 ;
  assign n5623 = \u13_icc_r_reg[8]/NET0131  & ~n5621 ;
  assign n5624 = ~n5622 & n5623 ;
  assign n5625 = \u26_ps_cnt_reg[0]/NET0131  & ~\u26_ps_cnt_reg[1]/NET0131  ;
  assign n5626 = ~\u26_ps_cnt_reg[2]/NET0131  & ~\u26_ps_cnt_reg[3]/NET0131  ;
  assign n5627 = \u26_ps_cnt_reg[4]/NET0131  & \u26_ps_cnt_reg[5]/NET0131  ;
  assign n5628 = n5626 & n5627 ;
  assign n5629 = n5625 & n5628 ;
  assign n5630 = ~\u13_ac97_rst_force_reg/P0001  & ~n5629 ;
  assign n5631 = ~\u26_ps_cnt_reg[0]/NET0131  & n5630 ;
  assign n5632 = ~\u26_ps_cnt_reg[0]/NET0131  & \u26_ps_cnt_reg[1]/NET0131  ;
  assign n5633 = ~n5625 & ~n5632 ;
  assign n5634 = n5630 & ~n5633 ;
  assign n5635 = \u26_ps_cnt_reg[0]/NET0131  & \u26_ps_cnt_reg[1]/NET0131  ;
  assign n5636 = \u26_ps_cnt_reg[2]/NET0131  & n5635 ;
  assign n5637 = ~\u26_ps_cnt_reg[2]/NET0131  & ~n5635 ;
  assign n5638 = ~n5636 & ~n5637 ;
  assign n5639 = n5630 & n5638 ;
  assign n5640 = ~\u26_ps_cnt_reg[3]/NET0131  & ~n5636 ;
  assign n5641 = \u26_ps_cnt_reg[3]/NET0131  & n5636 ;
  assign n5642 = ~n5640 & ~n5641 ;
  assign n5643 = n5630 & n5642 ;
  assign n5645 = ~\u26_ps_cnt_reg[4]/NET0131  & ~n5641 ;
  assign n5644 = \u26_ps_cnt_reg[4]/NET0131  & n5641 ;
  assign n5646 = n5630 & ~n5644 ;
  assign n5647 = ~n5645 & n5646 ;
  assign n5649 = \u26_ps_cnt_reg[5]/NET0131  & n5644 ;
  assign n5648 = ~\u26_ps_cnt_reg[5]/NET0131  & ~n5644 ;
  assign n5650 = n5630 & ~n5648 ;
  assign n5651 = ~n5649 & n5650 ;
  assign n5652 = n3063 & n3064 ;
  assign n5654 = \u11_wp_reg[0]/NET0131  & n5652 ;
  assign n5653 = ~\u11_wp_reg[0]/NET0131  & ~n5652 ;
  assign n5655 = \u13_icc_r_reg[16]/NET0131  & ~n5653 ;
  assign n5656 = ~n5654 & n5655 ;
  assign n5657 = n3310 & n3311 ;
  assign n5659 = \u9_wp_reg[0]/NET0131  & n5657 ;
  assign n5658 = ~\u9_wp_reg[0]/NET0131  & ~n5657 ;
  assign n5660 = \u13_icc_r_reg[0]/NET0131  & ~n5658 ;
  assign n5661 = ~n5659 & n5660 ;
  assign n5662 = n3500 & n3501 ;
  assign n5664 = \u10_wp_reg[0]/NET0131  & n5662 ;
  assign n5663 = ~\u10_wp_reg[0]/NET0131  & ~n5662 ;
  assign n5665 = \u13_icc_r_reg[8]/NET0131  & ~n5663 ;
  assign n5666 = ~n5664 & n5665 ;
  assign n5667 = ~\u10_wp_reg[1]/P0001  & \u10_wp_reg[2]/P0001  ;
  assign n5668 = n3503 & n5667 ;
  assign n5669 = \u10_mem_reg[2][18]/P0001  & ~n5668 ;
  assign n5670 = \u1_slt4_reg[6]/P0001  & n3501 ;
  assign n5671 = ~\u13_icc_r_reg[10]/NET0131  & \u13_icc_r_reg[11]/NET0131  ;
  assign n5672 = \u1_slt4_reg[18]/P0001  & n5671 ;
  assign n5673 = ~n5670 & ~n5672 ;
  assign n5674 = n5668 & ~n5673 ;
  assign n5675 = ~n5669 & ~n5674 ;
  assign n5676 = \u10_mem_reg[2][19]/P0001  & ~n5668 ;
  assign n5677 = \u1_slt4_reg[7]/P0001  & n3501 ;
  assign n5678 = \u1_slt4_reg[19]/P0001  & n5671 ;
  assign n5679 = ~n5677 & ~n5678 ;
  assign n5680 = n5668 & ~n5679 ;
  assign n5681 = ~n5676 & ~n5680 ;
  assign n5682 = \u10_mem_reg[2][20]/P0001  & ~n5668 ;
  assign n5683 = \u1_slt4_reg[8]/P0001  & n3501 ;
  assign n5684 = n5668 & n5683 ;
  assign n5685 = ~n5682 & ~n5684 ;
  assign n5686 = \u10_mem_reg[2][21]/P0001  & ~n5668 ;
  assign n5687 = \u1_slt4_reg[9]/P0001  & n3501 ;
  assign n5688 = n5668 & n5687 ;
  assign n5689 = ~n5686 & ~n5688 ;
  assign n5690 = \u10_mem_reg[2][22]/P0001  & ~n5668 ;
  assign n5691 = \u1_slt4_reg[10]/P0001  & n3501 ;
  assign n5692 = n5668 & n5691 ;
  assign n5693 = ~n5690 & ~n5692 ;
  assign n5694 = \u10_mem_reg[2][23]/P0001  & ~n5668 ;
  assign n5695 = \u1_slt4_reg[11]/P0001  & n3501 ;
  assign n5696 = n5668 & n5695 ;
  assign n5697 = ~n5694 & ~n5696 ;
  assign n5698 = ~\u9_wp_reg[1]/P0001  & ~\u9_wp_reg[2]/P0001  ;
  assign n5699 = n3313 & n5698 ;
  assign n5700 = \u1_slt3_reg[6]/P0001  & n3311 ;
  assign n5701 = ~\u13_icc_r_reg[2]/NET0131  & \u13_icc_r_reg[3]/NET0131  ;
  assign n5702 = \u1_slt3_reg[18]/P0001  & n5701 ;
  assign n5703 = ~n5700 & ~n5702 ;
  assign n5704 = n5699 & ~n5703 ;
  assign n5705 = \u9_mem_reg[0][18]/P0001  & ~n5699 ;
  assign n5706 = ~n5704 & ~n5705 ;
  assign n5707 = \u1_slt3_reg[7]/P0001  & n3311 ;
  assign n5708 = \u1_slt3_reg[19]/P0001  & n5701 ;
  assign n5709 = ~n5707 & ~n5708 ;
  assign n5710 = n5699 & ~n5709 ;
  assign n5711 = \u9_mem_reg[0][19]/P0001  & ~n5699 ;
  assign n5712 = ~n5710 & ~n5711 ;
  assign n5713 = \u10_mem_reg[2][24]/P0001  & ~n5668 ;
  assign n5714 = \u1_slt4_reg[12]/P0001  & n3501 ;
  assign n5715 = n5668 & n5714 ;
  assign n5716 = ~n5713 & ~n5715 ;
  assign n5717 = \u10_mem_reg[2][25]/P0001  & ~n5668 ;
  assign n5718 = \u1_slt4_reg[13]/P0001  & n3501 ;
  assign n5719 = n5668 & n5718 ;
  assign n5720 = ~n5717 & ~n5719 ;
  assign n5721 = \u10_mem_reg[2][26]/P0001  & ~n5668 ;
  assign n5722 = \u1_slt4_reg[14]/P0001  & n3501 ;
  assign n5723 = n5668 & n5722 ;
  assign n5724 = ~n5721 & ~n5723 ;
  assign n5725 = \u10_mem_reg[2][27]/P0001  & ~n5668 ;
  assign n5726 = \u1_slt4_reg[15]/P0001  & n3501 ;
  assign n5727 = n5668 & n5726 ;
  assign n5728 = ~n5725 & ~n5727 ;
  assign n5729 = \u10_mem_reg[2][28]/P0001  & ~n5668 ;
  assign n5730 = \u1_slt4_reg[16]/P0001  & n3501 ;
  assign n5731 = n5668 & n5730 ;
  assign n5732 = ~n5729 & ~n5731 ;
  assign n5733 = ~\u9_wp_reg[2]/P0001  & n3314 ;
  assign n5734 = ~n5703 & n5733 ;
  assign n5735 = \u9_mem_reg[1][18]/P0001  & ~n5733 ;
  assign n5736 = ~n5734 & ~n5735 ;
  assign n5737 = ~n5709 & n5733 ;
  assign n5738 = \u9_mem_reg[1][19]/P0001  & ~n5733 ;
  assign n5739 = ~n5737 & ~n5738 ;
  assign n5740 = \u9_mem_reg[1][20]/P0001  & ~n5733 ;
  assign n5741 = \u1_slt3_reg[8]/P0001  & n3311 ;
  assign n5742 = n5733 & n5741 ;
  assign n5743 = ~n5740 & ~n5742 ;
  assign n5744 = \u9_mem_reg[1][21]/P0001  & ~n5733 ;
  assign n5745 = \u1_slt3_reg[9]/P0001  & n3311 ;
  assign n5746 = n5733 & n5745 ;
  assign n5747 = ~n5744 & ~n5746 ;
  assign n5748 = \u10_mem_reg[2][29]/P0001  & ~n5668 ;
  assign n5749 = \u1_slt4_reg[17]/P0001  & n3501 ;
  assign n5750 = n5668 & n5749 ;
  assign n5751 = ~n5748 & ~n5750 ;
  assign n5752 = \u9_mem_reg[1][22]/P0001  & ~n5733 ;
  assign n5753 = \u1_slt3_reg[10]/P0001  & n3311 ;
  assign n5754 = n5733 & n5753 ;
  assign n5755 = ~n5752 & ~n5754 ;
  assign n5756 = \u9_mem_reg[1][23]/P0001  & ~n5733 ;
  assign n5757 = \u1_slt3_reg[11]/P0001  & n3311 ;
  assign n5758 = n5733 & n5757 ;
  assign n5759 = ~n5756 & ~n5758 ;
  assign n5760 = \u9_mem_reg[1][24]/P0001  & ~n5733 ;
  assign n5761 = \u1_slt3_reg[12]/P0001  & n3311 ;
  assign n5762 = n5733 & n5761 ;
  assign n5763 = ~n5760 & ~n5762 ;
  assign n5764 = \u9_mem_reg[1][25]/P0001  & ~n5733 ;
  assign n5765 = \u1_slt3_reg[13]/P0001  & n3311 ;
  assign n5766 = n5733 & n5765 ;
  assign n5767 = ~n5764 & ~n5766 ;
  assign n5768 = \u9_mem_reg[1][26]/P0001  & ~n5733 ;
  assign n5769 = \u1_slt3_reg[14]/P0001  & n3311 ;
  assign n5770 = n5733 & n5769 ;
  assign n5771 = ~n5768 & ~n5770 ;
  assign n5772 = \u9_mem_reg[1][27]/P0001  & ~n5733 ;
  assign n5773 = \u1_slt3_reg[15]/P0001  & n3311 ;
  assign n5774 = n5733 & n5773 ;
  assign n5775 = ~n5772 & ~n5774 ;
  assign n5776 = \u9_mem_reg[1][28]/P0001  & ~n5733 ;
  assign n5777 = \u1_slt3_reg[16]/P0001  & n3311 ;
  assign n5778 = n5733 & n5777 ;
  assign n5779 = ~n5776 & ~n5778 ;
  assign n5780 = \u9_mem_reg[1][29]/P0001  & ~n5733 ;
  assign n5781 = \u1_slt3_reg[17]/P0001  & n3311 ;
  assign n5782 = n5733 & n5781 ;
  assign n5783 = ~n5780 & ~n5782 ;
  assign n5784 = \u9_mem_reg[1][30]/P0001  & ~n5733 ;
  assign n5785 = \u1_slt3_reg[18]/P0001  & n3311 ;
  assign n5786 = n5733 & n5785 ;
  assign n5787 = ~n5784 & ~n5786 ;
  assign n5788 = \u9_mem_reg[1][31]/P0001  & ~n5733 ;
  assign n5789 = \u1_slt3_reg[19]/P0001  & n3311 ;
  assign n5790 = n5733 & n5789 ;
  assign n5791 = ~n5788 & ~n5790 ;
  assign n5792 = \u10_mem_reg[2][30]/P0001  & ~n5668 ;
  assign n5793 = \u1_slt4_reg[18]/P0001  & n3501 ;
  assign n5794 = n5668 & n5793 ;
  assign n5795 = ~n5792 & ~n5794 ;
  assign n5796 = \u10_mem_reg[2][31]/P0001  & ~n5668 ;
  assign n5797 = \u1_slt4_reg[19]/P0001  & n3501 ;
  assign n5798 = n5668 & n5797 ;
  assign n5799 = ~n5796 & ~n5798 ;
  assign n5800 = ~\u9_wp_reg[1]/P0001  & \u9_wp_reg[2]/P0001  ;
  assign n5801 = n3313 & n5800 ;
  assign n5802 = \u9_mem_reg[2][18]/P0001  & ~n5801 ;
  assign n5803 = ~n5703 & n5801 ;
  assign n5804 = ~n5802 & ~n5803 ;
  assign n5805 = \u9_mem_reg[2][19]/P0001  & ~n5801 ;
  assign n5806 = ~n5709 & n5801 ;
  assign n5807 = ~n5805 & ~n5806 ;
  assign n5808 = \u9_mem_reg[2][20]/P0001  & ~n5801 ;
  assign n5809 = n5741 & n5801 ;
  assign n5810 = ~n5808 & ~n5809 ;
  assign n5811 = \u9_mem_reg[2][21]/P0001  & ~n5801 ;
  assign n5812 = n5745 & n5801 ;
  assign n5813 = ~n5811 & ~n5812 ;
  assign n5814 = \u9_mem_reg[2][22]/P0001  & ~n5801 ;
  assign n5815 = n5753 & n5801 ;
  assign n5816 = ~n5814 & ~n5815 ;
  assign n5817 = \u9_mem_reg[2][23]/P0001  & ~n5801 ;
  assign n5818 = n5757 & n5801 ;
  assign n5819 = ~n5817 & ~n5818 ;
  assign n5820 = \u9_mem_reg[2][24]/P0001  & ~n5801 ;
  assign n5821 = n5761 & n5801 ;
  assign n5822 = ~n5820 & ~n5821 ;
  assign n5823 = \u9_mem_reg[2][25]/P0001  & ~n5801 ;
  assign n5824 = n5765 & n5801 ;
  assign n5825 = ~n5823 & ~n5824 ;
  assign n5826 = \u9_mem_reg[2][26]/P0001  & ~n5801 ;
  assign n5827 = n5769 & n5801 ;
  assign n5828 = ~n5826 & ~n5827 ;
  assign n5829 = \u9_mem_reg[2][27]/P0001  & ~n5801 ;
  assign n5830 = n5773 & n5801 ;
  assign n5831 = ~n5829 & ~n5830 ;
  assign n5832 = \u9_mem_reg[2][28]/P0001  & ~n5801 ;
  assign n5833 = n5777 & n5801 ;
  assign n5834 = ~n5832 & ~n5833 ;
  assign n5835 = \u9_mem_reg[2][29]/P0001  & ~n5801 ;
  assign n5836 = n5781 & n5801 ;
  assign n5837 = ~n5835 & ~n5836 ;
  assign n5838 = \u9_mem_reg[2][30]/P0001  & ~n5801 ;
  assign n5839 = n5785 & n5801 ;
  assign n5840 = ~n5838 & ~n5839 ;
  assign n5841 = \u9_mem_reg[2][31]/P0001  & ~n5801 ;
  assign n5842 = n5789 & n5801 ;
  assign n5843 = ~n5841 & ~n5842 ;
  assign n5844 = n3315 & ~n5703 ;
  assign n5845 = \u9_mem_reg[3][18]/P0001  & ~n3315 ;
  assign n5846 = ~n5844 & ~n5845 ;
  assign n5847 = n3315 & ~n5709 ;
  assign n5848 = \u9_mem_reg[3][19]/P0001  & ~n3315 ;
  assign n5849 = ~n5847 & ~n5848 ;
  assign n5850 = \u9_mem_reg[3][20]/P0001  & ~n3315 ;
  assign n5851 = n3315 & n5741 ;
  assign n5852 = ~n5850 & ~n5851 ;
  assign n5853 = \u9_mem_reg[3][21]/P0001  & ~n3315 ;
  assign n5854 = n3315 & n5745 ;
  assign n5855 = ~n5853 & ~n5854 ;
  assign n5856 = \u9_mem_reg[3][22]/P0001  & ~n3315 ;
  assign n5857 = n3315 & n5753 ;
  assign n5858 = ~n5856 & ~n5857 ;
  assign n5859 = \u9_mem_reg[3][23]/P0001  & ~n3315 ;
  assign n5860 = n3315 & n5757 ;
  assign n5861 = ~n5859 & ~n5860 ;
  assign n5862 = \u9_mem_reg[3][24]/P0001  & ~n3315 ;
  assign n5863 = n3315 & n5761 ;
  assign n5864 = ~n5862 & ~n5863 ;
  assign n5865 = \u9_mem_reg[3][25]/P0001  & ~n3315 ;
  assign n5866 = n3315 & n5765 ;
  assign n5867 = ~n5865 & ~n5866 ;
  assign n5868 = \u9_mem_reg[3][26]/P0001  & ~n3315 ;
  assign n5869 = n3315 & n5769 ;
  assign n5870 = ~n5868 & ~n5869 ;
  assign n5871 = \u9_mem_reg[3][27]/P0001  & ~n3315 ;
  assign n5872 = n3315 & n5773 ;
  assign n5873 = ~n5871 & ~n5872 ;
  assign n5874 = \u9_mem_reg[3][28]/P0001  & ~n3315 ;
  assign n5875 = n3315 & n5777 ;
  assign n5876 = ~n5874 & ~n5875 ;
  assign n5877 = \u9_mem_reg[3][29]/P0001  & ~n3315 ;
  assign n5878 = n3315 & n5781 ;
  assign n5879 = ~n5877 & ~n5878 ;
  assign n5880 = \u9_mem_reg[3][30]/P0001  & ~n3315 ;
  assign n5881 = n3315 & n5785 ;
  assign n5882 = ~n5880 & ~n5881 ;
  assign n5883 = \u9_mem_reg[3][31]/P0001  & ~n3315 ;
  assign n5884 = n3315 & n5789 ;
  assign n5885 = ~n5883 & ~n5884 ;
  assign n5886 = n3505 & ~n5673 ;
  assign n5887 = \u10_mem_reg[3][18]/P0001  & ~n3505 ;
  assign n5888 = ~n5886 & ~n5887 ;
  assign n5889 = n3505 & ~n5679 ;
  assign n5890 = \u10_mem_reg[3][19]/P0001  & ~n3505 ;
  assign n5891 = ~n5889 & ~n5890 ;
  assign n5892 = \u10_mem_reg[3][20]/P0001  & ~n3505 ;
  assign n5893 = n3505 & n5683 ;
  assign n5894 = ~n5892 & ~n5893 ;
  assign n5895 = \u10_mem_reg[3][21]/P0001  & ~n3505 ;
  assign n5896 = n3505 & n5687 ;
  assign n5897 = ~n5895 & ~n5896 ;
  assign n5898 = \u10_mem_reg[3][22]/P0001  & ~n3505 ;
  assign n5899 = n3505 & n5691 ;
  assign n5900 = ~n5898 & ~n5899 ;
  assign n5901 = \u10_mem_reg[3][23]/P0001  & ~n3505 ;
  assign n5902 = n3505 & n5695 ;
  assign n5903 = ~n5901 & ~n5902 ;
  assign n5904 = \u10_mem_reg[3][24]/P0001  & ~n3505 ;
  assign n5905 = n3505 & n5714 ;
  assign n5906 = ~n5904 & ~n5905 ;
  assign n5907 = \u10_mem_reg[3][25]/P0001  & ~n3505 ;
  assign n5908 = n3505 & n5718 ;
  assign n5909 = ~n5907 & ~n5908 ;
  assign n5910 = \u10_mem_reg[3][26]/P0001  & ~n3505 ;
  assign n5911 = n3505 & n5722 ;
  assign n5912 = ~n5910 & ~n5911 ;
  assign n5913 = \u10_mem_reg[3][27]/P0001  & ~n3505 ;
  assign n5914 = n3505 & n5726 ;
  assign n5915 = ~n5913 & ~n5914 ;
  assign n5916 = \u10_mem_reg[3][28]/P0001  & ~n3505 ;
  assign n5917 = n3505 & n5730 ;
  assign n5918 = ~n5916 & ~n5917 ;
  assign n5919 = \u10_mem_reg[3][29]/P0001  & ~n3505 ;
  assign n5920 = n3505 & n5749 ;
  assign n5921 = ~n5919 & ~n5920 ;
  assign n5922 = \u10_mem_reg[3][30]/P0001  & ~n3505 ;
  assign n5923 = n3505 & n5793 ;
  assign n5924 = ~n5922 & ~n5923 ;
  assign n5925 = \u10_mem_reg[3][31]/P0001  & ~n3505 ;
  assign n5926 = n3505 & n5797 ;
  assign n5927 = ~n5925 & ~n5926 ;
  assign n5928 = ~\u10_wp_reg[1]/P0001  & ~\u10_wp_reg[2]/P0001  ;
  assign n5929 = n3503 & n5928 ;
  assign n5930 = \u10_mem_reg[0][18]/P0001  & ~n5929 ;
  assign n5931 = ~n5673 & n5929 ;
  assign n5932 = ~n5930 & ~n5931 ;
  assign n5933 = ~\u11_wp_reg[1]/P0001  & ~\u11_wp_reg[2]/P0001  ;
  assign n5934 = n3066 & n5933 ;
  assign n5935 = \u1_slt6_reg[6]/P0001  & n3064 ;
  assign n5936 = ~\u13_icc_r_reg[18]/NET0131  & \u13_icc_r_reg[19]/NET0131  ;
  assign n5937 = \u1_slt6_reg[18]/P0001  & n5936 ;
  assign n5938 = ~n5935 & ~n5937 ;
  assign n5939 = n5934 & ~n5938 ;
  assign n5940 = \u11_mem_reg[0][18]/P0001  & ~n5934 ;
  assign n5941 = ~n5939 & ~n5940 ;
  assign n5942 = \u1_slt6_reg[7]/P0001  & n3064 ;
  assign n5943 = \u1_slt6_reg[19]/P0001  & n5936 ;
  assign n5944 = ~n5942 & ~n5943 ;
  assign n5945 = n5934 & ~n5944 ;
  assign n5946 = \u11_mem_reg[0][19]/P0001  & ~n5934 ;
  assign n5947 = ~n5945 & ~n5946 ;
  assign n5948 = \u10_mem_reg[0][19]/P0001  & ~n5929 ;
  assign n5949 = ~n5679 & n5929 ;
  assign n5950 = ~n5948 & ~n5949 ;
  assign n5951 = ~\u11_wp_reg[2]/P0001  & n3067 ;
  assign n5952 = ~n5938 & n5951 ;
  assign n5953 = \u11_mem_reg[1][18]/P0001  & ~n5951 ;
  assign n5954 = ~n5952 & ~n5953 ;
  assign n5955 = ~n5944 & n5951 ;
  assign n5956 = \u11_mem_reg[1][19]/P0001  & ~n5951 ;
  assign n5957 = ~n5955 & ~n5956 ;
  assign n5958 = \u11_mem_reg[1][20]/P0001  & ~n5951 ;
  assign n5959 = \u1_slt6_reg[8]/P0001  & n3064 ;
  assign n5960 = n5951 & n5959 ;
  assign n5961 = ~n5958 & ~n5960 ;
  assign n5962 = \u11_mem_reg[1][21]/P0001  & ~n5951 ;
  assign n5963 = \u1_slt6_reg[9]/P0001  & n3064 ;
  assign n5964 = n5951 & n5963 ;
  assign n5965 = ~n5962 & ~n5964 ;
  assign n5966 = \u11_mem_reg[1][22]/P0001  & ~n5951 ;
  assign n5967 = \u1_slt6_reg[10]/P0001  & n3064 ;
  assign n5968 = n5951 & n5967 ;
  assign n5969 = ~n5966 & ~n5968 ;
  assign n5970 = \u11_mem_reg[1][23]/P0001  & ~n5951 ;
  assign n5971 = \u1_slt6_reg[11]/P0001  & n3064 ;
  assign n5972 = n5951 & n5971 ;
  assign n5973 = ~n5970 & ~n5972 ;
  assign n5974 = \u11_mem_reg[1][24]/P0001  & ~n5951 ;
  assign n5975 = \u1_slt6_reg[12]/P0001  & n3064 ;
  assign n5976 = n5951 & n5975 ;
  assign n5977 = ~n5974 & ~n5976 ;
  assign n5978 = \u11_mem_reg[1][25]/P0001  & ~n5951 ;
  assign n5979 = \u1_slt6_reg[13]/P0001  & n3064 ;
  assign n5980 = n5951 & n5979 ;
  assign n5981 = ~n5978 & ~n5980 ;
  assign n5982 = \u11_mem_reg[1][26]/P0001  & ~n5951 ;
  assign n5983 = \u1_slt6_reg[14]/P0001  & n3064 ;
  assign n5984 = n5951 & n5983 ;
  assign n5985 = ~n5982 & ~n5984 ;
  assign n5986 = \u11_mem_reg[1][27]/P0001  & ~n5951 ;
  assign n5987 = \u1_slt6_reg[15]/P0001  & n3064 ;
  assign n5988 = n5951 & n5987 ;
  assign n5989 = ~n5986 & ~n5988 ;
  assign n5990 = \u11_mem_reg[1][28]/P0001  & ~n5951 ;
  assign n5991 = \u1_slt6_reg[16]/P0001  & n3064 ;
  assign n5992 = n5951 & n5991 ;
  assign n5993 = ~n5990 & ~n5992 ;
  assign n5994 = \u11_mem_reg[1][29]/P0001  & ~n5951 ;
  assign n5995 = \u1_slt6_reg[17]/P0001  & n3064 ;
  assign n5996 = n5951 & n5995 ;
  assign n5997 = ~n5994 & ~n5996 ;
  assign n5998 = \u11_mem_reg[1][30]/P0001  & ~n5951 ;
  assign n5999 = \u1_slt6_reg[18]/P0001  & n3064 ;
  assign n6000 = n5951 & n5999 ;
  assign n6001 = ~n5998 & ~n6000 ;
  assign n6002 = \u11_mem_reg[1][31]/P0001  & ~n5951 ;
  assign n6003 = \u1_slt6_reg[19]/P0001  & n3064 ;
  assign n6004 = n5951 & n6003 ;
  assign n6005 = ~n6002 & ~n6004 ;
  assign n6006 = ~\u11_wp_reg[1]/P0001  & \u11_wp_reg[2]/P0001  ;
  assign n6007 = n3066 & n6006 ;
  assign n6008 = \u11_mem_reg[2][18]/P0001  & ~n6007 ;
  assign n6009 = ~n5938 & n6007 ;
  assign n6010 = ~n6008 & ~n6009 ;
  assign n6011 = \u11_mem_reg[2][19]/P0001  & ~n6007 ;
  assign n6012 = ~n5944 & n6007 ;
  assign n6013 = ~n6011 & ~n6012 ;
  assign n6014 = \u11_mem_reg[2][20]/P0001  & ~n6007 ;
  assign n6015 = n5959 & n6007 ;
  assign n6016 = ~n6014 & ~n6015 ;
  assign n6017 = \u11_mem_reg[2][21]/P0001  & ~n6007 ;
  assign n6018 = n5963 & n6007 ;
  assign n6019 = ~n6017 & ~n6018 ;
  assign n6020 = \u11_mem_reg[2][22]/P0001  & ~n6007 ;
  assign n6021 = n5967 & n6007 ;
  assign n6022 = ~n6020 & ~n6021 ;
  assign n6023 = \u11_mem_reg[2][23]/P0001  & ~n6007 ;
  assign n6024 = n5971 & n6007 ;
  assign n6025 = ~n6023 & ~n6024 ;
  assign n6026 = \u11_mem_reg[2][24]/P0001  & ~n6007 ;
  assign n6027 = n5975 & n6007 ;
  assign n6028 = ~n6026 & ~n6027 ;
  assign n6029 = \u11_mem_reg[2][25]/P0001  & ~n6007 ;
  assign n6030 = n5979 & n6007 ;
  assign n6031 = ~n6029 & ~n6030 ;
  assign n6032 = ~\u10_wp_reg[2]/P0001  & n3504 ;
  assign n6033 = ~n5673 & n6032 ;
  assign n6034 = \u10_mem_reg[1][18]/P0001  & ~n6032 ;
  assign n6035 = ~n6033 & ~n6034 ;
  assign n6036 = \u11_mem_reg[2][26]/P0001  & ~n6007 ;
  assign n6037 = n5983 & n6007 ;
  assign n6038 = ~n6036 & ~n6037 ;
  assign n6039 = \u11_mem_reg[2][27]/P0001  & ~n6007 ;
  assign n6040 = n5987 & n6007 ;
  assign n6041 = ~n6039 & ~n6040 ;
  assign n6042 = ~n5679 & n6032 ;
  assign n6043 = \u10_mem_reg[1][19]/P0001  & ~n6032 ;
  assign n6044 = ~n6042 & ~n6043 ;
  assign n6045 = \u11_mem_reg[2][28]/P0001  & ~n6007 ;
  assign n6046 = n5991 & n6007 ;
  assign n6047 = ~n6045 & ~n6046 ;
  assign n6048 = \u11_mem_reg[2][29]/P0001  & ~n6007 ;
  assign n6049 = n5995 & n6007 ;
  assign n6050 = ~n6048 & ~n6049 ;
  assign n6051 = \u11_mem_reg[2][30]/P0001  & ~n6007 ;
  assign n6052 = n5999 & n6007 ;
  assign n6053 = ~n6051 & ~n6052 ;
  assign n6054 = \u10_mem_reg[1][20]/P0001  & ~n6032 ;
  assign n6055 = n5683 & n6032 ;
  assign n6056 = ~n6054 & ~n6055 ;
  assign n6057 = \u11_mem_reg[2][31]/P0001  & ~n6007 ;
  assign n6058 = n6003 & n6007 ;
  assign n6059 = ~n6057 & ~n6058 ;
  assign n6060 = \u10_mem_reg[1][21]/P0001  & ~n6032 ;
  assign n6061 = n5687 & n6032 ;
  assign n6062 = ~n6060 & ~n6061 ;
  assign n6063 = \u10_mem_reg[1][22]/P0001  & ~n6032 ;
  assign n6064 = n5691 & n6032 ;
  assign n6065 = ~n6063 & ~n6064 ;
  assign n6066 = \u10_mem_reg[1][23]/P0001  & ~n6032 ;
  assign n6067 = n5695 & n6032 ;
  assign n6068 = ~n6066 & ~n6067 ;
  assign n6069 = \u10_mem_reg[1][24]/P0001  & ~n6032 ;
  assign n6070 = n5714 & n6032 ;
  assign n6071 = ~n6069 & ~n6070 ;
  assign n6072 = \u10_mem_reg[1][25]/P0001  & ~n6032 ;
  assign n6073 = n5718 & n6032 ;
  assign n6074 = ~n6072 & ~n6073 ;
  assign n6075 = \u10_mem_reg[1][26]/P0001  & ~n6032 ;
  assign n6076 = n5722 & n6032 ;
  assign n6077 = ~n6075 & ~n6076 ;
  assign n6078 = \u10_mem_reg[1][27]/P0001  & ~n6032 ;
  assign n6079 = n5726 & n6032 ;
  assign n6080 = ~n6078 & ~n6079 ;
  assign n6081 = \u10_mem_reg[1][28]/P0001  & ~n6032 ;
  assign n6082 = n5730 & n6032 ;
  assign n6083 = ~n6081 & ~n6082 ;
  assign n6084 = \u10_mem_reg[1][29]/P0001  & ~n6032 ;
  assign n6085 = n5749 & n6032 ;
  assign n6086 = ~n6084 & ~n6085 ;
  assign n6087 = n3068 & ~n5938 ;
  assign n6088 = \u11_mem_reg[3][18]/P0001  & ~n3068 ;
  assign n6089 = ~n6087 & ~n6088 ;
  assign n6090 = n3068 & ~n5944 ;
  assign n6091 = \u11_mem_reg[3][19]/P0001  & ~n3068 ;
  assign n6092 = ~n6090 & ~n6091 ;
  assign n6093 = \u11_mem_reg[3][20]/P0001  & ~n3068 ;
  assign n6094 = n3068 & n5959 ;
  assign n6095 = ~n6093 & ~n6094 ;
  assign n6096 = \u10_mem_reg[1][30]/P0001  & ~n6032 ;
  assign n6097 = n5793 & n6032 ;
  assign n6098 = ~n6096 & ~n6097 ;
  assign n6099 = \u11_mem_reg[3][21]/P0001  & ~n3068 ;
  assign n6100 = n3068 & n5963 ;
  assign n6101 = ~n6099 & ~n6100 ;
  assign n6102 = \u11_mem_reg[3][22]/P0001  & ~n3068 ;
  assign n6103 = n3068 & n5967 ;
  assign n6104 = ~n6102 & ~n6103 ;
  assign n6105 = \u10_mem_reg[1][31]/P0001  & ~n6032 ;
  assign n6106 = n5797 & n6032 ;
  assign n6107 = ~n6105 & ~n6106 ;
  assign n6108 = \u11_mem_reg[3][23]/P0001  & ~n3068 ;
  assign n6109 = n3068 & n5971 ;
  assign n6110 = ~n6108 & ~n6109 ;
  assign n6111 = \u11_mem_reg[3][24]/P0001  & ~n3068 ;
  assign n6112 = n3068 & n5975 ;
  assign n6113 = ~n6111 & ~n6112 ;
  assign n6114 = \u11_mem_reg[3][25]/P0001  & ~n3068 ;
  assign n6115 = n3068 & n5979 ;
  assign n6116 = ~n6114 & ~n6115 ;
  assign n6117 = \u11_mem_reg[3][26]/P0001  & ~n3068 ;
  assign n6118 = n3068 & n5983 ;
  assign n6119 = ~n6117 & ~n6118 ;
  assign n6120 = \u11_mem_reg[3][27]/P0001  & ~n3068 ;
  assign n6121 = n3068 & n5987 ;
  assign n6122 = ~n6120 & ~n6121 ;
  assign n6123 = \u11_mem_reg[3][28]/P0001  & ~n3068 ;
  assign n6124 = n3068 & n5991 ;
  assign n6125 = ~n6123 & ~n6124 ;
  assign n6126 = \u11_mem_reg[3][29]/P0001  & ~n3068 ;
  assign n6127 = n3068 & n5995 ;
  assign n6128 = ~n6126 & ~n6127 ;
  assign n6129 = \u11_mem_reg[3][30]/P0001  & ~n3068 ;
  assign n6130 = n3068 & n5999 ;
  assign n6131 = ~n6129 & ~n6130 ;
  assign n6132 = \u11_mem_reg[3][31]/P0001  & ~n3068 ;
  assign n6133 = n3068 & n6003 ;
  assign n6134 = ~n6132 & ~n6133 ;
  assign n6135 = \u15_valid_r_reg/P0001  & ~\valid_s_reg/NET0131  ;
  assign n6136 = \u15_crac_wr_reg/NET0131  & n6135 ;
  assign n6137 = ~\u13_ints_r_reg[1]/NET0131  & ~n6136 ;
  assign n6138 = ~n2743 & ~n6137 ;
  assign n6139 = \wb_addr_i[5]_pad  & ~\wb_addr_i[6]_pad  ;
  assign n6140 = \wb_addr_i[3]_pad  & \wb_addr_i[4]_pad  ;
  assign n6141 = n6139 & n6140 ;
  assign n6142 = ~\wb_addr_i[2]_pad  & ~\wb_addr_i[3]_pad  ;
  assign n6143 = ~\wb_addr_i[4]_pad  & n6142 ;
  assign n6144 = ~\wb_addr_i[5]_pad  & \wb_addr_i[6]_pad  ;
  assign n6145 = n6143 & n6144 ;
  assign n6146 = ~n6141 & ~n6145 ;
  assign n6159 = \wb_addr_i[4]_pad  & n6142 ;
  assign n6160 = \u15_crac_din_reg[1]/NET0131  & n6159 ;
  assign n6155 = suspended_o_pad & n6143 ;
  assign n6156 = \wb_addr_i[2]_pad  & \wb_addr_i[3]_pad  ;
  assign n6157 = ~\wb_addr_i[4]_pad  & n6156 ;
  assign n6158 = \u13_icc_r_reg[1]/NET0131  & n6157 ;
  assign n6163 = ~n6155 & ~n6158 ;
  assign n6164 = ~n6160 & n6163 ;
  assign n6147 = ~\wb_addr_i[4]_pad  & n2740 ;
  assign n6148 = \u13_occ1_r_reg[1]/NET0131  & n6147 ;
  assign n6149 = \u13_ints_r_reg[1]/NET0131  & n2741 ;
  assign n6161 = ~n6148 & ~n6149 ;
  assign n6150 = \wb_addr_i[2]_pad  & ~\wb_addr_i[3]_pad  ;
  assign n6151 = ~\wb_addr_i[4]_pad  & n6150 ;
  assign n6152 = \u13_occ0_r_reg[1]/NET0131  & n6151 ;
  assign n6153 = \wb_addr_i[4]_pad  & n6150 ;
  assign n6154 = \u13_intm_r_reg[1]/NET0131  & n6153 ;
  assign n6162 = ~n6152 & ~n6154 ;
  assign n6165 = n6161 & n6162 ;
  assign n6166 = n6164 & n6165 ;
  assign n6167 = n6146 & ~n6166 ;
  assign n6172 = \u11_dout_reg[1]/P0001  & n6145 ;
  assign n6168 = ~\wb_addr_i[2]_pad  & n6141 ;
  assign n6169 = \u9_dout_reg[1]/P0001  & n6168 ;
  assign n6170 = \wb_addr_i[2]_pad  & n6141 ;
  assign n6171 = \u10_dout_reg[1]/P0001  & n6170 ;
  assign n6173 = ~n6169 & ~n6171 ;
  assign n6174 = ~n6172 & n6173 ;
  assign n6175 = ~n6167 & n6174 ;
  assign n6177 = ~\u26_cnt_reg[0]/NET0131  & ~\u26_cnt_reg[1]/NET0131  ;
  assign n6178 = \u26_cnt_reg[2]/NET0131  & n6177 ;
  assign n6179 = n5629 & ~n6178 ;
  assign n6180 = ~\u26_cnt_reg[0]/NET0131  & ~n6179 ;
  assign n6176 = \u26_cnt_reg[0]/NET0131  & n5629 ;
  assign n6181 = ~\u13_ac97_rst_force_reg/P0001  & ~n6176 ;
  assign n6182 = ~n6180 & n6181 ;
  assign n6184 = \u26_cnt_reg[1]/NET0131  & n6176 ;
  assign n6183 = ~\u26_cnt_reg[1]/NET0131  & ~n6176 ;
  assign n6185 = ~\u13_ac97_rst_force_reg/P0001  & ~n6183 ;
  assign n6186 = ~n6184 & n6185 ;
  assign n6188 = \u26_cnt_reg[2]/NET0131  & n6184 ;
  assign n6187 = ~\u26_cnt_reg[2]/NET0131  & ~n6184 ;
  assign n6189 = ~\u13_ac97_rst_force_reg/P0001  & ~n6187 ;
  assign n6190 = ~n6188 & n6189 ;
  assign n6191 = \u3_empty_reg/NET0131  & n2787 ;
  assign n6192 = ~\u17_int_set_reg[1]/NET0131  & ~n6191 ;
  assign n6193 = \u4_empty_reg/NET0131  & n2759 ;
  assign n6194 = ~\u18_int_set_reg[1]/NET0131  & ~n6193 ;
  assign n6195 = \u5_empty_reg/NET0131  & n2770 ;
  assign n6196 = ~\u19_int_set_reg[1]/NET0131  & ~n6195 ;
  assign n6197 = \u6_empty_reg/NET0131  & n2795 ;
  assign n6198 = ~\u20_int_set_reg[1]/NET0131  & ~n6197 ;
  assign n6199 = \u7_empty_reg/NET0131  & n2808 ;
  assign n6200 = ~\u21_int_set_reg[1]/NET0131  & ~n6199 ;
  assign n6201 = \u8_empty_reg/NET0131  & n2159 ;
  assign n6202 = ~\u22_int_set_reg[1]/NET0131  & ~n6201 ;
  assign n6203 = \u9_full_reg/NET0131  & n3310 ;
  assign n6204 = ~\u23_int_set_reg[2]/NET0131  & ~n6203 ;
  assign n6205 = \u10_full_reg/NET0131  & n3500 ;
  assign n6206 = ~\u24_int_set_reg[2]/NET0131  & ~n6205 ;
  assign n6207 = \u11_full_reg/NET0131  & n3063 ;
  assign n6208 = ~\u25_int_set_reg[2]/NET0131  & ~n6207 ;
  assign n6209 = ~\ac97_reset_pad_o__pad  & ~n6178 ;
  assign n6210 = ~\u13_ac97_rst_force_reg/P0001  & ~n6209 ;
  assign n6211 = ~\u13_crac_r_reg[7]/NET0131  & \u15_crac_we_r_reg/P0001  ;
  assign n6212 = \u15_crac_wr_reg/NET0131  & ~n6135 ;
  assign n6213 = ~n6211 & ~n6212 ;
  assign n6214 = \u13_crac_r_reg[7]/NET0131  & \u15_crac_we_r_reg/P0001  ;
  assign n6215 = ~\u15_valid_r_reg/P0001  & \valid_s_reg/NET0131  ;
  assign n6216 = \u15_rdd1_reg/NET0131  & n6215 ;
  assign n6217 = \u15_crac_rd_reg/NET0131  & ~n6216 ;
  assign n6218 = ~n6214 & ~n6217 ;
  assign n6219 = \u2_ld_reg/P0001  & \u8_dout_reg[2]/P0001  ;
  assign n6220 = \u0_slt9_r_reg[1]/P0001  & ~\u2_ld_reg/P0001  ;
  assign n6221 = ~n6219 & ~n6220 ;
  assign n6225 = ~\u3_rp_reg[1]/NET0131  & \u3_wp_reg[0]/P0001  ;
  assign n6226 = \u3_rp_reg[2]/NET0131  & ~\u3_wp_reg[1]/NET0131  ;
  assign n6227 = ~\u3_rp_reg[2]/NET0131  & \u3_wp_reg[1]/NET0131  ;
  assign n6228 = ~n6226 & ~n6227 ;
  assign n6229 = ~n6225 & n6228 ;
  assign n6222 = ~\u3_rp_reg[3]/NET0131  & ~\u3_wp_reg[2]/P0001  ;
  assign n6223 = \u3_rp_reg[3]/NET0131  & \u3_wp_reg[2]/P0001  ;
  assign n6224 = ~n6222 & ~n6223 ;
  assign n6230 = \u3_rp_reg[1]/NET0131  & ~\u3_wp_reg[0]/P0001  ;
  assign n6231 = \u12_o3_we_reg/P0001  & ~n6230 ;
  assign n6232 = n6224 & n6231 ;
  assign n6233 = n6229 & n6232 ;
  assign n6234 = ~\u17_int_set_reg[2]/NET0131  & ~n6233 ;
  assign n6236 = ~\u4_rp_reg[1]/NET0131  & \u4_wp_reg[0]/P0001  ;
  assign n6237 = \u4_rp_reg[2]/NET0131  & ~\u4_wp_reg[1]/NET0131  ;
  assign n6238 = ~\u4_rp_reg[2]/NET0131  & \u4_wp_reg[1]/NET0131  ;
  assign n6239 = ~n6237 & ~n6238 ;
  assign n6240 = ~n6236 & n6239 ;
  assign n6241 = ~\u4_rp_reg[3]/NET0131  & ~\u4_wp_reg[2]/P0001  ;
  assign n6242 = \u4_rp_reg[3]/NET0131  & \u4_wp_reg[2]/P0001  ;
  assign n6243 = ~n6241 & ~n6242 ;
  assign n6235 = \u4_rp_reg[1]/NET0131  & ~\u4_wp_reg[0]/P0001  ;
  assign n6244 = \u12_o4_we_reg/P0001  & ~n6235 ;
  assign n6245 = n6243 & n6244 ;
  assign n6246 = n6240 & n6245 ;
  assign n6247 = ~\u18_int_set_reg[2]/NET0131  & ~n6246 ;
  assign n6249 = ~\u5_rp_reg[1]/NET0131  & \u5_wp_reg[0]/P0001  ;
  assign n6250 = \u5_rp_reg[2]/NET0131  & ~\u5_wp_reg[1]/NET0131  ;
  assign n6251 = ~\u5_rp_reg[2]/NET0131  & \u5_wp_reg[1]/NET0131  ;
  assign n6252 = ~n6250 & ~n6251 ;
  assign n6253 = ~n6249 & n6252 ;
  assign n6254 = ~\u5_rp_reg[3]/NET0131  & ~\u5_wp_reg[2]/P0001  ;
  assign n6255 = \u5_rp_reg[3]/NET0131  & \u5_wp_reg[2]/P0001  ;
  assign n6256 = ~n6254 & ~n6255 ;
  assign n6248 = \u5_rp_reg[1]/NET0131  & ~\u5_wp_reg[0]/P0001  ;
  assign n6257 = \u12_o6_we_reg/P0001  & ~n6248 ;
  assign n6258 = n6256 & n6257 ;
  assign n6259 = n6253 & n6258 ;
  assign n6260 = ~\u19_int_set_reg[2]/NET0131  & ~n6259 ;
  assign n6261 = ~\u6_rp_reg[1]/NET0131  & \u6_wp_reg[0]/P0001  ;
  assign n6262 = \u6_rp_reg[1]/NET0131  & ~\u6_wp_reg[0]/P0001  ;
  assign n6263 = ~n6261 & ~n6262 ;
  assign n6264 = \u6_rp_reg[2]/NET0131  & ~\u6_wp_reg[1]/NET0131  ;
  assign n6265 = ~\u6_rp_reg[2]/NET0131  & \u6_wp_reg[1]/NET0131  ;
  assign n6266 = ~n6264 & ~n6265 ;
  assign n6267 = n6263 & n6266 ;
  assign n6268 = ~\u6_rp_reg[3]/NET0131  & ~\u6_wp_reg[2]/P0001  ;
  assign n6269 = \u6_rp_reg[3]/NET0131  & \u6_wp_reg[2]/P0001  ;
  assign n6270 = ~n6268 & ~n6269 ;
  assign n6271 = \u12_o7_we_reg/P0001  & n6270 ;
  assign n6272 = n6267 & n6271 ;
  assign n6273 = ~\u20_int_set_reg[2]/NET0131  & ~n6272 ;
  assign n6277 = ~\u7_rp_reg[1]/NET0131  & \u7_wp_reg[0]/P0001  ;
  assign n6278 = \u7_rp_reg[2]/NET0131  & ~\u7_wp_reg[1]/NET0131  ;
  assign n6279 = ~\u7_rp_reg[2]/NET0131  & \u7_wp_reg[1]/NET0131  ;
  assign n6280 = ~n6278 & ~n6279 ;
  assign n6281 = ~n6277 & n6280 ;
  assign n6274 = ~\u7_rp_reg[3]/NET0131  & ~\u7_wp_reg[2]/P0001  ;
  assign n6275 = \u7_rp_reg[3]/NET0131  & \u7_wp_reg[2]/P0001  ;
  assign n6276 = ~n6274 & ~n6275 ;
  assign n6282 = \u7_rp_reg[1]/NET0131  & ~\u7_wp_reg[0]/P0001  ;
  assign n6283 = \u12_o8_we_reg/P0001  & ~n6282 ;
  assign n6284 = n6276 & n6283 ;
  assign n6285 = n6281 & n6284 ;
  assign n6286 = ~\u21_int_set_reg[2]/NET0131  & ~n6285 ;
  assign n6287 = ~\u8_rp_reg[1]/NET0131  & \u8_wp_reg[0]/P0001  ;
  assign n6288 = \u8_rp_reg[1]/NET0131  & ~\u8_wp_reg[0]/P0001  ;
  assign n6289 = ~n6287 & ~n6288 ;
  assign n6290 = \u8_rp_reg[2]/NET0131  & ~\u8_wp_reg[1]/NET0131  ;
  assign n6291 = ~\u8_rp_reg[2]/NET0131  & \u8_wp_reg[1]/NET0131  ;
  assign n6292 = ~n6290 & ~n6291 ;
  assign n6293 = n6289 & n6292 ;
  assign n6294 = ~\u8_rp_reg[3]/NET0131  & ~\u8_wp_reg[2]/P0001  ;
  assign n6295 = \u8_rp_reg[3]/NET0131  & \u8_wp_reg[2]/P0001  ;
  assign n6296 = ~n6294 & ~n6295 ;
  assign n6297 = \u12_o9_we_reg/P0001  & n6296 ;
  assign n6298 = n6293 & n6297 ;
  assign n6299 = ~\u22_int_set_reg[2]/NET0131  & ~n6298 ;
  assign n6300 = \u12_o9_we_reg/P0001  & \u8_wp_reg[0]/P0001  ;
  assign n6301 = \u8_wp_reg[1]/NET0131  & n6300 ;
  assign n6303 = \u8_wp_reg[2]/P0001  & n6301 ;
  assign n6302 = ~\u8_wp_reg[2]/P0001  & ~n6301 ;
  assign n6304 = \u13_occ1_r_reg[8]/NET0131  & ~n6302 ;
  assign n6305 = ~n6303 & n6304 ;
  assign n6306 = \u12_o4_we_reg/P0001  & \u4_wp_reg[0]/P0001  ;
  assign n6307 = \u4_wp_reg[1]/NET0131  & n6306 ;
  assign n6309 = \u4_wp_reg[2]/P0001  & n6307 ;
  assign n6308 = ~\u4_wp_reg[2]/P0001  & ~n6307 ;
  assign n6310 = \u13_occ0_r_reg[8]/NET0131  & ~n6308 ;
  assign n6311 = ~n6309 & n6310 ;
  assign n6312 = \u12_o6_we_reg/P0001  & \u5_wp_reg[0]/P0001  ;
  assign n6313 = \u5_wp_reg[1]/NET0131  & n6312 ;
  assign n6315 = \u5_wp_reg[2]/P0001  & n6313 ;
  assign n6314 = ~\u5_wp_reg[2]/P0001  & ~n6313 ;
  assign n6316 = \u13_occ0_r_reg[16]/NET0131  & ~n6314 ;
  assign n6317 = ~n6315 & n6316 ;
  assign n6318 = \u12_o3_we_reg/P0001  & \u3_wp_reg[0]/P0001  ;
  assign n6319 = \u3_wp_reg[1]/NET0131  & n6318 ;
  assign n6321 = \u3_wp_reg[2]/P0001  & n6319 ;
  assign n6320 = ~\u3_wp_reg[2]/P0001  & ~n6319 ;
  assign n6322 = \u13_occ0_r_reg[0]/NET0131  & ~n6320 ;
  assign n6323 = ~n6321 & n6322 ;
  assign n6324 = \u12_o7_we_reg/P0001  & \u6_wp_reg[0]/P0001  ;
  assign n6325 = \u6_wp_reg[1]/NET0131  & n6324 ;
  assign n6327 = \u6_wp_reg[2]/P0001  & n6325 ;
  assign n6326 = ~\u6_wp_reg[2]/P0001  & ~n6325 ;
  assign n6328 = \u13_occ0_r_reg[24]/NET0131  & ~n6326 ;
  assign n6329 = ~n6327 & n6328 ;
  assign n6330 = \u12_o8_we_reg/P0001  & \u7_wp_reg[0]/P0001  ;
  assign n6331 = \u7_wp_reg[1]/NET0131  & n6330 ;
  assign n6333 = \u7_wp_reg[2]/P0001  & n6331 ;
  assign n6332 = ~\u7_wp_reg[2]/P0001  & ~n6331 ;
  assign n6334 = \u13_occ1_r_reg[0]/NET0131  & ~n6332 ;
  assign n6335 = ~n6333 & n6334 ;
  assign n6336 = ~\u11_wp_reg[0]/NET0131  & n3063 ;
  assign n6337 = ~\u9_wp_reg[0]/NET0131  & n3310 ;
  assign n6338 = ~\u10_wp_reg[0]/NET0131  & n3500 ;
  assign n6339 = \u14_u0_en_out_l_reg/NET0131  & \valid_s_reg/NET0131  ;
  assign n6342 = \u13_occ0_r_reg[0]/NET0131  & ~\u14_u0_full_empty_r_reg/P0001  ;
  assign n6343 = \u1_slt0_reg[15]/P0001  & n6342 ;
  assign n6340 = ~\u14_u0_en_out_l_reg/NET0131  & ~\valid_s_reg/NET0131  ;
  assign n6341 = \u13_occ0_r_reg[1]/NET0131  & \u1_slt1_reg[11]/P0001  ;
  assign n6344 = ~n6340 & ~n6341 ;
  assign n6345 = n6343 & n6344 ;
  assign n6346 = ~n6339 & ~n6345 ;
  assign n6349 = \u13_occ0_r_reg[8]/NET0131  & ~\u14_u1_full_empty_r_reg/P0001  ;
  assign n6350 = \u1_slt0_reg[15]/P0001  & n6349 ;
  assign n6347 = ~\u14_u1_en_out_l_reg/NET0131  & ~\valid_s_reg/NET0131  ;
  assign n6348 = \u13_occ0_r_reg[9]/NET0131  & \u1_slt1_reg[10]/P0001  ;
  assign n6351 = ~n6347 & ~n6348 ;
  assign n6352 = n6350 & n6351 ;
  assign n6353 = ~n2758 & ~n6352 ;
  assign n6356 = \u13_occ0_r_reg[16]/NET0131  & ~\u14_u2_full_empty_r_reg/P0001  ;
  assign n6357 = \u1_slt0_reg[15]/P0001  & n6356 ;
  assign n6354 = ~\u14_u2_en_out_l_reg/NET0131  & ~\valid_s_reg/NET0131  ;
  assign n6355 = \u13_occ0_r_reg[17]/NET0131  & \u1_slt1_reg[8]/P0001  ;
  assign n6358 = ~n6354 & ~n6355 ;
  assign n6359 = n6357 & n6358 ;
  assign n6360 = ~n2769 & ~n6359 ;
  assign n6363 = \u13_occ0_r_reg[24]/NET0131  & ~\u14_u3_full_empty_r_reg/P0001  ;
  assign n6364 = \u1_slt0_reg[15]/P0001  & n6363 ;
  assign n6361 = ~\u14_u3_en_out_l_reg/NET0131  & ~\valid_s_reg/NET0131  ;
  assign n6362 = \u13_occ0_r_reg[25]/NET0131  & \u1_slt1_reg[7]/P0001  ;
  assign n6365 = ~n6361 & ~n6362 ;
  assign n6366 = n6364 & n6365 ;
  assign n6367 = ~n2794 & ~n6366 ;
  assign n6370 = \u13_occ1_r_reg[0]/NET0131  & ~\u14_u4_full_empty_r_reg/P0001  ;
  assign n6371 = \u1_slt0_reg[15]/P0001  & n6370 ;
  assign n6368 = ~\u14_u4_en_out_l_reg/NET0131  & ~\valid_s_reg/NET0131  ;
  assign n6369 = \u13_occ1_r_reg[1]/NET0131  & \u1_slt1_reg[6]/P0001  ;
  assign n6372 = ~n6368 & ~n6369 ;
  assign n6373 = n6371 & n6372 ;
  assign n6374 = ~n2807 & ~n6373 ;
  assign n6377 = \u13_occ1_r_reg[8]/NET0131  & ~\u14_u5_full_empty_r_reg/P0001  ;
  assign n6378 = \u1_slt0_reg[15]/P0001  & n6377 ;
  assign n6375 = ~\u14_u5_en_out_l_reg/NET0131  & ~\valid_s_reg/NET0131  ;
  assign n6376 = \u13_occ1_r_reg[9]/NET0131  & \u1_slt1_reg[5]/P0001  ;
  assign n6379 = ~n6375 & ~n6376 ;
  assign n6380 = n6378 & n6379 ;
  assign n6381 = ~n2158 & ~n6380 ;
  assign n6384 = \u13_icc_r_reg[0]/NET0131  & ~\u14_u6_full_empty_r_reg/P0001  ;
  assign n6385 = \u1_slt0_reg[15]/P0001  & n6384 ;
  assign n6382 = ~\in_valid_s_reg[0]/NET0131  & ~\u14_u6_en_out_l_reg/NET0131  ;
  assign n6383 = \u13_icc_r_reg[1]/NET0131  & ~\u1_slt0_reg[12]/P0001  ;
  assign n6386 = ~n6382 & ~n6383 ;
  assign n6387 = n6385 & n6386 ;
  assign n6388 = ~n3309 & ~n6387 ;
  assign n6391 = \u13_icc_r_reg[8]/NET0131  & ~\u14_u7_full_empty_r_reg/P0001  ;
  assign n6392 = \u1_slt0_reg[15]/P0001  & n6391 ;
  assign n6389 = ~\in_valid_s_reg[1]/NET0131  & ~\u14_u7_en_out_l_reg/NET0131  ;
  assign n6390 = \u13_icc_r_reg[9]/NET0131  & ~\u1_slt0_reg[11]/P0001  ;
  assign n6393 = ~n6389 & ~n6390 ;
  assign n6394 = n6392 & n6393 ;
  assign n6395 = ~n3499 & ~n6394 ;
  assign n6398 = \u13_icc_r_reg[16]/NET0131  & ~\u14_u8_full_empty_r_reg/P0001  ;
  assign n6399 = \u1_slt0_reg[15]/P0001  & n6398 ;
  assign n6396 = ~\in_valid_s_reg[2]/NET0131  & ~\u14_u8_en_out_l_reg/NET0131  ;
  assign n6397 = \u13_icc_r_reg[17]/NET0131  & ~\u1_slt0_reg[9]/P0001  ;
  assign n6400 = ~n6396 & ~n6397 ;
  assign n6401 = n6399 & n6400 ;
  assign n6402 = ~n3062 & ~n6401 ;
  assign n6403 = \u12_o9_we_reg/P0001  & ~\u8_wp_reg[0]/P0001  ;
  assign n6404 = ~\u12_o9_we_reg/P0001  & \u8_wp_reg[0]/P0001  ;
  assign n6405 = ~n6403 & ~n6404 ;
  assign n6406 = \u13_occ1_r_reg[8]/NET0131  & ~n6405 ;
  assign n6407 = \u12_o3_we_reg/P0001  & ~\u3_wp_reg[0]/P0001  ;
  assign n6408 = ~\u12_o3_we_reg/P0001  & \u3_wp_reg[0]/P0001  ;
  assign n6409 = ~n6407 & ~n6408 ;
  assign n6410 = \u13_occ0_r_reg[0]/NET0131  & ~n6409 ;
  assign n6411 = \u12_o4_we_reg/P0001  & ~\u4_wp_reg[0]/P0001  ;
  assign n6412 = ~\u12_o4_we_reg/P0001  & \u4_wp_reg[0]/P0001  ;
  assign n6413 = ~n6411 & ~n6412 ;
  assign n6414 = \u13_occ0_r_reg[8]/NET0131  & ~n6413 ;
  assign n6415 = \u12_o6_we_reg/P0001  & ~\u5_wp_reg[0]/P0001  ;
  assign n6416 = ~\u12_o6_we_reg/P0001  & \u5_wp_reg[0]/P0001  ;
  assign n6417 = ~n6415 & ~n6416 ;
  assign n6418 = \u13_occ0_r_reg[16]/NET0131  & ~n6417 ;
  assign n6419 = \u12_o7_we_reg/P0001  & ~\u6_wp_reg[0]/P0001  ;
  assign n6420 = ~\u12_o7_we_reg/P0001  & \u6_wp_reg[0]/P0001  ;
  assign n6421 = ~n6419 & ~n6420 ;
  assign n6422 = \u13_occ0_r_reg[24]/NET0131  & ~n6421 ;
  assign n6423 = \u12_o8_we_reg/P0001  & ~\u7_wp_reg[0]/P0001  ;
  assign n6424 = ~\u12_o8_we_reg/P0001  & \u7_wp_reg[0]/P0001  ;
  assign n6425 = ~n6423 & ~n6424 ;
  assign n6426 = \u13_occ1_r_reg[0]/NET0131  & ~n6425 ;
  assign n6427 = ~\u8_wp_reg[1]/NET0131  & ~n6300 ;
  assign n6428 = \u13_occ1_r_reg[8]/NET0131  & ~n6301 ;
  assign n6429 = ~n6427 & n6428 ;
  assign n6430 = ~\u4_wp_reg[1]/NET0131  & ~n6306 ;
  assign n6431 = \u13_occ0_r_reg[8]/NET0131  & ~n6307 ;
  assign n6432 = ~n6430 & n6431 ;
  assign n6433 = ~\u5_wp_reg[1]/NET0131  & ~n6312 ;
  assign n6434 = \u13_occ0_r_reg[16]/NET0131  & ~n6313 ;
  assign n6435 = ~n6433 & n6434 ;
  assign n6436 = ~\u3_wp_reg[1]/NET0131  & ~n6318 ;
  assign n6437 = \u13_occ0_r_reg[0]/NET0131  & ~n6319 ;
  assign n6438 = ~n6436 & n6437 ;
  assign n6439 = ~\u6_wp_reg[1]/NET0131  & ~n6324 ;
  assign n6440 = \u13_occ0_r_reg[24]/NET0131  & ~n6325 ;
  assign n6441 = ~n6439 & n6440 ;
  assign n6442 = ~\u7_wp_reg[1]/NET0131  & ~n6330 ;
  assign n6443 = \u13_occ1_r_reg[0]/NET0131  & ~n6331 ;
  assign n6444 = ~n6442 & n6443 ;
  assign n6445 = ~\u15_rdd1_reg/NET0131  & ~n6135 ;
  assign n6446 = \u15_crac_rd_reg/NET0131  & ~n6445 ;
  assign n6447 = \u15_crac_rd_reg/NET0131  & n6135 ;
  assign n6448 = \u15_crac_rd_done_reg/P0001  & \u15_rdd3_reg/NET0131  ;
  assign n6449 = \u15_rdd2_reg/NET0131  & ~n6448 ;
  assign n6450 = ~n6447 & ~n6449 ;
  assign n6451 = \u15_rdd2_reg/NET0131  & n6215 ;
  assign n6452 = ~\u15_crac_rd_done_reg/P0001  & \u15_rdd3_reg/NET0131  ;
  assign n6453 = ~n6451 & ~n6452 ;
  assign n6454 = \u2_res_cnt_reg[0]/P0001  & n5629 ;
  assign n6455 = \u2_res_cnt_reg[1]/P0001  & n6454 ;
  assign n6456 = \u2_res_cnt_reg[2]/P0001  & n6455 ;
  assign n6458 = \u2_res_cnt_reg[3]/P0001  & n6456 ;
  assign n6457 = ~\u2_res_cnt_reg[3]/P0001  & ~n6456 ;
  assign n6459 = \u2_sync_resume_reg/NET0131  & ~n6457 ;
  assign n6460 = ~n6458 & n6459 ;
  assign n6461 = \u12_rf_we_reg/P0001  & n6143 ;
  assign n6462 = \u12_dout_reg[0]/P0001  & n6461 ;
  assign n6463 = \u12_dout_reg[1]/P0001  & n6461 ;
  assign n6464 = ~\u14_crac_valid_r_reg/P0001  & ~\valid_s_reg/NET0131  ;
  assign n6465 = ~\u15_crac_wr_reg/NET0131  & \valid_s_reg/NET0131  ;
  assign n6466 = ~\u15_crac_rd_reg/NET0131  & n6465 ;
  assign n6467 = ~n6464 & ~n6466 ;
  assign n6468 = \u15_rdd3_reg/NET0131  & n6215 ;
  assign n6469 = \u2_cnt_reg[0]/NET0131  & \u2_cnt_reg[1]/NET0131  ;
  assign n6470 = \u2_cnt_reg[2]/NET0131  & n6469 ;
  assign n6471 = \u2_cnt_reg[3]/NET0131  & n6470 ;
  assign n6472 = \u2_cnt_reg[4]/NET0131  & n6471 ;
  assign n6473 = \u2_cnt_reg[5]/NET0131  & \u2_cnt_reg[6]/NET0131  ;
  assign n6474 = n6472 & n6473 ;
  assign n6476 = ~\u2_cnt_reg[7]/NET0131  & n6474 ;
  assign n6475 = \u2_cnt_reg[7]/NET0131  & ~n6474 ;
  assign n6477 = ~suspended_o_pad & ~n6475 ;
  assign n6478 = ~n6476 & n6477 ;
  assign n6479 = \u2_to_cnt_reg[0]/NET0131  & \u2_to_cnt_reg[1]/NET0131  ;
  assign n6480 = \u2_to_cnt_reg[2]/NET0131  & n6479 ;
  assign n6482 = ~\u2_to_cnt_reg[3]/NET0131  & ~n6480 ;
  assign n6481 = \u2_to_cnt_reg[3]/NET0131  & n6480 ;
  assign n6483 = ~\u2_bit_clk_e_reg/P0001  & ~n6481 ;
  assign n6484 = ~n6482 & n6483 ;
  assign n6485 = \u8_wp_reg[1]/NET0131  & n6403 ;
  assign n6486 = \u8_mem_reg[2][5]/NET0131  & ~n6485 ;
  assign n6487 = \u12_dout_reg[5]/P0001  & n6485 ;
  assign n6488 = ~n6486 & ~n6487 ;
  assign n6489 = ~\u3_wp_reg[1]/NET0131  & n6318 ;
  assign n6490 = \u3_mem_reg[1][29]/NET0131  & ~n6489 ;
  assign n6491 = \u12_dout_reg[29]/P0001  & n6489 ;
  assign n6492 = ~n6490 & ~n6491 ;
  assign n6493 = \u8_mem_reg[2][6]/NET0131  & ~n6485 ;
  assign n6494 = \u12_dout_reg[6]/P0001  & n6485 ;
  assign n6495 = ~n6493 & ~n6494 ;
  assign n6496 = \u8_mem_reg[2][7]/NET0131  & ~n6485 ;
  assign n6497 = \u12_dout_reg[7]/P0001  & n6485 ;
  assign n6498 = ~n6496 & ~n6497 ;
  assign n6499 = \u3_mem_reg[1][2]/NET0131  & ~n6489 ;
  assign n6500 = \u12_dout_reg[2]/P0001  & n6489 ;
  assign n6501 = ~n6499 & ~n6500 ;
  assign n6502 = \u8_mem_reg[2][8]/NET0131  & ~n6485 ;
  assign n6503 = \u12_dout_reg[8]/P0001  & n6485 ;
  assign n6504 = ~n6502 & ~n6503 ;
  assign n6505 = \u8_mem_reg[2][9]/NET0131  & ~n6485 ;
  assign n6506 = \u12_dout_reg[9]/P0001  & n6485 ;
  assign n6507 = ~n6505 & ~n6506 ;
  assign n6508 = \u8_mem_reg[3][19]/NET0131  & ~n6301 ;
  assign n6509 = \u12_dout_reg[19]/P0001  & n6301 ;
  assign n6510 = ~n6508 & ~n6509 ;
  assign n6511 = \u8_mem_reg[3][0]/NET0131  & ~n6301 ;
  assign n6512 = \u12_dout_reg[0]/P0001  & n6301 ;
  assign n6513 = ~n6511 & ~n6512 ;
  assign n6514 = \u8_mem_reg[3][10]/NET0131  & ~n6301 ;
  assign n6515 = \u12_dout_reg[10]/P0001  & n6301 ;
  assign n6516 = ~n6514 & ~n6515 ;
  assign n6517 = \u3_mem_reg[1][31]/NET0131  & ~n6489 ;
  assign n6518 = \u12_dout_reg[31]/P0001  & n6489 ;
  assign n6519 = ~n6517 & ~n6518 ;
  assign n6520 = \u8_mem_reg[3][12]/NET0131  & ~n6301 ;
  assign n6521 = \u12_dout_reg[12]/P0001  & n6301 ;
  assign n6522 = ~n6520 & ~n6521 ;
  assign n6523 = \u3_mem_reg[1][3]/NET0131  & ~n6489 ;
  assign n6524 = \u12_dout_reg[3]/P0001  & n6489 ;
  assign n6525 = ~n6523 & ~n6524 ;
  assign n6526 = \u8_mem_reg[3][13]/NET0131  & ~n6301 ;
  assign n6527 = \u12_dout_reg[13]/P0001  & n6301 ;
  assign n6528 = ~n6526 & ~n6527 ;
  assign n6529 = \u8_mem_reg[3][14]/NET0131  & ~n6301 ;
  assign n6530 = \u12_dout_reg[14]/P0001  & n6301 ;
  assign n6531 = ~n6529 & ~n6530 ;
  assign n6532 = \u8_mem_reg[3][15]/NET0131  & ~n6301 ;
  assign n6533 = \u12_dout_reg[15]/P0001  & n6301 ;
  assign n6534 = ~n6532 & ~n6533 ;
  assign n6535 = \u3_mem_reg[1][4]/NET0131  & ~n6489 ;
  assign n6536 = \u12_dout_reg[4]/P0001  & n6489 ;
  assign n6537 = ~n6535 & ~n6536 ;
  assign n6538 = \u8_mem_reg[3][16]/NET0131  & ~n6301 ;
  assign n6539 = \u12_dout_reg[16]/P0001  & n6301 ;
  assign n6540 = ~n6538 & ~n6539 ;
  assign n6541 = \u3_mem_reg[1][5]/NET0131  & ~n6489 ;
  assign n6542 = \u12_dout_reg[5]/P0001  & n6489 ;
  assign n6543 = ~n6541 & ~n6542 ;
  assign n6544 = \u8_mem_reg[3][17]/NET0131  & ~n6301 ;
  assign n6545 = \u12_dout_reg[17]/P0001  & n6301 ;
  assign n6546 = ~n6544 & ~n6545 ;
  assign n6547 = \u8_mem_reg[3][18]/NET0131  & ~n6301 ;
  assign n6548 = \u12_dout_reg[18]/P0001  & n6301 ;
  assign n6549 = ~n6547 & ~n6548 ;
  assign n6550 = \u3_mem_reg[1][6]/NET0131  & ~n6489 ;
  assign n6551 = \u12_dout_reg[6]/P0001  & n6489 ;
  assign n6552 = ~n6550 & ~n6551 ;
  assign n6553 = \u8_mem_reg[3][1]/NET0131  & ~n6301 ;
  assign n6554 = \u12_dout_reg[1]/P0001  & n6301 ;
  assign n6555 = ~n6553 & ~n6554 ;
  assign n6556 = \u3_mem_reg[1][7]/NET0131  & ~n6489 ;
  assign n6557 = \u12_dout_reg[7]/P0001  & n6489 ;
  assign n6558 = ~n6556 & ~n6557 ;
  assign n6559 = \u8_mem_reg[3][20]/NET0131  & ~n6301 ;
  assign n6560 = \u12_dout_reg[20]/P0001  & n6301 ;
  assign n6561 = ~n6559 & ~n6560 ;
  assign n6562 = \u8_mem_reg[3][21]/NET0131  & ~n6301 ;
  assign n6563 = \u12_dout_reg[21]/P0001  & n6301 ;
  assign n6564 = ~n6562 & ~n6563 ;
  assign n6565 = \u3_mem_reg[1][8]/NET0131  & ~n6489 ;
  assign n6566 = \u12_dout_reg[8]/P0001  & n6489 ;
  assign n6567 = ~n6565 & ~n6566 ;
  assign n6568 = \u8_mem_reg[3][22]/NET0131  & ~n6301 ;
  assign n6569 = \u12_dout_reg[22]/P0001  & n6301 ;
  assign n6570 = ~n6568 & ~n6569 ;
  assign n6571 = \u8_mem_reg[3][23]/NET0131  & ~n6301 ;
  assign n6572 = \u12_dout_reg[23]/P0001  & n6301 ;
  assign n6573 = ~n6571 & ~n6572 ;
  assign n6574 = \u3_mem_reg[1][9]/NET0131  & ~n6489 ;
  assign n6575 = \u12_dout_reg[9]/P0001  & n6489 ;
  assign n6576 = ~n6574 & ~n6575 ;
  assign n6577 = \u8_mem_reg[3][24]/NET0131  & ~n6301 ;
  assign n6578 = \u12_dout_reg[24]/P0001  & n6301 ;
  assign n6579 = ~n6577 & ~n6578 ;
  assign n6580 = \u8_mem_reg[3][25]/NET0131  & ~n6301 ;
  assign n6581 = \u12_dout_reg[25]/P0001  & n6301 ;
  assign n6582 = ~n6580 & ~n6581 ;
  assign n6583 = \u3_wp_reg[1]/NET0131  & n6407 ;
  assign n6584 = \u3_mem_reg[2][0]/NET0131  & ~n6583 ;
  assign n6585 = \u12_dout_reg[0]/P0001  & n6583 ;
  assign n6586 = ~n6584 & ~n6585 ;
  assign n6587 = \u8_mem_reg[3][27]/NET0131  & ~n6301 ;
  assign n6588 = \u12_dout_reg[27]/P0001  & n6301 ;
  assign n6589 = ~n6587 & ~n6588 ;
  assign n6590 = \u3_mem_reg[2][10]/NET0131  & ~n6583 ;
  assign n6591 = \u12_dout_reg[10]/P0001  & n6583 ;
  assign n6592 = ~n6590 & ~n6591 ;
  assign n6593 = \u8_mem_reg[3][29]/NET0131  & ~n6301 ;
  assign n6594 = \u12_dout_reg[29]/P0001  & n6301 ;
  assign n6595 = ~n6593 & ~n6594 ;
  assign n6596 = \u3_mem_reg[2][11]/NET0131  & ~n6583 ;
  assign n6597 = \u12_dout_reg[11]/P0001  & n6583 ;
  assign n6598 = ~n6596 & ~n6597 ;
  assign n6599 = \u8_mem_reg[3][2]/NET0131  & ~n6301 ;
  assign n6600 = \u12_dout_reg[2]/P0001  & n6301 ;
  assign n6601 = ~n6599 & ~n6600 ;
  assign n6602 = \u8_mem_reg[3][30]/NET0131  & ~n6301 ;
  assign n6603 = \u12_dout_reg[30]/P0001  & n6301 ;
  assign n6604 = ~n6602 & ~n6603 ;
  assign n6605 = \u3_mem_reg[2][12]/NET0131  & ~n6583 ;
  assign n6606 = \u12_dout_reg[12]/P0001  & n6583 ;
  assign n6607 = ~n6605 & ~n6606 ;
  assign n6608 = \u8_mem_reg[3][3]/NET0131  & ~n6301 ;
  assign n6609 = \u12_dout_reg[3]/P0001  & n6301 ;
  assign n6610 = ~n6608 & ~n6609 ;
  assign n6611 = \u3_mem_reg[2][13]/NET0131  & ~n6583 ;
  assign n6612 = \u12_dout_reg[13]/P0001  & n6583 ;
  assign n6613 = ~n6611 & ~n6612 ;
  assign n6614 = \u8_mem_reg[3][5]/NET0131  & ~n6301 ;
  assign n6615 = \u12_dout_reg[5]/P0001  & n6301 ;
  assign n6616 = ~n6614 & ~n6615 ;
  assign n6617 = \u8_mem_reg[3][7]/NET0131  & ~n6301 ;
  assign n6618 = \u12_dout_reg[7]/P0001  & n6301 ;
  assign n6619 = ~n6617 & ~n6618 ;
  assign n6620 = \u3_mem_reg[2][15]/NET0131  & ~n6583 ;
  assign n6621 = \u12_dout_reg[15]/P0001  & n6583 ;
  assign n6622 = ~n6620 & ~n6621 ;
  assign n6623 = \u8_mem_reg[3][9]/NET0131  & ~n6301 ;
  assign n6624 = \u12_dout_reg[9]/P0001  & n6301 ;
  assign n6625 = ~n6623 & ~n6624 ;
  assign n6626 = \u3_mem_reg[2][16]/NET0131  & ~n6583 ;
  assign n6627 = \u12_dout_reg[16]/P0001  & n6583 ;
  assign n6628 = ~n6626 & ~n6627 ;
  assign n6629 = ~\u8_wp_reg[1]/NET0131  & n6300 ;
  assign n6630 = \u8_mem_reg[1][4]/NET0131  & ~n6629 ;
  assign n6631 = \u12_dout_reg[4]/P0001  & n6629 ;
  assign n6632 = ~n6630 & ~n6631 ;
  assign n6633 = \u3_mem_reg[2][18]/NET0131  & ~n6583 ;
  assign n6634 = \u12_dout_reg[18]/P0001  & n6583 ;
  assign n6635 = ~n6633 & ~n6634 ;
  assign n6636 = \u3_mem_reg[2][19]/NET0131  & ~n6583 ;
  assign n6637 = \u12_dout_reg[19]/P0001  & n6583 ;
  assign n6638 = ~n6636 & ~n6637 ;
  assign n6639 = \u3_mem_reg[2][1]/NET0131  & ~n6583 ;
  assign n6640 = \u12_dout_reg[1]/P0001  & n6583 ;
  assign n6641 = ~n6639 & ~n6640 ;
  assign n6642 = \u3_mem_reg[1][30]/NET0131  & ~n6489 ;
  assign n6643 = \u12_dout_reg[30]/P0001  & n6489 ;
  assign n6644 = ~n6642 & ~n6643 ;
  assign n6645 = \u3_mem_reg[2][21]/NET0131  & ~n6583 ;
  assign n6646 = \u12_dout_reg[21]/P0001  & n6583 ;
  assign n6647 = ~n6645 & ~n6646 ;
  assign n6648 = \u3_mem_reg[2][22]/NET0131  & ~n6583 ;
  assign n6649 = \u12_dout_reg[22]/P0001  & n6583 ;
  assign n6650 = ~n6648 & ~n6649 ;
  assign n6651 = \u3_mem_reg[2][24]/NET0131  & ~n6583 ;
  assign n6652 = \u12_dout_reg[24]/P0001  & n6583 ;
  assign n6653 = ~n6651 & ~n6652 ;
  assign n6654 = \u3_mem_reg[2][26]/NET0131  & ~n6583 ;
  assign n6655 = \u12_dout_reg[26]/P0001  & n6583 ;
  assign n6656 = ~n6654 & ~n6655 ;
  assign n6657 = \u3_mem_reg[2][27]/NET0131  & ~n6583 ;
  assign n6658 = \u12_dout_reg[27]/P0001  & n6583 ;
  assign n6659 = ~n6657 & ~n6658 ;
  assign n6660 = \u3_mem_reg[2][28]/NET0131  & ~n6583 ;
  assign n6661 = \u12_dout_reg[28]/P0001  & n6583 ;
  assign n6662 = ~n6660 & ~n6661 ;
  assign n6663 = \u3_mem_reg[2][29]/NET0131  & ~n6583 ;
  assign n6664 = \u12_dout_reg[29]/P0001  & n6583 ;
  assign n6665 = ~n6663 & ~n6664 ;
  assign n6666 = \u3_mem_reg[2][2]/NET0131  & ~n6583 ;
  assign n6667 = \u12_dout_reg[2]/P0001  & n6583 ;
  assign n6668 = ~n6666 & ~n6667 ;
  assign n6669 = \u3_mem_reg[2][30]/NET0131  & ~n6583 ;
  assign n6670 = \u12_dout_reg[30]/P0001  & n6583 ;
  assign n6671 = ~n6669 & ~n6670 ;
  assign n6672 = \u3_mem_reg[2][31]/NET0131  & ~n6583 ;
  assign n6673 = \u12_dout_reg[31]/P0001  & n6583 ;
  assign n6674 = ~n6672 & ~n6673 ;
  assign n6675 = \u3_mem_reg[2][3]/NET0131  & ~n6583 ;
  assign n6676 = \u12_dout_reg[3]/P0001  & n6583 ;
  assign n6677 = ~n6675 & ~n6676 ;
  assign n6678 = \u3_mem_reg[2][4]/NET0131  & ~n6583 ;
  assign n6679 = \u12_dout_reg[4]/P0001  & n6583 ;
  assign n6680 = ~n6678 & ~n6679 ;
  assign n6681 = \u3_mem_reg[2][5]/NET0131  & ~n6583 ;
  assign n6682 = \u12_dout_reg[5]/P0001  & n6583 ;
  assign n6683 = ~n6681 & ~n6682 ;
  assign n6684 = \u3_mem_reg[2][6]/NET0131  & ~n6583 ;
  assign n6685 = \u12_dout_reg[6]/P0001  & n6583 ;
  assign n6686 = ~n6684 & ~n6685 ;
  assign n6687 = \u3_mem_reg[2][7]/NET0131  & ~n6583 ;
  assign n6688 = \u12_dout_reg[7]/P0001  & n6583 ;
  assign n6689 = ~n6687 & ~n6688 ;
  assign n6690 = \u3_mem_reg[2][8]/NET0131  & ~n6583 ;
  assign n6691 = \u12_dout_reg[8]/P0001  & n6583 ;
  assign n6692 = ~n6690 & ~n6691 ;
  assign n6693 = \u3_mem_reg[2][9]/NET0131  & ~n6583 ;
  assign n6694 = \u12_dout_reg[9]/P0001  & n6583 ;
  assign n6695 = ~n6693 & ~n6694 ;
  assign n6696 = \u3_mem_reg[3][0]/NET0131  & ~n6319 ;
  assign n6697 = \u12_dout_reg[0]/P0001  & n6319 ;
  assign n6698 = ~n6696 & ~n6697 ;
  assign n6699 = \u3_mem_reg[3][10]/NET0131  & ~n6319 ;
  assign n6700 = \u12_dout_reg[10]/P0001  & n6319 ;
  assign n6701 = ~n6699 & ~n6700 ;
  assign n6702 = \u3_mem_reg[3][11]/NET0131  & ~n6319 ;
  assign n6703 = \u12_dout_reg[11]/P0001  & n6319 ;
  assign n6704 = ~n6702 & ~n6703 ;
  assign n6705 = \u3_mem_reg[3][12]/NET0131  & ~n6319 ;
  assign n6706 = \u12_dout_reg[12]/P0001  & n6319 ;
  assign n6707 = ~n6705 & ~n6706 ;
  assign n6708 = \u3_mem_reg[3][13]/NET0131  & ~n6319 ;
  assign n6709 = \u12_dout_reg[13]/P0001  & n6319 ;
  assign n6710 = ~n6708 & ~n6709 ;
  assign n6711 = \u3_mem_reg[3][14]/NET0131  & ~n6319 ;
  assign n6712 = \u12_dout_reg[14]/P0001  & n6319 ;
  assign n6713 = ~n6711 & ~n6712 ;
  assign n6714 = \u3_mem_reg[3][15]/NET0131  & ~n6319 ;
  assign n6715 = \u12_dout_reg[15]/P0001  & n6319 ;
  assign n6716 = ~n6714 & ~n6715 ;
  assign n6717 = \u3_mem_reg[3][16]/NET0131  & ~n6319 ;
  assign n6718 = \u12_dout_reg[16]/P0001  & n6319 ;
  assign n6719 = ~n6717 & ~n6718 ;
  assign n6720 = \u3_mem_reg[3][17]/NET0131  & ~n6319 ;
  assign n6721 = \u12_dout_reg[17]/P0001  & n6319 ;
  assign n6722 = ~n6720 & ~n6721 ;
  assign n6723 = \u3_mem_reg[3][18]/NET0131  & ~n6319 ;
  assign n6724 = \u12_dout_reg[18]/P0001  & n6319 ;
  assign n6725 = ~n6723 & ~n6724 ;
  assign n6726 = \u3_mem_reg[3][19]/NET0131  & ~n6319 ;
  assign n6727 = \u12_dout_reg[19]/P0001  & n6319 ;
  assign n6728 = ~n6726 & ~n6727 ;
  assign n6729 = \u3_mem_reg[3][1]/NET0131  & ~n6319 ;
  assign n6730 = \u12_dout_reg[1]/P0001  & n6319 ;
  assign n6731 = ~n6729 & ~n6730 ;
  assign n6732 = \u3_mem_reg[3][21]/NET0131  & ~n6319 ;
  assign n6733 = \u12_dout_reg[21]/P0001  & n6319 ;
  assign n6734 = ~n6732 & ~n6733 ;
  assign n6735 = \u3_mem_reg[3][22]/NET0131  & ~n6319 ;
  assign n6736 = \u12_dout_reg[22]/P0001  & n6319 ;
  assign n6737 = ~n6735 & ~n6736 ;
  assign n6738 = \u3_mem_reg[3][23]/NET0131  & ~n6319 ;
  assign n6739 = \u12_dout_reg[23]/P0001  & n6319 ;
  assign n6740 = ~n6738 & ~n6739 ;
  assign n6741 = \u3_mem_reg[3][24]/NET0131  & ~n6319 ;
  assign n6742 = \u12_dout_reg[24]/P0001  & n6319 ;
  assign n6743 = ~n6741 & ~n6742 ;
  assign n6744 = \u3_mem_reg[3][26]/NET0131  & ~n6319 ;
  assign n6745 = \u12_dout_reg[26]/P0001  & n6319 ;
  assign n6746 = ~n6744 & ~n6745 ;
  assign n6747 = \u3_mem_reg[3][27]/NET0131  & ~n6319 ;
  assign n6748 = \u12_dout_reg[27]/P0001  & n6319 ;
  assign n6749 = ~n6747 & ~n6748 ;
  assign n6750 = \u8_mem_reg[3][28]/NET0131  & ~n6301 ;
  assign n6751 = \u12_dout_reg[28]/P0001  & n6301 ;
  assign n6752 = ~n6750 & ~n6751 ;
  assign n6753 = \u3_mem_reg[3][28]/NET0131  & ~n6319 ;
  assign n6754 = \u12_dout_reg[28]/P0001  & n6319 ;
  assign n6755 = ~n6753 & ~n6754 ;
  assign n6756 = \u3_mem_reg[3][29]/NET0131  & ~n6319 ;
  assign n6757 = \u12_dout_reg[29]/P0001  & n6319 ;
  assign n6758 = ~n6756 & ~n6757 ;
  assign n6759 = \u3_mem_reg[3][2]/NET0131  & ~n6319 ;
  assign n6760 = \u12_dout_reg[2]/P0001  & n6319 ;
  assign n6761 = ~n6759 & ~n6760 ;
  assign n6762 = \u3_mem_reg[3][30]/NET0131  & ~n6319 ;
  assign n6763 = \u12_dout_reg[30]/P0001  & n6319 ;
  assign n6764 = ~n6762 & ~n6763 ;
  assign n6765 = \u3_mem_reg[3][31]/NET0131  & ~n6319 ;
  assign n6766 = \u12_dout_reg[31]/P0001  & n6319 ;
  assign n6767 = ~n6765 & ~n6766 ;
  assign n6768 = \u3_mem_reg[3][4]/NET0131  & ~n6319 ;
  assign n6769 = \u12_dout_reg[4]/P0001  & n6319 ;
  assign n6770 = ~n6768 & ~n6769 ;
  assign n6771 = \u3_mem_reg[3][5]/NET0131  & ~n6319 ;
  assign n6772 = \u12_dout_reg[5]/P0001  & n6319 ;
  assign n6773 = ~n6771 & ~n6772 ;
  assign n6774 = \u3_mem_reg[1][1]/NET0131  & ~n6489 ;
  assign n6775 = \u12_dout_reg[1]/P0001  & n6489 ;
  assign n6776 = ~n6774 & ~n6775 ;
  assign n6777 = \u3_mem_reg[3][6]/NET0131  & ~n6319 ;
  assign n6778 = \u12_dout_reg[6]/P0001  & n6319 ;
  assign n6779 = ~n6777 & ~n6778 ;
  assign n6780 = \u3_mem_reg[3][7]/NET0131  & ~n6319 ;
  assign n6781 = \u12_dout_reg[7]/P0001  & n6319 ;
  assign n6782 = ~n6780 & ~n6781 ;
  assign n6783 = \u3_mem_reg[3][8]/NET0131  & ~n6319 ;
  assign n6784 = \u12_dout_reg[8]/P0001  & n6319 ;
  assign n6785 = ~n6783 & ~n6784 ;
  assign n6786 = \u3_mem_reg[3][9]/NET0131  & ~n6319 ;
  assign n6787 = \u12_dout_reg[9]/P0001  & n6319 ;
  assign n6788 = ~n6786 & ~n6787 ;
  assign n6789 = \u8_mem_reg[1][31]/NET0131  & ~n6629 ;
  assign n6790 = \u12_dout_reg[31]/P0001  & n6629 ;
  assign n6791 = ~n6789 & ~n6790 ;
  assign n6792 = \u8_mem_reg[3][26]/NET0131  & ~n6301 ;
  assign n6793 = \u12_dout_reg[26]/P0001  & n6301 ;
  assign n6794 = ~n6792 & ~n6793 ;
  assign n6795 = \u8_mem_reg[2][3]/NET0131  & ~n6485 ;
  assign n6796 = \u12_dout_reg[3]/P0001  & n6485 ;
  assign n6797 = ~n6795 & ~n6796 ;
  assign n6798 = \u3_mem_reg[3][25]/NET0131  & ~n6319 ;
  assign n6799 = \u12_dout_reg[25]/P0001  & n6319 ;
  assign n6800 = ~n6798 & ~n6799 ;
  assign n6801 = \u3_mem_reg[1][27]/NET0131  & ~n6489 ;
  assign n6802 = \u12_dout_reg[27]/P0001  & n6489 ;
  assign n6803 = ~n6801 & ~n6802 ;
  assign n6804 = \u3_mem_reg[2][23]/NET0131  & ~n6583 ;
  assign n6805 = \u12_dout_reg[23]/P0001  & n6583 ;
  assign n6806 = ~n6804 & ~n6805 ;
  assign n6807 = ~\u4_wp_reg[1]/NET0131  & n6306 ;
  assign n6808 = \u4_mem_reg[1][0]/NET0131  & ~n6807 ;
  assign n6809 = \u12_dout_reg[0]/P0001  & n6807 ;
  assign n6810 = ~n6808 & ~n6809 ;
  assign n6811 = \u4_mem_reg[1][10]/NET0131  & ~n6807 ;
  assign n6812 = \u12_dout_reg[10]/P0001  & n6807 ;
  assign n6813 = ~n6811 & ~n6812 ;
  assign n6814 = \u4_mem_reg[1][11]/NET0131  & ~n6807 ;
  assign n6815 = \u12_dout_reg[11]/P0001  & n6807 ;
  assign n6816 = ~n6814 & ~n6815 ;
  assign n6817 = \u4_mem_reg[1][12]/NET0131  & ~n6807 ;
  assign n6818 = \u12_dout_reg[12]/P0001  & n6807 ;
  assign n6819 = ~n6817 & ~n6818 ;
  assign n6820 = \u4_mem_reg[1][13]/NET0131  & ~n6807 ;
  assign n6821 = \u12_dout_reg[13]/P0001  & n6807 ;
  assign n6822 = ~n6820 & ~n6821 ;
  assign n6823 = \u4_mem_reg[1][14]/NET0131  & ~n6807 ;
  assign n6824 = \u12_dout_reg[14]/P0001  & n6807 ;
  assign n6825 = ~n6823 & ~n6824 ;
  assign n6826 = \u4_mem_reg[1][15]/NET0131  & ~n6807 ;
  assign n6827 = \u12_dout_reg[15]/P0001  & n6807 ;
  assign n6828 = ~n6826 & ~n6827 ;
  assign n6829 = \u4_mem_reg[1][16]/NET0131  & ~n6807 ;
  assign n6830 = \u12_dout_reg[16]/P0001  & n6807 ;
  assign n6831 = ~n6829 & ~n6830 ;
  assign n6832 = \u4_mem_reg[1][17]/NET0131  & ~n6807 ;
  assign n6833 = \u12_dout_reg[17]/P0001  & n6807 ;
  assign n6834 = ~n6832 & ~n6833 ;
  assign n6835 = \u4_mem_reg[1][18]/NET0131  & ~n6807 ;
  assign n6836 = \u12_dout_reg[18]/P0001  & n6807 ;
  assign n6837 = ~n6835 & ~n6836 ;
  assign n6838 = \u4_mem_reg[1][19]/NET0131  & ~n6807 ;
  assign n6839 = \u12_dout_reg[19]/P0001  & n6807 ;
  assign n6840 = ~n6838 & ~n6839 ;
  assign n6841 = \u4_mem_reg[1][1]/NET0131  & ~n6807 ;
  assign n6842 = \u12_dout_reg[1]/P0001  & n6807 ;
  assign n6843 = ~n6841 & ~n6842 ;
  assign n6844 = \u4_mem_reg[1][20]/NET0131  & ~n6807 ;
  assign n6845 = \u12_dout_reg[20]/P0001  & n6807 ;
  assign n6846 = ~n6844 & ~n6845 ;
  assign n6847 = \u4_mem_reg[1][21]/NET0131  & ~n6807 ;
  assign n6848 = \u12_dout_reg[21]/P0001  & n6807 ;
  assign n6849 = ~n6847 & ~n6848 ;
  assign n6850 = \u4_mem_reg[1][22]/NET0131  & ~n6807 ;
  assign n6851 = \u12_dout_reg[22]/P0001  & n6807 ;
  assign n6852 = ~n6850 & ~n6851 ;
  assign n6853 = \u4_mem_reg[1][23]/NET0131  & ~n6807 ;
  assign n6854 = \u12_dout_reg[23]/P0001  & n6807 ;
  assign n6855 = ~n6853 & ~n6854 ;
  assign n6856 = \u4_mem_reg[1][24]/NET0131  & ~n6807 ;
  assign n6857 = \u12_dout_reg[24]/P0001  & n6807 ;
  assign n6858 = ~n6856 & ~n6857 ;
  assign n6859 = \u4_mem_reg[1][25]/NET0131  & ~n6807 ;
  assign n6860 = \u12_dout_reg[25]/P0001  & n6807 ;
  assign n6861 = ~n6859 & ~n6860 ;
  assign n6862 = \u4_mem_reg[1][26]/NET0131  & ~n6807 ;
  assign n6863 = \u12_dout_reg[26]/P0001  & n6807 ;
  assign n6864 = ~n6862 & ~n6863 ;
  assign n6865 = \u4_mem_reg[1][27]/NET0131  & ~n6807 ;
  assign n6866 = \u12_dout_reg[27]/P0001  & n6807 ;
  assign n6867 = ~n6865 & ~n6866 ;
  assign n6868 = \u4_mem_reg[1][28]/NET0131  & ~n6807 ;
  assign n6869 = \u12_dout_reg[28]/P0001  & n6807 ;
  assign n6870 = ~n6868 & ~n6869 ;
  assign n6871 = \u4_mem_reg[1][29]/NET0131  & ~n6807 ;
  assign n6872 = \u12_dout_reg[29]/P0001  & n6807 ;
  assign n6873 = ~n6871 & ~n6872 ;
  assign n6874 = \u4_mem_reg[1][2]/NET0131  & ~n6807 ;
  assign n6875 = \u12_dout_reg[2]/P0001  & n6807 ;
  assign n6876 = ~n6874 & ~n6875 ;
  assign n6877 = \u4_mem_reg[1][30]/NET0131  & ~n6807 ;
  assign n6878 = \u12_dout_reg[30]/P0001  & n6807 ;
  assign n6879 = ~n6877 & ~n6878 ;
  assign n6880 = \u4_mem_reg[1][31]/NET0131  & ~n6807 ;
  assign n6881 = \u12_dout_reg[31]/P0001  & n6807 ;
  assign n6882 = ~n6880 & ~n6881 ;
  assign n6883 = \u4_mem_reg[1][3]/NET0131  & ~n6807 ;
  assign n6884 = \u12_dout_reg[3]/P0001  & n6807 ;
  assign n6885 = ~n6883 & ~n6884 ;
  assign n6886 = \u4_mem_reg[1][4]/NET0131  & ~n6807 ;
  assign n6887 = \u12_dout_reg[4]/P0001  & n6807 ;
  assign n6888 = ~n6886 & ~n6887 ;
  assign n6889 = \u4_mem_reg[1][5]/NET0131  & ~n6807 ;
  assign n6890 = \u12_dout_reg[5]/P0001  & n6807 ;
  assign n6891 = ~n6889 & ~n6890 ;
  assign n6892 = \u4_mem_reg[1][6]/NET0131  & ~n6807 ;
  assign n6893 = \u12_dout_reg[6]/P0001  & n6807 ;
  assign n6894 = ~n6892 & ~n6893 ;
  assign n6895 = \u4_mem_reg[1][7]/NET0131  & ~n6807 ;
  assign n6896 = \u12_dout_reg[7]/P0001  & n6807 ;
  assign n6897 = ~n6895 & ~n6896 ;
  assign n6898 = \u4_mem_reg[1][8]/NET0131  & ~n6807 ;
  assign n6899 = \u12_dout_reg[8]/P0001  & n6807 ;
  assign n6900 = ~n6898 & ~n6899 ;
  assign n6901 = \u4_mem_reg[1][9]/NET0131  & ~n6807 ;
  assign n6902 = \u12_dout_reg[9]/P0001  & n6807 ;
  assign n6903 = ~n6901 & ~n6902 ;
  assign n6904 = \u4_wp_reg[1]/NET0131  & n6411 ;
  assign n6905 = \u4_mem_reg[2][0]/NET0131  & ~n6904 ;
  assign n6906 = \u12_dout_reg[0]/P0001  & n6904 ;
  assign n6907 = ~n6905 & ~n6906 ;
  assign n6908 = \u4_mem_reg[2][10]/NET0131  & ~n6904 ;
  assign n6909 = \u12_dout_reg[10]/P0001  & n6904 ;
  assign n6910 = ~n6908 & ~n6909 ;
  assign n6911 = \u4_mem_reg[2][11]/NET0131  & ~n6904 ;
  assign n6912 = \u12_dout_reg[11]/P0001  & n6904 ;
  assign n6913 = ~n6911 & ~n6912 ;
  assign n6914 = \u4_mem_reg[2][12]/NET0131  & ~n6904 ;
  assign n6915 = \u12_dout_reg[12]/P0001  & n6904 ;
  assign n6916 = ~n6914 & ~n6915 ;
  assign n6917 = \u4_mem_reg[2][13]/NET0131  & ~n6904 ;
  assign n6918 = \u12_dout_reg[13]/P0001  & n6904 ;
  assign n6919 = ~n6917 & ~n6918 ;
  assign n6920 = \u4_mem_reg[2][14]/NET0131  & ~n6904 ;
  assign n6921 = \u12_dout_reg[14]/P0001  & n6904 ;
  assign n6922 = ~n6920 & ~n6921 ;
  assign n6923 = \u4_mem_reg[2][15]/NET0131  & ~n6904 ;
  assign n6924 = \u12_dout_reg[15]/P0001  & n6904 ;
  assign n6925 = ~n6923 & ~n6924 ;
  assign n6926 = \u4_mem_reg[2][16]/NET0131  & ~n6904 ;
  assign n6927 = \u12_dout_reg[16]/P0001  & n6904 ;
  assign n6928 = ~n6926 & ~n6927 ;
  assign n6929 = \u4_mem_reg[2][17]/NET0131  & ~n6904 ;
  assign n6930 = \u12_dout_reg[17]/P0001  & n6904 ;
  assign n6931 = ~n6929 & ~n6930 ;
  assign n6932 = \u4_mem_reg[2][18]/NET0131  & ~n6904 ;
  assign n6933 = \u12_dout_reg[18]/P0001  & n6904 ;
  assign n6934 = ~n6932 & ~n6933 ;
  assign n6935 = \u4_mem_reg[2][19]/NET0131  & ~n6904 ;
  assign n6936 = \u12_dout_reg[19]/P0001  & n6904 ;
  assign n6937 = ~n6935 & ~n6936 ;
  assign n6938 = \u4_mem_reg[2][1]/NET0131  & ~n6904 ;
  assign n6939 = \u12_dout_reg[1]/P0001  & n6904 ;
  assign n6940 = ~n6938 & ~n6939 ;
  assign n6941 = \u4_mem_reg[2][20]/NET0131  & ~n6904 ;
  assign n6942 = \u12_dout_reg[20]/P0001  & n6904 ;
  assign n6943 = ~n6941 & ~n6942 ;
  assign n6944 = \u4_mem_reg[2][21]/NET0131  & ~n6904 ;
  assign n6945 = \u12_dout_reg[21]/P0001  & n6904 ;
  assign n6946 = ~n6944 & ~n6945 ;
  assign n6947 = \u4_mem_reg[2][22]/NET0131  & ~n6904 ;
  assign n6948 = \u12_dout_reg[22]/P0001  & n6904 ;
  assign n6949 = ~n6947 & ~n6948 ;
  assign n6950 = \u4_mem_reg[2][23]/NET0131  & ~n6904 ;
  assign n6951 = \u12_dout_reg[23]/P0001  & n6904 ;
  assign n6952 = ~n6950 & ~n6951 ;
  assign n6953 = \u4_mem_reg[2][24]/NET0131  & ~n6904 ;
  assign n6954 = \u12_dout_reg[24]/P0001  & n6904 ;
  assign n6955 = ~n6953 & ~n6954 ;
  assign n6956 = \u4_mem_reg[2][25]/NET0131  & ~n6904 ;
  assign n6957 = \u12_dout_reg[25]/P0001  & n6904 ;
  assign n6958 = ~n6956 & ~n6957 ;
  assign n6959 = \u4_mem_reg[2][26]/NET0131  & ~n6904 ;
  assign n6960 = \u12_dout_reg[26]/P0001  & n6904 ;
  assign n6961 = ~n6959 & ~n6960 ;
  assign n6962 = \u4_mem_reg[2][27]/NET0131  & ~n6904 ;
  assign n6963 = \u12_dout_reg[27]/P0001  & n6904 ;
  assign n6964 = ~n6962 & ~n6963 ;
  assign n6965 = \u4_mem_reg[2][28]/NET0131  & ~n6904 ;
  assign n6966 = \u12_dout_reg[28]/P0001  & n6904 ;
  assign n6967 = ~n6965 & ~n6966 ;
  assign n6968 = \u4_mem_reg[2][29]/NET0131  & ~n6904 ;
  assign n6969 = \u12_dout_reg[29]/P0001  & n6904 ;
  assign n6970 = ~n6968 & ~n6969 ;
  assign n6971 = \u4_mem_reg[2][2]/NET0131  & ~n6904 ;
  assign n6972 = \u12_dout_reg[2]/P0001  & n6904 ;
  assign n6973 = ~n6971 & ~n6972 ;
  assign n6974 = \u4_mem_reg[2][30]/NET0131  & ~n6904 ;
  assign n6975 = \u12_dout_reg[30]/P0001  & n6904 ;
  assign n6976 = ~n6974 & ~n6975 ;
  assign n6977 = \u4_mem_reg[2][31]/NET0131  & ~n6904 ;
  assign n6978 = \u12_dout_reg[31]/P0001  & n6904 ;
  assign n6979 = ~n6977 & ~n6978 ;
  assign n6980 = \u4_mem_reg[2][3]/NET0131  & ~n6904 ;
  assign n6981 = \u12_dout_reg[3]/P0001  & n6904 ;
  assign n6982 = ~n6980 & ~n6981 ;
  assign n6983 = \u4_mem_reg[2][4]/NET0131  & ~n6904 ;
  assign n6984 = \u12_dout_reg[4]/P0001  & n6904 ;
  assign n6985 = ~n6983 & ~n6984 ;
  assign n6986 = \u4_mem_reg[2][5]/NET0131  & ~n6904 ;
  assign n6987 = \u12_dout_reg[5]/P0001  & n6904 ;
  assign n6988 = ~n6986 & ~n6987 ;
  assign n6989 = \u4_mem_reg[2][6]/NET0131  & ~n6904 ;
  assign n6990 = \u12_dout_reg[6]/P0001  & n6904 ;
  assign n6991 = ~n6989 & ~n6990 ;
  assign n6992 = \u4_mem_reg[2][7]/NET0131  & ~n6904 ;
  assign n6993 = \u12_dout_reg[7]/P0001  & n6904 ;
  assign n6994 = ~n6992 & ~n6993 ;
  assign n6995 = \u4_mem_reg[2][8]/NET0131  & ~n6904 ;
  assign n6996 = \u12_dout_reg[8]/P0001  & n6904 ;
  assign n6997 = ~n6995 & ~n6996 ;
  assign n6998 = \u4_mem_reg[2][9]/NET0131  & ~n6904 ;
  assign n6999 = \u12_dout_reg[9]/P0001  & n6904 ;
  assign n7000 = ~n6998 & ~n6999 ;
  assign n7001 = \u4_mem_reg[3][0]/NET0131  & ~n6307 ;
  assign n7002 = \u12_dout_reg[0]/P0001  & n6307 ;
  assign n7003 = ~n7001 & ~n7002 ;
  assign n7004 = \u4_mem_reg[3][10]/NET0131  & ~n6307 ;
  assign n7005 = \u12_dout_reg[10]/P0001  & n6307 ;
  assign n7006 = ~n7004 & ~n7005 ;
  assign n7007 = \u4_mem_reg[3][11]/NET0131  & ~n6307 ;
  assign n7008 = \u12_dout_reg[11]/P0001  & n6307 ;
  assign n7009 = ~n7007 & ~n7008 ;
  assign n7010 = \u4_mem_reg[3][12]/NET0131  & ~n6307 ;
  assign n7011 = \u12_dout_reg[12]/P0001  & n6307 ;
  assign n7012 = ~n7010 & ~n7011 ;
  assign n7013 = \u4_mem_reg[3][13]/NET0131  & ~n6307 ;
  assign n7014 = \u12_dout_reg[13]/P0001  & n6307 ;
  assign n7015 = ~n7013 & ~n7014 ;
  assign n7016 = \u4_mem_reg[3][14]/NET0131  & ~n6307 ;
  assign n7017 = \u12_dout_reg[14]/P0001  & n6307 ;
  assign n7018 = ~n7016 & ~n7017 ;
  assign n7019 = \u4_mem_reg[3][15]/NET0131  & ~n6307 ;
  assign n7020 = \u12_dout_reg[15]/P0001  & n6307 ;
  assign n7021 = ~n7019 & ~n7020 ;
  assign n7022 = \u4_mem_reg[3][16]/NET0131  & ~n6307 ;
  assign n7023 = \u12_dout_reg[16]/P0001  & n6307 ;
  assign n7024 = ~n7022 & ~n7023 ;
  assign n7025 = \u4_mem_reg[3][17]/NET0131  & ~n6307 ;
  assign n7026 = \u12_dout_reg[17]/P0001  & n6307 ;
  assign n7027 = ~n7025 & ~n7026 ;
  assign n7028 = \u4_mem_reg[3][18]/NET0131  & ~n6307 ;
  assign n7029 = \u12_dout_reg[18]/P0001  & n6307 ;
  assign n7030 = ~n7028 & ~n7029 ;
  assign n7031 = \u4_mem_reg[3][19]/NET0131  & ~n6307 ;
  assign n7032 = \u12_dout_reg[19]/P0001  & n6307 ;
  assign n7033 = ~n7031 & ~n7032 ;
  assign n7034 = \u4_mem_reg[3][1]/NET0131  & ~n6307 ;
  assign n7035 = \u12_dout_reg[1]/P0001  & n6307 ;
  assign n7036 = ~n7034 & ~n7035 ;
  assign n7037 = \u4_mem_reg[3][20]/NET0131  & ~n6307 ;
  assign n7038 = \u12_dout_reg[20]/P0001  & n6307 ;
  assign n7039 = ~n7037 & ~n7038 ;
  assign n7040 = \u4_mem_reg[3][21]/NET0131  & ~n6307 ;
  assign n7041 = \u12_dout_reg[21]/P0001  & n6307 ;
  assign n7042 = ~n7040 & ~n7041 ;
  assign n7043 = \u4_mem_reg[3][22]/NET0131  & ~n6307 ;
  assign n7044 = \u12_dout_reg[22]/P0001  & n6307 ;
  assign n7045 = ~n7043 & ~n7044 ;
  assign n7046 = \u4_mem_reg[3][23]/NET0131  & ~n6307 ;
  assign n7047 = \u12_dout_reg[23]/P0001  & n6307 ;
  assign n7048 = ~n7046 & ~n7047 ;
  assign n7049 = \u4_mem_reg[3][24]/NET0131  & ~n6307 ;
  assign n7050 = \u12_dout_reg[24]/P0001  & n6307 ;
  assign n7051 = ~n7049 & ~n7050 ;
  assign n7052 = \u4_mem_reg[3][25]/NET0131  & ~n6307 ;
  assign n7053 = \u12_dout_reg[25]/P0001  & n6307 ;
  assign n7054 = ~n7052 & ~n7053 ;
  assign n7055 = \u4_mem_reg[3][26]/NET0131  & ~n6307 ;
  assign n7056 = \u12_dout_reg[26]/P0001  & n6307 ;
  assign n7057 = ~n7055 & ~n7056 ;
  assign n7058 = \u4_mem_reg[3][27]/NET0131  & ~n6307 ;
  assign n7059 = \u12_dout_reg[27]/P0001  & n6307 ;
  assign n7060 = ~n7058 & ~n7059 ;
  assign n7061 = \u4_mem_reg[3][28]/NET0131  & ~n6307 ;
  assign n7062 = \u12_dout_reg[28]/P0001  & n6307 ;
  assign n7063 = ~n7061 & ~n7062 ;
  assign n7064 = \u4_mem_reg[3][29]/NET0131  & ~n6307 ;
  assign n7065 = \u12_dout_reg[29]/P0001  & n6307 ;
  assign n7066 = ~n7064 & ~n7065 ;
  assign n7067 = \u4_mem_reg[3][2]/NET0131  & ~n6307 ;
  assign n7068 = \u12_dout_reg[2]/P0001  & n6307 ;
  assign n7069 = ~n7067 & ~n7068 ;
  assign n7070 = \u4_mem_reg[3][30]/NET0131  & ~n6307 ;
  assign n7071 = \u12_dout_reg[30]/P0001  & n6307 ;
  assign n7072 = ~n7070 & ~n7071 ;
  assign n7073 = \u4_mem_reg[3][31]/NET0131  & ~n6307 ;
  assign n7074 = \u12_dout_reg[31]/P0001  & n6307 ;
  assign n7075 = ~n7073 & ~n7074 ;
  assign n7076 = \u4_mem_reg[3][3]/NET0131  & ~n6307 ;
  assign n7077 = \u12_dout_reg[3]/P0001  & n6307 ;
  assign n7078 = ~n7076 & ~n7077 ;
  assign n7079 = \u4_mem_reg[3][4]/NET0131  & ~n6307 ;
  assign n7080 = \u12_dout_reg[4]/P0001  & n6307 ;
  assign n7081 = ~n7079 & ~n7080 ;
  assign n7082 = \u4_mem_reg[3][5]/NET0131  & ~n6307 ;
  assign n7083 = \u12_dout_reg[5]/P0001  & n6307 ;
  assign n7084 = ~n7082 & ~n7083 ;
  assign n7085 = \u4_mem_reg[3][6]/NET0131  & ~n6307 ;
  assign n7086 = \u12_dout_reg[6]/P0001  & n6307 ;
  assign n7087 = ~n7085 & ~n7086 ;
  assign n7088 = \u4_mem_reg[3][7]/NET0131  & ~n6307 ;
  assign n7089 = \u12_dout_reg[7]/P0001  & n6307 ;
  assign n7090 = ~n7088 & ~n7089 ;
  assign n7091 = \u4_mem_reg[3][8]/NET0131  & ~n6307 ;
  assign n7092 = \u12_dout_reg[8]/P0001  & n6307 ;
  assign n7093 = ~n7091 & ~n7092 ;
  assign n7094 = \u4_mem_reg[3][9]/NET0131  & ~n6307 ;
  assign n7095 = \u12_dout_reg[9]/P0001  & n6307 ;
  assign n7096 = ~n7094 & ~n7095 ;
  assign n7097 = \u3_mem_reg[2][14]/NET0131  & ~n6583 ;
  assign n7098 = \u12_dout_reg[14]/P0001  & n6583 ;
  assign n7099 = ~n7097 & ~n7098 ;
  assign n7100 = ~\u5_wp_reg[1]/NET0131  & n6312 ;
  assign n7101 = \u5_mem_reg[1][0]/NET0131  & ~n7100 ;
  assign n7102 = \u12_dout_reg[0]/P0001  & n7100 ;
  assign n7103 = ~n7101 & ~n7102 ;
  assign n7104 = \u5_mem_reg[1][10]/NET0131  & ~n7100 ;
  assign n7105 = \u12_dout_reg[10]/P0001  & n7100 ;
  assign n7106 = ~n7104 & ~n7105 ;
  assign n7107 = \u5_mem_reg[1][11]/NET0131  & ~n7100 ;
  assign n7108 = \u12_dout_reg[11]/P0001  & n7100 ;
  assign n7109 = ~n7107 & ~n7108 ;
  assign n7110 = \u5_mem_reg[1][12]/NET0131  & ~n7100 ;
  assign n7111 = \u12_dout_reg[12]/P0001  & n7100 ;
  assign n7112 = ~n7110 & ~n7111 ;
  assign n7113 = \u5_mem_reg[1][13]/NET0131  & ~n7100 ;
  assign n7114 = \u12_dout_reg[13]/P0001  & n7100 ;
  assign n7115 = ~n7113 & ~n7114 ;
  assign n7116 = \u5_mem_reg[1][14]/NET0131  & ~n7100 ;
  assign n7117 = \u12_dout_reg[14]/P0001  & n7100 ;
  assign n7118 = ~n7116 & ~n7117 ;
  assign n7119 = \u5_mem_reg[1][15]/NET0131  & ~n7100 ;
  assign n7120 = \u12_dout_reg[15]/P0001  & n7100 ;
  assign n7121 = ~n7119 & ~n7120 ;
  assign n7122 = \u5_mem_reg[1][16]/NET0131  & ~n7100 ;
  assign n7123 = \u12_dout_reg[16]/P0001  & n7100 ;
  assign n7124 = ~n7122 & ~n7123 ;
  assign n7125 = \u5_mem_reg[1][17]/NET0131  & ~n7100 ;
  assign n7126 = \u12_dout_reg[17]/P0001  & n7100 ;
  assign n7127 = ~n7125 & ~n7126 ;
  assign n7128 = \u5_mem_reg[1][18]/NET0131  & ~n7100 ;
  assign n7129 = \u12_dout_reg[18]/P0001  & n7100 ;
  assign n7130 = ~n7128 & ~n7129 ;
  assign n7131 = \u5_mem_reg[1][19]/NET0131  & ~n7100 ;
  assign n7132 = \u12_dout_reg[19]/P0001  & n7100 ;
  assign n7133 = ~n7131 & ~n7132 ;
  assign n7134 = \u5_mem_reg[1][1]/NET0131  & ~n7100 ;
  assign n7135 = \u12_dout_reg[1]/P0001  & n7100 ;
  assign n7136 = ~n7134 & ~n7135 ;
  assign n7137 = \u5_mem_reg[1][20]/NET0131  & ~n7100 ;
  assign n7138 = \u12_dout_reg[20]/P0001  & n7100 ;
  assign n7139 = ~n7137 & ~n7138 ;
  assign n7140 = \u5_mem_reg[1][21]/NET0131  & ~n7100 ;
  assign n7141 = \u12_dout_reg[21]/P0001  & n7100 ;
  assign n7142 = ~n7140 & ~n7141 ;
  assign n7143 = \u5_mem_reg[1][22]/NET0131  & ~n7100 ;
  assign n7144 = \u12_dout_reg[22]/P0001  & n7100 ;
  assign n7145 = ~n7143 & ~n7144 ;
  assign n7146 = \u5_mem_reg[1][23]/NET0131  & ~n7100 ;
  assign n7147 = \u12_dout_reg[23]/P0001  & n7100 ;
  assign n7148 = ~n7146 & ~n7147 ;
  assign n7149 = \u5_mem_reg[1][24]/NET0131  & ~n7100 ;
  assign n7150 = \u12_dout_reg[24]/P0001  & n7100 ;
  assign n7151 = ~n7149 & ~n7150 ;
  assign n7152 = \u5_mem_reg[1][25]/NET0131  & ~n7100 ;
  assign n7153 = \u12_dout_reg[25]/P0001  & n7100 ;
  assign n7154 = ~n7152 & ~n7153 ;
  assign n7155 = \u5_mem_reg[1][26]/NET0131  & ~n7100 ;
  assign n7156 = \u12_dout_reg[26]/P0001  & n7100 ;
  assign n7157 = ~n7155 & ~n7156 ;
  assign n7158 = \u5_mem_reg[1][27]/NET0131  & ~n7100 ;
  assign n7159 = \u12_dout_reg[27]/P0001  & n7100 ;
  assign n7160 = ~n7158 & ~n7159 ;
  assign n7161 = \u5_mem_reg[1][28]/NET0131  & ~n7100 ;
  assign n7162 = \u12_dout_reg[28]/P0001  & n7100 ;
  assign n7163 = ~n7161 & ~n7162 ;
  assign n7164 = \u5_mem_reg[1][29]/NET0131  & ~n7100 ;
  assign n7165 = \u12_dout_reg[29]/P0001  & n7100 ;
  assign n7166 = ~n7164 & ~n7165 ;
  assign n7167 = \u5_mem_reg[1][2]/NET0131  & ~n7100 ;
  assign n7168 = \u12_dout_reg[2]/P0001  & n7100 ;
  assign n7169 = ~n7167 & ~n7168 ;
  assign n7170 = \u5_mem_reg[1][30]/NET0131  & ~n7100 ;
  assign n7171 = \u12_dout_reg[30]/P0001  & n7100 ;
  assign n7172 = ~n7170 & ~n7171 ;
  assign n7173 = \u5_mem_reg[1][31]/NET0131  & ~n7100 ;
  assign n7174 = \u12_dout_reg[31]/P0001  & n7100 ;
  assign n7175 = ~n7173 & ~n7174 ;
  assign n7176 = \u5_mem_reg[1][3]/NET0131  & ~n7100 ;
  assign n7177 = \u12_dout_reg[3]/P0001  & n7100 ;
  assign n7178 = ~n7176 & ~n7177 ;
  assign n7179 = \u5_mem_reg[1][4]/NET0131  & ~n7100 ;
  assign n7180 = \u12_dout_reg[4]/P0001  & n7100 ;
  assign n7181 = ~n7179 & ~n7180 ;
  assign n7182 = \u5_mem_reg[1][5]/NET0131  & ~n7100 ;
  assign n7183 = \u12_dout_reg[5]/P0001  & n7100 ;
  assign n7184 = ~n7182 & ~n7183 ;
  assign n7185 = \u5_mem_reg[1][6]/NET0131  & ~n7100 ;
  assign n7186 = \u12_dout_reg[6]/P0001  & n7100 ;
  assign n7187 = ~n7185 & ~n7186 ;
  assign n7188 = \u5_mem_reg[1][7]/NET0131  & ~n7100 ;
  assign n7189 = \u12_dout_reg[7]/P0001  & n7100 ;
  assign n7190 = ~n7188 & ~n7189 ;
  assign n7191 = \u5_mem_reg[1][8]/NET0131  & ~n7100 ;
  assign n7192 = \u12_dout_reg[8]/P0001  & n7100 ;
  assign n7193 = ~n7191 & ~n7192 ;
  assign n7194 = \u5_mem_reg[1][9]/NET0131  & ~n7100 ;
  assign n7195 = \u12_dout_reg[9]/P0001  & n7100 ;
  assign n7196 = ~n7194 & ~n7195 ;
  assign n7197 = \u5_wp_reg[1]/NET0131  & n6415 ;
  assign n7198 = \u5_mem_reg[2][0]/NET0131  & ~n7197 ;
  assign n7199 = \u12_dout_reg[0]/P0001  & n7197 ;
  assign n7200 = ~n7198 & ~n7199 ;
  assign n7201 = \u5_mem_reg[2][10]/NET0131  & ~n7197 ;
  assign n7202 = \u12_dout_reg[10]/P0001  & n7197 ;
  assign n7203 = ~n7201 & ~n7202 ;
  assign n7204 = \u5_mem_reg[2][11]/NET0131  & ~n7197 ;
  assign n7205 = \u12_dout_reg[11]/P0001  & n7197 ;
  assign n7206 = ~n7204 & ~n7205 ;
  assign n7207 = \u5_mem_reg[2][12]/NET0131  & ~n7197 ;
  assign n7208 = \u12_dout_reg[12]/P0001  & n7197 ;
  assign n7209 = ~n7207 & ~n7208 ;
  assign n7210 = \u5_mem_reg[2][13]/NET0131  & ~n7197 ;
  assign n7211 = \u12_dout_reg[13]/P0001  & n7197 ;
  assign n7212 = ~n7210 & ~n7211 ;
  assign n7213 = \u5_mem_reg[2][14]/NET0131  & ~n7197 ;
  assign n7214 = \u12_dout_reg[14]/P0001  & n7197 ;
  assign n7215 = ~n7213 & ~n7214 ;
  assign n7216 = \u5_mem_reg[2][15]/NET0131  & ~n7197 ;
  assign n7217 = \u12_dout_reg[15]/P0001  & n7197 ;
  assign n7218 = ~n7216 & ~n7217 ;
  assign n7219 = \u5_mem_reg[2][16]/NET0131  & ~n7197 ;
  assign n7220 = \u12_dout_reg[16]/P0001  & n7197 ;
  assign n7221 = ~n7219 & ~n7220 ;
  assign n7222 = \u5_mem_reg[2][17]/NET0131  & ~n7197 ;
  assign n7223 = \u12_dout_reg[17]/P0001  & n7197 ;
  assign n7224 = ~n7222 & ~n7223 ;
  assign n7225 = \u5_mem_reg[2][18]/NET0131  & ~n7197 ;
  assign n7226 = \u12_dout_reg[18]/P0001  & n7197 ;
  assign n7227 = ~n7225 & ~n7226 ;
  assign n7228 = \u5_mem_reg[2][19]/NET0131  & ~n7197 ;
  assign n7229 = \u12_dout_reg[19]/P0001  & n7197 ;
  assign n7230 = ~n7228 & ~n7229 ;
  assign n7231 = \u5_mem_reg[2][1]/NET0131  & ~n7197 ;
  assign n7232 = \u12_dout_reg[1]/P0001  & n7197 ;
  assign n7233 = ~n7231 & ~n7232 ;
  assign n7234 = \u5_mem_reg[2][20]/NET0131  & ~n7197 ;
  assign n7235 = \u12_dout_reg[20]/P0001  & n7197 ;
  assign n7236 = ~n7234 & ~n7235 ;
  assign n7237 = \u5_mem_reg[2][21]/NET0131  & ~n7197 ;
  assign n7238 = \u12_dout_reg[21]/P0001  & n7197 ;
  assign n7239 = ~n7237 & ~n7238 ;
  assign n7240 = \u5_mem_reg[2][22]/NET0131  & ~n7197 ;
  assign n7241 = \u12_dout_reg[22]/P0001  & n7197 ;
  assign n7242 = ~n7240 & ~n7241 ;
  assign n7243 = \u5_mem_reg[2][23]/NET0131  & ~n7197 ;
  assign n7244 = \u12_dout_reg[23]/P0001  & n7197 ;
  assign n7245 = ~n7243 & ~n7244 ;
  assign n7246 = \u5_mem_reg[2][24]/NET0131  & ~n7197 ;
  assign n7247 = \u12_dout_reg[24]/P0001  & n7197 ;
  assign n7248 = ~n7246 & ~n7247 ;
  assign n7249 = \u5_mem_reg[2][25]/NET0131  & ~n7197 ;
  assign n7250 = \u12_dout_reg[25]/P0001  & n7197 ;
  assign n7251 = ~n7249 & ~n7250 ;
  assign n7252 = \u5_mem_reg[2][26]/NET0131  & ~n7197 ;
  assign n7253 = \u12_dout_reg[26]/P0001  & n7197 ;
  assign n7254 = ~n7252 & ~n7253 ;
  assign n7255 = \u5_mem_reg[2][27]/NET0131  & ~n7197 ;
  assign n7256 = \u12_dout_reg[27]/P0001  & n7197 ;
  assign n7257 = ~n7255 & ~n7256 ;
  assign n7258 = \u5_mem_reg[2][28]/NET0131  & ~n7197 ;
  assign n7259 = \u12_dout_reg[28]/P0001  & n7197 ;
  assign n7260 = ~n7258 & ~n7259 ;
  assign n7261 = \u5_mem_reg[2][29]/NET0131  & ~n7197 ;
  assign n7262 = \u12_dout_reg[29]/P0001  & n7197 ;
  assign n7263 = ~n7261 & ~n7262 ;
  assign n7264 = \u5_mem_reg[2][2]/NET0131  & ~n7197 ;
  assign n7265 = \u12_dout_reg[2]/P0001  & n7197 ;
  assign n7266 = ~n7264 & ~n7265 ;
  assign n7267 = \u5_mem_reg[2][30]/NET0131  & ~n7197 ;
  assign n7268 = \u12_dout_reg[30]/P0001  & n7197 ;
  assign n7269 = ~n7267 & ~n7268 ;
  assign n7270 = \u5_mem_reg[2][31]/NET0131  & ~n7197 ;
  assign n7271 = \u12_dout_reg[31]/P0001  & n7197 ;
  assign n7272 = ~n7270 & ~n7271 ;
  assign n7273 = \u5_mem_reg[2][3]/NET0131  & ~n7197 ;
  assign n7274 = \u12_dout_reg[3]/P0001  & n7197 ;
  assign n7275 = ~n7273 & ~n7274 ;
  assign n7276 = \u5_mem_reg[2][4]/NET0131  & ~n7197 ;
  assign n7277 = \u12_dout_reg[4]/P0001  & n7197 ;
  assign n7278 = ~n7276 & ~n7277 ;
  assign n7279 = \u5_mem_reg[2][5]/NET0131  & ~n7197 ;
  assign n7280 = \u12_dout_reg[5]/P0001  & n7197 ;
  assign n7281 = ~n7279 & ~n7280 ;
  assign n7282 = \u5_mem_reg[2][6]/NET0131  & ~n7197 ;
  assign n7283 = \u12_dout_reg[6]/P0001  & n7197 ;
  assign n7284 = ~n7282 & ~n7283 ;
  assign n7285 = \u5_mem_reg[2][7]/NET0131  & ~n7197 ;
  assign n7286 = \u12_dout_reg[7]/P0001  & n7197 ;
  assign n7287 = ~n7285 & ~n7286 ;
  assign n7288 = \u5_mem_reg[2][8]/NET0131  & ~n7197 ;
  assign n7289 = \u12_dout_reg[8]/P0001  & n7197 ;
  assign n7290 = ~n7288 & ~n7289 ;
  assign n7291 = \u5_mem_reg[2][9]/NET0131  & ~n7197 ;
  assign n7292 = \u12_dout_reg[9]/P0001  & n7197 ;
  assign n7293 = ~n7291 & ~n7292 ;
  assign n7294 = \u5_mem_reg[3][0]/NET0131  & ~n6313 ;
  assign n7295 = \u12_dout_reg[0]/P0001  & n6313 ;
  assign n7296 = ~n7294 & ~n7295 ;
  assign n7297 = \u5_mem_reg[3][10]/NET0131  & ~n6313 ;
  assign n7298 = \u12_dout_reg[10]/P0001  & n6313 ;
  assign n7299 = ~n7297 & ~n7298 ;
  assign n7300 = \u5_mem_reg[3][11]/NET0131  & ~n6313 ;
  assign n7301 = \u12_dout_reg[11]/P0001  & n6313 ;
  assign n7302 = ~n7300 & ~n7301 ;
  assign n7303 = \u5_mem_reg[3][12]/NET0131  & ~n6313 ;
  assign n7304 = \u12_dout_reg[12]/P0001  & n6313 ;
  assign n7305 = ~n7303 & ~n7304 ;
  assign n7306 = \u5_mem_reg[3][13]/NET0131  & ~n6313 ;
  assign n7307 = \u12_dout_reg[13]/P0001  & n6313 ;
  assign n7308 = ~n7306 & ~n7307 ;
  assign n7309 = \u5_mem_reg[3][14]/NET0131  & ~n6313 ;
  assign n7310 = \u12_dout_reg[14]/P0001  & n6313 ;
  assign n7311 = ~n7309 & ~n7310 ;
  assign n7312 = \u5_mem_reg[3][15]/NET0131  & ~n6313 ;
  assign n7313 = \u12_dout_reg[15]/P0001  & n6313 ;
  assign n7314 = ~n7312 & ~n7313 ;
  assign n7315 = \u5_mem_reg[3][16]/NET0131  & ~n6313 ;
  assign n7316 = \u12_dout_reg[16]/P0001  & n6313 ;
  assign n7317 = ~n7315 & ~n7316 ;
  assign n7318 = \u5_mem_reg[3][17]/NET0131  & ~n6313 ;
  assign n7319 = \u12_dout_reg[17]/P0001  & n6313 ;
  assign n7320 = ~n7318 & ~n7319 ;
  assign n7321 = \u5_mem_reg[3][18]/NET0131  & ~n6313 ;
  assign n7322 = \u12_dout_reg[18]/P0001  & n6313 ;
  assign n7323 = ~n7321 & ~n7322 ;
  assign n7324 = \u5_mem_reg[3][19]/NET0131  & ~n6313 ;
  assign n7325 = \u12_dout_reg[19]/P0001  & n6313 ;
  assign n7326 = ~n7324 & ~n7325 ;
  assign n7327 = \u5_mem_reg[3][1]/NET0131  & ~n6313 ;
  assign n7328 = \u12_dout_reg[1]/P0001  & n6313 ;
  assign n7329 = ~n7327 & ~n7328 ;
  assign n7330 = \u5_mem_reg[3][20]/NET0131  & ~n6313 ;
  assign n7331 = \u12_dout_reg[20]/P0001  & n6313 ;
  assign n7332 = ~n7330 & ~n7331 ;
  assign n7333 = \u5_mem_reg[3][21]/NET0131  & ~n6313 ;
  assign n7334 = \u12_dout_reg[21]/P0001  & n6313 ;
  assign n7335 = ~n7333 & ~n7334 ;
  assign n7336 = \u5_mem_reg[3][22]/NET0131  & ~n6313 ;
  assign n7337 = \u12_dout_reg[22]/P0001  & n6313 ;
  assign n7338 = ~n7336 & ~n7337 ;
  assign n7339 = \u5_mem_reg[3][23]/NET0131  & ~n6313 ;
  assign n7340 = \u12_dout_reg[23]/P0001  & n6313 ;
  assign n7341 = ~n7339 & ~n7340 ;
  assign n7342 = \u5_mem_reg[3][24]/NET0131  & ~n6313 ;
  assign n7343 = \u12_dout_reg[24]/P0001  & n6313 ;
  assign n7344 = ~n7342 & ~n7343 ;
  assign n7345 = \u5_mem_reg[3][25]/NET0131  & ~n6313 ;
  assign n7346 = \u12_dout_reg[25]/P0001  & n6313 ;
  assign n7347 = ~n7345 & ~n7346 ;
  assign n7348 = \u5_mem_reg[3][26]/NET0131  & ~n6313 ;
  assign n7349 = \u12_dout_reg[26]/P0001  & n6313 ;
  assign n7350 = ~n7348 & ~n7349 ;
  assign n7351 = \u5_mem_reg[3][27]/NET0131  & ~n6313 ;
  assign n7352 = \u12_dout_reg[27]/P0001  & n6313 ;
  assign n7353 = ~n7351 & ~n7352 ;
  assign n7354 = \u5_mem_reg[3][28]/NET0131  & ~n6313 ;
  assign n7355 = \u12_dout_reg[28]/P0001  & n6313 ;
  assign n7356 = ~n7354 & ~n7355 ;
  assign n7357 = \u5_mem_reg[3][29]/NET0131  & ~n6313 ;
  assign n7358 = \u12_dout_reg[29]/P0001  & n6313 ;
  assign n7359 = ~n7357 & ~n7358 ;
  assign n7360 = \u5_mem_reg[3][2]/NET0131  & ~n6313 ;
  assign n7361 = \u12_dout_reg[2]/P0001  & n6313 ;
  assign n7362 = ~n7360 & ~n7361 ;
  assign n7363 = \u5_mem_reg[3][30]/NET0131  & ~n6313 ;
  assign n7364 = \u12_dout_reg[30]/P0001  & n6313 ;
  assign n7365 = ~n7363 & ~n7364 ;
  assign n7366 = \u5_mem_reg[3][31]/NET0131  & ~n6313 ;
  assign n7367 = \u12_dout_reg[31]/P0001  & n6313 ;
  assign n7368 = ~n7366 & ~n7367 ;
  assign n7369 = \u5_mem_reg[3][3]/NET0131  & ~n6313 ;
  assign n7370 = \u12_dout_reg[3]/P0001  & n6313 ;
  assign n7371 = ~n7369 & ~n7370 ;
  assign n7372 = \u5_mem_reg[3][4]/NET0131  & ~n6313 ;
  assign n7373 = \u12_dout_reg[4]/P0001  & n6313 ;
  assign n7374 = ~n7372 & ~n7373 ;
  assign n7375 = \u5_mem_reg[3][5]/NET0131  & ~n6313 ;
  assign n7376 = \u12_dout_reg[5]/P0001  & n6313 ;
  assign n7377 = ~n7375 & ~n7376 ;
  assign n7378 = \u5_mem_reg[3][6]/NET0131  & ~n6313 ;
  assign n7379 = \u12_dout_reg[6]/P0001  & n6313 ;
  assign n7380 = ~n7378 & ~n7379 ;
  assign n7381 = \u5_mem_reg[3][7]/NET0131  & ~n6313 ;
  assign n7382 = \u12_dout_reg[7]/P0001  & n6313 ;
  assign n7383 = ~n7381 & ~n7382 ;
  assign n7384 = \u5_mem_reg[3][8]/NET0131  & ~n6313 ;
  assign n7385 = \u12_dout_reg[8]/P0001  & n6313 ;
  assign n7386 = ~n7384 & ~n7385 ;
  assign n7387 = \u5_mem_reg[3][9]/NET0131  & ~n6313 ;
  assign n7388 = \u12_dout_reg[9]/P0001  & n6313 ;
  assign n7389 = ~n7387 & ~n7388 ;
  assign n7390 = \u8_mem_reg[3][6]/NET0131  & ~n6301 ;
  assign n7391 = \u12_dout_reg[6]/P0001  & n6301 ;
  assign n7392 = ~n7390 & ~n7391 ;
  assign n7393 = \u8_mem_reg[1][28]/NET0131  & ~n6629 ;
  assign n7394 = \u12_dout_reg[28]/P0001  & n6629 ;
  assign n7395 = ~n7393 & ~n7394 ;
  assign n7396 = \u3_mem_reg[2][20]/NET0131  & ~n6583 ;
  assign n7397 = \u12_dout_reg[20]/P0001  & n6583 ;
  assign n7398 = ~n7396 & ~n7397 ;
  assign n7399 = \u8_mem_reg[3][31]/NET0131  & ~n6301 ;
  assign n7400 = \u12_dout_reg[31]/P0001  & n6301 ;
  assign n7401 = ~n7399 & ~n7400 ;
  assign n7402 = ~\u6_wp_reg[1]/NET0131  & n6324 ;
  assign n7403 = \u6_mem_reg[1][0]/NET0131  & ~n7402 ;
  assign n7404 = \u12_dout_reg[0]/P0001  & n7402 ;
  assign n7405 = ~n7403 & ~n7404 ;
  assign n7406 = \u6_mem_reg[1][10]/NET0131  & ~n7402 ;
  assign n7407 = \u12_dout_reg[10]/P0001  & n7402 ;
  assign n7408 = ~n7406 & ~n7407 ;
  assign n7409 = \u6_mem_reg[1][11]/NET0131  & ~n7402 ;
  assign n7410 = \u12_dout_reg[11]/P0001  & n7402 ;
  assign n7411 = ~n7409 & ~n7410 ;
  assign n7412 = \u6_mem_reg[1][12]/NET0131  & ~n7402 ;
  assign n7413 = \u12_dout_reg[12]/P0001  & n7402 ;
  assign n7414 = ~n7412 & ~n7413 ;
  assign n7415 = \u6_mem_reg[1][13]/NET0131  & ~n7402 ;
  assign n7416 = \u12_dout_reg[13]/P0001  & n7402 ;
  assign n7417 = ~n7415 & ~n7416 ;
  assign n7418 = \u6_mem_reg[1][14]/NET0131  & ~n7402 ;
  assign n7419 = \u12_dout_reg[14]/P0001  & n7402 ;
  assign n7420 = ~n7418 & ~n7419 ;
  assign n7421 = \u6_mem_reg[1][15]/NET0131  & ~n7402 ;
  assign n7422 = \u12_dout_reg[15]/P0001  & n7402 ;
  assign n7423 = ~n7421 & ~n7422 ;
  assign n7424 = \u6_mem_reg[1][16]/NET0131  & ~n7402 ;
  assign n7425 = \u12_dout_reg[16]/P0001  & n7402 ;
  assign n7426 = ~n7424 & ~n7425 ;
  assign n7427 = \u6_mem_reg[1][17]/NET0131  & ~n7402 ;
  assign n7428 = \u12_dout_reg[17]/P0001  & n7402 ;
  assign n7429 = ~n7427 & ~n7428 ;
  assign n7430 = \u6_mem_reg[1][18]/NET0131  & ~n7402 ;
  assign n7431 = \u12_dout_reg[18]/P0001  & n7402 ;
  assign n7432 = ~n7430 & ~n7431 ;
  assign n7433 = \u6_mem_reg[1][19]/NET0131  & ~n7402 ;
  assign n7434 = \u12_dout_reg[19]/P0001  & n7402 ;
  assign n7435 = ~n7433 & ~n7434 ;
  assign n7436 = \u6_mem_reg[1][1]/NET0131  & ~n7402 ;
  assign n7437 = \u12_dout_reg[1]/P0001  & n7402 ;
  assign n7438 = ~n7436 & ~n7437 ;
  assign n7439 = \u6_mem_reg[1][20]/NET0131  & ~n7402 ;
  assign n7440 = \u12_dout_reg[20]/P0001  & n7402 ;
  assign n7441 = ~n7439 & ~n7440 ;
  assign n7442 = \u6_mem_reg[1][21]/NET0131  & ~n7402 ;
  assign n7443 = \u12_dout_reg[21]/P0001  & n7402 ;
  assign n7444 = ~n7442 & ~n7443 ;
  assign n7445 = \u6_mem_reg[1][22]/NET0131  & ~n7402 ;
  assign n7446 = \u12_dout_reg[22]/P0001  & n7402 ;
  assign n7447 = ~n7445 & ~n7446 ;
  assign n7448 = \u6_mem_reg[1][23]/NET0131  & ~n7402 ;
  assign n7449 = \u12_dout_reg[23]/P0001  & n7402 ;
  assign n7450 = ~n7448 & ~n7449 ;
  assign n7451 = \u6_mem_reg[1][24]/NET0131  & ~n7402 ;
  assign n7452 = \u12_dout_reg[24]/P0001  & n7402 ;
  assign n7453 = ~n7451 & ~n7452 ;
  assign n7454 = \u6_mem_reg[1][25]/NET0131  & ~n7402 ;
  assign n7455 = \u12_dout_reg[25]/P0001  & n7402 ;
  assign n7456 = ~n7454 & ~n7455 ;
  assign n7457 = \u6_mem_reg[1][26]/NET0131  & ~n7402 ;
  assign n7458 = \u12_dout_reg[26]/P0001  & n7402 ;
  assign n7459 = ~n7457 & ~n7458 ;
  assign n7460 = \u6_mem_reg[1][27]/NET0131  & ~n7402 ;
  assign n7461 = \u12_dout_reg[27]/P0001  & n7402 ;
  assign n7462 = ~n7460 & ~n7461 ;
  assign n7463 = \u6_mem_reg[1][28]/NET0131  & ~n7402 ;
  assign n7464 = \u12_dout_reg[28]/P0001  & n7402 ;
  assign n7465 = ~n7463 & ~n7464 ;
  assign n7466 = \u6_mem_reg[1][29]/NET0131  & ~n7402 ;
  assign n7467 = \u12_dout_reg[29]/P0001  & n7402 ;
  assign n7468 = ~n7466 & ~n7467 ;
  assign n7469 = \u6_mem_reg[1][2]/NET0131  & ~n7402 ;
  assign n7470 = \u12_dout_reg[2]/P0001  & n7402 ;
  assign n7471 = ~n7469 & ~n7470 ;
  assign n7472 = \u6_mem_reg[1][30]/NET0131  & ~n7402 ;
  assign n7473 = \u12_dout_reg[30]/P0001  & n7402 ;
  assign n7474 = ~n7472 & ~n7473 ;
  assign n7475 = \u6_mem_reg[1][31]/NET0131  & ~n7402 ;
  assign n7476 = \u12_dout_reg[31]/P0001  & n7402 ;
  assign n7477 = ~n7475 & ~n7476 ;
  assign n7478 = \u6_mem_reg[1][3]/NET0131  & ~n7402 ;
  assign n7479 = \u12_dout_reg[3]/P0001  & n7402 ;
  assign n7480 = ~n7478 & ~n7479 ;
  assign n7481 = \u6_mem_reg[1][4]/NET0131  & ~n7402 ;
  assign n7482 = \u12_dout_reg[4]/P0001  & n7402 ;
  assign n7483 = ~n7481 & ~n7482 ;
  assign n7484 = \u6_mem_reg[1][5]/NET0131  & ~n7402 ;
  assign n7485 = \u12_dout_reg[5]/P0001  & n7402 ;
  assign n7486 = ~n7484 & ~n7485 ;
  assign n7487 = \u6_mem_reg[1][6]/NET0131  & ~n7402 ;
  assign n7488 = \u12_dout_reg[6]/P0001  & n7402 ;
  assign n7489 = ~n7487 & ~n7488 ;
  assign n7490 = \u6_mem_reg[1][7]/NET0131  & ~n7402 ;
  assign n7491 = \u12_dout_reg[7]/P0001  & n7402 ;
  assign n7492 = ~n7490 & ~n7491 ;
  assign n7493 = \u6_mem_reg[1][8]/NET0131  & ~n7402 ;
  assign n7494 = \u12_dout_reg[8]/P0001  & n7402 ;
  assign n7495 = ~n7493 & ~n7494 ;
  assign n7496 = \u6_mem_reg[1][9]/NET0131  & ~n7402 ;
  assign n7497 = \u12_dout_reg[9]/P0001  & n7402 ;
  assign n7498 = ~n7496 & ~n7497 ;
  assign n7499 = \u6_wp_reg[1]/NET0131  & n6419 ;
  assign n7500 = \u6_mem_reg[2][0]/NET0131  & ~n7499 ;
  assign n7501 = \u12_dout_reg[0]/P0001  & n7499 ;
  assign n7502 = ~n7500 & ~n7501 ;
  assign n7503 = \u6_mem_reg[2][10]/NET0131  & ~n7499 ;
  assign n7504 = \u12_dout_reg[10]/P0001  & n7499 ;
  assign n7505 = ~n7503 & ~n7504 ;
  assign n7506 = \u6_mem_reg[2][11]/NET0131  & ~n7499 ;
  assign n7507 = \u12_dout_reg[11]/P0001  & n7499 ;
  assign n7508 = ~n7506 & ~n7507 ;
  assign n7509 = \u6_mem_reg[2][12]/NET0131  & ~n7499 ;
  assign n7510 = \u12_dout_reg[12]/P0001  & n7499 ;
  assign n7511 = ~n7509 & ~n7510 ;
  assign n7512 = \u6_mem_reg[2][13]/NET0131  & ~n7499 ;
  assign n7513 = \u12_dout_reg[13]/P0001  & n7499 ;
  assign n7514 = ~n7512 & ~n7513 ;
  assign n7515 = \u6_mem_reg[2][14]/NET0131  & ~n7499 ;
  assign n7516 = \u12_dout_reg[14]/P0001  & n7499 ;
  assign n7517 = ~n7515 & ~n7516 ;
  assign n7518 = \u6_mem_reg[2][15]/NET0131  & ~n7499 ;
  assign n7519 = \u12_dout_reg[15]/P0001  & n7499 ;
  assign n7520 = ~n7518 & ~n7519 ;
  assign n7521 = \u6_mem_reg[2][16]/NET0131  & ~n7499 ;
  assign n7522 = \u12_dout_reg[16]/P0001  & n7499 ;
  assign n7523 = ~n7521 & ~n7522 ;
  assign n7524 = \u6_mem_reg[2][17]/NET0131  & ~n7499 ;
  assign n7525 = \u12_dout_reg[17]/P0001  & n7499 ;
  assign n7526 = ~n7524 & ~n7525 ;
  assign n7527 = \u6_mem_reg[2][18]/NET0131  & ~n7499 ;
  assign n7528 = \u12_dout_reg[18]/P0001  & n7499 ;
  assign n7529 = ~n7527 & ~n7528 ;
  assign n7530 = \u6_mem_reg[2][19]/NET0131  & ~n7499 ;
  assign n7531 = \u12_dout_reg[19]/P0001  & n7499 ;
  assign n7532 = ~n7530 & ~n7531 ;
  assign n7533 = \u6_mem_reg[2][1]/NET0131  & ~n7499 ;
  assign n7534 = \u12_dout_reg[1]/P0001  & n7499 ;
  assign n7535 = ~n7533 & ~n7534 ;
  assign n7536 = \u6_mem_reg[2][20]/NET0131  & ~n7499 ;
  assign n7537 = \u12_dout_reg[20]/P0001  & n7499 ;
  assign n7538 = ~n7536 & ~n7537 ;
  assign n7539 = \u6_mem_reg[2][21]/NET0131  & ~n7499 ;
  assign n7540 = \u12_dout_reg[21]/P0001  & n7499 ;
  assign n7541 = ~n7539 & ~n7540 ;
  assign n7542 = \u6_mem_reg[2][22]/NET0131  & ~n7499 ;
  assign n7543 = \u12_dout_reg[22]/P0001  & n7499 ;
  assign n7544 = ~n7542 & ~n7543 ;
  assign n7545 = \u6_mem_reg[2][23]/NET0131  & ~n7499 ;
  assign n7546 = \u12_dout_reg[23]/P0001  & n7499 ;
  assign n7547 = ~n7545 & ~n7546 ;
  assign n7548 = \u6_mem_reg[2][24]/NET0131  & ~n7499 ;
  assign n7549 = \u12_dout_reg[24]/P0001  & n7499 ;
  assign n7550 = ~n7548 & ~n7549 ;
  assign n7551 = \u6_mem_reg[2][25]/NET0131  & ~n7499 ;
  assign n7552 = \u12_dout_reg[25]/P0001  & n7499 ;
  assign n7553 = ~n7551 & ~n7552 ;
  assign n7554 = \u6_mem_reg[2][26]/NET0131  & ~n7499 ;
  assign n7555 = \u12_dout_reg[26]/P0001  & n7499 ;
  assign n7556 = ~n7554 & ~n7555 ;
  assign n7557 = \u6_mem_reg[2][27]/NET0131  & ~n7499 ;
  assign n7558 = \u12_dout_reg[27]/P0001  & n7499 ;
  assign n7559 = ~n7557 & ~n7558 ;
  assign n7560 = \u6_mem_reg[2][28]/NET0131  & ~n7499 ;
  assign n7561 = \u12_dout_reg[28]/P0001  & n7499 ;
  assign n7562 = ~n7560 & ~n7561 ;
  assign n7563 = \u6_mem_reg[2][29]/NET0131  & ~n7499 ;
  assign n7564 = \u12_dout_reg[29]/P0001  & n7499 ;
  assign n7565 = ~n7563 & ~n7564 ;
  assign n7566 = \u6_mem_reg[2][2]/NET0131  & ~n7499 ;
  assign n7567 = \u12_dout_reg[2]/P0001  & n7499 ;
  assign n7568 = ~n7566 & ~n7567 ;
  assign n7569 = \u6_mem_reg[2][30]/NET0131  & ~n7499 ;
  assign n7570 = \u12_dout_reg[30]/P0001  & n7499 ;
  assign n7571 = ~n7569 & ~n7570 ;
  assign n7572 = \u6_mem_reg[2][31]/NET0131  & ~n7499 ;
  assign n7573 = \u12_dout_reg[31]/P0001  & n7499 ;
  assign n7574 = ~n7572 & ~n7573 ;
  assign n7575 = \u6_mem_reg[2][3]/NET0131  & ~n7499 ;
  assign n7576 = \u12_dout_reg[3]/P0001  & n7499 ;
  assign n7577 = ~n7575 & ~n7576 ;
  assign n7578 = \u6_mem_reg[2][4]/NET0131  & ~n7499 ;
  assign n7579 = \u12_dout_reg[4]/P0001  & n7499 ;
  assign n7580 = ~n7578 & ~n7579 ;
  assign n7581 = \u6_mem_reg[2][5]/NET0131  & ~n7499 ;
  assign n7582 = \u12_dout_reg[5]/P0001  & n7499 ;
  assign n7583 = ~n7581 & ~n7582 ;
  assign n7584 = \u6_mem_reg[2][6]/NET0131  & ~n7499 ;
  assign n7585 = \u12_dout_reg[6]/P0001  & n7499 ;
  assign n7586 = ~n7584 & ~n7585 ;
  assign n7587 = \u6_mem_reg[2][7]/NET0131  & ~n7499 ;
  assign n7588 = \u12_dout_reg[7]/P0001  & n7499 ;
  assign n7589 = ~n7587 & ~n7588 ;
  assign n7590 = \u6_mem_reg[2][8]/NET0131  & ~n7499 ;
  assign n7591 = \u12_dout_reg[8]/P0001  & n7499 ;
  assign n7592 = ~n7590 & ~n7591 ;
  assign n7593 = \u6_mem_reg[2][9]/NET0131  & ~n7499 ;
  assign n7594 = \u12_dout_reg[9]/P0001  & n7499 ;
  assign n7595 = ~n7593 & ~n7594 ;
  assign n7596 = \u6_mem_reg[3][0]/NET0131  & ~n6325 ;
  assign n7597 = \u12_dout_reg[0]/P0001  & n6325 ;
  assign n7598 = ~n7596 & ~n7597 ;
  assign n7599 = \u6_mem_reg[3][10]/NET0131  & ~n6325 ;
  assign n7600 = \u12_dout_reg[10]/P0001  & n6325 ;
  assign n7601 = ~n7599 & ~n7600 ;
  assign n7602 = \u6_mem_reg[3][11]/NET0131  & ~n6325 ;
  assign n7603 = \u12_dout_reg[11]/P0001  & n6325 ;
  assign n7604 = ~n7602 & ~n7603 ;
  assign n7605 = \u6_mem_reg[3][12]/NET0131  & ~n6325 ;
  assign n7606 = \u12_dout_reg[12]/P0001  & n6325 ;
  assign n7607 = ~n7605 & ~n7606 ;
  assign n7608 = \u6_mem_reg[3][13]/NET0131  & ~n6325 ;
  assign n7609 = \u12_dout_reg[13]/P0001  & n6325 ;
  assign n7610 = ~n7608 & ~n7609 ;
  assign n7611 = \u6_mem_reg[3][14]/NET0131  & ~n6325 ;
  assign n7612 = \u12_dout_reg[14]/P0001  & n6325 ;
  assign n7613 = ~n7611 & ~n7612 ;
  assign n7614 = \u6_mem_reg[3][15]/NET0131  & ~n6325 ;
  assign n7615 = \u12_dout_reg[15]/P0001  & n6325 ;
  assign n7616 = ~n7614 & ~n7615 ;
  assign n7617 = \u6_mem_reg[3][16]/NET0131  & ~n6325 ;
  assign n7618 = \u12_dout_reg[16]/P0001  & n6325 ;
  assign n7619 = ~n7617 & ~n7618 ;
  assign n7620 = \u6_mem_reg[3][17]/NET0131  & ~n6325 ;
  assign n7621 = \u12_dout_reg[17]/P0001  & n6325 ;
  assign n7622 = ~n7620 & ~n7621 ;
  assign n7623 = \u6_mem_reg[3][18]/NET0131  & ~n6325 ;
  assign n7624 = \u12_dout_reg[18]/P0001  & n6325 ;
  assign n7625 = ~n7623 & ~n7624 ;
  assign n7626 = \u6_mem_reg[3][19]/NET0131  & ~n6325 ;
  assign n7627 = \u12_dout_reg[19]/P0001  & n6325 ;
  assign n7628 = ~n7626 & ~n7627 ;
  assign n7629 = \u6_mem_reg[3][1]/NET0131  & ~n6325 ;
  assign n7630 = \u12_dout_reg[1]/P0001  & n6325 ;
  assign n7631 = ~n7629 & ~n7630 ;
  assign n7632 = \u6_mem_reg[3][20]/NET0131  & ~n6325 ;
  assign n7633 = \u12_dout_reg[20]/P0001  & n6325 ;
  assign n7634 = ~n7632 & ~n7633 ;
  assign n7635 = \u6_mem_reg[3][21]/NET0131  & ~n6325 ;
  assign n7636 = \u12_dout_reg[21]/P0001  & n6325 ;
  assign n7637 = ~n7635 & ~n7636 ;
  assign n7638 = \u6_mem_reg[3][22]/NET0131  & ~n6325 ;
  assign n7639 = \u12_dout_reg[22]/P0001  & n6325 ;
  assign n7640 = ~n7638 & ~n7639 ;
  assign n7641 = \u6_mem_reg[3][23]/NET0131  & ~n6325 ;
  assign n7642 = \u12_dout_reg[23]/P0001  & n6325 ;
  assign n7643 = ~n7641 & ~n7642 ;
  assign n7644 = \u6_mem_reg[3][24]/NET0131  & ~n6325 ;
  assign n7645 = \u12_dout_reg[24]/P0001  & n6325 ;
  assign n7646 = ~n7644 & ~n7645 ;
  assign n7647 = \u6_mem_reg[3][25]/NET0131  & ~n6325 ;
  assign n7648 = \u12_dout_reg[25]/P0001  & n6325 ;
  assign n7649 = ~n7647 & ~n7648 ;
  assign n7650 = \u6_mem_reg[3][26]/NET0131  & ~n6325 ;
  assign n7651 = \u12_dout_reg[26]/P0001  & n6325 ;
  assign n7652 = ~n7650 & ~n7651 ;
  assign n7653 = \u6_mem_reg[3][27]/NET0131  & ~n6325 ;
  assign n7654 = \u12_dout_reg[27]/P0001  & n6325 ;
  assign n7655 = ~n7653 & ~n7654 ;
  assign n7656 = \u6_mem_reg[3][28]/NET0131  & ~n6325 ;
  assign n7657 = \u12_dout_reg[28]/P0001  & n6325 ;
  assign n7658 = ~n7656 & ~n7657 ;
  assign n7659 = \u6_mem_reg[3][29]/NET0131  & ~n6325 ;
  assign n7660 = \u12_dout_reg[29]/P0001  & n6325 ;
  assign n7661 = ~n7659 & ~n7660 ;
  assign n7662 = \u6_mem_reg[3][2]/NET0131  & ~n6325 ;
  assign n7663 = \u12_dout_reg[2]/P0001  & n6325 ;
  assign n7664 = ~n7662 & ~n7663 ;
  assign n7665 = \u6_mem_reg[3][30]/NET0131  & ~n6325 ;
  assign n7666 = \u12_dout_reg[30]/P0001  & n6325 ;
  assign n7667 = ~n7665 & ~n7666 ;
  assign n7668 = \u6_mem_reg[3][31]/NET0131  & ~n6325 ;
  assign n7669 = \u12_dout_reg[31]/P0001  & n6325 ;
  assign n7670 = ~n7668 & ~n7669 ;
  assign n7671 = \u6_mem_reg[3][3]/NET0131  & ~n6325 ;
  assign n7672 = \u12_dout_reg[3]/P0001  & n6325 ;
  assign n7673 = ~n7671 & ~n7672 ;
  assign n7674 = \u6_mem_reg[3][4]/NET0131  & ~n6325 ;
  assign n7675 = \u12_dout_reg[4]/P0001  & n6325 ;
  assign n7676 = ~n7674 & ~n7675 ;
  assign n7677 = \u6_mem_reg[3][5]/NET0131  & ~n6325 ;
  assign n7678 = \u12_dout_reg[5]/P0001  & n6325 ;
  assign n7679 = ~n7677 & ~n7678 ;
  assign n7680 = \u6_mem_reg[3][6]/NET0131  & ~n6325 ;
  assign n7681 = \u12_dout_reg[6]/P0001  & n6325 ;
  assign n7682 = ~n7680 & ~n7681 ;
  assign n7683 = \u6_mem_reg[3][7]/NET0131  & ~n6325 ;
  assign n7684 = \u12_dout_reg[7]/P0001  & n6325 ;
  assign n7685 = ~n7683 & ~n7684 ;
  assign n7686 = \u6_mem_reg[3][8]/NET0131  & ~n6325 ;
  assign n7687 = \u12_dout_reg[8]/P0001  & n6325 ;
  assign n7688 = ~n7686 & ~n7687 ;
  assign n7689 = \u6_mem_reg[3][9]/NET0131  & ~n6325 ;
  assign n7690 = \u12_dout_reg[9]/P0001  & n6325 ;
  assign n7691 = ~n7689 & ~n7690 ;
  assign n7692 = \u8_mem_reg[1][6]/NET0131  & ~n6629 ;
  assign n7693 = \u12_dout_reg[6]/P0001  & n6629 ;
  assign n7694 = ~n7692 & ~n7693 ;
  assign n7695 = \u3_mem_reg[2][25]/NET0131  & ~n6583 ;
  assign n7696 = \u12_dout_reg[25]/P0001  & n6583 ;
  assign n7697 = ~n7695 & ~n7696 ;
  assign n7698 = \u8_mem_reg[3][4]/NET0131  & ~n6301 ;
  assign n7699 = \u12_dout_reg[4]/P0001  & n6301 ;
  assign n7700 = ~n7698 & ~n7699 ;
  assign n7701 = \u3_mem_reg[3][3]/NET0131  & ~n6319 ;
  assign n7702 = \u12_dout_reg[3]/P0001  & n6319 ;
  assign n7703 = ~n7701 & ~n7702 ;
  assign n7704 = \u8_mem_reg[3][8]/NET0131  & ~n6301 ;
  assign n7705 = \u12_dout_reg[8]/P0001  & n6301 ;
  assign n7706 = ~n7704 & ~n7705 ;
  assign n7707 = \u3_mem_reg[1][14]/NET0131  & ~n6489 ;
  assign n7708 = \u12_dout_reg[14]/P0001  & n6489 ;
  assign n7709 = ~n7707 & ~n7708 ;
  assign n7710 = ~\u7_wp_reg[1]/NET0131  & n6330 ;
  assign n7711 = \u7_mem_reg[1][0]/NET0131  & ~n7710 ;
  assign n7712 = \u12_dout_reg[0]/P0001  & n7710 ;
  assign n7713 = ~n7711 & ~n7712 ;
  assign n7714 = \u7_mem_reg[1][10]/NET0131  & ~n7710 ;
  assign n7715 = \u12_dout_reg[10]/P0001  & n7710 ;
  assign n7716 = ~n7714 & ~n7715 ;
  assign n7717 = \u7_mem_reg[1][11]/NET0131  & ~n7710 ;
  assign n7718 = \u12_dout_reg[11]/P0001  & n7710 ;
  assign n7719 = ~n7717 & ~n7718 ;
  assign n7720 = \u3_mem_reg[1][23]/NET0131  & ~n6489 ;
  assign n7721 = \u12_dout_reg[23]/P0001  & n6489 ;
  assign n7722 = ~n7720 & ~n7721 ;
  assign n7723 = \u7_mem_reg[1][12]/NET0131  & ~n7710 ;
  assign n7724 = \u12_dout_reg[12]/P0001  & n7710 ;
  assign n7725 = ~n7723 & ~n7724 ;
  assign n7726 = \u7_mem_reg[1][13]/NET0131  & ~n7710 ;
  assign n7727 = \u12_dout_reg[13]/P0001  & n7710 ;
  assign n7728 = ~n7726 & ~n7727 ;
  assign n7729 = \u7_mem_reg[1][14]/NET0131  & ~n7710 ;
  assign n7730 = \u12_dout_reg[14]/P0001  & n7710 ;
  assign n7731 = ~n7729 & ~n7730 ;
  assign n7732 = \u7_mem_reg[1][15]/NET0131  & ~n7710 ;
  assign n7733 = \u12_dout_reg[15]/P0001  & n7710 ;
  assign n7734 = ~n7732 & ~n7733 ;
  assign n7735 = \u7_mem_reg[1][16]/NET0131  & ~n7710 ;
  assign n7736 = \u12_dout_reg[16]/P0001  & n7710 ;
  assign n7737 = ~n7735 & ~n7736 ;
  assign n7738 = \u7_mem_reg[1][17]/NET0131  & ~n7710 ;
  assign n7739 = \u12_dout_reg[17]/P0001  & n7710 ;
  assign n7740 = ~n7738 & ~n7739 ;
  assign n7741 = \u7_mem_reg[1][18]/NET0131  & ~n7710 ;
  assign n7742 = \u12_dout_reg[18]/P0001  & n7710 ;
  assign n7743 = ~n7741 & ~n7742 ;
  assign n7744 = \u7_mem_reg[1][19]/NET0131  & ~n7710 ;
  assign n7745 = \u12_dout_reg[19]/P0001  & n7710 ;
  assign n7746 = ~n7744 & ~n7745 ;
  assign n7747 = \u7_mem_reg[1][1]/NET0131  & ~n7710 ;
  assign n7748 = \u12_dout_reg[1]/P0001  & n7710 ;
  assign n7749 = ~n7747 & ~n7748 ;
  assign n7750 = \u7_mem_reg[1][20]/NET0131  & ~n7710 ;
  assign n7751 = \u12_dout_reg[20]/P0001  & n7710 ;
  assign n7752 = ~n7750 & ~n7751 ;
  assign n7753 = \u7_mem_reg[1][21]/NET0131  & ~n7710 ;
  assign n7754 = \u12_dout_reg[21]/P0001  & n7710 ;
  assign n7755 = ~n7753 & ~n7754 ;
  assign n7756 = \u7_mem_reg[1][22]/NET0131  & ~n7710 ;
  assign n7757 = \u12_dout_reg[22]/P0001  & n7710 ;
  assign n7758 = ~n7756 & ~n7757 ;
  assign n7759 = \u7_mem_reg[1][23]/NET0131  & ~n7710 ;
  assign n7760 = \u12_dout_reg[23]/P0001  & n7710 ;
  assign n7761 = ~n7759 & ~n7760 ;
  assign n7762 = \u7_mem_reg[1][24]/NET0131  & ~n7710 ;
  assign n7763 = \u12_dout_reg[24]/P0001  & n7710 ;
  assign n7764 = ~n7762 & ~n7763 ;
  assign n7765 = \u7_mem_reg[1][25]/NET0131  & ~n7710 ;
  assign n7766 = \u12_dout_reg[25]/P0001  & n7710 ;
  assign n7767 = ~n7765 & ~n7766 ;
  assign n7768 = \u7_mem_reg[1][26]/NET0131  & ~n7710 ;
  assign n7769 = \u12_dout_reg[26]/P0001  & n7710 ;
  assign n7770 = ~n7768 & ~n7769 ;
  assign n7771 = \u7_mem_reg[1][27]/NET0131  & ~n7710 ;
  assign n7772 = \u12_dout_reg[27]/P0001  & n7710 ;
  assign n7773 = ~n7771 & ~n7772 ;
  assign n7774 = \u7_mem_reg[1][28]/NET0131  & ~n7710 ;
  assign n7775 = \u12_dout_reg[28]/P0001  & n7710 ;
  assign n7776 = ~n7774 & ~n7775 ;
  assign n7777 = \u7_mem_reg[1][29]/NET0131  & ~n7710 ;
  assign n7778 = \u12_dout_reg[29]/P0001  & n7710 ;
  assign n7779 = ~n7777 & ~n7778 ;
  assign n7780 = \u7_mem_reg[1][2]/NET0131  & ~n7710 ;
  assign n7781 = \u12_dout_reg[2]/P0001  & n7710 ;
  assign n7782 = ~n7780 & ~n7781 ;
  assign n7783 = \u7_mem_reg[1][30]/NET0131  & ~n7710 ;
  assign n7784 = \u12_dout_reg[30]/P0001  & n7710 ;
  assign n7785 = ~n7783 & ~n7784 ;
  assign n7786 = \u7_mem_reg[1][31]/NET0131  & ~n7710 ;
  assign n7787 = \u12_dout_reg[31]/P0001  & n7710 ;
  assign n7788 = ~n7786 & ~n7787 ;
  assign n7789 = \u7_mem_reg[1][3]/NET0131  & ~n7710 ;
  assign n7790 = \u12_dout_reg[3]/P0001  & n7710 ;
  assign n7791 = ~n7789 & ~n7790 ;
  assign n7792 = \u7_mem_reg[1][4]/NET0131  & ~n7710 ;
  assign n7793 = \u12_dout_reg[4]/P0001  & n7710 ;
  assign n7794 = ~n7792 & ~n7793 ;
  assign n7795 = \u7_mem_reg[1][5]/NET0131  & ~n7710 ;
  assign n7796 = \u12_dout_reg[5]/P0001  & n7710 ;
  assign n7797 = ~n7795 & ~n7796 ;
  assign n7798 = \u7_mem_reg[1][6]/NET0131  & ~n7710 ;
  assign n7799 = \u12_dout_reg[6]/P0001  & n7710 ;
  assign n7800 = ~n7798 & ~n7799 ;
  assign n7801 = \u7_mem_reg[1][7]/NET0131  & ~n7710 ;
  assign n7802 = \u12_dout_reg[7]/P0001  & n7710 ;
  assign n7803 = ~n7801 & ~n7802 ;
  assign n7804 = \u7_mem_reg[1][8]/NET0131  & ~n7710 ;
  assign n7805 = \u12_dout_reg[8]/P0001  & n7710 ;
  assign n7806 = ~n7804 & ~n7805 ;
  assign n7807 = \u3_mem_reg[3][20]/NET0131  & ~n6319 ;
  assign n7808 = \u12_dout_reg[20]/P0001  & n6319 ;
  assign n7809 = ~n7807 & ~n7808 ;
  assign n7810 = \u7_mem_reg[1][9]/NET0131  & ~n7710 ;
  assign n7811 = \u12_dout_reg[9]/P0001  & n7710 ;
  assign n7812 = ~n7810 & ~n7811 ;
  assign n7813 = \u7_wp_reg[1]/NET0131  & n6423 ;
  assign n7814 = \u7_mem_reg[2][0]/NET0131  & ~n7813 ;
  assign n7815 = \u12_dout_reg[0]/P0001  & n7813 ;
  assign n7816 = ~n7814 & ~n7815 ;
  assign n7817 = \u7_mem_reg[2][10]/NET0131  & ~n7813 ;
  assign n7818 = \u12_dout_reg[10]/P0001  & n7813 ;
  assign n7819 = ~n7817 & ~n7818 ;
  assign n7820 = \u7_mem_reg[2][11]/NET0131  & ~n7813 ;
  assign n7821 = \u12_dout_reg[11]/P0001  & n7813 ;
  assign n7822 = ~n7820 & ~n7821 ;
  assign n7823 = \u7_mem_reg[2][12]/NET0131  & ~n7813 ;
  assign n7824 = \u12_dout_reg[12]/P0001  & n7813 ;
  assign n7825 = ~n7823 & ~n7824 ;
  assign n7826 = \u7_mem_reg[2][13]/NET0131  & ~n7813 ;
  assign n7827 = \u12_dout_reg[13]/P0001  & n7813 ;
  assign n7828 = ~n7826 & ~n7827 ;
  assign n7829 = \u7_mem_reg[2][14]/NET0131  & ~n7813 ;
  assign n7830 = \u12_dout_reg[14]/P0001  & n7813 ;
  assign n7831 = ~n7829 & ~n7830 ;
  assign n7832 = \u7_mem_reg[2][15]/NET0131  & ~n7813 ;
  assign n7833 = \u12_dout_reg[15]/P0001  & n7813 ;
  assign n7834 = ~n7832 & ~n7833 ;
  assign n7835 = \u7_mem_reg[2][16]/NET0131  & ~n7813 ;
  assign n7836 = \u12_dout_reg[16]/P0001  & n7813 ;
  assign n7837 = ~n7835 & ~n7836 ;
  assign n7838 = \u7_mem_reg[2][17]/NET0131  & ~n7813 ;
  assign n7839 = \u12_dout_reg[17]/P0001  & n7813 ;
  assign n7840 = ~n7838 & ~n7839 ;
  assign n7841 = \u7_mem_reg[2][18]/NET0131  & ~n7813 ;
  assign n7842 = \u12_dout_reg[18]/P0001  & n7813 ;
  assign n7843 = ~n7841 & ~n7842 ;
  assign n7844 = \u7_mem_reg[2][19]/NET0131  & ~n7813 ;
  assign n7845 = \u12_dout_reg[19]/P0001  & n7813 ;
  assign n7846 = ~n7844 & ~n7845 ;
  assign n7847 = \u7_mem_reg[2][1]/NET0131  & ~n7813 ;
  assign n7848 = \u12_dout_reg[1]/P0001  & n7813 ;
  assign n7849 = ~n7847 & ~n7848 ;
  assign n7850 = \u7_mem_reg[2][20]/NET0131  & ~n7813 ;
  assign n7851 = \u12_dout_reg[20]/P0001  & n7813 ;
  assign n7852 = ~n7850 & ~n7851 ;
  assign n7853 = \u7_mem_reg[2][21]/NET0131  & ~n7813 ;
  assign n7854 = \u12_dout_reg[21]/P0001  & n7813 ;
  assign n7855 = ~n7853 & ~n7854 ;
  assign n7856 = \u7_mem_reg[2][22]/NET0131  & ~n7813 ;
  assign n7857 = \u12_dout_reg[22]/P0001  & n7813 ;
  assign n7858 = ~n7856 & ~n7857 ;
  assign n7859 = \u7_mem_reg[2][23]/NET0131  & ~n7813 ;
  assign n7860 = \u12_dout_reg[23]/P0001  & n7813 ;
  assign n7861 = ~n7859 & ~n7860 ;
  assign n7862 = \u7_mem_reg[2][24]/NET0131  & ~n7813 ;
  assign n7863 = \u12_dout_reg[24]/P0001  & n7813 ;
  assign n7864 = ~n7862 & ~n7863 ;
  assign n7865 = \u7_mem_reg[2][25]/NET0131  & ~n7813 ;
  assign n7866 = \u12_dout_reg[25]/P0001  & n7813 ;
  assign n7867 = ~n7865 & ~n7866 ;
  assign n7868 = \u7_mem_reg[2][26]/NET0131  & ~n7813 ;
  assign n7869 = \u12_dout_reg[26]/P0001  & n7813 ;
  assign n7870 = ~n7868 & ~n7869 ;
  assign n7871 = \u7_mem_reg[2][27]/NET0131  & ~n7813 ;
  assign n7872 = \u12_dout_reg[27]/P0001  & n7813 ;
  assign n7873 = ~n7871 & ~n7872 ;
  assign n7874 = \u7_mem_reg[2][28]/NET0131  & ~n7813 ;
  assign n7875 = \u12_dout_reg[28]/P0001  & n7813 ;
  assign n7876 = ~n7874 & ~n7875 ;
  assign n7877 = \u7_mem_reg[2][29]/NET0131  & ~n7813 ;
  assign n7878 = \u12_dout_reg[29]/P0001  & n7813 ;
  assign n7879 = ~n7877 & ~n7878 ;
  assign n7880 = \u7_mem_reg[2][2]/NET0131  & ~n7813 ;
  assign n7881 = \u12_dout_reg[2]/P0001  & n7813 ;
  assign n7882 = ~n7880 & ~n7881 ;
  assign n7883 = \u7_mem_reg[2][30]/NET0131  & ~n7813 ;
  assign n7884 = \u12_dout_reg[30]/P0001  & n7813 ;
  assign n7885 = ~n7883 & ~n7884 ;
  assign n7886 = \u7_mem_reg[2][31]/NET0131  & ~n7813 ;
  assign n7887 = \u12_dout_reg[31]/P0001  & n7813 ;
  assign n7888 = ~n7886 & ~n7887 ;
  assign n7889 = \u7_mem_reg[2][3]/NET0131  & ~n7813 ;
  assign n7890 = \u12_dout_reg[3]/P0001  & n7813 ;
  assign n7891 = ~n7889 & ~n7890 ;
  assign n7892 = \u7_mem_reg[2][4]/NET0131  & ~n7813 ;
  assign n7893 = \u12_dout_reg[4]/P0001  & n7813 ;
  assign n7894 = ~n7892 & ~n7893 ;
  assign n7895 = \u7_mem_reg[2][5]/NET0131  & ~n7813 ;
  assign n7896 = \u12_dout_reg[5]/P0001  & n7813 ;
  assign n7897 = ~n7895 & ~n7896 ;
  assign n7898 = \u7_mem_reg[2][6]/NET0131  & ~n7813 ;
  assign n7899 = \u12_dout_reg[6]/P0001  & n7813 ;
  assign n7900 = ~n7898 & ~n7899 ;
  assign n7901 = \u7_mem_reg[2][7]/NET0131  & ~n7813 ;
  assign n7902 = \u12_dout_reg[7]/P0001  & n7813 ;
  assign n7903 = ~n7901 & ~n7902 ;
  assign n7904 = \u7_mem_reg[2][8]/NET0131  & ~n7813 ;
  assign n7905 = \u12_dout_reg[8]/P0001  & n7813 ;
  assign n7906 = ~n7904 & ~n7905 ;
  assign n7907 = \u7_mem_reg[2][9]/NET0131  & ~n7813 ;
  assign n7908 = \u12_dout_reg[9]/P0001  & n7813 ;
  assign n7909 = ~n7907 & ~n7908 ;
  assign n7910 = \u7_mem_reg[3][0]/NET0131  & ~n6331 ;
  assign n7911 = \u12_dout_reg[0]/P0001  & n6331 ;
  assign n7912 = ~n7910 & ~n7911 ;
  assign n7913 = \u7_mem_reg[3][10]/NET0131  & ~n6331 ;
  assign n7914 = \u12_dout_reg[10]/P0001  & n6331 ;
  assign n7915 = ~n7913 & ~n7914 ;
  assign n7916 = \u7_mem_reg[3][11]/NET0131  & ~n6331 ;
  assign n7917 = \u12_dout_reg[11]/P0001  & n6331 ;
  assign n7918 = ~n7916 & ~n7917 ;
  assign n7919 = \u7_mem_reg[3][12]/NET0131  & ~n6331 ;
  assign n7920 = \u12_dout_reg[12]/P0001  & n6331 ;
  assign n7921 = ~n7919 & ~n7920 ;
  assign n7922 = \u7_mem_reg[3][13]/NET0131  & ~n6331 ;
  assign n7923 = \u12_dout_reg[13]/P0001  & n6331 ;
  assign n7924 = ~n7922 & ~n7923 ;
  assign n7925 = \u7_mem_reg[3][14]/NET0131  & ~n6331 ;
  assign n7926 = \u12_dout_reg[14]/P0001  & n6331 ;
  assign n7927 = ~n7925 & ~n7926 ;
  assign n7928 = \u7_mem_reg[3][15]/NET0131  & ~n6331 ;
  assign n7929 = \u12_dout_reg[15]/P0001  & n6331 ;
  assign n7930 = ~n7928 & ~n7929 ;
  assign n7931 = \u7_mem_reg[3][16]/NET0131  & ~n6331 ;
  assign n7932 = \u12_dout_reg[16]/P0001  & n6331 ;
  assign n7933 = ~n7931 & ~n7932 ;
  assign n7934 = \u7_mem_reg[3][17]/NET0131  & ~n6331 ;
  assign n7935 = \u12_dout_reg[17]/P0001  & n6331 ;
  assign n7936 = ~n7934 & ~n7935 ;
  assign n7937 = \u7_mem_reg[3][18]/NET0131  & ~n6331 ;
  assign n7938 = \u12_dout_reg[18]/P0001  & n6331 ;
  assign n7939 = ~n7937 & ~n7938 ;
  assign n7940 = \u7_mem_reg[3][19]/NET0131  & ~n6331 ;
  assign n7941 = \u12_dout_reg[19]/P0001  & n6331 ;
  assign n7942 = ~n7940 & ~n7941 ;
  assign n7943 = \u7_mem_reg[3][1]/NET0131  & ~n6331 ;
  assign n7944 = \u12_dout_reg[1]/P0001  & n6331 ;
  assign n7945 = ~n7943 & ~n7944 ;
  assign n7946 = \u7_mem_reg[3][20]/NET0131  & ~n6331 ;
  assign n7947 = \u12_dout_reg[20]/P0001  & n6331 ;
  assign n7948 = ~n7946 & ~n7947 ;
  assign n7949 = \u7_mem_reg[3][21]/NET0131  & ~n6331 ;
  assign n7950 = \u12_dout_reg[21]/P0001  & n6331 ;
  assign n7951 = ~n7949 & ~n7950 ;
  assign n7952 = \u7_mem_reg[3][22]/NET0131  & ~n6331 ;
  assign n7953 = \u12_dout_reg[22]/P0001  & n6331 ;
  assign n7954 = ~n7952 & ~n7953 ;
  assign n7955 = \u7_mem_reg[3][23]/NET0131  & ~n6331 ;
  assign n7956 = \u12_dout_reg[23]/P0001  & n6331 ;
  assign n7957 = ~n7955 & ~n7956 ;
  assign n7958 = \u7_mem_reg[3][24]/NET0131  & ~n6331 ;
  assign n7959 = \u12_dout_reg[24]/P0001  & n6331 ;
  assign n7960 = ~n7958 & ~n7959 ;
  assign n7961 = \u7_mem_reg[3][25]/NET0131  & ~n6331 ;
  assign n7962 = \u12_dout_reg[25]/P0001  & n6331 ;
  assign n7963 = ~n7961 & ~n7962 ;
  assign n7964 = \u7_mem_reg[3][26]/NET0131  & ~n6331 ;
  assign n7965 = \u12_dout_reg[26]/P0001  & n6331 ;
  assign n7966 = ~n7964 & ~n7965 ;
  assign n7967 = \u7_mem_reg[3][27]/NET0131  & ~n6331 ;
  assign n7968 = \u12_dout_reg[27]/P0001  & n6331 ;
  assign n7969 = ~n7967 & ~n7968 ;
  assign n7970 = \u7_mem_reg[3][28]/NET0131  & ~n6331 ;
  assign n7971 = \u12_dout_reg[28]/P0001  & n6331 ;
  assign n7972 = ~n7970 & ~n7971 ;
  assign n7973 = \u7_mem_reg[3][29]/NET0131  & ~n6331 ;
  assign n7974 = \u12_dout_reg[29]/P0001  & n6331 ;
  assign n7975 = ~n7973 & ~n7974 ;
  assign n7976 = \u7_mem_reg[3][2]/NET0131  & ~n6331 ;
  assign n7977 = \u12_dout_reg[2]/P0001  & n6331 ;
  assign n7978 = ~n7976 & ~n7977 ;
  assign n7979 = \u7_mem_reg[3][30]/NET0131  & ~n6331 ;
  assign n7980 = \u12_dout_reg[30]/P0001  & n6331 ;
  assign n7981 = ~n7979 & ~n7980 ;
  assign n7982 = \u7_mem_reg[3][31]/NET0131  & ~n6331 ;
  assign n7983 = \u12_dout_reg[31]/P0001  & n6331 ;
  assign n7984 = ~n7982 & ~n7983 ;
  assign n7985 = \u7_mem_reg[3][3]/NET0131  & ~n6331 ;
  assign n7986 = \u12_dout_reg[3]/P0001  & n6331 ;
  assign n7987 = ~n7985 & ~n7986 ;
  assign n7988 = \u7_mem_reg[3][4]/NET0131  & ~n6331 ;
  assign n7989 = \u12_dout_reg[4]/P0001  & n6331 ;
  assign n7990 = ~n7988 & ~n7989 ;
  assign n7991 = \u7_mem_reg[3][5]/NET0131  & ~n6331 ;
  assign n7992 = \u12_dout_reg[5]/P0001  & n6331 ;
  assign n7993 = ~n7991 & ~n7992 ;
  assign n7994 = \u7_mem_reg[3][6]/NET0131  & ~n6331 ;
  assign n7995 = \u12_dout_reg[6]/P0001  & n6331 ;
  assign n7996 = ~n7994 & ~n7995 ;
  assign n7997 = \u7_mem_reg[3][7]/NET0131  & ~n6331 ;
  assign n7998 = \u12_dout_reg[7]/P0001  & n6331 ;
  assign n7999 = ~n7997 & ~n7998 ;
  assign n8000 = \u7_mem_reg[3][8]/NET0131  & ~n6331 ;
  assign n8001 = \u12_dout_reg[8]/P0001  & n6331 ;
  assign n8002 = ~n8000 & ~n8001 ;
  assign n8003 = \u7_mem_reg[3][9]/NET0131  & ~n6331 ;
  assign n8004 = \u12_dout_reg[9]/P0001  & n6331 ;
  assign n8005 = ~n8003 & ~n8004 ;
  assign n8006 = \u3_mem_reg[2][17]/NET0131  & ~n6583 ;
  assign n8007 = \u12_dout_reg[17]/P0001  & n6583 ;
  assign n8008 = ~n8006 & ~n8007 ;
  assign n8009 = \u8_mem_reg[1][0]/NET0131  & ~n6629 ;
  assign n8010 = \u12_dout_reg[0]/P0001  & n6629 ;
  assign n8011 = ~n8009 & ~n8010 ;
  assign n8012 = \u8_mem_reg[1][10]/NET0131  & ~n6629 ;
  assign n8013 = \u12_dout_reg[10]/P0001  & n6629 ;
  assign n8014 = ~n8012 & ~n8013 ;
  assign n8015 = \u8_mem_reg[1][11]/NET0131  & ~n6629 ;
  assign n8016 = \u12_dout_reg[11]/P0001  & n6629 ;
  assign n8017 = ~n8015 & ~n8016 ;
  assign n8018 = \u8_mem_reg[1][12]/NET0131  & ~n6629 ;
  assign n8019 = \u12_dout_reg[12]/P0001  & n6629 ;
  assign n8020 = ~n8018 & ~n8019 ;
  assign n8021 = \u8_mem_reg[1][13]/NET0131  & ~n6629 ;
  assign n8022 = \u12_dout_reg[13]/P0001  & n6629 ;
  assign n8023 = ~n8021 & ~n8022 ;
  assign n8024 = \u8_mem_reg[1][14]/NET0131  & ~n6629 ;
  assign n8025 = \u12_dout_reg[14]/P0001  & n6629 ;
  assign n8026 = ~n8024 & ~n8025 ;
  assign n8027 = \u8_mem_reg[1][15]/NET0131  & ~n6629 ;
  assign n8028 = \u12_dout_reg[15]/P0001  & n6629 ;
  assign n8029 = ~n8027 & ~n8028 ;
  assign n8030 = \u8_mem_reg[1][16]/NET0131  & ~n6629 ;
  assign n8031 = \u12_dout_reg[16]/P0001  & n6629 ;
  assign n8032 = ~n8030 & ~n8031 ;
  assign n8033 = \u8_mem_reg[1][17]/NET0131  & ~n6629 ;
  assign n8034 = \u12_dout_reg[17]/P0001  & n6629 ;
  assign n8035 = ~n8033 & ~n8034 ;
  assign n8036 = \u8_mem_reg[1][18]/NET0131  & ~n6629 ;
  assign n8037 = \u12_dout_reg[18]/P0001  & n6629 ;
  assign n8038 = ~n8036 & ~n8037 ;
  assign n8039 = \u8_mem_reg[1][19]/NET0131  & ~n6629 ;
  assign n8040 = \u12_dout_reg[19]/P0001  & n6629 ;
  assign n8041 = ~n8039 & ~n8040 ;
  assign n8042 = \u8_mem_reg[1][1]/NET0131  & ~n6629 ;
  assign n8043 = \u12_dout_reg[1]/P0001  & n6629 ;
  assign n8044 = ~n8042 & ~n8043 ;
  assign n8045 = \u8_mem_reg[1][20]/NET0131  & ~n6629 ;
  assign n8046 = \u12_dout_reg[20]/P0001  & n6629 ;
  assign n8047 = ~n8045 & ~n8046 ;
  assign n8048 = \u8_mem_reg[1][21]/NET0131  & ~n6629 ;
  assign n8049 = \u12_dout_reg[21]/P0001  & n6629 ;
  assign n8050 = ~n8048 & ~n8049 ;
  assign n8051 = \u8_mem_reg[1][22]/NET0131  & ~n6629 ;
  assign n8052 = \u12_dout_reg[22]/P0001  & n6629 ;
  assign n8053 = ~n8051 & ~n8052 ;
  assign n8054 = \u8_mem_reg[1][23]/NET0131  & ~n6629 ;
  assign n8055 = \u12_dout_reg[23]/P0001  & n6629 ;
  assign n8056 = ~n8054 & ~n8055 ;
  assign n8057 = \u8_mem_reg[1][24]/NET0131  & ~n6629 ;
  assign n8058 = \u12_dout_reg[24]/P0001  & n6629 ;
  assign n8059 = ~n8057 & ~n8058 ;
  assign n8060 = \u8_mem_reg[1][25]/NET0131  & ~n6629 ;
  assign n8061 = \u12_dout_reg[25]/P0001  & n6629 ;
  assign n8062 = ~n8060 & ~n8061 ;
  assign n8063 = \u3_mem_reg[1][0]/NET0131  & ~n6489 ;
  assign n8064 = \u12_dout_reg[0]/P0001  & n6489 ;
  assign n8065 = ~n8063 & ~n8064 ;
  assign n8066 = \u8_mem_reg[1][26]/NET0131  & ~n6629 ;
  assign n8067 = \u12_dout_reg[26]/P0001  & n6629 ;
  assign n8068 = ~n8066 & ~n8067 ;
  assign n8069 = \u8_mem_reg[1][27]/NET0131  & ~n6629 ;
  assign n8070 = \u12_dout_reg[27]/P0001  & n6629 ;
  assign n8071 = ~n8069 & ~n8070 ;
  assign n8072 = \u3_mem_reg[1][10]/NET0131  & ~n6489 ;
  assign n8073 = \u12_dout_reg[10]/P0001  & n6489 ;
  assign n8074 = ~n8072 & ~n8073 ;
  assign n8075 = \u8_mem_reg[1][29]/NET0131  & ~n6629 ;
  assign n8076 = \u12_dout_reg[29]/P0001  & n6629 ;
  assign n8077 = ~n8075 & ~n8076 ;
  assign n8078 = \u3_mem_reg[1][11]/NET0131  & ~n6489 ;
  assign n8079 = \u12_dout_reg[11]/P0001  & n6489 ;
  assign n8080 = ~n8078 & ~n8079 ;
  assign n8081 = \u8_mem_reg[1][2]/NET0131  & ~n6629 ;
  assign n8082 = \u12_dout_reg[2]/P0001  & n6629 ;
  assign n8083 = ~n8081 & ~n8082 ;
  assign n8084 = \u8_mem_reg[1][30]/NET0131  & ~n6629 ;
  assign n8085 = \u12_dout_reg[30]/P0001  & n6629 ;
  assign n8086 = ~n8084 & ~n8085 ;
  assign n8087 = \u3_mem_reg[1][12]/NET0131  & ~n6489 ;
  assign n8088 = \u12_dout_reg[12]/P0001  & n6489 ;
  assign n8089 = ~n8087 & ~n8088 ;
  assign n8090 = \u8_mem_reg[3][11]/NET0131  & ~n6301 ;
  assign n8091 = \u12_dout_reg[11]/P0001  & n6301 ;
  assign n8092 = ~n8090 & ~n8091 ;
  assign n8093 = \u8_mem_reg[1][3]/NET0131  & ~n6629 ;
  assign n8094 = \u12_dout_reg[3]/P0001  & n6629 ;
  assign n8095 = ~n8093 & ~n8094 ;
  assign n8096 = \u3_mem_reg[1][13]/NET0131  & ~n6489 ;
  assign n8097 = \u12_dout_reg[13]/P0001  & n6489 ;
  assign n8098 = ~n8096 & ~n8097 ;
  assign n8099 = \u8_mem_reg[1][5]/NET0131  & ~n6629 ;
  assign n8100 = \u12_dout_reg[5]/P0001  & n6629 ;
  assign n8101 = ~n8099 & ~n8100 ;
  assign n8102 = \u8_mem_reg[1][7]/NET0131  & ~n6629 ;
  assign n8103 = \u12_dout_reg[7]/P0001  & n6629 ;
  assign n8104 = ~n8102 & ~n8103 ;
  assign n8105 = \u3_mem_reg[1][15]/NET0131  & ~n6489 ;
  assign n8106 = \u12_dout_reg[15]/P0001  & n6489 ;
  assign n8107 = ~n8105 & ~n8106 ;
  assign n8108 = \u8_mem_reg[1][8]/NET0131  & ~n6629 ;
  assign n8109 = \u12_dout_reg[8]/P0001  & n6629 ;
  assign n8110 = ~n8108 & ~n8109 ;
  assign n8111 = \u8_mem_reg[1][9]/NET0131  & ~n6629 ;
  assign n8112 = \u12_dout_reg[9]/P0001  & n6629 ;
  assign n8113 = ~n8111 & ~n8112 ;
  assign n8114 = \u3_mem_reg[1][16]/NET0131  & ~n6489 ;
  assign n8115 = \u12_dout_reg[16]/P0001  & n6489 ;
  assign n8116 = ~n8114 & ~n8115 ;
  assign n8117 = \u8_mem_reg[2][0]/NET0131  & ~n6485 ;
  assign n8118 = \u12_dout_reg[0]/P0001  & n6485 ;
  assign n8119 = ~n8117 & ~n8118 ;
  assign n8120 = \u8_mem_reg[2][10]/NET0131  & ~n6485 ;
  assign n8121 = \u12_dout_reg[10]/P0001  & n6485 ;
  assign n8122 = ~n8120 & ~n8121 ;
  assign n8123 = \u3_mem_reg[1][17]/NET0131  & ~n6489 ;
  assign n8124 = \u12_dout_reg[17]/P0001  & n6489 ;
  assign n8125 = ~n8123 & ~n8124 ;
  assign n8126 = \u8_mem_reg[2][11]/NET0131  & ~n6485 ;
  assign n8127 = \u12_dout_reg[11]/P0001  & n6485 ;
  assign n8128 = ~n8126 & ~n8127 ;
  assign n8129 = \u8_mem_reg[2][12]/NET0131  & ~n6485 ;
  assign n8130 = \u12_dout_reg[12]/P0001  & n6485 ;
  assign n8131 = ~n8129 & ~n8130 ;
  assign n8132 = \u3_mem_reg[1][18]/NET0131  & ~n6489 ;
  assign n8133 = \u12_dout_reg[18]/P0001  & n6489 ;
  assign n8134 = ~n8132 & ~n8133 ;
  assign n8135 = \u8_mem_reg[2][13]/NET0131  & ~n6485 ;
  assign n8136 = \u12_dout_reg[13]/P0001  & n6485 ;
  assign n8137 = ~n8135 & ~n8136 ;
  assign n8138 = \u8_mem_reg[2][14]/NET0131  & ~n6485 ;
  assign n8139 = \u12_dout_reg[14]/P0001  & n6485 ;
  assign n8140 = ~n8138 & ~n8139 ;
  assign n8141 = \u3_mem_reg[1][19]/NET0131  & ~n6489 ;
  assign n8142 = \u12_dout_reg[19]/P0001  & n6489 ;
  assign n8143 = ~n8141 & ~n8142 ;
  assign n8144 = \u8_mem_reg[2][15]/NET0131  & ~n6485 ;
  assign n8145 = \u12_dout_reg[15]/P0001  & n6485 ;
  assign n8146 = ~n8144 & ~n8145 ;
  assign n8147 = \u8_mem_reg[2][16]/NET0131  & ~n6485 ;
  assign n8148 = \u12_dout_reg[16]/P0001  & n6485 ;
  assign n8149 = ~n8147 & ~n8148 ;
  assign n8150 = \u8_mem_reg[2][17]/NET0131  & ~n6485 ;
  assign n8151 = \u12_dout_reg[17]/P0001  & n6485 ;
  assign n8152 = ~n8150 & ~n8151 ;
  assign n8153 = \u8_mem_reg[2][18]/NET0131  & ~n6485 ;
  assign n8154 = \u12_dout_reg[18]/P0001  & n6485 ;
  assign n8155 = ~n8153 & ~n8154 ;
  assign n8156 = \u3_mem_reg[1][20]/NET0131  & ~n6489 ;
  assign n8157 = \u12_dout_reg[20]/P0001  & n6489 ;
  assign n8158 = ~n8156 & ~n8157 ;
  assign n8159 = \u8_mem_reg[2][19]/NET0131  & ~n6485 ;
  assign n8160 = \u12_dout_reg[19]/P0001  & n6485 ;
  assign n8161 = ~n8159 & ~n8160 ;
  assign n8162 = \u8_mem_reg[2][1]/NET0131  & ~n6485 ;
  assign n8163 = \u12_dout_reg[1]/P0001  & n6485 ;
  assign n8164 = ~n8162 & ~n8163 ;
  assign n8165 = \u3_mem_reg[1][21]/NET0131  & ~n6489 ;
  assign n8166 = \u12_dout_reg[21]/P0001  & n6489 ;
  assign n8167 = ~n8165 & ~n8166 ;
  assign n8168 = \u8_mem_reg[2][20]/NET0131  & ~n6485 ;
  assign n8169 = \u12_dout_reg[20]/P0001  & n6485 ;
  assign n8170 = ~n8168 & ~n8169 ;
  assign n8171 = \u8_mem_reg[2][21]/NET0131  & ~n6485 ;
  assign n8172 = \u12_dout_reg[21]/P0001  & n6485 ;
  assign n8173 = ~n8171 & ~n8172 ;
  assign n8174 = \u3_mem_reg[1][22]/NET0131  & ~n6489 ;
  assign n8175 = \u12_dout_reg[22]/P0001  & n6489 ;
  assign n8176 = ~n8174 & ~n8175 ;
  assign n8177 = \u8_mem_reg[2][22]/NET0131  & ~n6485 ;
  assign n8178 = \u12_dout_reg[22]/P0001  & n6485 ;
  assign n8179 = ~n8177 & ~n8178 ;
  assign n8180 = \u8_mem_reg[2][23]/NET0131  & ~n6485 ;
  assign n8181 = \u12_dout_reg[23]/P0001  & n6485 ;
  assign n8182 = ~n8180 & ~n8181 ;
  assign n8183 = \u8_mem_reg[2][24]/NET0131  & ~n6485 ;
  assign n8184 = \u12_dout_reg[24]/P0001  & n6485 ;
  assign n8185 = ~n8183 & ~n8184 ;
  assign n8186 = \u8_mem_reg[2][25]/NET0131  & ~n6485 ;
  assign n8187 = \u12_dout_reg[25]/P0001  & n6485 ;
  assign n8188 = ~n8186 & ~n8187 ;
  assign n8189 = \u3_mem_reg[1][24]/NET0131  & ~n6489 ;
  assign n8190 = \u12_dout_reg[24]/P0001  & n6489 ;
  assign n8191 = ~n8189 & ~n8190 ;
  assign n8192 = \u8_mem_reg[2][26]/NET0131  & ~n6485 ;
  assign n8193 = \u12_dout_reg[26]/P0001  & n6485 ;
  assign n8194 = ~n8192 & ~n8193 ;
  assign n8195 = \u8_mem_reg[2][27]/NET0131  & ~n6485 ;
  assign n8196 = \u12_dout_reg[27]/P0001  & n6485 ;
  assign n8197 = ~n8195 & ~n8196 ;
  assign n8198 = \u3_mem_reg[1][25]/NET0131  & ~n6489 ;
  assign n8199 = \u12_dout_reg[25]/P0001  & n6489 ;
  assign n8200 = ~n8198 & ~n8199 ;
  assign n8201 = \u8_mem_reg[2][28]/NET0131  & ~n6485 ;
  assign n8202 = \u12_dout_reg[28]/P0001  & n6485 ;
  assign n8203 = ~n8201 & ~n8202 ;
  assign n8204 = \u8_mem_reg[2][29]/NET0131  & ~n6485 ;
  assign n8205 = \u12_dout_reg[29]/P0001  & n6485 ;
  assign n8206 = ~n8204 & ~n8205 ;
  assign n8207 = \u3_mem_reg[1][26]/NET0131  & ~n6489 ;
  assign n8208 = \u12_dout_reg[26]/P0001  & n6489 ;
  assign n8209 = ~n8207 & ~n8208 ;
  assign n8210 = \u8_mem_reg[2][2]/NET0131  & ~n6485 ;
  assign n8211 = \u12_dout_reg[2]/P0001  & n6485 ;
  assign n8212 = ~n8210 & ~n8211 ;
  assign n8213 = \u8_mem_reg[2][30]/NET0131  & ~n6485 ;
  assign n8214 = \u12_dout_reg[30]/P0001  & n6485 ;
  assign n8215 = ~n8213 & ~n8214 ;
  assign n8216 = \u8_mem_reg[2][31]/NET0131  & ~n6485 ;
  assign n8217 = \u12_dout_reg[31]/P0001  & n6485 ;
  assign n8218 = ~n8216 & ~n8217 ;
  assign n8219 = \u3_mem_reg[1][28]/NET0131  & ~n6489 ;
  assign n8220 = \u12_dout_reg[28]/P0001  & n6489 ;
  assign n8221 = ~n8219 & ~n8220 ;
  assign n8222 = \u8_mem_reg[2][4]/NET0131  & ~n6485 ;
  assign n8223 = \u12_dout_reg[4]/P0001  & n6485 ;
  assign n8224 = ~n8222 & ~n8223 ;
  assign n8225 = ~\u3_wp_reg[1]/NET0131  & n6407 ;
  assign n8226 = ~\u4_wp_reg[1]/NET0131  & n6411 ;
  assign n8227 = ~\u5_wp_reg[1]/NET0131  & n6415 ;
  assign n8228 = ~\u6_wp_reg[1]/NET0131  & n6419 ;
  assign n8229 = ~\u7_wp_reg[1]/NET0131  & n6423 ;
  assign n8230 = ~\u8_wp_reg[1]/NET0131  & n6403 ;
  assign n8231 = \u13_ints_r_reg[0]/NET0131  & n2741 ;
  assign n8232 = \u13_occ0_r_reg[0]/NET0131  & n6151 ;
  assign n8237 = ~n8231 & ~n8232 ;
  assign n8233 = \u13_intm_r_reg[0]/NET0131  & n6153 ;
  assign n8234 = \u13_icc_r_reg[0]/NET0131  & n6157 ;
  assign n8238 = ~n8233 & ~n8234 ;
  assign n8235 = \u13_occ1_r_reg[0]/NET0131  & n6147 ;
  assign n8236 = \u15_crac_din_reg[0]/NET0131  & n6159 ;
  assign n8239 = ~n8235 & ~n8236 ;
  assign n8240 = n8238 & n8239 ;
  assign n8241 = n8237 & n8240 ;
  assign n8242 = n6146 & ~n8241 ;
  assign n8245 = \u11_dout_reg[0]/P0001  & n6145 ;
  assign n8243 = \u9_dout_reg[0]/P0001  & n6168 ;
  assign n8244 = \u10_dout_reg[0]/P0001  & n6170 ;
  assign n8246 = ~n8243 & ~n8244 ;
  assign n8247 = ~n8245 & n8246 ;
  assign n8248 = ~n8242 & n8247 ;
  assign n8249 = \u13_ints_r_reg[10]/NET0131  & n2741 ;
  assign n8250 = \u13_occ0_r_reg[10]/NET0131  & n6151 ;
  assign n8255 = ~n8249 & ~n8250 ;
  assign n8251 = \u13_intm_r_reg[10]/NET0131  & n6153 ;
  assign n8252 = \u13_icc_r_reg[10]/NET0131  & n6157 ;
  assign n8256 = ~n8251 & ~n8252 ;
  assign n8253 = \u13_occ1_r_reg[10]/NET0131  & n6147 ;
  assign n8254 = \u15_crac_din_reg[10]/NET0131  & n6159 ;
  assign n8257 = ~n8253 & ~n8254 ;
  assign n8258 = n8256 & n8257 ;
  assign n8259 = n8255 & n8258 ;
  assign n8260 = n6146 & ~n8259 ;
  assign n8263 = \u11_dout_reg[10]/P0001  & n6145 ;
  assign n8261 = \u9_dout_reg[10]/P0001  & n6168 ;
  assign n8262 = \u10_dout_reg[10]/P0001  & n6170 ;
  assign n8264 = ~n8261 & ~n8262 ;
  assign n8265 = ~n8263 & n8264 ;
  assign n8266 = ~n8260 & n8265 ;
  assign n8267 = \u13_ints_r_reg[11]/NET0131  & n2741 ;
  assign n8268 = \u13_occ0_r_reg[11]/NET0131  & n6151 ;
  assign n8273 = ~n8267 & ~n8268 ;
  assign n8269 = \u13_intm_r_reg[11]/NET0131  & n6153 ;
  assign n8270 = \u13_icc_r_reg[11]/NET0131  & n6157 ;
  assign n8274 = ~n8269 & ~n8270 ;
  assign n8271 = \u13_occ1_r_reg[11]/NET0131  & n6147 ;
  assign n8272 = \u15_crac_din_reg[11]/NET0131  & n6159 ;
  assign n8275 = ~n8271 & ~n8272 ;
  assign n8276 = n8274 & n8275 ;
  assign n8277 = n8273 & n8276 ;
  assign n8278 = n6146 & ~n8277 ;
  assign n8281 = \u11_dout_reg[11]/P0001  & n6145 ;
  assign n8279 = \u9_dout_reg[11]/P0001  & n6168 ;
  assign n8280 = \u10_dout_reg[11]/P0001  & n6170 ;
  assign n8282 = ~n8279 & ~n8280 ;
  assign n8283 = ~n8281 & n8282 ;
  assign n8284 = ~n8278 & n8283 ;
  assign n8285 = \u13_ints_r_reg[12]/NET0131  & n2741 ;
  assign n8286 = \u13_occ0_r_reg[12]/NET0131  & n6151 ;
  assign n8291 = ~n8285 & ~n8286 ;
  assign n8287 = \u13_intm_r_reg[12]/NET0131  & n6153 ;
  assign n8288 = \u13_icc_r_reg[12]/NET0131  & n6157 ;
  assign n8292 = ~n8287 & ~n8288 ;
  assign n8289 = \u13_occ1_r_reg[12]/NET0131  & n6147 ;
  assign n8290 = \u15_crac_din_reg[12]/NET0131  & n6159 ;
  assign n8293 = ~n8289 & ~n8290 ;
  assign n8294 = n8292 & n8293 ;
  assign n8295 = n8291 & n8294 ;
  assign n8296 = n6146 & ~n8295 ;
  assign n8299 = \u11_dout_reg[12]/P0001  & n6145 ;
  assign n8297 = \u9_dout_reg[12]/P0001  & n6168 ;
  assign n8298 = \u10_dout_reg[12]/P0001  & n6170 ;
  assign n8300 = ~n8297 & ~n8298 ;
  assign n8301 = ~n8299 & n8300 ;
  assign n8302 = ~n8296 & n8301 ;
  assign n8303 = \u13_ints_r_reg[13]/NET0131  & n2741 ;
  assign n8304 = \u13_occ0_r_reg[13]/NET0131  & n6151 ;
  assign n8309 = ~n8303 & ~n8304 ;
  assign n8305 = \u13_intm_r_reg[13]/NET0131  & n6153 ;
  assign n8306 = \u13_icc_r_reg[13]/NET0131  & n6157 ;
  assign n8310 = ~n8305 & ~n8306 ;
  assign n8307 = \u13_occ1_r_reg[13]/NET0131  & n6147 ;
  assign n8308 = \u15_crac_din_reg[13]/NET0131  & n6159 ;
  assign n8311 = ~n8307 & ~n8308 ;
  assign n8312 = n8310 & n8311 ;
  assign n8313 = n8309 & n8312 ;
  assign n8314 = n6146 & ~n8313 ;
  assign n8317 = \u11_dout_reg[13]/P0001  & n6145 ;
  assign n8315 = \u9_dout_reg[13]/P0001  & n6168 ;
  assign n8316 = \u10_dout_reg[13]/P0001  & n6170 ;
  assign n8318 = ~n8315 & ~n8316 ;
  assign n8319 = ~n8317 & n8318 ;
  assign n8320 = ~n8314 & n8319 ;
  assign n8321 = \u13_ints_r_reg[14]/NET0131  & n2741 ;
  assign n8322 = \u13_occ0_r_reg[14]/NET0131  & n6151 ;
  assign n8327 = ~n8321 & ~n8322 ;
  assign n8323 = \u13_intm_r_reg[14]/NET0131  & n6153 ;
  assign n8324 = \u13_icc_r_reg[14]/NET0131  & n6157 ;
  assign n8328 = ~n8323 & ~n8324 ;
  assign n8325 = \u13_occ1_r_reg[14]/NET0131  & n6147 ;
  assign n8326 = \u15_crac_din_reg[14]/NET0131  & n6159 ;
  assign n8329 = ~n8325 & ~n8326 ;
  assign n8330 = n8328 & n8329 ;
  assign n8331 = n8327 & n8330 ;
  assign n8332 = n6146 & ~n8331 ;
  assign n8335 = \u11_dout_reg[14]/P0001  & n6145 ;
  assign n8333 = \u9_dout_reg[14]/P0001  & n6168 ;
  assign n8334 = \u10_dout_reg[14]/P0001  & n6170 ;
  assign n8336 = ~n8333 & ~n8334 ;
  assign n8337 = ~n8335 & n8336 ;
  assign n8338 = ~n8332 & n8337 ;
  assign n8339 = \u13_intm_r_reg[15]/NET0131  & n6153 ;
  assign n8340 = \u13_occ1_r_reg[15]/NET0131  & n6147 ;
  assign n8345 = ~n8339 & ~n8340 ;
  assign n8341 = \u13_occ0_r_reg[15]/NET0131  & n6151 ;
  assign n8342 = \u13_icc_r_reg[15]/NET0131  & n6157 ;
  assign n8346 = ~n8341 & ~n8342 ;
  assign n8343 = \u13_ints_r_reg[15]/NET0131  & n2741 ;
  assign n8344 = \u15_crac_din_reg[15]/NET0131  & n6159 ;
  assign n8347 = ~n8343 & ~n8344 ;
  assign n8348 = n8346 & n8347 ;
  assign n8349 = n8345 & n8348 ;
  assign n8350 = n6146 & ~n8349 ;
  assign n8353 = \u11_dout_reg[15]/P0001  & n6145 ;
  assign n8351 = \u9_dout_reg[15]/P0001  & n6168 ;
  assign n8352 = \u10_dout_reg[15]/P0001  & n6170 ;
  assign n8354 = ~n8351 & ~n8352 ;
  assign n8355 = ~n8353 & n8354 ;
  assign n8356 = ~n8350 & n8355 ;
  assign n8357 = \u13_ints_r_reg[2]/NET0131  & n2741 ;
  assign n8358 = \u13_occ0_r_reg[2]/NET0131  & n6151 ;
  assign n8363 = ~n8357 & ~n8358 ;
  assign n8359 = \u13_intm_r_reg[2]/NET0131  & n6153 ;
  assign n8360 = \u13_icc_r_reg[2]/NET0131  & n6157 ;
  assign n8364 = ~n8359 & ~n8360 ;
  assign n8361 = \u13_occ1_r_reg[2]/NET0131  & n6147 ;
  assign n8362 = \u15_crac_din_reg[2]/NET0131  & n6159 ;
  assign n8365 = ~n8361 & ~n8362 ;
  assign n8366 = n8364 & n8365 ;
  assign n8367 = n8363 & n8366 ;
  assign n8368 = n6146 & ~n8367 ;
  assign n8371 = \u11_dout_reg[2]/P0001  & n6145 ;
  assign n8369 = \u9_dout_reg[2]/P0001  & n6168 ;
  assign n8370 = \u10_dout_reg[2]/P0001  & n6170 ;
  assign n8372 = ~n8369 & ~n8370 ;
  assign n8373 = ~n8371 & n8372 ;
  assign n8374 = ~n8368 & n8373 ;
  assign n8375 = \u13_ints_r_reg[3]/NET0131  & n2741 ;
  assign n8376 = \u13_occ0_r_reg[3]/NET0131  & n6151 ;
  assign n8381 = ~n8375 & ~n8376 ;
  assign n8377 = \u13_intm_r_reg[3]/NET0131  & n6153 ;
  assign n8378 = \u13_icc_r_reg[3]/NET0131  & n6157 ;
  assign n8382 = ~n8377 & ~n8378 ;
  assign n8379 = \u13_occ1_r_reg[3]/NET0131  & n6147 ;
  assign n8380 = \u15_crac_din_reg[3]/NET0131  & n6159 ;
  assign n8383 = ~n8379 & ~n8380 ;
  assign n8384 = n8382 & n8383 ;
  assign n8385 = n8381 & n8384 ;
  assign n8386 = n6146 & ~n8385 ;
  assign n8389 = \u11_dout_reg[3]/P0001  & n6145 ;
  assign n8387 = \u9_dout_reg[3]/P0001  & n6168 ;
  assign n8388 = \u10_dout_reg[3]/P0001  & n6170 ;
  assign n8390 = ~n8387 & ~n8388 ;
  assign n8391 = ~n8389 & n8390 ;
  assign n8392 = ~n8386 & n8391 ;
  assign n8393 = \u13_ints_r_reg[4]/NET0131  & n2741 ;
  assign n8394 = \u13_occ0_r_reg[4]/NET0131  & n6151 ;
  assign n8399 = ~n8393 & ~n8394 ;
  assign n8395 = \u13_intm_r_reg[4]/NET0131  & n6153 ;
  assign n8396 = \u13_icc_r_reg[4]/NET0131  & n6157 ;
  assign n8400 = ~n8395 & ~n8396 ;
  assign n8397 = \u13_occ1_r_reg[4]/NET0131  & n6147 ;
  assign n8398 = \u15_crac_din_reg[4]/NET0131  & n6159 ;
  assign n8401 = ~n8397 & ~n8398 ;
  assign n8402 = n8400 & n8401 ;
  assign n8403 = n8399 & n8402 ;
  assign n8404 = n6146 & ~n8403 ;
  assign n8407 = \u11_dout_reg[4]/P0001  & n6145 ;
  assign n8405 = \u9_dout_reg[4]/P0001  & n6168 ;
  assign n8406 = \u10_dout_reg[4]/P0001  & n6170 ;
  assign n8408 = ~n8405 & ~n8406 ;
  assign n8409 = ~n8407 & n8408 ;
  assign n8410 = ~n8404 & n8409 ;
  assign n8411 = \u13_ints_r_reg[5]/NET0131  & n2741 ;
  assign n8412 = \u13_occ0_r_reg[5]/NET0131  & n6151 ;
  assign n8417 = ~n8411 & ~n8412 ;
  assign n8413 = \u13_intm_r_reg[5]/NET0131  & n6153 ;
  assign n8414 = \u13_icc_r_reg[5]/NET0131  & n6157 ;
  assign n8418 = ~n8413 & ~n8414 ;
  assign n8415 = \u13_occ1_r_reg[5]/NET0131  & n6147 ;
  assign n8416 = \u15_crac_din_reg[5]/NET0131  & n6159 ;
  assign n8419 = ~n8415 & ~n8416 ;
  assign n8420 = n8418 & n8419 ;
  assign n8421 = n8417 & n8420 ;
  assign n8422 = n6146 & ~n8421 ;
  assign n8425 = \u11_dout_reg[5]/P0001  & n6145 ;
  assign n8423 = \u9_dout_reg[5]/P0001  & n6168 ;
  assign n8424 = \u10_dout_reg[5]/P0001  & n6170 ;
  assign n8426 = ~n8423 & ~n8424 ;
  assign n8427 = ~n8425 & n8426 ;
  assign n8428 = ~n8422 & n8427 ;
  assign n8429 = \u13_ints_r_reg[6]/NET0131  & n2741 ;
  assign n8430 = \u13_occ0_r_reg[6]/NET0131  & n6151 ;
  assign n8435 = ~n8429 & ~n8430 ;
  assign n8431 = \u13_intm_r_reg[6]/NET0131  & n6153 ;
  assign n8432 = \u13_icc_r_reg[6]/NET0131  & n6157 ;
  assign n8436 = ~n8431 & ~n8432 ;
  assign n8433 = \u13_occ1_r_reg[6]/NET0131  & n6147 ;
  assign n8434 = \u15_crac_din_reg[6]/NET0131  & n6159 ;
  assign n8437 = ~n8433 & ~n8434 ;
  assign n8438 = n8436 & n8437 ;
  assign n8439 = n8435 & n8438 ;
  assign n8440 = n6146 & ~n8439 ;
  assign n8443 = \u11_dout_reg[6]/P0001  & n6145 ;
  assign n8441 = \u9_dout_reg[6]/P0001  & n6168 ;
  assign n8442 = \u10_dout_reg[6]/P0001  & n6170 ;
  assign n8444 = ~n8441 & ~n8442 ;
  assign n8445 = ~n8443 & n8444 ;
  assign n8446 = ~n8440 & n8445 ;
  assign n8447 = \u13_intm_r_reg[7]/NET0131  & n6153 ;
  assign n8448 = \u13_occ1_r_reg[7]/NET0131  & n6147 ;
  assign n8453 = ~n8447 & ~n8448 ;
  assign n8449 = \u13_occ0_r_reg[7]/NET0131  & n6151 ;
  assign n8450 = \u13_icc_r_reg[7]/NET0131  & n6157 ;
  assign n8454 = ~n8449 & ~n8450 ;
  assign n8451 = \u13_ints_r_reg[7]/NET0131  & n2741 ;
  assign n8452 = \u15_crac_din_reg[7]/NET0131  & n6159 ;
  assign n8455 = ~n8451 & ~n8452 ;
  assign n8456 = n8454 & n8455 ;
  assign n8457 = n8453 & n8456 ;
  assign n8458 = n6146 & ~n8457 ;
  assign n8461 = \u11_dout_reg[7]/P0001  & n6145 ;
  assign n8459 = \u9_dout_reg[7]/P0001  & n6168 ;
  assign n8460 = \u10_dout_reg[7]/P0001  & n6170 ;
  assign n8462 = ~n8459 & ~n8460 ;
  assign n8463 = ~n8461 & n8462 ;
  assign n8464 = ~n8458 & n8463 ;
  assign n8465 = \u13_ints_r_reg[8]/NET0131  & n2741 ;
  assign n8466 = \u13_occ0_r_reg[8]/NET0131  & n6151 ;
  assign n8471 = ~n8465 & ~n8466 ;
  assign n8467 = \u13_intm_r_reg[8]/NET0131  & n6153 ;
  assign n8468 = \u13_icc_r_reg[8]/NET0131  & n6157 ;
  assign n8472 = ~n8467 & ~n8468 ;
  assign n8469 = \u13_occ1_r_reg[8]/NET0131  & n6147 ;
  assign n8470 = \u15_crac_din_reg[8]/NET0131  & n6159 ;
  assign n8473 = ~n8469 & ~n8470 ;
  assign n8474 = n8472 & n8473 ;
  assign n8475 = n8471 & n8474 ;
  assign n8476 = n6146 & ~n8475 ;
  assign n8479 = \u11_dout_reg[8]/P0001  & n6145 ;
  assign n8477 = \u9_dout_reg[8]/P0001  & n6168 ;
  assign n8478 = \u10_dout_reg[8]/P0001  & n6170 ;
  assign n8480 = ~n8477 & ~n8478 ;
  assign n8481 = ~n8479 & n8480 ;
  assign n8482 = ~n8476 & n8481 ;
  assign n8483 = \u13_ints_r_reg[9]/NET0131  & n2741 ;
  assign n8484 = \u13_occ0_r_reg[9]/NET0131  & n6151 ;
  assign n8489 = ~n8483 & ~n8484 ;
  assign n8485 = \u13_intm_r_reg[9]/NET0131  & n6153 ;
  assign n8486 = \u13_icc_r_reg[9]/NET0131  & n6157 ;
  assign n8490 = ~n8485 & ~n8486 ;
  assign n8487 = \u13_occ1_r_reg[9]/NET0131  & n6147 ;
  assign n8488 = \u15_crac_din_reg[9]/NET0131  & n6159 ;
  assign n8491 = ~n8487 & ~n8488 ;
  assign n8492 = n8490 & n8491 ;
  assign n8493 = n8489 & n8492 ;
  assign n8494 = n6146 & ~n8493 ;
  assign n8497 = \u11_dout_reg[9]/P0001  & n6145 ;
  assign n8495 = \u9_dout_reg[9]/P0001  & n6168 ;
  assign n8496 = \u10_dout_reg[9]/P0001  & n6170 ;
  assign n8498 = ~n8495 & ~n8496 ;
  assign n8499 = ~n8497 & n8498 ;
  assign n8500 = ~n8494 & n8499 ;
  assign n8501 = \u12_rf_we_reg/P0001  & n6159 ;
  assign n8502 = \u12_rf_we_reg/P0001  & n6157 ;
  assign n8503 = \u12_rf_we_reg/P0001  & n6153 ;
  assign n8504 = \u12_rf_we_reg/P0001  & n6151 ;
  assign n8505 = \u12_rf_we_reg/P0001  & n6147 ;
  assign n8506 = ~\u2_cnt_reg[4]/NET0131  & ~n6471 ;
  assign n8507 = ~n6472 & ~n8506 ;
  assign n8508 = ~suspended_o_pad & ~n8507 ;
  assign n8511 = n2765 & ~n6243 ;
  assign n8512 = ~n2760 & ~n6240 ;
  assign n8513 = ~n8511 & n8512 ;
  assign n8514 = \u4_rp_reg[0]/P0001  & ~n8513 ;
  assign n8517 = ~n6235 & ~n6239 ;
  assign n8509 = ~n6235 & ~n6236 ;
  assign n8510 = ~\u4_rp_reg[0]/P0001  & ~n8509 ;
  assign n8515 = \u4_rp_reg[0]/P0001  & n2765 ;
  assign n8516 = n6243 & ~n8515 ;
  assign n8518 = ~n8510 & ~n8516 ;
  assign n8519 = ~n8517 & n8518 ;
  assign n8520 = ~n8514 & n8519 ;
  assign n8523 = n2776 & ~n6256 ;
  assign n8524 = ~n2771 & ~n6253 ;
  assign n8525 = ~n8523 & n8524 ;
  assign n8526 = \u5_rp_reg[0]/P0001  & ~n8525 ;
  assign n8529 = ~n6248 & ~n6252 ;
  assign n8521 = ~n6248 & ~n6249 ;
  assign n8522 = ~\u5_rp_reg[0]/P0001  & ~n8521 ;
  assign n8527 = \u5_rp_reg[0]/P0001  & n2776 ;
  assign n8528 = n6256 & ~n8527 ;
  assign n8530 = ~n8522 & ~n8528 ;
  assign n8531 = ~n8529 & n8530 ;
  assign n8532 = ~n8526 & n8531 ;
  assign n8533 = ~\u14_crac_wr_r_reg/P0001  & ~\valid_s_reg/NET0131  ;
  assign n8534 = ~n6465 & ~n8533 ;
  assign n8537 = n6261 & n6266 ;
  assign n8538 = n6262 & ~n6266 ;
  assign n8539 = ~n8537 & ~n8538 ;
  assign n8540 = ~n2796 & ~n8539 ;
  assign n8541 = \u6_rp_reg[0]/P0001  & ~n8540 ;
  assign n8542 = ~\u6_rp_reg[0]/P0001  & ~n6267 ;
  assign n8535 = \u6_rp_reg[0]/P0001  & n2801 ;
  assign n8536 = ~n6270 & n8535 ;
  assign n8543 = n6270 & ~n8535 ;
  assign n8544 = ~n8536 & ~n8543 ;
  assign n8545 = ~n8542 & n8544 ;
  assign n8546 = ~n8541 & n8545 ;
  assign n8551 = ~n6277 & ~n6282 ;
  assign n8552 = \u7_rp_reg[1]/NET0131  & n6280 ;
  assign n8553 = \u7_rp_reg[0]/P0001  & ~n8552 ;
  assign n8554 = ~n8551 & ~n8553 ;
  assign n8555 = ~n2805 & ~n8551 ;
  assign n8556 = \u7_rp_reg[0]/P0001  & ~n8555 ;
  assign n8547 = \u7_rp_reg[0]/P0001  & n2981 ;
  assign n8548 = ~n6276 & ~n8547 ;
  assign n8549 = n6276 & n8547 ;
  assign n8550 = ~n8548 & ~n8549 ;
  assign n8557 = \u7_rp_reg[0]/P0001  & \u7_rp_reg[1]/NET0131  ;
  assign n8558 = ~n6280 & ~n8557 ;
  assign n8559 = ~n8550 & ~n8558 ;
  assign n8560 = ~n8556 & n8559 ;
  assign n8561 = ~n8554 & n8560 ;
  assign n8566 = ~n6225 & ~n6230 ;
  assign n8567 = \u3_rp_reg[1]/NET0131  & n6228 ;
  assign n8568 = \u3_rp_reg[0]/P0001  & ~n8567 ;
  assign n8569 = ~n8566 & ~n8568 ;
  assign n8570 = ~n2784 & ~n8566 ;
  assign n8571 = \u3_rp_reg[0]/P0001  & ~n8570 ;
  assign n8562 = \u3_rp_reg[0]/P0001  & n3009 ;
  assign n8563 = ~n6224 & ~n8562 ;
  assign n8564 = n6224 & n8562 ;
  assign n8565 = ~n8563 & ~n8564 ;
  assign n8572 = \u3_rp_reg[0]/P0001  & \u3_rp_reg[1]/NET0131  ;
  assign n8573 = ~n6228 & ~n8572 ;
  assign n8574 = ~n8565 & ~n8573 ;
  assign n8575 = ~n8571 & n8574 ;
  assign n8576 = ~n8569 & n8575 ;
  assign n8579 = n6287 & n6292 ;
  assign n8580 = n6288 & ~n6292 ;
  assign n8581 = ~n8579 & ~n8580 ;
  assign n8582 = ~n2160 & ~n8581 ;
  assign n8583 = \u8_rp_reg[0]/P0001  & ~n8582 ;
  assign n8584 = ~\u8_rp_reg[0]/P0001  & ~n6293 ;
  assign n8577 = \u8_rp_reg[0]/P0001  & n2163 ;
  assign n8578 = ~n6296 & n8577 ;
  assign n8585 = n6296 & ~n8577 ;
  assign n8586 = ~n8578 & ~n8585 ;
  assign n8587 = ~n8584 & n8586 ;
  assign n8588 = ~n8583 & n8587 ;
  assign n8589 = \u2_ld_reg/P0001  & \u8_dout_reg[1]/P0001  ;
  assign n8590 = \u0_slt9_r_reg[0]/P0001  & ~\u2_ld_reg/P0001  ;
  assign n8591 = ~n8589 & ~n8590 ;
  assign n8592 = \u12_i3_re_reg/NET0131  & \u9_rp_reg[0]/P0001  ;
  assign n8594 = \u9_rp_reg[1]/P0001  & n8592 ;
  assign n8593 = ~\u9_rp_reg[1]/P0001  & ~n8592 ;
  assign n8595 = \u13_icc_r_reg[0]/NET0131  & ~n8593 ;
  assign n8596 = ~n8594 & n8595 ;
  assign n8597 = \u10_rp_reg[0]/P0001  & \u12_i4_re_reg/P0001  ;
  assign n8599 = \u10_rp_reg[1]/P0001  & n8597 ;
  assign n8598 = ~\u10_rp_reg[1]/P0001  & ~n8597 ;
  assign n8600 = \u13_icc_r_reg[8]/NET0131  & ~n8598 ;
  assign n8601 = ~n8599 & n8600 ;
  assign n8602 = \u11_rp_reg[0]/P0001  & \u12_i6_re_reg/NET0131  ;
  assign n8604 = \u11_rp_reg[1]/P0001  & n8602 ;
  assign n8603 = ~\u11_rp_reg[1]/P0001  & ~n8602 ;
  assign n8605 = \u13_icc_r_reg[16]/NET0131  & ~n8603 ;
  assign n8606 = ~n8604 & n8605 ;
  assign n8608 = \u9_rp_reg[2]/P0001  & n8594 ;
  assign n8607 = ~\u9_rp_reg[2]/P0001  & ~n8594 ;
  assign n8609 = \u13_icc_r_reg[0]/NET0131  & ~n8607 ;
  assign n8610 = ~n8608 & n8609 ;
  assign n8612 = \u11_rp_reg[2]/P0001  & n8604 ;
  assign n8611 = ~\u11_rp_reg[2]/P0001  & ~n8604 ;
  assign n8613 = \u13_icc_r_reg[16]/NET0131  & ~n8611 ;
  assign n8614 = ~n8612 & n8613 ;
  assign n8616 = \u10_rp_reg[2]/P0001  & n8599 ;
  assign n8615 = ~\u10_rp_reg[2]/P0001  & ~n8599 ;
  assign n8617 = \u13_icc_r_reg[8]/NET0131  & ~n8615 ;
  assign n8618 = ~n8616 & n8617 ;
  assign n8619 = ~\u2_res_cnt_reg[2]/P0001  & ~n6455 ;
  assign n8620 = \u2_sync_resume_reg/NET0131  & ~n6456 ;
  assign n8621 = ~n8619 & n8620 ;
  assign n8622 = ~\u11_rp_reg[0]/P0001  & ~\u12_i6_re_reg/NET0131  ;
  assign n8623 = \u13_icc_r_reg[16]/NET0131  & ~n8602 ;
  assign n8624 = ~n8622 & n8623 ;
  assign n8625 = \u13_crac_r_reg[0]/NET0131  & n6159 ;
  assign n8626 = \u13_intm_r_reg[16]/NET0131  & n6153 ;
  assign n8630 = ~n8625 & ~n8626 ;
  assign n8629 = \u13_ints_r_reg[16]/NET0131  & n2741 ;
  assign n8627 = \u13_icc_r_reg[16]/NET0131  & n6157 ;
  assign n8628 = \u13_occ0_r_reg[16]/NET0131  & n6151 ;
  assign n8631 = ~n8627 & ~n8628 ;
  assign n8632 = ~n8629 & n8631 ;
  assign n8633 = n8630 & n8632 ;
  assign n8634 = n6146 & ~n8633 ;
  assign n8637 = \u11_dout_reg[16]/P0001  & n6145 ;
  assign n8635 = \u9_dout_reg[16]/P0001  & n6168 ;
  assign n8636 = \u10_dout_reg[16]/P0001  & n6170 ;
  assign n8638 = ~n8635 & ~n8636 ;
  assign n8639 = ~n8637 & n8638 ;
  assign n8640 = ~n8634 & n8639 ;
  assign n8641 = \u13_icc_r_reg[17]/NET0131  & n6157 ;
  assign n8642 = \u13_intm_r_reg[17]/NET0131  & n6153 ;
  assign n8646 = ~n8641 & ~n8642 ;
  assign n8645 = \u13_ints_r_reg[17]/NET0131  & n2741 ;
  assign n8643 = \u13_crac_r_reg[1]/NET0131  & n6159 ;
  assign n8644 = \u13_occ0_r_reg[17]/NET0131  & n6151 ;
  assign n8647 = ~n8643 & ~n8644 ;
  assign n8648 = ~n8645 & n8647 ;
  assign n8649 = n8646 & n8648 ;
  assign n8650 = n6146 & ~n8649 ;
  assign n8653 = \u11_dout_reg[17]/P0001  & n6145 ;
  assign n8651 = \u9_dout_reg[17]/P0001  & n6168 ;
  assign n8652 = \u10_dout_reg[17]/P0001  & n6170 ;
  assign n8654 = ~n8651 & ~n8652 ;
  assign n8655 = ~n8653 & n8654 ;
  assign n8656 = ~n8650 & n8655 ;
  assign n8657 = \u13_crac_r_reg[3]/NET0131  & n6159 ;
  assign n8658 = \u13_intm_r_reg[19]/NET0131  & n6153 ;
  assign n8662 = ~n8657 & ~n8658 ;
  assign n8661 = \u13_ints_r_reg[19]/NET0131  & n2741 ;
  assign n8659 = \u13_icc_r_reg[19]/NET0131  & n6157 ;
  assign n8660 = \u13_occ0_r_reg[19]/NET0131  & n6151 ;
  assign n8663 = ~n8659 & ~n8660 ;
  assign n8664 = ~n8661 & n8663 ;
  assign n8665 = n8662 & n8664 ;
  assign n8666 = n6146 & ~n8665 ;
  assign n8669 = \u11_dout_reg[19]/P0001  & n6145 ;
  assign n8667 = \u9_dout_reg[19]/P0001  & n6168 ;
  assign n8668 = \u10_dout_reg[19]/P0001  & n6170 ;
  assign n8670 = ~n8667 & ~n8668 ;
  assign n8671 = ~n8669 & n8670 ;
  assign n8672 = ~n8666 & n8671 ;
  assign n8673 = ~\u12_i3_re_reg/NET0131  & ~\u9_rp_reg[0]/P0001  ;
  assign n8674 = \u13_icc_r_reg[0]/NET0131  & ~n8592 ;
  assign n8675 = ~n8673 & n8674 ;
  assign n8676 = \u13_icc_r_reg[20]/NET0131  & n6157 ;
  assign n8677 = \u13_intm_r_reg[20]/NET0131  & n6153 ;
  assign n8681 = ~n8676 & ~n8677 ;
  assign n8680 = \u13_ints_r_reg[20]/NET0131  & n2741 ;
  assign n8678 = \u13_crac_r_reg[4]/NET0131  & n6159 ;
  assign n8679 = \u13_occ0_r_reg[20]/NET0131  & n6151 ;
  assign n8682 = ~n8678 & ~n8679 ;
  assign n8683 = ~n8680 & n8682 ;
  assign n8684 = n8681 & n8683 ;
  assign n8685 = n6146 & ~n8684 ;
  assign n8688 = \u11_dout_reg[20]/P0001  & n6145 ;
  assign n8686 = \u9_dout_reg[20]/P0001  & n6168 ;
  assign n8687 = \u10_dout_reg[20]/P0001  & n6170 ;
  assign n8689 = ~n8686 & ~n8687 ;
  assign n8690 = ~n8688 & n8689 ;
  assign n8691 = ~n8685 & n8690 ;
  assign n8692 = \u13_icc_r_reg[21]/NET0131  & n6157 ;
  assign n8693 = \u13_intm_r_reg[21]/NET0131  & n6153 ;
  assign n8697 = ~n8692 & ~n8693 ;
  assign n8696 = \u13_ints_r_reg[21]/NET0131  & n2741 ;
  assign n8694 = \u13_crac_r_reg[5]/NET0131  & n6159 ;
  assign n8695 = \u13_occ0_r_reg[21]/NET0131  & n6151 ;
  assign n8698 = ~n8694 & ~n8695 ;
  assign n8699 = ~n8696 & n8698 ;
  assign n8700 = n8697 & n8699 ;
  assign n8701 = n6146 & ~n8700 ;
  assign n8704 = \u11_dout_reg[21]/P0001  & n6145 ;
  assign n8702 = \u9_dout_reg[21]/P0001  & n6168 ;
  assign n8703 = \u10_dout_reg[21]/P0001  & n6170 ;
  assign n8705 = ~n8702 & ~n8703 ;
  assign n8706 = ~n8704 & n8705 ;
  assign n8707 = ~n8701 & n8706 ;
  assign n8708 = \u13_icc_r_reg[22]/NET0131  & n6157 ;
  assign n8709 = \u13_intm_r_reg[22]/NET0131  & n6153 ;
  assign n8713 = ~n8708 & ~n8709 ;
  assign n8712 = \u13_ints_r_reg[22]/NET0131  & n2741 ;
  assign n8710 = \u13_crac_r_reg[6]/NET0131  & n6159 ;
  assign n8711 = \u13_occ0_r_reg[22]/NET0131  & n6151 ;
  assign n8714 = ~n8710 & ~n8711 ;
  assign n8715 = ~n8712 & n8714 ;
  assign n8716 = n8713 & n8715 ;
  assign n8717 = n6146 & ~n8716 ;
  assign n8720 = \u11_dout_reg[22]/P0001  & n6145 ;
  assign n8718 = \u9_dout_reg[22]/P0001  & n6168 ;
  assign n8719 = \u10_dout_reg[22]/P0001  & n6170 ;
  assign n8721 = ~n8718 & ~n8719 ;
  assign n8722 = ~n8720 & n8721 ;
  assign n8723 = ~n8717 & n8722 ;
  assign n8724 = \u13_ints_r_reg[23]/NET0131  & n2741 ;
  assign n8725 = \u13_intm_r_reg[23]/NET0131  & n6153 ;
  assign n8728 = ~n8724 & ~n8725 ;
  assign n8726 = \u13_occ0_r_reg[23]/NET0131  & n6151 ;
  assign n8727 = \u13_icc_r_reg[23]/NET0131  & n6157 ;
  assign n8729 = ~n8726 & ~n8727 ;
  assign n8730 = n8728 & n8729 ;
  assign n8731 = n6146 & ~n8730 ;
  assign n8734 = \u10_dout_reg[23]/P0001  & n6170 ;
  assign n8732 = \u9_dout_reg[23]/P0001  & n6168 ;
  assign n8733 = \u11_dout_reg[23]/P0001  & n6145 ;
  assign n8735 = ~n8732 & ~n8733 ;
  assign n8736 = ~n8734 & n8735 ;
  assign n8737 = ~n8731 & n8736 ;
  assign n8738 = ~\u10_rp_reg[0]/P0001  & ~\u12_i4_re_reg/P0001  ;
  assign n8739 = \u13_icc_r_reg[8]/NET0131  & ~n8597 ;
  assign n8740 = ~n8738 & n8739 ;
  assign n8741 = \u13_crac_r_reg[2]/NET0131  & n6159 ;
  assign n8742 = \u13_intm_r_reg[18]/NET0131  & n6153 ;
  assign n8746 = ~n8741 & ~n8742 ;
  assign n8745 = \u13_ints_r_reg[18]/NET0131  & n2741 ;
  assign n8743 = \u13_icc_r_reg[18]/NET0131  & n6157 ;
  assign n8744 = \u13_occ0_r_reg[18]/NET0131  & n6151 ;
  assign n8747 = ~n8743 & ~n8744 ;
  assign n8748 = ~n8745 & n8747 ;
  assign n8749 = n8746 & n8748 ;
  assign n8750 = n6146 & ~n8749 ;
  assign n8753 = \u11_dout_reg[18]/P0001  & n6145 ;
  assign n8751 = \u9_dout_reg[18]/P0001  & n6168 ;
  assign n8752 = \u10_dout_reg[18]/P0001  & n6170 ;
  assign n8754 = ~n8751 & ~n8752 ;
  assign n8755 = ~n8753 & n8754 ;
  assign n8756 = ~n8750 & n8755 ;
  assign n8758 = ~\u2_to_cnt_reg[4]/NET0131  & ~n6481 ;
  assign n8757 = \u2_to_cnt_reg[4]/NET0131  & n6481 ;
  assign n8759 = ~\u2_bit_clk_e_reg/P0001  & ~n8757 ;
  assign n8760 = ~n8758 & n8759 ;
  assign n8762 = \u2_to_cnt_reg[5]/NET0131  & n8757 ;
  assign n8761 = ~\u2_to_cnt_reg[5]/NET0131  & ~n8757 ;
  assign n8763 = ~\u2_bit_clk_e_reg/P0001  & ~n8761 ;
  assign n8764 = ~n8762 & n8763 ;
  assign n8765 = ~\u2_to_cnt_reg[2]/NET0131  & ~n6479 ;
  assign n8766 = ~\u2_bit_clk_e_reg/P0001  & ~n6480 ;
  assign n8767 = ~n8765 & n8766 ;
  assign n8768 = \u12_i3_re_reg/NET0131  & \u9_empty_reg/P0001  ;
  assign n8769 = ~\u23_int_set_reg[1]/NET0131  & ~n8768 ;
  assign n8770 = \u10_empty_reg/P0001  & \u12_i4_re_reg/P0001  ;
  assign n8771 = ~\u24_int_set_reg[1]/NET0131  & ~n8770 ;
  assign n8772 = \u11_empty_reg/P0001  & \u12_i6_re_reg/NET0131  ;
  assign n8773 = ~\u25_int_set_reg[1]/NET0131  & ~n8772 ;
  assign n8774 = ~\u2_res_cnt_reg[0]/P0001  & ~n5629 ;
  assign n8775 = \u2_sync_resume_reg/NET0131  & ~n6454 ;
  assign n8776 = ~n8774 & n8775 ;
  assign n8777 = wb_we_i_pad & n2735 ;
  assign n8778 = \u12_we1_reg/P0001  & n8777 ;
  assign n8779 = ~\u12_we2_reg/P0001  & n8778 ;
  assign n8780 = n6139 & n8779 ;
  assign n8781 = n6143 & n8780 ;
  assign n8782 = n6151 & n8780 ;
  assign n8783 = n6147 & n8780 ;
  assign n8784 = n6159 & n8780 ;
  assign n8785 = n6153 & n8780 ;
  assign n8788 = \u13_ints_r_reg[24]/NET0131  & n2741 ;
  assign n8786 = \u13_occ0_r_reg[24]/NET0131  & n6151 ;
  assign n8787 = \u13_intm_r_reg[24]/NET0131  & n6153 ;
  assign n8789 = ~n8786 & ~n8787 ;
  assign n8790 = ~n8788 & n8789 ;
  assign n8791 = n6146 & ~n8790 ;
  assign n8794 = \u10_dout_reg[24]/P0001  & n6170 ;
  assign n8792 = \u9_dout_reg[24]/P0001  & n6168 ;
  assign n8793 = \u11_dout_reg[24]/P0001  & n6145 ;
  assign n8795 = ~n8792 & ~n8793 ;
  assign n8796 = ~n8794 & n8795 ;
  assign n8797 = ~n8791 & n8796 ;
  assign n8800 = \u13_ints_r_reg[25]/NET0131  & n2741 ;
  assign n8798 = \u13_occ0_r_reg[25]/NET0131  & n6151 ;
  assign n8799 = \u13_intm_r_reg[25]/NET0131  & n6153 ;
  assign n8801 = ~n8798 & ~n8799 ;
  assign n8802 = ~n8800 & n8801 ;
  assign n8803 = n6146 & ~n8802 ;
  assign n8806 = \u10_dout_reg[25]/P0001  & n6170 ;
  assign n8804 = \u9_dout_reg[25]/P0001  & n6168 ;
  assign n8805 = \u11_dout_reg[25]/P0001  & n6145 ;
  assign n8807 = ~n8804 & ~n8805 ;
  assign n8808 = ~n8806 & n8807 ;
  assign n8809 = ~n8803 & n8808 ;
  assign n8812 = \u13_ints_r_reg[26]/NET0131  & n2741 ;
  assign n8810 = \u13_occ0_r_reg[26]/NET0131  & n6151 ;
  assign n8811 = \u13_intm_r_reg[26]/NET0131  & n6153 ;
  assign n8813 = ~n8810 & ~n8811 ;
  assign n8814 = ~n8812 & n8813 ;
  assign n8815 = n6146 & ~n8814 ;
  assign n8818 = \u10_dout_reg[26]/P0001  & n6170 ;
  assign n8816 = \u9_dout_reg[26]/P0001  & n6168 ;
  assign n8817 = \u11_dout_reg[26]/P0001  & n6145 ;
  assign n8819 = ~n8816 & ~n8817 ;
  assign n8820 = ~n8818 & n8819 ;
  assign n8821 = ~n8815 & n8820 ;
  assign n8824 = \u13_ints_r_reg[27]/NET0131  & n2741 ;
  assign n8822 = \u13_occ0_r_reg[27]/NET0131  & n6151 ;
  assign n8823 = \u13_intm_r_reg[27]/NET0131  & n6153 ;
  assign n8825 = ~n8822 & ~n8823 ;
  assign n8826 = ~n8824 & n8825 ;
  assign n8827 = n6146 & ~n8826 ;
  assign n8830 = \u10_dout_reg[27]/P0001  & n6170 ;
  assign n8828 = \u9_dout_reg[27]/P0001  & n6168 ;
  assign n8829 = \u11_dout_reg[27]/P0001  & n6145 ;
  assign n8831 = ~n8828 & ~n8829 ;
  assign n8832 = ~n8830 & n8831 ;
  assign n8833 = ~n8827 & n8832 ;
  assign n8836 = \u13_ints_r_reg[28]/NET0131  & n2741 ;
  assign n8834 = \u13_occ0_r_reg[28]/NET0131  & n6151 ;
  assign n8835 = \u13_intm_r_reg[28]/NET0131  & n6153 ;
  assign n8837 = ~n8834 & ~n8835 ;
  assign n8838 = ~n8836 & n8837 ;
  assign n8839 = n6146 & ~n8838 ;
  assign n8842 = \u10_dout_reg[28]/P0001  & n6170 ;
  assign n8840 = \u9_dout_reg[28]/P0001  & n6168 ;
  assign n8841 = \u11_dout_reg[28]/P0001  & n6145 ;
  assign n8843 = ~n8840 & ~n8841 ;
  assign n8844 = ~n8842 & n8843 ;
  assign n8845 = ~n8839 & n8844 ;
  assign n8846 = \u13_occ0_r_reg[29]/NET0131  & n6151 ;
  assign n8847 = \u11_dout_reg[29]/P0001  & n6145 ;
  assign n8850 = ~n8846 & ~n8847 ;
  assign n8848 = \u9_dout_reg[29]/P0001  & n6168 ;
  assign n8849 = \u10_dout_reg[29]/P0001  & n6170 ;
  assign n8851 = ~n8848 & ~n8849 ;
  assign n8852 = n8850 & n8851 ;
  assign n8853 = \u13_occ0_r_reg[30]/NET0131  & n6151 ;
  assign n8854 = \u11_dout_reg[30]/P0001  & n6145 ;
  assign n8857 = ~n8853 & ~n8854 ;
  assign n8855 = \u9_dout_reg[30]/P0001  & n6168 ;
  assign n8856 = \u10_dout_reg[30]/P0001  & n6170 ;
  assign n8858 = ~n8855 & ~n8856 ;
  assign n8859 = n8857 & n8858 ;
  assign n8862 = \u10_dout_reg[31]/P0001  & n6170 ;
  assign n8860 = \u13_crac_r_reg[7]/NET0131  & n6159 ;
  assign n8861 = \u13_occ0_r_reg[31]/NET0131  & n6151 ;
  assign n8865 = ~n8860 & ~n8861 ;
  assign n8866 = ~n8862 & n8865 ;
  assign n8863 = \u11_dout_reg[31]/P0001  & n6145 ;
  assign n8864 = \u9_dout_reg[31]/P0001  & n6168 ;
  assign n8867 = ~n8863 & ~n8864 ;
  assign n8868 = n8866 & n8867 ;
  assign n8869 = ~\u2_res_cnt_reg[1]/P0001  & ~n6454 ;
  assign n8870 = \u2_sync_resume_reg/NET0131  & ~n6455 ;
  assign n8871 = ~n8869 & n8870 ;
  assign n8872 = ~\u2_cnt_reg[3]/NET0131  & ~n6470 ;
  assign n8873 = ~n6471 & ~n8872 ;
  assign n8874 = ~suspended_o_pad & ~n8873 ;
  assign n8893 = \u13_intm_r_reg[9]/NET0131  & \u13_ints_r_reg[9]/NET0131  ;
  assign n8894 = \u13_intm_r_reg[10]/NET0131  & \u13_ints_r_reg[10]/NET0131  ;
  assign n8913 = ~n8893 & ~n8894 ;
  assign n8895 = \u13_intm_r_reg[4]/NET0131  & \u13_ints_r_reg[4]/NET0131  ;
  assign n8896 = \u13_intm_r_reg[21]/NET0131  & \u13_ints_r_reg[21]/NET0131  ;
  assign n8914 = ~n8895 & ~n8896 ;
  assign n8920 = n8913 & n8914 ;
  assign n8889 = \u13_intm_r_reg[22]/NET0131  & \u13_ints_r_reg[22]/NET0131  ;
  assign n8890 = \u13_intm_r_reg[12]/NET0131  & \u13_ints_r_reg[12]/NET0131  ;
  assign n8911 = ~n8889 & ~n8890 ;
  assign n8891 = \u13_intm_r_reg[19]/NET0131  & \u13_ints_r_reg[19]/NET0131  ;
  assign n8892 = \u13_intm_r_reg[27]/NET0131  & \u13_ints_r_reg[27]/NET0131  ;
  assign n8912 = ~n8891 & ~n8892 ;
  assign n8921 = n8911 & n8912 ;
  assign n8927 = n8920 & n8921 ;
  assign n8903 = \u13_intm_r_reg[3]/NET0131  & \u13_ints_r_reg[3]/NET0131  ;
  assign n8901 = \u13_intm_r_reg[25]/NET0131  & \u13_ints_r_reg[25]/NET0131  ;
  assign n8902 = \u13_intm_r_reg[18]/NET0131  & \u13_ints_r_reg[18]/NET0131  ;
  assign n8917 = ~n8901 & ~n8902 ;
  assign n8918 = ~n8903 & n8917 ;
  assign n8897 = \u13_intm_r_reg[17]/NET0131  & \u13_ints_r_reg[17]/NET0131  ;
  assign n8898 = \u13_intm_r_reg[16]/NET0131  & \u13_ints_r_reg[16]/NET0131  ;
  assign n8915 = ~n8897 & ~n8898 ;
  assign n8899 = \u13_intm_r_reg[20]/NET0131  & \u13_ints_r_reg[20]/NET0131  ;
  assign n8900 = \u13_intm_r_reg[2]/NET0131  & \u13_ints_r_reg[2]/NET0131  ;
  assign n8916 = ~n8899 & ~n8900 ;
  assign n8919 = n8915 & n8916 ;
  assign n8928 = n8918 & n8919 ;
  assign n8929 = n8927 & n8928 ;
  assign n8875 = \u13_intm_r_reg[26]/NET0131  & \u13_ints_r_reg[26]/NET0131  ;
  assign n8876 = \u13_intm_r_reg[15]/NET0131  & \u13_ints_r_reg[15]/NET0131  ;
  assign n8904 = ~n8875 & ~n8876 ;
  assign n8877 = \u13_intm_r_reg[0]/NET0131  & \u13_ints_r_reg[0]/NET0131  ;
  assign n8878 = \u13_intm_r_reg[28]/NET0131  & \u13_ints_r_reg[28]/NET0131  ;
  assign n8905 = ~n8877 & ~n8878 ;
  assign n8879 = \u13_intm_r_reg[1]/NET0131  & \u13_ints_r_reg[1]/NET0131  ;
  assign n8880 = \u13_intm_r_reg[13]/NET0131  & \u13_ints_r_reg[13]/NET0131  ;
  assign n8906 = ~n8879 & ~n8880 ;
  assign n8924 = n8905 & n8906 ;
  assign n8925 = n8904 & n8924 ;
  assign n8885 = \u13_intm_r_reg[7]/NET0131  & \u13_ints_r_reg[7]/NET0131  ;
  assign n8886 = \u13_intm_r_reg[23]/NET0131  & \u13_ints_r_reg[23]/NET0131  ;
  assign n8909 = ~n8885 & ~n8886 ;
  assign n8887 = \u13_intm_r_reg[24]/NET0131  & \u13_ints_r_reg[24]/NET0131  ;
  assign n8888 = \u13_intm_r_reg[14]/NET0131  & \u13_ints_r_reg[14]/NET0131  ;
  assign n8910 = ~n8887 & ~n8888 ;
  assign n8922 = n8909 & n8910 ;
  assign n8881 = \u13_intm_r_reg[11]/NET0131  & \u13_ints_r_reg[11]/NET0131  ;
  assign n8882 = \u13_intm_r_reg[6]/NET0131  & \u13_ints_r_reg[6]/NET0131  ;
  assign n8907 = ~n8881 & ~n8882 ;
  assign n8883 = \u13_intm_r_reg[5]/NET0131  & \u13_ints_r_reg[5]/NET0131  ;
  assign n8884 = \u13_intm_r_reg[8]/NET0131  & \u13_ints_r_reg[8]/NET0131  ;
  assign n8908 = ~n8883 & ~n8884 ;
  assign n8923 = n8907 & n8908 ;
  assign n8926 = n8922 & n8923 ;
  assign n8930 = n8925 & n8926 ;
  assign n8931 = n8929 & n8930 ;
  assign n8932 = n6157 & n8780 ;
  assign n8933 = ~n2738 & ~n8779 ;
  assign n8934 = ~wb_ack_o_pad & wb_cyc_i_pad ;
  assign n8935 = ~n8933 & n8934 ;
  assign n8936 = ~n6287 & ~n6292 ;
  assign n8937 = ~n8579 & ~n8936 ;
  assign n8938 = n6225 & ~n6228 ;
  assign n8939 = ~n6229 & ~n8938 ;
  assign n8940 = n6236 & ~n6239 ;
  assign n8941 = ~n6240 & ~n8940 ;
  assign n8942 = n6249 & ~n6252 ;
  assign n8943 = ~n6253 & ~n8942 ;
  assign n8944 = ~n6261 & ~n6266 ;
  assign n8945 = ~n8537 & ~n8944 ;
  assign n8946 = n6277 & ~n6280 ;
  assign n8947 = ~n6281 & ~n8946 ;
  assign n8948 = n2739 & n8779 ;
  assign n8949 = \u2_ld_reg/P0001  & \u8_dout_reg[0]/P0001  ;
  assign n8950 = \u11_rp_reg[0]/P0001  & ~\u11_wp_reg[1]/P0001  ;
  assign n8951 = \u11_rp_reg[1]/P0001  & ~\u11_wp_reg[2]/P0001  ;
  assign n8952 = ~\u11_rp_reg[1]/P0001  & \u11_wp_reg[2]/P0001  ;
  assign n8953 = ~n8951 & ~n8952 ;
  assign n8954 = n8950 & n8953 ;
  assign n8955 = ~n8950 & ~n8953 ;
  assign n8956 = ~n8954 & ~n8955 ;
  assign n8957 = \u9_rp_reg[0]/P0001  & ~\u9_wp_reg[1]/P0001  ;
  assign n8958 = \u9_rp_reg[1]/P0001  & ~\u9_wp_reg[2]/P0001  ;
  assign n8959 = ~\u9_rp_reg[1]/P0001  & \u9_wp_reg[2]/P0001  ;
  assign n8960 = ~n8958 & ~n8959 ;
  assign n8961 = n8957 & n8960 ;
  assign n8962 = ~n8957 & ~n8960 ;
  assign n8963 = ~n8961 & ~n8962 ;
  assign n8964 = \u10_rp_reg[0]/P0001  & ~\u10_wp_reg[1]/P0001  ;
  assign n8965 = \u10_rp_reg[1]/P0001  & ~\u10_wp_reg[2]/P0001  ;
  assign n8966 = ~\u10_rp_reg[1]/P0001  & \u10_wp_reg[2]/P0001  ;
  assign n8967 = ~n8965 & ~n8966 ;
  assign n8968 = n8964 & n8967 ;
  assign n8969 = ~n8964 & ~n8967 ;
  assign n8970 = ~n8968 & ~n8969 ;
  assign n8971 = ~\u13_ints_r_reg[0]/NET0131  & ~\u15_crac_rd_done_reg/P0001  ;
  assign n8972 = ~n2743 & ~n8971 ;
  assign n8973 = ~\u13_ints_r_reg[10]/NET0131  & ~\u19_int_set_reg[2]/NET0131  ;
  assign n8974 = ~n2743 & ~n8973 ;
  assign n8975 = ~\u13_ints_r_reg[12]/NET0131  & ~\u20_int_set_reg[1]/NET0131  ;
  assign n8976 = ~n2743 & ~n8975 ;
  assign n8977 = ~\u13_ints_r_reg[13]/NET0131  & ~\u20_int_set_reg[2]/NET0131  ;
  assign n8978 = ~n2743 & ~n8977 ;
  assign n8979 = ~\u13_ints_r_reg[15]/NET0131  & ~\u21_int_set_reg[1]/NET0131  ;
  assign n8980 = ~n2743 & ~n8979 ;
  assign n8981 = ~\u13_ints_r_reg[16]/NET0131  & ~\u21_int_set_reg[2]/NET0131  ;
  assign n8982 = ~n2743 & ~n8981 ;
  assign n8983 = ~\u13_ints_r_reg[18]/NET0131  & ~\u22_int_set_reg[1]/NET0131  ;
  assign n8984 = ~n2743 & ~n8983 ;
  assign n8985 = ~\u13_ints_r_reg[19]/NET0131  & ~\u22_int_set_reg[2]/NET0131  ;
  assign n8986 = ~n2743 & ~n8985 ;
  assign n8987 = ~\u13_ints_r_reg[21]/NET0131  & ~\u23_int_set_reg[1]/NET0131  ;
  assign n8988 = ~n2743 & ~n8987 ;
  assign n8989 = ~\u13_ints_r_reg[22]/NET0131  & ~\u23_int_set_reg[2]/NET0131  ;
  assign n8990 = ~n2743 & ~n8989 ;
  assign n8991 = ~\u13_ints_r_reg[24]/NET0131  & ~\u24_int_set_reg[1]/NET0131  ;
  assign n8992 = ~n2743 & ~n8991 ;
  assign n8993 = ~\u13_ints_r_reg[25]/NET0131  & ~\u24_int_set_reg[2]/NET0131  ;
  assign n8994 = ~n2743 & ~n8993 ;
  assign n8995 = ~\u13_ints_r_reg[27]/NET0131  & ~\u25_int_set_reg[1]/NET0131  ;
  assign n8996 = ~n2743 & ~n8995 ;
  assign n8997 = ~\u13_ints_r_reg[28]/NET0131  & ~\u25_int_set_reg[2]/NET0131  ;
  assign n8998 = ~n2743 & ~n8997 ;
  assign n8999 = ~\u13_ints_r_reg[3]/NET0131  & ~\u17_int_set_reg[1]/NET0131  ;
  assign n9000 = ~n2743 & ~n8999 ;
  assign n9001 = ~\u13_ints_r_reg[4]/NET0131  & ~\u17_int_set_reg[2]/NET0131  ;
  assign n9002 = ~n2743 & ~n9001 ;
  assign n9003 = ~\u13_ints_r_reg[6]/NET0131  & ~\u18_int_set_reg[1]/NET0131  ;
  assign n9004 = ~n2743 & ~n9003 ;
  assign n9005 = ~\u13_ints_r_reg[7]/NET0131  & ~\u18_int_set_reg[2]/NET0131  ;
  assign n9006 = ~n2743 & ~n9005 ;
  assign n9007 = ~\u13_ints_r_reg[9]/NET0131  & ~\u19_int_set_reg[1]/NET0131  ;
  assign n9008 = ~n2743 & ~n9007 ;
  assign n9012 = ~\u9_rp_reg[0]/P0001  & \u9_wp_reg[1]/P0001  ;
  assign n9013 = ~n8957 & ~n9012 ;
  assign n9014 = n8960 & n9013 ;
  assign n9009 = ~\u9_rp_reg[2]/P0001  & ~\u9_wp_reg[3]/P0001  ;
  assign n9010 = \u9_rp_reg[2]/P0001  & \u9_wp_reg[3]/P0001  ;
  assign n9011 = ~n9009 & ~n9010 ;
  assign n9015 = n3312 & ~n9011 ;
  assign n9016 = n9014 & n9015 ;
  assign n9017 = ~\wb_addr_i[29]_pad  & ~\wb_addr_i[30]_pad  ;
  assign n9018 = ~\wb_addr_i[31]_pad  & n9017 ;
  assign n9019 = n8777 & n9018 ;
  assign n9020 = ~n8779 & n9019 ;
  assign n9021 = \u2_cnt_reg[0]/NET0131  & ~\u2_cnt_reg[4]/NET0131  ;
  assign n9022 = ~\u2_cnt_reg[1]/NET0131  & \u2_cnt_reg[6]/NET0131  ;
  assign n9023 = n9021 & n9022 ;
  assign n9024 = ~\u2_cnt_reg[2]/NET0131  & ~\u2_cnt_reg[3]/NET0131  ;
  assign n9025 = \u2_cnt_reg[5]/NET0131  & ~\u2_cnt_reg[7]/NET0131  ;
  assign n9026 = n9024 & n9025 ;
  assign n9027 = n9023 & n9026 ;
  assign n9031 = ~\u10_rp_reg[0]/P0001  & \u10_wp_reg[1]/P0001  ;
  assign n9032 = ~n8964 & ~n9031 ;
  assign n9033 = n8967 & n9032 ;
  assign n9028 = ~\u10_rp_reg[2]/P0001  & ~\u10_wp_reg[3]/P0001  ;
  assign n9029 = \u10_rp_reg[2]/P0001  & \u10_wp_reg[3]/P0001  ;
  assign n9030 = ~n9028 & ~n9029 ;
  assign n9034 = n3502 & ~n9030 ;
  assign n9035 = n9033 & n9034 ;
  assign n9039 = ~\u11_rp_reg[0]/P0001  & \u11_wp_reg[1]/P0001  ;
  assign n9040 = ~n8950 & ~n9039 ;
  assign n9041 = n8953 & n9040 ;
  assign n9036 = ~\u11_rp_reg[2]/P0001  & ~\u11_wp_reg[3]/P0001  ;
  assign n9037 = \u11_rp_reg[2]/P0001  & \u11_wp_reg[3]/P0001  ;
  assign n9038 = ~n9036 & ~n9037 ;
  assign n9042 = n3065 & ~n9038 ;
  assign n9043 = n9041 & n9042 ;
  assign n9044 = ~\u2_cnt_reg[5]/NET0131  & ~n6472 ;
  assign n9045 = \u2_cnt_reg[5]/NET0131  & n6472 ;
  assign n9046 = ~n9044 & ~n9045 ;
  assign n9047 = ~suspended_o_pad & ~n9046 ;
  assign n9048 = ~\u2_cnt_reg[6]/NET0131  & ~n9045 ;
  assign n9049 = ~n6474 & ~n9048 ;
  assign n9050 = ~suspended_o_pad & ~n9049 ;
  assign n9054 = ~\u2_cnt_reg[4]/NET0131  & ~\u2_cnt_reg[5]/NET0131  ;
  assign n9055 = ~\u2_cnt_reg[6]/NET0131  & n9054 ;
  assign n9051 = ~\u2_cnt_reg[1]/NET0131  & ~\u2_cnt_reg[2]/NET0131  ;
  assign n9052 = \u2_cnt_reg[0]/NET0131  & \u2_cnt_reg[3]/NET0131  ;
  assign n9053 = n9051 & n9052 ;
  assign n9056 = \u2_cnt_reg[7]/NET0131  & n9053 ;
  assign n9057 = n9055 & n9056 ;
  assign n9058 = ~\u2_cnt_reg[6]/NET0131  & ~\u2_cnt_reg[7]/NET0131  ;
  assign n9059 = n9054 & n9058 ;
  assign n9060 = ~\u2_to_cnt_reg[2]/NET0131  & ~\u2_to_cnt_reg[3]/NET0131  ;
  assign n9061 = ~\u2_to_cnt_reg[4]/NET0131  & \u2_to_cnt_reg[5]/NET0131  ;
  assign n9062 = n9060 & n9061 ;
  assign n9063 = \u2_to_cnt_reg[0]/NET0131  & ~\u2_to_cnt_reg[1]/NET0131  ;
  assign n9064 = n9062 & n9063 ;
  assign n9065 = \u2_to_cnt_reg[0]/NET0131  & ~n9064 ;
  assign n9066 = ~\u2_bit_clk_e_reg/P0001  & ~n9065 ;
  assign n9067 = \u2_to_cnt_reg[0]/NET0131  & ~n9062 ;
  assign n9068 = ~\u2_to_cnt_reg[1]/NET0131  & ~n9067 ;
  assign n9069 = ~\u2_bit_clk_e_reg/P0001  & ~n6479 ;
  assign n9070 = ~n9068 & n9069 ;
  assign n9071 = n9030 & n9033 ;
  assign n9072 = n9038 & n9041 ;
  assign n9073 = \u2_cnt_reg[2]/NET0131  & \u2_cnt_reg[3]/NET0131  ;
  assign n9074 = ~\u2_cnt_reg[5]/NET0131  & ~\u2_cnt_reg[7]/NET0131  ;
  assign n9075 = n9073 & n9074 ;
  assign n9076 = n9023 & n9075 ;
  assign n9077 = n9011 & n9014 ;
  assign n9078 = ~\u2_cnt_reg[1]/NET0131  & ~\u2_cnt_reg[3]/NET0131  ;
  assign n9079 = ~\u2_cnt_reg[2]/NET0131  & n9078 ;
  assign n9080 = ~\u2_cnt_reg[4]/NET0131  & n9079 ;
  assign n9081 = n6473 & ~n9080 ;
  assign n9082 = ~\u2_cnt_reg[7]/NET0131  & ~n9081 ;
  assign n9083 = n2738 & n6168 ;
  assign n9084 = n2738 & n6170 ;
  assign n9085 = \u2_cnt_reg[3]/NET0131  & ~n9051 ;
  assign n9086 = \u2_cnt_reg[4]/NET0131  & \u2_cnt_reg[5]/NET0131  ;
  assign n9087 = n9085 & n9086 ;
  assign n9088 = n9058 & ~n9087 ;
  assign n9089 = ~suspended_o_pad & \u2_cnt_reg[0]/NET0131  ;
  assign n9090 = ~\u2_cnt_reg[0]/NET0131  & ~\u2_cnt_reg[1]/NET0131  ;
  assign n9091 = ~n6469 & ~n9090 ;
  assign n9092 = ~suspended_o_pad & ~n9091 ;
  assign n9093 = ~\u2_cnt_reg[2]/NET0131  & ~n6469 ;
  assign n9094 = ~n6470 & ~n9093 ;
  assign n9095 = ~suspended_o_pad & ~n9094 ;
  assign n9096 = n9055 & ~n9085 ;
  assign n9097 = \u2_cnt_reg[7]/NET0131  & ~n9096 ;
  assign n9098 = ~\u2_cnt_reg[0]/NET0131  & n9059 ;
  assign n9099 = n9079 & n9098 ;
  assign n9100 = \u2_cnt_reg[2]/NET0131  & \u2_cnt_reg[5]/NET0131  ;
  assign n9101 = n9021 & n9100 ;
  assign n9102 = n9058 & n9078 ;
  assign n9103 = n9101 & n9102 ;
  assign n9104 = n2738 & n6145 ;
  assign n9105 = \u2_cnt_reg[1]/NET0131  & n9073 ;
  assign n9106 = n9054 & ~n9105 ;
  assign n9107 = \u2_cnt_reg[6]/NET0131  & ~n9106 ;
  assign n9108 = ~\u2_cnt_reg[7]/NET0131  & ~n9107 ;
  assign n9109 = \u2_cnt_reg[4]/NET0131  & n9058 ;
  assign n9110 = \u2_cnt_reg[5]/NET0131  & n9053 ;
  assign n9111 = n9109 & n9110 ;
  assign n9112 = \u9_rp_reg[0]/P0001  & ~\u9_rp_reg[1]/P0001  ;
  assign n9113 = \u9_mem_reg[1][0]/P0001  & n9112 ;
  assign n9114 = ~\u9_rp_reg[0]/P0001  & ~\u9_rp_reg[1]/P0001  ;
  assign n9115 = \u9_mem_reg[0][0]/P0001  & n9114 ;
  assign n9120 = ~n9113 & ~n9115 ;
  assign n9116 = \u9_rp_reg[0]/P0001  & \u9_rp_reg[1]/P0001  ;
  assign n9117 = \u9_mem_reg[3][0]/P0001  & n9116 ;
  assign n9118 = ~\u9_rp_reg[0]/P0001  & \u9_rp_reg[1]/P0001  ;
  assign n9119 = \u9_mem_reg[2][0]/P0001  & n9118 ;
  assign n9121 = ~n9117 & ~n9119 ;
  assign n9122 = n9120 & n9121 ;
  assign n9123 = \u9_mem_reg[2][10]/P0001  & n9118 ;
  assign n9124 = \u9_mem_reg[0][10]/P0001  & n9114 ;
  assign n9127 = ~n9123 & ~n9124 ;
  assign n9125 = \u9_mem_reg[3][10]/P0001  & n9116 ;
  assign n9126 = \u9_mem_reg[1][10]/P0001  & n9112 ;
  assign n9128 = ~n9125 & ~n9126 ;
  assign n9129 = n9127 & n9128 ;
  assign n9130 = \u9_mem_reg[1][11]/P0001  & n9112 ;
  assign n9131 = \u9_mem_reg[0][11]/P0001  & n9114 ;
  assign n9134 = ~n9130 & ~n9131 ;
  assign n9132 = \u9_mem_reg[3][11]/P0001  & n9116 ;
  assign n9133 = \u9_mem_reg[2][11]/P0001  & n9118 ;
  assign n9135 = ~n9132 & ~n9133 ;
  assign n9136 = n9134 & n9135 ;
  assign n9137 = \u9_mem_reg[1][12]/P0001  & n9112 ;
  assign n9138 = \u9_mem_reg[0][12]/P0001  & n9114 ;
  assign n9141 = ~n9137 & ~n9138 ;
  assign n9139 = \u9_mem_reg[3][12]/P0001  & n9116 ;
  assign n9140 = \u9_mem_reg[2][12]/P0001  & n9118 ;
  assign n9142 = ~n9139 & ~n9140 ;
  assign n9143 = n9141 & n9142 ;
  assign n9144 = \u9_mem_reg[1][13]/P0001  & n9112 ;
  assign n9145 = \u9_mem_reg[0][13]/P0001  & n9114 ;
  assign n9148 = ~n9144 & ~n9145 ;
  assign n9146 = \u9_mem_reg[3][13]/P0001  & n9116 ;
  assign n9147 = \u9_mem_reg[2][13]/P0001  & n9118 ;
  assign n9149 = ~n9146 & ~n9147 ;
  assign n9150 = n9148 & n9149 ;
  assign n9151 = \u9_mem_reg[1][14]/P0001  & n9112 ;
  assign n9152 = \u9_mem_reg[0][14]/P0001  & n9114 ;
  assign n9155 = ~n9151 & ~n9152 ;
  assign n9153 = \u9_mem_reg[3][14]/P0001  & n9116 ;
  assign n9154 = \u9_mem_reg[2][14]/P0001  & n9118 ;
  assign n9156 = ~n9153 & ~n9154 ;
  assign n9157 = n9155 & n9156 ;
  assign n9158 = \u9_mem_reg[1][15]/P0001  & n9112 ;
  assign n9159 = \u9_mem_reg[0][15]/P0001  & n9114 ;
  assign n9162 = ~n9158 & ~n9159 ;
  assign n9160 = \u9_mem_reg[3][15]/P0001  & n9116 ;
  assign n9161 = \u9_mem_reg[2][15]/P0001  & n9118 ;
  assign n9163 = ~n9160 & ~n9161 ;
  assign n9164 = n9162 & n9163 ;
  assign n9165 = \u9_mem_reg[2][16]/P0001  & n9118 ;
  assign n9166 = \u9_mem_reg[1][16]/P0001  & n9112 ;
  assign n9169 = ~n9165 & ~n9166 ;
  assign n9167 = \u9_mem_reg[3][16]/P0001  & n9116 ;
  assign n9168 = \u9_mem_reg[0][16]/P0001  & n9114 ;
  assign n9170 = ~n9167 & ~n9168 ;
  assign n9171 = n9169 & n9170 ;
  assign n9172 = \u9_mem_reg[1][17]/P0001  & n9112 ;
  assign n9173 = \u9_mem_reg[0][17]/P0001  & n9114 ;
  assign n9176 = ~n9172 & ~n9173 ;
  assign n9174 = \u9_mem_reg[3][17]/P0001  & n9116 ;
  assign n9175 = \u9_mem_reg[2][17]/P0001  & n9118 ;
  assign n9177 = ~n9174 & ~n9175 ;
  assign n9178 = n9176 & n9177 ;
  assign n9179 = \u9_mem_reg[1][18]/P0001  & n9112 ;
  assign n9180 = \u9_mem_reg[2][18]/P0001  & n9118 ;
  assign n9183 = ~n9179 & ~n9180 ;
  assign n9181 = \u9_mem_reg[3][18]/P0001  & n9116 ;
  assign n9182 = \u9_mem_reg[0][18]/P0001  & n9114 ;
  assign n9184 = ~n9181 & ~n9182 ;
  assign n9185 = n9183 & n9184 ;
  assign n9186 = \u9_mem_reg[2][19]/P0001  & n9118 ;
  assign n9187 = \u9_mem_reg[1][19]/P0001  & n9112 ;
  assign n9190 = ~n9186 & ~n9187 ;
  assign n9188 = \u9_mem_reg[3][19]/P0001  & n9116 ;
  assign n9189 = \u9_mem_reg[0][19]/P0001  & n9114 ;
  assign n9191 = ~n9188 & ~n9189 ;
  assign n9192 = n9190 & n9191 ;
  assign n9193 = \u9_mem_reg[1][1]/P0001  & n9112 ;
  assign n9194 = \u9_mem_reg[0][1]/P0001  & n9114 ;
  assign n9197 = ~n9193 & ~n9194 ;
  assign n9195 = \u9_mem_reg[3][1]/P0001  & n9116 ;
  assign n9196 = \u9_mem_reg[2][1]/P0001  & n9118 ;
  assign n9198 = ~n9195 & ~n9196 ;
  assign n9199 = n9197 & n9198 ;
  assign n9200 = \u9_mem_reg[0][20]/P0001  & n9114 ;
  assign n9201 = \u9_mem_reg[2][20]/P0001  & n9118 ;
  assign n9204 = ~n9200 & ~n9201 ;
  assign n9202 = \u9_mem_reg[3][20]/P0001  & n9116 ;
  assign n9203 = \u9_mem_reg[1][20]/P0001  & n9112 ;
  assign n9205 = ~n9202 & ~n9203 ;
  assign n9206 = n9204 & n9205 ;
  assign n9207 = \u9_mem_reg[2][21]/P0001  & n9118 ;
  assign n9208 = \u9_mem_reg[1][21]/P0001  & n9112 ;
  assign n9211 = ~n9207 & ~n9208 ;
  assign n9209 = \u9_mem_reg[3][21]/P0001  & n9116 ;
  assign n9210 = \u9_mem_reg[0][21]/P0001  & n9114 ;
  assign n9212 = ~n9209 & ~n9210 ;
  assign n9213 = n9211 & n9212 ;
  assign n9214 = \u9_mem_reg[2][22]/P0001  & n9118 ;
  assign n9215 = \u9_mem_reg[1][22]/P0001  & n9112 ;
  assign n9218 = ~n9214 & ~n9215 ;
  assign n9216 = \u9_mem_reg[3][22]/P0001  & n9116 ;
  assign n9217 = \u9_mem_reg[0][22]/P0001  & n9114 ;
  assign n9219 = ~n9216 & ~n9217 ;
  assign n9220 = n9218 & n9219 ;
  assign n9221 = \u9_mem_reg[1][23]/P0001  & n9112 ;
  assign n9222 = \u9_mem_reg[2][23]/P0001  & n9118 ;
  assign n9225 = ~n9221 & ~n9222 ;
  assign n9223 = \u9_mem_reg[3][23]/P0001  & n9116 ;
  assign n9224 = \u9_mem_reg[0][23]/P0001  & n9114 ;
  assign n9226 = ~n9223 & ~n9224 ;
  assign n9227 = n9225 & n9226 ;
  assign n9228 = \u9_mem_reg[2][24]/P0001  & n9118 ;
  assign n9229 = \u9_mem_reg[1][24]/P0001  & n9112 ;
  assign n9232 = ~n9228 & ~n9229 ;
  assign n9230 = \u9_mem_reg[3][24]/P0001  & n9116 ;
  assign n9231 = \u9_mem_reg[0][24]/P0001  & n9114 ;
  assign n9233 = ~n9230 & ~n9231 ;
  assign n9234 = n9232 & n9233 ;
  assign n9235 = \u9_mem_reg[2][26]/P0001  & n9118 ;
  assign n9236 = \u9_mem_reg[1][26]/P0001  & n9112 ;
  assign n9239 = ~n9235 & ~n9236 ;
  assign n9237 = \u9_mem_reg[3][26]/P0001  & n9116 ;
  assign n9238 = \u9_mem_reg[0][26]/P0001  & n9114 ;
  assign n9240 = ~n9237 & ~n9238 ;
  assign n9241 = n9239 & n9240 ;
  assign n9242 = \u9_mem_reg[2][27]/P0001  & n9118 ;
  assign n9243 = \u9_mem_reg[1][27]/P0001  & n9112 ;
  assign n9246 = ~n9242 & ~n9243 ;
  assign n9244 = \u9_mem_reg[3][27]/P0001  & n9116 ;
  assign n9245 = \u9_mem_reg[0][27]/P0001  & n9114 ;
  assign n9247 = ~n9244 & ~n9245 ;
  assign n9248 = n9246 & n9247 ;
  assign n9249 = \u9_mem_reg[2][28]/P0001  & n9118 ;
  assign n9250 = \u9_mem_reg[1][28]/P0001  & n9112 ;
  assign n9253 = ~n9249 & ~n9250 ;
  assign n9251 = \u9_mem_reg[3][28]/P0001  & n9116 ;
  assign n9252 = \u9_mem_reg[0][28]/P0001  & n9114 ;
  assign n9254 = ~n9251 & ~n9252 ;
  assign n9255 = n9253 & n9254 ;
  assign n9256 = \u9_mem_reg[1][29]/P0001  & n9112 ;
  assign n9257 = \u9_mem_reg[2][29]/P0001  & n9118 ;
  assign n9260 = ~n9256 & ~n9257 ;
  assign n9258 = \u9_mem_reg[3][29]/P0001  & n9116 ;
  assign n9259 = \u9_mem_reg[0][29]/P0001  & n9114 ;
  assign n9261 = ~n9258 & ~n9259 ;
  assign n9262 = n9260 & n9261 ;
  assign n9263 = \u9_mem_reg[1][2]/P0001  & n9112 ;
  assign n9264 = \u9_mem_reg[0][2]/P0001  & n9114 ;
  assign n9267 = ~n9263 & ~n9264 ;
  assign n9265 = \u9_mem_reg[3][2]/P0001  & n9116 ;
  assign n9266 = \u9_mem_reg[2][2]/P0001  & n9118 ;
  assign n9268 = ~n9265 & ~n9266 ;
  assign n9269 = n9267 & n9268 ;
  assign n9270 = \u9_mem_reg[2][30]/P0001  & n9118 ;
  assign n9271 = \u9_mem_reg[1][30]/P0001  & n9112 ;
  assign n9274 = ~n9270 & ~n9271 ;
  assign n9272 = \u9_mem_reg[3][30]/P0001  & n9116 ;
  assign n9273 = \u9_mem_reg[0][30]/P0001  & n9114 ;
  assign n9275 = ~n9272 & ~n9273 ;
  assign n9276 = n9274 & n9275 ;
  assign n9277 = \u9_mem_reg[2][31]/P0001  & n9118 ;
  assign n9278 = \u9_mem_reg[1][31]/P0001  & n9112 ;
  assign n9281 = ~n9277 & ~n9278 ;
  assign n9279 = \u9_mem_reg[3][31]/P0001  & n9116 ;
  assign n9280 = \u9_mem_reg[0][31]/P0001  & n9114 ;
  assign n9282 = ~n9279 & ~n9280 ;
  assign n9283 = n9281 & n9282 ;
  assign n9284 = \u9_mem_reg[1][3]/P0001  & n9112 ;
  assign n9285 = \u9_mem_reg[0][3]/P0001  & n9114 ;
  assign n9288 = ~n9284 & ~n9285 ;
  assign n9286 = \u9_mem_reg[3][3]/P0001  & n9116 ;
  assign n9287 = \u9_mem_reg[2][3]/P0001  & n9118 ;
  assign n9289 = ~n9286 & ~n9287 ;
  assign n9290 = n9288 & n9289 ;
  assign n9291 = \u9_mem_reg[1][5]/P0001  & n9112 ;
  assign n9292 = \u9_mem_reg[0][5]/P0001  & n9114 ;
  assign n9295 = ~n9291 & ~n9292 ;
  assign n9293 = \u9_mem_reg[3][5]/P0001  & n9116 ;
  assign n9294 = \u9_mem_reg[2][5]/P0001  & n9118 ;
  assign n9296 = ~n9293 & ~n9294 ;
  assign n9297 = n9295 & n9296 ;
  assign n9298 = \u9_mem_reg[2][6]/P0001  & n9118 ;
  assign n9299 = \u9_mem_reg[1][6]/P0001  & n9112 ;
  assign n9302 = ~n9298 & ~n9299 ;
  assign n9300 = \u9_mem_reg[3][6]/P0001  & n9116 ;
  assign n9301 = \u9_mem_reg[0][6]/P0001  & n9114 ;
  assign n9303 = ~n9300 & ~n9301 ;
  assign n9304 = n9302 & n9303 ;
  assign n9305 = \u9_mem_reg[2][7]/P0001  & n9118 ;
  assign n9306 = \u9_mem_reg[0][7]/P0001  & n9114 ;
  assign n9309 = ~n9305 & ~n9306 ;
  assign n9307 = \u9_mem_reg[3][7]/P0001  & n9116 ;
  assign n9308 = \u9_mem_reg[1][7]/P0001  & n9112 ;
  assign n9310 = ~n9307 & ~n9308 ;
  assign n9311 = n9309 & n9310 ;
  assign n9312 = ~\u10_rp_reg[0]/P0001  & \u10_rp_reg[1]/P0001  ;
  assign n9313 = \u10_mem_reg[2][0]/P0001  & n9312 ;
  assign n9314 = ~\u10_rp_reg[0]/P0001  & ~\u10_rp_reg[1]/P0001  ;
  assign n9315 = \u10_mem_reg[0][0]/P0001  & n9314 ;
  assign n9320 = ~n9313 & ~n9315 ;
  assign n9316 = \u10_rp_reg[0]/P0001  & \u10_rp_reg[1]/P0001  ;
  assign n9317 = \u10_mem_reg[3][0]/P0001  & n9316 ;
  assign n9318 = \u10_rp_reg[0]/P0001  & ~\u10_rp_reg[1]/P0001  ;
  assign n9319 = \u10_mem_reg[1][0]/P0001  & n9318 ;
  assign n9321 = ~n9317 & ~n9319 ;
  assign n9322 = n9320 & n9321 ;
  assign n9323 = \u9_mem_reg[1][25]/P0001  & n9112 ;
  assign n9324 = \u9_mem_reg[2][25]/P0001  & n9118 ;
  assign n9327 = ~n9323 & ~n9324 ;
  assign n9325 = \u9_mem_reg[3][25]/P0001  & n9116 ;
  assign n9326 = \u9_mem_reg[0][25]/P0001  & n9114 ;
  assign n9328 = ~n9325 & ~n9326 ;
  assign n9329 = n9327 & n9328 ;
  assign n9330 = \u10_mem_reg[1][11]/P0001  & n9318 ;
  assign n9331 = \u10_mem_reg[0][11]/P0001  & n9314 ;
  assign n9334 = ~n9330 & ~n9331 ;
  assign n9332 = \u10_mem_reg[3][11]/P0001  & n9316 ;
  assign n9333 = \u10_mem_reg[2][11]/P0001  & n9312 ;
  assign n9335 = ~n9332 & ~n9333 ;
  assign n9336 = n9334 & n9335 ;
  assign n9337 = \u10_mem_reg[1][12]/P0001  & n9318 ;
  assign n9338 = \u10_mem_reg[0][12]/P0001  & n9314 ;
  assign n9341 = ~n9337 & ~n9338 ;
  assign n9339 = \u10_mem_reg[3][12]/P0001  & n9316 ;
  assign n9340 = \u10_mem_reg[2][12]/P0001  & n9312 ;
  assign n9342 = ~n9339 & ~n9340 ;
  assign n9343 = n9341 & n9342 ;
  assign n9344 = \u10_mem_reg[2][13]/P0001  & n9312 ;
  assign n9345 = \u10_mem_reg[0][13]/P0001  & n9314 ;
  assign n9348 = ~n9344 & ~n9345 ;
  assign n9346 = \u10_mem_reg[3][13]/P0001  & n9316 ;
  assign n9347 = \u10_mem_reg[1][13]/P0001  & n9318 ;
  assign n9349 = ~n9346 & ~n9347 ;
  assign n9350 = n9348 & n9349 ;
  assign n9351 = \u10_mem_reg[2][15]/P0001  & n9312 ;
  assign n9352 = \u10_mem_reg[0][15]/P0001  & n9314 ;
  assign n9355 = ~n9351 & ~n9352 ;
  assign n9353 = \u10_mem_reg[3][15]/P0001  & n9316 ;
  assign n9354 = \u10_mem_reg[1][15]/P0001  & n9318 ;
  assign n9356 = ~n9353 & ~n9354 ;
  assign n9357 = n9355 & n9356 ;
  assign n9358 = \u10_mem_reg[1][16]/P0001  & n9318 ;
  assign n9359 = \u10_mem_reg[0][16]/P0001  & n9314 ;
  assign n9362 = ~n9358 & ~n9359 ;
  assign n9360 = \u10_mem_reg[3][16]/P0001  & n9316 ;
  assign n9361 = \u10_mem_reg[2][16]/P0001  & n9312 ;
  assign n9363 = ~n9360 & ~n9361 ;
  assign n9364 = n9362 & n9363 ;
  assign n9365 = \u10_mem_reg[2][17]/P0001  & n9312 ;
  assign n9366 = \u10_mem_reg[1][17]/P0001  & n9318 ;
  assign n9369 = ~n9365 & ~n9366 ;
  assign n9367 = \u10_mem_reg[3][17]/P0001  & n9316 ;
  assign n9368 = \u10_mem_reg[0][17]/P0001  & n9314 ;
  assign n9370 = ~n9367 & ~n9368 ;
  assign n9371 = n9369 & n9370 ;
  assign n9372 = \u10_mem_reg[1][18]/P0001  & n9318 ;
  assign n9373 = \u10_mem_reg[2][18]/P0001  & n9312 ;
  assign n9376 = ~n9372 & ~n9373 ;
  assign n9374 = \u10_mem_reg[3][18]/P0001  & n9316 ;
  assign n9375 = \u10_mem_reg[0][18]/P0001  & n9314 ;
  assign n9377 = ~n9374 & ~n9375 ;
  assign n9378 = n9376 & n9377 ;
  assign n9379 = \u10_mem_reg[0][19]/P0001  & n9314 ;
  assign n9380 = \u10_mem_reg[2][19]/P0001  & n9312 ;
  assign n9383 = ~n9379 & ~n9380 ;
  assign n9381 = \u10_mem_reg[3][19]/P0001  & n9316 ;
  assign n9382 = \u10_mem_reg[1][19]/P0001  & n9318 ;
  assign n9384 = ~n9381 & ~n9382 ;
  assign n9385 = n9383 & n9384 ;
  assign n9386 = \u10_mem_reg[2][1]/P0001  & n9312 ;
  assign n9387 = \u10_mem_reg[0][1]/P0001  & n9314 ;
  assign n9390 = ~n9386 & ~n9387 ;
  assign n9388 = \u10_mem_reg[3][1]/P0001  & n9316 ;
  assign n9389 = \u10_mem_reg[1][1]/P0001  & n9318 ;
  assign n9391 = ~n9388 & ~n9389 ;
  assign n9392 = n9390 & n9391 ;
  assign n9393 = \u11_rp_reg[0]/P0001  & ~\u11_rp_reg[1]/P0001  ;
  assign n9394 = \u11_mem_reg[1][6]/P0001  & n9393 ;
  assign n9395 = ~\u11_rp_reg[0]/P0001  & ~\u11_rp_reg[1]/P0001  ;
  assign n9396 = \u11_mem_reg[0][6]/P0001  & n9395 ;
  assign n9401 = ~n9394 & ~n9396 ;
  assign n9397 = \u11_rp_reg[0]/P0001  & \u11_rp_reg[1]/P0001  ;
  assign n9398 = \u11_mem_reg[3][6]/P0001  & n9397 ;
  assign n9399 = ~\u11_rp_reg[0]/P0001  & \u11_rp_reg[1]/P0001  ;
  assign n9400 = \u11_mem_reg[2][6]/P0001  & n9399 ;
  assign n9402 = ~n9398 & ~n9400 ;
  assign n9403 = n9401 & n9402 ;
  assign n9404 = \u10_mem_reg[0][20]/P0001  & n9314 ;
  assign n9405 = \u10_mem_reg[2][20]/P0001  & n9312 ;
  assign n9408 = ~n9404 & ~n9405 ;
  assign n9406 = \u10_mem_reg[3][20]/P0001  & n9316 ;
  assign n9407 = \u10_mem_reg[1][20]/P0001  & n9318 ;
  assign n9409 = ~n9406 & ~n9407 ;
  assign n9410 = n9408 & n9409 ;
  assign n9411 = \u10_mem_reg[0][21]/P0001  & n9314 ;
  assign n9412 = \u10_mem_reg[2][21]/P0001  & n9312 ;
  assign n9415 = ~n9411 & ~n9412 ;
  assign n9413 = \u10_mem_reg[3][21]/P0001  & n9316 ;
  assign n9414 = \u10_mem_reg[1][21]/P0001  & n9318 ;
  assign n9416 = ~n9413 & ~n9414 ;
  assign n9417 = n9415 & n9416 ;
  assign n9418 = \u10_mem_reg[1][22]/P0001  & n9318 ;
  assign n9419 = \u10_mem_reg[2][22]/P0001  & n9312 ;
  assign n9422 = ~n9418 & ~n9419 ;
  assign n9420 = \u10_mem_reg[3][22]/P0001  & n9316 ;
  assign n9421 = \u10_mem_reg[0][22]/P0001  & n9314 ;
  assign n9423 = ~n9420 & ~n9421 ;
  assign n9424 = n9422 & n9423 ;
  assign n9425 = \u10_mem_reg[0][23]/P0001  & n9314 ;
  assign n9426 = \u10_mem_reg[2][23]/P0001  & n9312 ;
  assign n9429 = ~n9425 & ~n9426 ;
  assign n9427 = \u10_mem_reg[3][23]/P0001  & n9316 ;
  assign n9428 = \u10_mem_reg[1][23]/P0001  & n9318 ;
  assign n9430 = ~n9427 & ~n9428 ;
  assign n9431 = n9429 & n9430 ;
  assign n9432 = \u10_mem_reg[2][24]/P0001  & n9312 ;
  assign n9433 = \u10_mem_reg[1][24]/P0001  & n9318 ;
  assign n9436 = ~n9432 & ~n9433 ;
  assign n9434 = \u10_mem_reg[3][24]/P0001  & n9316 ;
  assign n9435 = \u10_mem_reg[0][24]/P0001  & n9314 ;
  assign n9437 = ~n9434 & ~n9435 ;
  assign n9438 = n9436 & n9437 ;
  assign n9439 = \u10_mem_reg[1][25]/P0001  & n9318 ;
  assign n9440 = \u10_mem_reg[2][25]/P0001  & n9312 ;
  assign n9443 = ~n9439 & ~n9440 ;
  assign n9441 = \u10_mem_reg[3][25]/P0001  & n9316 ;
  assign n9442 = \u10_mem_reg[0][25]/P0001  & n9314 ;
  assign n9444 = ~n9441 & ~n9442 ;
  assign n9445 = n9443 & n9444 ;
  assign n9446 = \u10_mem_reg[2][26]/P0001  & n9312 ;
  assign n9447 = \u10_mem_reg[1][26]/P0001  & n9318 ;
  assign n9450 = ~n9446 & ~n9447 ;
  assign n9448 = \u10_mem_reg[3][26]/P0001  & n9316 ;
  assign n9449 = \u10_mem_reg[0][26]/P0001  & n9314 ;
  assign n9451 = ~n9448 & ~n9449 ;
  assign n9452 = n9450 & n9451 ;
  assign n9453 = \u10_mem_reg[0][27]/P0001  & n9314 ;
  assign n9454 = \u10_mem_reg[2][27]/P0001  & n9312 ;
  assign n9457 = ~n9453 & ~n9454 ;
  assign n9455 = \u10_mem_reg[3][27]/P0001  & n9316 ;
  assign n9456 = \u10_mem_reg[1][27]/P0001  & n9318 ;
  assign n9458 = ~n9455 & ~n9456 ;
  assign n9459 = n9457 & n9458 ;
  assign n9460 = \u9_mem_reg[1][4]/P0001  & n9112 ;
  assign n9461 = \u9_mem_reg[0][4]/P0001  & n9114 ;
  assign n9464 = ~n9460 & ~n9461 ;
  assign n9462 = \u9_mem_reg[3][4]/P0001  & n9116 ;
  assign n9463 = \u9_mem_reg[2][4]/P0001  & n9118 ;
  assign n9465 = ~n9462 & ~n9463 ;
  assign n9466 = n9464 & n9465 ;
  assign n9467 = \u10_mem_reg[0][28]/P0001  & n9314 ;
  assign n9468 = \u10_mem_reg[2][28]/P0001  & n9312 ;
  assign n9471 = ~n9467 & ~n9468 ;
  assign n9469 = \u10_mem_reg[3][28]/P0001  & n9316 ;
  assign n9470 = \u10_mem_reg[1][28]/P0001  & n9318 ;
  assign n9472 = ~n9469 & ~n9470 ;
  assign n9473 = n9471 & n9472 ;
  assign n9474 = \u10_mem_reg[2][29]/P0001  & n9312 ;
  assign n9475 = \u10_mem_reg[1][29]/P0001  & n9318 ;
  assign n9478 = ~n9474 & ~n9475 ;
  assign n9476 = \u10_mem_reg[3][29]/P0001  & n9316 ;
  assign n9477 = \u10_mem_reg[0][29]/P0001  & n9314 ;
  assign n9479 = ~n9476 & ~n9477 ;
  assign n9480 = n9478 & n9479 ;
  assign n9481 = \u11_mem_reg[1][0]/P0001  & n9393 ;
  assign n9482 = \u11_mem_reg[0][0]/P0001  & n9395 ;
  assign n9485 = ~n9481 & ~n9482 ;
  assign n9483 = \u11_mem_reg[3][0]/P0001  & n9397 ;
  assign n9484 = \u11_mem_reg[2][0]/P0001  & n9399 ;
  assign n9486 = ~n9483 & ~n9484 ;
  assign n9487 = n9485 & n9486 ;
  assign n9488 = \u11_mem_reg[1][10]/P0001  & n9393 ;
  assign n9489 = \u11_mem_reg[0][10]/P0001  & n9395 ;
  assign n9492 = ~n9488 & ~n9489 ;
  assign n9490 = \u11_mem_reg[3][10]/P0001  & n9397 ;
  assign n9491 = \u11_mem_reg[2][10]/P0001  & n9399 ;
  assign n9493 = ~n9490 & ~n9491 ;
  assign n9494 = n9492 & n9493 ;
  assign n9495 = \u10_mem_reg[0][30]/P0001  & n9314 ;
  assign n9496 = \u10_mem_reg[2][30]/P0001  & n9312 ;
  assign n9499 = ~n9495 & ~n9496 ;
  assign n9497 = \u10_mem_reg[3][30]/P0001  & n9316 ;
  assign n9498 = \u10_mem_reg[1][30]/P0001  & n9318 ;
  assign n9500 = ~n9497 & ~n9498 ;
  assign n9501 = n9499 & n9500 ;
  assign n9502 = \u11_mem_reg[1][11]/P0001  & n9393 ;
  assign n9503 = \u11_mem_reg[0][11]/P0001  & n9395 ;
  assign n9506 = ~n9502 & ~n9503 ;
  assign n9504 = \u11_mem_reg[3][11]/P0001  & n9397 ;
  assign n9505 = \u11_mem_reg[2][11]/P0001  & n9399 ;
  assign n9507 = ~n9504 & ~n9505 ;
  assign n9508 = n9506 & n9507 ;
  assign n9509 = \u11_mem_reg[1][12]/P0001  & n9393 ;
  assign n9510 = \u11_mem_reg[0][12]/P0001  & n9395 ;
  assign n9513 = ~n9509 & ~n9510 ;
  assign n9511 = \u11_mem_reg[3][12]/P0001  & n9397 ;
  assign n9512 = \u11_mem_reg[2][12]/P0001  & n9399 ;
  assign n9514 = ~n9511 & ~n9512 ;
  assign n9515 = n9513 & n9514 ;
  assign n9516 = \u11_mem_reg[1][13]/P0001  & n9393 ;
  assign n9517 = \u11_mem_reg[0][13]/P0001  & n9395 ;
  assign n9520 = ~n9516 & ~n9517 ;
  assign n9518 = \u11_mem_reg[3][13]/P0001  & n9397 ;
  assign n9519 = \u11_mem_reg[2][13]/P0001  & n9399 ;
  assign n9521 = ~n9518 & ~n9519 ;
  assign n9522 = n9520 & n9521 ;
  assign n9523 = \u11_mem_reg[2][14]/P0001  & n9399 ;
  assign n9524 = \u11_mem_reg[0][14]/P0001  & n9395 ;
  assign n9527 = ~n9523 & ~n9524 ;
  assign n9525 = \u11_mem_reg[3][14]/P0001  & n9397 ;
  assign n9526 = \u11_mem_reg[1][14]/P0001  & n9393 ;
  assign n9528 = ~n9525 & ~n9526 ;
  assign n9529 = n9527 & n9528 ;
  assign n9530 = \u10_mem_reg[2][3]/P0001  & n9312 ;
  assign n9531 = \u10_mem_reg[1][3]/P0001  & n9318 ;
  assign n9534 = ~n9530 & ~n9531 ;
  assign n9532 = \u10_mem_reg[3][3]/P0001  & n9316 ;
  assign n9533 = \u10_mem_reg[0][3]/P0001  & n9314 ;
  assign n9535 = ~n9532 & ~n9533 ;
  assign n9536 = n9534 & n9535 ;
  assign n9537 = \u11_mem_reg[1][15]/P0001  & n9393 ;
  assign n9538 = \u11_mem_reg[0][15]/P0001  & n9395 ;
  assign n9541 = ~n9537 & ~n9538 ;
  assign n9539 = \u11_mem_reg[3][15]/P0001  & n9397 ;
  assign n9540 = \u11_mem_reg[2][15]/P0001  & n9399 ;
  assign n9542 = ~n9539 & ~n9540 ;
  assign n9543 = n9541 & n9542 ;
  assign n9544 = \u11_mem_reg[1][16]/P0001  & n9393 ;
  assign n9545 = \u11_mem_reg[0][16]/P0001  & n9395 ;
  assign n9548 = ~n9544 & ~n9545 ;
  assign n9546 = \u11_mem_reg[3][16]/P0001  & n9397 ;
  assign n9547 = \u11_mem_reg[2][16]/P0001  & n9399 ;
  assign n9549 = ~n9546 & ~n9547 ;
  assign n9550 = n9548 & n9549 ;
  assign n9551 = \u10_mem_reg[2][4]/P0001  & n9312 ;
  assign n9552 = \u10_mem_reg[1][4]/P0001  & n9318 ;
  assign n9555 = ~n9551 & ~n9552 ;
  assign n9553 = \u10_mem_reg[3][4]/P0001  & n9316 ;
  assign n9554 = \u10_mem_reg[0][4]/P0001  & n9314 ;
  assign n9556 = ~n9553 & ~n9554 ;
  assign n9557 = n9555 & n9556 ;
  assign n9558 = \u11_mem_reg[1][17]/P0001  & n9393 ;
  assign n9559 = \u11_mem_reg[0][17]/P0001  & n9395 ;
  assign n9562 = ~n9558 & ~n9559 ;
  assign n9560 = \u11_mem_reg[3][17]/P0001  & n9397 ;
  assign n9561 = \u11_mem_reg[2][17]/P0001  & n9399 ;
  assign n9563 = ~n9560 & ~n9561 ;
  assign n9564 = n9562 & n9563 ;
  assign n9565 = \u11_mem_reg[2][18]/P0001  & n9399 ;
  assign n9566 = \u11_mem_reg[1][18]/P0001  & n9393 ;
  assign n9569 = ~n9565 & ~n9566 ;
  assign n9567 = \u11_mem_reg[3][18]/P0001  & n9397 ;
  assign n9568 = \u11_mem_reg[0][18]/P0001  & n9395 ;
  assign n9570 = ~n9567 & ~n9568 ;
  assign n9571 = n9569 & n9570 ;
  assign n9572 = \u10_mem_reg[2][5]/P0001  & n9312 ;
  assign n9573 = \u10_mem_reg[0][5]/P0001  & n9314 ;
  assign n9576 = ~n9572 & ~n9573 ;
  assign n9574 = \u10_mem_reg[3][5]/P0001  & n9316 ;
  assign n9575 = \u10_mem_reg[1][5]/P0001  & n9318 ;
  assign n9577 = ~n9574 & ~n9575 ;
  assign n9578 = n9576 & n9577 ;
  assign n9579 = \u11_mem_reg[2][19]/P0001  & n9399 ;
  assign n9580 = \u11_mem_reg[1][19]/P0001  & n9393 ;
  assign n9583 = ~n9579 & ~n9580 ;
  assign n9581 = \u11_mem_reg[3][19]/P0001  & n9397 ;
  assign n9582 = \u11_mem_reg[0][19]/P0001  & n9395 ;
  assign n9584 = ~n9581 & ~n9582 ;
  assign n9585 = n9583 & n9584 ;
  assign n9586 = \u11_mem_reg[1][1]/P0001  & n9393 ;
  assign n9587 = \u11_mem_reg[0][1]/P0001  & n9395 ;
  assign n9590 = ~n9586 & ~n9587 ;
  assign n9588 = \u11_mem_reg[3][1]/P0001  & n9397 ;
  assign n9589 = \u11_mem_reg[2][1]/P0001  & n9399 ;
  assign n9591 = ~n9588 & ~n9589 ;
  assign n9592 = n9590 & n9591 ;
  assign n9593 = \u10_mem_reg[2][6]/P0001  & n9312 ;
  assign n9594 = \u10_mem_reg[1][6]/P0001  & n9318 ;
  assign n9597 = ~n9593 & ~n9594 ;
  assign n9595 = \u10_mem_reg[3][6]/P0001  & n9316 ;
  assign n9596 = \u10_mem_reg[0][6]/P0001  & n9314 ;
  assign n9598 = ~n9595 & ~n9596 ;
  assign n9599 = n9597 & n9598 ;
  assign n9600 = \u11_mem_reg[2][20]/P0001  & n9399 ;
  assign n9601 = \u11_mem_reg[1][20]/P0001  & n9393 ;
  assign n9604 = ~n9600 & ~n9601 ;
  assign n9602 = \u11_mem_reg[3][20]/P0001  & n9397 ;
  assign n9603 = \u11_mem_reg[0][20]/P0001  & n9395 ;
  assign n9605 = ~n9602 & ~n9603 ;
  assign n9606 = n9604 & n9605 ;
  assign n9607 = \u11_mem_reg[1][21]/P0001  & n9393 ;
  assign n9608 = \u11_mem_reg[2][21]/P0001  & n9399 ;
  assign n9611 = ~n9607 & ~n9608 ;
  assign n9609 = \u11_mem_reg[3][21]/P0001  & n9397 ;
  assign n9610 = \u11_mem_reg[0][21]/P0001  & n9395 ;
  assign n9612 = ~n9609 & ~n9610 ;
  assign n9613 = n9611 & n9612 ;
  assign n9614 = \u10_mem_reg[2][7]/P0001  & n9312 ;
  assign n9615 = \u10_mem_reg[1][7]/P0001  & n9318 ;
  assign n9618 = ~n9614 & ~n9615 ;
  assign n9616 = \u10_mem_reg[3][7]/P0001  & n9316 ;
  assign n9617 = \u10_mem_reg[0][7]/P0001  & n9314 ;
  assign n9619 = ~n9616 & ~n9617 ;
  assign n9620 = n9618 & n9619 ;
  assign n9621 = \u11_mem_reg[2][22]/P0001  & n9399 ;
  assign n9622 = \u11_mem_reg[1][22]/P0001  & n9393 ;
  assign n9625 = ~n9621 & ~n9622 ;
  assign n9623 = \u11_mem_reg[3][22]/P0001  & n9397 ;
  assign n9624 = \u11_mem_reg[0][22]/P0001  & n9395 ;
  assign n9626 = ~n9623 & ~n9624 ;
  assign n9627 = n9625 & n9626 ;
  assign n9628 = \u11_mem_reg[2][23]/P0001  & n9399 ;
  assign n9629 = \u11_mem_reg[1][23]/P0001  & n9393 ;
  assign n9632 = ~n9628 & ~n9629 ;
  assign n9630 = \u11_mem_reg[3][23]/P0001  & n9397 ;
  assign n9631 = \u11_mem_reg[0][23]/P0001  & n9395 ;
  assign n9633 = ~n9630 & ~n9631 ;
  assign n9634 = n9632 & n9633 ;
  assign n9635 = \u10_mem_reg[2][8]/P0001  & n9312 ;
  assign n9636 = \u10_mem_reg[0][8]/P0001  & n9314 ;
  assign n9639 = ~n9635 & ~n9636 ;
  assign n9637 = \u10_mem_reg[3][8]/P0001  & n9316 ;
  assign n9638 = \u10_mem_reg[1][8]/P0001  & n9318 ;
  assign n9640 = ~n9637 & ~n9638 ;
  assign n9641 = n9639 & n9640 ;
  assign n9642 = \u11_mem_reg[2][24]/P0001  & n9399 ;
  assign n9643 = \u11_mem_reg[1][24]/P0001  & n9393 ;
  assign n9646 = ~n9642 & ~n9643 ;
  assign n9644 = \u11_mem_reg[3][24]/P0001  & n9397 ;
  assign n9645 = \u11_mem_reg[0][24]/P0001  & n9395 ;
  assign n9647 = ~n9644 & ~n9645 ;
  assign n9648 = n9646 & n9647 ;
  assign n9649 = \u11_mem_reg[2][25]/P0001  & n9399 ;
  assign n9650 = \u11_mem_reg[1][25]/P0001  & n9393 ;
  assign n9653 = ~n9649 & ~n9650 ;
  assign n9651 = \u11_mem_reg[3][25]/P0001  & n9397 ;
  assign n9652 = \u11_mem_reg[0][25]/P0001  & n9395 ;
  assign n9654 = ~n9651 & ~n9652 ;
  assign n9655 = n9653 & n9654 ;
  assign n9656 = \u10_mem_reg[1][9]/P0001  & n9318 ;
  assign n9657 = \u10_mem_reg[0][9]/P0001  & n9314 ;
  assign n9660 = ~n9656 & ~n9657 ;
  assign n9658 = \u10_mem_reg[3][9]/P0001  & n9316 ;
  assign n9659 = \u10_mem_reg[2][9]/P0001  & n9312 ;
  assign n9661 = ~n9658 & ~n9659 ;
  assign n9662 = n9660 & n9661 ;
  assign n9663 = \u11_mem_reg[2][26]/P0001  & n9399 ;
  assign n9664 = \u11_mem_reg[1][26]/P0001  & n9393 ;
  assign n9667 = ~n9663 & ~n9664 ;
  assign n9665 = \u11_mem_reg[3][26]/P0001  & n9397 ;
  assign n9666 = \u11_mem_reg[0][26]/P0001  & n9395 ;
  assign n9668 = ~n9665 & ~n9666 ;
  assign n9669 = n9667 & n9668 ;
  assign n9670 = \u11_mem_reg[2][27]/P0001  & n9399 ;
  assign n9671 = \u11_mem_reg[1][27]/P0001  & n9393 ;
  assign n9674 = ~n9670 & ~n9671 ;
  assign n9672 = \u11_mem_reg[3][27]/P0001  & n9397 ;
  assign n9673 = \u11_mem_reg[0][27]/P0001  & n9395 ;
  assign n9675 = ~n9672 & ~n9673 ;
  assign n9676 = n9674 & n9675 ;
  assign n9677 = \u11_mem_reg[2][28]/P0001  & n9399 ;
  assign n9678 = \u11_mem_reg[1][28]/P0001  & n9393 ;
  assign n9681 = ~n9677 & ~n9678 ;
  assign n9679 = \u11_mem_reg[3][28]/P0001  & n9397 ;
  assign n9680 = \u11_mem_reg[0][28]/P0001  & n9395 ;
  assign n9682 = ~n9679 & ~n9680 ;
  assign n9683 = n9681 & n9682 ;
  assign n9684 = \u10_mem_reg[3][14]/P0001  & n9316 ;
  assign n9685 = \u10_mem_reg[2][14]/P0001  & n9312 ;
  assign n9688 = ~n9684 & ~n9685 ;
  assign n9686 = \u10_mem_reg[0][14]/P0001  & n9314 ;
  assign n9687 = \u10_mem_reg[1][14]/P0001  & n9318 ;
  assign n9689 = ~n9686 & ~n9687 ;
  assign n9690 = n9688 & n9689 ;
  assign n9691 = \u11_mem_reg[2][29]/P0001  & n9399 ;
  assign n9692 = \u11_mem_reg[1][29]/P0001  & n9393 ;
  assign n9695 = ~n9691 & ~n9692 ;
  assign n9693 = \u11_mem_reg[3][29]/P0001  & n9397 ;
  assign n9694 = \u11_mem_reg[0][29]/P0001  & n9395 ;
  assign n9696 = ~n9693 & ~n9694 ;
  assign n9697 = n9695 & n9696 ;
  assign n9698 = \u11_mem_reg[1][2]/P0001  & n9393 ;
  assign n9699 = \u11_mem_reg[0][2]/P0001  & n9395 ;
  assign n9702 = ~n9698 & ~n9699 ;
  assign n9700 = \u11_mem_reg[3][2]/P0001  & n9397 ;
  assign n9701 = \u11_mem_reg[2][2]/P0001  & n9399 ;
  assign n9703 = ~n9700 & ~n9701 ;
  assign n9704 = n9702 & n9703 ;
  assign n9705 = \u11_mem_reg[2][30]/P0001  & n9399 ;
  assign n9706 = \u11_mem_reg[1][30]/P0001  & n9393 ;
  assign n9709 = ~n9705 & ~n9706 ;
  assign n9707 = \u11_mem_reg[3][30]/P0001  & n9397 ;
  assign n9708 = \u11_mem_reg[0][30]/P0001  & n9395 ;
  assign n9710 = ~n9707 & ~n9708 ;
  assign n9711 = n9709 & n9710 ;
  assign n9712 = \u11_mem_reg[2][31]/P0001  & n9399 ;
  assign n9713 = \u11_mem_reg[1][31]/P0001  & n9393 ;
  assign n9716 = ~n9712 & ~n9713 ;
  assign n9714 = \u11_mem_reg[3][31]/P0001  & n9397 ;
  assign n9715 = \u11_mem_reg[0][31]/P0001  & n9395 ;
  assign n9717 = ~n9714 & ~n9715 ;
  assign n9718 = n9716 & n9717 ;
  assign n9719 = \u11_mem_reg[1][3]/P0001  & n9393 ;
  assign n9720 = \u11_mem_reg[0][3]/P0001  & n9395 ;
  assign n9723 = ~n9719 & ~n9720 ;
  assign n9721 = \u11_mem_reg[3][3]/P0001  & n9397 ;
  assign n9722 = \u11_mem_reg[2][3]/P0001  & n9399 ;
  assign n9724 = ~n9721 & ~n9722 ;
  assign n9725 = n9723 & n9724 ;
  assign n9726 = \u11_mem_reg[1][4]/P0001  & n9393 ;
  assign n9727 = \u11_mem_reg[0][4]/P0001  & n9395 ;
  assign n9730 = ~n9726 & ~n9727 ;
  assign n9728 = \u11_mem_reg[3][4]/P0001  & n9397 ;
  assign n9729 = \u11_mem_reg[2][4]/P0001  & n9399 ;
  assign n9731 = ~n9728 & ~n9729 ;
  assign n9732 = n9730 & n9731 ;
  assign n9733 = \u11_mem_reg[1][5]/P0001  & n9393 ;
  assign n9734 = \u11_mem_reg[0][5]/P0001  & n9395 ;
  assign n9737 = ~n9733 & ~n9734 ;
  assign n9735 = \u11_mem_reg[3][5]/P0001  & n9397 ;
  assign n9736 = \u11_mem_reg[2][5]/P0001  & n9399 ;
  assign n9738 = ~n9735 & ~n9736 ;
  assign n9739 = n9737 & n9738 ;
  assign n9740 = \u11_mem_reg[2][7]/P0001  & n9399 ;
  assign n9741 = \u11_mem_reg[0][7]/P0001  & n9395 ;
  assign n9744 = ~n9740 & ~n9741 ;
  assign n9742 = \u11_mem_reg[3][7]/P0001  & n9397 ;
  assign n9743 = \u11_mem_reg[1][7]/P0001  & n9393 ;
  assign n9745 = ~n9742 & ~n9743 ;
  assign n9746 = n9744 & n9745 ;
  assign n9747 = \u11_mem_reg[1][8]/P0001  & n9393 ;
  assign n9748 = \u11_mem_reg[0][8]/P0001  & n9395 ;
  assign n9751 = ~n9747 & ~n9748 ;
  assign n9749 = \u11_mem_reg[3][8]/P0001  & n9397 ;
  assign n9750 = \u11_mem_reg[2][8]/P0001  & n9399 ;
  assign n9752 = ~n9749 & ~n9750 ;
  assign n9753 = n9751 & n9752 ;
  assign n9754 = \u11_mem_reg[1][9]/P0001  & n9393 ;
  assign n9755 = \u11_mem_reg[0][9]/P0001  & n9395 ;
  assign n9758 = ~n9754 & ~n9755 ;
  assign n9756 = \u11_mem_reg[3][9]/P0001  & n9397 ;
  assign n9757 = \u11_mem_reg[2][9]/P0001  & n9399 ;
  assign n9759 = ~n9756 & ~n9757 ;
  assign n9760 = n9758 & n9759 ;
  assign n9761 = \u10_mem_reg[2][10]/P0001  & n9312 ;
  assign n9762 = \u10_mem_reg[0][10]/P0001  & n9314 ;
  assign n9765 = ~n9761 & ~n9762 ;
  assign n9763 = \u10_mem_reg[3][10]/P0001  & n9316 ;
  assign n9764 = \u10_mem_reg[1][10]/P0001  & n9318 ;
  assign n9766 = ~n9763 & ~n9764 ;
  assign n9767 = n9765 & n9766 ;
  assign n9768 = \u10_mem_reg[2][2]/P0001  & n9312 ;
  assign n9769 = \u10_mem_reg[1][2]/P0001  & n9318 ;
  assign n9772 = ~n9768 & ~n9769 ;
  assign n9770 = \u10_mem_reg[3][2]/P0001  & n9316 ;
  assign n9771 = \u10_mem_reg[0][2]/P0001  & n9314 ;
  assign n9773 = ~n9770 & ~n9771 ;
  assign n9774 = n9772 & n9773 ;
  assign n9775 = \u9_mem_reg[1][8]/P0001  & n9112 ;
  assign n9776 = \u9_mem_reg[0][8]/P0001  & n9114 ;
  assign n9779 = ~n9775 & ~n9776 ;
  assign n9777 = \u9_mem_reg[3][8]/P0001  & n9116 ;
  assign n9778 = \u9_mem_reg[2][8]/P0001  & n9118 ;
  assign n9780 = ~n9777 & ~n9778 ;
  assign n9781 = n9779 & n9780 ;
  assign n9782 = \u10_mem_reg[1][31]/P0001  & n9318 ;
  assign n9783 = \u10_mem_reg[2][31]/P0001  & n9312 ;
  assign n9786 = ~n9782 & ~n9783 ;
  assign n9784 = \u10_mem_reg[3][31]/P0001  & n9316 ;
  assign n9785 = \u10_mem_reg[0][31]/P0001  & n9314 ;
  assign n9787 = ~n9784 & ~n9785 ;
  assign n9788 = n9786 & n9787 ;
  assign n9789 = \u9_mem_reg[1][9]/P0001  & n9112 ;
  assign n9790 = \u9_mem_reg[0][9]/P0001  & n9114 ;
  assign n9793 = ~n9789 & ~n9790 ;
  assign n9791 = \u9_mem_reg[3][9]/P0001  & n9116 ;
  assign n9792 = \u9_mem_reg[2][9]/P0001  & n9118 ;
  assign n9794 = ~n9791 & ~n9792 ;
  assign n9795 = n9793 & n9794 ;
  assign n9799 = \u10_din_tmp1_reg[3]/P0001  & n3501 ;
  assign n9796 = \u13_icc_r_reg[10]/NET0131  & ~\u13_icc_r_reg[11]/NET0131  ;
  assign n9797 = \u1_slt4_reg[5]/P0001  & n9796 ;
  assign n9798 = \u1_slt4_reg[3]/P0001  & n5671 ;
  assign n9800 = ~n9797 & ~n9798 ;
  assign n9801 = ~n9799 & n9800 ;
  assign n9802 = n2737 & n9018 ;
  assign n9806 = \u9_din_tmp1_reg[1]/P0001  & n3311 ;
  assign n9803 = \u1_slt3_reg[1]/P0001  & n5701 ;
  assign n9804 = \u13_icc_r_reg[2]/NET0131  & ~\u13_icc_r_reg[3]/NET0131  ;
  assign n9805 = \u1_slt3_reg[3]/P0001  & n9804 ;
  assign n9807 = ~n9803 & ~n9805 ;
  assign n9808 = ~n9806 & n9807 ;
  assign n9811 = \u9_din_tmp1_reg[2]/P0001  & n3311 ;
  assign n9809 = \u1_slt3_reg[2]/P0001  & n5701 ;
  assign n9810 = \u1_slt3_reg[4]/P0001  & n9804 ;
  assign n9812 = ~n9809 & ~n9810 ;
  assign n9813 = ~n9811 & n9812 ;
  assign n9816 = \u9_din_tmp1_reg[8]/P0001  & n3311 ;
  assign n9814 = \u1_slt3_reg[8]/P0001  & n5701 ;
  assign n9815 = \u1_slt3_reg[10]/P0001  & n9804 ;
  assign n9817 = ~n9814 & ~n9815 ;
  assign n9818 = ~n9816 & n9817 ;
  assign n9821 = \u1_slt3_reg[19]/P0001  & n9804 ;
  assign n9819 = \u1_slt3_reg[17]/P0001  & n5701 ;
  assign n9820 = \u1_slt3_reg[5]/P0001  & n3311 ;
  assign n9822 = ~n9819 & ~n9820 ;
  assign n9823 = ~n9821 & n9822 ;
  assign n9826 = \u1_slt3_reg[18]/P0001  & n9804 ;
  assign n9824 = \u1_slt3_reg[16]/P0001  & n5701 ;
  assign n9825 = \u1_slt3_reg[4]/P0001  & n3311 ;
  assign n9827 = ~n9824 & ~n9825 ;
  assign n9828 = ~n9826 & n9827 ;
  assign n9831 = \u9_din_tmp1_reg[15]/P0001  & n3311 ;
  assign n9829 = \u1_slt3_reg[15]/P0001  & n5701 ;
  assign n9830 = \u1_slt3_reg[17]/P0001  & n9804 ;
  assign n9832 = ~n9829 & ~n9830 ;
  assign n9833 = ~n9831 & n9832 ;
  assign n9836 = \u9_din_tmp1_reg[14]/P0001  & n3311 ;
  assign n9834 = \u1_slt3_reg[14]/P0001  & n5701 ;
  assign n9835 = \u1_slt3_reg[16]/P0001  & n9804 ;
  assign n9837 = ~n9834 & ~n9835 ;
  assign n9838 = ~n9836 & n9837 ;
  assign n9841 = \u9_din_tmp1_reg[13]/P0001  & n3311 ;
  assign n9839 = \u1_slt3_reg[13]/P0001  & n5701 ;
  assign n9840 = \u1_slt3_reg[15]/P0001  & n9804 ;
  assign n9842 = ~n9839 & ~n9840 ;
  assign n9843 = ~n9841 & n9842 ;
  assign n9846 = \u9_din_tmp1_reg[12]/P0001  & n3311 ;
  assign n9844 = \u1_slt3_reg[12]/P0001  & n5701 ;
  assign n9845 = \u1_slt3_reg[14]/P0001  & n9804 ;
  assign n9847 = ~n9844 & ~n9845 ;
  assign n9848 = ~n9846 & n9847 ;
  assign n9851 = \u9_din_tmp1_reg[11]/P0001  & n3311 ;
  assign n9849 = \u1_slt3_reg[13]/P0001  & n9804 ;
  assign n9850 = \u1_slt3_reg[11]/P0001  & n5701 ;
  assign n9852 = ~n9849 & ~n9850 ;
  assign n9853 = ~n9851 & n9852 ;
  assign n9856 = \u9_din_tmp1_reg[9]/P0001  & n3311 ;
  assign n9854 = \u1_slt3_reg[9]/P0001  & n5701 ;
  assign n9855 = \u1_slt3_reg[11]/P0001  & n9804 ;
  assign n9857 = ~n9854 & ~n9855 ;
  assign n9858 = ~n9856 & n9857 ;
  assign n9861 = \u9_din_tmp1_reg[3]/P0001  & n3311 ;
  assign n9859 = \u1_slt3_reg[3]/P0001  & n5701 ;
  assign n9860 = \u1_slt3_reg[5]/P0001  & n9804 ;
  assign n9862 = ~n9859 & ~n9860 ;
  assign n9863 = ~n9861 & n9862 ;
  assign n9866 = \u9_din_tmp1_reg[10]/P0001  & n3311 ;
  assign n9864 = \u1_slt3_reg[12]/P0001  & n9804 ;
  assign n9865 = \u1_slt3_reg[10]/P0001  & n5701 ;
  assign n9867 = ~n9864 & ~n9865 ;
  assign n9868 = ~n9866 & n9867 ;
  assign n9872 = \u11_din_tmp1_reg[11]/P0001  & n3064 ;
  assign n9869 = \u13_icc_r_reg[18]/NET0131  & ~\u13_icc_r_reg[19]/NET0131  ;
  assign n9870 = \u1_slt6_reg[13]/P0001  & n9869 ;
  assign n9871 = \u1_slt6_reg[11]/P0001  & n5936 ;
  assign n9873 = ~n9870 & ~n9871 ;
  assign n9874 = ~n9872 & n9873 ;
  assign n9877 = \u10_din_tmp1_reg[9]/P0001  & n3501 ;
  assign n9875 = \u1_slt4_reg[9]/P0001  & n5671 ;
  assign n9876 = \u1_slt4_reg[11]/P0001  & n9796 ;
  assign n9878 = ~n9875 & ~n9876 ;
  assign n9879 = ~n9877 & n9878 ;
  assign n9882 = \u9_din_tmp1_reg[6]/P0001  & n3311 ;
  assign n9880 = \u1_slt3_reg[6]/P0001  & n5701 ;
  assign n9881 = \u1_slt3_reg[8]/P0001  & n9804 ;
  assign n9883 = ~n9880 & ~n9881 ;
  assign n9884 = ~n9882 & n9883 ;
  assign n9887 = \u10_din_tmp1_reg[0]/P0001  & n3501 ;
  assign n9885 = \u1_slt4_reg[0]/P0001  & n5671 ;
  assign n9886 = \u1_slt4_reg[2]/P0001  & n9796 ;
  assign n9888 = ~n9885 & ~n9886 ;
  assign n9889 = ~n9887 & n9888 ;
  assign n9892 = \u10_din_tmp1_reg[10]/P0001  & n3501 ;
  assign n9890 = \u1_slt4_reg[12]/P0001  & n9796 ;
  assign n9891 = \u1_slt4_reg[10]/P0001  & n5671 ;
  assign n9893 = ~n9890 & ~n9891 ;
  assign n9894 = ~n9892 & n9893 ;
  assign n9897 = \u10_din_tmp1_reg[11]/P0001  & n3501 ;
  assign n9895 = \u1_slt4_reg[13]/P0001  & n9796 ;
  assign n9896 = \u1_slt4_reg[11]/P0001  & n5671 ;
  assign n9898 = ~n9895 & ~n9896 ;
  assign n9899 = ~n9897 & n9898 ;
  assign n9902 = \u10_din_tmp1_reg[12]/P0001  & n3501 ;
  assign n9900 = \u1_slt4_reg[14]/P0001  & n9796 ;
  assign n9901 = \u1_slt4_reg[12]/P0001  & n5671 ;
  assign n9903 = ~n9900 & ~n9901 ;
  assign n9904 = ~n9902 & n9903 ;
  assign n9907 = \u9_din_tmp1_reg[7]/P0001  & n3311 ;
  assign n9905 = \u1_slt3_reg[7]/P0001  & n5701 ;
  assign n9906 = \u1_slt3_reg[9]/P0001  & n9804 ;
  assign n9908 = ~n9905 & ~n9906 ;
  assign n9909 = ~n9907 & n9908 ;
  assign n9912 = \u10_din_tmp1_reg[13]/P0001  & n3501 ;
  assign n9910 = \u1_slt4_reg[15]/P0001  & n9796 ;
  assign n9911 = \u1_slt4_reg[13]/P0001  & n5671 ;
  assign n9913 = ~n9910 & ~n9911 ;
  assign n9914 = ~n9912 & n9913 ;
  assign n9917 = \u9_din_tmp1_reg[5]/P0001  & n3311 ;
  assign n9915 = \u1_slt3_reg[5]/P0001  & n5701 ;
  assign n9916 = \u1_slt3_reg[7]/P0001  & n9804 ;
  assign n9918 = ~n9915 & ~n9916 ;
  assign n9919 = ~n9917 & n9918 ;
  assign n9922 = \u11_din_tmp1_reg[0]/P0001  & n3064 ;
  assign n9920 = \u1_slt6_reg[0]/P0001  & n5936 ;
  assign n9921 = \u1_slt6_reg[2]/P0001  & n9869 ;
  assign n9923 = ~n9920 & ~n9921 ;
  assign n9924 = ~n9922 & n9923 ;
  assign n9927 = \u11_din_tmp1_reg[10]/P0001  & n3064 ;
  assign n9925 = \u1_slt6_reg[12]/P0001  & n9869 ;
  assign n9926 = \u1_slt6_reg[10]/P0001  & n5936 ;
  assign n9928 = ~n9925 & ~n9926 ;
  assign n9929 = ~n9927 & n9928 ;
  assign n9932 = \u10_din_tmp1_reg[15]/P0001  & n3501 ;
  assign n9930 = \u1_slt4_reg[17]/P0001  & n9796 ;
  assign n9931 = \u1_slt4_reg[15]/P0001  & n5671 ;
  assign n9933 = ~n9930 & ~n9931 ;
  assign n9934 = ~n9932 & n9933 ;
  assign n9937 = \u11_din_tmp1_reg[12]/P0001  & n3064 ;
  assign n9935 = \u1_slt6_reg[14]/P0001  & n9869 ;
  assign n9936 = \u1_slt6_reg[12]/P0001  & n5936 ;
  assign n9938 = ~n9935 & ~n9936 ;
  assign n9939 = ~n9937 & n9938 ;
  assign n9942 = \u11_din_tmp1_reg[13]/P0001  & n3064 ;
  assign n9940 = \u1_slt6_reg[15]/P0001  & n9869 ;
  assign n9941 = \u1_slt6_reg[13]/P0001  & n5936 ;
  assign n9943 = ~n9940 & ~n9941 ;
  assign n9944 = ~n9942 & n9943 ;
  assign n9947 = \u1_slt4_reg[16]/P0001  & n5671 ;
  assign n9945 = \u1_slt4_reg[18]/P0001  & n9796 ;
  assign n9946 = \u1_slt4_reg[4]/P0001  & n3501 ;
  assign n9948 = ~n9945 & ~n9946 ;
  assign n9949 = ~n9947 & n9948 ;
  assign n9952 = \u11_din_tmp1_reg[14]/P0001  & n3064 ;
  assign n9950 = \u1_slt6_reg[16]/P0001  & n9869 ;
  assign n9951 = \u1_slt6_reg[14]/P0001  & n5936 ;
  assign n9953 = ~n9950 & ~n9951 ;
  assign n9954 = ~n9952 & n9953 ;
  assign n9957 = \u1_slt4_reg[17]/P0001  & n5671 ;
  assign n9955 = \u1_slt4_reg[19]/P0001  & n9796 ;
  assign n9956 = \u1_slt4_reg[5]/P0001  & n3501 ;
  assign n9958 = ~n9955 & ~n9956 ;
  assign n9959 = ~n9957 & n9958 ;
  assign n9962 = \u1_slt6_reg[17]/P0001  & n5936 ;
  assign n9960 = \u1_slt6_reg[19]/P0001  & n9869 ;
  assign n9961 = \u1_slt6_reg[5]/P0001  & n3064 ;
  assign n9963 = ~n9960 & ~n9961 ;
  assign n9964 = ~n9962 & n9963 ;
  assign n9967 = \u11_din_tmp1_reg[1]/P0001  & n3064 ;
  assign n9965 = \u1_slt6_reg[1]/P0001  & n5936 ;
  assign n9966 = \u1_slt6_reg[3]/P0001  & n9869 ;
  assign n9968 = ~n9965 & ~n9966 ;
  assign n9969 = ~n9967 & n9968 ;
  assign n9972 = \u10_din_tmp1_reg[1]/P0001  & n3501 ;
  assign n9970 = \u1_slt4_reg[1]/P0001  & n5671 ;
  assign n9971 = \u1_slt4_reg[3]/P0001  & n9796 ;
  assign n9973 = ~n9970 & ~n9971 ;
  assign n9974 = ~n9972 & n9973 ;
  assign n9977 = \u10_din_tmp1_reg[14]/P0001  & n3501 ;
  assign n9975 = \u1_slt4_reg[16]/P0001  & n9796 ;
  assign n9976 = \u1_slt4_reg[14]/P0001  & n5671 ;
  assign n9978 = ~n9975 & ~n9976 ;
  assign n9979 = ~n9977 & n9978 ;
  assign n9982 = \u11_din_tmp1_reg[2]/P0001  & n3064 ;
  assign n9980 = \u1_slt6_reg[4]/P0001  & n9869 ;
  assign n9981 = \u1_slt6_reg[2]/P0001  & n5936 ;
  assign n9983 = ~n9980 & ~n9981 ;
  assign n9984 = ~n9982 & n9983 ;
  assign n9987 = \u1_slt6_reg[16]/P0001  & n5936 ;
  assign n9985 = \u1_slt6_reg[18]/P0001  & n9869 ;
  assign n9986 = \u1_slt6_reg[4]/P0001  & n3064 ;
  assign n9988 = ~n9985 & ~n9986 ;
  assign n9989 = ~n9987 & n9988 ;
  assign n9992 = \u11_din_tmp1_reg[3]/P0001  & n3064 ;
  assign n9990 = \u1_slt6_reg[5]/P0001  & n9869 ;
  assign n9991 = \u1_slt6_reg[3]/P0001  & n5936 ;
  assign n9993 = ~n9990 & ~n9991 ;
  assign n9994 = ~n9992 & n9993 ;
  assign n9997 = \u11_din_tmp1_reg[4]/P0001  & n3064 ;
  assign n9995 = \u1_slt6_reg[6]/P0001  & n9869 ;
  assign n9996 = \u1_slt6_reg[4]/P0001  & n5936 ;
  assign n9998 = ~n9995 & ~n9996 ;
  assign n9999 = ~n9997 & n9998 ;
  assign n10002 = \u11_din_tmp1_reg[5]/P0001  & n3064 ;
  assign n10000 = \u1_slt6_reg[7]/P0001  & n9869 ;
  assign n10001 = \u1_slt6_reg[5]/P0001  & n5936 ;
  assign n10003 = ~n10000 & ~n10001 ;
  assign n10004 = ~n10002 & n10003 ;
  assign n10007 = \u11_din_tmp1_reg[6]/P0001  & n3064 ;
  assign n10005 = \u1_slt6_reg[8]/P0001  & n9869 ;
  assign n10006 = \u1_slt6_reg[6]/P0001  & n5936 ;
  assign n10008 = ~n10005 & ~n10006 ;
  assign n10009 = ~n10007 & n10008 ;
  assign n10012 = \u11_din_tmp1_reg[7]/P0001  & n3064 ;
  assign n10010 = \u1_slt6_reg[9]/P0001  & n9869 ;
  assign n10011 = \u1_slt6_reg[7]/P0001  & n5936 ;
  assign n10013 = ~n10010 & ~n10011 ;
  assign n10014 = ~n10012 & n10013 ;
  assign n10017 = \u11_din_tmp1_reg[8]/P0001  & n3064 ;
  assign n10015 = \u1_slt6_reg[10]/P0001  & n9869 ;
  assign n10016 = \u1_slt6_reg[8]/P0001  & n5936 ;
  assign n10018 = ~n10015 & ~n10016 ;
  assign n10019 = ~n10017 & n10018 ;
  assign n10022 = \u11_din_tmp1_reg[9]/P0001  & n3064 ;
  assign n10020 = \u1_slt6_reg[9]/P0001  & n5936 ;
  assign n10021 = \u1_slt6_reg[11]/P0001  & n9869 ;
  assign n10023 = ~n10020 & ~n10021 ;
  assign n10024 = ~n10022 & n10023 ;
  assign n10027 = \u10_din_tmp1_reg[2]/P0001  & n3501 ;
  assign n10025 = \u1_slt4_reg[4]/P0001  & n9796 ;
  assign n10026 = \u1_slt4_reg[2]/P0001  & n5671 ;
  assign n10028 = ~n10025 & ~n10026 ;
  assign n10029 = ~n10027 & n10028 ;
  assign n10032 = \u10_din_tmp1_reg[4]/P0001  & n3501 ;
  assign n10030 = \u1_slt4_reg[6]/P0001  & n9796 ;
  assign n10031 = \u1_slt4_reg[4]/P0001  & n5671 ;
  assign n10033 = ~n10030 & ~n10031 ;
  assign n10034 = ~n10032 & n10033 ;
  assign n10037 = \u10_din_tmp1_reg[5]/P0001  & n3501 ;
  assign n10035 = \u1_slt4_reg[7]/P0001  & n9796 ;
  assign n10036 = \u1_slt4_reg[5]/P0001  & n5671 ;
  assign n10038 = ~n10035 & ~n10036 ;
  assign n10039 = ~n10037 & n10038 ;
  assign n10042 = \u10_din_tmp1_reg[6]/P0001  & n3501 ;
  assign n10040 = \u1_slt4_reg[8]/P0001  & n9796 ;
  assign n10041 = \u1_slt4_reg[6]/P0001  & n5671 ;
  assign n10043 = ~n10040 & ~n10041 ;
  assign n10044 = ~n10042 & n10043 ;
  assign n10047 = \u10_din_tmp1_reg[7]/P0001  & n3501 ;
  assign n10045 = \u1_slt4_reg[9]/P0001  & n9796 ;
  assign n10046 = \u1_slt4_reg[7]/P0001  & n5671 ;
  assign n10048 = ~n10045 & ~n10046 ;
  assign n10049 = ~n10047 & n10048 ;
  assign n10052 = \u10_din_tmp1_reg[8]/P0001  & n3501 ;
  assign n10050 = \u1_slt4_reg[10]/P0001  & n9796 ;
  assign n10051 = \u1_slt4_reg[8]/P0001  & n5671 ;
  assign n10053 = ~n10050 & ~n10051 ;
  assign n10054 = ~n10052 & n10053 ;
  assign n10057 = \u11_din_tmp1_reg[15]/P0001  & n3064 ;
  assign n10055 = \u1_slt6_reg[17]/P0001  & n9869 ;
  assign n10056 = \u1_slt6_reg[15]/P0001  & n5936 ;
  assign n10058 = ~n10055 & ~n10056 ;
  assign n10059 = ~n10057 & n10058 ;
  assign n10062 = \u9_din_tmp1_reg[0]/P0001  & n3311 ;
  assign n10060 = \u1_slt3_reg[0]/P0001  & n5701 ;
  assign n10061 = \u1_slt3_reg[2]/P0001  & n9804 ;
  assign n10063 = ~n10060 & ~n10061 ;
  assign n10064 = ~n10062 & n10063 ;
  assign n10067 = \u9_din_tmp1_reg[4]/P0001  & n3311 ;
  assign n10065 = \u1_slt3_reg[4]/P0001  & n5701 ;
  assign n10066 = \u1_slt3_reg[6]/P0001  & n9804 ;
  assign n10068 = ~n10065 & ~n10066 ;
  assign n10069 = ~n10067 & n10068 ;
  assign n10070 = \u2_cnt_reg[0]/NET0131  & ~\u2_cnt_reg[5]/NET0131  ;
  assign n10071 = n9079 & n10070 ;
  assign n10072 = n9109 & n10071 ;
  assign n10073 = \u11_mem_reg[0][24]/P0001  & ~n5933 ;
  assign n10074 = n5933 & n5975 ;
  assign n10075 = ~n10073 & ~n10074 ;
  assign n10076 = \u10_mem_reg[0][20]/P0001  & ~n5928 ;
  assign n10077 = n5683 & n5928 ;
  assign n10078 = ~n10076 & ~n10077 ;
  assign n10079 = \u9_mem_reg[0][31]/P0001  & ~n5698 ;
  assign n10080 = n5698 & n5789 ;
  assign n10081 = ~n10079 & ~n10080 ;
  assign n10082 = \u9_mem_reg[0][20]/P0001  & ~n5698 ;
  assign n10083 = n5698 & n5741 ;
  assign n10084 = ~n10082 & ~n10083 ;
  assign n10085 = \u9_mem_reg[0][21]/P0001  & ~n5698 ;
  assign n10086 = n5698 & n5745 ;
  assign n10087 = ~n10085 & ~n10086 ;
  assign n10088 = \u9_mem_reg[0][23]/P0001  & ~n5698 ;
  assign n10089 = n5698 & n5757 ;
  assign n10090 = ~n10088 & ~n10089 ;
  assign n10091 = \u9_mem_reg[0][24]/P0001  & ~n5698 ;
  assign n10092 = n5698 & n5761 ;
  assign n10093 = ~n10091 & ~n10092 ;
  assign n10094 = \u9_mem_reg[0][25]/P0001  & ~n5698 ;
  assign n10095 = n5698 & n5765 ;
  assign n10096 = ~n10094 & ~n10095 ;
  assign n10097 = \u9_mem_reg[0][26]/P0001  & ~n5698 ;
  assign n10098 = n5698 & n5769 ;
  assign n10099 = ~n10097 & ~n10098 ;
  assign n10100 = \u9_mem_reg[0][27]/P0001  & ~n5698 ;
  assign n10101 = n5698 & n5773 ;
  assign n10102 = ~n10100 & ~n10101 ;
  assign n10103 = \u9_mem_reg[0][28]/P0001  & ~n5698 ;
  assign n10104 = n5698 & n5777 ;
  assign n10105 = ~n10103 & ~n10104 ;
  assign n10106 = \u9_mem_reg[0][29]/P0001  & ~n5698 ;
  assign n10107 = n5698 & n5781 ;
  assign n10108 = ~n10106 & ~n10107 ;
  assign n10109 = \u9_mem_reg[0][30]/P0001  & ~n5698 ;
  assign n10110 = n5698 & n5785 ;
  assign n10111 = ~n10109 & ~n10110 ;
  assign n10112 = \u11_mem_reg[0][21]/P0001  & ~n5933 ;
  assign n10113 = n5933 & n5963 ;
  assign n10114 = ~n10112 & ~n10113 ;
  assign n10115 = \u10_mem_reg[0][22]/P0001  & ~n5928 ;
  assign n10116 = n5691 & n5928 ;
  assign n10117 = ~n10115 & ~n10116 ;
  assign n10118 = \u11_mem_reg[0][27]/P0001  & ~n5933 ;
  assign n10119 = n5933 & n5987 ;
  assign n10120 = ~n10118 & ~n10119 ;
  assign n10121 = \u11_mem_reg[0][31]/P0001  & ~n5933 ;
  assign n10122 = n5933 & n6003 ;
  assign n10123 = ~n10121 & ~n10122 ;
  assign n10124 = \u11_mem_reg[0][29]/P0001  & ~n5933 ;
  assign n10125 = n5933 & n5995 ;
  assign n10126 = ~n10124 & ~n10125 ;
  assign n10127 = \u11_mem_reg[0][20]/P0001  & ~n5933 ;
  assign n10128 = n5933 & n5959 ;
  assign n10129 = ~n10127 & ~n10128 ;
  assign n10130 = \u11_mem_reg[0][22]/P0001  & ~n5933 ;
  assign n10131 = n5933 & n5967 ;
  assign n10132 = ~n10130 & ~n10131 ;
  assign n10133 = \u11_mem_reg[0][23]/P0001  & ~n5933 ;
  assign n10134 = n5933 & n5971 ;
  assign n10135 = ~n10133 & ~n10134 ;
  assign n10136 = \u11_mem_reg[0][25]/P0001  & ~n5933 ;
  assign n10137 = n5933 & n5979 ;
  assign n10138 = ~n10136 & ~n10137 ;
  assign n10139 = \u10_mem_reg[0][21]/P0001  & ~n5928 ;
  assign n10140 = n5687 & n5928 ;
  assign n10141 = ~n10139 & ~n10140 ;
  assign n10142 = \u11_mem_reg[0][26]/P0001  & ~n5933 ;
  assign n10143 = n5933 & n5983 ;
  assign n10144 = ~n10142 & ~n10143 ;
  assign n10145 = \u10_mem_reg[0][23]/P0001  & ~n5928 ;
  assign n10146 = n5695 & n5928 ;
  assign n10147 = ~n10145 & ~n10146 ;
  assign n10148 = \u11_mem_reg[0][30]/P0001  & ~n5933 ;
  assign n10149 = n5933 & n5999 ;
  assign n10150 = ~n10148 & ~n10149 ;
  assign n10151 = \u10_mem_reg[0][24]/P0001  & ~n5928 ;
  assign n10152 = n5714 & n5928 ;
  assign n10153 = ~n10151 & ~n10152 ;
  assign n10154 = \u10_mem_reg[0][25]/P0001  & ~n5928 ;
  assign n10155 = n5718 & n5928 ;
  assign n10156 = ~n10154 & ~n10155 ;
  assign n10157 = \u10_mem_reg[0][26]/P0001  & ~n5928 ;
  assign n10158 = n5722 & n5928 ;
  assign n10159 = ~n10157 & ~n10158 ;
  assign n10160 = \u10_mem_reg[0][27]/P0001  & ~n5928 ;
  assign n10161 = n5726 & n5928 ;
  assign n10162 = ~n10160 & ~n10161 ;
  assign n10163 = \u10_mem_reg[0][28]/P0001  & ~n5928 ;
  assign n10164 = n5730 & n5928 ;
  assign n10165 = ~n10163 & ~n10164 ;
  assign n10166 = \u11_mem_reg[0][28]/P0001  & ~n5933 ;
  assign n10167 = n5933 & n5991 ;
  assign n10168 = ~n10166 & ~n10167 ;
  assign n10169 = \u10_mem_reg[0][30]/P0001  & ~n5928 ;
  assign n10170 = n5793 & n5928 ;
  assign n10171 = ~n10169 & ~n10170 ;
  assign n10172 = \u10_mem_reg[0][31]/P0001  & ~n5928 ;
  assign n10173 = n5797 & n5928 ;
  assign n10174 = ~n10172 & ~n10173 ;
  assign n10175 = \u10_mem_reg[0][29]/P0001  & ~n5928 ;
  assign n10176 = n5749 & n5928 ;
  assign n10177 = ~n10175 & ~n10176 ;
  assign n10178 = \u9_mem_reg[0][22]/P0001  & ~n5698 ;
  assign n10179 = n5698 & n5753 ;
  assign n10180 = ~n10178 & ~n10179 ;
  assign n10181 = \u2_bit_clk_r1_reg/P0001  & ~\u2_bit_clk_r_reg/P0001  ;
  assign n10182 = ~\u2_bit_clk_r1_reg/P0001  & \u2_bit_clk_r_reg/P0001  ;
  assign n10183 = ~n10181 & ~n10182 ;
  assign n10184 = ~\dma_ack_i[6]_pad  & \dma_req_o[6]_pad  ;
  assign n10185 = ~\dma_ack_i[6]_pad  & \u13_icc_r_reg[6]/NET0131  ;
  assign n10186 = n4429 & n10185 ;
  assign n10187 = \u16_u6_dma_req_r1_reg/P0001  & n10186 ;
  assign n10188 = ~n10184 & ~n10187 ;
  assign n10189 = ~\dma_ack_i[7]_pad  & \dma_req_o[7]_pad  ;
  assign n10190 = ~\dma_ack_i[7]_pad  & \u13_icc_r_reg[14]/NET0131  ;
  assign n10191 = n4462 & n10190 ;
  assign n10192 = \u16_u7_dma_req_r1_reg/P0001  & n10191 ;
  assign n10193 = ~n10189 & ~n10192 ;
  assign n10194 = ~\u2_sync_beat_reg/P0001  & ~\u2_sync_resume_reg/NET0131  ;
  assign n10195 = \u3_empty_reg/NET0131  & ~\valid_s_reg/NET0131  ;
  assign n10196 = \u14_u0_full_empty_r_reg/P0001  & \valid_s_reg/NET0131  ;
  assign n10197 = ~n10195 & ~n10196 ;
  assign n10198 = \u4_empty_reg/NET0131  & ~\valid_s_reg/NET0131  ;
  assign n10199 = \u14_u1_full_empty_r_reg/P0001  & \valid_s_reg/NET0131  ;
  assign n10200 = ~n10198 & ~n10199 ;
  assign n10201 = \u5_empty_reg/NET0131  & ~\valid_s_reg/NET0131  ;
  assign n10202 = \u14_u2_full_empty_r_reg/P0001  & \valid_s_reg/NET0131  ;
  assign n10203 = ~n10201 & ~n10202 ;
  assign n10204 = \u6_empty_reg/NET0131  & ~\valid_s_reg/NET0131  ;
  assign n10205 = \u14_u3_full_empty_r_reg/P0001  & \valid_s_reg/NET0131  ;
  assign n10206 = ~n10204 & ~n10205 ;
  assign n10207 = \u7_empty_reg/NET0131  & ~\valid_s_reg/NET0131  ;
  assign n10208 = \u14_u4_full_empty_r_reg/P0001  & \valid_s_reg/NET0131  ;
  assign n10209 = ~n10207 & ~n10208 ;
  assign n10210 = \u8_empty_reg/NET0131  & ~\valid_s_reg/NET0131  ;
  assign n10211 = \u14_u5_full_empty_r_reg/P0001  & \valid_s_reg/NET0131  ;
  assign n10212 = ~n10210 & ~n10211 ;
  assign n10213 = ~\in_valid_s_reg[0]/NET0131  & \u9_full_reg/NET0131  ;
  assign n10214 = \in_valid_s_reg[0]/NET0131  & \u14_u6_full_empty_r_reg/P0001  ;
  assign n10215 = ~n10213 & ~n10214 ;
  assign n10216 = ~\in_valid_s_reg[1]/NET0131  & \u10_full_reg/NET0131  ;
  assign n10217 = \in_valid_s_reg[1]/NET0131  & \u14_u7_full_empty_r_reg/P0001  ;
  assign n10218 = ~n10216 & ~n10217 ;
  assign n10219 = ~\in_valid_s_reg[2]/NET0131  & \u11_full_reg/NET0131  ;
  assign n10220 = \in_valid_s_reg[2]/NET0131  & \u14_u8_full_empty_r_reg/P0001  ;
  assign n10221 = ~n10219 & ~n10220 ;
  assign n10222 = \u1_sr_reg[11]/P0001  & \u2_out_le_reg[0]/P0001  ;
  assign n10223 = \u1_slt0_reg[11]/P0001  & ~\u2_out_le_reg[0]/P0001  ;
  assign n10224 = ~n10222 & ~n10223 ;
  assign n10225 = \u1_sr_reg[12]/P0001  & \u2_out_le_reg[0]/P0001  ;
  assign n10226 = \u1_slt0_reg[12]/P0001  & ~\u2_out_le_reg[0]/P0001  ;
  assign n10227 = ~n10225 & ~n10226 ;
  assign n10228 = \u1_sr_reg[15]/P0001  & \u2_out_le_reg[0]/P0001  ;
  assign n10229 = \u1_slt0_reg[15]/P0001  & ~\u2_out_le_reg[0]/P0001  ;
  assign n10230 = ~n10228 & ~n10229 ;
  assign n10231 = \u1_sr_reg[9]/P0001  & \u2_out_le_reg[0]/P0001  ;
  assign n10232 = \u1_slt0_reg[9]/P0001  & ~\u2_out_le_reg[0]/P0001  ;
  assign n10233 = ~n10231 & ~n10232 ;
  assign n10234 = \u1_sr_reg[10]/P0001  & \u2_out_le_reg[1]/P0001  ;
  assign n10235 = \u1_slt1_reg[10]/P0001  & ~\u2_out_le_reg[1]/P0001  ;
  assign n10236 = ~n10234 & ~n10235 ;
  assign n10237 = \u1_sr_reg[11]/P0001  & \u2_out_le_reg[1]/P0001  ;
  assign n10238 = \u1_slt1_reg[11]/P0001  & ~\u2_out_le_reg[1]/P0001  ;
  assign n10239 = ~n10237 & ~n10238 ;
  assign n10240 = \u1_sr_reg[5]/P0001  & \u2_out_le_reg[1]/P0001  ;
  assign n10241 = \u1_slt1_reg[5]/P0001  & ~\u2_out_le_reg[1]/P0001  ;
  assign n10242 = ~n10240 & ~n10241 ;
  assign n10243 = \u1_sr_reg[6]/P0001  & \u2_out_le_reg[1]/P0001  ;
  assign n10244 = \u1_slt1_reg[6]/P0001  & ~\u2_out_le_reg[1]/P0001  ;
  assign n10245 = ~n10243 & ~n10244 ;
  assign n10246 = \u1_sr_reg[7]/P0001  & \u2_out_le_reg[1]/P0001  ;
  assign n10247 = \u1_slt1_reg[7]/P0001  & ~\u2_out_le_reg[1]/P0001  ;
  assign n10248 = ~n10246 & ~n10247 ;
  assign n10249 = \u1_sr_reg[8]/P0001  & \u2_out_le_reg[1]/P0001  ;
  assign n10250 = \u1_slt1_reg[8]/P0001  & ~\u2_out_le_reg[1]/P0001  ;
  assign n10251 = ~n10249 & ~n10250 ;
  assign \_al_n1  = ~1'b0 ;
  assign \g16/_0_  = ~n2157 ;
  assign \g23/_0_  = n2168 ;
  assign \g29500/_0_  = n2178 ;
  assign \g29503/_3_  = ~n2181 ;
  assign \g29505/_3_  = n2183 ;
  assign \g29507/_3_  = ~n2186 ;
  assign \g29509/_3_  = ~n2189 ;
  assign \g29511/_0_  = n2190 ;
  assign \g29513/_3_  = ~n2193 ;
  assign \g29515/_3_  = ~n2196 ;
  assign \g29517/_3_  = ~n2199 ;
  assign \g29519/_0_  = ~n2202 ;
  assign \g29522/_0_  = n2203 ;
  assign \g29524/_0_  = n2204 ;
  assign \g29526/_0_  = n2205 ;
  assign \g29528/_0_  = n2206 ;
  assign \g29530/_0_  = n2207 ;
  assign \g29532/_0_  = n2208 ;
  assign \g29534/_3_  = ~n2211 ;
  assign \g29536/_3_  = ~n2214 ;
  assign \g29538/_3_  = ~n2217 ;
  assign \g29540/_3_  = ~n2220 ;
  assign \g29542/_3_  = ~n2223 ;
  assign \g29544/_3_  = ~n2226 ;
  assign \g29546/_3_  = ~n2229 ;
  assign \g29548/_3_  = ~n2232 ;
  assign \g29550/_0_  = n2233 ;
  assign \g29552/_0_  = n2234 ;
  assign \g29554/_0_  = n2235 ;
  assign \g29556/_0_  = n2236 ;
  assign \g29558/_0_  = n2237 ;
  assign \g29560/_0_  = n2238 ;
  assign \g29562/_0_  = n2239 ;
  assign \g29564/_0_  = n2240 ;
  assign \g29566/_0_  = n2241 ;
  assign \g29568/_0_  = n2242 ;
  assign \g29570/_0_  = n2243 ;
  assign \g29572/_0_  = n2244 ;
  assign \g29574/_3_  = ~n2247 ;
  assign \g29576/_3_  = ~n2250 ;
  assign \g29578/_3_  = ~n2253 ;
  assign \g29580/_3_  = ~n2256 ;
  assign \g29582/_3_  = ~n2259 ;
  assign \g29584/_3_  = ~n2262 ;
  assign \g29586/_3_  = ~n2265 ;
  assign \g29588/_3_  = ~n2268 ;
  assign \g29590/_3_  = ~n2271 ;
  assign \g29592/_3_  = ~n2274 ;
  assign \g29594/_3_  = ~n2277 ;
  assign \g29596/_3_  = ~n2280 ;
  assign \g29598/_3_  = ~n2283 ;
  assign \g29600/_3_  = ~n2286 ;
  assign \g29602/_3_  = ~n2289 ;
  assign \g29604/_3_  = ~n2292 ;
  assign \g29606/_0_  = n2293 ;
  assign \g29608/_0_  = n2294 ;
  assign \g29610/_0_  = n2295 ;
  assign \g29612/_0_  = n2296 ;
  assign \g29614/_3_  = ~n2299 ;
  assign \g29616/_3_  = ~n2302 ;
  assign \g29618/_3_  = ~n2305 ;
  assign \g29620/_3_  = ~n2308 ;
  assign \g29622/_3_  = ~n2311 ;
  assign \g29624/_3_  = ~n2314 ;
  assign \g29626/_3_  = ~n2317 ;
  assign \g29628/_3_  = ~n2320 ;
  assign \g29630/_3_  = ~n2323 ;
  assign \g29632/_3_  = ~n2326 ;
  assign \g29634/_3_  = ~n2329 ;
  assign \g29636/_3_  = ~n2332 ;
  assign \g29638/_3_  = ~n2335 ;
  assign \g29640/_3_  = ~n2338 ;
  assign \g29642/_3_  = ~n2341 ;
  assign \g29644/_3_  = ~n2344 ;
  assign \g29646/_3_  = ~n2347 ;
  assign \g29648/_3_  = ~n2350 ;
  assign \g29650/_3_  = ~n2353 ;
  assign \g29652/_3_  = ~n2356 ;
  assign \g29654/_3_  = ~n2359 ;
  assign \g29656/_3_  = ~n2362 ;
  assign \g29658/_3_  = ~n2365 ;
  assign \g29660/_3_  = ~n2368 ;
  assign \g29662/_3_  = ~n2371 ;
  assign \g29664/_3_  = ~n2374 ;
  assign \g29666/_3_  = ~n2377 ;
  assign \g29668/_3_  = ~n2380 ;
  assign \g29670/_3_  = ~n2383 ;
  assign \g29672/_3_  = ~n2386 ;
  assign \g29674/_3_  = ~n2389 ;
  assign \g29676/_3_  = ~n2392 ;
  assign \g29678/_3_  = ~n2395 ;
  assign \g29680/_3_  = ~n2398 ;
  assign \g29682/_3_  = ~n2401 ;
  assign \g29684/_3_  = ~n2404 ;
  assign \g29686/_3_  = ~n2407 ;
  assign \g29688/_3_  = ~n2410 ;
  assign \g29690/_3_  = ~n2413 ;
  assign \g29692/_3_  = ~n2416 ;
  assign \g29694/_0_  = n2417 ;
  assign \g29696/_0_  = n2418 ;
  assign \g29698/_0_  = n2419 ;
  assign \g29700/_0_  = n2420 ;
  assign \g29702/_0_  = n2421 ;
  assign \g29704/_0_  = n2422 ;
  assign \g29706/_0_  = n2423 ;
  assign \g29708/_0_  = n2424 ;
  assign \g29710/_0_  = n2425 ;
  assign \g29712/_0_  = n2426 ;
  assign \g29714/_0_  = n2427 ;
  assign \g29716/_0_  = n2428 ;
  assign \g29718/_0_  = n2429 ;
  assign \g29720/_0_  = n2430 ;
  assign \g29722/_0_  = n2431 ;
  assign \g29724/_0_  = n2432 ;
  assign \g29726/_0_  = n2433 ;
  assign \g29728/_0_  = n2434 ;
  assign \g29730/_0_  = n2435 ;
  assign \g29732/_0_  = n2436 ;
  assign \g29734/_3_  = ~n2439 ;
  assign \g29736/_3_  = ~n2442 ;
  assign \g29738/_3_  = ~n2445 ;
  assign \g29740/_3_  = ~n2448 ;
  assign \g29742/_3_  = ~n2451 ;
  assign \g29744/_3_  = ~n2454 ;
  assign \g29746/_3_  = ~n2457 ;
  assign \g29748/_3_  = ~n2460 ;
  assign \g29750/_3_  = ~n2463 ;
  assign \g29752/_3_  = ~n2466 ;
  assign \g29754/_3_  = ~n2469 ;
  assign \g29756/_3_  = ~n2472 ;
  assign \g29758/_3_  = ~n2475 ;
  assign \g29760/_3_  = ~n2478 ;
  assign \g29762/_3_  = ~n2481 ;
  assign \g29764/_3_  = ~n2484 ;
  assign \g29766/_3_  = ~n2487 ;
  assign \g29768/_3_  = ~n2490 ;
  assign \g29770/_3_  = ~n2493 ;
  assign \g29772/_3_  = ~n2496 ;
  assign \g29774/_3_  = ~n2499 ;
  assign \g29776/_3_  = ~n2502 ;
  assign \g29778/_3_  = ~n2505 ;
  assign \g29780/_3_  = ~n2508 ;
  assign \g29782/_3_  = ~n2511 ;
  assign \g29784/_3_  = ~n2514 ;
  assign \g29786/_3_  = ~n2517 ;
  assign \g29788/_3_  = ~n2520 ;
  assign \g29790/_3_  = ~n2523 ;
  assign \g29792/_3_  = ~n2526 ;
  assign \g29794/_3_  = ~n2529 ;
  assign \g29796/_3_  = ~n2532 ;
  assign \g29798/_3_  = ~n2535 ;
  assign \g29800/_3_  = ~n2538 ;
  assign \g29802/_3_  = ~n2541 ;
  assign \g29804/_3_  = ~n2544 ;
  assign \g29806/_3_  = ~n2547 ;
  assign \g29808/_3_  = ~n2550 ;
  assign \g29810/_3_  = ~n2553 ;
  assign \g29812/_3_  = ~n2556 ;
  assign \g29814/_3_  = ~n2559 ;
  assign \g29816/_3_  = ~n2562 ;
  assign \g29818/_3_  = ~n2565 ;
  assign \g29820/_3_  = ~n2568 ;
  assign \g29822/_3_  = ~n2571 ;
  assign \g29824/_3_  = ~n2574 ;
  assign \g29826/_3_  = ~n2577 ;
  assign \g29828/_3_  = ~n2580 ;
  assign \g29830/_3_  = ~n2583 ;
  assign \g29832/_3_  = ~n2586 ;
  assign \g29834/_3_  = ~n2589 ;
  assign \g29836/_3_  = ~n2592 ;
  assign \g29838/_3_  = ~n2595 ;
  assign \g29840/_3_  = ~n2598 ;
  assign \g29842/_3_  = ~n2601 ;
  assign \g29844/_3_  = ~n2604 ;
  assign \g29846/_3_  = ~n2607 ;
  assign \g29848/_3_  = ~n2610 ;
  assign \g29850/_3_  = ~n2613 ;
  assign \g29852/_3_  = ~n2616 ;
  assign \g29854/_3_  = ~n2619 ;
  assign \g29856/_3_  = ~n2622 ;
  assign \g29858/_3_  = ~n2625 ;
  assign \g29860/_3_  = ~n2628 ;
  assign \g29862/_3_  = ~n2631 ;
  assign \g29864/_3_  = ~n2634 ;
  assign \g29866/_3_  = ~n2637 ;
  assign \g29868/_3_  = ~n2640 ;
  assign \g29870/_3_  = ~n2643 ;
  assign \g29872/_3_  = ~n2646 ;
  assign \g29874/_3_  = ~n2649 ;
  assign \g29876/_3_  = ~n2652 ;
  assign \g29878/_3_  = ~n2655 ;
  assign \g29880/_3_  = ~n2658 ;
  assign \g29904/_0_  = ~n2670 ;
  assign \g29905/_0_  = ~n2682 ;
  assign \g29906/_0_  = ~n2694 ;
  assign \g29907/_0_  = ~n2706 ;
  assign \g29908/_0_  = ~n2718 ;
  assign \g29909/_0_  = ~n2730 ;
  assign \g29914/_3_  = ~n2733 ;
  assign \g29952/_0_  = n2744 ;
  assign \g29953/_0_  = n2746 ;
  assign \g29954/_0_  = n2748 ;
  assign \g29955/_0_  = n2750 ;
  assign \g29956/_0_  = n2752 ;
  assign \g29957/_0_  = n2754 ;
  assign \g29975/_0_  = n2668 ;
  assign \g29976/_0_  = n2680 ;
  assign \g29977/_0_  = n2692 ;
  assign \g29978/_0_  = n2704 ;
  assign \g29979/_0_  = n2716 ;
  assign \g29980/_0_  = n2728 ;
  assign \g29989/_3_  = ~n2757 ;
  assign \g30020/_0_  = n2768 ;
  assign \g30021/_0_  = n2779 ;
  assign \g30045/_0_  = n2783 ;
  assign \g30046/_0_  = n2793 ;
  assign \g30047/_0_  = n2804 ;
  assign \g30048/_0_  = n2814 ;
  assign \g30049/_0_  = n2666 ;
  assign \g30050/_0_  = n2678 ;
  assign \g30051/_0_  = n2690 ;
  assign \g30052/_0_  = n2702 ;
  assign \g30053/_0_  = n2714 ;
  assign \g30054/_0_  = n2726 ;
  assign \g30062/_0_  = n2818 ;
  assign \g30063/_0_  = n2822 ;
  assign \g30064/_0_  = n2824 ;
  assign \g30065/_0_  = n2826 ;
  assign \g30066/_0_  = n2828 ;
  assign \g30067/_0_  = n2832 ;
  assign \g30068/_0_  = n2836 ;
  assign \g30069/_0_  = n2840 ;
  assign \g30070/_0_  = n2843 ;
  assign \g30071/_0_  = n2846 ;
  assign \g30072/_0_  = n2849 ;
  assign \g30073/_0_  = n2852 ;
  assign \g30074/_0_  = n2855 ;
  assign \g30075/_0_  = n2858 ;
  assign \g30136/_3_  = ~n2861 ;
  assign \g30707/_0_  = n2867 ;
  assign \g30708/_0_  = n2872 ;
  assign \g30711/_0_  = n2877 ;
  assign \g30714/_0_  = n2882 ;
  assign \g30715/_0_  = n2887 ;
  assign \g30720/_0_  = n2892 ;
  assign \g30725/_0_  = n2897 ;
  assign \g30741/_0_  = ~n2914 ;
  assign \g30742/_0_  = ~n2924 ;
  assign \g30743/_0_  = ~n2941 ;
  assign \g30744/_0_  = ~n2951 ;
  assign \g30745/_0_  = ~n2968 ;
  assign \g30746/_0_  = ~n2978 ;
  assign \g30747/_0_  = ~n2996 ;
  assign \g30748/_0_  = ~n3006 ;
  assign \g30749/_0_  = ~n3024 ;
  assign \g30750/_0_  = ~n3041 ;
  assign \g30751/_0_  = ~n3051 ;
  assign \g30752/_0_  = ~n3061 ;
  assign \g30789/_0_  = n3071 ;
  assign \g30790/_0_  = n3112 ;
  assign \g30791/_0_  = n3152 ;
  assign \g30792/_0_  = n3178 ;
  assign \g30793/_0_  = n3204 ;
  assign \g30794/_0_  = n3230 ;
  assign \g30795/_0_  = n3256 ;
  assign \g30796/_0_  = n3282 ;
  assign \g30797/_0_  = n3308 ;
  assign \g30798/_0_  = n3318 ;
  assign \g30799/_0_  = n3344 ;
  assign \g30800/_0_  = n3370 ;
  assign \g30801/_0_  = n3384 ;
  assign \g30802/_0_  = n3398 ;
  assign \g30803/_0_  = n3417 ;
  assign \g30804/_0_  = n3436 ;
  assign \g30805/_0_  = n3448 ;
  assign \g30806/_0_  = n3460 ;
  assign \g30807/_0_  = n3479 ;
  assign \g30808/_0_  = n3498 ;
  assign \g30809/_0_  = n3508 ;
  assign \g30810/_0_  = n3549 ;
  assign \g30811/_0_  = n3589 ;
  assign \g30812/_0_  = n3615 ;
  assign \g30813/_0_  = n3641 ;
  assign \g30814/_0_  = n3667 ;
  assign \g30815/_0_  = n3693 ;
  assign \g30816/_0_  = n3719 ;
  assign \g30817/_0_  = n3745 ;
  assign \g30818/_0_  = n3771 ;
  assign \g30819/_0_  = n3797 ;
  assign \g30820/_0_  = n3811 ;
  assign \g30821/_0_  = n3825 ;
  assign \g30822/_0_  = n3844 ;
  assign \g30823/_0_  = n3863 ;
  assign \g30824/_0_  = n3875 ;
  assign \g30825/_0_  = n3887 ;
  assign \g30826/_0_  = n3906 ;
  assign \g30827/_0_  = n3925 ;
  assign \g30828/_0_  = n3966 ;
  assign \g30829/_0_  = n4006 ;
  assign \g30830/_0_  = n4032 ;
  assign \g30831/_0_  = n4058 ;
  assign \g30832/_0_  = n4084 ;
  assign \g30833/_0_  = n4110 ;
  assign \g30834/_0_  = n4136 ;
  assign \g30835/_0_  = n4162 ;
  assign \g30836/_0_  = n4188 ;
  assign \g30837/_0_  = n4214 ;
  assign \g30838/_0_  = n4228 ;
  assign \g30839/_0_  = n4242 ;
  assign \g30840/_0_  = n4261 ;
  assign \g30841/_0_  = n4280 ;
  assign \g30842/_0_  = n4292 ;
  assign \g30843/_0_  = n4304 ;
  assign \g30844/_0_  = n4323 ;
  assign \g30845/_0_  = n4342 ;
  assign \g30846/_0_  = n4383 ;
  assign \g30847/_0_  = n4422 ;
  assign \g30848/_0_  = n4429 ;
  assign \g30849/_0_  = n4455 ;
  assign \g30850/_0_  = n4462 ;
  assign \g30851/_0_  = n4488 ;
  assign \g30852/_0_  = n4514 ;
  assign \g30853/_0_  = n2153 ;
  assign \g30854/_0_  = n4539 ;
  assign \g30855/_0_  = n4565 ;
  assign \g30856/_0_  = n4591 ;
  assign \g30857/_0_  = n4617 ;
  assign \g30858/_0_  = n4643 ;
  assign \g30859/_0_  = n4657 ;
  assign \g30860/_0_  = n4671 ;
  assign \g30861/_0_  = n4690 ;
  assign \g30862/_0_  = n4709 ;
  assign \g30863/_0_  = n4721 ;
  assign \g30864/_0_  = n4733 ;
  assign \g30865/_0_  = n4752 ;
  assign \g30866/_0_  = n4771 ;
  assign \g30867/_0_  = n4812 ;
  assign \g30868/_0_  = n4852 ;
  assign \g30869/_0_  = n4878 ;
  assign \g30870/_0_  = n4903 ;
  assign \g30871/_0_  = n4929 ;
  assign \g30872/_0_  = n4955 ;
  assign \g30873/_0_  = n4981 ;
  assign \g30874/_0_  = n5006 ;
  assign \g30875/_0_  = n5032 ;
  assign \g30876/_0_  = n5073 ;
  assign \g30877/_0_  = n5099 ;
  assign \g30878/_0_  = n5139 ;
  assign \g30879/_0_  = n5165 ;
  assign \g30880/_0_  = n5179 ;
  assign \g30881/_0_  = n5205 ;
  assign \g30882/_0_  = n5219 ;
  assign \g30883/_0_  = n5245 ;
  assign \g30884/_0_  = n5264 ;
  assign \g30885/_0_  = n5290 ;
  assign \g30886/_0_  = n5309 ;
  assign \g30887/_0_  = n5335 ;
  assign \g30888/_0_  = n5361 ;
  assign \g30889/_0_  = n5373 ;
  assign \g30890/_0_  = n5385 ;
  assign \g30891/_0_  = n5411 ;
  assign \g30892/_0_  = n5430 ;
  assign \g30893/_0_  = n5456 ;
  assign \g30894/_0_  = n5475 ;
  assign \g30895/_0_  = n5489 ;
  assign \g30896/_0_  = n5503 ;
  assign \g30897/_0_  = n5522 ;
  assign \g30898/_0_  = n5541 ;
  assign \g30899/_0_  = n5553 ;
  assign \g30900/_0_  = n5565 ;
  assign \g30901/_0_  = n5584 ;
  assign \g30902/_0_  = n5603 ;
  assign \g30906/_0_  = n5606 ;
  assign \g30907/_0_  = n5609 ;
  assign \g30908/_0_  = n5612 ;
  assign \g30909/_0_  = n5616 ;
  assign \g30910/_0_  = n5620 ;
  assign \g30911/_0_  = n5624 ;
  assign \g30918/_0_  = n5631 ;
  assign \g30919/_0_  = n5634 ;
  assign \g30920/_0_  = n5639 ;
  assign \g30921/_0_  = n5643 ;
  assign \g30922/_0_  = n5647 ;
  assign \g30923/_0_  = n5651 ;
  assign \g30924/_0_  = n5656 ;
  assign \g30925/_0_  = n5661 ;
  assign \g30926/_0_  = n5666 ;
  assign \g30946/_0_  = ~n5675 ;
  assign \g30947/_0_  = ~n5681 ;
  assign \g30948/_0_  = ~n5685 ;
  assign \g30949/_0_  = ~n5689 ;
  assign \g30950/_0_  = ~n5693 ;
  assign \g30951/_0_  = ~n5697 ;
  assign \g30952/_0_  = ~n5706 ;
  assign \g30953/_0_  = ~n5712 ;
  assign \g30954/_0_  = ~n5716 ;
  assign \g30955/_0_  = ~n5720 ;
  assign \g30956/_0_  = ~n5724 ;
  assign \g30957/_0_  = ~n5728 ;
  assign \g30958/_0_  = ~n5732 ;
  assign \g30959/_0_  = ~n5736 ;
  assign \g30960/_0_  = ~n5739 ;
  assign \g30961/_0_  = ~n5743 ;
  assign \g30962/_0_  = ~n5747 ;
  assign \g30963/_0_  = ~n5751 ;
  assign \g30964/_0_  = ~n5755 ;
  assign \g30965/_0_  = ~n5759 ;
  assign \g30966/_0_  = ~n5763 ;
  assign \g30967/_0_  = ~n5767 ;
  assign \g30968/_0_  = ~n5771 ;
  assign \g30969/_0_  = ~n5775 ;
  assign \g30970/_0_  = ~n5779 ;
  assign \g30971/_0_  = ~n5783 ;
  assign \g30972/_0_  = ~n5787 ;
  assign \g30973/_0_  = ~n5791 ;
  assign \g30974/_0_  = ~n5795 ;
  assign \g30975/_0_  = ~n5799 ;
  assign \g30976/_0_  = ~n5804 ;
  assign \g30977/_0_  = ~n5807 ;
  assign \g30978/_0_  = ~n5810 ;
  assign \g30979/_0_  = ~n5813 ;
  assign \g30980/_0_  = ~n5816 ;
  assign \g30981/_0_  = ~n5819 ;
  assign \g30982/_0_  = ~n5822 ;
  assign \g30983/_0_  = ~n5825 ;
  assign \g30984/_0_  = ~n5828 ;
  assign \g30985/_0_  = ~n5831 ;
  assign \g30986/_0_  = ~n5834 ;
  assign \g30987/_0_  = ~n5837 ;
  assign \g30988/_0_  = ~n5840 ;
  assign \g30989/_0_  = ~n5843 ;
  assign \g30990/_0_  = ~n5846 ;
  assign \g30991/_0_  = ~n5849 ;
  assign \g30992/_0_  = ~n5852 ;
  assign \g30993/_0_  = ~n5855 ;
  assign \g30994/_0_  = ~n5858 ;
  assign \g30995/_0_  = ~n5861 ;
  assign \g30996/_0_  = ~n5864 ;
  assign \g30997/_0_  = ~n5867 ;
  assign \g30998/_0_  = ~n5870 ;
  assign \g30999/_0_  = ~n5873 ;
  assign \g31000/_0_  = ~n5876 ;
  assign \g31001/_0_  = ~n5879 ;
  assign \g31002/_0_  = ~n5882 ;
  assign \g31003/_0_  = ~n5885 ;
  assign \g31004/_0_  = ~n5888 ;
  assign \g31005/_0_  = ~n5891 ;
  assign \g31006/_0_  = ~n5894 ;
  assign \g31007/_0_  = ~n5897 ;
  assign \g31008/_0_  = ~n5900 ;
  assign \g31009/_0_  = ~n5903 ;
  assign \g31010/_0_  = ~n5906 ;
  assign \g31011/_0_  = ~n5909 ;
  assign \g31012/_0_  = ~n5912 ;
  assign \g31013/_0_  = ~n5915 ;
  assign \g31014/_0_  = ~n5918 ;
  assign \g31015/_0_  = ~n5921 ;
  assign \g31016/_0_  = ~n5924 ;
  assign \g31017/_0_  = ~n5927 ;
  assign \g31018/_0_  = ~n5932 ;
  assign \g31019/_0_  = ~n5941 ;
  assign \g31020/_0_  = ~n5947 ;
  assign \g31021/_0_  = ~n5950 ;
  assign \g31022/_0_  = ~n5954 ;
  assign \g31023/_0_  = ~n5957 ;
  assign \g31024/_0_  = ~n5961 ;
  assign \g31025/_0_  = ~n5965 ;
  assign \g31026/_0_  = ~n5969 ;
  assign \g31027/_0_  = ~n5973 ;
  assign \g31028/_0_  = ~n5977 ;
  assign \g31029/_0_  = ~n5981 ;
  assign \g31030/_0_  = ~n5985 ;
  assign \g31031/_0_  = ~n5989 ;
  assign \g31032/_0_  = ~n5993 ;
  assign \g31033/_0_  = ~n5997 ;
  assign \g31034/_0_  = ~n6001 ;
  assign \g31035/_0_  = ~n6005 ;
  assign \g31036/_0_  = ~n6010 ;
  assign \g31037/_0_  = ~n6013 ;
  assign \g31038/_0_  = ~n6016 ;
  assign \g31039/_0_  = ~n6019 ;
  assign \g31040/_0_  = ~n6022 ;
  assign \g31041/_0_  = ~n6025 ;
  assign \g31042/_0_  = ~n6028 ;
  assign \g31043/_0_  = ~n6031 ;
  assign \g31044/_0_  = ~n6035 ;
  assign \g31045/_0_  = ~n6038 ;
  assign \g31046/_0_  = ~n6041 ;
  assign \g31047/_0_  = ~n6044 ;
  assign \g31048/_0_  = ~n6047 ;
  assign \g31049/_0_  = ~n6050 ;
  assign \g31050/_0_  = ~n6053 ;
  assign \g31051/_0_  = ~n6056 ;
  assign \g31052/_0_  = ~n6059 ;
  assign \g31053/_0_  = ~n6062 ;
  assign \g31054/_0_  = ~n6065 ;
  assign \g31055/_0_  = ~n6068 ;
  assign \g31056/_0_  = ~n6071 ;
  assign \g31057/_0_  = ~n6074 ;
  assign \g31058/_0_  = ~n6077 ;
  assign \g31059/_0_  = ~n6080 ;
  assign \g31060/_0_  = ~n6083 ;
  assign \g31061/_0_  = ~n6086 ;
  assign \g31062/_0_  = ~n6089 ;
  assign \g31063/_0_  = ~n6092 ;
  assign \g31064/_0_  = ~n6095 ;
  assign \g31065/_0_  = ~n6098 ;
  assign \g31066/_0_  = ~n6101 ;
  assign \g31067/_0_  = ~n6104 ;
  assign \g31068/_0_  = ~n6107 ;
  assign \g31069/_0_  = ~n6110 ;
  assign \g31070/_0_  = ~n6113 ;
  assign \g31071/_0_  = ~n6116 ;
  assign \g31072/_0_  = ~n6119 ;
  assign \g31073/_0_  = ~n6122 ;
  assign \g31074/_0_  = ~n6125 ;
  assign \g31075/_0_  = ~n6128 ;
  assign \g31076/_0_  = ~n6131 ;
  assign \g31077/_0_  = ~n6134 ;
  assign \g31084/u3_syn_4  = n3068 ;
  assign \g31085/u3_syn_4  = n5668 ;
  assign \g31096/u3_syn_4  = n5733 ;
  assign \g31115/u3_syn_4  = n5801 ;
  assign \g31136/u3_syn_4  = n3315 ;
  assign \g31158/u3_syn_4  = n3505 ;
  assign \g31176/u3_syn_4  = n5951 ;
  assign \g31193/u3_syn_4  = n6032 ;
  assign \g31195/u3_syn_4  = n6007 ;
  assign \g31247/u3_syn_4  = n5699 ;
  assign \g31280/u3_syn_4  = n5929 ;
  assign \g31285/u3_syn_4  = n5934 ;
  assign \g31568/_0_  = n6138 ;
  assign \g31631/_0_  = ~n6175 ;
  assign \g31672/_0_  = n6182 ;
  assign \g31731/_0_  = n6186 ;
  assign \g31732/_0_  = n6190 ;
  assign \g31742/_2_  = ~n6192 ;
  assign \g31744/_2_  = ~n6194 ;
  assign \g31746/_2_  = ~n6196 ;
  assign \g31748/_2_  = ~n6198 ;
  assign \g31751/_2_  = ~n6200 ;
  assign \g31754/_2_  = ~n6202 ;
  assign \g31756/_2_  = ~n6204 ;
  assign \g31758/_2_  = ~n6206 ;
  assign \g31760/_2_  = ~n6208 ;
  assign \g31761/_0_  = n6210 ;
  assign \g31789/_0_  = ~n6213 ;
  assign \g31807/_3_  = ~n6218 ;
  assign \g31825/_3_  = ~n6221 ;
  assign \g32607/_0_  = ~n6234 ;
  assign \g32608/_0_  = ~n6247 ;
  assign \g32609/_0_  = ~n6260 ;
  assign \g32610/_0_  = ~n6273 ;
  assign \g32611/_0_  = ~n6286 ;
  assign \g32612/_0_  = ~n6299 ;
  assign \g32613/_0_  = n6305 ;
  assign \g32614/_0_  = n6311 ;
  assign \g32615/_0_  = n6317 ;
  assign \g32616/_0_  = n6323 ;
  assign \g32617/_0_  = n6329 ;
  assign \g32618/_0_  = n6335 ;
  assign \g32645/_0__syn_2  = n6336 ;
  assign \g32687/_0__syn_2  = n6337 ;
  assign \g32749/_0__syn_2  = n6338 ;
  assign \g32757/_0_  = ~n6346 ;
  assign \g32758/_0_  = ~n6353 ;
  assign \g32759/_0_  = ~n6360 ;
  assign \g32760/_0_  = ~n6367 ;
  assign \g32761/_0_  = ~n6374 ;
  assign \g32762/_0_  = ~n6381 ;
  assign \g32763/_0_  = ~n6388 ;
  assign \g32764/_0_  = ~n6395 ;
  assign \g32765/_0_  = ~n6402 ;
  assign \g32769/_0_  = n6406 ;
  assign \g32835/_1_  = n3313 ;
  assign \g32839/_0_  = n6410 ;
  assign \g32844/_0_  = n6414 ;
  assign \g32901/_1_  = n3503 ;
  assign \g32902/_0_  = n6418 ;
  assign \g32963/_1_  = n3066 ;
  assign \g32972/_0_  = n6422 ;
  assign \g32977/_0_  = n6426 ;
  assign \g32979/_0_  = n6429 ;
  assign \g32980/_0_  = n6432 ;
  assign \g32981/_0_  = n6435 ;
  assign \g32982/_0_  = n6438 ;
  assign \g32983/_0_  = n6441 ;
  assign \g32987/_0_  = n6444 ;
  assign \g33018/_0_  = n6446 ;
  assign \g33019/_0_  = ~n6450 ;
  assign \g33088/_0_  = ~n6453 ;
  assign \g33261/_0_  = n6460 ;
  assign \g33264/_0_  = n6462 ;
  assign \g33275/_0_  = n6463 ;
  assign \g33276/_0_  = n6467 ;
  assign \g33277/_0_  = n6468 ;
  assign \g33371/_0_  = ~n6478 ;
  assign \g33382/_0_  = n6484 ;
  assign \g33401/_0_  = ~n6488 ;
  assign \g33402/_0_  = ~n6492 ;
  assign \g33403/_0_  = ~n6495 ;
  assign \g33404/_0_  = ~n6498 ;
  assign \g33405/_0_  = ~n6501 ;
  assign \g33406/_0_  = ~n6504 ;
  assign \g33407/_0_  = ~n6507 ;
  assign \g33408/_0_  = ~n6510 ;
  assign \g33409/_0_  = ~n6513 ;
  assign \g33410/_0_  = ~n6516 ;
  assign \g33411/_0_  = ~n6519 ;
  assign \g33412/_0_  = ~n6522 ;
  assign \g33413/_0_  = ~n6525 ;
  assign \g33414/_0_  = ~n6528 ;
  assign \g33415/_0_  = ~n6531 ;
  assign \g33416/_0_  = ~n6534 ;
  assign \g33417/_0_  = ~n6537 ;
  assign \g33418/_0_  = ~n6540 ;
  assign \g33419/_0_  = ~n6543 ;
  assign \g33420/_0_  = ~n6546 ;
  assign \g33421/_0_  = ~n6549 ;
  assign \g33422/_0_  = ~n6552 ;
  assign \g33423/_0_  = ~n6555 ;
  assign \g33424/_0_  = ~n6558 ;
  assign \g33425/_0_  = ~n6561 ;
  assign \g33426/_0_  = ~n6564 ;
  assign \g33427/_0_  = ~n6567 ;
  assign \g33428/_0_  = ~n6570 ;
  assign \g33429/_0_  = ~n6573 ;
  assign \g33430/_0_  = ~n6576 ;
  assign \g33431/_0_  = ~n6579 ;
  assign \g33432/_0_  = ~n6582 ;
  assign \g33433/_0_  = ~n6586 ;
  assign \g33434/_0_  = ~n6589 ;
  assign \g33435/_0_  = ~n6592 ;
  assign \g33436/_0_  = ~n6595 ;
  assign \g33437/_0_  = ~n6598 ;
  assign \g33438/_0_  = ~n6601 ;
  assign \g33439/_0_  = ~n6604 ;
  assign \g33440/_0_  = ~n6607 ;
  assign \g33441/_0_  = ~n6610 ;
  assign \g33442/_0_  = ~n6613 ;
  assign \g33443/_0_  = ~n6616 ;
  assign \g33444/_0_  = ~n6619 ;
  assign \g33445/_0_  = ~n6622 ;
  assign \g33446/_0_  = ~n6625 ;
  assign \g33447/_0_  = ~n6628 ;
  assign \g33448/_0_  = ~n6632 ;
  assign \g33449/_0_  = ~n6635 ;
  assign \g33450/_0_  = ~n6638 ;
  assign \g33451/_0_  = ~n6641 ;
  assign \g33452/_0_  = ~n6644 ;
  assign \g33453/_0_  = ~n6647 ;
  assign \g33454/_0_  = ~n6650 ;
  assign \g33455/_0_  = ~n6653 ;
  assign \g33456/_0_  = ~n6656 ;
  assign \g33457/_0_  = ~n6659 ;
  assign \g33458/_0_  = ~n6662 ;
  assign \g33459/_0_  = ~n6665 ;
  assign \g33460/_0_  = ~n6668 ;
  assign \g33461/_0_  = ~n6671 ;
  assign \g33462/_0_  = ~n6674 ;
  assign \g33463/_0_  = ~n6677 ;
  assign \g33464/_0_  = ~n6680 ;
  assign \g33465/_0_  = ~n6683 ;
  assign \g33466/_0_  = ~n6686 ;
  assign \g33467/_0_  = ~n6689 ;
  assign \g33468/_0_  = ~n6692 ;
  assign \g33469/_0_  = ~n6695 ;
  assign \g33470/_0_  = ~n6698 ;
  assign \g33471/_0_  = ~n6701 ;
  assign \g33472/_0_  = ~n6704 ;
  assign \g33473/_0_  = ~n6707 ;
  assign \g33474/_0_  = ~n6710 ;
  assign \g33475/_0_  = ~n6713 ;
  assign \g33476/_0_  = ~n6716 ;
  assign \g33477/_0_  = ~n6719 ;
  assign \g33478/_0_  = ~n6722 ;
  assign \g33479/_0_  = ~n6725 ;
  assign \g33480/_0_  = ~n6728 ;
  assign \g33481/_0_  = ~n6731 ;
  assign \g33482/_0_  = ~n6734 ;
  assign \g33483/_0_  = ~n6737 ;
  assign \g33484/_0_  = ~n6740 ;
  assign \g33485/_0_  = ~n6743 ;
  assign \g33486/_0_  = ~n6746 ;
  assign \g33487/_0_  = ~n6749 ;
  assign \g33488/_0_  = ~n6752 ;
  assign \g33489/_0_  = ~n6755 ;
  assign \g33490/_0_  = ~n6758 ;
  assign \g33491/_0_  = ~n6761 ;
  assign \g33492/_0_  = ~n6764 ;
  assign \g33493/_0_  = ~n6767 ;
  assign \g33494/_0_  = ~n6770 ;
  assign \g33495/_0_  = ~n6773 ;
  assign \g33496/_0_  = ~n6776 ;
  assign \g33497/_0_  = ~n6779 ;
  assign \g33498/_0_  = ~n6782 ;
  assign \g33499/_0_  = ~n6785 ;
  assign \g33500/_0_  = ~n6788 ;
  assign \g33501/_0_  = ~n6791 ;
  assign \g33502/_0_  = ~n6794 ;
  assign \g33503/_0_  = ~n6797 ;
  assign \g33504/_0_  = ~n6800 ;
  assign \g33505/_0_  = ~n6803 ;
  assign \g33506/_0_  = ~n6806 ;
  assign \g33507/_0_  = ~n6810 ;
  assign \g33508/_0_  = ~n6813 ;
  assign \g33509/_0_  = ~n6816 ;
  assign \g33510/_0_  = ~n6819 ;
  assign \g33511/_0_  = ~n6822 ;
  assign \g33512/_0_  = ~n6825 ;
  assign \g33513/_0_  = ~n6828 ;
  assign \g33514/_0_  = ~n6831 ;
  assign \g33515/_0_  = ~n6834 ;
  assign \g33516/_0_  = ~n6837 ;
  assign \g33517/_0_  = ~n6840 ;
  assign \g33518/_0_  = ~n6843 ;
  assign \g33519/_0_  = ~n6846 ;
  assign \g33520/_0_  = ~n6849 ;
  assign \g33521/_0_  = ~n6852 ;
  assign \g33522/_0_  = ~n6855 ;
  assign \g33523/_0_  = ~n6858 ;
  assign \g33524/_0_  = ~n6861 ;
  assign \g33525/_0_  = ~n6864 ;
  assign \g33526/_0_  = ~n6867 ;
  assign \g33527/_0_  = ~n6870 ;
  assign \g33528/_0_  = ~n6873 ;
  assign \g33529/_0_  = ~n6876 ;
  assign \g33530/_0_  = ~n6879 ;
  assign \g33531/_0_  = ~n6882 ;
  assign \g33532/_0_  = ~n6885 ;
  assign \g33533/_0_  = ~n6888 ;
  assign \g33534/_0_  = ~n6891 ;
  assign \g33535/_0_  = ~n6894 ;
  assign \g33536/_0_  = ~n6897 ;
  assign \g33537/_0_  = ~n6900 ;
  assign \g33538/_0_  = ~n6903 ;
  assign \g33539/_0_  = ~n6907 ;
  assign \g33540/_0_  = ~n6910 ;
  assign \g33541/_0_  = ~n6913 ;
  assign \g33542/_0_  = ~n6916 ;
  assign \g33543/_0_  = ~n6919 ;
  assign \g33544/_0_  = ~n6922 ;
  assign \g33545/_0_  = ~n6925 ;
  assign \g33546/_0_  = ~n6928 ;
  assign \g33547/_0_  = ~n6931 ;
  assign \g33548/_0_  = ~n6934 ;
  assign \g33549/_0_  = ~n6937 ;
  assign \g33550/_0_  = ~n6940 ;
  assign \g33551/_0_  = ~n6943 ;
  assign \g33552/_0_  = ~n6946 ;
  assign \g33553/_0_  = ~n6949 ;
  assign \g33554/_0_  = ~n6952 ;
  assign \g33555/_0_  = ~n6955 ;
  assign \g33556/_0_  = ~n6958 ;
  assign \g33557/_0_  = ~n6961 ;
  assign \g33558/_0_  = ~n6964 ;
  assign \g33559/_0_  = ~n6967 ;
  assign \g33560/_0_  = ~n6970 ;
  assign \g33561/_0_  = ~n6973 ;
  assign \g33562/_0_  = ~n6976 ;
  assign \g33563/_0_  = ~n6979 ;
  assign \g33564/_0_  = ~n6982 ;
  assign \g33565/_0_  = ~n6985 ;
  assign \g33566/_0_  = ~n6988 ;
  assign \g33567/_0_  = ~n6991 ;
  assign \g33568/_0_  = ~n6994 ;
  assign \g33569/_0_  = ~n6997 ;
  assign \g33570/_0_  = ~n7000 ;
  assign \g33571/_0_  = ~n7003 ;
  assign \g33572/_0_  = ~n7006 ;
  assign \g33573/_0_  = ~n7009 ;
  assign \g33574/_0_  = ~n7012 ;
  assign \g33575/_0_  = ~n7015 ;
  assign \g33576/_0_  = ~n7018 ;
  assign \g33577/_0_  = ~n7021 ;
  assign \g33578/_0_  = ~n7024 ;
  assign \g33579/_0_  = ~n7027 ;
  assign \g33580/_0_  = ~n7030 ;
  assign \g33581/_0_  = ~n7033 ;
  assign \g33582/_0_  = ~n7036 ;
  assign \g33583/_0_  = ~n7039 ;
  assign \g33584/_0_  = ~n7042 ;
  assign \g33585/_0_  = ~n7045 ;
  assign \g33586/_0_  = ~n7048 ;
  assign \g33587/_0_  = ~n7051 ;
  assign \g33588/_0_  = ~n7054 ;
  assign \g33589/_0_  = ~n7057 ;
  assign \g33590/_0_  = ~n7060 ;
  assign \g33591/_0_  = ~n7063 ;
  assign \g33592/_0_  = ~n7066 ;
  assign \g33593/_0_  = ~n7069 ;
  assign \g33594/_0_  = ~n7072 ;
  assign \g33595/_0_  = ~n7075 ;
  assign \g33596/_0_  = ~n7078 ;
  assign \g33597/_0_  = ~n7081 ;
  assign \g33598/_0_  = ~n7084 ;
  assign \g33599/_0_  = ~n7087 ;
  assign \g33600/_0_  = ~n7090 ;
  assign \g33601/_0_  = ~n7093 ;
  assign \g33602/_0_  = ~n7096 ;
  assign \g33603/_0_  = ~n7099 ;
  assign \g33604/_0_  = ~n7103 ;
  assign \g33605/_0_  = ~n7106 ;
  assign \g33606/_0_  = ~n7109 ;
  assign \g33607/_0_  = ~n7112 ;
  assign \g33608/_0_  = ~n7115 ;
  assign \g33609/_0_  = ~n7118 ;
  assign \g33610/_0_  = ~n7121 ;
  assign \g33611/_0_  = ~n7124 ;
  assign \g33612/_0_  = ~n7127 ;
  assign \g33613/_0_  = ~n7130 ;
  assign \g33614/_0_  = ~n7133 ;
  assign \g33615/_0_  = ~n7136 ;
  assign \g33616/_0_  = ~n7139 ;
  assign \g33617/_0_  = ~n7142 ;
  assign \g33618/_0_  = ~n7145 ;
  assign \g33619/_0_  = ~n7148 ;
  assign \g33620/_0_  = ~n7151 ;
  assign \g33621/_0_  = ~n7154 ;
  assign \g33622/_0_  = ~n7157 ;
  assign \g33623/_0_  = ~n7160 ;
  assign \g33624/_0_  = ~n7163 ;
  assign \g33625/_0_  = ~n7166 ;
  assign \g33626/_0_  = ~n7169 ;
  assign \g33627/_0_  = ~n7172 ;
  assign \g33628/_0_  = ~n7175 ;
  assign \g33629/_0_  = ~n7178 ;
  assign \g33630/_0_  = ~n7181 ;
  assign \g33631/_0_  = ~n7184 ;
  assign \g33632/_0_  = ~n7187 ;
  assign \g33633/_0_  = ~n7190 ;
  assign \g33634/_0_  = ~n7193 ;
  assign \g33635/_0_  = ~n7196 ;
  assign \g33636/_0_  = ~n7200 ;
  assign \g33637/_0_  = ~n7203 ;
  assign \g33638/_0_  = ~n7206 ;
  assign \g33639/_0_  = ~n7209 ;
  assign \g33640/_0_  = ~n7212 ;
  assign \g33641/_0_  = ~n7215 ;
  assign \g33642/_0_  = ~n7218 ;
  assign \g33643/_0_  = ~n7221 ;
  assign \g33644/_0_  = ~n7224 ;
  assign \g33645/_0_  = ~n7227 ;
  assign \g33646/_0_  = ~n7230 ;
  assign \g33647/_0_  = ~n7233 ;
  assign \g33648/_0_  = ~n7236 ;
  assign \g33649/_0_  = ~n7239 ;
  assign \g33650/_0_  = ~n7242 ;
  assign \g33651/_0_  = ~n7245 ;
  assign \g33652/_0_  = ~n7248 ;
  assign \g33653/_0_  = ~n7251 ;
  assign \g33654/_0_  = ~n7254 ;
  assign \g33655/_0_  = ~n7257 ;
  assign \g33656/_0_  = ~n7260 ;
  assign \g33657/_0_  = ~n7263 ;
  assign \g33658/_0_  = ~n7266 ;
  assign \g33659/_0_  = ~n7269 ;
  assign \g33660/_0_  = ~n7272 ;
  assign \g33661/_0_  = ~n7275 ;
  assign \g33662/_0_  = ~n7278 ;
  assign \g33663/_0_  = ~n7281 ;
  assign \g33664/_0_  = ~n7284 ;
  assign \g33665/_0_  = ~n7287 ;
  assign \g33666/_0_  = ~n7290 ;
  assign \g33667/_0_  = ~n7293 ;
  assign \g33668/_0_  = ~n7296 ;
  assign \g33669/_0_  = ~n7299 ;
  assign \g33670/_0_  = ~n7302 ;
  assign \g33671/_0_  = ~n7305 ;
  assign \g33672/_0_  = ~n7308 ;
  assign \g33673/_0_  = ~n7311 ;
  assign \g33674/_0_  = ~n7314 ;
  assign \g33675/_0_  = ~n7317 ;
  assign \g33676/_0_  = ~n7320 ;
  assign \g33677/_0_  = ~n7323 ;
  assign \g33678/_0_  = ~n7326 ;
  assign \g33679/_0_  = ~n7329 ;
  assign \g33680/_0_  = ~n7332 ;
  assign \g33681/_0_  = ~n7335 ;
  assign \g33682/_0_  = ~n7338 ;
  assign \g33683/_0_  = ~n7341 ;
  assign \g33684/_0_  = ~n7344 ;
  assign \g33685/_0_  = ~n7347 ;
  assign \g33686/_0_  = ~n7350 ;
  assign \g33687/_0_  = ~n7353 ;
  assign \g33688/_0_  = ~n7356 ;
  assign \g33689/_0_  = ~n7359 ;
  assign \g33690/_0_  = ~n7362 ;
  assign \g33691/_0_  = ~n7365 ;
  assign \g33692/_0_  = ~n7368 ;
  assign \g33693/_0_  = ~n7371 ;
  assign \g33694/_0_  = ~n7374 ;
  assign \g33695/_0_  = ~n7377 ;
  assign \g33696/_0_  = ~n7380 ;
  assign \g33697/_0_  = ~n7383 ;
  assign \g33698/_0_  = ~n7386 ;
  assign \g33699/_0_  = ~n7389 ;
  assign \g33700/_0_  = ~n7392 ;
  assign \g33701/_0_  = ~n7395 ;
  assign \g33702/_0_  = ~n7398 ;
  assign \g33703/_0_  = ~n7401 ;
  assign \g33704/_0_  = ~n7405 ;
  assign \g33705/_0_  = ~n7408 ;
  assign \g33706/_0_  = ~n7411 ;
  assign \g33707/_0_  = ~n7414 ;
  assign \g33708/_0_  = ~n7417 ;
  assign \g33709/_0_  = ~n7420 ;
  assign \g33710/_0_  = ~n7423 ;
  assign \g33711/_0_  = ~n7426 ;
  assign \g33712/_0_  = ~n7429 ;
  assign \g33713/_0_  = ~n7432 ;
  assign \g33714/_0_  = ~n7435 ;
  assign \g33715/_0_  = ~n7438 ;
  assign \g33716/_0_  = ~n7441 ;
  assign \g33717/_0_  = ~n7444 ;
  assign \g33718/_0_  = ~n7447 ;
  assign \g33719/_0_  = ~n7450 ;
  assign \g33720/_0_  = ~n7453 ;
  assign \g33721/_0_  = ~n7456 ;
  assign \g33722/_0_  = ~n7459 ;
  assign \g33723/_0_  = ~n7462 ;
  assign \g33724/_0_  = ~n7465 ;
  assign \g33725/_0_  = ~n7468 ;
  assign \g33726/_0_  = ~n7471 ;
  assign \g33727/_0_  = ~n7474 ;
  assign \g33728/_0_  = ~n7477 ;
  assign \g33729/_0_  = ~n7480 ;
  assign \g33730/_0_  = ~n7483 ;
  assign \g33731/_0_  = ~n7486 ;
  assign \g33732/_0_  = ~n7489 ;
  assign \g33733/_0_  = ~n7492 ;
  assign \g33734/_0_  = ~n7495 ;
  assign \g33735/_0_  = ~n7498 ;
  assign \g33736/_0_  = ~n7502 ;
  assign \g33737/_0_  = ~n7505 ;
  assign \g33738/_0_  = ~n7508 ;
  assign \g33739/_0_  = ~n7511 ;
  assign \g33740/_0_  = ~n7514 ;
  assign \g33741/_0_  = ~n7517 ;
  assign \g33742/_0_  = ~n7520 ;
  assign \g33743/_0_  = ~n7523 ;
  assign \g33744/_0_  = ~n7526 ;
  assign \g33745/_0_  = ~n7529 ;
  assign \g33746/_0_  = ~n7532 ;
  assign \g33747/_0_  = ~n7535 ;
  assign \g33748/_0_  = ~n7538 ;
  assign \g33749/_0_  = ~n7541 ;
  assign \g33750/_0_  = ~n7544 ;
  assign \g33751/_0_  = ~n7547 ;
  assign \g33752/_0_  = ~n7550 ;
  assign \g33753/_0_  = ~n7553 ;
  assign \g33754/_0_  = ~n7556 ;
  assign \g33755/_0_  = ~n7559 ;
  assign \g33756/_0_  = ~n7562 ;
  assign \g33757/_0_  = ~n7565 ;
  assign \g33758/_0_  = ~n7568 ;
  assign \g33759/_0_  = ~n7571 ;
  assign \g33760/_0_  = ~n7574 ;
  assign \g33761/_0_  = ~n7577 ;
  assign \g33762/_0_  = ~n7580 ;
  assign \g33763/_0_  = ~n7583 ;
  assign \g33764/_0_  = ~n7586 ;
  assign \g33765/_0_  = ~n7589 ;
  assign \g33766/_0_  = ~n7592 ;
  assign \g33767/_0_  = ~n7595 ;
  assign \g33768/_0_  = ~n7598 ;
  assign \g33769/_0_  = ~n7601 ;
  assign \g33770/_0_  = ~n7604 ;
  assign \g33771/_0_  = ~n7607 ;
  assign \g33772/_0_  = ~n7610 ;
  assign \g33773/_0_  = ~n7613 ;
  assign \g33774/_0_  = ~n7616 ;
  assign \g33775/_0_  = ~n7619 ;
  assign \g33776/_0_  = ~n7622 ;
  assign \g33777/_0_  = ~n7625 ;
  assign \g33778/_0_  = ~n7628 ;
  assign \g33779/_0_  = ~n7631 ;
  assign \g33780/_0_  = ~n7634 ;
  assign \g33781/_0_  = ~n7637 ;
  assign \g33782/_0_  = ~n7640 ;
  assign \g33783/_0_  = ~n7643 ;
  assign \g33784/_0_  = ~n7646 ;
  assign \g33785/_0_  = ~n7649 ;
  assign \g33786/_0_  = ~n7652 ;
  assign \g33787/_0_  = ~n7655 ;
  assign \g33788/_0_  = ~n7658 ;
  assign \g33789/_0_  = ~n7661 ;
  assign \g33790/_0_  = ~n7664 ;
  assign \g33791/_0_  = ~n7667 ;
  assign \g33792/_0_  = ~n7670 ;
  assign \g33793/_0_  = ~n7673 ;
  assign \g33794/_0_  = ~n7676 ;
  assign \g33795/_0_  = ~n7679 ;
  assign \g33796/_0_  = ~n7682 ;
  assign \g33797/_0_  = ~n7685 ;
  assign \g33798/_0_  = ~n7688 ;
  assign \g33799/_0_  = ~n7691 ;
  assign \g33800/_0_  = ~n7694 ;
  assign \g33801/_0_  = ~n7697 ;
  assign \g33802/_0_  = ~n7700 ;
  assign \g33803/_0_  = ~n7703 ;
  assign \g33804/_0_  = ~n7706 ;
  assign \g33805/_0_  = ~n7709 ;
  assign \g33806/_0_  = ~n7713 ;
  assign \g33807/_0_  = ~n7716 ;
  assign \g33808/_0_  = ~n7719 ;
  assign \g33809/_0_  = ~n7722 ;
  assign \g33810/_0_  = ~n7725 ;
  assign \g33811/_0_  = ~n7728 ;
  assign \g33812/_0_  = ~n7731 ;
  assign \g33813/_0_  = ~n7734 ;
  assign \g33814/_0_  = ~n7737 ;
  assign \g33815/_0_  = ~n7740 ;
  assign \g33816/_0_  = ~n7743 ;
  assign \g33817/_0_  = ~n7746 ;
  assign \g33818/_0_  = ~n7749 ;
  assign \g33819/_0_  = ~n7752 ;
  assign \g33820/_0_  = ~n7755 ;
  assign \g33821/_0_  = ~n7758 ;
  assign \g33822/_0_  = ~n7761 ;
  assign \g33823/_0_  = ~n7764 ;
  assign \g33824/_0_  = ~n7767 ;
  assign \g33825/_0_  = ~n7770 ;
  assign \g33826/_0_  = ~n7773 ;
  assign \g33827/_0_  = ~n7776 ;
  assign \g33828/_0_  = ~n7779 ;
  assign \g33829/_0_  = ~n7782 ;
  assign \g33830/_0_  = ~n7785 ;
  assign \g33831/_0_  = ~n7788 ;
  assign \g33832/_0_  = ~n7791 ;
  assign \g33833/_0_  = ~n7794 ;
  assign \g33834/_0_  = ~n7797 ;
  assign \g33835/_0_  = ~n7800 ;
  assign \g33836/_0_  = ~n7803 ;
  assign \g33837/_0_  = ~n7806 ;
  assign \g33838/_0_  = ~n7809 ;
  assign \g33839/_0_  = ~n7812 ;
  assign \g33840/_0_  = ~n7816 ;
  assign \g33841/_0_  = ~n7819 ;
  assign \g33842/_0_  = ~n7822 ;
  assign \g33843/_0_  = ~n7825 ;
  assign \g33844/_0_  = ~n7828 ;
  assign \g33845/_0_  = ~n7831 ;
  assign \g33846/_0_  = ~n7834 ;
  assign \g33847/_0_  = ~n7837 ;
  assign \g33848/_0_  = ~n7840 ;
  assign \g33849/_0_  = ~n7843 ;
  assign \g33850/_0_  = ~n7846 ;
  assign \g33851/_0_  = ~n7849 ;
  assign \g33852/_0_  = ~n7852 ;
  assign \g33853/_0_  = ~n7855 ;
  assign \g33854/_0_  = ~n7858 ;
  assign \g33855/_0_  = ~n7861 ;
  assign \g33856/_0_  = ~n7864 ;
  assign \g33857/_0_  = ~n7867 ;
  assign \g33858/_0_  = ~n7870 ;
  assign \g33859/_0_  = ~n7873 ;
  assign \g33860/_0_  = ~n7876 ;
  assign \g33861/_0_  = ~n7879 ;
  assign \g33862/_0_  = ~n7882 ;
  assign \g33863/_0_  = ~n7885 ;
  assign \g33864/_0_  = ~n7888 ;
  assign \g33865/_0_  = ~n7891 ;
  assign \g33866/_0_  = ~n7894 ;
  assign \g33867/_0_  = ~n7897 ;
  assign \g33868/_0_  = ~n7900 ;
  assign \g33869/_0_  = ~n7903 ;
  assign \g33870/_0_  = ~n7906 ;
  assign \g33871/_0_  = ~n7909 ;
  assign \g33872/_0_  = ~n7912 ;
  assign \g33873/_0_  = ~n7915 ;
  assign \g33874/_0_  = ~n7918 ;
  assign \g33875/_0_  = ~n7921 ;
  assign \g33876/_0_  = ~n7924 ;
  assign \g33877/_0_  = ~n7927 ;
  assign \g33878/_0_  = ~n7930 ;
  assign \g33879/_0_  = ~n7933 ;
  assign \g33880/_0_  = ~n7936 ;
  assign \g33881/_0_  = ~n7939 ;
  assign \g33882/_0_  = ~n7942 ;
  assign \g33883/_0_  = ~n7945 ;
  assign \g33884/_0_  = ~n7948 ;
  assign \g33885/_0_  = ~n7951 ;
  assign \g33886/_0_  = ~n7954 ;
  assign \g33887/_0_  = ~n7957 ;
  assign \g33888/_0_  = ~n7960 ;
  assign \g33889/_0_  = ~n7963 ;
  assign \g33890/_0_  = ~n7966 ;
  assign \g33891/_0_  = ~n7969 ;
  assign \g33892/_0_  = ~n7972 ;
  assign \g33893/_0_  = ~n7975 ;
  assign \g33894/_0_  = ~n7978 ;
  assign \g33895/_0_  = ~n7981 ;
  assign \g33896/_0_  = ~n7984 ;
  assign \g33897/_0_  = ~n7987 ;
  assign \g33898/_0_  = ~n7990 ;
  assign \g33899/_0_  = ~n7993 ;
  assign \g33900/_0_  = ~n7996 ;
  assign \g33901/_0_  = ~n7999 ;
  assign \g33902/_0_  = ~n8002 ;
  assign \g33903/_0_  = ~n8005 ;
  assign \g33904/_0_  = ~n8008 ;
  assign \g33905/_0_  = ~n8011 ;
  assign \g33906/_0_  = ~n8014 ;
  assign \g33907/_0_  = ~n8017 ;
  assign \g33908/_0_  = ~n8020 ;
  assign \g33909/_0_  = ~n8023 ;
  assign \g33910/_0_  = ~n8026 ;
  assign \g33911/_0_  = ~n8029 ;
  assign \g33912/_0_  = ~n8032 ;
  assign \g33913/_0_  = ~n8035 ;
  assign \g33914/_0_  = ~n8038 ;
  assign \g33915/_0_  = ~n8041 ;
  assign \g33916/_0_  = ~n8044 ;
  assign \g33917/_0_  = ~n8047 ;
  assign \g33918/_0_  = ~n8050 ;
  assign \g33919/_0_  = ~n8053 ;
  assign \g33920/_0_  = ~n8056 ;
  assign \g33921/_0_  = ~n8059 ;
  assign \g33922/_0_  = ~n8062 ;
  assign \g33923/_0_  = ~n8065 ;
  assign \g33924/_0_  = ~n8068 ;
  assign \g33925/_0_  = ~n8071 ;
  assign \g33926/_0_  = ~n8074 ;
  assign \g33927/_0_  = ~n8077 ;
  assign \g33928/_0_  = ~n8080 ;
  assign \g33929/_0_  = ~n8083 ;
  assign \g33930/_0_  = ~n8086 ;
  assign \g33931/_0_  = ~n8089 ;
  assign \g33932/_0_  = ~n8092 ;
  assign \g33933/_0_  = ~n8095 ;
  assign \g33934/_0_  = ~n8098 ;
  assign \g33935/_0_  = ~n8101 ;
  assign \g33936/_0_  = ~n8104 ;
  assign \g33937/_0_  = ~n8107 ;
  assign \g33938/_0_  = ~n8110 ;
  assign \g33939/_0_  = ~n8113 ;
  assign \g33940/_0_  = ~n8116 ;
  assign \g33941/_0_  = ~n8119 ;
  assign \g33942/_0_  = ~n8122 ;
  assign \g33943/_0_  = ~n8125 ;
  assign \g33944/_0_  = ~n8128 ;
  assign \g33945/_0_  = ~n8131 ;
  assign \g33946/_0_  = ~n8134 ;
  assign \g33947/_0_  = ~n8137 ;
  assign \g33948/_0_  = ~n8140 ;
  assign \g33949/_0_  = ~n8143 ;
  assign \g33950/_0_  = ~n8146 ;
  assign \g33951/_0_  = ~n8149 ;
  assign \g33952/_0_  = ~n8152 ;
  assign \g33953/_0_  = ~n8155 ;
  assign \g33954/_0_  = ~n8158 ;
  assign \g33955/_0_  = ~n8161 ;
  assign \g33956/_0_  = ~n8164 ;
  assign \g33957/_0_  = ~n8167 ;
  assign \g33958/_0_  = ~n8170 ;
  assign \g33959/_0_  = ~n8173 ;
  assign \g33960/_0_  = ~n8176 ;
  assign \g33961/_0_  = ~n8179 ;
  assign \g33962/_0_  = ~n8182 ;
  assign \g33963/_0_  = ~n8185 ;
  assign \g33964/_0_  = ~n8188 ;
  assign \g33965/_0_  = ~n8191 ;
  assign \g33966/_0_  = ~n8194 ;
  assign \g33967/_0_  = ~n8197 ;
  assign \g33968/_0_  = ~n8200 ;
  assign \g33969/_0_  = ~n8203 ;
  assign \g33970/_0_  = ~n8206 ;
  assign \g33971/_0_  = ~n8209 ;
  assign \g33972/_0_  = ~n8212 ;
  assign \g33973/_0_  = ~n8215 ;
  assign \g33974/_0_  = ~n8218 ;
  assign \g33975/_0_  = ~n8221 ;
  assign \g33976/_0_  = ~n8224 ;
  assign \g33977/u3_syn_4  = n8225 ;
  assign \g33981/u3_syn_4  = n8226 ;
  assign \g34014/u3_syn_4  = n8227 ;
  assign \g34047/u3_syn_4  = n8228 ;
  assign \g34084/u3_syn_4  = n8229 ;
  assign \g34123/u3_syn_4  = n8230 ;
  assign \g34306/_0_  = ~n8248 ;
  assign \g34316/_0_  = ~n8266 ;
  assign \g34324/_0_  = ~n8284 ;
  assign \g34326/_0_  = ~n8302 ;
  assign \g34328/_0_  = ~n8320 ;
  assign \g34331/_0_  = ~n8338 ;
  assign \g34333/_0_  = ~n8356 ;
  assign \g34344/_0_  = ~n8374 ;
  assign \g34347/_0_  = ~n8392 ;
  assign \g34351/_0_  = ~n8410 ;
  assign \g34361/_0_  = ~n8428 ;
  assign \g34368/_0_  = ~n8446 ;
  assign \g34377/_0_  = ~n8464 ;
  assign \g34385/_0_  = ~n8482 ;
  assign \g34393/_0_  = ~n8500 ;
  assign \g34414/_1_  = n8501 ;
  assign \g34451/_1_  = n8502 ;
  assign \g34476/_1_  = n8503 ;
  assign \g34487/_0_  = n8504 ;
  assign \g34490/_1_  = n8505 ;
  assign \g34715/_0_  = ~n8508 ;
  assign \g34878/_0_  = n8520 ;
  assign \g34882/_0_  = n8532 ;
  assign \g34883/_0_  = n8534 ;
  assign \g34893/_0_  = n8546 ;
  assign \g34896/_0_  = n8561 ;
  assign \g34898/_0_  = n8576 ;
  assign \g34899/_0_  = n8588 ;
  assign \g34916/_3_  = ~n8591 ;
  assign \g35264/_0_  = n8596 ;
  assign \g35265/_0_  = n8601 ;
  assign \g35266/_0_  = n8606 ;
  assign \g35267/_0_  = n8610 ;
  assign \g35268/_0_  = n8614 ;
  assign \g35269/_0_  = n8618 ;
  assign \g35270/_0_  = n8621 ;
  assign \g35271/_0_  = n8624 ;
  assign \g35272/_0_  = ~n8640 ;
  assign \g35273/_0_  = ~n8656 ;
  assign \g35274/_0_  = ~n8672 ;
  assign \g35275/_0_  = n8675 ;
  assign \g35276/_0_  = ~n8691 ;
  assign \g35277/_0_  = ~n8707 ;
  assign \g35278/_0_  = ~n8723 ;
  assign \g35279/_0_  = ~n8737 ;
  assign \g35283/_0_  = n8740 ;
  assign \g35287/_0_  = n3062 ;
  assign \g35294/_0_  = n6339 ;
  assign \g35300/_0_  = n2758 ;
  assign \g35304/_0_  = n2769 ;
  assign \g35308/_0_  = n2794 ;
  assign \g35312/_0_  = n2807 ;
  assign \g35316/_0_  = n2158 ;
  assign \g35318/_0_  = n3309 ;
  assign \g35326/_0_  = ~n8756 ;
  assign \g35334/_0_  = n3499 ;
  assign \g35336/_0_  = n8760 ;
  assign \g35337/_0_  = n8764 ;
  assign \g35338/_0_  = n8767 ;
  assign \g35357/_0_  = ~n8769 ;
  assign \g35358/_0_  = ~n8771 ;
  assign \g35359/_0_  = ~n8773 ;
  assign \g35419/_0_  = n8776 ;
  assign \g35438/_0_  = n8781 ;
  assign \g35439/_0_  = n8782 ;
  assign \g35440/_0_  = n8783 ;
  assign \g35441/_0_  = n8784 ;
  assign \g35442/_0_  = n8785 ;
  assign \g35444/_0_  = ~n8797 ;
  assign \g35445/_0_  = ~n8809 ;
  assign \g35446/_0_  = ~n8821 ;
  assign \g35447/_0_  = ~n8833 ;
  assign \g35448/_0_  = ~n8845 ;
  assign \g35449/_0_  = ~n8852 ;
  assign \g35450/_0_  = ~n8859 ;
  assign \g35451/_0_  = ~n8868 ;
  assign \g35452/_0_  = n8871 ;
  assign \g35463/_0_  = ~n8874 ;
  assign \g35464/_0_  = ~n8931 ;
  assign \g35466/_0_  = n8932 ;
  assign \g35485/_2_  = n8935 ;
  assign \g35495/_0_  = n8937 ;
  assign \g35496/_0_  = ~n8939 ;
  assign \g35499/_0_  = ~n8941 ;
  assign \g35500/_0_  = ~n8943 ;
  assign \g35501/_0_  = n8945 ;
  assign \g35502/_0_  = ~n8947 ;
  assign \g35563/_0_  = n8948 ;
  assign \g35633/_0_  = n8949 ;
  assign \g35717/_0_  = n8956 ;
  assign \g35718/_0_  = n8963 ;
  assign \g35719/_0_  = n8970 ;
  assign \g35809/_0_  = n8972 ;
  assign \g35810/_0_  = n8974 ;
  assign \g35811/_0_  = n8976 ;
  assign \g35812/_0_  = n8978 ;
  assign \g35813/_0_  = n8980 ;
  assign \g35814/_0_  = n8982 ;
  assign \g35815/_0_  = n8984 ;
  assign \g35816/_0_  = n8986 ;
  assign \g35817/_0_  = n8988 ;
  assign \g35818/_0_  = n8990 ;
  assign \g35819/_0_  = n8992 ;
  assign \g35820/_0_  = n8994 ;
  assign \g35821/_0_  = n8996 ;
  assign \g35822/_0_  = n8998 ;
  assign \g35823/_0_  = n9000 ;
  assign \g35824/_0_  = n9002 ;
  assign \g35825/_0_  = n9004 ;
  assign \g35826/_0_  = n9006 ;
  assign \g35827/_0_  = n9008 ;
  assign \g35830/_0_  = n9016 ;
  assign \g35833/_0_  = n9020 ;
  assign \g35835/_0_  = n9027 ;
  assign \g35836/_0_  = n9035 ;
  assign \g35837/_0_  = n9043 ;
  assign \g35839/_0_  = ~n9047 ;
  assign \g35840/_0_  = ~n9050 ;
  assign \g35841/_0_  = n9057 ;
  assign \g35843/_0_  = n9059 ;
  assign \g35844/_0_  = n9066 ;
  assign \g35845/_0_  = n9070 ;
  assign \g35853/_0_  = n9071 ;
  assign \g35854/_0_  = n9072 ;
  assign \g35855/_0_  = n9076 ;
  assign \g35856/_0_  = n9077 ;
  assign \g36306/_0_  = ~n9082 ;
  assign \g36414/_0_  = n9083 ;
  assign \g36415/_0_  = n9084 ;
  assign \g36449/_0_  = ~n9088 ;
  assign \g36550/_0_  = ~n9089 ;
  assign \g36551/_0_  = ~n9092 ;
  assign \g36553/_0_  = ~n9095 ;
  assign \g36560/_0_  = n9097 ;
  assign \g36562/_3_  = n9099 ;
  assign \g36563/_0_  = n9103 ;
  assign \g36612/_0_  = n9104 ;
  assign \g36614/_2_  = ~n9108 ;
  assign \g36695/_0_  = n9111 ;
  assign \g36784/_0_  = ~n9122 ;
  assign \g36785/_0_  = ~n9129 ;
  assign \g36786/_0_  = ~n9136 ;
  assign \g36787/_0_  = ~n9143 ;
  assign \g36788/_0_  = ~n9150 ;
  assign \g36789/_0_  = ~n9157 ;
  assign \g36790/_0_  = ~n9164 ;
  assign \g36791/_0_  = ~n9171 ;
  assign \g36792/_0_  = ~n9178 ;
  assign \g36793/_0_  = ~n9185 ;
  assign \g36794/_0_  = ~n9192 ;
  assign \g36796/_0_  = ~n9199 ;
  assign \g36797/_0_  = ~n9206 ;
  assign \g36798/_0_  = ~n9213 ;
  assign \g36799/_0_  = ~n9220 ;
  assign \g36800/_0_  = ~n9227 ;
  assign \g36801/_0_  = ~n9234 ;
  assign \g36802/_0_  = ~n9241 ;
  assign \g36803/_0_  = ~n9248 ;
  assign \g36804/_0_  = ~n9255 ;
  assign \g36805/_0_  = ~n9262 ;
  assign \g36806/_0_  = ~n9269 ;
  assign \g36807/_0_  = ~n9276 ;
  assign \g36808/_0_  = ~n9283 ;
  assign \g36809/_0_  = ~n9290 ;
  assign \g36810/_0_  = ~n9297 ;
  assign \g36811/_0_  = ~n9304 ;
  assign \g36813/_0_  = ~n9311 ;
  assign \g36814/_0_  = ~n9322 ;
  assign \g36815/_0_  = ~n9329 ;
  assign \g36820/_0_  = ~n9336 ;
  assign \g36825/_0_  = ~n9343 ;
  assign \g36832/_0_  = ~n9350 ;
  assign \g36846/_0_  = ~n9357 ;
  assign \g36855/_0_  = ~n9364 ;
  assign \g36857/_0_  = ~n9371 ;
  assign \g36859/_0_  = ~n9378 ;
  assign \g36860/_0_  = ~n9385 ;
  assign \g36861/_0_  = ~n9392 ;
  assign \g36862/_0_  = ~n9403 ;
  assign \g36863/_0_  = ~n9410 ;
  assign \g36864/_0_  = ~n9417 ;
  assign \g36867/_0_  = ~n9424 ;
  assign \g36870/_0_  = ~n9431 ;
  assign \g36871/_0_  = ~n9438 ;
  assign \g36877/_0_  = ~n9445 ;
  assign \g36879/_0_  = ~n9452 ;
  assign \g36892/_0_  = ~n9459 ;
  assign \g36893/_0_  = ~n9466 ;
  assign \g36901/_0_  = ~n9473 ;
  assign \g36909/_0_  = ~n9480 ;
  assign \g36914/_0_  = ~n9487 ;
  assign \g36919/_0_  = ~n9494 ;
  assign \g36922/_0_  = ~n9501 ;
  assign \g36923/_0_  = ~n9508 ;
  assign \g36927/_0_  = ~n9515 ;
  assign \g36930/_0_  = ~n9522 ;
  assign \g36931/_0_  = ~n9529 ;
  assign \g36933/_0_  = ~n9536 ;
  assign \g36934/_0_  = ~n9543 ;
  assign \g36935/_0_  = ~n9550 ;
  assign \g36936/_0_  = ~n9557 ;
  assign \g36937/_0_  = ~n9564 ;
  assign \g36938/_0_  = ~n9571 ;
  assign \g36939/_0_  = ~n9578 ;
  assign \g36940/_0_  = ~n9585 ;
  assign \g36941/_0_  = ~n9592 ;
  assign \g36943/_0_  = ~n9599 ;
  assign \g36944/_0_  = ~n9606 ;
  assign \g36945/_0_  = ~n9613 ;
  assign \g36946/_0_  = ~n9620 ;
  assign \g36947/_0_  = ~n9627 ;
  assign \g36948/_0_  = ~n9634 ;
  assign \g36949/_0_  = ~n9641 ;
  assign \g36950/_0_  = ~n9648 ;
  assign \g36951/_0_  = ~n9655 ;
  assign \g36952/_0_  = ~n9662 ;
  assign \g36953/_0_  = ~n9669 ;
  assign \g36954/_0_  = ~n9676 ;
  assign \g36957/_0_  = ~n9683 ;
  assign \g36958/_0_  = ~n9690 ;
  assign \g36959/_0_  = ~n9697 ;
  assign \g36960/_0_  = ~n9704 ;
  assign \g36961/_0_  = ~n9711 ;
  assign \g36962/_0_  = ~n9718 ;
  assign \g36963/_0_  = ~n9725 ;
  assign \g36970/_0_  = ~n9732 ;
  assign \g36977/_0_  = ~n9739 ;
  assign \g36986/_0_  = ~n9746 ;
  assign \g36991/_0_  = ~n9753 ;
  assign \g36994/_0_  = ~n9760 ;
  assign \g37015/_0_  = ~n9767 ;
  assign \g37057/_0_  = ~n9774 ;
  assign \g37073/_0_  = ~n9781 ;
  assign \g37128/_0_  = ~n9788 ;
  assign \g37129/_0_  = ~n9795 ;
  assign \g37138/_0_  = ~n9801 ;
  assign \g37139/_0_  = n9802 ;
  assign \g37140/_0_  = ~n9808 ;
  assign \g37141/_0_  = ~n9813 ;
  assign \g37142/_0_  = ~n9818 ;
  assign \g37143/_0_  = ~n9823 ;
  assign \g37144/_0_  = ~n9828 ;
  assign \g37145/_0_  = ~n9833 ;
  assign \g37146/_0_  = ~n9838 ;
  assign \g37147/_0_  = ~n9843 ;
  assign \g37148/_0_  = ~n9848 ;
  assign \g37149/_0_  = ~n9853 ;
  assign \g37150/_0_  = ~n9858 ;
  assign \g37151/_0_  = ~n9863 ;
  assign \g37152/_0_  = ~n9868 ;
  assign \g37153/_0_  = ~n9874 ;
  assign \g37154/_0_  = ~n9879 ;
  assign \g37155/_0_  = ~n9884 ;
  assign \g37156/_0_  = ~n9889 ;
  assign \g37157/_0_  = ~n9894 ;
  assign \g37158/_0_  = ~n9899 ;
  assign \g37159/_0_  = ~n9904 ;
  assign \g37160/_0_  = ~n9909 ;
  assign \g37161/_0_  = ~n9914 ;
  assign \g37162/_0_  = ~n9919 ;
  assign \g37163/_0_  = ~n9924 ;
  assign \g37164/_0_  = ~n9929 ;
  assign \g37165/_0_  = ~n9934 ;
  assign \g37166/_0_  = ~n9939 ;
  assign \g37167/_0_  = ~n9944 ;
  assign \g37168/_0_  = ~n9949 ;
  assign \g37169/_0_  = ~n9954 ;
  assign \g37170/_0_  = ~n9959 ;
  assign \g37171/_0_  = ~n9964 ;
  assign \g37172/_0_  = ~n9969 ;
  assign \g37173/_0_  = ~n9974 ;
  assign \g37174/_0_  = ~n9979 ;
  assign \g37175/_0_  = ~n9984 ;
  assign \g37176/_0_  = ~n9989 ;
  assign \g37177/_0_  = ~n9994 ;
  assign \g37178/_0_  = ~n9999 ;
  assign \g37179/_0_  = ~n10004 ;
  assign \g37180/_0_  = ~n10009 ;
  assign \g37181/_0_  = ~n10014 ;
  assign \g37182/_0_  = ~n10019 ;
  assign \g37183/_0_  = ~n10024 ;
  assign \g37184/_0_  = ~n10029 ;
  assign \g37185/_0_  = ~n10034 ;
  assign \g37187/_0_  = ~n10039 ;
  assign \g37188/_0_  = ~n10044 ;
  assign \g37190/_0_  = ~n10049 ;
  assign \g37191/_0_  = ~n10054 ;
  assign \g37192/_0_  = ~n10059 ;
  assign \g37193/_0_  = ~n10064 ;
  assign \g37194/_0_  = ~n10069 ;
  assign \g37372/_3_  = n10072 ;
  assign \g37377/_0_  = ~n10075 ;
  assign \g37378/_0_  = ~n10078 ;
  assign \g37379/_0_  = ~n10081 ;
  assign \g37380/_0_  = ~n10084 ;
  assign \g37381/_0_  = ~n10087 ;
  assign \g37382/_0_  = ~n10090 ;
  assign \g37383/_0_  = ~n10093 ;
  assign \g37384/_0_  = ~n10096 ;
  assign \g37385/_0_  = ~n10099 ;
  assign \g37386/_0_  = ~n10102 ;
  assign \g37387/_0_  = ~n10105 ;
  assign \g37388/_0_  = ~n10108 ;
  assign \g37389/_0_  = ~n10111 ;
  assign \g37390/_0_  = ~n10114 ;
  assign \g37391/_0_  = ~n10117 ;
  assign \g37392/_0_  = ~n10120 ;
  assign \g37393/_0_  = ~n10123 ;
  assign \g37394/_0_  = ~n10126 ;
  assign \g37395/_0_  = ~n10129 ;
  assign \g37396/_0_  = ~n10132 ;
  assign \g37397/_0_  = ~n10135 ;
  assign \g37398/_0_  = ~n10138 ;
  assign \g37399/_0_  = ~n10141 ;
  assign \g37400/_0_  = ~n10144 ;
  assign \g37401/_0_  = ~n10147 ;
  assign \g37402/_0_  = ~n10150 ;
  assign \g37403/_0_  = ~n10153 ;
  assign \g37404/_0_  = ~n10156 ;
  assign \g37405/_0_  = ~n10159 ;
  assign \g37406/_0_  = ~n10162 ;
  assign \g37407/_0_  = ~n10165 ;
  assign \g37408/_0_  = ~n10168 ;
  assign \g37409/_0_  = ~n10171 ;
  assign \g37410/_0_  = ~n10174 ;
  assign \g37411/_0_  = ~n10177 ;
  assign \g37412/_0_  = ~n10180 ;
  assign \g37413/_0_  = ~n10183 ;
  assign \g37576/_3_  = n9064 ;
  assign \g37590/_2_  = n2738 ;
  assign \g40278/_0_  = n8778 ;
  assign \g40379/_0_  = n8521 ;
  assign \g40389/_2_  = n9013 ;
  assign \g40390/_2_  = n9032 ;
  assign \g40391/_0_  = n6289 ;
  assign \g40393/_2_  = n9040 ;
  assign \g40395/_0_  = n8551 ;
  assign \g40397/_0_  = n8509 ;
  assign \g40400/_0_  = n6263 ;
  assign \g40402/_0_  = n8566 ;
  assign \g45458/_0_  = n2155 ;
  assign \g45675/_0_  = ~n10188 ;
  assign \g45677/_0_  = n10186 ;
  assign \g45678/_0_  = ~n10193 ;
  assign \g45682/_0_  = n10191 ;
  assign sync_pad_o_pad = ~n10194 ;
  assign \u14_u0_full_empty_r_reg/P0001_reg_syn_3  = ~n10197 ;
  assign \u14_u1_full_empty_r_reg/P0001_reg_syn_3  = ~n10200 ;
  assign \u14_u2_full_empty_r_reg/P0001_reg_syn_3  = ~n10203 ;
  assign \u14_u3_full_empty_r_reg/P0001_reg_syn_3  = ~n10206 ;
  assign \u14_u4_full_empty_r_reg/P0001_reg_syn_3  = ~n10209 ;
  assign \u14_u5_full_empty_r_reg/P0001_reg_syn_3  = ~n10212 ;
  assign \u14_u6_full_empty_r_reg/P0001_reg_syn_3  = ~n10215 ;
  assign \u14_u7_full_empty_r_reg/P0001_reg_syn_3  = ~n10218 ;
  assign \u14_u8_full_empty_r_reg/P0001_reg_syn_3  = ~n10221 ;
  assign \u1_slt0_reg[11]/P0001_reg_syn_3  = ~n10224 ;
  assign \u1_slt0_reg[12]/P0001_reg_syn_3  = ~n10227 ;
  assign \u1_slt0_reg[15]/P0001_reg_syn_3  = ~n10230 ;
  assign \u1_slt0_reg[9]/P0001_reg_syn_3  = ~n10233 ;
  assign \u1_slt1_reg[10]/P0001_reg_syn_3  = ~n10236 ;
  assign \u1_slt1_reg[11]/P0001_reg_syn_3  = ~n10239 ;
  assign \u1_slt1_reg[5]/P0001_reg_syn_3  = ~n10242 ;
  assign \u1_slt1_reg[6]/P0001_reg_syn_3  = ~n10245 ;
  assign \u1_slt1_reg[7]/P0001_reg_syn_3  = ~n10248 ;
  assign \u1_slt1_reg[8]/P0001_reg_syn_3  = ~n10251 ;
  assign wb_err_o_pad = 1'b0 ;
endmodule
