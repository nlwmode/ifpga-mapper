module top (\a[0] , \a[1] , \a[2] , \a[3] , \a[4] , \a[5] , \a[6] , \a[7] , \a[8] , \a[9] , \a[10] , \a[11] , \a[12] , \a[13] , \a[14] , \a[15] , \a[16] , \a[17] , \a[18] , \a[19] , \a[20] , \a[21] , \a[22] , \a[23] , \a[24] , \a[25] , \a[26] , \a[27] , \a[28] , \a[29] , \a[30] , \a[31] , \a[32] , \a[33] , \a[34] , \a[35] , \a[36] , \a[37] , \a[38] , \a[39] , \a[40] , \a[41] , \a[42] , \a[43] , \a[44] , \a[45] , \a[46] , \a[47] , \a[48] , \a[49] , \a[50] , \a[51] , \a[52] , \a[53] , \a[54] , \a[55] , \a[56] , \a[57] , \a[58] , \a[59] , \a[60] , \a[61] , \a[62] , \a[63] , \a[64] , \a[65] , \a[66] , \a[67] , \a[68] , \a[69] , \a[70] , \a[71] , \a[72] , \a[73] , \a[74] , \a[75] , \a[76] , \a[77] , \a[78] , \a[79] , \a[80] , \a[81] , \a[82] , \a[83] , \a[84] , \a[85] , \a[86] , \a[87] , \a[88] , \a[89] , \a[90] , \a[91] , \a[92] , \a[93] , \a[94] , \a[95] , \a[96] , \a[97] , \a[98] , \a[99] , \a[100] , \a[101] , \a[102] , \a[103] , \a[104] , \a[105] , \a[106] , \a[107] , \a[108] , \a[109] , \a[110] , \a[111] , \a[112] , \a[113] , \a[114] , \a[115] , \a[116] , \a[117] , \a[118] , \a[119] , \a[120] , \a[121] , \a[122] , \a[123] , \a[124] , \a[125] , \a[126] , \a[127] , \shift[0] , \shift[1] , \shift[2] , \shift[3] , \shift[4] , \shift[5] , \shift[6] , \result[0] , \result[1] , \result[2] , \result[3] , \result[4] , \result[5] , \result[6] , \result[7] , \result[8] , \result[9] , \result[10] , \result[11] , \result[12] , \result[13] , \result[14] , \result[15] , \result[16] , \result[17] , \result[18] , \result[19] , \result[20] , \result[21] , \result[22] , \result[23] , \result[24] , \result[25] , \result[26] , \result[27] , \result[28] , \result[29] , \result[30] , \result[31] , \result[32] , \result[33] , \result[34] , \result[35] , \result[36] , \result[37] , \result[38] , \result[39] , \result[40] , \result[41] , \result[42] , \result[43] , \result[44] , \result[45] , \result[46] , \result[47] , \result[48] , \result[49] , \result[50] , \result[51] , \result[52] , \result[53] , \result[54] , \result[55] , \result[56] , \result[57] , \result[58] , \result[59] , \result[60] , \result[61] , \result[62] , \result[63] , \result[64] , \result[65] , \result[66] , \result[67] , \result[68] , \result[69] , \result[70] , \result[71] , \result[72] , \result[73] , \result[74] , \result[75] , \result[76] , \result[77] , \result[78] , \result[79] , \result[80] , \result[81] , \result[82] , \result[83] , \result[84] , \result[85] , \result[86] , \result[87] , \result[88] , \result[89] , \result[90] , \result[91] , \result[92] , \result[93] , \result[94] , \result[95] , \result[96] , \result[97] , \result[98] , \result[99] , \result[100] , \result[101] , \result[102] , \result[103] , \result[104] , \result[105] , \result[106] , \result[107] , \result[108] , \result[109] , \result[110] , \result[111] , \result[112] , \result[113] , \result[114] , \result[115] , \result[116] , \result[117] , \result[118] , \result[119] , \result[120] , \result[121] , \result[122] , \result[123] , \result[124] , \result[125] , \result[126] , \result[127] );
	input \a[0]  ;
	input \a[1]  ;
	input \a[2]  ;
	input \a[3]  ;
	input \a[4]  ;
	input \a[5]  ;
	input \a[6]  ;
	input \a[7]  ;
	input \a[8]  ;
	input \a[9]  ;
	input \a[10]  ;
	input \a[11]  ;
	input \a[12]  ;
	input \a[13]  ;
	input \a[14]  ;
	input \a[15]  ;
	input \a[16]  ;
	input \a[17]  ;
	input \a[18]  ;
	input \a[19]  ;
	input \a[20]  ;
	input \a[21]  ;
	input \a[22]  ;
	input \a[23]  ;
	input \a[24]  ;
	input \a[25]  ;
	input \a[26]  ;
	input \a[27]  ;
	input \a[28]  ;
	input \a[29]  ;
	input \a[30]  ;
	input \a[31]  ;
	input \a[32]  ;
	input \a[33]  ;
	input \a[34]  ;
	input \a[35]  ;
	input \a[36]  ;
	input \a[37]  ;
	input \a[38]  ;
	input \a[39]  ;
	input \a[40]  ;
	input \a[41]  ;
	input \a[42]  ;
	input \a[43]  ;
	input \a[44]  ;
	input \a[45]  ;
	input \a[46]  ;
	input \a[47]  ;
	input \a[48]  ;
	input \a[49]  ;
	input \a[50]  ;
	input \a[51]  ;
	input \a[52]  ;
	input \a[53]  ;
	input \a[54]  ;
	input \a[55]  ;
	input \a[56]  ;
	input \a[57]  ;
	input \a[58]  ;
	input \a[59]  ;
	input \a[60]  ;
	input \a[61]  ;
	input \a[62]  ;
	input \a[63]  ;
	input \a[64]  ;
	input \a[65]  ;
	input \a[66]  ;
	input \a[67]  ;
	input \a[68]  ;
	input \a[69]  ;
	input \a[70]  ;
	input \a[71]  ;
	input \a[72]  ;
	input \a[73]  ;
	input \a[74]  ;
	input \a[75]  ;
	input \a[76]  ;
	input \a[77]  ;
	input \a[78]  ;
	input \a[79]  ;
	input \a[80]  ;
	input \a[81]  ;
	input \a[82]  ;
	input \a[83]  ;
	input \a[84]  ;
	input \a[85]  ;
	input \a[86]  ;
	input \a[87]  ;
	input \a[88]  ;
	input \a[89]  ;
	input \a[90]  ;
	input \a[91]  ;
	input \a[92]  ;
	input \a[93]  ;
	input \a[94]  ;
	input \a[95]  ;
	input \a[96]  ;
	input \a[97]  ;
	input \a[98]  ;
	input \a[99]  ;
	input \a[100]  ;
	input \a[101]  ;
	input \a[102]  ;
	input \a[103]  ;
	input \a[104]  ;
	input \a[105]  ;
	input \a[106]  ;
	input \a[107]  ;
	input \a[108]  ;
	input \a[109]  ;
	input \a[110]  ;
	input \a[111]  ;
	input \a[112]  ;
	input \a[113]  ;
	input \a[114]  ;
	input \a[115]  ;
	input \a[116]  ;
	input \a[117]  ;
	input \a[118]  ;
	input \a[119]  ;
	input \a[120]  ;
	input \a[121]  ;
	input \a[122]  ;
	input \a[123]  ;
	input \a[124]  ;
	input \a[125]  ;
	input \a[126]  ;
	input \a[127]  ;
	input \shift[0]  ;
	input \shift[1]  ;
	input \shift[2]  ;
	input \shift[3]  ;
	input \shift[4]  ;
	input \shift[5]  ;
	input \shift[6]  ;
	output \result[0]  ;
	output \result[1]  ;
	output \result[2]  ;
	output \result[3]  ;
	output \result[4]  ;
	output \result[5]  ;
	output \result[6]  ;
	output \result[7]  ;
	output \result[8]  ;
	output \result[9]  ;
	output \result[10]  ;
	output \result[11]  ;
	output \result[12]  ;
	output \result[13]  ;
	output \result[14]  ;
	output \result[15]  ;
	output \result[16]  ;
	output \result[17]  ;
	output \result[18]  ;
	output \result[19]  ;
	output \result[20]  ;
	output \result[21]  ;
	output \result[22]  ;
	output \result[23]  ;
	output \result[24]  ;
	output \result[25]  ;
	output \result[26]  ;
	output \result[27]  ;
	output \result[28]  ;
	output \result[29]  ;
	output \result[30]  ;
	output \result[31]  ;
	output \result[32]  ;
	output \result[33]  ;
	output \result[34]  ;
	output \result[35]  ;
	output \result[36]  ;
	output \result[37]  ;
	output \result[38]  ;
	output \result[39]  ;
	output \result[40]  ;
	output \result[41]  ;
	output \result[42]  ;
	output \result[43]  ;
	output \result[44]  ;
	output \result[45]  ;
	output \result[46]  ;
	output \result[47]  ;
	output \result[48]  ;
	output \result[49]  ;
	output \result[50]  ;
	output \result[51]  ;
	output \result[52]  ;
	output \result[53]  ;
	output \result[54]  ;
	output \result[55]  ;
	output \result[56]  ;
	output \result[57]  ;
	output \result[58]  ;
	output \result[59]  ;
	output \result[60]  ;
	output \result[61]  ;
	output \result[62]  ;
	output \result[63]  ;
	output \result[64]  ;
	output \result[65]  ;
	output \result[66]  ;
	output \result[67]  ;
	output \result[68]  ;
	output \result[69]  ;
	output \result[70]  ;
	output \result[71]  ;
	output \result[72]  ;
	output \result[73]  ;
	output \result[74]  ;
	output \result[75]  ;
	output \result[76]  ;
	output \result[77]  ;
	output \result[78]  ;
	output \result[79]  ;
	output \result[80]  ;
	output \result[81]  ;
	output \result[82]  ;
	output \result[83]  ;
	output \result[84]  ;
	output \result[85]  ;
	output \result[86]  ;
	output \result[87]  ;
	output \result[88]  ;
	output \result[89]  ;
	output \result[90]  ;
	output \result[91]  ;
	output \result[92]  ;
	output \result[93]  ;
	output \result[94]  ;
	output \result[95]  ;
	output \result[96]  ;
	output \result[97]  ;
	output \result[98]  ;
	output \result[99]  ;
	output \result[100]  ;
	output \result[101]  ;
	output \result[102]  ;
	output \result[103]  ;
	output \result[104]  ;
	output \result[105]  ;
	output \result[106]  ;
	output \result[107]  ;
	output \result[108]  ;
	output \result[109]  ;
	output \result[110]  ;
	output \result[111]  ;
	output \result[112]  ;
	output \result[113]  ;
	output \result[114]  ;
	output \result[115]  ;
	output \result[116]  ;
	output \result[117]  ;
	output \result[118]  ;
	output \result[119]  ;
	output \result[120]  ;
	output \result[121]  ;
	output \result[122]  ;
	output \result[123]  ;
	output \result[124]  ;
	output \result[125]  ;
	output \result[126]  ;
	output \result[127]  ;
	wire _w1676_ ;
	wire _w1675_ ;
	wire _w1674_ ;
	wire _w1673_ ;
	wire _w1672_ ;
	wire _w1671_ ;
	wire _w1670_ ;
	wire _w1669_ ;
	wire _w1668_ ;
	wire _w1667_ ;
	wire _w1666_ ;
	wire _w1665_ ;
	wire _w1664_ ;
	wire _w1663_ ;
	wire _w1662_ ;
	wire _w1661_ ;
	wire _w1660_ ;
	wire _w1659_ ;
	wire _w1658_ ;
	wire _w1657_ ;
	wire _w1656_ ;
	wire _w1655_ ;
	wire _w1654_ ;
	wire _w1653_ ;
	wire _w1652_ ;
	wire _w1651_ ;
	wire _w1650_ ;
	wire _w1649_ ;
	wire _w1648_ ;
	wire _w1647_ ;
	wire _w1646_ ;
	wire _w1645_ ;
	wire _w1644_ ;
	wire _w1643_ ;
	wire _w1642_ ;
	wire _w1641_ ;
	wire _w1640_ ;
	wire _w1639_ ;
	wire _w1638_ ;
	wire _w1637_ ;
	wire _w1636_ ;
	wire _w1635_ ;
	wire _w1634_ ;
	wire _w1633_ ;
	wire _w1632_ ;
	wire _w1631_ ;
	wire _w1630_ ;
	wire _w1629_ ;
	wire _w1628_ ;
	wire _w1627_ ;
	wire _w1626_ ;
	wire _w1625_ ;
	wire _w1624_ ;
	wire _w1623_ ;
	wire _w1622_ ;
	wire _w1621_ ;
	wire _w1620_ ;
	wire _w1619_ ;
	wire _w1618_ ;
	wire _w1617_ ;
	wire _w1616_ ;
	wire _w1615_ ;
	wire _w1614_ ;
	wire _w1613_ ;
	wire _w1612_ ;
	wire _w1611_ ;
	wire _w1610_ ;
	wire _w1609_ ;
	wire _w1608_ ;
	wire _w1607_ ;
	wire _w1606_ ;
	wire _w1605_ ;
	wire _w1604_ ;
	wire _w1603_ ;
	wire _w1602_ ;
	wire _w1601_ ;
	wire _w1600_ ;
	wire _w1599_ ;
	wire _w1598_ ;
	wire _w1597_ ;
	wire _w1596_ ;
	wire _w1595_ ;
	wire _w1594_ ;
	wire _w1593_ ;
	wire _w1592_ ;
	wire _w1591_ ;
	wire _w1590_ ;
	wire _w1589_ ;
	wire _w1588_ ;
	wire _w1587_ ;
	wire _w1586_ ;
	wire _w1585_ ;
	wire _w1584_ ;
	wire _w1583_ ;
	wire _w1582_ ;
	wire _w1581_ ;
	wire _w1580_ ;
	wire _w1579_ ;
	wire _w1578_ ;
	wire _w1577_ ;
	wire _w1576_ ;
	wire _w1575_ ;
	wire _w1574_ ;
	wire _w1573_ ;
	wire _w1572_ ;
	wire _w1571_ ;
	wire _w1570_ ;
	wire _w1569_ ;
	wire _w1568_ ;
	wire _w1567_ ;
	wire _w1566_ ;
	wire _w1565_ ;
	wire _w1564_ ;
	wire _w1563_ ;
	wire _w1562_ ;
	wire _w1561_ ;
	wire _w1560_ ;
	wire _w1559_ ;
	wire _w1558_ ;
	wire _w1557_ ;
	wire _w1556_ ;
	wire _w1555_ ;
	wire _w1554_ ;
	wire _w1553_ ;
	wire _w1552_ ;
	wire _w1551_ ;
	wire _w1550_ ;
	wire _w1549_ ;
	wire _w1548_ ;
	wire _w1547_ ;
	wire _w1546_ ;
	wire _w1545_ ;
	wire _w1544_ ;
	wire _w1543_ ;
	wire _w1542_ ;
	wire _w1541_ ;
	wire _w1540_ ;
	wire _w1539_ ;
	wire _w1538_ ;
	wire _w1537_ ;
	wire _w1536_ ;
	wire _w1535_ ;
	wire _w1534_ ;
	wire _w1533_ ;
	wire _w1532_ ;
	wire _w1531_ ;
	wire _w1530_ ;
	wire _w1529_ ;
	wire _w1528_ ;
	wire _w1527_ ;
	wire _w1526_ ;
	wire _w1525_ ;
	wire _w1524_ ;
	wire _w1523_ ;
	wire _w1522_ ;
	wire _w1521_ ;
	wire _w1520_ ;
	wire _w1519_ ;
	wire _w1518_ ;
	wire _w1517_ ;
	wire _w1516_ ;
	wire _w1515_ ;
	wire _w1514_ ;
	wire _w1513_ ;
	wire _w1512_ ;
	wire _w1511_ ;
	wire _w1510_ ;
	wire _w1509_ ;
	wire _w1508_ ;
	wire _w1507_ ;
	wire _w1506_ ;
	wire _w1505_ ;
	wire _w1504_ ;
	wire _w1503_ ;
	wire _w1502_ ;
	wire _w1501_ ;
	wire _w1500_ ;
	wire _w1499_ ;
	wire _w1498_ ;
	wire _w1497_ ;
	wire _w1496_ ;
	wire _w1495_ ;
	wire _w1494_ ;
	wire _w1493_ ;
	wire _w1492_ ;
	wire _w1491_ ;
	wire _w1490_ ;
	wire _w1489_ ;
	wire _w1488_ ;
	wire _w1487_ ;
	wire _w1486_ ;
	wire _w1485_ ;
	wire _w1484_ ;
	wire _w1483_ ;
	wire _w1482_ ;
	wire _w1481_ ;
	wire _w1480_ ;
	wire _w1479_ ;
	wire _w1478_ ;
	wire _w1477_ ;
	wire _w1476_ ;
	wire _w1475_ ;
	wire _w1474_ ;
	wire _w1473_ ;
	wire _w1472_ ;
	wire _w1471_ ;
	wire _w1470_ ;
	wire _w1469_ ;
	wire _w1468_ ;
	wire _w1467_ ;
	wire _w1466_ ;
	wire _w1465_ ;
	wire _w1464_ ;
	wire _w1463_ ;
	wire _w1462_ ;
	wire _w1461_ ;
	wire _w1460_ ;
	wire _w1459_ ;
	wire _w1458_ ;
	wire _w1457_ ;
	wire _w1456_ ;
	wire _w1455_ ;
	wire _w1454_ ;
	wire _w1453_ ;
	wire _w1452_ ;
	wire _w1451_ ;
	wire _w1450_ ;
	wire _w1449_ ;
	wire _w1448_ ;
	wire _w1447_ ;
	wire _w1446_ ;
	wire _w1445_ ;
	wire _w1444_ ;
	wire _w1443_ ;
	wire _w1442_ ;
	wire _w1441_ ;
	wire _w1440_ ;
	wire _w1439_ ;
	wire _w1438_ ;
	wire _w1437_ ;
	wire _w1436_ ;
	wire _w1435_ ;
	wire _w1434_ ;
	wire _w1433_ ;
	wire _w1432_ ;
	wire _w1431_ ;
	wire _w1430_ ;
	wire _w1429_ ;
	wire _w1428_ ;
	wire _w1427_ ;
	wire _w1426_ ;
	wire _w1425_ ;
	wire _w1424_ ;
	wire _w1423_ ;
	wire _w1422_ ;
	wire _w1421_ ;
	wire _w1420_ ;
	wire _w1419_ ;
	wire _w1418_ ;
	wire _w1417_ ;
	wire _w1416_ ;
	wire _w1415_ ;
	wire _w1414_ ;
	wire _w1413_ ;
	wire _w1412_ ;
	wire _w1411_ ;
	wire _w1410_ ;
	wire _w1409_ ;
	wire _w1408_ ;
	wire _w1407_ ;
	wire _w1406_ ;
	wire _w1405_ ;
	wire _w1404_ ;
	wire _w1403_ ;
	wire _w1402_ ;
	wire _w1401_ ;
	wire _w1400_ ;
	wire _w1399_ ;
	wire _w1398_ ;
	wire _w1397_ ;
	wire _w1396_ ;
	wire _w1395_ ;
	wire _w1394_ ;
	wire _w1393_ ;
	wire _w1392_ ;
	wire _w1391_ ;
	wire _w1390_ ;
	wire _w1389_ ;
	wire _w1388_ ;
	wire _w1387_ ;
	wire _w1386_ ;
	wire _w1385_ ;
	wire _w1384_ ;
	wire _w1383_ ;
	wire _w1382_ ;
	wire _w1381_ ;
	wire _w1380_ ;
	wire _w1379_ ;
	wire _w1378_ ;
	wire _w1377_ ;
	wire _w1376_ ;
	wire _w1375_ ;
	wire _w1374_ ;
	wire _w1373_ ;
	wire _w1372_ ;
	wire _w1371_ ;
	wire _w1370_ ;
	wire _w1369_ ;
	wire _w1368_ ;
	wire _w1367_ ;
	wire _w1366_ ;
	wire _w1365_ ;
	wire _w1364_ ;
	wire _w1363_ ;
	wire _w1362_ ;
	wire _w1361_ ;
	wire _w1360_ ;
	wire _w1359_ ;
	wire _w1358_ ;
	wire _w1357_ ;
	wire _w1356_ ;
	wire _w1355_ ;
	wire _w1354_ ;
	wire _w1353_ ;
	wire _w1352_ ;
	wire _w1351_ ;
	wire _w1350_ ;
	wire _w1349_ ;
	wire _w1348_ ;
	wire _w1347_ ;
	wire _w1346_ ;
	wire _w1345_ ;
	wire _w1344_ ;
	wire _w1343_ ;
	wire _w1342_ ;
	wire _w1341_ ;
	wire _w1340_ ;
	wire _w1339_ ;
	wire _w1338_ ;
	wire _w1337_ ;
	wire _w1336_ ;
	wire _w1335_ ;
	wire _w1334_ ;
	wire _w1333_ ;
	wire _w1332_ ;
	wire _w1331_ ;
	wire _w1330_ ;
	wire _w1329_ ;
	wire _w1328_ ;
	wire _w1327_ ;
	wire _w1326_ ;
	wire _w1325_ ;
	wire _w1324_ ;
	wire _w1323_ ;
	wire _w1322_ ;
	wire _w1321_ ;
	wire _w1320_ ;
	wire _w1319_ ;
	wire _w1318_ ;
	wire _w1317_ ;
	wire _w1316_ ;
	wire _w1315_ ;
	wire _w1314_ ;
	wire _w1313_ ;
	wire _w1312_ ;
	wire _w1311_ ;
	wire _w1310_ ;
	wire _w1309_ ;
	wire _w1308_ ;
	wire _w1307_ ;
	wire _w1306_ ;
	wire _w1305_ ;
	wire _w1304_ ;
	wire _w1303_ ;
	wire _w1302_ ;
	wire _w1301_ ;
	wire _w1300_ ;
	wire _w1299_ ;
	wire _w1298_ ;
	wire _w1297_ ;
	wire _w1296_ ;
	wire _w1295_ ;
	wire _w1294_ ;
	wire _w1293_ ;
	wire _w1292_ ;
	wire _w1291_ ;
	wire _w1290_ ;
	wire _w1289_ ;
	wire _w1288_ ;
	wire _w1287_ ;
	wire _w1286_ ;
	wire _w1285_ ;
	wire _w1284_ ;
	wire _w1283_ ;
	wire _w1282_ ;
	wire _w1281_ ;
	wire _w1280_ ;
	wire _w1279_ ;
	wire _w1278_ ;
	wire _w1277_ ;
	wire _w1276_ ;
	wire _w1275_ ;
	wire _w1274_ ;
	wire _w1273_ ;
	wire _w1272_ ;
	wire _w1271_ ;
	wire _w1270_ ;
	wire _w1269_ ;
	wire _w1268_ ;
	wire _w1267_ ;
	wire _w1266_ ;
	wire _w1265_ ;
	wire _w1264_ ;
	wire _w1263_ ;
	wire _w1262_ ;
	wire _w1261_ ;
	wire _w1260_ ;
	wire _w1259_ ;
	wire _w1258_ ;
	wire _w1257_ ;
	wire _w1256_ ;
	wire _w1255_ ;
	wire _w1254_ ;
	wire _w1253_ ;
	wire _w1252_ ;
	wire _w1251_ ;
	wire _w1250_ ;
	wire _w1249_ ;
	wire _w1248_ ;
	wire _w1247_ ;
	wire _w1246_ ;
	wire _w677_ ;
	wire _w676_ ;
	wire _w675_ ;
	wire _w674_ ;
	wire _w673_ ;
	wire _w672_ ;
	wire _w671_ ;
	wire _w670_ ;
	wire _w669_ ;
	wire _w668_ ;
	wire _w667_ ;
	wire _w666_ ;
	wire _w665_ ;
	wire _w664_ ;
	wire _w663_ ;
	wire _w662_ ;
	wire _w661_ ;
	wire _w660_ ;
	wire _w659_ ;
	wire _w658_ ;
	wire _w657_ ;
	wire _w656_ ;
	wire _w655_ ;
	wire _w654_ ;
	wire _w653_ ;
	wire _w652_ ;
	wire _w651_ ;
	wire _w650_ ;
	wire _w649_ ;
	wire _w648_ ;
	wire _w647_ ;
	wire _w646_ ;
	wire _w645_ ;
	wire _w644_ ;
	wire _w643_ ;
	wire _w642_ ;
	wire _w641_ ;
	wire _w640_ ;
	wire _w639_ ;
	wire _w638_ ;
	wire _w637_ ;
	wire _w636_ ;
	wire _w635_ ;
	wire _w634_ ;
	wire _w633_ ;
	wire _w632_ ;
	wire _w631_ ;
	wire _w630_ ;
	wire _w629_ ;
	wire _w628_ ;
	wire _w627_ ;
	wire _w626_ ;
	wire _w625_ ;
	wire _w624_ ;
	wire _w623_ ;
	wire _w622_ ;
	wire _w621_ ;
	wire _w620_ ;
	wire _w619_ ;
	wire _w618_ ;
	wire _w617_ ;
	wire _w616_ ;
	wire _w615_ ;
	wire _w614_ ;
	wire _w613_ ;
	wire _w612_ ;
	wire _w611_ ;
	wire _w610_ ;
	wire _w609_ ;
	wire _w608_ ;
	wire _w607_ ;
	wire _w606_ ;
	wire _w605_ ;
	wire _w604_ ;
	wire _w603_ ;
	wire _w602_ ;
	wire _w601_ ;
	wire _w600_ ;
	wire _w599_ ;
	wire _w598_ ;
	wire _w597_ ;
	wire _w596_ ;
	wire _w595_ ;
	wire _w594_ ;
	wire _w593_ ;
	wire _w592_ ;
	wire _w591_ ;
	wire _w590_ ;
	wire _w589_ ;
	wire _w588_ ;
	wire _w587_ ;
	wire _w586_ ;
	wire _w585_ ;
	wire _w584_ ;
	wire _w583_ ;
	wire _w582_ ;
	wire _w581_ ;
	wire _w580_ ;
	wire _w579_ ;
	wire _w578_ ;
	wire _w577_ ;
	wire _w576_ ;
	wire _w575_ ;
	wire _w574_ ;
	wire _w573_ ;
	wire _w572_ ;
	wire _w571_ ;
	wire _w570_ ;
	wire _w569_ ;
	wire _w568_ ;
	wire _w567_ ;
	wire _w566_ ;
	wire _w565_ ;
	wire _w564_ ;
	wire _w563_ ;
	wire _w562_ ;
	wire _w561_ ;
	wire _w560_ ;
	wire _w559_ ;
	wire _w558_ ;
	wire _w557_ ;
	wire _w556_ ;
	wire _w555_ ;
	wire _w554_ ;
	wire _w553_ ;
	wire _w552_ ;
	wire _w551_ ;
	wire _w550_ ;
	wire _w549_ ;
	wire _w548_ ;
	wire _w547_ ;
	wire _w546_ ;
	wire _w545_ ;
	wire _w544_ ;
	wire _w543_ ;
	wire _w542_ ;
	wire _w541_ ;
	wire _w540_ ;
	wire _w539_ ;
	wire _w538_ ;
	wire _w537_ ;
	wire _w536_ ;
	wire _w535_ ;
	wire _w534_ ;
	wire _w533_ ;
	wire _w532_ ;
	wire _w531_ ;
	wire _w530_ ;
	wire _w529_ ;
	wire _w528_ ;
	wire _w527_ ;
	wire _w526_ ;
	wire _w525_ ;
	wire _w524_ ;
	wire _w523_ ;
	wire _w522_ ;
	wire _w521_ ;
	wire _w520_ ;
	wire _w519_ ;
	wire _w518_ ;
	wire _w517_ ;
	wire _w516_ ;
	wire _w515_ ;
	wire _w514_ ;
	wire _w513_ ;
	wire _w512_ ;
	wire _w511_ ;
	wire _w510_ ;
	wire _w509_ ;
	wire _w508_ ;
	wire _w507_ ;
	wire _w506_ ;
	wire _w505_ ;
	wire _w504_ ;
	wire _w503_ ;
	wire _w502_ ;
	wire _w501_ ;
	wire _w500_ ;
	wire _w499_ ;
	wire _w498_ ;
	wire _w497_ ;
	wire _w496_ ;
	wire _w495_ ;
	wire _w494_ ;
	wire _w493_ ;
	wire _w492_ ;
	wire _w491_ ;
	wire _w490_ ;
	wire _w489_ ;
	wire _w488_ ;
	wire _w487_ ;
	wire _w486_ ;
	wire _w485_ ;
	wire _w484_ ;
	wire _w483_ ;
	wire _w482_ ;
	wire _w481_ ;
	wire _w480_ ;
	wire _w479_ ;
	wire _w478_ ;
	wire _w477_ ;
	wire _w476_ ;
	wire _w475_ ;
	wire _w474_ ;
	wire _w473_ ;
	wire _w472_ ;
	wire _w471_ ;
	wire _w470_ ;
	wire _w469_ ;
	wire _w468_ ;
	wire _w467_ ;
	wire _w466_ ;
	wire _w465_ ;
	wire _w464_ ;
	wire _w463_ ;
	wire _w462_ ;
	wire _w461_ ;
	wire _w460_ ;
	wire _w459_ ;
	wire _w458_ ;
	wire _w457_ ;
	wire _w456_ ;
	wire _w455_ ;
	wire _w454_ ;
	wire _w453_ ;
	wire _w452_ ;
	wire _w451_ ;
	wire _w450_ ;
	wire _w449_ ;
	wire _w448_ ;
	wire _w447_ ;
	wire _w446_ ;
	wire _w445_ ;
	wire _w444_ ;
	wire _w443_ ;
	wire _w442_ ;
	wire _w441_ ;
	wire _w440_ ;
	wire _w439_ ;
	wire _w438_ ;
	wire _w437_ ;
	wire _w436_ ;
	wire _w435_ ;
	wire _w434_ ;
	wire _w433_ ;
	wire _w432_ ;
	wire _w431_ ;
	wire _w430_ ;
	wire _w429_ ;
	wire _w428_ ;
	wire _w427_ ;
	wire _w426_ ;
	wire _w425_ ;
	wire _w424_ ;
	wire _w423_ ;
	wire _w422_ ;
	wire _w421_ ;
	wire _w420_ ;
	wire _w419_ ;
	wire _w418_ ;
	wire _w417_ ;
	wire _w416_ ;
	wire _w415_ ;
	wire _w414_ ;
	wire _w413_ ;
	wire _w412_ ;
	wire _w411_ ;
	wire _w410_ ;
	wire _w409_ ;
	wire _w408_ ;
	wire _w407_ ;
	wire _w406_ ;
	wire _w405_ ;
	wire _w404_ ;
	wire _w403_ ;
	wire _w402_ ;
	wire _w401_ ;
	wire _w400_ ;
	wire _w399_ ;
	wire _w398_ ;
	wire _w397_ ;
	wire _w396_ ;
	wire _w395_ ;
	wire _w394_ ;
	wire _w263_ ;
	wire _w262_ ;
	wire _w261_ ;
	wire _w260_ ;
	wire _w259_ ;
	wire _w258_ ;
	wire _w257_ ;
	wire _w256_ ;
	wire _w255_ ;
	wire _w254_ ;
	wire _w253_ ;
	wire _w252_ ;
	wire _w251_ ;
	wire _w250_ ;
	wire _w249_ ;
	wire _w248_ ;
	wire _w247_ ;
	wire _w246_ ;
	wire _w245_ ;
	wire _w244_ ;
	wire _w243_ ;
	wire _w242_ ;
	wire _w241_ ;
	wire _w240_ ;
	wire _w239_ ;
	wire _w238_ ;
	wire _w237_ ;
	wire _w236_ ;
	wire _w235_ ;
	wire _w234_ ;
	wire _w233_ ;
	wire _w232_ ;
	wire _w231_ ;
	wire _w230_ ;
	wire _w229_ ;
	wire _w228_ ;
	wire _w227_ ;
	wire _w226_ ;
	wire _w225_ ;
	wire _w224_ ;
	wire _w223_ ;
	wire _w222_ ;
	wire _w221_ ;
	wire _w220_ ;
	wire _w219_ ;
	wire _w218_ ;
	wire _w217_ ;
	wire _w216_ ;
	wire _w215_ ;
	wire _w214_ ;
	wire _w213_ ;
	wire _w212_ ;
	wire _w211_ ;
	wire _w210_ ;
	wire _w209_ ;
	wire _w208_ ;
	wire _w207_ ;
	wire _w206_ ;
	wire _w205_ ;
	wire _w204_ ;
	wire _w203_ ;
	wire _w202_ ;
	wire _w201_ ;
	wire _w200_ ;
	wire _w199_ ;
	wire _w198_ ;
	wire _w197_ ;
	wire _w196_ ;
	wire _w165_ ;
	wire _w164_ ;
	wire _w163_ ;
	wire _w162_ ;
	wire _w161_ ;
	wire _w160_ ;
	wire _w159_ ;
	wire _w158_ ;
	wire _w157_ ;
	wire _w156_ ;
	wire _w155_ ;
	wire _w154_ ;
	wire _w153_ ;
	wire _w152_ ;
	wire _w151_ ;
	wire _w150_ ;
	wire _w137_ ;
	wire _w138_ ;
	wire _w139_ ;
	wire _w140_ ;
	wire _w141_ ;
	wire _w142_ ;
	wire _w143_ ;
	wire _w144_ ;
	wire _w145_ ;
	wire _w146_ ;
	wire _w147_ ;
	wire _w148_ ;
	wire _w149_ ;
	wire _w166_ ;
	wire _w167_ ;
	wire _w168_ ;
	wire _w169_ ;
	wire _w170_ ;
	wire _w171_ ;
	wire _w172_ ;
	wire _w173_ ;
	wire _w174_ ;
	wire _w175_ ;
	wire _w176_ ;
	wire _w177_ ;
	wire _w178_ ;
	wire _w179_ ;
	wire _w180_ ;
	wire _w181_ ;
	wire _w182_ ;
	wire _w183_ ;
	wire _w184_ ;
	wire _w185_ ;
	wire _w186_ ;
	wire _w187_ ;
	wire _w188_ ;
	wire _w189_ ;
	wire _w190_ ;
	wire _w191_ ;
	wire _w192_ ;
	wire _w193_ ;
	wire _w194_ ;
	wire _w195_ ;
	wire _w264_ ;
	wire _w265_ ;
	wire _w266_ ;
	wire _w267_ ;
	wire _w268_ ;
	wire _w269_ ;
	wire _w270_ ;
	wire _w271_ ;
	wire _w272_ ;
	wire _w273_ ;
	wire _w274_ ;
	wire _w275_ ;
	wire _w276_ ;
	wire _w277_ ;
	wire _w278_ ;
	wire _w279_ ;
	wire _w280_ ;
	wire _w281_ ;
	wire _w282_ ;
	wire _w283_ ;
	wire _w284_ ;
	wire _w285_ ;
	wire _w286_ ;
	wire _w287_ ;
	wire _w288_ ;
	wire _w289_ ;
	wire _w290_ ;
	wire _w291_ ;
	wire _w292_ ;
	wire _w293_ ;
	wire _w294_ ;
	wire _w295_ ;
	wire _w296_ ;
	wire _w297_ ;
	wire _w298_ ;
	wire _w299_ ;
	wire _w300_ ;
	wire _w301_ ;
	wire _w302_ ;
	wire _w303_ ;
	wire _w304_ ;
	wire _w305_ ;
	wire _w306_ ;
	wire _w307_ ;
	wire _w308_ ;
	wire _w309_ ;
	wire _w310_ ;
	wire _w311_ ;
	wire _w312_ ;
	wire _w313_ ;
	wire _w314_ ;
	wire _w315_ ;
	wire _w316_ ;
	wire _w317_ ;
	wire _w318_ ;
	wire _w319_ ;
	wire _w320_ ;
	wire _w321_ ;
	wire _w322_ ;
	wire _w323_ ;
	wire _w324_ ;
	wire _w325_ ;
	wire _w326_ ;
	wire _w327_ ;
	wire _w328_ ;
	wire _w329_ ;
	wire _w330_ ;
	wire _w331_ ;
	wire _w332_ ;
	wire _w333_ ;
	wire _w334_ ;
	wire _w335_ ;
	wire _w336_ ;
	wire _w337_ ;
	wire _w338_ ;
	wire _w339_ ;
	wire _w340_ ;
	wire _w341_ ;
	wire _w342_ ;
	wire _w343_ ;
	wire _w344_ ;
	wire _w345_ ;
	wire _w346_ ;
	wire _w347_ ;
	wire _w348_ ;
	wire _w349_ ;
	wire _w350_ ;
	wire _w351_ ;
	wire _w352_ ;
	wire _w353_ ;
	wire _w354_ ;
	wire _w355_ ;
	wire _w356_ ;
	wire _w357_ ;
	wire _w358_ ;
	wire _w359_ ;
	wire _w360_ ;
	wire _w361_ ;
	wire _w362_ ;
	wire _w363_ ;
	wire _w364_ ;
	wire _w365_ ;
	wire _w366_ ;
	wire _w367_ ;
	wire _w368_ ;
	wire _w369_ ;
	wire _w370_ ;
	wire _w371_ ;
	wire _w372_ ;
	wire _w373_ ;
	wire _w374_ ;
	wire _w375_ ;
	wire _w376_ ;
	wire _w377_ ;
	wire _w378_ ;
	wire _w379_ ;
	wire _w380_ ;
	wire _w381_ ;
	wire _w382_ ;
	wire _w383_ ;
	wire _w384_ ;
	wire _w385_ ;
	wire _w386_ ;
	wire _w387_ ;
	wire _w388_ ;
	wire _w389_ ;
	wire _w390_ ;
	wire _w391_ ;
	wire _w392_ ;
	wire _w393_ ;
	wire _w678_ ;
	wire _w679_ ;
	wire _w680_ ;
	wire _w681_ ;
	wire _w682_ ;
	wire _w683_ ;
	wire _w684_ ;
	wire _w685_ ;
	wire _w686_ ;
	wire _w687_ ;
	wire _w688_ ;
	wire _w689_ ;
	wire _w690_ ;
	wire _w691_ ;
	wire _w692_ ;
	wire _w693_ ;
	wire _w694_ ;
	wire _w695_ ;
	wire _w696_ ;
	wire _w697_ ;
	wire _w698_ ;
	wire _w699_ ;
	wire _w700_ ;
	wire _w701_ ;
	wire _w702_ ;
	wire _w703_ ;
	wire _w704_ ;
	wire _w705_ ;
	wire _w706_ ;
	wire _w707_ ;
	wire _w708_ ;
	wire _w709_ ;
	wire _w710_ ;
	wire _w711_ ;
	wire _w712_ ;
	wire _w713_ ;
	wire _w714_ ;
	wire _w715_ ;
	wire _w716_ ;
	wire _w717_ ;
	wire _w718_ ;
	wire _w719_ ;
	wire _w720_ ;
	wire _w721_ ;
	wire _w722_ ;
	wire _w723_ ;
	wire _w724_ ;
	wire _w725_ ;
	wire _w726_ ;
	wire _w727_ ;
	wire _w728_ ;
	wire _w729_ ;
	wire _w730_ ;
	wire _w731_ ;
	wire _w732_ ;
	wire _w733_ ;
	wire _w734_ ;
	wire _w735_ ;
	wire _w736_ ;
	wire _w737_ ;
	wire _w738_ ;
	wire _w739_ ;
	wire _w740_ ;
	wire _w741_ ;
	wire _w742_ ;
	wire _w743_ ;
	wire _w744_ ;
	wire _w745_ ;
	wire _w746_ ;
	wire _w747_ ;
	wire _w748_ ;
	wire _w749_ ;
	wire _w750_ ;
	wire _w751_ ;
	wire _w752_ ;
	wire _w753_ ;
	wire _w754_ ;
	wire _w755_ ;
	wire _w756_ ;
	wire _w757_ ;
	wire _w758_ ;
	wire _w759_ ;
	wire _w760_ ;
	wire _w761_ ;
	wire _w762_ ;
	wire _w763_ ;
	wire _w764_ ;
	wire _w765_ ;
	wire _w766_ ;
	wire _w767_ ;
	wire _w768_ ;
	wire _w769_ ;
	wire _w770_ ;
	wire _w771_ ;
	wire _w772_ ;
	wire _w773_ ;
	wire _w774_ ;
	wire _w775_ ;
	wire _w776_ ;
	wire _w777_ ;
	wire _w778_ ;
	wire _w779_ ;
	wire _w780_ ;
	wire _w781_ ;
	wire _w782_ ;
	wire _w783_ ;
	wire _w784_ ;
	wire _w785_ ;
	wire _w786_ ;
	wire _w787_ ;
	wire _w788_ ;
	wire _w789_ ;
	wire _w790_ ;
	wire _w791_ ;
	wire _w792_ ;
	wire _w793_ ;
	wire _w794_ ;
	wire _w795_ ;
	wire _w796_ ;
	wire _w797_ ;
	wire _w798_ ;
	wire _w799_ ;
	wire _w800_ ;
	wire _w801_ ;
	wire _w802_ ;
	wire _w803_ ;
	wire _w804_ ;
	wire _w805_ ;
	wire _w806_ ;
	wire _w807_ ;
	wire _w808_ ;
	wire _w809_ ;
	wire _w810_ ;
	wire _w811_ ;
	wire _w812_ ;
	wire _w813_ ;
	wire _w814_ ;
	wire _w815_ ;
	wire _w816_ ;
	wire _w817_ ;
	wire _w818_ ;
	wire _w819_ ;
	wire _w820_ ;
	wire _w821_ ;
	wire _w822_ ;
	wire _w823_ ;
	wire _w824_ ;
	wire _w825_ ;
	wire _w826_ ;
	wire _w827_ ;
	wire _w828_ ;
	wire _w829_ ;
	wire _w830_ ;
	wire _w831_ ;
	wire _w832_ ;
	wire _w833_ ;
	wire _w834_ ;
	wire _w835_ ;
	wire _w836_ ;
	wire _w837_ ;
	wire _w838_ ;
	wire _w839_ ;
	wire _w840_ ;
	wire _w841_ ;
	wire _w842_ ;
	wire _w843_ ;
	wire _w844_ ;
	wire _w845_ ;
	wire _w846_ ;
	wire _w847_ ;
	wire _w848_ ;
	wire _w849_ ;
	wire _w850_ ;
	wire _w851_ ;
	wire _w852_ ;
	wire _w853_ ;
	wire _w854_ ;
	wire _w855_ ;
	wire _w856_ ;
	wire _w857_ ;
	wire _w858_ ;
	wire _w859_ ;
	wire _w860_ ;
	wire _w861_ ;
	wire _w862_ ;
	wire _w863_ ;
	wire _w864_ ;
	wire _w865_ ;
	wire _w866_ ;
	wire _w867_ ;
	wire _w868_ ;
	wire _w869_ ;
	wire _w870_ ;
	wire _w871_ ;
	wire _w872_ ;
	wire _w873_ ;
	wire _w874_ ;
	wire _w875_ ;
	wire _w876_ ;
	wire _w877_ ;
	wire _w878_ ;
	wire _w879_ ;
	wire _w880_ ;
	wire _w881_ ;
	wire _w882_ ;
	wire _w883_ ;
	wire _w884_ ;
	wire _w885_ ;
	wire _w886_ ;
	wire _w887_ ;
	wire _w888_ ;
	wire _w889_ ;
	wire _w890_ ;
	wire _w891_ ;
	wire _w892_ ;
	wire _w893_ ;
	wire _w894_ ;
	wire _w895_ ;
	wire _w896_ ;
	wire _w897_ ;
	wire _w898_ ;
	wire _w899_ ;
	wire _w900_ ;
	wire _w901_ ;
	wire _w902_ ;
	wire _w903_ ;
	wire _w904_ ;
	wire _w905_ ;
	wire _w906_ ;
	wire _w907_ ;
	wire _w908_ ;
	wire _w909_ ;
	wire _w910_ ;
	wire _w911_ ;
	wire _w912_ ;
	wire _w913_ ;
	wire _w914_ ;
	wire _w915_ ;
	wire _w916_ ;
	wire _w917_ ;
	wire _w918_ ;
	wire _w919_ ;
	wire _w920_ ;
	wire _w921_ ;
	wire _w922_ ;
	wire _w923_ ;
	wire _w924_ ;
	wire _w925_ ;
	wire _w926_ ;
	wire _w927_ ;
	wire _w928_ ;
	wire _w929_ ;
	wire _w930_ ;
	wire _w931_ ;
	wire _w932_ ;
	wire _w933_ ;
	wire _w934_ ;
	wire _w935_ ;
	wire _w936_ ;
	wire _w937_ ;
	wire _w938_ ;
	wire _w939_ ;
	wire _w940_ ;
	wire _w941_ ;
	wire _w942_ ;
	wire _w943_ ;
	wire _w944_ ;
	wire _w945_ ;
	wire _w946_ ;
	wire _w947_ ;
	wire _w948_ ;
	wire _w949_ ;
	wire _w950_ ;
	wire _w951_ ;
	wire _w952_ ;
	wire _w953_ ;
	wire _w954_ ;
	wire _w955_ ;
	wire _w956_ ;
	wire _w957_ ;
	wire _w958_ ;
	wire _w959_ ;
	wire _w960_ ;
	wire _w961_ ;
	wire _w962_ ;
	wire _w963_ ;
	wire _w964_ ;
	wire _w965_ ;
	wire _w966_ ;
	wire _w967_ ;
	wire _w968_ ;
	wire _w969_ ;
	wire _w970_ ;
	wire _w971_ ;
	wire _w972_ ;
	wire _w973_ ;
	wire _w974_ ;
	wire _w975_ ;
	wire _w976_ ;
	wire _w977_ ;
	wire _w978_ ;
	wire _w979_ ;
	wire _w980_ ;
	wire _w981_ ;
	wire _w982_ ;
	wire _w983_ ;
	wire _w984_ ;
	wire _w985_ ;
	wire _w986_ ;
	wire _w987_ ;
	wire _w988_ ;
	wire _w989_ ;
	wire _w990_ ;
	wire _w991_ ;
	wire _w992_ ;
	wire _w993_ ;
	wire _w994_ ;
	wire _w995_ ;
	wire _w996_ ;
	wire _w997_ ;
	wire _w998_ ;
	wire _w999_ ;
	wire _w1000_ ;
	wire _w1001_ ;
	wire _w1002_ ;
	wire _w1003_ ;
	wire _w1004_ ;
	wire _w1005_ ;
	wire _w1006_ ;
	wire _w1007_ ;
	wire _w1008_ ;
	wire _w1009_ ;
	wire _w1010_ ;
	wire _w1011_ ;
	wire _w1012_ ;
	wire _w1013_ ;
	wire _w1014_ ;
	wire _w1015_ ;
	wire _w1016_ ;
	wire _w1017_ ;
	wire _w1018_ ;
	wire _w1019_ ;
	wire _w1020_ ;
	wire _w1021_ ;
	wire _w1022_ ;
	wire _w1023_ ;
	wire _w1024_ ;
	wire _w1025_ ;
	wire _w1026_ ;
	wire _w1027_ ;
	wire _w1028_ ;
	wire _w1029_ ;
	wire _w1030_ ;
	wire _w1031_ ;
	wire _w1032_ ;
	wire _w1033_ ;
	wire _w1034_ ;
	wire _w1035_ ;
	wire _w1036_ ;
	wire _w1037_ ;
	wire _w1038_ ;
	wire _w1039_ ;
	wire _w1040_ ;
	wire _w1041_ ;
	wire _w1042_ ;
	wire _w1043_ ;
	wire _w1044_ ;
	wire _w1045_ ;
	wire _w1046_ ;
	wire _w1047_ ;
	wire _w1048_ ;
	wire _w1049_ ;
	wire _w1050_ ;
	wire _w1051_ ;
	wire _w1052_ ;
	wire _w1053_ ;
	wire _w1054_ ;
	wire _w1055_ ;
	wire _w1056_ ;
	wire _w1057_ ;
	wire _w1058_ ;
	wire _w1059_ ;
	wire _w1060_ ;
	wire _w1061_ ;
	wire _w1062_ ;
	wire _w1063_ ;
	wire _w1064_ ;
	wire _w1065_ ;
	wire _w1066_ ;
	wire _w1067_ ;
	wire _w1068_ ;
	wire _w1069_ ;
	wire _w1070_ ;
	wire _w1071_ ;
	wire _w1072_ ;
	wire _w1073_ ;
	wire _w1074_ ;
	wire _w1075_ ;
	wire _w1076_ ;
	wire _w1077_ ;
	wire _w1078_ ;
	wire _w1079_ ;
	wire _w1080_ ;
	wire _w1081_ ;
	wire _w1082_ ;
	wire _w1083_ ;
	wire _w1084_ ;
	wire _w1085_ ;
	wire _w1086_ ;
	wire _w1087_ ;
	wire _w1088_ ;
	wire _w1089_ ;
	wire _w1090_ ;
	wire _w1091_ ;
	wire _w1092_ ;
	wire _w1093_ ;
	wire _w1094_ ;
	wire _w1095_ ;
	wire _w1096_ ;
	wire _w1097_ ;
	wire _w1098_ ;
	wire _w1099_ ;
	wire _w1100_ ;
	wire _w1101_ ;
	wire _w1102_ ;
	wire _w1103_ ;
	wire _w1104_ ;
	wire _w1105_ ;
	wire _w1106_ ;
	wire _w1107_ ;
	wire _w1108_ ;
	wire _w1109_ ;
	wire _w1110_ ;
	wire _w1111_ ;
	wire _w1112_ ;
	wire _w1113_ ;
	wire _w1114_ ;
	wire _w1115_ ;
	wire _w1116_ ;
	wire _w1117_ ;
	wire _w1118_ ;
	wire _w1119_ ;
	wire _w1120_ ;
	wire _w1121_ ;
	wire _w1122_ ;
	wire _w1123_ ;
	wire _w1124_ ;
	wire _w1125_ ;
	wire _w1126_ ;
	wire _w1127_ ;
	wire _w1128_ ;
	wire _w1129_ ;
	wire _w1130_ ;
	wire _w1131_ ;
	wire _w1132_ ;
	wire _w1133_ ;
	wire _w1134_ ;
	wire _w1135_ ;
	wire _w1136_ ;
	wire _w1137_ ;
	wire _w1138_ ;
	wire _w1139_ ;
	wire _w1140_ ;
	wire _w1141_ ;
	wire _w1142_ ;
	wire _w1143_ ;
	wire _w1144_ ;
	wire _w1145_ ;
	wire _w1146_ ;
	wire _w1147_ ;
	wire _w1148_ ;
	wire _w1149_ ;
	wire _w1150_ ;
	wire _w1151_ ;
	wire _w1152_ ;
	wire _w1153_ ;
	wire _w1154_ ;
	wire _w1155_ ;
	wire _w1156_ ;
	wire _w1157_ ;
	wire _w1158_ ;
	wire _w1159_ ;
	wire _w1160_ ;
	wire _w1161_ ;
	wire _w1162_ ;
	wire _w1163_ ;
	wire _w1164_ ;
	wire _w1165_ ;
	wire _w1166_ ;
	wire _w1167_ ;
	wire _w1168_ ;
	wire _w1169_ ;
	wire _w1170_ ;
	wire _w1171_ ;
	wire _w1172_ ;
	wire _w1173_ ;
	wire _w1174_ ;
	wire _w1175_ ;
	wire _w1176_ ;
	wire _w1177_ ;
	wire _w1178_ ;
	wire _w1179_ ;
	wire _w1180_ ;
	wire _w1181_ ;
	wire _w1182_ ;
	wire _w1183_ ;
	wire _w1184_ ;
	wire _w1185_ ;
	wire _w1186_ ;
	wire _w1187_ ;
	wire _w1188_ ;
	wire _w1189_ ;
	wire _w1190_ ;
	wire _w1191_ ;
	wire _w1192_ ;
	wire _w1193_ ;
	wire _w1194_ ;
	wire _w1195_ ;
	wire _w1196_ ;
	wire _w1197_ ;
	wire _w1198_ ;
	wire _w1199_ ;
	wire _w1200_ ;
	wire _w1201_ ;
	wire _w1202_ ;
	wire _w1203_ ;
	wire _w1204_ ;
	wire _w1205_ ;
	wire _w1206_ ;
	wire _w1207_ ;
	wire _w1208_ ;
	wire _w1209_ ;
	wire _w1210_ ;
	wire _w1211_ ;
	wire _w1212_ ;
	wire _w1213_ ;
	wire _w1214_ ;
	wire _w1215_ ;
	wire _w1216_ ;
	wire _w1217_ ;
	wire _w1218_ ;
	wire _w1219_ ;
	wire _w1220_ ;
	wire _w1221_ ;
	wire _w1222_ ;
	wire _w1223_ ;
	wire _w1224_ ;
	wire _w1225_ ;
	wire _w1226_ ;
	wire _w1227_ ;
	wire _w1228_ ;
	wire _w1229_ ;
	wire _w1230_ ;
	wire _w1231_ ;
	wire _w1232_ ;
	wire _w1233_ ;
	wire _w1234_ ;
	wire _w1235_ ;
	wire _w1236_ ;
	wire _w1237_ ;
	wire _w1238_ ;
	wire _w1239_ ;
	wire _w1240_ ;
	wire _w1241_ ;
	wire _w1242_ ;
	wire _w1243_ ;
	wire _w1244_ ;
	wire _w1245_ ;
	LUT2 #(
		.INIT('h1)
	) name0 (
		\shift[2] ,
		\shift[3] ,
		_w137_
	);
	LUT4 #(
		.INIT('hac00)
	) name1 (
		\a[77] ,
		\a[78] ,
		\shift[0] ,
		\shift[1] ,
		_w138_
	);
	LUT4 #(
		.INIT('h00ac)
	) name2 (
		\a[79] ,
		\a[80] ,
		\shift[0] ,
		\shift[1] ,
		_w139_
	);
	LUT3 #(
		.INIT('ha8)
	) name3 (
		_w137_,
		_w138_,
		_w139_,
		_w140_
	);
	LUT2 #(
		.INIT('h2)
	) name4 (
		\shift[2] ,
		\shift[3] ,
		_w141_
	);
	LUT4 #(
		.INIT('hac00)
	) name5 (
		\a[73] ,
		\a[74] ,
		\shift[0] ,
		\shift[1] ,
		_w142_
	);
	LUT4 #(
		.INIT('h00ac)
	) name6 (
		\a[75] ,
		\a[76] ,
		\shift[0] ,
		\shift[1] ,
		_w143_
	);
	LUT3 #(
		.INIT('ha8)
	) name7 (
		_w141_,
		_w142_,
		_w143_,
		_w144_
	);
	LUT2 #(
		.INIT('h8)
	) name8 (
		\shift[2] ,
		\shift[3] ,
		_w145_
	);
	LUT4 #(
		.INIT('hac00)
	) name9 (
		\a[65] ,
		\a[66] ,
		\shift[0] ,
		\shift[1] ,
		_w146_
	);
	LUT4 #(
		.INIT('h00ac)
	) name10 (
		\a[67] ,
		\a[68] ,
		\shift[0] ,
		\shift[1] ,
		_w147_
	);
	LUT3 #(
		.INIT('ha8)
	) name11 (
		_w145_,
		_w146_,
		_w147_,
		_w148_
	);
	LUT2 #(
		.INIT('h4)
	) name12 (
		\shift[2] ,
		\shift[3] ,
		_w149_
	);
	LUT4 #(
		.INIT('hac00)
	) name13 (
		\a[69] ,
		\a[70] ,
		\shift[0] ,
		\shift[1] ,
		_w150_
	);
	LUT4 #(
		.INIT('h00ac)
	) name14 (
		\a[71] ,
		\a[72] ,
		\shift[0] ,
		\shift[1] ,
		_w151_
	);
	LUT3 #(
		.INIT('ha8)
	) name15 (
		_w149_,
		_w150_,
		_w151_,
		_w152_
	);
	LUT4 #(
		.INIT('h0001)
	) name16 (
		_w140_,
		_w144_,
		_w148_,
		_w152_,
		_w153_
	);
	LUT4 #(
		.INIT('hac00)
	) name17 (
		\a[93] ,
		\a[94] ,
		\shift[0] ,
		\shift[1] ,
		_w154_
	);
	LUT4 #(
		.INIT('h00ac)
	) name18 (
		\a[95] ,
		\a[96] ,
		\shift[0] ,
		\shift[1] ,
		_w155_
	);
	LUT3 #(
		.INIT('ha8)
	) name19 (
		_w137_,
		_w154_,
		_w155_,
		_w156_
	);
	LUT4 #(
		.INIT('hac00)
	) name20 (
		\a[89] ,
		\a[90] ,
		\shift[0] ,
		\shift[1] ,
		_w157_
	);
	LUT4 #(
		.INIT('h00ac)
	) name21 (
		\a[91] ,
		\a[92] ,
		\shift[0] ,
		\shift[1] ,
		_w158_
	);
	LUT3 #(
		.INIT('ha8)
	) name22 (
		_w141_,
		_w157_,
		_w158_,
		_w159_
	);
	LUT4 #(
		.INIT('hac00)
	) name23 (
		\a[81] ,
		\a[82] ,
		\shift[0] ,
		\shift[1] ,
		_w160_
	);
	LUT4 #(
		.INIT('h00ac)
	) name24 (
		\a[83] ,
		\a[84] ,
		\shift[0] ,
		\shift[1] ,
		_w161_
	);
	LUT3 #(
		.INIT('ha8)
	) name25 (
		_w145_,
		_w160_,
		_w161_,
		_w162_
	);
	LUT4 #(
		.INIT('hac00)
	) name26 (
		\a[85] ,
		\a[86] ,
		\shift[0] ,
		\shift[1] ,
		_w163_
	);
	LUT4 #(
		.INIT('h00ac)
	) name27 (
		\a[87] ,
		\a[88] ,
		\shift[0] ,
		\shift[1] ,
		_w164_
	);
	LUT3 #(
		.INIT('ha8)
	) name28 (
		_w149_,
		_w163_,
		_w164_,
		_w165_
	);
	LUT4 #(
		.INIT('h0001)
	) name29 (
		_w156_,
		_w159_,
		_w162_,
		_w165_,
		_w166_
	);
	LUT4 #(
		.INIT('hf7b3)
	) name30 (
		\shift[4] ,
		\shift[5] ,
		_w153_,
		_w166_,
		_w167_
	);
	LUT4 #(
		.INIT('hac00)
	) name31 (
		\a[125] ,
		\a[126] ,
		\shift[0] ,
		\shift[1] ,
		_w168_
	);
	LUT4 #(
		.INIT('h00ca)
	) name32 (
		\a[0] ,
		\a[127] ,
		\shift[0] ,
		\shift[1] ,
		_w169_
	);
	LUT3 #(
		.INIT('ha8)
	) name33 (
		_w137_,
		_w168_,
		_w169_,
		_w170_
	);
	LUT4 #(
		.INIT('hac00)
	) name34 (
		\a[121] ,
		\a[122] ,
		\shift[0] ,
		\shift[1] ,
		_w171_
	);
	LUT4 #(
		.INIT('h00ac)
	) name35 (
		\a[123] ,
		\a[124] ,
		\shift[0] ,
		\shift[1] ,
		_w172_
	);
	LUT3 #(
		.INIT('ha8)
	) name36 (
		_w141_,
		_w171_,
		_w172_,
		_w173_
	);
	LUT4 #(
		.INIT('hac00)
	) name37 (
		\a[113] ,
		\a[114] ,
		\shift[0] ,
		\shift[1] ,
		_w174_
	);
	LUT4 #(
		.INIT('h00ac)
	) name38 (
		\a[115] ,
		\a[116] ,
		\shift[0] ,
		\shift[1] ,
		_w175_
	);
	LUT3 #(
		.INIT('ha8)
	) name39 (
		_w145_,
		_w174_,
		_w175_,
		_w176_
	);
	LUT4 #(
		.INIT('hac00)
	) name40 (
		\a[117] ,
		\a[118] ,
		\shift[0] ,
		\shift[1] ,
		_w177_
	);
	LUT4 #(
		.INIT('h00ac)
	) name41 (
		\a[119] ,
		\a[120] ,
		\shift[0] ,
		\shift[1] ,
		_w178_
	);
	LUT3 #(
		.INIT('ha8)
	) name42 (
		_w149_,
		_w177_,
		_w178_,
		_w179_
	);
	LUT4 #(
		.INIT('h0001)
	) name43 (
		_w170_,
		_w173_,
		_w176_,
		_w179_,
		_w180_
	);
	LUT4 #(
		.INIT('hac00)
	) name44 (
		\a[109] ,
		\a[110] ,
		\shift[0] ,
		\shift[1] ,
		_w181_
	);
	LUT4 #(
		.INIT('h00ac)
	) name45 (
		\a[111] ,
		\a[112] ,
		\shift[0] ,
		\shift[1] ,
		_w182_
	);
	LUT3 #(
		.INIT('ha8)
	) name46 (
		_w137_,
		_w181_,
		_w182_,
		_w183_
	);
	LUT4 #(
		.INIT('hac00)
	) name47 (
		\a[105] ,
		\a[106] ,
		\shift[0] ,
		\shift[1] ,
		_w184_
	);
	LUT4 #(
		.INIT('h00ac)
	) name48 (
		\a[107] ,
		\a[108] ,
		\shift[0] ,
		\shift[1] ,
		_w185_
	);
	LUT3 #(
		.INIT('ha8)
	) name49 (
		_w141_,
		_w184_,
		_w185_,
		_w186_
	);
	LUT4 #(
		.INIT('hac00)
	) name50 (
		\a[97] ,
		\a[98] ,
		\shift[0] ,
		\shift[1] ,
		_w187_
	);
	LUT4 #(
		.INIT('h00ac)
	) name51 (
		\a[99] ,
		\a[100] ,
		\shift[0] ,
		\shift[1] ,
		_w188_
	);
	LUT3 #(
		.INIT('ha8)
	) name52 (
		_w145_,
		_w187_,
		_w188_,
		_w189_
	);
	LUT4 #(
		.INIT('hac00)
	) name53 (
		\a[101] ,
		\a[102] ,
		\shift[0] ,
		\shift[1] ,
		_w190_
	);
	LUT4 #(
		.INIT('h00ac)
	) name54 (
		\a[103] ,
		\a[104] ,
		\shift[0] ,
		\shift[1] ,
		_w191_
	);
	LUT3 #(
		.INIT('ha8)
	) name55 (
		_w149_,
		_w190_,
		_w191_,
		_w192_
	);
	LUT4 #(
		.INIT('h0001)
	) name56 (
		_w183_,
		_w186_,
		_w189_,
		_w192_,
		_w193_
	);
	LUT4 #(
		.INIT('hfedc)
	) name57 (
		\shift[4] ,
		\shift[5] ,
		_w180_,
		_w193_,
		_w194_
	);
	LUT3 #(
		.INIT('h15)
	) name58 (
		\shift[6] ,
		_w167_,
		_w194_,
		_w195_
	);
	LUT4 #(
		.INIT('hac00)
	) name59 (
		\a[13] ,
		\a[14] ,
		\shift[0] ,
		\shift[1] ,
		_w196_
	);
	LUT4 #(
		.INIT('h00ac)
	) name60 (
		\a[15] ,
		\a[16] ,
		\shift[0] ,
		\shift[1] ,
		_w197_
	);
	LUT3 #(
		.INIT('ha8)
	) name61 (
		_w137_,
		_w196_,
		_w197_,
		_w198_
	);
	LUT4 #(
		.INIT('hac00)
	) name62 (
		\a[9] ,
		\a[10] ,
		\shift[0] ,
		\shift[1] ,
		_w199_
	);
	LUT4 #(
		.INIT('h00ac)
	) name63 (
		\a[11] ,
		\a[12] ,
		\shift[0] ,
		\shift[1] ,
		_w200_
	);
	LUT3 #(
		.INIT('ha8)
	) name64 (
		_w141_,
		_w199_,
		_w200_,
		_w201_
	);
	LUT4 #(
		.INIT('hac00)
	) name65 (
		\a[1] ,
		\a[2] ,
		\shift[0] ,
		\shift[1] ,
		_w202_
	);
	LUT4 #(
		.INIT('h00ac)
	) name66 (
		\a[3] ,
		\a[4] ,
		\shift[0] ,
		\shift[1] ,
		_w203_
	);
	LUT3 #(
		.INIT('ha8)
	) name67 (
		_w145_,
		_w202_,
		_w203_,
		_w204_
	);
	LUT4 #(
		.INIT('hac00)
	) name68 (
		\a[5] ,
		\a[6] ,
		\shift[0] ,
		\shift[1] ,
		_w205_
	);
	LUT4 #(
		.INIT('h00ac)
	) name69 (
		\a[7] ,
		\a[8] ,
		\shift[0] ,
		\shift[1] ,
		_w206_
	);
	LUT3 #(
		.INIT('ha8)
	) name70 (
		_w149_,
		_w205_,
		_w206_,
		_w207_
	);
	LUT4 #(
		.INIT('h0001)
	) name71 (
		_w198_,
		_w201_,
		_w204_,
		_w207_,
		_w208_
	);
	LUT4 #(
		.INIT('hac00)
	) name72 (
		\a[29] ,
		\a[30] ,
		\shift[0] ,
		\shift[1] ,
		_w209_
	);
	LUT4 #(
		.INIT('h00ac)
	) name73 (
		\a[31] ,
		\a[32] ,
		\shift[0] ,
		\shift[1] ,
		_w210_
	);
	LUT3 #(
		.INIT('ha8)
	) name74 (
		_w137_,
		_w209_,
		_w210_,
		_w211_
	);
	LUT4 #(
		.INIT('hac00)
	) name75 (
		\a[25] ,
		\a[26] ,
		\shift[0] ,
		\shift[1] ,
		_w212_
	);
	LUT4 #(
		.INIT('h00ac)
	) name76 (
		\a[27] ,
		\a[28] ,
		\shift[0] ,
		\shift[1] ,
		_w213_
	);
	LUT3 #(
		.INIT('ha8)
	) name77 (
		_w141_,
		_w212_,
		_w213_,
		_w214_
	);
	LUT4 #(
		.INIT('hac00)
	) name78 (
		\a[17] ,
		\a[18] ,
		\shift[0] ,
		\shift[1] ,
		_w215_
	);
	LUT4 #(
		.INIT('h00ac)
	) name79 (
		\a[19] ,
		\a[20] ,
		\shift[0] ,
		\shift[1] ,
		_w216_
	);
	LUT3 #(
		.INIT('ha8)
	) name80 (
		_w145_,
		_w215_,
		_w216_,
		_w217_
	);
	LUT4 #(
		.INIT('hac00)
	) name81 (
		\a[21] ,
		\a[22] ,
		\shift[0] ,
		\shift[1] ,
		_w218_
	);
	LUT4 #(
		.INIT('h00ac)
	) name82 (
		\a[23] ,
		\a[24] ,
		\shift[0] ,
		\shift[1] ,
		_w219_
	);
	LUT3 #(
		.INIT('ha8)
	) name83 (
		_w149_,
		_w218_,
		_w219_,
		_w220_
	);
	LUT4 #(
		.INIT('h0001)
	) name84 (
		_w211_,
		_w214_,
		_w217_,
		_w220_,
		_w221_
	);
	LUT4 #(
		.INIT('hf7b3)
	) name85 (
		\shift[4] ,
		\shift[5] ,
		_w208_,
		_w221_,
		_w222_
	);
	LUT4 #(
		.INIT('hac00)
	) name86 (
		\a[61] ,
		\a[62] ,
		\shift[0] ,
		\shift[1] ,
		_w223_
	);
	LUT4 #(
		.INIT('h00ac)
	) name87 (
		\a[63] ,
		\a[64] ,
		\shift[0] ,
		\shift[1] ,
		_w224_
	);
	LUT3 #(
		.INIT('ha8)
	) name88 (
		_w137_,
		_w223_,
		_w224_,
		_w225_
	);
	LUT4 #(
		.INIT('hac00)
	) name89 (
		\a[57] ,
		\a[58] ,
		\shift[0] ,
		\shift[1] ,
		_w226_
	);
	LUT4 #(
		.INIT('h00ac)
	) name90 (
		\a[59] ,
		\a[60] ,
		\shift[0] ,
		\shift[1] ,
		_w227_
	);
	LUT3 #(
		.INIT('ha8)
	) name91 (
		_w141_,
		_w226_,
		_w227_,
		_w228_
	);
	LUT4 #(
		.INIT('hac00)
	) name92 (
		\a[49] ,
		\a[50] ,
		\shift[0] ,
		\shift[1] ,
		_w229_
	);
	LUT4 #(
		.INIT('h00ac)
	) name93 (
		\a[51] ,
		\a[52] ,
		\shift[0] ,
		\shift[1] ,
		_w230_
	);
	LUT3 #(
		.INIT('ha8)
	) name94 (
		_w145_,
		_w229_,
		_w230_,
		_w231_
	);
	LUT4 #(
		.INIT('hac00)
	) name95 (
		\a[53] ,
		\a[54] ,
		\shift[0] ,
		\shift[1] ,
		_w232_
	);
	LUT4 #(
		.INIT('h00ac)
	) name96 (
		\a[55] ,
		\a[56] ,
		\shift[0] ,
		\shift[1] ,
		_w233_
	);
	LUT3 #(
		.INIT('ha8)
	) name97 (
		_w149_,
		_w232_,
		_w233_,
		_w234_
	);
	LUT4 #(
		.INIT('h0001)
	) name98 (
		_w225_,
		_w228_,
		_w231_,
		_w234_,
		_w235_
	);
	LUT4 #(
		.INIT('hac00)
	) name99 (
		\a[45] ,
		\a[46] ,
		\shift[0] ,
		\shift[1] ,
		_w236_
	);
	LUT4 #(
		.INIT('h00ac)
	) name100 (
		\a[47] ,
		\a[48] ,
		\shift[0] ,
		\shift[1] ,
		_w237_
	);
	LUT3 #(
		.INIT('ha8)
	) name101 (
		_w137_,
		_w236_,
		_w237_,
		_w238_
	);
	LUT4 #(
		.INIT('hac00)
	) name102 (
		\a[41] ,
		\a[42] ,
		\shift[0] ,
		\shift[1] ,
		_w239_
	);
	LUT4 #(
		.INIT('h00ac)
	) name103 (
		\a[43] ,
		\a[44] ,
		\shift[0] ,
		\shift[1] ,
		_w240_
	);
	LUT3 #(
		.INIT('ha8)
	) name104 (
		_w141_,
		_w239_,
		_w240_,
		_w241_
	);
	LUT4 #(
		.INIT('hac00)
	) name105 (
		\a[33] ,
		\a[34] ,
		\shift[0] ,
		\shift[1] ,
		_w242_
	);
	LUT4 #(
		.INIT('h00ac)
	) name106 (
		\a[35] ,
		\a[36] ,
		\shift[0] ,
		\shift[1] ,
		_w243_
	);
	LUT3 #(
		.INIT('ha8)
	) name107 (
		_w145_,
		_w242_,
		_w243_,
		_w244_
	);
	LUT4 #(
		.INIT('ha00c)
	) name108 (
		\a[37] ,
		\a[40] ,
		\shift[0] ,
		\shift[1] ,
		_w245_
	);
	LUT4 #(
		.INIT('hf53f)
	) name109 (
		\a[38] ,
		\a[39] ,
		\shift[0] ,
		\shift[1] ,
		_w246_
	);
	LUT3 #(
		.INIT('h8a)
	) name110 (
		_w149_,
		_w245_,
		_w246_,
		_w247_
	);
	LUT4 #(
		.INIT('h0001)
	) name111 (
		_w238_,
		_w241_,
		_w244_,
		_w247_,
		_w248_
	);
	LUT4 #(
		.INIT('hfedc)
	) name112 (
		\shift[4] ,
		\shift[5] ,
		_w235_,
		_w248_,
		_w249_
	);
	LUT3 #(
		.INIT('h2a)
	) name113 (
		\shift[6] ,
		_w222_,
		_w249_,
		_w250_
	);
	LUT2 #(
		.INIT('he)
	) name114 (
		_w195_,
		_w250_,
		_w251_
	);
	LUT4 #(
		.INIT('ha00c)
	) name115 (
		\a[78] ,
		\a[81] ,
		\shift[0] ,
		\shift[1] ,
		_w252_
	);
	LUT4 #(
		.INIT('hf53f)
	) name116 (
		\a[79] ,
		\a[80] ,
		\shift[0] ,
		\shift[1] ,
		_w253_
	);
	LUT3 #(
		.INIT('h8a)
	) name117 (
		_w137_,
		_w252_,
		_w253_,
		_w254_
	);
	LUT4 #(
		.INIT('ha00c)
	) name118 (
		\a[74] ,
		\a[77] ,
		\shift[0] ,
		\shift[1] ,
		_w255_
	);
	LUT4 #(
		.INIT('hf53f)
	) name119 (
		\a[75] ,
		\a[76] ,
		\shift[0] ,
		\shift[1] ,
		_w256_
	);
	LUT3 #(
		.INIT('h8a)
	) name120 (
		_w141_,
		_w255_,
		_w256_,
		_w257_
	);
	LUT4 #(
		.INIT('ha00c)
	) name121 (
		\a[66] ,
		\a[69] ,
		\shift[0] ,
		\shift[1] ,
		_w258_
	);
	LUT4 #(
		.INIT('hf53f)
	) name122 (
		\a[67] ,
		\a[68] ,
		\shift[0] ,
		\shift[1] ,
		_w259_
	);
	LUT3 #(
		.INIT('h8a)
	) name123 (
		_w145_,
		_w258_,
		_w259_,
		_w260_
	);
	LUT4 #(
		.INIT('ha00c)
	) name124 (
		\a[70] ,
		\a[73] ,
		\shift[0] ,
		\shift[1] ,
		_w261_
	);
	LUT4 #(
		.INIT('hf53f)
	) name125 (
		\a[71] ,
		\a[72] ,
		\shift[0] ,
		\shift[1] ,
		_w262_
	);
	LUT3 #(
		.INIT('h8a)
	) name126 (
		_w149_,
		_w261_,
		_w262_,
		_w263_
	);
	LUT4 #(
		.INIT('h0001)
	) name127 (
		_w254_,
		_w257_,
		_w260_,
		_w263_,
		_w264_
	);
	LUT4 #(
		.INIT('ha00c)
	) name128 (
		\a[94] ,
		\a[97] ,
		\shift[0] ,
		\shift[1] ,
		_w265_
	);
	LUT4 #(
		.INIT('hf53f)
	) name129 (
		\a[95] ,
		\a[96] ,
		\shift[0] ,
		\shift[1] ,
		_w266_
	);
	LUT3 #(
		.INIT('h8a)
	) name130 (
		_w137_,
		_w265_,
		_w266_,
		_w267_
	);
	LUT4 #(
		.INIT('ha00c)
	) name131 (
		\a[90] ,
		\a[93] ,
		\shift[0] ,
		\shift[1] ,
		_w268_
	);
	LUT4 #(
		.INIT('hf53f)
	) name132 (
		\a[91] ,
		\a[92] ,
		\shift[0] ,
		\shift[1] ,
		_w269_
	);
	LUT3 #(
		.INIT('h8a)
	) name133 (
		_w141_,
		_w268_,
		_w269_,
		_w270_
	);
	LUT4 #(
		.INIT('ha00c)
	) name134 (
		\a[82] ,
		\a[85] ,
		\shift[0] ,
		\shift[1] ,
		_w271_
	);
	LUT4 #(
		.INIT('hf53f)
	) name135 (
		\a[83] ,
		\a[84] ,
		\shift[0] ,
		\shift[1] ,
		_w272_
	);
	LUT3 #(
		.INIT('h8a)
	) name136 (
		_w145_,
		_w271_,
		_w272_,
		_w273_
	);
	LUT4 #(
		.INIT('ha00c)
	) name137 (
		\a[86] ,
		\a[89] ,
		\shift[0] ,
		\shift[1] ,
		_w274_
	);
	LUT4 #(
		.INIT('hf53f)
	) name138 (
		\a[87] ,
		\a[88] ,
		\shift[0] ,
		\shift[1] ,
		_w275_
	);
	LUT3 #(
		.INIT('h8a)
	) name139 (
		_w149_,
		_w274_,
		_w275_,
		_w276_
	);
	LUT4 #(
		.INIT('h0001)
	) name140 (
		_w267_,
		_w270_,
		_w273_,
		_w276_,
		_w277_
	);
	LUT4 #(
		.INIT('hf7b3)
	) name141 (
		\shift[4] ,
		\shift[5] ,
		_w264_,
		_w277_,
		_w278_
	);
	LUT4 #(
		.INIT('hc00a)
	) name142 (
		\a[1] ,
		\a[126] ,
		\shift[0] ,
		\shift[1] ,
		_w279_
	);
	LUT4 #(
		.INIT('hf35f)
	) name143 (
		\a[0] ,
		\a[127] ,
		\shift[0] ,
		\shift[1] ,
		_w280_
	);
	LUT3 #(
		.INIT('h8a)
	) name144 (
		_w137_,
		_w279_,
		_w280_,
		_w281_
	);
	LUT4 #(
		.INIT('ha00c)
	) name145 (
		\a[122] ,
		\a[125] ,
		\shift[0] ,
		\shift[1] ,
		_w282_
	);
	LUT4 #(
		.INIT('hf53f)
	) name146 (
		\a[123] ,
		\a[124] ,
		\shift[0] ,
		\shift[1] ,
		_w283_
	);
	LUT3 #(
		.INIT('h8a)
	) name147 (
		_w141_,
		_w282_,
		_w283_,
		_w284_
	);
	LUT4 #(
		.INIT('ha00c)
	) name148 (
		\a[114] ,
		\a[117] ,
		\shift[0] ,
		\shift[1] ,
		_w285_
	);
	LUT4 #(
		.INIT('hf53f)
	) name149 (
		\a[115] ,
		\a[116] ,
		\shift[0] ,
		\shift[1] ,
		_w286_
	);
	LUT3 #(
		.INIT('h8a)
	) name150 (
		_w145_,
		_w285_,
		_w286_,
		_w287_
	);
	LUT4 #(
		.INIT('ha00c)
	) name151 (
		\a[118] ,
		\a[121] ,
		\shift[0] ,
		\shift[1] ,
		_w288_
	);
	LUT4 #(
		.INIT('hf53f)
	) name152 (
		\a[119] ,
		\a[120] ,
		\shift[0] ,
		\shift[1] ,
		_w289_
	);
	LUT3 #(
		.INIT('h8a)
	) name153 (
		_w149_,
		_w288_,
		_w289_,
		_w290_
	);
	LUT4 #(
		.INIT('h0001)
	) name154 (
		_w281_,
		_w284_,
		_w287_,
		_w290_,
		_w291_
	);
	LUT4 #(
		.INIT('ha00c)
	) name155 (
		\a[110] ,
		\a[113] ,
		\shift[0] ,
		\shift[1] ,
		_w292_
	);
	LUT4 #(
		.INIT('hf53f)
	) name156 (
		\a[111] ,
		\a[112] ,
		\shift[0] ,
		\shift[1] ,
		_w293_
	);
	LUT3 #(
		.INIT('h8a)
	) name157 (
		_w137_,
		_w292_,
		_w293_,
		_w294_
	);
	LUT4 #(
		.INIT('ha00c)
	) name158 (
		\a[106] ,
		\a[109] ,
		\shift[0] ,
		\shift[1] ,
		_w295_
	);
	LUT4 #(
		.INIT('hf53f)
	) name159 (
		\a[107] ,
		\a[108] ,
		\shift[0] ,
		\shift[1] ,
		_w296_
	);
	LUT3 #(
		.INIT('h8a)
	) name160 (
		_w141_,
		_w295_,
		_w296_,
		_w297_
	);
	LUT4 #(
		.INIT('ha00c)
	) name161 (
		\a[98] ,
		\a[101] ,
		\shift[0] ,
		\shift[1] ,
		_w298_
	);
	LUT4 #(
		.INIT('hf53f)
	) name162 (
		\a[99] ,
		\a[100] ,
		\shift[0] ,
		\shift[1] ,
		_w299_
	);
	LUT3 #(
		.INIT('h8a)
	) name163 (
		_w145_,
		_w298_,
		_w299_,
		_w300_
	);
	LUT4 #(
		.INIT('ha00c)
	) name164 (
		\a[102] ,
		\a[105] ,
		\shift[0] ,
		\shift[1] ,
		_w301_
	);
	LUT4 #(
		.INIT('hf53f)
	) name165 (
		\a[103] ,
		\a[104] ,
		\shift[0] ,
		\shift[1] ,
		_w302_
	);
	LUT3 #(
		.INIT('h8a)
	) name166 (
		_w149_,
		_w301_,
		_w302_,
		_w303_
	);
	LUT4 #(
		.INIT('h0001)
	) name167 (
		_w294_,
		_w297_,
		_w300_,
		_w303_,
		_w304_
	);
	LUT4 #(
		.INIT('hfedc)
	) name168 (
		\shift[4] ,
		\shift[5] ,
		_w291_,
		_w304_,
		_w305_
	);
	LUT3 #(
		.INIT('h15)
	) name169 (
		\shift[6] ,
		_w278_,
		_w305_,
		_w306_
	);
	LUT4 #(
		.INIT('ha00c)
	) name170 (
		\a[62] ,
		\a[65] ,
		\shift[0] ,
		\shift[1] ,
		_w307_
	);
	LUT4 #(
		.INIT('hf53f)
	) name171 (
		\a[63] ,
		\a[64] ,
		\shift[0] ,
		\shift[1] ,
		_w308_
	);
	LUT3 #(
		.INIT('h8a)
	) name172 (
		_w137_,
		_w307_,
		_w308_,
		_w309_
	);
	LUT4 #(
		.INIT('ha00c)
	) name173 (
		\a[58] ,
		\a[61] ,
		\shift[0] ,
		\shift[1] ,
		_w310_
	);
	LUT4 #(
		.INIT('hf53f)
	) name174 (
		\a[59] ,
		\a[60] ,
		\shift[0] ,
		\shift[1] ,
		_w311_
	);
	LUT3 #(
		.INIT('h8a)
	) name175 (
		_w141_,
		_w310_,
		_w311_,
		_w312_
	);
	LUT4 #(
		.INIT('ha00c)
	) name176 (
		\a[50] ,
		\a[53] ,
		\shift[0] ,
		\shift[1] ,
		_w313_
	);
	LUT4 #(
		.INIT('hf53f)
	) name177 (
		\a[51] ,
		\a[52] ,
		\shift[0] ,
		\shift[1] ,
		_w314_
	);
	LUT3 #(
		.INIT('h8a)
	) name178 (
		_w145_,
		_w313_,
		_w314_,
		_w315_
	);
	LUT4 #(
		.INIT('ha00c)
	) name179 (
		\a[54] ,
		\a[57] ,
		\shift[0] ,
		\shift[1] ,
		_w316_
	);
	LUT4 #(
		.INIT('hf53f)
	) name180 (
		\a[55] ,
		\a[56] ,
		\shift[0] ,
		\shift[1] ,
		_w317_
	);
	LUT3 #(
		.INIT('h8a)
	) name181 (
		_w149_,
		_w316_,
		_w317_,
		_w318_
	);
	LUT4 #(
		.INIT('h0001)
	) name182 (
		_w309_,
		_w312_,
		_w315_,
		_w318_,
		_w319_
	);
	LUT4 #(
		.INIT('ha00c)
	) name183 (
		\a[14] ,
		\a[17] ,
		\shift[0] ,
		\shift[1] ,
		_w320_
	);
	LUT4 #(
		.INIT('hf53f)
	) name184 (
		\a[15] ,
		\a[16] ,
		\shift[0] ,
		\shift[1] ,
		_w321_
	);
	LUT3 #(
		.INIT('h8a)
	) name185 (
		_w137_,
		_w320_,
		_w321_,
		_w322_
	);
	LUT4 #(
		.INIT('ha00c)
	) name186 (
		\a[10] ,
		\a[13] ,
		\shift[0] ,
		\shift[1] ,
		_w323_
	);
	LUT4 #(
		.INIT('hf53f)
	) name187 (
		\a[11] ,
		\a[12] ,
		\shift[0] ,
		\shift[1] ,
		_w324_
	);
	LUT3 #(
		.INIT('h8a)
	) name188 (
		_w141_,
		_w323_,
		_w324_,
		_w325_
	);
	LUT4 #(
		.INIT('ha00c)
	) name189 (
		\a[2] ,
		\a[5] ,
		\shift[0] ,
		\shift[1] ,
		_w326_
	);
	LUT4 #(
		.INIT('hf53f)
	) name190 (
		\a[3] ,
		\a[4] ,
		\shift[0] ,
		\shift[1] ,
		_w327_
	);
	LUT3 #(
		.INIT('h8a)
	) name191 (
		_w145_,
		_w326_,
		_w327_,
		_w328_
	);
	LUT4 #(
		.INIT('ha00c)
	) name192 (
		\a[6] ,
		\a[9] ,
		\shift[0] ,
		\shift[1] ,
		_w329_
	);
	LUT4 #(
		.INIT('hf53f)
	) name193 (
		\a[7] ,
		\a[8] ,
		\shift[0] ,
		\shift[1] ,
		_w330_
	);
	LUT3 #(
		.INIT('h8a)
	) name194 (
		_w149_,
		_w329_,
		_w330_,
		_w331_
	);
	LUT4 #(
		.INIT('h0001)
	) name195 (
		_w322_,
		_w325_,
		_w328_,
		_w331_,
		_w332_
	);
	LUT4 #(
		.INIT('hfe76)
	) name196 (
		\shift[4] ,
		\shift[5] ,
		_w319_,
		_w332_,
		_w333_
	);
	LUT4 #(
		.INIT('ha00c)
	) name197 (
		\a[46] ,
		\a[49] ,
		\shift[0] ,
		\shift[1] ,
		_w334_
	);
	LUT4 #(
		.INIT('hf53f)
	) name198 (
		\a[47] ,
		\a[48] ,
		\shift[0] ,
		\shift[1] ,
		_w335_
	);
	LUT3 #(
		.INIT('h8a)
	) name199 (
		_w137_,
		_w334_,
		_w335_,
		_w336_
	);
	LUT4 #(
		.INIT('hac00)
	) name200 (
		\a[42] ,
		\a[43] ,
		\shift[0] ,
		\shift[1] ,
		_w337_
	);
	LUT4 #(
		.INIT('h00ac)
	) name201 (
		\a[44] ,
		\a[45] ,
		\shift[0] ,
		\shift[1] ,
		_w338_
	);
	LUT3 #(
		.INIT('ha8)
	) name202 (
		_w141_,
		_w337_,
		_w338_,
		_w339_
	);
	LUT4 #(
		.INIT('ha00c)
	) name203 (
		\a[34] ,
		\a[37] ,
		\shift[0] ,
		\shift[1] ,
		_w340_
	);
	LUT4 #(
		.INIT('hf53f)
	) name204 (
		\a[35] ,
		\a[36] ,
		\shift[0] ,
		\shift[1] ,
		_w341_
	);
	LUT3 #(
		.INIT('h8a)
	) name205 (
		_w145_,
		_w340_,
		_w341_,
		_w342_
	);
	LUT4 #(
		.INIT('h00ac)
	) name206 (
		\a[40] ,
		\a[41] ,
		\shift[0] ,
		\shift[1] ,
		_w343_
	);
	LUT4 #(
		.INIT('hac00)
	) name207 (
		\a[38] ,
		\a[39] ,
		\shift[0] ,
		\shift[1] ,
		_w344_
	);
	LUT3 #(
		.INIT('ha8)
	) name208 (
		_w149_,
		_w343_,
		_w344_,
		_w345_
	);
	LUT4 #(
		.INIT('h0001)
	) name209 (
		_w336_,
		_w339_,
		_w342_,
		_w345_,
		_w346_
	);
	LUT4 #(
		.INIT('ha00c)
	) name210 (
		\a[30] ,
		\a[33] ,
		\shift[0] ,
		\shift[1] ,
		_w347_
	);
	LUT4 #(
		.INIT('hf53f)
	) name211 (
		\a[31] ,
		\a[32] ,
		\shift[0] ,
		\shift[1] ,
		_w348_
	);
	LUT3 #(
		.INIT('h8a)
	) name212 (
		_w137_,
		_w347_,
		_w348_,
		_w349_
	);
	LUT4 #(
		.INIT('ha00c)
	) name213 (
		\a[26] ,
		\a[29] ,
		\shift[0] ,
		\shift[1] ,
		_w350_
	);
	LUT4 #(
		.INIT('hf53f)
	) name214 (
		\a[27] ,
		\a[28] ,
		\shift[0] ,
		\shift[1] ,
		_w351_
	);
	LUT3 #(
		.INIT('h8a)
	) name215 (
		_w141_,
		_w350_,
		_w351_,
		_w352_
	);
	LUT4 #(
		.INIT('ha00c)
	) name216 (
		\a[18] ,
		\a[21] ,
		\shift[0] ,
		\shift[1] ,
		_w353_
	);
	LUT4 #(
		.INIT('hf53f)
	) name217 (
		\a[19] ,
		\a[20] ,
		\shift[0] ,
		\shift[1] ,
		_w354_
	);
	LUT3 #(
		.INIT('h8a)
	) name218 (
		_w145_,
		_w353_,
		_w354_,
		_w355_
	);
	LUT4 #(
		.INIT('ha00c)
	) name219 (
		\a[22] ,
		\a[25] ,
		\shift[0] ,
		\shift[1] ,
		_w356_
	);
	LUT4 #(
		.INIT('hf53f)
	) name220 (
		\a[23] ,
		\a[24] ,
		\shift[0] ,
		\shift[1] ,
		_w357_
	);
	LUT3 #(
		.INIT('h8a)
	) name221 (
		_w149_,
		_w356_,
		_w357_,
		_w358_
	);
	LUT4 #(
		.INIT('h0001)
	) name222 (
		_w349_,
		_w352_,
		_w355_,
		_w358_,
		_w359_
	);
	LUT4 #(
		.INIT('hfdb9)
	) name223 (
		\shift[4] ,
		\shift[5] ,
		_w346_,
		_w359_,
		_w360_
	);
	LUT3 #(
		.INIT('h2a)
	) name224 (
		\shift[6] ,
		_w333_,
		_w360_,
		_w361_
	);
	LUT2 #(
		.INIT('he)
	) name225 (
		_w306_,
		_w361_,
		_w362_
	);
	LUT4 #(
		.INIT('hac00)
	) name226 (
		\a[79] ,
		\a[80] ,
		\shift[0] ,
		\shift[1] ,
		_w363_
	);
	LUT4 #(
		.INIT('h00ac)
	) name227 (
		\a[81] ,
		\a[82] ,
		\shift[0] ,
		\shift[1] ,
		_w364_
	);
	LUT3 #(
		.INIT('ha8)
	) name228 (
		_w137_,
		_w363_,
		_w364_,
		_w365_
	);
	LUT4 #(
		.INIT('hac00)
	) name229 (
		\a[75] ,
		\a[76] ,
		\shift[0] ,
		\shift[1] ,
		_w366_
	);
	LUT4 #(
		.INIT('h00ac)
	) name230 (
		\a[77] ,
		\a[78] ,
		\shift[0] ,
		\shift[1] ,
		_w367_
	);
	LUT3 #(
		.INIT('ha8)
	) name231 (
		_w141_,
		_w366_,
		_w367_,
		_w368_
	);
	LUT4 #(
		.INIT('hac00)
	) name232 (
		\a[67] ,
		\a[68] ,
		\shift[0] ,
		\shift[1] ,
		_w369_
	);
	LUT4 #(
		.INIT('h00ac)
	) name233 (
		\a[69] ,
		\a[70] ,
		\shift[0] ,
		\shift[1] ,
		_w370_
	);
	LUT3 #(
		.INIT('ha8)
	) name234 (
		_w145_,
		_w369_,
		_w370_,
		_w371_
	);
	LUT4 #(
		.INIT('hac00)
	) name235 (
		\a[71] ,
		\a[72] ,
		\shift[0] ,
		\shift[1] ,
		_w372_
	);
	LUT4 #(
		.INIT('h00ac)
	) name236 (
		\a[73] ,
		\a[74] ,
		\shift[0] ,
		\shift[1] ,
		_w373_
	);
	LUT3 #(
		.INIT('ha8)
	) name237 (
		_w149_,
		_w372_,
		_w373_,
		_w374_
	);
	LUT4 #(
		.INIT('h0001)
	) name238 (
		_w365_,
		_w368_,
		_w371_,
		_w374_,
		_w375_
	);
	LUT4 #(
		.INIT('hac00)
	) name239 (
		\a[95] ,
		\a[96] ,
		\shift[0] ,
		\shift[1] ,
		_w376_
	);
	LUT4 #(
		.INIT('h00ac)
	) name240 (
		\a[97] ,
		\a[98] ,
		\shift[0] ,
		\shift[1] ,
		_w377_
	);
	LUT3 #(
		.INIT('ha8)
	) name241 (
		_w137_,
		_w376_,
		_w377_,
		_w378_
	);
	LUT4 #(
		.INIT('hac00)
	) name242 (
		\a[91] ,
		\a[92] ,
		\shift[0] ,
		\shift[1] ,
		_w379_
	);
	LUT4 #(
		.INIT('h00ac)
	) name243 (
		\a[93] ,
		\a[94] ,
		\shift[0] ,
		\shift[1] ,
		_w380_
	);
	LUT3 #(
		.INIT('ha8)
	) name244 (
		_w141_,
		_w379_,
		_w380_,
		_w381_
	);
	LUT4 #(
		.INIT('hac00)
	) name245 (
		\a[83] ,
		\a[84] ,
		\shift[0] ,
		\shift[1] ,
		_w382_
	);
	LUT4 #(
		.INIT('h00ac)
	) name246 (
		\a[85] ,
		\a[86] ,
		\shift[0] ,
		\shift[1] ,
		_w383_
	);
	LUT3 #(
		.INIT('ha8)
	) name247 (
		_w145_,
		_w382_,
		_w383_,
		_w384_
	);
	LUT4 #(
		.INIT('hac00)
	) name248 (
		\a[87] ,
		\a[88] ,
		\shift[0] ,
		\shift[1] ,
		_w385_
	);
	LUT4 #(
		.INIT('h00ac)
	) name249 (
		\a[89] ,
		\a[90] ,
		\shift[0] ,
		\shift[1] ,
		_w386_
	);
	LUT3 #(
		.INIT('ha8)
	) name250 (
		_w149_,
		_w385_,
		_w386_,
		_w387_
	);
	LUT4 #(
		.INIT('h0001)
	) name251 (
		_w378_,
		_w381_,
		_w384_,
		_w387_,
		_w388_
	);
	LUT4 #(
		.INIT('hf7b3)
	) name252 (
		\shift[4] ,
		\shift[5] ,
		_w375_,
		_w388_,
		_w389_
	);
	LUT4 #(
		.INIT('hca00)
	) name253 (
		\a[0] ,
		\a[127] ,
		\shift[0] ,
		\shift[1] ,
		_w390_
	);
	LUT4 #(
		.INIT('h00ac)
	) name254 (
		\a[1] ,
		\a[2] ,
		\shift[0] ,
		\shift[1] ,
		_w391_
	);
	LUT3 #(
		.INIT('ha8)
	) name255 (
		_w137_,
		_w390_,
		_w391_,
		_w392_
	);
	LUT4 #(
		.INIT('hac00)
	) name256 (
		\a[123] ,
		\a[124] ,
		\shift[0] ,
		\shift[1] ,
		_w393_
	);
	LUT4 #(
		.INIT('h00ac)
	) name257 (
		\a[125] ,
		\a[126] ,
		\shift[0] ,
		\shift[1] ,
		_w394_
	);
	LUT3 #(
		.INIT('ha8)
	) name258 (
		_w141_,
		_w393_,
		_w394_,
		_w395_
	);
	LUT4 #(
		.INIT('hac00)
	) name259 (
		\a[115] ,
		\a[116] ,
		\shift[0] ,
		\shift[1] ,
		_w396_
	);
	LUT4 #(
		.INIT('h00ac)
	) name260 (
		\a[117] ,
		\a[118] ,
		\shift[0] ,
		\shift[1] ,
		_w397_
	);
	LUT3 #(
		.INIT('ha8)
	) name261 (
		_w145_,
		_w396_,
		_w397_,
		_w398_
	);
	LUT4 #(
		.INIT('hac00)
	) name262 (
		\a[119] ,
		\a[120] ,
		\shift[0] ,
		\shift[1] ,
		_w399_
	);
	LUT4 #(
		.INIT('h00ac)
	) name263 (
		\a[121] ,
		\a[122] ,
		\shift[0] ,
		\shift[1] ,
		_w400_
	);
	LUT3 #(
		.INIT('ha8)
	) name264 (
		_w149_,
		_w399_,
		_w400_,
		_w401_
	);
	LUT4 #(
		.INIT('h0001)
	) name265 (
		_w392_,
		_w395_,
		_w398_,
		_w401_,
		_w402_
	);
	LUT4 #(
		.INIT('hac00)
	) name266 (
		\a[111] ,
		\a[112] ,
		\shift[0] ,
		\shift[1] ,
		_w403_
	);
	LUT4 #(
		.INIT('h00ac)
	) name267 (
		\a[113] ,
		\a[114] ,
		\shift[0] ,
		\shift[1] ,
		_w404_
	);
	LUT3 #(
		.INIT('ha8)
	) name268 (
		_w137_,
		_w403_,
		_w404_,
		_w405_
	);
	LUT4 #(
		.INIT('hac00)
	) name269 (
		\a[107] ,
		\a[108] ,
		\shift[0] ,
		\shift[1] ,
		_w406_
	);
	LUT4 #(
		.INIT('h00ac)
	) name270 (
		\a[109] ,
		\a[110] ,
		\shift[0] ,
		\shift[1] ,
		_w407_
	);
	LUT3 #(
		.INIT('ha8)
	) name271 (
		_w141_,
		_w406_,
		_w407_,
		_w408_
	);
	LUT4 #(
		.INIT('hac00)
	) name272 (
		\a[99] ,
		\a[100] ,
		\shift[0] ,
		\shift[1] ,
		_w409_
	);
	LUT4 #(
		.INIT('h00ac)
	) name273 (
		\a[101] ,
		\a[102] ,
		\shift[0] ,
		\shift[1] ,
		_w410_
	);
	LUT3 #(
		.INIT('ha8)
	) name274 (
		_w145_,
		_w409_,
		_w410_,
		_w411_
	);
	LUT4 #(
		.INIT('hac00)
	) name275 (
		\a[103] ,
		\a[104] ,
		\shift[0] ,
		\shift[1] ,
		_w412_
	);
	LUT4 #(
		.INIT('h00ac)
	) name276 (
		\a[105] ,
		\a[106] ,
		\shift[0] ,
		\shift[1] ,
		_w413_
	);
	LUT3 #(
		.INIT('ha8)
	) name277 (
		_w149_,
		_w412_,
		_w413_,
		_w414_
	);
	LUT4 #(
		.INIT('h0001)
	) name278 (
		_w405_,
		_w408_,
		_w411_,
		_w414_,
		_w415_
	);
	LUT4 #(
		.INIT('hfedc)
	) name279 (
		\shift[4] ,
		\shift[5] ,
		_w402_,
		_w415_,
		_w416_
	);
	LUT3 #(
		.INIT('h15)
	) name280 (
		\shift[6] ,
		_w389_,
		_w416_,
		_w417_
	);
	LUT4 #(
		.INIT('hac00)
	) name281 (
		\a[63] ,
		\a[64] ,
		\shift[0] ,
		\shift[1] ,
		_w418_
	);
	LUT4 #(
		.INIT('h00ac)
	) name282 (
		\a[65] ,
		\a[66] ,
		\shift[0] ,
		\shift[1] ,
		_w419_
	);
	LUT3 #(
		.INIT('ha8)
	) name283 (
		_w137_,
		_w418_,
		_w419_,
		_w420_
	);
	LUT4 #(
		.INIT('hac00)
	) name284 (
		\a[59] ,
		\a[60] ,
		\shift[0] ,
		\shift[1] ,
		_w421_
	);
	LUT4 #(
		.INIT('h00ac)
	) name285 (
		\a[61] ,
		\a[62] ,
		\shift[0] ,
		\shift[1] ,
		_w422_
	);
	LUT3 #(
		.INIT('ha8)
	) name286 (
		_w141_,
		_w421_,
		_w422_,
		_w423_
	);
	LUT4 #(
		.INIT('hac00)
	) name287 (
		\a[51] ,
		\a[52] ,
		\shift[0] ,
		\shift[1] ,
		_w424_
	);
	LUT4 #(
		.INIT('h00ac)
	) name288 (
		\a[53] ,
		\a[54] ,
		\shift[0] ,
		\shift[1] ,
		_w425_
	);
	LUT3 #(
		.INIT('ha8)
	) name289 (
		_w145_,
		_w424_,
		_w425_,
		_w426_
	);
	LUT4 #(
		.INIT('hac00)
	) name290 (
		\a[55] ,
		\a[56] ,
		\shift[0] ,
		\shift[1] ,
		_w427_
	);
	LUT4 #(
		.INIT('h00ac)
	) name291 (
		\a[57] ,
		\a[58] ,
		\shift[0] ,
		\shift[1] ,
		_w428_
	);
	LUT3 #(
		.INIT('ha8)
	) name292 (
		_w149_,
		_w427_,
		_w428_,
		_w429_
	);
	LUT4 #(
		.INIT('h0001)
	) name293 (
		_w420_,
		_w423_,
		_w426_,
		_w429_,
		_w430_
	);
	LUT4 #(
		.INIT('hac00)
	) name294 (
		\a[15] ,
		\a[16] ,
		\shift[0] ,
		\shift[1] ,
		_w431_
	);
	LUT4 #(
		.INIT('h00ac)
	) name295 (
		\a[17] ,
		\a[18] ,
		\shift[0] ,
		\shift[1] ,
		_w432_
	);
	LUT3 #(
		.INIT('ha8)
	) name296 (
		_w137_,
		_w431_,
		_w432_,
		_w433_
	);
	LUT4 #(
		.INIT('hac00)
	) name297 (
		\a[11] ,
		\a[12] ,
		\shift[0] ,
		\shift[1] ,
		_w434_
	);
	LUT4 #(
		.INIT('h00ac)
	) name298 (
		\a[13] ,
		\a[14] ,
		\shift[0] ,
		\shift[1] ,
		_w435_
	);
	LUT3 #(
		.INIT('ha8)
	) name299 (
		_w141_,
		_w434_,
		_w435_,
		_w436_
	);
	LUT4 #(
		.INIT('hac00)
	) name300 (
		\a[3] ,
		\a[4] ,
		\shift[0] ,
		\shift[1] ,
		_w437_
	);
	LUT4 #(
		.INIT('h00ac)
	) name301 (
		\a[5] ,
		\a[6] ,
		\shift[0] ,
		\shift[1] ,
		_w438_
	);
	LUT3 #(
		.INIT('ha8)
	) name302 (
		_w145_,
		_w437_,
		_w438_,
		_w439_
	);
	LUT4 #(
		.INIT('hac00)
	) name303 (
		\a[7] ,
		\a[8] ,
		\shift[0] ,
		\shift[1] ,
		_w440_
	);
	LUT4 #(
		.INIT('h00ac)
	) name304 (
		\a[9] ,
		\a[10] ,
		\shift[0] ,
		\shift[1] ,
		_w441_
	);
	LUT3 #(
		.INIT('ha8)
	) name305 (
		_w149_,
		_w440_,
		_w441_,
		_w442_
	);
	LUT4 #(
		.INIT('h0001)
	) name306 (
		_w433_,
		_w436_,
		_w439_,
		_w442_,
		_w443_
	);
	LUT4 #(
		.INIT('hfe76)
	) name307 (
		\shift[4] ,
		\shift[5] ,
		_w430_,
		_w443_,
		_w444_
	);
	LUT4 #(
		.INIT('hac00)
	) name308 (
		\a[47] ,
		\a[48] ,
		\shift[0] ,
		\shift[1] ,
		_w445_
	);
	LUT4 #(
		.INIT('h00ac)
	) name309 (
		\a[49] ,
		\a[50] ,
		\shift[0] ,
		\shift[1] ,
		_w446_
	);
	LUT3 #(
		.INIT('ha8)
	) name310 (
		_w137_,
		_w445_,
		_w446_,
		_w447_
	);
	LUT4 #(
		.INIT('hac00)
	) name311 (
		\a[43] ,
		\a[44] ,
		\shift[0] ,
		\shift[1] ,
		_w448_
	);
	LUT4 #(
		.INIT('h00ac)
	) name312 (
		\a[45] ,
		\a[46] ,
		\shift[0] ,
		\shift[1] ,
		_w449_
	);
	LUT3 #(
		.INIT('ha8)
	) name313 (
		_w141_,
		_w448_,
		_w449_,
		_w450_
	);
	LUT4 #(
		.INIT('h00ac)
	) name314 (
		\a[37] ,
		\a[38] ,
		\shift[0] ,
		\shift[1] ,
		_w451_
	);
	LUT4 #(
		.INIT('hac00)
	) name315 (
		\a[35] ,
		\a[36] ,
		\shift[0] ,
		\shift[1] ,
		_w452_
	);
	LUT3 #(
		.INIT('ha8)
	) name316 (
		_w145_,
		_w451_,
		_w452_,
		_w453_
	);
	LUT4 #(
		.INIT('h00ac)
	) name317 (
		\a[41] ,
		\a[42] ,
		\shift[0] ,
		\shift[1] ,
		_w454_
	);
	LUT4 #(
		.INIT('hac00)
	) name318 (
		\a[39] ,
		\a[40] ,
		\shift[0] ,
		\shift[1] ,
		_w455_
	);
	LUT3 #(
		.INIT('ha8)
	) name319 (
		_w149_,
		_w454_,
		_w455_,
		_w456_
	);
	LUT4 #(
		.INIT('h0001)
	) name320 (
		_w447_,
		_w450_,
		_w453_,
		_w456_,
		_w457_
	);
	LUT4 #(
		.INIT('hac00)
	) name321 (
		\a[31] ,
		\a[32] ,
		\shift[0] ,
		\shift[1] ,
		_w458_
	);
	LUT4 #(
		.INIT('h00ac)
	) name322 (
		\a[33] ,
		\a[34] ,
		\shift[0] ,
		\shift[1] ,
		_w459_
	);
	LUT3 #(
		.INIT('ha8)
	) name323 (
		_w137_,
		_w458_,
		_w459_,
		_w460_
	);
	LUT4 #(
		.INIT('hac00)
	) name324 (
		\a[27] ,
		\a[28] ,
		\shift[0] ,
		\shift[1] ,
		_w461_
	);
	LUT4 #(
		.INIT('h00ac)
	) name325 (
		\a[29] ,
		\a[30] ,
		\shift[0] ,
		\shift[1] ,
		_w462_
	);
	LUT3 #(
		.INIT('ha8)
	) name326 (
		_w141_,
		_w461_,
		_w462_,
		_w463_
	);
	LUT4 #(
		.INIT('hac00)
	) name327 (
		\a[19] ,
		\a[20] ,
		\shift[0] ,
		\shift[1] ,
		_w464_
	);
	LUT4 #(
		.INIT('h00ac)
	) name328 (
		\a[21] ,
		\a[22] ,
		\shift[0] ,
		\shift[1] ,
		_w465_
	);
	LUT3 #(
		.INIT('ha8)
	) name329 (
		_w145_,
		_w464_,
		_w465_,
		_w466_
	);
	LUT4 #(
		.INIT('hac00)
	) name330 (
		\a[23] ,
		\a[24] ,
		\shift[0] ,
		\shift[1] ,
		_w467_
	);
	LUT4 #(
		.INIT('h00ac)
	) name331 (
		\a[25] ,
		\a[26] ,
		\shift[0] ,
		\shift[1] ,
		_w468_
	);
	LUT3 #(
		.INIT('ha8)
	) name332 (
		_w149_,
		_w467_,
		_w468_,
		_w469_
	);
	LUT4 #(
		.INIT('h0001)
	) name333 (
		_w460_,
		_w463_,
		_w466_,
		_w469_,
		_w470_
	);
	LUT4 #(
		.INIT('hfdb9)
	) name334 (
		\shift[4] ,
		\shift[5] ,
		_w457_,
		_w470_,
		_w471_
	);
	LUT3 #(
		.INIT('h2a)
	) name335 (
		\shift[6] ,
		_w444_,
		_w471_,
		_w472_
	);
	LUT2 #(
		.INIT('he)
	) name336 (
		_w417_,
		_w472_,
		_w473_
	);
	LUT4 #(
		.INIT('h0ac0)
	) name337 (
		\a[113] ,
		\a[114] ,
		\shift[0] ,
		\shift[1] ,
		_w474_
	);
	LUT4 #(
		.INIT('h5ff3)
	) name338 (
		\a[112] ,
		\a[115] ,
		\shift[0] ,
		\shift[1] ,
		_w475_
	);
	LUT3 #(
		.INIT('h8a)
	) name339 (
		_w137_,
		_w474_,
		_w475_,
		_w476_
	);
	LUT4 #(
		.INIT('h0ac0)
	) name340 (
		\a[109] ,
		\a[110] ,
		\shift[0] ,
		\shift[1] ,
		_w477_
	);
	LUT4 #(
		.INIT('h5ff3)
	) name341 (
		\a[108] ,
		\a[111] ,
		\shift[0] ,
		\shift[1] ,
		_w478_
	);
	LUT3 #(
		.INIT('h8a)
	) name342 (
		_w141_,
		_w477_,
		_w478_,
		_w479_
	);
	LUT4 #(
		.INIT('h0ac0)
	) name343 (
		\a[101] ,
		\a[102] ,
		\shift[0] ,
		\shift[1] ,
		_w480_
	);
	LUT4 #(
		.INIT('h5ff3)
	) name344 (
		\a[100] ,
		\a[103] ,
		\shift[0] ,
		\shift[1] ,
		_w481_
	);
	LUT3 #(
		.INIT('h8a)
	) name345 (
		_w145_,
		_w480_,
		_w481_,
		_w482_
	);
	LUT4 #(
		.INIT('h0ac0)
	) name346 (
		\a[105] ,
		\a[106] ,
		\shift[0] ,
		\shift[1] ,
		_w483_
	);
	LUT4 #(
		.INIT('h5ff3)
	) name347 (
		\a[104] ,
		\a[107] ,
		\shift[0] ,
		\shift[1] ,
		_w484_
	);
	LUT3 #(
		.INIT('h8a)
	) name348 (
		_w149_,
		_w483_,
		_w484_,
		_w485_
	);
	LUT4 #(
		.INIT('h0001)
	) name349 (
		_w476_,
		_w479_,
		_w482_,
		_w485_,
		_w486_
	);
	LUT4 #(
		.INIT('h0ac0)
	) name350 (
		\a[97] ,
		\a[98] ,
		\shift[0] ,
		\shift[1] ,
		_w487_
	);
	LUT4 #(
		.INIT('h5ff3)
	) name351 (
		\a[96] ,
		\a[99] ,
		\shift[0] ,
		\shift[1] ,
		_w488_
	);
	LUT3 #(
		.INIT('h8a)
	) name352 (
		_w137_,
		_w487_,
		_w488_,
		_w489_
	);
	LUT4 #(
		.INIT('h0ac0)
	) name353 (
		\a[93] ,
		\a[94] ,
		\shift[0] ,
		\shift[1] ,
		_w490_
	);
	LUT4 #(
		.INIT('h5ff3)
	) name354 (
		\a[92] ,
		\a[95] ,
		\shift[0] ,
		\shift[1] ,
		_w491_
	);
	LUT3 #(
		.INIT('h8a)
	) name355 (
		_w141_,
		_w490_,
		_w491_,
		_w492_
	);
	LUT4 #(
		.INIT('h0ac0)
	) name356 (
		\a[85] ,
		\a[86] ,
		\shift[0] ,
		\shift[1] ,
		_w493_
	);
	LUT4 #(
		.INIT('h5ff3)
	) name357 (
		\a[84] ,
		\a[87] ,
		\shift[0] ,
		\shift[1] ,
		_w494_
	);
	LUT3 #(
		.INIT('h8a)
	) name358 (
		_w145_,
		_w493_,
		_w494_,
		_w495_
	);
	LUT4 #(
		.INIT('h0ac0)
	) name359 (
		\a[89] ,
		\a[90] ,
		\shift[0] ,
		\shift[1] ,
		_w496_
	);
	LUT4 #(
		.INIT('h5ff3)
	) name360 (
		\a[88] ,
		\a[91] ,
		\shift[0] ,
		\shift[1] ,
		_w497_
	);
	LUT3 #(
		.INIT('h8a)
	) name361 (
		_w149_,
		_w496_,
		_w497_,
		_w498_
	);
	LUT4 #(
		.INIT('h0001)
	) name362 (
		_w489_,
		_w492_,
		_w495_,
		_w498_,
		_w499_
	);
	LUT4 #(
		.INIT('hfdb9)
	) name363 (
		\shift[4] ,
		\shift[5] ,
		_w486_,
		_w499_,
		_w500_
	);
	LUT4 #(
		.INIT('h0ac0)
	) name364 (
		\a[1] ,
		\a[2] ,
		\shift[0] ,
		\shift[1] ,
		_w501_
	);
	LUT4 #(
		.INIT('h5ff3)
	) name365 (
		\a[0] ,
		\a[3] ,
		\shift[0] ,
		\shift[1] ,
		_w502_
	);
	LUT3 #(
		.INIT('h8a)
	) name366 (
		_w137_,
		_w501_,
		_w502_,
		_w503_
	);
	LUT4 #(
		.INIT('h0ac0)
	) name367 (
		\a[125] ,
		\a[126] ,
		\shift[0] ,
		\shift[1] ,
		_w504_
	);
	LUT4 #(
		.INIT('h5ff3)
	) name368 (
		\a[124] ,
		\a[127] ,
		\shift[0] ,
		\shift[1] ,
		_w505_
	);
	LUT3 #(
		.INIT('h8a)
	) name369 (
		_w141_,
		_w504_,
		_w505_,
		_w506_
	);
	LUT4 #(
		.INIT('h0ac0)
	) name370 (
		\a[117] ,
		\a[118] ,
		\shift[0] ,
		\shift[1] ,
		_w507_
	);
	LUT4 #(
		.INIT('h5ff3)
	) name371 (
		\a[116] ,
		\a[119] ,
		\shift[0] ,
		\shift[1] ,
		_w508_
	);
	LUT3 #(
		.INIT('h8a)
	) name372 (
		_w145_,
		_w507_,
		_w508_,
		_w509_
	);
	LUT4 #(
		.INIT('h0ac0)
	) name373 (
		\a[121] ,
		\a[122] ,
		\shift[0] ,
		\shift[1] ,
		_w510_
	);
	LUT4 #(
		.INIT('h5ff3)
	) name374 (
		\a[120] ,
		\a[123] ,
		\shift[0] ,
		\shift[1] ,
		_w511_
	);
	LUT3 #(
		.INIT('h8a)
	) name375 (
		_w149_,
		_w510_,
		_w511_,
		_w512_
	);
	LUT4 #(
		.INIT('h0001)
	) name376 (
		_w503_,
		_w506_,
		_w509_,
		_w512_,
		_w513_
	);
	LUT4 #(
		.INIT('h0ac0)
	) name377 (
		\a[81] ,
		\a[82] ,
		\shift[0] ,
		\shift[1] ,
		_w514_
	);
	LUT4 #(
		.INIT('h5ff3)
	) name378 (
		\a[80] ,
		\a[83] ,
		\shift[0] ,
		\shift[1] ,
		_w515_
	);
	LUT3 #(
		.INIT('h8a)
	) name379 (
		_w137_,
		_w514_,
		_w515_,
		_w516_
	);
	LUT4 #(
		.INIT('h0ac0)
	) name380 (
		\a[77] ,
		\a[78] ,
		\shift[0] ,
		\shift[1] ,
		_w517_
	);
	LUT4 #(
		.INIT('h5ff3)
	) name381 (
		\a[76] ,
		\a[79] ,
		\shift[0] ,
		\shift[1] ,
		_w518_
	);
	LUT3 #(
		.INIT('h8a)
	) name382 (
		_w141_,
		_w517_,
		_w518_,
		_w519_
	);
	LUT4 #(
		.INIT('h0ac0)
	) name383 (
		\a[69] ,
		\a[70] ,
		\shift[0] ,
		\shift[1] ,
		_w520_
	);
	LUT4 #(
		.INIT('h5ff3)
	) name384 (
		\a[68] ,
		\a[71] ,
		\shift[0] ,
		\shift[1] ,
		_w521_
	);
	LUT3 #(
		.INIT('h8a)
	) name385 (
		_w145_,
		_w520_,
		_w521_,
		_w522_
	);
	LUT4 #(
		.INIT('h0ac0)
	) name386 (
		\a[73] ,
		\a[74] ,
		\shift[0] ,
		\shift[1] ,
		_w523_
	);
	LUT4 #(
		.INIT('h5ff3)
	) name387 (
		\a[72] ,
		\a[75] ,
		\shift[0] ,
		\shift[1] ,
		_w524_
	);
	LUT3 #(
		.INIT('h8a)
	) name388 (
		_w149_,
		_w523_,
		_w524_,
		_w525_
	);
	LUT4 #(
		.INIT('h0001)
	) name389 (
		_w516_,
		_w519_,
		_w522_,
		_w525_,
		_w526_
	);
	LUT4 #(
		.INIT('hfe76)
	) name390 (
		\shift[4] ,
		\shift[5] ,
		_w513_,
		_w526_,
		_w527_
	);
	LUT3 #(
		.INIT('h15)
	) name391 (
		\shift[6] ,
		_w500_,
		_w527_,
		_w528_
	);
	LUT4 #(
		.INIT('h0ac0)
	) name392 (
		\a[65] ,
		\a[66] ,
		\shift[0] ,
		\shift[1] ,
		_w529_
	);
	LUT4 #(
		.INIT('h5ff3)
	) name393 (
		\a[64] ,
		\a[67] ,
		\shift[0] ,
		\shift[1] ,
		_w530_
	);
	LUT3 #(
		.INIT('h8a)
	) name394 (
		_w137_,
		_w529_,
		_w530_,
		_w531_
	);
	LUT4 #(
		.INIT('h0ac0)
	) name395 (
		\a[61] ,
		\a[62] ,
		\shift[0] ,
		\shift[1] ,
		_w532_
	);
	LUT4 #(
		.INIT('h5ff3)
	) name396 (
		\a[60] ,
		\a[63] ,
		\shift[0] ,
		\shift[1] ,
		_w533_
	);
	LUT3 #(
		.INIT('h8a)
	) name397 (
		_w141_,
		_w532_,
		_w533_,
		_w534_
	);
	LUT4 #(
		.INIT('h0ac0)
	) name398 (
		\a[53] ,
		\a[54] ,
		\shift[0] ,
		\shift[1] ,
		_w535_
	);
	LUT4 #(
		.INIT('h5ff3)
	) name399 (
		\a[52] ,
		\a[55] ,
		\shift[0] ,
		\shift[1] ,
		_w536_
	);
	LUT3 #(
		.INIT('h8a)
	) name400 (
		_w145_,
		_w535_,
		_w536_,
		_w537_
	);
	LUT4 #(
		.INIT('h0ac0)
	) name401 (
		\a[57] ,
		\a[58] ,
		\shift[0] ,
		\shift[1] ,
		_w538_
	);
	LUT4 #(
		.INIT('h5ff3)
	) name402 (
		\a[56] ,
		\a[59] ,
		\shift[0] ,
		\shift[1] ,
		_w539_
	);
	LUT3 #(
		.INIT('h8a)
	) name403 (
		_w149_,
		_w538_,
		_w539_,
		_w540_
	);
	LUT4 #(
		.INIT('h0001)
	) name404 (
		_w531_,
		_w534_,
		_w537_,
		_w540_,
		_w541_
	);
	LUT4 #(
		.INIT('h0ac0)
	) name405 (
		\a[49] ,
		\a[50] ,
		\shift[0] ,
		\shift[1] ,
		_w542_
	);
	LUT4 #(
		.INIT('h5ff3)
	) name406 (
		\a[48] ,
		\a[51] ,
		\shift[0] ,
		\shift[1] ,
		_w543_
	);
	LUT3 #(
		.INIT('h8a)
	) name407 (
		_w137_,
		_w542_,
		_w543_,
		_w544_
	);
	LUT4 #(
		.INIT('hac00)
	) name408 (
		\a[44] ,
		\a[45] ,
		\shift[0] ,
		\shift[1] ,
		_w545_
	);
	LUT4 #(
		.INIT('h00ac)
	) name409 (
		\a[46] ,
		\a[47] ,
		\shift[0] ,
		\shift[1] ,
		_w546_
	);
	LUT3 #(
		.INIT('ha8)
	) name410 (
		_w141_,
		_w545_,
		_w546_,
		_w547_
	);
	LUT4 #(
		.INIT('h0ac0)
	) name411 (
		\a[37] ,
		\a[38] ,
		\shift[0] ,
		\shift[1] ,
		_w548_
	);
	LUT4 #(
		.INIT('h5ff3)
	) name412 (
		\a[36] ,
		\a[39] ,
		\shift[0] ,
		\shift[1] ,
		_w549_
	);
	LUT3 #(
		.INIT('h8a)
	) name413 (
		_w145_,
		_w548_,
		_w549_,
		_w550_
	);
	LUT4 #(
		.INIT('h0ac0)
	) name414 (
		\a[41] ,
		\a[42] ,
		\shift[0] ,
		\shift[1] ,
		_w551_
	);
	LUT4 #(
		.INIT('h5ff3)
	) name415 (
		\a[40] ,
		\a[43] ,
		\shift[0] ,
		\shift[1] ,
		_w552_
	);
	LUT3 #(
		.INIT('h8a)
	) name416 (
		_w149_,
		_w551_,
		_w552_,
		_w553_
	);
	LUT4 #(
		.INIT('h0001)
	) name417 (
		_w544_,
		_w547_,
		_w550_,
		_w553_,
		_w554_
	);
	LUT4 #(
		.INIT('hfedc)
	) name418 (
		\shift[4] ,
		\shift[5] ,
		_w541_,
		_w554_,
		_w555_
	);
	LUT4 #(
		.INIT('h0ac0)
	) name419 (
		\a[17] ,
		\a[18] ,
		\shift[0] ,
		\shift[1] ,
		_w556_
	);
	LUT4 #(
		.INIT('h5ff3)
	) name420 (
		\a[16] ,
		\a[19] ,
		\shift[0] ,
		\shift[1] ,
		_w557_
	);
	LUT3 #(
		.INIT('h8a)
	) name421 (
		_w137_,
		_w556_,
		_w557_,
		_w558_
	);
	LUT4 #(
		.INIT('h0ac0)
	) name422 (
		\a[13] ,
		\a[14] ,
		\shift[0] ,
		\shift[1] ,
		_w559_
	);
	LUT4 #(
		.INIT('h5ff3)
	) name423 (
		\a[12] ,
		\a[15] ,
		\shift[0] ,
		\shift[1] ,
		_w560_
	);
	LUT3 #(
		.INIT('h8a)
	) name424 (
		_w141_,
		_w559_,
		_w560_,
		_w561_
	);
	LUT4 #(
		.INIT('h0ac0)
	) name425 (
		\a[5] ,
		\a[6] ,
		\shift[0] ,
		\shift[1] ,
		_w562_
	);
	LUT4 #(
		.INIT('h5ff3)
	) name426 (
		\a[4] ,
		\a[7] ,
		\shift[0] ,
		\shift[1] ,
		_w563_
	);
	LUT3 #(
		.INIT('h8a)
	) name427 (
		_w145_,
		_w562_,
		_w563_,
		_w564_
	);
	LUT4 #(
		.INIT('h0ac0)
	) name428 (
		\a[9] ,
		\a[10] ,
		\shift[0] ,
		\shift[1] ,
		_w565_
	);
	LUT4 #(
		.INIT('h5ff3)
	) name429 (
		\a[8] ,
		\a[11] ,
		\shift[0] ,
		\shift[1] ,
		_w566_
	);
	LUT3 #(
		.INIT('h8a)
	) name430 (
		_w149_,
		_w565_,
		_w566_,
		_w567_
	);
	LUT4 #(
		.INIT('h0001)
	) name431 (
		_w558_,
		_w561_,
		_w564_,
		_w567_,
		_w568_
	);
	LUT4 #(
		.INIT('h0ac0)
	) name432 (
		\a[33] ,
		\a[34] ,
		\shift[0] ,
		\shift[1] ,
		_w569_
	);
	LUT4 #(
		.INIT('h5ff3)
	) name433 (
		\a[32] ,
		\a[35] ,
		\shift[0] ,
		\shift[1] ,
		_w570_
	);
	LUT3 #(
		.INIT('h8a)
	) name434 (
		_w137_,
		_w569_,
		_w570_,
		_w571_
	);
	LUT4 #(
		.INIT('h0ac0)
	) name435 (
		\a[29] ,
		\a[30] ,
		\shift[0] ,
		\shift[1] ,
		_w572_
	);
	LUT4 #(
		.INIT('h5ff3)
	) name436 (
		\a[28] ,
		\a[31] ,
		\shift[0] ,
		\shift[1] ,
		_w573_
	);
	LUT3 #(
		.INIT('h8a)
	) name437 (
		_w141_,
		_w572_,
		_w573_,
		_w574_
	);
	LUT4 #(
		.INIT('h0ac0)
	) name438 (
		\a[21] ,
		\a[22] ,
		\shift[0] ,
		\shift[1] ,
		_w575_
	);
	LUT4 #(
		.INIT('h5ff3)
	) name439 (
		\a[20] ,
		\a[23] ,
		\shift[0] ,
		\shift[1] ,
		_w576_
	);
	LUT3 #(
		.INIT('h8a)
	) name440 (
		_w145_,
		_w575_,
		_w576_,
		_w577_
	);
	LUT4 #(
		.INIT('h0ac0)
	) name441 (
		\a[25] ,
		\a[26] ,
		\shift[0] ,
		\shift[1] ,
		_w578_
	);
	LUT4 #(
		.INIT('h5ff3)
	) name442 (
		\a[24] ,
		\a[27] ,
		\shift[0] ,
		\shift[1] ,
		_w579_
	);
	LUT3 #(
		.INIT('h8a)
	) name443 (
		_w149_,
		_w578_,
		_w579_,
		_w580_
	);
	LUT4 #(
		.INIT('h0001)
	) name444 (
		_w571_,
		_w574_,
		_w577_,
		_w580_,
		_w581_
	);
	LUT4 #(
		.INIT('hf7b3)
	) name445 (
		\shift[4] ,
		\shift[5] ,
		_w568_,
		_w581_,
		_w582_
	);
	LUT3 #(
		.INIT('h2a)
	) name446 (
		\shift[6] ,
		_w555_,
		_w582_,
		_w583_
	);
	LUT2 #(
		.INIT('he)
	) name447 (
		_w528_,
		_w583_,
		_w584_
	);
	LUT3 #(
		.INIT('ha8)
	) name448 (
		_w137_,
		_w160_,
		_w161_,
		_w585_
	);
	LUT3 #(
		.INIT('he0)
	) name449 (
		_w138_,
		_w139_,
		_w141_,
		_w586_
	);
	LUT3 #(
		.INIT('ha8)
	) name450 (
		_w145_,
		_w150_,
		_w151_,
		_w587_
	);
	LUT3 #(
		.INIT('he0)
	) name451 (
		_w142_,
		_w143_,
		_w149_,
		_w588_
	);
	LUT4 #(
		.INIT('h0001)
	) name452 (
		_w585_,
		_w586_,
		_w587_,
		_w588_,
		_w589_
	);
	LUT3 #(
		.INIT('ha8)
	) name453 (
		_w137_,
		_w187_,
		_w188_,
		_w590_
	);
	LUT3 #(
		.INIT('ha8)
	) name454 (
		_w141_,
		_w154_,
		_w155_,
		_w591_
	);
	LUT3 #(
		.INIT('ha8)
	) name455 (
		_w145_,
		_w163_,
		_w164_,
		_w592_
	);
	LUT3 #(
		.INIT('ha8)
	) name456 (
		_w149_,
		_w157_,
		_w158_,
		_w593_
	);
	LUT4 #(
		.INIT('h0001)
	) name457 (
		_w590_,
		_w591_,
		_w592_,
		_w593_,
		_w594_
	);
	LUT4 #(
		.INIT('hf7b3)
	) name458 (
		\shift[4] ,
		\shift[5] ,
		_w589_,
		_w594_,
		_w595_
	);
	LUT3 #(
		.INIT('ha8)
	) name459 (
		_w137_,
		_w202_,
		_w203_,
		_w596_
	);
	LUT3 #(
		.INIT('ha8)
	) name460 (
		_w141_,
		_w168_,
		_w169_,
		_w597_
	);
	LUT3 #(
		.INIT('ha8)
	) name461 (
		_w145_,
		_w177_,
		_w178_,
		_w598_
	);
	LUT3 #(
		.INIT('ha8)
	) name462 (
		_w149_,
		_w171_,
		_w172_,
		_w599_
	);
	LUT4 #(
		.INIT('h0001)
	) name463 (
		_w596_,
		_w597_,
		_w598_,
		_w599_,
		_w600_
	);
	LUT3 #(
		.INIT('ha8)
	) name464 (
		_w137_,
		_w174_,
		_w175_,
		_w601_
	);
	LUT3 #(
		.INIT('ha8)
	) name465 (
		_w141_,
		_w181_,
		_w182_,
		_w602_
	);
	LUT3 #(
		.INIT('ha8)
	) name466 (
		_w145_,
		_w190_,
		_w191_,
		_w603_
	);
	LUT3 #(
		.INIT('ha8)
	) name467 (
		_w149_,
		_w184_,
		_w185_,
		_w604_
	);
	LUT4 #(
		.INIT('h0001)
	) name468 (
		_w601_,
		_w602_,
		_w603_,
		_w604_,
		_w605_
	);
	LUT4 #(
		.INIT('hfedc)
	) name469 (
		\shift[4] ,
		\shift[5] ,
		_w600_,
		_w605_,
		_w606_
	);
	LUT3 #(
		.INIT('h15)
	) name470 (
		\shift[6] ,
		_w595_,
		_w606_,
		_w607_
	);
	LUT3 #(
		.INIT('ha8)
	) name471 (
		_w137_,
		_w229_,
		_w230_,
		_w608_
	);
	LUT3 #(
		.INIT('ha8)
	) name472 (
		_w141_,
		_w236_,
		_w237_,
		_w609_
	);
	LUT3 #(
		.INIT('h8a)
	) name473 (
		_w145_,
		_w245_,
		_w246_,
		_w610_
	);
	LUT3 #(
		.INIT('ha8)
	) name474 (
		_w149_,
		_w239_,
		_w240_,
		_w611_
	);
	LUT4 #(
		.INIT('h0001)
	) name475 (
		_w608_,
		_w609_,
		_w610_,
		_w611_,
		_w612_
	);
	LUT3 #(
		.INIT('ha8)
	) name476 (
		_w137_,
		_w146_,
		_w147_,
		_w613_
	);
	LUT3 #(
		.INIT('ha8)
	) name477 (
		_w141_,
		_w223_,
		_w224_,
		_w614_
	);
	LUT3 #(
		.INIT('ha8)
	) name478 (
		_w145_,
		_w232_,
		_w233_,
		_w615_
	);
	LUT3 #(
		.INIT('ha8)
	) name479 (
		_w149_,
		_w226_,
		_w227_,
		_w616_
	);
	LUT4 #(
		.INIT('h0001)
	) name480 (
		_w613_,
		_w614_,
		_w615_,
		_w616_,
		_w617_
	);
	LUT4 #(
		.INIT('hfdec)
	) name481 (
		\shift[4] ,
		\shift[5] ,
		_w612_,
		_w617_,
		_w618_
	);
	LUT3 #(
		.INIT('ha8)
	) name482 (
		_w137_,
		_w242_,
		_w243_,
		_w619_
	);
	LUT3 #(
		.INIT('ha8)
	) name483 (
		_w141_,
		_w209_,
		_w210_,
		_w620_
	);
	LUT3 #(
		.INIT('ha8)
	) name484 (
		_w145_,
		_w218_,
		_w219_,
		_w621_
	);
	LUT3 #(
		.INIT('ha8)
	) name485 (
		_w149_,
		_w212_,
		_w213_,
		_w622_
	);
	LUT4 #(
		.INIT('h0001)
	) name486 (
		_w619_,
		_w620_,
		_w621_,
		_w622_,
		_w623_
	);
	LUT3 #(
		.INIT('ha8)
	) name487 (
		_w137_,
		_w215_,
		_w216_,
		_w624_
	);
	LUT3 #(
		.INIT('ha8)
	) name488 (
		_w141_,
		_w196_,
		_w197_,
		_w625_
	);
	LUT3 #(
		.INIT('ha8)
	) name489 (
		_w145_,
		_w205_,
		_w206_,
		_w626_
	);
	LUT3 #(
		.INIT('ha8)
	) name490 (
		_w149_,
		_w199_,
		_w200_,
		_w627_
	);
	LUT4 #(
		.INIT('h0001)
	) name491 (
		_w624_,
		_w625_,
		_w626_,
		_w627_,
		_w628_
	);
	LUT4 #(
		.INIT('hfb73)
	) name492 (
		\shift[4] ,
		\shift[5] ,
		_w623_,
		_w628_,
		_w629_
	);
	LUT3 #(
		.INIT('h2a)
	) name493 (
		\shift[6] ,
		_w618_,
		_w629_,
		_w630_
	);
	LUT2 #(
		.INIT('he)
	) name494 (
		_w607_,
		_w630_,
		_w631_
	);
	LUT3 #(
		.INIT('h8a)
	) name495 (
		_w137_,
		_w271_,
		_w272_,
		_w632_
	);
	LUT3 #(
		.INIT('h8a)
	) name496 (
		_w141_,
		_w252_,
		_w253_,
		_w633_
	);
	LUT3 #(
		.INIT('h8a)
	) name497 (
		_w145_,
		_w261_,
		_w262_,
		_w634_
	);
	LUT3 #(
		.INIT('h8a)
	) name498 (
		_w149_,
		_w255_,
		_w256_,
		_w635_
	);
	LUT4 #(
		.INIT('h0001)
	) name499 (
		_w632_,
		_w633_,
		_w634_,
		_w635_,
		_w636_
	);
	LUT3 #(
		.INIT('h8a)
	) name500 (
		_w137_,
		_w298_,
		_w299_,
		_w637_
	);
	LUT3 #(
		.INIT('h8a)
	) name501 (
		_w141_,
		_w265_,
		_w266_,
		_w638_
	);
	LUT3 #(
		.INIT('h8a)
	) name502 (
		_w145_,
		_w274_,
		_w275_,
		_w639_
	);
	LUT3 #(
		.INIT('h8a)
	) name503 (
		_w149_,
		_w268_,
		_w269_,
		_w640_
	);
	LUT4 #(
		.INIT('h0001)
	) name504 (
		_w637_,
		_w638_,
		_w639_,
		_w640_,
		_w641_
	);
	LUT4 #(
		.INIT('hf7b3)
	) name505 (
		\shift[4] ,
		\shift[5] ,
		_w636_,
		_w641_,
		_w642_
	);
	LUT3 #(
		.INIT('h8a)
	) name506 (
		_w137_,
		_w326_,
		_w327_,
		_w643_
	);
	LUT3 #(
		.INIT('h8a)
	) name507 (
		_w141_,
		_w279_,
		_w280_,
		_w644_
	);
	LUT3 #(
		.INIT('h8a)
	) name508 (
		_w145_,
		_w288_,
		_w289_,
		_w645_
	);
	LUT3 #(
		.INIT('h8a)
	) name509 (
		_w149_,
		_w282_,
		_w283_,
		_w646_
	);
	LUT4 #(
		.INIT('h0001)
	) name510 (
		_w643_,
		_w644_,
		_w645_,
		_w646_,
		_w647_
	);
	LUT3 #(
		.INIT('h8a)
	) name511 (
		_w137_,
		_w285_,
		_w286_,
		_w648_
	);
	LUT3 #(
		.INIT('h8a)
	) name512 (
		_w141_,
		_w292_,
		_w293_,
		_w649_
	);
	LUT3 #(
		.INIT('h8a)
	) name513 (
		_w145_,
		_w301_,
		_w302_,
		_w650_
	);
	LUT3 #(
		.INIT('h8a)
	) name514 (
		_w149_,
		_w295_,
		_w296_,
		_w651_
	);
	LUT4 #(
		.INIT('h0001)
	) name515 (
		_w648_,
		_w649_,
		_w650_,
		_w651_,
		_w652_
	);
	LUT4 #(
		.INIT('hfedc)
	) name516 (
		\shift[4] ,
		\shift[5] ,
		_w647_,
		_w652_,
		_w653_
	);
	LUT3 #(
		.INIT('h15)
	) name517 (
		\shift[6] ,
		_w642_,
		_w653_,
		_w654_
	);
	LUT3 #(
		.INIT('h8a)
	) name518 (
		_w137_,
		_w313_,
		_w314_,
		_w655_
	);
	LUT3 #(
		.INIT('h8a)
	) name519 (
		_w141_,
		_w334_,
		_w335_,
		_w656_
	);
	LUT3 #(
		.INIT('ha8)
	) name520 (
		_w145_,
		_w343_,
		_w344_,
		_w657_
	);
	LUT3 #(
		.INIT('ha8)
	) name521 (
		_w149_,
		_w337_,
		_w338_,
		_w658_
	);
	LUT4 #(
		.INIT('h0001)
	) name522 (
		_w655_,
		_w656_,
		_w657_,
		_w658_,
		_w659_
	);
	LUT3 #(
		.INIT('h8a)
	) name523 (
		_w137_,
		_w258_,
		_w259_,
		_w660_
	);
	LUT3 #(
		.INIT('h8a)
	) name524 (
		_w141_,
		_w307_,
		_w308_,
		_w661_
	);
	LUT3 #(
		.INIT('h8a)
	) name525 (
		_w145_,
		_w316_,
		_w317_,
		_w662_
	);
	LUT3 #(
		.INIT('h8a)
	) name526 (
		_w149_,
		_w310_,
		_w311_,
		_w663_
	);
	LUT4 #(
		.INIT('h0001)
	) name527 (
		_w660_,
		_w661_,
		_w662_,
		_w663_,
		_w664_
	);
	LUT4 #(
		.INIT('hfdec)
	) name528 (
		\shift[4] ,
		\shift[5] ,
		_w659_,
		_w664_,
		_w665_
	);
	LUT3 #(
		.INIT('h8a)
	) name529 (
		_w137_,
		_w340_,
		_w341_,
		_w666_
	);
	LUT3 #(
		.INIT('h8a)
	) name530 (
		_w141_,
		_w347_,
		_w348_,
		_w667_
	);
	LUT3 #(
		.INIT('h8a)
	) name531 (
		_w145_,
		_w356_,
		_w357_,
		_w668_
	);
	LUT3 #(
		.INIT('h8a)
	) name532 (
		_w149_,
		_w350_,
		_w351_,
		_w669_
	);
	LUT4 #(
		.INIT('h0001)
	) name533 (
		_w666_,
		_w667_,
		_w668_,
		_w669_,
		_w670_
	);
	LUT3 #(
		.INIT('h8a)
	) name534 (
		_w137_,
		_w353_,
		_w354_,
		_w671_
	);
	LUT3 #(
		.INIT('h8a)
	) name535 (
		_w141_,
		_w320_,
		_w321_,
		_w672_
	);
	LUT3 #(
		.INIT('h8a)
	) name536 (
		_w145_,
		_w329_,
		_w330_,
		_w673_
	);
	LUT3 #(
		.INIT('h8a)
	) name537 (
		_w149_,
		_w323_,
		_w324_,
		_w674_
	);
	LUT4 #(
		.INIT('h0001)
	) name538 (
		_w671_,
		_w672_,
		_w673_,
		_w674_,
		_w675_
	);
	LUT4 #(
		.INIT('hfb73)
	) name539 (
		\shift[4] ,
		\shift[5] ,
		_w670_,
		_w675_,
		_w676_
	);
	LUT3 #(
		.INIT('h2a)
	) name540 (
		\shift[6] ,
		_w665_,
		_w676_,
		_w677_
	);
	LUT2 #(
		.INIT('he)
	) name541 (
		_w654_,
		_w677_,
		_w678_
	);
	LUT3 #(
		.INIT('ha8)
	) name542 (
		_w137_,
		_w382_,
		_w383_,
		_w679_
	);
	LUT3 #(
		.INIT('ha8)
	) name543 (
		_w141_,
		_w363_,
		_w364_,
		_w680_
	);
	LUT3 #(
		.INIT('ha8)
	) name544 (
		_w145_,
		_w372_,
		_w373_,
		_w681_
	);
	LUT3 #(
		.INIT('ha8)
	) name545 (
		_w149_,
		_w366_,
		_w367_,
		_w682_
	);
	LUT4 #(
		.INIT('h0001)
	) name546 (
		_w679_,
		_w680_,
		_w681_,
		_w682_,
		_w683_
	);
	LUT3 #(
		.INIT('ha8)
	) name547 (
		_w137_,
		_w409_,
		_w410_,
		_w684_
	);
	LUT3 #(
		.INIT('ha8)
	) name548 (
		_w141_,
		_w376_,
		_w377_,
		_w685_
	);
	LUT3 #(
		.INIT('ha8)
	) name549 (
		_w145_,
		_w385_,
		_w386_,
		_w686_
	);
	LUT3 #(
		.INIT('ha8)
	) name550 (
		_w149_,
		_w379_,
		_w380_,
		_w687_
	);
	LUT4 #(
		.INIT('h0001)
	) name551 (
		_w684_,
		_w685_,
		_w686_,
		_w687_,
		_w688_
	);
	LUT4 #(
		.INIT('hf7b3)
	) name552 (
		\shift[4] ,
		\shift[5] ,
		_w683_,
		_w688_,
		_w689_
	);
	LUT3 #(
		.INIT('ha8)
	) name553 (
		_w137_,
		_w437_,
		_w438_,
		_w690_
	);
	LUT3 #(
		.INIT('ha8)
	) name554 (
		_w141_,
		_w390_,
		_w391_,
		_w691_
	);
	LUT3 #(
		.INIT('ha8)
	) name555 (
		_w145_,
		_w399_,
		_w400_,
		_w692_
	);
	LUT3 #(
		.INIT('ha8)
	) name556 (
		_w149_,
		_w393_,
		_w394_,
		_w693_
	);
	LUT4 #(
		.INIT('h0001)
	) name557 (
		_w690_,
		_w691_,
		_w692_,
		_w693_,
		_w694_
	);
	LUT3 #(
		.INIT('ha8)
	) name558 (
		_w137_,
		_w396_,
		_w397_,
		_w695_
	);
	LUT3 #(
		.INIT('ha8)
	) name559 (
		_w141_,
		_w403_,
		_w404_,
		_w696_
	);
	LUT3 #(
		.INIT('ha8)
	) name560 (
		_w145_,
		_w412_,
		_w413_,
		_w697_
	);
	LUT3 #(
		.INIT('ha8)
	) name561 (
		_w149_,
		_w406_,
		_w407_,
		_w698_
	);
	LUT4 #(
		.INIT('h0001)
	) name562 (
		_w695_,
		_w696_,
		_w697_,
		_w698_,
		_w699_
	);
	LUT4 #(
		.INIT('hfedc)
	) name563 (
		\shift[4] ,
		\shift[5] ,
		_w694_,
		_w699_,
		_w700_
	);
	LUT3 #(
		.INIT('h15)
	) name564 (
		\shift[6] ,
		_w689_,
		_w700_,
		_w701_
	);
	LUT3 #(
		.INIT('ha8)
	) name565 (
		_w137_,
		_w424_,
		_w425_,
		_w702_
	);
	LUT3 #(
		.INIT('ha8)
	) name566 (
		_w141_,
		_w445_,
		_w446_,
		_w703_
	);
	LUT3 #(
		.INIT('ha8)
	) name567 (
		_w145_,
		_w454_,
		_w455_,
		_w704_
	);
	LUT3 #(
		.INIT('ha8)
	) name568 (
		_w149_,
		_w448_,
		_w449_,
		_w705_
	);
	LUT4 #(
		.INIT('h0001)
	) name569 (
		_w702_,
		_w703_,
		_w704_,
		_w705_,
		_w706_
	);
	LUT3 #(
		.INIT('ha8)
	) name570 (
		_w137_,
		_w369_,
		_w370_,
		_w707_
	);
	LUT3 #(
		.INIT('ha8)
	) name571 (
		_w141_,
		_w418_,
		_w419_,
		_w708_
	);
	LUT3 #(
		.INIT('ha8)
	) name572 (
		_w145_,
		_w427_,
		_w428_,
		_w709_
	);
	LUT3 #(
		.INIT('ha8)
	) name573 (
		_w149_,
		_w421_,
		_w422_,
		_w710_
	);
	LUT4 #(
		.INIT('h0001)
	) name574 (
		_w707_,
		_w708_,
		_w709_,
		_w710_,
		_w711_
	);
	LUT4 #(
		.INIT('hfdec)
	) name575 (
		\shift[4] ,
		\shift[5] ,
		_w706_,
		_w711_,
		_w712_
	);
	LUT3 #(
		.INIT('ha8)
	) name576 (
		_w137_,
		_w451_,
		_w452_,
		_w713_
	);
	LUT3 #(
		.INIT('ha8)
	) name577 (
		_w141_,
		_w458_,
		_w459_,
		_w714_
	);
	LUT3 #(
		.INIT('ha8)
	) name578 (
		_w145_,
		_w467_,
		_w468_,
		_w715_
	);
	LUT3 #(
		.INIT('ha8)
	) name579 (
		_w149_,
		_w461_,
		_w462_,
		_w716_
	);
	LUT4 #(
		.INIT('h0001)
	) name580 (
		_w713_,
		_w714_,
		_w715_,
		_w716_,
		_w717_
	);
	LUT3 #(
		.INIT('ha8)
	) name581 (
		_w137_,
		_w464_,
		_w465_,
		_w718_
	);
	LUT3 #(
		.INIT('ha8)
	) name582 (
		_w141_,
		_w431_,
		_w432_,
		_w719_
	);
	LUT3 #(
		.INIT('ha8)
	) name583 (
		_w145_,
		_w440_,
		_w441_,
		_w720_
	);
	LUT3 #(
		.INIT('ha8)
	) name584 (
		_w149_,
		_w434_,
		_w435_,
		_w721_
	);
	LUT4 #(
		.INIT('h0001)
	) name585 (
		_w718_,
		_w719_,
		_w720_,
		_w721_,
		_w722_
	);
	LUT4 #(
		.INIT('hfb73)
	) name586 (
		\shift[4] ,
		\shift[5] ,
		_w717_,
		_w722_,
		_w723_
	);
	LUT3 #(
		.INIT('h2a)
	) name587 (
		\shift[6] ,
		_w712_,
		_w723_,
		_w724_
	);
	LUT2 #(
		.INIT('he)
	) name588 (
		_w701_,
		_w724_,
		_w725_
	);
	LUT3 #(
		.INIT('h8a)
	) name589 (
		_w137_,
		_w493_,
		_w494_,
		_w726_
	);
	LUT3 #(
		.INIT('h8a)
	) name590 (
		_w141_,
		_w514_,
		_w515_,
		_w727_
	);
	LUT3 #(
		.INIT('h8a)
	) name591 (
		_w145_,
		_w523_,
		_w524_,
		_w728_
	);
	LUT3 #(
		.INIT('h8a)
	) name592 (
		_w149_,
		_w517_,
		_w518_,
		_w729_
	);
	LUT4 #(
		.INIT('h0001)
	) name593 (
		_w726_,
		_w727_,
		_w728_,
		_w729_,
		_w730_
	);
	LUT3 #(
		.INIT('h8a)
	) name594 (
		_w137_,
		_w480_,
		_w481_,
		_w731_
	);
	LUT3 #(
		.INIT('h8a)
	) name595 (
		_w141_,
		_w487_,
		_w488_,
		_w732_
	);
	LUT3 #(
		.INIT('h8a)
	) name596 (
		_w145_,
		_w496_,
		_w497_,
		_w733_
	);
	LUT3 #(
		.INIT('h8a)
	) name597 (
		_w149_,
		_w490_,
		_w491_,
		_w734_
	);
	LUT4 #(
		.INIT('h0001)
	) name598 (
		_w731_,
		_w732_,
		_w733_,
		_w734_,
		_w735_
	);
	LUT4 #(
		.INIT('hf7b3)
	) name599 (
		\shift[4] ,
		\shift[5] ,
		_w730_,
		_w735_,
		_w736_
	);
	LUT3 #(
		.INIT('h8a)
	) name600 (
		_w137_,
		_w562_,
		_w563_,
		_w737_
	);
	LUT3 #(
		.INIT('h8a)
	) name601 (
		_w141_,
		_w501_,
		_w502_,
		_w738_
	);
	LUT3 #(
		.INIT('h8a)
	) name602 (
		_w145_,
		_w510_,
		_w511_,
		_w739_
	);
	LUT3 #(
		.INIT('h8a)
	) name603 (
		_w149_,
		_w504_,
		_w505_,
		_w740_
	);
	LUT4 #(
		.INIT('h0001)
	) name604 (
		_w737_,
		_w738_,
		_w739_,
		_w740_,
		_w741_
	);
	LUT3 #(
		.INIT('h8a)
	) name605 (
		_w137_,
		_w507_,
		_w508_,
		_w742_
	);
	LUT3 #(
		.INIT('h8a)
	) name606 (
		_w141_,
		_w474_,
		_w475_,
		_w743_
	);
	LUT3 #(
		.INIT('h8a)
	) name607 (
		_w145_,
		_w483_,
		_w484_,
		_w744_
	);
	LUT3 #(
		.INIT('h8a)
	) name608 (
		_w149_,
		_w477_,
		_w478_,
		_w745_
	);
	LUT4 #(
		.INIT('h0001)
	) name609 (
		_w742_,
		_w743_,
		_w744_,
		_w745_,
		_w746_
	);
	LUT4 #(
		.INIT('hfedc)
	) name610 (
		\shift[4] ,
		\shift[5] ,
		_w741_,
		_w746_,
		_w747_
	);
	LUT3 #(
		.INIT('h15)
	) name611 (
		\shift[6] ,
		_w736_,
		_w747_,
		_w748_
	);
	LUT3 #(
		.INIT('h8a)
	) name612 (
		_w141_,
		_w542_,
		_w543_,
		_w749_
	);
	LUT3 #(
		.INIT('ha8)
	) name613 (
		_w149_,
		_w545_,
		_w546_,
		_w750_
	);
	LUT3 #(
		.INIT('h8a)
	) name614 (
		_w145_,
		_w551_,
		_w552_,
		_w751_
	);
	LUT3 #(
		.INIT('h8a)
	) name615 (
		_w137_,
		_w535_,
		_w536_,
		_w752_
	);
	LUT4 #(
		.INIT('h0001)
	) name616 (
		_w749_,
		_w750_,
		_w751_,
		_w752_,
		_w753_
	);
	LUT3 #(
		.INIT('h8a)
	) name617 (
		_w137_,
		_w520_,
		_w521_,
		_w754_
	);
	LUT3 #(
		.INIT('h8a)
	) name618 (
		_w141_,
		_w529_,
		_w530_,
		_w755_
	);
	LUT3 #(
		.INIT('h8a)
	) name619 (
		_w145_,
		_w538_,
		_w539_,
		_w756_
	);
	LUT3 #(
		.INIT('h8a)
	) name620 (
		_w149_,
		_w532_,
		_w533_,
		_w757_
	);
	LUT4 #(
		.INIT('h0001)
	) name621 (
		_w754_,
		_w755_,
		_w756_,
		_w757_,
		_w758_
	);
	LUT4 #(
		.INIT('hfdec)
	) name622 (
		\shift[4] ,
		\shift[5] ,
		_w753_,
		_w758_,
		_w759_
	);
	LUT3 #(
		.INIT('h8a)
	) name623 (
		_w137_,
		_w548_,
		_w549_,
		_w760_
	);
	LUT3 #(
		.INIT('h8a)
	) name624 (
		_w141_,
		_w569_,
		_w570_,
		_w761_
	);
	LUT3 #(
		.INIT('h8a)
	) name625 (
		_w145_,
		_w578_,
		_w579_,
		_w762_
	);
	LUT3 #(
		.INIT('h8a)
	) name626 (
		_w149_,
		_w572_,
		_w573_,
		_w763_
	);
	LUT4 #(
		.INIT('h0001)
	) name627 (
		_w760_,
		_w761_,
		_w762_,
		_w763_,
		_w764_
	);
	LUT3 #(
		.INIT('h8a)
	) name628 (
		_w137_,
		_w575_,
		_w576_,
		_w765_
	);
	LUT3 #(
		.INIT('h8a)
	) name629 (
		_w141_,
		_w556_,
		_w557_,
		_w766_
	);
	LUT3 #(
		.INIT('h8a)
	) name630 (
		_w145_,
		_w565_,
		_w566_,
		_w767_
	);
	LUT3 #(
		.INIT('h8a)
	) name631 (
		_w149_,
		_w559_,
		_w560_,
		_w768_
	);
	LUT4 #(
		.INIT('h0001)
	) name632 (
		_w765_,
		_w766_,
		_w767_,
		_w768_,
		_w769_
	);
	LUT4 #(
		.INIT('hfb73)
	) name633 (
		\shift[4] ,
		\shift[5] ,
		_w764_,
		_w769_,
		_w770_
	);
	LUT3 #(
		.INIT('h2a)
	) name634 (
		\shift[6] ,
		_w759_,
		_w770_,
		_w771_
	);
	LUT2 #(
		.INIT('he)
	) name635 (
		_w748_,
		_w771_,
		_w772_
	);
	LUT3 #(
		.INIT('ha8)
	) name636 (
		_w137_,
		_w163_,
		_w164_,
		_w773_
	);
	LUT3 #(
		.INIT('ha8)
	) name637 (
		_w141_,
		_w160_,
		_w161_,
		_w774_
	);
	LUT3 #(
		.INIT('he0)
	) name638 (
		_w142_,
		_w143_,
		_w145_,
		_w775_
	);
	LUT3 #(
		.INIT('he0)
	) name639 (
		_w138_,
		_w139_,
		_w149_,
		_w776_
	);
	LUT4 #(
		.INIT('h0001)
	) name640 (
		_w773_,
		_w774_,
		_w775_,
		_w776_,
		_w777_
	);
	LUT3 #(
		.INIT('ha8)
	) name641 (
		_w137_,
		_w190_,
		_w191_,
		_w778_
	);
	LUT3 #(
		.INIT('ha8)
	) name642 (
		_w141_,
		_w187_,
		_w188_,
		_w779_
	);
	LUT3 #(
		.INIT('ha8)
	) name643 (
		_w145_,
		_w157_,
		_w158_,
		_w780_
	);
	LUT3 #(
		.INIT('ha8)
	) name644 (
		_w149_,
		_w154_,
		_w155_,
		_w781_
	);
	LUT4 #(
		.INIT('h0001)
	) name645 (
		_w778_,
		_w779_,
		_w780_,
		_w781_,
		_w782_
	);
	LUT4 #(
		.INIT('hf7b3)
	) name646 (
		\shift[4] ,
		\shift[5] ,
		_w777_,
		_w782_,
		_w783_
	);
	LUT3 #(
		.INIT('ha8)
	) name647 (
		_w137_,
		_w205_,
		_w206_,
		_w784_
	);
	LUT3 #(
		.INIT('ha8)
	) name648 (
		_w141_,
		_w202_,
		_w203_,
		_w785_
	);
	LUT3 #(
		.INIT('ha8)
	) name649 (
		_w145_,
		_w171_,
		_w172_,
		_w786_
	);
	LUT3 #(
		.INIT('ha8)
	) name650 (
		_w149_,
		_w168_,
		_w169_,
		_w787_
	);
	LUT4 #(
		.INIT('h0001)
	) name651 (
		_w784_,
		_w785_,
		_w786_,
		_w787_,
		_w788_
	);
	LUT3 #(
		.INIT('ha8)
	) name652 (
		_w137_,
		_w177_,
		_w178_,
		_w789_
	);
	LUT3 #(
		.INIT('ha8)
	) name653 (
		_w141_,
		_w174_,
		_w175_,
		_w790_
	);
	LUT3 #(
		.INIT('ha8)
	) name654 (
		_w145_,
		_w184_,
		_w185_,
		_w791_
	);
	LUT3 #(
		.INIT('ha8)
	) name655 (
		_w149_,
		_w181_,
		_w182_,
		_w792_
	);
	LUT4 #(
		.INIT('h0001)
	) name656 (
		_w789_,
		_w790_,
		_w791_,
		_w792_,
		_w793_
	);
	LUT4 #(
		.INIT('hfedc)
	) name657 (
		\shift[4] ,
		\shift[5] ,
		_w788_,
		_w793_,
		_w794_
	);
	LUT3 #(
		.INIT('h15)
	) name658 (
		\shift[6] ,
		_w783_,
		_w794_,
		_w795_
	);
	LUT3 #(
		.INIT('ha8)
	) name659 (
		_w137_,
		_w232_,
		_w233_,
		_w796_
	);
	LUT3 #(
		.INIT('ha8)
	) name660 (
		_w141_,
		_w229_,
		_w230_,
		_w797_
	);
	LUT3 #(
		.INIT('ha8)
	) name661 (
		_w145_,
		_w239_,
		_w240_,
		_w798_
	);
	LUT3 #(
		.INIT('ha8)
	) name662 (
		_w149_,
		_w236_,
		_w237_,
		_w799_
	);
	LUT4 #(
		.INIT('h0001)
	) name663 (
		_w796_,
		_w797_,
		_w798_,
		_w799_,
		_w800_
	);
	LUT3 #(
		.INIT('ha8)
	) name664 (
		_w137_,
		_w150_,
		_w151_,
		_w801_
	);
	LUT3 #(
		.INIT('ha8)
	) name665 (
		_w141_,
		_w146_,
		_w147_,
		_w802_
	);
	LUT3 #(
		.INIT('ha8)
	) name666 (
		_w145_,
		_w226_,
		_w227_,
		_w803_
	);
	LUT3 #(
		.INIT('ha8)
	) name667 (
		_w149_,
		_w223_,
		_w224_,
		_w804_
	);
	LUT4 #(
		.INIT('h0001)
	) name668 (
		_w801_,
		_w802_,
		_w803_,
		_w804_,
		_w805_
	);
	LUT4 #(
		.INIT('hfdec)
	) name669 (
		\shift[4] ,
		\shift[5] ,
		_w800_,
		_w805_,
		_w806_
	);
	LUT3 #(
		.INIT('h8a)
	) name670 (
		_w137_,
		_w245_,
		_w246_,
		_w807_
	);
	LUT3 #(
		.INIT('ha8)
	) name671 (
		_w141_,
		_w242_,
		_w243_,
		_w808_
	);
	LUT3 #(
		.INIT('ha8)
	) name672 (
		_w145_,
		_w212_,
		_w213_,
		_w809_
	);
	LUT3 #(
		.INIT('ha8)
	) name673 (
		_w149_,
		_w209_,
		_w210_,
		_w810_
	);
	LUT4 #(
		.INIT('h0001)
	) name674 (
		_w807_,
		_w808_,
		_w809_,
		_w810_,
		_w811_
	);
	LUT3 #(
		.INIT('ha8)
	) name675 (
		_w137_,
		_w218_,
		_w219_,
		_w812_
	);
	LUT3 #(
		.INIT('ha8)
	) name676 (
		_w141_,
		_w215_,
		_w216_,
		_w813_
	);
	LUT3 #(
		.INIT('ha8)
	) name677 (
		_w145_,
		_w199_,
		_w200_,
		_w814_
	);
	LUT3 #(
		.INIT('ha8)
	) name678 (
		_w149_,
		_w196_,
		_w197_,
		_w815_
	);
	LUT4 #(
		.INIT('h0001)
	) name679 (
		_w812_,
		_w813_,
		_w814_,
		_w815_,
		_w816_
	);
	LUT4 #(
		.INIT('hfb73)
	) name680 (
		\shift[4] ,
		\shift[5] ,
		_w811_,
		_w816_,
		_w817_
	);
	LUT3 #(
		.INIT('h2a)
	) name681 (
		\shift[6] ,
		_w806_,
		_w817_,
		_w818_
	);
	LUT2 #(
		.INIT('he)
	) name682 (
		_w795_,
		_w818_,
		_w819_
	);
	LUT3 #(
		.INIT('h8a)
	) name683 (
		_w137_,
		_w274_,
		_w275_,
		_w820_
	);
	LUT3 #(
		.INIT('h8a)
	) name684 (
		_w141_,
		_w271_,
		_w272_,
		_w821_
	);
	LUT3 #(
		.INIT('h8a)
	) name685 (
		_w145_,
		_w255_,
		_w256_,
		_w822_
	);
	LUT3 #(
		.INIT('h8a)
	) name686 (
		_w149_,
		_w252_,
		_w253_,
		_w823_
	);
	LUT4 #(
		.INIT('h0001)
	) name687 (
		_w820_,
		_w821_,
		_w822_,
		_w823_,
		_w824_
	);
	LUT3 #(
		.INIT('h8a)
	) name688 (
		_w137_,
		_w301_,
		_w302_,
		_w825_
	);
	LUT3 #(
		.INIT('h8a)
	) name689 (
		_w141_,
		_w298_,
		_w299_,
		_w826_
	);
	LUT3 #(
		.INIT('h8a)
	) name690 (
		_w145_,
		_w268_,
		_w269_,
		_w827_
	);
	LUT3 #(
		.INIT('h8a)
	) name691 (
		_w149_,
		_w265_,
		_w266_,
		_w828_
	);
	LUT4 #(
		.INIT('h0001)
	) name692 (
		_w825_,
		_w826_,
		_w827_,
		_w828_,
		_w829_
	);
	LUT4 #(
		.INIT('hf7b3)
	) name693 (
		\shift[4] ,
		\shift[5] ,
		_w824_,
		_w829_,
		_w830_
	);
	LUT3 #(
		.INIT('h8a)
	) name694 (
		_w137_,
		_w329_,
		_w330_,
		_w831_
	);
	LUT3 #(
		.INIT('h8a)
	) name695 (
		_w141_,
		_w326_,
		_w327_,
		_w832_
	);
	LUT3 #(
		.INIT('h8a)
	) name696 (
		_w145_,
		_w282_,
		_w283_,
		_w833_
	);
	LUT3 #(
		.INIT('h8a)
	) name697 (
		_w149_,
		_w279_,
		_w280_,
		_w834_
	);
	LUT4 #(
		.INIT('h0001)
	) name698 (
		_w831_,
		_w832_,
		_w833_,
		_w834_,
		_w835_
	);
	LUT3 #(
		.INIT('h8a)
	) name699 (
		_w137_,
		_w288_,
		_w289_,
		_w836_
	);
	LUT3 #(
		.INIT('h8a)
	) name700 (
		_w141_,
		_w285_,
		_w286_,
		_w837_
	);
	LUT3 #(
		.INIT('h8a)
	) name701 (
		_w145_,
		_w295_,
		_w296_,
		_w838_
	);
	LUT3 #(
		.INIT('h8a)
	) name702 (
		_w149_,
		_w292_,
		_w293_,
		_w839_
	);
	LUT4 #(
		.INIT('h0001)
	) name703 (
		_w836_,
		_w837_,
		_w838_,
		_w839_,
		_w840_
	);
	LUT4 #(
		.INIT('hfedc)
	) name704 (
		\shift[4] ,
		\shift[5] ,
		_w835_,
		_w840_,
		_w841_
	);
	LUT3 #(
		.INIT('h15)
	) name705 (
		\shift[6] ,
		_w830_,
		_w841_,
		_w842_
	);
	LUT3 #(
		.INIT('h8a)
	) name706 (
		_w137_,
		_w316_,
		_w317_,
		_w843_
	);
	LUT3 #(
		.INIT('h8a)
	) name707 (
		_w141_,
		_w313_,
		_w314_,
		_w844_
	);
	LUT3 #(
		.INIT('ha8)
	) name708 (
		_w145_,
		_w337_,
		_w338_,
		_w845_
	);
	LUT3 #(
		.INIT('h8a)
	) name709 (
		_w149_,
		_w334_,
		_w335_,
		_w846_
	);
	LUT4 #(
		.INIT('h0001)
	) name710 (
		_w843_,
		_w844_,
		_w845_,
		_w846_,
		_w847_
	);
	LUT3 #(
		.INIT('h8a)
	) name711 (
		_w137_,
		_w261_,
		_w262_,
		_w848_
	);
	LUT3 #(
		.INIT('h8a)
	) name712 (
		_w141_,
		_w258_,
		_w259_,
		_w849_
	);
	LUT3 #(
		.INIT('h8a)
	) name713 (
		_w145_,
		_w310_,
		_w311_,
		_w850_
	);
	LUT3 #(
		.INIT('h8a)
	) name714 (
		_w149_,
		_w307_,
		_w308_,
		_w851_
	);
	LUT4 #(
		.INIT('h0001)
	) name715 (
		_w848_,
		_w849_,
		_w850_,
		_w851_,
		_w852_
	);
	LUT4 #(
		.INIT('hfdec)
	) name716 (
		\shift[4] ,
		\shift[5] ,
		_w847_,
		_w852_,
		_w853_
	);
	LUT3 #(
		.INIT('ha8)
	) name717 (
		_w137_,
		_w343_,
		_w344_,
		_w854_
	);
	LUT3 #(
		.INIT('h8a)
	) name718 (
		_w141_,
		_w340_,
		_w341_,
		_w855_
	);
	LUT3 #(
		.INIT('h8a)
	) name719 (
		_w145_,
		_w350_,
		_w351_,
		_w856_
	);
	LUT3 #(
		.INIT('h8a)
	) name720 (
		_w149_,
		_w347_,
		_w348_,
		_w857_
	);
	LUT4 #(
		.INIT('h0001)
	) name721 (
		_w854_,
		_w855_,
		_w856_,
		_w857_,
		_w858_
	);
	LUT3 #(
		.INIT('h8a)
	) name722 (
		_w137_,
		_w356_,
		_w357_,
		_w859_
	);
	LUT3 #(
		.INIT('h8a)
	) name723 (
		_w141_,
		_w353_,
		_w354_,
		_w860_
	);
	LUT3 #(
		.INIT('h8a)
	) name724 (
		_w145_,
		_w323_,
		_w324_,
		_w861_
	);
	LUT3 #(
		.INIT('h8a)
	) name725 (
		_w149_,
		_w320_,
		_w321_,
		_w862_
	);
	LUT4 #(
		.INIT('h0001)
	) name726 (
		_w859_,
		_w860_,
		_w861_,
		_w862_,
		_w863_
	);
	LUT4 #(
		.INIT('hfb73)
	) name727 (
		\shift[4] ,
		\shift[5] ,
		_w858_,
		_w863_,
		_w864_
	);
	LUT3 #(
		.INIT('h2a)
	) name728 (
		\shift[6] ,
		_w853_,
		_w864_,
		_w865_
	);
	LUT2 #(
		.INIT('he)
	) name729 (
		_w842_,
		_w865_,
		_w866_
	);
	LUT3 #(
		.INIT('ha8)
	) name730 (
		_w137_,
		_w385_,
		_w386_,
		_w867_
	);
	LUT3 #(
		.INIT('ha8)
	) name731 (
		_w141_,
		_w382_,
		_w383_,
		_w868_
	);
	LUT3 #(
		.INIT('ha8)
	) name732 (
		_w145_,
		_w366_,
		_w367_,
		_w869_
	);
	LUT3 #(
		.INIT('ha8)
	) name733 (
		_w149_,
		_w363_,
		_w364_,
		_w870_
	);
	LUT4 #(
		.INIT('h0001)
	) name734 (
		_w867_,
		_w868_,
		_w869_,
		_w870_,
		_w871_
	);
	LUT3 #(
		.INIT('ha8)
	) name735 (
		_w137_,
		_w412_,
		_w413_,
		_w872_
	);
	LUT3 #(
		.INIT('ha8)
	) name736 (
		_w141_,
		_w409_,
		_w410_,
		_w873_
	);
	LUT3 #(
		.INIT('ha8)
	) name737 (
		_w145_,
		_w379_,
		_w380_,
		_w874_
	);
	LUT3 #(
		.INIT('ha8)
	) name738 (
		_w149_,
		_w376_,
		_w377_,
		_w875_
	);
	LUT4 #(
		.INIT('h0001)
	) name739 (
		_w872_,
		_w873_,
		_w874_,
		_w875_,
		_w876_
	);
	LUT4 #(
		.INIT('hf7b3)
	) name740 (
		\shift[4] ,
		\shift[5] ,
		_w871_,
		_w876_,
		_w877_
	);
	LUT3 #(
		.INIT('ha8)
	) name741 (
		_w137_,
		_w440_,
		_w441_,
		_w878_
	);
	LUT3 #(
		.INIT('ha8)
	) name742 (
		_w141_,
		_w437_,
		_w438_,
		_w879_
	);
	LUT3 #(
		.INIT('ha8)
	) name743 (
		_w145_,
		_w393_,
		_w394_,
		_w880_
	);
	LUT3 #(
		.INIT('ha8)
	) name744 (
		_w149_,
		_w390_,
		_w391_,
		_w881_
	);
	LUT4 #(
		.INIT('h0001)
	) name745 (
		_w878_,
		_w879_,
		_w880_,
		_w881_,
		_w882_
	);
	LUT3 #(
		.INIT('ha8)
	) name746 (
		_w137_,
		_w399_,
		_w400_,
		_w883_
	);
	LUT3 #(
		.INIT('ha8)
	) name747 (
		_w141_,
		_w396_,
		_w397_,
		_w884_
	);
	LUT3 #(
		.INIT('ha8)
	) name748 (
		_w145_,
		_w406_,
		_w407_,
		_w885_
	);
	LUT3 #(
		.INIT('ha8)
	) name749 (
		_w149_,
		_w403_,
		_w404_,
		_w886_
	);
	LUT4 #(
		.INIT('h0001)
	) name750 (
		_w883_,
		_w884_,
		_w885_,
		_w886_,
		_w887_
	);
	LUT4 #(
		.INIT('hfedc)
	) name751 (
		\shift[4] ,
		\shift[5] ,
		_w882_,
		_w887_,
		_w888_
	);
	LUT3 #(
		.INIT('h15)
	) name752 (
		\shift[6] ,
		_w877_,
		_w888_,
		_w889_
	);
	LUT3 #(
		.INIT('ha8)
	) name753 (
		_w137_,
		_w427_,
		_w428_,
		_w890_
	);
	LUT3 #(
		.INIT('ha8)
	) name754 (
		_w141_,
		_w424_,
		_w425_,
		_w891_
	);
	LUT3 #(
		.INIT('ha8)
	) name755 (
		_w145_,
		_w448_,
		_w449_,
		_w892_
	);
	LUT3 #(
		.INIT('ha8)
	) name756 (
		_w149_,
		_w445_,
		_w446_,
		_w893_
	);
	LUT4 #(
		.INIT('h0001)
	) name757 (
		_w890_,
		_w891_,
		_w892_,
		_w893_,
		_w894_
	);
	LUT3 #(
		.INIT('ha8)
	) name758 (
		_w137_,
		_w372_,
		_w373_,
		_w895_
	);
	LUT3 #(
		.INIT('ha8)
	) name759 (
		_w141_,
		_w369_,
		_w370_,
		_w896_
	);
	LUT3 #(
		.INIT('ha8)
	) name760 (
		_w145_,
		_w421_,
		_w422_,
		_w897_
	);
	LUT3 #(
		.INIT('ha8)
	) name761 (
		_w149_,
		_w418_,
		_w419_,
		_w898_
	);
	LUT4 #(
		.INIT('h0001)
	) name762 (
		_w895_,
		_w896_,
		_w897_,
		_w898_,
		_w899_
	);
	LUT4 #(
		.INIT('hfdec)
	) name763 (
		\shift[4] ,
		\shift[5] ,
		_w894_,
		_w899_,
		_w900_
	);
	LUT3 #(
		.INIT('ha8)
	) name764 (
		_w137_,
		_w454_,
		_w455_,
		_w901_
	);
	LUT3 #(
		.INIT('ha8)
	) name765 (
		_w141_,
		_w451_,
		_w452_,
		_w902_
	);
	LUT3 #(
		.INIT('ha8)
	) name766 (
		_w145_,
		_w461_,
		_w462_,
		_w903_
	);
	LUT3 #(
		.INIT('ha8)
	) name767 (
		_w149_,
		_w458_,
		_w459_,
		_w904_
	);
	LUT4 #(
		.INIT('h0001)
	) name768 (
		_w901_,
		_w902_,
		_w903_,
		_w904_,
		_w905_
	);
	LUT3 #(
		.INIT('ha8)
	) name769 (
		_w137_,
		_w467_,
		_w468_,
		_w906_
	);
	LUT3 #(
		.INIT('ha8)
	) name770 (
		_w141_,
		_w464_,
		_w465_,
		_w907_
	);
	LUT3 #(
		.INIT('ha8)
	) name771 (
		_w145_,
		_w434_,
		_w435_,
		_w908_
	);
	LUT3 #(
		.INIT('ha8)
	) name772 (
		_w149_,
		_w431_,
		_w432_,
		_w909_
	);
	LUT4 #(
		.INIT('h0001)
	) name773 (
		_w906_,
		_w907_,
		_w908_,
		_w909_,
		_w910_
	);
	LUT4 #(
		.INIT('hfb73)
	) name774 (
		\shift[4] ,
		\shift[5] ,
		_w905_,
		_w910_,
		_w911_
	);
	LUT3 #(
		.INIT('h2a)
	) name775 (
		\shift[6] ,
		_w900_,
		_w911_,
		_w912_
	);
	LUT2 #(
		.INIT('he)
	) name776 (
		_w889_,
		_w912_,
		_w913_
	);
	LUT3 #(
		.INIT('h8a)
	) name777 (
		_w137_,
		_w496_,
		_w497_,
		_w914_
	);
	LUT3 #(
		.INIT('h8a)
	) name778 (
		_w141_,
		_w493_,
		_w494_,
		_w915_
	);
	LUT3 #(
		.INIT('h8a)
	) name779 (
		_w145_,
		_w517_,
		_w518_,
		_w916_
	);
	LUT3 #(
		.INIT('h8a)
	) name780 (
		_w149_,
		_w514_,
		_w515_,
		_w917_
	);
	LUT4 #(
		.INIT('h0001)
	) name781 (
		_w914_,
		_w915_,
		_w916_,
		_w917_,
		_w918_
	);
	LUT3 #(
		.INIT('h8a)
	) name782 (
		_w137_,
		_w483_,
		_w484_,
		_w919_
	);
	LUT3 #(
		.INIT('h8a)
	) name783 (
		_w141_,
		_w480_,
		_w481_,
		_w920_
	);
	LUT3 #(
		.INIT('h8a)
	) name784 (
		_w145_,
		_w490_,
		_w491_,
		_w921_
	);
	LUT3 #(
		.INIT('h8a)
	) name785 (
		_w149_,
		_w487_,
		_w488_,
		_w922_
	);
	LUT4 #(
		.INIT('h0001)
	) name786 (
		_w919_,
		_w920_,
		_w921_,
		_w922_,
		_w923_
	);
	LUT4 #(
		.INIT('hf7b3)
	) name787 (
		\shift[4] ,
		\shift[5] ,
		_w918_,
		_w923_,
		_w924_
	);
	LUT3 #(
		.INIT('h8a)
	) name788 (
		_w137_,
		_w565_,
		_w566_,
		_w925_
	);
	LUT3 #(
		.INIT('h8a)
	) name789 (
		_w141_,
		_w562_,
		_w563_,
		_w926_
	);
	LUT3 #(
		.INIT('h8a)
	) name790 (
		_w145_,
		_w504_,
		_w505_,
		_w927_
	);
	LUT3 #(
		.INIT('h8a)
	) name791 (
		_w149_,
		_w501_,
		_w502_,
		_w928_
	);
	LUT4 #(
		.INIT('h0001)
	) name792 (
		_w925_,
		_w926_,
		_w927_,
		_w928_,
		_w929_
	);
	LUT3 #(
		.INIT('h8a)
	) name793 (
		_w137_,
		_w510_,
		_w511_,
		_w930_
	);
	LUT3 #(
		.INIT('h8a)
	) name794 (
		_w141_,
		_w507_,
		_w508_,
		_w931_
	);
	LUT3 #(
		.INIT('h8a)
	) name795 (
		_w145_,
		_w477_,
		_w478_,
		_w932_
	);
	LUT3 #(
		.INIT('h8a)
	) name796 (
		_w149_,
		_w474_,
		_w475_,
		_w933_
	);
	LUT4 #(
		.INIT('h0001)
	) name797 (
		_w930_,
		_w931_,
		_w932_,
		_w933_,
		_w934_
	);
	LUT4 #(
		.INIT('hfedc)
	) name798 (
		\shift[4] ,
		\shift[5] ,
		_w929_,
		_w934_,
		_w935_
	);
	LUT3 #(
		.INIT('h15)
	) name799 (
		\shift[6] ,
		_w924_,
		_w935_,
		_w936_
	);
	LUT3 #(
		.INIT('h8a)
	) name800 (
		_w137_,
		_w538_,
		_w539_,
		_w937_
	);
	LUT3 #(
		.INIT('h8a)
	) name801 (
		_w149_,
		_w542_,
		_w543_,
		_w938_
	);
	LUT3 #(
		.INIT('ha8)
	) name802 (
		_w145_,
		_w545_,
		_w546_,
		_w939_
	);
	LUT3 #(
		.INIT('h8a)
	) name803 (
		_w141_,
		_w535_,
		_w536_,
		_w940_
	);
	LUT4 #(
		.INIT('h0001)
	) name804 (
		_w937_,
		_w938_,
		_w939_,
		_w940_,
		_w941_
	);
	LUT3 #(
		.INIT('h8a)
	) name805 (
		_w137_,
		_w523_,
		_w524_,
		_w942_
	);
	LUT3 #(
		.INIT('h8a)
	) name806 (
		_w141_,
		_w520_,
		_w521_,
		_w943_
	);
	LUT3 #(
		.INIT('h8a)
	) name807 (
		_w145_,
		_w532_,
		_w533_,
		_w944_
	);
	LUT3 #(
		.INIT('h8a)
	) name808 (
		_w149_,
		_w529_,
		_w530_,
		_w945_
	);
	LUT4 #(
		.INIT('h0001)
	) name809 (
		_w942_,
		_w943_,
		_w944_,
		_w945_,
		_w946_
	);
	LUT4 #(
		.INIT('hfdec)
	) name810 (
		\shift[4] ,
		\shift[5] ,
		_w941_,
		_w946_,
		_w947_
	);
	LUT3 #(
		.INIT('h8a)
	) name811 (
		_w137_,
		_w551_,
		_w552_,
		_w948_
	);
	LUT3 #(
		.INIT('h8a)
	) name812 (
		_w141_,
		_w548_,
		_w549_,
		_w949_
	);
	LUT3 #(
		.INIT('h8a)
	) name813 (
		_w145_,
		_w572_,
		_w573_,
		_w950_
	);
	LUT3 #(
		.INIT('h8a)
	) name814 (
		_w149_,
		_w569_,
		_w570_,
		_w951_
	);
	LUT4 #(
		.INIT('h0001)
	) name815 (
		_w948_,
		_w949_,
		_w950_,
		_w951_,
		_w952_
	);
	LUT3 #(
		.INIT('h8a)
	) name816 (
		_w137_,
		_w578_,
		_w579_,
		_w953_
	);
	LUT3 #(
		.INIT('h8a)
	) name817 (
		_w141_,
		_w575_,
		_w576_,
		_w954_
	);
	LUT3 #(
		.INIT('h8a)
	) name818 (
		_w145_,
		_w559_,
		_w560_,
		_w955_
	);
	LUT3 #(
		.INIT('h8a)
	) name819 (
		_w149_,
		_w556_,
		_w557_,
		_w956_
	);
	LUT4 #(
		.INIT('h0001)
	) name820 (
		_w953_,
		_w954_,
		_w955_,
		_w956_,
		_w957_
	);
	LUT4 #(
		.INIT('hfb73)
	) name821 (
		\shift[4] ,
		\shift[5] ,
		_w952_,
		_w957_,
		_w958_
	);
	LUT3 #(
		.INIT('h2a)
	) name822 (
		\shift[6] ,
		_w947_,
		_w958_,
		_w959_
	);
	LUT2 #(
		.INIT('he)
	) name823 (
		_w936_,
		_w959_,
		_w960_
	);
	LUT3 #(
		.INIT('ha8)
	) name824 (
		_w137_,
		_w157_,
		_w158_,
		_w961_
	);
	LUT3 #(
		.INIT('ha8)
	) name825 (
		_w141_,
		_w163_,
		_w164_,
		_w962_
	);
	LUT3 #(
		.INIT('he0)
	) name826 (
		_w138_,
		_w139_,
		_w145_,
		_w963_
	);
	LUT3 #(
		.INIT('ha8)
	) name827 (
		_w149_,
		_w160_,
		_w161_,
		_w964_
	);
	LUT4 #(
		.INIT('h0001)
	) name828 (
		_w961_,
		_w962_,
		_w963_,
		_w964_,
		_w965_
	);
	LUT3 #(
		.INIT('ha8)
	) name829 (
		_w137_,
		_w184_,
		_w185_,
		_w966_
	);
	LUT3 #(
		.INIT('ha8)
	) name830 (
		_w141_,
		_w190_,
		_w191_,
		_w967_
	);
	LUT3 #(
		.INIT('ha8)
	) name831 (
		_w145_,
		_w154_,
		_w155_,
		_w968_
	);
	LUT3 #(
		.INIT('ha8)
	) name832 (
		_w149_,
		_w187_,
		_w188_,
		_w969_
	);
	LUT4 #(
		.INIT('h0001)
	) name833 (
		_w966_,
		_w967_,
		_w968_,
		_w969_,
		_w970_
	);
	LUT4 #(
		.INIT('hf7b3)
	) name834 (
		\shift[4] ,
		\shift[5] ,
		_w965_,
		_w970_,
		_w971_
	);
	LUT3 #(
		.INIT('ha8)
	) name835 (
		_w137_,
		_w199_,
		_w200_,
		_w972_
	);
	LUT3 #(
		.INIT('ha8)
	) name836 (
		_w141_,
		_w205_,
		_w206_,
		_w973_
	);
	LUT3 #(
		.INIT('ha8)
	) name837 (
		_w145_,
		_w168_,
		_w169_,
		_w974_
	);
	LUT3 #(
		.INIT('ha8)
	) name838 (
		_w149_,
		_w202_,
		_w203_,
		_w975_
	);
	LUT4 #(
		.INIT('h0001)
	) name839 (
		_w972_,
		_w973_,
		_w974_,
		_w975_,
		_w976_
	);
	LUT3 #(
		.INIT('ha8)
	) name840 (
		_w137_,
		_w171_,
		_w172_,
		_w977_
	);
	LUT3 #(
		.INIT('ha8)
	) name841 (
		_w141_,
		_w177_,
		_w178_,
		_w978_
	);
	LUT3 #(
		.INIT('ha8)
	) name842 (
		_w145_,
		_w181_,
		_w182_,
		_w979_
	);
	LUT3 #(
		.INIT('ha8)
	) name843 (
		_w149_,
		_w174_,
		_w175_,
		_w980_
	);
	LUT4 #(
		.INIT('h0001)
	) name844 (
		_w977_,
		_w978_,
		_w979_,
		_w980_,
		_w981_
	);
	LUT4 #(
		.INIT('hfedc)
	) name845 (
		\shift[4] ,
		\shift[5] ,
		_w976_,
		_w981_,
		_w982_
	);
	LUT3 #(
		.INIT('h15)
	) name846 (
		\shift[6] ,
		_w971_,
		_w982_,
		_w983_
	);
	LUT3 #(
		.INIT('ha8)
	) name847 (
		_w137_,
		_w226_,
		_w227_,
		_w984_
	);
	LUT3 #(
		.INIT('ha8)
	) name848 (
		_w141_,
		_w232_,
		_w233_,
		_w985_
	);
	LUT3 #(
		.INIT('ha8)
	) name849 (
		_w145_,
		_w236_,
		_w237_,
		_w986_
	);
	LUT3 #(
		.INIT('ha8)
	) name850 (
		_w149_,
		_w229_,
		_w230_,
		_w987_
	);
	LUT4 #(
		.INIT('h0001)
	) name851 (
		_w984_,
		_w985_,
		_w986_,
		_w987_,
		_w988_
	);
	LUT3 #(
		.INIT('ha8)
	) name852 (
		_w137_,
		_w142_,
		_w143_,
		_w989_
	);
	LUT3 #(
		.INIT('ha8)
	) name853 (
		_w141_,
		_w150_,
		_w151_,
		_w990_
	);
	LUT3 #(
		.INIT('ha8)
	) name854 (
		_w145_,
		_w223_,
		_w224_,
		_w991_
	);
	LUT3 #(
		.INIT('he0)
	) name855 (
		_w146_,
		_w147_,
		_w149_,
		_w992_
	);
	LUT4 #(
		.INIT('h0001)
	) name856 (
		_w989_,
		_w990_,
		_w991_,
		_w992_,
		_w993_
	);
	LUT4 #(
		.INIT('hfdec)
	) name857 (
		\shift[4] ,
		\shift[5] ,
		_w988_,
		_w993_,
		_w994_
	);
	LUT3 #(
		.INIT('ha8)
	) name858 (
		_w137_,
		_w239_,
		_w240_,
		_w995_
	);
	LUT3 #(
		.INIT('h8a)
	) name859 (
		_w141_,
		_w245_,
		_w246_,
		_w996_
	);
	LUT3 #(
		.INIT('ha8)
	) name860 (
		_w145_,
		_w209_,
		_w210_,
		_w997_
	);
	LUT3 #(
		.INIT('ha8)
	) name861 (
		_w149_,
		_w242_,
		_w243_,
		_w998_
	);
	LUT4 #(
		.INIT('h0001)
	) name862 (
		_w995_,
		_w996_,
		_w997_,
		_w998_,
		_w999_
	);
	LUT3 #(
		.INIT('ha8)
	) name863 (
		_w137_,
		_w212_,
		_w213_,
		_w1000_
	);
	LUT3 #(
		.INIT('ha8)
	) name864 (
		_w141_,
		_w218_,
		_w219_,
		_w1001_
	);
	LUT3 #(
		.INIT('ha8)
	) name865 (
		_w145_,
		_w196_,
		_w197_,
		_w1002_
	);
	LUT3 #(
		.INIT('ha8)
	) name866 (
		_w149_,
		_w215_,
		_w216_,
		_w1003_
	);
	LUT4 #(
		.INIT('h0001)
	) name867 (
		_w1000_,
		_w1001_,
		_w1002_,
		_w1003_,
		_w1004_
	);
	LUT4 #(
		.INIT('hfb73)
	) name868 (
		\shift[4] ,
		\shift[5] ,
		_w999_,
		_w1004_,
		_w1005_
	);
	LUT3 #(
		.INIT('h2a)
	) name869 (
		\shift[6] ,
		_w994_,
		_w1005_,
		_w1006_
	);
	LUT2 #(
		.INIT('he)
	) name870 (
		_w983_,
		_w1006_,
		_w1007_
	);
	LUT3 #(
		.INIT('h8a)
	) name871 (
		_w137_,
		_w268_,
		_w269_,
		_w1008_
	);
	LUT3 #(
		.INIT('h8a)
	) name872 (
		_w141_,
		_w274_,
		_w275_,
		_w1009_
	);
	LUT3 #(
		.INIT('h8a)
	) name873 (
		_w145_,
		_w252_,
		_w253_,
		_w1010_
	);
	LUT3 #(
		.INIT('h8a)
	) name874 (
		_w149_,
		_w271_,
		_w272_,
		_w1011_
	);
	LUT4 #(
		.INIT('h0001)
	) name875 (
		_w1008_,
		_w1009_,
		_w1010_,
		_w1011_,
		_w1012_
	);
	LUT3 #(
		.INIT('h8a)
	) name876 (
		_w137_,
		_w295_,
		_w296_,
		_w1013_
	);
	LUT3 #(
		.INIT('h8a)
	) name877 (
		_w141_,
		_w301_,
		_w302_,
		_w1014_
	);
	LUT3 #(
		.INIT('h8a)
	) name878 (
		_w145_,
		_w265_,
		_w266_,
		_w1015_
	);
	LUT3 #(
		.INIT('h8a)
	) name879 (
		_w149_,
		_w298_,
		_w299_,
		_w1016_
	);
	LUT4 #(
		.INIT('h0001)
	) name880 (
		_w1013_,
		_w1014_,
		_w1015_,
		_w1016_,
		_w1017_
	);
	LUT4 #(
		.INIT('hf7b3)
	) name881 (
		\shift[4] ,
		\shift[5] ,
		_w1012_,
		_w1017_,
		_w1018_
	);
	LUT3 #(
		.INIT('h8a)
	) name882 (
		_w137_,
		_w323_,
		_w324_,
		_w1019_
	);
	LUT3 #(
		.INIT('h8a)
	) name883 (
		_w141_,
		_w329_,
		_w330_,
		_w1020_
	);
	LUT3 #(
		.INIT('h8a)
	) name884 (
		_w145_,
		_w279_,
		_w280_,
		_w1021_
	);
	LUT3 #(
		.INIT('h8a)
	) name885 (
		_w149_,
		_w326_,
		_w327_,
		_w1022_
	);
	LUT4 #(
		.INIT('h0001)
	) name886 (
		_w1019_,
		_w1020_,
		_w1021_,
		_w1022_,
		_w1023_
	);
	LUT3 #(
		.INIT('h8a)
	) name887 (
		_w137_,
		_w282_,
		_w283_,
		_w1024_
	);
	LUT3 #(
		.INIT('h8a)
	) name888 (
		_w141_,
		_w288_,
		_w289_,
		_w1025_
	);
	LUT3 #(
		.INIT('h8a)
	) name889 (
		_w145_,
		_w292_,
		_w293_,
		_w1026_
	);
	LUT3 #(
		.INIT('h8a)
	) name890 (
		_w149_,
		_w285_,
		_w286_,
		_w1027_
	);
	LUT4 #(
		.INIT('h0001)
	) name891 (
		_w1024_,
		_w1025_,
		_w1026_,
		_w1027_,
		_w1028_
	);
	LUT4 #(
		.INIT('hfedc)
	) name892 (
		\shift[4] ,
		\shift[5] ,
		_w1023_,
		_w1028_,
		_w1029_
	);
	LUT3 #(
		.INIT('h15)
	) name893 (
		\shift[6] ,
		_w1018_,
		_w1029_,
		_w1030_
	);
	LUT3 #(
		.INIT('h8a)
	) name894 (
		_w137_,
		_w310_,
		_w311_,
		_w1031_
	);
	LUT3 #(
		.INIT('h8a)
	) name895 (
		_w141_,
		_w316_,
		_w317_,
		_w1032_
	);
	LUT3 #(
		.INIT('h8a)
	) name896 (
		_w145_,
		_w334_,
		_w335_,
		_w1033_
	);
	LUT3 #(
		.INIT('h8a)
	) name897 (
		_w149_,
		_w313_,
		_w314_,
		_w1034_
	);
	LUT4 #(
		.INIT('h0001)
	) name898 (
		_w1031_,
		_w1032_,
		_w1033_,
		_w1034_,
		_w1035_
	);
	LUT3 #(
		.INIT('h8a)
	) name899 (
		_w137_,
		_w255_,
		_w256_,
		_w1036_
	);
	LUT3 #(
		.INIT('h8a)
	) name900 (
		_w141_,
		_w261_,
		_w262_,
		_w1037_
	);
	LUT3 #(
		.INIT('h8a)
	) name901 (
		_w145_,
		_w307_,
		_w308_,
		_w1038_
	);
	LUT3 #(
		.INIT('h8a)
	) name902 (
		_w149_,
		_w258_,
		_w259_,
		_w1039_
	);
	LUT4 #(
		.INIT('h0001)
	) name903 (
		_w1036_,
		_w1037_,
		_w1038_,
		_w1039_,
		_w1040_
	);
	LUT4 #(
		.INIT('hfdec)
	) name904 (
		\shift[4] ,
		\shift[5] ,
		_w1035_,
		_w1040_,
		_w1041_
	);
	LUT3 #(
		.INIT('ha8)
	) name905 (
		_w137_,
		_w337_,
		_w338_,
		_w1042_
	);
	LUT3 #(
		.INIT('ha8)
	) name906 (
		_w141_,
		_w343_,
		_w344_,
		_w1043_
	);
	LUT3 #(
		.INIT('h8a)
	) name907 (
		_w145_,
		_w347_,
		_w348_,
		_w1044_
	);
	LUT3 #(
		.INIT('h8a)
	) name908 (
		_w149_,
		_w340_,
		_w341_,
		_w1045_
	);
	LUT4 #(
		.INIT('h0001)
	) name909 (
		_w1042_,
		_w1043_,
		_w1044_,
		_w1045_,
		_w1046_
	);
	LUT3 #(
		.INIT('h8a)
	) name910 (
		_w137_,
		_w350_,
		_w351_,
		_w1047_
	);
	LUT3 #(
		.INIT('h8a)
	) name911 (
		_w141_,
		_w356_,
		_w357_,
		_w1048_
	);
	LUT3 #(
		.INIT('h8a)
	) name912 (
		_w145_,
		_w320_,
		_w321_,
		_w1049_
	);
	LUT3 #(
		.INIT('h8a)
	) name913 (
		_w149_,
		_w353_,
		_w354_,
		_w1050_
	);
	LUT4 #(
		.INIT('h0001)
	) name914 (
		_w1047_,
		_w1048_,
		_w1049_,
		_w1050_,
		_w1051_
	);
	LUT4 #(
		.INIT('hfb73)
	) name915 (
		\shift[4] ,
		\shift[5] ,
		_w1046_,
		_w1051_,
		_w1052_
	);
	LUT3 #(
		.INIT('h2a)
	) name916 (
		\shift[6] ,
		_w1041_,
		_w1052_,
		_w1053_
	);
	LUT2 #(
		.INIT('he)
	) name917 (
		_w1030_,
		_w1053_,
		_w1054_
	);
	LUT3 #(
		.INIT('ha8)
	) name918 (
		_w137_,
		_w379_,
		_w380_,
		_w1055_
	);
	LUT3 #(
		.INIT('ha8)
	) name919 (
		_w141_,
		_w385_,
		_w386_,
		_w1056_
	);
	LUT3 #(
		.INIT('ha8)
	) name920 (
		_w145_,
		_w363_,
		_w364_,
		_w1057_
	);
	LUT3 #(
		.INIT('ha8)
	) name921 (
		_w149_,
		_w382_,
		_w383_,
		_w1058_
	);
	LUT4 #(
		.INIT('h0001)
	) name922 (
		_w1055_,
		_w1056_,
		_w1057_,
		_w1058_,
		_w1059_
	);
	LUT3 #(
		.INIT('ha8)
	) name923 (
		_w137_,
		_w406_,
		_w407_,
		_w1060_
	);
	LUT3 #(
		.INIT('ha8)
	) name924 (
		_w141_,
		_w412_,
		_w413_,
		_w1061_
	);
	LUT3 #(
		.INIT('ha8)
	) name925 (
		_w145_,
		_w376_,
		_w377_,
		_w1062_
	);
	LUT3 #(
		.INIT('ha8)
	) name926 (
		_w149_,
		_w409_,
		_w410_,
		_w1063_
	);
	LUT4 #(
		.INIT('h0001)
	) name927 (
		_w1060_,
		_w1061_,
		_w1062_,
		_w1063_,
		_w1064_
	);
	LUT4 #(
		.INIT('hf7b3)
	) name928 (
		\shift[4] ,
		\shift[5] ,
		_w1059_,
		_w1064_,
		_w1065_
	);
	LUT3 #(
		.INIT('ha8)
	) name929 (
		_w137_,
		_w434_,
		_w435_,
		_w1066_
	);
	LUT3 #(
		.INIT('ha8)
	) name930 (
		_w141_,
		_w440_,
		_w441_,
		_w1067_
	);
	LUT3 #(
		.INIT('ha8)
	) name931 (
		_w145_,
		_w390_,
		_w391_,
		_w1068_
	);
	LUT3 #(
		.INIT('ha8)
	) name932 (
		_w149_,
		_w437_,
		_w438_,
		_w1069_
	);
	LUT4 #(
		.INIT('h0001)
	) name933 (
		_w1066_,
		_w1067_,
		_w1068_,
		_w1069_,
		_w1070_
	);
	LUT3 #(
		.INIT('ha8)
	) name934 (
		_w137_,
		_w393_,
		_w394_,
		_w1071_
	);
	LUT3 #(
		.INIT('ha8)
	) name935 (
		_w141_,
		_w399_,
		_w400_,
		_w1072_
	);
	LUT3 #(
		.INIT('ha8)
	) name936 (
		_w145_,
		_w403_,
		_w404_,
		_w1073_
	);
	LUT3 #(
		.INIT('ha8)
	) name937 (
		_w149_,
		_w396_,
		_w397_,
		_w1074_
	);
	LUT4 #(
		.INIT('h0001)
	) name938 (
		_w1071_,
		_w1072_,
		_w1073_,
		_w1074_,
		_w1075_
	);
	LUT4 #(
		.INIT('hfedc)
	) name939 (
		\shift[4] ,
		\shift[5] ,
		_w1070_,
		_w1075_,
		_w1076_
	);
	LUT3 #(
		.INIT('h15)
	) name940 (
		\shift[6] ,
		_w1065_,
		_w1076_,
		_w1077_
	);
	LUT3 #(
		.INIT('ha8)
	) name941 (
		_w137_,
		_w421_,
		_w422_,
		_w1078_
	);
	LUT3 #(
		.INIT('ha8)
	) name942 (
		_w141_,
		_w427_,
		_w428_,
		_w1079_
	);
	LUT3 #(
		.INIT('ha8)
	) name943 (
		_w145_,
		_w445_,
		_w446_,
		_w1080_
	);
	LUT3 #(
		.INIT('ha8)
	) name944 (
		_w149_,
		_w424_,
		_w425_,
		_w1081_
	);
	LUT4 #(
		.INIT('h0001)
	) name945 (
		_w1078_,
		_w1079_,
		_w1080_,
		_w1081_,
		_w1082_
	);
	LUT3 #(
		.INIT('ha8)
	) name946 (
		_w137_,
		_w366_,
		_w367_,
		_w1083_
	);
	LUT3 #(
		.INIT('ha8)
	) name947 (
		_w141_,
		_w372_,
		_w373_,
		_w1084_
	);
	LUT3 #(
		.INIT('ha8)
	) name948 (
		_w145_,
		_w418_,
		_w419_,
		_w1085_
	);
	LUT3 #(
		.INIT('ha8)
	) name949 (
		_w149_,
		_w369_,
		_w370_,
		_w1086_
	);
	LUT4 #(
		.INIT('h0001)
	) name950 (
		_w1083_,
		_w1084_,
		_w1085_,
		_w1086_,
		_w1087_
	);
	LUT4 #(
		.INIT('hfdec)
	) name951 (
		\shift[4] ,
		\shift[5] ,
		_w1082_,
		_w1087_,
		_w1088_
	);
	LUT3 #(
		.INIT('ha8)
	) name952 (
		_w137_,
		_w448_,
		_w449_,
		_w1089_
	);
	LUT3 #(
		.INIT('ha8)
	) name953 (
		_w141_,
		_w454_,
		_w455_,
		_w1090_
	);
	LUT3 #(
		.INIT('ha8)
	) name954 (
		_w145_,
		_w458_,
		_w459_,
		_w1091_
	);
	LUT3 #(
		.INIT('ha8)
	) name955 (
		_w149_,
		_w451_,
		_w452_,
		_w1092_
	);
	LUT4 #(
		.INIT('h0001)
	) name956 (
		_w1089_,
		_w1090_,
		_w1091_,
		_w1092_,
		_w1093_
	);
	LUT3 #(
		.INIT('ha8)
	) name957 (
		_w137_,
		_w461_,
		_w462_,
		_w1094_
	);
	LUT3 #(
		.INIT('ha8)
	) name958 (
		_w141_,
		_w467_,
		_w468_,
		_w1095_
	);
	LUT3 #(
		.INIT('ha8)
	) name959 (
		_w145_,
		_w431_,
		_w432_,
		_w1096_
	);
	LUT3 #(
		.INIT('ha8)
	) name960 (
		_w149_,
		_w464_,
		_w465_,
		_w1097_
	);
	LUT4 #(
		.INIT('h0001)
	) name961 (
		_w1094_,
		_w1095_,
		_w1096_,
		_w1097_,
		_w1098_
	);
	LUT4 #(
		.INIT('hfb73)
	) name962 (
		\shift[4] ,
		\shift[5] ,
		_w1093_,
		_w1098_,
		_w1099_
	);
	LUT3 #(
		.INIT('h2a)
	) name963 (
		\shift[6] ,
		_w1088_,
		_w1099_,
		_w1100_
	);
	LUT2 #(
		.INIT('he)
	) name964 (
		_w1077_,
		_w1100_,
		_w1101_
	);
	LUT3 #(
		.INIT('h8a)
	) name965 (
		_w137_,
		_w490_,
		_w491_,
		_w1102_
	);
	LUT3 #(
		.INIT('h8a)
	) name966 (
		_w141_,
		_w496_,
		_w497_,
		_w1103_
	);
	LUT3 #(
		.INIT('h8a)
	) name967 (
		_w145_,
		_w514_,
		_w515_,
		_w1104_
	);
	LUT3 #(
		.INIT('h8a)
	) name968 (
		_w149_,
		_w493_,
		_w494_,
		_w1105_
	);
	LUT4 #(
		.INIT('h0001)
	) name969 (
		_w1102_,
		_w1103_,
		_w1104_,
		_w1105_,
		_w1106_
	);
	LUT3 #(
		.INIT('h8a)
	) name970 (
		_w137_,
		_w477_,
		_w478_,
		_w1107_
	);
	LUT3 #(
		.INIT('h8a)
	) name971 (
		_w141_,
		_w483_,
		_w484_,
		_w1108_
	);
	LUT3 #(
		.INIT('h8a)
	) name972 (
		_w145_,
		_w487_,
		_w488_,
		_w1109_
	);
	LUT3 #(
		.INIT('h8a)
	) name973 (
		_w149_,
		_w480_,
		_w481_,
		_w1110_
	);
	LUT4 #(
		.INIT('h0001)
	) name974 (
		_w1107_,
		_w1108_,
		_w1109_,
		_w1110_,
		_w1111_
	);
	LUT4 #(
		.INIT('hf7b3)
	) name975 (
		\shift[4] ,
		\shift[5] ,
		_w1106_,
		_w1111_,
		_w1112_
	);
	LUT3 #(
		.INIT('h8a)
	) name976 (
		_w137_,
		_w559_,
		_w560_,
		_w1113_
	);
	LUT3 #(
		.INIT('h8a)
	) name977 (
		_w141_,
		_w565_,
		_w566_,
		_w1114_
	);
	LUT3 #(
		.INIT('h8a)
	) name978 (
		_w145_,
		_w501_,
		_w502_,
		_w1115_
	);
	LUT3 #(
		.INIT('h8a)
	) name979 (
		_w149_,
		_w562_,
		_w563_,
		_w1116_
	);
	LUT4 #(
		.INIT('h0001)
	) name980 (
		_w1113_,
		_w1114_,
		_w1115_,
		_w1116_,
		_w1117_
	);
	LUT3 #(
		.INIT('h8a)
	) name981 (
		_w137_,
		_w504_,
		_w505_,
		_w1118_
	);
	LUT3 #(
		.INIT('h8a)
	) name982 (
		_w141_,
		_w510_,
		_w511_,
		_w1119_
	);
	LUT3 #(
		.INIT('h8a)
	) name983 (
		_w145_,
		_w474_,
		_w475_,
		_w1120_
	);
	LUT3 #(
		.INIT('h8a)
	) name984 (
		_w149_,
		_w507_,
		_w508_,
		_w1121_
	);
	LUT4 #(
		.INIT('h0001)
	) name985 (
		_w1118_,
		_w1119_,
		_w1120_,
		_w1121_,
		_w1122_
	);
	LUT4 #(
		.INIT('hfedc)
	) name986 (
		\shift[4] ,
		\shift[5] ,
		_w1117_,
		_w1122_,
		_w1123_
	);
	LUT3 #(
		.INIT('h15)
	) name987 (
		\shift[6] ,
		_w1112_,
		_w1123_,
		_w1124_
	);
	LUT3 #(
		.INIT('h8a)
	) name988 (
		_w137_,
		_w532_,
		_w533_,
		_w1125_
	);
	LUT3 #(
		.INIT('h8a)
	) name989 (
		_w141_,
		_w538_,
		_w539_,
		_w1126_
	);
	LUT3 #(
		.INIT('h8a)
	) name990 (
		_w145_,
		_w542_,
		_w543_,
		_w1127_
	);
	LUT3 #(
		.INIT('h8a)
	) name991 (
		_w149_,
		_w535_,
		_w536_,
		_w1128_
	);
	LUT4 #(
		.INIT('h0001)
	) name992 (
		_w1125_,
		_w1126_,
		_w1127_,
		_w1128_,
		_w1129_
	);
	LUT3 #(
		.INIT('h8a)
	) name993 (
		_w137_,
		_w517_,
		_w518_,
		_w1130_
	);
	LUT3 #(
		.INIT('h8a)
	) name994 (
		_w141_,
		_w523_,
		_w524_,
		_w1131_
	);
	LUT3 #(
		.INIT('h8a)
	) name995 (
		_w145_,
		_w529_,
		_w530_,
		_w1132_
	);
	LUT3 #(
		.INIT('h8a)
	) name996 (
		_w149_,
		_w520_,
		_w521_,
		_w1133_
	);
	LUT4 #(
		.INIT('h0001)
	) name997 (
		_w1130_,
		_w1131_,
		_w1132_,
		_w1133_,
		_w1134_
	);
	LUT4 #(
		.INIT('hfdec)
	) name998 (
		\shift[4] ,
		\shift[5] ,
		_w1129_,
		_w1134_,
		_w1135_
	);
	LUT3 #(
		.INIT('ha8)
	) name999 (
		_w137_,
		_w545_,
		_w546_,
		_w1136_
	);
	LUT3 #(
		.INIT('h8a)
	) name1000 (
		_w141_,
		_w551_,
		_w552_,
		_w1137_
	);
	LUT3 #(
		.INIT('h8a)
	) name1001 (
		_w145_,
		_w569_,
		_w570_,
		_w1138_
	);
	LUT3 #(
		.INIT('h8a)
	) name1002 (
		_w149_,
		_w548_,
		_w549_,
		_w1139_
	);
	LUT4 #(
		.INIT('h0001)
	) name1003 (
		_w1136_,
		_w1137_,
		_w1138_,
		_w1139_,
		_w1140_
	);
	LUT3 #(
		.INIT('h8a)
	) name1004 (
		_w137_,
		_w572_,
		_w573_,
		_w1141_
	);
	LUT3 #(
		.INIT('h8a)
	) name1005 (
		_w141_,
		_w578_,
		_w579_,
		_w1142_
	);
	LUT3 #(
		.INIT('h8a)
	) name1006 (
		_w145_,
		_w556_,
		_w557_,
		_w1143_
	);
	LUT3 #(
		.INIT('h8a)
	) name1007 (
		_w149_,
		_w575_,
		_w576_,
		_w1144_
	);
	LUT4 #(
		.INIT('h0001)
	) name1008 (
		_w1141_,
		_w1142_,
		_w1143_,
		_w1144_,
		_w1145_
	);
	LUT4 #(
		.INIT('hfb73)
	) name1009 (
		\shift[4] ,
		\shift[5] ,
		_w1140_,
		_w1145_,
		_w1146_
	);
	LUT3 #(
		.INIT('h2a)
	) name1010 (
		\shift[6] ,
		_w1135_,
		_w1146_,
		_w1147_
	);
	LUT2 #(
		.INIT('he)
	) name1011 (
		_w1124_,
		_w1147_,
		_w1148_
	);
	LUT4 #(
		.INIT('hf7b3)
	) name1012 (
		\shift[4] ,
		\shift[5] ,
		_w166_,
		_w193_,
		_w1149_
	);
	LUT4 #(
		.INIT('hfdec)
	) name1013 (
		\shift[4] ,
		\shift[5] ,
		_w180_,
		_w208_,
		_w1150_
	);
	LUT3 #(
		.INIT('h15)
	) name1014 (
		\shift[6] ,
		_w1149_,
		_w1150_,
		_w1151_
	);
	LUT4 #(
		.INIT('hfe76)
	) name1015 (
		\shift[4] ,
		\shift[5] ,
		_w153_,
		_w221_,
		_w1152_
	);
	LUT4 #(
		.INIT('hfdb9)
	) name1016 (
		\shift[4] ,
		\shift[5] ,
		_w235_,
		_w248_,
		_w1153_
	);
	LUT3 #(
		.INIT('h2a)
	) name1017 (
		\shift[6] ,
		_w1152_,
		_w1153_,
		_w1154_
	);
	LUT2 #(
		.INIT('he)
	) name1018 (
		_w1151_,
		_w1154_,
		_w1155_
	);
	LUT4 #(
		.INIT('hf7b3)
	) name1019 (
		\shift[4] ,
		\shift[5] ,
		_w277_,
		_w304_,
		_w1156_
	);
	LUT4 #(
		.INIT('hfdec)
	) name1020 (
		\shift[4] ,
		\shift[5] ,
		_w291_,
		_w332_,
		_w1157_
	);
	LUT3 #(
		.INIT('h15)
	) name1021 (
		\shift[6] ,
		_w1156_,
		_w1157_,
		_w1158_
	);
	LUT4 #(
		.INIT('hfedc)
	) name1022 (
		\shift[4] ,
		\shift[5] ,
		_w264_,
		_w319_,
		_w1159_
	);
	LUT4 #(
		.INIT('hfb73)
	) name1023 (
		\shift[4] ,
		\shift[5] ,
		_w346_,
		_w359_,
		_w1160_
	);
	LUT3 #(
		.INIT('h2a)
	) name1024 (
		\shift[6] ,
		_w1159_,
		_w1160_,
		_w1161_
	);
	LUT2 #(
		.INIT('he)
	) name1025 (
		_w1158_,
		_w1161_,
		_w1162_
	);
	LUT4 #(
		.INIT('hf7b3)
	) name1026 (
		\shift[4] ,
		\shift[5] ,
		_w388_,
		_w415_,
		_w1163_
	);
	LUT4 #(
		.INIT('hfdec)
	) name1027 (
		\shift[4] ,
		\shift[5] ,
		_w402_,
		_w443_,
		_w1164_
	);
	LUT3 #(
		.INIT('h15)
	) name1028 (
		\shift[6] ,
		_w1163_,
		_w1164_,
		_w1165_
	);
	LUT4 #(
		.INIT('hfedc)
	) name1029 (
		\shift[4] ,
		\shift[5] ,
		_w375_,
		_w430_,
		_w1166_
	);
	LUT4 #(
		.INIT('hfb73)
	) name1030 (
		\shift[4] ,
		\shift[5] ,
		_w457_,
		_w470_,
		_w1167_
	);
	LUT3 #(
		.INIT('h2a)
	) name1031 (
		\shift[6] ,
		_w1166_,
		_w1167_,
		_w1168_
	);
	LUT2 #(
		.INIT('he)
	) name1032 (
		_w1165_,
		_w1168_,
		_w1169_
	);
	LUT4 #(
		.INIT('hfb73)
	) name1033 (
		\shift[4] ,
		\shift[5] ,
		_w486_,
		_w499_,
		_w1170_
	);
	LUT4 #(
		.INIT('hfdec)
	) name1034 (
		\shift[4] ,
		\shift[5] ,
		_w513_,
		_w568_,
		_w1171_
	);
	LUT3 #(
		.INIT('h15)
	) name1035 (
		\shift[6] ,
		_w1170_,
		_w1171_,
		_w1172_
	);
	LUT4 #(
		.INIT('hfedc)
	) name1036 (
		\shift[4] ,
		\shift[5] ,
		_w526_,
		_w541_,
		_w1173_
	);
	LUT4 #(
		.INIT('hfb73)
	) name1037 (
		\shift[4] ,
		\shift[5] ,
		_w554_,
		_w581_,
		_w1174_
	);
	LUT3 #(
		.INIT('h2a)
	) name1038 (
		\shift[6] ,
		_w1173_,
		_w1174_,
		_w1175_
	);
	LUT2 #(
		.INIT('he)
	) name1039 (
		_w1172_,
		_w1175_,
		_w1176_
	);
	LUT4 #(
		.INIT('hf7b3)
	) name1040 (
		\shift[4] ,
		\shift[5] ,
		_w594_,
		_w605_,
		_w1177_
	);
	LUT4 #(
		.INIT('hfdec)
	) name1041 (
		\shift[4] ,
		\shift[5] ,
		_w600_,
		_w628_,
		_w1178_
	);
	LUT3 #(
		.INIT('h15)
	) name1042 (
		\shift[6] ,
		_w1177_,
		_w1178_,
		_w1179_
	);
	LUT4 #(
		.INIT('hfeba)
	) name1043 (
		\shift[4] ,
		\shift[5] ,
		_w589_,
		_w612_,
		_w1180_
	);
	LUT4 #(
		.INIT('hfd75)
	) name1044 (
		\shift[4] ,
		\shift[5] ,
		_w617_,
		_w623_,
		_w1181_
	);
	LUT3 #(
		.INIT('h2a)
	) name1045 (
		\shift[6] ,
		_w1180_,
		_w1181_,
		_w1182_
	);
	LUT2 #(
		.INIT('he)
	) name1046 (
		_w1179_,
		_w1182_,
		_w1183_
	);
	LUT4 #(
		.INIT('hf7b3)
	) name1047 (
		\shift[4] ,
		\shift[5] ,
		_w641_,
		_w652_,
		_w1184_
	);
	LUT4 #(
		.INIT('hfdec)
	) name1048 (
		\shift[4] ,
		\shift[5] ,
		_w647_,
		_w675_,
		_w1185_
	);
	LUT3 #(
		.INIT('h15)
	) name1049 (
		\shift[6] ,
		_w1184_,
		_w1185_,
		_w1186_
	);
	LUT4 #(
		.INIT('hfeba)
	) name1050 (
		\shift[4] ,
		\shift[5] ,
		_w636_,
		_w659_,
		_w1187_
	);
	LUT4 #(
		.INIT('hfd75)
	) name1051 (
		\shift[4] ,
		\shift[5] ,
		_w664_,
		_w670_,
		_w1188_
	);
	LUT3 #(
		.INIT('h2a)
	) name1052 (
		\shift[6] ,
		_w1187_,
		_w1188_,
		_w1189_
	);
	LUT2 #(
		.INIT('he)
	) name1053 (
		_w1186_,
		_w1189_,
		_w1190_
	);
	LUT4 #(
		.INIT('hf7b3)
	) name1054 (
		\shift[4] ,
		\shift[5] ,
		_w688_,
		_w699_,
		_w1191_
	);
	LUT4 #(
		.INIT('hfdec)
	) name1055 (
		\shift[4] ,
		\shift[5] ,
		_w694_,
		_w722_,
		_w1192_
	);
	LUT3 #(
		.INIT('h15)
	) name1056 (
		\shift[6] ,
		_w1191_,
		_w1192_,
		_w1193_
	);
	LUT4 #(
		.INIT('hfeba)
	) name1057 (
		\shift[4] ,
		\shift[5] ,
		_w683_,
		_w706_,
		_w1194_
	);
	LUT4 #(
		.INIT('hfd75)
	) name1058 (
		\shift[4] ,
		\shift[5] ,
		_w711_,
		_w717_,
		_w1195_
	);
	LUT3 #(
		.INIT('h2a)
	) name1059 (
		\shift[6] ,
		_w1194_,
		_w1195_,
		_w1196_
	);
	LUT2 #(
		.INIT('he)
	) name1060 (
		_w1193_,
		_w1196_,
		_w1197_
	);
	LUT4 #(
		.INIT('hf7e6)
	) name1061 (
		\shift[4] ,
		\shift[5] ,
		_w735_,
		_w769_,
		_w1198_
	);
	LUT4 #(
		.INIT('hfdb9)
	) name1062 (
		\shift[4] ,
		\shift[5] ,
		_w741_,
		_w746_,
		_w1199_
	);
	LUT3 #(
		.INIT('h15)
	) name1063 (
		\shift[6] ,
		_w1198_,
		_w1199_,
		_w1200_
	);
	LUT4 #(
		.INIT('hfbd9)
	) name1064 (
		\shift[4] ,
		\shift[5] ,
		_w753_,
		_w758_,
		_w1201_
	);
	LUT4 #(
		.INIT('hfe76)
	) name1065 (
		\shift[4] ,
		\shift[5] ,
		_w730_,
		_w764_,
		_w1202_
	);
	LUT3 #(
		.INIT('h2a)
	) name1066 (
		\shift[6] ,
		_w1201_,
		_w1202_,
		_w1203_
	);
	LUT2 #(
		.INIT('he)
	) name1067 (
		_w1200_,
		_w1203_,
		_w1204_
	);
	LUT4 #(
		.INIT('hf7e6)
	) name1068 (
		\shift[4] ,
		\shift[5] ,
		_w782_,
		_w816_,
		_w1205_
	);
	LUT4 #(
		.INIT('hfdb9)
	) name1069 (
		\shift[4] ,
		\shift[5] ,
		_w788_,
		_w793_,
		_w1206_
	);
	LUT3 #(
		.INIT('h15)
	) name1070 (
		\shift[6] ,
		_w1205_,
		_w1206_,
		_w1207_
	);
	LUT4 #(
		.INIT('hfbd9)
	) name1071 (
		\shift[4] ,
		\shift[5] ,
		_w800_,
		_w805_,
		_w1208_
	);
	LUT4 #(
		.INIT('hfe76)
	) name1072 (
		\shift[4] ,
		\shift[5] ,
		_w777_,
		_w811_,
		_w1209_
	);
	LUT3 #(
		.INIT('h2a)
	) name1073 (
		\shift[6] ,
		_w1208_,
		_w1209_,
		_w1210_
	);
	LUT2 #(
		.INIT('he)
	) name1074 (
		_w1207_,
		_w1210_,
		_w1211_
	);
	LUT4 #(
		.INIT('hf7e6)
	) name1075 (
		\shift[4] ,
		\shift[5] ,
		_w829_,
		_w863_,
		_w1212_
	);
	LUT4 #(
		.INIT('hfdb9)
	) name1076 (
		\shift[4] ,
		\shift[5] ,
		_w835_,
		_w840_,
		_w1213_
	);
	LUT3 #(
		.INIT('h15)
	) name1077 (
		\shift[6] ,
		_w1212_,
		_w1213_,
		_w1214_
	);
	LUT4 #(
		.INIT('hfbd9)
	) name1078 (
		\shift[4] ,
		\shift[5] ,
		_w847_,
		_w852_,
		_w1215_
	);
	LUT4 #(
		.INIT('hfe76)
	) name1079 (
		\shift[4] ,
		\shift[5] ,
		_w824_,
		_w858_,
		_w1216_
	);
	LUT3 #(
		.INIT('h2a)
	) name1080 (
		\shift[6] ,
		_w1215_,
		_w1216_,
		_w1217_
	);
	LUT2 #(
		.INIT('he)
	) name1081 (
		_w1214_,
		_w1217_,
		_w1218_
	);
	LUT4 #(
		.INIT('hf7b3)
	) name1082 (
		\shift[4] ,
		\shift[5] ,
		_w876_,
		_w887_,
		_w1219_
	);
	LUT4 #(
		.INIT('hfdec)
	) name1083 (
		\shift[4] ,
		\shift[5] ,
		_w882_,
		_w910_,
		_w1220_
	);
	LUT3 #(
		.INIT('h15)
	) name1084 (
		\shift[6] ,
		_w1219_,
		_w1220_,
		_w1221_
	);
	LUT4 #(
		.INIT('hfbd9)
	) name1085 (
		\shift[4] ,
		\shift[5] ,
		_w894_,
		_w899_,
		_w1222_
	);
	LUT4 #(
		.INIT('hfe76)
	) name1086 (
		\shift[4] ,
		\shift[5] ,
		_w871_,
		_w905_,
		_w1223_
	);
	LUT3 #(
		.INIT('h2a)
	) name1087 (
		\shift[6] ,
		_w1222_,
		_w1223_,
		_w1224_
	);
	LUT2 #(
		.INIT('he)
	) name1088 (
		_w1221_,
		_w1224_,
		_w1225_
	);
	LUT4 #(
		.INIT('hf7b3)
	) name1089 (
		\shift[4] ,
		\shift[5] ,
		_w923_,
		_w934_,
		_w1226_
	);
	LUT4 #(
		.INIT('hfdec)
	) name1090 (
		\shift[4] ,
		\shift[5] ,
		_w929_,
		_w957_,
		_w1227_
	);
	LUT3 #(
		.INIT('h15)
	) name1091 (
		\shift[6] ,
		_w1226_,
		_w1227_,
		_w1228_
	);
	LUT4 #(
		.INIT('hfbd9)
	) name1092 (
		\shift[4] ,
		\shift[5] ,
		_w941_,
		_w946_,
		_w1229_
	);
	LUT4 #(
		.INIT('hfe76)
	) name1093 (
		\shift[4] ,
		\shift[5] ,
		_w918_,
		_w952_,
		_w1230_
	);
	LUT3 #(
		.INIT('h2a)
	) name1094 (
		\shift[6] ,
		_w1229_,
		_w1230_,
		_w1231_
	);
	LUT2 #(
		.INIT('he)
	) name1095 (
		_w1228_,
		_w1231_,
		_w1232_
	);
	LUT4 #(
		.INIT('hf7b3)
	) name1096 (
		\shift[4] ,
		\shift[5] ,
		_w970_,
		_w981_,
		_w1233_
	);
	LUT4 #(
		.INIT('hfdec)
	) name1097 (
		\shift[4] ,
		\shift[5] ,
		_w976_,
		_w1004_,
		_w1234_
	);
	LUT3 #(
		.INIT('h15)
	) name1098 (
		\shift[6] ,
		_w1233_,
		_w1234_,
		_w1235_
	);
	LUT4 #(
		.INIT('hfbd9)
	) name1099 (
		\shift[4] ,
		\shift[5] ,
		_w988_,
		_w993_,
		_w1236_
	);
	LUT4 #(
		.INIT('hfe76)
	) name1100 (
		\shift[4] ,
		\shift[5] ,
		_w965_,
		_w999_,
		_w1237_
	);
	LUT3 #(
		.INIT('h2a)
	) name1101 (
		\shift[6] ,
		_w1236_,
		_w1237_,
		_w1238_
	);
	LUT2 #(
		.INIT('he)
	) name1102 (
		_w1235_,
		_w1238_,
		_w1239_
	);
	LUT4 #(
		.INIT('hf7b3)
	) name1103 (
		\shift[4] ,
		\shift[5] ,
		_w1017_,
		_w1028_,
		_w1240_
	);
	LUT4 #(
		.INIT('hfdec)
	) name1104 (
		\shift[4] ,
		\shift[5] ,
		_w1023_,
		_w1051_,
		_w1241_
	);
	LUT3 #(
		.INIT('h15)
	) name1105 (
		\shift[6] ,
		_w1240_,
		_w1241_,
		_w1242_
	);
	LUT4 #(
		.INIT('hfbd9)
	) name1106 (
		\shift[4] ,
		\shift[5] ,
		_w1035_,
		_w1040_,
		_w1243_
	);
	LUT4 #(
		.INIT('hfe76)
	) name1107 (
		\shift[4] ,
		\shift[5] ,
		_w1012_,
		_w1046_,
		_w1244_
	);
	LUT3 #(
		.INIT('h2a)
	) name1108 (
		\shift[6] ,
		_w1243_,
		_w1244_,
		_w1245_
	);
	LUT2 #(
		.INIT('he)
	) name1109 (
		_w1242_,
		_w1245_,
		_w1246_
	);
	LUT4 #(
		.INIT('hf7b3)
	) name1110 (
		\shift[4] ,
		\shift[5] ,
		_w1064_,
		_w1075_,
		_w1247_
	);
	LUT4 #(
		.INIT('hfdec)
	) name1111 (
		\shift[4] ,
		\shift[5] ,
		_w1070_,
		_w1098_,
		_w1248_
	);
	LUT3 #(
		.INIT('h15)
	) name1112 (
		\shift[6] ,
		_w1247_,
		_w1248_,
		_w1249_
	);
	LUT4 #(
		.INIT('hfbd9)
	) name1113 (
		\shift[4] ,
		\shift[5] ,
		_w1082_,
		_w1087_,
		_w1250_
	);
	LUT4 #(
		.INIT('hfe76)
	) name1114 (
		\shift[4] ,
		\shift[5] ,
		_w1059_,
		_w1093_,
		_w1251_
	);
	LUT3 #(
		.INIT('h2a)
	) name1115 (
		\shift[6] ,
		_w1250_,
		_w1251_,
		_w1252_
	);
	LUT2 #(
		.INIT('he)
	) name1116 (
		_w1249_,
		_w1252_,
		_w1253_
	);
	LUT4 #(
		.INIT('hf7b3)
	) name1117 (
		\shift[4] ,
		\shift[5] ,
		_w1111_,
		_w1122_,
		_w1254_
	);
	LUT4 #(
		.INIT('hfdec)
	) name1118 (
		\shift[4] ,
		\shift[5] ,
		_w1117_,
		_w1145_,
		_w1255_
	);
	LUT3 #(
		.INIT('h15)
	) name1119 (
		\shift[6] ,
		_w1254_,
		_w1255_,
		_w1256_
	);
	LUT4 #(
		.INIT('hfbd9)
	) name1120 (
		\shift[4] ,
		\shift[5] ,
		_w1129_,
		_w1134_,
		_w1257_
	);
	LUT4 #(
		.INIT('hfe76)
	) name1121 (
		\shift[4] ,
		\shift[5] ,
		_w1106_,
		_w1140_,
		_w1258_
	);
	LUT3 #(
		.INIT('h2a)
	) name1122 (
		\shift[6] ,
		_w1257_,
		_w1258_,
		_w1259_
	);
	LUT2 #(
		.INIT('he)
	) name1123 (
		_w1256_,
		_w1259_,
		_w1260_
	);
	LUT4 #(
		.INIT('hfb73)
	) name1124 (
		\shift[4] ,
		\shift[5] ,
		_w180_,
		_w193_,
		_w1261_
	);
	LUT4 #(
		.INIT('hfdec)
	) name1125 (
		\shift[4] ,
		\shift[5] ,
		_w208_,
		_w221_,
		_w1262_
	);
	LUT3 #(
		.INIT('h15)
	) name1126 (
		\shift[6] ,
		_w1261_,
		_w1262_,
		_w1263_
	);
	LUT4 #(
		.INIT('hfdec)
	) name1127 (
		\shift[4] ,
		\shift[5] ,
		_w153_,
		_w166_,
		_w1264_
	);
	LUT4 #(
		.INIT('hfb73)
	) name1128 (
		\shift[4] ,
		\shift[5] ,
		_w235_,
		_w248_,
		_w1265_
	);
	LUT3 #(
		.INIT('h2a)
	) name1129 (
		\shift[6] ,
		_w1264_,
		_w1265_,
		_w1266_
	);
	LUT2 #(
		.INIT('he)
	) name1130 (
		_w1263_,
		_w1266_,
		_w1267_
	);
	LUT4 #(
		.INIT('hfb73)
	) name1131 (
		\shift[4] ,
		\shift[5] ,
		_w291_,
		_w304_,
		_w1268_
	);
	LUT4 #(
		.INIT('hfdec)
	) name1132 (
		\shift[4] ,
		\shift[5] ,
		_w332_,
		_w359_,
		_w1269_
	);
	LUT3 #(
		.INIT('h15)
	) name1133 (
		\shift[6] ,
		_w1268_,
		_w1269_,
		_w1270_
	);
	LUT4 #(
		.INIT('hfdb9)
	) name1134 (
		\shift[4] ,
		\shift[5] ,
		_w264_,
		_w319_,
		_w1271_
	);
	LUT4 #(
		.INIT('hfe76)
	) name1135 (
		\shift[4] ,
		\shift[5] ,
		_w277_,
		_w346_,
		_w1272_
	);
	LUT3 #(
		.INIT('h2a)
	) name1136 (
		\shift[6] ,
		_w1271_,
		_w1272_,
		_w1273_
	);
	LUT2 #(
		.INIT('he)
	) name1137 (
		_w1270_,
		_w1273_,
		_w1274_
	);
	LUT4 #(
		.INIT('hfb73)
	) name1138 (
		\shift[4] ,
		\shift[5] ,
		_w402_,
		_w415_,
		_w1275_
	);
	LUT4 #(
		.INIT('hfdec)
	) name1139 (
		\shift[4] ,
		\shift[5] ,
		_w443_,
		_w470_,
		_w1276_
	);
	LUT3 #(
		.INIT('h15)
	) name1140 (
		\shift[6] ,
		_w1275_,
		_w1276_,
		_w1277_
	);
	LUT4 #(
		.INIT('hfdb9)
	) name1141 (
		\shift[4] ,
		\shift[5] ,
		_w375_,
		_w430_,
		_w1278_
	);
	LUT4 #(
		.INIT('hfe76)
	) name1142 (
		\shift[4] ,
		\shift[5] ,
		_w388_,
		_w457_,
		_w1279_
	);
	LUT3 #(
		.INIT('h2a)
	) name1143 (
		\shift[6] ,
		_w1278_,
		_w1279_,
		_w1280_
	);
	LUT2 #(
		.INIT('he)
	) name1144 (
		_w1277_,
		_w1280_,
		_w1281_
	);
	LUT4 #(
		.INIT('hf7e6)
	) name1145 (
		\shift[4] ,
		\shift[5] ,
		_w486_,
		_w581_,
		_w1282_
	);
	LUT4 #(
		.INIT('hfbd9)
	) name1146 (
		\shift[4] ,
		\shift[5] ,
		_w513_,
		_w568_,
		_w1283_
	);
	LUT3 #(
		.INIT('h15)
	) name1147 (
		\shift[6] ,
		_w1282_,
		_w1283_,
		_w1284_
	);
	LUT4 #(
		.INIT('hfeba)
	) name1148 (
		\shift[4] ,
		\shift[5] ,
		_w499_,
		_w541_,
		_w1285_
	);
	LUT4 #(
		.INIT('hfd75)
	) name1149 (
		\shift[4] ,
		\shift[5] ,
		_w526_,
		_w554_,
		_w1286_
	);
	LUT3 #(
		.INIT('h2a)
	) name1150 (
		\shift[6] ,
		_w1285_,
		_w1286_,
		_w1287_
	);
	LUT2 #(
		.INIT('he)
	) name1151 (
		_w1284_,
		_w1287_,
		_w1288_
	);
	LUT4 #(
		.INIT('hfb73)
	) name1152 (
		\shift[4] ,
		\shift[5] ,
		_w600_,
		_w605_,
		_w1289_
	);
	LUT4 #(
		.INIT('hfedc)
	) name1153 (
		\shift[4] ,
		\shift[5] ,
		_w623_,
		_w628_,
		_w1290_
	);
	LUT3 #(
		.INIT('h15)
	) name1154 (
		\shift[6] ,
		_w1289_,
		_w1290_,
		_w1291_
	);
	LUT4 #(
		.INIT('hfdec)
	) name1155 (
		\shift[4] ,
		\shift[5] ,
		_w589_,
		_w594_,
		_w1292_
	);
	LUT4 #(
		.INIT('hf7b3)
	) name1156 (
		\shift[4] ,
		\shift[5] ,
		_w612_,
		_w617_,
		_w1293_
	);
	LUT3 #(
		.INIT('h2a)
	) name1157 (
		\shift[6] ,
		_w1292_,
		_w1293_,
		_w1294_
	);
	LUT2 #(
		.INIT('he)
	) name1158 (
		_w1291_,
		_w1294_,
		_w1295_
	);
	LUT4 #(
		.INIT('hfb73)
	) name1159 (
		\shift[4] ,
		\shift[5] ,
		_w647_,
		_w652_,
		_w1296_
	);
	LUT4 #(
		.INIT('hfedc)
	) name1160 (
		\shift[4] ,
		\shift[5] ,
		_w670_,
		_w675_,
		_w1297_
	);
	LUT3 #(
		.INIT('h15)
	) name1161 (
		\shift[6] ,
		_w1296_,
		_w1297_,
		_w1298_
	);
	LUT4 #(
		.INIT('hfdec)
	) name1162 (
		\shift[4] ,
		\shift[5] ,
		_w636_,
		_w641_,
		_w1299_
	);
	LUT4 #(
		.INIT('hf7b3)
	) name1163 (
		\shift[4] ,
		\shift[5] ,
		_w659_,
		_w664_,
		_w1300_
	);
	LUT3 #(
		.INIT('h2a)
	) name1164 (
		\shift[6] ,
		_w1299_,
		_w1300_,
		_w1301_
	);
	LUT2 #(
		.INIT('he)
	) name1165 (
		_w1298_,
		_w1301_,
		_w1302_
	);
	LUT4 #(
		.INIT('hfb73)
	) name1166 (
		\shift[4] ,
		\shift[5] ,
		_w694_,
		_w699_,
		_w1303_
	);
	LUT4 #(
		.INIT('hfedc)
	) name1167 (
		\shift[4] ,
		\shift[5] ,
		_w717_,
		_w722_,
		_w1304_
	);
	LUT3 #(
		.INIT('h15)
	) name1168 (
		\shift[6] ,
		_w1303_,
		_w1304_,
		_w1305_
	);
	LUT4 #(
		.INIT('hfdec)
	) name1169 (
		\shift[4] ,
		\shift[5] ,
		_w683_,
		_w688_,
		_w1306_
	);
	LUT4 #(
		.INIT('hf7b3)
	) name1170 (
		\shift[4] ,
		\shift[5] ,
		_w706_,
		_w711_,
		_w1307_
	);
	LUT3 #(
		.INIT('h2a)
	) name1171 (
		\shift[6] ,
		_w1306_,
		_w1307_,
		_w1308_
	);
	LUT2 #(
		.INIT('he)
	) name1172 (
		_w1305_,
		_w1308_,
		_w1309_
	);
	LUT4 #(
		.INIT('hfedc)
	) name1173 (
		\shift[4] ,
		\shift[5] ,
		_w764_,
		_w769_,
		_w1310_
	);
	LUT4 #(
		.INIT('hfb73)
	) name1174 (
		\shift[4] ,
		\shift[5] ,
		_w741_,
		_w746_,
		_w1311_
	);
	LUT3 #(
		.INIT('h15)
	) name1175 (
		\shift[6] ,
		_w1310_,
		_w1311_,
		_w1312_
	);
	LUT4 #(
		.INIT('hf7b3)
	) name1176 (
		\shift[4] ,
		\shift[5] ,
		_w753_,
		_w758_,
		_w1313_
	);
	LUT4 #(
		.INIT('hfdec)
	) name1177 (
		\shift[4] ,
		\shift[5] ,
		_w730_,
		_w735_,
		_w1314_
	);
	LUT3 #(
		.INIT('h2a)
	) name1178 (
		\shift[6] ,
		_w1313_,
		_w1314_,
		_w1315_
	);
	LUT2 #(
		.INIT('he)
	) name1179 (
		_w1312_,
		_w1315_,
		_w1316_
	);
	LUT4 #(
		.INIT('hfedc)
	) name1180 (
		\shift[4] ,
		\shift[5] ,
		_w811_,
		_w816_,
		_w1317_
	);
	LUT4 #(
		.INIT('hfb73)
	) name1181 (
		\shift[4] ,
		\shift[5] ,
		_w788_,
		_w793_,
		_w1318_
	);
	LUT3 #(
		.INIT('h15)
	) name1182 (
		\shift[6] ,
		_w1317_,
		_w1318_,
		_w1319_
	);
	LUT4 #(
		.INIT('hf7b3)
	) name1183 (
		\shift[4] ,
		\shift[5] ,
		_w800_,
		_w805_,
		_w1320_
	);
	LUT4 #(
		.INIT('hfdec)
	) name1184 (
		\shift[4] ,
		\shift[5] ,
		_w777_,
		_w782_,
		_w1321_
	);
	LUT3 #(
		.INIT('h2a)
	) name1185 (
		\shift[6] ,
		_w1320_,
		_w1321_,
		_w1322_
	);
	LUT2 #(
		.INIT('he)
	) name1186 (
		_w1319_,
		_w1322_,
		_w1323_
	);
	LUT4 #(
		.INIT('hfedc)
	) name1187 (
		\shift[4] ,
		\shift[5] ,
		_w858_,
		_w863_,
		_w1324_
	);
	LUT4 #(
		.INIT('hfb73)
	) name1188 (
		\shift[4] ,
		\shift[5] ,
		_w835_,
		_w840_,
		_w1325_
	);
	LUT3 #(
		.INIT('h15)
	) name1189 (
		\shift[6] ,
		_w1324_,
		_w1325_,
		_w1326_
	);
	LUT4 #(
		.INIT('hf7b3)
	) name1190 (
		\shift[4] ,
		\shift[5] ,
		_w847_,
		_w852_,
		_w1327_
	);
	LUT4 #(
		.INIT('hfdec)
	) name1191 (
		\shift[4] ,
		\shift[5] ,
		_w824_,
		_w829_,
		_w1328_
	);
	LUT3 #(
		.INIT('h2a)
	) name1192 (
		\shift[6] ,
		_w1327_,
		_w1328_,
		_w1329_
	);
	LUT2 #(
		.INIT('he)
	) name1193 (
		_w1326_,
		_w1329_,
		_w1330_
	);
	LUT4 #(
		.INIT('hfb73)
	) name1194 (
		\shift[4] ,
		\shift[5] ,
		_w882_,
		_w887_,
		_w1331_
	);
	LUT4 #(
		.INIT('hfedc)
	) name1195 (
		\shift[4] ,
		\shift[5] ,
		_w905_,
		_w910_,
		_w1332_
	);
	LUT3 #(
		.INIT('h15)
	) name1196 (
		\shift[6] ,
		_w1331_,
		_w1332_,
		_w1333_
	);
	LUT4 #(
		.INIT('hf7b3)
	) name1197 (
		\shift[4] ,
		\shift[5] ,
		_w894_,
		_w899_,
		_w1334_
	);
	LUT4 #(
		.INIT('hfdec)
	) name1198 (
		\shift[4] ,
		\shift[5] ,
		_w871_,
		_w876_,
		_w1335_
	);
	LUT3 #(
		.INIT('h2a)
	) name1199 (
		\shift[6] ,
		_w1334_,
		_w1335_,
		_w1336_
	);
	LUT2 #(
		.INIT('he)
	) name1200 (
		_w1333_,
		_w1336_,
		_w1337_
	);
	LUT4 #(
		.INIT('hfb73)
	) name1201 (
		\shift[4] ,
		\shift[5] ,
		_w929_,
		_w934_,
		_w1338_
	);
	LUT4 #(
		.INIT('hfedc)
	) name1202 (
		\shift[4] ,
		\shift[5] ,
		_w952_,
		_w957_,
		_w1339_
	);
	LUT3 #(
		.INIT('h15)
	) name1203 (
		\shift[6] ,
		_w1338_,
		_w1339_,
		_w1340_
	);
	LUT4 #(
		.INIT('hf7b3)
	) name1204 (
		\shift[4] ,
		\shift[5] ,
		_w941_,
		_w946_,
		_w1341_
	);
	LUT4 #(
		.INIT('hfdec)
	) name1205 (
		\shift[4] ,
		\shift[5] ,
		_w918_,
		_w923_,
		_w1342_
	);
	LUT3 #(
		.INIT('h2a)
	) name1206 (
		\shift[6] ,
		_w1341_,
		_w1342_,
		_w1343_
	);
	LUT2 #(
		.INIT('he)
	) name1207 (
		_w1340_,
		_w1343_,
		_w1344_
	);
	LUT4 #(
		.INIT('hfb73)
	) name1208 (
		\shift[4] ,
		\shift[5] ,
		_w976_,
		_w981_,
		_w1345_
	);
	LUT4 #(
		.INIT('hfedc)
	) name1209 (
		\shift[4] ,
		\shift[5] ,
		_w999_,
		_w1004_,
		_w1346_
	);
	LUT3 #(
		.INIT('h15)
	) name1210 (
		\shift[6] ,
		_w1345_,
		_w1346_,
		_w1347_
	);
	LUT4 #(
		.INIT('hf7b3)
	) name1211 (
		\shift[4] ,
		\shift[5] ,
		_w988_,
		_w993_,
		_w1348_
	);
	LUT4 #(
		.INIT('hfdec)
	) name1212 (
		\shift[4] ,
		\shift[5] ,
		_w965_,
		_w970_,
		_w1349_
	);
	LUT3 #(
		.INIT('h2a)
	) name1213 (
		\shift[6] ,
		_w1348_,
		_w1349_,
		_w1350_
	);
	LUT2 #(
		.INIT('he)
	) name1214 (
		_w1347_,
		_w1350_,
		_w1351_
	);
	LUT4 #(
		.INIT('hfb73)
	) name1215 (
		\shift[4] ,
		\shift[5] ,
		_w1023_,
		_w1028_,
		_w1352_
	);
	LUT4 #(
		.INIT('hfedc)
	) name1216 (
		\shift[4] ,
		\shift[5] ,
		_w1046_,
		_w1051_,
		_w1353_
	);
	LUT3 #(
		.INIT('h15)
	) name1217 (
		\shift[6] ,
		_w1352_,
		_w1353_,
		_w1354_
	);
	LUT4 #(
		.INIT('hf7b3)
	) name1218 (
		\shift[4] ,
		\shift[5] ,
		_w1035_,
		_w1040_,
		_w1355_
	);
	LUT4 #(
		.INIT('hfdec)
	) name1219 (
		\shift[4] ,
		\shift[5] ,
		_w1012_,
		_w1017_,
		_w1356_
	);
	LUT3 #(
		.INIT('h2a)
	) name1220 (
		\shift[6] ,
		_w1355_,
		_w1356_,
		_w1357_
	);
	LUT2 #(
		.INIT('he)
	) name1221 (
		_w1354_,
		_w1357_,
		_w1358_
	);
	LUT4 #(
		.INIT('hfb73)
	) name1222 (
		\shift[4] ,
		\shift[5] ,
		_w1070_,
		_w1075_,
		_w1359_
	);
	LUT4 #(
		.INIT('hfedc)
	) name1223 (
		\shift[4] ,
		\shift[5] ,
		_w1093_,
		_w1098_,
		_w1360_
	);
	LUT3 #(
		.INIT('h15)
	) name1224 (
		\shift[6] ,
		_w1359_,
		_w1360_,
		_w1361_
	);
	LUT4 #(
		.INIT('hf7b3)
	) name1225 (
		\shift[4] ,
		\shift[5] ,
		_w1082_,
		_w1087_,
		_w1362_
	);
	LUT4 #(
		.INIT('hfdec)
	) name1226 (
		\shift[4] ,
		\shift[5] ,
		_w1059_,
		_w1064_,
		_w1363_
	);
	LUT3 #(
		.INIT('h2a)
	) name1227 (
		\shift[6] ,
		_w1362_,
		_w1363_,
		_w1364_
	);
	LUT2 #(
		.INIT('he)
	) name1228 (
		_w1361_,
		_w1364_,
		_w1365_
	);
	LUT4 #(
		.INIT('hfb73)
	) name1229 (
		\shift[4] ,
		\shift[5] ,
		_w1117_,
		_w1122_,
		_w1366_
	);
	LUT4 #(
		.INIT('hfedc)
	) name1230 (
		\shift[4] ,
		\shift[5] ,
		_w1140_,
		_w1145_,
		_w1367_
	);
	LUT3 #(
		.INIT('h15)
	) name1231 (
		\shift[6] ,
		_w1366_,
		_w1367_,
		_w1368_
	);
	LUT4 #(
		.INIT('hf7b3)
	) name1232 (
		\shift[4] ,
		\shift[5] ,
		_w1129_,
		_w1134_,
		_w1369_
	);
	LUT4 #(
		.INIT('hfdec)
	) name1233 (
		\shift[4] ,
		\shift[5] ,
		_w1106_,
		_w1111_,
		_w1370_
	);
	LUT3 #(
		.INIT('h2a)
	) name1234 (
		\shift[6] ,
		_w1369_,
		_w1370_,
		_w1371_
	);
	LUT2 #(
		.INIT('he)
	) name1235 (
		_w1368_,
		_w1371_,
		_w1372_
	);
	LUT4 #(
		.INIT('hf7b3)
	) name1236 (
		\shift[4] ,
		\shift[5] ,
		_w180_,
		_w208_,
		_w1373_
	);
	LUT4 #(
		.INIT('hfdec)
	) name1237 (
		\shift[4] ,
		\shift[5] ,
		_w221_,
		_w248_,
		_w1374_
	);
	LUT3 #(
		.INIT('h15)
	) name1238 (
		\shift[6] ,
		_w1373_,
		_w1374_,
		_w1375_
	);
	LUT4 #(
		.INIT('hfbd9)
	) name1239 (
		\shift[4] ,
		\shift[5] ,
		_w153_,
		_w166_,
		_w1376_
	);
	LUT4 #(
		.INIT('hfe76)
	) name1240 (
		\shift[4] ,
		\shift[5] ,
		_w193_,
		_w235_,
		_w1377_
	);
	LUT3 #(
		.INIT('h2a)
	) name1241 (
		\shift[6] ,
		_w1376_,
		_w1377_,
		_w1378_
	);
	LUT2 #(
		.INIT('he)
	) name1242 (
		_w1375_,
		_w1378_,
		_w1379_
	);
	LUT4 #(
		.INIT('hf7b3)
	) name1243 (
		\shift[4] ,
		\shift[5] ,
		_w291_,
		_w332_,
		_w1380_
	);
	LUT4 #(
		.INIT('hfedc)
	) name1244 (
		\shift[4] ,
		\shift[5] ,
		_w346_,
		_w359_,
		_w1381_
	);
	LUT3 #(
		.INIT('h15)
	) name1245 (
		\shift[6] ,
		_w1380_,
		_w1381_,
		_w1382_
	);
	LUT4 #(
		.INIT('hfb73)
	) name1246 (
		\shift[4] ,
		\shift[5] ,
		_w264_,
		_w319_,
		_w1383_
	);
	LUT4 #(
		.INIT('hfdec)
	) name1247 (
		\shift[4] ,
		\shift[5] ,
		_w277_,
		_w304_,
		_w1384_
	);
	LUT3 #(
		.INIT('h2a)
	) name1248 (
		\shift[6] ,
		_w1383_,
		_w1384_,
		_w1385_
	);
	LUT2 #(
		.INIT('he)
	) name1249 (
		_w1382_,
		_w1385_,
		_w1386_
	);
	LUT4 #(
		.INIT('hf7b3)
	) name1250 (
		\shift[4] ,
		\shift[5] ,
		_w402_,
		_w443_,
		_w1387_
	);
	LUT4 #(
		.INIT('hfedc)
	) name1251 (
		\shift[4] ,
		\shift[5] ,
		_w457_,
		_w470_,
		_w1388_
	);
	LUT3 #(
		.INIT('h15)
	) name1252 (
		\shift[6] ,
		_w1387_,
		_w1388_,
		_w1389_
	);
	LUT4 #(
		.INIT('hfb73)
	) name1253 (
		\shift[4] ,
		\shift[5] ,
		_w375_,
		_w430_,
		_w1390_
	);
	LUT4 #(
		.INIT('hfdec)
	) name1254 (
		\shift[4] ,
		\shift[5] ,
		_w388_,
		_w415_,
		_w1391_
	);
	LUT3 #(
		.INIT('h2a)
	) name1255 (
		\shift[6] ,
		_w1390_,
		_w1391_,
		_w1392_
	);
	LUT2 #(
		.INIT('he)
	) name1256 (
		_w1389_,
		_w1392_,
		_w1393_
	);
	LUT4 #(
		.INIT('hfedc)
	) name1257 (
		\shift[4] ,
		\shift[5] ,
		_w554_,
		_w581_,
		_w1394_
	);
	LUT4 #(
		.INIT('hf7b3)
	) name1258 (
		\shift[4] ,
		\shift[5] ,
		_w513_,
		_w568_,
		_w1395_
	);
	LUT3 #(
		.INIT('h15)
	) name1259 (
		\shift[6] ,
		_w1394_,
		_w1395_,
		_w1396_
	);
	LUT4 #(
		.INIT('hfe76)
	) name1260 (
		\shift[4] ,
		\shift[5] ,
		_w486_,
		_w541_,
		_w1397_
	);
	LUT4 #(
		.INIT('hfdb9)
	) name1261 (
		\shift[4] ,
		\shift[5] ,
		_w499_,
		_w526_,
		_w1398_
	);
	LUT3 #(
		.INIT('h2a)
	) name1262 (
		\shift[6] ,
		_w1397_,
		_w1398_,
		_w1399_
	);
	LUT2 #(
		.INIT('he)
	) name1263 (
		_w1396_,
		_w1399_,
		_w1400_
	);
	LUT4 #(
		.INIT('hf7e6)
	) name1264 (
		\shift[4] ,
		\shift[5] ,
		_w600_,
		_w612_,
		_w1401_
	);
	LUT4 #(
		.INIT('hfdb9)
	) name1265 (
		\shift[4] ,
		\shift[5] ,
		_w623_,
		_w628_,
		_w1402_
	);
	LUT3 #(
		.INIT('h15)
	) name1266 (
		\shift[6] ,
		_w1401_,
		_w1402_,
		_w1403_
	);
	LUT4 #(
		.INIT('hfbd9)
	) name1267 (
		\shift[4] ,
		\shift[5] ,
		_w589_,
		_w594_,
		_w1404_
	);
	LUT4 #(
		.INIT('hfe76)
	) name1268 (
		\shift[4] ,
		\shift[5] ,
		_w605_,
		_w617_,
		_w1405_
	);
	LUT3 #(
		.INIT('h2a)
	) name1269 (
		\shift[6] ,
		_w1404_,
		_w1405_,
		_w1406_
	);
	LUT2 #(
		.INIT('he)
	) name1270 (
		_w1403_,
		_w1406_,
		_w1407_
	);
	LUT4 #(
		.INIT('hf7e6)
	) name1271 (
		\shift[4] ,
		\shift[5] ,
		_w647_,
		_w659_,
		_w1408_
	);
	LUT4 #(
		.INIT('hfdb9)
	) name1272 (
		\shift[4] ,
		\shift[5] ,
		_w670_,
		_w675_,
		_w1409_
	);
	LUT3 #(
		.INIT('h15)
	) name1273 (
		\shift[6] ,
		_w1408_,
		_w1409_,
		_w1410_
	);
	LUT4 #(
		.INIT('hfbd9)
	) name1274 (
		\shift[4] ,
		\shift[5] ,
		_w636_,
		_w641_,
		_w1411_
	);
	LUT4 #(
		.INIT('hfe76)
	) name1275 (
		\shift[4] ,
		\shift[5] ,
		_w652_,
		_w664_,
		_w1412_
	);
	LUT3 #(
		.INIT('h2a)
	) name1276 (
		\shift[6] ,
		_w1411_,
		_w1412_,
		_w1413_
	);
	LUT2 #(
		.INIT('he)
	) name1277 (
		_w1410_,
		_w1413_,
		_w1414_
	);
	LUT4 #(
		.INIT('hf7e6)
	) name1278 (
		\shift[4] ,
		\shift[5] ,
		_w694_,
		_w706_,
		_w1415_
	);
	LUT4 #(
		.INIT('hfdb9)
	) name1279 (
		\shift[4] ,
		\shift[5] ,
		_w717_,
		_w722_,
		_w1416_
	);
	LUT3 #(
		.INIT('h15)
	) name1280 (
		\shift[6] ,
		_w1415_,
		_w1416_,
		_w1417_
	);
	LUT4 #(
		.INIT('hfbd9)
	) name1281 (
		\shift[4] ,
		\shift[5] ,
		_w683_,
		_w688_,
		_w1418_
	);
	LUT4 #(
		.INIT('hfe76)
	) name1282 (
		\shift[4] ,
		\shift[5] ,
		_w699_,
		_w711_,
		_w1419_
	);
	LUT3 #(
		.INIT('h2a)
	) name1283 (
		\shift[6] ,
		_w1418_,
		_w1419_,
		_w1420_
	);
	LUT2 #(
		.INIT('he)
	) name1284 (
		_w1417_,
		_w1420_,
		_w1421_
	);
	LUT4 #(
		.INIT('hfeba)
	) name1285 (
		\shift[4] ,
		\shift[5] ,
		_w753_,
		_w769_,
		_w1422_
	);
	LUT4 #(
		.INIT('hf7d5)
	) name1286 (
		\shift[4] ,
		\shift[5] ,
		_w741_,
		_w764_,
		_w1423_
	);
	LUT3 #(
		.INIT('h15)
	) name1287 (
		\shift[6] ,
		_w1422_,
		_w1423_,
		_w1424_
	);
	LUT4 #(
		.INIT('hfb73)
	) name1288 (
		\shift[4] ,
		\shift[5] ,
		_w730_,
		_w758_,
		_w1425_
	);
	LUT4 #(
		.INIT('hfdec)
	) name1289 (
		\shift[4] ,
		\shift[5] ,
		_w735_,
		_w746_,
		_w1426_
	);
	LUT3 #(
		.INIT('h2a)
	) name1290 (
		\shift[6] ,
		_w1425_,
		_w1426_,
		_w1427_
	);
	LUT2 #(
		.INIT('he)
	) name1291 (
		_w1424_,
		_w1427_,
		_w1428_
	);
	LUT4 #(
		.INIT('hfeba)
	) name1292 (
		\shift[4] ,
		\shift[5] ,
		_w800_,
		_w816_,
		_w1429_
	);
	LUT4 #(
		.INIT('hf7d5)
	) name1293 (
		\shift[4] ,
		\shift[5] ,
		_w788_,
		_w811_,
		_w1430_
	);
	LUT3 #(
		.INIT('h15)
	) name1294 (
		\shift[6] ,
		_w1429_,
		_w1430_,
		_w1431_
	);
	LUT4 #(
		.INIT('hfb73)
	) name1295 (
		\shift[4] ,
		\shift[5] ,
		_w777_,
		_w805_,
		_w1432_
	);
	LUT4 #(
		.INIT('hfdec)
	) name1296 (
		\shift[4] ,
		\shift[5] ,
		_w782_,
		_w793_,
		_w1433_
	);
	LUT3 #(
		.INIT('h2a)
	) name1297 (
		\shift[6] ,
		_w1432_,
		_w1433_,
		_w1434_
	);
	LUT2 #(
		.INIT('he)
	) name1298 (
		_w1431_,
		_w1434_,
		_w1435_
	);
	LUT4 #(
		.INIT('hfeba)
	) name1299 (
		\shift[4] ,
		\shift[5] ,
		_w847_,
		_w863_,
		_w1436_
	);
	LUT4 #(
		.INIT('hf7d5)
	) name1300 (
		\shift[4] ,
		\shift[5] ,
		_w835_,
		_w858_,
		_w1437_
	);
	LUT3 #(
		.INIT('h15)
	) name1301 (
		\shift[6] ,
		_w1436_,
		_w1437_,
		_w1438_
	);
	LUT4 #(
		.INIT('hfb73)
	) name1302 (
		\shift[4] ,
		\shift[5] ,
		_w824_,
		_w852_,
		_w1439_
	);
	LUT4 #(
		.INIT('hfdec)
	) name1303 (
		\shift[4] ,
		\shift[5] ,
		_w829_,
		_w840_,
		_w1440_
	);
	LUT3 #(
		.INIT('h2a)
	) name1304 (
		\shift[6] ,
		_w1439_,
		_w1440_,
		_w1441_
	);
	LUT2 #(
		.INIT('he)
	) name1305 (
		_w1438_,
		_w1441_,
		_w1442_
	);
	LUT4 #(
		.INIT('hf7e6)
	) name1306 (
		\shift[4] ,
		\shift[5] ,
		_w882_,
		_w894_,
		_w1443_
	);
	LUT4 #(
		.INIT('hfdb9)
	) name1307 (
		\shift[4] ,
		\shift[5] ,
		_w905_,
		_w910_,
		_w1444_
	);
	LUT3 #(
		.INIT('h15)
	) name1308 (
		\shift[6] ,
		_w1443_,
		_w1444_,
		_w1445_
	);
	LUT4 #(
		.INIT('hfb73)
	) name1309 (
		\shift[4] ,
		\shift[5] ,
		_w871_,
		_w899_,
		_w1446_
	);
	LUT4 #(
		.INIT('hfdec)
	) name1310 (
		\shift[4] ,
		\shift[5] ,
		_w876_,
		_w887_,
		_w1447_
	);
	LUT3 #(
		.INIT('h2a)
	) name1311 (
		\shift[6] ,
		_w1446_,
		_w1447_,
		_w1448_
	);
	LUT2 #(
		.INIT('he)
	) name1312 (
		_w1445_,
		_w1448_,
		_w1449_
	);
	LUT4 #(
		.INIT('hf7e6)
	) name1313 (
		\shift[4] ,
		\shift[5] ,
		_w929_,
		_w941_,
		_w1450_
	);
	LUT4 #(
		.INIT('hfdb9)
	) name1314 (
		\shift[4] ,
		\shift[5] ,
		_w952_,
		_w957_,
		_w1451_
	);
	LUT3 #(
		.INIT('h15)
	) name1315 (
		\shift[6] ,
		_w1450_,
		_w1451_,
		_w1452_
	);
	LUT4 #(
		.INIT('hfb73)
	) name1316 (
		\shift[4] ,
		\shift[5] ,
		_w918_,
		_w946_,
		_w1453_
	);
	LUT4 #(
		.INIT('hfdec)
	) name1317 (
		\shift[4] ,
		\shift[5] ,
		_w923_,
		_w934_,
		_w1454_
	);
	LUT3 #(
		.INIT('h2a)
	) name1318 (
		\shift[6] ,
		_w1453_,
		_w1454_,
		_w1455_
	);
	LUT2 #(
		.INIT('he)
	) name1319 (
		_w1452_,
		_w1455_,
		_w1456_
	);
	LUT4 #(
		.INIT('hf7e6)
	) name1320 (
		\shift[4] ,
		\shift[5] ,
		_w976_,
		_w988_,
		_w1457_
	);
	LUT4 #(
		.INIT('hfdb9)
	) name1321 (
		\shift[4] ,
		\shift[5] ,
		_w999_,
		_w1004_,
		_w1458_
	);
	LUT3 #(
		.INIT('h15)
	) name1322 (
		\shift[6] ,
		_w1457_,
		_w1458_,
		_w1459_
	);
	LUT4 #(
		.INIT('hfb73)
	) name1323 (
		\shift[4] ,
		\shift[5] ,
		_w965_,
		_w993_,
		_w1460_
	);
	LUT4 #(
		.INIT('hfdec)
	) name1324 (
		\shift[4] ,
		\shift[5] ,
		_w970_,
		_w981_,
		_w1461_
	);
	LUT3 #(
		.INIT('h2a)
	) name1325 (
		\shift[6] ,
		_w1460_,
		_w1461_,
		_w1462_
	);
	LUT2 #(
		.INIT('he)
	) name1326 (
		_w1459_,
		_w1462_,
		_w1463_
	);
	LUT4 #(
		.INIT('hf7e6)
	) name1327 (
		\shift[4] ,
		\shift[5] ,
		_w1023_,
		_w1035_,
		_w1464_
	);
	LUT4 #(
		.INIT('hfdb9)
	) name1328 (
		\shift[4] ,
		\shift[5] ,
		_w1046_,
		_w1051_,
		_w1465_
	);
	LUT3 #(
		.INIT('h15)
	) name1329 (
		\shift[6] ,
		_w1464_,
		_w1465_,
		_w1466_
	);
	LUT4 #(
		.INIT('hfb73)
	) name1330 (
		\shift[4] ,
		\shift[5] ,
		_w1012_,
		_w1040_,
		_w1467_
	);
	LUT4 #(
		.INIT('hfdec)
	) name1331 (
		\shift[4] ,
		\shift[5] ,
		_w1017_,
		_w1028_,
		_w1468_
	);
	LUT3 #(
		.INIT('h2a)
	) name1332 (
		\shift[6] ,
		_w1467_,
		_w1468_,
		_w1469_
	);
	LUT2 #(
		.INIT('he)
	) name1333 (
		_w1466_,
		_w1469_,
		_w1470_
	);
	LUT4 #(
		.INIT('hf7e6)
	) name1334 (
		\shift[4] ,
		\shift[5] ,
		_w1070_,
		_w1082_,
		_w1471_
	);
	LUT4 #(
		.INIT('hfdb9)
	) name1335 (
		\shift[4] ,
		\shift[5] ,
		_w1093_,
		_w1098_,
		_w1472_
	);
	LUT3 #(
		.INIT('h15)
	) name1336 (
		\shift[6] ,
		_w1471_,
		_w1472_,
		_w1473_
	);
	LUT4 #(
		.INIT('hfb73)
	) name1337 (
		\shift[4] ,
		\shift[5] ,
		_w1059_,
		_w1087_,
		_w1474_
	);
	LUT4 #(
		.INIT('hfdec)
	) name1338 (
		\shift[4] ,
		\shift[5] ,
		_w1064_,
		_w1075_,
		_w1475_
	);
	LUT3 #(
		.INIT('h2a)
	) name1339 (
		\shift[6] ,
		_w1474_,
		_w1475_,
		_w1476_
	);
	LUT2 #(
		.INIT('he)
	) name1340 (
		_w1473_,
		_w1476_,
		_w1477_
	);
	LUT4 #(
		.INIT('hf7e6)
	) name1341 (
		\shift[4] ,
		\shift[5] ,
		_w1117_,
		_w1129_,
		_w1478_
	);
	LUT4 #(
		.INIT('hfdb9)
	) name1342 (
		\shift[4] ,
		\shift[5] ,
		_w1140_,
		_w1145_,
		_w1479_
	);
	LUT3 #(
		.INIT('h15)
	) name1343 (
		\shift[6] ,
		_w1478_,
		_w1479_,
		_w1480_
	);
	LUT4 #(
		.INIT('hfb73)
	) name1344 (
		\shift[4] ,
		\shift[5] ,
		_w1106_,
		_w1134_,
		_w1481_
	);
	LUT4 #(
		.INIT('hfdec)
	) name1345 (
		\shift[4] ,
		\shift[5] ,
		_w1111_,
		_w1122_,
		_w1482_
	);
	LUT3 #(
		.INIT('h2a)
	) name1346 (
		\shift[6] ,
		_w1481_,
		_w1482_,
		_w1483_
	);
	LUT2 #(
		.INIT('he)
	) name1347 (
		_w1480_,
		_w1483_,
		_w1484_
	);
	LUT3 #(
		.INIT('h15)
	) name1348 (
		\shift[6] ,
		_w222_,
		_w249_,
		_w1485_
	);
	LUT3 #(
		.INIT('h2a)
	) name1349 (
		\shift[6] ,
		_w167_,
		_w194_,
		_w1486_
	);
	LUT2 #(
		.INIT('he)
	) name1350 (
		_w1485_,
		_w1486_,
		_w1487_
	);
	LUT3 #(
		.INIT('h15)
	) name1351 (
		\shift[6] ,
		_w333_,
		_w360_,
		_w1488_
	);
	LUT3 #(
		.INIT('h2a)
	) name1352 (
		\shift[6] ,
		_w278_,
		_w305_,
		_w1489_
	);
	LUT2 #(
		.INIT('he)
	) name1353 (
		_w1488_,
		_w1489_,
		_w1490_
	);
	LUT3 #(
		.INIT('h15)
	) name1354 (
		\shift[6] ,
		_w444_,
		_w471_,
		_w1491_
	);
	LUT3 #(
		.INIT('h2a)
	) name1355 (
		\shift[6] ,
		_w389_,
		_w416_,
		_w1492_
	);
	LUT2 #(
		.INIT('he)
	) name1356 (
		_w1491_,
		_w1492_,
		_w1493_
	);
	LUT3 #(
		.INIT('h15)
	) name1357 (
		\shift[6] ,
		_w555_,
		_w582_,
		_w1494_
	);
	LUT3 #(
		.INIT('h2a)
	) name1358 (
		\shift[6] ,
		_w500_,
		_w527_,
		_w1495_
	);
	LUT2 #(
		.INIT('he)
	) name1359 (
		_w1494_,
		_w1495_,
		_w1496_
	);
	LUT3 #(
		.INIT('h15)
	) name1360 (
		\shift[6] ,
		_w618_,
		_w629_,
		_w1497_
	);
	LUT3 #(
		.INIT('h2a)
	) name1361 (
		\shift[6] ,
		_w595_,
		_w606_,
		_w1498_
	);
	LUT2 #(
		.INIT('he)
	) name1362 (
		_w1497_,
		_w1498_,
		_w1499_
	);
	LUT3 #(
		.INIT('h15)
	) name1363 (
		\shift[6] ,
		_w665_,
		_w676_,
		_w1500_
	);
	LUT3 #(
		.INIT('h2a)
	) name1364 (
		\shift[6] ,
		_w642_,
		_w653_,
		_w1501_
	);
	LUT2 #(
		.INIT('he)
	) name1365 (
		_w1500_,
		_w1501_,
		_w1502_
	);
	LUT3 #(
		.INIT('h15)
	) name1366 (
		\shift[6] ,
		_w712_,
		_w723_,
		_w1503_
	);
	LUT3 #(
		.INIT('h2a)
	) name1367 (
		\shift[6] ,
		_w689_,
		_w700_,
		_w1504_
	);
	LUT2 #(
		.INIT('he)
	) name1368 (
		_w1503_,
		_w1504_,
		_w1505_
	);
	LUT3 #(
		.INIT('h15)
	) name1369 (
		\shift[6] ,
		_w759_,
		_w770_,
		_w1506_
	);
	LUT3 #(
		.INIT('h2a)
	) name1370 (
		\shift[6] ,
		_w736_,
		_w747_,
		_w1507_
	);
	LUT2 #(
		.INIT('he)
	) name1371 (
		_w1506_,
		_w1507_,
		_w1508_
	);
	LUT3 #(
		.INIT('h15)
	) name1372 (
		\shift[6] ,
		_w806_,
		_w817_,
		_w1509_
	);
	LUT3 #(
		.INIT('h2a)
	) name1373 (
		\shift[6] ,
		_w783_,
		_w794_,
		_w1510_
	);
	LUT2 #(
		.INIT('he)
	) name1374 (
		_w1509_,
		_w1510_,
		_w1511_
	);
	LUT3 #(
		.INIT('h15)
	) name1375 (
		\shift[6] ,
		_w853_,
		_w864_,
		_w1512_
	);
	LUT3 #(
		.INIT('h2a)
	) name1376 (
		\shift[6] ,
		_w830_,
		_w841_,
		_w1513_
	);
	LUT2 #(
		.INIT('he)
	) name1377 (
		_w1512_,
		_w1513_,
		_w1514_
	);
	LUT3 #(
		.INIT('h15)
	) name1378 (
		\shift[6] ,
		_w900_,
		_w911_,
		_w1515_
	);
	LUT3 #(
		.INIT('h2a)
	) name1379 (
		\shift[6] ,
		_w877_,
		_w888_,
		_w1516_
	);
	LUT2 #(
		.INIT('he)
	) name1380 (
		_w1515_,
		_w1516_,
		_w1517_
	);
	LUT3 #(
		.INIT('h15)
	) name1381 (
		\shift[6] ,
		_w947_,
		_w958_,
		_w1518_
	);
	LUT3 #(
		.INIT('h2a)
	) name1382 (
		\shift[6] ,
		_w924_,
		_w935_,
		_w1519_
	);
	LUT2 #(
		.INIT('he)
	) name1383 (
		_w1518_,
		_w1519_,
		_w1520_
	);
	LUT3 #(
		.INIT('h15)
	) name1384 (
		\shift[6] ,
		_w994_,
		_w1005_,
		_w1521_
	);
	LUT3 #(
		.INIT('h2a)
	) name1385 (
		\shift[6] ,
		_w971_,
		_w982_,
		_w1522_
	);
	LUT2 #(
		.INIT('he)
	) name1386 (
		_w1521_,
		_w1522_,
		_w1523_
	);
	LUT3 #(
		.INIT('h15)
	) name1387 (
		\shift[6] ,
		_w1041_,
		_w1052_,
		_w1524_
	);
	LUT3 #(
		.INIT('h2a)
	) name1388 (
		\shift[6] ,
		_w1018_,
		_w1029_,
		_w1525_
	);
	LUT2 #(
		.INIT('he)
	) name1389 (
		_w1524_,
		_w1525_,
		_w1526_
	);
	LUT3 #(
		.INIT('h15)
	) name1390 (
		\shift[6] ,
		_w1088_,
		_w1099_,
		_w1527_
	);
	LUT3 #(
		.INIT('h2a)
	) name1391 (
		\shift[6] ,
		_w1065_,
		_w1076_,
		_w1528_
	);
	LUT2 #(
		.INIT('he)
	) name1392 (
		_w1527_,
		_w1528_,
		_w1529_
	);
	LUT3 #(
		.INIT('h15)
	) name1393 (
		\shift[6] ,
		_w1135_,
		_w1146_,
		_w1530_
	);
	LUT3 #(
		.INIT('h2a)
	) name1394 (
		\shift[6] ,
		_w1112_,
		_w1123_,
		_w1531_
	);
	LUT2 #(
		.INIT('he)
	) name1395 (
		_w1530_,
		_w1531_,
		_w1532_
	);
	LUT3 #(
		.INIT('h15)
	) name1396 (
		\shift[6] ,
		_w1152_,
		_w1153_,
		_w1533_
	);
	LUT3 #(
		.INIT('h2a)
	) name1397 (
		\shift[6] ,
		_w1149_,
		_w1150_,
		_w1534_
	);
	LUT2 #(
		.INIT('he)
	) name1398 (
		_w1533_,
		_w1534_,
		_w1535_
	);
	LUT3 #(
		.INIT('h15)
	) name1399 (
		\shift[6] ,
		_w1159_,
		_w1160_,
		_w1536_
	);
	LUT3 #(
		.INIT('h2a)
	) name1400 (
		\shift[6] ,
		_w1156_,
		_w1157_,
		_w1537_
	);
	LUT2 #(
		.INIT('he)
	) name1401 (
		_w1536_,
		_w1537_,
		_w1538_
	);
	LUT3 #(
		.INIT('h15)
	) name1402 (
		\shift[6] ,
		_w1166_,
		_w1167_,
		_w1539_
	);
	LUT3 #(
		.INIT('h2a)
	) name1403 (
		\shift[6] ,
		_w1163_,
		_w1164_,
		_w1540_
	);
	LUT2 #(
		.INIT('he)
	) name1404 (
		_w1539_,
		_w1540_,
		_w1541_
	);
	LUT3 #(
		.INIT('h15)
	) name1405 (
		\shift[6] ,
		_w1173_,
		_w1174_,
		_w1542_
	);
	LUT3 #(
		.INIT('h2a)
	) name1406 (
		\shift[6] ,
		_w1170_,
		_w1171_,
		_w1543_
	);
	LUT2 #(
		.INIT('he)
	) name1407 (
		_w1542_,
		_w1543_,
		_w1544_
	);
	LUT3 #(
		.INIT('h15)
	) name1408 (
		\shift[6] ,
		_w1180_,
		_w1181_,
		_w1545_
	);
	LUT3 #(
		.INIT('h2a)
	) name1409 (
		\shift[6] ,
		_w1177_,
		_w1178_,
		_w1546_
	);
	LUT2 #(
		.INIT('he)
	) name1410 (
		_w1545_,
		_w1546_,
		_w1547_
	);
	LUT3 #(
		.INIT('h15)
	) name1411 (
		\shift[6] ,
		_w1187_,
		_w1188_,
		_w1548_
	);
	LUT3 #(
		.INIT('h2a)
	) name1412 (
		\shift[6] ,
		_w1184_,
		_w1185_,
		_w1549_
	);
	LUT2 #(
		.INIT('he)
	) name1413 (
		_w1548_,
		_w1549_,
		_w1550_
	);
	LUT3 #(
		.INIT('h15)
	) name1414 (
		\shift[6] ,
		_w1194_,
		_w1195_,
		_w1551_
	);
	LUT3 #(
		.INIT('h2a)
	) name1415 (
		\shift[6] ,
		_w1191_,
		_w1192_,
		_w1552_
	);
	LUT2 #(
		.INIT('he)
	) name1416 (
		_w1551_,
		_w1552_,
		_w1553_
	);
	LUT3 #(
		.INIT('h15)
	) name1417 (
		\shift[6] ,
		_w1201_,
		_w1202_,
		_w1554_
	);
	LUT3 #(
		.INIT('h2a)
	) name1418 (
		\shift[6] ,
		_w1198_,
		_w1199_,
		_w1555_
	);
	LUT2 #(
		.INIT('he)
	) name1419 (
		_w1554_,
		_w1555_,
		_w1556_
	);
	LUT3 #(
		.INIT('h15)
	) name1420 (
		\shift[6] ,
		_w1208_,
		_w1209_,
		_w1557_
	);
	LUT3 #(
		.INIT('h2a)
	) name1421 (
		\shift[6] ,
		_w1205_,
		_w1206_,
		_w1558_
	);
	LUT2 #(
		.INIT('he)
	) name1422 (
		_w1557_,
		_w1558_,
		_w1559_
	);
	LUT3 #(
		.INIT('h15)
	) name1423 (
		\shift[6] ,
		_w1215_,
		_w1216_,
		_w1560_
	);
	LUT3 #(
		.INIT('h2a)
	) name1424 (
		\shift[6] ,
		_w1212_,
		_w1213_,
		_w1561_
	);
	LUT2 #(
		.INIT('he)
	) name1425 (
		_w1560_,
		_w1561_,
		_w1562_
	);
	LUT3 #(
		.INIT('h15)
	) name1426 (
		\shift[6] ,
		_w1222_,
		_w1223_,
		_w1563_
	);
	LUT3 #(
		.INIT('h2a)
	) name1427 (
		\shift[6] ,
		_w1219_,
		_w1220_,
		_w1564_
	);
	LUT2 #(
		.INIT('he)
	) name1428 (
		_w1563_,
		_w1564_,
		_w1565_
	);
	LUT3 #(
		.INIT('h15)
	) name1429 (
		\shift[6] ,
		_w1229_,
		_w1230_,
		_w1566_
	);
	LUT3 #(
		.INIT('h2a)
	) name1430 (
		\shift[6] ,
		_w1226_,
		_w1227_,
		_w1567_
	);
	LUT2 #(
		.INIT('he)
	) name1431 (
		_w1566_,
		_w1567_,
		_w1568_
	);
	LUT3 #(
		.INIT('h15)
	) name1432 (
		\shift[6] ,
		_w1236_,
		_w1237_,
		_w1569_
	);
	LUT3 #(
		.INIT('h2a)
	) name1433 (
		\shift[6] ,
		_w1233_,
		_w1234_,
		_w1570_
	);
	LUT2 #(
		.INIT('he)
	) name1434 (
		_w1569_,
		_w1570_,
		_w1571_
	);
	LUT3 #(
		.INIT('h15)
	) name1435 (
		\shift[6] ,
		_w1243_,
		_w1244_,
		_w1572_
	);
	LUT3 #(
		.INIT('h2a)
	) name1436 (
		\shift[6] ,
		_w1240_,
		_w1241_,
		_w1573_
	);
	LUT2 #(
		.INIT('he)
	) name1437 (
		_w1572_,
		_w1573_,
		_w1574_
	);
	LUT3 #(
		.INIT('h15)
	) name1438 (
		\shift[6] ,
		_w1250_,
		_w1251_,
		_w1575_
	);
	LUT3 #(
		.INIT('h2a)
	) name1439 (
		\shift[6] ,
		_w1247_,
		_w1248_,
		_w1576_
	);
	LUT2 #(
		.INIT('he)
	) name1440 (
		_w1575_,
		_w1576_,
		_w1577_
	);
	LUT3 #(
		.INIT('h15)
	) name1441 (
		\shift[6] ,
		_w1257_,
		_w1258_,
		_w1578_
	);
	LUT3 #(
		.INIT('h2a)
	) name1442 (
		\shift[6] ,
		_w1254_,
		_w1255_,
		_w1579_
	);
	LUT2 #(
		.INIT('he)
	) name1443 (
		_w1578_,
		_w1579_,
		_w1580_
	);
	LUT3 #(
		.INIT('h15)
	) name1444 (
		\shift[6] ,
		_w1264_,
		_w1265_,
		_w1581_
	);
	LUT3 #(
		.INIT('h2a)
	) name1445 (
		\shift[6] ,
		_w1261_,
		_w1262_,
		_w1582_
	);
	LUT2 #(
		.INIT('he)
	) name1446 (
		_w1581_,
		_w1582_,
		_w1583_
	);
	LUT3 #(
		.INIT('h15)
	) name1447 (
		\shift[6] ,
		_w1271_,
		_w1272_,
		_w1584_
	);
	LUT3 #(
		.INIT('h2a)
	) name1448 (
		\shift[6] ,
		_w1268_,
		_w1269_,
		_w1585_
	);
	LUT2 #(
		.INIT('he)
	) name1449 (
		_w1584_,
		_w1585_,
		_w1586_
	);
	LUT3 #(
		.INIT('h15)
	) name1450 (
		\shift[6] ,
		_w1278_,
		_w1279_,
		_w1587_
	);
	LUT3 #(
		.INIT('h2a)
	) name1451 (
		\shift[6] ,
		_w1275_,
		_w1276_,
		_w1588_
	);
	LUT2 #(
		.INIT('he)
	) name1452 (
		_w1587_,
		_w1588_,
		_w1589_
	);
	LUT3 #(
		.INIT('h15)
	) name1453 (
		\shift[6] ,
		_w1285_,
		_w1286_,
		_w1590_
	);
	LUT3 #(
		.INIT('h2a)
	) name1454 (
		\shift[6] ,
		_w1282_,
		_w1283_,
		_w1591_
	);
	LUT2 #(
		.INIT('he)
	) name1455 (
		_w1590_,
		_w1591_,
		_w1592_
	);
	LUT3 #(
		.INIT('h15)
	) name1456 (
		\shift[6] ,
		_w1292_,
		_w1293_,
		_w1593_
	);
	LUT3 #(
		.INIT('h2a)
	) name1457 (
		\shift[6] ,
		_w1289_,
		_w1290_,
		_w1594_
	);
	LUT2 #(
		.INIT('he)
	) name1458 (
		_w1593_,
		_w1594_,
		_w1595_
	);
	LUT3 #(
		.INIT('h15)
	) name1459 (
		\shift[6] ,
		_w1299_,
		_w1300_,
		_w1596_
	);
	LUT3 #(
		.INIT('h2a)
	) name1460 (
		\shift[6] ,
		_w1296_,
		_w1297_,
		_w1597_
	);
	LUT2 #(
		.INIT('he)
	) name1461 (
		_w1596_,
		_w1597_,
		_w1598_
	);
	LUT3 #(
		.INIT('h15)
	) name1462 (
		\shift[6] ,
		_w1306_,
		_w1307_,
		_w1599_
	);
	LUT3 #(
		.INIT('h2a)
	) name1463 (
		\shift[6] ,
		_w1303_,
		_w1304_,
		_w1600_
	);
	LUT2 #(
		.INIT('he)
	) name1464 (
		_w1599_,
		_w1600_,
		_w1601_
	);
	LUT3 #(
		.INIT('h15)
	) name1465 (
		\shift[6] ,
		_w1313_,
		_w1314_,
		_w1602_
	);
	LUT3 #(
		.INIT('h2a)
	) name1466 (
		\shift[6] ,
		_w1310_,
		_w1311_,
		_w1603_
	);
	LUT2 #(
		.INIT('he)
	) name1467 (
		_w1602_,
		_w1603_,
		_w1604_
	);
	LUT3 #(
		.INIT('h15)
	) name1468 (
		\shift[6] ,
		_w1320_,
		_w1321_,
		_w1605_
	);
	LUT3 #(
		.INIT('h2a)
	) name1469 (
		\shift[6] ,
		_w1317_,
		_w1318_,
		_w1606_
	);
	LUT2 #(
		.INIT('he)
	) name1470 (
		_w1605_,
		_w1606_,
		_w1607_
	);
	LUT3 #(
		.INIT('h15)
	) name1471 (
		\shift[6] ,
		_w1327_,
		_w1328_,
		_w1608_
	);
	LUT3 #(
		.INIT('h2a)
	) name1472 (
		\shift[6] ,
		_w1324_,
		_w1325_,
		_w1609_
	);
	LUT2 #(
		.INIT('he)
	) name1473 (
		_w1608_,
		_w1609_,
		_w1610_
	);
	LUT3 #(
		.INIT('h15)
	) name1474 (
		\shift[6] ,
		_w1334_,
		_w1335_,
		_w1611_
	);
	LUT3 #(
		.INIT('h2a)
	) name1475 (
		\shift[6] ,
		_w1331_,
		_w1332_,
		_w1612_
	);
	LUT2 #(
		.INIT('he)
	) name1476 (
		_w1611_,
		_w1612_,
		_w1613_
	);
	LUT3 #(
		.INIT('h15)
	) name1477 (
		\shift[6] ,
		_w1341_,
		_w1342_,
		_w1614_
	);
	LUT3 #(
		.INIT('h2a)
	) name1478 (
		\shift[6] ,
		_w1338_,
		_w1339_,
		_w1615_
	);
	LUT2 #(
		.INIT('he)
	) name1479 (
		_w1614_,
		_w1615_,
		_w1616_
	);
	LUT3 #(
		.INIT('h15)
	) name1480 (
		\shift[6] ,
		_w1348_,
		_w1349_,
		_w1617_
	);
	LUT3 #(
		.INIT('h2a)
	) name1481 (
		\shift[6] ,
		_w1345_,
		_w1346_,
		_w1618_
	);
	LUT2 #(
		.INIT('he)
	) name1482 (
		_w1617_,
		_w1618_,
		_w1619_
	);
	LUT3 #(
		.INIT('h15)
	) name1483 (
		\shift[6] ,
		_w1355_,
		_w1356_,
		_w1620_
	);
	LUT3 #(
		.INIT('h2a)
	) name1484 (
		\shift[6] ,
		_w1352_,
		_w1353_,
		_w1621_
	);
	LUT2 #(
		.INIT('he)
	) name1485 (
		_w1620_,
		_w1621_,
		_w1622_
	);
	LUT3 #(
		.INIT('h15)
	) name1486 (
		\shift[6] ,
		_w1362_,
		_w1363_,
		_w1623_
	);
	LUT3 #(
		.INIT('h2a)
	) name1487 (
		\shift[6] ,
		_w1359_,
		_w1360_,
		_w1624_
	);
	LUT2 #(
		.INIT('he)
	) name1488 (
		_w1623_,
		_w1624_,
		_w1625_
	);
	LUT3 #(
		.INIT('h15)
	) name1489 (
		\shift[6] ,
		_w1369_,
		_w1370_,
		_w1626_
	);
	LUT3 #(
		.INIT('h2a)
	) name1490 (
		\shift[6] ,
		_w1366_,
		_w1367_,
		_w1627_
	);
	LUT2 #(
		.INIT('he)
	) name1491 (
		_w1626_,
		_w1627_,
		_w1628_
	);
	LUT3 #(
		.INIT('h15)
	) name1492 (
		\shift[6] ,
		_w1376_,
		_w1377_,
		_w1629_
	);
	LUT3 #(
		.INIT('h2a)
	) name1493 (
		\shift[6] ,
		_w1373_,
		_w1374_,
		_w1630_
	);
	LUT2 #(
		.INIT('he)
	) name1494 (
		_w1629_,
		_w1630_,
		_w1631_
	);
	LUT3 #(
		.INIT('h15)
	) name1495 (
		\shift[6] ,
		_w1383_,
		_w1384_,
		_w1632_
	);
	LUT3 #(
		.INIT('h2a)
	) name1496 (
		\shift[6] ,
		_w1380_,
		_w1381_,
		_w1633_
	);
	LUT2 #(
		.INIT('he)
	) name1497 (
		_w1632_,
		_w1633_,
		_w1634_
	);
	LUT3 #(
		.INIT('h15)
	) name1498 (
		\shift[6] ,
		_w1390_,
		_w1391_,
		_w1635_
	);
	LUT3 #(
		.INIT('h2a)
	) name1499 (
		\shift[6] ,
		_w1387_,
		_w1388_,
		_w1636_
	);
	LUT2 #(
		.INIT('he)
	) name1500 (
		_w1635_,
		_w1636_,
		_w1637_
	);
	LUT3 #(
		.INIT('h15)
	) name1501 (
		\shift[6] ,
		_w1397_,
		_w1398_,
		_w1638_
	);
	LUT3 #(
		.INIT('h2a)
	) name1502 (
		\shift[6] ,
		_w1394_,
		_w1395_,
		_w1639_
	);
	LUT2 #(
		.INIT('he)
	) name1503 (
		_w1638_,
		_w1639_,
		_w1640_
	);
	LUT3 #(
		.INIT('h15)
	) name1504 (
		\shift[6] ,
		_w1404_,
		_w1405_,
		_w1641_
	);
	LUT3 #(
		.INIT('h2a)
	) name1505 (
		\shift[6] ,
		_w1401_,
		_w1402_,
		_w1642_
	);
	LUT2 #(
		.INIT('he)
	) name1506 (
		_w1641_,
		_w1642_,
		_w1643_
	);
	LUT3 #(
		.INIT('h15)
	) name1507 (
		\shift[6] ,
		_w1411_,
		_w1412_,
		_w1644_
	);
	LUT3 #(
		.INIT('h2a)
	) name1508 (
		\shift[6] ,
		_w1408_,
		_w1409_,
		_w1645_
	);
	LUT2 #(
		.INIT('he)
	) name1509 (
		_w1644_,
		_w1645_,
		_w1646_
	);
	LUT3 #(
		.INIT('h15)
	) name1510 (
		\shift[6] ,
		_w1418_,
		_w1419_,
		_w1647_
	);
	LUT3 #(
		.INIT('h2a)
	) name1511 (
		\shift[6] ,
		_w1415_,
		_w1416_,
		_w1648_
	);
	LUT2 #(
		.INIT('he)
	) name1512 (
		_w1647_,
		_w1648_,
		_w1649_
	);
	LUT3 #(
		.INIT('h15)
	) name1513 (
		\shift[6] ,
		_w1425_,
		_w1426_,
		_w1650_
	);
	LUT3 #(
		.INIT('h2a)
	) name1514 (
		\shift[6] ,
		_w1422_,
		_w1423_,
		_w1651_
	);
	LUT2 #(
		.INIT('he)
	) name1515 (
		_w1650_,
		_w1651_,
		_w1652_
	);
	LUT3 #(
		.INIT('h15)
	) name1516 (
		\shift[6] ,
		_w1432_,
		_w1433_,
		_w1653_
	);
	LUT3 #(
		.INIT('h2a)
	) name1517 (
		\shift[6] ,
		_w1429_,
		_w1430_,
		_w1654_
	);
	LUT2 #(
		.INIT('he)
	) name1518 (
		_w1653_,
		_w1654_,
		_w1655_
	);
	LUT3 #(
		.INIT('h15)
	) name1519 (
		\shift[6] ,
		_w1439_,
		_w1440_,
		_w1656_
	);
	LUT3 #(
		.INIT('h2a)
	) name1520 (
		\shift[6] ,
		_w1436_,
		_w1437_,
		_w1657_
	);
	LUT2 #(
		.INIT('he)
	) name1521 (
		_w1656_,
		_w1657_,
		_w1658_
	);
	LUT3 #(
		.INIT('h15)
	) name1522 (
		\shift[6] ,
		_w1446_,
		_w1447_,
		_w1659_
	);
	LUT3 #(
		.INIT('h2a)
	) name1523 (
		\shift[6] ,
		_w1443_,
		_w1444_,
		_w1660_
	);
	LUT2 #(
		.INIT('he)
	) name1524 (
		_w1659_,
		_w1660_,
		_w1661_
	);
	LUT3 #(
		.INIT('h15)
	) name1525 (
		\shift[6] ,
		_w1453_,
		_w1454_,
		_w1662_
	);
	LUT3 #(
		.INIT('h2a)
	) name1526 (
		\shift[6] ,
		_w1450_,
		_w1451_,
		_w1663_
	);
	LUT2 #(
		.INIT('he)
	) name1527 (
		_w1662_,
		_w1663_,
		_w1664_
	);
	LUT3 #(
		.INIT('h15)
	) name1528 (
		\shift[6] ,
		_w1460_,
		_w1461_,
		_w1665_
	);
	LUT3 #(
		.INIT('h2a)
	) name1529 (
		\shift[6] ,
		_w1457_,
		_w1458_,
		_w1666_
	);
	LUT2 #(
		.INIT('he)
	) name1530 (
		_w1665_,
		_w1666_,
		_w1667_
	);
	LUT3 #(
		.INIT('h15)
	) name1531 (
		\shift[6] ,
		_w1467_,
		_w1468_,
		_w1668_
	);
	LUT3 #(
		.INIT('h2a)
	) name1532 (
		\shift[6] ,
		_w1464_,
		_w1465_,
		_w1669_
	);
	LUT2 #(
		.INIT('he)
	) name1533 (
		_w1668_,
		_w1669_,
		_w1670_
	);
	LUT3 #(
		.INIT('h15)
	) name1534 (
		\shift[6] ,
		_w1474_,
		_w1475_,
		_w1671_
	);
	LUT3 #(
		.INIT('h2a)
	) name1535 (
		\shift[6] ,
		_w1471_,
		_w1472_,
		_w1672_
	);
	LUT2 #(
		.INIT('he)
	) name1536 (
		_w1671_,
		_w1672_,
		_w1673_
	);
	LUT3 #(
		.INIT('h15)
	) name1537 (
		\shift[6] ,
		_w1481_,
		_w1482_,
		_w1674_
	);
	LUT3 #(
		.INIT('h2a)
	) name1538 (
		\shift[6] ,
		_w1478_,
		_w1479_,
		_w1675_
	);
	LUT2 #(
		.INIT('he)
	) name1539 (
		_w1674_,
		_w1675_,
		_w1676_
	);
	assign \result[0]  = _w251_ ;
	assign \result[1]  = _w362_ ;
	assign \result[2]  = _w473_ ;
	assign \result[3]  = _w584_ ;
	assign \result[4]  = _w631_ ;
	assign \result[5]  = _w678_ ;
	assign \result[6]  = _w725_ ;
	assign \result[7]  = _w772_ ;
	assign \result[8]  = _w819_ ;
	assign \result[9]  = _w866_ ;
	assign \result[10]  = _w913_ ;
	assign \result[11]  = _w960_ ;
	assign \result[12]  = _w1007_ ;
	assign \result[13]  = _w1054_ ;
	assign \result[14]  = _w1101_ ;
	assign \result[15]  = _w1148_ ;
	assign \result[16]  = _w1155_ ;
	assign \result[17]  = _w1162_ ;
	assign \result[18]  = _w1169_ ;
	assign \result[19]  = _w1176_ ;
	assign \result[20]  = _w1183_ ;
	assign \result[21]  = _w1190_ ;
	assign \result[22]  = _w1197_ ;
	assign \result[23]  = _w1204_ ;
	assign \result[24]  = _w1211_ ;
	assign \result[25]  = _w1218_ ;
	assign \result[26]  = _w1225_ ;
	assign \result[27]  = _w1232_ ;
	assign \result[28]  = _w1239_ ;
	assign \result[29]  = _w1246_ ;
	assign \result[30]  = _w1253_ ;
	assign \result[31]  = _w1260_ ;
	assign \result[32]  = _w1267_ ;
	assign \result[33]  = _w1274_ ;
	assign \result[34]  = _w1281_ ;
	assign \result[35]  = _w1288_ ;
	assign \result[36]  = _w1295_ ;
	assign \result[37]  = _w1302_ ;
	assign \result[38]  = _w1309_ ;
	assign \result[39]  = _w1316_ ;
	assign \result[40]  = _w1323_ ;
	assign \result[41]  = _w1330_ ;
	assign \result[42]  = _w1337_ ;
	assign \result[43]  = _w1344_ ;
	assign \result[44]  = _w1351_ ;
	assign \result[45]  = _w1358_ ;
	assign \result[46]  = _w1365_ ;
	assign \result[47]  = _w1372_ ;
	assign \result[48]  = _w1379_ ;
	assign \result[49]  = _w1386_ ;
	assign \result[50]  = _w1393_ ;
	assign \result[51]  = _w1400_ ;
	assign \result[52]  = _w1407_ ;
	assign \result[53]  = _w1414_ ;
	assign \result[54]  = _w1421_ ;
	assign \result[55]  = _w1428_ ;
	assign \result[56]  = _w1435_ ;
	assign \result[57]  = _w1442_ ;
	assign \result[58]  = _w1449_ ;
	assign \result[59]  = _w1456_ ;
	assign \result[60]  = _w1463_ ;
	assign \result[61]  = _w1470_ ;
	assign \result[62]  = _w1477_ ;
	assign \result[63]  = _w1484_ ;
	assign \result[64]  = _w1487_ ;
	assign \result[65]  = _w1490_ ;
	assign \result[66]  = _w1493_ ;
	assign \result[67]  = _w1496_ ;
	assign \result[68]  = _w1499_ ;
	assign \result[69]  = _w1502_ ;
	assign \result[70]  = _w1505_ ;
	assign \result[71]  = _w1508_ ;
	assign \result[72]  = _w1511_ ;
	assign \result[73]  = _w1514_ ;
	assign \result[74]  = _w1517_ ;
	assign \result[75]  = _w1520_ ;
	assign \result[76]  = _w1523_ ;
	assign \result[77]  = _w1526_ ;
	assign \result[78]  = _w1529_ ;
	assign \result[79]  = _w1532_ ;
	assign \result[80]  = _w1535_ ;
	assign \result[81]  = _w1538_ ;
	assign \result[82]  = _w1541_ ;
	assign \result[83]  = _w1544_ ;
	assign \result[84]  = _w1547_ ;
	assign \result[85]  = _w1550_ ;
	assign \result[86]  = _w1553_ ;
	assign \result[87]  = _w1556_ ;
	assign \result[88]  = _w1559_ ;
	assign \result[89]  = _w1562_ ;
	assign \result[90]  = _w1565_ ;
	assign \result[91]  = _w1568_ ;
	assign \result[92]  = _w1571_ ;
	assign \result[93]  = _w1574_ ;
	assign \result[94]  = _w1577_ ;
	assign \result[95]  = _w1580_ ;
	assign \result[96]  = _w1583_ ;
	assign \result[97]  = _w1586_ ;
	assign \result[98]  = _w1589_ ;
	assign \result[99]  = _w1592_ ;
	assign \result[100]  = _w1595_ ;
	assign \result[101]  = _w1598_ ;
	assign \result[102]  = _w1601_ ;
	assign \result[103]  = _w1604_ ;
	assign \result[104]  = _w1607_ ;
	assign \result[105]  = _w1610_ ;
	assign \result[106]  = _w1613_ ;
	assign \result[107]  = _w1616_ ;
	assign \result[108]  = _w1619_ ;
	assign \result[109]  = _w1622_ ;
	assign \result[110]  = _w1625_ ;
	assign \result[111]  = _w1628_ ;
	assign \result[112]  = _w1631_ ;
	assign \result[113]  = _w1634_ ;
	assign \result[114]  = _w1637_ ;
	assign \result[115]  = _w1640_ ;
	assign \result[116]  = _w1643_ ;
	assign \result[117]  = _w1646_ ;
	assign \result[118]  = _w1649_ ;
	assign \result[119]  = _w1652_ ;
	assign \result[120]  = _w1655_ ;
	assign \result[121]  = _w1658_ ;
	assign \result[122]  = _w1661_ ;
	assign \result[123]  = _w1664_ ;
	assign \result[124]  = _w1667_ ;
	assign \result[125]  = _w1670_ ;
	assign \result[126]  = _w1673_ ;
	assign \result[127]  = _w1676_ ;
endmodule;