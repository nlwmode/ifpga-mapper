module top( \102GAT(31)_pad  , \105GAT(32)_pad  , \108GAT(33)_pad  , \112GAT(34)_pad  , \115GAT(35)_pad  , \11GAT(3)_pad  , \14GAT(4)_pad  , \17GAT(5)_pad  , \1GAT(0)_pad  , \21GAT(6)_pad  , \24GAT(7)_pad  , \27GAT(8)_pad  , \30GAT(9)_pad  , \34GAT(10)_pad  , \37GAT(11)_pad  , \40GAT(12)_pad  , \43GAT(13)_pad  , \47GAT(14)_pad  , \4GAT(1)_pad  , \50GAT(15)_pad  , \53GAT(16)_pad  , \56GAT(17)_pad  , \60GAT(18)_pad  , \63GAT(19)_pad  , \66GAT(20)_pad  , \69GAT(21)_pad  , \73GAT(22)_pad  , \76GAT(23)_pad  , \79GAT(24)_pad  , \82GAT(25)_pad  , \86GAT(26)_pad  , \89GAT(27)_pad  , \8GAT(2)_pad  , \92GAT(28)_pad  , \95GAT(29)_pad  , \99GAT(30)_pad  , \203GAT(82)  , \309GAT(131)  , \360GAT(162)  , \421GAT(188)_pad  , \430GAT(193)_pad  , \431GAT(194)_pad  , \432GAT(195)_pad  );
  input \102GAT(31)_pad  ;
  input \105GAT(32)_pad  ;
  input \108GAT(33)_pad  ;
  input \112GAT(34)_pad  ;
  input \115GAT(35)_pad  ;
  input \11GAT(3)_pad  ;
  input \14GAT(4)_pad  ;
  input \17GAT(5)_pad  ;
  input \1GAT(0)_pad  ;
  input \21GAT(6)_pad  ;
  input \24GAT(7)_pad  ;
  input \27GAT(8)_pad  ;
  input \30GAT(9)_pad  ;
  input \34GAT(10)_pad  ;
  input \37GAT(11)_pad  ;
  input \40GAT(12)_pad  ;
  input \43GAT(13)_pad  ;
  input \47GAT(14)_pad  ;
  input \4GAT(1)_pad  ;
  input \50GAT(15)_pad  ;
  input \53GAT(16)_pad  ;
  input \56GAT(17)_pad  ;
  input \60GAT(18)_pad  ;
  input \63GAT(19)_pad  ;
  input \66GAT(20)_pad  ;
  input \69GAT(21)_pad  ;
  input \73GAT(22)_pad  ;
  input \76GAT(23)_pad  ;
  input \79GAT(24)_pad  ;
  input \82GAT(25)_pad  ;
  input \86GAT(26)_pad  ;
  input \89GAT(27)_pad  ;
  input \8GAT(2)_pad  ;
  input \92GAT(28)_pad  ;
  input \95GAT(29)_pad  ;
  input \99GAT(30)_pad  ;
  output \203GAT(82)  ;
  output \309GAT(131)  ;
  output \360GAT(162)  ;
  output \421GAT(188)_pad  ;
  output \430GAT(193)_pad  ;
  output \431GAT(194)_pad  ;
  output \432GAT(195)_pad  ;
  wire n37 , n38 , n39 , n40 , n41 , n42 , n43 , n44 , n45 , n46 , n47 , n48 , n49 , n50 , n51 , n52 , n53 , n54 , n55 , n56 , n57 , n58 , n59 , n60 , n61 , n62 , n63 , n64 , n65 , n66 , n67 , n68 , n69 , n70 , n71 , n72 , n73 , n74 , n75 , n76 , n77 , n78 , n79 , n80 , n81 , n82 , n83 , n84 , n85 , n86 , n87 , n88 , n89 , n90 , n91 , n92 , n93 , n94 , n95 , n96 , n97 , n98 , n99 , n100 , n101 , n102 , n103 , n104 , n105 , n106 , n107 , n108 , n109 , n110 , n111 , n112 , n113 , n114 , n115 , n116 , n117 , n118 , n119 , n120 , n121 , n122 , n123 , n124 , n125 , n126 , n127 , n128 , n129 , n130 , n131 , n132 , n133 , n134 , n135 , n136 , n137 , n138 , n139 , n140 , n141 , n142 , n143 , n144 , n145 , n146 , n147 , n148 , n149 , n150 , n151 , n152 , n153 , n154 , n155 , n156 , n157 , n158 , n159 , n160 , n161 , n162 , n163 , n164 , n165 ;
  assign n45 = ~\89GAT(27)_pad  & \95GAT(29)_pad  ;
  assign n43 = ~\11GAT(3)_pad  & \17GAT(5)_pad  ;
  assign n44 = ~\1GAT(0)_pad  & \4GAT(1)_pad  ;
  assign n49 = ~n43 & ~n44 ;
  assign n50 = ~n45 & n49 ;
  assign n37 = ~\50GAT(15)_pad  & \56GAT(17)_pad  ;
  assign n38 = ~\24GAT(7)_pad  & \30GAT(9)_pad  ;
  assign n46 = ~n37 & ~n38 ;
  assign n39 = ~\63GAT(19)_pad  & \69GAT(21)_pad  ;
  assign n40 = ~\102GAT(31)_pad  & \108GAT(33)_pad  ;
  assign n47 = ~n39 & ~n40 ;
  assign n41 = ~\76GAT(23)_pad  & \82GAT(25)_pad  ;
  assign n42 = ~\37GAT(11)_pad  & \43GAT(13)_pad  ;
  assign n48 = ~n41 & ~n42 ;
  assign n51 = n47 & n48 ;
  assign n52 = n46 & n51 ;
  assign n53 = n50 & n52 ;
  assign n78 = \76GAT(23)_pad  & ~n53 ;
  assign n79 = ~\76GAT(23)_pad  & n53 ;
  assign n80 = ~n78 & ~n79 ;
  assign n81 = \82GAT(25)_pad  & ~\86GAT(26)_pad  ;
  assign n82 = n80 & n81 ;
  assign n72 = \37GAT(11)_pad  & ~n53 ;
  assign n73 = \43GAT(13)_pad  & ~n72 ;
  assign n74 = ~\47GAT(14)_pad  & n73 ;
  assign n75 = \63GAT(19)_pad  & ~n53 ;
  assign n76 = \69GAT(21)_pad  & ~n75 ;
  assign n77 = ~\73GAT(22)_pad  & n76 ;
  assign n86 = ~n74 & ~n77 ;
  assign n87 = ~n82 & n86 ;
  assign n54 = \1GAT(0)_pad  & ~n53 ;
  assign n55 = \4GAT(1)_pad  & ~n54 ;
  assign n56 = ~\8GAT(2)_pad  & n55 ;
  assign n57 = \50GAT(15)_pad  & ~n53 ;
  assign n58 = \56GAT(17)_pad  & ~n57 ;
  assign n59 = ~\60GAT(18)_pad  & n58 ;
  assign n83 = ~n56 & ~n59 ;
  assign n60 = \89GAT(27)_pad  & ~n53 ;
  assign n61 = \95GAT(29)_pad  & ~n60 ;
  assign n62 = ~\99GAT(30)_pad  & n61 ;
  assign n63 = \24GAT(7)_pad  & ~n53 ;
  assign n64 = \30GAT(9)_pad  & ~n63 ;
  assign n65 = ~\34GAT(10)_pad  & n64 ;
  assign n84 = ~n62 & ~n65 ;
  assign n66 = \11GAT(3)_pad  & ~n53 ;
  assign n67 = \17GAT(5)_pad  & ~n66 ;
  assign n68 = ~\21GAT(6)_pad  & n67 ;
  assign n69 = \102GAT(31)_pad  & ~n53 ;
  assign n70 = \108GAT(33)_pad  & ~n69 ;
  assign n71 = ~\112GAT(34)_pad  & n70 ;
  assign n85 = ~n68 & ~n71 ;
  assign n88 = n84 & n85 ;
  assign n89 = n83 & n88 ;
  assign n90 = n87 & n89 ;
  assign n115 = \86GAT(26)_pad  & ~n90 ;
  assign n116 = \82GAT(25)_pad  & ~n115 ;
  assign n117 = n82 & n90 ;
  assign n118 = ~\92GAT(28)_pad  & n80 ;
  assign n119 = ~n117 & n118 ;
  assign n120 = n116 & n119 ;
  assign n109 = \99GAT(30)_pad  & ~n90 ;
  assign n110 = n61 & ~n109 ;
  assign n111 = ~\105GAT(32)_pad  & n110 ;
  assign n112 = \60GAT(18)_pad  & ~n90 ;
  assign n113 = n58 & ~n112 ;
  assign n114 = ~\66GAT(20)_pad  & n113 ;
  assign n124 = ~n111 & ~n114 ;
  assign n125 = ~n120 & n124 ;
  assign n91 = \34GAT(10)_pad  & ~n90 ;
  assign n92 = n64 & ~n91 ;
  assign n93 = ~\40GAT(12)_pad  & n92 ;
  assign n94 = \21GAT(6)_pad  & ~n90 ;
  assign n95 = n67 & ~n94 ;
  assign n96 = ~\27GAT(8)_pad  & n95 ;
  assign n121 = ~n93 & ~n96 ;
  assign n97 = \73GAT(22)_pad  & ~n90 ;
  assign n98 = n76 & ~n97 ;
  assign n99 = ~\79GAT(24)_pad  & n98 ;
  assign n100 = \112GAT(34)_pad  & ~n90 ;
  assign n101 = n70 & ~n100 ;
  assign n102 = ~\115GAT(35)_pad  & n101 ;
  assign n122 = ~n99 & ~n102 ;
  assign n103 = \47GAT(14)_pad  & ~n90 ;
  assign n104 = n73 & ~n103 ;
  assign n105 = ~\53GAT(16)_pad  & n104 ;
  assign n106 = \8GAT(2)_pad  & ~n90 ;
  assign n107 = n55 & ~n106 ;
  assign n108 = ~\14GAT(4)_pad  & n107 ;
  assign n123 = ~n105 & ~n108 ;
  assign n126 = n122 & n123 ;
  assign n127 = n121 & n126 ;
  assign n128 = n125 & n127 ;
  assign n129 = \66GAT(20)_pad  & ~n128 ;
  assign n130 = n113 & ~n129 ;
  assign n131 = \53GAT(16)_pad  & ~n128 ;
  assign n132 = n104 & ~n131 ;
  assign n133 = ~n130 & ~n132 ;
  assign n134 = \40GAT(12)_pad  & ~n128 ;
  assign n135 = n92 & ~n134 ;
  assign n136 = \27GAT(8)_pad  & ~n128 ;
  assign n137 = n95 & ~n136 ;
  assign n138 = ~n135 & ~n137 ;
  assign n139 = n133 & n138 ;
  assign n140 = \105GAT(32)_pad  & ~n128 ;
  assign n141 = n110 & ~n140 ;
  assign n142 = \115GAT(35)_pad  & ~n128 ;
  assign n143 = n101 & ~n142 ;
  assign n149 = ~n141 & ~n143 ;
  assign n144 = \92GAT(28)_pad  & ~n128 ;
  assign n145 = ~n78 & n116 ;
  assign n146 = ~n144 & n145 ;
  assign n147 = \79GAT(24)_pad  & ~n128 ;
  assign n148 = n98 & ~n147 ;
  assign n150 = ~n146 & ~n148 ;
  assign n151 = n149 & n150 ;
  assign n152 = n139 & n151 ;
  assign n153 = \14GAT(4)_pad  & ~n128 ;
  assign n154 = n107 & ~n153 ;
  assign n155 = ~n152 & ~n154 ;
  assign n156 = ~n135 & n148 ;
  assign n157 = ~n146 & ~n156 ;
  assign n158 = n133 & ~n157 ;
  assign n159 = n138 & ~n158 ;
  assign n160 = n141 & ~n146 ;
  assign n161 = ~n132 & ~n160 ;
  assign n162 = ~n135 & ~n161 ;
  assign n163 = n133 & n156 ;
  assign n164 = ~n137 & ~n163 ;
  assign n165 = ~n162 & n164 ;
  assign \203GAT(82)  = ~n53 ;
  assign \309GAT(131)  = ~n90 ;
  assign \360GAT(162)  = ~n128 ;
  assign \421GAT(188)_pad  = n155 ;
  assign \430GAT(193)_pad  = ~n139 ;
  assign \431GAT(194)_pad  = ~n159 ;
  assign \432GAT(195)_pad  = ~n165 ;
endmodule
