module top( \DATA_0_0_pad  , \DATA_0_10_pad  , \DATA_0_11_pad  , \DATA_0_12_pad  , \DATA_0_13_pad  , \DATA_0_14_pad  , \DATA_0_15_pad  , \DATA_0_16_pad  , \DATA_0_17_pad  , \DATA_0_18_pad  , \DATA_0_19_pad  , \DATA_0_1_pad  , \DATA_0_20_pad  , \DATA_0_21_pad  , \DATA_0_22_pad  , \DATA_0_23_pad  , \DATA_0_24_pad  , \DATA_0_25_pad  , \DATA_0_26_pad  , \DATA_0_27_pad  , \DATA_0_28_pad  , \DATA_0_29_pad  , \DATA_0_2_pad  , \DATA_0_30_pad  , \DATA_0_31_pad  , \DATA_0_3_pad  , \DATA_0_4_pad  , \DATA_0_5_pad  , \DATA_0_6_pad  , \DATA_0_7_pad  , \DATA_0_8_pad  , \DATA_0_9_pad  , RESET_pad , \TM0_pad  , \TM1_pad  , \WX10829_reg/NET0131  , \WX10831_reg/NET0131  , \WX10833_reg/NET0131  , \WX10835_reg/NET0131  , \WX10837_reg/NET0131  , \WX10839_reg/NET0131  , \WX10841_reg/NET0131  , \WX10843_reg/NET0131  , \WX10845_reg/NET0131  , \WX10847_reg/NET0131  , \WX10849_reg/NET0131  , \WX10851_reg/NET0131  , \WX10853_reg/NET0131  , \WX10855_reg/NET0131  , \WX10857_reg/NET0131  , \WX10859_reg/NET0131  , \WX10861_reg/NET0131  , \WX10863_reg/NET0131  , \WX10865_reg/NET0131  , \WX10867_reg/NET0131  , \WX10869_reg/NET0131  , \WX10871_reg/NET0131  , \WX10873_reg/NET0131  , \WX10875_reg/NET0131  , \WX10877_reg/NET0131  , \WX10879_reg/NET0131  , \WX10881_reg/NET0131  , \WX10883_reg/NET0131  , \WX10885_reg/NET0131  , \WX10887_reg/NET0131  , \WX10889_reg/NET0131  , \WX10891_reg/NET0131  , \WX10989_reg/NET0131  , \WX10991_reg/NET0131  , \WX10993_reg/NET0131  , \WX10995_reg/NET0131  , \WX10997_reg/NET0131  , \WX10999_reg/NET0131  , \WX11001_reg/NET0131  , \WX11003_reg/NET0131  , \WX11005_reg/NET0131  , \WX11007_reg/NET0131  , \WX11009_reg/NET0131  , \WX11011_reg/NET0131  , \WX11013_reg/NET0131  , \WX11015_reg/NET0131  , \WX11017_reg/NET0131  , \WX11019_reg/NET0131  , \WX11021_reg/NET0131  , \WX11023_reg/NET0131  , \WX11025_reg/NET0131  , \WX11027_reg/NET0131  , \WX11029_reg/NET0131  , \WX11031_reg/NET0131  , \WX11033_reg/NET0131  , \WX11035_reg/NET0131  , \WX11037_reg/NET0131  , \WX11039_reg/NET0131  , \WX11041_reg/NET0131  , \WX11043_reg/NET0131  , \WX11045_reg/NET0131  , \WX11047_reg/NET0131  , \WX11049_reg/NET0131  , \WX11051_reg/NET0131  , \WX11053_reg/NET0131  , \WX11055_reg/NET0131  , \WX11057_reg/NET0131  , \WX11059_reg/NET0131  , \WX11061_reg/NET0131  , \WX11063_reg/NET0131  , \WX11065_reg/NET0131  , \WX11067_reg/NET0131  , \WX11069_reg/NET0131  , \WX11071_reg/NET0131  , \WX11073_reg/NET0131  , \WX11075_reg/NET0131  , \WX11077_reg/NET0131  , \WX11079_reg/NET0131  , \WX11081_reg/NET0131  , \WX11083_reg/NET0131  , \WX11085_reg/NET0131  , \WX11087_reg/NET0131  , \WX11089_reg/NET0131  , \WX11091_reg/NET0131  , \WX11093_reg/NET0131  , \WX11095_reg/NET0131  , \WX11097_reg/NET0131  , \WX11099_reg/NET0131  , \WX11101_reg/NET0131  , \WX11103_reg/NET0131  , \WX11105_reg/NET0131  , \WX11107_reg/NET0131  , \WX11109_reg/NET0131  , \WX11111_reg/NET0131  , \WX11113_reg/NET0131  , \WX11115_reg/NET0131  , \WX11117_reg/NET0131  , \WX11119_reg/NET0131  , \WX11121_reg/NET0131  , \WX11123_reg/NET0131  , \WX11125_reg/NET0131  , \WX11127_reg/NET0131  , \WX11129_reg/NET0131  , \WX11131_reg/NET0131  , \WX11133_reg/NET0131  , \WX11135_reg/NET0131  , \WX11137_reg/NET0131  , \WX11139_reg/NET0131  , \WX11141_reg/NET0131  , \WX11143_reg/NET0131  , \WX11145_reg/NET0131  , \WX11147_reg/NET0131  , \WX11149_reg/NET0131  , \WX11151_reg/NET0131  , \WX11153_reg/NET0131  , \WX11155_reg/NET0131  , \WX11157_reg/NET0131  , \WX11159_reg/NET0131  , \WX11161_reg/NET0131  , \WX11163_reg/NET0131  , \WX11165_reg/NET0131  , \WX11167_reg/NET0131  , \WX11169_reg/NET0131  , \WX11171_reg/NET0131  , \WX11173_reg/NET0131  , \WX11175_reg/NET0131  , \WX11177_reg/NET0131  , \WX11179_reg/NET0131  , \WX11181_reg/NET0131  , \WX11183_reg/NET0131  , \WX11185_reg/NET0131  , \WX11187_reg/NET0131  , \WX11189_reg/NET0131  , \WX11191_reg/NET0131  , \WX11193_reg/NET0131  , \WX11195_reg/NET0131  , \WX11197_reg/NET0131  , \WX11199_reg/NET0131  , \WX11201_reg/NET0131  , \WX11203_reg/NET0131  , \WX11205_reg/NET0131  , \WX11207_reg/NET0131  , \WX11209_reg/NET0131  , \WX11211_reg/NET0131  , \WX11213_reg/NET0131  , \WX11215_reg/NET0131  , \WX11217_reg/NET0131  , \WX11219_reg/NET0131  , \WX11221_reg/NET0131  , \WX11223_reg/NET0131  , \WX11225_reg/NET0131  , \WX11227_reg/NET0131  , \WX11229_reg/NET0131  , \WX11231_reg/NET0131  , \WX11233_reg/NET0131  , \WX11235_reg/NET0131  , \WX11237_reg/NET0131  , \WX11239_reg/NET0131  , \WX11241_reg/NET0131  , \WX11243_reg/NET0131  , \WX1938_reg/NET0131  , \WX1940_reg/NET0131  , \WX1942_reg/NET0131  , \WX1944_reg/NET0131  , \WX1946_reg/NET0131  , \WX1948_reg/NET0131  , \WX1950_reg/NET0131  , \WX1952_reg/NET0131  , \WX1954_reg/NET0131  , \WX1956_reg/NET0131  , \WX1958_reg/NET0131  , \WX1960_reg/NET0131  , \WX1962_reg/NET0131  , \WX1964_reg/NET0131  , \WX1966_reg/NET0131  , \WX1968_reg/NET0131  , \WX1970_reg/NET0131  , \WX1972_reg/NET0131  , \WX1974_reg/NET0131  , \WX1976_reg/NET0131  , \WX1978_reg/NET0131  , \WX1980_reg/NET0131  , \WX1982_reg/NET0131  , \WX1984_reg/NET0131  , \WX1986_reg/NET0131  , \WX1988_reg/NET0131  , \WX1990_reg/NET0131  , \WX1992_reg/NET0131  , \WX1994_reg/NET0131  , \WX1996_reg/NET0131  , \WX1998_reg/NET0131  , \WX2000_reg/NET0131  , \WX2002_reg/NET0131  , \WX2004_reg/NET0131  , \WX2006_reg/NET0131  , \WX2008_reg/NET0131  , \WX2010_reg/NET0131  , \WX2012_reg/NET0131  , \WX2014_reg/NET0131  , \WX2016_reg/NET0131  , \WX2018_reg/NET0131  , \WX2020_reg/NET0131  , \WX2022_reg/NET0131  , \WX2024_reg/NET0131  , \WX2026_reg/NET0131  , \WX2028_reg/NET0131  , \WX2030_reg/NET0131  , \WX2032_reg/NET0131  , \WX2034_reg/NET0131  , \WX2036_reg/NET0131  , \WX2038_reg/NET0131  , \WX2040_reg/NET0131  , \WX2042_reg/NET0131  , \WX2044_reg/NET0131  , \WX2046_reg/NET0131  , \WX2048_reg/NET0131  , \WX2050_reg/NET0131  , \WX2052_reg/NET0131  , \WX2054_reg/NET0131  , \WX2056_reg/NET0131  , \WX2058_reg/NET0131  , \WX2060_reg/NET0131  , \WX2062_reg/NET0131  , \WX2064_reg/NET0131  , \WX2066_reg/NET0131  , \WX2068_reg/NET0131  , \WX2070_reg/NET0131  , \WX2072_reg/NET0131  , \WX2074_reg/NET0131  , \WX2076_reg/NET0131  , \WX2078_reg/NET0131  , \WX2080_reg/NET0131  , \WX2082_reg/NET0131  , \WX2084_reg/NET0131  , \WX2086_reg/NET0131  , \WX2088_reg/NET0131  , \WX2090_reg/NET0131  , \WX2092_reg/NET0131  , \WX2094_reg/NET0131  , \WX2096_reg/NET0131  , \WX2098_reg/NET0131  , \WX2100_reg/NET0131  , \WX2102_reg/NET0131  , \WX2104_reg/NET0131  , \WX2106_reg/NET0131  , \WX2108_reg/NET0131  , \WX2110_reg/NET0131  , \WX2112_reg/NET0131  , \WX2114_reg/NET0131  , \WX2116_reg/NET0131  , \WX2118_reg/NET0131  , \WX2120_reg/NET0131  , \WX2122_reg/NET0131  , \WX2124_reg/NET0131  , \WX2126_reg/NET0131  , \WX2128_reg/NET0131  , \WX2130_reg/NET0131  , \WX2132_reg/NET0131  , \WX2134_reg/NET0131  , \WX2136_reg/NET0131  , \WX2138_reg/NET0131  , \WX2140_reg/NET0131  , \WX2142_reg/NET0131  , \WX2144_reg/NET0131  , \WX2146_reg/NET0131  , \WX2148_reg/NET0131  , \WX2150_reg/NET0131  , \WX2152_reg/NET0131  , \WX2154_reg/NET0131  , \WX2156_reg/NET0131  , \WX2158_reg/NET0131  , \WX2160_reg/NET0131  , \WX2162_reg/NET0131  , \WX2164_reg/NET0131  , \WX2166_reg/NET0131  , \WX2168_reg/NET0131  , \WX2170_reg/NET0131  , \WX2172_reg/NET0131  , \WX2174_reg/NET0131  , \WX2176_reg/NET0131  , \WX2178_reg/NET0131  , \WX2180_reg/NET0131  , \WX2182_reg/NET0131  , \WX2184_reg/NET0131  , \WX2186_reg/NET0131  , \WX2188_reg/NET0131  , \WX2190_reg/NET0131  , \WX2192_reg/NET0131  , \WX3231_reg/NET0131  , \WX3233_reg/NET0131  , \WX3235_reg/NET0131  , \WX3237_reg/NET0131  , \WX3239_reg/NET0131  , \WX3241_reg/NET0131  , \WX3243_reg/NET0131  , \WX3245_reg/NET0131  , \WX3247_reg/NET0131  , \WX3249_reg/NET0131  , \WX3251_reg/NET0131  , \WX3253_reg/NET0131  , \WX3255_reg/NET0131  , \WX3257_reg/NET0131  , \WX3259_reg/NET0131  , \WX3261_reg/NET0131  , \WX3263_reg/NET0131  , \WX3265_reg/NET0131  , \WX3267_reg/NET0131  , \WX3269_reg/NET0131  , \WX3271_reg/NET0131  , \WX3273_reg/NET0131  , \WX3275_reg/NET0131  , \WX3277_reg/NET0131  , \WX3279_reg/NET0131  , \WX3281_reg/NET0131  , \WX3283_reg/NET0131  , \WX3285_reg/NET0131  , \WX3287_reg/NET0131  , \WX3289_reg/NET0131  , \WX3291_reg/NET0131  , \WX3293_reg/NET0131  , \WX3295_reg/NET0131  , \WX3297_reg/NET0131  , \WX3299_reg/NET0131  , \WX3301_reg/NET0131  , \WX3303_reg/NET0131  , \WX3305_reg/NET0131  , \WX3307_reg/NET0131  , \WX3309_reg/NET0131  , \WX3311_reg/NET0131  , \WX3313_reg/NET0131  , \WX3315_reg/NET0131  , \WX3317_reg/NET0131  , \WX3319_reg/NET0131  , \WX3321_reg/NET0131  , \WX3323_reg/NET0131  , \WX3325_reg/NET0131  , \WX3327_reg/NET0131  , \WX3329_reg/NET0131  , \WX3331_reg/NET0131  , \WX3333_reg/NET0131  , \WX3335_reg/NET0131  , \WX3337_reg/NET0131  , \WX3339_reg/NET0131  , \WX3341_reg/NET0131  , \WX3343_reg/NET0131  , \WX3345_reg/NET0131  , \WX3347_reg/NET0131  , \WX3349_reg/NET0131  , \WX3351_reg/NET0131  , \WX3353_reg/NET0131  , \WX3355_reg/NET0131  , \WX3357_reg/NET0131  , \WX3359_reg/NET0131  , \WX3361_reg/NET0131  , \WX3363_reg/NET0131  , \WX3365_reg/NET0131  , \WX3367_reg/NET0131  , \WX3369_reg/NET0131  , \WX3371_reg/NET0131  , \WX3373_reg/NET0131  , \WX3375_reg/NET0131  , \WX3377_reg/NET0131  , \WX3379_reg/NET0131  , \WX3381_reg/NET0131  , \WX3383_reg/NET0131  , \WX3385_reg/NET0131  , \WX3387_reg/NET0131  , \WX3389_reg/NET0131  , \WX3391_reg/NET0131  , \WX3393_reg/NET0131  , \WX3395_reg/NET0131  , \WX3397_reg/NET0131  , \WX3399_reg/NET0131  , \WX3401_reg/NET0131  , \WX3403_reg/NET0131  , \WX3405_reg/NET0131  , \WX3407_reg/NET0131  , \WX3409_reg/NET0131  , \WX3411_reg/NET0131  , \WX3413_reg/NET0131  , \WX3415_reg/NET0131  , \WX3417_reg/NET0131  , \WX3419_reg/NET0131  , \WX3421_reg/NET0131  , \WX3423_reg/NET0131  , \WX3425_reg/NET0131  , \WX3427_reg/NET0131  , \WX3429_reg/NET0131  , \WX3431_reg/NET0131  , \WX3433_reg/NET0131  , \WX3435_reg/NET0131  , \WX3437_reg/NET0131  , \WX3439_reg/NET0131  , \WX3441_reg/NET0131  , \WX3443_reg/NET0131  , \WX3445_reg/NET0131  , \WX3447_reg/NET0131  , \WX3449_reg/NET0131  , \WX3451_reg/NET0131  , \WX3453_reg/NET0131  , \WX3455_reg/NET0131  , \WX3457_reg/NET0131  , \WX3459_reg/NET0131  , \WX3461_reg/NET0131  , \WX3463_reg/NET0131  , \WX3465_reg/NET0131  , \WX3467_reg/NET0131  , \WX3469_reg/NET0131  , \WX3471_reg/NET0131  , \WX3473_reg/NET0131  , \WX3475_reg/NET0131  , \WX3477_reg/NET0131  , \WX3479_reg/NET0131  , \WX3481_reg/NET0131  , \WX3483_reg/NET0131  , \WX3485_reg/NET0131  , \WX4524_reg/NET0131  , \WX4526_reg/NET0131  , \WX4528_reg/NET0131  , \WX4530_reg/NET0131  , \WX4532_reg/NET0131  , \WX4534_reg/NET0131  , \WX4536_reg/NET0131  , \WX4538_reg/NET0131  , \WX4540_reg/NET0131  , \WX4542_reg/NET0131  , \WX4544_reg/NET0131  , \WX4546_reg/NET0131  , \WX4548_reg/NET0131  , \WX4550_reg/NET0131  , \WX4552_reg/NET0131  , \WX4554_reg/NET0131  , \WX4556_reg/NET0131  , \WX4558_reg/NET0131  , \WX4560_reg/NET0131  , \WX4562_reg/NET0131  , \WX4564_reg/NET0131  , \WX4566_reg/NET0131  , \WX4568_reg/NET0131  , \WX4570_reg/NET0131  , \WX4572_reg/NET0131  , \WX4574_reg/NET0131  , \WX4576_reg/NET0131  , \WX4578_reg/NET0131  , \WX4580_reg/NET0131  , \WX4582_reg/NET0131  , \WX4584_reg/NET0131  , \WX4586_reg/NET0131  , \WX4588_reg/NET0131  , \WX4590_reg/NET0131  , \WX4592_reg/NET0131  , \WX4594_reg/NET0131  , \WX4596_reg/NET0131  , \WX4598_reg/NET0131  , \WX4600_reg/NET0131  , \WX4602_reg/NET0131  , \WX4604_reg/NET0131  , \WX4606_reg/NET0131  , \WX4608_reg/NET0131  , \WX4610_reg/NET0131  , \WX4612_reg/NET0131  , \WX4614_reg/NET0131  , \WX4616_reg/NET0131  , \WX4618_reg/NET0131  , \WX4620_reg/NET0131  , \WX4622_reg/NET0131  , \WX4624_reg/NET0131  , \WX4626_reg/NET0131  , \WX4628_reg/NET0131  , \WX4630_reg/NET0131  , \WX4632_reg/NET0131  , \WX4634_reg/NET0131  , \WX4636_reg/NET0131  , \WX4638_reg/NET0131  , \WX4640_reg/NET0131  , \WX4642_reg/NET0131  , \WX4644_reg/NET0131  , \WX4646_reg/NET0131  , \WX4648_reg/NET0131  , \WX4650_reg/NET0131  , \WX4652_reg/NET0131  , \WX4654_reg/NET0131  , \WX4656_reg/NET0131  , \WX4658_reg/NET0131  , \WX4660_reg/NET0131  , \WX4662_reg/NET0131  , \WX4664_reg/NET0131  , \WX4666_reg/NET0131  , \WX4668_reg/NET0131  , \WX4670_reg/NET0131  , \WX4672_reg/NET0131  , \WX4674_reg/NET0131  , \WX4676_reg/NET0131  , \WX4678_reg/NET0131  , \WX4680_reg/NET0131  , \WX4682_reg/NET0131  , \WX4684_reg/NET0131  , \WX4686_reg/NET0131  , \WX4688_reg/NET0131  , \WX4690_reg/NET0131  , \WX4692_reg/NET0131  , \WX4694_reg/NET0131  , \WX4696_reg/NET0131  , \WX4698_reg/NET0131  , \WX4700_reg/NET0131  , \WX4702_reg/NET0131  , \WX4704_reg/NET0131  , \WX4706_reg/NET0131  , \WX4708_reg/NET0131  , \WX4710_reg/NET0131  , \WX4712_reg/NET0131  , \WX4714_reg/NET0131  , \WX4716_reg/NET0131  , \WX4718_reg/NET0131  , \WX4720_reg/NET0131  , \WX4722_reg/NET0131  , \WX4724_reg/NET0131  , \WX4726_reg/NET0131  , \WX4728_reg/NET0131  , \WX4730_reg/NET0131  , \WX4732_reg/NET0131  , \WX4734_reg/NET0131  , \WX4736_reg/NET0131  , \WX4738_reg/NET0131  , \WX4740_reg/NET0131  , \WX4742_reg/NET0131  , \WX4744_reg/NET0131  , \WX4746_reg/NET0131  , \WX4748_reg/NET0131  , \WX4750_reg/NET0131  , \WX4752_reg/NET0131  , \WX4754_reg/NET0131  , \WX4756_reg/NET0131  , \WX4758_reg/NET0131  , \WX4760_reg/NET0131  , \WX4762_reg/NET0131  , \WX4764_reg/NET0131  , \WX4766_reg/NET0131  , \WX4768_reg/NET0131  , \WX4770_reg/NET0131  , \WX4772_reg/NET0131  , \WX4774_reg/NET0131  , \WX4776_reg/NET0131  , \WX4778_reg/NET0131  , \WX5817_reg/NET0131  , \WX5819_reg/NET0131  , \WX5821_reg/NET0131  , \WX5823_reg/NET0131  , \WX5825_reg/NET0131  , \WX5827_reg/NET0131  , \WX5829_reg/NET0131  , \WX5831_reg/NET0131  , \WX5833_reg/NET0131  , \WX5835_reg/NET0131  , \WX5837_reg/NET0131  , \WX5839_reg/NET0131  , \WX5841_reg/NET0131  , \WX5843_reg/NET0131  , \WX5845_reg/NET0131  , \WX5847_reg/NET0131  , \WX5849_reg/NET0131  , \WX5851_reg/NET0131  , \WX5853_reg/NET0131  , \WX5855_reg/NET0131  , \WX5857_reg/NET0131  , \WX5859_reg/NET0131  , \WX5861_reg/NET0131  , \WX5863_reg/NET0131  , \WX5865_reg/NET0131  , \WX5867_reg/NET0131  , \WX5869_reg/NET0131  , \WX5871_reg/NET0131  , \WX5873_reg/NET0131  , \WX5875_reg/NET0131  , \WX5877_reg/NET0131  , \WX5879_reg/NET0131  , \WX5881_reg/NET0131  , \WX5883_reg/NET0131  , \WX5885_reg/NET0131  , \WX5887_reg/NET0131  , \WX5889_reg/NET0131  , \WX5891_reg/NET0131  , \WX5893_reg/NET0131  , \WX5895_reg/NET0131  , \WX5897_reg/NET0131  , \WX5899_reg/NET0131  , \WX5901_reg/NET0131  , \WX5903_reg/NET0131  , \WX5905_reg/NET0131  , \WX5907_reg/NET0131  , \WX5909_reg/NET0131  , \WX5911_reg/NET0131  , \WX5913_reg/NET0131  , \WX5915_reg/NET0131  , \WX5917_reg/NET0131  , \WX5919_reg/NET0131  , \WX5921_reg/NET0131  , \WX5923_reg/NET0131  , \WX5925_reg/NET0131  , \WX5927_reg/NET0131  , \WX5929_reg/NET0131  , \WX5931_reg/NET0131  , \WX5933_reg/NET0131  , \WX5935_reg/NET0131  , \WX5937_reg/NET0131  , \WX5939_reg/NET0131  , \WX5941_reg/NET0131  , \WX5943_reg/NET0131  , \WX5945_reg/NET0131  , \WX5947_reg/NET0131  , \WX5949_reg/NET0131  , \WX5951_reg/NET0131  , \WX5953_reg/NET0131  , \WX5955_reg/NET0131  , \WX5957_reg/NET0131  , \WX5959_reg/NET0131  , \WX5961_reg/NET0131  , \WX5963_reg/NET0131  , \WX5965_reg/NET0131  , \WX5967_reg/NET0131  , \WX5969_reg/NET0131  , \WX5971_reg/NET0131  , \WX5973_reg/NET0131  , \WX5975_reg/NET0131  , \WX5977_reg/NET0131  , \WX5979_reg/NET0131  , \WX5981_reg/NET0131  , \WX5983_reg/NET0131  , \WX5985_reg/NET0131  , \WX5987_reg/NET0131  , \WX5989_reg/NET0131  , \WX5991_reg/NET0131  , \WX5993_reg/NET0131  , \WX5995_reg/NET0131  , \WX5997_reg/NET0131  , \WX5999_reg/NET0131  , \WX6001_reg/NET0131  , \WX6003_reg/NET0131  , \WX6005_reg/NET0131  , \WX6007_reg/NET0131  , \WX6009_reg/NET0131  , \WX6011_reg/NET0131  , \WX6013_reg/NET0131  , \WX6015_reg/NET0131  , \WX6017_reg/NET0131  , \WX6019_reg/NET0131  , \WX6021_reg/NET0131  , \WX6023_reg/NET0131  , \WX6025_reg/NET0131  , \WX6027_reg/NET0131  , \WX6029_reg/NET0131  , \WX6031_reg/NET0131  , \WX6033_reg/NET0131  , \WX6035_reg/NET0131  , \WX6037_reg/NET0131  , \WX6039_reg/NET0131  , \WX6041_reg/NET0131  , \WX6043_reg/NET0131  , \WX6045_reg/NET0131  , \WX6047_reg/NET0131  , \WX6049_reg/NET0131  , \WX6051_reg/NET0131  , \WX6053_reg/NET0131  , \WX6055_reg/NET0131  , \WX6057_reg/NET0131  , \WX6059_reg/NET0131  , \WX6061_reg/NET0131  , \WX6063_reg/NET0131  , \WX6065_reg/NET0131  , \WX6067_reg/NET0131  , \WX6069_reg/NET0131  , \WX6071_reg/NET0131  , \WX645_reg/NET0131  , \WX647_reg/NET0131  , \WX649_reg/NET0131  , \WX651_reg/NET0131  , \WX653_reg/NET0131  , \WX655_reg/NET0131  , \WX657_reg/NET0131  , \WX659_reg/NET0131  , \WX661_reg/NET0131  , \WX663_reg/NET0131  , \WX665_reg/NET0131  , \WX667_reg/NET0131  , \WX669_reg/NET0131  , \WX671_reg/NET0131  , \WX673_reg/NET0131  , \WX675_reg/NET0131  , \WX677_reg/NET0131  , \WX679_reg/NET0131  , \WX681_reg/NET0131  , \WX683_reg/NET0131  , \WX685_reg/NET0131  , \WX687_reg/NET0131  , \WX689_reg/NET0131  , \WX691_reg/NET0131  , \WX693_reg/NET0131  , \WX695_reg/NET0131  , \WX697_reg/NET0131  , \WX699_reg/NET0131  , \WX701_reg/NET0131  , \WX703_reg/NET0131  , \WX705_reg/NET0131  , \WX707_reg/NET0131  , \WX709_reg/NET0131  , \WX7110_reg/NET0131  , \WX7112_reg/NET0131  , \WX7114_reg/NET0131  , \WX7116_reg/NET0131  , \WX7118_reg/NET0131  , \WX711_reg/NET0131  , \WX7120_reg/NET0131  , \WX7122_reg/NET0131  , \WX7124_reg/NET0131  , \WX7126_reg/NET0131  , \WX7128_reg/NET0131  , \WX7130_reg/NET0131  , \WX7132_reg/NET0131  , \WX7134_reg/NET0131  , \WX7136_reg/NET0131  , \WX7138_reg/NET0131  , \WX713_reg/NET0131  , \WX7140_reg/NET0131  , \WX7142_reg/NET0131  , \WX7144_reg/NET0131  , \WX7146_reg/NET0131  , \WX7148_reg/NET0131  , \WX7150_reg/NET0131  , \WX7152_reg/NET0131  , \WX7154_reg/NET0131  , \WX7156_reg/NET0131  , \WX7158_reg/NET0131  , \WX715_reg/NET0131  , \WX7160_reg/NET0131  , \WX7162_reg/NET0131  , \WX7164_reg/NET0131  , \WX7166_reg/NET0131  , \WX7168_reg/NET0131  , \WX7170_reg/NET0131  , \WX7172_reg/NET0131  , \WX7174_reg/NET0131  , \WX7176_reg/NET0131  , \WX7178_reg/NET0131  , \WX717_reg/NET0131  , \WX7180_reg/NET0131  , \WX7182_reg/NET0131  , \WX7184_reg/NET0131  , \WX7186_reg/NET0131  , \WX7188_reg/NET0131  , \WX7190_reg/NET0131  , \WX7192_reg/NET0131  , \WX7194_reg/NET0131  , \WX7196_reg/NET0131  , \WX7198_reg/NET0131  , \WX719_reg/NET0131  , \WX7200_reg/NET0131  , \WX7202_reg/NET0131  , \WX7204_reg/NET0131  , \WX7206_reg/NET0131  , \WX7208_reg/NET0131  , \WX7210_reg/NET0131  , \WX7212_reg/NET0131  , \WX7214_reg/NET0131  , \WX7216_reg/NET0131  , \WX7218_reg/NET0131  , \WX721_reg/NET0131  , \WX7220_reg/NET0131  , \WX7222_reg/NET0131  , \WX7224_reg/NET0131  , \WX7226_reg/NET0131  , \WX7228_reg/NET0131  , \WX7230_reg/NET0131  , \WX7232_reg/NET0131  , \WX7234_reg/NET0131  , \WX7236_reg/NET0131  , \WX7238_reg/NET0131  , \WX723_reg/NET0131  , \WX7240_reg/NET0131  , \WX7242_reg/NET0131  , \WX7244_reg/NET0131  , \WX7246_reg/NET0131  , \WX7248_reg/NET0131  , \WX7250_reg/NET0131  , \WX7252_reg/NET0131  , \WX7254_reg/NET0131  , \WX7256_reg/NET0131  , \WX7258_reg/NET0131  , \WX725_reg/NET0131  , \WX7260_reg/NET0131  , \WX7262_reg/NET0131  , \WX7264_reg/NET0131  , \WX7266_reg/NET0131  , \WX7268_reg/NET0131  , \WX7270_reg/NET0131  , \WX7272_reg/NET0131  , \WX7274_reg/NET0131  , \WX7276_reg/NET0131  , \WX7278_reg/NET0131  , \WX727_reg/NET0131  , \WX7280_reg/NET0131  , \WX7282_reg/NET0131  , \WX7284_reg/NET0131  , \WX7286_reg/NET0131  , \WX7288_reg/NET0131  , \WX7290_reg/NET0131  , \WX7292_reg/NET0131  , \WX7294_reg/NET0131  , \WX7296_reg/NET0131  , \WX7298_reg/NET0131  , \WX729_reg/NET0131  , \WX7300_reg/NET0131  , \WX7302_reg/NET0131  , \WX7304_reg/NET0131  , \WX7306_reg/NET0131  , \WX7308_reg/NET0131  , \WX7310_reg/NET0131  , \WX7312_reg/NET0131  , \WX7314_reg/NET0131  , \WX7316_reg/NET0131  , \WX7318_reg/NET0131  , \WX731_reg/NET0131  , \WX7320_reg/NET0131  , \WX7322_reg/NET0131  , \WX7324_reg/NET0131  , \WX7326_reg/NET0131  , \WX7328_reg/NET0131  , \WX7330_reg/NET0131  , \WX7332_reg/NET0131  , \WX7334_reg/NET0131  , \WX7336_reg/NET0131  , \WX7338_reg/NET0131  , \WX733_reg/NET0131  , \WX7340_reg/NET0131  , \WX7342_reg/NET0131  , \WX7344_reg/NET0131  , \WX7346_reg/NET0131  , \WX7348_reg/NET0131  , \WX7350_reg/NET0131  , \WX7352_reg/NET0131  , \WX7354_reg/NET0131  , \WX7356_reg/NET0131  , \WX7358_reg/NET0131  , \WX735_reg/NET0131  , \WX7360_reg/NET0131  , \WX7362_reg/NET0131  , \WX7364_reg/NET0131  , \WX737_reg/NET0131  , \WX739_reg/NET0131  , \WX741_reg/NET0131  , \WX743_reg/NET0131  , \WX745_reg/NET0131  , \WX747_reg/NET0131  , \WX749_reg/NET0131  , \WX751_reg/NET0131  , \WX753_reg/NET0131  , \WX755_reg/NET0131  , \WX757_reg/NET0131  , \WX759_reg/NET0131  , \WX761_reg/NET0131  , \WX763_reg/NET0131  , \WX765_reg/NET0131  , \WX767_reg/NET0131  , \WX769_reg/NET0131  , \WX771_reg/NET0131  , \WX773_reg/NET0131  , \WX775_reg/NET0131  , \WX777_reg/NET0131  , \WX779_reg/NET0131  , \WX781_reg/NET0131  , \WX783_reg/NET0131  , \WX785_reg/NET0131  , \WX787_reg/NET0131  , \WX789_reg/NET0131  , \WX791_reg/NET0131  , \WX793_reg/NET0131  , \WX795_reg/NET0131  , \WX797_reg/NET0131  , \WX799_reg/NET0131  , \WX801_reg/NET0131  , \WX803_reg/NET0131  , \WX805_reg/NET0131  , \WX807_reg/NET0131  , \WX809_reg/NET0131  , \WX811_reg/NET0131  , \WX813_reg/NET0131  , \WX815_reg/NET0131  , \WX817_reg/NET0131  , \WX819_reg/NET0131  , \WX821_reg/NET0131  , \WX823_reg/NET0131  , \WX825_reg/NET0131  , \WX827_reg/NET0131  , \WX829_reg/NET0131  , \WX831_reg/NET0131  , \WX833_reg/NET0131  , \WX835_reg/NET0131  , \WX837_reg/NET0131  , \WX839_reg/NET0131  , \WX8403_reg/NET0131  , \WX8405_reg/NET0131  , \WX8407_reg/NET0131  , \WX8409_reg/NET0131  , \WX8411_reg/NET0131  , \WX8413_reg/NET0131  , \WX8415_reg/NET0131  , \WX8417_reg/NET0131  , \WX8419_reg/NET0131  , \WX841_reg/NET0131  , \WX8421_reg/NET0131  , \WX8423_reg/NET0131  , \WX8425_reg/NET0131  , \WX8427_reg/NET0131  , \WX8429_reg/NET0131  , \WX8431_reg/NET0131  , \WX8433_reg/NET0131  , \WX8435_reg/NET0131  , \WX8437_reg/NET0131  , \WX8439_reg/NET0131  , \WX843_reg/NET0131  , \WX8441_reg/NET0131  , \WX8443_reg/NET0131  , \WX8445_reg/NET0131  , \WX8447_reg/NET0131  , \WX8449_reg/NET0131  , \WX8451_reg/NET0131  , \WX8453_reg/NET0131  , \WX8455_reg/NET0131  , \WX8457_reg/NET0131  , \WX8459_reg/NET0131  , \WX845_reg/NET0131  , \WX8461_reg/NET0131  , \WX8463_reg/NET0131  , \WX8465_reg/NET0131  , \WX8467_reg/NET0131  , \WX8469_reg/NET0131  , \WX8471_reg/NET0131  , \WX8473_reg/NET0131  , \WX8475_reg/NET0131  , \WX8477_reg/NET0131  , \WX8479_reg/NET0131  , \WX847_reg/NET0131  , \WX8481_reg/NET0131  , \WX8483_reg/NET0131  , \WX8485_reg/NET0131  , \WX8487_reg/NET0131  , \WX8489_reg/NET0131  , \WX8491_reg/NET0131  , \WX8493_reg/NET0131  , \WX8495_reg/NET0131  , \WX8497_reg/NET0131  , \WX8499_reg/NET0131  , \WX849_reg/NET0131  , \WX8501_reg/NET0131  , \WX8503_reg/NET0131  , \WX8505_reg/NET0131  , \WX8507_reg/NET0131  , \WX8509_reg/NET0131  , \WX8511_reg/NET0131  , \WX8513_reg/NET0131  , \WX8515_reg/NET0131  , \WX8517_reg/NET0131  , \WX8519_reg/NET0131  , \WX851_reg/NET0131  , \WX8521_reg/NET0131  , \WX8523_reg/NET0131  , \WX8525_reg/NET0131  , \WX8527_reg/NET0131  , \WX8529_reg/NET0131  , \WX8531_reg/NET0131  , \WX8533_reg/NET0131  , \WX8535_reg/NET0131  , \WX8537_reg/NET0131  , \WX8539_reg/NET0131  , \WX853_reg/NET0131  , \WX8541_reg/NET0131  , \WX8543_reg/NET0131  , \WX8545_reg/NET0131  , \WX8547_reg/NET0131  , \WX8549_reg/NET0131  , \WX8551_reg/NET0131  , \WX8553_reg/NET0131  , \WX8555_reg/NET0131  , \WX8557_reg/NET0131  , \WX8559_reg/NET0131  , \WX855_reg/NET0131  , \WX8561_reg/NET0131  , \WX8563_reg/NET0131  , \WX8565_reg/NET0131  , \WX8567_reg/NET0131  , \WX8569_reg/NET0131  , \WX8571_reg/NET0131  , \WX8573_reg/NET0131  , \WX8575_reg/NET0131  , \WX8577_reg/NET0131  , \WX8579_reg/NET0131  , \WX857_reg/NET0131  , \WX8581_reg/NET0131  , \WX8583_reg/NET0131  , \WX8585_reg/NET0131  , \WX8587_reg/NET0131  , \WX8589_reg/NET0131  , \WX8591_reg/NET0131  , \WX8593_reg/NET0131  , \WX8595_reg/NET0131  , \WX8597_reg/NET0131  , \WX8599_reg/NET0131  , \WX859_reg/NET0131  , \WX8601_reg/NET0131  , \WX8603_reg/NET0131  , \WX8605_reg/NET0131  , \WX8607_reg/NET0131  , \WX8609_reg/NET0131  , \WX8611_reg/NET0131  , \WX8613_reg/NET0131  , \WX8615_reg/NET0131  , \WX8617_reg/NET0131  , \WX8619_reg/NET0131  , \WX861_reg/NET0131  , \WX8621_reg/NET0131  , \WX8623_reg/NET0131  , \WX8625_reg/NET0131  , \WX8627_reg/NET0131  , \WX8629_reg/NET0131  , \WX8631_reg/NET0131  , \WX8633_reg/NET0131  , \WX8635_reg/NET0131  , \WX8637_reg/NET0131  , \WX8639_reg/NET0131  , \WX863_reg/NET0131  , \WX8641_reg/NET0131  , \WX8643_reg/NET0131  , \WX8645_reg/NET0131  , \WX8647_reg/NET0131  , \WX8649_reg/NET0131  , \WX8651_reg/NET0131  , \WX8653_reg/NET0131  , \WX8655_reg/NET0131  , \WX8657_reg/NET0131  , \WX865_reg/NET0131  , \WX867_reg/NET0131  , \WX869_reg/NET0131  , \WX871_reg/NET0131  , \WX873_reg/NET0131  , \WX875_reg/NET0131  , \WX877_reg/NET0131  , \WX879_reg/NET0131  , \WX881_reg/NET0131  , \WX883_reg/NET0131  , \WX885_reg/NET0131  , \WX887_reg/NET0131  , \WX889_reg/NET0131  , \WX891_reg/NET0131  , \WX893_reg/NET0131  , \WX895_reg/NET0131  , \WX897_reg/NET0131  , \WX899_reg/NET0131  , \WX9696_reg/NET0131  , \WX9698_reg/NET0131  , \WX9700_reg/NET0131  , \WX9702_reg/NET0131  , \WX9704_reg/NET0131  , \WX9706_reg/NET0131  , \WX9708_reg/NET0131  , \WX9710_reg/NET0131  , \WX9712_reg/NET0131  , \WX9714_reg/NET0131  , \WX9716_reg/NET0131  , \WX9718_reg/NET0131  , \WX9720_reg/NET0131  , \WX9722_reg/NET0131  , \WX9724_reg/NET0131  , \WX9726_reg/NET0131  , \WX9728_reg/NET0131  , \WX9730_reg/NET0131  , \WX9732_reg/NET0131  , \WX9734_reg/NET0131  , \WX9736_reg/NET0131  , \WX9738_reg/NET0131  , \WX9740_reg/NET0131  , \WX9742_reg/NET0131  , \WX9744_reg/NET0131  , \WX9746_reg/NET0131  , \WX9748_reg/NET0131  , \WX9750_reg/NET0131  , \WX9752_reg/NET0131  , \WX9754_reg/NET0131  , \WX9756_reg/NET0131  , \WX9758_reg/NET0131  , \WX9760_reg/NET0131  , \WX9762_reg/NET0131  , \WX9764_reg/NET0131  , \WX9766_reg/NET0131  , \WX9768_reg/NET0131  , \WX9770_reg/NET0131  , \WX9772_reg/NET0131  , \WX9774_reg/NET0131  , \WX9776_reg/NET0131  , \WX9778_reg/NET0131  , \WX9780_reg/NET0131  , \WX9782_reg/NET0131  , \WX9784_reg/NET0131  , \WX9786_reg/NET0131  , \WX9788_reg/NET0131  , \WX9790_reg/NET0131  , \WX9792_reg/NET0131  , \WX9794_reg/NET0131  , \WX9796_reg/NET0131  , \WX9798_reg/NET0131  , \WX9800_reg/NET0131  , \WX9802_reg/NET0131  , \WX9804_reg/NET0131  , \WX9806_reg/NET0131  , \WX9808_reg/NET0131  , \WX9810_reg/NET0131  , \WX9812_reg/NET0131  , \WX9814_reg/NET0131  , \WX9816_reg/NET0131  , \WX9818_reg/NET0131  , \WX9820_reg/NET0131  , \WX9822_reg/NET0131  , \WX9824_reg/NET0131  , \WX9826_reg/NET0131  , \WX9828_reg/NET0131  , \WX9830_reg/NET0131  , \WX9832_reg/NET0131  , \WX9834_reg/NET0131  , \WX9836_reg/NET0131  , \WX9838_reg/NET0131  , \WX9840_reg/NET0131  , \WX9842_reg/NET0131  , \WX9844_reg/NET0131  , \WX9846_reg/NET0131  , \WX9848_reg/NET0131  , \WX9850_reg/NET0131  , \WX9852_reg/NET0131  , \WX9854_reg/NET0131  , \WX9856_reg/NET0131  , \WX9858_reg/NET0131  , \WX9860_reg/NET0131  , \WX9862_reg/NET0131  , \WX9864_reg/NET0131  , \WX9866_reg/NET0131  , \WX9868_reg/NET0131  , \WX9870_reg/NET0131  , \WX9872_reg/NET0131  , \WX9874_reg/NET0131  , \WX9876_reg/NET0131  , \WX9878_reg/NET0131  , \WX9880_reg/NET0131  , \WX9882_reg/NET0131  , \WX9884_reg/NET0131  , \WX9886_reg/NET0131  , \WX9888_reg/NET0131  , \WX9890_reg/NET0131  , \WX9892_reg/NET0131  , \WX9894_reg/NET0131  , \WX9896_reg/NET0131  , \WX9898_reg/NET0131  , \WX9900_reg/NET0131  , \WX9902_reg/NET0131  , \WX9904_reg/NET0131  , \WX9906_reg/NET0131  , \WX9908_reg/NET0131  , \WX9910_reg/NET0131  , \WX9912_reg/NET0131  , \WX9914_reg/NET0131  , \WX9916_reg/NET0131  , \WX9918_reg/NET0131  , \WX9920_reg/NET0131  , \WX9922_reg/NET0131  , \WX9924_reg/NET0131  , \WX9926_reg/NET0131  , \WX9928_reg/NET0131  , \WX9930_reg/NET0131  , \WX9932_reg/NET0131  , \WX9934_reg/NET0131  , \WX9936_reg/NET0131  , \WX9938_reg/NET0131  , \WX9940_reg/NET0131  , \WX9942_reg/NET0131  , \WX9944_reg/NET0131  , \WX9946_reg/NET0131  , \WX9948_reg/NET0131  , \WX9950_reg/NET0131  , \_2077__reg/NET0131  , \_2078__reg/NET0131  , \_2079__reg/NET0131  , \_2080__reg/NET0131  , \_2081__reg/NET0131  , \_2082__reg/NET0131  , \_2083__reg/NET0131  , \_2084__reg/NET0131  , \_2085__reg/NET0131  , \_2086__reg/NET0131  , \_2087__reg/NET0131  , \_2088__reg/NET0131  , \_2089__reg/NET0131  , \_2090__reg/NET0131  , \_2091__reg/NET0131  , \_2092__reg/NET0131  , \_2093__reg/NET0131  , \_2094__reg/NET0131  , \_2095__reg/NET0131  , \_2096__reg/NET0131  , \_2097__reg/NET0131  , \_2098__reg/NET0131  , \_2099__reg/NET0131  , \_2100__reg/NET0131  , \_2101__reg/NET0131  , \_2102__reg/NET0131  , \_2103__reg/NET0131  , \_2104__reg/NET0131  , \_2105__reg/NET0131  , \_2106__reg/NET0131  , \_2107__reg/NET0131  , \_2108__reg/NET0131  , \_2109__reg/NET0131  , \_2110__reg/NET0131  , \_2111__reg/NET0131  , \_2112__reg/NET0131  , \_2113__reg/NET0131  , \_2114__reg/NET0131  , \_2115__reg/NET0131  , \_2116__reg/NET0131  , \_2117__reg/NET0131  , \_2118__reg/NET0131  , \_2119__reg/NET0131  , \_2120__reg/NET0131  , \_2121__reg/NET0131  , \_2122__reg/NET0131  , \_2123__reg/NET0131  , \_2124__reg/NET0131  , \_2125__reg/NET0131  , \_2126__reg/NET0131  , \_2127__reg/NET0131  , \_2128__reg/NET0131  , \_2129__reg/NET0131  , \_2130__reg/NET0131  , \_2131__reg/NET0131  , \_2132__reg/NET0131  , \_2133__reg/NET0131  , \_2134__reg/NET0131  , \_2135__reg/NET0131  , \_2136__reg/NET0131  , \_2137__reg/NET0131  , \_2138__reg/NET0131  , \_2139__reg/NET0131  , \_2140__reg/NET0131  , \_2141__reg/NET0131  , \_2142__reg/NET0131  , \_2143__reg/NET0131  , \_2144__reg/NET0131  , \_2145__reg/NET0131  , \_2146__reg/NET0131  , \_2147__reg/NET0131  , \_2148__reg/NET0131  , \_2149__reg/NET0131  , \_2150__reg/NET0131  , \_2151__reg/NET0131  , \_2152__reg/NET0131  , \_2153__reg/NET0131  , \_2154__reg/NET0131  , \_2155__reg/NET0131  , \_2156__reg/NET0131  , \_2157__reg/NET0131  , \_2158__reg/NET0131  , \_2159__reg/NET0131  , \_2160__reg/NET0131  , \_2161__reg/NET0131  , \_2162__reg/NET0131  , \_2163__reg/NET0131  , \_2164__reg/NET0131  , \_2165__reg/NET0131  , \_2166__reg/NET0131  , \_2167__reg/NET0131  , \_2168__reg/NET0131  , \_2169__reg/NET0131  , \_2170__reg/NET0131  , \_2171__reg/NET0131  , \_2172__reg/NET0131  , \_2173__reg/NET0131  , \_2174__reg/NET0131  , \_2175__reg/NET0131  , \_2176__reg/NET0131  , \_2177__reg/NET0131  , \_2178__reg/NET0131  , \_2179__reg/NET0131  , \_2180__reg/NET0131  , \_2181__reg/NET0131  , \_2182__reg/NET0131  , \_2183__reg/NET0131  , \_2184__reg/NET0131  , \_2185__reg/NET0131  , \_2186__reg/NET0131  , \_2187__reg/NET0131  , \_2188__reg/NET0131  , \_2189__reg/NET0131  , \_2190__reg/NET0131  , \_2191__reg/NET0131  , \_2192__reg/NET0131  , \_2193__reg/NET0131  , \_2194__reg/NET0131  , \_2195__reg/NET0131  , \_2196__reg/NET0131  , \_2197__reg/NET0131  , \_2198__reg/NET0131  , \_2199__reg/NET0131  , \_2200__reg/NET0131  , \_2201__reg/NET0131  , \_2202__reg/NET0131  , \_2203__reg/NET0131  , \_2204__reg/NET0131  , \_2205__reg/NET0131  , \_2206__reg/NET0131  , \_2207__reg/NET0131  , \_2208__reg/NET0131  , \_2209__reg/NET0131  , \_2210__reg/NET0131  , \_2211__reg/NET0131  , \_2212__reg/NET0131  , \_2213__reg/NET0131  , \_2214__reg/NET0131  , \_2215__reg/NET0131  , \_2216__reg/NET0131  , \_2217__reg/NET0131  , \_2218__reg/NET0131  , \_2219__reg/NET0131  , \_2220__reg/NET0131  , \_2221__reg/NET0131  , \_2222__reg/NET0131  , \_2223__reg/NET0131  , \_2224__reg/NET0131  , \_2225__reg/NET0131  , \_2226__reg/NET0131  , \_2227__reg/NET0131  , \_2228__reg/NET0131  , \_2229__reg/NET0131  , \_2230__reg/NET0131  , \_2231__reg/NET0131  , \_2232__reg/NET0131  , \_2233__reg/NET0131  , \_2234__reg/NET0131  , \_2235__reg/NET0131  , \_2236__reg/NET0131  , \_2237__reg/NET0131  , \_2238__reg/NET0131  , \_2239__reg/NET0131  , \_2240__reg/NET0131  , \_2241__reg/NET0131  , \_2242__reg/NET0131  , \_2243__reg/NET0131  , \_2244__reg/NET0131  , \_2245__reg/NET0131  , \_2246__reg/NET0131  , \_2247__reg/NET0131  , \_2248__reg/NET0131  , \_2249__reg/NET0131  , \_2250__reg/NET0131  , \_2251__reg/NET0131  , \_2252__reg/NET0131  , \_2253__reg/NET0131  , \_2254__reg/NET0131  , \_2255__reg/NET0131  , \_2256__reg/NET0131  , \_2257__reg/NET0131  , \_2258__reg/NET0131  , \_2259__reg/NET0131  , \_2260__reg/NET0131  , \_2261__reg/NET0131  , \_2262__reg/NET0131  , \_2263__reg/NET0131  , \_2264__reg/NET0131  , \_2265__reg/NET0131  , \_2266__reg/NET0131  , \_2267__reg/NET0131  , \_2268__reg/NET0131  , \_2269__reg/NET0131  , \_2270__reg/NET0131  , \_2271__reg/NET0131  , \_2272__reg/NET0131  , \_2273__reg/NET0131  , \_2274__reg/NET0131  , \_2275__reg/NET0131  , \_2276__reg/NET0131  , \_2277__reg/NET0131  , \_2278__reg/NET0131  , \_2279__reg/NET0131  , \_2280__reg/NET0131  , \_2281__reg/NET0131  , \_2282__reg/NET0131  , \_2283__reg/NET0131  , \_2284__reg/NET0131  , \_2285__reg/NET0131  , \_2286__reg/NET0131  , \_2287__reg/NET0131  , \_2288__reg/NET0131  , \_2289__reg/NET0131  , \_2290__reg/NET0131  , \_2291__reg/NET0131  , \_2292__reg/NET0131  , \_2293__reg/NET0131  , \_2294__reg/NET0131  , \_2295__reg/NET0131  , \_2296__reg/NET0131  , \_2297__reg/NET0131  , \_2298__reg/NET0131  , \_2299__reg/NET0131  , \_2300__reg/NET0131  , \_2301__reg/NET0131  , \_2302__reg/NET0131  , \_2303__reg/NET0131  , \_2304__reg/NET0131  , \_2305__reg/NET0131  , \_2306__reg/NET0131  , \_2307__reg/NET0131  , \_2308__reg/NET0131  , \_2309__reg/NET0131  , \_2310__reg/NET0131  , \_2311__reg/NET0131  , \_2312__reg/NET0131  , \_2313__reg/NET0131  , \_2314__reg/NET0131  , \_2315__reg/NET0131  , \_2316__reg/NET0131  , \_2317__reg/NET0131  , \_2318__reg/NET0131  , \_2319__reg/NET0131  , \_2320__reg/NET0131  , \_2321__reg/NET0131  , \_2322__reg/NET0131  , \_2323__reg/NET0131  , \_2324__reg/NET0131  , \_2325__reg/NET0131  , \_2326__reg/NET0131  , \_2327__reg/NET0131  , \_2328__reg/NET0131  , \_2329__reg/NET0131  , \_2330__reg/NET0131  , \_2331__reg/NET0131  , \_2332__reg/NET0131  , \_2333__reg/NET0131  , \_2334__reg/NET0131  , \_2335__reg/NET0131  , \_2336__reg/NET0131  , \_2337__reg/NET0131  , \_2338__reg/NET0131  , \_2339__reg/NET0131  , \_2340__reg/NET0131  , \_2341__reg/NET0131  , \_2342__reg/NET0131  , \_2343__reg/NET0131  , \_2344__reg/NET0131  , \_2345__reg/NET0131  , \_2346__reg/NET0131  , \_2347__reg/NET0131  , \_2348__reg/NET0131  , \_2349__reg/NET0131  , \_2350__reg/NET0131  , \_2351__reg/NET0131  , \_2352__reg/NET0131  , \_2353__reg/NET0131  , \_2354__reg/NET0131  , \_2355__reg/NET0131  , \_2356__reg/NET0131  , \_2357__reg/NET0131  , \_2358__reg/NET0131  , \_2359__reg/NET0131  , \_2360__reg/NET0131  , \_2361__reg/NET0131  , \_2362__reg/NET0131  , \_2363__reg/NET0131  , \_2364__reg/NET0131  , \DATA_9_0_pad  , \DATA_9_10_pad  , \DATA_9_11_pad  , \DATA_9_12_pad  , \DATA_9_13_pad  , \DATA_9_14_pad  , \DATA_9_15_pad  , \DATA_9_16_pad  , \DATA_9_17_pad  , \DATA_9_18_pad  , \DATA_9_19_pad  , \DATA_9_1_pad  , \DATA_9_20_pad  , \DATA_9_21_pad  , \DATA_9_22_pad  , \DATA_9_23_pad  , \DATA_9_24_pad  , \DATA_9_25_pad  , \DATA_9_26_pad  , \DATA_9_27_pad  , \DATA_9_28_pad  , \DATA_9_29_pad  , \DATA_9_2_pad  , \DATA_9_30_pad  , \DATA_9_31_pad  , \DATA_9_3_pad  , \DATA_9_4_pad  , \DATA_9_5_pad  , \DATA_9_6_pad  , \DATA_9_7_pad  , \DATA_9_8_pad  , \DATA_9_9_pad  , \_al_n0  , \_al_n1  , \g19/_0_  , \g35/_0_  , \g36/_0_  , \g40/_0_  , \g55780/_0_  , \g55783/_0_  , \g55795/_0_  , \g55796/_0_  , \g55797/_0_  , \g55798/_0_  , \g55799/_0_  , \g55800/_0_  , \g55801/_0_  , \g55802/_0_  , \g55803/_0_  , \g55834/_0_  , \g55835/_0_  , \g55836/_0_  , \g55837/_0_  , \g55838/_0_  , \g55839/_0_  , \g55840/_0_  , \g55841/_0_  , \g55842/_0_  , \g55856/_0_  , \g55894/_0_  , \g55895/_0_  , \g55896/_0_  , \g55897/_0_  , \g55898/_0_  , \g55899/_0_  , \g55900/_0_  , \g55901/_0_  , \g55902/_0_  , \g55916/_0_  , \g55953/_0_  , \g55954/_0_  , \g55955/_0_  , \g55956/_0_  , \g55957/_0_  , \g55958/_0_  , \g55959/_0_  , \g55960/_0_  , \g55961/_0_  , \g55975/_0_  , \g56012/_0_  , \g56013/_0_  , \g56014/_0_  , \g56015/_0_  , \g56016/_0_  , \g56017/_0_  , \g56018/_0_  , \g56019/_0_  , \g56020/_0_  , \g56034/_0_  , \g56071/_0_  , \g56072/_0_  , \g56073/_0_  , \g56074/_0_  , \g56075/_0_  , \g56076/_0_  , \g56077/_0_  , \g56078/_0_  , \g56079/_0_  , \g56093/_0_  , \g56130/_0_  , \g56131/_0_  , \g56132/_0_  , \g56133/_0_  , \g56134/_0_  , \g56135/_0_  , \g56136/_0_  , \g56137/_0_  , \g56138/_0_  , \g56152/_0_  , \g56189/_0_  , \g56190/_0_  , \g56191/_0_  , \g56192/_0_  , \g56193/_0_  , \g56194/_0_  , \g56195/_0_  , \g56196/_0_  , \g56197/_0_  , \g56211/_0_  , \g56248/_0_  , \g56249/_0_  , \g56250/_0_  , \g56251/_0_  , \g56252/_0_  , \g56253/_0_  , \g56254/_0_  , \g56255/_0_  , \g56256/_0_  , \g56270/_0_  , \g56307/_0_  , \g56308/_0_  , \g56309/_0_  , \g56310/_0_  , \g56311/_0_  , \g56312/_0_  , \g56313/_0_  , \g56314/_0_  , \g56315/_0_  , \g56329/_0_  , \g56366/_0_  , \g56367/_0_  , \g56368/_0_  , \g56369/_0_  , \g56370/_0_  , \g56371/_0_  , \g56372/_0_  , \g56373/_0_  , \g56374/_0_  , \g56388/_0_  , \g56425/_0_  , \g56426/_0_  , \g56427/_0_  , \g56428/_0_  , \g56429/_0_  , \g56430/_0_  , \g56431/_0_  , \g56432/_0_  , \g56433/_0_  , \g56447/_0_  , \g56484/_0_  , \g56485/_0_  , \g56486/_0_  , \g56487/_0_  , \g56488/_0_  , \g56489/_0_  , \g56490/_0_  , \g56491/_0_  , \g56492/_0_  , \g56507/_0_  , \g56543/_0_  , \g56544/_0_  , \g56545/_0_  , \g56546/_0_  , \g56547/_0_  , \g56548/_0_  , \g56549/_0_  , \g56551/_0_  , \g56567/_0_  , \g56602/_0_  , \g56603/_0_  , \g56604/_0_  , \g56605/_0_  , \g56606/_0_  , \g56607/_0_  , \g56608/_0_  , \g56610/_0_  , \g56627/_0_  , \g56661/_0_  , \g56662/_0_  , \g56663/_0_  , \g56664/_0_  , \g56665/_0_  , \g56666/_0_  , \g56667/_0_  , \g56668/_0_  , \g56686/_0_  , \g56720/_0_  , \g56721/_0_  , \g56722/_0_  , \g56723/_0_  , \g56724/_0_  , \g56725/_0_  , \g56726/_0_  , \g56727/_0_  , \g56728/_0_  , \g56745/_0_  , \g56779/_0_  , \g56780/_0_  , \g56781/_0_  , \g56782/_0_  , \g56783/_0_  , \g56784/_0_  , \g56785/_0_  , \g56804/_0_  , \g56838/_0_  , \g56839/_0_  , \g56840/_0_  , \g56841/_0_  , \g56842/_0_  , \g56843/_0_  , \g56844/_0_  , \g56845/_0_  , \g56846/_0_  , \g56863/_0_  , \g56897/_0_  , \g56898/_0_  , \g56899/_0_  , \g56900/_0_  , \g56901/_0_  , \g56902/_0_  , \g56903/_0_  , \g56905/_0_  , \g56921/_0_  , \g56956/_0_  , \g56957/_0_  , \g56958/_0_  , \g56959/_0_  , \g56960/_0_  , \g56961/_0_  , \g56962/_0_  , \g56964/_0_  , \g56980/_0_  , \g57015/_0_  , \g57016/_0_  , \g57017/_0_  , \g57018/_0_  , \g57019/_0_  , \g57020/_0_  , \g57021/_0_  , \g57023/_0_  , \g57040/_0_  , \g57074/_0_  , \g57075/_0_  , \g57076/_0_  , \g57077/_0_  , \g57078/_0_  , \g57079/_0_  , \g57080/_0_  , \g57081/_0_  , \g57099/_0_  , \g57133/_0_  , \g57134/_0_  , \g57135/_0_  , \g57136/_0_  , \g57137/_0_  , \g57138/_0_  , \g57139/_0_  , \g57140/_0_  , \g57141/_0_  , \g57159/_0_  , \g57193/_0_  , \g57195/_0_  , \g57196/_0_  , \g57197/_0_  , \g57198/_0_  , \g57199/_0_  , \g57200/_0_  , \g57202/_0_  , \g57219/_0_  , \g57254/_0_  , \g57255/_0_  , \g57256/_0_  , \g57257/_0_  , \g57258/_0_  , \g57259/_0_  , \g57260/_0_  , \g57262/_0_  , \g57263/_0_  , \g57285/_0_  , \g57318/_0_  , \g57319/_0_  , \g57320/_0_  , \g57321/_0_  , \g57322/_0_  , \g57323/_0_  , \g57324/_0_  , \g57325/_0_  , \g57326/_0_  , \g57328/_0_  , \g57329/_0_  , \g57330/_0_  , \g57350/_0_  , \g57387/_0_  , \g57388/_0_  , \g57390/_0_  , \g57391/_0_  , \g57392/_0_  , \g57393/_0_  , \g57395/_0_  , \g57396/_0_  , \g57439/_0_  , \g57476/_0_  , \g57477/_0_  , \g57478/_0_  , \g57479/_0_  , \g57480/_0_  , \g57481/_0_  , \g57482/_0_  , \g57483/_0_  , \g57484/_0_  , \g57485/_0_  , \g57486/_0_  , \g57487/_0_  , \g57488/_0_  , \g57489/_0_  , \g57490/_0_  , \g57491/_0_  , \g57492/_0_  , \g57493/_0_  , \g57494/_0_  , \g57495/_0_  , \g57496/_0_  , \g57497/_0_  , \g57498/_0_  , \g57499/_0_  , \g57500/_0_  , \g57501/_0_  , \g57502/_0_  , \g57503/_0_  , \g57504/_0_  , \g57505/_0_  , \g57524/_0_  , \g57537/_0_  , \g57541/_0_  , \g57543/_0_  , \g58163/_0_  , \g58572/_0_  , \g58573/_0_  , \g58574/_0_  , \g58575/_0_  , \g58576/_0_  , \g58577/_0_  , \g58578/_0_  , \g58579/_0_  , \g58580/_0_  , \g58581/_0_  , \g58582/_0_  , \g58583/_0_  , \g58584/_0_  , \g58585/_0_  , \g58586/_0_  , \g58587/_0_  , \g58588/_0_  , \g58589/_0_  , \g58590/_0_  , \g58591/_0_  , \g58592/_0_  , \g58593/_0_  , \g58594/_0_  , \g58595/_0_  , \g58596/_0_  , \g58597/_0_  , \g58598/_0_  , \g58600/_0_  , \g58602/_0_  , \g58604/_0_  , \g58615/_0_  , \g59240/_0_  , \g59241/_0_  , \g59242/_0_  , \g59243/_0_  , \g59244/_0_  , \g59245/_0_  , \g59246/_0_  , \g59247/_0_  , \g59248/_0_  , \g59249/_0_  , \g59250/_0_  , \g59251/_0_  , \g59252/_0_  , \g59253/_0_  , \g59254/_0_  , \g59255/_0_  , \g59256/_0_  , \g59257/_0_  , \g59258/_0_  , \g59259/_0_  , \g59260/_0_  , \g59261/_0_  , \g59262/_0_  , \g59263/_0_  , \g59264/_0_  , \g59265/_0_  , \g59266/_0_  , \g59267/_0_  , \g59268/_0_  , \g59269/_0_  , \g59270/_0_  , \g59271/_0_  , \g59272/_0_  , \g59273/_0_  , \g59274/_0_  , \g59275/_0_  , \g59276/_0_  , \g59277/_0_  , \g59278/_0_  , \g59279/_0_  , \g59280/_0_  , \g59281/_0_  , \g59282/_0_  , \g59283/_0_  , \g59284/_0_  , \g59285/_0_  , \g59286/_0_  , \g59287/_0_  , \g59288/_0_  , \g59289/_0_  , \g59290/_0_  , \g59291/_0_  , \g59292/_0_  , \g59293/_0_  , \g59294/_0_  , \g59295/_0_  , \g59296/_0_  , \g59297/_0_  , \g59298/_0_  , \g59299/_0_  , \g59300/_0_  , \g59301/_0_  , \g59302/_0_  , \g59303/_0_  , \g59304/_0_  , \g59305/_0_  , \g59306/_0_  , \g59307/_0_  , \g59308/_0_  , \g59309/_0_  , \g59310/_0_  , \g59311/_0_  , \g59312/_0_  , \g59313/_0_  , \g59314/_0_  , \g59315/_0_  , \g59316/_0_  , \g59317/_0_  , \g59318/_0_  , \g59319/_0_  , \g59320/_0_  , \g59321/_0_  , \g59322/_0_  , \g59323/_0_  , \g59324/_0_  , \g59325/_0_  , \g59326/_0_  , \g59327/_0_  , \g59328/_0_  , \g59329/_0_  , \g59330/_0_  , \g59331/_0_  , \g59332/_0_  , \g59333/_0_  , \g59334/_0_  , \g59335/_0_  , \g59336/_0_  , \g59337/_0_  , \g59338/_0_  , \g59339/_0_  , \g59340/_0_  , \g59341/_0_  , \g59342/_0_  , \g59343/_0_  , \g59344/_0_  , \g59345/_0_  , \g59346/_0_  , \g59347/_0_  , \g59348/_0_  , \g59349/_0_  , \g59350/_0_  , \g59351/_0_  , \g59352/_0_  , \g59353/_0_  , \g59354/_0_  , \g59355/_0_  , \g59356/_0_  , \g59357/_0_  , \g59358/_0_  , \g59359/_0_  , \g59360/_0_  , \g59361/_0_  , \g59362/_0_  , \g59363/_0_  , \g59364/_0_  , \g59365/_0_  , \g59366/_0_  , \g59367/_0_  , \g59368/_0_  , \g59369/_0_  , \g59370/_0_  , \g59371/_0_  , \g59372/_0_  , \g59373/_0_  , \g59374/_0_  , \g59375/_0_  , \g59376/_0_  , \g59377/_0_  , \g59378/_0_  , \g59379/_0_  , \g59380/_0_  , \g59381/_0_  , \g59382/_0_  , \g59383/_0_  , \g59384/_0_  , \g59385/_0_  , \g59386/_0_  , \g59387/_0_  , \g59388/_0_  , \g59389/_0_  , \g59390/_0_  , \g59391/_0_  , \g59392/_0_  , \g59393/_0_  , \g59394/_0_  , \g59395/_0_  , \g59396/_0_  , \g59397/_0_  , \g59398/_0_  , \g59399/_0_  , \g59400/_0_  , \g59401/_0_  , \g59402/_0_  , \g59403/_0_  , \g59404/_0_  , \g59405/_0_  , \g59406/_0_  , \g59407/_0_  , \g59408/_0_  , \g59409/_0_  , \g59410/_0_  , \g59411/_0_  , \g59412/_0_  , \g59413/_0_  , \g59414/_0_  , \g59415/_0_  , \g59416/_0_  , \g59417/_0_  , \g59418/_0_  , \g59419/_0_  , \g59420/_0_  , \g59421/_0_  , \g59422/_0_  , \g59423/_0_  , \g59424/_0_  , \g59425/_0_  , \g59426/_0_  , \g59427/_0_  , \g59428/_0_  , \g59429/_0_  , \g59430/_0_  , \g59431/_0_  , \g59432/_0_  , \g59433/_0_  , \g59434/_0_  , \g59435/_0_  , \g59436/_0_  , \g59437/_0_  , \g59438/_0_  , \g59439/_0_  , \g59440/_0_  , \g59441/_0_  , \g59442/_0_  , \g59443/_0_  , \g59444/_0_  , \g59445/_0_  , \g59446/_0_  , \g59447/_0_  , \g59448/_0_  , \g59449/_0_  , \g59450/_0_  , \g59451/_0_  , \g59452/_0_  , \g59453/_0_  , \g59454/_0_  , \g59455/_0_  , \g59456/_0_  , \g59457/_0_  , \g59458/_0_  , \g59459/_0_  , \g59460/_0_  , \g59461/_0_  , \g59462/_0_  , \g59463/_0_  , \g59464/_0_  , \g59465/_0_  , \g59466/_0_  , \g59467/_0_  , \g59468/_0_  , \g59469/_0_  , \g59470/_0_  , \g59471/_0_  , \g59472/_0_  , \g59473/_0_  , \g59474/_0_  , \g59475/_0_  , \g59476/_0_  , \g59477/_0_  , \g59478/_0_  , \g59479/_0_  , \g59480/_0_  , \g59481/_0_  , \g59482/_0_  , \g59483/_0_  , \g59484/_0_  , \g59485/_0_  , \g59486/_0_  , \g59487/_0_  , \g59488/_0_  , \g59489/_0_  , \g59490/_0_  , \g59491/_0_  , \g59492/_0_  , \g59493/_0_  , \g59494/_0_  , \g59495/_0_  , \g59496/_0_  , \g59497/_0_  , \g59498/_0_  , \g59500/_0_  , \g59503/_0_  , \g59512/_0_  , \g61336/_0_  , \g61521/_0_  , \g61523/_0_  , \g61524/_0_  , \g61526/_0_  , \g61527/_0_  , \g61528/_0_  , \g61529/_0_  , \g61530/_0_  , \g61531/_0_  , \g61532/_0_  , \g61533/_0_  , \g61535/_0_  , \g61537/_0_  , \g61539/_0_  , \g61540/_0_  , \g61541/_0_  , \g61542/_0_  , \g61546/_0_  , \g61550/_0_  , \g61551/_0_  , \g61552/_0_  , \g61554/_0_  , \g61555/_0_  , \g61556/_0_  , \g61558/_0_  , \g61559/_0_  , \g61561/_0_  , \g61562/_0_  , \g61563/_0_  , \g61564/_0_  , \g61565/_0_  , \g61566/_0_  , \g61568/_0_  , \g61570/_0_  , \g61571/_0_  , \g61572/_0_  , \g61573/_0_  , \g61577/_0_  , \g61578/_0_  , \g61579/_0_  , \g61580/_0_  , \g61581/_0_  , \g61582/_0_  , \g61583/_0_  , \g61584/_0_  , \g61585/_0_  , \g61586/_0_  , \g61587/_0_  , \g61588/_0_  , \g61589/_0_  , \g61591/_0_  , \g61592/_0_  , \g61594/_0_  , \g61595/_0_  , \g61596/_0_  , \g61597/_0_  , \g61598/_0_  , \g61599/_0_  , \g61600/_0_  , \g61601/_0_  , \g61605/_0_  , \g61606/_0_  , \g61607/_0_  , \g61608/_0_  , \g61609/_0_  , \g61610/_0_  , \g61611/_0_  , \g61612/_0_  , \g61613/_0_  , \g61615/_0_  , \g61616/_0_  , \g61617/_0_  , \g61618/_0_  , \g61619/_0_  , \g61620/_0_  , \g61621/_0_  , \g61623/_0_  , \g61624/_0_  , \g61625/_0_  , \g61626/_0_  , \g61627/_0_  , \g61629/_0_  , \g61630/_0_  , \g61631/_0_  , \g61632/_0_  , \g61633/_0_  , \g61634/_0_  , \g61636/_0_  , \g61638/_0_  , \g61639/_0_  , \g61640/_0_  , \g61641/_0_  , \g61642/_0_  , \g61644/_0_  , \g61647/_0_  , \g61648/_0_  , \g61649/_0_  , \g61650/_0_  , \g61653/_0_  , \g61654/_0_  , \g61655/_0_  , \g61656/_0_  , \g61658/_0_  , \g61661/_0_  , \g61662/_0_  , \g61663/_0_  , \g61664/_0_  , \g61666/_0_  , \g61667/_0_  , \g61668/_0_  , \g61670/_0_  , \g61671/_0_  , \g61672/_0_  , \g61673/_0_  , \g61675/_0_  , \g61676/_0_  , \g61680/_0_  , \g61681/_0_  , \g61682/_0_  , \g61683/_0_  , \g61684/_0_  , \g61686/_0_  , \g61687/_0_  , \g61688/_0_  , \g61689/_0_  , \g61690/_0_  , \g61691/_0_  , \g61693/_0_  , \g61694/_0_  , \g61696/_0_  , \g61697/_0_  , \g61698/_0_  , \g61699/_0_  , \g61700/_0_  , \g61701/_0_  , \g61702/_0_  , \g61703/_0_  , \g61704/_0_  , \g61705/_0_  , \g61706/_0_  , \g61707/_0_  , \g61708/_0_  , \g61711/_0_  , \g61712/_0_  , \g61714/_0_  , \g61716/_0_  , \g61717/_0_  , \g61719/_0_  , \g61720/_0_  , \g61721/_0_  , \g61724/_0_  , \g61725/_0_  , \g61728/_0_  , \g61729/_0_  , \g61731/_0_  , \g61732/_0_  , \g61733/_0_  , \g61736/_0_  , \g61737/_0_  , \g61739/_0_  , \g61740/_0_  , \g61741/_0_  , \g61743/_0_  , \g61744/_0_  , \g61745/_0_  , \g61746/_0_  , \g61747/_0_  , \g61748/_0_  , \g61749/_0_  , \g61750/_0_  , \g61751/_0_  , \g61752/_0_  , \g61753/_0_  , \g61754/_0_  , \g61755/_0_  , \g61757/_0_  , \g61758/_0_  , \g61759/_0_  , \g61760/_0_  , \g61761/_0_  , \g61762/_0_  , \g61763/_0_  , \g61764/_0_  , \g61765/_0_  , \g61766/_0_  , \g61767/_0_  , \g61768/_0_  , \g61769/_0_  , \g61770/_0_  , \g61771/_0_  , \g61772/_0_  , \g61773/_0_  , \g61774/_0_  , \g61775/_0_  , \g61776/_0_  , \g61777/_0_  , \g61778/_0_  , \g61780/_0_  , \g61781/_0_  , \g61783/_0_  , \g61784/_0_  , \g61786/_0_  , \g61787/_0_  , \g61790/_0_  , \g61791/_0_  , \g61794/_0_  , \g61795/_0_  , \g61796/_0_  , \g61797/_0_  , \g61798/_0_  , \g61799/_0_  , \g61800/_0_  , \g61801/_0_  , \g61802/_0_  , \g61803/_0_  , \g61805/_0_  , \g61806/_0_  , \g61807/_0_  , \g61808/_0_  , \g61809/_0_  , \g61810/_0_  , \g61811/_0_  , \g61812/_0_  , \g61813/_0_  , \g61816/_0_  , \g61817/_0_  , \g61818/_0_  , \g61820/_0_  , \g61822/_0_  , \g61823/_0_  , \g61825/_0_  , \g61826/_0_  , \g61827/_0_  , \g61828/_0_  , \g61829/_0_  , \g61832/_0_  , \g61834/_0_  , \g61835/_0_  , \g61837/_0_  , \g61838/_0_  , \g61839/_0_  , \g61840/_0_  , \g61844/_0_  , \g61847/_0_  , \g61848/_0_  , \g61849/_0_  , \g61850/_0_  , \g61851/_0_  , \g61853/_0_  , \g61854/_0_  , \g61855/_0_  , \g61856/_0_  , \g61858/_0_  , \g61859/_0_  , \g61861/_0_  , \g61862/_0_  , \g61863/_0_  , \g61864/_0_  , \g61865/_0_  , \g61866/_0_  , \g61867/_0_  , \g61868/_0_  , \g61869/_0_  , \g61870/_0_  , \g61871/_0_  , \g61873/_0_  , \g61874/_0_  , \g61875/_0_  , \g61877/_0_  , \g61878/_0_  , \g61879/_0_  , \g61880/_0_  , \g61881/_0_  , \g61883/_0_  , \g61884/_0_  , \g61886/_0_  , \g61887/_0_  , \g61890/_0_  , \g61891/_0_  , \g61892/_0_  , \g61893/_0_  , \g61894/_0_  , \g61895/_0_  , \g61900/_0_  , \g61901/_0_  , \g61902/_0_  , \g61904/_0_  , \g61905/_0_  , \g61906/_0_  , \g61907/_0_  , \g61914/_0_  , \g61915/_0_  , \g61917/_0_  , \g61919/_0_  , \g61921/_0_  , \g61924/_0_  , \g61925/_0_  , \g61926/_0_  , \g61927/_0_  , \g61928/_0_  , \g61929/_0_  , \g61930/_0_  , \g61931/_0_  , \g61932/_0_  , \g61933/_0_  , \g61934/_0_  , \g61935/_0_  , \g61936/_0_  , \g61937/_0_  , \g61938/_0_  , \g61939/_0_  , \g61943/_0_  , \g61944/_0_  , \g61945/_0_  , \g61947/_0_  , \g61948/_0_  , \g61949/_0_  , \g61950/_0_  , \g61951/_0_  , \g61952/_0_  , \g61953/_0_  , \g61955/_0_  , \g61956/_0_  , \g61957/_0_  , \g61958/_0_  , \g61959/_0_  , \g61960/_0_  , \g61961/_0_  , \g61962/_0_  , \g61963/_0_  , \g61964/_0_  , \g61965/_0_  , \g61966/_0_  , \g61967/_0_  , \g61968/_0_  , \g61969/_0_  , \g61970/_0_  , \g61971/_0_  , \g61972/_0_  , \g61973/_0_  , \g61974/_0_  , \g61976/_0_  , \g61978/_0_  , \g61980/_0_  , \g61981/_0_  , \g61982/_0_  , \g61983/_0_  , \g61984/_0_  , \g61985/_0_  , \g61986/_0_  , \g61987/_0_  , \g61988/_0_  , \g61989/_0_  , \g61990/_0_  , \g61992/_0_  , \g61994/_0_  , \g61995/_0_  , \g61996/_0_  , \g61997/_0_  , \g61998/_0_  , \g62000/_0_  , \g62001/_0_  , \g62002/_0_  , \g62003/_0_  , \g62004/_0_  , \g62005/_0_  , \g62007/_0_  , \g62008/_0_  , \g62009/_0_  , \g62010/_0_  , \g62011/_0_  , \g62012/_0_  , \g62013/_0_  , \g62014/_0_  , \g62015/_0_  , \g62016/_0_  , \g62017/_0_  , \g62018/_0_  , \g62019/_0_  , \g62020/_0_  , \g62021/_0_  , \g62022/_0_  , \g62023/_0_  , \g62024/_0_  , \g62025/_0_  , \g62026/_0_  , \g62027/_0_  , \g62030/_0_  , \g62033/_0_  , \g62034/_0_  , \g62036/_0_  , \g62038/_0_  , \g62041/_0_  , \g62042/_0_  , \g62043/_0_  , \g62044/_0_  , \g62045/_0_  , \g62046/_0_  , \g62047/_0_  , \g62048/_0_  , \g62050/_0_  , \g62051/_0_  , \g62052/_0_  , \g62055/_0_  , \g62057/_0_  , \g62058/_0_  , \g62059/_0_  , \g62060/_0_  , \g62061/_0_  , \g62062/_0_  , \g62064/_0_  , \g62065/_0_  , \g62066/_0_  , \g62067/_0_  , \g62068/_0_  , \g62072/_0_  , \g62073/_0_  , \g62074/_0_  , \g62075/_0_  , \g62076/_0_  , \g62077/_0_  , \g62078/_0_  , \g62080/_0_  , \g62081/_0_  , \g62082/_0_  , \g62084/_0_  , \g62085/_0_  , \g62086/_0_  , \g62087/_0_  , \g62088/_0_  , \g62089/_0_  , \g62090/_0_  , \g62091/_0_  , \g62092/_0_  , \g62094/_0_  , \g62096/_0_  , \g62097/_0_  , \g62098/_0_  , \g62099/_0_  , \g62100/_0_  , \g62101/_0_  , \g62102/_0_  , \g62104/_0_  , \g62106/_0_  , \g62107/_0_  , \g62108/_0_  , \g62110/_0_  , \g62112/_0_  , \g62113/_0_  , \g62114/_0_  , \g62116/_0_  , \g62117/_0_  , \g62118/_0_  , \g62119/_0_  , \g62120/_0_  , \g62121/_0_  , \g62122/_0_  , \g62124/_0_  , \g62126/_0_  , \g62127/_0_  , \g62128/_0_  , \g62129/_0_  , \g62130/_0_  , \g62131/_0_  , \g62132/_0_  , \g62133/_0_  , \g62135/_0_  , \g62136/_0_  , \g62137/_0_  , \g62138/_0_  , \g62140/_0_  , \g62143/_0_  , \g62144/_0_  , \g62149/_0_  , \g62150/_0_  , \g62151/_0_  , \g62153/_0_  , \g62155/_0_  , \g62156/_0_  , \g62158/_0_  , \g62160/_0_  , \g62161/_0_  , \g62162/_0_  , \g62164/_0_  , \g62165/_0_  , \g62166/_0_  , \g62167/_0_  , \g62168/_0_  , \g62169/_0_  , \g62172/_0_  , \g62173/_0_  , \g62175/_0_  , \g62176/_0_  , \g62177/_0_  , \g62178/_0_  , \g62179/_0_  , \g62180/_0_  , \g62181/_0_  , \g62182/_0_  , \g62183/_0_  , \g62184/_0_  , \g62185/_0_  , \g62186/_0_  , \g62188/_0_  , \g62189/_0_  , \g62190/_0_  , \g62191/_0_  , \g62193/_0_  , \g62194/_0_  , \g62195/_0_  , \g62196/_0_  , \g62197/_0_  , \g62200/_0_  , \g62201/_0_  , \g62202/_0_  , \g62203/_0_  , \g62205/_0_  , \g62206/_0_  , \g62207/_0_  , \g62208/_0_  , \g62209/_0_  , \g62210/_0_  , \g62211/_0_  , \g62215/_0_  , \g62218/_0_  , \g62219/_0_  , \g62221/_0_  , \g62222/_0_  , \g62223/_0_  , \g62224/_0_  , \g62225/_0_  , \g62226/_0_  , \g62229/_0_  , \g62230/_0_  , \g62231/_0_  , \g62233/_0_  , \g62236/_0_  , \g62237/_0_  , \g62238/_0_  , \g62240/_0_  , \g62241/_0_  , \g62243/_0_  , \g62244/_0_  , \g62245/_0_  , \g62247/_0_  , \g62248/_0_  , \g62250/_0_  , \g62252/_0_  , \g62253/_0_  , \g62255/_0_  , \g62256/_0_  , \g62257/_0_  , \g62258/_0_  , \g62259/_0_  , \g62260/_0_  , \g62261/_0_  , \g62262/_0_  , \g62263/_0_  , \g62264/_0_  , \g62265/_0_  , \g62267/_0_  , \g62269/_0_  , \g62270/_0_  , \g62272/_0_  , \g62274/_0_  , \g62277/_0_  , \g62279/_0_  , \g62280/_0_  , \g62281/_0_  , \g62283/_0_  , \g62284/_0_  , \g62285/_0_  , \g62286/_0_  , \g62288/_0_  , \g62289/_0_  , \g62290/_0_  , \g62294/_0_  , \g62295/_0_  , \g62296/_0_  , \g62297/_0_  , \g62298/_0_  , \g62299/_0_  , \g62303/_0_  , \g62305/_0_  , \g62306/_0_  , \g62307/_0_  , \g62309/_0_  , \g62311/_0_  , \g62312/_0_  , \g62313/_0_  , \g62314/_0_  , \g62315/_0_  , \g62316/_0_  , \g62317/_0_  , \g62318/_0_  , \g62319/_0_  , \g62320/_0_  , \g62322/_0_  , \g62324/_0_  , \g62325/_0_  , \g62326/_0_  , \g62327/_0_  , \g62329/_0_  , \g62330/_0_  , \g62331/_0_  , \g62332/_0_  , \g62333/_0_  , \g62335/_0_  , \g62336/_0_  , \g62338/_0_  , \g62341/_0_  , \g62342/_0_  , \g62344/_0_  , \g62345/_0_  , \g62348/_0_  , \g62349/_0_  , \g62350/_0_  , \g62353/_0_  , \g62354/_0_  , \g62355/_0_  , \g62356/_0_  , \g62359/_0_  , \g62362/_0_  , \g62363/_0_  , \g62364/_0_  , \g62365/_0_  , \g62366/_0_  , \g62367/_0_  , \g62368/_0_  , \g62369/_0_  , \g62370/_0_  , \g62371/_0_  , \g62372/_0_  , \g62373/_0_  , \g62374/_0_  , \g62376/_0_  , \g62467/_0_  , \g62468/_0_  , \g62469/_0_  , \g62470/_0_  , \g62471/_0_  , \g62472/_0_  , \g62473/_0_  , \g62474/_0_  , \g62475/_0_  , \g62478/_0_  , \g62480/_0_  , \g62481/_0_  , \g62482/_0_  , \g62483/_0_  , \g62484/_0_  , \g62485/_0_  , \g62486/_0_  , \g62487/_0_  , \g62488/_0_  , \g62489/_0_  , \g62490/_0_  , \g62491/_0_  , \g62492/_0_  , \g62493/_0_  , \g62494/_0_  , \g62495/_0_  , \g62496/_0_  , \g62497/_0_  , \g62498/_0_  , \g62499/_0_  , \g62500/_0_  , \g62501/_0_  , \g62502/_0_  , \g62503/_0_  , \g62504/_0_  , \g62509/_0_  , \g62510/_0_  , \g62511/_0_  , \g62512/_0_  , \g62513/_0_  , \g62514/_0_  , \g62515/_0_  , \g62516/_0_  , \g62517/_0_  , \g62518/_0_  , \g62519/_0_  , \g62520/_0_  , \g62521/_0_  , \g62523/_0_  , \g62526/_0_  , \g62528/_0_  , \g62529/_0_  , \g62531/_0_  , \g62532/_0_  , \g62533/_0_  , \g62534/_0_  , \g62535/_0_  , \g62536/_0_  , \g62537/_0_  , \g62539/_0_  , \g62540/_0_  , \g62541/_0_  , \g62542/_0_  , \g62543/_0_  , \g62544/_0_  , \g62545/_0_  , \g62547/_0_  , \g62548/_0_  , \g62549/_0_  , \g62550/_0_  , \g62551/_0_  , \g62552/_0_  , \g62553/_0_  , \g62554/_0_  , \g62555/_0_  , \g62556/_0_  , \g62557/_0_  , \g62560/_0_  , \g62562/_0_  , \g62563/_0_  , \g62564/_0_  , \g62565/_0_  , \g62566/_0_  , \g62567/_0_  , \g62569/_0_  , \g62570/_0_  , \g62571/_0_  , \g62572/_0_  , \g62573/_0_  , \g62574/_0_  , \g62576/_0_  , \g62577/_0_  , \g62581/_0_  , \g62582/_0_  , \g62584/_0_  , \g62585/_0_  , \g62586/_0_  , \g62588/_0_  , \g62589/_0_  , \g62593/_0_  , \g62594/_0_  , \g62595/_0_  , \g62596/_0_  , \g62597/_0_  , \g62598/_0_  , \g62599/_0_  , \g62600/_0_  , \g62601/_0_  , \g62602/_0_  , \g62603/_0_  , \g62604/_0_  , \g62605/_0_  , \g62606/_0_  , \g62607/_0_  , \g62608/_0_  , \g62609/_0_  , \g62610/_0_  , \g62612/_0_  , \g62613/_0_  , \g62614/_0_  , \g62615/_0_  , \g62617/_0_  , \g62618/_0_  , \g62620/_0_  , \g62621/_0_  , \g62622/_0_  , \g62624/_0_  , \g62625/_0_  , \g62626/_0_  , \g62627/_0_  , \g62629/_0_  , \g62630/_0_  , \g62632/_0_  , \g62633/_0_  , \g62635/_0_  , \g62636/_0_  , \g62637/_0_  , \g62638/_0_  , \g62640/_0_  , \g62641/_0_  , \g62642/_0_  , \g62643/_0_  , \g62644/_0_  , \g62646/_0_  , \g62647/_0_  , \g62649/_0_  , \g62650/_0_  , \g62651/_0_  , \g62653/_0_  , \g62655/_0_  , \g62656/_0_  , \g62657/_0_  , \g62658/_0_  , \g62660/_0_  , \g62661/_0_  , \g62662/_0_  , \g62663/_0_  , \g62664/_0_  , \g62665/_0_  , \g62667/_0_  , \g62669/_0_  , \g62670/_0_  , \g62671/_0_  , \g62672/_0_  , \g62674/_0_  , \g62675/_0_  , \g62676/_0_  , \g62677/_0_  , \g62678/_0_  , \g62679/_0_  , \g62680/_0_  , \g62681/_0_  , \g62682/_0_  , \g62684/_0_  , \g62685/_0_  , \g62686/_0_  , \g62687/_0_  , \g62690/_0_  , \g62693/_0_  , \g62698/_0_  , \g62699/_0_  , \g62700/_0_  , \g62701/_0_  , \g62702/_0_  , \g62703/_0_  , \g62704/_0_  , \g62709/_0_  , \g62710/_0_  , \g62711/_0_  , \g62714/_0_  , \g62715/_0_  , \g62717/_0_  , \g62718/_0_  , \g62719/_0_  , \g62720/_0_  , \g62721/_0_  , \g62723/_0_  , \g62725/_0_  , \g62726/_0_  , \g62729/_0_  , \g62731/_0_  , \g62733/_0_  , \g62738/_0_  , \g62741/_0_  , \g62742/_0_  , \g62744/_0_  , \g62745/_0_  , \g62746/_0_  , \g62747/_0_  , \g62748/_0_  , \g62749/_0_  , \g62753/_0_  , \g62755/_0_  , \g62756/_0_  , \g62758/_0_  , \g62759/_0_  , \g62760/_0_  , \g62761/_0_  , \g62763/_0_  , \g62766/_0_  , \g62767/_0_  , \g62768/_0_  , \g65554/_0_  , \g65561/_0_  , \g65569/_0_  , \g65580/_0_  , \g65599/_0_  , \g65606/_0_  , \g65636/_0_  , \g65864/_0_  );
  input \DATA_0_0_pad  ;
  input \DATA_0_10_pad  ;
  input \DATA_0_11_pad  ;
  input \DATA_0_12_pad  ;
  input \DATA_0_13_pad  ;
  input \DATA_0_14_pad  ;
  input \DATA_0_15_pad  ;
  input \DATA_0_16_pad  ;
  input \DATA_0_17_pad  ;
  input \DATA_0_18_pad  ;
  input \DATA_0_19_pad  ;
  input \DATA_0_1_pad  ;
  input \DATA_0_20_pad  ;
  input \DATA_0_21_pad  ;
  input \DATA_0_22_pad  ;
  input \DATA_0_23_pad  ;
  input \DATA_0_24_pad  ;
  input \DATA_0_25_pad  ;
  input \DATA_0_26_pad  ;
  input \DATA_0_27_pad  ;
  input \DATA_0_28_pad  ;
  input \DATA_0_29_pad  ;
  input \DATA_0_2_pad  ;
  input \DATA_0_30_pad  ;
  input \DATA_0_31_pad  ;
  input \DATA_0_3_pad  ;
  input \DATA_0_4_pad  ;
  input \DATA_0_5_pad  ;
  input \DATA_0_6_pad  ;
  input \DATA_0_7_pad  ;
  input \DATA_0_8_pad  ;
  input \DATA_0_9_pad  ;
  input RESET_pad ;
  input \TM0_pad  ;
  input \TM1_pad  ;
  input \WX10829_reg/NET0131  ;
  input \WX10831_reg/NET0131  ;
  input \WX10833_reg/NET0131  ;
  input \WX10835_reg/NET0131  ;
  input \WX10837_reg/NET0131  ;
  input \WX10839_reg/NET0131  ;
  input \WX10841_reg/NET0131  ;
  input \WX10843_reg/NET0131  ;
  input \WX10845_reg/NET0131  ;
  input \WX10847_reg/NET0131  ;
  input \WX10849_reg/NET0131  ;
  input \WX10851_reg/NET0131  ;
  input \WX10853_reg/NET0131  ;
  input \WX10855_reg/NET0131  ;
  input \WX10857_reg/NET0131  ;
  input \WX10859_reg/NET0131  ;
  input \WX10861_reg/NET0131  ;
  input \WX10863_reg/NET0131  ;
  input \WX10865_reg/NET0131  ;
  input \WX10867_reg/NET0131  ;
  input \WX10869_reg/NET0131  ;
  input \WX10871_reg/NET0131  ;
  input \WX10873_reg/NET0131  ;
  input \WX10875_reg/NET0131  ;
  input \WX10877_reg/NET0131  ;
  input \WX10879_reg/NET0131  ;
  input \WX10881_reg/NET0131  ;
  input \WX10883_reg/NET0131  ;
  input \WX10885_reg/NET0131  ;
  input \WX10887_reg/NET0131  ;
  input \WX10889_reg/NET0131  ;
  input \WX10891_reg/NET0131  ;
  input \WX10989_reg/NET0131  ;
  input \WX10991_reg/NET0131  ;
  input \WX10993_reg/NET0131  ;
  input \WX10995_reg/NET0131  ;
  input \WX10997_reg/NET0131  ;
  input \WX10999_reg/NET0131  ;
  input \WX11001_reg/NET0131  ;
  input \WX11003_reg/NET0131  ;
  input \WX11005_reg/NET0131  ;
  input \WX11007_reg/NET0131  ;
  input \WX11009_reg/NET0131  ;
  input \WX11011_reg/NET0131  ;
  input \WX11013_reg/NET0131  ;
  input \WX11015_reg/NET0131  ;
  input \WX11017_reg/NET0131  ;
  input \WX11019_reg/NET0131  ;
  input \WX11021_reg/NET0131  ;
  input \WX11023_reg/NET0131  ;
  input \WX11025_reg/NET0131  ;
  input \WX11027_reg/NET0131  ;
  input \WX11029_reg/NET0131  ;
  input \WX11031_reg/NET0131  ;
  input \WX11033_reg/NET0131  ;
  input \WX11035_reg/NET0131  ;
  input \WX11037_reg/NET0131  ;
  input \WX11039_reg/NET0131  ;
  input \WX11041_reg/NET0131  ;
  input \WX11043_reg/NET0131  ;
  input \WX11045_reg/NET0131  ;
  input \WX11047_reg/NET0131  ;
  input \WX11049_reg/NET0131  ;
  input \WX11051_reg/NET0131  ;
  input \WX11053_reg/NET0131  ;
  input \WX11055_reg/NET0131  ;
  input \WX11057_reg/NET0131  ;
  input \WX11059_reg/NET0131  ;
  input \WX11061_reg/NET0131  ;
  input \WX11063_reg/NET0131  ;
  input \WX11065_reg/NET0131  ;
  input \WX11067_reg/NET0131  ;
  input \WX11069_reg/NET0131  ;
  input \WX11071_reg/NET0131  ;
  input \WX11073_reg/NET0131  ;
  input \WX11075_reg/NET0131  ;
  input \WX11077_reg/NET0131  ;
  input \WX11079_reg/NET0131  ;
  input \WX11081_reg/NET0131  ;
  input \WX11083_reg/NET0131  ;
  input \WX11085_reg/NET0131  ;
  input \WX11087_reg/NET0131  ;
  input \WX11089_reg/NET0131  ;
  input \WX11091_reg/NET0131  ;
  input \WX11093_reg/NET0131  ;
  input \WX11095_reg/NET0131  ;
  input \WX11097_reg/NET0131  ;
  input \WX11099_reg/NET0131  ;
  input \WX11101_reg/NET0131  ;
  input \WX11103_reg/NET0131  ;
  input \WX11105_reg/NET0131  ;
  input \WX11107_reg/NET0131  ;
  input \WX11109_reg/NET0131  ;
  input \WX11111_reg/NET0131  ;
  input \WX11113_reg/NET0131  ;
  input \WX11115_reg/NET0131  ;
  input \WX11117_reg/NET0131  ;
  input \WX11119_reg/NET0131  ;
  input \WX11121_reg/NET0131  ;
  input \WX11123_reg/NET0131  ;
  input \WX11125_reg/NET0131  ;
  input \WX11127_reg/NET0131  ;
  input \WX11129_reg/NET0131  ;
  input \WX11131_reg/NET0131  ;
  input \WX11133_reg/NET0131  ;
  input \WX11135_reg/NET0131  ;
  input \WX11137_reg/NET0131  ;
  input \WX11139_reg/NET0131  ;
  input \WX11141_reg/NET0131  ;
  input \WX11143_reg/NET0131  ;
  input \WX11145_reg/NET0131  ;
  input \WX11147_reg/NET0131  ;
  input \WX11149_reg/NET0131  ;
  input \WX11151_reg/NET0131  ;
  input \WX11153_reg/NET0131  ;
  input \WX11155_reg/NET0131  ;
  input \WX11157_reg/NET0131  ;
  input \WX11159_reg/NET0131  ;
  input \WX11161_reg/NET0131  ;
  input \WX11163_reg/NET0131  ;
  input \WX11165_reg/NET0131  ;
  input \WX11167_reg/NET0131  ;
  input \WX11169_reg/NET0131  ;
  input \WX11171_reg/NET0131  ;
  input \WX11173_reg/NET0131  ;
  input \WX11175_reg/NET0131  ;
  input \WX11177_reg/NET0131  ;
  input \WX11179_reg/NET0131  ;
  input \WX11181_reg/NET0131  ;
  input \WX11183_reg/NET0131  ;
  input \WX11185_reg/NET0131  ;
  input \WX11187_reg/NET0131  ;
  input \WX11189_reg/NET0131  ;
  input \WX11191_reg/NET0131  ;
  input \WX11193_reg/NET0131  ;
  input \WX11195_reg/NET0131  ;
  input \WX11197_reg/NET0131  ;
  input \WX11199_reg/NET0131  ;
  input \WX11201_reg/NET0131  ;
  input \WX11203_reg/NET0131  ;
  input \WX11205_reg/NET0131  ;
  input \WX11207_reg/NET0131  ;
  input \WX11209_reg/NET0131  ;
  input \WX11211_reg/NET0131  ;
  input \WX11213_reg/NET0131  ;
  input \WX11215_reg/NET0131  ;
  input \WX11217_reg/NET0131  ;
  input \WX11219_reg/NET0131  ;
  input \WX11221_reg/NET0131  ;
  input \WX11223_reg/NET0131  ;
  input \WX11225_reg/NET0131  ;
  input \WX11227_reg/NET0131  ;
  input \WX11229_reg/NET0131  ;
  input \WX11231_reg/NET0131  ;
  input \WX11233_reg/NET0131  ;
  input \WX11235_reg/NET0131  ;
  input \WX11237_reg/NET0131  ;
  input \WX11239_reg/NET0131  ;
  input \WX11241_reg/NET0131  ;
  input \WX11243_reg/NET0131  ;
  input \WX1938_reg/NET0131  ;
  input \WX1940_reg/NET0131  ;
  input \WX1942_reg/NET0131  ;
  input \WX1944_reg/NET0131  ;
  input \WX1946_reg/NET0131  ;
  input \WX1948_reg/NET0131  ;
  input \WX1950_reg/NET0131  ;
  input \WX1952_reg/NET0131  ;
  input \WX1954_reg/NET0131  ;
  input \WX1956_reg/NET0131  ;
  input \WX1958_reg/NET0131  ;
  input \WX1960_reg/NET0131  ;
  input \WX1962_reg/NET0131  ;
  input \WX1964_reg/NET0131  ;
  input \WX1966_reg/NET0131  ;
  input \WX1968_reg/NET0131  ;
  input \WX1970_reg/NET0131  ;
  input \WX1972_reg/NET0131  ;
  input \WX1974_reg/NET0131  ;
  input \WX1976_reg/NET0131  ;
  input \WX1978_reg/NET0131  ;
  input \WX1980_reg/NET0131  ;
  input \WX1982_reg/NET0131  ;
  input \WX1984_reg/NET0131  ;
  input \WX1986_reg/NET0131  ;
  input \WX1988_reg/NET0131  ;
  input \WX1990_reg/NET0131  ;
  input \WX1992_reg/NET0131  ;
  input \WX1994_reg/NET0131  ;
  input \WX1996_reg/NET0131  ;
  input \WX1998_reg/NET0131  ;
  input \WX2000_reg/NET0131  ;
  input \WX2002_reg/NET0131  ;
  input \WX2004_reg/NET0131  ;
  input \WX2006_reg/NET0131  ;
  input \WX2008_reg/NET0131  ;
  input \WX2010_reg/NET0131  ;
  input \WX2012_reg/NET0131  ;
  input \WX2014_reg/NET0131  ;
  input \WX2016_reg/NET0131  ;
  input \WX2018_reg/NET0131  ;
  input \WX2020_reg/NET0131  ;
  input \WX2022_reg/NET0131  ;
  input \WX2024_reg/NET0131  ;
  input \WX2026_reg/NET0131  ;
  input \WX2028_reg/NET0131  ;
  input \WX2030_reg/NET0131  ;
  input \WX2032_reg/NET0131  ;
  input \WX2034_reg/NET0131  ;
  input \WX2036_reg/NET0131  ;
  input \WX2038_reg/NET0131  ;
  input \WX2040_reg/NET0131  ;
  input \WX2042_reg/NET0131  ;
  input \WX2044_reg/NET0131  ;
  input \WX2046_reg/NET0131  ;
  input \WX2048_reg/NET0131  ;
  input \WX2050_reg/NET0131  ;
  input \WX2052_reg/NET0131  ;
  input \WX2054_reg/NET0131  ;
  input \WX2056_reg/NET0131  ;
  input \WX2058_reg/NET0131  ;
  input \WX2060_reg/NET0131  ;
  input \WX2062_reg/NET0131  ;
  input \WX2064_reg/NET0131  ;
  input \WX2066_reg/NET0131  ;
  input \WX2068_reg/NET0131  ;
  input \WX2070_reg/NET0131  ;
  input \WX2072_reg/NET0131  ;
  input \WX2074_reg/NET0131  ;
  input \WX2076_reg/NET0131  ;
  input \WX2078_reg/NET0131  ;
  input \WX2080_reg/NET0131  ;
  input \WX2082_reg/NET0131  ;
  input \WX2084_reg/NET0131  ;
  input \WX2086_reg/NET0131  ;
  input \WX2088_reg/NET0131  ;
  input \WX2090_reg/NET0131  ;
  input \WX2092_reg/NET0131  ;
  input \WX2094_reg/NET0131  ;
  input \WX2096_reg/NET0131  ;
  input \WX2098_reg/NET0131  ;
  input \WX2100_reg/NET0131  ;
  input \WX2102_reg/NET0131  ;
  input \WX2104_reg/NET0131  ;
  input \WX2106_reg/NET0131  ;
  input \WX2108_reg/NET0131  ;
  input \WX2110_reg/NET0131  ;
  input \WX2112_reg/NET0131  ;
  input \WX2114_reg/NET0131  ;
  input \WX2116_reg/NET0131  ;
  input \WX2118_reg/NET0131  ;
  input \WX2120_reg/NET0131  ;
  input \WX2122_reg/NET0131  ;
  input \WX2124_reg/NET0131  ;
  input \WX2126_reg/NET0131  ;
  input \WX2128_reg/NET0131  ;
  input \WX2130_reg/NET0131  ;
  input \WX2132_reg/NET0131  ;
  input \WX2134_reg/NET0131  ;
  input \WX2136_reg/NET0131  ;
  input \WX2138_reg/NET0131  ;
  input \WX2140_reg/NET0131  ;
  input \WX2142_reg/NET0131  ;
  input \WX2144_reg/NET0131  ;
  input \WX2146_reg/NET0131  ;
  input \WX2148_reg/NET0131  ;
  input \WX2150_reg/NET0131  ;
  input \WX2152_reg/NET0131  ;
  input \WX2154_reg/NET0131  ;
  input \WX2156_reg/NET0131  ;
  input \WX2158_reg/NET0131  ;
  input \WX2160_reg/NET0131  ;
  input \WX2162_reg/NET0131  ;
  input \WX2164_reg/NET0131  ;
  input \WX2166_reg/NET0131  ;
  input \WX2168_reg/NET0131  ;
  input \WX2170_reg/NET0131  ;
  input \WX2172_reg/NET0131  ;
  input \WX2174_reg/NET0131  ;
  input \WX2176_reg/NET0131  ;
  input \WX2178_reg/NET0131  ;
  input \WX2180_reg/NET0131  ;
  input \WX2182_reg/NET0131  ;
  input \WX2184_reg/NET0131  ;
  input \WX2186_reg/NET0131  ;
  input \WX2188_reg/NET0131  ;
  input \WX2190_reg/NET0131  ;
  input \WX2192_reg/NET0131  ;
  input \WX3231_reg/NET0131  ;
  input \WX3233_reg/NET0131  ;
  input \WX3235_reg/NET0131  ;
  input \WX3237_reg/NET0131  ;
  input \WX3239_reg/NET0131  ;
  input \WX3241_reg/NET0131  ;
  input \WX3243_reg/NET0131  ;
  input \WX3245_reg/NET0131  ;
  input \WX3247_reg/NET0131  ;
  input \WX3249_reg/NET0131  ;
  input \WX3251_reg/NET0131  ;
  input \WX3253_reg/NET0131  ;
  input \WX3255_reg/NET0131  ;
  input \WX3257_reg/NET0131  ;
  input \WX3259_reg/NET0131  ;
  input \WX3261_reg/NET0131  ;
  input \WX3263_reg/NET0131  ;
  input \WX3265_reg/NET0131  ;
  input \WX3267_reg/NET0131  ;
  input \WX3269_reg/NET0131  ;
  input \WX3271_reg/NET0131  ;
  input \WX3273_reg/NET0131  ;
  input \WX3275_reg/NET0131  ;
  input \WX3277_reg/NET0131  ;
  input \WX3279_reg/NET0131  ;
  input \WX3281_reg/NET0131  ;
  input \WX3283_reg/NET0131  ;
  input \WX3285_reg/NET0131  ;
  input \WX3287_reg/NET0131  ;
  input \WX3289_reg/NET0131  ;
  input \WX3291_reg/NET0131  ;
  input \WX3293_reg/NET0131  ;
  input \WX3295_reg/NET0131  ;
  input \WX3297_reg/NET0131  ;
  input \WX3299_reg/NET0131  ;
  input \WX3301_reg/NET0131  ;
  input \WX3303_reg/NET0131  ;
  input \WX3305_reg/NET0131  ;
  input \WX3307_reg/NET0131  ;
  input \WX3309_reg/NET0131  ;
  input \WX3311_reg/NET0131  ;
  input \WX3313_reg/NET0131  ;
  input \WX3315_reg/NET0131  ;
  input \WX3317_reg/NET0131  ;
  input \WX3319_reg/NET0131  ;
  input \WX3321_reg/NET0131  ;
  input \WX3323_reg/NET0131  ;
  input \WX3325_reg/NET0131  ;
  input \WX3327_reg/NET0131  ;
  input \WX3329_reg/NET0131  ;
  input \WX3331_reg/NET0131  ;
  input \WX3333_reg/NET0131  ;
  input \WX3335_reg/NET0131  ;
  input \WX3337_reg/NET0131  ;
  input \WX3339_reg/NET0131  ;
  input \WX3341_reg/NET0131  ;
  input \WX3343_reg/NET0131  ;
  input \WX3345_reg/NET0131  ;
  input \WX3347_reg/NET0131  ;
  input \WX3349_reg/NET0131  ;
  input \WX3351_reg/NET0131  ;
  input \WX3353_reg/NET0131  ;
  input \WX3355_reg/NET0131  ;
  input \WX3357_reg/NET0131  ;
  input \WX3359_reg/NET0131  ;
  input \WX3361_reg/NET0131  ;
  input \WX3363_reg/NET0131  ;
  input \WX3365_reg/NET0131  ;
  input \WX3367_reg/NET0131  ;
  input \WX3369_reg/NET0131  ;
  input \WX3371_reg/NET0131  ;
  input \WX3373_reg/NET0131  ;
  input \WX3375_reg/NET0131  ;
  input \WX3377_reg/NET0131  ;
  input \WX3379_reg/NET0131  ;
  input \WX3381_reg/NET0131  ;
  input \WX3383_reg/NET0131  ;
  input \WX3385_reg/NET0131  ;
  input \WX3387_reg/NET0131  ;
  input \WX3389_reg/NET0131  ;
  input \WX3391_reg/NET0131  ;
  input \WX3393_reg/NET0131  ;
  input \WX3395_reg/NET0131  ;
  input \WX3397_reg/NET0131  ;
  input \WX3399_reg/NET0131  ;
  input \WX3401_reg/NET0131  ;
  input \WX3403_reg/NET0131  ;
  input \WX3405_reg/NET0131  ;
  input \WX3407_reg/NET0131  ;
  input \WX3409_reg/NET0131  ;
  input \WX3411_reg/NET0131  ;
  input \WX3413_reg/NET0131  ;
  input \WX3415_reg/NET0131  ;
  input \WX3417_reg/NET0131  ;
  input \WX3419_reg/NET0131  ;
  input \WX3421_reg/NET0131  ;
  input \WX3423_reg/NET0131  ;
  input \WX3425_reg/NET0131  ;
  input \WX3427_reg/NET0131  ;
  input \WX3429_reg/NET0131  ;
  input \WX3431_reg/NET0131  ;
  input \WX3433_reg/NET0131  ;
  input \WX3435_reg/NET0131  ;
  input \WX3437_reg/NET0131  ;
  input \WX3439_reg/NET0131  ;
  input \WX3441_reg/NET0131  ;
  input \WX3443_reg/NET0131  ;
  input \WX3445_reg/NET0131  ;
  input \WX3447_reg/NET0131  ;
  input \WX3449_reg/NET0131  ;
  input \WX3451_reg/NET0131  ;
  input \WX3453_reg/NET0131  ;
  input \WX3455_reg/NET0131  ;
  input \WX3457_reg/NET0131  ;
  input \WX3459_reg/NET0131  ;
  input \WX3461_reg/NET0131  ;
  input \WX3463_reg/NET0131  ;
  input \WX3465_reg/NET0131  ;
  input \WX3467_reg/NET0131  ;
  input \WX3469_reg/NET0131  ;
  input \WX3471_reg/NET0131  ;
  input \WX3473_reg/NET0131  ;
  input \WX3475_reg/NET0131  ;
  input \WX3477_reg/NET0131  ;
  input \WX3479_reg/NET0131  ;
  input \WX3481_reg/NET0131  ;
  input \WX3483_reg/NET0131  ;
  input \WX3485_reg/NET0131  ;
  input \WX4524_reg/NET0131  ;
  input \WX4526_reg/NET0131  ;
  input \WX4528_reg/NET0131  ;
  input \WX4530_reg/NET0131  ;
  input \WX4532_reg/NET0131  ;
  input \WX4534_reg/NET0131  ;
  input \WX4536_reg/NET0131  ;
  input \WX4538_reg/NET0131  ;
  input \WX4540_reg/NET0131  ;
  input \WX4542_reg/NET0131  ;
  input \WX4544_reg/NET0131  ;
  input \WX4546_reg/NET0131  ;
  input \WX4548_reg/NET0131  ;
  input \WX4550_reg/NET0131  ;
  input \WX4552_reg/NET0131  ;
  input \WX4554_reg/NET0131  ;
  input \WX4556_reg/NET0131  ;
  input \WX4558_reg/NET0131  ;
  input \WX4560_reg/NET0131  ;
  input \WX4562_reg/NET0131  ;
  input \WX4564_reg/NET0131  ;
  input \WX4566_reg/NET0131  ;
  input \WX4568_reg/NET0131  ;
  input \WX4570_reg/NET0131  ;
  input \WX4572_reg/NET0131  ;
  input \WX4574_reg/NET0131  ;
  input \WX4576_reg/NET0131  ;
  input \WX4578_reg/NET0131  ;
  input \WX4580_reg/NET0131  ;
  input \WX4582_reg/NET0131  ;
  input \WX4584_reg/NET0131  ;
  input \WX4586_reg/NET0131  ;
  input \WX4588_reg/NET0131  ;
  input \WX4590_reg/NET0131  ;
  input \WX4592_reg/NET0131  ;
  input \WX4594_reg/NET0131  ;
  input \WX4596_reg/NET0131  ;
  input \WX4598_reg/NET0131  ;
  input \WX4600_reg/NET0131  ;
  input \WX4602_reg/NET0131  ;
  input \WX4604_reg/NET0131  ;
  input \WX4606_reg/NET0131  ;
  input \WX4608_reg/NET0131  ;
  input \WX4610_reg/NET0131  ;
  input \WX4612_reg/NET0131  ;
  input \WX4614_reg/NET0131  ;
  input \WX4616_reg/NET0131  ;
  input \WX4618_reg/NET0131  ;
  input \WX4620_reg/NET0131  ;
  input \WX4622_reg/NET0131  ;
  input \WX4624_reg/NET0131  ;
  input \WX4626_reg/NET0131  ;
  input \WX4628_reg/NET0131  ;
  input \WX4630_reg/NET0131  ;
  input \WX4632_reg/NET0131  ;
  input \WX4634_reg/NET0131  ;
  input \WX4636_reg/NET0131  ;
  input \WX4638_reg/NET0131  ;
  input \WX4640_reg/NET0131  ;
  input \WX4642_reg/NET0131  ;
  input \WX4644_reg/NET0131  ;
  input \WX4646_reg/NET0131  ;
  input \WX4648_reg/NET0131  ;
  input \WX4650_reg/NET0131  ;
  input \WX4652_reg/NET0131  ;
  input \WX4654_reg/NET0131  ;
  input \WX4656_reg/NET0131  ;
  input \WX4658_reg/NET0131  ;
  input \WX4660_reg/NET0131  ;
  input \WX4662_reg/NET0131  ;
  input \WX4664_reg/NET0131  ;
  input \WX4666_reg/NET0131  ;
  input \WX4668_reg/NET0131  ;
  input \WX4670_reg/NET0131  ;
  input \WX4672_reg/NET0131  ;
  input \WX4674_reg/NET0131  ;
  input \WX4676_reg/NET0131  ;
  input \WX4678_reg/NET0131  ;
  input \WX4680_reg/NET0131  ;
  input \WX4682_reg/NET0131  ;
  input \WX4684_reg/NET0131  ;
  input \WX4686_reg/NET0131  ;
  input \WX4688_reg/NET0131  ;
  input \WX4690_reg/NET0131  ;
  input \WX4692_reg/NET0131  ;
  input \WX4694_reg/NET0131  ;
  input \WX4696_reg/NET0131  ;
  input \WX4698_reg/NET0131  ;
  input \WX4700_reg/NET0131  ;
  input \WX4702_reg/NET0131  ;
  input \WX4704_reg/NET0131  ;
  input \WX4706_reg/NET0131  ;
  input \WX4708_reg/NET0131  ;
  input \WX4710_reg/NET0131  ;
  input \WX4712_reg/NET0131  ;
  input \WX4714_reg/NET0131  ;
  input \WX4716_reg/NET0131  ;
  input \WX4718_reg/NET0131  ;
  input \WX4720_reg/NET0131  ;
  input \WX4722_reg/NET0131  ;
  input \WX4724_reg/NET0131  ;
  input \WX4726_reg/NET0131  ;
  input \WX4728_reg/NET0131  ;
  input \WX4730_reg/NET0131  ;
  input \WX4732_reg/NET0131  ;
  input \WX4734_reg/NET0131  ;
  input \WX4736_reg/NET0131  ;
  input \WX4738_reg/NET0131  ;
  input \WX4740_reg/NET0131  ;
  input \WX4742_reg/NET0131  ;
  input \WX4744_reg/NET0131  ;
  input \WX4746_reg/NET0131  ;
  input \WX4748_reg/NET0131  ;
  input \WX4750_reg/NET0131  ;
  input \WX4752_reg/NET0131  ;
  input \WX4754_reg/NET0131  ;
  input \WX4756_reg/NET0131  ;
  input \WX4758_reg/NET0131  ;
  input \WX4760_reg/NET0131  ;
  input \WX4762_reg/NET0131  ;
  input \WX4764_reg/NET0131  ;
  input \WX4766_reg/NET0131  ;
  input \WX4768_reg/NET0131  ;
  input \WX4770_reg/NET0131  ;
  input \WX4772_reg/NET0131  ;
  input \WX4774_reg/NET0131  ;
  input \WX4776_reg/NET0131  ;
  input \WX4778_reg/NET0131  ;
  input \WX5817_reg/NET0131  ;
  input \WX5819_reg/NET0131  ;
  input \WX5821_reg/NET0131  ;
  input \WX5823_reg/NET0131  ;
  input \WX5825_reg/NET0131  ;
  input \WX5827_reg/NET0131  ;
  input \WX5829_reg/NET0131  ;
  input \WX5831_reg/NET0131  ;
  input \WX5833_reg/NET0131  ;
  input \WX5835_reg/NET0131  ;
  input \WX5837_reg/NET0131  ;
  input \WX5839_reg/NET0131  ;
  input \WX5841_reg/NET0131  ;
  input \WX5843_reg/NET0131  ;
  input \WX5845_reg/NET0131  ;
  input \WX5847_reg/NET0131  ;
  input \WX5849_reg/NET0131  ;
  input \WX5851_reg/NET0131  ;
  input \WX5853_reg/NET0131  ;
  input \WX5855_reg/NET0131  ;
  input \WX5857_reg/NET0131  ;
  input \WX5859_reg/NET0131  ;
  input \WX5861_reg/NET0131  ;
  input \WX5863_reg/NET0131  ;
  input \WX5865_reg/NET0131  ;
  input \WX5867_reg/NET0131  ;
  input \WX5869_reg/NET0131  ;
  input \WX5871_reg/NET0131  ;
  input \WX5873_reg/NET0131  ;
  input \WX5875_reg/NET0131  ;
  input \WX5877_reg/NET0131  ;
  input \WX5879_reg/NET0131  ;
  input \WX5881_reg/NET0131  ;
  input \WX5883_reg/NET0131  ;
  input \WX5885_reg/NET0131  ;
  input \WX5887_reg/NET0131  ;
  input \WX5889_reg/NET0131  ;
  input \WX5891_reg/NET0131  ;
  input \WX5893_reg/NET0131  ;
  input \WX5895_reg/NET0131  ;
  input \WX5897_reg/NET0131  ;
  input \WX5899_reg/NET0131  ;
  input \WX5901_reg/NET0131  ;
  input \WX5903_reg/NET0131  ;
  input \WX5905_reg/NET0131  ;
  input \WX5907_reg/NET0131  ;
  input \WX5909_reg/NET0131  ;
  input \WX5911_reg/NET0131  ;
  input \WX5913_reg/NET0131  ;
  input \WX5915_reg/NET0131  ;
  input \WX5917_reg/NET0131  ;
  input \WX5919_reg/NET0131  ;
  input \WX5921_reg/NET0131  ;
  input \WX5923_reg/NET0131  ;
  input \WX5925_reg/NET0131  ;
  input \WX5927_reg/NET0131  ;
  input \WX5929_reg/NET0131  ;
  input \WX5931_reg/NET0131  ;
  input \WX5933_reg/NET0131  ;
  input \WX5935_reg/NET0131  ;
  input \WX5937_reg/NET0131  ;
  input \WX5939_reg/NET0131  ;
  input \WX5941_reg/NET0131  ;
  input \WX5943_reg/NET0131  ;
  input \WX5945_reg/NET0131  ;
  input \WX5947_reg/NET0131  ;
  input \WX5949_reg/NET0131  ;
  input \WX5951_reg/NET0131  ;
  input \WX5953_reg/NET0131  ;
  input \WX5955_reg/NET0131  ;
  input \WX5957_reg/NET0131  ;
  input \WX5959_reg/NET0131  ;
  input \WX5961_reg/NET0131  ;
  input \WX5963_reg/NET0131  ;
  input \WX5965_reg/NET0131  ;
  input \WX5967_reg/NET0131  ;
  input \WX5969_reg/NET0131  ;
  input \WX5971_reg/NET0131  ;
  input \WX5973_reg/NET0131  ;
  input \WX5975_reg/NET0131  ;
  input \WX5977_reg/NET0131  ;
  input \WX5979_reg/NET0131  ;
  input \WX5981_reg/NET0131  ;
  input \WX5983_reg/NET0131  ;
  input \WX5985_reg/NET0131  ;
  input \WX5987_reg/NET0131  ;
  input \WX5989_reg/NET0131  ;
  input \WX5991_reg/NET0131  ;
  input \WX5993_reg/NET0131  ;
  input \WX5995_reg/NET0131  ;
  input \WX5997_reg/NET0131  ;
  input \WX5999_reg/NET0131  ;
  input \WX6001_reg/NET0131  ;
  input \WX6003_reg/NET0131  ;
  input \WX6005_reg/NET0131  ;
  input \WX6007_reg/NET0131  ;
  input \WX6009_reg/NET0131  ;
  input \WX6011_reg/NET0131  ;
  input \WX6013_reg/NET0131  ;
  input \WX6015_reg/NET0131  ;
  input \WX6017_reg/NET0131  ;
  input \WX6019_reg/NET0131  ;
  input \WX6021_reg/NET0131  ;
  input \WX6023_reg/NET0131  ;
  input \WX6025_reg/NET0131  ;
  input \WX6027_reg/NET0131  ;
  input \WX6029_reg/NET0131  ;
  input \WX6031_reg/NET0131  ;
  input \WX6033_reg/NET0131  ;
  input \WX6035_reg/NET0131  ;
  input \WX6037_reg/NET0131  ;
  input \WX6039_reg/NET0131  ;
  input \WX6041_reg/NET0131  ;
  input \WX6043_reg/NET0131  ;
  input \WX6045_reg/NET0131  ;
  input \WX6047_reg/NET0131  ;
  input \WX6049_reg/NET0131  ;
  input \WX6051_reg/NET0131  ;
  input \WX6053_reg/NET0131  ;
  input \WX6055_reg/NET0131  ;
  input \WX6057_reg/NET0131  ;
  input \WX6059_reg/NET0131  ;
  input \WX6061_reg/NET0131  ;
  input \WX6063_reg/NET0131  ;
  input \WX6065_reg/NET0131  ;
  input \WX6067_reg/NET0131  ;
  input \WX6069_reg/NET0131  ;
  input \WX6071_reg/NET0131  ;
  input \WX645_reg/NET0131  ;
  input \WX647_reg/NET0131  ;
  input \WX649_reg/NET0131  ;
  input \WX651_reg/NET0131  ;
  input \WX653_reg/NET0131  ;
  input \WX655_reg/NET0131  ;
  input \WX657_reg/NET0131  ;
  input \WX659_reg/NET0131  ;
  input \WX661_reg/NET0131  ;
  input \WX663_reg/NET0131  ;
  input \WX665_reg/NET0131  ;
  input \WX667_reg/NET0131  ;
  input \WX669_reg/NET0131  ;
  input \WX671_reg/NET0131  ;
  input \WX673_reg/NET0131  ;
  input \WX675_reg/NET0131  ;
  input \WX677_reg/NET0131  ;
  input \WX679_reg/NET0131  ;
  input \WX681_reg/NET0131  ;
  input \WX683_reg/NET0131  ;
  input \WX685_reg/NET0131  ;
  input \WX687_reg/NET0131  ;
  input \WX689_reg/NET0131  ;
  input \WX691_reg/NET0131  ;
  input \WX693_reg/NET0131  ;
  input \WX695_reg/NET0131  ;
  input \WX697_reg/NET0131  ;
  input \WX699_reg/NET0131  ;
  input \WX701_reg/NET0131  ;
  input \WX703_reg/NET0131  ;
  input \WX705_reg/NET0131  ;
  input \WX707_reg/NET0131  ;
  input \WX709_reg/NET0131  ;
  input \WX7110_reg/NET0131  ;
  input \WX7112_reg/NET0131  ;
  input \WX7114_reg/NET0131  ;
  input \WX7116_reg/NET0131  ;
  input \WX7118_reg/NET0131  ;
  input \WX711_reg/NET0131  ;
  input \WX7120_reg/NET0131  ;
  input \WX7122_reg/NET0131  ;
  input \WX7124_reg/NET0131  ;
  input \WX7126_reg/NET0131  ;
  input \WX7128_reg/NET0131  ;
  input \WX7130_reg/NET0131  ;
  input \WX7132_reg/NET0131  ;
  input \WX7134_reg/NET0131  ;
  input \WX7136_reg/NET0131  ;
  input \WX7138_reg/NET0131  ;
  input \WX713_reg/NET0131  ;
  input \WX7140_reg/NET0131  ;
  input \WX7142_reg/NET0131  ;
  input \WX7144_reg/NET0131  ;
  input \WX7146_reg/NET0131  ;
  input \WX7148_reg/NET0131  ;
  input \WX7150_reg/NET0131  ;
  input \WX7152_reg/NET0131  ;
  input \WX7154_reg/NET0131  ;
  input \WX7156_reg/NET0131  ;
  input \WX7158_reg/NET0131  ;
  input \WX715_reg/NET0131  ;
  input \WX7160_reg/NET0131  ;
  input \WX7162_reg/NET0131  ;
  input \WX7164_reg/NET0131  ;
  input \WX7166_reg/NET0131  ;
  input \WX7168_reg/NET0131  ;
  input \WX7170_reg/NET0131  ;
  input \WX7172_reg/NET0131  ;
  input \WX7174_reg/NET0131  ;
  input \WX7176_reg/NET0131  ;
  input \WX7178_reg/NET0131  ;
  input \WX717_reg/NET0131  ;
  input \WX7180_reg/NET0131  ;
  input \WX7182_reg/NET0131  ;
  input \WX7184_reg/NET0131  ;
  input \WX7186_reg/NET0131  ;
  input \WX7188_reg/NET0131  ;
  input \WX7190_reg/NET0131  ;
  input \WX7192_reg/NET0131  ;
  input \WX7194_reg/NET0131  ;
  input \WX7196_reg/NET0131  ;
  input \WX7198_reg/NET0131  ;
  input \WX719_reg/NET0131  ;
  input \WX7200_reg/NET0131  ;
  input \WX7202_reg/NET0131  ;
  input \WX7204_reg/NET0131  ;
  input \WX7206_reg/NET0131  ;
  input \WX7208_reg/NET0131  ;
  input \WX7210_reg/NET0131  ;
  input \WX7212_reg/NET0131  ;
  input \WX7214_reg/NET0131  ;
  input \WX7216_reg/NET0131  ;
  input \WX7218_reg/NET0131  ;
  input \WX721_reg/NET0131  ;
  input \WX7220_reg/NET0131  ;
  input \WX7222_reg/NET0131  ;
  input \WX7224_reg/NET0131  ;
  input \WX7226_reg/NET0131  ;
  input \WX7228_reg/NET0131  ;
  input \WX7230_reg/NET0131  ;
  input \WX7232_reg/NET0131  ;
  input \WX7234_reg/NET0131  ;
  input \WX7236_reg/NET0131  ;
  input \WX7238_reg/NET0131  ;
  input \WX723_reg/NET0131  ;
  input \WX7240_reg/NET0131  ;
  input \WX7242_reg/NET0131  ;
  input \WX7244_reg/NET0131  ;
  input \WX7246_reg/NET0131  ;
  input \WX7248_reg/NET0131  ;
  input \WX7250_reg/NET0131  ;
  input \WX7252_reg/NET0131  ;
  input \WX7254_reg/NET0131  ;
  input \WX7256_reg/NET0131  ;
  input \WX7258_reg/NET0131  ;
  input \WX725_reg/NET0131  ;
  input \WX7260_reg/NET0131  ;
  input \WX7262_reg/NET0131  ;
  input \WX7264_reg/NET0131  ;
  input \WX7266_reg/NET0131  ;
  input \WX7268_reg/NET0131  ;
  input \WX7270_reg/NET0131  ;
  input \WX7272_reg/NET0131  ;
  input \WX7274_reg/NET0131  ;
  input \WX7276_reg/NET0131  ;
  input \WX7278_reg/NET0131  ;
  input \WX727_reg/NET0131  ;
  input \WX7280_reg/NET0131  ;
  input \WX7282_reg/NET0131  ;
  input \WX7284_reg/NET0131  ;
  input \WX7286_reg/NET0131  ;
  input \WX7288_reg/NET0131  ;
  input \WX7290_reg/NET0131  ;
  input \WX7292_reg/NET0131  ;
  input \WX7294_reg/NET0131  ;
  input \WX7296_reg/NET0131  ;
  input \WX7298_reg/NET0131  ;
  input \WX729_reg/NET0131  ;
  input \WX7300_reg/NET0131  ;
  input \WX7302_reg/NET0131  ;
  input \WX7304_reg/NET0131  ;
  input \WX7306_reg/NET0131  ;
  input \WX7308_reg/NET0131  ;
  input \WX7310_reg/NET0131  ;
  input \WX7312_reg/NET0131  ;
  input \WX7314_reg/NET0131  ;
  input \WX7316_reg/NET0131  ;
  input \WX7318_reg/NET0131  ;
  input \WX731_reg/NET0131  ;
  input \WX7320_reg/NET0131  ;
  input \WX7322_reg/NET0131  ;
  input \WX7324_reg/NET0131  ;
  input \WX7326_reg/NET0131  ;
  input \WX7328_reg/NET0131  ;
  input \WX7330_reg/NET0131  ;
  input \WX7332_reg/NET0131  ;
  input \WX7334_reg/NET0131  ;
  input \WX7336_reg/NET0131  ;
  input \WX7338_reg/NET0131  ;
  input \WX733_reg/NET0131  ;
  input \WX7340_reg/NET0131  ;
  input \WX7342_reg/NET0131  ;
  input \WX7344_reg/NET0131  ;
  input \WX7346_reg/NET0131  ;
  input \WX7348_reg/NET0131  ;
  input \WX7350_reg/NET0131  ;
  input \WX7352_reg/NET0131  ;
  input \WX7354_reg/NET0131  ;
  input \WX7356_reg/NET0131  ;
  input \WX7358_reg/NET0131  ;
  input \WX735_reg/NET0131  ;
  input \WX7360_reg/NET0131  ;
  input \WX7362_reg/NET0131  ;
  input \WX7364_reg/NET0131  ;
  input \WX737_reg/NET0131  ;
  input \WX739_reg/NET0131  ;
  input \WX741_reg/NET0131  ;
  input \WX743_reg/NET0131  ;
  input \WX745_reg/NET0131  ;
  input \WX747_reg/NET0131  ;
  input \WX749_reg/NET0131  ;
  input \WX751_reg/NET0131  ;
  input \WX753_reg/NET0131  ;
  input \WX755_reg/NET0131  ;
  input \WX757_reg/NET0131  ;
  input \WX759_reg/NET0131  ;
  input \WX761_reg/NET0131  ;
  input \WX763_reg/NET0131  ;
  input \WX765_reg/NET0131  ;
  input \WX767_reg/NET0131  ;
  input \WX769_reg/NET0131  ;
  input \WX771_reg/NET0131  ;
  input \WX773_reg/NET0131  ;
  input \WX775_reg/NET0131  ;
  input \WX777_reg/NET0131  ;
  input \WX779_reg/NET0131  ;
  input \WX781_reg/NET0131  ;
  input \WX783_reg/NET0131  ;
  input \WX785_reg/NET0131  ;
  input \WX787_reg/NET0131  ;
  input \WX789_reg/NET0131  ;
  input \WX791_reg/NET0131  ;
  input \WX793_reg/NET0131  ;
  input \WX795_reg/NET0131  ;
  input \WX797_reg/NET0131  ;
  input \WX799_reg/NET0131  ;
  input \WX801_reg/NET0131  ;
  input \WX803_reg/NET0131  ;
  input \WX805_reg/NET0131  ;
  input \WX807_reg/NET0131  ;
  input \WX809_reg/NET0131  ;
  input \WX811_reg/NET0131  ;
  input \WX813_reg/NET0131  ;
  input \WX815_reg/NET0131  ;
  input \WX817_reg/NET0131  ;
  input \WX819_reg/NET0131  ;
  input \WX821_reg/NET0131  ;
  input \WX823_reg/NET0131  ;
  input \WX825_reg/NET0131  ;
  input \WX827_reg/NET0131  ;
  input \WX829_reg/NET0131  ;
  input \WX831_reg/NET0131  ;
  input \WX833_reg/NET0131  ;
  input \WX835_reg/NET0131  ;
  input \WX837_reg/NET0131  ;
  input \WX839_reg/NET0131  ;
  input \WX8403_reg/NET0131  ;
  input \WX8405_reg/NET0131  ;
  input \WX8407_reg/NET0131  ;
  input \WX8409_reg/NET0131  ;
  input \WX8411_reg/NET0131  ;
  input \WX8413_reg/NET0131  ;
  input \WX8415_reg/NET0131  ;
  input \WX8417_reg/NET0131  ;
  input \WX8419_reg/NET0131  ;
  input \WX841_reg/NET0131  ;
  input \WX8421_reg/NET0131  ;
  input \WX8423_reg/NET0131  ;
  input \WX8425_reg/NET0131  ;
  input \WX8427_reg/NET0131  ;
  input \WX8429_reg/NET0131  ;
  input \WX8431_reg/NET0131  ;
  input \WX8433_reg/NET0131  ;
  input \WX8435_reg/NET0131  ;
  input \WX8437_reg/NET0131  ;
  input \WX8439_reg/NET0131  ;
  input \WX843_reg/NET0131  ;
  input \WX8441_reg/NET0131  ;
  input \WX8443_reg/NET0131  ;
  input \WX8445_reg/NET0131  ;
  input \WX8447_reg/NET0131  ;
  input \WX8449_reg/NET0131  ;
  input \WX8451_reg/NET0131  ;
  input \WX8453_reg/NET0131  ;
  input \WX8455_reg/NET0131  ;
  input \WX8457_reg/NET0131  ;
  input \WX8459_reg/NET0131  ;
  input \WX845_reg/NET0131  ;
  input \WX8461_reg/NET0131  ;
  input \WX8463_reg/NET0131  ;
  input \WX8465_reg/NET0131  ;
  input \WX8467_reg/NET0131  ;
  input \WX8469_reg/NET0131  ;
  input \WX8471_reg/NET0131  ;
  input \WX8473_reg/NET0131  ;
  input \WX8475_reg/NET0131  ;
  input \WX8477_reg/NET0131  ;
  input \WX8479_reg/NET0131  ;
  input \WX847_reg/NET0131  ;
  input \WX8481_reg/NET0131  ;
  input \WX8483_reg/NET0131  ;
  input \WX8485_reg/NET0131  ;
  input \WX8487_reg/NET0131  ;
  input \WX8489_reg/NET0131  ;
  input \WX8491_reg/NET0131  ;
  input \WX8493_reg/NET0131  ;
  input \WX8495_reg/NET0131  ;
  input \WX8497_reg/NET0131  ;
  input \WX8499_reg/NET0131  ;
  input \WX849_reg/NET0131  ;
  input \WX8501_reg/NET0131  ;
  input \WX8503_reg/NET0131  ;
  input \WX8505_reg/NET0131  ;
  input \WX8507_reg/NET0131  ;
  input \WX8509_reg/NET0131  ;
  input \WX8511_reg/NET0131  ;
  input \WX8513_reg/NET0131  ;
  input \WX8515_reg/NET0131  ;
  input \WX8517_reg/NET0131  ;
  input \WX8519_reg/NET0131  ;
  input \WX851_reg/NET0131  ;
  input \WX8521_reg/NET0131  ;
  input \WX8523_reg/NET0131  ;
  input \WX8525_reg/NET0131  ;
  input \WX8527_reg/NET0131  ;
  input \WX8529_reg/NET0131  ;
  input \WX8531_reg/NET0131  ;
  input \WX8533_reg/NET0131  ;
  input \WX8535_reg/NET0131  ;
  input \WX8537_reg/NET0131  ;
  input \WX8539_reg/NET0131  ;
  input \WX853_reg/NET0131  ;
  input \WX8541_reg/NET0131  ;
  input \WX8543_reg/NET0131  ;
  input \WX8545_reg/NET0131  ;
  input \WX8547_reg/NET0131  ;
  input \WX8549_reg/NET0131  ;
  input \WX8551_reg/NET0131  ;
  input \WX8553_reg/NET0131  ;
  input \WX8555_reg/NET0131  ;
  input \WX8557_reg/NET0131  ;
  input \WX8559_reg/NET0131  ;
  input \WX855_reg/NET0131  ;
  input \WX8561_reg/NET0131  ;
  input \WX8563_reg/NET0131  ;
  input \WX8565_reg/NET0131  ;
  input \WX8567_reg/NET0131  ;
  input \WX8569_reg/NET0131  ;
  input \WX8571_reg/NET0131  ;
  input \WX8573_reg/NET0131  ;
  input \WX8575_reg/NET0131  ;
  input \WX8577_reg/NET0131  ;
  input \WX8579_reg/NET0131  ;
  input \WX857_reg/NET0131  ;
  input \WX8581_reg/NET0131  ;
  input \WX8583_reg/NET0131  ;
  input \WX8585_reg/NET0131  ;
  input \WX8587_reg/NET0131  ;
  input \WX8589_reg/NET0131  ;
  input \WX8591_reg/NET0131  ;
  input \WX8593_reg/NET0131  ;
  input \WX8595_reg/NET0131  ;
  input \WX8597_reg/NET0131  ;
  input \WX8599_reg/NET0131  ;
  input \WX859_reg/NET0131  ;
  input \WX8601_reg/NET0131  ;
  input \WX8603_reg/NET0131  ;
  input \WX8605_reg/NET0131  ;
  input \WX8607_reg/NET0131  ;
  input \WX8609_reg/NET0131  ;
  input \WX8611_reg/NET0131  ;
  input \WX8613_reg/NET0131  ;
  input \WX8615_reg/NET0131  ;
  input \WX8617_reg/NET0131  ;
  input \WX8619_reg/NET0131  ;
  input \WX861_reg/NET0131  ;
  input \WX8621_reg/NET0131  ;
  input \WX8623_reg/NET0131  ;
  input \WX8625_reg/NET0131  ;
  input \WX8627_reg/NET0131  ;
  input \WX8629_reg/NET0131  ;
  input \WX8631_reg/NET0131  ;
  input \WX8633_reg/NET0131  ;
  input \WX8635_reg/NET0131  ;
  input \WX8637_reg/NET0131  ;
  input \WX8639_reg/NET0131  ;
  input \WX863_reg/NET0131  ;
  input \WX8641_reg/NET0131  ;
  input \WX8643_reg/NET0131  ;
  input \WX8645_reg/NET0131  ;
  input \WX8647_reg/NET0131  ;
  input \WX8649_reg/NET0131  ;
  input \WX8651_reg/NET0131  ;
  input \WX8653_reg/NET0131  ;
  input \WX8655_reg/NET0131  ;
  input \WX8657_reg/NET0131  ;
  input \WX865_reg/NET0131  ;
  input \WX867_reg/NET0131  ;
  input \WX869_reg/NET0131  ;
  input \WX871_reg/NET0131  ;
  input \WX873_reg/NET0131  ;
  input \WX875_reg/NET0131  ;
  input \WX877_reg/NET0131  ;
  input \WX879_reg/NET0131  ;
  input \WX881_reg/NET0131  ;
  input \WX883_reg/NET0131  ;
  input \WX885_reg/NET0131  ;
  input \WX887_reg/NET0131  ;
  input \WX889_reg/NET0131  ;
  input \WX891_reg/NET0131  ;
  input \WX893_reg/NET0131  ;
  input \WX895_reg/NET0131  ;
  input \WX897_reg/NET0131  ;
  input \WX899_reg/NET0131  ;
  input \WX9696_reg/NET0131  ;
  input \WX9698_reg/NET0131  ;
  input \WX9700_reg/NET0131  ;
  input \WX9702_reg/NET0131  ;
  input \WX9704_reg/NET0131  ;
  input \WX9706_reg/NET0131  ;
  input \WX9708_reg/NET0131  ;
  input \WX9710_reg/NET0131  ;
  input \WX9712_reg/NET0131  ;
  input \WX9714_reg/NET0131  ;
  input \WX9716_reg/NET0131  ;
  input \WX9718_reg/NET0131  ;
  input \WX9720_reg/NET0131  ;
  input \WX9722_reg/NET0131  ;
  input \WX9724_reg/NET0131  ;
  input \WX9726_reg/NET0131  ;
  input \WX9728_reg/NET0131  ;
  input \WX9730_reg/NET0131  ;
  input \WX9732_reg/NET0131  ;
  input \WX9734_reg/NET0131  ;
  input \WX9736_reg/NET0131  ;
  input \WX9738_reg/NET0131  ;
  input \WX9740_reg/NET0131  ;
  input \WX9742_reg/NET0131  ;
  input \WX9744_reg/NET0131  ;
  input \WX9746_reg/NET0131  ;
  input \WX9748_reg/NET0131  ;
  input \WX9750_reg/NET0131  ;
  input \WX9752_reg/NET0131  ;
  input \WX9754_reg/NET0131  ;
  input \WX9756_reg/NET0131  ;
  input \WX9758_reg/NET0131  ;
  input \WX9760_reg/NET0131  ;
  input \WX9762_reg/NET0131  ;
  input \WX9764_reg/NET0131  ;
  input \WX9766_reg/NET0131  ;
  input \WX9768_reg/NET0131  ;
  input \WX9770_reg/NET0131  ;
  input \WX9772_reg/NET0131  ;
  input \WX9774_reg/NET0131  ;
  input \WX9776_reg/NET0131  ;
  input \WX9778_reg/NET0131  ;
  input \WX9780_reg/NET0131  ;
  input \WX9782_reg/NET0131  ;
  input \WX9784_reg/NET0131  ;
  input \WX9786_reg/NET0131  ;
  input \WX9788_reg/NET0131  ;
  input \WX9790_reg/NET0131  ;
  input \WX9792_reg/NET0131  ;
  input \WX9794_reg/NET0131  ;
  input \WX9796_reg/NET0131  ;
  input \WX9798_reg/NET0131  ;
  input \WX9800_reg/NET0131  ;
  input \WX9802_reg/NET0131  ;
  input \WX9804_reg/NET0131  ;
  input \WX9806_reg/NET0131  ;
  input \WX9808_reg/NET0131  ;
  input \WX9810_reg/NET0131  ;
  input \WX9812_reg/NET0131  ;
  input \WX9814_reg/NET0131  ;
  input \WX9816_reg/NET0131  ;
  input \WX9818_reg/NET0131  ;
  input \WX9820_reg/NET0131  ;
  input \WX9822_reg/NET0131  ;
  input \WX9824_reg/NET0131  ;
  input \WX9826_reg/NET0131  ;
  input \WX9828_reg/NET0131  ;
  input \WX9830_reg/NET0131  ;
  input \WX9832_reg/NET0131  ;
  input \WX9834_reg/NET0131  ;
  input \WX9836_reg/NET0131  ;
  input \WX9838_reg/NET0131  ;
  input \WX9840_reg/NET0131  ;
  input \WX9842_reg/NET0131  ;
  input \WX9844_reg/NET0131  ;
  input \WX9846_reg/NET0131  ;
  input \WX9848_reg/NET0131  ;
  input \WX9850_reg/NET0131  ;
  input \WX9852_reg/NET0131  ;
  input \WX9854_reg/NET0131  ;
  input \WX9856_reg/NET0131  ;
  input \WX9858_reg/NET0131  ;
  input \WX9860_reg/NET0131  ;
  input \WX9862_reg/NET0131  ;
  input \WX9864_reg/NET0131  ;
  input \WX9866_reg/NET0131  ;
  input \WX9868_reg/NET0131  ;
  input \WX9870_reg/NET0131  ;
  input \WX9872_reg/NET0131  ;
  input \WX9874_reg/NET0131  ;
  input \WX9876_reg/NET0131  ;
  input \WX9878_reg/NET0131  ;
  input \WX9880_reg/NET0131  ;
  input \WX9882_reg/NET0131  ;
  input \WX9884_reg/NET0131  ;
  input \WX9886_reg/NET0131  ;
  input \WX9888_reg/NET0131  ;
  input \WX9890_reg/NET0131  ;
  input \WX9892_reg/NET0131  ;
  input \WX9894_reg/NET0131  ;
  input \WX9896_reg/NET0131  ;
  input \WX9898_reg/NET0131  ;
  input \WX9900_reg/NET0131  ;
  input \WX9902_reg/NET0131  ;
  input \WX9904_reg/NET0131  ;
  input \WX9906_reg/NET0131  ;
  input \WX9908_reg/NET0131  ;
  input \WX9910_reg/NET0131  ;
  input \WX9912_reg/NET0131  ;
  input \WX9914_reg/NET0131  ;
  input \WX9916_reg/NET0131  ;
  input \WX9918_reg/NET0131  ;
  input \WX9920_reg/NET0131  ;
  input \WX9922_reg/NET0131  ;
  input \WX9924_reg/NET0131  ;
  input \WX9926_reg/NET0131  ;
  input \WX9928_reg/NET0131  ;
  input \WX9930_reg/NET0131  ;
  input \WX9932_reg/NET0131  ;
  input \WX9934_reg/NET0131  ;
  input \WX9936_reg/NET0131  ;
  input \WX9938_reg/NET0131  ;
  input \WX9940_reg/NET0131  ;
  input \WX9942_reg/NET0131  ;
  input \WX9944_reg/NET0131  ;
  input \WX9946_reg/NET0131  ;
  input \WX9948_reg/NET0131  ;
  input \WX9950_reg/NET0131  ;
  input \_2077__reg/NET0131  ;
  input \_2078__reg/NET0131  ;
  input \_2079__reg/NET0131  ;
  input \_2080__reg/NET0131  ;
  input \_2081__reg/NET0131  ;
  input \_2082__reg/NET0131  ;
  input \_2083__reg/NET0131  ;
  input \_2084__reg/NET0131  ;
  input \_2085__reg/NET0131  ;
  input \_2086__reg/NET0131  ;
  input \_2087__reg/NET0131  ;
  input \_2088__reg/NET0131  ;
  input \_2089__reg/NET0131  ;
  input \_2090__reg/NET0131  ;
  input \_2091__reg/NET0131  ;
  input \_2092__reg/NET0131  ;
  input \_2093__reg/NET0131  ;
  input \_2094__reg/NET0131  ;
  input \_2095__reg/NET0131  ;
  input \_2096__reg/NET0131  ;
  input \_2097__reg/NET0131  ;
  input \_2098__reg/NET0131  ;
  input \_2099__reg/NET0131  ;
  input \_2100__reg/NET0131  ;
  input \_2101__reg/NET0131  ;
  input \_2102__reg/NET0131  ;
  input \_2103__reg/NET0131  ;
  input \_2104__reg/NET0131  ;
  input \_2105__reg/NET0131  ;
  input \_2106__reg/NET0131  ;
  input \_2107__reg/NET0131  ;
  input \_2108__reg/NET0131  ;
  input \_2109__reg/NET0131  ;
  input \_2110__reg/NET0131  ;
  input \_2111__reg/NET0131  ;
  input \_2112__reg/NET0131  ;
  input \_2113__reg/NET0131  ;
  input \_2114__reg/NET0131  ;
  input \_2115__reg/NET0131  ;
  input \_2116__reg/NET0131  ;
  input \_2117__reg/NET0131  ;
  input \_2118__reg/NET0131  ;
  input \_2119__reg/NET0131  ;
  input \_2120__reg/NET0131  ;
  input \_2121__reg/NET0131  ;
  input \_2122__reg/NET0131  ;
  input \_2123__reg/NET0131  ;
  input \_2124__reg/NET0131  ;
  input \_2125__reg/NET0131  ;
  input \_2126__reg/NET0131  ;
  input \_2127__reg/NET0131  ;
  input \_2128__reg/NET0131  ;
  input \_2129__reg/NET0131  ;
  input \_2130__reg/NET0131  ;
  input \_2131__reg/NET0131  ;
  input \_2132__reg/NET0131  ;
  input \_2133__reg/NET0131  ;
  input \_2134__reg/NET0131  ;
  input \_2135__reg/NET0131  ;
  input \_2136__reg/NET0131  ;
  input \_2137__reg/NET0131  ;
  input \_2138__reg/NET0131  ;
  input \_2139__reg/NET0131  ;
  input \_2140__reg/NET0131  ;
  input \_2141__reg/NET0131  ;
  input \_2142__reg/NET0131  ;
  input \_2143__reg/NET0131  ;
  input \_2144__reg/NET0131  ;
  input \_2145__reg/NET0131  ;
  input \_2146__reg/NET0131  ;
  input \_2147__reg/NET0131  ;
  input \_2148__reg/NET0131  ;
  input \_2149__reg/NET0131  ;
  input \_2150__reg/NET0131  ;
  input \_2151__reg/NET0131  ;
  input \_2152__reg/NET0131  ;
  input \_2153__reg/NET0131  ;
  input \_2154__reg/NET0131  ;
  input \_2155__reg/NET0131  ;
  input \_2156__reg/NET0131  ;
  input \_2157__reg/NET0131  ;
  input \_2158__reg/NET0131  ;
  input \_2159__reg/NET0131  ;
  input \_2160__reg/NET0131  ;
  input \_2161__reg/NET0131  ;
  input \_2162__reg/NET0131  ;
  input \_2163__reg/NET0131  ;
  input \_2164__reg/NET0131  ;
  input \_2165__reg/NET0131  ;
  input \_2166__reg/NET0131  ;
  input \_2167__reg/NET0131  ;
  input \_2168__reg/NET0131  ;
  input \_2169__reg/NET0131  ;
  input \_2170__reg/NET0131  ;
  input \_2171__reg/NET0131  ;
  input \_2172__reg/NET0131  ;
  input \_2173__reg/NET0131  ;
  input \_2174__reg/NET0131  ;
  input \_2175__reg/NET0131  ;
  input \_2176__reg/NET0131  ;
  input \_2177__reg/NET0131  ;
  input \_2178__reg/NET0131  ;
  input \_2179__reg/NET0131  ;
  input \_2180__reg/NET0131  ;
  input \_2181__reg/NET0131  ;
  input \_2182__reg/NET0131  ;
  input \_2183__reg/NET0131  ;
  input \_2184__reg/NET0131  ;
  input \_2185__reg/NET0131  ;
  input \_2186__reg/NET0131  ;
  input \_2187__reg/NET0131  ;
  input \_2188__reg/NET0131  ;
  input \_2189__reg/NET0131  ;
  input \_2190__reg/NET0131  ;
  input \_2191__reg/NET0131  ;
  input \_2192__reg/NET0131  ;
  input \_2193__reg/NET0131  ;
  input \_2194__reg/NET0131  ;
  input \_2195__reg/NET0131  ;
  input \_2196__reg/NET0131  ;
  input \_2197__reg/NET0131  ;
  input \_2198__reg/NET0131  ;
  input \_2199__reg/NET0131  ;
  input \_2200__reg/NET0131  ;
  input \_2201__reg/NET0131  ;
  input \_2202__reg/NET0131  ;
  input \_2203__reg/NET0131  ;
  input \_2204__reg/NET0131  ;
  input \_2205__reg/NET0131  ;
  input \_2206__reg/NET0131  ;
  input \_2207__reg/NET0131  ;
  input \_2208__reg/NET0131  ;
  input \_2209__reg/NET0131  ;
  input \_2210__reg/NET0131  ;
  input \_2211__reg/NET0131  ;
  input \_2212__reg/NET0131  ;
  input \_2213__reg/NET0131  ;
  input \_2214__reg/NET0131  ;
  input \_2215__reg/NET0131  ;
  input \_2216__reg/NET0131  ;
  input \_2217__reg/NET0131  ;
  input \_2218__reg/NET0131  ;
  input \_2219__reg/NET0131  ;
  input \_2220__reg/NET0131  ;
  input \_2221__reg/NET0131  ;
  input \_2222__reg/NET0131  ;
  input \_2223__reg/NET0131  ;
  input \_2224__reg/NET0131  ;
  input \_2225__reg/NET0131  ;
  input \_2226__reg/NET0131  ;
  input \_2227__reg/NET0131  ;
  input \_2228__reg/NET0131  ;
  input \_2229__reg/NET0131  ;
  input \_2230__reg/NET0131  ;
  input \_2231__reg/NET0131  ;
  input \_2232__reg/NET0131  ;
  input \_2233__reg/NET0131  ;
  input \_2234__reg/NET0131  ;
  input \_2235__reg/NET0131  ;
  input \_2236__reg/NET0131  ;
  input \_2237__reg/NET0131  ;
  input \_2238__reg/NET0131  ;
  input \_2239__reg/NET0131  ;
  input \_2240__reg/NET0131  ;
  input \_2241__reg/NET0131  ;
  input \_2242__reg/NET0131  ;
  input \_2243__reg/NET0131  ;
  input \_2244__reg/NET0131  ;
  input \_2245__reg/NET0131  ;
  input \_2246__reg/NET0131  ;
  input \_2247__reg/NET0131  ;
  input \_2248__reg/NET0131  ;
  input \_2249__reg/NET0131  ;
  input \_2250__reg/NET0131  ;
  input \_2251__reg/NET0131  ;
  input \_2252__reg/NET0131  ;
  input \_2253__reg/NET0131  ;
  input \_2254__reg/NET0131  ;
  input \_2255__reg/NET0131  ;
  input \_2256__reg/NET0131  ;
  input \_2257__reg/NET0131  ;
  input \_2258__reg/NET0131  ;
  input \_2259__reg/NET0131  ;
  input \_2260__reg/NET0131  ;
  input \_2261__reg/NET0131  ;
  input \_2262__reg/NET0131  ;
  input \_2263__reg/NET0131  ;
  input \_2264__reg/NET0131  ;
  input \_2265__reg/NET0131  ;
  input \_2266__reg/NET0131  ;
  input \_2267__reg/NET0131  ;
  input \_2268__reg/NET0131  ;
  input \_2269__reg/NET0131  ;
  input \_2270__reg/NET0131  ;
  input \_2271__reg/NET0131  ;
  input \_2272__reg/NET0131  ;
  input \_2273__reg/NET0131  ;
  input \_2274__reg/NET0131  ;
  input \_2275__reg/NET0131  ;
  input \_2276__reg/NET0131  ;
  input \_2277__reg/NET0131  ;
  input \_2278__reg/NET0131  ;
  input \_2279__reg/NET0131  ;
  input \_2280__reg/NET0131  ;
  input \_2281__reg/NET0131  ;
  input \_2282__reg/NET0131  ;
  input \_2283__reg/NET0131  ;
  input \_2284__reg/NET0131  ;
  input \_2285__reg/NET0131  ;
  input \_2286__reg/NET0131  ;
  input \_2287__reg/NET0131  ;
  input \_2288__reg/NET0131  ;
  input \_2289__reg/NET0131  ;
  input \_2290__reg/NET0131  ;
  input \_2291__reg/NET0131  ;
  input \_2292__reg/NET0131  ;
  input \_2293__reg/NET0131  ;
  input \_2294__reg/NET0131  ;
  input \_2295__reg/NET0131  ;
  input \_2296__reg/NET0131  ;
  input \_2297__reg/NET0131  ;
  input \_2298__reg/NET0131  ;
  input \_2299__reg/NET0131  ;
  input \_2300__reg/NET0131  ;
  input \_2301__reg/NET0131  ;
  input \_2302__reg/NET0131  ;
  input \_2303__reg/NET0131  ;
  input \_2304__reg/NET0131  ;
  input \_2305__reg/NET0131  ;
  input \_2306__reg/NET0131  ;
  input \_2307__reg/NET0131  ;
  input \_2308__reg/NET0131  ;
  input \_2309__reg/NET0131  ;
  input \_2310__reg/NET0131  ;
  input \_2311__reg/NET0131  ;
  input \_2312__reg/NET0131  ;
  input \_2313__reg/NET0131  ;
  input \_2314__reg/NET0131  ;
  input \_2315__reg/NET0131  ;
  input \_2316__reg/NET0131  ;
  input \_2317__reg/NET0131  ;
  input \_2318__reg/NET0131  ;
  input \_2319__reg/NET0131  ;
  input \_2320__reg/NET0131  ;
  input \_2321__reg/NET0131  ;
  input \_2322__reg/NET0131  ;
  input \_2323__reg/NET0131  ;
  input \_2324__reg/NET0131  ;
  input \_2325__reg/NET0131  ;
  input \_2326__reg/NET0131  ;
  input \_2327__reg/NET0131  ;
  input \_2328__reg/NET0131  ;
  input \_2329__reg/NET0131  ;
  input \_2330__reg/NET0131  ;
  input \_2331__reg/NET0131  ;
  input \_2332__reg/NET0131  ;
  input \_2333__reg/NET0131  ;
  input \_2334__reg/NET0131  ;
  input \_2335__reg/NET0131  ;
  input \_2336__reg/NET0131  ;
  input \_2337__reg/NET0131  ;
  input \_2338__reg/NET0131  ;
  input \_2339__reg/NET0131  ;
  input \_2340__reg/NET0131  ;
  input \_2341__reg/NET0131  ;
  input \_2342__reg/NET0131  ;
  input \_2343__reg/NET0131  ;
  input \_2344__reg/NET0131  ;
  input \_2345__reg/NET0131  ;
  input \_2346__reg/NET0131  ;
  input \_2347__reg/NET0131  ;
  input \_2348__reg/NET0131  ;
  input \_2349__reg/NET0131  ;
  input \_2350__reg/NET0131  ;
  input \_2351__reg/NET0131  ;
  input \_2352__reg/NET0131  ;
  input \_2353__reg/NET0131  ;
  input \_2354__reg/NET0131  ;
  input \_2355__reg/NET0131  ;
  input \_2356__reg/NET0131  ;
  input \_2357__reg/NET0131  ;
  input \_2358__reg/NET0131  ;
  input \_2359__reg/NET0131  ;
  input \_2360__reg/NET0131  ;
  input \_2361__reg/NET0131  ;
  input \_2362__reg/NET0131  ;
  input \_2363__reg/NET0131  ;
  input \_2364__reg/NET0131  ;
  output \DATA_9_0_pad  ;
  output \DATA_9_10_pad  ;
  output \DATA_9_11_pad  ;
  output \DATA_9_12_pad  ;
  output \DATA_9_13_pad  ;
  output \DATA_9_14_pad  ;
  output \DATA_9_15_pad  ;
  output \DATA_9_16_pad  ;
  output \DATA_9_17_pad  ;
  output \DATA_9_18_pad  ;
  output \DATA_9_19_pad  ;
  output \DATA_9_1_pad  ;
  output \DATA_9_20_pad  ;
  output \DATA_9_21_pad  ;
  output \DATA_9_22_pad  ;
  output \DATA_9_23_pad  ;
  output \DATA_9_24_pad  ;
  output \DATA_9_25_pad  ;
  output \DATA_9_26_pad  ;
  output \DATA_9_27_pad  ;
  output \DATA_9_28_pad  ;
  output \DATA_9_29_pad  ;
  output \DATA_9_2_pad  ;
  output \DATA_9_30_pad  ;
  output \DATA_9_31_pad  ;
  output \DATA_9_3_pad  ;
  output \DATA_9_4_pad  ;
  output \DATA_9_5_pad  ;
  output \DATA_9_6_pad  ;
  output \DATA_9_7_pad  ;
  output \DATA_9_8_pad  ;
  output \DATA_9_9_pad  ;
  output \_al_n0  ;
  output \_al_n1  ;
  output \g19/_0_  ;
  output \g35/_0_  ;
  output \g36/_0_  ;
  output \g40/_0_  ;
  output \g55780/_0_  ;
  output \g55783/_0_  ;
  output \g55795/_0_  ;
  output \g55796/_0_  ;
  output \g55797/_0_  ;
  output \g55798/_0_  ;
  output \g55799/_0_  ;
  output \g55800/_0_  ;
  output \g55801/_0_  ;
  output \g55802/_0_  ;
  output \g55803/_0_  ;
  output \g55834/_0_  ;
  output \g55835/_0_  ;
  output \g55836/_0_  ;
  output \g55837/_0_  ;
  output \g55838/_0_  ;
  output \g55839/_0_  ;
  output \g55840/_0_  ;
  output \g55841/_0_  ;
  output \g55842/_0_  ;
  output \g55856/_0_  ;
  output \g55894/_0_  ;
  output \g55895/_0_  ;
  output \g55896/_0_  ;
  output \g55897/_0_  ;
  output \g55898/_0_  ;
  output \g55899/_0_  ;
  output \g55900/_0_  ;
  output \g55901/_0_  ;
  output \g55902/_0_  ;
  output \g55916/_0_  ;
  output \g55953/_0_  ;
  output \g55954/_0_  ;
  output \g55955/_0_  ;
  output \g55956/_0_  ;
  output \g55957/_0_  ;
  output \g55958/_0_  ;
  output \g55959/_0_  ;
  output \g55960/_0_  ;
  output \g55961/_0_  ;
  output \g55975/_0_  ;
  output \g56012/_0_  ;
  output \g56013/_0_  ;
  output \g56014/_0_  ;
  output \g56015/_0_  ;
  output \g56016/_0_  ;
  output \g56017/_0_  ;
  output \g56018/_0_  ;
  output \g56019/_0_  ;
  output \g56020/_0_  ;
  output \g56034/_0_  ;
  output \g56071/_0_  ;
  output \g56072/_0_  ;
  output \g56073/_0_  ;
  output \g56074/_0_  ;
  output \g56075/_0_  ;
  output \g56076/_0_  ;
  output \g56077/_0_  ;
  output \g56078/_0_  ;
  output \g56079/_0_  ;
  output \g56093/_0_  ;
  output \g56130/_0_  ;
  output \g56131/_0_  ;
  output \g56132/_0_  ;
  output \g56133/_0_  ;
  output \g56134/_0_  ;
  output \g56135/_0_  ;
  output \g56136/_0_  ;
  output \g56137/_0_  ;
  output \g56138/_0_  ;
  output \g56152/_0_  ;
  output \g56189/_0_  ;
  output \g56190/_0_  ;
  output \g56191/_0_  ;
  output \g56192/_0_  ;
  output \g56193/_0_  ;
  output \g56194/_0_  ;
  output \g56195/_0_  ;
  output \g56196/_0_  ;
  output \g56197/_0_  ;
  output \g56211/_0_  ;
  output \g56248/_0_  ;
  output \g56249/_0_  ;
  output \g56250/_0_  ;
  output \g56251/_0_  ;
  output \g56252/_0_  ;
  output \g56253/_0_  ;
  output \g56254/_0_  ;
  output \g56255/_0_  ;
  output \g56256/_0_  ;
  output \g56270/_0_  ;
  output \g56307/_0_  ;
  output \g56308/_0_  ;
  output \g56309/_0_  ;
  output \g56310/_0_  ;
  output \g56311/_0_  ;
  output \g56312/_0_  ;
  output \g56313/_0_  ;
  output \g56314/_0_  ;
  output \g56315/_0_  ;
  output \g56329/_0_  ;
  output \g56366/_0_  ;
  output \g56367/_0_  ;
  output \g56368/_0_  ;
  output \g56369/_0_  ;
  output \g56370/_0_  ;
  output \g56371/_0_  ;
  output \g56372/_0_  ;
  output \g56373/_0_  ;
  output \g56374/_0_  ;
  output \g56388/_0_  ;
  output \g56425/_0_  ;
  output \g56426/_0_  ;
  output \g56427/_0_  ;
  output \g56428/_0_  ;
  output \g56429/_0_  ;
  output \g56430/_0_  ;
  output \g56431/_0_  ;
  output \g56432/_0_  ;
  output \g56433/_0_  ;
  output \g56447/_0_  ;
  output \g56484/_0_  ;
  output \g56485/_0_  ;
  output \g56486/_0_  ;
  output \g56487/_0_  ;
  output \g56488/_0_  ;
  output \g56489/_0_  ;
  output \g56490/_0_  ;
  output \g56491/_0_  ;
  output \g56492/_0_  ;
  output \g56507/_0_  ;
  output \g56543/_0_  ;
  output \g56544/_0_  ;
  output \g56545/_0_  ;
  output \g56546/_0_  ;
  output \g56547/_0_  ;
  output \g56548/_0_  ;
  output \g56549/_0_  ;
  output \g56551/_0_  ;
  output \g56567/_0_  ;
  output \g56602/_0_  ;
  output \g56603/_0_  ;
  output \g56604/_0_  ;
  output \g56605/_0_  ;
  output \g56606/_0_  ;
  output \g56607/_0_  ;
  output \g56608/_0_  ;
  output \g56610/_0_  ;
  output \g56627/_0_  ;
  output \g56661/_0_  ;
  output \g56662/_0_  ;
  output \g56663/_0_  ;
  output \g56664/_0_  ;
  output \g56665/_0_  ;
  output \g56666/_0_  ;
  output \g56667/_0_  ;
  output \g56668/_0_  ;
  output \g56686/_0_  ;
  output \g56720/_0_  ;
  output \g56721/_0_  ;
  output \g56722/_0_  ;
  output \g56723/_0_  ;
  output \g56724/_0_  ;
  output \g56725/_0_  ;
  output \g56726/_0_  ;
  output \g56727/_0_  ;
  output \g56728/_0_  ;
  output \g56745/_0_  ;
  output \g56779/_0_  ;
  output \g56780/_0_  ;
  output \g56781/_0_  ;
  output \g56782/_0_  ;
  output \g56783/_0_  ;
  output \g56784/_0_  ;
  output \g56785/_0_  ;
  output \g56804/_0_  ;
  output \g56838/_0_  ;
  output \g56839/_0_  ;
  output \g56840/_0_  ;
  output \g56841/_0_  ;
  output \g56842/_0_  ;
  output \g56843/_0_  ;
  output \g56844/_0_  ;
  output \g56845/_0_  ;
  output \g56846/_0_  ;
  output \g56863/_0_  ;
  output \g56897/_0_  ;
  output \g56898/_0_  ;
  output \g56899/_0_  ;
  output \g56900/_0_  ;
  output \g56901/_0_  ;
  output \g56902/_0_  ;
  output \g56903/_0_  ;
  output \g56905/_0_  ;
  output \g56921/_0_  ;
  output \g56956/_0_  ;
  output \g56957/_0_  ;
  output \g56958/_0_  ;
  output \g56959/_0_  ;
  output \g56960/_0_  ;
  output \g56961/_0_  ;
  output \g56962/_0_  ;
  output \g56964/_0_  ;
  output \g56980/_0_  ;
  output \g57015/_0_  ;
  output \g57016/_0_  ;
  output \g57017/_0_  ;
  output \g57018/_0_  ;
  output \g57019/_0_  ;
  output \g57020/_0_  ;
  output \g57021/_0_  ;
  output \g57023/_0_  ;
  output \g57040/_0_  ;
  output \g57074/_0_  ;
  output \g57075/_0_  ;
  output \g57076/_0_  ;
  output \g57077/_0_  ;
  output \g57078/_0_  ;
  output \g57079/_0_  ;
  output \g57080/_0_  ;
  output \g57081/_0_  ;
  output \g57099/_0_  ;
  output \g57133/_0_  ;
  output \g57134/_0_  ;
  output \g57135/_0_  ;
  output \g57136/_0_  ;
  output \g57137/_0_  ;
  output \g57138/_0_  ;
  output \g57139/_0_  ;
  output \g57140/_0_  ;
  output \g57141/_0_  ;
  output \g57159/_0_  ;
  output \g57193/_0_  ;
  output \g57195/_0_  ;
  output \g57196/_0_  ;
  output \g57197/_0_  ;
  output \g57198/_0_  ;
  output \g57199/_0_  ;
  output \g57200/_0_  ;
  output \g57202/_0_  ;
  output \g57219/_0_  ;
  output \g57254/_0_  ;
  output \g57255/_0_  ;
  output \g57256/_0_  ;
  output \g57257/_0_  ;
  output \g57258/_0_  ;
  output \g57259/_0_  ;
  output \g57260/_0_  ;
  output \g57262/_0_  ;
  output \g57263/_0_  ;
  output \g57285/_0_  ;
  output \g57318/_0_  ;
  output \g57319/_0_  ;
  output \g57320/_0_  ;
  output \g57321/_0_  ;
  output \g57322/_0_  ;
  output \g57323/_0_  ;
  output \g57324/_0_  ;
  output \g57325/_0_  ;
  output \g57326/_0_  ;
  output \g57328/_0_  ;
  output \g57329/_0_  ;
  output \g57330/_0_  ;
  output \g57350/_0_  ;
  output \g57387/_0_  ;
  output \g57388/_0_  ;
  output \g57390/_0_  ;
  output \g57391/_0_  ;
  output \g57392/_0_  ;
  output \g57393/_0_  ;
  output \g57395/_0_  ;
  output \g57396/_0_  ;
  output \g57439/_0_  ;
  output \g57476/_0_  ;
  output \g57477/_0_  ;
  output \g57478/_0_  ;
  output \g57479/_0_  ;
  output \g57480/_0_  ;
  output \g57481/_0_  ;
  output \g57482/_0_  ;
  output \g57483/_0_  ;
  output \g57484/_0_  ;
  output \g57485/_0_  ;
  output \g57486/_0_  ;
  output \g57487/_0_  ;
  output \g57488/_0_  ;
  output \g57489/_0_  ;
  output \g57490/_0_  ;
  output \g57491/_0_  ;
  output \g57492/_0_  ;
  output \g57493/_0_  ;
  output \g57494/_0_  ;
  output \g57495/_0_  ;
  output \g57496/_0_  ;
  output \g57497/_0_  ;
  output \g57498/_0_  ;
  output \g57499/_0_  ;
  output \g57500/_0_  ;
  output \g57501/_0_  ;
  output \g57502/_0_  ;
  output \g57503/_0_  ;
  output \g57504/_0_  ;
  output \g57505/_0_  ;
  output \g57524/_0_  ;
  output \g57537/_0_  ;
  output \g57541/_0_  ;
  output \g57543/_0_  ;
  output \g58163/_0_  ;
  output \g58572/_0_  ;
  output \g58573/_0_  ;
  output \g58574/_0_  ;
  output \g58575/_0_  ;
  output \g58576/_0_  ;
  output \g58577/_0_  ;
  output \g58578/_0_  ;
  output \g58579/_0_  ;
  output \g58580/_0_  ;
  output \g58581/_0_  ;
  output \g58582/_0_  ;
  output \g58583/_0_  ;
  output \g58584/_0_  ;
  output \g58585/_0_  ;
  output \g58586/_0_  ;
  output \g58587/_0_  ;
  output \g58588/_0_  ;
  output \g58589/_0_  ;
  output \g58590/_0_  ;
  output \g58591/_0_  ;
  output \g58592/_0_  ;
  output \g58593/_0_  ;
  output \g58594/_0_  ;
  output \g58595/_0_  ;
  output \g58596/_0_  ;
  output \g58597/_0_  ;
  output \g58598/_0_  ;
  output \g58600/_0_  ;
  output \g58602/_0_  ;
  output \g58604/_0_  ;
  output \g58615/_0_  ;
  output \g59240/_0_  ;
  output \g59241/_0_  ;
  output \g59242/_0_  ;
  output \g59243/_0_  ;
  output \g59244/_0_  ;
  output \g59245/_0_  ;
  output \g59246/_0_  ;
  output \g59247/_0_  ;
  output \g59248/_0_  ;
  output \g59249/_0_  ;
  output \g59250/_0_  ;
  output \g59251/_0_  ;
  output \g59252/_0_  ;
  output \g59253/_0_  ;
  output \g59254/_0_  ;
  output \g59255/_0_  ;
  output \g59256/_0_  ;
  output \g59257/_0_  ;
  output \g59258/_0_  ;
  output \g59259/_0_  ;
  output \g59260/_0_  ;
  output \g59261/_0_  ;
  output \g59262/_0_  ;
  output \g59263/_0_  ;
  output \g59264/_0_  ;
  output \g59265/_0_  ;
  output \g59266/_0_  ;
  output \g59267/_0_  ;
  output \g59268/_0_  ;
  output \g59269/_0_  ;
  output \g59270/_0_  ;
  output \g59271/_0_  ;
  output \g59272/_0_  ;
  output \g59273/_0_  ;
  output \g59274/_0_  ;
  output \g59275/_0_  ;
  output \g59276/_0_  ;
  output \g59277/_0_  ;
  output \g59278/_0_  ;
  output \g59279/_0_  ;
  output \g59280/_0_  ;
  output \g59281/_0_  ;
  output \g59282/_0_  ;
  output \g59283/_0_  ;
  output \g59284/_0_  ;
  output \g59285/_0_  ;
  output \g59286/_0_  ;
  output \g59287/_0_  ;
  output \g59288/_0_  ;
  output \g59289/_0_  ;
  output \g59290/_0_  ;
  output \g59291/_0_  ;
  output \g59292/_0_  ;
  output \g59293/_0_  ;
  output \g59294/_0_  ;
  output \g59295/_0_  ;
  output \g59296/_0_  ;
  output \g59297/_0_  ;
  output \g59298/_0_  ;
  output \g59299/_0_  ;
  output \g59300/_0_  ;
  output \g59301/_0_  ;
  output \g59302/_0_  ;
  output \g59303/_0_  ;
  output \g59304/_0_  ;
  output \g59305/_0_  ;
  output \g59306/_0_  ;
  output \g59307/_0_  ;
  output \g59308/_0_  ;
  output \g59309/_0_  ;
  output \g59310/_0_  ;
  output \g59311/_0_  ;
  output \g59312/_0_  ;
  output \g59313/_0_  ;
  output \g59314/_0_  ;
  output \g59315/_0_  ;
  output \g59316/_0_  ;
  output \g59317/_0_  ;
  output \g59318/_0_  ;
  output \g59319/_0_  ;
  output \g59320/_0_  ;
  output \g59321/_0_  ;
  output \g59322/_0_  ;
  output \g59323/_0_  ;
  output \g59324/_0_  ;
  output \g59325/_0_  ;
  output \g59326/_0_  ;
  output \g59327/_0_  ;
  output \g59328/_0_  ;
  output \g59329/_0_  ;
  output \g59330/_0_  ;
  output \g59331/_0_  ;
  output \g59332/_0_  ;
  output \g59333/_0_  ;
  output \g59334/_0_  ;
  output \g59335/_0_  ;
  output \g59336/_0_  ;
  output \g59337/_0_  ;
  output \g59338/_0_  ;
  output \g59339/_0_  ;
  output \g59340/_0_  ;
  output \g59341/_0_  ;
  output \g59342/_0_  ;
  output \g59343/_0_  ;
  output \g59344/_0_  ;
  output \g59345/_0_  ;
  output \g59346/_0_  ;
  output \g59347/_0_  ;
  output \g59348/_0_  ;
  output \g59349/_0_  ;
  output \g59350/_0_  ;
  output \g59351/_0_  ;
  output \g59352/_0_  ;
  output \g59353/_0_  ;
  output \g59354/_0_  ;
  output \g59355/_0_  ;
  output \g59356/_0_  ;
  output \g59357/_0_  ;
  output \g59358/_0_  ;
  output \g59359/_0_  ;
  output \g59360/_0_  ;
  output \g59361/_0_  ;
  output \g59362/_0_  ;
  output \g59363/_0_  ;
  output \g59364/_0_  ;
  output \g59365/_0_  ;
  output \g59366/_0_  ;
  output \g59367/_0_  ;
  output \g59368/_0_  ;
  output \g59369/_0_  ;
  output \g59370/_0_  ;
  output \g59371/_0_  ;
  output \g59372/_0_  ;
  output \g59373/_0_  ;
  output \g59374/_0_  ;
  output \g59375/_0_  ;
  output \g59376/_0_  ;
  output \g59377/_0_  ;
  output \g59378/_0_  ;
  output \g59379/_0_  ;
  output \g59380/_0_  ;
  output \g59381/_0_  ;
  output \g59382/_0_  ;
  output \g59383/_0_  ;
  output \g59384/_0_  ;
  output \g59385/_0_  ;
  output \g59386/_0_  ;
  output \g59387/_0_  ;
  output \g59388/_0_  ;
  output \g59389/_0_  ;
  output \g59390/_0_  ;
  output \g59391/_0_  ;
  output \g59392/_0_  ;
  output \g59393/_0_  ;
  output \g59394/_0_  ;
  output \g59395/_0_  ;
  output \g59396/_0_  ;
  output \g59397/_0_  ;
  output \g59398/_0_  ;
  output \g59399/_0_  ;
  output \g59400/_0_  ;
  output \g59401/_0_  ;
  output \g59402/_0_  ;
  output \g59403/_0_  ;
  output \g59404/_0_  ;
  output \g59405/_0_  ;
  output \g59406/_0_  ;
  output \g59407/_0_  ;
  output \g59408/_0_  ;
  output \g59409/_0_  ;
  output \g59410/_0_  ;
  output \g59411/_0_  ;
  output \g59412/_0_  ;
  output \g59413/_0_  ;
  output \g59414/_0_  ;
  output \g59415/_0_  ;
  output \g59416/_0_  ;
  output \g59417/_0_  ;
  output \g59418/_0_  ;
  output \g59419/_0_  ;
  output \g59420/_0_  ;
  output \g59421/_0_  ;
  output \g59422/_0_  ;
  output \g59423/_0_  ;
  output \g59424/_0_  ;
  output \g59425/_0_  ;
  output \g59426/_0_  ;
  output \g59427/_0_  ;
  output \g59428/_0_  ;
  output \g59429/_0_  ;
  output \g59430/_0_  ;
  output \g59431/_0_  ;
  output \g59432/_0_  ;
  output \g59433/_0_  ;
  output \g59434/_0_  ;
  output \g59435/_0_  ;
  output \g59436/_0_  ;
  output \g59437/_0_  ;
  output \g59438/_0_  ;
  output \g59439/_0_  ;
  output \g59440/_0_  ;
  output \g59441/_0_  ;
  output \g59442/_0_  ;
  output \g59443/_0_  ;
  output \g59444/_0_  ;
  output \g59445/_0_  ;
  output \g59446/_0_  ;
  output \g59447/_0_  ;
  output \g59448/_0_  ;
  output \g59449/_0_  ;
  output \g59450/_0_  ;
  output \g59451/_0_  ;
  output \g59452/_0_  ;
  output \g59453/_0_  ;
  output \g59454/_0_  ;
  output \g59455/_0_  ;
  output \g59456/_0_  ;
  output \g59457/_0_  ;
  output \g59458/_0_  ;
  output \g59459/_0_  ;
  output \g59460/_0_  ;
  output \g59461/_0_  ;
  output \g59462/_0_  ;
  output \g59463/_0_  ;
  output \g59464/_0_  ;
  output \g59465/_0_  ;
  output \g59466/_0_  ;
  output \g59467/_0_  ;
  output \g59468/_0_  ;
  output \g59469/_0_  ;
  output \g59470/_0_  ;
  output \g59471/_0_  ;
  output \g59472/_0_  ;
  output \g59473/_0_  ;
  output \g59474/_0_  ;
  output \g59475/_0_  ;
  output \g59476/_0_  ;
  output \g59477/_0_  ;
  output \g59478/_0_  ;
  output \g59479/_0_  ;
  output \g59480/_0_  ;
  output \g59481/_0_  ;
  output \g59482/_0_  ;
  output \g59483/_0_  ;
  output \g59484/_0_  ;
  output \g59485/_0_  ;
  output \g59486/_0_  ;
  output \g59487/_0_  ;
  output \g59488/_0_  ;
  output \g59489/_0_  ;
  output \g59490/_0_  ;
  output \g59491/_0_  ;
  output \g59492/_0_  ;
  output \g59493/_0_  ;
  output \g59494/_0_  ;
  output \g59495/_0_  ;
  output \g59496/_0_  ;
  output \g59497/_0_  ;
  output \g59498/_0_  ;
  output \g59500/_0_  ;
  output \g59503/_0_  ;
  output \g59512/_0_  ;
  output \g61336/_0_  ;
  output \g61521/_0_  ;
  output \g61523/_0_  ;
  output \g61524/_0_  ;
  output \g61526/_0_  ;
  output \g61527/_0_  ;
  output \g61528/_0_  ;
  output \g61529/_0_  ;
  output \g61530/_0_  ;
  output \g61531/_0_  ;
  output \g61532/_0_  ;
  output \g61533/_0_  ;
  output \g61535/_0_  ;
  output \g61537/_0_  ;
  output \g61539/_0_  ;
  output \g61540/_0_  ;
  output \g61541/_0_  ;
  output \g61542/_0_  ;
  output \g61546/_0_  ;
  output \g61550/_0_  ;
  output \g61551/_0_  ;
  output \g61552/_0_  ;
  output \g61554/_0_  ;
  output \g61555/_0_  ;
  output \g61556/_0_  ;
  output \g61558/_0_  ;
  output \g61559/_0_  ;
  output \g61561/_0_  ;
  output \g61562/_0_  ;
  output \g61563/_0_  ;
  output \g61564/_0_  ;
  output \g61565/_0_  ;
  output \g61566/_0_  ;
  output \g61568/_0_  ;
  output \g61570/_0_  ;
  output \g61571/_0_  ;
  output \g61572/_0_  ;
  output \g61573/_0_  ;
  output \g61577/_0_  ;
  output \g61578/_0_  ;
  output \g61579/_0_  ;
  output \g61580/_0_  ;
  output \g61581/_0_  ;
  output \g61582/_0_  ;
  output \g61583/_0_  ;
  output \g61584/_0_  ;
  output \g61585/_0_  ;
  output \g61586/_0_  ;
  output \g61587/_0_  ;
  output \g61588/_0_  ;
  output \g61589/_0_  ;
  output \g61591/_0_  ;
  output \g61592/_0_  ;
  output \g61594/_0_  ;
  output \g61595/_0_  ;
  output \g61596/_0_  ;
  output \g61597/_0_  ;
  output \g61598/_0_  ;
  output \g61599/_0_  ;
  output \g61600/_0_  ;
  output \g61601/_0_  ;
  output \g61605/_0_  ;
  output \g61606/_0_  ;
  output \g61607/_0_  ;
  output \g61608/_0_  ;
  output \g61609/_0_  ;
  output \g61610/_0_  ;
  output \g61611/_0_  ;
  output \g61612/_0_  ;
  output \g61613/_0_  ;
  output \g61615/_0_  ;
  output \g61616/_0_  ;
  output \g61617/_0_  ;
  output \g61618/_0_  ;
  output \g61619/_0_  ;
  output \g61620/_0_  ;
  output \g61621/_0_  ;
  output \g61623/_0_  ;
  output \g61624/_0_  ;
  output \g61625/_0_  ;
  output \g61626/_0_  ;
  output \g61627/_0_  ;
  output \g61629/_0_  ;
  output \g61630/_0_  ;
  output \g61631/_0_  ;
  output \g61632/_0_  ;
  output \g61633/_0_  ;
  output \g61634/_0_  ;
  output \g61636/_0_  ;
  output \g61638/_0_  ;
  output \g61639/_0_  ;
  output \g61640/_0_  ;
  output \g61641/_0_  ;
  output \g61642/_0_  ;
  output \g61644/_0_  ;
  output \g61647/_0_  ;
  output \g61648/_0_  ;
  output \g61649/_0_  ;
  output \g61650/_0_  ;
  output \g61653/_0_  ;
  output \g61654/_0_  ;
  output \g61655/_0_  ;
  output \g61656/_0_  ;
  output \g61658/_0_  ;
  output \g61661/_0_  ;
  output \g61662/_0_  ;
  output \g61663/_0_  ;
  output \g61664/_0_  ;
  output \g61666/_0_  ;
  output \g61667/_0_  ;
  output \g61668/_0_  ;
  output \g61670/_0_  ;
  output \g61671/_0_  ;
  output \g61672/_0_  ;
  output \g61673/_0_  ;
  output \g61675/_0_  ;
  output \g61676/_0_  ;
  output \g61680/_0_  ;
  output \g61681/_0_  ;
  output \g61682/_0_  ;
  output \g61683/_0_  ;
  output \g61684/_0_  ;
  output \g61686/_0_  ;
  output \g61687/_0_  ;
  output \g61688/_0_  ;
  output \g61689/_0_  ;
  output \g61690/_0_  ;
  output \g61691/_0_  ;
  output \g61693/_0_  ;
  output \g61694/_0_  ;
  output \g61696/_0_  ;
  output \g61697/_0_  ;
  output \g61698/_0_  ;
  output \g61699/_0_  ;
  output \g61700/_0_  ;
  output \g61701/_0_  ;
  output \g61702/_0_  ;
  output \g61703/_0_  ;
  output \g61704/_0_  ;
  output \g61705/_0_  ;
  output \g61706/_0_  ;
  output \g61707/_0_  ;
  output \g61708/_0_  ;
  output \g61711/_0_  ;
  output \g61712/_0_  ;
  output \g61714/_0_  ;
  output \g61716/_0_  ;
  output \g61717/_0_  ;
  output \g61719/_0_  ;
  output \g61720/_0_  ;
  output \g61721/_0_  ;
  output \g61724/_0_  ;
  output \g61725/_0_  ;
  output \g61728/_0_  ;
  output \g61729/_0_  ;
  output \g61731/_0_  ;
  output \g61732/_0_  ;
  output \g61733/_0_  ;
  output \g61736/_0_  ;
  output \g61737/_0_  ;
  output \g61739/_0_  ;
  output \g61740/_0_  ;
  output \g61741/_0_  ;
  output \g61743/_0_  ;
  output \g61744/_0_  ;
  output \g61745/_0_  ;
  output \g61746/_0_  ;
  output \g61747/_0_  ;
  output \g61748/_0_  ;
  output \g61749/_0_  ;
  output \g61750/_0_  ;
  output \g61751/_0_  ;
  output \g61752/_0_  ;
  output \g61753/_0_  ;
  output \g61754/_0_  ;
  output \g61755/_0_  ;
  output \g61757/_0_  ;
  output \g61758/_0_  ;
  output \g61759/_0_  ;
  output \g61760/_0_  ;
  output \g61761/_0_  ;
  output \g61762/_0_  ;
  output \g61763/_0_  ;
  output \g61764/_0_  ;
  output \g61765/_0_  ;
  output \g61766/_0_  ;
  output \g61767/_0_  ;
  output \g61768/_0_  ;
  output \g61769/_0_  ;
  output \g61770/_0_  ;
  output \g61771/_0_  ;
  output \g61772/_0_  ;
  output \g61773/_0_  ;
  output \g61774/_0_  ;
  output \g61775/_0_  ;
  output \g61776/_0_  ;
  output \g61777/_0_  ;
  output \g61778/_0_  ;
  output \g61780/_0_  ;
  output \g61781/_0_  ;
  output \g61783/_0_  ;
  output \g61784/_0_  ;
  output \g61786/_0_  ;
  output \g61787/_0_  ;
  output \g61790/_0_  ;
  output \g61791/_0_  ;
  output \g61794/_0_  ;
  output \g61795/_0_  ;
  output \g61796/_0_  ;
  output \g61797/_0_  ;
  output \g61798/_0_  ;
  output \g61799/_0_  ;
  output \g61800/_0_  ;
  output \g61801/_0_  ;
  output \g61802/_0_  ;
  output \g61803/_0_  ;
  output \g61805/_0_  ;
  output \g61806/_0_  ;
  output \g61807/_0_  ;
  output \g61808/_0_  ;
  output \g61809/_0_  ;
  output \g61810/_0_  ;
  output \g61811/_0_  ;
  output \g61812/_0_  ;
  output \g61813/_0_  ;
  output \g61816/_0_  ;
  output \g61817/_0_  ;
  output \g61818/_0_  ;
  output \g61820/_0_  ;
  output \g61822/_0_  ;
  output \g61823/_0_  ;
  output \g61825/_0_  ;
  output \g61826/_0_  ;
  output \g61827/_0_  ;
  output \g61828/_0_  ;
  output \g61829/_0_  ;
  output \g61832/_0_  ;
  output \g61834/_0_  ;
  output \g61835/_0_  ;
  output \g61837/_0_  ;
  output \g61838/_0_  ;
  output \g61839/_0_  ;
  output \g61840/_0_  ;
  output \g61844/_0_  ;
  output \g61847/_0_  ;
  output \g61848/_0_  ;
  output \g61849/_0_  ;
  output \g61850/_0_  ;
  output \g61851/_0_  ;
  output \g61853/_0_  ;
  output \g61854/_0_  ;
  output \g61855/_0_  ;
  output \g61856/_0_  ;
  output \g61858/_0_  ;
  output \g61859/_0_  ;
  output \g61861/_0_  ;
  output \g61862/_0_  ;
  output \g61863/_0_  ;
  output \g61864/_0_  ;
  output \g61865/_0_  ;
  output \g61866/_0_  ;
  output \g61867/_0_  ;
  output \g61868/_0_  ;
  output \g61869/_0_  ;
  output \g61870/_0_  ;
  output \g61871/_0_  ;
  output \g61873/_0_  ;
  output \g61874/_0_  ;
  output \g61875/_0_  ;
  output \g61877/_0_  ;
  output \g61878/_0_  ;
  output \g61879/_0_  ;
  output \g61880/_0_  ;
  output \g61881/_0_  ;
  output \g61883/_0_  ;
  output \g61884/_0_  ;
  output \g61886/_0_  ;
  output \g61887/_0_  ;
  output \g61890/_0_  ;
  output \g61891/_0_  ;
  output \g61892/_0_  ;
  output \g61893/_0_  ;
  output \g61894/_0_  ;
  output \g61895/_0_  ;
  output \g61900/_0_  ;
  output \g61901/_0_  ;
  output \g61902/_0_  ;
  output \g61904/_0_  ;
  output \g61905/_0_  ;
  output \g61906/_0_  ;
  output \g61907/_0_  ;
  output \g61914/_0_  ;
  output \g61915/_0_  ;
  output \g61917/_0_  ;
  output \g61919/_0_  ;
  output \g61921/_0_  ;
  output \g61924/_0_  ;
  output \g61925/_0_  ;
  output \g61926/_0_  ;
  output \g61927/_0_  ;
  output \g61928/_0_  ;
  output \g61929/_0_  ;
  output \g61930/_0_  ;
  output \g61931/_0_  ;
  output \g61932/_0_  ;
  output \g61933/_0_  ;
  output \g61934/_0_  ;
  output \g61935/_0_  ;
  output \g61936/_0_  ;
  output \g61937/_0_  ;
  output \g61938/_0_  ;
  output \g61939/_0_  ;
  output \g61943/_0_  ;
  output \g61944/_0_  ;
  output \g61945/_0_  ;
  output \g61947/_0_  ;
  output \g61948/_0_  ;
  output \g61949/_0_  ;
  output \g61950/_0_  ;
  output \g61951/_0_  ;
  output \g61952/_0_  ;
  output \g61953/_0_  ;
  output \g61955/_0_  ;
  output \g61956/_0_  ;
  output \g61957/_0_  ;
  output \g61958/_0_  ;
  output \g61959/_0_  ;
  output \g61960/_0_  ;
  output \g61961/_0_  ;
  output \g61962/_0_  ;
  output \g61963/_0_  ;
  output \g61964/_0_  ;
  output \g61965/_0_  ;
  output \g61966/_0_  ;
  output \g61967/_0_  ;
  output \g61968/_0_  ;
  output \g61969/_0_  ;
  output \g61970/_0_  ;
  output \g61971/_0_  ;
  output \g61972/_0_  ;
  output \g61973/_0_  ;
  output \g61974/_0_  ;
  output \g61976/_0_  ;
  output \g61978/_0_  ;
  output \g61980/_0_  ;
  output \g61981/_0_  ;
  output \g61982/_0_  ;
  output \g61983/_0_  ;
  output \g61984/_0_  ;
  output \g61985/_0_  ;
  output \g61986/_0_  ;
  output \g61987/_0_  ;
  output \g61988/_0_  ;
  output \g61989/_0_  ;
  output \g61990/_0_  ;
  output \g61992/_0_  ;
  output \g61994/_0_  ;
  output \g61995/_0_  ;
  output \g61996/_0_  ;
  output \g61997/_0_  ;
  output \g61998/_0_  ;
  output \g62000/_0_  ;
  output \g62001/_0_  ;
  output \g62002/_0_  ;
  output \g62003/_0_  ;
  output \g62004/_0_  ;
  output \g62005/_0_  ;
  output \g62007/_0_  ;
  output \g62008/_0_  ;
  output \g62009/_0_  ;
  output \g62010/_0_  ;
  output \g62011/_0_  ;
  output \g62012/_0_  ;
  output \g62013/_0_  ;
  output \g62014/_0_  ;
  output \g62015/_0_  ;
  output \g62016/_0_  ;
  output \g62017/_0_  ;
  output \g62018/_0_  ;
  output \g62019/_0_  ;
  output \g62020/_0_  ;
  output \g62021/_0_  ;
  output \g62022/_0_  ;
  output \g62023/_0_  ;
  output \g62024/_0_  ;
  output \g62025/_0_  ;
  output \g62026/_0_  ;
  output \g62027/_0_  ;
  output \g62030/_0_  ;
  output \g62033/_0_  ;
  output \g62034/_0_  ;
  output \g62036/_0_  ;
  output \g62038/_0_  ;
  output \g62041/_0_  ;
  output \g62042/_0_  ;
  output \g62043/_0_  ;
  output \g62044/_0_  ;
  output \g62045/_0_  ;
  output \g62046/_0_  ;
  output \g62047/_0_  ;
  output \g62048/_0_  ;
  output \g62050/_0_  ;
  output \g62051/_0_  ;
  output \g62052/_0_  ;
  output \g62055/_0_  ;
  output \g62057/_0_  ;
  output \g62058/_0_  ;
  output \g62059/_0_  ;
  output \g62060/_0_  ;
  output \g62061/_0_  ;
  output \g62062/_0_  ;
  output \g62064/_0_  ;
  output \g62065/_0_  ;
  output \g62066/_0_  ;
  output \g62067/_0_  ;
  output \g62068/_0_  ;
  output \g62072/_0_  ;
  output \g62073/_0_  ;
  output \g62074/_0_  ;
  output \g62075/_0_  ;
  output \g62076/_0_  ;
  output \g62077/_0_  ;
  output \g62078/_0_  ;
  output \g62080/_0_  ;
  output \g62081/_0_  ;
  output \g62082/_0_  ;
  output \g62084/_0_  ;
  output \g62085/_0_  ;
  output \g62086/_0_  ;
  output \g62087/_0_  ;
  output \g62088/_0_  ;
  output \g62089/_0_  ;
  output \g62090/_0_  ;
  output \g62091/_0_  ;
  output \g62092/_0_  ;
  output \g62094/_0_  ;
  output \g62096/_0_  ;
  output \g62097/_0_  ;
  output \g62098/_0_  ;
  output \g62099/_0_  ;
  output \g62100/_0_  ;
  output \g62101/_0_  ;
  output \g62102/_0_  ;
  output \g62104/_0_  ;
  output \g62106/_0_  ;
  output \g62107/_0_  ;
  output \g62108/_0_  ;
  output \g62110/_0_  ;
  output \g62112/_0_  ;
  output \g62113/_0_  ;
  output \g62114/_0_  ;
  output \g62116/_0_  ;
  output \g62117/_0_  ;
  output \g62118/_0_  ;
  output \g62119/_0_  ;
  output \g62120/_0_  ;
  output \g62121/_0_  ;
  output \g62122/_0_  ;
  output \g62124/_0_  ;
  output \g62126/_0_  ;
  output \g62127/_0_  ;
  output \g62128/_0_  ;
  output \g62129/_0_  ;
  output \g62130/_0_  ;
  output \g62131/_0_  ;
  output \g62132/_0_  ;
  output \g62133/_0_  ;
  output \g62135/_0_  ;
  output \g62136/_0_  ;
  output \g62137/_0_  ;
  output \g62138/_0_  ;
  output \g62140/_0_  ;
  output \g62143/_0_  ;
  output \g62144/_0_  ;
  output \g62149/_0_  ;
  output \g62150/_0_  ;
  output \g62151/_0_  ;
  output \g62153/_0_  ;
  output \g62155/_0_  ;
  output \g62156/_0_  ;
  output \g62158/_0_  ;
  output \g62160/_0_  ;
  output \g62161/_0_  ;
  output \g62162/_0_  ;
  output \g62164/_0_  ;
  output \g62165/_0_  ;
  output \g62166/_0_  ;
  output \g62167/_0_  ;
  output \g62168/_0_  ;
  output \g62169/_0_  ;
  output \g62172/_0_  ;
  output \g62173/_0_  ;
  output \g62175/_0_  ;
  output \g62176/_0_  ;
  output \g62177/_0_  ;
  output \g62178/_0_  ;
  output \g62179/_0_  ;
  output \g62180/_0_  ;
  output \g62181/_0_  ;
  output \g62182/_0_  ;
  output \g62183/_0_  ;
  output \g62184/_0_  ;
  output \g62185/_0_  ;
  output \g62186/_0_  ;
  output \g62188/_0_  ;
  output \g62189/_0_  ;
  output \g62190/_0_  ;
  output \g62191/_0_  ;
  output \g62193/_0_  ;
  output \g62194/_0_  ;
  output \g62195/_0_  ;
  output \g62196/_0_  ;
  output \g62197/_0_  ;
  output \g62200/_0_  ;
  output \g62201/_0_  ;
  output \g62202/_0_  ;
  output \g62203/_0_  ;
  output \g62205/_0_  ;
  output \g62206/_0_  ;
  output \g62207/_0_  ;
  output \g62208/_0_  ;
  output \g62209/_0_  ;
  output \g62210/_0_  ;
  output \g62211/_0_  ;
  output \g62215/_0_  ;
  output \g62218/_0_  ;
  output \g62219/_0_  ;
  output \g62221/_0_  ;
  output \g62222/_0_  ;
  output \g62223/_0_  ;
  output \g62224/_0_  ;
  output \g62225/_0_  ;
  output \g62226/_0_  ;
  output \g62229/_0_  ;
  output \g62230/_0_  ;
  output \g62231/_0_  ;
  output \g62233/_0_  ;
  output \g62236/_0_  ;
  output \g62237/_0_  ;
  output \g62238/_0_  ;
  output \g62240/_0_  ;
  output \g62241/_0_  ;
  output \g62243/_0_  ;
  output \g62244/_0_  ;
  output \g62245/_0_  ;
  output \g62247/_0_  ;
  output \g62248/_0_  ;
  output \g62250/_0_  ;
  output \g62252/_0_  ;
  output \g62253/_0_  ;
  output \g62255/_0_  ;
  output \g62256/_0_  ;
  output \g62257/_0_  ;
  output \g62258/_0_  ;
  output \g62259/_0_  ;
  output \g62260/_0_  ;
  output \g62261/_0_  ;
  output \g62262/_0_  ;
  output \g62263/_0_  ;
  output \g62264/_0_  ;
  output \g62265/_0_  ;
  output \g62267/_0_  ;
  output \g62269/_0_  ;
  output \g62270/_0_  ;
  output \g62272/_0_  ;
  output \g62274/_0_  ;
  output \g62277/_0_  ;
  output \g62279/_0_  ;
  output \g62280/_0_  ;
  output \g62281/_0_  ;
  output \g62283/_0_  ;
  output \g62284/_0_  ;
  output \g62285/_0_  ;
  output \g62286/_0_  ;
  output \g62288/_0_  ;
  output \g62289/_0_  ;
  output \g62290/_0_  ;
  output \g62294/_0_  ;
  output \g62295/_0_  ;
  output \g62296/_0_  ;
  output \g62297/_0_  ;
  output \g62298/_0_  ;
  output \g62299/_0_  ;
  output \g62303/_0_  ;
  output \g62305/_0_  ;
  output \g62306/_0_  ;
  output \g62307/_0_  ;
  output \g62309/_0_  ;
  output \g62311/_0_  ;
  output \g62312/_0_  ;
  output \g62313/_0_  ;
  output \g62314/_0_  ;
  output \g62315/_0_  ;
  output \g62316/_0_  ;
  output \g62317/_0_  ;
  output \g62318/_0_  ;
  output \g62319/_0_  ;
  output \g62320/_0_  ;
  output \g62322/_0_  ;
  output \g62324/_0_  ;
  output \g62325/_0_  ;
  output \g62326/_0_  ;
  output \g62327/_0_  ;
  output \g62329/_0_  ;
  output \g62330/_0_  ;
  output \g62331/_0_  ;
  output \g62332/_0_  ;
  output \g62333/_0_  ;
  output \g62335/_0_  ;
  output \g62336/_0_  ;
  output \g62338/_0_  ;
  output \g62341/_0_  ;
  output \g62342/_0_  ;
  output \g62344/_0_  ;
  output \g62345/_0_  ;
  output \g62348/_0_  ;
  output \g62349/_0_  ;
  output \g62350/_0_  ;
  output \g62353/_0_  ;
  output \g62354/_0_  ;
  output \g62355/_0_  ;
  output \g62356/_0_  ;
  output \g62359/_0_  ;
  output \g62362/_0_  ;
  output \g62363/_0_  ;
  output \g62364/_0_  ;
  output \g62365/_0_  ;
  output \g62366/_0_  ;
  output \g62367/_0_  ;
  output \g62368/_0_  ;
  output \g62369/_0_  ;
  output \g62370/_0_  ;
  output \g62371/_0_  ;
  output \g62372/_0_  ;
  output \g62373/_0_  ;
  output \g62374/_0_  ;
  output \g62376/_0_  ;
  output \g62467/_0_  ;
  output \g62468/_0_  ;
  output \g62469/_0_  ;
  output \g62470/_0_  ;
  output \g62471/_0_  ;
  output \g62472/_0_  ;
  output \g62473/_0_  ;
  output \g62474/_0_  ;
  output \g62475/_0_  ;
  output \g62478/_0_  ;
  output \g62480/_0_  ;
  output \g62481/_0_  ;
  output \g62482/_0_  ;
  output \g62483/_0_  ;
  output \g62484/_0_  ;
  output \g62485/_0_  ;
  output \g62486/_0_  ;
  output \g62487/_0_  ;
  output \g62488/_0_  ;
  output \g62489/_0_  ;
  output \g62490/_0_  ;
  output \g62491/_0_  ;
  output \g62492/_0_  ;
  output \g62493/_0_  ;
  output \g62494/_0_  ;
  output \g62495/_0_  ;
  output \g62496/_0_  ;
  output \g62497/_0_  ;
  output \g62498/_0_  ;
  output \g62499/_0_  ;
  output \g62500/_0_  ;
  output \g62501/_0_  ;
  output \g62502/_0_  ;
  output \g62503/_0_  ;
  output \g62504/_0_  ;
  output \g62509/_0_  ;
  output \g62510/_0_  ;
  output \g62511/_0_  ;
  output \g62512/_0_  ;
  output \g62513/_0_  ;
  output \g62514/_0_  ;
  output \g62515/_0_  ;
  output \g62516/_0_  ;
  output \g62517/_0_  ;
  output \g62518/_0_  ;
  output \g62519/_0_  ;
  output \g62520/_0_  ;
  output \g62521/_0_  ;
  output \g62523/_0_  ;
  output \g62526/_0_  ;
  output \g62528/_0_  ;
  output \g62529/_0_  ;
  output \g62531/_0_  ;
  output \g62532/_0_  ;
  output \g62533/_0_  ;
  output \g62534/_0_  ;
  output \g62535/_0_  ;
  output \g62536/_0_  ;
  output \g62537/_0_  ;
  output \g62539/_0_  ;
  output \g62540/_0_  ;
  output \g62541/_0_  ;
  output \g62542/_0_  ;
  output \g62543/_0_  ;
  output \g62544/_0_  ;
  output \g62545/_0_  ;
  output \g62547/_0_  ;
  output \g62548/_0_  ;
  output \g62549/_0_  ;
  output \g62550/_0_  ;
  output \g62551/_0_  ;
  output \g62552/_0_  ;
  output \g62553/_0_  ;
  output \g62554/_0_  ;
  output \g62555/_0_  ;
  output \g62556/_0_  ;
  output \g62557/_0_  ;
  output \g62560/_0_  ;
  output \g62562/_0_  ;
  output \g62563/_0_  ;
  output \g62564/_0_  ;
  output \g62565/_0_  ;
  output \g62566/_0_  ;
  output \g62567/_0_  ;
  output \g62569/_0_  ;
  output \g62570/_0_  ;
  output \g62571/_0_  ;
  output \g62572/_0_  ;
  output \g62573/_0_  ;
  output \g62574/_0_  ;
  output \g62576/_0_  ;
  output \g62577/_0_  ;
  output \g62581/_0_  ;
  output \g62582/_0_  ;
  output \g62584/_0_  ;
  output \g62585/_0_  ;
  output \g62586/_0_  ;
  output \g62588/_0_  ;
  output \g62589/_0_  ;
  output \g62593/_0_  ;
  output \g62594/_0_  ;
  output \g62595/_0_  ;
  output \g62596/_0_  ;
  output \g62597/_0_  ;
  output \g62598/_0_  ;
  output \g62599/_0_  ;
  output \g62600/_0_  ;
  output \g62601/_0_  ;
  output \g62602/_0_  ;
  output \g62603/_0_  ;
  output \g62604/_0_  ;
  output \g62605/_0_  ;
  output \g62606/_0_  ;
  output \g62607/_0_  ;
  output \g62608/_0_  ;
  output \g62609/_0_  ;
  output \g62610/_0_  ;
  output \g62612/_0_  ;
  output \g62613/_0_  ;
  output \g62614/_0_  ;
  output \g62615/_0_  ;
  output \g62617/_0_  ;
  output \g62618/_0_  ;
  output \g62620/_0_  ;
  output \g62621/_0_  ;
  output \g62622/_0_  ;
  output \g62624/_0_  ;
  output \g62625/_0_  ;
  output \g62626/_0_  ;
  output \g62627/_0_  ;
  output \g62629/_0_  ;
  output \g62630/_0_  ;
  output \g62632/_0_  ;
  output \g62633/_0_  ;
  output \g62635/_0_  ;
  output \g62636/_0_  ;
  output \g62637/_0_  ;
  output \g62638/_0_  ;
  output \g62640/_0_  ;
  output \g62641/_0_  ;
  output \g62642/_0_  ;
  output \g62643/_0_  ;
  output \g62644/_0_  ;
  output \g62646/_0_  ;
  output \g62647/_0_  ;
  output \g62649/_0_  ;
  output \g62650/_0_  ;
  output \g62651/_0_  ;
  output \g62653/_0_  ;
  output \g62655/_0_  ;
  output \g62656/_0_  ;
  output \g62657/_0_  ;
  output \g62658/_0_  ;
  output \g62660/_0_  ;
  output \g62661/_0_  ;
  output \g62662/_0_  ;
  output \g62663/_0_  ;
  output \g62664/_0_  ;
  output \g62665/_0_  ;
  output \g62667/_0_  ;
  output \g62669/_0_  ;
  output \g62670/_0_  ;
  output \g62671/_0_  ;
  output \g62672/_0_  ;
  output \g62674/_0_  ;
  output \g62675/_0_  ;
  output \g62676/_0_  ;
  output \g62677/_0_  ;
  output \g62678/_0_  ;
  output \g62679/_0_  ;
  output \g62680/_0_  ;
  output \g62681/_0_  ;
  output \g62682/_0_  ;
  output \g62684/_0_  ;
  output \g62685/_0_  ;
  output \g62686/_0_  ;
  output \g62687/_0_  ;
  output \g62690/_0_  ;
  output \g62693/_0_  ;
  output \g62698/_0_  ;
  output \g62699/_0_  ;
  output \g62700/_0_  ;
  output \g62701/_0_  ;
  output \g62702/_0_  ;
  output \g62703/_0_  ;
  output \g62704/_0_  ;
  output \g62709/_0_  ;
  output \g62710/_0_  ;
  output \g62711/_0_  ;
  output \g62714/_0_  ;
  output \g62715/_0_  ;
  output \g62717/_0_  ;
  output \g62718/_0_  ;
  output \g62719/_0_  ;
  output \g62720/_0_  ;
  output \g62721/_0_  ;
  output \g62723/_0_  ;
  output \g62725/_0_  ;
  output \g62726/_0_  ;
  output \g62729/_0_  ;
  output \g62731/_0_  ;
  output \g62733/_0_  ;
  output \g62738/_0_  ;
  output \g62741/_0_  ;
  output \g62742/_0_  ;
  output \g62744/_0_  ;
  output \g62745/_0_  ;
  output \g62746/_0_  ;
  output \g62747/_0_  ;
  output \g62748/_0_  ;
  output \g62749/_0_  ;
  output \g62753/_0_  ;
  output \g62755/_0_  ;
  output \g62756/_0_  ;
  output \g62758/_0_  ;
  output \g62759/_0_  ;
  output \g62760/_0_  ;
  output \g62761/_0_  ;
  output \g62763/_0_  ;
  output \g62766/_0_  ;
  output \g62767/_0_  ;
  output \g62768/_0_  ;
  output \g65554/_0_  ;
  output \g65561/_0_  ;
  output \g65569/_0_  ;
  output \g65580/_0_  ;
  output \g65599/_0_  ;
  output \g65606/_0_  ;
  output \g65636/_0_  ;
  output \g65864/_0_  ;
  wire n1508 , n1509 , n1510 , n1511 , n1512 , n1513 , n1514 , n1515 , n1516 , n1517 , n1518 , n1519 , n1520 , n1521 , n1522 , n1523 , n1524 , n1525 , n1526 , n1527 , n1528 , n1529 , n1530 , n1531 , n1532 , n1533 , n1534 , n1535 , n1536 , n1537 , n1538 , n1539 , n1540 , n1541 , n1542 , n1543 , n1544 , n1545 , n1546 , n1547 , n1548 , n1549 , n1550 , n1551 , n1552 , n1553 , n1554 , n1555 , n1556 , n1557 , n1558 , n1559 , n1560 , n1561 , n1562 , n1563 , n1564 , n1565 , n1566 , n1567 , n1568 , n1569 , n1570 , n1571 , n1572 , n1573 , n1574 , n1575 , n1576 , n1577 , n1578 , n1579 , n1580 , n1581 , n1582 , n1583 , n1584 , n1585 , n1586 , n1587 , n1588 , n1589 , n1590 , n1591 , n1592 , n1593 , n1594 , n1595 , n1596 , n1597 , n1598 , n1599 , n1600 , n1601 , n1602 , n1603 , n1604 , n1605 , n1606 , n1607 , n1608 , n1609 , n1610 , n1611 , n1612 , n1613 , n1614 , n1615 , n1616 , n1617 , n1618 , n1619 , n1620 , n1621 , n1622 , n1623 , n1624 , n1625 , n1626 , n1627 , n1628 , n1629 , n1630 , n1631 , n1632 , n1633 , n1634 , n1635 , n1636 , n1637 , n1638 , n1639 , n1640 , n1641 , n1642 , n1643 , n1644 , n1645 , n1646 , n1647 , n1648 , n1649 , n1650 , n1651 , n1652 , n1653 , n1654 , n1655 , n1656 , n1657 , n1658 , n1659 , n1660 , n1661 , n1662 , n1663 , n1664 , n1665 , n1666 , n1667 , n1668 , n1669 , n1670 , n1671 , n1672 , n1673 , n1674 , n1675 , n1676 , n1677 , n1678 , n1679 , n1680 , n1681 , n1682 , n1683 , n1684 , n1685 , n1686 , n1687 , n1688 , n1689 , n1690 , n1691 , n1692 , n1693 , n1694 , n1695 , n1696 , n1697 , n1698 , n1699 , n1700 , n1701 , n1702 , n1703 , n1704 , n1705 , n1706 , n1707 , n1708 , n1709 , n1710 , n1711 , n1712 , n1713 , n1714 , n1715 , n1716 , n1717 , n1718 , n1719 , n1720 , n1721 , n1722 , n1723 , n1724 , n1725 , n1726 , n1727 , n1728 , n1729 , n1730 , n1731 , n1732 , n1733 , n1734 , n1735 , n1736 , n1737 , n1738 , n1739 , n1740 , n1741 , n1742 , n1743 , n1744 , n1745 , n1746 , n1747 , n1748 , n1749 , n1750 , n1751 , n1752 , n1753 , n1754 , n1755 , n1756 , n1757 , n1758 , n1759 , n1760 , n1761 , n1762 , n1763 , n1764 , n1765 , n1766 , n1767 , n1768 , n1769 , n1770 , n1771 , n1772 , n1773 , n1774 , n1775 , n1776 , n1777 , n1778 , n1779 , n1780 , n1781 , n1782 , n1783 , n1784 , n1785 , n1786 , n1787 , n1788 , n1789 , n1790 , n1791 , n1792 , n1793 , n1794 , n1795 , n1796 , n1797 , n1798 , n1799 , n1800 , n1801 , n1802 , n1803 , n1804 , n1805 , n1806 , n1807 , n1808 , n1809 , n1810 , n1811 , n1812 , n1813 , n1814 , n1815 , n1816 , n1817 , n1818 , n1819 , n1820 , n1821 , n1822 , n1823 , n1824 , n1825 , n1826 , n1827 , n1828 , n1829 , n1830 , n1831 , n1832 , n1833 , n1834 , n1835 , n1836 , n1837 , n1838 , n1839 , n1840 , n1841 , n1842 , n1843 , n1844 , n1845 , n1846 , n1847 , n1848 , n1849 , n1850 , n1851 , n1852 , n1853 , n1854 , n1855 , n1856 , n1857 , n1858 , n1859 , n1860 , n1861 , n1862 , n1863 , n1864 , n1865 , n1866 , n1867 , n1868 , n1869 , n1870 , n1871 , n1872 , n1873 , n1874 , n1875 , n1876 , n1877 , n1878 , n1879 , n1880 , n1881 , n1882 , n1883 , n1884 , n1885 , n1886 , n1887 , n1888 , n1889 , n1890 , n1891 , n1892 , n1893 , n1894 , n1895 , n1896 , n1897 , n1898 , n1899 , n1900 , n1901 , n1902 , n1903 , n1904 , n1905 , n1906 , n1907 , n1908 , n1909 , n1910 , n1911 , n1912 , n1913 , n1914 , n1915 , n1916 , n1917 , n1918 , n1919 , n1920 , n1921 , n1922 , n1923 , n1924 , n1925 , n1926 , n1927 , n1928 , n1929 , n1930 , n1931 , n1932 , n1933 , n1934 , n1935 , n1936 , n1937 , n1938 , n1939 , n1940 , n1941 , n1942 , n1943 , n1944 , n1945 , n1946 , n1947 , n1948 , n1949 , n1950 , n1951 , n1952 , n1953 , n1954 , n1955 , n1956 , n1957 , n1958 , n1959 , n1960 , n1961 , n1962 , n1963 , n1964 , n1965 , n1966 , n1967 , n1968 , n1969 , n1970 , n1971 , n1972 , n1973 , n1974 , n1975 , n1976 , n1977 , n1978 , n1979 , n1980 , n1981 , n1982 , n1983 , n1984 , n1985 , n1986 , n1987 , n1988 , n1989 , n1990 , n1991 , n1992 , n1993 , n1994 , n1995 , n1996 , n1997 , n1998 , n1999 , n2000 , n2001 , n2002 , n2003 , n2004 , n2005 , n2006 , n2007 , n2008 , n2009 , n2010 , n2011 , n2012 , n2013 , n2014 , n2015 , n2016 , n2017 , n2018 , n2019 , n2020 , n2021 , n2022 , n2023 , n2024 , n2025 , n2026 , n2027 , n2028 , n2029 , n2030 , n2031 , n2032 , n2033 , n2034 , n2035 , n2036 , n2037 , n2038 , n2039 , n2040 , n2041 , n2042 , n2043 , n2044 , n2045 , n2046 , n2047 , n2048 , n2049 , n2050 , n2051 , n2052 , n2053 , n2054 , n2055 , n2056 , n2057 , n2058 , n2059 , n2060 , n2061 , n2062 , n2063 , n2064 , n2065 , n2066 , n2067 , n2068 , n2069 , n2070 , n2071 , n2072 , n2073 , n2074 , n2075 , n2076 , n2077 , n2078 , n2079 , n2080 , n2081 , n2082 , n2083 , n2084 , n2085 , n2086 , n2087 , n2088 , n2089 , n2090 , n2091 , n2092 , n2093 , n2094 , n2095 , n2096 , n2097 , n2098 , n2099 , n2100 , n2101 , n2102 , n2103 , n2104 , n2105 , n2106 , n2107 , n2108 , n2109 , n2110 , n2111 , n2112 , n2113 , n2114 , n2115 , n2116 , n2117 , n2118 , n2119 , n2120 , n2121 , n2122 , n2123 , n2124 , n2125 , n2126 , n2127 , n2128 , n2129 , n2130 , n2131 , n2132 , n2133 , n2134 , n2135 , n2136 , n2137 , n2138 , n2139 , n2140 , n2141 , n2142 , n2143 , n2144 , n2145 , n2146 , n2147 , n2148 , n2149 , n2150 , n2151 , n2152 , n2153 , n2154 , n2155 , n2156 , n2157 , n2158 , n2159 , n2160 , n2161 , n2162 , n2163 , n2164 , n2165 , n2166 , n2167 , n2168 , n2169 , n2170 , n2171 , n2172 , n2173 , n2174 , n2175 , n2176 , n2177 , n2178 , n2179 , n2180 , n2181 , n2182 , n2183 , n2184 , n2185 , n2186 , n2187 , n2188 , n2189 , n2190 , n2191 , n2192 , n2193 , n2194 , n2195 , n2196 , n2197 , n2198 , n2199 , n2200 , n2201 , n2202 , n2203 , n2204 , n2205 , n2206 , n2207 , n2208 , n2209 , n2210 , n2211 , n2212 , n2213 , n2214 , n2215 , n2216 , n2217 , n2218 , n2219 , n2220 , n2221 , n2222 , n2223 , n2224 , n2225 , n2226 , n2227 , n2228 , n2229 , n2230 , n2231 , n2232 , n2233 , n2234 , n2235 , n2236 , n2237 , n2238 , n2239 , n2240 , n2241 , n2242 , n2243 , n2244 , n2245 , n2246 , n2247 , n2248 , n2249 , n2250 , n2251 , n2252 , n2253 , n2254 , n2255 , n2256 , n2257 , n2258 , n2259 , n2260 , n2261 , n2262 , n2263 , n2264 , n2265 , n2266 , n2267 , n2268 , n2269 , n2270 , n2271 , n2272 , n2273 , n2274 , n2275 , n2276 , n2277 , n2278 , n2279 , n2280 , n2281 , n2282 , n2283 , n2284 , n2285 , n2286 , n2287 , n2288 , n2289 , n2290 , n2291 , n2292 , n2293 , n2294 , n2295 , n2296 , n2297 , n2298 , n2299 , n2300 , n2301 , n2302 , n2303 , n2304 , n2305 , n2306 , n2307 , n2308 , n2309 , n2310 , n2311 , n2312 , n2313 , n2314 , n2315 , n2316 , n2317 , n2318 , n2319 , n2320 , n2321 , n2322 , n2323 , n2324 , n2325 , n2326 , n2327 , n2328 , n2329 , n2330 , n2331 , n2332 , n2333 , n2334 , n2335 , n2336 , n2337 , n2338 , n2339 , n2340 , n2341 , n2342 , n2343 , n2344 , n2345 , n2346 , n2347 , n2348 , n2349 , n2350 , n2351 , n2352 , n2353 , n2354 , n2355 , n2356 , n2357 , n2358 , n2359 , n2360 , n2361 , n2362 , n2363 , n2364 , n2365 , n2366 , n2367 , n2368 , n2369 , n2370 , n2371 , n2372 , n2373 , n2374 , n2375 , n2376 , n2377 , n2378 , n2379 , n2380 , n2381 , n2382 , n2383 , n2384 , n2385 , n2386 , n2387 , n2388 , n2389 , n2390 , n2391 , n2392 , n2393 , n2394 , n2395 , n2396 , n2397 , n2398 , n2399 , n2400 , n2401 , n2402 , n2403 , n2404 , n2405 , n2406 , n2407 , n2408 , n2409 , n2410 , n2411 , n2412 , n2413 , n2414 , n2415 , n2416 , n2417 , n2418 , n2419 , n2420 , n2421 , n2422 , n2423 , n2424 , n2425 , n2426 , n2427 , n2428 , n2429 , n2430 , n2431 , n2432 , n2433 , n2434 , n2435 , n2436 , n2437 , n2438 , n2439 , n2440 , n2441 , n2442 , n2443 , n2444 , n2445 , n2446 , n2447 , n2448 , n2449 , n2450 , n2451 , n2452 , n2453 , n2454 , n2455 , n2456 , n2457 , n2458 , n2459 , n2460 , n2461 , n2462 , n2463 , n2464 , n2465 , n2466 , n2467 , n2468 , n2469 , n2470 , n2471 , n2472 , n2473 , n2474 , n2475 , n2476 , n2477 , n2478 , n2479 , n2480 , n2481 , n2482 , n2483 , n2484 , n2485 , n2486 , n2487 , n2488 , n2489 , n2490 , n2491 , n2492 , n2493 , n2494 , n2495 , n2496 , n2497 , n2498 , n2499 , n2500 , n2501 , n2502 , n2503 , n2504 , n2505 , n2506 , n2507 , n2508 , n2509 , n2510 , n2511 , n2512 , n2513 , n2514 , n2515 , n2516 , n2517 , n2518 , n2519 , n2520 , n2521 , n2522 , n2523 , n2524 , n2525 , n2526 , n2527 , n2528 , n2529 , n2530 , n2531 , n2532 , n2533 , n2534 , n2535 , n2536 , n2537 , n2538 , n2539 , n2540 , n2541 , n2542 , n2543 , n2544 , n2545 , n2546 , n2547 , n2548 , n2549 , n2550 , n2551 , n2552 , n2553 , n2554 , n2555 , n2556 , n2557 , n2558 , n2559 , n2560 , n2561 , n2562 , n2563 , n2564 , n2565 , n2566 , n2567 , n2568 , n2569 , n2570 , n2571 , n2572 , n2573 , n2574 , n2575 , n2576 , n2577 , n2578 , n2579 , n2580 , n2581 , n2582 , n2583 , n2584 , n2585 , n2586 , n2587 , n2588 , n2589 , n2590 , n2591 , n2592 , n2593 , n2594 , n2595 , n2596 , n2597 , n2598 , n2599 , n2600 , n2601 , n2602 , n2603 , n2604 , n2605 , n2606 , n2607 , n2608 , n2609 , n2610 , n2611 , n2612 , n2613 , n2614 , n2615 , n2616 , n2617 , n2618 , n2619 , n2620 , n2621 , n2622 , n2623 , n2624 , n2625 , n2626 , n2627 , n2628 , n2629 , n2630 , n2631 , n2632 , n2633 , n2634 , n2635 , n2636 , n2637 , n2638 , n2639 , n2640 , n2641 , n2642 , n2643 , n2644 , n2645 , n2646 , n2647 , n2648 , n2649 , n2650 , n2651 , n2652 , n2653 , n2654 , n2655 , n2656 , n2657 , n2658 , n2659 , n2660 , n2661 , n2662 , n2663 , n2664 , n2665 , n2666 , n2667 , n2668 , n2669 , n2670 , n2671 , n2672 , n2673 , n2674 , n2675 , n2676 , n2677 , n2678 , n2679 , n2680 , n2681 , n2682 , n2683 , n2684 , n2685 , n2686 , n2687 , n2688 , n2689 , n2690 , n2691 , n2692 , n2693 , n2694 , n2695 , n2696 , n2697 , n2698 , n2699 , n2700 , n2701 , n2702 , n2703 , n2704 , n2705 , n2706 , n2707 , n2708 , n2709 , n2710 , n2711 , n2712 , n2713 , n2714 , n2715 , n2716 , n2717 , n2718 , n2719 , n2720 , n2721 , n2722 , n2723 , n2724 , n2725 , n2726 , n2727 , n2728 , n2729 , n2730 , n2731 , n2732 , n2733 , n2734 , n2735 , n2736 , n2737 , n2738 , n2739 , n2740 , n2741 , n2742 , n2743 , n2744 , n2745 , n2746 , n2747 , n2748 , n2749 , n2750 , n2751 , n2752 , n2753 , n2754 , n2755 , n2756 , n2757 , n2758 , n2759 , n2760 , n2761 , n2762 , n2763 , n2764 , n2765 , n2766 , n2767 , n2768 , n2769 , n2770 , n2771 , n2772 , n2773 , n2774 , n2775 , n2776 , n2777 , n2778 , n2779 , n2780 , n2781 , n2782 , n2783 , n2784 , n2785 , n2786 , n2787 , n2788 , n2789 , n2790 , n2791 , n2792 , n2793 , n2794 , n2795 , n2796 , n2797 , n2798 , n2799 , n2800 , n2801 , n2802 , n2803 , n2804 , n2805 , n2806 , n2807 , n2808 , n2809 , n2810 , n2811 , n2812 , n2813 , n2814 , n2815 , n2816 , n2817 , n2818 , n2819 , n2820 , n2821 , n2822 , n2823 , n2824 , n2825 , n2826 , n2827 , n2828 , n2829 , n2830 , n2831 , n2832 , n2833 , n2834 , n2835 , n2836 , n2837 , n2838 , n2839 , n2840 , n2841 , n2842 , n2843 , n2844 , n2845 , n2846 , n2847 , n2848 , n2849 , n2850 , n2851 , n2852 , n2853 , n2854 , n2855 , n2856 , n2857 , n2858 , n2859 , n2860 , n2861 , n2862 , n2863 , n2864 , n2865 , n2866 , n2867 , n2868 , n2869 , n2870 , n2871 , n2872 , n2873 , n2874 , n2875 , n2876 , n2877 , n2878 , n2879 , n2880 , n2881 , n2882 , n2883 , n2884 , n2885 , n2886 , n2887 , n2888 , n2889 , n2890 , n2891 , n2892 , n2893 , n2894 , n2895 , n2896 , n2897 , n2898 , n2899 , n2900 , n2901 , n2902 , n2903 , n2904 , n2905 , n2906 , n2907 , n2908 , n2909 , n2910 , n2911 , n2912 , n2913 , n2914 , n2915 , n2916 , n2917 , n2918 , n2919 , n2920 , n2921 , n2922 , n2923 , n2924 , n2925 , n2926 , n2927 , n2928 , n2929 , n2930 , n2931 , n2932 , n2933 , n2934 , n2935 , n2936 , n2937 , n2938 , n2939 , n2940 , n2941 , n2942 , n2943 , n2944 , n2945 , n2946 , n2947 , n2948 , n2949 , n2950 , n2951 , n2952 , n2953 , n2954 , n2955 , n2956 , n2957 , n2958 , n2959 , n2960 , n2961 , n2962 , n2963 , n2964 , n2965 , n2966 , n2967 , n2968 , n2969 , n2970 , n2971 , n2972 , n2973 , n2974 , n2975 , n2976 , n2977 , n2978 , n2979 , n2980 , n2981 , n2982 , n2983 , n2984 , n2985 , n2986 , n2987 , n2988 , n2989 , n2990 , n2991 , n2992 , n2993 , n2994 , n2995 , n2996 , n2997 , n2998 , n2999 , n3000 , n3001 , n3002 , n3003 , n3004 , n3005 , n3006 , n3007 , n3008 , n3009 , n3010 , n3011 , n3012 , n3013 , n3014 , n3015 , n3016 , n3017 , n3018 , n3019 , n3020 , n3021 , n3022 , n3023 , n3024 , n3025 , n3026 , n3027 , n3028 , n3029 , n3030 , n3031 , n3032 , n3033 , n3034 , n3035 , n3036 , n3037 , n3038 , n3039 , n3040 , n3041 , n3042 , n3043 , n3044 , n3045 , n3046 , n3047 , n3048 , n3049 , n3050 , n3051 , n3052 , n3053 , n3054 , n3055 , n3056 , n3057 , n3058 , n3059 , n3060 , n3061 , n3062 , n3063 , n3064 , n3065 , n3066 , n3067 , n3068 , n3069 , n3070 , n3071 , n3072 , n3073 , n3074 , n3075 , n3076 , n3077 , n3078 , n3079 , n3080 , n3081 , n3082 , n3083 , n3084 , n3085 , n3086 , n3087 , n3088 , n3089 , n3090 , n3091 , n3092 , n3093 , n3094 , n3095 , n3096 , n3097 , n3098 , n3099 , n3100 , n3101 , n3102 , n3103 , n3104 , n3105 , n3106 , n3107 , n3108 , n3109 , n3110 , n3111 , n3112 , n3113 , n3114 , n3115 , n3116 , n3117 , n3118 , n3119 , n3120 , n3121 , n3122 , n3123 , n3124 , n3125 , n3126 , n3127 , n3128 , n3129 , n3130 , n3131 , n3132 , n3133 , n3134 , n3135 , n3136 , n3137 , n3138 , n3139 , n3140 , n3141 , n3142 , n3143 , n3144 , n3145 , n3146 , n3147 , n3148 , n3149 , n3150 , n3151 , n3152 , n3153 , n3154 , n3155 , n3156 , n3157 , n3158 , n3159 , n3160 , n3161 , n3162 , n3163 , n3164 , n3165 , n3166 , n3167 , n3168 , n3169 , n3170 , n3171 , n3172 , n3173 , n3174 , n3175 , n3176 , n3177 , n3178 , n3179 , n3180 , n3181 , n3182 , n3183 , n3184 , n3185 , n3186 , n3187 , n3188 , n3189 , n3190 , n3191 , n3192 , n3193 , n3194 , n3195 , n3196 , n3197 , n3198 , n3199 , n3200 , n3201 , n3202 , n3203 , n3204 , n3205 , n3206 , n3207 , n3208 , n3209 , n3210 , n3211 , n3212 , n3213 , n3214 , n3215 , n3216 , n3217 , n3218 , n3219 , n3220 , n3221 , n3222 , n3223 , n3224 , n3225 , n3226 , n3227 , n3228 , n3229 , n3230 , n3231 , n3232 , n3233 , n3234 , n3235 , n3236 , n3237 , n3238 , n3239 , n3240 , n3241 , n3242 , n3243 , n3244 , n3245 , n3246 , n3247 , n3248 , n3249 , n3250 , n3251 , n3252 , n3253 , n3254 , n3255 , n3256 , n3257 , n3258 , n3259 , n3260 , n3261 , n3262 , n3263 , n3264 , n3265 , n3266 , n3267 , n3268 , n3269 , n3270 , n3271 , n3272 , n3273 , n3274 , n3275 , n3276 , n3277 , n3278 , n3279 , n3280 , n3281 , n3282 , n3283 , n3284 , n3285 , n3286 , n3287 , n3288 , n3289 , n3290 , n3291 , n3292 , n3293 , n3294 , n3295 , n3296 , n3297 , n3298 , n3299 , n3300 , n3301 , n3302 , n3303 , n3304 , n3305 , n3306 , n3307 , n3308 , n3309 , n3310 , n3311 , n3312 , n3313 , n3314 , n3315 , n3316 , n3317 , n3318 , n3319 , n3320 , n3321 , n3322 , n3323 , n3324 , n3325 , n3326 , n3327 , n3328 , n3329 , n3330 , n3331 , n3332 , n3333 , n3334 , n3335 , n3336 , n3337 , n3338 , n3339 , n3340 , n3341 , n3342 , n3343 , n3344 , n3345 , n3346 , n3347 , n3348 , n3349 , n3350 , n3351 , n3352 , n3353 , n3354 , n3355 , n3356 , n3357 , n3358 , n3359 , n3360 , n3361 , n3362 , n3363 , n3364 , n3365 , n3366 , n3367 , n3368 , n3369 , n3370 , n3371 , n3372 , n3373 , n3374 , n3375 , n3376 , n3377 , n3378 , n3379 , n3380 , n3381 , n3382 , n3383 , n3384 , n3385 , n3386 , n3387 , n3388 , n3389 , n3390 , n3391 , n3392 , n3393 , n3394 , n3395 , n3396 , n3397 , n3398 , n3399 , n3400 , n3401 , n3402 , n3403 , n3404 , n3405 , n3406 , n3407 , n3408 , n3409 , n3410 , n3411 , n3412 , n3413 , n3414 , n3415 , n3416 , n3417 , n3418 , n3419 , n3420 , n3421 , n3422 , n3423 , n3424 , n3425 , n3426 , n3427 , n3428 , n3429 , n3430 , n3431 , n3432 , n3433 , n3434 , n3435 , n3436 , n3437 , n3438 , n3439 , n3440 , n3441 , n3442 , n3443 , n3444 , n3445 , n3446 , n3447 , n3448 , n3449 , n3450 , n3451 , n3452 , n3453 , n3454 , n3455 , n3456 , n3457 , n3458 , n3459 , n3460 , n3461 , n3462 , n3463 , n3464 , n3465 , n3466 , n3467 , n3468 , n3469 , n3470 , n3471 , n3472 , n3473 , n3474 , n3475 , n3476 , n3477 , n3478 , n3479 , n3480 , n3481 , n3482 , n3483 , n3484 , n3485 , n3486 , n3487 , n3488 , n3489 , n3490 , n3491 , n3492 , n3493 , n3494 , n3495 , n3496 , n3497 , n3498 , n3499 , n3500 , n3501 , n3502 , n3503 , n3504 , n3505 , n3506 , n3507 , n3508 , n3509 , n3510 , n3511 , n3512 , n3513 , n3514 , n3515 , n3516 , n3517 , n3518 , n3519 , n3520 , n3521 , n3522 , n3523 , n3524 , n3525 , n3526 , n3527 , n3528 , n3529 , n3530 , n3531 , n3532 , n3533 , n3534 , n3535 , n3536 , n3537 , n3538 , n3539 , n3540 , n3541 , n3542 , n3543 , n3544 , n3545 , n3546 , n3547 , n3548 , n3549 , n3550 , n3551 , n3552 , n3553 , n3554 , n3555 , n3556 , n3557 , n3558 , n3559 , n3560 , n3561 , n3562 , n3563 , n3564 , n3565 , n3566 , n3567 , n3568 , n3569 , n3570 , n3571 , n3572 , n3573 , n3574 , n3575 , n3576 , n3577 , n3578 , n3579 , n3580 , n3581 , n3582 , n3583 , n3584 , n3585 , n3586 , n3587 , n3588 , n3589 , n3590 , n3591 , n3592 , n3593 , n3594 , n3595 , n3596 , n3597 , n3598 , n3599 , n3600 , n3601 , n3602 , n3603 , n3604 , n3605 , n3606 , n3607 , n3608 , n3609 , n3610 , n3611 , n3612 , n3613 , n3614 , n3615 , n3616 , n3617 , n3618 , n3619 , n3620 , n3621 , n3622 , n3623 , n3624 , n3625 , n3626 , n3627 , n3628 , n3629 , n3630 , n3631 , n3632 , n3633 , n3634 , n3635 , n3636 , n3637 , n3638 , n3639 , n3640 , n3641 , n3642 , n3643 , n3644 , n3645 , n3646 , n3647 , n3648 , n3649 , n3650 , n3651 , n3652 , n3653 , n3654 , n3655 , n3656 , n3657 , n3658 , n3659 , n3660 , n3661 , n3662 , n3663 , n3664 , n3665 , n3666 , n3667 , n3668 , n3669 , n3670 , n3671 , n3672 , n3673 , n3674 , n3675 , n3676 , n3677 , n3678 , n3679 , n3680 , n3681 , n3682 , n3683 , n3684 , n3685 , n3686 , n3687 , n3688 , n3689 , n3690 , n3691 , n3692 , n3693 , n3694 , n3695 , n3696 , n3697 , n3698 , n3699 , n3700 , n3701 , n3702 , n3703 , n3704 , n3705 , n3706 , n3707 , n3708 , n3709 , n3710 , n3711 , n3712 , n3713 , n3714 , n3715 , n3716 , n3717 , n3718 , n3719 , n3720 , n3721 , n3722 , n3723 , n3724 , n3725 , n3726 , n3727 , n3728 , n3729 , n3730 , n3731 , n3732 , n3733 , n3734 , n3735 , n3736 , n3737 , n3738 , n3739 , n3740 , n3741 , n3742 , n3743 , n3744 , n3745 , n3746 , n3747 , n3748 , n3749 , n3750 , n3751 , n3752 , n3753 , n3754 , n3755 , n3756 , n3757 , n3758 , n3759 , n3760 , n3761 , n3762 , n3763 , n3764 , n3765 , n3766 , n3767 , n3768 , n3769 , n3770 , n3771 , n3772 , n3773 , n3774 , n3775 , n3776 , n3777 , n3778 , n3779 , n3780 , n3781 , n3782 , n3783 , n3784 , n3785 , n3786 , n3787 , n3788 , n3789 , n3790 , n3791 , n3792 , n3793 , n3794 , n3795 , n3796 , n3797 , n3798 , n3799 , n3800 , n3801 , n3802 , n3803 , n3804 , n3805 , n3806 , n3807 , n3808 , n3809 , n3810 , n3811 , n3812 , n3813 , n3814 , n3815 , n3816 , n3817 , n3818 , n3819 , n3820 , n3821 , n3822 , n3823 , n3824 , n3825 , n3826 , n3827 , n3828 , n3829 , n3830 , n3831 , n3832 , n3833 , n3834 , n3835 , n3836 , n3837 , n3838 , n3839 , n3840 , n3841 , n3842 , n3843 , n3844 , n3845 , n3846 , n3847 , n3848 , n3849 , n3850 , n3851 , n3852 , n3853 , n3854 , n3855 , n3856 , n3857 , n3858 , n3859 , n3860 , n3861 , n3862 , n3863 , n3864 , n3865 , n3866 , n3867 , n3868 , n3869 , n3870 , n3871 , n3872 , n3873 , n3874 , n3875 , n3876 , n3877 , n3878 , n3879 , n3880 , n3881 , n3882 , n3883 , n3884 , n3885 , n3886 , n3887 , n3888 , n3889 , n3890 , n3891 , n3892 , n3893 , n3894 , n3895 , n3896 , n3897 , n3898 , n3899 , n3900 , n3901 , n3902 , n3903 , n3904 , n3905 , n3906 , n3907 , n3908 , n3909 , n3910 , n3911 , n3912 , n3913 , n3914 , n3915 , n3916 , n3917 , n3918 , n3919 , n3920 , n3921 , n3922 , n3923 , n3924 , n3925 , n3926 , n3927 , n3928 , n3929 , n3930 , n3931 , n3932 , n3933 , n3934 , n3935 , n3936 , n3937 , n3938 , n3939 , n3940 , n3941 , n3942 , n3943 , n3944 , n3945 , n3946 , n3947 , n3948 , n3949 , n3950 , n3951 , n3952 , n3953 , n3954 , n3955 , n3956 , n3957 , n3958 , n3959 , n3960 , n3961 , n3962 , n3963 , n3964 , n3965 , n3966 , n3967 , n3968 , n3969 , n3970 , n3971 , n3972 , n3973 , n3974 , n3975 , n3976 , n3977 , n3978 , n3979 , n3980 , n3981 , n3982 , n3983 , n3984 , n3985 , n3986 , n3987 , n3988 , n3989 , n3990 , n3991 , n3992 , n3993 , n3994 , n3995 , n3996 , n3997 , n3998 , n3999 , n4000 , n4001 , n4002 , n4003 , n4004 , n4005 , n4006 , n4007 , n4008 , n4009 , n4010 , n4011 , n4012 , n4013 , n4014 , n4015 , n4016 , n4017 , n4018 , n4019 , n4020 , n4021 , n4022 , n4023 , n4024 , n4025 , n4026 , n4027 , n4028 , n4029 , n4030 , n4031 , n4032 , n4033 , n4034 , n4035 , n4036 , n4037 , n4038 , n4039 , n4040 , n4041 , n4042 , n4043 , n4044 , n4045 , n4046 , n4047 , n4048 , n4049 , n4050 , n4051 , n4052 , n4053 , n4054 , n4055 , n4056 , n4057 , n4058 , n4059 , n4060 , n4061 , n4062 , n4063 , n4064 , n4065 , n4066 , n4067 , n4068 , n4069 , n4070 , n4071 , n4072 , n4073 , n4074 , n4075 , n4076 , n4077 , n4078 , n4079 , n4080 , n4081 , n4082 , n4083 , n4084 , n4085 , n4086 , n4087 , n4088 , n4089 , n4090 , n4091 , n4092 , n4093 , n4094 , n4095 , n4096 , n4097 , n4098 , n4099 , n4100 , n4101 , n4102 , n4103 , n4104 , n4105 , n4106 , n4107 , n4108 , n4109 , n4110 , n4111 , n4112 , n4113 , n4114 , n4115 , n4116 , n4117 , n4118 , n4119 , n4120 , n4121 , n4122 , n4123 , n4124 , n4125 , n4126 , n4127 , n4128 , n4129 , n4130 , n4131 , n4132 , n4133 , n4134 , n4135 , n4136 , n4137 , n4138 , n4139 , n4140 , n4141 , n4142 , n4143 , n4144 , n4145 , n4146 , n4147 , n4148 , n4149 , n4150 , n4151 , n4152 , n4153 , n4154 , n4155 , n4156 , n4157 , n4158 , n4159 , n4160 , n4161 , n4162 , n4163 , n4164 , n4165 , n4166 , n4167 , n4168 , n4169 , n4170 , n4171 , n4172 , n4173 , n4174 , n4175 , n4176 , n4177 , n4178 , n4179 , n4180 , n4181 , n4182 , n4183 , n4184 , n4185 , n4186 , n4187 , n4188 , n4189 , n4190 , n4191 , n4192 , n4193 , n4194 , n4195 , n4196 , n4197 , n4198 , n4199 , n4200 , n4201 , n4202 , n4203 , n4204 , n4205 , n4206 , n4207 , n4208 , n4209 , n4210 , n4211 , n4212 , n4213 , n4214 , n4215 , n4216 , n4217 , n4218 , n4219 , n4220 , n4221 , n4222 , n4223 , n4224 , n4225 , n4226 , n4227 , n4228 , n4229 , n4230 , n4231 , n4232 , n4233 , n4234 , n4235 , n4236 , n4237 , n4238 , n4239 , n4240 , n4241 , n4242 , n4243 , n4244 , n4245 , n4246 , n4247 , n4248 , n4249 , n4250 , n4251 , n4252 , n4253 , n4254 , n4255 , n4256 , n4257 , n4258 , n4259 , n4260 , n4261 , n4262 , n4263 , n4264 , n4265 , n4266 , n4267 , n4268 , n4269 , n4270 , n4271 , n4272 , n4273 , n4274 , n4275 , n4276 , n4277 , n4278 , n4279 , n4280 , n4281 , n4282 , n4283 , n4284 , n4285 , n4286 , n4287 , n4288 , n4289 , n4290 , n4291 , n4292 , n4293 , n4294 , n4295 , n4296 , n4297 , n4298 , n4299 , n4300 , n4301 , n4302 , n4303 , n4304 , n4305 , n4306 , n4307 , n4308 , n4309 , n4310 , n4311 , n4312 , n4313 , n4314 , n4315 , n4316 , n4317 , n4318 , n4319 , n4320 , n4321 , n4322 , n4323 , n4324 , n4325 , n4326 , n4327 , n4328 , n4329 , n4330 , n4331 , n4332 , n4333 , n4334 , n4335 , n4336 , n4337 , n4338 , n4339 , n4340 , n4341 , n4342 , n4343 , n4344 , n4345 , n4346 , n4347 , n4348 , n4349 , n4350 , n4351 , n4352 , n4353 , n4354 , n4355 , n4356 , n4357 , n4358 , n4359 , n4360 , n4361 , n4362 , n4363 , n4364 , n4365 , n4366 , n4367 , n4368 , n4369 , n4370 , n4371 , n4372 , n4373 , n4374 , n4375 , n4376 , n4377 , n4378 , n4379 , n4380 , n4381 , n4382 , n4383 , n4384 , n4385 , n4386 , n4387 , n4388 , n4389 , n4390 , n4391 , n4392 , n4393 , n4394 , n4395 , n4396 , n4397 , n4398 , n4399 , n4400 , n4401 , n4402 , n4403 , n4404 , n4405 , n4406 , n4407 , n4408 , n4409 , n4410 , n4411 , n4412 , n4413 , n4414 , n4415 , n4416 , n4417 , n4418 , n4419 , n4420 , n4421 , n4422 , n4423 , n4424 , n4425 , n4426 , n4427 , n4428 , n4429 , n4430 , n4431 , n4432 , n4433 , n4434 , n4435 , n4436 , n4437 , n4438 , n4439 , n4440 , n4441 , n4442 , n4443 , n4444 , n4445 , n4446 , n4447 , n4448 , n4449 , n4450 , n4451 , n4452 , n4453 , n4454 , n4455 , n4456 , n4457 , n4458 , n4459 , n4460 , n4461 , n4462 , n4463 , n4464 , n4465 , n4466 , n4467 , n4468 , n4469 , n4470 , n4471 , n4472 , n4473 , n4474 , n4475 , n4476 , n4477 , n4478 , n4479 , n4480 , n4481 , n4482 , n4483 , n4484 , n4485 , n4486 , n4487 , n4488 , n4489 , n4490 , n4491 , n4492 , n4493 , n4494 , n4495 , n4496 , n4497 , n4498 , n4499 , n4500 , n4501 , n4502 , n4503 , n4504 , n4505 , n4506 , n4507 , n4508 , n4509 , n4510 , n4511 , n4512 , n4513 , n4514 , n4515 , n4516 , n4517 , n4518 , n4519 , n4520 , n4521 , n4522 , n4523 , n4524 , n4525 , n4526 , n4527 , n4528 , n4529 , n4530 , n4531 , n4532 , n4533 , n4534 , n4535 , n4536 , n4537 , n4538 , n4539 , n4540 , n4541 , n4542 , n4543 , n4544 , n4545 , n4546 , n4547 , n4548 , n4549 , n4550 , n4551 , n4552 , n4553 , n4554 , n4555 , n4556 , n4557 , n4558 , n4559 , n4560 , n4561 , n4562 , n4563 , n4564 , n4565 , n4566 , n4567 , n4568 , n4569 , n4570 , n4571 , n4572 , n4573 , n4574 , n4575 , n4576 , n4577 , n4578 , n4579 , n4580 , n4581 , n4582 , n4583 , n4584 , n4585 , n4586 , n4587 , n4588 , n4589 , n4590 , n4591 , n4592 , n4593 , n4594 , n4595 , n4596 , n4597 , n4598 , n4599 , n4600 , n4601 , n4602 , n4603 , n4604 , n4605 , n4606 , n4607 , n4608 , n4609 , n4610 , n4611 , n4612 , n4613 , n4614 , n4615 , n4616 , n4617 , n4618 , n4619 , n4620 , n4621 , n4622 , n4623 , n4624 , n4625 , n4626 , n4627 , n4628 , n4629 , n4630 , n4631 , n4632 , n4633 , n4634 , n4635 , n4636 , n4637 , n4638 , n4639 , n4640 , n4641 , n4642 , n4643 , n4644 , n4645 , n4646 , n4647 , n4648 , n4649 , n4650 , n4651 , n4652 , n4653 , n4654 , n4655 , n4656 , n4657 , n4658 , n4659 , n4660 , n4661 , n4662 , n4663 , n4664 , n4665 , n4666 , n4667 , n4668 , n4669 , n4670 , n4671 , n4672 , n4673 , n4674 , n4675 , n4676 , n4677 , n4678 , n4679 , n4680 , n4681 , n4682 , n4683 , n4684 , n4685 , n4686 , n4687 , n4688 , n4689 , n4690 , n4691 , n4692 , n4693 , n4694 , n4695 , n4696 , n4697 , n4698 , n4699 , n4700 , n4701 , n4702 , n4703 , n4704 , n4705 , n4706 , n4707 , n4708 , n4709 , n4710 , n4711 , n4712 , n4713 , n4714 , n4715 , n4716 , n4717 , n4718 , n4719 , n4720 , n4721 , n4722 , n4723 , n4724 , n4725 , n4726 , n4727 , n4728 , n4729 , n4730 , n4731 , n4732 , n4733 , n4734 , n4735 , n4736 , n4737 , n4738 , n4739 , n4740 , n4741 , n4742 , n4743 , n4744 , n4745 , n4746 , n4747 , n4748 , n4749 , n4750 , n4751 , n4752 , n4753 , n4754 , n4755 , n4756 , n4757 , n4758 , n4759 , n4760 , n4761 , n4762 , n4763 , n4764 , n4765 , n4766 , n4767 , n4768 , n4769 , n4770 , n4771 , n4772 , n4773 , n4774 , n4775 , n4776 , n4777 , n4778 , n4779 , n4780 , n4781 , n4782 , n4783 , n4784 , n4785 , n4786 , n4787 , n4788 , n4789 , n4790 , n4791 , n4792 , n4793 , n4794 , n4795 , n4796 , n4797 , n4798 , n4799 , n4800 , n4801 , n4802 , n4803 , n4804 , n4805 , n4806 , n4807 , n4808 , n4809 , n4810 , n4811 , n4812 , n4813 , n4814 , n4815 , n4816 , n4817 , n4818 , n4819 , n4820 , n4821 , n4822 , n4823 , n4824 , n4825 , n4826 , n4827 , n4828 , n4829 , n4830 , n4831 , n4832 , n4833 , n4834 , n4835 , n4836 , n4837 , n4838 , n4839 , n4840 , n4841 , n4842 , n4843 , n4844 , n4845 , n4846 , n4847 , n4848 , n4849 , n4850 , n4851 , n4852 , n4853 , n4854 , n4855 , n4856 , n4857 , n4858 , n4859 , n4860 , n4861 , n4862 , n4863 , n4864 , n4865 , n4866 , n4867 , n4868 , n4869 , n4870 , n4871 , n4872 , n4873 , n4874 , n4875 , n4876 , n4877 , n4878 , n4879 , n4880 , n4881 , n4882 , n4883 , n4884 , n4885 , n4886 , n4887 , n4888 , n4889 , n4890 , n4891 , n4892 , n4893 , n4894 , n4895 , n4896 , n4897 , n4898 , n4899 , n4900 , n4901 , n4902 , n4903 , n4904 , n4905 , n4906 , n4907 , n4908 , n4909 , n4910 , n4911 , n4912 , n4913 , n4914 , n4915 , n4916 , n4917 , n4918 , n4919 , n4920 , n4921 , n4922 , n4923 , n4924 , n4925 , n4926 , n4927 , n4928 , n4929 , n4930 , n4931 , n4932 , n4933 , n4934 , n4935 , n4936 , n4937 , n4938 , n4939 , n4940 , n4941 , n4942 , n4943 , n4944 , n4945 , n4946 , n4947 , n4948 , n4949 , n4950 , n4951 , n4952 , n4953 , n4954 , n4955 , n4956 , n4957 , n4958 , n4959 , n4960 , n4961 , n4962 , n4963 , n4964 , n4965 , n4966 , n4967 , n4968 , n4969 , n4970 , n4971 , n4972 , n4973 , n4974 , n4975 , n4976 , n4977 , n4978 , n4979 , n4980 , n4981 , n4982 , n4983 , n4984 , n4985 , n4986 , n4987 , n4988 , n4989 , n4990 , n4991 , n4992 , n4993 , n4994 , n4995 , n4996 , n4997 , n4998 , n4999 , n5000 , n5001 , n5002 , n5003 , n5004 , n5005 , n5006 , n5007 , n5008 , n5009 , n5010 , n5011 , n5012 , n5013 , n5014 , n5015 , n5016 , n5017 , n5018 , n5019 , n5020 , n5021 , n5022 , n5023 , n5024 , n5025 , n5026 , n5027 , n5028 , n5029 , n5030 , n5031 , n5032 , n5033 , n5034 , n5035 , n5036 , n5037 , n5038 , n5039 , n5040 , n5041 , n5042 , n5043 , n5044 , n5045 , n5046 , n5047 , n5048 , n5049 , n5050 , n5051 , n5052 , n5053 , n5054 , n5055 , n5056 , n5057 , n5058 , n5059 , n5060 , n5061 , n5062 , n5063 , n5064 , n5065 , n5066 , n5067 , n5068 , n5069 , n5070 , n5071 , n5072 , n5073 , n5074 , n5075 , n5076 , n5077 , n5078 , n5079 , n5080 , n5081 , n5082 , n5083 , n5084 , n5085 , n5086 , n5087 , n5088 , n5089 , n5090 , n5091 , n5092 , n5093 , n5094 , n5095 , n5096 , n5097 , n5098 , n5099 , n5100 , n5101 , n5102 , n5103 , n5104 , n5105 , n5106 , n5107 , n5108 , n5109 , n5110 , n5111 , n5112 , n5113 , n5114 , n5115 , n5116 , n5117 , n5118 , n5119 , n5120 , n5121 , n5122 , n5123 , n5124 , n5125 , n5126 , n5127 , n5128 , n5129 , n5130 , n5131 , n5132 , n5133 , n5134 , n5135 , n5136 , n5137 , n5138 , n5139 , n5140 , n5141 , n5142 , n5143 , n5144 , n5145 , n5146 , n5147 , n5148 , n5149 , n5150 , n5151 , n5152 , n5153 , n5154 , n5155 , n5156 , n5157 , n5158 , n5159 , n5160 , n5161 , n5162 , n5163 , n5164 , n5165 , n5166 , n5167 , n5168 , n5169 , n5170 , n5171 , n5172 , n5173 , n5174 , n5175 , n5176 , n5177 , n5178 , n5179 , n5180 , n5181 , n5182 , n5183 , n5184 , n5185 , n5186 , n5187 , n5188 , n5189 , n5190 , n5191 , n5192 , n5193 , n5194 , n5195 , n5196 , n5197 , n5198 , n5199 , n5200 , n5201 , n5202 , n5203 , n5204 , n5205 , n5206 , n5207 , n5208 , n5209 , n5210 , n5211 , n5212 , n5213 , n5214 , n5215 , n5216 , n5217 , n5218 , n5219 , n5220 , n5221 , n5222 , n5223 , n5224 , n5225 , n5226 , n5227 , n5228 , n5229 , n5230 , n5231 , n5232 , n5233 , n5234 , n5235 , n5236 , n5237 , n5238 , n5239 , n5240 , n5241 , n5242 , n5243 , n5244 , n5245 , n5246 , n5247 , n5248 , n5249 , n5250 , n5251 , n5252 , n5253 , n5254 , n5255 , n5256 , n5257 , n5258 , n5259 , n5260 , n5261 , n5262 , n5263 , n5264 , n5265 , n5266 , n5267 , n5268 , n5269 , n5270 , n5271 , n5272 , n5273 , n5274 , n5275 , n5276 , n5277 , n5278 , n5279 , n5280 , n5281 , n5282 , n5283 , n5284 , n5285 , n5286 , n5287 , n5288 , n5289 , n5290 , n5291 , n5292 , n5293 , n5294 , n5295 , n5296 , n5297 , n5298 , n5299 , n5300 , n5301 , n5302 , n5303 , n5304 , n5305 , n5306 , n5307 , n5308 , n5309 , n5310 , n5311 , n5312 , n5313 , n5314 , n5315 , n5316 , n5317 , n5318 , n5319 , n5320 , n5321 , n5322 , n5323 , n5324 , n5325 , n5326 , n5327 , n5328 , n5329 , n5330 , n5331 , n5332 , n5333 , n5334 , n5335 , n5336 , n5337 , n5338 , n5339 , n5340 , n5341 , n5342 , n5343 , n5344 , n5345 , n5346 , n5347 , n5348 , n5349 , n5350 , n5351 , n5352 , n5353 , n5354 , n5355 , n5356 , n5357 , n5358 , n5359 , n5360 , n5361 , n5362 , n5363 , n5364 , n5365 , n5366 , n5367 , n5368 , n5369 , n5370 , n5371 , n5372 , n5373 , n5374 , n5375 , n5376 , n5377 , n5378 , n5379 , n5380 , n5381 , n5382 , n5383 , n5384 , n5385 , n5386 , n5387 , n5388 , n5389 , n5390 , n5391 , n5392 , n5393 , n5394 , n5395 , n5396 , n5397 , n5398 , n5399 , n5400 , n5401 , n5402 , n5403 , n5404 , n5405 , n5406 , n5407 , n5408 , n5409 , n5410 , n5411 , n5412 , n5413 , n5414 , n5415 , n5416 , n5417 , n5418 , n5419 , n5420 , n5421 , n5422 , n5423 , n5424 , n5425 , n5426 , n5427 , n5428 , n5429 , n5430 , n5431 , n5432 , n5433 , n5434 , n5435 , n5436 , n5437 , n5438 , n5439 , n5440 , n5441 , n5442 , n5443 , n5444 , n5445 , n5446 , n5447 , n5448 , n5449 , n5450 , n5451 , n5452 , n5453 , n5454 , n5455 , n5456 , n5457 , n5458 , n5459 , n5460 , n5461 , n5462 , n5463 , n5464 , n5465 , n5466 , n5467 , n5468 , n5469 , n5470 , n5471 , n5472 , n5473 , n5474 , n5475 , n5476 , n5477 , n5478 , n5479 , n5480 , n5481 , n5482 , n5483 , n5484 , n5485 , n5486 , n5487 , n5488 , n5489 , n5490 , n5491 , n5492 , n5493 , n5494 , n5495 , n5496 , n5497 , n5498 , n5499 , n5500 , n5501 , n5502 , n5503 , n5504 , n5505 , n5506 , n5507 , n5508 , n5509 , n5510 , n5511 , n5512 , n5513 , n5514 , n5515 , n5516 , n5517 , n5518 , n5519 , n5520 , n5521 , n5522 , n5523 , n5524 , n5525 , n5526 , n5527 , n5528 , n5529 , n5530 , n5531 , n5532 , n5533 , n5534 , n5535 , n5536 , n5537 , n5538 , n5539 , n5540 , n5541 , n5542 , n5543 , n5544 , n5545 , n5546 , n5547 , n5548 , n5549 , n5550 , n5551 , n5552 , n5553 , n5554 , n5555 , n5556 , n5557 , n5558 , n5559 , n5560 , n5561 , n5562 , n5563 , n5564 , n5565 , n5566 , n5567 , n5568 , n5569 , n5570 , n5571 , n5572 , n5573 , n5574 , n5575 , n5576 , n5577 , n5578 , n5579 , n5580 , n5581 , n5582 , n5583 , n5584 , n5585 , n5586 , n5587 , n5588 , n5589 , n5590 , n5591 , n5592 , n5593 , n5594 , n5595 , n5596 , n5597 , n5598 , n5599 , n5600 , n5601 , n5602 , n5603 , n5604 , n5605 , n5606 , n5607 , n5608 , n5609 , n5610 , n5611 , n5612 , n5613 , n5614 , n5615 , n5616 , n5617 , n5618 , n5619 , n5620 , n5621 , n5622 , n5623 , n5624 , n5625 , n5626 , n5627 , n5628 , n5629 , n5630 , n5631 , n5632 , n5633 , n5634 , n5635 , n5636 , n5637 , n5638 , n5639 , n5640 , n5641 , n5642 , n5643 , n5644 , n5645 , n5646 , n5647 , n5648 , n5649 , n5650 , n5651 , n5652 , n5653 , n5654 , n5655 , n5656 , n5657 , n5658 , n5659 , n5660 , n5661 , n5662 , n5663 , n5664 , n5665 , n5666 , n5667 , n5668 , n5669 , n5670 , n5671 , n5672 , n5673 , n5674 , n5675 , n5676 , n5677 , n5678 , n5679 , n5680 , n5681 , n5682 , n5683 , n5684 , n5685 , n5686 , n5687 , n5688 , n5689 , n5690 , n5691 , n5692 , n5693 , n5694 , n5695 , n5696 , n5697 , n5698 , n5699 , n5700 , n5701 , n5702 , n5703 , n5704 , n5705 , n5706 , n5707 , n5708 , n5709 , n5710 , n5711 , n5712 , n5713 , n5714 , n5715 , n5716 , n5717 , n5718 , n5719 , n5720 , n5721 , n5722 , n5723 , n5724 , n5725 , n5726 , n5727 , n5728 , n5729 , n5730 , n5731 , n5732 , n5733 , n5734 , n5735 , n5736 , n5737 , n5738 , n5739 , n5740 , n5741 , n5742 , n5743 , n5744 , n5745 , n5746 , n5747 , n5748 , n5749 , n5750 , n5751 , n5752 , n5753 , n5754 , n5755 , n5756 , n5757 , n5758 , n5759 , n5760 , n5761 , n5762 , n5763 , n5764 , n5765 , n5766 , n5767 , n5768 , n5769 , n5770 , n5771 , n5772 , n5773 , n5774 , n5775 , n5776 , n5777 , n5778 , n5779 , n5780 , n5781 , n5782 , n5783 , n5784 , n5785 , n5786 , n5787 , n5788 , n5789 , n5790 , n5791 , n5792 , n5793 , n5794 , n5795 , n5796 , n5797 , n5798 , n5799 , n5800 , n5801 , n5802 , n5803 , n5804 , n5805 , n5806 , n5807 , n5808 , n5809 , n5810 , n5811 , n5812 , n5813 , n5814 , n5815 , n5816 , n5817 , n5818 , n5819 , n5820 , n5821 , n5822 , n5823 , n5824 , n5825 , n5826 , n5827 , n5828 , n5829 , n5830 , n5831 , n5832 , n5833 , n5834 , n5835 , n5836 , n5837 , n5838 , n5839 , n5840 , n5841 , n5842 , n5843 , n5844 , n5845 , n5846 , n5847 , n5848 , n5849 , n5850 , n5851 , n5852 , n5853 , n5854 , n5855 , n5856 , n5857 , n5858 , n5859 , n5860 , n5861 , n5862 , n5863 , n5864 , n5865 , n5866 , n5867 , n5868 , n5869 , n5870 , n5871 , n5872 , n5873 , n5874 , n5875 , n5876 , n5877 , n5878 , n5879 , n5880 , n5881 , n5882 , n5883 , n5884 , n5885 , n5886 , n5887 , n5888 , n5889 , n5890 , n5891 , n5892 , n5893 , n5894 , n5895 , n5896 , n5897 , n5898 , n5899 , n5900 , n5901 , n5902 , n5903 , n5904 , n5905 , n5906 , n5907 , n5908 , n5909 , n5910 , n5911 , n5912 , n5913 , n5914 , n5915 , n5916 , n5917 , n5918 , n5919 , n5920 , n5921 , n5922 , n5923 , n5924 , n5925 , n5926 , n5927 , n5928 , n5929 , n5930 , n5931 , n5932 , n5933 , n5934 , n5935 , n5936 , n5937 , n5938 , n5939 , n5940 , n5941 , n5942 , n5943 , n5944 , n5945 , n5946 , n5947 , n5948 , n5949 , n5950 , n5951 , n5952 , n5953 , n5954 , n5955 , n5956 , n5957 , n5958 , n5959 , n5960 , n5961 , n5962 , n5963 , n5964 , n5965 , n5966 , n5967 , n5968 , n5969 , n5970 , n5971 , n5972 , n5973 , n5974 , n5975 , n5976 , n5977 , n5978 , n5979 , n5980 , n5981 , n5982 , n5983 , n5984 , n5985 , n5986 , n5987 , n5988 , n5989 , n5990 , n5991 , n5992 , n5993 , n5994 , n5995 , n5996 , n5997 , n5998 , n5999 , n6000 , n6001 , n6002 , n6003 , n6004 , n6005 , n6006 , n6007 , n6008 , n6009 , n6010 , n6011 , n6012 , n6013 , n6014 , n6015 , n6016 , n6017 , n6018 , n6019 , n6020 , n6021 , n6022 , n6023 , n6024 , n6025 , n6026 , n6027 , n6028 , n6029 , n6030 , n6031 , n6032 , n6033 , n6034 , n6035 , n6036 , n6037 , n6038 , n6039 , n6040 , n6041 , n6042 , n6043 , n6044 , n6045 , n6046 , n6047 , n6048 , n6049 , n6050 , n6051 , n6052 , n6053 , n6054 , n6055 , n6056 , n6057 , n6058 , n6059 , n6060 , n6061 , n6062 , n6063 , n6064 , n6065 , n6066 , n6067 , n6068 , n6069 , n6070 , n6071 , n6072 , n6073 , n6074 , n6075 , n6076 , n6077 , n6078 , n6079 , n6080 , n6081 , n6082 , n6083 , n6084 , n6085 , n6086 , n6087 , n6088 , n6089 , n6090 , n6091 , n6092 , n6093 , n6094 , n6095 , n6096 , n6097 , n6098 , n6099 , n6100 , n6101 , n6102 , n6103 , n6104 , n6105 , n6106 , n6107 , n6108 , n6109 , n6110 , n6111 , n6112 , n6113 , n6114 , n6115 , n6116 , n6117 , n6118 , n6119 , n6120 , n6121 , n6122 , n6123 , n6124 , n6125 , n6126 , n6127 , n6128 , n6129 , n6130 , n6131 , n6132 , n6133 , n6134 , n6135 , n6136 , n6137 , n6138 , n6139 , n6140 , n6141 , n6142 , n6143 , n6144 , n6145 , n6146 , n6147 , n6148 , n6149 , n6150 , n6151 , n6152 , n6153 , n6154 , n6155 , n6156 , n6157 , n6158 , n6159 , n6160 , n6161 , n6162 , n6163 , n6164 , n6165 , n6166 , n6167 , n6168 , n6169 , n6170 , n6171 , n6172 , n6173 , n6174 , n6175 , n6176 , n6177 , n6178 , n6179 , n6180 , n6181 , n6182 , n6183 , n6184 , n6185 , n6186 , n6187 , n6188 , n6189 , n6190 , n6191 , n6192 , n6193 , n6194 , n6195 , n6196 , n6197 , n6198 , n6199 , n6200 , n6201 , n6202 , n6203 , n6204 , n6205 , n6206 , n6207 , n6208 , n6209 , n6210 , n6211 , n6212 , n6213 , n6214 , n6215 , n6216 , n6217 , n6218 , n6219 , n6220 , n6221 , n6222 , n6223 , n6224 , n6225 , n6226 , n6227 , n6228 , n6229 , n6230 , n6231 , n6232 , n6233 , n6234 , n6235 , n6236 , n6237 , n6238 , n6239 , n6240 , n6241 , n6242 , n6243 , n6244 , n6245 , n6246 , n6247 , n6248 , n6249 , n6250 , n6251 , n6252 , n6253 , n6254 , n6255 , n6256 , n6257 , n6258 , n6259 , n6260 , n6261 , n6262 , n6263 , n6264 , n6265 , n6266 , n6267 , n6268 , n6269 , n6270 , n6271 , n6272 , n6273 , n6274 , n6275 , n6276 , n6277 , n6278 , n6279 , n6280 , n6281 , n6282 , n6283 , n6284 , n6285 , n6286 , n6287 , n6288 , n6289 , n6290 , n6291 , n6292 , n6293 , n6294 , n6295 , n6296 , n6297 , n6298 , n6299 , n6300 , n6301 , n6302 , n6303 , n6304 , n6305 , n6306 , n6307 , n6308 , n6309 , n6310 , n6311 , n6312 , n6313 , n6314 , n6315 , n6316 , n6317 , n6318 , n6319 , n6320 , n6321 , n6322 , n6323 , n6324 , n6325 , n6326 , n6327 , n6328 , n6329 , n6330 , n6331 , n6332 , n6333 , n6334 , n6335 , n6336 , n6337 , n6338 , n6339 , n6340 , n6341 , n6342 , n6343 , n6344 , n6345 , n6346 , n6347 , n6348 , n6349 , n6350 , n6351 , n6352 , n6353 , n6354 , n6355 , n6356 , n6357 , n6358 , n6359 , n6360 , n6361 , n6362 , n6363 , n6364 , n6365 , n6366 , n6367 , n6368 , n6369 , n6370 , n6371 , n6372 , n6373 , n6374 , n6375 , n6376 , n6377 , n6378 , n6379 , n6380 , n6381 , n6382 , n6383 , n6384 , n6385 , n6386 , n6387 , n6388 , n6389 , n6390 , n6391 , n6392 , n6393 , n6394 , n6395 , n6396 , n6397 , n6398 , n6399 , n6400 , n6401 , n6402 , n6403 , n6404 , n6405 , n6406 , n6407 , n6408 , n6409 , n6410 , n6411 , n6412 , n6413 , n6414 , n6415 , n6416 , n6417 , n6418 , n6419 , n6420 , n6421 , n6422 , n6423 , n6424 , n6425 , n6426 , n6427 , n6428 , n6429 , n6430 , n6431 , n6432 , n6433 , n6434 , n6435 , n6436 , n6437 , n6438 , n6439 , n6440 , n6441 , n6442 , n6443 , n6444 , n6445 , n6446 , n6447 , n6448 , n6449 , n6450 , n6451 , n6452 , n6453 , n6454 , n6455 , n6456 , n6457 , n6458 , n6459 , n6460 , n6461 , n6462 , n6463 , n6464 , n6465 , n6466 , n6467 , n6468 , n6469 , n6470 , n6471 , n6472 , n6473 , n6474 , n6475 , n6476 , n6477 , n6478 , n6479 , n6480 , n6481 , n6482 , n6483 , n6484 , n6485 , n6486 , n6487 , n6488 , n6489 , n6490 , n6491 , n6492 , n6493 , n6494 , n6495 , n6496 , n6497 , n6498 , n6499 , n6500 , n6501 , n6502 , n6503 , n6504 , n6505 , n6506 , n6507 , n6508 , n6509 , n6510 , n6511 , n6512 , n6513 , n6514 , n6515 , n6516 , n6517 , n6518 , n6519 , n6520 , n6521 , n6522 , n6523 , n6524 , n6525 , n6526 , n6527 , n6528 , n6529 , n6530 , n6531 , n6532 , n6533 , n6534 , n6535 , n6536 , n6537 , n6538 , n6539 , n6540 , n6541 , n6542 , n6543 , n6544 , n6545 , n6546 , n6547 , n6548 , n6549 , n6550 , n6551 , n6552 , n6553 , n6554 , n6555 , n6556 , n6557 , n6558 , n6559 , n6560 , n6561 , n6562 , n6563 , n6564 , n6565 , n6566 , n6567 , n6568 , n6569 , n6570 , n6571 , n6572 , n6573 , n6574 , n6575 , n6576 , n6577 , n6578 , n6579 , n6580 , n6581 , n6582 , n6583 , n6584 , n6585 , n6586 , n6587 , n6588 , n6589 , n6590 , n6591 , n6592 , n6593 , n6594 , n6595 , n6596 , n6597 , n6598 , n6599 , n6600 , n6601 , n6602 , n6603 , n6604 , n6605 , n6606 , n6607 , n6608 , n6609 , n6610 , n6611 , n6612 , n6613 , n6614 , n6615 , n6616 , n6617 , n6618 , n6619 , n6620 , n6621 , n6622 , n6623 , n6624 , n6625 , n6626 , n6627 , n6628 , n6629 , n6630 , n6631 , n6632 , n6633 , n6634 , n6635 , n6636 , n6637 , n6638 , n6639 , n6640 , n6641 , n6642 , n6643 , n6644 , n6645 , n6646 , n6647 , n6648 , n6649 , n6650 , n6651 , n6652 , n6653 , n6654 , n6655 , n6656 , n6657 , n6658 , n6659 , n6660 , n6661 , n6662 , n6663 , n6664 , n6665 , n6666 , n6667 , n6668 , n6669 , n6670 , n6671 , n6672 , n6673 , n6674 , n6675 , n6676 , n6677 , n6678 , n6679 , n6680 , n6681 , n6682 , n6683 , n6684 , n6685 , n6686 , n6687 , n6688 , n6689 , n6690 , n6691 , n6692 , n6693 , n6694 , n6695 , n6696 , n6697 , n6698 , n6699 , n6700 , n6701 , n6702 , n6703 , n6704 , n6705 , n6706 , n6707 , n6708 , n6709 , n6710 , n6711 , n6712 , n6713 , n6714 , n6715 , n6716 , n6717 , n6718 , n6719 , n6720 , n6721 , n6722 , n6723 , n6724 , n6725 , n6726 , n6727 , n6728 , n6729 , n6730 , n6731 , n6732 , n6733 , n6734 , n6735 , n6736 , n6737 , n6738 , n6739 , n6740 , n6741 , n6742 , n6743 , n6744 , n6745 , n6746 , n6747 , n6748 , n6749 , n6750 , n6751 , n6752 , n6753 , n6754 , n6755 , n6756 , n6757 , n6758 , n6759 , n6760 , n6761 , n6762 , n6763 , n6764 , n6765 , n6766 , n6767 , n6768 , n6769 , n6770 , n6771 , n6772 , n6773 , n6774 , n6775 , n6776 , n6777 , n6778 , n6779 , n6780 , n6781 , n6782 , n6783 , n6784 , n6785 , n6786 , n6787 , n6788 , n6789 , n6790 , n6791 , n6792 , n6793 , n6794 , n6795 , n6796 , n6797 , n6798 , n6799 , n6800 , n6801 , n6802 , n6803 , n6804 , n6805 , n6806 , n6807 , n6808 , n6809 , n6810 , n6811 , n6812 , n6813 , n6814 , n6815 , n6816 , n6817 , n6818 , n6819 , n6820 , n6821 , n6822 , n6823 , n6824 , n6825 , n6826 , n6827 , n6828 , n6829 , n6830 , n6831 , n6832 , n6833 , n6834 , n6835 , n6836 , n6837 , n6838 , n6839 , n6840 , n6841 , n6842 , n6843 , n6844 , n6845 , n6846 , n6847 , n6848 , n6849 , n6850 , n6851 , n6852 , n6853 , n6854 , n6855 , n6856 , n6857 , n6858 , n6859 , n6860 , n6861 , n6862 , n6863 , n6864 , n6865 , n6866 , n6867 , n6868 , n6869 , n6870 , n6871 , n6872 , n6873 , n6874 , n6875 , n6876 , n6877 , n6878 , n6879 , n6880 , n6881 , n6882 , n6883 , n6884 , n6885 , n6886 , n6887 , n6888 , n6889 , n6890 , n6891 , n6892 , n6893 , n6894 , n6895 , n6896 , n6897 , n6898 , n6899 , n6900 , n6901 , n6902 , n6903 , n6904 , n6905 , n6906 , n6907 , n6908 , n6909 , n6910 , n6911 , n6912 , n6913 , n6914 , n6915 , n6916 , n6917 , n6918 , n6919 , n6920 , n6921 , n6922 , n6923 , n6924 , n6925 , n6926 , n6927 , n6928 , n6929 , n6930 , n6931 , n6932 , n6933 , n6934 , n6935 , n6936 , n6937 , n6938 , n6939 , n6940 , n6941 , n6942 , n6943 , n6944 , n6945 , n6946 , n6947 , n6948 , n6949 , n6950 , n6951 , n6952 , n6953 , n6954 , n6955 , n6956 , n6957 , n6958 , n6959 , n6960 , n6961 , n6962 , n6963 , n6964 , n6965 , n6966 , n6967 , n6968 , n6969 , n6970 , n6971 , n6972 , n6973 , n6974 , n6975 , n6976 , n6977 , n6978 , n6979 , n6980 , n6981 , n6982 , n6983 , n6984 , n6985 , n6986 , n6987 , n6988 , n6989 , n6990 , n6991 , n6992 , n6993 , n6994 , n6995 , n6996 , n6997 , n6998 , n6999 , n7000 , n7001 , n7002 , n7003 , n7004 , n7005 , n7006 , n7007 , n7008 , n7009 , n7010 , n7011 , n7012 , n7013 , n7014 , n7015 , n7016 , n7017 , n7018 , n7019 , n7020 , n7021 , n7022 , n7023 , n7024 , n7025 , n7026 , n7027 , n7028 , n7029 , n7030 , n7031 , n7032 , n7033 , n7034 , n7035 , n7036 , n7037 , n7038 , n7039 , n7040 , n7041 , n7042 , n7043 , n7044 , n7045 , n7046 , n7047 , n7048 , n7049 , n7050 , n7051 , n7052 , n7053 , n7054 , n7055 , n7056 , n7057 , n7058 , n7059 , n7060 , n7061 , n7062 , n7063 , n7064 , n7065 , n7066 , n7067 , n7068 , n7069 , n7070 , n7071 , n7072 , n7073 , n7074 , n7075 , n7076 , n7077 , n7078 , n7079 , n7080 , n7081 , n7082 , n7083 , n7084 , n7085 , n7086 , n7087 , n7088 , n7089 , n7090 , n7091 , n7092 , n7093 , n7094 , n7095 , n7096 , n7097 , n7098 , n7099 , n7100 , n7101 , n7102 , n7103 , n7104 , n7105 , n7106 , n7107 , n7108 , n7109 , n7110 , n7111 , n7112 , n7113 , n7114 , n7115 , n7116 , n7117 , n7118 , n7119 , n7120 , n7121 , n7122 , n7123 , n7124 , n7125 , n7126 , n7127 , n7128 , n7129 , n7130 , n7131 , n7132 , n7133 , n7134 , n7135 , n7136 , n7137 , n7138 , n7139 , n7140 , n7141 , n7142 , n7143 , n7144 , n7145 , n7146 , n7147 , n7148 , n7149 , n7150 , n7151 , n7152 , n7153 , n7154 , n7155 , n7156 , n7157 , n7158 , n7159 , n7160 , n7161 , n7162 , n7163 , n7164 , n7165 , n7166 , n7167 , n7168 , n7169 , n7170 , n7171 , n7172 , n7173 , n7174 , n7175 , n7176 , n7177 , n7178 , n7179 , n7180 , n7181 , n7182 , n7183 , n7184 , n7185 , n7186 , n7187 , n7188 , n7189 , n7190 , n7191 , n7192 , n7193 , n7194 , n7195 , n7196 , n7197 , n7198 , n7199 , n7200 , n7201 , n7202 , n7203 , n7204 , n7205 , n7206 , n7207 , n7208 , n7209 , n7210 , n7211 , n7212 , n7213 , n7214 , n7215 , n7216 , n7217 , n7218 , n7219 , n7220 , n7221 , n7222 , n7223 , n7224 , n7225 , n7226 , n7227 , n7228 , n7229 , n7230 , n7231 , n7232 , n7233 , n7234 , n7235 , n7236 , n7237 , n7238 , n7239 , n7240 , n7241 , n7242 , n7243 , n7244 , n7245 , n7246 , n7247 , n7248 , n7249 , n7250 , n7251 , n7252 , n7253 , n7254 , n7255 , n7256 , n7257 , n7258 , n7259 , n7260 , n7261 , n7262 , n7263 , n7264 , n7265 , n7266 , n7267 , n7268 , n7269 , n7270 , n7271 , n7272 , n7273 , n7274 , n7275 , n7276 , n7277 , n7278 , n7279 , n7280 , n7281 , n7282 , n7283 , n7284 , n7285 , n7286 , n7287 , n7288 , n7289 , n7290 , n7291 , n7292 , n7293 , n7294 , n7295 , n7296 , n7297 , n7298 , n7299 , n7300 , n7301 , n7302 , n7303 , n7304 , n7305 , n7306 , n7307 , n7308 , n7309 , n7310 , n7311 , n7312 , n7313 , n7314 , n7315 , n7316 , n7317 , n7318 , n7319 , n7320 , n7321 , n7322 , n7323 , n7324 , n7325 , n7326 , n7327 , n7328 , n7329 , n7330 , n7331 , n7332 , n7333 , n7334 , n7335 , n7336 , n7337 , n7338 , n7339 , n7340 , n7341 , n7342 , n7343 , n7344 , n7345 , n7346 , n7347 , n7348 , n7349 , n7350 , n7351 , n7352 , n7353 , n7354 , n7355 , n7356 , n7357 , n7358 , n7359 , n7360 , n7361 , n7362 , n7363 , n7364 , n7365 , n7366 , n7367 , n7368 , n7369 , n7370 , n7371 , n7372 , n7373 , n7374 , n7375 , n7376 , n7377 , n7378 , n7379 , n7380 , n7381 , n7382 , n7383 , n7384 , n7385 , n7386 , n7387 , n7388 , n7389 , n7390 , n7391 , n7392 , n7393 , n7394 , n7395 , n7396 , n7397 , n7398 , n7399 , n7400 , n7401 , n7402 , n7403 , n7404 , n7405 , n7406 , n7407 , n7408 , n7409 , n7410 , n7411 , n7412 , n7413 , n7414 , n7415 , n7416 , n7417 , n7418 , n7419 , n7420 , n7421 , n7422 , n7423 , n7424 , n7425 , n7426 , n7427 , n7428 , n7429 , n7430 , n7431 , n7432 , n7433 , n7434 , n7435 , n7436 , n7437 , n7438 , n7439 , n7440 , n7441 , n7442 , n7443 , n7444 , n7445 , n7446 , n7447 , n7448 , n7449 , n7450 , n7451 , n7452 , n7453 , n7454 , n7455 , n7456 , n7457 , n7458 , n7459 , n7460 , n7461 , n7462 , n7463 , n7464 , n7465 , n7466 , n7467 , n7468 , n7469 , n7470 , n7471 , n7472 , n7473 , n7474 , n7475 , n7476 , n7477 , n7478 , n7479 , n7480 , n7481 , n7482 , n7483 , n7484 , n7485 , n7486 , n7487 , n7488 , n7489 , n7490 , n7491 , n7492 , n7493 , n7494 , n7495 , n7496 , n7497 , n7498 , n7499 , n7500 , n7501 , n7502 , n7503 , n7504 , n7505 , n7506 , n7507 , n7508 , n7509 , n7510 , n7511 , n7512 , n7513 , n7514 , n7515 , n7516 , n7517 , n7518 , n7519 , n7520 , n7521 , n7522 , n7523 , n7524 , n7525 , n7526 , n7527 , n7528 , n7529 , n7530 , n7531 , n7532 , n7533 , n7534 , n7535 , n7536 , n7537 , n7538 , n7539 , n7540 , n7541 , n7542 , n7543 , n7544 , n7545 , n7546 , n7547 , n7548 , n7549 , n7550 , n7551 , n7552 , n7553 , n7554 , n7555 , n7556 , n7557 , n7558 , n7559 , n7560 , n7561 , n7562 , n7563 , n7564 , n7565 , n7566 , n7567 , n7568 , n7569 , n7570 , n7571 , n7572 , n7573 , n7574 , n7575 , n7576 , n7577 , n7578 , n7579 , n7580 , n7581 , n7582 , n7583 , n7584 , n7585 , n7586 , n7587 , n7588 , n7589 , n7590 , n7591 , n7592 , n7593 , n7594 , n7595 , n7596 , n7597 , n7598 , n7599 , n7600 , n7601 , n7602 , n7603 , n7604 , n7605 , n7606 , n7607 , n7608 , n7609 , n7610 , n7611 , n7612 , n7613 , n7614 , n7615 , n7616 , n7617 , n7618 , n7619 , n7620 , n7621 , n7622 , n7623 , n7624 , n7625 , n7626 , n7627 , n7628 , n7629 , n7630 , n7631 , n7632 , n7633 , n7634 , n7635 , n7636 , n7637 , n7638 , n7639 , n7640 , n7641 , n7642 , n7643 , n7644 , n7645 , n7646 , n7647 , n7648 , n7649 , n7650 , n7651 , n7652 , n7653 , n7654 , n7655 , n7656 , n7657 , n7658 , n7659 , n7660 , n7661 , n7662 , n7663 , n7664 , n7665 , n7666 , n7667 , n7668 , n7669 , n7670 , n7671 , n7672 , n7673 , n7674 , n7675 , n7676 , n7677 , n7678 , n7679 , n7680 , n7681 , n7682 , n7683 , n7684 , n7685 , n7686 , n7687 , n7688 , n7689 , n7690 , n7691 , n7692 , n7693 , n7694 , n7695 , n7696 , n7697 , n7698 , n7699 , n7700 , n7701 , n7702 , n7703 , n7704 , n7705 , n7706 , n7707 , n7708 , n7709 , n7710 , n7711 , n7712 , n7713 , n7714 , n7715 , n7716 , n7717 , n7718 , n7719 , n7720 , n7721 , n7722 , n7723 , n7724 , n7725 , n7726 , n7727 , n7728 , n7729 , n7730 , n7731 , n7732 , n7733 , n7734 , n7735 , n7736 , n7737 , n7738 , n7739 , n7740 , n7741 , n7742 , n7743 , n7744 , n7745 , n7746 , n7747 , n7748 , n7749 , n7750 , n7751 , n7752 , n7753 , n7754 , n7755 , n7756 , n7757 , n7758 , n7759 , n7760 , n7761 , n7762 , n7763 , n7764 , n7765 , n7766 , n7767 , n7768 , n7769 , n7770 , n7771 , n7772 , n7773 , n7774 , n7775 , n7776 , n7777 , n7778 , n7779 , n7780 , n7781 , n7782 , n7783 , n7784 , n7785 , n7786 , n7787 , n7788 , n7789 , n7790 , n7791 , n7792 , n7793 , n7794 , n7795 , n7796 , n7797 , n7798 , n7799 , n7800 , n7801 , n7802 , n7803 , n7804 , n7805 , n7806 , n7807 , n7808 , n7809 , n7810 , n7811 , n7812 , n7813 , n7814 , n7815 , n7816 , n7817 , n7818 , n7819 , n7820 , n7821 , n7822 , n7823 , n7824 , n7825 , n7826 , n7827 , n7828 , n7829 , n7830 , n7831 , n7832 , n7833 , n7834 , n7835 , n7836 , n7837 , n7838 , n7839 , n7840 , n7841 , n7842 , n7843 , n7844 , n7845 , n7846 , n7847 , n7848 , n7849 , n7850 , n7851 , n7852 , n7853 , n7854 , n7855 , n7856 , n7857 , n7858 , n7859 , n7860 , n7861 , n7862 , n7863 , n7864 , n7865 , n7866 , n7867 , n7868 , n7869 , n7870 , n7871 , n7872 , n7873 , n7874 , n7875 , n7876 , n7877 , n7878 , n7879 , n7880 , n7881 , n7882 , n7883 , n7884 , n7885 , n7886 , n7887 , n7888 , n7889 , n7890 , n7891 , n7892 , n7893 , n7894 , n7895 , n7896 , n7897 , n7898 , n7899 , n7900 , n7901 , n7902 , n7903 , n7904 , n7905 , n7906 , n7907 , n7908 , n7909 , n7910 , n7911 , n7912 , n7913 , n7914 , n7915 , n7916 , n7917 , n7918 , n7919 , n7920 , n7921 , n7922 , n7923 , n7924 , n7925 , n7926 , n7927 , n7928 , n7929 , n7930 , n7931 , n7932 , n7933 , n7934 , n7935 , n7936 , n7937 , n7938 , n7939 , n7940 , n7941 , n7942 , n7943 , n7944 , n7945 , n7946 , n7947 , n7948 , n7949 , n7950 , n7951 , n7952 , n7953 , n7954 , n7955 , n7956 , n7957 , n7958 , n7959 , n7960 , n7961 , n7962 , n7963 , n7964 , n7965 , n7966 , n7967 , n7968 , n7969 , n7970 , n7971 , n7972 , n7973 , n7974 , n7975 , n7976 , n7977 , n7978 , n7979 , n7980 , n7981 , n7982 , n7983 , n7984 , n7985 , n7986 , n7987 , n7988 , n7989 , n7990 , n7991 , n7992 , n7993 , n7994 , n7995 , n7996 , n7997 , n7998 , n7999 , n8000 , n8001 , n8002 , n8003 , n8004 , n8005 , n8006 , n8007 , n8008 , n8009 , n8010 , n8011 , n8012 , n8013 , n8014 , n8015 , n8016 , n8017 , n8018 , n8019 , n8020 , n8021 , n8022 , n8023 , n8024 , n8025 , n8026 , n8027 , n8028 , n8029 , n8030 , n8031 , n8032 , n8033 , n8034 , n8035 , n8036 , n8037 , n8038 , n8039 , n8040 , n8041 , n8042 , n8043 , n8044 , n8045 , n8046 , n8047 , n8048 , n8049 , n8050 , n8051 , n8052 , n8053 , n8054 , n8055 , n8056 , n8057 , n8058 , n8059 , n8060 , n8061 , n8062 , n8063 , n8064 , n8065 , n8066 , n8067 , n8068 , n8069 , n8070 , n8071 , n8072 , n8073 , n8074 , n8075 , n8076 , n8077 , n8078 , n8079 , n8080 , n8081 , n8082 , n8083 , n8084 , n8085 , n8086 , n8087 , n8088 , n8089 , n8090 , n8091 , n8092 , n8093 , n8094 , n8095 , n8096 , n8097 , n8098 , n8099 , n8100 , n8101 , n8102 , n8103 , n8104 , n8105 , n8106 , n8107 , n8108 , n8109 , n8110 , n8111 , n8112 , n8113 , n8114 , n8115 , n8116 , n8117 , n8118 , n8119 , n8120 , n8121 , n8122 , n8123 , n8124 , n8125 , n8126 , n8127 , n8128 , n8129 , n8130 , n8131 , n8132 , n8133 , n8134 , n8135 , n8136 , n8137 , n8138 , n8139 , n8140 , n8141 , n8142 , n8143 , n8144 , n8145 , n8146 , n8147 , n8148 , n8149 , n8150 , n8151 , n8152 , n8153 , n8154 , n8155 , n8156 , n8157 , n8158 , n8159 , n8160 , n8161 , n8162 , n8163 , n8164 , n8165 , n8166 , n8167 , n8168 , n8169 , n8170 , n8171 , n8172 , n8173 , n8174 , n8175 , n8176 , n8177 , n8178 , n8179 , n8180 , n8181 , n8182 , n8183 , n8184 , n8185 , n8186 , n8187 , n8188 , n8189 , n8190 , n8191 , n8192 , n8193 , n8194 , n8195 , n8196 , n8197 , n8198 , n8199 , n8200 , n8201 , n8202 , n8203 , n8204 , n8205 , n8206 , n8207 , n8208 , n8209 , n8210 , n8211 , n8212 , n8213 , n8214 , n8215 , n8216 , n8217 , n8218 , n8219 , n8220 , n8221 , n8222 , n8223 , n8224 , n8225 , n8226 , n8227 , n8228 , n8229 , n8230 , n8231 , n8232 , n8233 , n8234 , n8235 , n8236 , n8237 , n8238 , n8239 , n8240 , n8241 , n8242 , n8243 , n8244 , n8245 , n8246 , n8247 , n8248 , n8249 , n8250 , n8251 , n8252 , n8253 , n8254 , n8255 , n8256 , n8257 , n8258 , n8259 , n8260 , n8261 , n8262 , n8263 , n8264 , n8265 , n8266 , n8267 , n8268 , n8269 , n8270 , n8271 , n8272 , n8273 , n8274 , n8275 , n8276 , n8277 , n8278 , n8279 , n8280 , n8281 , n8282 , n8283 , n8284 , n8285 , n8286 , n8287 , n8288 , n8289 , n8290 , n8291 , n8292 , n8293 , n8294 , n8295 , n8296 , n8297 , n8298 , n8299 , n8300 , n8301 , n8302 , n8303 , n8304 , n8305 , n8306 , n8307 , n8308 , n8309 , n8310 , n8311 , n8312 , n8313 , n8314 , n8315 , n8316 , n8317 , n8318 , n8319 , n8320 , n8321 , n8322 , n8323 , n8324 , n8325 , n8326 , n8327 , n8328 , n8329 , n8330 , n8331 , n8332 , n8333 , n8334 , n8335 , n8336 , n8337 , n8338 , n8339 , n8340 , n8341 , n8342 , n8343 , n8344 , n8345 , n8346 , n8347 , n8348 , n8349 , n8350 , n8351 , n8352 , n8353 , n8354 , n8355 , n8356 , n8357 , n8358 , n8359 , n8360 , n8361 , n8362 , n8363 , n8364 , n8365 , n8366 , n8367 , n8368 , n8369 , n8370 , n8371 , n8372 , n8373 , n8374 , n8375 , n8376 , n8377 , n8378 , n8379 , n8380 , n8381 , n8382 , n8383 , n8384 , n8385 , n8386 , n8387 , n8388 , n8389 , n8390 , n8391 , n8392 , n8393 , n8394 , n8395 , n8396 , n8397 , n8398 , n8399 , n8400 , n8401 , n8402 , n8403 , n8404 , n8405 , n8406 , n8407 , n8408 , n8409 , n8410 , n8411 , n8412 , n8413 , n8414 , n8415 , n8416 , n8417 , n8418 , n8419 , n8420 , n8421 , n8422 , n8423 , n8424 , n8425 , n8426 , n8427 , n8428 , n8429 , n8430 , n8431 , n8432 , n8433 , n8434 , n8435 , n8436 , n8437 , n8438 , n8439 , n8440 , n8441 , n8442 , n8443 , n8444 , n8445 , n8446 , n8447 , n8448 , n8449 , n8450 , n8451 , n8452 , n8453 , n8454 , n8455 , n8456 , n8457 , n8458 , n8459 , n8460 , n8461 , n8462 , n8463 , n8464 , n8465 , n8466 , n8467 , n8468 , n8469 , n8470 , n8471 , n8472 , n8473 , n8474 , n8475 , n8476 , n8477 , n8478 , n8479 , n8480 , n8481 , n8482 , n8483 , n8484 , n8485 , n8486 , n8487 , n8488 , n8489 , n8490 , n8491 , n8492 , n8493 , n8494 , n8495 , n8496 , n8497 , n8498 , n8499 , n8500 , n8501 , n8502 , n8503 , n8504 , n8505 , n8506 , n8507 , n8508 , n8509 , n8510 , n8511 , n8512 , n8513 , n8514 , n8515 , n8516 , n8517 , n8518 , n8519 , n8520 , n8521 , n8522 , n8523 , n8524 , n8525 , n8526 , n8527 , n8528 , n8529 , n8530 , n8531 , n8532 , n8533 , n8534 , n8535 , n8536 , n8537 , n8538 , n8539 , n8540 , n8541 , n8542 , n8543 , n8544 , n8545 , n8546 , n8547 , n8548 , n8549 , n8550 , n8551 , n8552 , n8553 , n8554 , n8555 , n8556 , n8557 , n8558 , n8559 , n8560 , n8561 , n8562 , n8563 , n8564 , n8565 , n8566 , n8567 , n8568 , n8569 , n8570 , n8571 , n8572 , n8573 , n8574 , n8575 , n8576 , n8577 , n8578 , n8579 , n8580 , n8581 , n8582 , n8583 , n8584 , n8585 , n8586 , n8587 , n8588 , n8589 , n8590 , n8591 , n8592 , n8593 , n8594 , n8595 , n8596 , n8597 , n8598 , n8599 , n8600 , n8601 , n8602 , n8603 , n8604 , n8605 , n8606 , n8607 , n8608 , n8609 , n8610 , n8611 , n8612 , n8613 , n8614 , n8615 , n8616 , n8617 , n8618 , n8619 , n8620 , n8621 , n8622 , n8623 , n8624 , n8625 , n8626 , n8627 , n8628 , n8629 , n8630 , n8631 , n8632 , n8633 , n8634 , n8635 , n8636 , n8637 , n8638 , n8639 , n8640 , n8641 , n8642 , n8643 , n8644 , n8645 , n8646 , n8647 , n8648 , n8649 , n8650 , n8651 , n8652 , n8653 , n8654 , n8655 , n8656 , n8657 , n8658 , n8659 , n8660 , n8661 , n8662 , n8663 , n8664 , n8665 , n8666 , n8667 , n8668 , n8669 , n8670 , n8671 , n8672 , n8673 , n8674 , n8675 , n8676 , n8677 , n8678 , n8679 , n8680 , n8681 , n8682 , n8683 , n8684 , n8685 , n8686 , n8687 , n8688 , n8689 , n8690 , n8691 , n8692 , n8693 , n8694 , n8695 , n8696 , n8697 , n8698 , n8699 , n8700 , n8701 , n8702 , n8703 , n8704 , n8705 , n8706 , n8707 , n8708 , n8709 , n8710 ;
  assign n1508 = \TM0_pad  & ~\WX10891_reg/NET0131  ;
  assign n1509 = \WX835_reg/NET0131  & ~\WX899_reg/NET0131  ;
  assign n1510 = ~\WX835_reg/NET0131  & \WX899_reg/NET0131  ;
  assign n1511 = ~n1509 & ~n1510 ;
  assign n1512 = \WX707_reg/NET0131  & ~\WX771_reg/NET0131  ;
  assign n1513 = ~\WX707_reg/NET0131  & \WX771_reg/NET0131  ;
  assign n1514 = ~n1512 & ~n1513 ;
  assign n1515 = n1511 & n1514 ;
  assign n1516 = ~n1511 & ~n1514 ;
  assign n1517 = ~n1515 & ~n1516 ;
  assign n1518 = n1508 & n1517 ;
  assign n1519 = ~n1508 & ~n1517 ;
  assign n1520 = ~n1518 & ~n1519 ;
  assign n1521 = \TM0_pad  & ~\WX10871_reg/NET0131  ;
  assign n1522 = \WX815_reg/NET0131  & ~\WX879_reg/NET0131  ;
  assign n1523 = ~\WX815_reg/NET0131  & \WX879_reg/NET0131  ;
  assign n1524 = ~n1522 & ~n1523 ;
  assign n1525 = \WX687_reg/NET0131  & ~\WX751_reg/NET0131  ;
  assign n1526 = ~\WX687_reg/NET0131  & \WX751_reg/NET0131  ;
  assign n1527 = ~n1525 & ~n1526 ;
  assign n1528 = n1524 & n1527 ;
  assign n1529 = ~n1524 & ~n1527 ;
  assign n1530 = ~n1528 & ~n1529 ;
  assign n1531 = n1521 & n1530 ;
  assign n1532 = ~n1521 & ~n1530 ;
  assign n1533 = ~n1531 & ~n1532 ;
  assign n1534 = \TM0_pad  & ~\WX10869_reg/NET0131  ;
  assign n1535 = \WX813_reg/NET0131  & ~\WX877_reg/NET0131  ;
  assign n1536 = ~\WX813_reg/NET0131  & \WX877_reg/NET0131  ;
  assign n1537 = ~n1535 & ~n1536 ;
  assign n1538 = \WX685_reg/NET0131  & ~\WX749_reg/NET0131  ;
  assign n1539 = ~\WX685_reg/NET0131  & \WX749_reg/NET0131  ;
  assign n1540 = ~n1538 & ~n1539 ;
  assign n1541 = n1537 & n1540 ;
  assign n1542 = ~n1537 & ~n1540 ;
  assign n1543 = ~n1541 & ~n1542 ;
  assign n1544 = n1534 & n1543 ;
  assign n1545 = ~n1534 & ~n1543 ;
  assign n1546 = ~n1544 & ~n1545 ;
  assign n1547 = \TM0_pad  & ~\WX10867_reg/NET0131  ;
  assign n1548 = \WX811_reg/NET0131  & ~\WX875_reg/NET0131  ;
  assign n1549 = ~\WX811_reg/NET0131  & \WX875_reg/NET0131  ;
  assign n1550 = ~n1548 & ~n1549 ;
  assign n1551 = \WX683_reg/NET0131  & ~\WX747_reg/NET0131  ;
  assign n1552 = ~\WX683_reg/NET0131  & \WX747_reg/NET0131  ;
  assign n1553 = ~n1551 & ~n1552 ;
  assign n1554 = n1550 & n1553 ;
  assign n1555 = ~n1550 & ~n1553 ;
  assign n1556 = ~n1554 & ~n1555 ;
  assign n1557 = n1547 & n1556 ;
  assign n1558 = ~n1547 & ~n1556 ;
  assign n1559 = ~n1557 & ~n1558 ;
  assign n1560 = \TM0_pad  & ~\WX10865_reg/NET0131  ;
  assign n1561 = \WX809_reg/NET0131  & ~\WX873_reg/NET0131  ;
  assign n1562 = ~\WX809_reg/NET0131  & \WX873_reg/NET0131  ;
  assign n1563 = ~n1561 & ~n1562 ;
  assign n1564 = \WX681_reg/NET0131  & ~\WX745_reg/NET0131  ;
  assign n1565 = ~\WX681_reg/NET0131  & \WX745_reg/NET0131  ;
  assign n1566 = ~n1564 & ~n1565 ;
  assign n1567 = n1563 & n1566 ;
  assign n1568 = ~n1563 & ~n1566 ;
  assign n1569 = ~n1567 & ~n1568 ;
  assign n1570 = n1560 & n1569 ;
  assign n1571 = ~n1560 & ~n1569 ;
  assign n1572 = ~n1570 & ~n1571 ;
  assign n1573 = \TM0_pad  & ~\WX10863_reg/NET0131  ;
  assign n1574 = \WX807_reg/NET0131  & ~\WX871_reg/NET0131  ;
  assign n1575 = ~\WX807_reg/NET0131  & \WX871_reg/NET0131  ;
  assign n1576 = ~n1574 & ~n1575 ;
  assign n1577 = \WX679_reg/NET0131  & ~\WX743_reg/NET0131  ;
  assign n1578 = ~\WX679_reg/NET0131  & \WX743_reg/NET0131  ;
  assign n1579 = ~n1577 & ~n1578 ;
  assign n1580 = n1576 & n1579 ;
  assign n1581 = ~n1576 & ~n1579 ;
  assign n1582 = ~n1580 & ~n1581 ;
  assign n1583 = n1573 & n1582 ;
  assign n1584 = ~n1573 & ~n1582 ;
  assign n1585 = ~n1583 & ~n1584 ;
  assign n1586 = \TM0_pad  & ~\WX10861_reg/NET0131  ;
  assign n1587 = \WX805_reg/NET0131  & ~\WX869_reg/NET0131  ;
  assign n1588 = ~\WX805_reg/NET0131  & \WX869_reg/NET0131  ;
  assign n1589 = ~n1587 & ~n1588 ;
  assign n1590 = \WX677_reg/NET0131  & ~\WX741_reg/NET0131  ;
  assign n1591 = ~\WX677_reg/NET0131  & \WX741_reg/NET0131  ;
  assign n1592 = ~n1590 & ~n1591 ;
  assign n1593 = n1589 & n1592 ;
  assign n1594 = ~n1589 & ~n1592 ;
  assign n1595 = ~n1593 & ~n1594 ;
  assign n1596 = n1586 & n1595 ;
  assign n1597 = ~n1586 & ~n1595 ;
  assign n1598 = ~n1596 & ~n1597 ;
  assign n1599 = \WX803_reg/NET0131  & ~\WX867_reg/NET0131  ;
  assign n1600 = ~\WX803_reg/NET0131  & \WX867_reg/NET0131  ;
  assign n1601 = ~n1599 & ~n1600 ;
  assign n1602 = \WX739_reg/NET0131  & ~n1601 ;
  assign n1603 = ~\WX739_reg/NET0131  & n1601 ;
  assign n1604 = ~n1602 & ~n1603 ;
  assign n1605 = \TM0_pad  & \WX10859_reg/NET0131  ;
  assign n1606 = ~\TM1_pad  & ~\WX675_reg/NET0131  ;
  assign n1607 = \TM1_pad  & \WX675_reg/NET0131  ;
  assign n1608 = ~n1606 & ~n1607 ;
  assign n1609 = n1605 & ~n1608 ;
  assign n1610 = ~n1605 & n1608 ;
  assign n1611 = ~n1609 & ~n1610 ;
  assign n1612 = n1604 & n1611 ;
  assign n1613 = ~n1604 & ~n1611 ;
  assign n1614 = ~n1612 & ~n1613 ;
  assign n1615 = \WX801_reg/NET0131  & ~\WX865_reg/NET0131  ;
  assign n1616 = ~\WX801_reg/NET0131  & \WX865_reg/NET0131  ;
  assign n1617 = ~n1615 & ~n1616 ;
  assign n1618 = \WX737_reg/NET0131  & ~n1617 ;
  assign n1619 = ~\WX737_reg/NET0131  & n1617 ;
  assign n1620 = ~n1618 & ~n1619 ;
  assign n1621 = \TM0_pad  & \WX10857_reg/NET0131  ;
  assign n1622 = ~\TM1_pad  & ~\WX673_reg/NET0131  ;
  assign n1623 = \TM1_pad  & \WX673_reg/NET0131  ;
  assign n1624 = ~n1622 & ~n1623 ;
  assign n1625 = n1621 & ~n1624 ;
  assign n1626 = ~n1621 & n1624 ;
  assign n1627 = ~n1625 & ~n1626 ;
  assign n1628 = n1620 & n1627 ;
  assign n1629 = ~n1620 & ~n1627 ;
  assign n1630 = ~n1628 & ~n1629 ;
  assign n1631 = \WX799_reg/NET0131  & ~\WX863_reg/NET0131  ;
  assign n1632 = ~\WX799_reg/NET0131  & \WX863_reg/NET0131  ;
  assign n1633 = ~n1631 & ~n1632 ;
  assign n1634 = \WX735_reg/NET0131  & ~n1633 ;
  assign n1635 = ~\WX735_reg/NET0131  & n1633 ;
  assign n1636 = ~n1634 & ~n1635 ;
  assign n1637 = \TM0_pad  & \WX10855_reg/NET0131  ;
  assign n1638 = ~\TM1_pad  & ~\WX671_reg/NET0131  ;
  assign n1639 = \TM1_pad  & \WX671_reg/NET0131  ;
  assign n1640 = ~n1638 & ~n1639 ;
  assign n1641 = n1637 & ~n1640 ;
  assign n1642 = ~n1637 & n1640 ;
  assign n1643 = ~n1641 & ~n1642 ;
  assign n1644 = n1636 & n1643 ;
  assign n1645 = ~n1636 & ~n1643 ;
  assign n1646 = ~n1644 & ~n1645 ;
  assign n1647 = \WX797_reg/NET0131  & ~\WX861_reg/NET0131  ;
  assign n1648 = ~\WX797_reg/NET0131  & \WX861_reg/NET0131  ;
  assign n1649 = ~n1647 & ~n1648 ;
  assign n1650 = \WX733_reg/NET0131  & ~n1649 ;
  assign n1651 = ~\WX733_reg/NET0131  & n1649 ;
  assign n1652 = ~n1650 & ~n1651 ;
  assign n1653 = \TM0_pad  & \WX10853_reg/NET0131  ;
  assign n1654 = ~\TM1_pad  & ~\WX669_reg/NET0131  ;
  assign n1655 = \TM1_pad  & \WX669_reg/NET0131  ;
  assign n1656 = ~n1654 & ~n1655 ;
  assign n1657 = n1653 & ~n1656 ;
  assign n1658 = ~n1653 & n1656 ;
  assign n1659 = ~n1657 & ~n1658 ;
  assign n1660 = n1652 & n1659 ;
  assign n1661 = ~n1652 & ~n1659 ;
  assign n1662 = ~n1660 & ~n1661 ;
  assign n1663 = \TM0_pad  & ~\WX10889_reg/NET0131  ;
  assign n1664 = \WX833_reg/NET0131  & ~\WX897_reg/NET0131  ;
  assign n1665 = ~\WX833_reg/NET0131  & \WX897_reg/NET0131  ;
  assign n1666 = ~n1664 & ~n1665 ;
  assign n1667 = \WX705_reg/NET0131  & ~\WX769_reg/NET0131  ;
  assign n1668 = ~\WX705_reg/NET0131  & \WX769_reg/NET0131  ;
  assign n1669 = ~n1667 & ~n1668 ;
  assign n1670 = n1666 & n1669 ;
  assign n1671 = ~n1666 & ~n1669 ;
  assign n1672 = ~n1670 & ~n1671 ;
  assign n1673 = n1663 & n1672 ;
  assign n1674 = ~n1663 & ~n1672 ;
  assign n1675 = ~n1673 & ~n1674 ;
  assign n1676 = \WX795_reg/NET0131  & ~\WX859_reg/NET0131  ;
  assign n1677 = ~\WX795_reg/NET0131  & \WX859_reg/NET0131  ;
  assign n1678 = ~n1676 & ~n1677 ;
  assign n1679 = \WX731_reg/NET0131  & ~n1678 ;
  assign n1680 = ~\WX731_reg/NET0131  & n1678 ;
  assign n1681 = ~n1679 & ~n1680 ;
  assign n1682 = \TM0_pad  & \WX10851_reg/NET0131  ;
  assign n1683 = ~\TM1_pad  & ~\WX667_reg/NET0131  ;
  assign n1684 = \TM1_pad  & \WX667_reg/NET0131  ;
  assign n1685 = ~n1683 & ~n1684 ;
  assign n1686 = n1682 & ~n1685 ;
  assign n1687 = ~n1682 & n1685 ;
  assign n1688 = ~n1686 & ~n1687 ;
  assign n1689 = n1681 & n1688 ;
  assign n1690 = ~n1681 & ~n1688 ;
  assign n1691 = ~n1689 & ~n1690 ;
  assign n1692 = \WX793_reg/NET0131  & ~\WX857_reg/NET0131  ;
  assign n1693 = ~\WX793_reg/NET0131  & \WX857_reg/NET0131  ;
  assign n1694 = ~n1692 & ~n1693 ;
  assign n1695 = \WX729_reg/NET0131  & ~n1694 ;
  assign n1696 = ~\WX729_reg/NET0131  & n1694 ;
  assign n1697 = ~n1695 & ~n1696 ;
  assign n1698 = \TM0_pad  & \WX10849_reg/NET0131  ;
  assign n1699 = ~\TM1_pad  & ~\WX665_reg/NET0131  ;
  assign n1700 = \TM1_pad  & \WX665_reg/NET0131  ;
  assign n1701 = ~n1699 & ~n1700 ;
  assign n1702 = n1698 & ~n1701 ;
  assign n1703 = ~n1698 & n1701 ;
  assign n1704 = ~n1702 & ~n1703 ;
  assign n1705 = n1697 & n1704 ;
  assign n1706 = ~n1697 & ~n1704 ;
  assign n1707 = ~n1705 & ~n1706 ;
  assign n1708 = \WX791_reg/NET0131  & ~\WX855_reg/NET0131  ;
  assign n1709 = ~\WX791_reg/NET0131  & \WX855_reg/NET0131  ;
  assign n1710 = ~n1708 & ~n1709 ;
  assign n1711 = \WX727_reg/NET0131  & ~n1710 ;
  assign n1712 = ~\WX727_reg/NET0131  & n1710 ;
  assign n1713 = ~n1711 & ~n1712 ;
  assign n1714 = \TM0_pad  & \WX10847_reg/NET0131  ;
  assign n1715 = ~\TM1_pad  & ~\WX663_reg/NET0131  ;
  assign n1716 = \TM1_pad  & \WX663_reg/NET0131  ;
  assign n1717 = ~n1715 & ~n1716 ;
  assign n1718 = n1714 & ~n1717 ;
  assign n1719 = ~n1714 & n1717 ;
  assign n1720 = ~n1718 & ~n1719 ;
  assign n1721 = n1713 & n1720 ;
  assign n1722 = ~n1713 & ~n1720 ;
  assign n1723 = ~n1721 & ~n1722 ;
  assign n1724 = \WX789_reg/NET0131  & ~\WX853_reg/NET0131  ;
  assign n1725 = ~\WX789_reg/NET0131  & \WX853_reg/NET0131  ;
  assign n1726 = ~n1724 & ~n1725 ;
  assign n1727 = \WX725_reg/NET0131  & ~n1726 ;
  assign n1728 = ~\WX725_reg/NET0131  & n1726 ;
  assign n1729 = ~n1727 & ~n1728 ;
  assign n1730 = \TM0_pad  & \WX10845_reg/NET0131  ;
  assign n1731 = ~\TM1_pad  & ~\WX661_reg/NET0131  ;
  assign n1732 = \TM1_pad  & \WX661_reg/NET0131  ;
  assign n1733 = ~n1731 & ~n1732 ;
  assign n1734 = n1730 & ~n1733 ;
  assign n1735 = ~n1730 & n1733 ;
  assign n1736 = ~n1734 & ~n1735 ;
  assign n1737 = n1729 & n1736 ;
  assign n1738 = ~n1729 & ~n1736 ;
  assign n1739 = ~n1737 & ~n1738 ;
  assign n1740 = \WX787_reg/NET0131  & ~\WX851_reg/NET0131  ;
  assign n1741 = ~\WX787_reg/NET0131  & \WX851_reg/NET0131  ;
  assign n1742 = ~n1740 & ~n1741 ;
  assign n1743 = \WX723_reg/NET0131  & ~n1742 ;
  assign n1744 = ~\WX723_reg/NET0131  & n1742 ;
  assign n1745 = ~n1743 & ~n1744 ;
  assign n1746 = \TM0_pad  & \WX10843_reg/NET0131  ;
  assign n1747 = ~\TM1_pad  & ~\WX659_reg/NET0131  ;
  assign n1748 = \TM1_pad  & \WX659_reg/NET0131  ;
  assign n1749 = ~n1747 & ~n1748 ;
  assign n1750 = n1746 & ~n1749 ;
  assign n1751 = ~n1746 & n1749 ;
  assign n1752 = ~n1750 & ~n1751 ;
  assign n1753 = n1745 & n1752 ;
  assign n1754 = ~n1745 & ~n1752 ;
  assign n1755 = ~n1753 & ~n1754 ;
  assign n1756 = \WX785_reg/NET0131  & ~\WX849_reg/NET0131  ;
  assign n1757 = ~\WX785_reg/NET0131  & \WX849_reg/NET0131  ;
  assign n1758 = ~n1756 & ~n1757 ;
  assign n1759 = \WX721_reg/NET0131  & ~n1758 ;
  assign n1760 = ~\WX721_reg/NET0131  & n1758 ;
  assign n1761 = ~n1759 & ~n1760 ;
  assign n1762 = \TM0_pad  & \WX10841_reg/NET0131  ;
  assign n1763 = ~\TM1_pad  & ~\WX657_reg/NET0131  ;
  assign n1764 = \TM1_pad  & \WX657_reg/NET0131  ;
  assign n1765 = ~n1763 & ~n1764 ;
  assign n1766 = n1762 & ~n1765 ;
  assign n1767 = ~n1762 & n1765 ;
  assign n1768 = ~n1766 & ~n1767 ;
  assign n1769 = n1761 & n1768 ;
  assign n1770 = ~n1761 & ~n1768 ;
  assign n1771 = ~n1769 & ~n1770 ;
  assign n1772 = \WX783_reg/NET0131  & ~\WX847_reg/NET0131  ;
  assign n1773 = ~\WX783_reg/NET0131  & \WX847_reg/NET0131  ;
  assign n1774 = ~n1772 & ~n1773 ;
  assign n1775 = \WX719_reg/NET0131  & ~n1774 ;
  assign n1776 = ~\WX719_reg/NET0131  & n1774 ;
  assign n1777 = ~n1775 & ~n1776 ;
  assign n1778 = \TM0_pad  & \WX10839_reg/NET0131  ;
  assign n1779 = ~\TM1_pad  & ~\WX655_reg/NET0131  ;
  assign n1780 = \TM1_pad  & \WX655_reg/NET0131  ;
  assign n1781 = ~n1779 & ~n1780 ;
  assign n1782 = n1778 & ~n1781 ;
  assign n1783 = ~n1778 & n1781 ;
  assign n1784 = ~n1782 & ~n1783 ;
  assign n1785 = n1777 & n1784 ;
  assign n1786 = ~n1777 & ~n1784 ;
  assign n1787 = ~n1785 & ~n1786 ;
  assign n1788 = \WX781_reg/NET0131  & ~\WX845_reg/NET0131  ;
  assign n1789 = ~\WX781_reg/NET0131  & \WX845_reg/NET0131  ;
  assign n1790 = ~n1788 & ~n1789 ;
  assign n1791 = \WX717_reg/NET0131  & ~n1790 ;
  assign n1792 = ~\WX717_reg/NET0131  & n1790 ;
  assign n1793 = ~n1791 & ~n1792 ;
  assign n1794 = \TM0_pad  & \WX10837_reg/NET0131  ;
  assign n1795 = ~\TM1_pad  & ~\WX653_reg/NET0131  ;
  assign n1796 = \TM1_pad  & \WX653_reg/NET0131  ;
  assign n1797 = ~n1795 & ~n1796 ;
  assign n1798 = n1794 & ~n1797 ;
  assign n1799 = ~n1794 & n1797 ;
  assign n1800 = ~n1798 & ~n1799 ;
  assign n1801 = n1793 & n1800 ;
  assign n1802 = ~n1793 & ~n1800 ;
  assign n1803 = ~n1801 & ~n1802 ;
  assign n1804 = \WX779_reg/NET0131  & ~\WX843_reg/NET0131  ;
  assign n1805 = ~\WX779_reg/NET0131  & \WX843_reg/NET0131  ;
  assign n1806 = ~n1804 & ~n1805 ;
  assign n1807 = \WX715_reg/NET0131  & ~n1806 ;
  assign n1808 = ~\WX715_reg/NET0131  & n1806 ;
  assign n1809 = ~n1807 & ~n1808 ;
  assign n1810 = \TM0_pad  & \WX10835_reg/NET0131  ;
  assign n1811 = ~\TM1_pad  & ~\WX651_reg/NET0131  ;
  assign n1812 = \TM1_pad  & \WX651_reg/NET0131  ;
  assign n1813 = ~n1811 & ~n1812 ;
  assign n1814 = n1810 & ~n1813 ;
  assign n1815 = ~n1810 & n1813 ;
  assign n1816 = ~n1814 & ~n1815 ;
  assign n1817 = n1809 & n1816 ;
  assign n1818 = ~n1809 & ~n1816 ;
  assign n1819 = ~n1817 & ~n1818 ;
  assign n1820 = \WX777_reg/NET0131  & ~\WX841_reg/NET0131  ;
  assign n1821 = ~\WX777_reg/NET0131  & \WX841_reg/NET0131  ;
  assign n1822 = ~n1820 & ~n1821 ;
  assign n1823 = \WX713_reg/NET0131  & ~n1822 ;
  assign n1824 = ~\WX713_reg/NET0131  & n1822 ;
  assign n1825 = ~n1823 & ~n1824 ;
  assign n1826 = \TM0_pad  & \WX10833_reg/NET0131  ;
  assign n1827 = ~\TM1_pad  & ~\WX649_reg/NET0131  ;
  assign n1828 = \TM1_pad  & \WX649_reg/NET0131  ;
  assign n1829 = ~n1827 & ~n1828 ;
  assign n1830 = n1826 & ~n1829 ;
  assign n1831 = ~n1826 & n1829 ;
  assign n1832 = ~n1830 & ~n1831 ;
  assign n1833 = n1825 & n1832 ;
  assign n1834 = ~n1825 & ~n1832 ;
  assign n1835 = ~n1833 & ~n1834 ;
  assign n1836 = \TM0_pad  & ~\WX10887_reg/NET0131  ;
  assign n1837 = \WX831_reg/NET0131  & ~\WX895_reg/NET0131  ;
  assign n1838 = ~\WX831_reg/NET0131  & \WX895_reg/NET0131  ;
  assign n1839 = ~n1837 & ~n1838 ;
  assign n1840 = \WX703_reg/NET0131  & ~\WX767_reg/NET0131  ;
  assign n1841 = ~\WX703_reg/NET0131  & \WX767_reg/NET0131  ;
  assign n1842 = ~n1840 & ~n1841 ;
  assign n1843 = n1839 & n1842 ;
  assign n1844 = ~n1839 & ~n1842 ;
  assign n1845 = ~n1843 & ~n1844 ;
  assign n1846 = n1836 & n1845 ;
  assign n1847 = ~n1836 & ~n1845 ;
  assign n1848 = ~n1846 & ~n1847 ;
  assign n1849 = \WX775_reg/NET0131  & ~\WX839_reg/NET0131  ;
  assign n1850 = ~\WX775_reg/NET0131  & \WX839_reg/NET0131  ;
  assign n1851 = ~n1849 & ~n1850 ;
  assign n1852 = \WX711_reg/NET0131  & ~n1851 ;
  assign n1853 = ~\WX711_reg/NET0131  & n1851 ;
  assign n1854 = ~n1852 & ~n1853 ;
  assign n1855 = \TM0_pad  & \WX10831_reg/NET0131  ;
  assign n1856 = ~\TM1_pad  & ~\WX647_reg/NET0131  ;
  assign n1857 = \TM1_pad  & \WX647_reg/NET0131  ;
  assign n1858 = ~n1856 & ~n1857 ;
  assign n1859 = n1855 & ~n1858 ;
  assign n1860 = ~n1855 & n1858 ;
  assign n1861 = ~n1859 & ~n1860 ;
  assign n1862 = n1854 & n1861 ;
  assign n1863 = ~n1854 & ~n1861 ;
  assign n1864 = ~n1862 & ~n1863 ;
  assign n1865 = \WX773_reg/NET0131  & ~\WX837_reg/NET0131  ;
  assign n1866 = ~\WX773_reg/NET0131  & \WX837_reg/NET0131  ;
  assign n1867 = ~n1865 & ~n1866 ;
  assign n1868 = \WX709_reg/NET0131  & ~n1867 ;
  assign n1869 = ~\WX709_reg/NET0131  & n1867 ;
  assign n1870 = ~n1868 & ~n1869 ;
  assign n1871 = \TM0_pad  & \WX10829_reg/NET0131  ;
  assign n1872 = ~\TM1_pad  & ~\WX645_reg/NET0131  ;
  assign n1873 = \TM1_pad  & \WX645_reg/NET0131  ;
  assign n1874 = ~n1872 & ~n1873 ;
  assign n1875 = n1871 & ~n1874 ;
  assign n1876 = ~n1871 & n1874 ;
  assign n1877 = ~n1875 & ~n1876 ;
  assign n1878 = n1870 & n1877 ;
  assign n1879 = ~n1870 & ~n1877 ;
  assign n1880 = ~n1878 & ~n1879 ;
  assign n1881 = \TM0_pad  & ~\WX10885_reg/NET0131  ;
  assign n1882 = \WX829_reg/NET0131  & ~\WX893_reg/NET0131  ;
  assign n1883 = ~\WX829_reg/NET0131  & \WX893_reg/NET0131  ;
  assign n1884 = ~n1882 & ~n1883 ;
  assign n1885 = \WX701_reg/NET0131  & ~\WX765_reg/NET0131  ;
  assign n1886 = ~\WX701_reg/NET0131  & \WX765_reg/NET0131  ;
  assign n1887 = ~n1885 & ~n1886 ;
  assign n1888 = n1884 & n1887 ;
  assign n1889 = ~n1884 & ~n1887 ;
  assign n1890 = ~n1888 & ~n1889 ;
  assign n1891 = n1881 & n1890 ;
  assign n1892 = ~n1881 & ~n1890 ;
  assign n1893 = ~n1891 & ~n1892 ;
  assign n1894 = \TM0_pad  & ~\WX10883_reg/NET0131  ;
  assign n1895 = \WX827_reg/NET0131  & ~\WX891_reg/NET0131  ;
  assign n1896 = ~\WX827_reg/NET0131  & \WX891_reg/NET0131  ;
  assign n1897 = ~n1895 & ~n1896 ;
  assign n1898 = \WX699_reg/NET0131  & ~\WX763_reg/NET0131  ;
  assign n1899 = ~\WX699_reg/NET0131  & \WX763_reg/NET0131  ;
  assign n1900 = ~n1898 & ~n1899 ;
  assign n1901 = n1897 & n1900 ;
  assign n1902 = ~n1897 & ~n1900 ;
  assign n1903 = ~n1901 & ~n1902 ;
  assign n1904 = n1894 & n1903 ;
  assign n1905 = ~n1894 & ~n1903 ;
  assign n1906 = ~n1904 & ~n1905 ;
  assign n1907 = \TM0_pad  & ~\WX10881_reg/NET0131  ;
  assign n1908 = \WX825_reg/NET0131  & ~\WX889_reg/NET0131  ;
  assign n1909 = ~\WX825_reg/NET0131  & \WX889_reg/NET0131  ;
  assign n1910 = ~n1908 & ~n1909 ;
  assign n1911 = \WX697_reg/NET0131  & ~\WX761_reg/NET0131  ;
  assign n1912 = ~\WX697_reg/NET0131  & \WX761_reg/NET0131  ;
  assign n1913 = ~n1911 & ~n1912 ;
  assign n1914 = n1910 & n1913 ;
  assign n1915 = ~n1910 & ~n1913 ;
  assign n1916 = ~n1914 & ~n1915 ;
  assign n1917 = n1907 & n1916 ;
  assign n1918 = ~n1907 & ~n1916 ;
  assign n1919 = ~n1917 & ~n1918 ;
  assign n1920 = \TM0_pad  & ~\WX10879_reg/NET0131  ;
  assign n1921 = \WX823_reg/NET0131  & ~\WX887_reg/NET0131  ;
  assign n1922 = ~\WX823_reg/NET0131  & \WX887_reg/NET0131  ;
  assign n1923 = ~n1921 & ~n1922 ;
  assign n1924 = \WX695_reg/NET0131  & ~\WX759_reg/NET0131  ;
  assign n1925 = ~\WX695_reg/NET0131  & \WX759_reg/NET0131  ;
  assign n1926 = ~n1924 & ~n1925 ;
  assign n1927 = n1923 & n1926 ;
  assign n1928 = ~n1923 & ~n1926 ;
  assign n1929 = ~n1927 & ~n1928 ;
  assign n1930 = n1920 & n1929 ;
  assign n1931 = ~n1920 & ~n1929 ;
  assign n1932 = ~n1930 & ~n1931 ;
  assign n1933 = \TM0_pad  & ~\WX10877_reg/NET0131  ;
  assign n1934 = \WX821_reg/NET0131  & ~\WX885_reg/NET0131  ;
  assign n1935 = ~\WX821_reg/NET0131  & \WX885_reg/NET0131  ;
  assign n1936 = ~n1934 & ~n1935 ;
  assign n1937 = \WX693_reg/NET0131  & ~\WX757_reg/NET0131  ;
  assign n1938 = ~\WX693_reg/NET0131  & \WX757_reg/NET0131  ;
  assign n1939 = ~n1937 & ~n1938 ;
  assign n1940 = n1936 & n1939 ;
  assign n1941 = ~n1936 & ~n1939 ;
  assign n1942 = ~n1940 & ~n1941 ;
  assign n1943 = n1933 & n1942 ;
  assign n1944 = ~n1933 & ~n1942 ;
  assign n1945 = ~n1943 & ~n1944 ;
  assign n1946 = \TM0_pad  & ~\WX10875_reg/NET0131  ;
  assign n1947 = \WX819_reg/NET0131  & ~\WX883_reg/NET0131  ;
  assign n1948 = ~\WX819_reg/NET0131  & \WX883_reg/NET0131  ;
  assign n1949 = ~n1947 & ~n1948 ;
  assign n1950 = \WX691_reg/NET0131  & ~\WX755_reg/NET0131  ;
  assign n1951 = ~\WX691_reg/NET0131  & \WX755_reg/NET0131  ;
  assign n1952 = ~n1950 & ~n1951 ;
  assign n1953 = n1949 & n1952 ;
  assign n1954 = ~n1949 & ~n1952 ;
  assign n1955 = ~n1953 & ~n1954 ;
  assign n1956 = n1946 & n1955 ;
  assign n1957 = ~n1946 & ~n1955 ;
  assign n1958 = ~n1956 & ~n1957 ;
  assign n1959 = \TM0_pad  & ~\WX10873_reg/NET0131  ;
  assign n1960 = \WX817_reg/NET0131  & ~\WX881_reg/NET0131  ;
  assign n1961 = ~\WX817_reg/NET0131  & \WX881_reg/NET0131  ;
  assign n1962 = ~n1960 & ~n1961 ;
  assign n1963 = \WX689_reg/NET0131  & ~\WX753_reg/NET0131  ;
  assign n1964 = ~\WX689_reg/NET0131  & \WX753_reg/NET0131  ;
  assign n1965 = ~n1963 & ~n1964 ;
  assign n1966 = n1962 & n1965 ;
  assign n1967 = ~n1962 & ~n1965 ;
  assign n1968 = ~n1966 & ~n1967 ;
  assign n1969 = n1959 & n1968 ;
  assign n1970 = ~n1959 & ~n1968 ;
  assign n1971 = ~n1969 & ~n1970 ;
  assign n1972 = ~\TM0_pad  & ~n1595 ;
  assign n1973 = RESET_pad & \TM1_pad  ;
  assign n1974 = ~n1586 & n1973 ;
  assign n1975 = ~n1972 & n1974 ;
  assign n1978 = \WX2098_reg/NET0131  & ~\WX2162_reg/NET0131  ;
  assign n1979 = ~\WX2098_reg/NET0131  & \WX2162_reg/NET0131  ;
  assign n1980 = ~n1978 & ~n1979 ;
  assign n1981 = \WX1970_reg/NET0131  & ~\WX2034_reg/NET0131  ;
  assign n1982 = ~\WX1970_reg/NET0131  & \WX2034_reg/NET0131  ;
  assign n1983 = ~n1981 & ~n1982 ;
  assign n1985 = n1980 & ~n1983 ;
  assign n1984 = ~n1980 & n1983 ;
  assign n1986 = ~\TM0_pad  & ~n1984 ;
  assign n1987 = ~n1985 & n1986 ;
  assign n1976 = RESET_pad & ~\TM1_pad  ;
  assign n1977 = \TM0_pad  & ~\_2092__reg/NET0131  ;
  assign n1988 = n1976 & ~n1977 ;
  assign n1989 = ~n1987 & n1988 ;
  assign n1990 = ~n1975 & ~n1989 ;
  assign n1991 = \WX9830_reg/NET0131  & ~\WX9894_reg/NET0131  ;
  assign n1992 = ~\WX9830_reg/NET0131  & \WX9894_reg/NET0131  ;
  assign n1993 = ~n1991 & ~n1992 ;
  assign n1994 = \WX9766_reg/NET0131  & ~n1993 ;
  assign n1995 = ~\WX9766_reg/NET0131  & n1993 ;
  assign n1996 = ~n1994 & ~n1995 ;
  assign n1997 = \TM1_pad  & ~\WX9702_reg/NET0131  ;
  assign n1998 = ~\TM1_pad  & \WX9702_reg/NET0131  ;
  assign n1999 = ~n1997 & ~n1998 ;
  assign n2001 = n1996 & ~n1999 ;
  assign n2000 = ~n1996 & n1999 ;
  assign n2002 = ~\TM0_pad  & ~n2000 ;
  assign n2003 = ~n2001 & n2002 ;
  assign n2004 = ~n1810 & ~n2003 ;
  assign n2005 = n1973 & ~n2004 ;
  assign n2006 = \TM0_pad  & \_2329__reg/NET0131  ;
  assign n2007 = \WX11123_reg/NET0131  & ~\WX11187_reg/NET0131  ;
  assign n2008 = ~\WX11123_reg/NET0131  & \WX11187_reg/NET0131  ;
  assign n2009 = ~n2007 & ~n2008 ;
  assign n2010 = \WX11059_reg/NET0131  & ~n2009 ;
  assign n2011 = ~\WX11059_reg/NET0131  & n2009 ;
  assign n2012 = ~n2010 & ~n2011 ;
  assign n2013 = \TM1_pad  & ~\WX10995_reg/NET0131  ;
  assign n2014 = ~\TM1_pad  & \WX10995_reg/NET0131  ;
  assign n2015 = ~n2013 & ~n2014 ;
  assign n2017 = n2012 & ~n2015 ;
  assign n2016 = ~n2012 & n2015 ;
  assign n2018 = ~\TM0_pad  & ~n2016 ;
  assign n2019 = ~n2017 & n2018 ;
  assign n2020 = ~n2006 & ~n2019 ;
  assign n2021 = n1976 & ~n2020 ;
  assign n2022 = ~n2005 & ~n2021 ;
  assign n2023 = ~n1946 & n1973 ;
  assign n2024 = \WX11163_reg/NET0131  & ~\WX11227_reg/NET0131  ;
  assign n2025 = ~\WX11163_reg/NET0131  & \WX11227_reg/NET0131  ;
  assign n2026 = ~n2024 & ~n2025 ;
  assign n2027 = \WX11035_reg/NET0131  & ~\WX11099_reg/NET0131  ;
  assign n2028 = ~\WX11035_reg/NET0131  & \WX11099_reg/NET0131  ;
  assign n2029 = ~n2027 & ~n2028 ;
  assign n2031 = n2026 & ~n2029 ;
  assign n2030 = ~n2026 & n2029 ;
  assign n2032 = ~\TM0_pad  & ~n2030 ;
  assign n2033 = ~n2031 & n2032 ;
  assign n2034 = n2023 & ~n2033 ;
  assign n2036 = \TM0_pad  & ~\_2341__reg/NET0131  ;
  assign n2035 = ~\DATA_0_8_pad  & ~\TM0_pad  ;
  assign n2037 = n1976 & ~n2035 ;
  assign n2038 = ~n2036 & n2037 ;
  assign n2039 = ~n2034 & ~n2038 ;
  assign n2040 = ~n1560 & n1973 ;
  assign n2041 = \WX11153_reg/NET0131  & ~\WX11217_reg/NET0131  ;
  assign n2042 = ~\WX11153_reg/NET0131  & \WX11217_reg/NET0131  ;
  assign n2043 = ~n2041 & ~n2042 ;
  assign n2044 = \WX11025_reg/NET0131  & ~\WX11089_reg/NET0131  ;
  assign n2045 = ~\WX11025_reg/NET0131  & \WX11089_reg/NET0131  ;
  assign n2046 = ~n2044 & ~n2045 ;
  assign n2048 = n2043 & ~n2046 ;
  assign n2047 = ~n2043 & n2046 ;
  assign n2049 = ~\TM0_pad  & ~n2047 ;
  assign n2050 = ~n2048 & n2049 ;
  assign n2051 = n2040 & ~n2050 ;
  assign n2053 = \TM0_pad  & ~\_2346__reg/NET0131  ;
  assign n2052 = ~\DATA_0_13_pad  & ~\TM0_pad  ;
  assign n2054 = n1976 & ~n2052 ;
  assign n2055 = ~n2053 & n2054 ;
  assign n2056 = ~n2051 & ~n2055 ;
  assign n2057 = ~\TM0_pad  & ~n1864 ;
  assign n2058 = ~n1855 & ~n2057 ;
  assign n2059 = n1973 & ~n2058 ;
  assign n2060 = \TM0_pad  & \_2107__reg/NET0131  ;
  assign n2061 = \WX2068_reg/NET0131  & ~\WX2132_reg/NET0131  ;
  assign n2062 = ~\WX2068_reg/NET0131  & \WX2132_reg/NET0131  ;
  assign n2063 = ~n2061 & ~n2062 ;
  assign n2064 = \WX2004_reg/NET0131  & ~n2063 ;
  assign n2065 = ~\WX2004_reg/NET0131  & n2063 ;
  assign n2066 = ~n2064 & ~n2065 ;
  assign n2067 = \TM1_pad  & ~\WX1940_reg/NET0131  ;
  assign n2068 = ~\TM1_pad  & \WX1940_reg/NET0131  ;
  assign n2069 = ~n2067 & ~n2068 ;
  assign n2071 = n2066 & ~n2069 ;
  assign n2070 = ~n2066 & n2069 ;
  assign n2072 = ~\TM0_pad  & ~n2070 ;
  assign n2073 = ~n2071 & n2072 ;
  assign n2074 = ~n2060 & ~n2073 ;
  assign n2075 = n1976 & ~n2074 ;
  assign n2076 = ~n2059 & ~n2075 ;
  assign n2077 = ~\TM0_pad  & ~n1835 ;
  assign n2078 = ~n1826 & ~n2077 ;
  assign n2079 = n1973 & ~n2078 ;
  assign n2080 = \TM0_pad  & \_2106__reg/NET0131  ;
  assign n2081 = \WX2070_reg/NET0131  & ~\WX2134_reg/NET0131  ;
  assign n2082 = ~\WX2070_reg/NET0131  & \WX2134_reg/NET0131  ;
  assign n2083 = ~n2081 & ~n2082 ;
  assign n2084 = \WX2006_reg/NET0131  & ~n2083 ;
  assign n2085 = ~\WX2006_reg/NET0131  & n2083 ;
  assign n2086 = ~n2084 & ~n2085 ;
  assign n2087 = \TM1_pad  & ~\WX1942_reg/NET0131  ;
  assign n2088 = ~\TM1_pad  & \WX1942_reg/NET0131  ;
  assign n2089 = ~n2087 & ~n2088 ;
  assign n2091 = n2086 & ~n2089 ;
  assign n2090 = ~n2086 & n2089 ;
  assign n2092 = ~\TM0_pad  & ~n2090 ;
  assign n2093 = ~n2091 & n2092 ;
  assign n2094 = ~n2080 & ~n2093 ;
  assign n2095 = n1976 & ~n2094 ;
  assign n2096 = ~n2079 & ~n2095 ;
  assign n2097 = \WX3391_reg/NET0131  & ~\WX3455_reg/NET0131  ;
  assign n2098 = ~\WX3391_reg/NET0131  & \WX3455_reg/NET0131  ;
  assign n2099 = ~n2097 & ~n2098 ;
  assign n2100 = \WX3263_reg/NET0131  & ~\WX3327_reg/NET0131  ;
  assign n2101 = ~\WX3263_reg/NET0131  & \WX3327_reg/NET0131  ;
  assign n2102 = ~n2100 & ~n2101 ;
  assign n2104 = n2099 & ~n2102 ;
  assign n2103 = ~n2099 & n2102 ;
  assign n2105 = ~\TM0_pad  & ~n2103 ;
  assign n2106 = ~n2104 & n2105 ;
  assign n2107 = n1974 & ~n2106 ;
  assign n2109 = \WX4684_reg/NET0131  & ~\WX4748_reg/NET0131  ;
  assign n2110 = ~\WX4684_reg/NET0131  & \WX4748_reg/NET0131  ;
  assign n2111 = ~n2109 & ~n2110 ;
  assign n2112 = \WX4556_reg/NET0131  & ~\WX4620_reg/NET0131  ;
  assign n2113 = ~\WX4556_reg/NET0131  & \WX4620_reg/NET0131  ;
  assign n2114 = ~n2112 & ~n2113 ;
  assign n2116 = n2111 & ~n2114 ;
  assign n2115 = ~n2111 & n2114 ;
  assign n2117 = ~\TM0_pad  & ~n2115 ;
  assign n2118 = ~n2116 & n2117 ;
  assign n2108 = \TM0_pad  & ~\_2156__reg/NET0131  ;
  assign n2119 = n1976 & ~n2108 ;
  assign n2120 = ~n2118 & n2119 ;
  assign n2121 = ~n2107 & ~n2120 ;
  assign n2122 = \TM0_pad  & \_2139__reg/NET0131  ;
  assign n2123 = \WX3361_reg/NET0131  & ~\WX3425_reg/NET0131  ;
  assign n2124 = ~\WX3361_reg/NET0131  & \WX3425_reg/NET0131  ;
  assign n2125 = ~n2123 & ~n2124 ;
  assign n2126 = \WX3297_reg/NET0131  & ~n2125 ;
  assign n2127 = ~\WX3297_reg/NET0131  & n2125 ;
  assign n2128 = ~n2126 & ~n2127 ;
  assign n2129 = \TM1_pad  & ~\WX3233_reg/NET0131  ;
  assign n2130 = ~\TM1_pad  & \WX3233_reg/NET0131  ;
  assign n2131 = ~n2129 & ~n2130 ;
  assign n2133 = n2128 & ~n2131 ;
  assign n2132 = ~n2128 & n2131 ;
  assign n2134 = ~\TM0_pad  & ~n2132 ;
  assign n2135 = ~n2133 & n2134 ;
  assign n2136 = ~n2122 & ~n2135 ;
  assign n2137 = n1976 & ~n2136 ;
  assign n2138 = ~n1855 & ~n2073 ;
  assign n2139 = n1973 & ~n2138 ;
  assign n2140 = ~n2137 & ~n2139 ;
  assign n2141 = \TM0_pad  & \_2288__reg/NET0131  ;
  assign n2142 = \WX9848_reg/NET0131  & ~\WX9912_reg/NET0131  ;
  assign n2143 = ~\WX9848_reg/NET0131  & \WX9912_reg/NET0131  ;
  assign n2144 = ~n2142 & ~n2143 ;
  assign n2145 = \WX9784_reg/NET0131  & ~n2144 ;
  assign n2146 = ~\WX9784_reg/NET0131  & n2144 ;
  assign n2147 = ~n2145 & ~n2146 ;
  assign n2148 = \TM1_pad  & ~\WX9720_reg/NET0131  ;
  assign n2149 = ~\TM1_pad  & \WX9720_reg/NET0131  ;
  assign n2150 = ~n2148 & ~n2149 ;
  assign n2152 = n2147 & ~n2150 ;
  assign n2151 = ~n2147 & n2150 ;
  assign n2153 = ~\TM0_pad  & ~n2151 ;
  assign n2154 = ~n2152 & n2153 ;
  assign n2155 = ~n2141 & ~n2154 ;
  assign n2156 = n1976 & ~n2155 ;
  assign n2157 = \WX8555_reg/NET0131  & ~\WX8619_reg/NET0131  ;
  assign n2158 = ~\WX8555_reg/NET0131  & \WX8619_reg/NET0131  ;
  assign n2159 = ~n2157 & ~n2158 ;
  assign n2160 = \WX8491_reg/NET0131  & ~n2159 ;
  assign n2161 = ~\WX8491_reg/NET0131  & n2159 ;
  assign n2162 = ~n2160 & ~n2161 ;
  assign n2163 = \TM1_pad  & ~\WX8427_reg/NET0131  ;
  assign n2164 = ~\TM1_pad  & \WX8427_reg/NET0131  ;
  assign n2165 = ~n2163 & ~n2164 ;
  assign n2167 = n2162 & ~n2165 ;
  assign n2166 = ~n2162 & n2165 ;
  assign n2168 = ~\TM0_pad  & ~n2166 ;
  assign n2169 = ~n2167 & n2168 ;
  assign n2170 = ~n1653 & ~n2169 ;
  assign n2171 = n1973 & ~n2170 ;
  assign n2172 = ~n2156 & ~n2171 ;
  assign n2173 = \TM0_pad  & \_2321__reg/NET0131  ;
  assign n2174 = \WX11139_reg/NET0131  & ~\WX11203_reg/NET0131  ;
  assign n2175 = ~\WX11139_reg/NET0131  & \WX11203_reg/NET0131  ;
  assign n2176 = ~n2174 & ~n2175 ;
  assign n2177 = \WX11075_reg/NET0131  & ~n2176 ;
  assign n2178 = ~\WX11075_reg/NET0131  & n2176 ;
  assign n2179 = ~n2177 & ~n2178 ;
  assign n2180 = \TM1_pad  & ~\WX11011_reg/NET0131  ;
  assign n2181 = ~\TM1_pad  & \WX11011_reg/NET0131  ;
  assign n2182 = ~n2180 & ~n2181 ;
  assign n2184 = n2179 & ~n2182 ;
  assign n2183 = ~n2179 & n2182 ;
  assign n2185 = ~\TM0_pad  & ~n2183 ;
  assign n2186 = ~n2184 & n2185 ;
  assign n2187 = ~n2173 & ~n2186 ;
  assign n2188 = n1976 & ~n2187 ;
  assign n2189 = \WX9846_reg/NET0131  & ~\WX9910_reg/NET0131  ;
  assign n2190 = ~\WX9846_reg/NET0131  & \WX9910_reg/NET0131  ;
  assign n2191 = ~n2189 & ~n2190 ;
  assign n2192 = \WX9782_reg/NET0131  & ~n2191 ;
  assign n2193 = ~\WX9782_reg/NET0131  & n2191 ;
  assign n2194 = ~n2192 & ~n2193 ;
  assign n2195 = \TM1_pad  & ~\WX9718_reg/NET0131  ;
  assign n2196 = ~\TM1_pad  & \WX9718_reg/NET0131  ;
  assign n2197 = ~n2195 & ~n2196 ;
  assign n2199 = n2194 & ~n2197 ;
  assign n2198 = ~n2194 & n2197 ;
  assign n2200 = ~\TM0_pad  & ~n2198 ;
  assign n2201 = ~n2199 & n2200 ;
  assign n2202 = ~n1682 & ~n2201 ;
  assign n2203 = n1973 & ~n2202 ;
  assign n2204 = ~n2188 & ~n2203 ;
  assign n2205 = \TM0_pad  & \_2189__reg/NET0131  ;
  assign n2206 = \WX5975_reg/NET0131  & ~\WX6039_reg/NET0131  ;
  assign n2207 = ~\WX5975_reg/NET0131  & \WX6039_reg/NET0131  ;
  assign n2208 = ~n2206 & ~n2207 ;
  assign n2209 = \WX5911_reg/NET0131  & ~n2208 ;
  assign n2210 = ~\WX5911_reg/NET0131  & n2208 ;
  assign n2211 = ~n2209 & ~n2210 ;
  assign n2212 = \TM1_pad  & ~\WX5847_reg/NET0131  ;
  assign n2213 = ~\TM1_pad  & \WX5847_reg/NET0131  ;
  assign n2214 = ~n2212 & ~n2213 ;
  assign n2216 = n2211 & ~n2214 ;
  assign n2215 = ~n2211 & n2214 ;
  assign n2217 = ~\TM0_pad  & ~n2215 ;
  assign n2218 = ~n2216 & n2217 ;
  assign n2219 = ~n2205 & ~n2218 ;
  assign n2220 = n1976 & ~n2219 ;
  assign n2221 = \WX4682_reg/NET0131  & ~\WX4746_reg/NET0131  ;
  assign n2222 = ~\WX4682_reg/NET0131  & \WX4746_reg/NET0131  ;
  assign n2223 = ~n2221 & ~n2222 ;
  assign n2224 = \WX4618_reg/NET0131  & ~n2223 ;
  assign n2225 = ~\WX4618_reg/NET0131  & n2223 ;
  assign n2226 = ~n2224 & ~n2225 ;
  assign n2227 = \TM1_pad  & ~\WX4554_reg/NET0131  ;
  assign n2228 = ~\TM1_pad  & \WX4554_reg/NET0131  ;
  assign n2229 = ~n2227 & ~n2228 ;
  assign n2231 = n2226 & ~n2229 ;
  assign n2230 = ~n2226 & n2229 ;
  assign n2232 = ~\TM0_pad  & ~n2230 ;
  assign n2233 = ~n2231 & n2232 ;
  assign n2234 = ~n1605 & ~n2233 ;
  assign n2235 = n1973 & ~n2234 ;
  assign n2236 = ~n2220 & ~n2235 ;
  assign n2237 = \TM0_pad  & \_2222__reg/NET0131  ;
  assign n2238 = \WX7266_reg/NET0131  & ~\WX7330_reg/NET0131  ;
  assign n2239 = ~\WX7266_reg/NET0131  & \WX7330_reg/NET0131  ;
  assign n2240 = ~n2238 & ~n2239 ;
  assign n2241 = \WX7202_reg/NET0131  & ~n2240 ;
  assign n2242 = ~\WX7202_reg/NET0131  & n2240 ;
  assign n2243 = ~n2241 & ~n2242 ;
  assign n2244 = \TM1_pad  & ~\WX7138_reg/NET0131  ;
  assign n2245 = ~\TM1_pad  & \WX7138_reg/NET0131  ;
  assign n2246 = ~n2244 & ~n2245 ;
  assign n2248 = n2243 & ~n2246 ;
  assign n2247 = ~n2243 & n2246 ;
  assign n2249 = ~\TM0_pad  & ~n2247 ;
  assign n2250 = ~n2248 & n2249 ;
  assign n2251 = ~n2237 & ~n2250 ;
  assign n2252 = n1976 & ~n2251 ;
  assign n2253 = \WX5973_reg/NET0131  & ~\WX6037_reg/NET0131  ;
  assign n2254 = ~\WX5973_reg/NET0131  & \WX6037_reg/NET0131  ;
  assign n2255 = ~n2253 & ~n2254 ;
  assign n2256 = \WX5909_reg/NET0131  & ~n2255 ;
  assign n2257 = ~\WX5909_reg/NET0131  & n2255 ;
  assign n2258 = ~n2256 & ~n2257 ;
  assign n2259 = \TM1_pad  & ~\WX5845_reg/NET0131  ;
  assign n2260 = ~\TM1_pad  & \WX5845_reg/NET0131  ;
  assign n2261 = ~n2259 & ~n2260 ;
  assign n2263 = n2258 & ~n2261 ;
  assign n2262 = ~n2258 & n2261 ;
  assign n2264 = ~\TM0_pad  & ~n2262 ;
  assign n2265 = ~n2263 & n2264 ;
  assign n2266 = ~n1621 & ~n2265 ;
  assign n2267 = n1973 & ~n2266 ;
  assign n2268 = ~n2252 & ~n2267 ;
  assign n2269 = \TM0_pad  & \_2255__reg/NET0131  ;
  assign n2270 = \WX8557_reg/NET0131  & ~\WX8621_reg/NET0131  ;
  assign n2271 = ~\WX8557_reg/NET0131  & \WX8621_reg/NET0131  ;
  assign n2272 = ~n2270 & ~n2271 ;
  assign n2273 = \WX8493_reg/NET0131  & ~n2272 ;
  assign n2274 = ~\WX8493_reg/NET0131  & n2272 ;
  assign n2275 = ~n2273 & ~n2274 ;
  assign n2276 = \TM1_pad  & ~\WX8429_reg/NET0131  ;
  assign n2277 = ~\TM1_pad  & \WX8429_reg/NET0131  ;
  assign n2278 = ~n2276 & ~n2277 ;
  assign n2280 = n2275 & ~n2278 ;
  assign n2279 = ~n2275 & n2278 ;
  assign n2281 = ~\TM0_pad  & ~n2279 ;
  assign n2282 = ~n2280 & n2281 ;
  assign n2283 = ~n2269 & ~n2282 ;
  assign n2284 = n1976 & ~n2283 ;
  assign n2285 = \WX7264_reg/NET0131  & ~\WX7328_reg/NET0131  ;
  assign n2286 = ~\WX7264_reg/NET0131  & \WX7328_reg/NET0131  ;
  assign n2287 = ~n2285 & ~n2286 ;
  assign n2288 = \WX7200_reg/NET0131  & ~n2287 ;
  assign n2289 = ~\WX7200_reg/NET0131  & n2287 ;
  assign n2290 = ~n2288 & ~n2289 ;
  assign n2291 = \TM1_pad  & ~\WX7136_reg/NET0131  ;
  assign n2292 = ~\TM1_pad  & \WX7136_reg/NET0131  ;
  assign n2293 = ~n2291 & ~n2292 ;
  assign n2295 = n2290 & ~n2293 ;
  assign n2294 = ~n2290 & n2293 ;
  assign n2296 = ~\TM0_pad  & ~n2294 ;
  assign n2297 = ~n2295 & n2296 ;
  assign n2298 = ~n1637 & ~n2297 ;
  assign n2299 = n1973 & ~n2298 ;
  assign n2300 = ~n2284 & ~n2299 ;
  assign n2301 = ~\TM0_pad  & ~n1819 ;
  assign n2302 = ~n1810 & ~n2301 ;
  assign n2303 = n1973 & ~n2302 ;
  assign n2304 = \TM0_pad  & \_2105__reg/NET0131  ;
  assign n2305 = \WX2072_reg/NET0131  & ~\WX2136_reg/NET0131  ;
  assign n2306 = ~\WX2072_reg/NET0131  & \WX2136_reg/NET0131  ;
  assign n2307 = ~n2305 & ~n2306 ;
  assign n2308 = \WX2008_reg/NET0131  & ~n2307 ;
  assign n2309 = ~\WX2008_reg/NET0131  & n2307 ;
  assign n2310 = ~n2308 & ~n2309 ;
  assign n2311 = \TM1_pad  & ~\WX1944_reg/NET0131  ;
  assign n2312 = ~\TM1_pad  & \WX1944_reg/NET0131  ;
  assign n2313 = ~n2311 & ~n2312 ;
  assign n2315 = n2310 & ~n2313 ;
  assign n2314 = ~n2310 & n2313 ;
  assign n2316 = ~\TM0_pad  & ~n2314 ;
  assign n2317 = ~n2315 & n2316 ;
  assign n2318 = ~n2304 & ~n2317 ;
  assign n2319 = n1976 & ~n2318 ;
  assign n2320 = ~n2303 & ~n2319 ;
  assign n2321 = \WX11119_reg/NET0131  & ~\WX11183_reg/NET0131  ;
  assign n2322 = ~\WX11119_reg/NET0131  & \WX11183_reg/NET0131  ;
  assign n2323 = ~n2321 & ~n2322 ;
  assign n2324 = \WX11055_reg/NET0131  & ~n2323 ;
  assign n2325 = ~\WX11055_reg/NET0131  & n2323 ;
  assign n2326 = ~n2324 & ~n2325 ;
  assign n2327 = \TM1_pad  & ~\WX10991_reg/NET0131  ;
  assign n2328 = ~\TM1_pad  & \WX10991_reg/NET0131  ;
  assign n2329 = ~n2327 & ~n2328 ;
  assign n2331 = n2326 & ~n2329 ;
  assign n2330 = ~n2326 & n2329 ;
  assign n2332 = ~\TM0_pad  & ~n2330 ;
  assign n2333 = ~n2331 & n2332 ;
  assign n2334 = ~n1855 & ~n2333 ;
  assign n2335 = n1973 & ~n2334 ;
  assign n2337 = \TM0_pad  & ~\_2363__reg/NET0131  ;
  assign n2336 = ~\DATA_0_30_pad  & ~\TM0_pad  ;
  assign n2338 = n1976 & ~n2336 ;
  assign n2339 = ~n2337 & n2338 ;
  assign n2340 = ~n2335 & ~n2339 ;
  assign n2341 = ~n1573 & n1973 ;
  assign n2342 = \WX3393_reg/NET0131  & ~\WX3457_reg/NET0131  ;
  assign n2343 = ~\WX3393_reg/NET0131  & \WX3457_reg/NET0131  ;
  assign n2344 = ~n2342 & ~n2343 ;
  assign n2345 = \WX3265_reg/NET0131  & ~\WX3329_reg/NET0131  ;
  assign n2346 = ~\WX3265_reg/NET0131  & \WX3329_reg/NET0131  ;
  assign n2347 = ~n2345 & ~n2346 ;
  assign n2349 = n2344 & ~n2347 ;
  assign n2348 = ~n2344 & n2347 ;
  assign n2350 = ~\TM0_pad  & ~n2348 ;
  assign n2351 = ~n2349 & n2350 ;
  assign n2352 = n2341 & ~n2351 ;
  assign n2354 = \WX4686_reg/NET0131  & ~\WX4750_reg/NET0131  ;
  assign n2355 = ~\WX4686_reg/NET0131  & \WX4750_reg/NET0131  ;
  assign n2356 = ~n2354 & ~n2355 ;
  assign n2357 = \WX4558_reg/NET0131  & ~\WX4622_reg/NET0131  ;
  assign n2358 = ~\WX4558_reg/NET0131  & \WX4622_reg/NET0131  ;
  assign n2359 = ~n2357 & ~n2358 ;
  assign n2361 = n2356 & ~n2359 ;
  assign n2360 = ~n2356 & n2359 ;
  assign n2362 = ~\TM0_pad  & ~n2360 ;
  assign n2363 = ~n2361 & n2362 ;
  assign n2353 = \TM0_pad  & ~\_2155__reg/NET0131  ;
  assign n2364 = n1976 & ~n2353 ;
  assign n2365 = ~n2363 & n2364 ;
  assign n2366 = ~n2352 & ~n2365 ;
  assign n2367 = \TM0_pad  & \_2287__reg/NET0131  ;
  assign n2368 = \WX9850_reg/NET0131  & ~\WX9914_reg/NET0131  ;
  assign n2369 = ~\WX9850_reg/NET0131  & \WX9914_reg/NET0131  ;
  assign n2370 = ~n2368 & ~n2369 ;
  assign n2371 = \WX9786_reg/NET0131  & ~n2370 ;
  assign n2372 = ~\WX9786_reg/NET0131  & n2370 ;
  assign n2373 = ~n2371 & ~n2372 ;
  assign n2374 = \TM1_pad  & ~\WX9722_reg/NET0131  ;
  assign n2375 = ~\TM1_pad  & \WX9722_reg/NET0131  ;
  assign n2376 = ~n2374 & ~n2375 ;
  assign n2378 = n2373 & ~n2376 ;
  assign n2377 = ~n2373 & n2376 ;
  assign n2379 = ~\TM0_pad  & ~n2377 ;
  assign n2380 = ~n2378 & n2379 ;
  assign n2381 = ~n2367 & ~n2380 ;
  assign n2382 = n1976 & ~n2381 ;
  assign n2383 = ~n1637 & ~n2282 ;
  assign n2384 = n1973 & ~n2383 ;
  assign n2385 = ~n2382 & ~n2384 ;
  assign n2386 = \TM0_pad  & \_2138__reg/NET0131  ;
  assign n2387 = \WX3363_reg/NET0131  & ~\WX3427_reg/NET0131  ;
  assign n2388 = ~\WX3363_reg/NET0131  & \WX3427_reg/NET0131  ;
  assign n2389 = ~n2387 & ~n2388 ;
  assign n2390 = \WX3299_reg/NET0131  & ~n2389 ;
  assign n2391 = ~\WX3299_reg/NET0131  & n2389 ;
  assign n2392 = ~n2390 & ~n2391 ;
  assign n2393 = \TM1_pad  & ~\WX3235_reg/NET0131  ;
  assign n2394 = ~\TM1_pad  & \WX3235_reg/NET0131  ;
  assign n2395 = ~n2393 & ~n2394 ;
  assign n2397 = n2392 & ~n2395 ;
  assign n2396 = ~n2392 & n2395 ;
  assign n2398 = ~\TM0_pad  & ~n2396 ;
  assign n2399 = ~n2397 & n2398 ;
  assign n2400 = ~n2386 & ~n2399 ;
  assign n2401 = n1976 & ~n2400 ;
  assign n2402 = ~n1826 & ~n2093 ;
  assign n2403 = n1973 & ~n2402 ;
  assign n2404 = ~n2401 & ~n2403 ;
  assign n2405 = \TM0_pad  & \_2320__reg/NET0131  ;
  assign n2406 = \WX11141_reg/NET0131  & ~\WX11205_reg/NET0131  ;
  assign n2407 = ~\WX11141_reg/NET0131  & \WX11205_reg/NET0131  ;
  assign n2408 = ~n2406 & ~n2407 ;
  assign n2409 = \WX11077_reg/NET0131  & ~n2408 ;
  assign n2410 = ~\WX11077_reg/NET0131  & n2408 ;
  assign n2411 = ~n2409 & ~n2410 ;
  assign n2412 = \TM1_pad  & ~\WX11013_reg/NET0131  ;
  assign n2413 = ~\TM1_pad  & \WX11013_reg/NET0131  ;
  assign n2414 = ~n2412 & ~n2413 ;
  assign n2416 = n2411 & ~n2414 ;
  assign n2415 = ~n2411 & n2414 ;
  assign n2417 = ~\TM0_pad  & ~n2415 ;
  assign n2418 = ~n2416 & n2417 ;
  assign n2419 = ~n2405 & ~n2418 ;
  assign n2420 = n1976 & ~n2419 ;
  assign n2421 = ~n1653 & ~n2154 ;
  assign n2422 = n1973 & ~n2421 ;
  assign n2423 = ~n2420 & ~n2422 ;
  assign n2424 = n1974 & ~n2118 ;
  assign n2426 = \WX5977_reg/NET0131  & ~\WX6041_reg/NET0131  ;
  assign n2427 = ~\WX5977_reg/NET0131  & \WX6041_reg/NET0131  ;
  assign n2428 = ~n2426 & ~n2427 ;
  assign n2429 = \WX5849_reg/NET0131  & ~\WX5913_reg/NET0131  ;
  assign n2430 = ~\WX5849_reg/NET0131  & \WX5913_reg/NET0131  ;
  assign n2431 = ~n2429 & ~n2430 ;
  assign n2433 = n2428 & ~n2431 ;
  assign n2432 = ~n2428 & n2431 ;
  assign n2434 = ~\TM0_pad  & ~n2432 ;
  assign n2435 = ~n2433 & n2434 ;
  assign n2425 = \TM0_pad  & ~\_2188__reg/NET0131  ;
  assign n2436 = n1976 & ~n2425 ;
  assign n2437 = ~n2435 & n2436 ;
  assign n2438 = ~n2424 & ~n2437 ;
  assign n2439 = \TM0_pad  & \_2221__reg/NET0131  ;
  assign n2440 = \WX7268_reg/NET0131  & ~\WX7332_reg/NET0131  ;
  assign n2441 = ~\WX7268_reg/NET0131  & \WX7332_reg/NET0131  ;
  assign n2442 = ~n2440 & ~n2441 ;
  assign n2443 = \WX7204_reg/NET0131  & ~n2442 ;
  assign n2444 = ~\WX7204_reg/NET0131  & n2442 ;
  assign n2445 = ~n2443 & ~n2444 ;
  assign n2446 = \TM1_pad  & ~\WX7140_reg/NET0131  ;
  assign n2447 = ~\TM1_pad  & \WX7140_reg/NET0131  ;
  assign n2448 = ~n2446 & ~n2447 ;
  assign n2450 = n2445 & ~n2448 ;
  assign n2449 = ~n2445 & n2448 ;
  assign n2451 = ~\TM0_pad  & ~n2449 ;
  assign n2452 = ~n2450 & n2451 ;
  assign n2453 = ~n2439 & ~n2452 ;
  assign n2454 = n1976 & ~n2453 ;
  assign n2455 = ~n1605 & ~n2218 ;
  assign n2456 = n1973 & ~n2455 ;
  assign n2457 = ~n2454 & ~n2456 ;
  assign n2458 = \TM0_pad  & \_2254__reg/NET0131  ;
  assign n2459 = \WX8559_reg/NET0131  & ~\WX8623_reg/NET0131  ;
  assign n2460 = ~\WX8559_reg/NET0131  & \WX8623_reg/NET0131  ;
  assign n2461 = ~n2459 & ~n2460 ;
  assign n2462 = \WX8495_reg/NET0131  & ~n2461 ;
  assign n2463 = ~\WX8495_reg/NET0131  & n2461 ;
  assign n2464 = ~n2462 & ~n2463 ;
  assign n2465 = \TM1_pad  & ~\WX8431_reg/NET0131  ;
  assign n2466 = ~\TM1_pad  & \WX8431_reg/NET0131  ;
  assign n2467 = ~n2465 & ~n2466 ;
  assign n2469 = n2464 & ~n2467 ;
  assign n2468 = ~n2464 & n2467 ;
  assign n2470 = ~\TM0_pad  & ~n2468 ;
  assign n2471 = ~n2469 & n2470 ;
  assign n2472 = ~n2458 & ~n2471 ;
  assign n2473 = n1976 & ~n2472 ;
  assign n2474 = ~n1621 & ~n2250 ;
  assign n2475 = n1973 & ~n2474 ;
  assign n2476 = ~n2473 & ~n2475 ;
  assign n2477 = ~\TM0_pad  & ~n1803 ;
  assign n2478 = ~n1794 & ~n2477 ;
  assign n2479 = n1973 & ~n2478 ;
  assign n2480 = \TM0_pad  & \_2104__reg/NET0131  ;
  assign n2481 = \WX2074_reg/NET0131  & ~\WX2138_reg/NET0131  ;
  assign n2482 = ~\WX2074_reg/NET0131  & \WX2138_reg/NET0131  ;
  assign n2483 = ~n2481 & ~n2482 ;
  assign n2484 = \WX2010_reg/NET0131  & ~n2483 ;
  assign n2485 = ~\WX2010_reg/NET0131  & n2483 ;
  assign n2486 = ~n2484 & ~n2485 ;
  assign n2487 = \TM1_pad  & ~\WX1946_reg/NET0131  ;
  assign n2488 = ~\TM1_pad  & \WX1946_reg/NET0131  ;
  assign n2489 = ~n2487 & ~n2488 ;
  assign n2491 = n2486 & ~n2489 ;
  assign n2490 = ~n2486 & n2489 ;
  assign n2492 = ~\TM0_pad  & ~n2490 ;
  assign n2493 = ~n2491 & n2492 ;
  assign n2494 = ~n2480 & ~n2493 ;
  assign n2495 = n1976 & ~n2494 ;
  assign n2496 = ~n2479 & ~n2495 ;
  assign n2497 = \WX11121_reg/NET0131  & ~\WX11185_reg/NET0131  ;
  assign n2498 = ~\WX11121_reg/NET0131  & \WX11185_reg/NET0131  ;
  assign n2499 = ~n2497 & ~n2498 ;
  assign n2500 = \WX11057_reg/NET0131  & ~n2499 ;
  assign n2501 = ~\WX11057_reg/NET0131  & n2499 ;
  assign n2502 = ~n2500 & ~n2501 ;
  assign n2503 = \TM1_pad  & ~\WX10993_reg/NET0131  ;
  assign n2504 = ~\TM1_pad  & \WX10993_reg/NET0131  ;
  assign n2505 = ~n2503 & ~n2504 ;
  assign n2507 = n2502 & ~n2505 ;
  assign n2506 = ~n2502 & n2505 ;
  assign n2508 = ~\TM0_pad  & ~n2506 ;
  assign n2509 = ~n2507 & n2508 ;
  assign n2510 = ~n1826 & ~n2509 ;
  assign n2511 = n1973 & ~n2510 ;
  assign n2513 = \TM0_pad  & ~\_2362__reg/NET0131  ;
  assign n2512 = ~\DATA_0_29_pad  & ~\TM0_pad  ;
  assign n2514 = n1976 & ~n2512 ;
  assign n2515 = ~n2513 & n2514 ;
  assign n2516 = ~n2511 & ~n2515 ;
  assign n2517 = RESET_pad & \WX10831_reg/NET0131  ;
  assign n2518 = \WX3395_reg/NET0131  & ~\WX3459_reg/NET0131  ;
  assign n2519 = ~\WX3395_reg/NET0131  & \WX3459_reg/NET0131  ;
  assign n2520 = ~n2518 & ~n2519 ;
  assign n2521 = \WX3267_reg/NET0131  & ~\WX3331_reg/NET0131  ;
  assign n2522 = ~\WX3267_reg/NET0131  & \WX3331_reg/NET0131  ;
  assign n2523 = ~n2521 & ~n2522 ;
  assign n2525 = n2520 & ~n2523 ;
  assign n2524 = ~n2520 & n2523 ;
  assign n2526 = ~\TM0_pad  & ~n2524 ;
  assign n2527 = ~n2525 & n2526 ;
  assign n2528 = n2040 & ~n2527 ;
  assign n2530 = \WX4688_reg/NET0131  & ~\WX4752_reg/NET0131  ;
  assign n2531 = ~\WX4688_reg/NET0131  & \WX4752_reg/NET0131  ;
  assign n2532 = ~n2530 & ~n2531 ;
  assign n2533 = \WX4560_reg/NET0131  & ~\WX4624_reg/NET0131  ;
  assign n2534 = ~\WX4560_reg/NET0131  & \WX4624_reg/NET0131  ;
  assign n2535 = ~n2533 & ~n2534 ;
  assign n2537 = n2532 & ~n2535 ;
  assign n2536 = ~n2532 & n2535 ;
  assign n2538 = ~\TM0_pad  & ~n2536 ;
  assign n2539 = ~n2537 & n2538 ;
  assign n2529 = \TM0_pad  & ~\_2154__reg/NET0131  ;
  assign n2540 = n1976 & ~n2529 ;
  assign n2541 = ~n2539 & n2540 ;
  assign n2542 = ~n2528 & ~n2541 ;
  assign n2543 = \TM0_pad  & \_2286__reg/NET0131  ;
  assign n2544 = \WX9852_reg/NET0131  & ~\WX9916_reg/NET0131  ;
  assign n2545 = ~\WX9852_reg/NET0131  & \WX9916_reg/NET0131  ;
  assign n2546 = ~n2544 & ~n2545 ;
  assign n2547 = \WX9788_reg/NET0131  & ~n2546 ;
  assign n2548 = ~\WX9788_reg/NET0131  & n2546 ;
  assign n2549 = ~n2547 & ~n2548 ;
  assign n2550 = \TM1_pad  & ~\WX9724_reg/NET0131  ;
  assign n2551 = ~\TM1_pad  & \WX9724_reg/NET0131  ;
  assign n2552 = ~n2550 & ~n2551 ;
  assign n2554 = n2549 & ~n2552 ;
  assign n2553 = ~n2549 & n2552 ;
  assign n2555 = ~\TM0_pad  & ~n2553 ;
  assign n2556 = ~n2554 & n2555 ;
  assign n2557 = ~n2543 & ~n2556 ;
  assign n2558 = n1976 & ~n2557 ;
  assign n2559 = ~n1621 & ~n2471 ;
  assign n2560 = n1973 & ~n2559 ;
  assign n2561 = ~n2558 & ~n2560 ;
  assign n2562 = \TM0_pad  & \_2137__reg/NET0131  ;
  assign n2563 = \WX3365_reg/NET0131  & ~\WX3429_reg/NET0131  ;
  assign n2564 = ~\WX3365_reg/NET0131  & \WX3429_reg/NET0131  ;
  assign n2565 = ~n2563 & ~n2564 ;
  assign n2566 = \WX3301_reg/NET0131  & ~n2565 ;
  assign n2567 = ~\WX3301_reg/NET0131  & n2565 ;
  assign n2568 = ~n2566 & ~n2567 ;
  assign n2569 = \TM1_pad  & ~\WX3237_reg/NET0131  ;
  assign n2570 = ~\TM1_pad  & \WX3237_reg/NET0131  ;
  assign n2571 = ~n2569 & ~n2570 ;
  assign n2573 = n2568 & ~n2571 ;
  assign n2572 = ~n2568 & n2571 ;
  assign n2574 = ~\TM0_pad  & ~n2572 ;
  assign n2575 = ~n2573 & n2574 ;
  assign n2576 = ~n2562 & ~n2575 ;
  assign n2577 = n1976 & ~n2576 ;
  assign n2578 = ~n1810 & ~n2317 ;
  assign n2579 = n1973 & ~n2578 ;
  assign n2580 = ~n2577 & ~n2579 ;
  assign n2581 = \TM0_pad  & \_2319__reg/NET0131  ;
  assign n2582 = \WX11143_reg/NET0131  & ~\WX11207_reg/NET0131  ;
  assign n2583 = ~\WX11143_reg/NET0131  & \WX11207_reg/NET0131  ;
  assign n2584 = ~n2582 & ~n2583 ;
  assign n2585 = \WX11079_reg/NET0131  & ~n2584 ;
  assign n2586 = ~\WX11079_reg/NET0131  & n2584 ;
  assign n2587 = ~n2585 & ~n2586 ;
  assign n2588 = \TM1_pad  & ~\WX11015_reg/NET0131  ;
  assign n2589 = ~\TM1_pad  & \WX11015_reg/NET0131  ;
  assign n2590 = ~n2588 & ~n2589 ;
  assign n2592 = n2587 & ~n2590 ;
  assign n2591 = ~n2587 & n2590 ;
  assign n2593 = ~\TM0_pad  & ~n2591 ;
  assign n2594 = ~n2592 & n2593 ;
  assign n2595 = ~n2581 & ~n2594 ;
  assign n2596 = n1976 & ~n2595 ;
  assign n2597 = ~n1637 & ~n2380 ;
  assign n2598 = n1973 & ~n2597 ;
  assign n2599 = ~n2596 & ~n2598 ;
  assign n2600 = n2341 & ~n2363 ;
  assign n2602 = \WX5979_reg/NET0131  & ~\WX6043_reg/NET0131  ;
  assign n2603 = ~\WX5979_reg/NET0131  & \WX6043_reg/NET0131  ;
  assign n2604 = ~n2602 & ~n2603 ;
  assign n2605 = \WX5851_reg/NET0131  & ~\WX5915_reg/NET0131  ;
  assign n2606 = ~\WX5851_reg/NET0131  & \WX5915_reg/NET0131  ;
  assign n2607 = ~n2605 & ~n2606 ;
  assign n2609 = n2604 & ~n2607 ;
  assign n2608 = ~n2604 & n2607 ;
  assign n2610 = ~\TM0_pad  & ~n2608 ;
  assign n2611 = ~n2609 & n2610 ;
  assign n2601 = \TM0_pad  & ~\_2187__reg/NET0131  ;
  assign n2612 = n1976 & ~n2601 ;
  assign n2613 = ~n2611 & n2612 ;
  assign n2614 = ~n2600 & ~n2613 ;
  assign n2615 = n1974 & ~n2435 ;
  assign n2617 = \WX7270_reg/NET0131  & ~\WX7334_reg/NET0131  ;
  assign n2618 = ~\WX7270_reg/NET0131  & \WX7334_reg/NET0131  ;
  assign n2619 = ~n2617 & ~n2618 ;
  assign n2620 = \WX7142_reg/NET0131  & ~\WX7206_reg/NET0131  ;
  assign n2621 = ~\WX7142_reg/NET0131  & \WX7206_reg/NET0131  ;
  assign n2622 = ~n2620 & ~n2621 ;
  assign n2624 = n2619 & ~n2622 ;
  assign n2623 = ~n2619 & n2622 ;
  assign n2625 = ~\TM0_pad  & ~n2623 ;
  assign n2626 = ~n2624 & n2625 ;
  assign n2616 = \TM0_pad  & ~\_2220__reg/NET0131  ;
  assign n2627 = n1976 & ~n2616 ;
  assign n2628 = ~n2626 & n2627 ;
  assign n2629 = ~n2615 & ~n2628 ;
  assign n2630 = \TM0_pad  & \_2253__reg/NET0131  ;
  assign n2631 = \WX8561_reg/NET0131  & ~\WX8625_reg/NET0131  ;
  assign n2632 = ~\WX8561_reg/NET0131  & \WX8625_reg/NET0131  ;
  assign n2633 = ~n2631 & ~n2632 ;
  assign n2634 = \WX8497_reg/NET0131  & ~n2633 ;
  assign n2635 = ~\WX8497_reg/NET0131  & n2633 ;
  assign n2636 = ~n2634 & ~n2635 ;
  assign n2637 = \TM1_pad  & ~\WX8433_reg/NET0131  ;
  assign n2638 = ~\TM1_pad  & \WX8433_reg/NET0131  ;
  assign n2639 = ~n2637 & ~n2638 ;
  assign n2641 = n2636 & ~n2639 ;
  assign n2640 = ~n2636 & n2639 ;
  assign n2642 = ~\TM0_pad  & ~n2640 ;
  assign n2643 = ~n2641 & n2642 ;
  assign n2644 = ~n2630 & ~n2643 ;
  assign n2645 = n1976 & ~n2644 ;
  assign n2646 = ~n1605 & ~n2452 ;
  assign n2647 = n1973 & ~n2646 ;
  assign n2648 = ~n2645 & ~n2647 ;
  assign n2649 = ~\TM0_pad  & ~n1787 ;
  assign n2650 = ~n1778 & ~n2649 ;
  assign n2651 = n1973 & ~n2650 ;
  assign n2652 = \TM0_pad  & \_2103__reg/NET0131  ;
  assign n2653 = \WX2076_reg/NET0131  & ~\WX2140_reg/NET0131  ;
  assign n2654 = ~\WX2076_reg/NET0131  & \WX2140_reg/NET0131  ;
  assign n2655 = ~n2653 & ~n2654 ;
  assign n2656 = \WX2012_reg/NET0131  & ~n2655 ;
  assign n2657 = ~\WX2012_reg/NET0131  & n2655 ;
  assign n2658 = ~n2656 & ~n2657 ;
  assign n2659 = \TM1_pad  & ~\WX1948_reg/NET0131  ;
  assign n2660 = ~\TM1_pad  & \WX1948_reg/NET0131  ;
  assign n2661 = ~n2659 & ~n2660 ;
  assign n2663 = n2658 & ~n2661 ;
  assign n2662 = ~n2658 & n2661 ;
  assign n2664 = ~\TM0_pad  & ~n2662 ;
  assign n2665 = ~n2663 & n2664 ;
  assign n2666 = ~n2652 & ~n2665 ;
  assign n2667 = n1976 & ~n2666 ;
  assign n2668 = ~n2651 & ~n2667 ;
  assign n2669 = ~n1810 & ~n2019 ;
  assign n2670 = n1973 & ~n2669 ;
  assign n2672 = \TM0_pad  & ~\_2361__reg/NET0131  ;
  assign n2671 = ~\DATA_0_28_pad  & ~\TM0_pad  ;
  assign n2673 = n1976 & ~n2671 ;
  assign n2674 = ~n2672 & n2673 ;
  assign n2675 = ~n2670 & ~n2674 ;
  assign n2676 = RESET_pad & \WX10833_reg/NET0131  ;
  assign n2677 = ~n1547 & n1973 ;
  assign n2678 = \WX3397_reg/NET0131  & ~\WX3461_reg/NET0131  ;
  assign n2679 = ~\WX3397_reg/NET0131  & \WX3461_reg/NET0131  ;
  assign n2680 = ~n2678 & ~n2679 ;
  assign n2681 = \WX3269_reg/NET0131  & ~\WX3333_reg/NET0131  ;
  assign n2682 = ~\WX3269_reg/NET0131  & \WX3333_reg/NET0131  ;
  assign n2683 = ~n2681 & ~n2682 ;
  assign n2685 = n2680 & ~n2683 ;
  assign n2684 = ~n2680 & n2683 ;
  assign n2686 = ~\TM0_pad  & ~n2684 ;
  assign n2687 = ~n2685 & n2686 ;
  assign n2688 = n2677 & ~n2687 ;
  assign n2690 = \WX4690_reg/NET0131  & ~\WX4754_reg/NET0131  ;
  assign n2691 = ~\WX4690_reg/NET0131  & \WX4754_reg/NET0131  ;
  assign n2692 = ~n2690 & ~n2691 ;
  assign n2693 = \WX4562_reg/NET0131  & ~\WX4626_reg/NET0131  ;
  assign n2694 = ~\WX4562_reg/NET0131  & \WX4626_reg/NET0131  ;
  assign n2695 = ~n2693 & ~n2694 ;
  assign n2697 = n2692 & ~n2695 ;
  assign n2696 = ~n2692 & n2695 ;
  assign n2698 = ~\TM0_pad  & ~n2696 ;
  assign n2699 = ~n2697 & n2698 ;
  assign n2689 = \TM0_pad  & ~\_2153__reg/NET0131  ;
  assign n2700 = n1976 & ~n2689 ;
  assign n2701 = ~n2699 & n2700 ;
  assign n2702 = ~n2688 & ~n2701 ;
  assign n2703 = \TM0_pad  & \_2285__reg/NET0131  ;
  assign n2704 = \WX9854_reg/NET0131  & ~\WX9918_reg/NET0131  ;
  assign n2705 = ~\WX9854_reg/NET0131  & \WX9918_reg/NET0131  ;
  assign n2706 = ~n2704 & ~n2705 ;
  assign n2707 = \WX9790_reg/NET0131  & ~n2706 ;
  assign n2708 = ~\WX9790_reg/NET0131  & n2706 ;
  assign n2709 = ~n2707 & ~n2708 ;
  assign n2710 = \TM1_pad  & ~\WX9726_reg/NET0131  ;
  assign n2711 = ~\TM1_pad  & \WX9726_reg/NET0131  ;
  assign n2712 = ~n2710 & ~n2711 ;
  assign n2714 = n2709 & ~n2712 ;
  assign n2713 = ~n2709 & n2712 ;
  assign n2715 = ~\TM0_pad  & ~n2713 ;
  assign n2716 = ~n2714 & n2715 ;
  assign n2717 = ~n2703 & ~n2716 ;
  assign n2718 = n1976 & ~n2717 ;
  assign n2719 = ~n1605 & ~n2643 ;
  assign n2720 = n1973 & ~n2719 ;
  assign n2721 = ~n2718 & ~n2720 ;
  assign n2722 = \TM0_pad  & \_2136__reg/NET0131  ;
  assign n2723 = \WX3367_reg/NET0131  & ~\WX3431_reg/NET0131  ;
  assign n2724 = ~\WX3367_reg/NET0131  & \WX3431_reg/NET0131  ;
  assign n2725 = ~n2723 & ~n2724 ;
  assign n2726 = \WX3303_reg/NET0131  & ~n2725 ;
  assign n2727 = ~\WX3303_reg/NET0131  & n2725 ;
  assign n2728 = ~n2726 & ~n2727 ;
  assign n2729 = \TM1_pad  & ~\WX3239_reg/NET0131  ;
  assign n2730 = ~\TM1_pad  & \WX3239_reg/NET0131  ;
  assign n2731 = ~n2729 & ~n2730 ;
  assign n2733 = n2728 & ~n2731 ;
  assign n2732 = ~n2728 & n2731 ;
  assign n2734 = ~\TM0_pad  & ~n2732 ;
  assign n2735 = ~n2733 & n2734 ;
  assign n2736 = ~n2722 & ~n2735 ;
  assign n2737 = n1976 & ~n2736 ;
  assign n2738 = ~n1794 & ~n2493 ;
  assign n2739 = n1973 & ~n2738 ;
  assign n2740 = ~n2737 & ~n2739 ;
  assign n2741 = \TM0_pad  & \_2318__reg/NET0131  ;
  assign n2742 = \WX11145_reg/NET0131  & ~\WX11209_reg/NET0131  ;
  assign n2743 = ~\WX11145_reg/NET0131  & \WX11209_reg/NET0131  ;
  assign n2744 = ~n2742 & ~n2743 ;
  assign n2745 = \WX11081_reg/NET0131  & ~n2744 ;
  assign n2746 = ~\WX11081_reg/NET0131  & n2744 ;
  assign n2747 = ~n2745 & ~n2746 ;
  assign n2748 = \TM1_pad  & ~\WX11017_reg/NET0131  ;
  assign n2749 = ~\TM1_pad  & \WX11017_reg/NET0131  ;
  assign n2750 = ~n2748 & ~n2749 ;
  assign n2752 = n2747 & ~n2750 ;
  assign n2751 = ~n2747 & n2750 ;
  assign n2753 = ~\TM0_pad  & ~n2751 ;
  assign n2754 = ~n2752 & n2753 ;
  assign n2755 = ~n2741 & ~n2754 ;
  assign n2756 = n1976 & ~n2755 ;
  assign n2757 = ~n1621 & ~n2556 ;
  assign n2758 = n1973 & ~n2757 ;
  assign n2759 = ~n2756 & ~n2758 ;
  assign n2760 = n2040 & ~n2539 ;
  assign n2762 = \WX5981_reg/NET0131  & ~\WX6045_reg/NET0131  ;
  assign n2763 = ~\WX5981_reg/NET0131  & \WX6045_reg/NET0131  ;
  assign n2764 = ~n2762 & ~n2763 ;
  assign n2765 = \WX5853_reg/NET0131  & ~\WX5917_reg/NET0131  ;
  assign n2766 = ~\WX5853_reg/NET0131  & \WX5917_reg/NET0131  ;
  assign n2767 = ~n2765 & ~n2766 ;
  assign n2769 = n2764 & ~n2767 ;
  assign n2768 = ~n2764 & n2767 ;
  assign n2770 = ~\TM0_pad  & ~n2768 ;
  assign n2771 = ~n2769 & n2770 ;
  assign n2761 = \TM0_pad  & ~\_2186__reg/NET0131  ;
  assign n2772 = n1976 & ~n2761 ;
  assign n2773 = ~n2771 & n2772 ;
  assign n2774 = ~n2760 & ~n2773 ;
  assign n2775 = n2341 & ~n2611 ;
  assign n2777 = \WX7272_reg/NET0131  & ~\WX7336_reg/NET0131  ;
  assign n2778 = ~\WX7272_reg/NET0131  & \WX7336_reg/NET0131  ;
  assign n2779 = ~n2777 & ~n2778 ;
  assign n2780 = \WX7144_reg/NET0131  & ~\WX7208_reg/NET0131  ;
  assign n2781 = ~\WX7144_reg/NET0131  & \WX7208_reg/NET0131  ;
  assign n2782 = ~n2780 & ~n2781 ;
  assign n2784 = n2779 & ~n2782 ;
  assign n2783 = ~n2779 & n2782 ;
  assign n2785 = ~\TM0_pad  & ~n2783 ;
  assign n2786 = ~n2784 & n2785 ;
  assign n2776 = \TM0_pad  & ~\_2219__reg/NET0131  ;
  assign n2787 = n1976 & ~n2776 ;
  assign n2788 = ~n2786 & n2787 ;
  assign n2789 = ~n2775 & ~n2788 ;
  assign n2790 = n1974 & ~n2626 ;
  assign n2792 = \WX8563_reg/NET0131  & ~\WX8627_reg/NET0131  ;
  assign n2793 = ~\WX8563_reg/NET0131  & \WX8627_reg/NET0131  ;
  assign n2794 = ~n2792 & ~n2793 ;
  assign n2795 = \WX8435_reg/NET0131  & ~\WX8499_reg/NET0131  ;
  assign n2796 = ~\WX8435_reg/NET0131  & \WX8499_reg/NET0131  ;
  assign n2797 = ~n2795 & ~n2796 ;
  assign n2799 = n2794 & ~n2797 ;
  assign n2798 = ~n2794 & n2797 ;
  assign n2800 = ~\TM0_pad  & ~n2798 ;
  assign n2801 = ~n2799 & n2800 ;
  assign n2791 = \TM0_pad  & ~\_2252__reg/NET0131  ;
  assign n2802 = n1976 & ~n2791 ;
  assign n2803 = ~n2801 & n2802 ;
  assign n2804 = ~n2790 & ~n2803 ;
  assign n2805 = ~\TM0_pad  & ~n1771 ;
  assign n2806 = ~n1762 & ~n2805 ;
  assign n2807 = n1973 & ~n2806 ;
  assign n2808 = \TM0_pad  & \_2102__reg/NET0131  ;
  assign n2809 = \WX2078_reg/NET0131  & ~\WX2142_reg/NET0131  ;
  assign n2810 = ~\WX2078_reg/NET0131  & \WX2142_reg/NET0131  ;
  assign n2811 = ~n2809 & ~n2810 ;
  assign n2812 = \WX2014_reg/NET0131  & ~n2811 ;
  assign n2813 = ~\WX2014_reg/NET0131  & n2811 ;
  assign n2814 = ~n2812 & ~n2813 ;
  assign n2815 = \TM1_pad  & ~\WX1950_reg/NET0131  ;
  assign n2816 = ~\TM1_pad  & \WX1950_reg/NET0131  ;
  assign n2817 = ~n2815 & ~n2816 ;
  assign n2819 = n2814 & ~n2817 ;
  assign n2818 = ~n2814 & n2817 ;
  assign n2820 = ~\TM0_pad  & ~n2818 ;
  assign n2821 = ~n2819 & n2820 ;
  assign n2822 = ~n2808 & ~n2821 ;
  assign n2823 = n1976 & ~n2822 ;
  assign n2824 = ~n2807 & ~n2823 ;
  assign n2825 = \WX11125_reg/NET0131  & ~\WX11189_reg/NET0131  ;
  assign n2826 = ~\WX11125_reg/NET0131  & \WX11189_reg/NET0131  ;
  assign n2827 = ~n2825 & ~n2826 ;
  assign n2828 = \WX11061_reg/NET0131  & ~n2827 ;
  assign n2829 = ~\WX11061_reg/NET0131  & n2827 ;
  assign n2830 = ~n2828 & ~n2829 ;
  assign n2831 = \TM1_pad  & ~\WX10997_reg/NET0131  ;
  assign n2832 = ~\TM1_pad  & \WX10997_reg/NET0131  ;
  assign n2833 = ~n2831 & ~n2832 ;
  assign n2835 = n2830 & ~n2833 ;
  assign n2834 = ~n2830 & n2833 ;
  assign n2836 = ~\TM0_pad  & ~n2834 ;
  assign n2837 = ~n2835 & n2836 ;
  assign n2838 = ~n1794 & ~n2837 ;
  assign n2839 = n1973 & ~n2838 ;
  assign n2841 = \TM0_pad  & ~\_2360__reg/NET0131  ;
  assign n2840 = ~\DATA_0_27_pad  & ~\TM0_pad  ;
  assign n2842 = n1976 & ~n2840 ;
  assign n2843 = ~n2841 & n2842 ;
  assign n2844 = ~n2839 & ~n2843 ;
  assign n2845 = RESET_pad & \WX10835_reg/NET0131  ;
  assign n2846 = ~n1534 & n1973 ;
  assign n2847 = \WX3399_reg/NET0131  & ~\WX3463_reg/NET0131  ;
  assign n2848 = ~\WX3399_reg/NET0131  & \WX3463_reg/NET0131  ;
  assign n2849 = ~n2847 & ~n2848 ;
  assign n2850 = \WX3271_reg/NET0131  & ~\WX3335_reg/NET0131  ;
  assign n2851 = ~\WX3271_reg/NET0131  & \WX3335_reg/NET0131  ;
  assign n2852 = ~n2850 & ~n2851 ;
  assign n2854 = n2849 & ~n2852 ;
  assign n2853 = ~n2849 & n2852 ;
  assign n2855 = ~\TM0_pad  & ~n2853 ;
  assign n2856 = ~n2854 & n2855 ;
  assign n2857 = n2846 & ~n2856 ;
  assign n2859 = \WX4692_reg/NET0131  & ~\WX4756_reg/NET0131  ;
  assign n2860 = ~\WX4692_reg/NET0131  & \WX4756_reg/NET0131  ;
  assign n2861 = ~n2859 & ~n2860 ;
  assign n2862 = \WX4564_reg/NET0131  & ~\WX4628_reg/NET0131  ;
  assign n2863 = ~\WX4564_reg/NET0131  & \WX4628_reg/NET0131  ;
  assign n2864 = ~n2862 & ~n2863 ;
  assign n2866 = n2861 & ~n2864 ;
  assign n2865 = ~n2861 & n2864 ;
  assign n2867 = ~\TM0_pad  & ~n2865 ;
  assign n2868 = ~n2866 & n2867 ;
  assign n2858 = \TM0_pad  & ~\_2152__reg/NET0131  ;
  assign n2869 = n1976 & ~n2858 ;
  assign n2870 = ~n2868 & n2869 ;
  assign n2871 = ~n2857 & ~n2870 ;
  assign n2872 = n1974 & ~n2801 ;
  assign n2874 = \WX9856_reg/NET0131  & ~\WX9920_reg/NET0131  ;
  assign n2875 = ~\WX9856_reg/NET0131  & \WX9920_reg/NET0131  ;
  assign n2876 = ~n2874 & ~n2875 ;
  assign n2877 = \WX9728_reg/NET0131  & ~\WX9792_reg/NET0131  ;
  assign n2878 = ~\WX9728_reg/NET0131  & \WX9792_reg/NET0131  ;
  assign n2879 = ~n2877 & ~n2878 ;
  assign n2881 = n2876 & ~n2879 ;
  assign n2880 = ~n2876 & n2879 ;
  assign n2882 = ~\TM0_pad  & ~n2880 ;
  assign n2883 = ~n2881 & n2882 ;
  assign n2873 = \TM0_pad  & ~\_2284__reg/NET0131  ;
  assign n2884 = n1976 & ~n2873 ;
  assign n2885 = ~n2883 & n2884 ;
  assign n2886 = ~n2872 & ~n2885 ;
  assign n2887 = \TM0_pad  & \_2135__reg/NET0131  ;
  assign n2888 = \WX3369_reg/NET0131  & ~\WX3433_reg/NET0131  ;
  assign n2889 = ~\WX3369_reg/NET0131  & \WX3433_reg/NET0131  ;
  assign n2890 = ~n2888 & ~n2889 ;
  assign n2891 = \WX3305_reg/NET0131  & ~n2890 ;
  assign n2892 = ~\WX3305_reg/NET0131  & n2890 ;
  assign n2893 = ~n2891 & ~n2892 ;
  assign n2894 = \TM1_pad  & ~\WX3241_reg/NET0131  ;
  assign n2895 = ~\TM1_pad  & \WX3241_reg/NET0131  ;
  assign n2896 = ~n2894 & ~n2895 ;
  assign n2898 = n2893 & ~n2896 ;
  assign n2897 = ~n2893 & n2896 ;
  assign n2899 = ~\TM0_pad  & ~n2897 ;
  assign n2900 = ~n2898 & n2899 ;
  assign n2901 = ~n2887 & ~n2900 ;
  assign n2902 = n1976 & ~n2901 ;
  assign n2903 = ~n1778 & ~n2665 ;
  assign n2904 = n1973 & ~n2903 ;
  assign n2905 = ~n2902 & ~n2904 ;
  assign n2906 = \TM0_pad  & \_2317__reg/NET0131  ;
  assign n2907 = \WX11147_reg/NET0131  & ~\WX11211_reg/NET0131  ;
  assign n2908 = ~\WX11147_reg/NET0131  & \WX11211_reg/NET0131  ;
  assign n2909 = ~n2907 & ~n2908 ;
  assign n2910 = \WX11083_reg/NET0131  & ~n2909 ;
  assign n2911 = ~\WX11083_reg/NET0131  & n2909 ;
  assign n2912 = ~n2910 & ~n2911 ;
  assign n2913 = \TM1_pad  & ~\WX11019_reg/NET0131  ;
  assign n2914 = ~\TM1_pad  & \WX11019_reg/NET0131  ;
  assign n2915 = ~n2913 & ~n2914 ;
  assign n2917 = n2912 & ~n2915 ;
  assign n2916 = ~n2912 & n2915 ;
  assign n2918 = ~\TM0_pad  & ~n2916 ;
  assign n2919 = ~n2917 & n2918 ;
  assign n2920 = ~n2906 & ~n2919 ;
  assign n2921 = n1976 & ~n2920 ;
  assign n2922 = ~n1605 & ~n2716 ;
  assign n2923 = n1973 & ~n2922 ;
  assign n2924 = ~n2921 & ~n2923 ;
  assign n2925 = n2677 & ~n2699 ;
  assign n2927 = \WX5983_reg/NET0131  & ~\WX6047_reg/NET0131  ;
  assign n2928 = ~\WX5983_reg/NET0131  & \WX6047_reg/NET0131  ;
  assign n2929 = ~n2927 & ~n2928 ;
  assign n2930 = \WX5855_reg/NET0131  & ~\WX5919_reg/NET0131  ;
  assign n2931 = ~\WX5855_reg/NET0131  & \WX5919_reg/NET0131  ;
  assign n2932 = ~n2930 & ~n2931 ;
  assign n2934 = n2929 & ~n2932 ;
  assign n2933 = ~n2929 & n2932 ;
  assign n2935 = ~\TM0_pad  & ~n2933 ;
  assign n2936 = ~n2934 & n2935 ;
  assign n2926 = \TM0_pad  & ~\_2185__reg/NET0131  ;
  assign n2937 = n1976 & ~n2926 ;
  assign n2938 = ~n2936 & n2937 ;
  assign n2939 = ~n2925 & ~n2938 ;
  assign n2940 = n2040 & ~n2771 ;
  assign n2942 = \WX7274_reg/NET0131  & ~\WX7338_reg/NET0131  ;
  assign n2943 = ~\WX7274_reg/NET0131  & \WX7338_reg/NET0131  ;
  assign n2944 = ~n2942 & ~n2943 ;
  assign n2945 = \WX7146_reg/NET0131  & ~\WX7210_reg/NET0131  ;
  assign n2946 = ~\WX7146_reg/NET0131  & \WX7210_reg/NET0131  ;
  assign n2947 = ~n2945 & ~n2946 ;
  assign n2949 = n2944 & ~n2947 ;
  assign n2948 = ~n2944 & n2947 ;
  assign n2950 = ~\TM0_pad  & ~n2948 ;
  assign n2951 = ~n2949 & n2950 ;
  assign n2941 = \TM0_pad  & ~\_2218__reg/NET0131  ;
  assign n2952 = n1976 & ~n2941 ;
  assign n2953 = ~n2951 & n2952 ;
  assign n2954 = ~n2940 & ~n2953 ;
  assign n2955 = n2341 & ~n2786 ;
  assign n2957 = \WX8565_reg/NET0131  & ~\WX8629_reg/NET0131  ;
  assign n2958 = ~\WX8565_reg/NET0131  & \WX8629_reg/NET0131  ;
  assign n2959 = ~n2957 & ~n2958 ;
  assign n2960 = \WX8437_reg/NET0131  & ~\WX8501_reg/NET0131  ;
  assign n2961 = ~\WX8437_reg/NET0131  & \WX8501_reg/NET0131  ;
  assign n2962 = ~n2960 & ~n2961 ;
  assign n2964 = n2959 & ~n2962 ;
  assign n2963 = ~n2959 & n2962 ;
  assign n2965 = ~\TM0_pad  & ~n2963 ;
  assign n2966 = ~n2964 & n2965 ;
  assign n2956 = \TM0_pad  & ~\_2251__reg/NET0131  ;
  assign n2967 = n1976 & ~n2956 ;
  assign n2968 = ~n2966 & n2967 ;
  assign n2969 = ~n2955 & ~n2968 ;
  assign n2970 = ~\TM0_pad  & ~n1755 ;
  assign n2971 = ~n1746 & ~n2970 ;
  assign n2972 = n1973 & ~n2971 ;
  assign n2973 = \TM0_pad  & \_2101__reg/NET0131  ;
  assign n2974 = \WX2080_reg/NET0131  & ~\WX2144_reg/NET0131  ;
  assign n2975 = ~\WX2080_reg/NET0131  & \WX2144_reg/NET0131  ;
  assign n2976 = ~n2974 & ~n2975 ;
  assign n2977 = \WX2016_reg/NET0131  & ~n2976 ;
  assign n2978 = ~\WX2016_reg/NET0131  & n2976 ;
  assign n2979 = ~n2977 & ~n2978 ;
  assign n2980 = \TM1_pad  & ~\WX1952_reg/NET0131  ;
  assign n2981 = ~\TM1_pad  & \WX1952_reg/NET0131  ;
  assign n2982 = ~n2980 & ~n2981 ;
  assign n2984 = n2979 & ~n2982 ;
  assign n2983 = ~n2979 & n2982 ;
  assign n2985 = ~\TM0_pad  & ~n2983 ;
  assign n2986 = ~n2984 & n2985 ;
  assign n2987 = ~n2973 & ~n2986 ;
  assign n2988 = n1976 & ~n2987 ;
  assign n2989 = ~n2972 & ~n2988 ;
  assign n2990 = \WX11127_reg/NET0131  & ~\WX11191_reg/NET0131  ;
  assign n2991 = ~\WX11127_reg/NET0131  & \WX11191_reg/NET0131  ;
  assign n2992 = ~n2990 & ~n2991 ;
  assign n2993 = \WX11063_reg/NET0131  & ~n2992 ;
  assign n2994 = ~\WX11063_reg/NET0131  & n2992 ;
  assign n2995 = ~n2993 & ~n2994 ;
  assign n2996 = \TM1_pad  & ~\WX10999_reg/NET0131  ;
  assign n2997 = ~\TM1_pad  & \WX10999_reg/NET0131  ;
  assign n2998 = ~n2996 & ~n2997 ;
  assign n3000 = n2995 & ~n2998 ;
  assign n2999 = ~n2995 & n2998 ;
  assign n3001 = ~\TM0_pad  & ~n2999 ;
  assign n3002 = ~n3000 & n3001 ;
  assign n3003 = ~n1778 & ~n3002 ;
  assign n3004 = n1973 & ~n3003 ;
  assign n3006 = \TM0_pad  & ~\_2359__reg/NET0131  ;
  assign n3005 = ~\DATA_0_26_pad  & ~\TM0_pad  ;
  assign n3007 = n1976 & ~n3005 ;
  assign n3008 = ~n3006 & n3007 ;
  assign n3009 = ~n3004 & ~n3008 ;
  assign n3010 = RESET_pad & \WX10837_reg/NET0131  ;
  assign n3011 = ~n1521 & n1973 ;
  assign n3012 = \WX3401_reg/NET0131  & ~\WX3465_reg/NET0131  ;
  assign n3013 = ~\WX3401_reg/NET0131  & \WX3465_reg/NET0131  ;
  assign n3014 = ~n3012 & ~n3013 ;
  assign n3015 = \WX3273_reg/NET0131  & ~\WX3337_reg/NET0131  ;
  assign n3016 = ~\WX3273_reg/NET0131  & \WX3337_reg/NET0131  ;
  assign n3017 = ~n3015 & ~n3016 ;
  assign n3019 = n3014 & ~n3017 ;
  assign n3018 = ~n3014 & n3017 ;
  assign n3020 = ~\TM0_pad  & ~n3018 ;
  assign n3021 = ~n3019 & n3020 ;
  assign n3022 = n3011 & ~n3021 ;
  assign n3024 = \WX4694_reg/NET0131  & ~\WX4758_reg/NET0131  ;
  assign n3025 = ~\WX4694_reg/NET0131  & \WX4758_reg/NET0131  ;
  assign n3026 = ~n3024 & ~n3025 ;
  assign n3027 = \WX4566_reg/NET0131  & ~\WX4630_reg/NET0131  ;
  assign n3028 = ~\WX4566_reg/NET0131  & \WX4630_reg/NET0131  ;
  assign n3029 = ~n3027 & ~n3028 ;
  assign n3031 = n3026 & ~n3029 ;
  assign n3030 = ~n3026 & n3029 ;
  assign n3032 = ~\TM0_pad  & ~n3030 ;
  assign n3033 = ~n3031 & n3032 ;
  assign n3023 = \TM0_pad  & ~\_2151__reg/NET0131  ;
  assign n3034 = n1976 & ~n3023 ;
  assign n3035 = ~n3033 & n3034 ;
  assign n3036 = ~n3022 & ~n3035 ;
  assign n3037 = n2341 & ~n2966 ;
  assign n3039 = \WX9858_reg/NET0131  & ~\WX9922_reg/NET0131  ;
  assign n3040 = ~\WX9858_reg/NET0131  & \WX9922_reg/NET0131  ;
  assign n3041 = ~n3039 & ~n3040 ;
  assign n3042 = \WX9730_reg/NET0131  & ~\WX9794_reg/NET0131  ;
  assign n3043 = ~\WX9730_reg/NET0131  & \WX9794_reg/NET0131  ;
  assign n3044 = ~n3042 & ~n3043 ;
  assign n3046 = n3041 & ~n3044 ;
  assign n3045 = ~n3041 & n3044 ;
  assign n3047 = ~\TM0_pad  & ~n3045 ;
  assign n3048 = ~n3046 & n3047 ;
  assign n3038 = \TM0_pad  & ~\_2283__reg/NET0131  ;
  assign n3049 = n1976 & ~n3038 ;
  assign n3050 = ~n3048 & n3049 ;
  assign n3051 = ~n3037 & ~n3050 ;
  assign n3052 = \TM0_pad  & \_2134__reg/NET0131  ;
  assign n3053 = \WX3371_reg/NET0131  & ~\WX3435_reg/NET0131  ;
  assign n3054 = ~\WX3371_reg/NET0131  & \WX3435_reg/NET0131  ;
  assign n3055 = ~n3053 & ~n3054 ;
  assign n3056 = \WX3307_reg/NET0131  & ~n3055 ;
  assign n3057 = ~\WX3307_reg/NET0131  & n3055 ;
  assign n3058 = ~n3056 & ~n3057 ;
  assign n3059 = \TM1_pad  & ~\WX3243_reg/NET0131  ;
  assign n3060 = ~\TM1_pad  & \WX3243_reg/NET0131  ;
  assign n3061 = ~n3059 & ~n3060 ;
  assign n3063 = n3058 & ~n3061 ;
  assign n3062 = ~n3058 & n3061 ;
  assign n3064 = ~\TM0_pad  & ~n3062 ;
  assign n3065 = ~n3063 & n3064 ;
  assign n3066 = ~n3052 & ~n3065 ;
  assign n3067 = n1976 & ~n3066 ;
  assign n3068 = ~n1762 & ~n2821 ;
  assign n3069 = n1973 & ~n3068 ;
  assign n3070 = ~n3067 & ~n3069 ;
  assign n3071 = n1974 & ~n2883 ;
  assign n3073 = \WX11149_reg/NET0131  & ~\WX11213_reg/NET0131  ;
  assign n3074 = ~\WX11149_reg/NET0131  & \WX11213_reg/NET0131  ;
  assign n3075 = ~n3073 & ~n3074 ;
  assign n3076 = \WX11021_reg/NET0131  & ~\WX11085_reg/NET0131  ;
  assign n3077 = ~\WX11021_reg/NET0131  & \WX11085_reg/NET0131  ;
  assign n3078 = ~n3076 & ~n3077 ;
  assign n3080 = n3075 & ~n3078 ;
  assign n3079 = ~n3075 & n3078 ;
  assign n3081 = ~\TM0_pad  & ~n3079 ;
  assign n3082 = ~n3080 & n3081 ;
  assign n3072 = \TM0_pad  & ~\_2316__reg/NET0131  ;
  assign n3083 = n1976 & ~n3072 ;
  assign n3084 = ~n3082 & n3083 ;
  assign n3085 = ~n3071 & ~n3084 ;
  assign n3086 = n2846 & ~n2868 ;
  assign n3088 = \WX5985_reg/NET0131  & ~\WX6049_reg/NET0131  ;
  assign n3089 = ~\WX5985_reg/NET0131  & \WX6049_reg/NET0131  ;
  assign n3090 = ~n3088 & ~n3089 ;
  assign n3091 = \WX5857_reg/NET0131  & ~\WX5921_reg/NET0131  ;
  assign n3092 = ~\WX5857_reg/NET0131  & \WX5921_reg/NET0131  ;
  assign n3093 = ~n3091 & ~n3092 ;
  assign n3095 = n3090 & ~n3093 ;
  assign n3094 = ~n3090 & n3093 ;
  assign n3096 = ~\TM0_pad  & ~n3094 ;
  assign n3097 = ~n3095 & n3096 ;
  assign n3087 = \TM0_pad  & ~\_2184__reg/NET0131  ;
  assign n3098 = n1976 & ~n3087 ;
  assign n3099 = ~n3097 & n3098 ;
  assign n3100 = ~n3086 & ~n3099 ;
  assign n3101 = n2677 & ~n2936 ;
  assign n3103 = \WX7276_reg/NET0131  & ~\WX7340_reg/NET0131  ;
  assign n3104 = ~\WX7276_reg/NET0131  & \WX7340_reg/NET0131  ;
  assign n3105 = ~n3103 & ~n3104 ;
  assign n3106 = \WX7148_reg/NET0131  & ~\WX7212_reg/NET0131  ;
  assign n3107 = ~\WX7148_reg/NET0131  & \WX7212_reg/NET0131  ;
  assign n3108 = ~n3106 & ~n3107 ;
  assign n3110 = n3105 & ~n3108 ;
  assign n3109 = ~n3105 & n3108 ;
  assign n3111 = ~\TM0_pad  & ~n3109 ;
  assign n3112 = ~n3110 & n3111 ;
  assign n3102 = \TM0_pad  & ~\_2217__reg/NET0131  ;
  assign n3113 = n1976 & ~n3102 ;
  assign n3114 = ~n3112 & n3113 ;
  assign n3115 = ~n3101 & ~n3114 ;
  assign n3116 = n2040 & ~n2951 ;
  assign n3118 = \WX8567_reg/NET0131  & ~\WX8631_reg/NET0131  ;
  assign n3119 = ~\WX8567_reg/NET0131  & \WX8631_reg/NET0131  ;
  assign n3120 = ~n3118 & ~n3119 ;
  assign n3121 = \WX8439_reg/NET0131  & ~\WX8503_reg/NET0131  ;
  assign n3122 = ~\WX8439_reg/NET0131  & \WX8503_reg/NET0131  ;
  assign n3123 = ~n3121 & ~n3122 ;
  assign n3125 = n3120 & ~n3123 ;
  assign n3124 = ~n3120 & n3123 ;
  assign n3126 = ~\TM0_pad  & ~n3124 ;
  assign n3127 = ~n3125 & n3126 ;
  assign n3117 = \TM0_pad  & ~\_2250__reg/NET0131  ;
  assign n3128 = n1976 & ~n3117 ;
  assign n3129 = ~n3127 & n3128 ;
  assign n3130 = ~n3116 & ~n3129 ;
  assign n3131 = ~\TM0_pad  & ~n1739 ;
  assign n3132 = ~n1730 & ~n3131 ;
  assign n3133 = n1973 & ~n3132 ;
  assign n3134 = \TM0_pad  & \_2100__reg/NET0131  ;
  assign n3135 = \WX2082_reg/NET0131  & ~\WX2146_reg/NET0131  ;
  assign n3136 = ~\WX2082_reg/NET0131  & \WX2146_reg/NET0131  ;
  assign n3137 = ~n3135 & ~n3136 ;
  assign n3138 = \WX2018_reg/NET0131  & ~n3137 ;
  assign n3139 = ~\WX2018_reg/NET0131  & n3137 ;
  assign n3140 = ~n3138 & ~n3139 ;
  assign n3141 = \TM1_pad  & ~\WX1954_reg/NET0131  ;
  assign n3142 = ~\TM1_pad  & \WX1954_reg/NET0131  ;
  assign n3143 = ~n3141 & ~n3142 ;
  assign n3145 = n3140 & ~n3143 ;
  assign n3144 = ~n3140 & n3143 ;
  assign n3146 = ~\TM0_pad  & ~n3144 ;
  assign n3147 = ~n3145 & n3146 ;
  assign n3148 = ~n3134 & ~n3147 ;
  assign n3149 = n1976 & ~n3148 ;
  assign n3150 = ~n3133 & ~n3149 ;
  assign n3151 = \WX11129_reg/NET0131  & ~\WX11193_reg/NET0131  ;
  assign n3152 = ~\WX11129_reg/NET0131  & \WX11193_reg/NET0131  ;
  assign n3153 = ~n3151 & ~n3152 ;
  assign n3154 = \WX11065_reg/NET0131  & ~n3153 ;
  assign n3155 = ~\WX11065_reg/NET0131  & n3153 ;
  assign n3156 = ~n3154 & ~n3155 ;
  assign n3157 = \TM1_pad  & ~\WX11001_reg/NET0131  ;
  assign n3158 = ~\TM1_pad  & \WX11001_reg/NET0131  ;
  assign n3159 = ~n3157 & ~n3158 ;
  assign n3161 = n3156 & ~n3159 ;
  assign n3160 = ~n3156 & n3159 ;
  assign n3162 = ~\TM0_pad  & ~n3160 ;
  assign n3163 = ~n3161 & n3162 ;
  assign n3164 = ~n1762 & ~n3163 ;
  assign n3165 = n1973 & ~n3164 ;
  assign n3167 = \TM0_pad  & ~\_2358__reg/NET0131  ;
  assign n3166 = ~\DATA_0_25_pad  & ~\TM0_pad  ;
  assign n3168 = n1976 & ~n3166 ;
  assign n3169 = ~n3167 & n3168 ;
  assign n3170 = ~n3165 & ~n3169 ;
  assign n3171 = RESET_pad & \WX10839_reg/NET0131  ;
  assign n3172 = ~n1959 & n1973 ;
  assign n3173 = \WX3403_reg/NET0131  & ~\WX3467_reg/NET0131  ;
  assign n3174 = ~\WX3403_reg/NET0131  & \WX3467_reg/NET0131  ;
  assign n3175 = ~n3173 & ~n3174 ;
  assign n3176 = \WX3275_reg/NET0131  & ~\WX3339_reg/NET0131  ;
  assign n3177 = ~\WX3275_reg/NET0131  & \WX3339_reg/NET0131  ;
  assign n3178 = ~n3176 & ~n3177 ;
  assign n3180 = n3175 & ~n3178 ;
  assign n3179 = ~n3175 & n3178 ;
  assign n3181 = ~\TM0_pad  & ~n3179 ;
  assign n3182 = ~n3180 & n3181 ;
  assign n3183 = n3172 & ~n3182 ;
  assign n3185 = \WX4696_reg/NET0131  & ~\WX4760_reg/NET0131  ;
  assign n3186 = ~\WX4696_reg/NET0131  & \WX4760_reg/NET0131  ;
  assign n3187 = ~n3185 & ~n3186 ;
  assign n3188 = \WX4568_reg/NET0131  & ~\WX4632_reg/NET0131  ;
  assign n3189 = ~\WX4568_reg/NET0131  & \WX4632_reg/NET0131  ;
  assign n3190 = ~n3188 & ~n3189 ;
  assign n3192 = n3187 & ~n3190 ;
  assign n3191 = ~n3187 & n3190 ;
  assign n3193 = ~\TM0_pad  & ~n3191 ;
  assign n3194 = ~n3192 & n3193 ;
  assign n3184 = \TM0_pad  & ~\_2150__reg/NET0131  ;
  assign n3195 = n1976 & ~n3184 ;
  assign n3196 = ~n3194 & n3195 ;
  assign n3197 = ~n3183 & ~n3196 ;
  assign n3198 = n2040 & ~n3127 ;
  assign n3200 = \WX9860_reg/NET0131  & ~\WX9924_reg/NET0131  ;
  assign n3201 = ~\WX9860_reg/NET0131  & \WX9924_reg/NET0131  ;
  assign n3202 = ~n3200 & ~n3201 ;
  assign n3203 = \WX9732_reg/NET0131  & ~\WX9796_reg/NET0131  ;
  assign n3204 = ~\WX9732_reg/NET0131  & \WX9796_reg/NET0131  ;
  assign n3205 = ~n3203 & ~n3204 ;
  assign n3207 = n3202 & ~n3205 ;
  assign n3206 = ~n3202 & n3205 ;
  assign n3208 = ~\TM0_pad  & ~n3206 ;
  assign n3209 = ~n3207 & n3208 ;
  assign n3199 = \TM0_pad  & ~\_2282__reg/NET0131  ;
  assign n3210 = n1976 & ~n3199 ;
  assign n3211 = ~n3209 & n3210 ;
  assign n3212 = ~n3198 & ~n3211 ;
  assign n3213 = n2341 & ~n3048 ;
  assign n3215 = \WX11151_reg/NET0131  & ~\WX11215_reg/NET0131  ;
  assign n3216 = ~\WX11151_reg/NET0131  & \WX11215_reg/NET0131  ;
  assign n3217 = ~n3215 & ~n3216 ;
  assign n3218 = \WX11023_reg/NET0131  & ~\WX11087_reg/NET0131  ;
  assign n3219 = ~\WX11023_reg/NET0131  & \WX11087_reg/NET0131  ;
  assign n3220 = ~n3218 & ~n3219 ;
  assign n3222 = n3217 & ~n3220 ;
  assign n3221 = ~n3217 & n3220 ;
  assign n3223 = ~\TM0_pad  & ~n3221 ;
  assign n3224 = ~n3222 & n3223 ;
  assign n3214 = \TM0_pad  & ~\_2315__reg/NET0131  ;
  assign n3225 = n1976 & ~n3214 ;
  assign n3226 = ~n3224 & n3225 ;
  assign n3227 = ~n3213 & ~n3226 ;
  assign n3228 = \TM0_pad  & \_2133__reg/NET0131  ;
  assign n3229 = \WX3373_reg/NET0131  & ~\WX3437_reg/NET0131  ;
  assign n3230 = ~\WX3373_reg/NET0131  & \WX3437_reg/NET0131  ;
  assign n3231 = ~n3229 & ~n3230 ;
  assign n3232 = \WX3309_reg/NET0131  & ~n3231 ;
  assign n3233 = ~\WX3309_reg/NET0131  & n3231 ;
  assign n3234 = ~n3232 & ~n3233 ;
  assign n3235 = \TM1_pad  & ~\WX3245_reg/NET0131  ;
  assign n3236 = ~\TM1_pad  & \WX3245_reg/NET0131  ;
  assign n3237 = ~n3235 & ~n3236 ;
  assign n3239 = n3234 & ~n3237 ;
  assign n3238 = ~n3234 & n3237 ;
  assign n3240 = ~\TM0_pad  & ~n3238 ;
  assign n3241 = ~n3239 & n3240 ;
  assign n3242 = ~n3228 & ~n3241 ;
  assign n3243 = n1976 & ~n3242 ;
  assign n3244 = ~n1746 & ~n2986 ;
  assign n3245 = n1973 & ~n3244 ;
  assign n3246 = ~n3243 & ~n3245 ;
  assign n3247 = n3011 & ~n3033 ;
  assign n3249 = \WX5987_reg/NET0131  & ~\WX6051_reg/NET0131  ;
  assign n3250 = ~\WX5987_reg/NET0131  & \WX6051_reg/NET0131  ;
  assign n3251 = ~n3249 & ~n3250 ;
  assign n3252 = \WX5859_reg/NET0131  & ~\WX5923_reg/NET0131  ;
  assign n3253 = ~\WX5859_reg/NET0131  & \WX5923_reg/NET0131  ;
  assign n3254 = ~n3252 & ~n3253 ;
  assign n3256 = n3251 & ~n3254 ;
  assign n3255 = ~n3251 & n3254 ;
  assign n3257 = ~\TM0_pad  & ~n3255 ;
  assign n3258 = ~n3256 & n3257 ;
  assign n3248 = \TM0_pad  & ~\_2183__reg/NET0131  ;
  assign n3259 = n1976 & ~n3248 ;
  assign n3260 = ~n3258 & n3259 ;
  assign n3261 = ~n3247 & ~n3260 ;
  assign n3262 = n2846 & ~n3097 ;
  assign n3264 = \WX7278_reg/NET0131  & ~\WX7342_reg/NET0131  ;
  assign n3265 = ~\WX7278_reg/NET0131  & \WX7342_reg/NET0131  ;
  assign n3266 = ~n3264 & ~n3265 ;
  assign n3267 = \WX7150_reg/NET0131  & ~\WX7214_reg/NET0131  ;
  assign n3268 = ~\WX7150_reg/NET0131  & \WX7214_reg/NET0131  ;
  assign n3269 = ~n3267 & ~n3268 ;
  assign n3271 = n3266 & ~n3269 ;
  assign n3270 = ~n3266 & n3269 ;
  assign n3272 = ~\TM0_pad  & ~n3270 ;
  assign n3273 = ~n3271 & n3272 ;
  assign n3263 = \TM0_pad  & ~\_2216__reg/NET0131  ;
  assign n3274 = n1976 & ~n3263 ;
  assign n3275 = ~n3273 & n3274 ;
  assign n3276 = ~n3262 & ~n3275 ;
  assign n3277 = n2677 & ~n3112 ;
  assign n3279 = \WX8569_reg/NET0131  & ~\WX8633_reg/NET0131  ;
  assign n3280 = ~\WX8569_reg/NET0131  & \WX8633_reg/NET0131  ;
  assign n3281 = ~n3279 & ~n3280 ;
  assign n3282 = \WX8441_reg/NET0131  & ~\WX8505_reg/NET0131  ;
  assign n3283 = ~\WX8441_reg/NET0131  & \WX8505_reg/NET0131  ;
  assign n3284 = ~n3282 & ~n3283 ;
  assign n3286 = n3281 & ~n3284 ;
  assign n3285 = ~n3281 & n3284 ;
  assign n3287 = ~\TM0_pad  & ~n3285 ;
  assign n3288 = ~n3286 & n3287 ;
  assign n3278 = \TM0_pad  & ~\_2249__reg/NET0131  ;
  assign n3289 = n1976 & ~n3278 ;
  assign n3290 = ~n3288 & n3289 ;
  assign n3291 = ~n3277 & ~n3290 ;
  assign n3292 = ~\TM0_pad  & ~n1723 ;
  assign n3293 = ~n1714 & ~n3292 ;
  assign n3294 = n1973 & ~n3293 ;
  assign n3295 = \TM0_pad  & \_2099__reg/NET0131  ;
  assign n3296 = \WX2084_reg/NET0131  & ~\WX2148_reg/NET0131  ;
  assign n3297 = ~\WX2084_reg/NET0131  & \WX2148_reg/NET0131  ;
  assign n3298 = ~n3296 & ~n3297 ;
  assign n3299 = \WX2020_reg/NET0131  & ~n3298 ;
  assign n3300 = ~\WX2020_reg/NET0131  & n3298 ;
  assign n3301 = ~n3299 & ~n3300 ;
  assign n3302 = \TM1_pad  & ~\WX1956_reg/NET0131  ;
  assign n3303 = ~\TM1_pad  & \WX1956_reg/NET0131  ;
  assign n3304 = ~n3302 & ~n3303 ;
  assign n3306 = n3301 & ~n3304 ;
  assign n3305 = ~n3301 & n3304 ;
  assign n3307 = ~\TM0_pad  & ~n3305 ;
  assign n3308 = ~n3306 & n3307 ;
  assign n3309 = ~n3295 & ~n3308 ;
  assign n3310 = n1976 & ~n3309 ;
  assign n3311 = ~n3294 & ~n3310 ;
  assign n3312 = \WX11131_reg/NET0131  & ~\WX11195_reg/NET0131  ;
  assign n3313 = ~\WX11131_reg/NET0131  & \WX11195_reg/NET0131  ;
  assign n3314 = ~n3312 & ~n3313 ;
  assign n3315 = \WX11067_reg/NET0131  & ~n3314 ;
  assign n3316 = ~\WX11067_reg/NET0131  & n3314 ;
  assign n3317 = ~n3315 & ~n3316 ;
  assign n3318 = \TM1_pad  & ~\WX11003_reg/NET0131  ;
  assign n3319 = ~\TM1_pad  & \WX11003_reg/NET0131  ;
  assign n3320 = ~n3318 & ~n3319 ;
  assign n3322 = n3317 & ~n3320 ;
  assign n3321 = ~n3317 & n3320 ;
  assign n3323 = ~\TM0_pad  & ~n3321 ;
  assign n3324 = ~n3322 & n3323 ;
  assign n3325 = ~n1746 & ~n3324 ;
  assign n3326 = n1973 & ~n3325 ;
  assign n3328 = \TM0_pad  & ~\_2357__reg/NET0131  ;
  assign n3327 = ~\DATA_0_24_pad  & ~\TM0_pad  ;
  assign n3329 = n1976 & ~n3327 ;
  assign n3330 = ~n3328 & n3329 ;
  assign n3331 = ~n3326 & ~n3330 ;
  assign n3332 = RESET_pad & \WX10841_reg/NET0131  ;
  assign n3333 = \WX3405_reg/NET0131  & ~\WX3469_reg/NET0131  ;
  assign n3334 = ~\WX3405_reg/NET0131  & \WX3469_reg/NET0131  ;
  assign n3335 = ~n3333 & ~n3334 ;
  assign n3336 = \WX3277_reg/NET0131  & ~\WX3341_reg/NET0131  ;
  assign n3337 = ~\WX3277_reg/NET0131  & \WX3341_reg/NET0131  ;
  assign n3338 = ~n3336 & ~n3337 ;
  assign n3340 = n3335 & ~n3338 ;
  assign n3339 = ~n3335 & n3338 ;
  assign n3341 = ~\TM0_pad  & ~n3339 ;
  assign n3342 = ~n3340 & n3341 ;
  assign n3343 = n2023 & ~n3342 ;
  assign n3345 = \WX4698_reg/NET0131  & ~\WX4762_reg/NET0131  ;
  assign n3346 = ~\WX4698_reg/NET0131  & \WX4762_reg/NET0131  ;
  assign n3347 = ~n3345 & ~n3346 ;
  assign n3348 = \WX4570_reg/NET0131  & ~\WX4634_reg/NET0131  ;
  assign n3349 = ~\WX4570_reg/NET0131  & \WX4634_reg/NET0131  ;
  assign n3350 = ~n3348 & ~n3349 ;
  assign n3352 = n3347 & ~n3350 ;
  assign n3351 = ~n3347 & n3350 ;
  assign n3353 = ~\TM0_pad  & ~n3351 ;
  assign n3354 = ~n3352 & n3353 ;
  assign n3344 = \TM0_pad  & ~\_2149__reg/NET0131  ;
  assign n3355 = n1976 & ~n3344 ;
  assign n3356 = ~n3354 & n3355 ;
  assign n3357 = ~n3343 & ~n3356 ;
  assign n3358 = n2677 & ~n3288 ;
  assign n3360 = \WX9862_reg/NET0131  & ~\WX9926_reg/NET0131  ;
  assign n3361 = ~\WX9862_reg/NET0131  & \WX9926_reg/NET0131  ;
  assign n3362 = ~n3360 & ~n3361 ;
  assign n3363 = \WX9734_reg/NET0131  & ~\WX9798_reg/NET0131  ;
  assign n3364 = ~\WX9734_reg/NET0131  & \WX9798_reg/NET0131  ;
  assign n3365 = ~n3363 & ~n3364 ;
  assign n3367 = n3362 & ~n3365 ;
  assign n3366 = ~n3362 & n3365 ;
  assign n3368 = ~\TM0_pad  & ~n3366 ;
  assign n3369 = ~n3367 & n3368 ;
  assign n3359 = \TM0_pad  & ~\_2281__reg/NET0131  ;
  assign n3370 = n1976 & ~n3359 ;
  assign n3371 = ~n3369 & n3370 ;
  assign n3372 = ~n3358 & ~n3371 ;
  assign n3373 = n2040 & ~n3209 ;
  assign n3374 = \TM0_pad  & ~\_2314__reg/NET0131  ;
  assign n3375 = n1976 & ~n3374 ;
  assign n3376 = ~n2050 & n3375 ;
  assign n3377 = ~n3373 & ~n3376 ;
  assign n3378 = \TM0_pad  & \_2132__reg/NET0131  ;
  assign n3379 = \WX3375_reg/NET0131  & ~\WX3439_reg/NET0131  ;
  assign n3380 = ~\WX3375_reg/NET0131  & \WX3439_reg/NET0131  ;
  assign n3381 = ~n3379 & ~n3380 ;
  assign n3382 = \WX3311_reg/NET0131  & ~n3381 ;
  assign n3383 = ~\WX3311_reg/NET0131  & n3381 ;
  assign n3384 = ~n3382 & ~n3383 ;
  assign n3385 = \TM1_pad  & ~\WX3247_reg/NET0131  ;
  assign n3386 = ~\TM1_pad  & \WX3247_reg/NET0131  ;
  assign n3387 = ~n3385 & ~n3386 ;
  assign n3389 = n3384 & ~n3387 ;
  assign n3388 = ~n3384 & n3387 ;
  assign n3390 = ~\TM0_pad  & ~n3388 ;
  assign n3391 = ~n3389 & n3390 ;
  assign n3392 = ~n3378 & ~n3391 ;
  assign n3393 = n1976 & ~n3392 ;
  assign n3394 = ~n1730 & ~n3147 ;
  assign n3395 = n1973 & ~n3394 ;
  assign n3396 = ~n3393 & ~n3395 ;
  assign n3397 = n3172 & ~n3194 ;
  assign n3399 = \WX5989_reg/NET0131  & ~\WX6053_reg/NET0131  ;
  assign n3400 = ~\WX5989_reg/NET0131  & \WX6053_reg/NET0131  ;
  assign n3401 = ~n3399 & ~n3400 ;
  assign n3402 = \WX5861_reg/NET0131  & ~\WX5925_reg/NET0131  ;
  assign n3403 = ~\WX5861_reg/NET0131  & \WX5925_reg/NET0131  ;
  assign n3404 = ~n3402 & ~n3403 ;
  assign n3406 = n3401 & ~n3404 ;
  assign n3405 = ~n3401 & n3404 ;
  assign n3407 = ~\TM0_pad  & ~n3405 ;
  assign n3408 = ~n3406 & n3407 ;
  assign n3398 = \TM0_pad  & ~\_2182__reg/NET0131  ;
  assign n3409 = n1976 & ~n3398 ;
  assign n3410 = ~n3408 & n3409 ;
  assign n3411 = ~n3397 & ~n3410 ;
  assign n3412 = n3011 & ~n3258 ;
  assign n3414 = \WX7280_reg/NET0131  & ~\WX7344_reg/NET0131  ;
  assign n3415 = ~\WX7280_reg/NET0131  & \WX7344_reg/NET0131  ;
  assign n3416 = ~n3414 & ~n3415 ;
  assign n3417 = \WX7152_reg/NET0131  & ~\WX7216_reg/NET0131  ;
  assign n3418 = ~\WX7152_reg/NET0131  & \WX7216_reg/NET0131  ;
  assign n3419 = ~n3417 & ~n3418 ;
  assign n3421 = n3416 & ~n3419 ;
  assign n3420 = ~n3416 & n3419 ;
  assign n3422 = ~\TM0_pad  & ~n3420 ;
  assign n3423 = ~n3421 & n3422 ;
  assign n3413 = \TM0_pad  & ~\_2215__reg/NET0131  ;
  assign n3424 = n1976 & ~n3413 ;
  assign n3425 = ~n3423 & n3424 ;
  assign n3426 = ~n3412 & ~n3425 ;
  assign n3427 = n2846 & ~n3273 ;
  assign n3429 = \WX8571_reg/NET0131  & ~\WX8635_reg/NET0131  ;
  assign n3430 = ~\WX8571_reg/NET0131  & \WX8635_reg/NET0131  ;
  assign n3431 = ~n3429 & ~n3430 ;
  assign n3432 = \WX8443_reg/NET0131  & ~\WX8507_reg/NET0131  ;
  assign n3433 = ~\WX8443_reg/NET0131  & \WX8507_reg/NET0131  ;
  assign n3434 = ~n3432 & ~n3433 ;
  assign n3436 = n3431 & ~n3434 ;
  assign n3435 = ~n3431 & n3434 ;
  assign n3437 = ~\TM0_pad  & ~n3435 ;
  assign n3438 = ~n3436 & n3437 ;
  assign n3428 = \TM0_pad  & ~\_2248__reg/NET0131  ;
  assign n3439 = n1976 & ~n3428 ;
  assign n3440 = ~n3438 & n3439 ;
  assign n3441 = ~n3427 & ~n3440 ;
  assign n3442 = ~\TM0_pad  & ~n1707 ;
  assign n3443 = ~n1698 & ~n3442 ;
  assign n3444 = n1973 & ~n3443 ;
  assign n3445 = \TM0_pad  & \_2098__reg/NET0131  ;
  assign n3446 = \WX2086_reg/NET0131  & ~\WX2150_reg/NET0131  ;
  assign n3447 = ~\WX2086_reg/NET0131  & \WX2150_reg/NET0131  ;
  assign n3448 = ~n3446 & ~n3447 ;
  assign n3449 = \WX2022_reg/NET0131  & ~n3448 ;
  assign n3450 = ~\WX2022_reg/NET0131  & n3448 ;
  assign n3451 = ~n3449 & ~n3450 ;
  assign n3452 = \TM1_pad  & ~\WX1958_reg/NET0131  ;
  assign n3453 = ~\TM1_pad  & \WX1958_reg/NET0131  ;
  assign n3454 = ~n3452 & ~n3453 ;
  assign n3456 = n3451 & ~n3454 ;
  assign n3455 = ~n3451 & n3454 ;
  assign n3457 = ~\TM0_pad  & ~n3455 ;
  assign n3458 = ~n3456 & n3457 ;
  assign n3459 = ~n3445 & ~n3458 ;
  assign n3460 = n1976 & ~n3459 ;
  assign n3461 = ~n3444 & ~n3460 ;
  assign n3462 = \WX11133_reg/NET0131  & ~\WX11197_reg/NET0131  ;
  assign n3463 = ~\WX11133_reg/NET0131  & \WX11197_reg/NET0131  ;
  assign n3464 = ~n3462 & ~n3463 ;
  assign n3465 = \WX11069_reg/NET0131  & ~n3464 ;
  assign n3466 = ~\WX11069_reg/NET0131  & n3464 ;
  assign n3467 = ~n3465 & ~n3466 ;
  assign n3468 = \TM1_pad  & ~\WX11005_reg/NET0131  ;
  assign n3469 = ~\TM1_pad  & \WX11005_reg/NET0131  ;
  assign n3470 = ~n3468 & ~n3469 ;
  assign n3472 = n3467 & ~n3470 ;
  assign n3471 = ~n3467 & n3470 ;
  assign n3473 = ~\TM0_pad  & ~n3471 ;
  assign n3474 = ~n3472 & n3473 ;
  assign n3475 = ~n1730 & ~n3474 ;
  assign n3476 = n1973 & ~n3475 ;
  assign n3478 = \TM0_pad  & ~\_2356__reg/NET0131  ;
  assign n3477 = ~\DATA_0_23_pad  & ~\TM0_pad  ;
  assign n3479 = n1976 & ~n3477 ;
  assign n3480 = ~n3478 & n3479 ;
  assign n3481 = ~n3476 & ~n3480 ;
  assign n3482 = RESET_pad & \WX10843_reg/NET0131  ;
  assign n3483 = ~n1933 & n1973 ;
  assign n3484 = \WX3407_reg/NET0131  & ~\WX3471_reg/NET0131  ;
  assign n3485 = ~\WX3407_reg/NET0131  & \WX3471_reg/NET0131  ;
  assign n3486 = ~n3484 & ~n3485 ;
  assign n3487 = \WX3279_reg/NET0131  & ~\WX3343_reg/NET0131  ;
  assign n3488 = ~\WX3279_reg/NET0131  & \WX3343_reg/NET0131  ;
  assign n3489 = ~n3487 & ~n3488 ;
  assign n3491 = n3486 & ~n3489 ;
  assign n3490 = ~n3486 & n3489 ;
  assign n3492 = ~\TM0_pad  & ~n3490 ;
  assign n3493 = ~n3491 & n3492 ;
  assign n3494 = n3483 & ~n3493 ;
  assign n3496 = \WX4700_reg/NET0131  & ~\WX4764_reg/NET0131  ;
  assign n3497 = ~\WX4700_reg/NET0131  & \WX4764_reg/NET0131  ;
  assign n3498 = ~n3496 & ~n3497 ;
  assign n3499 = \WX4572_reg/NET0131  & ~\WX4636_reg/NET0131  ;
  assign n3500 = ~\WX4572_reg/NET0131  & \WX4636_reg/NET0131  ;
  assign n3501 = ~n3499 & ~n3500 ;
  assign n3503 = n3498 & ~n3501 ;
  assign n3502 = ~n3498 & n3501 ;
  assign n3504 = ~\TM0_pad  & ~n3502 ;
  assign n3505 = ~n3503 & n3504 ;
  assign n3495 = \TM0_pad  & ~\_2148__reg/NET0131  ;
  assign n3506 = n1976 & ~n3495 ;
  assign n3507 = ~n3505 & n3506 ;
  assign n3508 = ~n3494 & ~n3507 ;
  assign n3509 = n2846 & ~n3438 ;
  assign n3511 = \WX9864_reg/NET0131  & ~\WX9928_reg/NET0131  ;
  assign n3512 = ~\WX9864_reg/NET0131  & \WX9928_reg/NET0131  ;
  assign n3513 = ~n3511 & ~n3512 ;
  assign n3514 = \WX9736_reg/NET0131  & ~\WX9800_reg/NET0131  ;
  assign n3515 = ~\WX9736_reg/NET0131  & \WX9800_reg/NET0131  ;
  assign n3516 = ~n3514 & ~n3515 ;
  assign n3518 = n3513 & ~n3516 ;
  assign n3517 = ~n3513 & n3516 ;
  assign n3519 = ~\TM0_pad  & ~n3517 ;
  assign n3520 = ~n3518 & n3519 ;
  assign n3510 = \TM0_pad  & ~\_2280__reg/NET0131  ;
  assign n3521 = n1976 & ~n3510 ;
  assign n3522 = ~n3520 & n3521 ;
  assign n3523 = ~n3509 & ~n3522 ;
  assign n3524 = n2677 & ~n3369 ;
  assign n3526 = \WX11155_reg/NET0131  & ~\WX11219_reg/NET0131  ;
  assign n3527 = ~\WX11155_reg/NET0131  & \WX11219_reg/NET0131  ;
  assign n3528 = ~n3526 & ~n3527 ;
  assign n3529 = \WX11027_reg/NET0131  & ~\WX11091_reg/NET0131  ;
  assign n3530 = ~\WX11027_reg/NET0131  & \WX11091_reg/NET0131  ;
  assign n3531 = ~n3529 & ~n3530 ;
  assign n3533 = n3528 & ~n3531 ;
  assign n3532 = ~n3528 & n3531 ;
  assign n3534 = ~\TM0_pad  & ~n3532 ;
  assign n3535 = ~n3533 & n3534 ;
  assign n3525 = \TM0_pad  & ~\_2313__reg/NET0131  ;
  assign n3536 = n1976 & ~n3525 ;
  assign n3537 = ~n3535 & n3536 ;
  assign n3538 = ~n3524 & ~n3537 ;
  assign n3539 = \TM0_pad  & \_2131__reg/NET0131  ;
  assign n3540 = \WX3377_reg/NET0131  & ~\WX3441_reg/NET0131  ;
  assign n3541 = ~\WX3377_reg/NET0131  & \WX3441_reg/NET0131  ;
  assign n3542 = ~n3540 & ~n3541 ;
  assign n3543 = \WX3313_reg/NET0131  & ~n3542 ;
  assign n3544 = ~\WX3313_reg/NET0131  & n3542 ;
  assign n3545 = ~n3543 & ~n3544 ;
  assign n3546 = \TM1_pad  & ~\WX3249_reg/NET0131  ;
  assign n3547 = ~\TM1_pad  & \WX3249_reg/NET0131  ;
  assign n3548 = ~n3546 & ~n3547 ;
  assign n3550 = n3545 & ~n3548 ;
  assign n3549 = ~n3545 & n3548 ;
  assign n3551 = ~\TM0_pad  & ~n3549 ;
  assign n3552 = ~n3550 & n3551 ;
  assign n3553 = ~n3539 & ~n3552 ;
  assign n3554 = n1976 & ~n3553 ;
  assign n3555 = ~n1714 & ~n3308 ;
  assign n3556 = n1973 & ~n3555 ;
  assign n3557 = ~n3554 & ~n3556 ;
  assign n3558 = n2023 & ~n3354 ;
  assign n3560 = \WX5991_reg/NET0131  & ~\WX6055_reg/NET0131  ;
  assign n3561 = ~\WX5991_reg/NET0131  & \WX6055_reg/NET0131  ;
  assign n3562 = ~n3560 & ~n3561 ;
  assign n3563 = \WX5863_reg/NET0131  & ~\WX5927_reg/NET0131  ;
  assign n3564 = ~\WX5863_reg/NET0131  & \WX5927_reg/NET0131  ;
  assign n3565 = ~n3563 & ~n3564 ;
  assign n3567 = n3562 & ~n3565 ;
  assign n3566 = ~n3562 & n3565 ;
  assign n3568 = ~\TM0_pad  & ~n3566 ;
  assign n3569 = ~n3567 & n3568 ;
  assign n3559 = \TM0_pad  & ~\_2181__reg/NET0131  ;
  assign n3570 = n1976 & ~n3559 ;
  assign n3571 = ~n3569 & n3570 ;
  assign n3572 = ~n3558 & ~n3571 ;
  assign n3573 = n3172 & ~n3408 ;
  assign n3575 = \WX7282_reg/NET0131  & ~\WX7346_reg/NET0131  ;
  assign n3576 = ~\WX7282_reg/NET0131  & \WX7346_reg/NET0131  ;
  assign n3577 = ~n3575 & ~n3576 ;
  assign n3578 = \WX7154_reg/NET0131  & ~\WX7218_reg/NET0131  ;
  assign n3579 = ~\WX7154_reg/NET0131  & \WX7218_reg/NET0131  ;
  assign n3580 = ~n3578 & ~n3579 ;
  assign n3582 = n3577 & ~n3580 ;
  assign n3581 = ~n3577 & n3580 ;
  assign n3583 = ~\TM0_pad  & ~n3581 ;
  assign n3584 = ~n3582 & n3583 ;
  assign n3574 = \TM0_pad  & ~\_2214__reg/NET0131  ;
  assign n3585 = n1976 & ~n3574 ;
  assign n3586 = ~n3584 & n3585 ;
  assign n3587 = ~n3573 & ~n3586 ;
  assign n3588 = n3011 & ~n3423 ;
  assign n3590 = \WX8573_reg/NET0131  & ~\WX8637_reg/NET0131  ;
  assign n3591 = ~\WX8573_reg/NET0131  & \WX8637_reg/NET0131  ;
  assign n3592 = ~n3590 & ~n3591 ;
  assign n3593 = \WX8445_reg/NET0131  & ~\WX8509_reg/NET0131  ;
  assign n3594 = ~\WX8445_reg/NET0131  & \WX8509_reg/NET0131  ;
  assign n3595 = ~n3593 & ~n3594 ;
  assign n3597 = n3592 & ~n3595 ;
  assign n3596 = ~n3592 & n3595 ;
  assign n3598 = ~\TM0_pad  & ~n3596 ;
  assign n3599 = ~n3597 & n3598 ;
  assign n3589 = \TM0_pad  & ~\_2247__reg/NET0131  ;
  assign n3600 = n1976 & ~n3589 ;
  assign n3601 = ~n3599 & n3600 ;
  assign n3602 = ~n3588 & ~n3601 ;
  assign n3603 = ~\TM0_pad  & ~n1691 ;
  assign n3604 = ~n1682 & ~n3603 ;
  assign n3605 = n1973 & ~n3604 ;
  assign n3606 = \TM0_pad  & \_2097__reg/NET0131  ;
  assign n3607 = \WX2088_reg/NET0131  & ~\WX2152_reg/NET0131  ;
  assign n3608 = ~\WX2088_reg/NET0131  & \WX2152_reg/NET0131  ;
  assign n3609 = ~n3607 & ~n3608 ;
  assign n3610 = \WX2024_reg/NET0131  & ~n3609 ;
  assign n3611 = ~\WX2024_reg/NET0131  & n3609 ;
  assign n3612 = ~n3610 & ~n3611 ;
  assign n3613 = \TM1_pad  & ~\WX1960_reg/NET0131  ;
  assign n3614 = ~\TM1_pad  & \WX1960_reg/NET0131  ;
  assign n3615 = ~n3613 & ~n3614 ;
  assign n3617 = n3612 & ~n3615 ;
  assign n3616 = ~n3612 & n3615 ;
  assign n3618 = ~\TM0_pad  & ~n3616 ;
  assign n3619 = ~n3617 & n3618 ;
  assign n3620 = ~n3606 & ~n3619 ;
  assign n3621 = n1976 & ~n3620 ;
  assign n3622 = ~n3605 & ~n3621 ;
  assign n3623 = \WX11135_reg/NET0131  & ~\WX11199_reg/NET0131  ;
  assign n3624 = ~\WX11135_reg/NET0131  & \WX11199_reg/NET0131  ;
  assign n3625 = ~n3623 & ~n3624 ;
  assign n3626 = \WX11071_reg/NET0131  & ~n3625 ;
  assign n3627 = ~\WX11071_reg/NET0131  & n3625 ;
  assign n3628 = ~n3626 & ~n3627 ;
  assign n3629 = \TM1_pad  & ~\WX11007_reg/NET0131  ;
  assign n3630 = ~\TM1_pad  & \WX11007_reg/NET0131  ;
  assign n3631 = ~n3629 & ~n3630 ;
  assign n3633 = n3628 & ~n3631 ;
  assign n3632 = ~n3628 & n3631 ;
  assign n3634 = ~\TM0_pad  & ~n3632 ;
  assign n3635 = ~n3633 & n3634 ;
  assign n3636 = ~n1714 & ~n3635 ;
  assign n3637 = n1973 & ~n3636 ;
  assign n3639 = \TM0_pad  & ~\_2355__reg/NET0131  ;
  assign n3638 = ~\DATA_0_22_pad  & ~\TM0_pad  ;
  assign n3640 = n1976 & ~n3638 ;
  assign n3641 = ~n3639 & n3640 ;
  assign n3642 = ~n3637 & ~n3641 ;
  assign n3643 = RESET_pad & \WX10845_reg/NET0131  ;
  assign n3644 = ~n1920 & n1973 ;
  assign n3645 = \WX3409_reg/NET0131  & ~\WX3473_reg/NET0131  ;
  assign n3646 = ~\WX3409_reg/NET0131  & \WX3473_reg/NET0131  ;
  assign n3647 = ~n3645 & ~n3646 ;
  assign n3648 = \WX3281_reg/NET0131  & ~\WX3345_reg/NET0131  ;
  assign n3649 = ~\WX3281_reg/NET0131  & \WX3345_reg/NET0131  ;
  assign n3650 = ~n3648 & ~n3649 ;
  assign n3652 = n3647 & ~n3650 ;
  assign n3651 = ~n3647 & n3650 ;
  assign n3653 = ~\TM0_pad  & ~n3651 ;
  assign n3654 = ~n3652 & n3653 ;
  assign n3655 = n3644 & ~n3654 ;
  assign n3657 = \WX4702_reg/NET0131  & ~\WX4766_reg/NET0131  ;
  assign n3658 = ~\WX4702_reg/NET0131  & \WX4766_reg/NET0131  ;
  assign n3659 = ~n3657 & ~n3658 ;
  assign n3660 = \WX4574_reg/NET0131  & ~\WX4638_reg/NET0131  ;
  assign n3661 = ~\WX4574_reg/NET0131  & \WX4638_reg/NET0131  ;
  assign n3662 = ~n3660 & ~n3661 ;
  assign n3664 = n3659 & ~n3662 ;
  assign n3663 = ~n3659 & n3662 ;
  assign n3665 = ~\TM0_pad  & ~n3663 ;
  assign n3666 = ~n3664 & n3665 ;
  assign n3656 = \TM0_pad  & ~\_2147__reg/NET0131  ;
  assign n3667 = n1976 & ~n3656 ;
  assign n3668 = ~n3666 & n3667 ;
  assign n3669 = ~n3655 & ~n3668 ;
  assign n3670 = n3011 & ~n3599 ;
  assign n3672 = \WX9866_reg/NET0131  & ~\WX9930_reg/NET0131  ;
  assign n3673 = ~\WX9866_reg/NET0131  & \WX9930_reg/NET0131  ;
  assign n3674 = ~n3672 & ~n3673 ;
  assign n3675 = \WX9738_reg/NET0131  & ~\WX9802_reg/NET0131  ;
  assign n3676 = ~\WX9738_reg/NET0131  & \WX9802_reg/NET0131  ;
  assign n3677 = ~n3675 & ~n3676 ;
  assign n3679 = n3674 & ~n3677 ;
  assign n3678 = ~n3674 & n3677 ;
  assign n3680 = ~\TM0_pad  & ~n3678 ;
  assign n3681 = ~n3679 & n3680 ;
  assign n3671 = \TM0_pad  & ~\_2279__reg/NET0131  ;
  assign n3682 = n1976 & ~n3671 ;
  assign n3683 = ~n3681 & n3682 ;
  assign n3684 = ~n3670 & ~n3683 ;
  assign n3685 = n2846 & ~n3520 ;
  assign n3687 = \WX11157_reg/NET0131  & ~\WX11221_reg/NET0131  ;
  assign n3688 = ~\WX11157_reg/NET0131  & \WX11221_reg/NET0131  ;
  assign n3689 = ~n3687 & ~n3688 ;
  assign n3690 = \WX11029_reg/NET0131  & ~\WX11093_reg/NET0131  ;
  assign n3691 = ~\WX11029_reg/NET0131  & \WX11093_reg/NET0131  ;
  assign n3692 = ~n3690 & ~n3691 ;
  assign n3694 = n3689 & ~n3692 ;
  assign n3693 = ~n3689 & n3692 ;
  assign n3695 = ~\TM0_pad  & ~n3693 ;
  assign n3696 = ~n3694 & n3695 ;
  assign n3686 = \TM0_pad  & ~\_2312__reg/NET0131  ;
  assign n3697 = n1976 & ~n3686 ;
  assign n3698 = ~n3696 & n3697 ;
  assign n3699 = ~n3685 & ~n3698 ;
  assign n3700 = \TM0_pad  & \_2130__reg/NET0131  ;
  assign n3701 = \WX3379_reg/NET0131  & ~\WX3443_reg/NET0131  ;
  assign n3702 = ~\WX3379_reg/NET0131  & \WX3443_reg/NET0131  ;
  assign n3703 = ~n3701 & ~n3702 ;
  assign n3704 = \WX3315_reg/NET0131  & ~n3703 ;
  assign n3705 = ~\WX3315_reg/NET0131  & n3703 ;
  assign n3706 = ~n3704 & ~n3705 ;
  assign n3707 = \TM1_pad  & ~\WX3251_reg/NET0131  ;
  assign n3708 = ~\TM1_pad  & \WX3251_reg/NET0131  ;
  assign n3709 = ~n3707 & ~n3708 ;
  assign n3711 = n3706 & ~n3709 ;
  assign n3710 = ~n3706 & n3709 ;
  assign n3712 = ~\TM0_pad  & ~n3710 ;
  assign n3713 = ~n3711 & n3712 ;
  assign n3714 = ~n3700 & ~n3713 ;
  assign n3715 = n1976 & ~n3714 ;
  assign n3716 = ~n1698 & ~n3458 ;
  assign n3717 = n1973 & ~n3716 ;
  assign n3718 = ~n3715 & ~n3717 ;
  assign n3719 = n3483 & ~n3505 ;
  assign n3721 = \WX5993_reg/NET0131  & ~\WX6057_reg/NET0131  ;
  assign n3722 = ~\WX5993_reg/NET0131  & \WX6057_reg/NET0131  ;
  assign n3723 = ~n3721 & ~n3722 ;
  assign n3724 = \WX5865_reg/NET0131  & ~\WX5929_reg/NET0131  ;
  assign n3725 = ~\WX5865_reg/NET0131  & \WX5929_reg/NET0131  ;
  assign n3726 = ~n3724 & ~n3725 ;
  assign n3728 = n3723 & ~n3726 ;
  assign n3727 = ~n3723 & n3726 ;
  assign n3729 = ~\TM0_pad  & ~n3727 ;
  assign n3730 = ~n3728 & n3729 ;
  assign n3720 = \TM0_pad  & ~\_2180__reg/NET0131  ;
  assign n3731 = n1976 & ~n3720 ;
  assign n3732 = ~n3730 & n3731 ;
  assign n3733 = ~n3719 & ~n3732 ;
  assign n3734 = n2023 & ~n3569 ;
  assign n3736 = \WX7284_reg/NET0131  & ~\WX7348_reg/NET0131  ;
  assign n3737 = ~\WX7284_reg/NET0131  & \WX7348_reg/NET0131  ;
  assign n3738 = ~n3736 & ~n3737 ;
  assign n3739 = \WX7156_reg/NET0131  & ~\WX7220_reg/NET0131  ;
  assign n3740 = ~\WX7156_reg/NET0131  & \WX7220_reg/NET0131  ;
  assign n3741 = ~n3739 & ~n3740 ;
  assign n3743 = n3738 & ~n3741 ;
  assign n3742 = ~n3738 & n3741 ;
  assign n3744 = ~\TM0_pad  & ~n3742 ;
  assign n3745 = ~n3743 & n3744 ;
  assign n3735 = \TM0_pad  & ~\_2213__reg/NET0131  ;
  assign n3746 = n1976 & ~n3735 ;
  assign n3747 = ~n3745 & n3746 ;
  assign n3748 = ~n3734 & ~n3747 ;
  assign n3749 = n3172 & ~n3584 ;
  assign n3751 = \WX8575_reg/NET0131  & ~\WX8639_reg/NET0131  ;
  assign n3752 = ~\WX8575_reg/NET0131  & \WX8639_reg/NET0131  ;
  assign n3753 = ~n3751 & ~n3752 ;
  assign n3754 = \WX8447_reg/NET0131  & ~\WX8511_reg/NET0131  ;
  assign n3755 = ~\WX8447_reg/NET0131  & \WX8511_reg/NET0131  ;
  assign n3756 = ~n3754 & ~n3755 ;
  assign n3758 = n3753 & ~n3756 ;
  assign n3757 = ~n3753 & n3756 ;
  assign n3759 = ~\TM0_pad  & ~n3757 ;
  assign n3760 = ~n3758 & n3759 ;
  assign n3750 = \TM0_pad  & ~\_2246__reg/NET0131  ;
  assign n3761 = n1976 & ~n3750 ;
  assign n3762 = ~n3760 & n3761 ;
  assign n3763 = ~n3749 & ~n3762 ;
  assign n3764 = ~\TM0_pad  & ~n1662 ;
  assign n3765 = ~n1653 & ~n3764 ;
  assign n3766 = n1973 & ~n3765 ;
  assign n3767 = \TM0_pad  & \_2096__reg/NET0131  ;
  assign n3768 = \WX2090_reg/NET0131  & ~\WX2154_reg/NET0131  ;
  assign n3769 = ~\WX2090_reg/NET0131  & \WX2154_reg/NET0131  ;
  assign n3770 = ~n3768 & ~n3769 ;
  assign n3771 = \WX2026_reg/NET0131  & ~n3770 ;
  assign n3772 = ~\WX2026_reg/NET0131  & n3770 ;
  assign n3773 = ~n3771 & ~n3772 ;
  assign n3774 = \TM1_pad  & ~\WX1962_reg/NET0131  ;
  assign n3775 = ~\TM1_pad  & \WX1962_reg/NET0131  ;
  assign n3776 = ~n3774 & ~n3775 ;
  assign n3778 = n3773 & ~n3776 ;
  assign n3777 = ~n3773 & n3776 ;
  assign n3779 = ~\TM0_pad  & ~n3777 ;
  assign n3780 = ~n3778 & n3779 ;
  assign n3781 = ~n3767 & ~n3780 ;
  assign n3782 = n1976 & ~n3781 ;
  assign n3783 = ~n3766 & ~n3782 ;
  assign n3784 = \WX11137_reg/NET0131  & ~\WX11201_reg/NET0131  ;
  assign n3785 = ~\WX11137_reg/NET0131  & \WX11201_reg/NET0131  ;
  assign n3786 = ~n3784 & ~n3785 ;
  assign n3787 = \WX11073_reg/NET0131  & ~n3786 ;
  assign n3788 = ~\WX11073_reg/NET0131  & n3786 ;
  assign n3789 = ~n3787 & ~n3788 ;
  assign n3790 = \TM1_pad  & ~\WX11009_reg/NET0131  ;
  assign n3791 = ~\TM1_pad  & \WX11009_reg/NET0131  ;
  assign n3792 = ~n3790 & ~n3791 ;
  assign n3794 = n3789 & ~n3792 ;
  assign n3793 = ~n3789 & n3792 ;
  assign n3795 = ~\TM0_pad  & ~n3793 ;
  assign n3796 = ~n3794 & n3795 ;
  assign n3797 = ~n1698 & ~n3796 ;
  assign n3798 = n1973 & ~n3797 ;
  assign n3800 = \TM0_pad  & ~\_2354__reg/NET0131  ;
  assign n3799 = ~\DATA_0_21_pad  & ~\TM0_pad  ;
  assign n3801 = n1976 & ~n3799 ;
  assign n3802 = ~n3800 & n3801 ;
  assign n3803 = ~n3798 & ~n3802 ;
  assign n3804 = RESET_pad & \WX10847_reg/NET0131  ;
  assign n3805 = ~n1907 & n1973 ;
  assign n3806 = \WX3411_reg/NET0131  & ~\WX3475_reg/NET0131  ;
  assign n3807 = ~\WX3411_reg/NET0131  & \WX3475_reg/NET0131  ;
  assign n3808 = ~n3806 & ~n3807 ;
  assign n3809 = \WX3283_reg/NET0131  & ~\WX3347_reg/NET0131  ;
  assign n3810 = ~\WX3283_reg/NET0131  & \WX3347_reg/NET0131  ;
  assign n3811 = ~n3809 & ~n3810 ;
  assign n3813 = n3808 & ~n3811 ;
  assign n3812 = ~n3808 & n3811 ;
  assign n3814 = ~\TM0_pad  & ~n3812 ;
  assign n3815 = ~n3813 & n3814 ;
  assign n3816 = n3805 & ~n3815 ;
  assign n3818 = \WX4704_reg/NET0131  & ~\WX4768_reg/NET0131  ;
  assign n3819 = ~\WX4704_reg/NET0131  & \WX4768_reg/NET0131  ;
  assign n3820 = ~n3818 & ~n3819 ;
  assign n3821 = \WX4576_reg/NET0131  & ~\WX4640_reg/NET0131  ;
  assign n3822 = ~\WX4576_reg/NET0131  & \WX4640_reg/NET0131  ;
  assign n3823 = ~n3821 & ~n3822 ;
  assign n3825 = n3820 & ~n3823 ;
  assign n3824 = ~n3820 & n3823 ;
  assign n3826 = ~\TM0_pad  & ~n3824 ;
  assign n3827 = ~n3825 & n3826 ;
  assign n3817 = \TM0_pad  & ~\_2146__reg/NET0131  ;
  assign n3828 = n1976 & ~n3817 ;
  assign n3829 = ~n3827 & n3828 ;
  assign n3830 = ~n3816 & ~n3829 ;
  assign n3831 = n3172 & ~n3760 ;
  assign n3833 = \WX9868_reg/NET0131  & ~\WX9932_reg/NET0131  ;
  assign n3834 = ~\WX9868_reg/NET0131  & \WX9932_reg/NET0131  ;
  assign n3835 = ~n3833 & ~n3834 ;
  assign n3836 = \WX9740_reg/NET0131  & ~\WX9804_reg/NET0131  ;
  assign n3837 = ~\WX9740_reg/NET0131  & \WX9804_reg/NET0131  ;
  assign n3838 = ~n3836 & ~n3837 ;
  assign n3840 = n3835 & ~n3838 ;
  assign n3839 = ~n3835 & n3838 ;
  assign n3841 = ~\TM0_pad  & ~n3839 ;
  assign n3842 = ~n3840 & n3841 ;
  assign n3832 = \TM0_pad  & ~\_2278__reg/NET0131  ;
  assign n3843 = n1976 & ~n3832 ;
  assign n3844 = ~n3842 & n3843 ;
  assign n3845 = ~n3831 & ~n3844 ;
  assign n3846 = n3011 & ~n3681 ;
  assign n3848 = \WX11159_reg/NET0131  & ~\WX11223_reg/NET0131  ;
  assign n3849 = ~\WX11159_reg/NET0131  & \WX11223_reg/NET0131  ;
  assign n3850 = ~n3848 & ~n3849 ;
  assign n3851 = \WX11031_reg/NET0131  & ~\WX11095_reg/NET0131  ;
  assign n3852 = ~\WX11031_reg/NET0131  & \WX11095_reg/NET0131  ;
  assign n3853 = ~n3851 & ~n3852 ;
  assign n3855 = n3850 & ~n3853 ;
  assign n3854 = ~n3850 & n3853 ;
  assign n3856 = ~\TM0_pad  & ~n3854 ;
  assign n3857 = ~n3855 & n3856 ;
  assign n3847 = \TM0_pad  & ~\_2311__reg/NET0131  ;
  assign n3858 = n1976 & ~n3847 ;
  assign n3859 = ~n3857 & n3858 ;
  assign n3860 = ~n3846 & ~n3859 ;
  assign n3861 = \TM0_pad  & \_2129__reg/NET0131  ;
  assign n3862 = \WX3381_reg/NET0131  & ~\WX3445_reg/NET0131  ;
  assign n3863 = ~\WX3381_reg/NET0131  & \WX3445_reg/NET0131  ;
  assign n3864 = ~n3862 & ~n3863 ;
  assign n3865 = \WX3317_reg/NET0131  & ~n3864 ;
  assign n3866 = ~\WX3317_reg/NET0131  & n3864 ;
  assign n3867 = ~n3865 & ~n3866 ;
  assign n3868 = \TM1_pad  & ~\WX3253_reg/NET0131  ;
  assign n3869 = ~\TM1_pad  & \WX3253_reg/NET0131  ;
  assign n3870 = ~n3868 & ~n3869 ;
  assign n3872 = n3867 & ~n3870 ;
  assign n3871 = ~n3867 & n3870 ;
  assign n3873 = ~\TM0_pad  & ~n3871 ;
  assign n3874 = ~n3872 & n3873 ;
  assign n3875 = ~n3861 & ~n3874 ;
  assign n3876 = n1976 & ~n3875 ;
  assign n3877 = ~n1682 & ~n3619 ;
  assign n3878 = n1973 & ~n3877 ;
  assign n3879 = ~n3876 & ~n3878 ;
  assign n3880 = n3644 & ~n3666 ;
  assign n3882 = \WX5995_reg/NET0131  & ~\WX6059_reg/NET0131  ;
  assign n3883 = ~\WX5995_reg/NET0131  & \WX6059_reg/NET0131  ;
  assign n3884 = ~n3882 & ~n3883 ;
  assign n3885 = \WX5867_reg/NET0131  & ~\WX5931_reg/NET0131  ;
  assign n3886 = ~\WX5867_reg/NET0131  & \WX5931_reg/NET0131  ;
  assign n3887 = ~n3885 & ~n3886 ;
  assign n3889 = n3884 & ~n3887 ;
  assign n3888 = ~n3884 & n3887 ;
  assign n3890 = ~\TM0_pad  & ~n3888 ;
  assign n3891 = ~n3889 & n3890 ;
  assign n3881 = \TM0_pad  & ~\_2179__reg/NET0131  ;
  assign n3892 = n1976 & ~n3881 ;
  assign n3893 = ~n3891 & n3892 ;
  assign n3894 = ~n3880 & ~n3893 ;
  assign n3895 = n3483 & ~n3730 ;
  assign n3897 = \WX7286_reg/NET0131  & ~\WX7350_reg/NET0131  ;
  assign n3898 = ~\WX7286_reg/NET0131  & \WX7350_reg/NET0131  ;
  assign n3899 = ~n3897 & ~n3898 ;
  assign n3900 = \WX7158_reg/NET0131  & ~\WX7222_reg/NET0131  ;
  assign n3901 = ~\WX7158_reg/NET0131  & \WX7222_reg/NET0131  ;
  assign n3902 = ~n3900 & ~n3901 ;
  assign n3904 = n3899 & ~n3902 ;
  assign n3903 = ~n3899 & n3902 ;
  assign n3905 = ~\TM0_pad  & ~n3903 ;
  assign n3906 = ~n3904 & n3905 ;
  assign n3896 = \TM0_pad  & ~\_2212__reg/NET0131  ;
  assign n3907 = n1976 & ~n3896 ;
  assign n3908 = ~n3906 & n3907 ;
  assign n3909 = ~n3895 & ~n3908 ;
  assign n3910 = n2023 & ~n3745 ;
  assign n3912 = \WX8577_reg/NET0131  & ~\WX8641_reg/NET0131  ;
  assign n3913 = ~\WX8577_reg/NET0131  & \WX8641_reg/NET0131  ;
  assign n3914 = ~n3912 & ~n3913 ;
  assign n3915 = \WX8449_reg/NET0131  & ~\WX8513_reg/NET0131  ;
  assign n3916 = ~\WX8449_reg/NET0131  & \WX8513_reg/NET0131  ;
  assign n3917 = ~n3915 & ~n3916 ;
  assign n3919 = n3914 & ~n3917 ;
  assign n3918 = ~n3914 & n3917 ;
  assign n3920 = ~\TM0_pad  & ~n3918 ;
  assign n3921 = ~n3919 & n3920 ;
  assign n3911 = \TM0_pad  & ~\_2245__reg/NET0131  ;
  assign n3922 = n1976 & ~n3911 ;
  assign n3923 = ~n3921 & n3922 ;
  assign n3924 = ~n3910 & ~n3923 ;
  assign n3925 = ~\TM0_pad  & ~n1646 ;
  assign n3926 = ~n1637 & ~n3925 ;
  assign n3927 = n1973 & ~n3926 ;
  assign n3928 = \TM0_pad  & \_2095__reg/NET0131  ;
  assign n3929 = \WX2092_reg/NET0131  & ~\WX2156_reg/NET0131  ;
  assign n3930 = ~\WX2092_reg/NET0131  & \WX2156_reg/NET0131  ;
  assign n3931 = ~n3929 & ~n3930 ;
  assign n3932 = \WX2028_reg/NET0131  & ~n3931 ;
  assign n3933 = ~\WX2028_reg/NET0131  & n3931 ;
  assign n3934 = ~n3932 & ~n3933 ;
  assign n3935 = \TM1_pad  & ~\WX1964_reg/NET0131  ;
  assign n3936 = ~\TM1_pad  & \WX1964_reg/NET0131  ;
  assign n3937 = ~n3935 & ~n3936 ;
  assign n3939 = n3934 & ~n3937 ;
  assign n3938 = ~n3934 & n3937 ;
  assign n3940 = ~\TM0_pad  & ~n3938 ;
  assign n3941 = ~n3939 & n3940 ;
  assign n3942 = ~n3928 & ~n3941 ;
  assign n3943 = n1976 & ~n3942 ;
  assign n3944 = ~n3927 & ~n3943 ;
  assign n3945 = ~n1682 & ~n2186 ;
  assign n3946 = n1973 & ~n3945 ;
  assign n3948 = \TM0_pad  & ~\_2353__reg/NET0131  ;
  assign n3947 = ~\DATA_0_20_pad  & ~\TM0_pad  ;
  assign n3949 = n1976 & ~n3947 ;
  assign n3950 = ~n3948 & n3949 ;
  assign n3951 = ~n3946 & ~n3950 ;
  assign n3952 = RESET_pad & \WX10849_reg/NET0131  ;
  assign n3953 = ~n1894 & n1973 ;
  assign n3954 = \WX3413_reg/NET0131  & ~\WX3477_reg/NET0131  ;
  assign n3955 = ~\WX3413_reg/NET0131  & \WX3477_reg/NET0131  ;
  assign n3956 = ~n3954 & ~n3955 ;
  assign n3957 = \WX3285_reg/NET0131  & ~\WX3349_reg/NET0131  ;
  assign n3958 = ~\WX3285_reg/NET0131  & \WX3349_reg/NET0131  ;
  assign n3959 = ~n3957 & ~n3958 ;
  assign n3961 = n3956 & ~n3959 ;
  assign n3960 = ~n3956 & n3959 ;
  assign n3962 = ~\TM0_pad  & ~n3960 ;
  assign n3963 = ~n3961 & n3962 ;
  assign n3964 = n3953 & ~n3963 ;
  assign n3966 = \WX4706_reg/NET0131  & ~\WX4770_reg/NET0131  ;
  assign n3967 = ~\WX4706_reg/NET0131  & \WX4770_reg/NET0131  ;
  assign n3968 = ~n3966 & ~n3967 ;
  assign n3969 = \WX4578_reg/NET0131  & ~\WX4642_reg/NET0131  ;
  assign n3970 = ~\WX4578_reg/NET0131  & \WX4642_reg/NET0131  ;
  assign n3971 = ~n3969 & ~n3970 ;
  assign n3973 = n3968 & ~n3971 ;
  assign n3972 = ~n3968 & n3971 ;
  assign n3974 = ~\TM0_pad  & ~n3972 ;
  assign n3975 = ~n3973 & n3974 ;
  assign n3965 = \TM0_pad  & ~\_2145__reg/NET0131  ;
  assign n3976 = n1976 & ~n3965 ;
  assign n3977 = ~n3975 & n3976 ;
  assign n3978 = ~n3964 & ~n3977 ;
  assign n3979 = n2023 & ~n3921 ;
  assign n3981 = \WX9870_reg/NET0131  & ~\WX9934_reg/NET0131  ;
  assign n3982 = ~\WX9870_reg/NET0131  & \WX9934_reg/NET0131  ;
  assign n3983 = ~n3981 & ~n3982 ;
  assign n3984 = \WX9742_reg/NET0131  & ~\WX9806_reg/NET0131  ;
  assign n3985 = ~\WX9742_reg/NET0131  & \WX9806_reg/NET0131  ;
  assign n3986 = ~n3984 & ~n3985 ;
  assign n3988 = n3983 & ~n3986 ;
  assign n3987 = ~n3983 & n3986 ;
  assign n3989 = ~\TM0_pad  & ~n3987 ;
  assign n3990 = ~n3988 & n3989 ;
  assign n3980 = \TM0_pad  & ~\_2277__reg/NET0131  ;
  assign n3991 = n1976 & ~n3980 ;
  assign n3992 = ~n3990 & n3991 ;
  assign n3993 = ~n3979 & ~n3992 ;
  assign n3994 = n3172 & ~n3842 ;
  assign n3996 = \WX11161_reg/NET0131  & ~\WX11225_reg/NET0131  ;
  assign n3997 = ~\WX11161_reg/NET0131  & \WX11225_reg/NET0131  ;
  assign n3998 = ~n3996 & ~n3997 ;
  assign n3999 = \WX11033_reg/NET0131  & ~\WX11097_reg/NET0131  ;
  assign n4000 = ~\WX11033_reg/NET0131  & \WX11097_reg/NET0131  ;
  assign n4001 = ~n3999 & ~n4000 ;
  assign n4003 = n3998 & ~n4001 ;
  assign n4002 = ~n3998 & n4001 ;
  assign n4004 = ~\TM0_pad  & ~n4002 ;
  assign n4005 = ~n4003 & n4004 ;
  assign n3995 = \TM0_pad  & ~\_2310__reg/NET0131  ;
  assign n4006 = n1976 & ~n3995 ;
  assign n4007 = ~n4005 & n4006 ;
  assign n4008 = ~n3994 & ~n4007 ;
  assign n4009 = \TM0_pad  & \_2128__reg/NET0131  ;
  assign n4010 = \WX3383_reg/NET0131  & ~\WX3447_reg/NET0131  ;
  assign n4011 = ~\WX3383_reg/NET0131  & \WX3447_reg/NET0131  ;
  assign n4012 = ~n4010 & ~n4011 ;
  assign n4013 = \WX3319_reg/NET0131  & ~n4012 ;
  assign n4014 = ~\WX3319_reg/NET0131  & n4012 ;
  assign n4015 = ~n4013 & ~n4014 ;
  assign n4016 = \TM1_pad  & ~\WX3255_reg/NET0131  ;
  assign n4017 = ~\TM1_pad  & \WX3255_reg/NET0131  ;
  assign n4018 = ~n4016 & ~n4017 ;
  assign n4020 = n4015 & ~n4018 ;
  assign n4019 = ~n4015 & n4018 ;
  assign n4021 = ~\TM0_pad  & ~n4019 ;
  assign n4022 = ~n4020 & n4021 ;
  assign n4023 = ~n4009 & ~n4022 ;
  assign n4024 = n1976 & ~n4023 ;
  assign n4025 = ~n1653 & ~n3780 ;
  assign n4026 = n1973 & ~n4025 ;
  assign n4027 = ~n4024 & ~n4026 ;
  assign n4028 = n3805 & ~n3827 ;
  assign n4030 = \WX5997_reg/NET0131  & ~\WX6061_reg/NET0131  ;
  assign n4031 = ~\WX5997_reg/NET0131  & \WX6061_reg/NET0131  ;
  assign n4032 = ~n4030 & ~n4031 ;
  assign n4033 = \WX5869_reg/NET0131  & ~\WX5933_reg/NET0131  ;
  assign n4034 = ~\WX5869_reg/NET0131  & \WX5933_reg/NET0131  ;
  assign n4035 = ~n4033 & ~n4034 ;
  assign n4037 = n4032 & ~n4035 ;
  assign n4036 = ~n4032 & n4035 ;
  assign n4038 = ~\TM0_pad  & ~n4036 ;
  assign n4039 = ~n4037 & n4038 ;
  assign n4029 = \TM0_pad  & ~\_2178__reg/NET0131  ;
  assign n4040 = n1976 & ~n4029 ;
  assign n4041 = ~n4039 & n4040 ;
  assign n4042 = ~n4028 & ~n4041 ;
  assign n4043 = n3644 & ~n3891 ;
  assign n4045 = \WX7288_reg/NET0131  & ~\WX7352_reg/NET0131  ;
  assign n4046 = ~\WX7288_reg/NET0131  & \WX7352_reg/NET0131  ;
  assign n4047 = ~n4045 & ~n4046 ;
  assign n4048 = \WX7160_reg/NET0131  & ~\WX7224_reg/NET0131  ;
  assign n4049 = ~\WX7160_reg/NET0131  & \WX7224_reg/NET0131  ;
  assign n4050 = ~n4048 & ~n4049 ;
  assign n4052 = n4047 & ~n4050 ;
  assign n4051 = ~n4047 & n4050 ;
  assign n4053 = ~\TM0_pad  & ~n4051 ;
  assign n4054 = ~n4052 & n4053 ;
  assign n4044 = \TM0_pad  & ~\_2211__reg/NET0131  ;
  assign n4055 = n1976 & ~n4044 ;
  assign n4056 = ~n4054 & n4055 ;
  assign n4057 = ~n4043 & ~n4056 ;
  assign n4058 = n3483 & ~n3906 ;
  assign n4060 = \WX8579_reg/NET0131  & ~\WX8643_reg/NET0131  ;
  assign n4061 = ~\WX8579_reg/NET0131  & \WX8643_reg/NET0131  ;
  assign n4062 = ~n4060 & ~n4061 ;
  assign n4063 = \WX8451_reg/NET0131  & ~\WX8515_reg/NET0131  ;
  assign n4064 = ~\WX8451_reg/NET0131  & \WX8515_reg/NET0131  ;
  assign n4065 = ~n4063 & ~n4064 ;
  assign n4067 = n4062 & ~n4065 ;
  assign n4066 = ~n4062 & n4065 ;
  assign n4068 = ~\TM0_pad  & ~n4066 ;
  assign n4069 = ~n4067 & n4068 ;
  assign n4059 = \TM0_pad  & ~\_2244__reg/NET0131  ;
  assign n4070 = n1976 & ~n4059 ;
  assign n4071 = ~n4069 & n4070 ;
  assign n4072 = ~n4058 & ~n4071 ;
  assign n4073 = \TM0_pad  & \_2094__reg/NET0131  ;
  assign n4074 = \WX2094_reg/NET0131  & ~\WX2158_reg/NET0131  ;
  assign n4075 = ~\WX2094_reg/NET0131  & \WX2158_reg/NET0131  ;
  assign n4076 = ~n4074 & ~n4075 ;
  assign n4077 = \WX2030_reg/NET0131  & ~n4076 ;
  assign n4078 = ~\WX2030_reg/NET0131  & n4076 ;
  assign n4079 = ~n4077 & ~n4078 ;
  assign n4080 = \TM1_pad  & ~\WX1966_reg/NET0131  ;
  assign n4081 = ~\TM1_pad  & \WX1966_reg/NET0131  ;
  assign n4082 = ~n4080 & ~n4081 ;
  assign n4084 = n4079 & ~n4082 ;
  assign n4083 = ~n4079 & n4082 ;
  assign n4085 = ~\TM0_pad  & ~n4083 ;
  assign n4086 = ~n4084 & n4085 ;
  assign n4087 = ~n4073 & ~n4086 ;
  assign n4088 = n1976 & ~n4087 ;
  assign n4089 = ~\TM0_pad  & ~n1630 ;
  assign n4090 = ~n1621 & ~n4089 ;
  assign n4091 = n1973 & ~n4090 ;
  assign n4092 = ~n4088 & ~n4091 ;
  assign n4093 = ~n1653 & ~n2418 ;
  assign n4094 = n1973 & ~n4093 ;
  assign n4096 = \TM0_pad  & ~\_2352__reg/NET0131  ;
  assign n4095 = ~\DATA_0_19_pad  & ~\TM0_pad  ;
  assign n4097 = n1976 & ~n4095 ;
  assign n4098 = ~n4096 & n4097 ;
  assign n4099 = ~n4094 & ~n4098 ;
  assign n4100 = RESET_pad & \WX10851_reg/NET0131  ;
  assign n4101 = ~n1881 & n1973 ;
  assign n4102 = \WX3415_reg/NET0131  & ~\WX3479_reg/NET0131  ;
  assign n4103 = ~\WX3415_reg/NET0131  & \WX3479_reg/NET0131  ;
  assign n4104 = ~n4102 & ~n4103 ;
  assign n4105 = \WX3287_reg/NET0131  & ~\WX3351_reg/NET0131  ;
  assign n4106 = ~\WX3287_reg/NET0131  & \WX3351_reg/NET0131  ;
  assign n4107 = ~n4105 & ~n4106 ;
  assign n4109 = n4104 & ~n4107 ;
  assign n4108 = ~n4104 & n4107 ;
  assign n4110 = ~\TM0_pad  & ~n4108 ;
  assign n4111 = ~n4109 & n4110 ;
  assign n4112 = n4101 & ~n4111 ;
  assign n4114 = \WX4708_reg/NET0131  & ~\WX4772_reg/NET0131  ;
  assign n4115 = ~\WX4708_reg/NET0131  & \WX4772_reg/NET0131  ;
  assign n4116 = ~n4114 & ~n4115 ;
  assign n4117 = \WX4580_reg/NET0131  & ~\WX4644_reg/NET0131  ;
  assign n4118 = ~\WX4580_reg/NET0131  & \WX4644_reg/NET0131  ;
  assign n4119 = ~n4117 & ~n4118 ;
  assign n4121 = n4116 & ~n4119 ;
  assign n4120 = ~n4116 & n4119 ;
  assign n4122 = ~\TM0_pad  & ~n4120 ;
  assign n4123 = ~n4121 & n4122 ;
  assign n4113 = \TM0_pad  & ~\_2144__reg/NET0131  ;
  assign n4124 = n1976 & ~n4113 ;
  assign n4125 = ~n4123 & n4124 ;
  assign n4126 = ~n4112 & ~n4125 ;
  assign n4127 = n3483 & ~n4069 ;
  assign n4129 = \WX9872_reg/NET0131  & ~\WX9936_reg/NET0131  ;
  assign n4130 = ~\WX9872_reg/NET0131  & \WX9936_reg/NET0131  ;
  assign n4131 = ~n4129 & ~n4130 ;
  assign n4132 = \WX9744_reg/NET0131  & ~\WX9808_reg/NET0131  ;
  assign n4133 = ~\WX9744_reg/NET0131  & \WX9808_reg/NET0131  ;
  assign n4134 = ~n4132 & ~n4133 ;
  assign n4136 = n4131 & ~n4134 ;
  assign n4135 = ~n4131 & n4134 ;
  assign n4137 = ~\TM0_pad  & ~n4135 ;
  assign n4138 = ~n4136 & n4137 ;
  assign n4128 = \TM0_pad  & ~\_2276__reg/NET0131  ;
  assign n4139 = n1976 & ~n4128 ;
  assign n4140 = ~n4138 & n4139 ;
  assign n4141 = ~n4127 & ~n4140 ;
  assign n4142 = n2023 & ~n3990 ;
  assign n4143 = \TM0_pad  & ~\_2309__reg/NET0131  ;
  assign n4144 = n1976 & ~n4143 ;
  assign n4145 = ~n2033 & n4144 ;
  assign n4146 = ~n4142 & ~n4145 ;
  assign n4147 = \TM0_pad  & \_2127__reg/NET0131  ;
  assign n4148 = \WX3385_reg/NET0131  & ~\WX3449_reg/NET0131  ;
  assign n4149 = ~\WX3385_reg/NET0131  & \WX3449_reg/NET0131  ;
  assign n4150 = ~n4148 & ~n4149 ;
  assign n4151 = \WX3321_reg/NET0131  & ~n4150 ;
  assign n4152 = ~\WX3321_reg/NET0131  & n4150 ;
  assign n4153 = ~n4151 & ~n4152 ;
  assign n4154 = \TM1_pad  & ~\WX3257_reg/NET0131  ;
  assign n4155 = ~\TM1_pad  & \WX3257_reg/NET0131  ;
  assign n4156 = ~n4154 & ~n4155 ;
  assign n4158 = n4153 & ~n4156 ;
  assign n4157 = ~n4153 & n4156 ;
  assign n4159 = ~\TM0_pad  & ~n4157 ;
  assign n4160 = ~n4158 & n4159 ;
  assign n4161 = ~n4147 & ~n4160 ;
  assign n4162 = n1976 & ~n4161 ;
  assign n4163 = ~n1637 & ~n3941 ;
  assign n4164 = n1973 & ~n4163 ;
  assign n4165 = ~n4162 & ~n4164 ;
  assign n4166 = n3953 & ~n3975 ;
  assign n4168 = \WX5999_reg/NET0131  & ~\WX6063_reg/NET0131  ;
  assign n4169 = ~\WX5999_reg/NET0131  & \WX6063_reg/NET0131  ;
  assign n4170 = ~n4168 & ~n4169 ;
  assign n4171 = \WX5871_reg/NET0131  & ~\WX5935_reg/NET0131  ;
  assign n4172 = ~\WX5871_reg/NET0131  & \WX5935_reg/NET0131  ;
  assign n4173 = ~n4171 & ~n4172 ;
  assign n4175 = n4170 & ~n4173 ;
  assign n4174 = ~n4170 & n4173 ;
  assign n4176 = ~\TM0_pad  & ~n4174 ;
  assign n4177 = ~n4175 & n4176 ;
  assign n4167 = \TM0_pad  & ~\_2177__reg/NET0131  ;
  assign n4178 = n1976 & ~n4167 ;
  assign n4179 = ~n4177 & n4178 ;
  assign n4180 = ~n4166 & ~n4179 ;
  assign n4181 = n3805 & ~n4039 ;
  assign n4183 = \WX7290_reg/NET0131  & ~\WX7354_reg/NET0131  ;
  assign n4184 = ~\WX7290_reg/NET0131  & \WX7354_reg/NET0131  ;
  assign n4185 = ~n4183 & ~n4184 ;
  assign n4186 = \WX7162_reg/NET0131  & ~\WX7226_reg/NET0131  ;
  assign n4187 = ~\WX7162_reg/NET0131  & \WX7226_reg/NET0131  ;
  assign n4188 = ~n4186 & ~n4187 ;
  assign n4190 = n4185 & ~n4188 ;
  assign n4189 = ~n4185 & n4188 ;
  assign n4191 = ~\TM0_pad  & ~n4189 ;
  assign n4192 = ~n4190 & n4191 ;
  assign n4182 = \TM0_pad  & ~\_2210__reg/NET0131  ;
  assign n4193 = n1976 & ~n4182 ;
  assign n4194 = ~n4192 & n4193 ;
  assign n4195 = ~n4181 & ~n4194 ;
  assign n4196 = n3644 & ~n4054 ;
  assign n4198 = \WX8581_reg/NET0131  & ~\WX8645_reg/NET0131  ;
  assign n4199 = ~\WX8581_reg/NET0131  & \WX8645_reg/NET0131  ;
  assign n4200 = ~n4198 & ~n4199 ;
  assign n4201 = \WX8453_reg/NET0131  & ~\WX8517_reg/NET0131  ;
  assign n4202 = ~\WX8453_reg/NET0131  & \WX8517_reg/NET0131  ;
  assign n4203 = ~n4201 & ~n4202 ;
  assign n4205 = n4200 & ~n4203 ;
  assign n4204 = ~n4200 & n4203 ;
  assign n4206 = ~\TM0_pad  & ~n4204 ;
  assign n4207 = ~n4205 & n4206 ;
  assign n4197 = \TM0_pad  & ~\_2243__reg/NET0131  ;
  assign n4208 = n1976 & ~n4197 ;
  assign n4209 = ~n4207 & n4208 ;
  assign n4210 = ~n4196 & ~n4209 ;
  assign n4211 = ~\TM0_pad  & ~n1614 ;
  assign n4212 = ~n1605 & ~n4211 ;
  assign n4213 = n1973 & ~n4212 ;
  assign n4214 = \TM0_pad  & \_2093__reg/NET0131  ;
  assign n4215 = \WX2096_reg/NET0131  & ~\WX2160_reg/NET0131  ;
  assign n4216 = ~\WX2096_reg/NET0131  & \WX2160_reg/NET0131  ;
  assign n4217 = ~n4215 & ~n4216 ;
  assign n4218 = \WX2032_reg/NET0131  & ~n4217 ;
  assign n4219 = ~\WX2032_reg/NET0131  & n4217 ;
  assign n4220 = ~n4218 & ~n4219 ;
  assign n4221 = \TM1_pad  & ~\WX1968_reg/NET0131  ;
  assign n4222 = ~\TM1_pad  & \WX1968_reg/NET0131  ;
  assign n4223 = ~n4221 & ~n4222 ;
  assign n4225 = n4220 & ~n4223 ;
  assign n4224 = ~n4220 & n4223 ;
  assign n4226 = ~\TM0_pad  & ~n4224 ;
  assign n4227 = ~n4225 & n4226 ;
  assign n4228 = ~n4214 & ~n4227 ;
  assign n4229 = n1976 & ~n4228 ;
  assign n4230 = ~n4213 & ~n4229 ;
  assign n4231 = ~n1637 & ~n2594 ;
  assign n4232 = n1973 & ~n4231 ;
  assign n4234 = \TM0_pad  & ~\_2351__reg/NET0131  ;
  assign n4233 = ~\DATA_0_18_pad  & ~\TM0_pad  ;
  assign n4235 = n1976 & ~n4233 ;
  assign n4236 = ~n4234 & n4235 ;
  assign n4237 = ~n4232 & ~n4236 ;
  assign n4238 = RESET_pad & \WX10853_reg/NET0131  ;
  assign n4239 = ~n1836 & n1973 ;
  assign n4240 = \WX3417_reg/NET0131  & ~\WX3481_reg/NET0131  ;
  assign n4241 = ~\WX3417_reg/NET0131  & \WX3481_reg/NET0131  ;
  assign n4242 = ~n4240 & ~n4241 ;
  assign n4243 = \WX3289_reg/NET0131  & ~\WX3353_reg/NET0131  ;
  assign n4244 = ~\WX3289_reg/NET0131  & \WX3353_reg/NET0131  ;
  assign n4245 = ~n4243 & ~n4244 ;
  assign n4247 = n4242 & ~n4245 ;
  assign n4246 = ~n4242 & n4245 ;
  assign n4248 = ~\TM0_pad  & ~n4246 ;
  assign n4249 = ~n4247 & n4248 ;
  assign n4250 = n4239 & ~n4249 ;
  assign n4252 = \WX4710_reg/NET0131  & ~\WX4774_reg/NET0131  ;
  assign n4253 = ~\WX4710_reg/NET0131  & \WX4774_reg/NET0131  ;
  assign n4254 = ~n4252 & ~n4253 ;
  assign n4255 = \WX4582_reg/NET0131  & ~\WX4646_reg/NET0131  ;
  assign n4256 = ~\WX4582_reg/NET0131  & \WX4646_reg/NET0131  ;
  assign n4257 = ~n4255 & ~n4256 ;
  assign n4259 = n4254 & ~n4257 ;
  assign n4258 = ~n4254 & n4257 ;
  assign n4260 = ~\TM0_pad  & ~n4258 ;
  assign n4261 = ~n4259 & n4260 ;
  assign n4251 = \TM0_pad  & ~\_2143__reg/NET0131  ;
  assign n4262 = n1976 & ~n4251 ;
  assign n4263 = ~n4261 & n4262 ;
  assign n4264 = ~n4250 & ~n4263 ;
  assign n4265 = n3644 & ~n4207 ;
  assign n4267 = \WX9874_reg/NET0131  & ~\WX9938_reg/NET0131  ;
  assign n4268 = ~\WX9874_reg/NET0131  & \WX9938_reg/NET0131  ;
  assign n4269 = ~n4267 & ~n4268 ;
  assign n4270 = \WX9746_reg/NET0131  & ~\WX9810_reg/NET0131  ;
  assign n4271 = ~\WX9746_reg/NET0131  & \WX9810_reg/NET0131  ;
  assign n4272 = ~n4270 & ~n4271 ;
  assign n4274 = n4269 & ~n4272 ;
  assign n4273 = ~n4269 & n4272 ;
  assign n4275 = ~\TM0_pad  & ~n4273 ;
  assign n4276 = ~n4274 & n4275 ;
  assign n4266 = \TM0_pad  & ~\_2275__reg/NET0131  ;
  assign n4277 = n1976 & ~n4266 ;
  assign n4278 = ~n4276 & n4277 ;
  assign n4279 = ~n4265 & ~n4278 ;
  assign n4280 = n3483 & ~n4138 ;
  assign n4282 = \WX11165_reg/NET0131  & ~\WX11229_reg/NET0131  ;
  assign n4283 = ~\WX11165_reg/NET0131  & \WX11229_reg/NET0131  ;
  assign n4284 = ~n4282 & ~n4283 ;
  assign n4285 = \WX11037_reg/NET0131  & ~\WX11101_reg/NET0131  ;
  assign n4286 = ~\WX11037_reg/NET0131  & \WX11101_reg/NET0131  ;
  assign n4287 = ~n4285 & ~n4286 ;
  assign n4289 = n4284 & ~n4287 ;
  assign n4288 = ~n4284 & n4287 ;
  assign n4290 = ~\TM0_pad  & ~n4288 ;
  assign n4291 = ~n4289 & n4290 ;
  assign n4281 = \TM0_pad  & ~\_2308__reg/NET0131  ;
  assign n4292 = n1976 & ~n4281 ;
  assign n4293 = ~n4291 & n4292 ;
  assign n4294 = ~n4280 & ~n4293 ;
  assign n4295 = n4101 & ~n4123 ;
  assign n4297 = \WX6001_reg/NET0131  & ~\WX6065_reg/NET0131  ;
  assign n4298 = ~\WX6001_reg/NET0131  & \WX6065_reg/NET0131  ;
  assign n4299 = ~n4297 & ~n4298 ;
  assign n4300 = \WX5873_reg/NET0131  & ~\WX5937_reg/NET0131  ;
  assign n4301 = ~\WX5873_reg/NET0131  & \WX5937_reg/NET0131  ;
  assign n4302 = ~n4300 & ~n4301 ;
  assign n4304 = n4299 & ~n4302 ;
  assign n4303 = ~n4299 & n4302 ;
  assign n4305 = ~\TM0_pad  & ~n4303 ;
  assign n4306 = ~n4304 & n4305 ;
  assign n4296 = \TM0_pad  & ~\_2176__reg/NET0131  ;
  assign n4307 = n1976 & ~n4296 ;
  assign n4308 = ~n4306 & n4307 ;
  assign n4309 = ~n4295 & ~n4308 ;
  assign n4310 = \TM0_pad  & \_2126__reg/NET0131  ;
  assign n4311 = \WX3387_reg/NET0131  & ~\WX3451_reg/NET0131  ;
  assign n4312 = ~\WX3387_reg/NET0131  & \WX3451_reg/NET0131  ;
  assign n4313 = ~n4311 & ~n4312 ;
  assign n4314 = \WX3323_reg/NET0131  & ~n4313 ;
  assign n4315 = ~\WX3323_reg/NET0131  & n4313 ;
  assign n4316 = ~n4314 & ~n4315 ;
  assign n4317 = \TM1_pad  & ~\WX3259_reg/NET0131  ;
  assign n4318 = ~\TM1_pad  & \WX3259_reg/NET0131  ;
  assign n4319 = ~n4317 & ~n4318 ;
  assign n4321 = n4316 & ~n4319 ;
  assign n4320 = ~n4316 & n4319 ;
  assign n4322 = ~\TM0_pad  & ~n4320 ;
  assign n4323 = ~n4321 & n4322 ;
  assign n4324 = ~n4310 & ~n4323 ;
  assign n4325 = n1976 & ~n4324 ;
  assign n4326 = ~n1621 & ~n4086 ;
  assign n4327 = n1973 & ~n4326 ;
  assign n4328 = ~n4325 & ~n4327 ;
  assign n4329 = n3953 & ~n4177 ;
  assign n4331 = \WX7292_reg/NET0131  & ~\WX7356_reg/NET0131  ;
  assign n4332 = ~\WX7292_reg/NET0131  & \WX7356_reg/NET0131  ;
  assign n4333 = ~n4331 & ~n4332 ;
  assign n4334 = \WX7164_reg/NET0131  & ~\WX7228_reg/NET0131  ;
  assign n4335 = ~\WX7164_reg/NET0131  & \WX7228_reg/NET0131  ;
  assign n4336 = ~n4334 & ~n4335 ;
  assign n4338 = n4333 & ~n4336 ;
  assign n4337 = ~n4333 & n4336 ;
  assign n4339 = ~\TM0_pad  & ~n4337 ;
  assign n4340 = ~n4338 & n4339 ;
  assign n4330 = \TM0_pad  & ~\_2209__reg/NET0131  ;
  assign n4341 = n1976 & ~n4330 ;
  assign n4342 = ~n4340 & n4341 ;
  assign n4343 = ~n4329 & ~n4342 ;
  assign n4344 = n3805 & ~n4192 ;
  assign n4346 = \WX8583_reg/NET0131  & ~\WX8647_reg/NET0131  ;
  assign n4347 = ~\WX8583_reg/NET0131  & \WX8647_reg/NET0131  ;
  assign n4348 = ~n4346 & ~n4347 ;
  assign n4349 = \WX8455_reg/NET0131  & ~\WX8519_reg/NET0131  ;
  assign n4350 = ~\WX8455_reg/NET0131  & \WX8519_reg/NET0131  ;
  assign n4351 = ~n4349 & ~n4350 ;
  assign n4353 = n4348 & ~n4351 ;
  assign n4352 = ~n4348 & n4351 ;
  assign n4354 = ~\TM0_pad  & ~n4352 ;
  assign n4355 = ~n4353 & n4354 ;
  assign n4345 = \TM0_pad  & ~\_2242__reg/NET0131  ;
  assign n4356 = n1976 & ~n4345 ;
  assign n4357 = ~n4355 & n4356 ;
  assign n4358 = ~n4344 & ~n4357 ;
  assign n4359 = ~n1621 & ~n2754 ;
  assign n4360 = n1973 & ~n4359 ;
  assign n4362 = \TM0_pad  & ~\_2350__reg/NET0131  ;
  assign n4361 = ~\DATA_0_17_pad  & ~\TM0_pad  ;
  assign n4363 = n1976 & ~n4361 ;
  assign n4364 = ~n4362 & n4363 ;
  assign n4365 = ~n4360 & ~n4364 ;
  assign n4366 = RESET_pad & \WX10855_reg/NET0131  ;
  assign n4367 = n3953 & ~n4340 ;
  assign n4369 = \WX8585_reg/NET0131  & ~\WX8649_reg/NET0131  ;
  assign n4370 = ~\WX8585_reg/NET0131  & \WX8649_reg/NET0131  ;
  assign n4371 = ~n4369 & ~n4370 ;
  assign n4372 = \WX8457_reg/NET0131  & ~\WX8521_reg/NET0131  ;
  assign n4373 = ~\WX8457_reg/NET0131  & \WX8521_reg/NET0131  ;
  assign n4374 = ~n4372 & ~n4373 ;
  assign n4376 = n4371 & ~n4374 ;
  assign n4375 = ~n4371 & n4374 ;
  assign n4377 = ~\TM0_pad  & ~n4375 ;
  assign n4378 = ~n4376 & n4377 ;
  assign n4368 = \TM0_pad  & ~\_2241__reg/NET0131  ;
  assign n4379 = n1976 & ~n4368 ;
  assign n4380 = ~n4378 & n4379 ;
  assign n4381 = ~n4367 & ~n4380 ;
  assign n4382 = ~n1663 & n1973 ;
  assign n4383 = \WX3419_reg/NET0131  & ~\WX3483_reg/NET0131  ;
  assign n4384 = ~\WX3419_reg/NET0131  & \WX3483_reg/NET0131  ;
  assign n4385 = ~n4383 & ~n4384 ;
  assign n4386 = \WX3291_reg/NET0131  & ~\WX3355_reg/NET0131  ;
  assign n4387 = ~\WX3291_reg/NET0131  & \WX3355_reg/NET0131  ;
  assign n4388 = ~n4386 & ~n4387 ;
  assign n4390 = n4385 & ~n4388 ;
  assign n4389 = ~n4385 & n4388 ;
  assign n4391 = ~\TM0_pad  & ~n4389 ;
  assign n4392 = ~n4390 & n4391 ;
  assign n4393 = n4382 & ~n4392 ;
  assign n4395 = \WX4712_reg/NET0131  & ~\WX4776_reg/NET0131  ;
  assign n4396 = ~\WX4712_reg/NET0131  & \WX4776_reg/NET0131  ;
  assign n4397 = ~n4395 & ~n4396 ;
  assign n4398 = \WX4584_reg/NET0131  & ~\WX4648_reg/NET0131  ;
  assign n4399 = ~\WX4584_reg/NET0131  & \WX4648_reg/NET0131  ;
  assign n4400 = ~n4398 & ~n4399 ;
  assign n4402 = n4397 & ~n4400 ;
  assign n4401 = ~n4397 & n4400 ;
  assign n4403 = ~\TM0_pad  & ~n4401 ;
  assign n4404 = ~n4402 & n4403 ;
  assign n4394 = \TM0_pad  & ~\_2142__reg/NET0131  ;
  assign n4405 = n1976 & ~n4394 ;
  assign n4406 = ~n4404 & n4405 ;
  assign n4407 = ~n4393 & ~n4406 ;
  assign n4408 = n3805 & ~n4355 ;
  assign n4410 = \WX9876_reg/NET0131  & ~\WX9940_reg/NET0131  ;
  assign n4411 = ~\WX9876_reg/NET0131  & \WX9940_reg/NET0131  ;
  assign n4412 = ~n4410 & ~n4411 ;
  assign n4413 = \WX9748_reg/NET0131  & ~\WX9812_reg/NET0131  ;
  assign n4414 = ~\WX9748_reg/NET0131  & \WX9812_reg/NET0131  ;
  assign n4415 = ~n4413 & ~n4414 ;
  assign n4417 = n4412 & ~n4415 ;
  assign n4416 = ~n4412 & n4415 ;
  assign n4418 = ~\TM0_pad  & ~n4416 ;
  assign n4419 = ~n4417 & n4418 ;
  assign n4409 = \TM0_pad  & ~\_2274__reg/NET0131  ;
  assign n4420 = n1976 & ~n4409 ;
  assign n4421 = ~n4419 & n4420 ;
  assign n4422 = ~n4408 & ~n4421 ;
  assign n4423 = n3644 & ~n4276 ;
  assign n4425 = \WX11167_reg/NET0131  & ~\WX11231_reg/NET0131  ;
  assign n4426 = ~\WX11167_reg/NET0131  & \WX11231_reg/NET0131  ;
  assign n4427 = ~n4425 & ~n4426 ;
  assign n4428 = \WX11039_reg/NET0131  & ~\WX11103_reg/NET0131  ;
  assign n4429 = ~\WX11039_reg/NET0131  & \WX11103_reg/NET0131  ;
  assign n4430 = ~n4428 & ~n4429 ;
  assign n4432 = n4427 & ~n4430 ;
  assign n4431 = ~n4427 & n4430 ;
  assign n4433 = ~\TM0_pad  & ~n4431 ;
  assign n4434 = ~n4432 & n4433 ;
  assign n4424 = \TM0_pad  & ~\_2307__reg/NET0131  ;
  assign n4435 = n1976 & ~n4424 ;
  assign n4436 = ~n4434 & n4435 ;
  assign n4437 = ~n4423 & ~n4436 ;
  assign n4438 = n4239 & ~n4261 ;
  assign n4440 = \WX6003_reg/NET0131  & ~\WX6067_reg/NET0131  ;
  assign n4441 = ~\WX6003_reg/NET0131  & \WX6067_reg/NET0131  ;
  assign n4442 = ~n4440 & ~n4441 ;
  assign n4443 = \WX5875_reg/NET0131  & ~\WX5939_reg/NET0131  ;
  assign n4444 = ~\WX5875_reg/NET0131  & \WX5939_reg/NET0131  ;
  assign n4445 = ~n4443 & ~n4444 ;
  assign n4447 = n4442 & ~n4445 ;
  assign n4446 = ~n4442 & n4445 ;
  assign n4448 = ~\TM0_pad  & ~n4446 ;
  assign n4449 = ~n4447 & n4448 ;
  assign n4439 = \TM0_pad  & ~\_2175__reg/NET0131  ;
  assign n4450 = n1976 & ~n4439 ;
  assign n4451 = ~n4449 & n4450 ;
  assign n4452 = ~n4438 & ~n4451 ;
  assign n4453 = \TM0_pad  & \_2125__reg/NET0131  ;
  assign n4454 = \WX3389_reg/NET0131  & ~\WX3453_reg/NET0131  ;
  assign n4455 = ~\WX3389_reg/NET0131  & \WX3453_reg/NET0131  ;
  assign n4456 = ~n4454 & ~n4455 ;
  assign n4457 = \WX3325_reg/NET0131  & ~n4456 ;
  assign n4458 = ~\WX3325_reg/NET0131  & n4456 ;
  assign n4459 = ~n4457 & ~n4458 ;
  assign n4460 = \TM1_pad  & ~\WX3261_reg/NET0131  ;
  assign n4461 = ~\TM1_pad  & \WX3261_reg/NET0131  ;
  assign n4462 = ~n4460 & ~n4461 ;
  assign n4464 = n4459 & ~n4462 ;
  assign n4463 = ~n4459 & n4462 ;
  assign n4465 = ~\TM0_pad  & ~n4463 ;
  assign n4466 = ~n4464 & n4465 ;
  assign n4467 = ~n4453 & ~n4466 ;
  assign n4468 = n1976 & ~n4467 ;
  assign n4469 = ~n1605 & ~n4227 ;
  assign n4470 = n1973 & ~n4469 ;
  assign n4471 = ~n4468 & ~n4470 ;
  assign n4472 = n4101 & ~n4306 ;
  assign n4474 = \WX7294_reg/NET0131  & ~\WX7358_reg/NET0131  ;
  assign n4475 = ~\WX7294_reg/NET0131  & \WX7358_reg/NET0131  ;
  assign n4476 = ~n4474 & ~n4475 ;
  assign n4477 = \WX7166_reg/NET0131  & ~\WX7230_reg/NET0131  ;
  assign n4478 = ~\WX7166_reg/NET0131  & \WX7230_reg/NET0131  ;
  assign n4479 = ~n4477 & ~n4478 ;
  assign n4481 = n4476 & ~n4479 ;
  assign n4480 = ~n4476 & n4479 ;
  assign n4482 = ~\TM0_pad  & ~n4480 ;
  assign n4483 = ~n4481 & n4482 ;
  assign n4473 = \TM0_pad  & ~\_2208__reg/NET0131  ;
  assign n4484 = n1976 & ~n4473 ;
  assign n4485 = ~n4483 & n4484 ;
  assign n4486 = ~n4472 & ~n4485 ;
  assign n4487 = ~n1605 & ~n2919 ;
  assign n4488 = n1973 & ~n4487 ;
  assign n4490 = \TM0_pad  & ~\_2349__reg/NET0131  ;
  assign n4489 = ~\DATA_0_16_pad  & ~\TM0_pad  ;
  assign n4491 = n1976 & ~n4489 ;
  assign n4492 = ~n4490 & n4491 ;
  assign n4493 = ~n4488 & ~n4492 ;
  assign n4494 = RESET_pad & \WX10857_reg/NET0131  ;
  assign n4495 = n4101 & ~n4483 ;
  assign n4497 = \WX8587_reg/NET0131  & ~\WX8651_reg/NET0131  ;
  assign n4498 = ~\WX8587_reg/NET0131  & \WX8651_reg/NET0131  ;
  assign n4499 = ~n4497 & ~n4498 ;
  assign n4500 = \WX8459_reg/NET0131  & ~\WX8523_reg/NET0131  ;
  assign n4501 = ~\WX8459_reg/NET0131  & \WX8523_reg/NET0131  ;
  assign n4502 = ~n4500 & ~n4501 ;
  assign n4504 = n4499 & ~n4502 ;
  assign n4503 = ~n4499 & n4502 ;
  assign n4505 = ~\TM0_pad  & ~n4503 ;
  assign n4506 = ~n4504 & n4505 ;
  assign n4496 = \TM0_pad  & ~\_2240__reg/NET0131  ;
  assign n4507 = n1976 & ~n4496 ;
  assign n4508 = ~n4506 & n4507 ;
  assign n4509 = ~n4495 & ~n4508 ;
  assign n4510 = ~n1508 & n1973 ;
  assign n4511 = \WX3421_reg/NET0131  & ~\WX3485_reg/NET0131  ;
  assign n4512 = ~\WX3421_reg/NET0131  & \WX3485_reg/NET0131  ;
  assign n4513 = ~n4511 & ~n4512 ;
  assign n4514 = \WX3293_reg/NET0131  & ~\WX3357_reg/NET0131  ;
  assign n4515 = ~\WX3293_reg/NET0131  & \WX3357_reg/NET0131  ;
  assign n4516 = ~n4514 & ~n4515 ;
  assign n4518 = n4513 & ~n4516 ;
  assign n4517 = ~n4513 & n4516 ;
  assign n4519 = ~\TM0_pad  & ~n4517 ;
  assign n4520 = ~n4518 & n4519 ;
  assign n4521 = n4510 & ~n4520 ;
  assign n4523 = \WX4714_reg/NET0131  & ~\WX4778_reg/NET0131  ;
  assign n4524 = ~\WX4714_reg/NET0131  & \WX4778_reg/NET0131  ;
  assign n4525 = ~n4523 & ~n4524 ;
  assign n4526 = \WX4586_reg/NET0131  & ~\WX4650_reg/NET0131  ;
  assign n4527 = ~\WX4586_reg/NET0131  & \WX4650_reg/NET0131  ;
  assign n4528 = ~n4526 & ~n4527 ;
  assign n4530 = n4525 & ~n4528 ;
  assign n4529 = ~n4525 & n4528 ;
  assign n4531 = ~\TM0_pad  & ~n4529 ;
  assign n4532 = ~n4530 & n4531 ;
  assign n4522 = \TM0_pad  & ~\_2141__reg/NET0131  ;
  assign n4533 = n1976 & ~n4522 ;
  assign n4534 = ~n4532 & n4533 ;
  assign n4535 = ~n4521 & ~n4534 ;
  assign n4536 = n3953 & ~n4378 ;
  assign n4538 = \WX9878_reg/NET0131  & ~\WX9942_reg/NET0131  ;
  assign n4539 = ~\WX9878_reg/NET0131  & \WX9942_reg/NET0131  ;
  assign n4540 = ~n4538 & ~n4539 ;
  assign n4541 = \WX9750_reg/NET0131  & ~\WX9814_reg/NET0131  ;
  assign n4542 = ~\WX9750_reg/NET0131  & \WX9814_reg/NET0131  ;
  assign n4543 = ~n4541 & ~n4542 ;
  assign n4545 = n4540 & ~n4543 ;
  assign n4544 = ~n4540 & n4543 ;
  assign n4546 = ~\TM0_pad  & ~n4544 ;
  assign n4547 = ~n4545 & n4546 ;
  assign n4537 = \TM0_pad  & ~\_2273__reg/NET0131  ;
  assign n4548 = n1976 & ~n4537 ;
  assign n4549 = ~n4547 & n4548 ;
  assign n4550 = ~n4536 & ~n4549 ;
  assign n4551 = n3805 & ~n4419 ;
  assign n4553 = \WX11169_reg/NET0131  & ~\WX11233_reg/NET0131  ;
  assign n4554 = ~\WX11169_reg/NET0131  & \WX11233_reg/NET0131  ;
  assign n4555 = ~n4553 & ~n4554 ;
  assign n4556 = \WX11041_reg/NET0131  & ~\WX11105_reg/NET0131  ;
  assign n4557 = ~\WX11041_reg/NET0131  & \WX11105_reg/NET0131  ;
  assign n4558 = ~n4556 & ~n4557 ;
  assign n4560 = n4555 & ~n4558 ;
  assign n4559 = ~n4555 & n4558 ;
  assign n4561 = ~\TM0_pad  & ~n4559 ;
  assign n4562 = ~n4560 & n4561 ;
  assign n4552 = \TM0_pad  & ~\_2306__reg/NET0131  ;
  assign n4563 = n1976 & ~n4552 ;
  assign n4564 = ~n4562 & n4563 ;
  assign n4565 = ~n4551 & ~n4564 ;
  assign n4566 = n4382 & ~n4404 ;
  assign n4568 = \WX6005_reg/NET0131  & ~\WX6069_reg/NET0131  ;
  assign n4569 = ~\WX6005_reg/NET0131  & \WX6069_reg/NET0131  ;
  assign n4570 = ~n4568 & ~n4569 ;
  assign n4571 = \WX5877_reg/NET0131  & ~\WX5941_reg/NET0131  ;
  assign n4572 = ~\WX5877_reg/NET0131  & \WX5941_reg/NET0131  ;
  assign n4573 = ~n4571 & ~n4572 ;
  assign n4575 = n4570 & ~n4573 ;
  assign n4574 = ~n4570 & n4573 ;
  assign n4576 = ~\TM0_pad  & ~n4574 ;
  assign n4577 = ~n4575 & n4576 ;
  assign n4567 = \TM0_pad  & ~\_2174__reg/NET0131  ;
  assign n4578 = n1976 & ~n4567 ;
  assign n4579 = ~n4577 & n4578 ;
  assign n4580 = ~n4566 & ~n4579 ;
  assign n4581 = n1974 & ~n1987 ;
  assign n4582 = \TM0_pad  & ~\_2124__reg/NET0131  ;
  assign n4583 = n1976 & ~n4582 ;
  assign n4584 = ~n2106 & n4583 ;
  assign n4585 = ~n4581 & ~n4584 ;
  assign n4586 = n4239 & ~n4449 ;
  assign n4588 = \WX7296_reg/NET0131  & ~\WX7360_reg/NET0131  ;
  assign n4589 = ~\WX7296_reg/NET0131  & \WX7360_reg/NET0131  ;
  assign n4590 = ~n4588 & ~n4589 ;
  assign n4591 = \WX7168_reg/NET0131  & ~\WX7232_reg/NET0131  ;
  assign n4592 = ~\WX7168_reg/NET0131  & \WX7232_reg/NET0131  ;
  assign n4593 = ~n4591 & ~n4592 ;
  assign n4595 = n4590 & ~n4593 ;
  assign n4594 = ~n4590 & n4593 ;
  assign n4596 = ~\TM0_pad  & ~n4594 ;
  assign n4597 = ~n4595 & n4596 ;
  assign n4587 = \TM0_pad  & ~\_2207__reg/NET0131  ;
  assign n4598 = n1976 & ~n4587 ;
  assign n4599 = ~n4597 & n4598 ;
  assign n4600 = ~n4586 & ~n4599 ;
  assign n4601 = ~\TM0_pad  & ~n1569 ;
  assign n4602 = n2040 & ~n4601 ;
  assign n4604 = \WX2102_reg/NET0131  & ~\WX2166_reg/NET0131  ;
  assign n4605 = ~\WX2102_reg/NET0131  & \WX2166_reg/NET0131  ;
  assign n4606 = ~n4604 & ~n4605 ;
  assign n4607 = \WX1974_reg/NET0131  & ~\WX2038_reg/NET0131  ;
  assign n4608 = ~\WX1974_reg/NET0131  & \WX2038_reg/NET0131  ;
  assign n4609 = ~n4607 & ~n4608 ;
  assign n4611 = n4606 & ~n4609 ;
  assign n4610 = ~n4606 & n4609 ;
  assign n4612 = ~\TM0_pad  & ~n4610 ;
  assign n4613 = ~n4611 & n4612 ;
  assign n4603 = \TM0_pad  & ~\_2090__reg/NET0131  ;
  assign n4614 = n1976 & ~n4603 ;
  assign n4615 = ~n4613 & n4614 ;
  assign n4616 = ~n4602 & ~n4615 ;
  assign n4617 = RESET_pad & \WX10859_reg/NET0131  ;
  assign n4618 = n4239 & ~n4597 ;
  assign n4620 = \WX8589_reg/NET0131  & ~\WX8653_reg/NET0131  ;
  assign n4621 = ~\WX8589_reg/NET0131  & \WX8653_reg/NET0131  ;
  assign n4622 = ~n4620 & ~n4621 ;
  assign n4623 = \WX8461_reg/NET0131  & ~\WX8525_reg/NET0131  ;
  assign n4624 = ~\WX8461_reg/NET0131  & \WX8525_reg/NET0131  ;
  assign n4625 = ~n4623 & ~n4624 ;
  assign n4627 = n4622 & ~n4625 ;
  assign n4626 = ~n4622 & n4625 ;
  assign n4628 = ~\TM0_pad  & ~n4626 ;
  assign n4629 = ~n4627 & n4628 ;
  assign n4619 = \TM0_pad  & ~\_2239__reg/NET0131  ;
  assign n4630 = n1976 & ~n4619 ;
  assign n4631 = ~n4629 & n4630 ;
  assign n4632 = ~n4618 & ~n4631 ;
  assign n4633 = n4101 & ~n4506 ;
  assign n4635 = \WX9880_reg/NET0131  & ~\WX9944_reg/NET0131  ;
  assign n4636 = ~\WX9880_reg/NET0131  & \WX9944_reg/NET0131  ;
  assign n4637 = ~n4635 & ~n4636 ;
  assign n4638 = \WX9752_reg/NET0131  & ~\WX9816_reg/NET0131  ;
  assign n4639 = ~\WX9752_reg/NET0131  & \WX9816_reg/NET0131  ;
  assign n4640 = ~n4638 & ~n4639 ;
  assign n4642 = n4637 & ~n4640 ;
  assign n4641 = ~n4637 & n4640 ;
  assign n4643 = ~\TM0_pad  & ~n4641 ;
  assign n4644 = ~n4642 & n4643 ;
  assign n4634 = \TM0_pad  & ~\_2272__reg/NET0131  ;
  assign n4645 = n1976 & ~n4634 ;
  assign n4646 = ~n4644 & n4645 ;
  assign n4647 = ~n4633 & ~n4646 ;
  assign n4648 = n3953 & ~n4547 ;
  assign n4650 = \WX11171_reg/NET0131  & ~\WX11235_reg/NET0131  ;
  assign n4651 = ~\WX11171_reg/NET0131  & \WX11235_reg/NET0131  ;
  assign n4652 = ~n4650 & ~n4651 ;
  assign n4653 = \WX11043_reg/NET0131  & ~\WX11107_reg/NET0131  ;
  assign n4654 = ~\WX11043_reg/NET0131  & \WX11107_reg/NET0131  ;
  assign n4655 = ~n4653 & ~n4654 ;
  assign n4657 = n4652 & ~n4655 ;
  assign n4656 = ~n4652 & n4655 ;
  assign n4658 = ~\TM0_pad  & ~n4656 ;
  assign n4659 = ~n4657 & n4658 ;
  assign n4649 = \TM0_pad  & ~\_2305__reg/NET0131  ;
  assign n4660 = n1976 & ~n4649 ;
  assign n4661 = ~n4659 & n4660 ;
  assign n4662 = ~n4648 & ~n4661 ;
  assign n4663 = n4510 & ~n4532 ;
  assign n4665 = \WX6007_reg/NET0131  & ~\WX6071_reg/NET0131  ;
  assign n4666 = ~\WX6007_reg/NET0131  & \WX6071_reg/NET0131  ;
  assign n4667 = ~n4665 & ~n4666 ;
  assign n4668 = \WX5879_reg/NET0131  & ~\WX5943_reg/NET0131  ;
  assign n4669 = ~\WX5879_reg/NET0131  & \WX5943_reg/NET0131  ;
  assign n4670 = ~n4668 & ~n4669 ;
  assign n4672 = n4667 & ~n4670 ;
  assign n4671 = ~n4667 & n4670 ;
  assign n4673 = ~\TM0_pad  & ~n4671 ;
  assign n4674 = ~n4672 & n4673 ;
  assign n4664 = \TM0_pad  & ~\_2173__reg/NET0131  ;
  assign n4675 = n1976 & ~n4664 ;
  assign n4676 = ~n4674 & n4675 ;
  assign n4677 = ~n4663 & ~n4676 ;
  assign n4678 = \WX2100_reg/NET0131  & ~\WX2164_reg/NET0131  ;
  assign n4679 = ~\WX2100_reg/NET0131  & \WX2164_reg/NET0131  ;
  assign n4680 = ~n4678 & ~n4679 ;
  assign n4681 = \WX1972_reg/NET0131  & ~\WX2036_reg/NET0131  ;
  assign n4682 = ~\WX1972_reg/NET0131  & \WX2036_reg/NET0131  ;
  assign n4683 = ~n4681 & ~n4682 ;
  assign n4685 = n4680 & ~n4683 ;
  assign n4684 = ~n4680 & n4683 ;
  assign n4686 = ~\TM0_pad  & ~n4684 ;
  assign n4687 = ~n4685 & n4686 ;
  assign n4688 = n2341 & ~n4687 ;
  assign n4689 = \TM0_pad  & ~\_2123__reg/NET0131  ;
  assign n4690 = n1976 & ~n4689 ;
  assign n4691 = ~n2351 & n4690 ;
  assign n4692 = ~n4688 & ~n4691 ;
  assign n4693 = n4382 & ~n4577 ;
  assign n4695 = \WX7298_reg/NET0131  & ~\WX7362_reg/NET0131  ;
  assign n4696 = ~\WX7298_reg/NET0131  & \WX7362_reg/NET0131  ;
  assign n4697 = ~n4695 & ~n4696 ;
  assign n4698 = \WX7170_reg/NET0131  & ~\WX7234_reg/NET0131  ;
  assign n4699 = ~\WX7170_reg/NET0131  & \WX7234_reg/NET0131  ;
  assign n4700 = ~n4698 & ~n4699 ;
  assign n4702 = n4697 & ~n4700 ;
  assign n4701 = ~n4697 & n4700 ;
  assign n4703 = ~\TM0_pad  & ~n4701 ;
  assign n4704 = ~n4702 & n4703 ;
  assign n4694 = \TM0_pad  & ~\_2206__reg/NET0131  ;
  assign n4705 = n1976 & ~n4694 ;
  assign n4706 = ~n4704 & n4705 ;
  assign n4707 = ~n4693 & ~n4706 ;
  assign n4708 = \TM0_pad  & \_2172__reg/NET0131  ;
  assign n4709 = \WX4652_reg/NET0131  & ~\WX4716_reg/NET0131  ;
  assign n4710 = ~\WX4652_reg/NET0131  & \WX4716_reg/NET0131  ;
  assign n4711 = ~n4709 & ~n4710 ;
  assign n4712 = \WX4588_reg/NET0131  & ~n4711 ;
  assign n4713 = ~\WX4588_reg/NET0131  & n4711 ;
  assign n4714 = ~n4712 & ~n4713 ;
  assign n4715 = \TM1_pad  & ~\WX4524_reg/NET0131  ;
  assign n4716 = ~\TM1_pad  & \WX4524_reg/NET0131  ;
  assign n4717 = ~n4715 & ~n4716 ;
  assign n4719 = n4714 & ~n4717 ;
  assign n4718 = ~n4714 & n4717 ;
  assign n4720 = ~\TM0_pad  & ~n4718 ;
  assign n4721 = ~n4719 & n4720 ;
  assign n4722 = ~n4708 & ~n4721 ;
  assign n4723 = n1976 & ~n4722 ;
  assign n4724 = \WX3359_reg/NET0131  & ~\WX3423_reg/NET0131  ;
  assign n4725 = ~\WX3359_reg/NET0131  & \WX3423_reg/NET0131  ;
  assign n4726 = ~n4724 & ~n4725 ;
  assign n4727 = \WX3295_reg/NET0131  & ~n4726 ;
  assign n4728 = ~\WX3295_reg/NET0131  & n4726 ;
  assign n4729 = ~n4727 & ~n4728 ;
  assign n4730 = \TM1_pad  & ~\WX3231_reg/NET0131  ;
  assign n4731 = ~\TM1_pad  & \WX3231_reg/NET0131  ;
  assign n4732 = ~n4730 & ~n4731 ;
  assign n4734 = n4729 & ~n4732 ;
  assign n4733 = ~n4729 & n4732 ;
  assign n4735 = ~\TM0_pad  & ~n4733 ;
  assign n4736 = ~n4734 & n4735 ;
  assign n4737 = ~n1871 & ~n4736 ;
  assign n4738 = n1973 & ~n4737 ;
  assign n4739 = ~n4723 & ~n4738 ;
  assign n4740 = ~\TM0_pad  & ~n1556 ;
  assign n4741 = n2677 & ~n4740 ;
  assign n4743 = \WX2104_reg/NET0131  & ~\WX2168_reg/NET0131  ;
  assign n4744 = ~\WX2104_reg/NET0131  & \WX2168_reg/NET0131  ;
  assign n4745 = ~n4743 & ~n4744 ;
  assign n4746 = \WX1976_reg/NET0131  & ~\WX2040_reg/NET0131  ;
  assign n4747 = ~\WX1976_reg/NET0131  & \WX2040_reg/NET0131  ;
  assign n4748 = ~n4746 & ~n4747 ;
  assign n4750 = n4745 & ~n4748 ;
  assign n4749 = ~n4745 & n4748 ;
  assign n4751 = ~\TM0_pad  & ~n4749 ;
  assign n4752 = ~n4750 & n4751 ;
  assign n4742 = \TM0_pad  & ~\_2089__reg/NET0131  ;
  assign n4753 = n1976 & ~n4742 ;
  assign n4754 = ~n4752 & n4753 ;
  assign n4755 = ~n4741 & ~n4754 ;
  assign n4756 = n2341 & ~n3224 ;
  assign n4758 = \TM0_pad  & ~\_2347__reg/NET0131  ;
  assign n4757 = ~\DATA_0_14_pad  & ~\TM0_pad  ;
  assign n4759 = n1976 & ~n4757 ;
  assign n4760 = ~n4758 & n4759 ;
  assign n4761 = ~n4756 & ~n4760 ;
  assign n4762 = RESET_pad & \WX10861_reg/NET0131  ;
  assign n4763 = n4382 & ~n4704 ;
  assign n4765 = \WX8591_reg/NET0131  & ~\WX8655_reg/NET0131  ;
  assign n4766 = ~\WX8591_reg/NET0131  & \WX8655_reg/NET0131  ;
  assign n4767 = ~n4765 & ~n4766 ;
  assign n4768 = \WX8463_reg/NET0131  & ~\WX8527_reg/NET0131  ;
  assign n4769 = ~\WX8463_reg/NET0131  & \WX8527_reg/NET0131  ;
  assign n4770 = ~n4768 & ~n4769 ;
  assign n4772 = n4767 & ~n4770 ;
  assign n4771 = ~n4767 & n4770 ;
  assign n4773 = ~\TM0_pad  & ~n4771 ;
  assign n4774 = ~n4772 & n4773 ;
  assign n4764 = \TM0_pad  & ~\_2238__reg/NET0131  ;
  assign n4775 = n1976 & ~n4764 ;
  assign n4776 = ~n4774 & n4775 ;
  assign n4777 = ~n4763 & ~n4776 ;
  assign n4778 = n4239 & ~n4629 ;
  assign n4780 = \WX9882_reg/NET0131  & ~\WX9946_reg/NET0131  ;
  assign n4781 = ~\WX9882_reg/NET0131  & \WX9946_reg/NET0131  ;
  assign n4782 = ~n4780 & ~n4781 ;
  assign n4783 = \WX9754_reg/NET0131  & ~\WX9818_reg/NET0131  ;
  assign n4784 = ~\WX9754_reg/NET0131  & \WX9818_reg/NET0131  ;
  assign n4785 = ~n4783 & ~n4784 ;
  assign n4787 = n4782 & ~n4785 ;
  assign n4786 = ~n4782 & n4785 ;
  assign n4788 = ~\TM0_pad  & ~n4786 ;
  assign n4789 = ~n4787 & n4788 ;
  assign n4779 = \TM0_pad  & ~\_2271__reg/NET0131  ;
  assign n4790 = n1976 & ~n4779 ;
  assign n4791 = ~n4789 & n4790 ;
  assign n4792 = ~n4778 & ~n4791 ;
  assign n4793 = \TM0_pad  & \_2204__reg/NET0131  ;
  assign n4794 = \WX5945_reg/NET0131  & ~\WX6009_reg/NET0131  ;
  assign n4795 = ~\WX5945_reg/NET0131  & \WX6009_reg/NET0131  ;
  assign n4796 = ~n4794 & ~n4795 ;
  assign n4797 = \WX5881_reg/NET0131  & ~n4796 ;
  assign n4798 = ~\WX5881_reg/NET0131  & n4796 ;
  assign n4799 = ~n4797 & ~n4798 ;
  assign n4800 = \TM1_pad  & ~\WX5817_reg/NET0131  ;
  assign n4801 = ~\TM1_pad  & \WX5817_reg/NET0131  ;
  assign n4802 = ~n4800 & ~n4801 ;
  assign n4804 = n4799 & ~n4802 ;
  assign n4803 = ~n4799 & n4802 ;
  assign n4805 = ~\TM0_pad  & ~n4803 ;
  assign n4806 = ~n4804 & n4805 ;
  assign n4807 = ~n4793 & ~n4806 ;
  assign n4808 = n1976 & ~n4807 ;
  assign n4809 = ~n1871 & ~n4721 ;
  assign n4810 = n1973 & ~n4809 ;
  assign n4811 = ~n4808 & ~n4810 ;
  assign n4812 = n4101 & ~n4644 ;
  assign n4814 = \WX11173_reg/NET0131  & ~\WX11237_reg/NET0131  ;
  assign n4815 = ~\WX11173_reg/NET0131  & \WX11237_reg/NET0131  ;
  assign n4816 = ~n4814 & ~n4815 ;
  assign n4817 = \WX11045_reg/NET0131  & ~\WX11109_reg/NET0131  ;
  assign n4818 = ~\WX11045_reg/NET0131  & \WX11109_reg/NET0131  ;
  assign n4819 = ~n4817 & ~n4818 ;
  assign n4821 = n4816 & ~n4819 ;
  assign n4820 = ~n4816 & n4819 ;
  assign n4822 = ~\TM0_pad  & ~n4820 ;
  assign n4823 = ~n4821 & n4822 ;
  assign n4813 = \TM0_pad  & ~\_2304__reg/NET0131  ;
  assign n4824 = n1976 & ~n4813 ;
  assign n4825 = ~n4823 & n4824 ;
  assign n4826 = ~n4812 & ~n4825 ;
  assign n4827 = n2040 & ~n4613 ;
  assign n4828 = \TM0_pad  & ~\_2122__reg/NET0131  ;
  assign n4829 = n1976 & ~n4828 ;
  assign n4830 = ~n2527 & n4829 ;
  assign n4831 = ~n4827 & ~n4830 ;
  assign n4832 = n4510 & ~n4674 ;
  assign n4834 = \WX7300_reg/NET0131  & ~\WX7364_reg/NET0131  ;
  assign n4835 = ~\WX7300_reg/NET0131  & \WX7364_reg/NET0131  ;
  assign n4836 = ~n4834 & ~n4835 ;
  assign n4837 = \WX7172_reg/NET0131  & ~\WX7236_reg/NET0131  ;
  assign n4838 = ~\WX7172_reg/NET0131  & \WX7236_reg/NET0131  ;
  assign n4839 = ~n4837 & ~n4838 ;
  assign n4841 = n4836 & ~n4839 ;
  assign n4840 = ~n4836 & n4839 ;
  assign n4842 = ~\TM0_pad  & ~n4840 ;
  assign n4843 = ~n4841 & n4842 ;
  assign n4833 = \TM0_pad  & ~\_2205__reg/NET0131  ;
  assign n4844 = n1976 & ~n4833 ;
  assign n4845 = ~n4843 & n4844 ;
  assign n4846 = ~n4832 & ~n4845 ;
  assign n4847 = \TM0_pad  & \_2171__reg/NET0131  ;
  assign n4848 = \WX4654_reg/NET0131  & ~\WX4718_reg/NET0131  ;
  assign n4849 = ~\WX4654_reg/NET0131  & \WX4718_reg/NET0131  ;
  assign n4850 = ~n4848 & ~n4849 ;
  assign n4851 = \WX4590_reg/NET0131  & ~n4850 ;
  assign n4852 = ~\WX4590_reg/NET0131  & n4850 ;
  assign n4853 = ~n4851 & ~n4852 ;
  assign n4854 = \TM1_pad  & ~\WX4526_reg/NET0131  ;
  assign n4855 = ~\TM1_pad  & \WX4526_reg/NET0131  ;
  assign n4856 = ~n4854 & ~n4855 ;
  assign n4858 = n4853 & ~n4856 ;
  assign n4857 = ~n4853 & n4856 ;
  assign n4859 = ~\TM0_pad  & ~n4857 ;
  assign n4860 = ~n4858 & n4859 ;
  assign n4861 = ~n4847 & ~n4860 ;
  assign n4862 = n1976 & ~n4861 ;
  assign n4863 = ~n1855 & ~n2135 ;
  assign n4864 = n1973 & ~n4863 ;
  assign n4865 = ~n4862 & ~n4864 ;
  assign n4866 = RESET_pad & \WX10863_reg/NET0131  ;
  assign n4867 = n4510 & ~n4843 ;
  assign n4869 = \WX8593_reg/NET0131  & ~\WX8657_reg/NET0131  ;
  assign n4870 = ~\WX8593_reg/NET0131  & \WX8657_reg/NET0131  ;
  assign n4871 = ~n4869 & ~n4870 ;
  assign n4872 = \WX8465_reg/NET0131  & ~\WX8529_reg/NET0131  ;
  assign n4873 = ~\WX8465_reg/NET0131  & \WX8529_reg/NET0131  ;
  assign n4874 = ~n4872 & ~n4873 ;
  assign n4876 = n4871 & ~n4874 ;
  assign n4875 = ~n4871 & n4874 ;
  assign n4877 = ~\TM0_pad  & ~n4875 ;
  assign n4878 = ~n4876 & n4877 ;
  assign n4868 = \TM0_pad  & ~\_2237__reg/NET0131  ;
  assign n4879 = n1976 & ~n4868 ;
  assign n4880 = ~n4878 & n4879 ;
  assign n4881 = ~n4867 & ~n4880 ;
  assign n4882 = n4382 & ~n4774 ;
  assign n4884 = \WX9884_reg/NET0131  & ~\WX9948_reg/NET0131  ;
  assign n4885 = ~\WX9884_reg/NET0131  & \WX9948_reg/NET0131  ;
  assign n4886 = ~n4884 & ~n4885 ;
  assign n4887 = \WX9756_reg/NET0131  & ~\WX9820_reg/NET0131  ;
  assign n4888 = ~\WX9756_reg/NET0131  & \WX9820_reg/NET0131  ;
  assign n4889 = ~n4887 & ~n4888 ;
  assign n4891 = n4886 & ~n4889 ;
  assign n4890 = ~n4886 & n4889 ;
  assign n4892 = ~\TM0_pad  & ~n4890 ;
  assign n4893 = ~n4891 & n4892 ;
  assign n4883 = \TM0_pad  & ~\_2270__reg/NET0131  ;
  assign n4894 = n1976 & ~n4883 ;
  assign n4895 = ~n4893 & n4894 ;
  assign n4896 = ~n4882 & ~n4895 ;
  assign n4897 = \TM0_pad  & \_2203__reg/NET0131  ;
  assign n4898 = \WX5947_reg/NET0131  & ~\WX6011_reg/NET0131  ;
  assign n4899 = ~\WX5947_reg/NET0131  & \WX6011_reg/NET0131  ;
  assign n4900 = ~n4898 & ~n4899 ;
  assign n4901 = \WX5883_reg/NET0131  & ~n4900 ;
  assign n4902 = ~\WX5883_reg/NET0131  & n4900 ;
  assign n4903 = ~n4901 & ~n4902 ;
  assign n4904 = \TM1_pad  & ~\WX5819_reg/NET0131  ;
  assign n4905 = ~\TM1_pad  & \WX5819_reg/NET0131  ;
  assign n4906 = ~n4904 & ~n4905 ;
  assign n4908 = n4903 & ~n4906 ;
  assign n4907 = ~n4903 & n4906 ;
  assign n4909 = ~\TM0_pad  & ~n4907 ;
  assign n4910 = ~n4908 & n4909 ;
  assign n4911 = ~n4897 & ~n4910 ;
  assign n4912 = n1976 & ~n4911 ;
  assign n4913 = ~n1855 & ~n4860 ;
  assign n4914 = n1973 & ~n4913 ;
  assign n4915 = ~n4912 & ~n4914 ;
  assign n4916 = n4239 & ~n4789 ;
  assign n4918 = \WX11175_reg/NET0131  & ~\WX11239_reg/NET0131  ;
  assign n4919 = ~\WX11175_reg/NET0131  & \WX11239_reg/NET0131  ;
  assign n4920 = ~n4918 & ~n4919 ;
  assign n4921 = \WX11047_reg/NET0131  & ~\WX11111_reg/NET0131  ;
  assign n4922 = ~\WX11047_reg/NET0131  & \WX11111_reg/NET0131  ;
  assign n4923 = ~n4921 & ~n4922 ;
  assign n4925 = n4920 & ~n4923 ;
  assign n4924 = ~n4920 & n4923 ;
  assign n4926 = ~\TM0_pad  & ~n4924 ;
  assign n4927 = ~n4925 & n4926 ;
  assign n4917 = \TM0_pad  & ~\_2303__reg/NET0131  ;
  assign n4928 = n1976 & ~n4917 ;
  assign n4929 = ~n4927 & n4928 ;
  assign n4930 = ~n4916 & ~n4929 ;
  assign n4931 = \TM0_pad  & \_2236__reg/NET0131  ;
  assign n4932 = \WX7238_reg/NET0131  & ~\WX7302_reg/NET0131  ;
  assign n4933 = ~\WX7238_reg/NET0131  & \WX7302_reg/NET0131  ;
  assign n4934 = ~n4932 & ~n4933 ;
  assign n4935 = \WX7174_reg/NET0131  & ~n4934 ;
  assign n4936 = ~\WX7174_reg/NET0131  & n4934 ;
  assign n4937 = ~n4935 & ~n4936 ;
  assign n4938 = \TM1_pad  & ~\WX7110_reg/NET0131  ;
  assign n4939 = ~\TM1_pad  & \WX7110_reg/NET0131  ;
  assign n4940 = ~n4938 & ~n4939 ;
  assign n4942 = n4937 & ~n4940 ;
  assign n4941 = ~n4937 & n4940 ;
  assign n4943 = ~\TM0_pad  & ~n4941 ;
  assign n4944 = ~n4942 & n4943 ;
  assign n4945 = ~n4931 & ~n4944 ;
  assign n4946 = n1976 & ~n4945 ;
  assign n4947 = ~n1871 & ~n4806 ;
  assign n4948 = n1973 & ~n4947 ;
  assign n4949 = ~n4946 & ~n4948 ;
  assign n4950 = n2677 & ~n4752 ;
  assign n4951 = \TM0_pad  & ~\_2121__reg/NET0131  ;
  assign n4952 = n1976 & ~n4951 ;
  assign n4953 = ~n2687 & n4952 ;
  assign n4954 = ~n4950 & ~n4953 ;
  assign n4955 = \TM0_pad  & \_2170__reg/NET0131  ;
  assign n4956 = \WX4656_reg/NET0131  & ~\WX4720_reg/NET0131  ;
  assign n4957 = ~\WX4656_reg/NET0131  & \WX4720_reg/NET0131  ;
  assign n4958 = ~n4956 & ~n4957 ;
  assign n4959 = \WX4592_reg/NET0131  & ~n4958 ;
  assign n4960 = ~\WX4592_reg/NET0131  & n4958 ;
  assign n4961 = ~n4959 & ~n4960 ;
  assign n4962 = \TM1_pad  & ~\WX4528_reg/NET0131  ;
  assign n4963 = ~\TM1_pad  & \WX4528_reg/NET0131  ;
  assign n4964 = ~n4962 & ~n4963 ;
  assign n4966 = n4961 & ~n4964 ;
  assign n4965 = ~n4961 & n4964 ;
  assign n4967 = ~\TM0_pad  & ~n4965 ;
  assign n4968 = ~n4966 & n4967 ;
  assign n4969 = ~n4955 & ~n4968 ;
  assign n4970 = n1976 & ~n4969 ;
  assign n4971 = ~n1826 & ~n2399 ;
  assign n4972 = n1973 & ~n4971 ;
  assign n4973 = ~n4970 & ~n4972 ;
  assign n4974 = ~\TM0_pad  & ~n1530 ;
  assign n4975 = n3011 & ~n4974 ;
  assign n4977 = \WX2108_reg/NET0131  & ~\WX2172_reg/NET0131  ;
  assign n4978 = ~\WX2108_reg/NET0131  & \WX2172_reg/NET0131  ;
  assign n4979 = ~n4977 & ~n4978 ;
  assign n4980 = \WX1980_reg/NET0131  & ~\WX2044_reg/NET0131  ;
  assign n4981 = ~\WX1980_reg/NET0131  & \WX2044_reg/NET0131  ;
  assign n4982 = ~n4980 & ~n4981 ;
  assign n4984 = n4979 & ~n4982 ;
  assign n4983 = ~n4979 & n4982 ;
  assign n4985 = ~\TM0_pad  & ~n4983 ;
  assign n4986 = ~n4984 & n4985 ;
  assign n4976 = \TM0_pad  & ~\_2087__reg/NET0131  ;
  assign n4987 = n1976 & ~n4976 ;
  assign n4988 = ~n4986 & n4987 ;
  assign n4989 = ~n4975 & ~n4988 ;
  assign n4990 = n2677 & ~n3535 ;
  assign n4992 = \TM0_pad  & ~\_2345__reg/NET0131  ;
  assign n4991 = ~\DATA_0_12_pad  & ~\TM0_pad  ;
  assign n4993 = n1976 & ~n4991 ;
  assign n4994 = ~n4992 & n4993 ;
  assign n4995 = ~n4990 & ~n4994 ;
  assign n4996 = RESET_pad & \WX10865_reg/NET0131  ;
  assign n4997 = n4510 & ~n4878 ;
  assign n4999 = \WX9886_reg/NET0131  & ~\WX9950_reg/NET0131  ;
  assign n5000 = ~\WX9886_reg/NET0131  & \WX9950_reg/NET0131  ;
  assign n5001 = ~n4999 & ~n5000 ;
  assign n5002 = \WX9758_reg/NET0131  & ~\WX9822_reg/NET0131  ;
  assign n5003 = ~\WX9758_reg/NET0131  & \WX9822_reg/NET0131  ;
  assign n5004 = ~n5002 & ~n5003 ;
  assign n5006 = n5001 & ~n5004 ;
  assign n5005 = ~n5001 & n5004 ;
  assign n5007 = ~\TM0_pad  & ~n5005 ;
  assign n5008 = ~n5006 & n5007 ;
  assign n4998 = \TM0_pad  & ~\_2269__reg/NET0131  ;
  assign n5009 = n1976 & ~n4998 ;
  assign n5010 = ~n5008 & n5009 ;
  assign n5011 = ~n4997 & ~n5010 ;
  assign n5012 = \TM0_pad  & \_2202__reg/NET0131  ;
  assign n5013 = \WX5949_reg/NET0131  & ~\WX6013_reg/NET0131  ;
  assign n5014 = ~\WX5949_reg/NET0131  & \WX6013_reg/NET0131  ;
  assign n5015 = ~n5013 & ~n5014 ;
  assign n5016 = \WX5885_reg/NET0131  & ~n5015 ;
  assign n5017 = ~\WX5885_reg/NET0131  & n5015 ;
  assign n5018 = ~n5016 & ~n5017 ;
  assign n5019 = \TM1_pad  & ~\WX5821_reg/NET0131  ;
  assign n5020 = ~\TM1_pad  & \WX5821_reg/NET0131  ;
  assign n5021 = ~n5019 & ~n5020 ;
  assign n5023 = n5018 & ~n5021 ;
  assign n5022 = ~n5018 & n5021 ;
  assign n5024 = ~\TM0_pad  & ~n5022 ;
  assign n5025 = ~n5023 & n5024 ;
  assign n5026 = ~n5012 & ~n5025 ;
  assign n5027 = n1976 & ~n5026 ;
  assign n5028 = ~n1826 & ~n4968 ;
  assign n5029 = n1973 & ~n5028 ;
  assign n5030 = ~n5027 & ~n5029 ;
  assign n5031 = n4382 & ~n4893 ;
  assign n5033 = \WX11177_reg/NET0131  & ~\WX11241_reg/NET0131  ;
  assign n5034 = ~\WX11177_reg/NET0131  & \WX11241_reg/NET0131  ;
  assign n5035 = ~n5033 & ~n5034 ;
  assign n5036 = \WX11049_reg/NET0131  & ~\WX11113_reg/NET0131  ;
  assign n5037 = ~\WX11049_reg/NET0131  & \WX11113_reg/NET0131  ;
  assign n5038 = ~n5036 & ~n5037 ;
  assign n5040 = n5035 & ~n5038 ;
  assign n5039 = ~n5035 & n5038 ;
  assign n5041 = ~\TM0_pad  & ~n5039 ;
  assign n5042 = ~n5040 & n5041 ;
  assign n5032 = \TM0_pad  & ~\_2302__reg/NET0131  ;
  assign n5043 = n1976 & ~n5032 ;
  assign n5044 = ~n5042 & n5043 ;
  assign n5045 = ~n5031 & ~n5044 ;
  assign n5046 = \TM0_pad  & \_2235__reg/NET0131  ;
  assign n5047 = \TM1_pad  & ~\WX7112_reg/NET0131  ;
  assign n5048 = ~\TM1_pad  & \WX7112_reg/NET0131  ;
  assign n5049 = ~n5047 & ~n5048 ;
  assign n5050 = ~\WX7176_reg/NET0131  & ~n5049 ;
  assign n5051 = \WX7176_reg/NET0131  & n5049 ;
  assign n5052 = ~n5050 & ~n5051 ;
  assign n5053 = \WX7240_reg/NET0131  & ~\WX7304_reg/NET0131  ;
  assign n5054 = ~\WX7240_reg/NET0131  & \WX7304_reg/NET0131  ;
  assign n5055 = ~n5053 & ~n5054 ;
  assign n5057 = n5052 & n5055 ;
  assign n5056 = ~n5052 & ~n5055 ;
  assign n5058 = ~\TM0_pad  & ~n5056 ;
  assign n5059 = ~n5057 & n5058 ;
  assign n5060 = ~n5046 & ~n5059 ;
  assign n5061 = n1976 & ~n5060 ;
  assign n5062 = ~n1855 & ~n4910 ;
  assign n5063 = n1973 & ~n5062 ;
  assign n5064 = ~n5061 & ~n5063 ;
  assign n5065 = \WX2106_reg/NET0131  & ~\WX2170_reg/NET0131  ;
  assign n5066 = ~\WX2106_reg/NET0131  & \WX2170_reg/NET0131  ;
  assign n5067 = ~n5065 & ~n5066 ;
  assign n5068 = \WX1978_reg/NET0131  & ~\WX2042_reg/NET0131  ;
  assign n5069 = ~\WX1978_reg/NET0131  & \WX2042_reg/NET0131  ;
  assign n5070 = ~n5068 & ~n5069 ;
  assign n5072 = n5067 & ~n5070 ;
  assign n5071 = ~n5067 & n5070 ;
  assign n5073 = ~\TM0_pad  & ~n5071 ;
  assign n5074 = ~n5072 & n5073 ;
  assign n5075 = n2846 & ~n5074 ;
  assign n5076 = \TM0_pad  & ~\_2120__reg/NET0131  ;
  assign n5077 = n1976 & ~n5076 ;
  assign n5078 = ~n2856 & n5077 ;
  assign n5079 = ~n5075 & ~n5078 ;
  assign n5080 = \TM0_pad  & \_2268__reg/NET0131  ;
  assign n5081 = \WX8531_reg/NET0131  & ~\WX8595_reg/NET0131  ;
  assign n5082 = ~\WX8531_reg/NET0131  & \WX8595_reg/NET0131  ;
  assign n5083 = ~n5081 & ~n5082 ;
  assign n5084 = \WX8467_reg/NET0131  & ~n5083 ;
  assign n5085 = ~\WX8467_reg/NET0131  & n5083 ;
  assign n5086 = ~n5084 & ~n5085 ;
  assign n5087 = \TM1_pad  & ~\WX8403_reg/NET0131  ;
  assign n5088 = ~\TM1_pad  & \WX8403_reg/NET0131  ;
  assign n5089 = ~n5087 & ~n5088 ;
  assign n5091 = n5086 & ~n5089 ;
  assign n5090 = ~n5086 & n5089 ;
  assign n5092 = ~\TM0_pad  & ~n5090 ;
  assign n5093 = ~n5091 & n5092 ;
  assign n5094 = ~n5080 & ~n5093 ;
  assign n5095 = n1976 & ~n5094 ;
  assign n5096 = ~n1871 & ~n4944 ;
  assign n5097 = n1973 & ~n5096 ;
  assign n5098 = ~n5095 & ~n5097 ;
  assign n5099 = \TM0_pad  & \_2169__reg/NET0131  ;
  assign n5100 = \WX4658_reg/NET0131  & ~\WX4722_reg/NET0131  ;
  assign n5101 = ~\WX4658_reg/NET0131  & \WX4722_reg/NET0131  ;
  assign n5102 = ~n5100 & ~n5101 ;
  assign n5103 = \WX4594_reg/NET0131  & ~n5102 ;
  assign n5104 = ~\WX4594_reg/NET0131  & n5102 ;
  assign n5105 = ~n5103 & ~n5104 ;
  assign n5106 = \TM1_pad  & ~\WX4530_reg/NET0131  ;
  assign n5107 = ~\TM1_pad  & \WX4530_reg/NET0131  ;
  assign n5108 = ~n5106 & ~n5107 ;
  assign n5110 = n5105 & ~n5108 ;
  assign n5109 = ~n5105 & n5108 ;
  assign n5111 = ~\TM0_pad  & ~n5109 ;
  assign n5112 = ~n5110 & n5111 ;
  assign n5113 = ~n5099 & ~n5112 ;
  assign n5114 = n1976 & ~n5113 ;
  assign n5115 = ~n1810 & ~n2575 ;
  assign n5116 = n1973 & ~n5115 ;
  assign n5117 = ~n5114 & ~n5116 ;
  assign n5118 = n2846 & ~n3696 ;
  assign n5120 = \TM0_pad  & ~\_2344__reg/NET0131  ;
  assign n5119 = ~\DATA_0_11_pad  & ~\TM0_pad  ;
  assign n5121 = n1976 & ~n5119 ;
  assign n5122 = ~n5120 & n5121 ;
  assign n5123 = ~n5118 & ~n5122 ;
  assign n5124 = RESET_pad & \WX10867_reg/NET0131  ;
  assign n5125 = \TM0_pad  & \_2300__reg/NET0131  ;
  assign n5126 = \WX9824_reg/NET0131  & ~\WX9888_reg/NET0131  ;
  assign n5127 = ~\WX9824_reg/NET0131  & \WX9888_reg/NET0131  ;
  assign n5128 = ~n5126 & ~n5127 ;
  assign n5129 = \WX9760_reg/NET0131  & ~n5128 ;
  assign n5130 = ~\WX9760_reg/NET0131  & n5128 ;
  assign n5131 = ~n5129 & ~n5130 ;
  assign n5132 = \TM1_pad  & ~\WX9696_reg/NET0131  ;
  assign n5133 = ~\TM1_pad  & \WX9696_reg/NET0131  ;
  assign n5134 = ~n5132 & ~n5133 ;
  assign n5136 = n5131 & ~n5134 ;
  assign n5135 = ~n5131 & n5134 ;
  assign n5137 = ~\TM0_pad  & ~n5135 ;
  assign n5138 = ~n5136 & n5137 ;
  assign n5139 = ~n5125 & ~n5138 ;
  assign n5140 = n1976 & ~n5139 ;
  assign n5141 = ~n1871 & ~n5093 ;
  assign n5142 = n1973 & ~n5141 ;
  assign n5143 = ~n5140 & ~n5142 ;
  assign n5144 = \TM0_pad  & \_2201__reg/NET0131  ;
  assign n5145 = \WX5951_reg/NET0131  & ~\WX6015_reg/NET0131  ;
  assign n5146 = ~\WX5951_reg/NET0131  & \WX6015_reg/NET0131  ;
  assign n5147 = ~n5145 & ~n5146 ;
  assign n5148 = \WX5887_reg/NET0131  & ~n5147 ;
  assign n5149 = ~\WX5887_reg/NET0131  & n5147 ;
  assign n5150 = ~n5148 & ~n5149 ;
  assign n5151 = \TM1_pad  & ~\WX5823_reg/NET0131  ;
  assign n5152 = ~\TM1_pad  & \WX5823_reg/NET0131  ;
  assign n5153 = ~n5151 & ~n5152 ;
  assign n5155 = n5150 & ~n5153 ;
  assign n5154 = ~n5150 & n5153 ;
  assign n5156 = ~\TM0_pad  & ~n5154 ;
  assign n5157 = ~n5155 & n5156 ;
  assign n5158 = ~n5144 & ~n5157 ;
  assign n5159 = n1976 & ~n5158 ;
  assign n5160 = ~n1810 & ~n5112 ;
  assign n5161 = n1973 & ~n5160 ;
  assign n5162 = ~n5159 & ~n5161 ;
  assign n5163 = n4510 & ~n5008 ;
  assign n5165 = \WX11179_reg/NET0131  & ~\WX11243_reg/NET0131  ;
  assign n5166 = ~\WX11179_reg/NET0131  & \WX11243_reg/NET0131  ;
  assign n5167 = ~n5165 & ~n5166 ;
  assign n5168 = \WX11051_reg/NET0131  & ~\WX11115_reg/NET0131  ;
  assign n5169 = ~\WX11051_reg/NET0131  & \WX11115_reg/NET0131  ;
  assign n5170 = ~n5168 & ~n5169 ;
  assign n5172 = n5167 & ~n5170 ;
  assign n5171 = ~n5167 & n5170 ;
  assign n5173 = ~\TM0_pad  & ~n5171 ;
  assign n5174 = ~n5172 & n5173 ;
  assign n5164 = \TM0_pad  & ~\_2301__reg/NET0131  ;
  assign n5175 = n1976 & ~n5164 ;
  assign n5176 = ~n5174 & n5175 ;
  assign n5177 = ~n5163 & ~n5176 ;
  assign n5178 = \TM0_pad  & \_2234__reg/NET0131  ;
  assign n5179 = \WX7242_reg/NET0131  & ~\WX7306_reg/NET0131  ;
  assign n5180 = ~\WX7242_reg/NET0131  & \WX7306_reg/NET0131  ;
  assign n5181 = ~n5179 & ~n5180 ;
  assign n5182 = \WX7178_reg/NET0131  & ~n5181 ;
  assign n5183 = ~\WX7178_reg/NET0131  & n5181 ;
  assign n5184 = ~n5182 & ~n5183 ;
  assign n5185 = \TM1_pad  & ~\WX7114_reg/NET0131  ;
  assign n5186 = ~\TM1_pad  & \WX7114_reg/NET0131  ;
  assign n5187 = ~n5185 & ~n5186 ;
  assign n5189 = n5184 & ~n5187 ;
  assign n5188 = ~n5184 & n5187 ;
  assign n5190 = ~\TM0_pad  & ~n5188 ;
  assign n5191 = ~n5189 & n5190 ;
  assign n5192 = ~n5178 & ~n5191 ;
  assign n5193 = n1976 & ~n5192 ;
  assign n5194 = ~n1826 & ~n5025 ;
  assign n5195 = n1973 & ~n5194 ;
  assign n5196 = ~n5193 & ~n5195 ;
  assign n5197 = n3011 & ~n4986 ;
  assign n5198 = \TM0_pad  & ~\_2119__reg/NET0131  ;
  assign n5199 = n1976 & ~n5198 ;
  assign n5200 = ~n3021 & n5199 ;
  assign n5201 = ~n5197 & ~n5200 ;
  assign n5202 = \TM0_pad  & \_2267__reg/NET0131  ;
  assign n5203 = \WX8533_reg/NET0131  & ~\WX8597_reg/NET0131  ;
  assign n5204 = ~\WX8533_reg/NET0131  & \WX8597_reg/NET0131  ;
  assign n5205 = ~n5203 & ~n5204 ;
  assign n5206 = \WX8469_reg/NET0131  & ~n5205 ;
  assign n5207 = ~\WX8469_reg/NET0131  & n5205 ;
  assign n5208 = ~n5206 & ~n5207 ;
  assign n5209 = \TM1_pad  & ~\WX8405_reg/NET0131  ;
  assign n5210 = ~\TM1_pad  & \WX8405_reg/NET0131  ;
  assign n5211 = ~n5209 & ~n5210 ;
  assign n5213 = n5208 & ~n5211 ;
  assign n5212 = ~n5208 & n5211 ;
  assign n5214 = ~\TM0_pad  & ~n5212 ;
  assign n5215 = ~n5213 & n5214 ;
  assign n5216 = ~n5202 & ~n5215 ;
  assign n5217 = n1976 & ~n5216 ;
  assign n5218 = ~n1855 & ~n5059 ;
  assign n5219 = n1973 & ~n5218 ;
  assign n5220 = ~n5217 & ~n5219 ;
  assign n5221 = \TM0_pad  & \_2168__reg/NET0131  ;
  assign n5222 = \WX4660_reg/NET0131  & ~\WX4724_reg/NET0131  ;
  assign n5223 = ~\WX4660_reg/NET0131  & \WX4724_reg/NET0131  ;
  assign n5224 = ~n5222 & ~n5223 ;
  assign n5225 = \WX4596_reg/NET0131  & ~n5224 ;
  assign n5226 = ~\WX4596_reg/NET0131  & n5224 ;
  assign n5227 = ~n5225 & ~n5226 ;
  assign n5228 = \TM1_pad  & ~\WX4532_reg/NET0131  ;
  assign n5229 = ~\TM1_pad  & \WX4532_reg/NET0131  ;
  assign n5230 = ~n5228 & ~n5229 ;
  assign n5232 = n5227 & ~n5230 ;
  assign n5231 = ~n5227 & n5230 ;
  assign n5233 = ~\TM0_pad  & ~n5231 ;
  assign n5234 = ~n5232 & n5233 ;
  assign n5235 = ~n5221 & ~n5234 ;
  assign n5236 = n1976 & ~n5235 ;
  assign n5237 = ~n1794 & ~n2735 ;
  assign n5238 = n1973 & ~n5237 ;
  assign n5239 = ~n5236 & ~n5238 ;
  assign n5240 = n3011 & ~n3857 ;
  assign n5242 = \TM0_pad  & ~\_2343__reg/NET0131  ;
  assign n5241 = ~\DATA_0_10_pad  & ~\TM0_pad  ;
  assign n5243 = n1976 & ~n5241 ;
  assign n5244 = ~n5242 & n5243 ;
  assign n5245 = ~n5240 & ~n5244 ;
  assign n5246 = RESET_pad & \WX10869_reg/NET0131  ;
  assign n5247 = \TM0_pad  & \_2299__reg/NET0131  ;
  assign n5248 = \WX9826_reg/NET0131  & ~\WX9890_reg/NET0131  ;
  assign n5249 = ~\WX9826_reg/NET0131  & \WX9890_reg/NET0131  ;
  assign n5250 = ~n5248 & ~n5249 ;
  assign n5251 = \WX9762_reg/NET0131  & ~n5250 ;
  assign n5252 = ~\WX9762_reg/NET0131  & n5250 ;
  assign n5253 = ~n5251 & ~n5252 ;
  assign n5254 = \TM1_pad  & ~\WX9698_reg/NET0131  ;
  assign n5255 = ~\TM1_pad  & \WX9698_reg/NET0131  ;
  assign n5256 = ~n5254 & ~n5255 ;
  assign n5258 = n5253 & ~n5256 ;
  assign n5257 = ~n5253 & n5256 ;
  assign n5259 = ~\TM0_pad  & ~n5257 ;
  assign n5260 = ~n5258 & n5259 ;
  assign n5261 = ~n5247 & ~n5260 ;
  assign n5262 = n1976 & ~n5261 ;
  assign n5263 = ~n1855 & ~n5215 ;
  assign n5264 = n1973 & ~n5263 ;
  assign n5265 = ~n5262 & ~n5264 ;
  assign n5266 = \TM0_pad  & \_2332__reg/NET0131  ;
  assign n5267 = \TM1_pad  & ~\WX10989_reg/NET0131  ;
  assign n5268 = ~\TM1_pad  & \WX10989_reg/NET0131  ;
  assign n5269 = ~n5267 & ~n5268 ;
  assign n5270 = ~\WX11053_reg/NET0131  & ~n5269 ;
  assign n5271 = \WX11053_reg/NET0131  & n5269 ;
  assign n5272 = ~n5270 & ~n5271 ;
  assign n5273 = \WX11117_reg/NET0131  & ~\WX11181_reg/NET0131  ;
  assign n5274 = ~\WX11117_reg/NET0131  & \WX11181_reg/NET0131  ;
  assign n5275 = ~n5273 & ~n5274 ;
  assign n5277 = ~n5272 & ~n5275 ;
  assign n5276 = n5272 & n5275 ;
  assign n5278 = ~\TM0_pad  & ~n5276 ;
  assign n5279 = ~n5277 & n5278 ;
  assign n5280 = ~n5266 & ~n5279 ;
  assign n5281 = n1976 & ~n5280 ;
  assign n5282 = ~n1871 & ~n5138 ;
  assign n5283 = n1973 & ~n5282 ;
  assign n5284 = ~n5281 & ~n5283 ;
  assign n5285 = \TM0_pad  & \_2200__reg/NET0131  ;
  assign n5286 = \WX5953_reg/NET0131  & ~\WX6017_reg/NET0131  ;
  assign n5287 = ~\WX5953_reg/NET0131  & \WX6017_reg/NET0131  ;
  assign n5288 = ~n5286 & ~n5287 ;
  assign n5289 = \WX5889_reg/NET0131  & ~n5288 ;
  assign n5290 = ~\WX5889_reg/NET0131  & n5288 ;
  assign n5291 = ~n5289 & ~n5290 ;
  assign n5292 = \TM1_pad  & ~\WX5825_reg/NET0131  ;
  assign n5293 = ~\TM1_pad  & \WX5825_reg/NET0131  ;
  assign n5294 = ~n5292 & ~n5293 ;
  assign n5296 = n5291 & ~n5294 ;
  assign n5295 = ~n5291 & n5294 ;
  assign n5297 = ~\TM0_pad  & ~n5295 ;
  assign n5298 = ~n5296 & n5297 ;
  assign n5299 = ~n5285 & ~n5298 ;
  assign n5300 = n1976 & ~n5299 ;
  assign n5301 = ~n1794 & ~n5234 ;
  assign n5302 = n1973 & ~n5301 ;
  assign n5303 = ~n5300 & ~n5302 ;
  assign n5304 = \TM0_pad  & \_2233__reg/NET0131  ;
  assign n5305 = \WX7244_reg/NET0131  & ~\WX7308_reg/NET0131  ;
  assign n5306 = ~\WX7244_reg/NET0131  & \WX7308_reg/NET0131  ;
  assign n5307 = ~n5305 & ~n5306 ;
  assign n5308 = \WX7180_reg/NET0131  & ~n5307 ;
  assign n5309 = ~\WX7180_reg/NET0131  & n5307 ;
  assign n5310 = ~n5308 & ~n5309 ;
  assign n5311 = \TM1_pad  & ~\WX7116_reg/NET0131  ;
  assign n5312 = ~\TM1_pad  & \WX7116_reg/NET0131  ;
  assign n5313 = ~n5311 & ~n5312 ;
  assign n5315 = n5310 & ~n5313 ;
  assign n5314 = ~n5310 & n5313 ;
  assign n5316 = ~\TM0_pad  & ~n5314 ;
  assign n5317 = ~n5315 & n5316 ;
  assign n5318 = ~n5304 & ~n5317 ;
  assign n5319 = n1976 & ~n5318 ;
  assign n5320 = ~n1810 & ~n5157 ;
  assign n5321 = n1973 & ~n5320 ;
  assign n5322 = ~n5319 & ~n5321 ;
  assign n5323 = \WX2110_reg/NET0131  & ~\WX2174_reg/NET0131  ;
  assign n5324 = ~\WX2110_reg/NET0131  & \WX2174_reg/NET0131  ;
  assign n5325 = ~n5323 & ~n5324 ;
  assign n5326 = \WX1982_reg/NET0131  & ~\WX2046_reg/NET0131  ;
  assign n5327 = ~\WX1982_reg/NET0131  & \WX2046_reg/NET0131  ;
  assign n5328 = ~n5326 & ~n5327 ;
  assign n5330 = n5325 & ~n5328 ;
  assign n5329 = ~n5325 & n5328 ;
  assign n5331 = ~\TM0_pad  & ~n5329 ;
  assign n5332 = ~n5330 & n5331 ;
  assign n5333 = n3172 & ~n5332 ;
  assign n5334 = \TM0_pad  & ~\_2118__reg/NET0131  ;
  assign n5335 = n1976 & ~n5334 ;
  assign n5336 = ~n3182 & n5335 ;
  assign n5337 = ~n5333 & ~n5336 ;
  assign n5338 = \TM0_pad  & \_2266__reg/NET0131  ;
  assign n5339 = \WX8535_reg/NET0131  & ~\WX8599_reg/NET0131  ;
  assign n5340 = ~\WX8535_reg/NET0131  & \WX8599_reg/NET0131  ;
  assign n5341 = ~n5339 & ~n5340 ;
  assign n5342 = \WX8471_reg/NET0131  & ~n5341 ;
  assign n5343 = ~\WX8471_reg/NET0131  & n5341 ;
  assign n5344 = ~n5342 & ~n5343 ;
  assign n5345 = \TM1_pad  & ~\WX8407_reg/NET0131  ;
  assign n5346 = ~\TM1_pad  & \WX8407_reg/NET0131  ;
  assign n5347 = ~n5345 & ~n5346 ;
  assign n5349 = n5344 & ~n5347 ;
  assign n5348 = ~n5344 & n5347 ;
  assign n5350 = ~\TM0_pad  & ~n5348 ;
  assign n5351 = ~n5349 & n5350 ;
  assign n5352 = ~n5338 & ~n5351 ;
  assign n5353 = n1976 & ~n5352 ;
  assign n5354 = ~n1826 & ~n5191 ;
  assign n5355 = n1973 & ~n5354 ;
  assign n5356 = ~n5353 & ~n5355 ;
  assign n5357 = \TM0_pad  & \_2167__reg/NET0131  ;
  assign n5358 = \WX4662_reg/NET0131  & ~\WX4726_reg/NET0131  ;
  assign n5359 = ~\WX4662_reg/NET0131  & \WX4726_reg/NET0131  ;
  assign n5360 = ~n5358 & ~n5359 ;
  assign n5361 = \WX4598_reg/NET0131  & ~n5360 ;
  assign n5362 = ~\WX4598_reg/NET0131  & n5360 ;
  assign n5363 = ~n5361 & ~n5362 ;
  assign n5364 = \TM1_pad  & ~\WX4534_reg/NET0131  ;
  assign n5365 = ~\TM1_pad  & \WX4534_reg/NET0131  ;
  assign n5366 = ~n5364 & ~n5365 ;
  assign n5368 = n5363 & ~n5366 ;
  assign n5367 = ~n5363 & n5366 ;
  assign n5369 = ~\TM0_pad  & ~n5367 ;
  assign n5370 = ~n5368 & n5369 ;
  assign n5371 = ~n5357 & ~n5370 ;
  assign n5372 = n1976 & ~n5371 ;
  assign n5373 = ~n1778 & ~n2900 ;
  assign n5374 = n1973 & ~n5373 ;
  assign n5375 = ~n5372 & ~n5374 ;
  assign n5376 = n3172 & ~n4005 ;
  assign n5378 = \TM0_pad  & ~\_2342__reg/NET0131  ;
  assign n5377 = ~\DATA_0_9_pad  & ~\TM0_pad  ;
  assign n5379 = n1976 & ~n5377 ;
  assign n5380 = ~n5378 & n5379 ;
  assign n5381 = ~n5376 & ~n5380 ;
  assign n5382 = RESET_pad & \WX10871_reg/NET0131  ;
  assign n5383 = \TM0_pad  & \_2298__reg/NET0131  ;
  assign n5384 = \WX9828_reg/NET0131  & ~\WX9892_reg/NET0131  ;
  assign n5385 = ~\WX9828_reg/NET0131  & \WX9892_reg/NET0131  ;
  assign n5386 = ~n5384 & ~n5385 ;
  assign n5387 = \WX9764_reg/NET0131  & ~n5386 ;
  assign n5388 = ~\WX9764_reg/NET0131  & n5386 ;
  assign n5389 = ~n5387 & ~n5388 ;
  assign n5390 = \TM1_pad  & ~\WX9700_reg/NET0131  ;
  assign n5391 = ~\TM1_pad  & \WX9700_reg/NET0131  ;
  assign n5392 = ~n5390 & ~n5391 ;
  assign n5394 = n5389 & ~n5392 ;
  assign n5393 = ~n5389 & n5392 ;
  assign n5395 = ~\TM0_pad  & ~n5393 ;
  assign n5396 = ~n5394 & n5395 ;
  assign n5397 = ~n5383 & ~n5396 ;
  assign n5398 = n1976 & ~n5397 ;
  assign n5399 = ~n1826 & ~n5351 ;
  assign n5400 = n1973 & ~n5399 ;
  assign n5401 = ~n5398 & ~n5400 ;
  assign n5402 = \TM0_pad  & \_2331__reg/NET0131  ;
  assign n5403 = ~n2333 & ~n5402 ;
  assign n5404 = n1976 & ~n5403 ;
  assign n5405 = ~n1855 & ~n5260 ;
  assign n5406 = n1973 & ~n5405 ;
  assign n5407 = ~n5404 & ~n5406 ;
  assign n5408 = \TM0_pad  & \_2199__reg/NET0131  ;
  assign n5409 = \WX5955_reg/NET0131  & ~\WX6019_reg/NET0131  ;
  assign n5410 = ~\WX5955_reg/NET0131  & \WX6019_reg/NET0131  ;
  assign n5411 = ~n5409 & ~n5410 ;
  assign n5412 = \WX5891_reg/NET0131  & ~n5411 ;
  assign n5413 = ~\WX5891_reg/NET0131  & n5411 ;
  assign n5414 = ~n5412 & ~n5413 ;
  assign n5415 = \TM1_pad  & ~\WX5827_reg/NET0131  ;
  assign n5416 = ~\TM1_pad  & \WX5827_reg/NET0131  ;
  assign n5417 = ~n5415 & ~n5416 ;
  assign n5419 = n5414 & ~n5417 ;
  assign n5418 = ~n5414 & n5417 ;
  assign n5420 = ~\TM0_pad  & ~n5418 ;
  assign n5421 = ~n5419 & n5420 ;
  assign n5422 = ~n5408 & ~n5421 ;
  assign n5423 = n1976 & ~n5422 ;
  assign n5424 = ~n1778 & ~n5370 ;
  assign n5425 = n1973 & ~n5424 ;
  assign n5426 = ~n5423 & ~n5425 ;
  assign n5427 = \TM0_pad  & \_2232__reg/NET0131  ;
  assign n5428 = \WX7246_reg/NET0131  & ~\WX7310_reg/NET0131  ;
  assign n5429 = ~\WX7246_reg/NET0131  & \WX7310_reg/NET0131  ;
  assign n5430 = ~n5428 & ~n5429 ;
  assign n5431 = \WX7182_reg/NET0131  & ~n5430 ;
  assign n5432 = ~\WX7182_reg/NET0131  & n5430 ;
  assign n5433 = ~n5431 & ~n5432 ;
  assign n5434 = \TM1_pad  & ~\WX7118_reg/NET0131  ;
  assign n5435 = ~\TM1_pad  & \WX7118_reg/NET0131  ;
  assign n5436 = ~n5434 & ~n5435 ;
  assign n5438 = n5433 & ~n5436 ;
  assign n5437 = ~n5433 & n5436 ;
  assign n5439 = ~\TM0_pad  & ~n5437 ;
  assign n5440 = ~n5438 & n5439 ;
  assign n5441 = ~n5427 & ~n5440 ;
  assign n5442 = n1976 & ~n5441 ;
  assign n5443 = ~n1794 & ~n5298 ;
  assign n5444 = n1973 & ~n5443 ;
  assign n5445 = ~n5442 & ~n5444 ;
  assign n5446 = \WX2112_reg/NET0131  & ~\WX2176_reg/NET0131  ;
  assign n5447 = ~\WX2112_reg/NET0131  & \WX2176_reg/NET0131  ;
  assign n5448 = ~n5446 & ~n5447 ;
  assign n5449 = \WX1984_reg/NET0131  & ~\WX2048_reg/NET0131  ;
  assign n5450 = ~\WX1984_reg/NET0131  & \WX2048_reg/NET0131  ;
  assign n5451 = ~n5449 & ~n5450 ;
  assign n5453 = n5448 & ~n5451 ;
  assign n5452 = ~n5448 & n5451 ;
  assign n5454 = ~\TM0_pad  & ~n5452 ;
  assign n5455 = ~n5453 & n5454 ;
  assign n5456 = n2023 & ~n5455 ;
  assign n5457 = \TM0_pad  & ~\_2117__reg/NET0131  ;
  assign n5458 = n1976 & ~n5457 ;
  assign n5459 = ~n3342 & n5458 ;
  assign n5460 = ~n5456 & ~n5459 ;
  assign n5461 = \TM0_pad  & \_2265__reg/NET0131  ;
  assign n5462 = \WX8537_reg/NET0131  & ~\WX8601_reg/NET0131  ;
  assign n5463 = ~\WX8537_reg/NET0131  & \WX8601_reg/NET0131  ;
  assign n5464 = ~n5462 & ~n5463 ;
  assign n5465 = \WX8473_reg/NET0131  & ~n5464 ;
  assign n5466 = ~\WX8473_reg/NET0131  & n5464 ;
  assign n5467 = ~n5465 & ~n5466 ;
  assign n5468 = \TM1_pad  & ~\WX8409_reg/NET0131  ;
  assign n5469 = ~\TM1_pad  & \WX8409_reg/NET0131  ;
  assign n5470 = ~n5468 & ~n5469 ;
  assign n5472 = n5467 & ~n5470 ;
  assign n5471 = ~n5467 & n5470 ;
  assign n5473 = ~\TM0_pad  & ~n5471 ;
  assign n5474 = ~n5472 & n5473 ;
  assign n5475 = ~n5461 & ~n5474 ;
  assign n5476 = n1976 & ~n5475 ;
  assign n5477 = ~n1810 & ~n5317 ;
  assign n5478 = n1973 & ~n5477 ;
  assign n5479 = ~n5476 & ~n5478 ;
  assign n5480 = \TM0_pad  & \_2166__reg/NET0131  ;
  assign n5481 = \WX4664_reg/NET0131  & ~\WX4728_reg/NET0131  ;
  assign n5482 = ~\WX4664_reg/NET0131  & \WX4728_reg/NET0131  ;
  assign n5483 = ~n5481 & ~n5482 ;
  assign n5484 = \WX4600_reg/NET0131  & ~n5483 ;
  assign n5485 = ~\WX4600_reg/NET0131  & n5483 ;
  assign n5486 = ~n5484 & ~n5485 ;
  assign n5487 = \TM1_pad  & ~\WX4536_reg/NET0131  ;
  assign n5488 = ~\TM1_pad  & \WX4536_reg/NET0131  ;
  assign n5489 = ~n5487 & ~n5488 ;
  assign n5491 = n5486 & ~n5489 ;
  assign n5490 = ~n5486 & n5489 ;
  assign n5492 = ~\TM0_pad  & ~n5490 ;
  assign n5493 = ~n5491 & n5492 ;
  assign n5494 = ~n5480 & ~n5493 ;
  assign n5495 = n1976 & ~n5494 ;
  assign n5496 = ~n1762 & ~n3065 ;
  assign n5497 = n1973 & ~n5496 ;
  assign n5498 = ~n5495 & ~n5497 ;
  assign n5499 = ~\TM0_pad  & ~n1929 ;
  assign n5500 = n3644 & ~n5499 ;
  assign n5502 = \WX2116_reg/NET0131  & ~\WX2180_reg/NET0131  ;
  assign n5503 = ~\WX2116_reg/NET0131  & \WX2180_reg/NET0131  ;
  assign n5504 = ~n5502 & ~n5503 ;
  assign n5505 = \WX1988_reg/NET0131  & ~\WX2052_reg/NET0131  ;
  assign n5506 = ~\WX1988_reg/NET0131  & \WX2052_reg/NET0131  ;
  assign n5507 = ~n5505 & ~n5506 ;
  assign n5509 = n5504 & ~n5507 ;
  assign n5508 = ~n5504 & n5507 ;
  assign n5510 = ~\TM0_pad  & ~n5508 ;
  assign n5511 = ~n5509 & n5510 ;
  assign n5501 = \TM0_pad  & ~\_2083__reg/NET0131  ;
  assign n5512 = n1976 & ~n5501 ;
  assign n5513 = ~n5511 & n5512 ;
  assign n5514 = ~n5500 & ~n5513 ;
  assign n5515 = RESET_pad & \WX10873_reg/NET0131  ;
  assign n5516 = \TM0_pad  & \_2297__reg/NET0131  ;
  assign n5517 = ~n2003 & ~n5516 ;
  assign n5518 = n1976 & ~n5517 ;
  assign n5519 = ~n1810 & ~n5474 ;
  assign n5520 = n1973 & ~n5519 ;
  assign n5521 = ~n5518 & ~n5520 ;
  assign n5522 = \TM0_pad  & \_2330__reg/NET0131  ;
  assign n5523 = ~n2509 & ~n5522 ;
  assign n5524 = n1976 & ~n5523 ;
  assign n5525 = ~n1826 & ~n5396 ;
  assign n5526 = n1973 & ~n5525 ;
  assign n5527 = ~n5524 & ~n5526 ;
  assign n5528 = \TM0_pad  & \_2198__reg/NET0131  ;
  assign n5529 = \WX5957_reg/NET0131  & ~\WX6021_reg/NET0131  ;
  assign n5530 = ~\WX5957_reg/NET0131  & \WX6021_reg/NET0131  ;
  assign n5531 = ~n5529 & ~n5530 ;
  assign n5532 = \WX5893_reg/NET0131  & ~n5531 ;
  assign n5533 = ~\WX5893_reg/NET0131  & n5531 ;
  assign n5534 = ~n5532 & ~n5533 ;
  assign n5535 = \TM1_pad  & ~\WX5829_reg/NET0131  ;
  assign n5536 = ~\TM1_pad  & \WX5829_reg/NET0131  ;
  assign n5537 = ~n5535 & ~n5536 ;
  assign n5539 = n5534 & ~n5537 ;
  assign n5538 = ~n5534 & n5537 ;
  assign n5540 = ~\TM0_pad  & ~n5538 ;
  assign n5541 = ~n5539 & n5540 ;
  assign n5542 = ~n5528 & ~n5541 ;
  assign n5543 = n1976 & ~n5542 ;
  assign n5544 = ~n1762 & ~n5493 ;
  assign n5545 = n1973 & ~n5544 ;
  assign n5546 = ~n5543 & ~n5545 ;
  assign n5547 = \TM0_pad  & \_2231__reg/NET0131  ;
  assign n5548 = \WX7248_reg/NET0131  & ~\WX7312_reg/NET0131  ;
  assign n5549 = ~\WX7248_reg/NET0131  & \WX7312_reg/NET0131  ;
  assign n5550 = ~n5548 & ~n5549 ;
  assign n5551 = \WX7184_reg/NET0131  & ~n5550 ;
  assign n5552 = ~\WX7184_reg/NET0131  & n5550 ;
  assign n5553 = ~n5551 & ~n5552 ;
  assign n5554 = \TM1_pad  & ~\WX7120_reg/NET0131  ;
  assign n5555 = ~\TM1_pad  & \WX7120_reg/NET0131  ;
  assign n5556 = ~n5554 & ~n5555 ;
  assign n5558 = n5553 & ~n5556 ;
  assign n5557 = ~n5553 & n5556 ;
  assign n5559 = ~\TM0_pad  & ~n5557 ;
  assign n5560 = ~n5558 & n5559 ;
  assign n5561 = ~n5547 & ~n5560 ;
  assign n5562 = n1976 & ~n5561 ;
  assign n5563 = ~n1778 & ~n5421 ;
  assign n5564 = n1973 & ~n5563 ;
  assign n5565 = ~n5562 & ~n5564 ;
  assign n5566 = \WX2114_reg/NET0131  & ~\WX2178_reg/NET0131  ;
  assign n5567 = ~\WX2114_reg/NET0131  & \WX2178_reg/NET0131  ;
  assign n5568 = ~n5566 & ~n5567 ;
  assign n5569 = \WX1986_reg/NET0131  & ~\WX2050_reg/NET0131  ;
  assign n5570 = ~\WX1986_reg/NET0131  & \WX2050_reg/NET0131  ;
  assign n5571 = ~n5569 & ~n5570 ;
  assign n5573 = n5568 & ~n5571 ;
  assign n5572 = ~n5568 & n5571 ;
  assign n5574 = ~\TM0_pad  & ~n5572 ;
  assign n5575 = ~n5573 & n5574 ;
  assign n5576 = n3483 & ~n5575 ;
  assign n5577 = \TM0_pad  & ~\_2116__reg/NET0131  ;
  assign n5578 = n1976 & ~n5577 ;
  assign n5579 = ~n3493 & n5578 ;
  assign n5580 = ~n5576 & ~n5579 ;
  assign n5581 = \TM0_pad  & \_2264__reg/NET0131  ;
  assign n5582 = \WX8539_reg/NET0131  & ~\WX8603_reg/NET0131  ;
  assign n5583 = ~\WX8539_reg/NET0131  & \WX8603_reg/NET0131  ;
  assign n5584 = ~n5582 & ~n5583 ;
  assign n5585 = \WX8475_reg/NET0131  & ~n5584 ;
  assign n5586 = ~\WX8475_reg/NET0131  & n5584 ;
  assign n5587 = ~n5585 & ~n5586 ;
  assign n5588 = \TM1_pad  & ~\WX8411_reg/NET0131  ;
  assign n5589 = ~\TM1_pad  & \WX8411_reg/NET0131  ;
  assign n5590 = ~n5588 & ~n5589 ;
  assign n5592 = n5587 & ~n5590 ;
  assign n5591 = ~n5587 & n5590 ;
  assign n5593 = ~\TM0_pad  & ~n5591 ;
  assign n5594 = ~n5592 & n5593 ;
  assign n5595 = ~n5581 & ~n5594 ;
  assign n5596 = n1976 & ~n5595 ;
  assign n5597 = ~n1794 & ~n5440 ;
  assign n5598 = n1973 & ~n5597 ;
  assign n5599 = ~n5596 & ~n5598 ;
  assign n5600 = \TM0_pad  & \_2165__reg/NET0131  ;
  assign n5601 = \WX4666_reg/NET0131  & ~\WX4730_reg/NET0131  ;
  assign n5602 = ~\WX4666_reg/NET0131  & \WX4730_reg/NET0131  ;
  assign n5603 = ~n5601 & ~n5602 ;
  assign n5604 = \WX4602_reg/NET0131  & ~n5603 ;
  assign n5605 = ~\WX4602_reg/NET0131  & n5603 ;
  assign n5606 = ~n5604 & ~n5605 ;
  assign n5607 = \TM1_pad  & ~\WX4538_reg/NET0131  ;
  assign n5608 = ~\TM1_pad  & \WX4538_reg/NET0131  ;
  assign n5609 = ~n5607 & ~n5608 ;
  assign n5611 = n5606 & ~n5609 ;
  assign n5610 = ~n5606 & n5609 ;
  assign n5612 = ~\TM0_pad  & ~n5610 ;
  assign n5613 = ~n5611 & n5612 ;
  assign n5614 = ~n5600 & ~n5613 ;
  assign n5615 = n1976 & ~n5614 ;
  assign n5616 = ~n1746 & ~n3241 ;
  assign n5617 = n1973 & ~n5616 ;
  assign n5618 = ~n5615 & ~n5617 ;
  assign n5619 = ~\TM0_pad  & ~n1916 ;
  assign n5620 = n3805 & ~n5619 ;
  assign n5622 = \WX2118_reg/NET0131  & ~\WX2182_reg/NET0131  ;
  assign n5623 = ~\WX2118_reg/NET0131  & \WX2182_reg/NET0131  ;
  assign n5624 = ~n5622 & ~n5623 ;
  assign n5625 = \WX1990_reg/NET0131  & ~\WX2054_reg/NET0131  ;
  assign n5626 = ~\WX1990_reg/NET0131  & \WX2054_reg/NET0131  ;
  assign n5627 = ~n5625 & ~n5626 ;
  assign n5629 = n5624 & ~n5627 ;
  assign n5628 = ~n5624 & n5627 ;
  assign n5630 = ~\TM0_pad  & ~n5628 ;
  assign n5631 = ~n5629 & n5630 ;
  assign n5621 = \TM0_pad  & ~\_2082__reg/NET0131  ;
  assign n5632 = n1976 & ~n5621 ;
  assign n5633 = ~n5631 & n5632 ;
  assign n5634 = ~n5620 & ~n5633 ;
  assign n5635 = n3483 & ~n4291 ;
  assign n5637 = \TM0_pad  & ~\_2340__reg/NET0131  ;
  assign n5636 = ~\DATA_0_7_pad  & ~\TM0_pad  ;
  assign n5638 = n1976 & ~n5636 ;
  assign n5639 = ~n5637 & n5638 ;
  assign n5640 = ~n5635 & ~n5639 ;
  assign n5641 = RESET_pad & \WX10875_reg/NET0131  ;
  assign n5642 = \TM0_pad  & \_2296__reg/NET0131  ;
  assign n5643 = \WX9832_reg/NET0131  & ~\WX9896_reg/NET0131  ;
  assign n5644 = ~\WX9832_reg/NET0131  & \WX9896_reg/NET0131  ;
  assign n5645 = ~n5643 & ~n5644 ;
  assign n5646 = \WX9768_reg/NET0131  & ~n5645 ;
  assign n5647 = ~\WX9768_reg/NET0131  & n5645 ;
  assign n5648 = ~n5646 & ~n5647 ;
  assign n5649 = \TM1_pad  & ~\WX9704_reg/NET0131  ;
  assign n5650 = ~\TM1_pad  & \WX9704_reg/NET0131  ;
  assign n5651 = ~n5649 & ~n5650 ;
  assign n5653 = n5648 & ~n5651 ;
  assign n5652 = ~n5648 & n5651 ;
  assign n5654 = ~\TM0_pad  & ~n5652 ;
  assign n5655 = ~n5653 & n5654 ;
  assign n5656 = ~n5642 & ~n5655 ;
  assign n5657 = n1976 & ~n5656 ;
  assign n5658 = ~n1794 & ~n5594 ;
  assign n5659 = n1973 & ~n5658 ;
  assign n5660 = ~n5657 & ~n5659 ;
  assign n5661 = \TM0_pad  & \_2197__reg/NET0131  ;
  assign n5662 = \WX5959_reg/NET0131  & ~\WX6023_reg/NET0131  ;
  assign n5663 = ~\WX5959_reg/NET0131  & \WX6023_reg/NET0131  ;
  assign n5664 = ~n5662 & ~n5663 ;
  assign n5665 = \WX5895_reg/NET0131  & ~n5664 ;
  assign n5666 = ~\WX5895_reg/NET0131  & n5664 ;
  assign n5667 = ~n5665 & ~n5666 ;
  assign n5668 = \TM1_pad  & ~\WX5831_reg/NET0131  ;
  assign n5669 = ~\TM1_pad  & \WX5831_reg/NET0131  ;
  assign n5670 = ~n5668 & ~n5669 ;
  assign n5672 = n5667 & ~n5670 ;
  assign n5671 = ~n5667 & n5670 ;
  assign n5673 = ~\TM0_pad  & ~n5671 ;
  assign n5674 = ~n5672 & n5673 ;
  assign n5675 = ~n5661 & ~n5674 ;
  assign n5676 = n1976 & ~n5675 ;
  assign n5677 = ~n1746 & ~n5613 ;
  assign n5678 = n1973 & ~n5677 ;
  assign n5679 = ~n5676 & ~n5678 ;
  assign n5680 = \TM0_pad  & \_2230__reg/NET0131  ;
  assign n5681 = \WX7250_reg/NET0131  & ~\WX7314_reg/NET0131  ;
  assign n5682 = ~\WX7250_reg/NET0131  & \WX7314_reg/NET0131  ;
  assign n5683 = ~n5681 & ~n5682 ;
  assign n5684 = \WX7186_reg/NET0131  & ~n5683 ;
  assign n5685 = ~\WX7186_reg/NET0131  & n5683 ;
  assign n5686 = ~n5684 & ~n5685 ;
  assign n5687 = \TM1_pad  & ~\WX7122_reg/NET0131  ;
  assign n5688 = ~\TM1_pad  & \WX7122_reg/NET0131  ;
  assign n5689 = ~n5687 & ~n5688 ;
  assign n5691 = n5686 & ~n5689 ;
  assign n5690 = ~n5686 & n5689 ;
  assign n5692 = ~\TM0_pad  & ~n5690 ;
  assign n5693 = ~n5691 & n5692 ;
  assign n5694 = ~n5680 & ~n5693 ;
  assign n5695 = n1976 & ~n5694 ;
  assign n5696 = ~n1762 & ~n5541 ;
  assign n5697 = n1973 & ~n5696 ;
  assign n5698 = ~n5695 & ~n5697 ;
  assign n5699 = n3644 & ~n5511 ;
  assign n5700 = \TM0_pad  & ~\_2115__reg/NET0131  ;
  assign n5701 = n1976 & ~n5700 ;
  assign n5702 = ~n3654 & n5701 ;
  assign n5703 = ~n5699 & ~n5702 ;
  assign n5704 = \TM0_pad  & \_2263__reg/NET0131  ;
  assign n5705 = \WX8541_reg/NET0131  & ~\WX8605_reg/NET0131  ;
  assign n5706 = ~\WX8541_reg/NET0131  & \WX8605_reg/NET0131  ;
  assign n5707 = ~n5705 & ~n5706 ;
  assign n5708 = \WX8477_reg/NET0131  & ~n5707 ;
  assign n5709 = ~\WX8477_reg/NET0131  & n5707 ;
  assign n5710 = ~n5708 & ~n5709 ;
  assign n5711 = \TM1_pad  & ~\WX8413_reg/NET0131  ;
  assign n5712 = ~\TM1_pad  & \WX8413_reg/NET0131  ;
  assign n5713 = ~n5711 & ~n5712 ;
  assign n5715 = n5710 & ~n5713 ;
  assign n5714 = ~n5710 & n5713 ;
  assign n5716 = ~\TM0_pad  & ~n5714 ;
  assign n5717 = ~n5715 & n5716 ;
  assign n5718 = ~n5704 & ~n5717 ;
  assign n5719 = n1976 & ~n5718 ;
  assign n5720 = ~n1778 & ~n5560 ;
  assign n5721 = n1973 & ~n5720 ;
  assign n5722 = ~n5719 & ~n5721 ;
  assign n5723 = \TM0_pad  & \_2164__reg/NET0131  ;
  assign n5724 = \WX4668_reg/NET0131  & ~\WX4732_reg/NET0131  ;
  assign n5725 = ~\WX4668_reg/NET0131  & \WX4732_reg/NET0131  ;
  assign n5726 = ~n5724 & ~n5725 ;
  assign n5727 = \WX4604_reg/NET0131  & ~n5726 ;
  assign n5728 = ~\WX4604_reg/NET0131  & n5726 ;
  assign n5729 = ~n5727 & ~n5728 ;
  assign n5730 = \TM1_pad  & ~\WX4540_reg/NET0131  ;
  assign n5731 = ~\TM1_pad  & \WX4540_reg/NET0131  ;
  assign n5732 = ~n5730 & ~n5731 ;
  assign n5734 = n5729 & ~n5732 ;
  assign n5733 = ~n5729 & n5732 ;
  assign n5735 = ~\TM0_pad  & ~n5733 ;
  assign n5736 = ~n5734 & n5735 ;
  assign n5737 = ~n5723 & ~n5736 ;
  assign n5738 = n1976 & ~n5737 ;
  assign n5739 = ~n1730 & ~n3391 ;
  assign n5740 = n1973 & ~n5739 ;
  assign n5741 = ~n5738 & ~n5740 ;
  assign n5742 = ~\TM0_pad  & ~n1880 ;
  assign n5743 = ~n1871 & ~n5742 ;
  assign n5744 = n1973 & ~n5743 ;
  assign n5745 = \TM0_pad  & \_2108__reg/NET0131  ;
  assign n5746 = \TM1_pad  & ~\WX1938_reg/NET0131  ;
  assign n5747 = ~\TM1_pad  & \WX1938_reg/NET0131  ;
  assign n5748 = ~n5746 & ~n5747 ;
  assign n5749 = ~\WX2002_reg/NET0131  & ~n5748 ;
  assign n5750 = \WX2002_reg/NET0131  & n5748 ;
  assign n5751 = ~n5749 & ~n5750 ;
  assign n5752 = \WX2066_reg/NET0131  & ~\WX2130_reg/NET0131  ;
  assign n5753 = ~\WX2066_reg/NET0131  & \WX2130_reg/NET0131  ;
  assign n5754 = ~n5752 & ~n5753 ;
  assign n5756 = ~n5751 & ~n5754 ;
  assign n5755 = n5751 & n5754 ;
  assign n5757 = ~\TM0_pad  & ~n5755 ;
  assign n5758 = ~n5756 & n5757 ;
  assign n5759 = ~n5745 & ~n5758 ;
  assign n5760 = n1976 & ~n5759 ;
  assign n5761 = ~n5744 & ~n5760 ;
  assign n5762 = n3644 & ~n4434 ;
  assign n5764 = \TM0_pad  & ~\_2339__reg/NET0131  ;
  assign n5763 = ~\DATA_0_6_pad  & ~\TM0_pad  ;
  assign n5765 = n1976 & ~n5763 ;
  assign n5766 = ~n5764 & n5765 ;
  assign n5767 = ~n5762 & ~n5766 ;
  assign n5768 = RESET_pad & \WX10877_reg/NET0131  ;
  assign n5769 = \TM0_pad  & \_2163__reg/NET0131  ;
  assign n5770 = \WX4670_reg/NET0131  & ~\WX4734_reg/NET0131  ;
  assign n5771 = ~\WX4670_reg/NET0131  & \WX4734_reg/NET0131  ;
  assign n5772 = ~n5770 & ~n5771 ;
  assign n5773 = \WX4606_reg/NET0131  & ~n5772 ;
  assign n5774 = ~\WX4606_reg/NET0131  & n5772 ;
  assign n5775 = ~n5773 & ~n5774 ;
  assign n5776 = \TM1_pad  & ~\WX4542_reg/NET0131  ;
  assign n5777 = ~\TM1_pad  & \WX4542_reg/NET0131  ;
  assign n5778 = ~n5776 & ~n5777 ;
  assign n5780 = n5775 & ~n5778 ;
  assign n5779 = ~n5775 & n5778 ;
  assign n5781 = ~\TM0_pad  & ~n5779 ;
  assign n5782 = ~n5780 & n5781 ;
  assign n5783 = ~n5769 & ~n5782 ;
  assign n5784 = n1976 & ~n5783 ;
  assign n5785 = ~n1714 & ~n3552 ;
  assign n5786 = n1973 & ~n5785 ;
  assign n5787 = ~n5784 & ~n5786 ;
  assign n5788 = \TM0_pad  & \_2295__reg/NET0131  ;
  assign n5789 = \WX9834_reg/NET0131  & ~\WX9898_reg/NET0131  ;
  assign n5790 = ~\WX9834_reg/NET0131  & \WX9898_reg/NET0131  ;
  assign n5791 = ~n5789 & ~n5790 ;
  assign n5792 = \WX9770_reg/NET0131  & ~n5791 ;
  assign n5793 = ~\WX9770_reg/NET0131  & n5791 ;
  assign n5794 = ~n5792 & ~n5793 ;
  assign n5795 = \TM1_pad  & ~\WX9706_reg/NET0131  ;
  assign n5796 = ~\TM1_pad  & \WX9706_reg/NET0131  ;
  assign n5797 = ~n5795 & ~n5796 ;
  assign n5799 = n5794 & ~n5797 ;
  assign n5798 = ~n5794 & n5797 ;
  assign n5800 = ~\TM0_pad  & ~n5798 ;
  assign n5801 = ~n5799 & n5800 ;
  assign n5802 = ~n5788 & ~n5801 ;
  assign n5803 = n1976 & ~n5802 ;
  assign n5804 = ~n1778 & ~n5717 ;
  assign n5805 = n1973 & ~n5804 ;
  assign n5806 = ~n5803 & ~n5805 ;
  assign n5807 = \TM0_pad  & \_2328__reg/NET0131  ;
  assign n5808 = ~n2837 & ~n5807 ;
  assign n5809 = n1976 & ~n5808 ;
  assign n5810 = ~n1794 & ~n5655 ;
  assign n5811 = n1973 & ~n5810 ;
  assign n5812 = ~n5809 & ~n5811 ;
  assign n5813 = \TM0_pad  & \_2196__reg/NET0131  ;
  assign n5814 = \WX5961_reg/NET0131  & ~\WX6025_reg/NET0131  ;
  assign n5815 = ~\WX5961_reg/NET0131  & \WX6025_reg/NET0131  ;
  assign n5816 = ~n5814 & ~n5815 ;
  assign n5817 = \WX5897_reg/NET0131  & ~n5816 ;
  assign n5818 = ~\WX5897_reg/NET0131  & n5816 ;
  assign n5819 = ~n5817 & ~n5818 ;
  assign n5820 = \TM1_pad  & ~\WX5833_reg/NET0131  ;
  assign n5821 = ~\TM1_pad  & \WX5833_reg/NET0131  ;
  assign n5822 = ~n5820 & ~n5821 ;
  assign n5824 = n5819 & ~n5822 ;
  assign n5823 = ~n5819 & n5822 ;
  assign n5825 = ~\TM0_pad  & ~n5823 ;
  assign n5826 = ~n5824 & n5825 ;
  assign n5827 = ~n5813 & ~n5826 ;
  assign n5828 = n1976 & ~n5827 ;
  assign n5829 = ~n1730 & ~n5736 ;
  assign n5830 = n1973 & ~n5829 ;
  assign n5831 = ~n5828 & ~n5830 ;
  assign n5832 = \TM0_pad  & \_2229__reg/NET0131  ;
  assign n5833 = \WX7252_reg/NET0131  & ~\WX7316_reg/NET0131  ;
  assign n5834 = ~\WX7252_reg/NET0131  & \WX7316_reg/NET0131  ;
  assign n5835 = ~n5833 & ~n5834 ;
  assign n5836 = \WX7188_reg/NET0131  & ~n5835 ;
  assign n5837 = ~\WX7188_reg/NET0131  & n5835 ;
  assign n5838 = ~n5836 & ~n5837 ;
  assign n5839 = \TM1_pad  & ~\WX7124_reg/NET0131  ;
  assign n5840 = ~\TM1_pad  & \WX7124_reg/NET0131  ;
  assign n5841 = ~n5839 & ~n5840 ;
  assign n5843 = n5838 & ~n5841 ;
  assign n5842 = ~n5838 & n5841 ;
  assign n5844 = ~\TM0_pad  & ~n5842 ;
  assign n5845 = ~n5843 & n5844 ;
  assign n5846 = ~n5832 & ~n5845 ;
  assign n5847 = n1976 & ~n5846 ;
  assign n5848 = ~n1746 & ~n5674 ;
  assign n5849 = n1973 & ~n5848 ;
  assign n5850 = ~n5847 & ~n5849 ;
  assign n5851 = n3805 & ~n5631 ;
  assign n5852 = \TM0_pad  & ~\_2114__reg/NET0131  ;
  assign n5853 = n1976 & ~n5852 ;
  assign n5854 = ~n3815 & n5853 ;
  assign n5855 = ~n5851 & ~n5854 ;
  assign n5856 = \TM0_pad  & \_2262__reg/NET0131  ;
  assign n5857 = \WX8543_reg/NET0131  & ~\WX8607_reg/NET0131  ;
  assign n5858 = ~\WX8543_reg/NET0131  & \WX8607_reg/NET0131  ;
  assign n5859 = ~n5857 & ~n5858 ;
  assign n5860 = \WX8479_reg/NET0131  & ~n5859 ;
  assign n5861 = ~\WX8479_reg/NET0131  & n5859 ;
  assign n5862 = ~n5860 & ~n5861 ;
  assign n5863 = \TM1_pad  & ~\WX8415_reg/NET0131  ;
  assign n5864 = ~\TM1_pad  & \WX8415_reg/NET0131  ;
  assign n5865 = ~n5863 & ~n5864 ;
  assign n5867 = n5862 & ~n5865 ;
  assign n5866 = ~n5862 & n5865 ;
  assign n5868 = ~\TM0_pad  & ~n5866 ;
  assign n5869 = ~n5867 & n5868 ;
  assign n5870 = ~n5856 & ~n5869 ;
  assign n5871 = n1976 & ~n5870 ;
  assign n5872 = ~n1762 & ~n5693 ;
  assign n5873 = n1973 & ~n5872 ;
  assign n5874 = ~n5871 & ~n5873 ;
  assign n5875 = ~\TM0_pad  & ~n1890 ;
  assign n5876 = n4101 & ~n5875 ;
  assign n5878 = \WX2122_reg/NET0131  & ~\WX2186_reg/NET0131  ;
  assign n5879 = ~\WX2122_reg/NET0131  & \WX2186_reg/NET0131  ;
  assign n5880 = ~n5878 & ~n5879 ;
  assign n5881 = \WX1994_reg/NET0131  & ~\WX2058_reg/NET0131  ;
  assign n5882 = ~\WX1994_reg/NET0131  & \WX2058_reg/NET0131  ;
  assign n5883 = ~n5881 & ~n5882 ;
  assign n5885 = n5880 & ~n5883 ;
  assign n5884 = ~n5880 & n5883 ;
  assign n5886 = ~\TM0_pad  & ~n5884 ;
  assign n5887 = ~n5885 & n5886 ;
  assign n5877 = \TM0_pad  & ~\_2080__reg/NET0131  ;
  assign n5888 = n1976 & ~n5877 ;
  assign n5889 = ~n5887 & n5888 ;
  assign n5890 = ~n5876 & ~n5889 ;
  assign n5891 = n3805 & ~n4562 ;
  assign n5893 = \TM0_pad  & ~\_2338__reg/NET0131  ;
  assign n5892 = ~\DATA_0_5_pad  & ~\TM0_pad  ;
  assign n5894 = n1976 & ~n5892 ;
  assign n5895 = ~n5893 & n5894 ;
  assign n5896 = ~n5891 & ~n5895 ;
  assign n5897 = RESET_pad & \WX10879_reg/NET0131  ;
  assign n5898 = \TM0_pad  & \_2162__reg/NET0131  ;
  assign n5899 = \WX4672_reg/NET0131  & ~\WX4736_reg/NET0131  ;
  assign n5900 = ~\WX4672_reg/NET0131  & \WX4736_reg/NET0131  ;
  assign n5901 = ~n5899 & ~n5900 ;
  assign n5902 = \WX4608_reg/NET0131  & ~n5901 ;
  assign n5903 = ~\WX4608_reg/NET0131  & n5901 ;
  assign n5904 = ~n5902 & ~n5903 ;
  assign n5905 = \TM1_pad  & ~\WX4544_reg/NET0131  ;
  assign n5906 = ~\TM1_pad  & \WX4544_reg/NET0131  ;
  assign n5907 = ~n5905 & ~n5906 ;
  assign n5909 = n5904 & ~n5907 ;
  assign n5908 = ~n5904 & n5907 ;
  assign n5910 = ~\TM0_pad  & ~n5908 ;
  assign n5911 = ~n5909 & n5910 ;
  assign n5912 = ~n5898 & ~n5911 ;
  assign n5913 = n1976 & ~n5912 ;
  assign n5914 = ~n1698 & ~n3713 ;
  assign n5915 = n1973 & ~n5914 ;
  assign n5916 = ~n5913 & ~n5915 ;
  assign n5917 = \TM0_pad  & \_2294__reg/NET0131  ;
  assign n5918 = \WX9836_reg/NET0131  & ~\WX9900_reg/NET0131  ;
  assign n5919 = ~\WX9836_reg/NET0131  & \WX9900_reg/NET0131  ;
  assign n5920 = ~n5918 & ~n5919 ;
  assign n5921 = \WX9772_reg/NET0131  & ~n5920 ;
  assign n5922 = ~\WX9772_reg/NET0131  & n5920 ;
  assign n5923 = ~n5921 & ~n5922 ;
  assign n5924 = \TM1_pad  & ~\WX9708_reg/NET0131  ;
  assign n5925 = ~\TM1_pad  & \WX9708_reg/NET0131  ;
  assign n5926 = ~n5924 & ~n5925 ;
  assign n5928 = n5923 & ~n5926 ;
  assign n5927 = ~n5923 & n5926 ;
  assign n5929 = ~\TM0_pad  & ~n5927 ;
  assign n5930 = ~n5928 & n5929 ;
  assign n5931 = ~n5917 & ~n5930 ;
  assign n5932 = n1976 & ~n5931 ;
  assign n5933 = ~n1762 & ~n5869 ;
  assign n5934 = n1973 & ~n5933 ;
  assign n5935 = ~n5932 & ~n5934 ;
  assign n5936 = \TM0_pad  & \_2140__reg/NET0131  ;
  assign n5937 = ~n4736 & ~n5936 ;
  assign n5938 = n1976 & ~n5937 ;
  assign n5939 = ~n1871 & ~n5758 ;
  assign n5940 = n1973 & ~n5939 ;
  assign n5941 = ~n5938 & ~n5940 ;
  assign n5942 = \TM0_pad  & \_2327__reg/NET0131  ;
  assign n5943 = ~n3002 & ~n5942 ;
  assign n5944 = n1976 & ~n5943 ;
  assign n5945 = ~n1778 & ~n5801 ;
  assign n5946 = n1973 & ~n5945 ;
  assign n5947 = ~n5944 & ~n5946 ;
  assign n5948 = \TM0_pad  & \_2195__reg/NET0131  ;
  assign n5949 = \WX5963_reg/NET0131  & ~\WX6027_reg/NET0131  ;
  assign n5950 = ~\WX5963_reg/NET0131  & \WX6027_reg/NET0131  ;
  assign n5951 = ~n5949 & ~n5950 ;
  assign n5952 = \WX5899_reg/NET0131  & ~n5951 ;
  assign n5953 = ~\WX5899_reg/NET0131  & n5951 ;
  assign n5954 = ~n5952 & ~n5953 ;
  assign n5955 = \TM1_pad  & ~\WX5835_reg/NET0131  ;
  assign n5956 = ~\TM1_pad  & \WX5835_reg/NET0131  ;
  assign n5957 = ~n5955 & ~n5956 ;
  assign n5959 = n5954 & ~n5957 ;
  assign n5958 = ~n5954 & n5957 ;
  assign n5960 = ~\TM0_pad  & ~n5958 ;
  assign n5961 = ~n5959 & n5960 ;
  assign n5962 = ~n5948 & ~n5961 ;
  assign n5963 = n1976 & ~n5962 ;
  assign n5964 = ~n1714 & ~n5782 ;
  assign n5965 = n1973 & ~n5964 ;
  assign n5966 = ~n5963 & ~n5965 ;
  assign n5967 = \TM0_pad  & \_2228__reg/NET0131  ;
  assign n5968 = \WX7254_reg/NET0131  & ~\WX7318_reg/NET0131  ;
  assign n5969 = ~\WX7254_reg/NET0131  & \WX7318_reg/NET0131  ;
  assign n5970 = ~n5968 & ~n5969 ;
  assign n5971 = \WX7190_reg/NET0131  & ~n5970 ;
  assign n5972 = ~\WX7190_reg/NET0131  & n5970 ;
  assign n5973 = ~n5971 & ~n5972 ;
  assign n5974 = \TM1_pad  & ~\WX7126_reg/NET0131  ;
  assign n5975 = ~\TM1_pad  & \WX7126_reg/NET0131  ;
  assign n5976 = ~n5974 & ~n5975 ;
  assign n5978 = n5973 & ~n5976 ;
  assign n5977 = ~n5973 & n5976 ;
  assign n5979 = ~\TM0_pad  & ~n5977 ;
  assign n5980 = ~n5978 & n5979 ;
  assign n5981 = ~n5967 & ~n5980 ;
  assign n5982 = n1976 & ~n5981 ;
  assign n5983 = ~n1730 & ~n5826 ;
  assign n5984 = n1973 & ~n5983 ;
  assign n5985 = ~n5982 & ~n5984 ;
  assign n5986 = \WX2120_reg/NET0131  & ~\WX2184_reg/NET0131  ;
  assign n5987 = ~\WX2120_reg/NET0131  & \WX2184_reg/NET0131  ;
  assign n5988 = ~n5986 & ~n5987 ;
  assign n5989 = \WX1992_reg/NET0131  & ~\WX2056_reg/NET0131  ;
  assign n5990 = ~\WX1992_reg/NET0131  & \WX2056_reg/NET0131  ;
  assign n5991 = ~n5989 & ~n5990 ;
  assign n5993 = n5988 & ~n5991 ;
  assign n5992 = ~n5988 & n5991 ;
  assign n5994 = ~\TM0_pad  & ~n5992 ;
  assign n5995 = ~n5993 & n5994 ;
  assign n5996 = n3953 & ~n5995 ;
  assign n5997 = \TM0_pad  & ~\_2113__reg/NET0131  ;
  assign n5998 = n1976 & ~n5997 ;
  assign n5999 = ~n3963 & n5998 ;
  assign n6000 = ~n5996 & ~n5999 ;
  assign n6001 = \TM0_pad  & \_2261__reg/NET0131  ;
  assign n6002 = \WX8545_reg/NET0131  & ~\WX8609_reg/NET0131  ;
  assign n6003 = ~\WX8545_reg/NET0131  & \WX8609_reg/NET0131  ;
  assign n6004 = ~n6002 & ~n6003 ;
  assign n6005 = \WX8481_reg/NET0131  & ~n6004 ;
  assign n6006 = ~\WX8481_reg/NET0131  & n6004 ;
  assign n6007 = ~n6005 & ~n6006 ;
  assign n6008 = \TM1_pad  & ~\WX8417_reg/NET0131  ;
  assign n6009 = ~\TM1_pad  & \WX8417_reg/NET0131  ;
  assign n6010 = ~n6008 & ~n6009 ;
  assign n6012 = n6007 & ~n6010 ;
  assign n6011 = ~n6007 & n6010 ;
  assign n6013 = ~\TM0_pad  & ~n6011 ;
  assign n6014 = ~n6012 & n6013 ;
  assign n6015 = ~n6001 & ~n6014 ;
  assign n6016 = n1976 & ~n6015 ;
  assign n6017 = ~n1746 & ~n5845 ;
  assign n6018 = n1973 & ~n6017 ;
  assign n6019 = ~n6016 & ~n6018 ;
  assign n6020 = ~\TM0_pad  & ~n1845 ;
  assign n6021 = n4239 & ~n6020 ;
  assign n6023 = \WX2124_reg/NET0131  & ~\WX2188_reg/NET0131  ;
  assign n6024 = ~\WX2124_reg/NET0131  & \WX2188_reg/NET0131  ;
  assign n6025 = ~n6023 & ~n6024 ;
  assign n6026 = \WX1996_reg/NET0131  & ~\WX2060_reg/NET0131  ;
  assign n6027 = ~\WX1996_reg/NET0131  & \WX2060_reg/NET0131  ;
  assign n6028 = ~n6026 & ~n6027 ;
  assign n6030 = n6025 & ~n6028 ;
  assign n6029 = ~n6025 & n6028 ;
  assign n6031 = ~\TM0_pad  & ~n6029 ;
  assign n6032 = ~n6030 & n6031 ;
  assign n6022 = \TM0_pad  & ~\_2079__reg/NET0131  ;
  assign n6033 = n1976 & ~n6022 ;
  assign n6034 = ~n6032 & n6033 ;
  assign n6035 = ~n6021 & ~n6034 ;
  assign n6036 = ~\TM0_pad  & ~n1517 ;
  assign n6037 = n4510 & ~n6036 ;
  assign n6039 = \WX2128_reg/NET0131  & ~\WX2192_reg/NET0131  ;
  assign n6040 = ~\WX2128_reg/NET0131  & \WX2192_reg/NET0131  ;
  assign n6041 = ~n6039 & ~n6040 ;
  assign n6042 = \WX2000_reg/NET0131  & ~\WX2064_reg/NET0131  ;
  assign n6043 = ~\WX2000_reg/NET0131  & \WX2064_reg/NET0131  ;
  assign n6044 = ~n6042 & ~n6043 ;
  assign n6046 = n6041 & ~n6044 ;
  assign n6045 = ~n6041 & n6044 ;
  assign n6047 = ~\TM0_pad  & ~n6045 ;
  assign n6048 = ~n6046 & n6047 ;
  assign n6038 = \TM0_pad  & ~\_2077__reg/NET0131  ;
  assign n6049 = n1976 & ~n6038 ;
  assign n6050 = ~n6048 & n6049 ;
  assign n6051 = ~n6037 & ~n6050 ;
  assign n6052 = ~n1871 & ~n5279 ;
  assign n6053 = n1973 & ~n6052 ;
  assign n6055 = \TM0_pad  & ~\_2364__reg/NET0131  ;
  assign n6054 = ~\DATA_0_31_pad  & ~\TM0_pad  ;
  assign n6056 = n1976 & ~n6054 ;
  assign n6057 = ~n6055 & n6056 ;
  assign n6058 = ~n6053 & ~n6057 ;
  assign n6059 = n3953 & ~n4659 ;
  assign n6061 = \TM0_pad  & ~\_2337__reg/NET0131  ;
  assign n6060 = ~\DATA_0_4_pad  & ~\TM0_pad  ;
  assign n6062 = n1976 & ~n6060 ;
  assign n6063 = ~n6061 & n6062 ;
  assign n6064 = ~n6059 & ~n6063 ;
  assign n6065 = RESET_pad & \WX10881_reg/NET0131  ;
  assign n6066 = \TM0_pad  & \_2161__reg/NET0131  ;
  assign n6067 = \WX4674_reg/NET0131  & ~\WX4738_reg/NET0131  ;
  assign n6068 = ~\WX4674_reg/NET0131  & \WX4738_reg/NET0131  ;
  assign n6069 = ~n6067 & ~n6068 ;
  assign n6070 = \WX4610_reg/NET0131  & ~n6069 ;
  assign n6071 = ~\WX4610_reg/NET0131  & n6069 ;
  assign n6072 = ~n6070 & ~n6071 ;
  assign n6073 = \TM1_pad  & ~\WX4546_reg/NET0131  ;
  assign n6074 = ~\TM1_pad  & \WX4546_reg/NET0131  ;
  assign n6075 = ~n6073 & ~n6074 ;
  assign n6077 = n6072 & ~n6075 ;
  assign n6076 = ~n6072 & n6075 ;
  assign n6078 = ~\TM0_pad  & ~n6076 ;
  assign n6079 = ~n6077 & n6078 ;
  assign n6080 = ~n6066 & ~n6079 ;
  assign n6081 = n1976 & ~n6080 ;
  assign n6082 = ~n1682 & ~n3874 ;
  assign n6083 = n1973 & ~n6082 ;
  assign n6084 = ~n6081 & ~n6083 ;
  assign n6085 = \TM0_pad  & \_2293__reg/NET0131  ;
  assign n6086 = \WX9838_reg/NET0131  & ~\WX9902_reg/NET0131  ;
  assign n6087 = ~\WX9838_reg/NET0131  & \WX9902_reg/NET0131  ;
  assign n6088 = ~n6086 & ~n6087 ;
  assign n6089 = \WX9774_reg/NET0131  & ~n6088 ;
  assign n6090 = ~\WX9774_reg/NET0131  & n6088 ;
  assign n6091 = ~n6089 & ~n6090 ;
  assign n6092 = \TM1_pad  & ~\WX9710_reg/NET0131  ;
  assign n6093 = ~\TM1_pad  & \WX9710_reg/NET0131  ;
  assign n6094 = ~n6092 & ~n6093 ;
  assign n6096 = n6091 & ~n6094 ;
  assign n6095 = ~n6091 & n6094 ;
  assign n6097 = ~\TM0_pad  & ~n6095 ;
  assign n6098 = ~n6096 & n6097 ;
  assign n6099 = ~n6085 & ~n6098 ;
  assign n6100 = n1976 & ~n6099 ;
  assign n6101 = ~n1746 & ~n6014 ;
  assign n6102 = n1973 & ~n6101 ;
  assign n6103 = ~n6100 & ~n6102 ;
  assign n6104 = \TM0_pad  & \_2326__reg/NET0131  ;
  assign n6105 = ~n3163 & ~n6104 ;
  assign n6106 = n1976 & ~n6105 ;
  assign n6107 = ~n1762 & ~n5930 ;
  assign n6108 = n1973 & ~n6107 ;
  assign n6109 = ~n6106 & ~n6108 ;
  assign n6110 = \TM0_pad  & \_2194__reg/NET0131  ;
  assign n6111 = \WX5965_reg/NET0131  & ~\WX6029_reg/NET0131  ;
  assign n6112 = ~\WX5965_reg/NET0131  & \WX6029_reg/NET0131  ;
  assign n6113 = ~n6111 & ~n6112 ;
  assign n6114 = \WX5901_reg/NET0131  & ~n6113 ;
  assign n6115 = ~\WX5901_reg/NET0131  & n6113 ;
  assign n6116 = ~n6114 & ~n6115 ;
  assign n6117 = \TM1_pad  & ~\WX5837_reg/NET0131  ;
  assign n6118 = ~\TM1_pad  & \WX5837_reg/NET0131  ;
  assign n6119 = ~n6117 & ~n6118 ;
  assign n6121 = n6116 & ~n6119 ;
  assign n6120 = ~n6116 & n6119 ;
  assign n6122 = ~\TM0_pad  & ~n6120 ;
  assign n6123 = ~n6121 & n6122 ;
  assign n6124 = ~n6110 & ~n6123 ;
  assign n6125 = n1976 & ~n6124 ;
  assign n6126 = ~n1698 & ~n5911 ;
  assign n6127 = n1973 & ~n6126 ;
  assign n6128 = ~n6125 & ~n6127 ;
  assign n6129 = \TM0_pad  & \_2227__reg/NET0131  ;
  assign n6130 = \WX7256_reg/NET0131  & ~\WX7320_reg/NET0131  ;
  assign n6131 = ~\WX7256_reg/NET0131  & \WX7320_reg/NET0131  ;
  assign n6132 = ~n6130 & ~n6131 ;
  assign n6133 = \WX7192_reg/NET0131  & ~n6132 ;
  assign n6134 = ~\WX7192_reg/NET0131  & n6132 ;
  assign n6135 = ~n6133 & ~n6134 ;
  assign n6136 = \TM1_pad  & ~\WX7128_reg/NET0131  ;
  assign n6137 = ~\TM1_pad  & \WX7128_reg/NET0131  ;
  assign n6138 = ~n6136 & ~n6137 ;
  assign n6140 = n6135 & ~n6138 ;
  assign n6139 = ~n6135 & n6138 ;
  assign n6141 = ~\TM0_pad  & ~n6139 ;
  assign n6142 = ~n6140 & n6141 ;
  assign n6143 = ~n6129 & ~n6142 ;
  assign n6144 = n1976 & ~n6143 ;
  assign n6145 = ~n1714 & ~n5961 ;
  assign n6146 = n1973 & ~n6145 ;
  assign n6147 = ~n6144 & ~n6146 ;
  assign n6148 = n4101 & ~n5887 ;
  assign n6149 = \TM0_pad  & ~\_2112__reg/NET0131  ;
  assign n6150 = n1976 & ~n6149 ;
  assign n6151 = ~n4111 & n6150 ;
  assign n6152 = ~n6148 & ~n6151 ;
  assign n6153 = \TM0_pad  & \_2260__reg/NET0131  ;
  assign n6154 = \WX8547_reg/NET0131  & ~\WX8611_reg/NET0131  ;
  assign n6155 = ~\WX8547_reg/NET0131  & \WX8611_reg/NET0131  ;
  assign n6156 = ~n6154 & ~n6155 ;
  assign n6157 = \WX8483_reg/NET0131  & ~n6156 ;
  assign n6158 = ~\WX8483_reg/NET0131  & n6156 ;
  assign n6159 = ~n6157 & ~n6158 ;
  assign n6160 = \TM1_pad  & ~\WX8419_reg/NET0131  ;
  assign n6161 = ~\TM1_pad  & \WX8419_reg/NET0131  ;
  assign n6162 = ~n6160 & ~n6161 ;
  assign n6164 = n6159 & ~n6162 ;
  assign n6163 = ~n6159 & n6162 ;
  assign n6165 = ~\TM0_pad  & ~n6163 ;
  assign n6166 = ~n6164 & n6165 ;
  assign n6167 = ~n6153 & ~n6166 ;
  assign n6168 = n1976 & ~n6167 ;
  assign n6169 = ~n1730 & ~n5980 ;
  assign n6170 = n1973 & ~n6169 ;
  assign n6171 = ~n6168 & ~n6170 ;
  assign n6172 = n4101 & ~n4823 ;
  assign n6174 = \TM0_pad  & ~\_2336__reg/NET0131  ;
  assign n6173 = ~\DATA_0_3_pad  & ~\TM0_pad  ;
  assign n6175 = n1976 & ~n6173 ;
  assign n6176 = ~n6174 & n6175 ;
  assign n6177 = ~n6172 & ~n6176 ;
  assign n6178 = RESET_pad & \WX10883_reg/NET0131  ;
  assign n6179 = \TM0_pad  & \_2160__reg/NET0131  ;
  assign n6180 = \TM1_pad  & ~\WX4548_reg/NET0131  ;
  assign n6181 = ~\TM1_pad  & \WX4548_reg/NET0131  ;
  assign n6182 = ~n6180 & ~n6181 ;
  assign n6183 = ~\WX4612_reg/NET0131  & ~n6182 ;
  assign n6184 = \WX4612_reg/NET0131  & n6182 ;
  assign n6185 = ~n6183 & ~n6184 ;
  assign n6186 = \WX4676_reg/NET0131  & ~\WX4740_reg/NET0131  ;
  assign n6187 = ~\WX4676_reg/NET0131  & \WX4740_reg/NET0131  ;
  assign n6188 = ~n6186 & ~n6187 ;
  assign n6190 = n6185 & n6188 ;
  assign n6189 = ~n6185 & ~n6188 ;
  assign n6191 = ~\TM0_pad  & ~n6189 ;
  assign n6192 = ~n6190 & n6191 ;
  assign n6193 = ~n6179 & ~n6192 ;
  assign n6194 = n1976 & ~n6193 ;
  assign n6195 = ~n1653 & ~n4022 ;
  assign n6196 = n1973 & ~n6195 ;
  assign n6197 = ~n6194 & ~n6196 ;
  assign n6198 = \TM0_pad  & \_2159__reg/NET0131  ;
  assign n6199 = \WX4678_reg/NET0131  & ~\WX4742_reg/NET0131  ;
  assign n6200 = ~\WX4678_reg/NET0131  & \WX4742_reg/NET0131  ;
  assign n6201 = ~n6199 & ~n6200 ;
  assign n6202 = \WX4614_reg/NET0131  & ~n6201 ;
  assign n6203 = ~\WX4614_reg/NET0131  & n6201 ;
  assign n6204 = ~n6202 & ~n6203 ;
  assign n6205 = \TM1_pad  & ~\WX4550_reg/NET0131  ;
  assign n6206 = ~\TM1_pad  & \WX4550_reg/NET0131  ;
  assign n6207 = ~n6205 & ~n6206 ;
  assign n6209 = n6204 & ~n6207 ;
  assign n6208 = ~n6204 & n6207 ;
  assign n6210 = ~\TM0_pad  & ~n6208 ;
  assign n6211 = ~n6209 & n6210 ;
  assign n6212 = ~n6198 & ~n6211 ;
  assign n6213 = n1976 & ~n6212 ;
  assign n6214 = ~n1637 & ~n4160 ;
  assign n6215 = n1973 & ~n6214 ;
  assign n6216 = ~n6213 & ~n6215 ;
  assign n6217 = \TM0_pad  & \_2158__reg/NET0131  ;
  assign n6218 = \WX4680_reg/NET0131  & ~\WX4744_reg/NET0131  ;
  assign n6219 = ~\WX4680_reg/NET0131  & \WX4744_reg/NET0131  ;
  assign n6220 = ~n6218 & ~n6219 ;
  assign n6221 = \WX4616_reg/NET0131  & ~n6220 ;
  assign n6222 = ~\WX4616_reg/NET0131  & n6220 ;
  assign n6223 = ~n6221 & ~n6222 ;
  assign n6224 = \TM1_pad  & ~\WX4552_reg/NET0131  ;
  assign n6225 = ~\TM1_pad  & \WX4552_reg/NET0131  ;
  assign n6226 = ~n6224 & ~n6225 ;
  assign n6228 = n6223 & ~n6226 ;
  assign n6227 = ~n6223 & n6226 ;
  assign n6229 = ~\TM0_pad  & ~n6227 ;
  assign n6230 = ~n6228 & n6229 ;
  assign n6231 = ~n6217 & ~n6230 ;
  assign n6232 = n1976 & ~n6231 ;
  assign n6233 = ~n1621 & ~n4323 ;
  assign n6234 = n1973 & ~n6233 ;
  assign n6235 = ~n6232 & ~n6234 ;
  assign n6236 = \TM0_pad  & \_2157__reg/NET0131  ;
  assign n6237 = ~n2233 & ~n6236 ;
  assign n6238 = n1976 & ~n6237 ;
  assign n6239 = ~n1605 & ~n4466 ;
  assign n6240 = n1973 & ~n6239 ;
  assign n6241 = ~n6238 & ~n6240 ;
  assign n6242 = \TM0_pad  & \_2292__reg/NET0131  ;
  assign n6243 = \WX9840_reg/NET0131  & ~\WX9904_reg/NET0131  ;
  assign n6244 = ~\WX9840_reg/NET0131  & \WX9904_reg/NET0131  ;
  assign n6245 = ~n6243 & ~n6244 ;
  assign n6246 = \WX9776_reg/NET0131  & ~n6245 ;
  assign n6247 = ~\WX9776_reg/NET0131  & n6245 ;
  assign n6248 = ~n6246 & ~n6247 ;
  assign n6249 = \TM1_pad  & ~\WX9712_reg/NET0131  ;
  assign n6250 = ~\TM1_pad  & \WX9712_reg/NET0131  ;
  assign n6251 = ~n6249 & ~n6250 ;
  assign n6253 = n6248 & ~n6251 ;
  assign n6252 = ~n6248 & n6251 ;
  assign n6254 = ~\TM0_pad  & ~n6252 ;
  assign n6255 = ~n6253 & n6254 ;
  assign n6256 = ~n6242 & ~n6255 ;
  assign n6257 = n1976 & ~n6256 ;
  assign n6258 = ~n1730 & ~n6166 ;
  assign n6259 = n1973 & ~n6258 ;
  assign n6260 = ~n6257 & ~n6259 ;
  assign n6261 = \TM0_pad  & \_2291__reg/NET0131  ;
  assign n6262 = \WX9842_reg/NET0131  & ~\WX9906_reg/NET0131  ;
  assign n6263 = ~\WX9842_reg/NET0131  & \WX9906_reg/NET0131  ;
  assign n6264 = ~n6262 & ~n6263 ;
  assign n6265 = \WX9778_reg/NET0131  & ~n6264 ;
  assign n6266 = ~\WX9778_reg/NET0131  & n6264 ;
  assign n6267 = ~n6265 & ~n6266 ;
  assign n6268 = \TM1_pad  & ~\WX9714_reg/NET0131  ;
  assign n6269 = ~\TM1_pad  & \WX9714_reg/NET0131  ;
  assign n6270 = ~n6268 & ~n6269 ;
  assign n6272 = n6267 & ~n6270 ;
  assign n6271 = ~n6267 & n6270 ;
  assign n6273 = ~\TM0_pad  & ~n6271 ;
  assign n6274 = ~n6272 & n6273 ;
  assign n6275 = ~n6261 & ~n6274 ;
  assign n6276 = n1976 & ~n6275 ;
  assign n6277 = \WX8549_reg/NET0131  & ~\WX8613_reg/NET0131  ;
  assign n6278 = ~\WX8549_reg/NET0131  & \WX8613_reg/NET0131  ;
  assign n6279 = ~n6277 & ~n6278 ;
  assign n6280 = \WX8485_reg/NET0131  & ~n6279 ;
  assign n6281 = ~\WX8485_reg/NET0131  & n6279 ;
  assign n6282 = ~n6280 & ~n6281 ;
  assign n6283 = \TM1_pad  & ~\WX8421_reg/NET0131  ;
  assign n6284 = ~\TM1_pad  & \WX8421_reg/NET0131  ;
  assign n6285 = ~n6283 & ~n6284 ;
  assign n6287 = n6282 & ~n6285 ;
  assign n6286 = ~n6282 & n6285 ;
  assign n6288 = ~\TM0_pad  & ~n6286 ;
  assign n6289 = ~n6287 & n6288 ;
  assign n6290 = ~n1714 & ~n6289 ;
  assign n6291 = n1973 & ~n6290 ;
  assign n6292 = ~n6276 & ~n6291 ;
  assign n6293 = \TM0_pad  & \_2290__reg/NET0131  ;
  assign n6294 = \WX9844_reg/NET0131  & ~\WX9908_reg/NET0131  ;
  assign n6295 = ~\WX9844_reg/NET0131  & \WX9908_reg/NET0131  ;
  assign n6296 = ~n6294 & ~n6295 ;
  assign n6297 = \WX9780_reg/NET0131  & ~n6296 ;
  assign n6298 = ~\WX9780_reg/NET0131  & n6296 ;
  assign n6299 = ~n6297 & ~n6298 ;
  assign n6300 = \TM1_pad  & ~\WX9716_reg/NET0131  ;
  assign n6301 = ~\TM1_pad  & \WX9716_reg/NET0131  ;
  assign n6302 = ~n6300 & ~n6301 ;
  assign n6304 = n6299 & ~n6302 ;
  assign n6303 = ~n6299 & n6302 ;
  assign n6305 = ~\TM0_pad  & ~n6303 ;
  assign n6306 = ~n6304 & n6305 ;
  assign n6307 = ~n6293 & ~n6306 ;
  assign n6308 = n1976 & ~n6307 ;
  assign n6309 = \WX8551_reg/NET0131  & ~\WX8615_reg/NET0131  ;
  assign n6310 = ~\WX8551_reg/NET0131  & \WX8615_reg/NET0131  ;
  assign n6311 = ~n6309 & ~n6310 ;
  assign n6312 = \WX8487_reg/NET0131  & ~n6311 ;
  assign n6313 = ~\WX8487_reg/NET0131  & n6311 ;
  assign n6314 = ~n6312 & ~n6313 ;
  assign n6315 = \TM1_pad  & ~\WX8423_reg/NET0131  ;
  assign n6316 = ~\TM1_pad  & \WX8423_reg/NET0131  ;
  assign n6317 = ~n6315 & ~n6316 ;
  assign n6319 = n6314 & ~n6317 ;
  assign n6318 = ~n6314 & n6317 ;
  assign n6320 = ~\TM0_pad  & ~n6318 ;
  assign n6321 = ~n6319 & n6320 ;
  assign n6322 = ~n1698 & ~n6321 ;
  assign n6323 = n1973 & ~n6322 ;
  assign n6324 = ~n6308 & ~n6323 ;
  assign n6325 = \TM0_pad  & \_2289__reg/NET0131  ;
  assign n6326 = ~n2201 & ~n6325 ;
  assign n6327 = n1976 & ~n6326 ;
  assign n6328 = \WX8553_reg/NET0131  & ~\WX8617_reg/NET0131  ;
  assign n6329 = ~\WX8553_reg/NET0131  & \WX8617_reg/NET0131  ;
  assign n6330 = ~n6328 & ~n6329 ;
  assign n6331 = \WX8489_reg/NET0131  & ~n6330 ;
  assign n6332 = ~\WX8489_reg/NET0131  & n6330 ;
  assign n6333 = ~n6331 & ~n6332 ;
  assign n6334 = \TM1_pad  & ~\WX8425_reg/NET0131  ;
  assign n6335 = ~\TM1_pad  & \WX8425_reg/NET0131  ;
  assign n6336 = ~n6334 & ~n6335 ;
  assign n6338 = n6333 & ~n6336 ;
  assign n6337 = ~n6333 & n6336 ;
  assign n6339 = ~\TM0_pad  & ~n6337 ;
  assign n6340 = ~n6338 & n6339 ;
  assign n6341 = ~n1682 & ~n6340 ;
  assign n6342 = n1973 & ~n6341 ;
  assign n6343 = ~n6327 & ~n6342 ;
  assign n6344 = \TM0_pad  & \_2325__reg/NET0131  ;
  assign n6345 = ~n3324 & ~n6344 ;
  assign n6346 = n1976 & ~n6345 ;
  assign n6347 = ~n1746 & ~n6098 ;
  assign n6348 = n1973 & ~n6347 ;
  assign n6349 = ~n6346 & ~n6348 ;
  assign n6350 = \TM0_pad  & \_2324__reg/NET0131  ;
  assign n6351 = ~n3474 & ~n6350 ;
  assign n6352 = n1976 & ~n6351 ;
  assign n6353 = ~n1730 & ~n6255 ;
  assign n6354 = n1973 & ~n6353 ;
  assign n6355 = ~n6352 & ~n6354 ;
  assign n6356 = \TM0_pad  & \_2323__reg/NET0131  ;
  assign n6357 = ~n3635 & ~n6356 ;
  assign n6358 = n1976 & ~n6357 ;
  assign n6359 = ~n1714 & ~n6274 ;
  assign n6360 = n1973 & ~n6359 ;
  assign n6361 = ~n6358 & ~n6360 ;
  assign n6362 = \TM0_pad  & \_2322__reg/NET0131  ;
  assign n6363 = ~n3796 & ~n6362 ;
  assign n6364 = n1976 & ~n6363 ;
  assign n6365 = ~n1698 & ~n6306 ;
  assign n6366 = n1973 & ~n6365 ;
  assign n6367 = ~n6364 & ~n6366 ;
  assign n6368 = \TM0_pad  & \_2193__reg/NET0131  ;
  assign n6369 = \WX5967_reg/NET0131  & ~\WX6031_reg/NET0131  ;
  assign n6370 = ~\WX5967_reg/NET0131  & \WX6031_reg/NET0131  ;
  assign n6371 = ~n6369 & ~n6370 ;
  assign n6372 = \WX5903_reg/NET0131  & ~n6371 ;
  assign n6373 = ~\WX5903_reg/NET0131  & n6371 ;
  assign n6374 = ~n6372 & ~n6373 ;
  assign n6375 = \TM1_pad  & ~\WX5839_reg/NET0131  ;
  assign n6376 = ~\TM1_pad  & \WX5839_reg/NET0131  ;
  assign n6377 = ~n6375 & ~n6376 ;
  assign n6379 = n6374 & ~n6377 ;
  assign n6378 = ~n6374 & n6377 ;
  assign n6380 = ~\TM0_pad  & ~n6378 ;
  assign n6381 = ~n6379 & n6380 ;
  assign n6382 = ~n6368 & ~n6381 ;
  assign n6383 = n1976 & ~n6382 ;
  assign n6384 = ~n1682 & ~n6079 ;
  assign n6385 = n1973 & ~n6384 ;
  assign n6386 = ~n6383 & ~n6385 ;
  assign n6387 = \TM0_pad  & \_2192__reg/NET0131  ;
  assign n6388 = \WX5969_reg/NET0131  & ~\WX6033_reg/NET0131  ;
  assign n6389 = ~\WX5969_reg/NET0131  & \WX6033_reg/NET0131  ;
  assign n6390 = ~n6388 & ~n6389 ;
  assign n6391 = \WX5905_reg/NET0131  & ~n6390 ;
  assign n6392 = ~\WX5905_reg/NET0131  & n6390 ;
  assign n6393 = ~n6391 & ~n6392 ;
  assign n6394 = \TM1_pad  & ~\WX5841_reg/NET0131  ;
  assign n6395 = ~\TM1_pad  & \WX5841_reg/NET0131  ;
  assign n6396 = ~n6394 & ~n6395 ;
  assign n6398 = n6393 & ~n6396 ;
  assign n6397 = ~n6393 & n6396 ;
  assign n6399 = ~\TM0_pad  & ~n6397 ;
  assign n6400 = ~n6398 & n6399 ;
  assign n6401 = ~n6387 & ~n6400 ;
  assign n6402 = n1976 & ~n6401 ;
  assign n6403 = ~n1653 & ~n6192 ;
  assign n6404 = n1973 & ~n6403 ;
  assign n6405 = ~n6402 & ~n6404 ;
  assign n6406 = \TM0_pad  & \_2191__reg/NET0131  ;
  assign n6407 = \WX5971_reg/NET0131  & ~\WX6035_reg/NET0131  ;
  assign n6408 = ~\WX5971_reg/NET0131  & \WX6035_reg/NET0131  ;
  assign n6409 = ~n6407 & ~n6408 ;
  assign n6410 = \WX5907_reg/NET0131  & ~n6409 ;
  assign n6411 = ~\WX5907_reg/NET0131  & n6409 ;
  assign n6412 = ~n6410 & ~n6411 ;
  assign n6413 = \TM1_pad  & ~\WX5843_reg/NET0131  ;
  assign n6414 = ~\TM1_pad  & \WX5843_reg/NET0131  ;
  assign n6415 = ~n6413 & ~n6414 ;
  assign n6417 = n6412 & ~n6415 ;
  assign n6416 = ~n6412 & n6415 ;
  assign n6418 = ~\TM0_pad  & ~n6416 ;
  assign n6419 = ~n6417 & n6418 ;
  assign n6420 = ~n6406 & ~n6419 ;
  assign n6421 = n1976 & ~n6420 ;
  assign n6422 = ~n1637 & ~n6211 ;
  assign n6423 = n1973 & ~n6422 ;
  assign n6424 = ~n6421 & ~n6423 ;
  assign n6425 = \TM0_pad  & \_2190__reg/NET0131  ;
  assign n6426 = ~n2265 & ~n6425 ;
  assign n6427 = n1976 & ~n6426 ;
  assign n6428 = ~n1621 & ~n6230 ;
  assign n6429 = n1973 & ~n6428 ;
  assign n6430 = ~n6427 & ~n6429 ;
  assign n6431 = \TM0_pad  & \_2226__reg/NET0131  ;
  assign n6432 = \WX7258_reg/NET0131  & ~\WX7322_reg/NET0131  ;
  assign n6433 = ~\WX7258_reg/NET0131  & \WX7322_reg/NET0131  ;
  assign n6434 = ~n6432 & ~n6433 ;
  assign n6435 = \WX7194_reg/NET0131  & ~n6434 ;
  assign n6436 = ~\WX7194_reg/NET0131  & n6434 ;
  assign n6437 = ~n6435 & ~n6436 ;
  assign n6438 = \TM1_pad  & ~\WX7130_reg/NET0131  ;
  assign n6439 = ~\TM1_pad  & \WX7130_reg/NET0131  ;
  assign n6440 = ~n6438 & ~n6439 ;
  assign n6442 = n6437 & ~n6440 ;
  assign n6441 = ~n6437 & n6440 ;
  assign n6443 = ~\TM0_pad  & ~n6441 ;
  assign n6444 = ~n6442 & n6443 ;
  assign n6445 = ~n6431 & ~n6444 ;
  assign n6446 = n1976 & ~n6445 ;
  assign n6447 = ~n1698 & ~n6123 ;
  assign n6448 = n1973 & ~n6447 ;
  assign n6449 = ~n6446 & ~n6448 ;
  assign n6450 = \TM0_pad  & \_2225__reg/NET0131  ;
  assign n6451 = \WX7260_reg/NET0131  & ~\WX7324_reg/NET0131  ;
  assign n6452 = ~\WX7260_reg/NET0131  & \WX7324_reg/NET0131  ;
  assign n6453 = ~n6451 & ~n6452 ;
  assign n6454 = \WX7196_reg/NET0131  & ~n6453 ;
  assign n6455 = ~\WX7196_reg/NET0131  & n6453 ;
  assign n6456 = ~n6454 & ~n6455 ;
  assign n6457 = \TM1_pad  & ~\WX7132_reg/NET0131  ;
  assign n6458 = ~\TM1_pad  & \WX7132_reg/NET0131  ;
  assign n6459 = ~n6457 & ~n6458 ;
  assign n6461 = n6456 & ~n6459 ;
  assign n6460 = ~n6456 & n6459 ;
  assign n6462 = ~\TM0_pad  & ~n6460 ;
  assign n6463 = ~n6461 & n6462 ;
  assign n6464 = ~n6450 & ~n6463 ;
  assign n6465 = n1976 & ~n6464 ;
  assign n6466 = ~n1682 & ~n6381 ;
  assign n6467 = n1973 & ~n6466 ;
  assign n6468 = ~n6465 & ~n6467 ;
  assign n6469 = \TM0_pad  & \_2224__reg/NET0131  ;
  assign n6470 = \WX7262_reg/NET0131  & ~\WX7326_reg/NET0131  ;
  assign n6471 = ~\WX7262_reg/NET0131  & \WX7326_reg/NET0131  ;
  assign n6472 = ~n6470 & ~n6471 ;
  assign n6473 = \WX7198_reg/NET0131  & ~n6472 ;
  assign n6474 = ~\WX7198_reg/NET0131  & n6472 ;
  assign n6475 = ~n6473 & ~n6474 ;
  assign n6476 = \TM1_pad  & ~\WX7134_reg/NET0131  ;
  assign n6477 = ~\TM1_pad  & \WX7134_reg/NET0131  ;
  assign n6478 = ~n6476 & ~n6477 ;
  assign n6480 = n6475 & ~n6478 ;
  assign n6479 = ~n6475 & n6478 ;
  assign n6481 = ~\TM0_pad  & ~n6479 ;
  assign n6482 = ~n6480 & n6481 ;
  assign n6483 = ~n6469 & ~n6482 ;
  assign n6484 = n1976 & ~n6483 ;
  assign n6485 = ~n1653 & ~n6400 ;
  assign n6486 = n1973 & ~n6485 ;
  assign n6487 = ~n6484 & ~n6486 ;
  assign n6488 = \TM0_pad  & \_2223__reg/NET0131  ;
  assign n6489 = ~n2297 & ~n6488 ;
  assign n6490 = n1976 & ~n6489 ;
  assign n6491 = ~n1637 & ~n6419 ;
  assign n6492 = n1973 & ~n6491 ;
  assign n6493 = ~n6490 & ~n6492 ;
  assign n6494 = n4239 & ~n6032 ;
  assign n6495 = \TM0_pad  & ~\_2111__reg/NET0131  ;
  assign n6496 = n1976 & ~n6495 ;
  assign n6497 = ~n4249 & n6496 ;
  assign n6498 = ~n6494 & ~n6497 ;
  assign n6499 = \WX2126_reg/NET0131  & ~\WX2190_reg/NET0131  ;
  assign n6500 = ~\WX2126_reg/NET0131  & \WX2190_reg/NET0131  ;
  assign n6501 = ~n6499 & ~n6500 ;
  assign n6502 = \WX1998_reg/NET0131  & ~\WX2062_reg/NET0131  ;
  assign n6503 = ~\WX1998_reg/NET0131  & \WX2062_reg/NET0131  ;
  assign n6504 = ~n6502 & ~n6503 ;
  assign n6506 = n6501 & ~n6504 ;
  assign n6505 = ~n6501 & n6504 ;
  assign n6507 = ~\TM0_pad  & ~n6505 ;
  assign n6508 = ~n6506 & n6507 ;
  assign n6509 = n4382 & ~n6508 ;
  assign n6510 = \TM0_pad  & ~\_2110__reg/NET0131  ;
  assign n6511 = n1976 & ~n6510 ;
  assign n6512 = ~n4392 & n6511 ;
  assign n6513 = ~n6509 & ~n6512 ;
  assign n6514 = n4510 & ~n6048 ;
  assign n6515 = \TM0_pad  & ~\_2109__reg/NET0131  ;
  assign n6516 = n1976 & ~n6515 ;
  assign n6517 = ~n4520 & n6516 ;
  assign n6518 = ~n6514 & ~n6517 ;
  assign n6519 = \TM0_pad  & \_2259__reg/NET0131  ;
  assign n6520 = ~n6289 & ~n6519 ;
  assign n6521 = n1976 & ~n6520 ;
  assign n6522 = ~n1714 & ~n6142 ;
  assign n6523 = n1973 & ~n6522 ;
  assign n6524 = ~n6521 & ~n6523 ;
  assign n6525 = \TM0_pad  & \_2258__reg/NET0131  ;
  assign n6526 = ~n6321 & ~n6525 ;
  assign n6527 = n1976 & ~n6526 ;
  assign n6528 = ~n1698 & ~n6444 ;
  assign n6529 = n1973 & ~n6528 ;
  assign n6530 = ~n6527 & ~n6529 ;
  assign n6531 = \TM0_pad  & \_2257__reg/NET0131  ;
  assign n6532 = ~n6340 & ~n6531 ;
  assign n6533 = n1976 & ~n6532 ;
  assign n6534 = ~n1682 & ~n6463 ;
  assign n6535 = n1973 & ~n6534 ;
  assign n6536 = ~n6533 & ~n6535 ;
  assign n6537 = \TM0_pad  & \_2256__reg/NET0131  ;
  assign n6538 = ~n2169 & ~n6537 ;
  assign n6539 = n1976 & ~n6538 ;
  assign n6540 = ~n1653 & ~n6482 ;
  assign n6541 = n1973 & ~n6540 ;
  assign n6542 = ~n6539 & ~n6541 ;
  assign n6543 = n4239 & ~n4927 ;
  assign n6545 = \TM0_pad  & ~\_2335__reg/NET0131  ;
  assign n6544 = ~\DATA_0_2_pad  & ~\TM0_pad  ;
  assign n6546 = n1976 & ~n6544 ;
  assign n6547 = ~n6545 & n6546 ;
  assign n6548 = ~n6543 & ~n6547 ;
  assign n6549 = n4382 & ~n5042 ;
  assign n6551 = \TM0_pad  & ~\_2334__reg/NET0131  ;
  assign n6550 = ~\DATA_0_1_pad  & ~\TM0_pad  ;
  assign n6552 = n1976 & ~n6550 ;
  assign n6553 = ~n6551 & n6552 ;
  assign n6554 = ~n6549 & ~n6553 ;
  assign n6555 = n4510 & ~n5174 ;
  assign n6557 = \TM0_pad  & ~\_2333__reg/NET0131  ;
  assign n6556 = ~\DATA_0_0_pad  & ~\TM0_pad  ;
  assign n6558 = n1976 & ~n6556 ;
  assign n6559 = ~n6557 & n6558 ;
  assign n6560 = ~n6555 & ~n6559 ;
  assign n6561 = RESET_pad & \WX10885_reg/NET0131  ;
  assign n6562 = ~\WX837_reg/NET0131  & ~\_2107__reg/NET0131  ;
  assign n6563 = \WX837_reg/NET0131  & \_2107__reg/NET0131  ;
  assign n6564 = ~n6562 & ~n6563 ;
  assign n6565 = RESET_pad & ~n6564 ;
  assign n6566 = ~\WX2130_reg/NET0131  & ~\_2139__reg/NET0131  ;
  assign n6567 = \WX2130_reg/NET0131  & \_2139__reg/NET0131  ;
  assign n6568 = ~n6566 & ~n6567 ;
  assign n6569 = RESET_pad & ~n6568 ;
  assign n6570 = ~\WX11181_reg/NET0131  & ~\_2363__reg/NET0131  ;
  assign n6571 = \WX11181_reg/NET0131  & \_2363__reg/NET0131  ;
  assign n6572 = ~n6570 & ~n6571 ;
  assign n6573 = RESET_pad & ~n6572 ;
  assign n6574 = RESET_pad & \WX10887_reg/NET0131  ;
  assign n6575 = ~\WX891_reg/NET0131  & ~\_2108__reg/NET0131  ;
  assign n6576 = \WX891_reg/NET0131  & \_2108__reg/NET0131  ;
  assign n6577 = ~n6575 & ~n6576 ;
  assign n6579 = ~\_2080__reg/NET0131  & n6577 ;
  assign n6578 = \_2080__reg/NET0131  & ~n6577 ;
  assign n6580 = RESET_pad & ~n6578 ;
  assign n6581 = ~n6579 & n6580 ;
  assign n6582 = ~\WX877_reg/NET0131  & ~\_2108__reg/NET0131  ;
  assign n6583 = \WX877_reg/NET0131  & \_2108__reg/NET0131  ;
  assign n6584 = ~n6582 & ~n6583 ;
  assign n6586 = ~\_2087__reg/NET0131  & n6584 ;
  assign n6585 = \_2087__reg/NET0131  & ~n6584 ;
  assign n6587 = RESET_pad & ~n6585 ;
  assign n6588 = ~n6586 & n6587 ;
  assign n6589 = ~\WX867_reg/NET0131  & ~\_2108__reg/NET0131  ;
  assign n6590 = \WX867_reg/NET0131  & \_2108__reg/NET0131  ;
  assign n6591 = ~n6589 & ~n6590 ;
  assign n6593 = ~\_2092__reg/NET0131  & n6591 ;
  assign n6592 = \_2092__reg/NET0131  & ~n6591 ;
  assign n6594 = RESET_pad & ~n6592 ;
  assign n6595 = ~n6593 & n6594 ;
  assign n6596 = ~\WX2184_reg/NET0131  & ~\_2140__reg/NET0131  ;
  assign n6597 = \WX2184_reg/NET0131  & \_2140__reg/NET0131  ;
  assign n6598 = ~n6596 & ~n6597 ;
  assign n6600 = ~\_2112__reg/NET0131  & n6598 ;
  assign n6599 = \_2112__reg/NET0131  & ~n6598 ;
  assign n6601 = RESET_pad & ~n6599 ;
  assign n6602 = ~n6600 & n6601 ;
  assign n6603 = ~\WX2170_reg/NET0131  & ~\_2140__reg/NET0131  ;
  assign n6604 = \WX2170_reg/NET0131  & \_2140__reg/NET0131  ;
  assign n6605 = ~n6603 & ~n6604 ;
  assign n6607 = ~\_2119__reg/NET0131  & n6605 ;
  assign n6606 = \_2119__reg/NET0131  & ~n6605 ;
  assign n6608 = RESET_pad & ~n6606 ;
  assign n6609 = ~n6607 & n6608 ;
  assign n6610 = ~\WX2160_reg/NET0131  & ~\_2140__reg/NET0131  ;
  assign n6611 = \WX2160_reg/NET0131  & \_2140__reg/NET0131  ;
  assign n6612 = ~n6610 & ~n6611 ;
  assign n6614 = ~\_2124__reg/NET0131  & n6612 ;
  assign n6613 = \_2124__reg/NET0131  & ~n6612 ;
  assign n6615 = RESET_pad & ~n6613 ;
  assign n6616 = ~n6614 & n6615 ;
  assign n6617 = ~\WX3477_reg/NET0131  & ~\_2172__reg/NET0131  ;
  assign n6618 = \WX3477_reg/NET0131  & \_2172__reg/NET0131  ;
  assign n6619 = ~n6617 & ~n6618 ;
  assign n6621 = ~\_2144__reg/NET0131  & n6619 ;
  assign n6620 = \_2144__reg/NET0131  & ~n6619 ;
  assign n6622 = RESET_pad & ~n6620 ;
  assign n6623 = ~n6621 & n6622 ;
  assign n6624 = ~\WX3463_reg/NET0131  & ~\_2172__reg/NET0131  ;
  assign n6625 = \WX3463_reg/NET0131  & \_2172__reg/NET0131  ;
  assign n6626 = ~n6624 & ~n6625 ;
  assign n6628 = ~\_2151__reg/NET0131  & n6626 ;
  assign n6627 = \_2151__reg/NET0131  & ~n6626 ;
  assign n6629 = RESET_pad & ~n6627 ;
  assign n6630 = ~n6628 & n6629 ;
  assign n6631 = ~\WX3453_reg/NET0131  & ~\_2172__reg/NET0131  ;
  assign n6632 = \WX3453_reg/NET0131  & \_2172__reg/NET0131  ;
  assign n6633 = ~n6631 & ~n6632 ;
  assign n6635 = ~\_2156__reg/NET0131  & n6633 ;
  assign n6634 = \_2156__reg/NET0131  & ~n6633 ;
  assign n6636 = RESET_pad & ~n6634 ;
  assign n6637 = ~n6635 & n6636 ;
  assign n6638 = ~\WX4770_reg/NET0131  & ~\_2204__reg/NET0131  ;
  assign n6639 = \WX4770_reg/NET0131  & \_2204__reg/NET0131  ;
  assign n6640 = ~n6638 & ~n6639 ;
  assign n6642 = ~\_2176__reg/NET0131  & n6640 ;
  assign n6641 = \_2176__reg/NET0131  & ~n6640 ;
  assign n6643 = RESET_pad & ~n6641 ;
  assign n6644 = ~n6642 & n6643 ;
  assign n6645 = ~\WX4756_reg/NET0131  & ~\_2204__reg/NET0131  ;
  assign n6646 = \WX4756_reg/NET0131  & \_2204__reg/NET0131  ;
  assign n6647 = ~n6645 & ~n6646 ;
  assign n6649 = ~\_2183__reg/NET0131  & n6647 ;
  assign n6648 = \_2183__reg/NET0131  & ~n6647 ;
  assign n6650 = RESET_pad & ~n6648 ;
  assign n6651 = ~n6649 & n6650 ;
  assign n6652 = ~\WX4746_reg/NET0131  & ~\_2204__reg/NET0131  ;
  assign n6653 = \WX4746_reg/NET0131  & \_2204__reg/NET0131  ;
  assign n6654 = ~n6652 & ~n6653 ;
  assign n6656 = ~\_2188__reg/NET0131  & n6654 ;
  assign n6655 = \_2188__reg/NET0131  & ~n6654 ;
  assign n6657 = RESET_pad & ~n6655 ;
  assign n6658 = ~n6656 & n6657 ;
  assign n6659 = ~\WX6063_reg/NET0131  & ~\_2236__reg/NET0131  ;
  assign n6660 = \WX6063_reg/NET0131  & \_2236__reg/NET0131  ;
  assign n6661 = ~n6659 & ~n6660 ;
  assign n6663 = ~\_2208__reg/NET0131  & n6661 ;
  assign n6662 = \_2208__reg/NET0131  & ~n6661 ;
  assign n6664 = RESET_pad & ~n6662 ;
  assign n6665 = ~n6663 & n6664 ;
  assign n6666 = ~\WX6049_reg/NET0131  & ~\_2236__reg/NET0131  ;
  assign n6667 = \WX6049_reg/NET0131  & \_2236__reg/NET0131  ;
  assign n6668 = ~n6666 & ~n6667 ;
  assign n6670 = ~\_2215__reg/NET0131  & n6668 ;
  assign n6669 = \_2215__reg/NET0131  & ~n6668 ;
  assign n6671 = RESET_pad & ~n6669 ;
  assign n6672 = ~n6670 & n6671 ;
  assign n6673 = ~\WX6039_reg/NET0131  & ~\_2236__reg/NET0131  ;
  assign n6674 = \WX6039_reg/NET0131  & \_2236__reg/NET0131  ;
  assign n6675 = ~n6673 & ~n6674 ;
  assign n6677 = ~\_2220__reg/NET0131  & n6675 ;
  assign n6676 = \_2220__reg/NET0131  & ~n6675 ;
  assign n6678 = RESET_pad & ~n6676 ;
  assign n6679 = ~n6677 & n6678 ;
  assign n6680 = ~\WX7356_reg/NET0131  & ~\_2268__reg/NET0131  ;
  assign n6681 = \WX7356_reg/NET0131  & \_2268__reg/NET0131  ;
  assign n6682 = ~n6680 & ~n6681 ;
  assign n6684 = ~\_2240__reg/NET0131  & n6682 ;
  assign n6683 = \_2240__reg/NET0131  & ~n6682 ;
  assign n6685 = RESET_pad & ~n6683 ;
  assign n6686 = ~n6684 & n6685 ;
  assign n6687 = ~\WX7342_reg/NET0131  & ~\_2268__reg/NET0131  ;
  assign n6688 = \WX7342_reg/NET0131  & \_2268__reg/NET0131  ;
  assign n6689 = ~n6687 & ~n6688 ;
  assign n6691 = ~\_2247__reg/NET0131  & n6689 ;
  assign n6690 = \_2247__reg/NET0131  & ~n6689 ;
  assign n6692 = RESET_pad & ~n6690 ;
  assign n6693 = ~n6691 & n6692 ;
  assign n6694 = ~\WX7332_reg/NET0131  & ~\_2268__reg/NET0131  ;
  assign n6695 = \WX7332_reg/NET0131  & \_2268__reg/NET0131  ;
  assign n6696 = ~n6694 & ~n6695 ;
  assign n6698 = ~\_2252__reg/NET0131  & n6696 ;
  assign n6697 = \_2252__reg/NET0131  & ~n6696 ;
  assign n6699 = RESET_pad & ~n6697 ;
  assign n6700 = ~n6698 & n6699 ;
  assign n6701 = ~\WX8649_reg/NET0131  & ~\_2300__reg/NET0131  ;
  assign n6702 = \WX8649_reg/NET0131  & \_2300__reg/NET0131  ;
  assign n6703 = ~n6701 & ~n6702 ;
  assign n6705 = ~\_2272__reg/NET0131  & n6703 ;
  assign n6704 = \_2272__reg/NET0131  & ~n6703 ;
  assign n6706 = RESET_pad & ~n6704 ;
  assign n6707 = ~n6705 & n6706 ;
  assign n6708 = ~\WX8635_reg/NET0131  & ~\_2300__reg/NET0131  ;
  assign n6709 = \WX8635_reg/NET0131  & \_2300__reg/NET0131  ;
  assign n6710 = ~n6708 & ~n6709 ;
  assign n6712 = ~\_2279__reg/NET0131  & n6710 ;
  assign n6711 = \_2279__reg/NET0131  & ~n6710 ;
  assign n6713 = RESET_pad & ~n6711 ;
  assign n6714 = ~n6712 & n6713 ;
  assign n6715 = ~\WX8625_reg/NET0131  & ~\_2300__reg/NET0131  ;
  assign n6716 = \WX8625_reg/NET0131  & \_2300__reg/NET0131  ;
  assign n6717 = ~n6715 & ~n6716 ;
  assign n6719 = ~\_2284__reg/NET0131  & n6717 ;
  assign n6718 = \_2284__reg/NET0131  & ~n6717 ;
  assign n6720 = RESET_pad & ~n6718 ;
  assign n6721 = ~n6719 & n6720 ;
  assign n6722 = ~\WX9942_reg/NET0131  & ~\_2332__reg/NET0131  ;
  assign n6723 = \WX9942_reg/NET0131  & \_2332__reg/NET0131  ;
  assign n6724 = ~n6722 & ~n6723 ;
  assign n6726 = ~\_2304__reg/NET0131  & n6724 ;
  assign n6725 = \_2304__reg/NET0131  & ~n6724 ;
  assign n6727 = RESET_pad & ~n6725 ;
  assign n6728 = ~n6726 & n6727 ;
  assign n6729 = ~\WX9928_reg/NET0131  & ~\_2332__reg/NET0131  ;
  assign n6730 = \WX9928_reg/NET0131  & \_2332__reg/NET0131  ;
  assign n6731 = ~n6729 & ~n6730 ;
  assign n6733 = ~\_2311__reg/NET0131  & n6731 ;
  assign n6732 = \_2311__reg/NET0131  & ~n6731 ;
  assign n6734 = RESET_pad & ~n6732 ;
  assign n6735 = ~n6733 & n6734 ;
  assign n6736 = ~\WX9918_reg/NET0131  & ~\_2332__reg/NET0131  ;
  assign n6737 = \WX9918_reg/NET0131  & \_2332__reg/NET0131  ;
  assign n6738 = ~n6736 & ~n6737 ;
  assign n6740 = ~\_2316__reg/NET0131  & n6738 ;
  assign n6739 = \_2316__reg/NET0131  & ~n6738 ;
  assign n6741 = RESET_pad & ~n6739 ;
  assign n6742 = ~n6740 & n6741 ;
  assign n6743 = ~\WX11235_reg/NET0131  & ~\_2364__reg/NET0131  ;
  assign n6744 = \WX11235_reg/NET0131  & \_2364__reg/NET0131  ;
  assign n6745 = ~n6743 & ~n6744 ;
  assign n6747 = ~\_2336__reg/NET0131  & n6745 ;
  assign n6746 = \_2336__reg/NET0131  & ~n6745 ;
  assign n6748 = RESET_pad & ~n6746 ;
  assign n6749 = ~n6747 & n6748 ;
  assign n6750 = ~\WX11221_reg/NET0131  & ~\_2364__reg/NET0131  ;
  assign n6751 = \WX11221_reg/NET0131  & \_2364__reg/NET0131  ;
  assign n6752 = ~n6750 & ~n6751 ;
  assign n6754 = ~\_2343__reg/NET0131  & n6752 ;
  assign n6753 = \_2343__reg/NET0131  & ~n6752 ;
  assign n6755 = RESET_pad & ~n6753 ;
  assign n6756 = ~n6754 & n6755 ;
  assign n6757 = ~\WX11211_reg/NET0131  & ~\_2364__reg/NET0131  ;
  assign n6758 = \WX11211_reg/NET0131  & \_2364__reg/NET0131  ;
  assign n6759 = ~n6757 & ~n6758 ;
  assign n6761 = ~\_2348__reg/NET0131  & n6759 ;
  assign n6760 = \_2348__reg/NET0131  & ~n6759 ;
  assign n6762 = RESET_pad & ~n6760 ;
  assign n6763 = ~n6761 & n6762 ;
  assign n6764 = RESET_pad & \WX11117_reg/NET0131  ;
  assign n6765 = RESET_pad & \WX773_reg/NET0131  ;
  assign n6766 = RESET_pad & \WX10889_reg/NET0131  ;
  assign n6767 = RESET_pad & \WX2066_reg/NET0131  ;
  assign n6768 = ~\WX3475_reg/NET0131  & ~\_2145__reg/NET0131  ;
  assign n6769 = \WX3475_reg/NET0131  & \_2145__reg/NET0131  ;
  assign n6770 = ~n6768 & ~n6769 ;
  assign n6771 = RESET_pad & ~n6770 ;
  assign n6772 = ~\WX3427_reg/NET0131  & ~\_2169__reg/NET0131  ;
  assign n6773 = \WX3427_reg/NET0131  & \_2169__reg/NET0131  ;
  assign n6774 = ~n6772 & ~n6773 ;
  assign n6775 = RESET_pad & ~n6774 ;
  assign n6776 = ~\WX2132_reg/NET0131  & ~\_2138__reg/NET0131  ;
  assign n6777 = \WX2132_reg/NET0131  & \_2138__reg/NET0131  ;
  assign n6778 = ~n6776 & ~n6777 ;
  assign n6779 = RESET_pad & ~n6778 ;
  assign n6780 = ~\WX11215_reg/NET0131  & ~\_2346__reg/NET0131  ;
  assign n6781 = \WX11215_reg/NET0131  & \_2346__reg/NET0131  ;
  assign n6782 = ~n6780 & ~n6781 ;
  assign n6783 = RESET_pad & ~n6782 ;
  assign n6784 = ~\WX8599_reg/NET0131  & ~\_2297__reg/NET0131  ;
  assign n6785 = \WX8599_reg/NET0131  & \_2297__reg/NET0131  ;
  assign n6786 = ~n6784 & ~n6785 ;
  assign n6787 = RESET_pad & ~n6786 ;
  assign n6788 = ~\WX6043_reg/NET0131  & ~\_2218__reg/NET0131  ;
  assign n6789 = \WX6043_reg/NET0131  & \_2218__reg/NET0131  ;
  assign n6790 = ~n6788 & ~n6789 ;
  assign n6791 = RESET_pad & ~n6790 ;
  assign n6792 = ~\WX3461_reg/NET0131  & ~\_2152__reg/NET0131  ;
  assign n6793 = \WX3461_reg/NET0131  & \_2152__reg/NET0131  ;
  assign n6794 = ~n6792 & ~n6793 ;
  assign n6795 = RESET_pad & ~n6794 ;
  assign n6796 = ~\WX857_reg/NET0131  & ~\_2097__reg/NET0131  ;
  assign n6797 = \WX857_reg/NET0131  & \_2097__reg/NET0131  ;
  assign n6798 = ~n6796 & ~n6797 ;
  assign n6799 = RESET_pad & ~n6798 ;
  assign n6800 = ~\WX9934_reg/NET0131  & ~\_2308__reg/NET0131  ;
  assign n6801 = \WX9934_reg/NET0131  & \_2308__reg/NET0131  ;
  assign n6802 = ~n6800 & ~n6801 ;
  assign n6803 = RESET_pad & ~n6802 ;
  assign n6804 = ~\WX7312_reg/NET0131  & ~\_2262__reg/NET0131  ;
  assign n6805 = \WX7312_reg/NET0131  & \_2262__reg/NET0131  ;
  assign n6806 = ~n6804 & ~n6805 ;
  assign n6807 = RESET_pad & ~n6806 ;
  assign n6808 = ~\WX7338_reg/NET0131  & ~\_2249__reg/NET0131  ;
  assign n6809 = \WX7338_reg/NET0131  & \_2249__reg/NET0131  ;
  assign n6810 = ~n6808 & ~n6809 ;
  assign n6811 = RESET_pad & ~n6810 ;
  assign n6812 = ~\WX8605_reg/NET0131  & ~\_2294__reg/NET0131  ;
  assign n6813 = \WX8605_reg/NET0131  & \_2294__reg/NET0131  ;
  assign n6814 = ~n6812 & ~n6813 ;
  assign n6815 = RESET_pad & ~n6814 ;
  assign n6816 = ~\WX8601_reg/NET0131  & ~\_2296__reg/NET0131  ;
  assign n6817 = \WX8601_reg/NET0131  & \_2296__reg/NET0131  ;
  assign n6818 = ~n6816 & ~n6817 ;
  assign n6819 = RESET_pad & ~n6818 ;
  assign n6820 = ~\WX8603_reg/NET0131  & ~\_2295__reg/NET0131  ;
  assign n6821 = \WX8603_reg/NET0131  & \_2295__reg/NET0131  ;
  assign n6822 = ~n6820 & ~n6821 ;
  assign n6823 = RESET_pad & ~n6822 ;
  assign n6824 = ~\WX6037_reg/NET0131  & ~\_2221__reg/NET0131  ;
  assign n6825 = \WX6037_reg/NET0131  & \_2221__reg/NET0131  ;
  assign n6826 = ~n6824 & ~n6825 ;
  assign n6827 = RESET_pad & ~n6826 ;
  assign n6828 = ~\WX8619_reg/NET0131  & ~\_2287__reg/NET0131  ;
  assign n6829 = \WX8619_reg/NET0131  & \_2287__reg/NET0131  ;
  assign n6830 = ~n6828 & ~n6829 ;
  assign n6831 = RESET_pad & ~n6830 ;
  assign n6832 = ~\WX7362_reg/NET0131  & ~\_2237__reg/NET0131  ;
  assign n6833 = \WX7362_reg/NET0131  & \_2237__reg/NET0131  ;
  assign n6834 = ~n6832 & ~n6833 ;
  assign n6835 = RESET_pad & ~n6834 ;
  assign n6836 = ~\WX3425_reg/NET0131  & ~\_2170__reg/NET0131  ;
  assign n6837 = \WX3425_reg/NET0131  & \_2170__reg/NET0131  ;
  assign n6838 = ~n6836 & ~n6837 ;
  assign n6839 = RESET_pad & ~n6838 ;
  assign n6840 = ~\WX4728_reg/NET0131  & ~\_2197__reg/NET0131  ;
  assign n6841 = \WX4728_reg/NET0131  & \_2197__reg/NET0131  ;
  assign n6842 = ~n6840 & ~n6841 ;
  assign n6843 = RESET_pad & ~n6842 ;
  assign n6844 = ~\WX3485_reg/NET0131  & ~\_2172__reg/NET0131  ;
  assign n6845 = \WX3485_reg/NET0131  & \_2172__reg/NET0131  ;
  assign n6846 = ~n6844 & ~n6845 ;
  assign n6847 = RESET_pad & ~n6846 ;
  assign n6848 = ~\WX7328_reg/NET0131  & ~\_2254__reg/NET0131  ;
  assign n6849 = \WX7328_reg/NET0131  & \_2254__reg/NET0131  ;
  assign n6850 = ~n6848 & ~n6849 ;
  assign n6851 = RESET_pad & ~n6850 ;
  assign n6852 = ~\WX9930_reg/NET0131  & ~\_2310__reg/NET0131  ;
  assign n6853 = \WX9930_reg/NET0131  & \_2310__reg/NET0131  ;
  assign n6854 = ~n6852 & ~n6853 ;
  assign n6855 = RESET_pad & ~n6854 ;
  assign n6856 = ~\WX2148_reg/NET0131  & ~\_2130__reg/NET0131  ;
  assign n6857 = \WX2148_reg/NET0131  & \_2130__reg/NET0131  ;
  assign n6858 = ~n6856 & ~n6857 ;
  assign n6859 = RESET_pad & ~n6858 ;
  assign n6860 = ~\WX7340_reg/NET0131  & ~\_2248__reg/NET0131  ;
  assign n6861 = \WX7340_reg/NET0131  & \_2248__reg/NET0131  ;
  assign n6862 = ~n6860 & ~n6861 ;
  assign n6863 = RESET_pad & ~n6862 ;
  assign n6864 = ~\WX6061_reg/NET0131  & ~\_2209__reg/NET0131  ;
  assign n6865 = \WX6061_reg/NET0131  & \_2209__reg/NET0131  ;
  assign n6866 = ~n6864 & ~n6865 ;
  assign n6867 = RESET_pad & ~n6866 ;
  assign n6868 = ~\WX8657_reg/NET0131  & ~\_2300__reg/NET0131  ;
  assign n6869 = \WX8657_reg/NET0131  & \_2300__reg/NET0131  ;
  assign n6870 = ~n6868 & ~n6869 ;
  assign n6871 = RESET_pad & ~n6870 ;
  assign n6872 = ~\WX2172_reg/NET0131  & ~\_2118__reg/NET0131  ;
  assign n6873 = \WX2172_reg/NET0131  & \_2118__reg/NET0131  ;
  assign n6874 = ~n6872 & ~n6873 ;
  assign n6875 = RESET_pad & ~n6874 ;
  assign n6876 = ~\WX8607_reg/NET0131  & ~\_2293__reg/NET0131  ;
  assign n6877 = \WX8607_reg/NET0131  & \_2293__reg/NET0131  ;
  assign n6878 = ~n6876 & ~n6877 ;
  assign n6879 = RESET_pad & ~n6878 ;
  assign n6880 = ~\WX899_reg/NET0131  & ~\_2108__reg/NET0131  ;
  assign n6881 = \WX899_reg/NET0131  & \_2108__reg/NET0131  ;
  assign n6882 = ~n6880 & ~n6881 ;
  assign n6883 = RESET_pad & ~n6882 ;
  assign n6884 = ~\WX897_reg/NET0131  & ~\_2077__reg/NET0131  ;
  assign n6885 = \WX897_reg/NET0131  & \_2077__reg/NET0131  ;
  assign n6886 = ~n6884 & ~n6885 ;
  assign n6887 = RESET_pad & ~n6886 ;
  assign n6888 = ~\WX895_reg/NET0131  & ~\_2078__reg/NET0131  ;
  assign n6889 = \WX895_reg/NET0131  & \_2078__reg/NET0131  ;
  assign n6890 = ~n6888 & ~n6889 ;
  assign n6891 = RESET_pad & ~n6890 ;
  assign n6892 = ~\WX893_reg/NET0131  & ~\_2079__reg/NET0131  ;
  assign n6893 = \WX893_reg/NET0131  & \_2079__reg/NET0131  ;
  assign n6894 = ~n6892 & ~n6893 ;
  assign n6895 = RESET_pad & ~n6894 ;
  assign n6896 = ~\WX889_reg/NET0131  & ~\_2081__reg/NET0131  ;
  assign n6897 = \WX889_reg/NET0131  & \_2081__reg/NET0131  ;
  assign n6898 = ~n6896 & ~n6897 ;
  assign n6899 = RESET_pad & ~n6898 ;
  assign n6900 = ~\WX887_reg/NET0131  & ~\_2082__reg/NET0131  ;
  assign n6901 = \WX887_reg/NET0131  & \_2082__reg/NET0131  ;
  assign n6902 = ~n6900 & ~n6901 ;
  assign n6903 = RESET_pad & ~n6902 ;
  assign n6904 = ~\WX883_reg/NET0131  & ~\_2084__reg/NET0131  ;
  assign n6905 = \WX883_reg/NET0131  & \_2084__reg/NET0131  ;
  assign n6906 = ~n6904 & ~n6905 ;
  assign n6907 = RESET_pad & ~n6906 ;
  assign n6908 = ~\WX881_reg/NET0131  & ~\_2085__reg/NET0131  ;
  assign n6909 = \WX881_reg/NET0131  & \_2085__reg/NET0131  ;
  assign n6910 = ~n6908 & ~n6909 ;
  assign n6911 = RESET_pad & ~n6910 ;
  assign n6912 = ~\WX875_reg/NET0131  & ~\_2088__reg/NET0131  ;
  assign n6913 = \WX875_reg/NET0131  & \_2088__reg/NET0131  ;
  assign n6914 = ~n6912 & ~n6913 ;
  assign n6915 = RESET_pad & ~n6914 ;
  assign n6916 = ~\WX873_reg/NET0131  & ~\_2089__reg/NET0131  ;
  assign n6917 = \WX873_reg/NET0131  & \_2089__reg/NET0131  ;
  assign n6918 = ~n6916 & ~n6917 ;
  assign n6919 = RESET_pad & ~n6918 ;
  assign n6920 = ~\WX869_reg/NET0131  & ~\_2091__reg/NET0131  ;
  assign n6921 = \WX869_reg/NET0131  & \_2091__reg/NET0131  ;
  assign n6922 = ~n6920 & ~n6921 ;
  assign n6923 = RESET_pad & ~n6922 ;
  assign n6924 = ~\WX865_reg/NET0131  & ~\_2093__reg/NET0131  ;
  assign n6925 = \WX865_reg/NET0131  & \_2093__reg/NET0131  ;
  assign n6926 = ~n6924 & ~n6925 ;
  assign n6927 = RESET_pad & ~n6926 ;
  assign n6928 = ~\WX863_reg/NET0131  & ~\_2094__reg/NET0131  ;
  assign n6929 = \WX863_reg/NET0131  & \_2094__reg/NET0131  ;
  assign n6930 = ~n6928 & ~n6929 ;
  assign n6931 = RESET_pad & ~n6930 ;
  assign n6932 = ~\WX855_reg/NET0131  & ~\_2098__reg/NET0131  ;
  assign n6933 = \WX855_reg/NET0131  & \_2098__reg/NET0131  ;
  assign n6934 = ~n6932 & ~n6933 ;
  assign n6935 = RESET_pad & ~n6934 ;
  assign n6936 = ~\WX851_reg/NET0131  & ~\_2100__reg/NET0131  ;
  assign n6937 = \WX851_reg/NET0131  & \_2100__reg/NET0131  ;
  assign n6938 = ~n6936 & ~n6937 ;
  assign n6939 = RESET_pad & ~n6938 ;
  assign n6940 = ~\WX845_reg/NET0131  & ~\_2103__reg/NET0131  ;
  assign n6941 = \WX845_reg/NET0131  & \_2103__reg/NET0131  ;
  assign n6942 = ~n6940 & ~n6941 ;
  assign n6943 = RESET_pad & ~n6942 ;
  assign n6944 = ~\WX843_reg/NET0131  & ~\_2104__reg/NET0131  ;
  assign n6945 = \WX843_reg/NET0131  & \_2104__reg/NET0131  ;
  assign n6946 = ~n6944 & ~n6945 ;
  assign n6947 = RESET_pad & ~n6946 ;
  assign n6948 = ~\WX841_reg/NET0131  & ~\_2105__reg/NET0131  ;
  assign n6949 = \WX841_reg/NET0131  & \_2105__reg/NET0131  ;
  assign n6950 = ~n6948 & ~n6949 ;
  assign n6951 = RESET_pad & ~n6950 ;
  assign n6952 = ~\WX839_reg/NET0131  & ~\_2106__reg/NET0131  ;
  assign n6953 = \WX839_reg/NET0131  & \_2106__reg/NET0131  ;
  assign n6954 = ~n6952 & ~n6953 ;
  assign n6955 = RESET_pad & ~n6954 ;
  assign n6956 = ~\WX2192_reg/NET0131  & ~\_2140__reg/NET0131  ;
  assign n6957 = \WX2192_reg/NET0131  & \_2140__reg/NET0131  ;
  assign n6958 = ~n6956 & ~n6957 ;
  assign n6959 = RESET_pad & ~n6958 ;
  assign n6960 = ~\WX2190_reg/NET0131  & ~\_2109__reg/NET0131  ;
  assign n6961 = \WX2190_reg/NET0131  & \_2109__reg/NET0131  ;
  assign n6962 = ~n6960 & ~n6961 ;
  assign n6963 = RESET_pad & ~n6962 ;
  assign n6964 = ~\WX2188_reg/NET0131  & ~\_2110__reg/NET0131  ;
  assign n6965 = \WX2188_reg/NET0131  & \_2110__reg/NET0131  ;
  assign n6966 = ~n6964 & ~n6965 ;
  assign n6967 = RESET_pad & ~n6966 ;
  assign n6968 = ~\WX2186_reg/NET0131  & ~\_2111__reg/NET0131  ;
  assign n6969 = \WX2186_reg/NET0131  & \_2111__reg/NET0131  ;
  assign n6970 = ~n6968 & ~n6969 ;
  assign n6971 = RESET_pad & ~n6970 ;
  assign n6972 = ~\WX2182_reg/NET0131  & ~\_2113__reg/NET0131  ;
  assign n6973 = \WX2182_reg/NET0131  & \_2113__reg/NET0131  ;
  assign n6974 = ~n6972 & ~n6973 ;
  assign n6975 = RESET_pad & ~n6974 ;
  assign n6976 = ~\WX2180_reg/NET0131  & ~\_2114__reg/NET0131  ;
  assign n6977 = \WX2180_reg/NET0131  & \_2114__reg/NET0131  ;
  assign n6978 = ~n6976 & ~n6977 ;
  assign n6979 = RESET_pad & ~n6978 ;
  assign n6980 = ~\WX2174_reg/NET0131  & ~\_2117__reg/NET0131  ;
  assign n6981 = \WX2174_reg/NET0131  & \_2117__reg/NET0131  ;
  assign n6982 = ~n6980 & ~n6981 ;
  assign n6983 = RESET_pad & ~n6982 ;
  assign n6984 = ~\WX2168_reg/NET0131  & ~\_2120__reg/NET0131  ;
  assign n6985 = \WX2168_reg/NET0131  & \_2120__reg/NET0131  ;
  assign n6986 = ~n6984 & ~n6985 ;
  assign n6987 = RESET_pad & ~n6986 ;
  assign n6988 = ~\WX2166_reg/NET0131  & ~\_2121__reg/NET0131  ;
  assign n6989 = \WX2166_reg/NET0131  & \_2121__reg/NET0131  ;
  assign n6990 = ~n6988 & ~n6989 ;
  assign n6991 = RESET_pad & ~n6990 ;
  assign n6992 = ~\WX2164_reg/NET0131  & ~\_2122__reg/NET0131  ;
  assign n6993 = \WX2164_reg/NET0131  & \_2122__reg/NET0131  ;
  assign n6994 = ~n6992 & ~n6993 ;
  assign n6995 = RESET_pad & ~n6994 ;
  assign n6996 = ~\WX2162_reg/NET0131  & ~\_2123__reg/NET0131  ;
  assign n6997 = \WX2162_reg/NET0131  & \_2123__reg/NET0131  ;
  assign n6998 = ~n6996 & ~n6997 ;
  assign n6999 = RESET_pad & ~n6998 ;
  assign n7000 = ~\WX2158_reg/NET0131  & ~\_2125__reg/NET0131  ;
  assign n7001 = \WX2158_reg/NET0131  & \_2125__reg/NET0131  ;
  assign n7002 = ~n7000 & ~n7001 ;
  assign n7003 = RESET_pad & ~n7002 ;
  assign n7004 = ~\WX2156_reg/NET0131  & ~\_2126__reg/NET0131  ;
  assign n7005 = \WX2156_reg/NET0131  & \_2126__reg/NET0131  ;
  assign n7006 = ~n7004 & ~n7005 ;
  assign n7007 = RESET_pad & ~n7006 ;
  assign n7008 = ~\WX2154_reg/NET0131  & ~\_2127__reg/NET0131  ;
  assign n7009 = \WX2154_reg/NET0131  & \_2127__reg/NET0131  ;
  assign n7010 = ~n7008 & ~n7009 ;
  assign n7011 = RESET_pad & ~n7010 ;
  assign n7012 = ~\WX2146_reg/NET0131  & ~\_2131__reg/NET0131  ;
  assign n7013 = \WX2146_reg/NET0131  & \_2131__reg/NET0131  ;
  assign n7014 = ~n7012 & ~n7013 ;
  assign n7015 = RESET_pad & ~n7014 ;
  assign n7016 = ~\WX2144_reg/NET0131  & ~\_2132__reg/NET0131  ;
  assign n7017 = \WX2144_reg/NET0131  & \_2132__reg/NET0131  ;
  assign n7018 = ~n7016 & ~n7017 ;
  assign n7019 = RESET_pad & ~n7018 ;
  assign n7020 = ~\WX2142_reg/NET0131  & ~\_2133__reg/NET0131  ;
  assign n7021 = \WX2142_reg/NET0131  & \_2133__reg/NET0131  ;
  assign n7022 = ~n7020 & ~n7021 ;
  assign n7023 = RESET_pad & ~n7022 ;
  assign n7024 = ~\WX2138_reg/NET0131  & ~\_2135__reg/NET0131  ;
  assign n7025 = \WX2138_reg/NET0131  & \_2135__reg/NET0131  ;
  assign n7026 = ~n7024 & ~n7025 ;
  assign n7027 = RESET_pad & ~n7026 ;
  assign n7028 = ~\WX2134_reg/NET0131  & ~\_2137__reg/NET0131  ;
  assign n7029 = \WX2134_reg/NET0131  & \_2137__reg/NET0131  ;
  assign n7030 = ~n7028 & ~n7029 ;
  assign n7031 = RESET_pad & ~n7030 ;
  assign n7032 = ~\WX7348_reg/NET0131  & ~\_2244__reg/NET0131  ;
  assign n7033 = \WX7348_reg/NET0131  & \_2244__reg/NET0131  ;
  assign n7034 = ~n7032 & ~n7033 ;
  assign n7035 = RESET_pad & ~n7034 ;
  assign n7036 = ~\WX3483_reg/NET0131  & ~\_2141__reg/NET0131  ;
  assign n7037 = \WX3483_reg/NET0131  & \_2141__reg/NET0131  ;
  assign n7038 = ~n7036 & ~n7037 ;
  assign n7039 = RESET_pad & ~n7038 ;
  assign n7040 = ~\WX3481_reg/NET0131  & ~\_2142__reg/NET0131  ;
  assign n7041 = \WX3481_reg/NET0131  & \_2142__reg/NET0131  ;
  assign n7042 = ~n7040 & ~n7041 ;
  assign n7043 = RESET_pad & ~n7042 ;
  assign n7044 = ~\WX3479_reg/NET0131  & ~\_2143__reg/NET0131  ;
  assign n7045 = \WX3479_reg/NET0131  & \_2143__reg/NET0131  ;
  assign n7046 = ~n7044 & ~n7045 ;
  assign n7047 = RESET_pad & ~n7046 ;
  assign n7048 = ~\WX3473_reg/NET0131  & ~\_2146__reg/NET0131  ;
  assign n7049 = \WX3473_reg/NET0131  & \_2146__reg/NET0131  ;
  assign n7050 = ~n7048 & ~n7049 ;
  assign n7051 = RESET_pad & ~n7050 ;
  assign n7052 = ~\WX3471_reg/NET0131  & ~\_2147__reg/NET0131  ;
  assign n7053 = \WX3471_reg/NET0131  & \_2147__reg/NET0131  ;
  assign n7054 = ~n7052 & ~n7053 ;
  assign n7055 = RESET_pad & ~n7054 ;
  assign n7056 = ~\WX3469_reg/NET0131  & ~\_2148__reg/NET0131  ;
  assign n7057 = \WX3469_reg/NET0131  & \_2148__reg/NET0131  ;
  assign n7058 = ~n7056 & ~n7057 ;
  assign n7059 = RESET_pad & ~n7058 ;
  assign n7060 = ~\WX3465_reg/NET0131  & ~\_2150__reg/NET0131  ;
  assign n7061 = \WX3465_reg/NET0131  & \_2150__reg/NET0131  ;
  assign n7062 = ~n7060 & ~n7061 ;
  assign n7063 = RESET_pad & ~n7062 ;
  assign n7064 = ~\WX3459_reg/NET0131  & ~\_2153__reg/NET0131  ;
  assign n7065 = \WX3459_reg/NET0131  & \_2153__reg/NET0131  ;
  assign n7066 = ~n7064 & ~n7065 ;
  assign n7067 = RESET_pad & ~n7066 ;
  assign n7068 = ~\WX3457_reg/NET0131  & ~\_2154__reg/NET0131  ;
  assign n7069 = \WX3457_reg/NET0131  & \_2154__reg/NET0131  ;
  assign n7070 = ~n7068 & ~n7069 ;
  assign n7071 = RESET_pad & ~n7070 ;
  assign n7072 = ~\WX3455_reg/NET0131  & ~\_2155__reg/NET0131  ;
  assign n7073 = \WX3455_reg/NET0131  & \_2155__reg/NET0131  ;
  assign n7074 = ~n7072 & ~n7073 ;
  assign n7075 = RESET_pad & ~n7074 ;
  assign n7076 = ~\WX3451_reg/NET0131  & ~\_2157__reg/NET0131  ;
  assign n7077 = \WX3451_reg/NET0131  & \_2157__reg/NET0131  ;
  assign n7078 = ~n7076 & ~n7077 ;
  assign n7079 = RESET_pad & ~n7078 ;
  assign n7080 = ~\WX3449_reg/NET0131  & ~\_2158__reg/NET0131  ;
  assign n7081 = \WX3449_reg/NET0131  & \_2158__reg/NET0131  ;
  assign n7082 = ~n7080 & ~n7081 ;
  assign n7083 = RESET_pad & ~n7082 ;
  assign n7084 = ~\WX3445_reg/NET0131  & ~\_2160__reg/NET0131  ;
  assign n7085 = \WX3445_reg/NET0131  & \_2160__reg/NET0131  ;
  assign n7086 = ~n7084 & ~n7085 ;
  assign n7087 = RESET_pad & ~n7086 ;
  assign n7088 = ~\WX3443_reg/NET0131  & ~\_2161__reg/NET0131  ;
  assign n7089 = \WX3443_reg/NET0131  & \_2161__reg/NET0131  ;
  assign n7090 = ~n7088 & ~n7089 ;
  assign n7091 = RESET_pad & ~n7090 ;
  assign n7092 = ~\WX3441_reg/NET0131  & ~\_2162__reg/NET0131  ;
  assign n7093 = \WX3441_reg/NET0131  & \_2162__reg/NET0131  ;
  assign n7094 = ~n7092 & ~n7093 ;
  assign n7095 = RESET_pad & ~n7094 ;
  assign n7096 = ~\WX3439_reg/NET0131  & ~\_2163__reg/NET0131  ;
  assign n7097 = \WX3439_reg/NET0131  & \_2163__reg/NET0131  ;
  assign n7098 = ~n7096 & ~n7097 ;
  assign n7099 = RESET_pad & ~n7098 ;
  assign n7100 = ~\WX3437_reg/NET0131  & ~\_2164__reg/NET0131  ;
  assign n7101 = \WX3437_reg/NET0131  & \_2164__reg/NET0131  ;
  assign n7102 = ~n7100 & ~n7101 ;
  assign n7103 = RESET_pad & ~n7102 ;
  assign n7104 = ~\WX3435_reg/NET0131  & ~\_2165__reg/NET0131  ;
  assign n7105 = \WX3435_reg/NET0131  & \_2165__reg/NET0131  ;
  assign n7106 = ~n7104 & ~n7105 ;
  assign n7107 = RESET_pad & ~n7106 ;
  assign n7108 = ~\WX3433_reg/NET0131  & ~\_2166__reg/NET0131  ;
  assign n7109 = \WX3433_reg/NET0131  & \_2166__reg/NET0131  ;
  assign n7110 = ~n7108 & ~n7109 ;
  assign n7111 = RESET_pad & ~n7110 ;
  assign n7112 = ~\WX3431_reg/NET0131  & ~\_2167__reg/NET0131  ;
  assign n7113 = \WX3431_reg/NET0131  & \_2167__reg/NET0131  ;
  assign n7114 = ~n7112 & ~n7113 ;
  assign n7115 = RESET_pad & ~n7114 ;
  assign n7116 = ~\WX3429_reg/NET0131  & ~\_2168__reg/NET0131  ;
  assign n7117 = \WX3429_reg/NET0131  & \_2168__reg/NET0131  ;
  assign n7118 = ~n7116 & ~n7117 ;
  assign n7119 = RESET_pad & ~n7118 ;
  assign n7120 = ~\WX3423_reg/NET0131  & ~\_2171__reg/NET0131  ;
  assign n7121 = \WX3423_reg/NET0131  & \_2171__reg/NET0131  ;
  assign n7122 = ~n7120 & ~n7121 ;
  assign n7123 = RESET_pad & ~n7122 ;
  assign n7124 = ~\WX4778_reg/NET0131  & ~\_2204__reg/NET0131  ;
  assign n7125 = \WX4778_reg/NET0131  & \_2204__reg/NET0131  ;
  assign n7126 = ~n7124 & ~n7125 ;
  assign n7127 = RESET_pad & ~n7126 ;
  assign n7128 = ~\WX4776_reg/NET0131  & ~\_2173__reg/NET0131  ;
  assign n7129 = \WX4776_reg/NET0131  & \_2173__reg/NET0131  ;
  assign n7130 = ~n7128 & ~n7129 ;
  assign n7131 = RESET_pad & ~n7130 ;
  assign n7132 = ~\WX4774_reg/NET0131  & ~\_2174__reg/NET0131  ;
  assign n7133 = \WX4774_reg/NET0131  & \_2174__reg/NET0131  ;
  assign n7134 = ~n7132 & ~n7133 ;
  assign n7135 = RESET_pad & ~n7134 ;
  assign n7136 = ~\WX4772_reg/NET0131  & ~\_2175__reg/NET0131  ;
  assign n7137 = \WX4772_reg/NET0131  & \_2175__reg/NET0131  ;
  assign n7138 = ~n7136 & ~n7137 ;
  assign n7139 = RESET_pad & ~n7138 ;
  assign n7140 = ~\WX7316_reg/NET0131  & ~\_2260__reg/NET0131  ;
  assign n7141 = \WX7316_reg/NET0131  & \_2260__reg/NET0131  ;
  assign n7142 = ~n7140 & ~n7141 ;
  assign n7143 = RESET_pad & ~n7142 ;
  assign n7144 = ~\WX4768_reg/NET0131  & ~\_2177__reg/NET0131  ;
  assign n7145 = \WX4768_reg/NET0131  & \_2177__reg/NET0131  ;
  assign n7146 = ~n7144 & ~n7145 ;
  assign n7147 = RESET_pad & ~n7146 ;
  assign n7148 = ~\WX4766_reg/NET0131  & ~\_2178__reg/NET0131  ;
  assign n7149 = \WX4766_reg/NET0131  & \_2178__reg/NET0131  ;
  assign n7150 = ~n7148 & ~n7149 ;
  assign n7151 = RESET_pad & ~n7150 ;
  assign n7152 = ~\WX4764_reg/NET0131  & ~\_2179__reg/NET0131  ;
  assign n7153 = \WX4764_reg/NET0131  & \_2179__reg/NET0131  ;
  assign n7154 = ~n7152 & ~n7153 ;
  assign n7155 = RESET_pad & ~n7154 ;
  assign n7156 = ~\WX4760_reg/NET0131  & ~\_2181__reg/NET0131  ;
  assign n7157 = \WX4760_reg/NET0131  & \_2181__reg/NET0131  ;
  assign n7158 = ~n7156 & ~n7157 ;
  assign n7159 = RESET_pad & ~n7158 ;
  assign n7160 = ~\WX4758_reg/NET0131  & ~\_2182__reg/NET0131  ;
  assign n7161 = \WX4758_reg/NET0131  & \_2182__reg/NET0131  ;
  assign n7162 = ~n7160 & ~n7161 ;
  assign n7163 = RESET_pad & ~n7162 ;
  assign n7164 = ~\WX4754_reg/NET0131  & ~\_2184__reg/NET0131  ;
  assign n7165 = \WX4754_reg/NET0131  & \_2184__reg/NET0131  ;
  assign n7166 = ~n7164 & ~n7165 ;
  assign n7167 = RESET_pad & ~n7166 ;
  assign n7168 = ~\WX4752_reg/NET0131  & ~\_2185__reg/NET0131  ;
  assign n7169 = \WX4752_reg/NET0131  & \_2185__reg/NET0131  ;
  assign n7170 = ~n7168 & ~n7169 ;
  assign n7171 = RESET_pad & ~n7170 ;
  assign n7172 = ~\WX4750_reg/NET0131  & ~\_2186__reg/NET0131  ;
  assign n7173 = \WX4750_reg/NET0131  & \_2186__reg/NET0131  ;
  assign n7174 = ~n7172 & ~n7173 ;
  assign n7175 = RESET_pad & ~n7174 ;
  assign n7176 = ~\WX4748_reg/NET0131  & ~\_2187__reg/NET0131  ;
  assign n7177 = \WX4748_reg/NET0131  & \_2187__reg/NET0131  ;
  assign n7178 = ~n7176 & ~n7177 ;
  assign n7179 = RESET_pad & ~n7178 ;
  assign n7180 = ~\WX4744_reg/NET0131  & ~\_2189__reg/NET0131  ;
  assign n7181 = \WX4744_reg/NET0131  & \_2189__reg/NET0131  ;
  assign n7182 = ~n7180 & ~n7181 ;
  assign n7183 = RESET_pad & ~n7182 ;
  assign n7184 = ~\WX4742_reg/NET0131  & ~\_2190__reg/NET0131  ;
  assign n7185 = \WX4742_reg/NET0131  & \_2190__reg/NET0131  ;
  assign n7186 = ~n7184 & ~n7185 ;
  assign n7187 = RESET_pad & ~n7186 ;
  assign n7188 = ~\WX4740_reg/NET0131  & ~\_2191__reg/NET0131  ;
  assign n7189 = \WX4740_reg/NET0131  & \_2191__reg/NET0131  ;
  assign n7190 = ~n7188 & ~n7189 ;
  assign n7191 = RESET_pad & ~n7190 ;
  assign n7192 = ~\WX4738_reg/NET0131  & ~\_2192__reg/NET0131  ;
  assign n7193 = \WX4738_reg/NET0131  & \_2192__reg/NET0131  ;
  assign n7194 = ~n7192 & ~n7193 ;
  assign n7195 = RESET_pad & ~n7194 ;
  assign n7196 = ~\WX4736_reg/NET0131  & ~\_2193__reg/NET0131  ;
  assign n7197 = \WX4736_reg/NET0131  & \_2193__reg/NET0131  ;
  assign n7198 = ~n7196 & ~n7197 ;
  assign n7199 = RESET_pad & ~n7198 ;
  assign n7200 = ~\WX4734_reg/NET0131  & ~\_2194__reg/NET0131  ;
  assign n7201 = \WX4734_reg/NET0131  & \_2194__reg/NET0131  ;
  assign n7202 = ~n7200 & ~n7201 ;
  assign n7203 = RESET_pad & ~n7202 ;
  assign n7204 = ~\WX4732_reg/NET0131  & ~\_2195__reg/NET0131  ;
  assign n7205 = \WX4732_reg/NET0131  & \_2195__reg/NET0131  ;
  assign n7206 = ~n7204 & ~n7205 ;
  assign n7207 = RESET_pad & ~n7206 ;
  assign n7208 = ~\WX4730_reg/NET0131  & ~\_2196__reg/NET0131  ;
  assign n7209 = \WX4730_reg/NET0131  & \_2196__reg/NET0131  ;
  assign n7210 = ~n7208 & ~n7209 ;
  assign n7211 = RESET_pad & ~n7210 ;
  assign n7212 = ~\WX4724_reg/NET0131  & ~\_2199__reg/NET0131  ;
  assign n7213 = \WX4724_reg/NET0131  & \_2199__reg/NET0131  ;
  assign n7214 = ~n7212 & ~n7213 ;
  assign n7215 = RESET_pad & ~n7214 ;
  assign n7216 = ~\WX4722_reg/NET0131  & ~\_2200__reg/NET0131  ;
  assign n7217 = \WX4722_reg/NET0131  & \_2200__reg/NET0131  ;
  assign n7218 = ~n7216 & ~n7217 ;
  assign n7219 = RESET_pad & ~n7218 ;
  assign n7220 = ~\WX4720_reg/NET0131  & ~\_2201__reg/NET0131  ;
  assign n7221 = \WX4720_reg/NET0131  & \_2201__reg/NET0131  ;
  assign n7222 = ~n7220 & ~n7221 ;
  assign n7223 = RESET_pad & ~n7222 ;
  assign n7224 = ~\WX4718_reg/NET0131  & ~\_2202__reg/NET0131  ;
  assign n7225 = \WX4718_reg/NET0131  & \_2202__reg/NET0131  ;
  assign n7226 = ~n7224 & ~n7225 ;
  assign n7227 = RESET_pad & ~n7226 ;
  assign n7228 = ~\WX4716_reg/NET0131  & ~\_2203__reg/NET0131  ;
  assign n7229 = \WX4716_reg/NET0131  & \_2203__reg/NET0131  ;
  assign n7230 = ~n7228 & ~n7229 ;
  assign n7231 = RESET_pad & ~n7230 ;
  assign n7232 = ~\WX6071_reg/NET0131  & ~\_2236__reg/NET0131  ;
  assign n7233 = \WX6071_reg/NET0131  & \_2236__reg/NET0131  ;
  assign n7234 = ~n7232 & ~n7233 ;
  assign n7235 = RESET_pad & ~n7234 ;
  assign n7236 = ~\WX6067_reg/NET0131  & ~\_2206__reg/NET0131  ;
  assign n7237 = \WX6067_reg/NET0131  & \_2206__reg/NET0131  ;
  assign n7238 = ~n7236 & ~n7237 ;
  assign n7239 = RESET_pad & ~n7238 ;
  assign n7240 = ~\WX6065_reg/NET0131  & ~\_2207__reg/NET0131  ;
  assign n7241 = \WX6065_reg/NET0131  & \_2207__reg/NET0131  ;
  assign n7242 = ~n7240 & ~n7241 ;
  assign n7243 = RESET_pad & ~n7242 ;
  assign n7244 = ~\WX6059_reg/NET0131  & ~\_2210__reg/NET0131  ;
  assign n7245 = \WX6059_reg/NET0131  & \_2210__reg/NET0131  ;
  assign n7246 = ~n7244 & ~n7245 ;
  assign n7247 = RESET_pad & ~n7246 ;
  assign n7248 = ~\WX6057_reg/NET0131  & ~\_2211__reg/NET0131  ;
  assign n7249 = \WX6057_reg/NET0131  & \_2211__reg/NET0131  ;
  assign n7250 = ~n7248 & ~n7249 ;
  assign n7251 = RESET_pad & ~n7250 ;
  assign n7252 = ~\WX6055_reg/NET0131  & ~\_2212__reg/NET0131  ;
  assign n7253 = \WX6055_reg/NET0131  & \_2212__reg/NET0131  ;
  assign n7254 = ~n7252 & ~n7253 ;
  assign n7255 = RESET_pad & ~n7254 ;
  assign n7256 = ~\WX6053_reg/NET0131  & ~\_2213__reg/NET0131  ;
  assign n7257 = \WX6053_reg/NET0131  & \_2213__reg/NET0131  ;
  assign n7258 = ~n7256 & ~n7257 ;
  assign n7259 = RESET_pad & ~n7258 ;
  assign n7260 = ~\WX6051_reg/NET0131  & ~\_2214__reg/NET0131  ;
  assign n7261 = \WX6051_reg/NET0131  & \_2214__reg/NET0131  ;
  assign n7262 = ~n7260 & ~n7261 ;
  assign n7263 = RESET_pad & ~n7262 ;
  assign n7264 = ~\WX6047_reg/NET0131  & ~\_2216__reg/NET0131  ;
  assign n7265 = \WX6047_reg/NET0131  & \_2216__reg/NET0131  ;
  assign n7266 = ~n7264 & ~n7265 ;
  assign n7267 = RESET_pad & ~n7266 ;
  assign n7268 = ~\WX6045_reg/NET0131  & ~\_2217__reg/NET0131  ;
  assign n7269 = \WX6045_reg/NET0131  & \_2217__reg/NET0131  ;
  assign n7270 = ~n7268 & ~n7269 ;
  assign n7271 = RESET_pad & ~n7270 ;
  assign n7272 = ~\WX6035_reg/NET0131  & ~\_2222__reg/NET0131  ;
  assign n7273 = \WX6035_reg/NET0131  & \_2222__reg/NET0131  ;
  assign n7274 = ~n7272 & ~n7273 ;
  assign n7275 = RESET_pad & ~n7274 ;
  assign n7276 = ~\WX6033_reg/NET0131  & ~\_2223__reg/NET0131  ;
  assign n7277 = \WX6033_reg/NET0131  & \_2223__reg/NET0131  ;
  assign n7278 = ~n7276 & ~n7277 ;
  assign n7279 = RESET_pad & ~n7278 ;
  assign n7280 = ~\WX6031_reg/NET0131  & ~\_2224__reg/NET0131  ;
  assign n7281 = \WX6031_reg/NET0131  & \_2224__reg/NET0131  ;
  assign n7282 = ~n7280 & ~n7281 ;
  assign n7283 = RESET_pad & ~n7282 ;
  assign n7284 = ~\WX6029_reg/NET0131  & ~\_2225__reg/NET0131  ;
  assign n7285 = \WX6029_reg/NET0131  & \_2225__reg/NET0131  ;
  assign n7286 = ~n7284 & ~n7285 ;
  assign n7287 = RESET_pad & ~n7286 ;
  assign n7288 = ~\WX6023_reg/NET0131  & ~\_2228__reg/NET0131  ;
  assign n7289 = \WX6023_reg/NET0131  & \_2228__reg/NET0131  ;
  assign n7290 = ~n7288 & ~n7289 ;
  assign n7291 = RESET_pad & ~n7290 ;
  assign n7292 = ~\WX6021_reg/NET0131  & ~\_2229__reg/NET0131  ;
  assign n7293 = \WX6021_reg/NET0131  & \_2229__reg/NET0131  ;
  assign n7294 = ~n7292 & ~n7293 ;
  assign n7295 = RESET_pad & ~n7294 ;
  assign n7296 = ~\WX6019_reg/NET0131  & ~\_2230__reg/NET0131  ;
  assign n7297 = \WX6019_reg/NET0131  & \_2230__reg/NET0131  ;
  assign n7298 = ~n7296 & ~n7297 ;
  assign n7299 = RESET_pad & ~n7298 ;
  assign n7300 = ~\WX6015_reg/NET0131  & ~\_2232__reg/NET0131  ;
  assign n7301 = \WX6015_reg/NET0131  & \_2232__reg/NET0131  ;
  assign n7302 = ~n7300 & ~n7301 ;
  assign n7303 = RESET_pad & ~n7302 ;
  assign n7304 = ~\WX6011_reg/NET0131  & ~\_2234__reg/NET0131  ;
  assign n7305 = \WX6011_reg/NET0131  & \_2234__reg/NET0131  ;
  assign n7306 = ~n7304 & ~n7305 ;
  assign n7307 = RESET_pad & ~n7306 ;
  assign n7308 = ~\WX6009_reg/NET0131  & ~\_2235__reg/NET0131  ;
  assign n7309 = \WX6009_reg/NET0131  & \_2235__reg/NET0131  ;
  assign n7310 = ~n7308 & ~n7309 ;
  assign n7311 = RESET_pad & ~n7310 ;
  assign n7312 = ~\WX7364_reg/NET0131  & ~\_2268__reg/NET0131  ;
  assign n7313 = \WX7364_reg/NET0131  & \_2268__reg/NET0131  ;
  assign n7314 = ~n7312 & ~n7313 ;
  assign n7315 = RESET_pad & ~n7314 ;
  assign n7316 = ~\WX7360_reg/NET0131  & ~\_2238__reg/NET0131  ;
  assign n7317 = \WX7360_reg/NET0131  & \_2238__reg/NET0131  ;
  assign n7318 = ~n7316 & ~n7317 ;
  assign n7319 = RESET_pad & ~n7318 ;
  assign n7320 = ~\WX7358_reg/NET0131  & ~\_2239__reg/NET0131  ;
  assign n7321 = \WX7358_reg/NET0131  & \_2239__reg/NET0131  ;
  assign n7322 = ~n7320 & ~n7321 ;
  assign n7323 = RESET_pad & ~n7322 ;
  assign n7324 = ~\WX7354_reg/NET0131  & ~\_2241__reg/NET0131  ;
  assign n7325 = \WX7354_reg/NET0131  & \_2241__reg/NET0131  ;
  assign n7326 = ~n7324 & ~n7325 ;
  assign n7327 = RESET_pad & ~n7326 ;
  assign n7328 = ~\WX7352_reg/NET0131  & ~\_2242__reg/NET0131  ;
  assign n7329 = \WX7352_reg/NET0131  & \_2242__reg/NET0131  ;
  assign n7330 = ~n7328 & ~n7329 ;
  assign n7331 = RESET_pad & ~n7330 ;
  assign n7332 = ~\WX6025_reg/NET0131  & ~\_2227__reg/NET0131  ;
  assign n7333 = \WX6025_reg/NET0131  & \_2227__reg/NET0131  ;
  assign n7334 = ~n7332 & ~n7333 ;
  assign n7335 = RESET_pad & ~n7334 ;
  assign n7336 = ~\WX8647_reg/NET0131  & ~\_2273__reg/NET0131  ;
  assign n7337 = \WX8647_reg/NET0131  & \_2273__reg/NET0131  ;
  assign n7338 = ~n7336 & ~n7337 ;
  assign n7339 = RESET_pad & ~n7338 ;
  assign n7340 = ~\WX7336_reg/NET0131  & ~\_2250__reg/NET0131  ;
  assign n7341 = \WX7336_reg/NET0131  & \_2250__reg/NET0131  ;
  assign n7342 = ~n7340 & ~n7341 ;
  assign n7343 = RESET_pad & ~n7342 ;
  assign n7344 = ~\WX7330_reg/NET0131  & ~\_2253__reg/NET0131  ;
  assign n7345 = \WX7330_reg/NET0131  & \_2253__reg/NET0131  ;
  assign n7346 = ~n7344 & ~n7345 ;
  assign n7347 = RESET_pad & ~n7346 ;
  assign n7348 = ~\WX7326_reg/NET0131  & ~\_2255__reg/NET0131  ;
  assign n7349 = \WX7326_reg/NET0131  & \_2255__reg/NET0131  ;
  assign n7350 = ~n7348 & ~n7349 ;
  assign n7351 = RESET_pad & ~n7350 ;
  assign n7352 = ~\WX7322_reg/NET0131  & ~\_2257__reg/NET0131  ;
  assign n7353 = \WX7322_reg/NET0131  & \_2257__reg/NET0131  ;
  assign n7354 = ~n7352 & ~n7353 ;
  assign n7355 = RESET_pad & ~n7354 ;
  assign n7356 = ~\WX7320_reg/NET0131  & ~\_2258__reg/NET0131  ;
  assign n7357 = \WX7320_reg/NET0131  & \_2258__reg/NET0131  ;
  assign n7358 = ~n7356 & ~n7357 ;
  assign n7359 = RESET_pad & ~n7358 ;
  assign n7360 = ~\WX7318_reg/NET0131  & ~\_2259__reg/NET0131  ;
  assign n7361 = \WX7318_reg/NET0131  & \_2259__reg/NET0131  ;
  assign n7362 = ~n7360 & ~n7361 ;
  assign n7363 = RESET_pad & ~n7362 ;
  assign n7364 = ~\WX6069_reg/NET0131  & ~\_2205__reg/NET0131  ;
  assign n7365 = \WX6069_reg/NET0131  & \_2205__reg/NET0131  ;
  assign n7366 = ~n7364 & ~n7365 ;
  assign n7367 = RESET_pad & ~n7366 ;
  assign n7368 = ~\WX7314_reg/NET0131  & ~\_2261__reg/NET0131  ;
  assign n7369 = \WX7314_reg/NET0131  & \_2261__reg/NET0131  ;
  assign n7370 = ~n7368 & ~n7369 ;
  assign n7371 = RESET_pad & ~n7370 ;
  assign n7372 = ~\WX6017_reg/NET0131  & ~\_2231__reg/NET0131  ;
  assign n7373 = \WX6017_reg/NET0131  & \_2231__reg/NET0131  ;
  assign n7374 = ~n7372 & ~n7373 ;
  assign n7375 = RESET_pad & ~n7374 ;
  assign n7376 = ~\WX6027_reg/NET0131  & ~\_2226__reg/NET0131  ;
  assign n7377 = \WX6027_reg/NET0131  & \_2226__reg/NET0131  ;
  assign n7378 = ~n7376 & ~n7377 ;
  assign n7379 = RESET_pad & ~n7378 ;
  assign n7380 = ~\WX7306_reg/NET0131  & ~\_2265__reg/NET0131  ;
  assign n7381 = \WX7306_reg/NET0131  & \_2265__reg/NET0131  ;
  assign n7382 = ~n7380 & ~n7381 ;
  assign n7383 = RESET_pad & ~n7382 ;
  assign n7384 = ~\WX7302_reg/NET0131  & ~\_2267__reg/NET0131  ;
  assign n7385 = \WX7302_reg/NET0131  & \_2267__reg/NET0131  ;
  assign n7386 = ~n7384 & ~n7385 ;
  assign n7387 = RESET_pad & ~n7386 ;
  assign n7388 = ~\WX8655_reg/NET0131  & ~\_2269__reg/NET0131  ;
  assign n7389 = \WX8655_reg/NET0131  & \_2269__reg/NET0131  ;
  assign n7390 = ~n7388 & ~n7389 ;
  assign n7391 = RESET_pad & ~n7390 ;
  assign n7392 = ~\WX8653_reg/NET0131  & ~\_2270__reg/NET0131  ;
  assign n7393 = \WX8653_reg/NET0131  & \_2270__reg/NET0131  ;
  assign n7394 = ~n7392 & ~n7393 ;
  assign n7395 = RESET_pad & ~n7394 ;
  assign n7396 = ~\WX8651_reg/NET0131  & ~\_2271__reg/NET0131  ;
  assign n7397 = \WX8651_reg/NET0131  & \_2271__reg/NET0131  ;
  assign n7398 = ~n7396 & ~n7397 ;
  assign n7399 = RESET_pad & ~n7398 ;
  assign n7400 = ~\WX8645_reg/NET0131  & ~\_2274__reg/NET0131  ;
  assign n7401 = \WX8645_reg/NET0131  & \_2274__reg/NET0131  ;
  assign n7402 = ~n7400 & ~n7401 ;
  assign n7403 = RESET_pad & ~n7402 ;
  assign n7404 = ~\WX8641_reg/NET0131  & ~\_2276__reg/NET0131  ;
  assign n7405 = \WX8641_reg/NET0131  & \_2276__reg/NET0131  ;
  assign n7406 = ~n7404 & ~n7405 ;
  assign n7407 = RESET_pad & ~n7406 ;
  assign n7408 = ~\WX8637_reg/NET0131  & ~\_2278__reg/NET0131  ;
  assign n7409 = \WX8637_reg/NET0131  & \_2278__reg/NET0131  ;
  assign n7410 = ~n7408 & ~n7409 ;
  assign n7411 = RESET_pad & ~n7410 ;
  assign n7412 = ~\WX8631_reg/NET0131  & ~\_2281__reg/NET0131  ;
  assign n7413 = \WX8631_reg/NET0131  & \_2281__reg/NET0131  ;
  assign n7414 = ~n7412 & ~n7413 ;
  assign n7415 = RESET_pad & ~n7414 ;
  assign n7416 = ~\WX8629_reg/NET0131  & ~\_2282__reg/NET0131  ;
  assign n7417 = \WX8629_reg/NET0131  & \_2282__reg/NET0131  ;
  assign n7418 = ~n7416 & ~n7417 ;
  assign n7419 = RESET_pad & ~n7418 ;
  assign n7420 = ~\WX8627_reg/NET0131  & ~\_2283__reg/NET0131  ;
  assign n7421 = \WX8627_reg/NET0131  & \_2283__reg/NET0131  ;
  assign n7422 = ~n7420 & ~n7421 ;
  assign n7423 = RESET_pad & ~n7422 ;
  assign n7424 = ~\WX8621_reg/NET0131  & ~\_2286__reg/NET0131  ;
  assign n7425 = \WX8621_reg/NET0131  & \_2286__reg/NET0131  ;
  assign n7426 = ~n7424 & ~n7425 ;
  assign n7427 = RESET_pad & ~n7426 ;
  assign n7428 = ~\WX8617_reg/NET0131  & ~\_2288__reg/NET0131  ;
  assign n7429 = \WX8617_reg/NET0131  & \_2288__reg/NET0131  ;
  assign n7430 = ~n7428 & ~n7429 ;
  assign n7431 = RESET_pad & ~n7430 ;
  assign n7432 = ~\WX8615_reg/NET0131  & ~\_2289__reg/NET0131  ;
  assign n7433 = \WX8615_reg/NET0131  & \_2289__reg/NET0131  ;
  assign n7434 = ~n7432 & ~n7433 ;
  assign n7435 = RESET_pad & ~n7434 ;
  assign n7436 = ~\WX8613_reg/NET0131  & ~\_2290__reg/NET0131  ;
  assign n7437 = \WX8613_reg/NET0131  & \_2290__reg/NET0131  ;
  assign n7438 = ~n7436 & ~n7437 ;
  assign n7439 = RESET_pad & ~n7438 ;
  assign n7440 = ~\WX8611_reg/NET0131  & ~\_2291__reg/NET0131  ;
  assign n7441 = \WX8611_reg/NET0131  & \_2291__reg/NET0131  ;
  assign n7442 = ~n7440 & ~n7441 ;
  assign n7443 = RESET_pad & ~n7442 ;
  assign n7444 = ~\WX8609_reg/NET0131  & ~\_2292__reg/NET0131  ;
  assign n7445 = \WX8609_reg/NET0131  & \_2292__reg/NET0131  ;
  assign n7446 = ~n7444 & ~n7445 ;
  assign n7447 = RESET_pad & ~n7446 ;
  assign n7448 = ~\WX8597_reg/NET0131  & ~\_2298__reg/NET0131  ;
  assign n7449 = \WX8597_reg/NET0131  & \_2298__reg/NET0131  ;
  assign n7450 = ~n7448 & ~n7449 ;
  assign n7451 = RESET_pad & ~n7450 ;
  assign n7452 = ~\WX8595_reg/NET0131  & ~\_2299__reg/NET0131  ;
  assign n7453 = \WX8595_reg/NET0131  & \_2299__reg/NET0131  ;
  assign n7454 = ~n7452 & ~n7453 ;
  assign n7455 = RESET_pad & ~n7454 ;
  assign n7456 = ~\WX9950_reg/NET0131  & ~\_2332__reg/NET0131  ;
  assign n7457 = \WX9950_reg/NET0131  & \_2332__reg/NET0131  ;
  assign n7458 = ~n7456 & ~n7457 ;
  assign n7459 = RESET_pad & ~n7458 ;
  assign n7460 = ~\WX9948_reg/NET0131  & ~\_2301__reg/NET0131  ;
  assign n7461 = \WX9948_reg/NET0131  & \_2301__reg/NET0131  ;
  assign n7462 = ~n7460 & ~n7461 ;
  assign n7463 = RESET_pad & ~n7462 ;
  assign n7464 = ~\WX9946_reg/NET0131  & ~\_2302__reg/NET0131  ;
  assign n7465 = \WX9946_reg/NET0131  & \_2302__reg/NET0131  ;
  assign n7466 = ~n7464 & ~n7465 ;
  assign n7467 = RESET_pad & ~n7466 ;
  assign n7468 = ~\WX9940_reg/NET0131  & ~\_2305__reg/NET0131  ;
  assign n7469 = \WX9940_reg/NET0131  & \_2305__reg/NET0131  ;
  assign n7470 = ~n7468 & ~n7469 ;
  assign n7471 = RESET_pad & ~n7470 ;
  assign n7472 = ~\WX9938_reg/NET0131  & ~\_2306__reg/NET0131  ;
  assign n7473 = \WX9938_reg/NET0131  & \_2306__reg/NET0131  ;
  assign n7474 = ~n7472 & ~n7473 ;
  assign n7475 = RESET_pad & ~n7474 ;
  assign n7476 = ~\WX9932_reg/NET0131  & ~\_2309__reg/NET0131  ;
  assign n7477 = \WX9932_reg/NET0131  & \_2309__reg/NET0131  ;
  assign n7478 = ~n7476 & ~n7477 ;
  assign n7479 = RESET_pad & ~n7478 ;
  assign n7480 = ~\WX9926_reg/NET0131  & ~\_2312__reg/NET0131  ;
  assign n7481 = \WX9926_reg/NET0131  & \_2312__reg/NET0131  ;
  assign n7482 = ~n7480 & ~n7481 ;
  assign n7483 = RESET_pad & ~n7482 ;
  assign n7484 = ~\WX9922_reg/NET0131  & ~\_2314__reg/NET0131  ;
  assign n7485 = \WX9922_reg/NET0131  & \_2314__reg/NET0131  ;
  assign n7486 = ~n7484 & ~n7485 ;
  assign n7487 = RESET_pad & ~n7486 ;
  assign n7488 = ~\WX9920_reg/NET0131  & ~\_2315__reg/NET0131  ;
  assign n7489 = \WX9920_reg/NET0131  & \_2315__reg/NET0131  ;
  assign n7490 = ~n7488 & ~n7489 ;
  assign n7491 = RESET_pad & ~n7490 ;
  assign n7492 = ~\WX9916_reg/NET0131  & ~\_2317__reg/NET0131  ;
  assign n7493 = \WX9916_reg/NET0131  & \_2317__reg/NET0131  ;
  assign n7494 = ~n7492 & ~n7493 ;
  assign n7495 = RESET_pad & ~n7494 ;
  assign n7496 = ~\WX9914_reg/NET0131  & ~\_2318__reg/NET0131  ;
  assign n7497 = \WX9914_reg/NET0131  & \_2318__reg/NET0131  ;
  assign n7498 = ~n7496 & ~n7497 ;
  assign n7499 = RESET_pad & ~n7498 ;
  assign n7500 = ~\WX9912_reg/NET0131  & ~\_2319__reg/NET0131  ;
  assign n7501 = \WX9912_reg/NET0131  & \_2319__reg/NET0131  ;
  assign n7502 = ~n7500 & ~n7501 ;
  assign n7503 = RESET_pad & ~n7502 ;
  assign n7504 = ~\WX9910_reg/NET0131  & ~\_2320__reg/NET0131  ;
  assign n7505 = \WX9910_reg/NET0131  & \_2320__reg/NET0131  ;
  assign n7506 = ~n7504 & ~n7505 ;
  assign n7507 = RESET_pad & ~n7506 ;
  assign n7508 = ~\WX9908_reg/NET0131  & ~\_2321__reg/NET0131  ;
  assign n7509 = \WX9908_reg/NET0131  & \_2321__reg/NET0131  ;
  assign n7510 = ~n7508 & ~n7509 ;
  assign n7511 = RESET_pad & ~n7510 ;
  assign n7512 = ~\WX9906_reg/NET0131  & ~\_2322__reg/NET0131  ;
  assign n7513 = \WX9906_reg/NET0131  & \_2322__reg/NET0131  ;
  assign n7514 = ~n7512 & ~n7513 ;
  assign n7515 = RESET_pad & ~n7514 ;
  assign n7516 = ~\WX9904_reg/NET0131  & ~\_2323__reg/NET0131  ;
  assign n7517 = \WX9904_reg/NET0131  & \_2323__reg/NET0131  ;
  assign n7518 = ~n7516 & ~n7517 ;
  assign n7519 = RESET_pad & ~n7518 ;
  assign n7520 = ~\WX9902_reg/NET0131  & ~\_2324__reg/NET0131  ;
  assign n7521 = \WX9902_reg/NET0131  & \_2324__reg/NET0131  ;
  assign n7522 = ~n7520 & ~n7521 ;
  assign n7523 = RESET_pad & ~n7522 ;
  assign n7524 = ~\WX9900_reg/NET0131  & ~\_2325__reg/NET0131  ;
  assign n7525 = \WX9900_reg/NET0131  & \_2325__reg/NET0131  ;
  assign n7526 = ~n7524 & ~n7525 ;
  assign n7527 = RESET_pad & ~n7526 ;
  assign n7528 = ~\WX9898_reg/NET0131  & ~\_2326__reg/NET0131  ;
  assign n7529 = \WX9898_reg/NET0131  & \_2326__reg/NET0131  ;
  assign n7530 = ~n7528 & ~n7529 ;
  assign n7531 = RESET_pad & ~n7530 ;
  assign n7532 = ~\WX9896_reg/NET0131  & ~\_2327__reg/NET0131  ;
  assign n7533 = \WX9896_reg/NET0131  & \_2327__reg/NET0131  ;
  assign n7534 = ~n7532 & ~n7533 ;
  assign n7535 = RESET_pad & ~n7534 ;
  assign n7536 = ~\WX9894_reg/NET0131  & ~\_2328__reg/NET0131  ;
  assign n7537 = \WX9894_reg/NET0131  & \_2328__reg/NET0131  ;
  assign n7538 = ~n7536 & ~n7537 ;
  assign n7539 = RESET_pad & ~n7538 ;
  assign n7540 = ~\WX9892_reg/NET0131  & ~\_2329__reg/NET0131  ;
  assign n7541 = \WX9892_reg/NET0131  & \_2329__reg/NET0131  ;
  assign n7542 = ~n7540 & ~n7541 ;
  assign n7543 = RESET_pad & ~n7542 ;
  assign n7544 = ~\WX9888_reg/NET0131  & ~\_2331__reg/NET0131  ;
  assign n7545 = \WX9888_reg/NET0131  & \_2331__reg/NET0131  ;
  assign n7546 = ~n7544 & ~n7545 ;
  assign n7547 = RESET_pad & ~n7546 ;
  assign n7548 = ~\WX11243_reg/NET0131  & ~\_2364__reg/NET0131  ;
  assign n7549 = \WX11243_reg/NET0131  & \_2364__reg/NET0131  ;
  assign n7550 = ~n7548 & ~n7549 ;
  assign n7551 = RESET_pad & ~n7550 ;
  assign n7552 = ~\WX11241_reg/NET0131  & ~\_2333__reg/NET0131  ;
  assign n7553 = \WX11241_reg/NET0131  & \_2333__reg/NET0131  ;
  assign n7554 = ~n7552 & ~n7553 ;
  assign n7555 = RESET_pad & ~n7554 ;
  assign n7556 = ~\WX11239_reg/NET0131  & ~\_2334__reg/NET0131  ;
  assign n7557 = \WX11239_reg/NET0131  & \_2334__reg/NET0131  ;
  assign n7558 = ~n7556 & ~n7557 ;
  assign n7559 = RESET_pad & ~n7558 ;
  assign n7560 = ~\WX11237_reg/NET0131  & ~\_2335__reg/NET0131  ;
  assign n7561 = \WX11237_reg/NET0131  & \_2335__reg/NET0131  ;
  assign n7562 = ~n7560 & ~n7561 ;
  assign n7563 = RESET_pad & ~n7562 ;
  assign n7564 = ~\WX11233_reg/NET0131  & ~\_2337__reg/NET0131  ;
  assign n7565 = \WX11233_reg/NET0131  & \_2337__reg/NET0131  ;
  assign n7566 = ~n7564 & ~n7565 ;
  assign n7567 = RESET_pad & ~n7566 ;
  assign n7568 = ~\WX11231_reg/NET0131  & ~\_2338__reg/NET0131  ;
  assign n7569 = \WX11231_reg/NET0131  & \_2338__reg/NET0131  ;
  assign n7570 = ~n7568 & ~n7569 ;
  assign n7571 = RESET_pad & ~n7570 ;
  assign n7572 = ~\WX11229_reg/NET0131  & ~\_2339__reg/NET0131  ;
  assign n7573 = \WX11229_reg/NET0131  & \_2339__reg/NET0131  ;
  assign n7574 = ~n7572 & ~n7573 ;
  assign n7575 = RESET_pad & ~n7574 ;
  assign n7576 = ~\WX11227_reg/NET0131  & ~\_2340__reg/NET0131  ;
  assign n7577 = \WX11227_reg/NET0131  & \_2340__reg/NET0131  ;
  assign n7578 = ~n7576 & ~n7577 ;
  assign n7579 = RESET_pad & ~n7578 ;
  assign n7580 = ~\WX11225_reg/NET0131  & ~\_2341__reg/NET0131  ;
  assign n7581 = \WX11225_reg/NET0131  & \_2341__reg/NET0131  ;
  assign n7582 = ~n7580 & ~n7581 ;
  assign n7583 = RESET_pad & ~n7582 ;
  assign n7584 = ~\WX11223_reg/NET0131  & ~\_2342__reg/NET0131  ;
  assign n7585 = \WX11223_reg/NET0131  & \_2342__reg/NET0131  ;
  assign n7586 = ~n7584 & ~n7585 ;
  assign n7587 = RESET_pad & ~n7586 ;
  assign n7588 = ~\WX11219_reg/NET0131  & ~\_2344__reg/NET0131  ;
  assign n7589 = \WX11219_reg/NET0131  & \_2344__reg/NET0131  ;
  assign n7590 = ~n7588 & ~n7589 ;
  assign n7591 = RESET_pad & ~n7590 ;
  assign n7592 = ~\WX11217_reg/NET0131  & ~\_2345__reg/NET0131  ;
  assign n7593 = \WX11217_reg/NET0131  & \_2345__reg/NET0131  ;
  assign n7594 = ~n7592 & ~n7593 ;
  assign n7595 = RESET_pad & ~n7594 ;
  assign n7596 = ~\WX11213_reg/NET0131  & ~\_2347__reg/NET0131  ;
  assign n7597 = \WX11213_reg/NET0131  & \_2347__reg/NET0131  ;
  assign n7598 = ~n7596 & ~n7597 ;
  assign n7599 = RESET_pad & ~n7598 ;
  assign n7600 = ~\WX11209_reg/NET0131  & ~\_2349__reg/NET0131  ;
  assign n7601 = \WX11209_reg/NET0131  & \_2349__reg/NET0131  ;
  assign n7602 = ~n7600 & ~n7601 ;
  assign n7603 = RESET_pad & ~n7602 ;
  assign n7604 = ~\WX11207_reg/NET0131  & ~\_2350__reg/NET0131  ;
  assign n7605 = \WX11207_reg/NET0131  & \_2350__reg/NET0131  ;
  assign n7606 = ~n7604 & ~n7605 ;
  assign n7607 = RESET_pad & ~n7606 ;
  assign n7608 = ~\WX11205_reg/NET0131  & ~\_2351__reg/NET0131  ;
  assign n7609 = \WX11205_reg/NET0131  & \_2351__reg/NET0131  ;
  assign n7610 = ~n7608 & ~n7609 ;
  assign n7611 = RESET_pad & ~n7610 ;
  assign n7612 = ~\WX11203_reg/NET0131  & ~\_2352__reg/NET0131  ;
  assign n7613 = \WX11203_reg/NET0131  & \_2352__reg/NET0131  ;
  assign n7614 = ~n7612 & ~n7613 ;
  assign n7615 = RESET_pad & ~n7614 ;
  assign n7616 = ~\WX11201_reg/NET0131  & ~\_2353__reg/NET0131  ;
  assign n7617 = \WX11201_reg/NET0131  & \_2353__reg/NET0131  ;
  assign n7618 = ~n7616 & ~n7617 ;
  assign n7619 = RESET_pad & ~n7618 ;
  assign n7620 = ~\WX11199_reg/NET0131  & ~\_2354__reg/NET0131  ;
  assign n7621 = \WX11199_reg/NET0131  & \_2354__reg/NET0131  ;
  assign n7622 = ~n7620 & ~n7621 ;
  assign n7623 = RESET_pad & ~n7622 ;
  assign n7624 = ~\WX11197_reg/NET0131  & ~\_2355__reg/NET0131  ;
  assign n7625 = \WX11197_reg/NET0131  & \_2355__reg/NET0131  ;
  assign n7626 = ~n7624 & ~n7625 ;
  assign n7627 = RESET_pad & ~n7626 ;
  assign n7628 = ~\WX11195_reg/NET0131  & ~\_2356__reg/NET0131  ;
  assign n7629 = \WX11195_reg/NET0131  & \_2356__reg/NET0131  ;
  assign n7630 = ~n7628 & ~n7629 ;
  assign n7631 = RESET_pad & ~n7630 ;
  assign n7632 = ~\WX11193_reg/NET0131  & ~\_2357__reg/NET0131  ;
  assign n7633 = \WX11193_reg/NET0131  & \_2357__reg/NET0131  ;
  assign n7634 = ~n7632 & ~n7633 ;
  assign n7635 = RESET_pad & ~n7634 ;
  assign n7636 = ~\WX11191_reg/NET0131  & ~\_2358__reg/NET0131  ;
  assign n7637 = \WX11191_reg/NET0131  & \_2358__reg/NET0131  ;
  assign n7638 = ~n7636 & ~n7637 ;
  assign n7639 = RESET_pad & ~n7638 ;
  assign n7640 = ~\WX11189_reg/NET0131  & ~\_2359__reg/NET0131  ;
  assign n7641 = \WX11189_reg/NET0131  & \_2359__reg/NET0131  ;
  assign n7642 = ~n7640 & ~n7641 ;
  assign n7643 = RESET_pad & ~n7642 ;
  assign n7644 = ~\WX11187_reg/NET0131  & ~\_2360__reg/NET0131  ;
  assign n7645 = \WX11187_reg/NET0131  & \_2360__reg/NET0131  ;
  assign n7646 = ~n7644 & ~n7645 ;
  assign n7647 = RESET_pad & ~n7646 ;
  assign n7648 = ~\WX11183_reg/NET0131  & ~\_2362__reg/NET0131  ;
  assign n7649 = \WX11183_reg/NET0131  & \_2362__reg/NET0131  ;
  assign n7650 = ~n7648 & ~n7649 ;
  assign n7651 = RESET_pad & ~n7650 ;
  assign n7652 = ~\WX2150_reg/NET0131  & ~\_2129__reg/NET0131  ;
  assign n7653 = \WX2150_reg/NET0131  & \_2129__reg/NET0131  ;
  assign n7654 = ~n7652 & ~n7653 ;
  assign n7655 = RESET_pad & ~n7654 ;
  assign n7656 = ~\WX7304_reg/NET0131  & ~\_2266__reg/NET0131  ;
  assign n7657 = \WX7304_reg/NET0131  & \_2266__reg/NET0131  ;
  assign n7658 = ~n7656 & ~n7657 ;
  assign n7659 = RESET_pad & ~n7658 ;
  assign n7660 = ~\WX2136_reg/NET0131  & ~\_2136__reg/NET0131  ;
  assign n7661 = \WX2136_reg/NET0131  & \_2136__reg/NET0131  ;
  assign n7662 = ~n7660 & ~n7661 ;
  assign n7663 = RESET_pad & ~n7662 ;
  assign n7664 = ~\WX3467_reg/NET0131  & ~\_2149__reg/NET0131  ;
  assign n7665 = \WX3467_reg/NET0131  & \_2149__reg/NET0131  ;
  assign n7666 = ~n7664 & ~n7665 ;
  assign n7667 = RESET_pad & ~n7666 ;
  assign n7668 = ~\WX8633_reg/NET0131  & ~\_2280__reg/NET0131  ;
  assign n7669 = \WX8633_reg/NET0131  & \_2280__reg/NET0131  ;
  assign n7670 = ~n7668 & ~n7669 ;
  assign n7671 = RESET_pad & ~n7670 ;
  assign n7672 = ~\WX853_reg/NET0131  & ~\_2099__reg/NET0131  ;
  assign n7673 = \WX853_reg/NET0131  & \_2099__reg/NET0131  ;
  assign n7674 = ~n7672 & ~n7673 ;
  assign n7675 = RESET_pad & ~n7674 ;
  assign n7676 = ~\WX859_reg/NET0131  & ~\_2096__reg/NET0131  ;
  assign n7677 = \WX859_reg/NET0131  & \_2096__reg/NET0131  ;
  assign n7678 = ~n7676 & ~n7677 ;
  assign n7679 = RESET_pad & ~n7678 ;
  assign n7680 = ~\WX7310_reg/NET0131  & ~\_2263__reg/NET0131  ;
  assign n7681 = \WX7310_reg/NET0131  & \_2263__reg/NET0131  ;
  assign n7682 = ~n7680 & ~n7681 ;
  assign n7683 = RESET_pad & ~n7682 ;
  assign n7684 = ~\WX9936_reg/NET0131  & ~\_2307__reg/NET0131  ;
  assign n7685 = \WX9936_reg/NET0131  & \_2307__reg/NET0131  ;
  assign n7686 = ~n7684 & ~n7685 ;
  assign n7687 = RESET_pad & ~n7686 ;
  assign n7688 = ~\WX849_reg/NET0131  & ~\_2101__reg/NET0131  ;
  assign n7689 = \WX849_reg/NET0131  & \_2101__reg/NET0131  ;
  assign n7690 = ~n7688 & ~n7689 ;
  assign n7691 = RESET_pad & ~n7690 ;
  assign n7692 = ~\WX2140_reg/NET0131  & ~\_2134__reg/NET0131  ;
  assign n7693 = \WX2140_reg/NET0131  & \_2134__reg/NET0131  ;
  assign n7694 = ~n7692 & ~n7693 ;
  assign n7695 = RESET_pad & ~n7694 ;
  assign n7696 = ~\WX2178_reg/NET0131  & ~\_2115__reg/NET0131  ;
  assign n7697 = \WX2178_reg/NET0131  & \_2115__reg/NET0131  ;
  assign n7698 = ~n7696 & ~n7697 ;
  assign n7699 = RESET_pad & ~n7698 ;
  assign n7700 = ~\WX8623_reg/NET0131  & ~\_2285__reg/NET0131  ;
  assign n7701 = \WX8623_reg/NET0131  & \_2285__reg/NET0131  ;
  assign n7702 = ~n7700 & ~n7701 ;
  assign n7703 = RESET_pad & ~n7702 ;
  assign n7704 = ~\WX2176_reg/NET0131  & ~\_2116__reg/NET0131  ;
  assign n7705 = \WX2176_reg/NET0131  & \_2116__reg/NET0131  ;
  assign n7706 = ~n7704 & ~n7705 ;
  assign n7707 = RESET_pad & ~n7706 ;
  assign n7708 = ~\WX7346_reg/NET0131  & ~\_2245__reg/NET0131  ;
  assign n7709 = \WX7346_reg/NET0131  & \_2245__reg/NET0131  ;
  assign n7710 = ~n7708 & ~n7709 ;
  assign n7711 = RESET_pad & ~n7710 ;
  assign n7712 = ~\WX6041_reg/NET0131  & ~\_2219__reg/NET0131  ;
  assign n7713 = \WX6041_reg/NET0131  & \_2219__reg/NET0131  ;
  assign n7714 = ~n7712 & ~n7713 ;
  assign n7715 = RESET_pad & ~n7714 ;
  assign n7716 = ~\WX7350_reg/NET0131  & ~\_2243__reg/NET0131  ;
  assign n7717 = \WX7350_reg/NET0131  & \_2243__reg/NET0131  ;
  assign n7718 = ~n7716 & ~n7717 ;
  assign n7719 = RESET_pad & ~n7718 ;
  assign n7720 = ~\WX4762_reg/NET0131  & ~\_2180__reg/NET0131  ;
  assign n7721 = \WX4762_reg/NET0131  & \_2180__reg/NET0131  ;
  assign n7722 = ~n7720 & ~n7721 ;
  assign n7723 = RESET_pad & ~n7722 ;
  assign n7724 = ~\WX871_reg/NET0131  & ~\_2090__reg/NET0131  ;
  assign n7725 = \WX871_reg/NET0131  & \_2090__reg/NET0131  ;
  assign n7726 = ~n7724 & ~n7725 ;
  assign n7727 = RESET_pad & ~n7726 ;
  assign n7728 = ~\WX885_reg/NET0131  & ~\_2083__reg/NET0131  ;
  assign n7729 = \WX885_reg/NET0131  & \_2083__reg/NET0131  ;
  assign n7730 = ~n7728 & ~n7729 ;
  assign n7731 = RESET_pad & ~n7730 ;
  assign n7732 = ~\WX11185_reg/NET0131  & ~\_2361__reg/NET0131  ;
  assign n7733 = \WX11185_reg/NET0131  & \_2361__reg/NET0131  ;
  assign n7734 = ~n7732 & ~n7733 ;
  assign n7735 = RESET_pad & ~n7734 ;
  assign n7736 = ~\WX9890_reg/NET0131  & ~\_2330__reg/NET0131  ;
  assign n7737 = \WX9890_reg/NET0131  & \_2330__reg/NET0131  ;
  assign n7738 = ~n7736 & ~n7737 ;
  assign n7739 = RESET_pad & ~n7738 ;
  assign n7740 = ~\WX9944_reg/NET0131  & ~\_2303__reg/NET0131  ;
  assign n7741 = \WX9944_reg/NET0131  & \_2303__reg/NET0131  ;
  assign n7742 = ~n7740 & ~n7741 ;
  assign n7743 = RESET_pad & ~n7742 ;
  assign n7744 = ~\WX7344_reg/NET0131  & ~\_2246__reg/NET0131  ;
  assign n7745 = \WX7344_reg/NET0131  & \_2246__reg/NET0131  ;
  assign n7746 = ~n7744 & ~n7745 ;
  assign n7747 = RESET_pad & ~n7746 ;
  assign n7748 = ~\WX7324_reg/NET0131  & ~\_2256__reg/NET0131  ;
  assign n7749 = \WX7324_reg/NET0131  & \_2256__reg/NET0131  ;
  assign n7750 = ~n7748 & ~n7749 ;
  assign n7751 = RESET_pad & ~n7750 ;
  assign n7752 = ~\WX6013_reg/NET0131  & ~\_2233__reg/NET0131  ;
  assign n7753 = \WX6013_reg/NET0131  & \_2233__reg/NET0131  ;
  assign n7754 = ~n7752 & ~n7753 ;
  assign n7755 = RESET_pad & ~n7754 ;
  assign n7756 = ~\WX2152_reg/NET0131  & ~\_2128__reg/NET0131  ;
  assign n7757 = \WX2152_reg/NET0131  & \_2128__reg/NET0131  ;
  assign n7758 = ~n7756 & ~n7757 ;
  assign n7759 = RESET_pad & ~n7758 ;
  assign n7760 = ~\WX847_reg/NET0131  & ~\_2102__reg/NET0131  ;
  assign n7761 = \WX847_reg/NET0131  & \_2102__reg/NET0131  ;
  assign n7762 = ~n7760 & ~n7761 ;
  assign n7763 = RESET_pad & ~n7762 ;
  assign n7764 = ~\WX3447_reg/NET0131  & ~\_2159__reg/NET0131  ;
  assign n7765 = \WX3447_reg/NET0131  & \_2159__reg/NET0131  ;
  assign n7766 = ~n7764 & ~n7765 ;
  assign n7767 = RESET_pad & ~n7766 ;
  assign n7768 = ~\WX9924_reg/NET0131  & ~\_2313__reg/NET0131  ;
  assign n7769 = \WX9924_reg/NET0131  & \_2313__reg/NET0131  ;
  assign n7770 = ~n7768 & ~n7769 ;
  assign n7771 = RESET_pad & ~n7770 ;
  assign n7772 = ~\WX861_reg/NET0131  & ~\_2095__reg/NET0131  ;
  assign n7773 = \WX861_reg/NET0131  & \_2095__reg/NET0131  ;
  assign n7774 = ~n7772 & ~n7773 ;
  assign n7775 = RESET_pad & ~n7774 ;
  assign n7776 = ~\WX8639_reg/NET0131  & ~\_2277__reg/NET0131  ;
  assign n7777 = \WX8639_reg/NET0131  & \_2277__reg/NET0131  ;
  assign n7778 = ~n7776 & ~n7777 ;
  assign n7779 = RESET_pad & ~n7778 ;
  assign n7780 = ~\WX7308_reg/NET0131  & ~\_2264__reg/NET0131  ;
  assign n7781 = \WX7308_reg/NET0131  & \_2264__reg/NET0131  ;
  assign n7782 = ~n7780 & ~n7781 ;
  assign n7783 = RESET_pad & ~n7782 ;
  assign n7784 = ~\WX879_reg/NET0131  & ~\_2086__reg/NET0131  ;
  assign n7785 = \WX879_reg/NET0131  & \_2086__reg/NET0131  ;
  assign n7786 = ~n7784 & ~n7785 ;
  assign n7787 = RESET_pad & ~n7786 ;
  assign n7788 = ~\WX7334_reg/NET0131  & ~\_2251__reg/NET0131  ;
  assign n7789 = \WX7334_reg/NET0131  & \_2251__reg/NET0131  ;
  assign n7790 = ~n7788 & ~n7789 ;
  assign n7791 = RESET_pad & ~n7790 ;
  assign n7792 = ~\WX8643_reg/NET0131  & ~\_2275__reg/NET0131  ;
  assign n7793 = \WX8643_reg/NET0131  & \_2275__reg/NET0131  ;
  assign n7794 = ~n7792 & ~n7793 ;
  assign n7795 = RESET_pad & ~n7794 ;
  assign n7796 = ~\WX4726_reg/NET0131  & ~\_2198__reg/NET0131  ;
  assign n7797 = \WX4726_reg/NET0131  & \_2198__reg/NET0131  ;
  assign n7798 = ~n7796 & ~n7797 ;
  assign n7799 = RESET_pad & ~n7798 ;
  assign n7800 = RESET_pad & \WX11053_reg/NET0131  ;
  assign n7801 = RESET_pad & \WX709_reg/NET0131  ;
  assign n7802 = RESET_pad & \WX10891_reg/NET0131  ;
  assign n7803 = RESET_pad & \WX2002_reg/NET0131  ;
  assign n7804 = RESET_pad & ~\WX10829_reg/NET0131  ;
  assign n7805 = RESET_pad & \WX11059_reg/NET0131  ;
  assign n7806 = RESET_pad & \WX3271_reg/NET0131  ;
  assign n7807 = RESET_pad & \WX11033_reg/NET0131  ;
  assign n7808 = RESET_pad & \WX7252_reg/NET0131  ;
  assign n7809 = RESET_pad & \WX3257_reg/NET0131  ;
  assign n7810 = RESET_pad & \WX3403_reg/NET0131  ;
  assign n7811 = RESET_pad & \WX11115_reg/NET0131  ;
  assign n7812 = RESET_pad & \WX11049_reg/NET0131  ;
  assign n7813 = RESET_pad & \WX9714_reg/NET0131  ;
  assign n7814 = RESET_pad & \WX2004_reg/NET0131  ;
  assign n7815 = RESET_pad & \WX11037_reg/NET0131  ;
  assign n7816 = RESET_pad & \WX9852_reg/NET0131  ;
  assign n7817 = RESET_pad & \WX9702_reg/NET0131  ;
  assign n7818 = RESET_pad & \WX9876_reg/NET0131  ;
  assign n7819 = RESET_pad & \WX11121_reg/NET0131  ;
  assign n7820 = RESET_pad & \WX7114_reg/NET0131  ;
  assign n7821 = RESET_pad & \WX1986_reg/NET0131  ;
  assign n7822 = RESET_pad & \WX9802_reg/NET0131  ;
  assign n7823 = RESET_pad & \WX9824_reg/NET0131  ;
  assign n7824 = RESET_pad & \WX7220_reg/NET0131  ;
  assign n7825 = RESET_pad & \WX9806_reg/NET0131  ;
  assign n7826 = RESET_pad & \WX11073_reg/NET0131  ;
  assign n7827 = RESET_pad & \WX9878_reg/NET0131  ;
  assign n7828 = RESET_pad & \WX11111_reg/NET0131  ;
  assign n7829 = RESET_pad & \WX11169_reg/NET0131  ;
  assign n7830 = RESET_pad & \WX1998_reg/NET0131  ;
  assign n7831 = RESET_pad & \WX9850_reg/NET0131  ;
  assign n7832 = RESET_pad & \WX11079_reg/NET0131  ;
  assign n7833 = RESET_pad & \WX7110_reg/NET0131  ;
  assign n7834 = RESET_pad & \WX7240_reg/NET0131  ;
  assign n7835 = RESET_pad & \WX1954_reg/NET0131  ;
  assign n7836 = RESET_pad & \WX11081_reg/NET0131  ;
  assign n7837 = RESET_pad & \WX11083_reg/NET0131  ;
  assign n7838 = RESET_pad & \WX3339_reg/NET0131  ;
  assign n7839 = RESET_pad & \WX8491_reg/NET0131  ;
  assign n7840 = RESET_pad & \WX11175_reg/NET0131  ;
  assign n7841 = RESET_pad & \WX11089_reg/NET0131  ;
  assign n7842 = RESET_pad & \WX9770_reg/NET0131  ;
  assign n7843 = RESET_pad & \WX2068_reg/NET0131  ;
  assign n7844 = RESET_pad & \WX823_reg/NET0131  ;
  assign n7845 = RESET_pad & \WX5941_reg/NET0131  ;
  assign n7846 = RESET_pad & \WX11093_reg/NET0131  ;
  assign n7847 = RESET_pad & \WX5919_reg/NET0131  ;
  assign n7848 = RESET_pad & \WX7160_reg/NET0131  ;
  assign n7849 = RESET_pad & \WX791_reg/NET0131  ;
  assign n7850 = RESET_pad & \WX11095_reg/NET0131  ;
  assign n7851 = RESET_pad & \WX3349_reg/NET0131  ;
  assign n7852 = RESET_pad & \WX9708_reg/NET0131  ;
  assign n7853 = RESET_pad & \WX769_reg/NET0131  ;
  assign n7854 = RESET_pad & \WX11153_reg/NET0131  ;
  assign n7855 = RESET_pad & \WX7182_reg/NET0131  ;
  assign n7856 = RESET_pad & \WX7238_reg/NET0131  ;
  assign n7857 = RESET_pad & \WX11103_reg/NET0131  ;
  assign n7858 = RESET_pad & \WX5925_reg/NET0131  ;
  assign n7859 = RESET_pad & \WX7196_reg/NET0131  ;
  assign n7860 = RESET_pad & \WX7204_reg/NET0131  ;
  assign n7861 = RESET_pad & \WX3279_reg/NET0131  ;
  assign n7862 = RESET_pad & \WX5953_reg/NET0131  ;
  assign n7863 = RESET_pad & \WX3285_reg/NET0131  ;
  assign n7864 = RESET_pad & \WX4594_reg/NET0131  ;
  assign n7865 = RESET_pad & \WX777_reg/NET0131  ;
  assign n7866 = RESET_pad & \WX7164_reg/NET0131  ;
  assign n7867 = RESET_pad & \WX11167_reg/NET0131  ;
  assign n7868 = RESET_pad & \WX719_reg/NET0131  ;
  assign n7869 = RESET_pad & \WX707_reg/NET0131  ;
  assign n7870 = RESET_pad & \WX7294_reg/NET0131  ;
  assign n7871 = RESET_pad & \WX11113_reg/NET0131  ;
  assign n7872 = RESET_pad & \WX1988_reg/NET0131  ;
  assign n7873 = RESET_pad & \WX7234_reg/NET0131  ;
  assign n7874 = RESET_pad & \WX9712_reg/NET0131  ;
  assign n7875 = RESET_pad & \WX5929_reg/NET0131  ;
  assign n7876 = RESET_pad & \WX7244_reg/NET0131  ;
  assign n7877 = RESET_pad & \WX7248_reg/NET0131  ;
  assign n7878 = RESET_pad & \WX9882_reg/NET0131  ;
  assign n7879 = RESET_pad & \WX4550_reg/NET0131  ;
  assign n7880 = RESET_pad & \WX665_reg/NET0131  ;
  assign n7881 = RESET_pad & \WX7232_reg/NET0131  ;
  assign n7882 = RESET_pad & \WX705_reg/NET0131  ;
  assign n7883 = RESET_pad & \WX2064_reg/NET0131  ;
  assign n7884 = RESET_pad & \WX5927_reg/NET0131  ;
  assign n7885 = RESET_pad & \WX9822_reg/NET0131  ;
  assign n7886 = RESET_pad & \WX7276_reg/NET0131  ;
  assign n7887 = RESET_pad & \WX3277_reg/NET0131  ;
  assign n7888 = RESET_pad & \WX7284_reg/NET0131  ;
  assign n7889 = RESET_pad & \WX11177_reg/NET0131  ;
  assign n7890 = RESET_pad & \WX645_reg/NET0131  ;
  assign n7891 = RESET_pad & \WX11133_reg/NET0131  ;
  assign n7892 = RESET_pad & \WX1992_reg/NET0131  ;
  assign n7893 = RESET_pad & \WX11135_reg/NET0131  ;
  assign n7894 = RESET_pad & \WX11137_reg/NET0131  ;
  assign n7895 = RESET_pad & \WX2072_reg/NET0131  ;
  assign n7896 = RESET_pad & \WX11161_reg/NET0131  ;
  assign n7897 = RESET_pad & \WX5933_reg/NET0131  ;
  assign n7898 = RESET_pad & \WX3379_reg/NET0131  ;
  assign n7899 = RESET_pad & \WX4556_reg/NET0131  ;
  assign n7900 = RESET_pad & \WX11143_reg/NET0131  ;
  assign n7901 = RESET_pad & \WX9750_reg/NET0131  ;
  assign n7902 = RESET_pad & \WX9786_reg/NET0131  ;
  assign n7903 = RESET_pad & \WX7230_reg/NET0131  ;
  assign n7904 = RESET_pad & \WX3237_reg/NET0131  ;
  assign n7905 = RESET_pad & \WX11041_reg/NET0131  ;
  assign n7906 = RESET_pad & \WX5939_reg/NET0131  ;
  assign n7907 = RESET_pad & \WX9716_reg/NET0131  ;
  assign n7908 = RESET_pad & \WX5871_reg/NET0131  ;
  assign n7909 = RESET_pad & \WX757_reg/NET0131  ;
  assign n7910 = RESET_pad & \WX11045_reg/NET0131  ;
  assign n7911 = RESET_pad & \WX9744_reg/NET0131  ;
  assign n7912 = RESET_pad & \WX9762_reg/NET0131  ;
  assign n7913 = RESET_pad & \WX4558_reg/NET0131  ;
  assign n7914 = RESET_pad & \WX3273_reg/NET0131  ;
  assign n7915 = RESET_pad & \WX5945_reg/NET0131  ;
  assign n7916 = RESET_pad & \WX9860_reg/NET0131  ;
  assign n7917 = RESET_pad & \WX7228_reg/NET0131  ;
  assign n7918 = RESET_pad & \WX7226_reg/NET0131  ;
  assign n7919 = RESET_pad & \WX4542_reg/NET0131  ;
  assign n7920 = RESET_pad & \WX9808_reg/NET0131  ;
  assign n7921 = RESET_pad & \WX11109_reg/NET0131  ;
  assign n7922 = RESET_pad & \WX8423_reg/NET0131  ;
  assign n7923 = RESET_pad & \WX3327_reg/NET0131  ;
  assign n7924 = RESET_pad & \WX807_reg/NET0131  ;
  assign n7925 = RESET_pad & \WX8533_reg/NET0131  ;
  assign n7926 = RESET_pad & \WX7222_reg/NET0131  ;
  assign n7927 = RESET_pad & \WX9856_reg/NET0131  ;
  assign n7928 = RESET_pad & \WX1984_reg/NET0131  ;
  assign n7929 = RESET_pad & \WX7118_reg/NET0131  ;
  assign n7930 = RESET_pad & \WX7218_reg/NET0131  ;
  assign n7931 = RESET_pad & \WX7224_reg/NET0131  ;
  assign n7932 = RESET_pad & \WX4544_reg/NET0131  ;
  assign n7933 = RESET_pad & \WX4560_reg/NET0131  ;
  assign n7934 = RESET_pad & \WX667_reg/NET0131  ;
  assign n7935 = RESET_pad & \WX7214_reg/NET0131  ;
  assign n7936 = RESET_pad & \WX3319_reg/NET0131  ;
  assign n7937 = RESET_pad & \WX663_reg/NET0131  ;
  assign n7938 = RESET_pad & \WX4598_reg/NET0131  ;
  assign n7939 = RESET_pad & \WX9820_reg/NET0131  ;
  assign n7940 = RESET_pad & \WX5979_reg/NET0131  ;
  assign n7941 = RESET_pad & \WX11107_reg/NET0131  ;
  assign n7942 = RESET_pad & \WX9698_reg/NET0131  ;
  assign n7943 = RESET_pad & \WX7198_reg/NET0131  ;
  assign n7944 = RESET_pad & \WX3365_reg/NET0131  ;
  assign n7945 = RESET_pad & \WX11131_reg/NET0131  ;
  assign n7946 = RESET_pad & \WX3361_reg/NET0131  ;
  assign n7947 = RESET_pad & \WX11163_reg/NET0131  ;
  assign n7948 = RESET_pad & \WX8517_reg/NET0131  ;
  assign n7949 = RESET_pad & \WX9772_reg/NET0131  ;
  assign n7950 = RESET_pad & \WX11105_reg/NET0131  ;
  assign n7951 = RESET_pad & \WX11123_reg/NET0131  ;
  assign n7952 = RESET_pad & \WX3351_reg/NET0131  ;
  assign n7953 = RESET_pad & \WX4562_reg/NET0131  ;
  assign n7954 = RESET_pad & \WX4540_reg/NET0131  ;
  assign n7955 = RESET_pad & \WX5879_reg/NET0131  ;
  assign n7956 = RESET_pad & \WX5875_reg/NET0131  ;
  assign n7957 = RESET_pad & \WX5991_reg/NET0131  ;
  assign n7958 = RESET_pad & \WX2056_reg/NET0131  ;
  assign n7959 = RESET_pad & \WX3263_reg/NET0131  ;
  assign n7960 = RESET_pad & \WX7166_reg/NET0131  ;
  assign n7961 = RESET_pad & \WX7190_reg/NET0131  ;
  assign n7962 = RESET_pad & \WX1972_reg/NET0131  ;
  assign n7963 = RESET_pad & \WX661_reg/NET0131  ;
  assign n7964 = RESET_pad & \WX9774_reg/NET0131  ;
  assign n7965 = RESET_pad & \WX1994_reg/NET0131  ;
  assign n7966 = RESET_pad & \WX7256_reg/NET0131  ;
  assign n7967 = RESET_pad & \WX5985_reg/NET0131  ;
  assign n7968 = RESET_pad & \WX7192_reg/NET0131  ;
  assign n7969 = RESET_pad & \WX7194_reg/NET0131  ;
  assign n7970 = RESET_pad & \WX8445_reg/NET0131  ;
  assign n7971 = RESET_pad & \WX5999_reg/NET0131  ;
  assign n7972 = RESET_pad & \WX1966_reg/NET0131  ;
  assign n7973 = RESET_pad & \WX9726_reg/NET0131  ;
  assign n7974 = RESET_pad & \WX9704_reg/NET0131  ;
  assign n7975 = RESET_pad & \WX7186_reg/NET0131  ;
  assign n7976 = RESET_pad & \WX8441_reg/NET0131  ;
  assign n7977 = RESET_pad & \WX5923_reg/NET0131  ;
  assign n7978 = RESET_pad & \WX2128_reg/NET0131  ;
  assign n7979 = RESET_pad & \WX2126_reg/NET0131  ;
  assign n7980 = RESET_pad & \WX7180_reg/NET0131  ;
  assign n7981 = RESET_pad & \WX721_reg/NET0131  ;
  assign n7982 = RESET_pad & \WX7278_reg/NET0131  ;
  assign n7983 = RESET_pad & \WX835_reg/NET0131  ;
  assign n7984 = RESET_pad & \WX5997_reg/NET0131  ;
  assign n7985 = RESET_pad & \WX3363_reg/NET0131  ;
  assign n7986 = RESET_pad & \WX5921_reg/NET0131  ;
  assign n7987 = RESET_pad & \WX659_reg/NET0131  ;
  assign n7988 = RESET_pad & \WX3259_reg/NET0131  ;
  assign n7989 = RESET_pad & \WX9780_reg/NET0131  ;
  assign n7990 = RESET_pad & \WX1956_reg/NET0131  ;
  assign n7991 = RESET_pad & \WX11099_reg/NET0131  ;
  assign n7992 = RESET_pad & \WX2088_reg/NET0131  ;
  assign n7993 = RESET_pad & \WX9800_reg/NET0131  ;
  assign n7994 = RESET_pad & \WX767_reg/NET0131  ;
  assign n7995 = RESET_pad & \WX7280_reg/NET0131  ;
  assign n7996 = RESET_pad & \WX8519_reg/NET0131  ;
  assign n7997 = RESET_pad & \WX771_reg/NET0131  ;
  assign n7998 = RESET_pad & \WX781_reg/NET0131  ;
  assign n7999 = RESET_pad & \WX1958_reg/NET0131  ;
  assign n8000 = RESET_pad & \WX3289_reg/NET0131  ;
  assign n8001 = RESET_pad & \WX4638_reg/NET0131  ;
  assign n8002 = RESET_pad & \WX687_reg/NET0131  ;
  assign n8003 = RESET_pad & \WX2112_reg/NET0131  ;
  assign n8004 = RESET_pad & \WX9730_reg/NET0131  ;
  assign n8005 = RESET_pad & \WX9754_reg/NET0131  ;
  assign n8006 = RESET_pad & \WX787_reg/NET0131  ;
  assign n8007 = RESET_pad & \WX731_reg/NET0131  ;
  assign n8008 = RESET_pad & \WX3415_reg/NET0131  ;
  assign n8009 = RESET_pad & \WX3255_reg/NET0131  ;
  assign n8010 = RESET_pad & \WX2122_reg/NET0131  ;
  assign n8011 = RESET_pad & \WX8529_reg/NET0131  ;
  assign n8012 = RESET_pad & \WX9832_reg/NET0131  ;
  assign n8013 = RESET_pad & \WX8449_reg/NET0131  ;
  assign n8014 = RESET_pad & \WX727_reg/NET0131  ;
  assign n8015 = RESET_pad & \WX7158_reg/NET0131  ;
  assign n8016 = RESET_pad & \WX11011_reg/NET0131  ;
  assign n8017 = RESET_pad & \WX7152_reg/NET0131  ;
  assign n8018 = RESET_pad & \WX4676_reg/NET0131  ;
  assign n8019 = RESET_pad & \WX7156_reg/NET0131  ;
  assign n8020 = RESET_pad & \WX7154_reg/NET0131  ;
  assign n8021 = RESET_pad & \WX657_reg/NET0131  ;
  assign n8022 = RESET_pad & \WX9816_reg/NET0131  ;
  assign n8023 = RESET_pad & \WX831_reg/NET0131  ;
  assign n8024 = RESET_pad & \WX7134_reg/NET0131  ;
  assign n8025 = RESET_pad & \WX7246_reg/NET0131  ;
  assign n8026 = RESET_pad & \WX7144_reg/NET0131  ;
  assign n8027 = RESET_pad & \WX9736_reg/NET0131  ;
  assign n8028 = RESET_pad & \WX1946_reg/NET0131  ;
  assign n8029 = RESET_pad & \WX7150_reg/NET0131  ;
  assign n8030 = RESET_pad & \WX2000_reg/NET0131  ;
  assign n8031 = RESET_pad & \WX761_reg/NET0131  ;
  assign n8032 = RESET_pad & \WX9842_reg/NET0131  ;
  assign n8033 = RESET_pad & \WX819_reg/NET0131  ;
  assign n8034 = RESET_pad & \WX7148_reg/NET0131  ;
  assign n8035 = RESET_pad & \WX3321_reg/NET0131  ;
  assign n8036 = RESET_pad & \WX4634_reg/NET0131  ;
  assign n8037 = RESET_pad & \WX11087_reg/NET0131  ;
  assign n8038 = RESET_pad & \WX7124_reg/NET0131  ;
  assign n8039 = RESET_pad & \WX3301_reg/NET0131  ;
  assign n8040 = RESET_pad & \WX3409_reg/NET0131  ;
  assign n8041 = RESET_pad & \WX9778_reg/NET0131  ;
  assign n8042 = RESET_pad & \WX7272_reg/NET0131  ;
  assign n8043 = RESET_pad & \WX7138_reg/NET0131  ;
  assign n8044 = RESET_pad & \WX2118_reg/NET0131  ;
  assign n8045 = RESET_pad & \WX4626_reg/NET0131  ;
  assign n8046 = RESET_pad & \WX5949_reg/NET0131  ;
  assign n8047 = RESET_pad & \WX693_reg/NET0131  ;
  assign n8048 = RESET_pad & \WX3265_reg/NET0131  ;
  assign n8049 = RESET_pad & \WX11141_reg/NET0131  ;
  assign n8050 = RESET_pad & \WX5947_reg/NET0131  ;
  assign n8051 = RESET_pad & \WX2114_reg/NET0131  ;
  assign n8052 = RESET_pad & \WX4584_reg/NET0131  ;
  assign n8053 = RESET_pad & \WX735_reg/NET0131  ;
  assign n8054 = RESET_pad & \WX3267_reg/NET0131  ;
  assign n8055 = RESET_pad & \WX7120_reg/NET0131  ;
  assign n8056 = RESET_pad & \WX7132_reg/NET0131  ;
  assign n8057 = RESET_pad & \WX3357_reg/NET0131  ;
  assign n8058 = RESET_pad & \WX3281_reg/NET0131  ;
  assign n8059 = RESET_pad & \WX3247_reg/NET0131  ;
  assign n8060 = RESET_pad & \WX9798_reg/NET0131  ;
  assign n8061 = RESET_pad & \WX11119_reg/NET0131  ;
  assign n8062 = RESET_pad & \WX7126_reg/NET0131  ;
  assign n8063 = RESET_pad & \WX5937_reg/NET0131  ;
  assign n8064 = RESET_pad & \WX7128_reg/NET0131  ;
  assign n8065 = RESET_pad & \WX3347_reg/NET0131  ;
  assign n8066 = RESET_pad & \WX2060_reg/NET0131  ;
  assign n8067 = RESET_pad & \WX7130_reg/NET0131  ;
  assign n8068 = RESET_pad & \WX9742_reg/NET0131  ;
  assign n8069 = RESET_pad & \WX11085_reg/NET0131  ;
  assign n8070 = RESET_pad & \WX11043_reg/NET0131  ;
  assign n8071 = RESET_pad & \WX3283_reg/NET0131  ;
  assign n8072 = RESET_pad & \WX755_reg/NET0131  ;
  assign n8073 = RESET_pad & \WX8447_reg/NET0131  ;
  assign n8074 = RESET_pad & \WX669_reg/NET0131  ;
  assign n8075 = RESET_pad & \WX4564_reg/NET0131  ;
  assign n8076 = RESET_pad & \WX685_reg/NET0131  ;
  assign n8077 = RESET_pad & \WX11067_reg/NET0131  ;
  assign n8078 = RESET_pad & \WX8453_reg/NET0131  ;
  assign n8079 = RESET_pad & \WX4538_reg/NET0131  ;
  assign n8080 = RESET_pad & \WX5959_reg/NET0131  ;
  assign n8081 = RESET_pad & \WX3355_reg/NET0131  ;
  assign n8082 = RESET_pad & \WX4588_reg/NET0131  ;
  assign n8083 = RESET_pad & \WX9724_reg/NET0131  ;
  assign n8084 = RESET_pad & \WX5965_reg/NET0131  ;
  assign n8085 = RESET_pad & \WX11147_reg/NET0131  ;
  assign n8086 = RESET_pad & \WX7122_reg/NET0131  ;
  assign n8087 = RESET_pad & \WX695_reg/NET0131  ;
  assign n8088 = RESET_pad & \WX4636_reg/NET0131  ;
  assign n8089 = RESET_pad & \WX4628_reg/NET0131  ;
  assign n8090 = RESET_pad & \WX8551_reg/NET0131  ;
  assign n8091 = RESET_pad & \WX9872_reg/NET0131  ;
  assign n8092 = RESET_pad & \WX5861_reg/NET0131  ;
  assign n8093 = RESET_pad & \WX8407_reg/NET0131  ;
  assign n8094 = RESET_pad & \WX8547_reg/NET0131  ;
  assign n8095 = RESET_pad & \WX9862_reg/NET0131  ;
  assign n8096 = RESET_pad & \WX4570_reg/NET0131  ;
  assign n8097 = RESET_pad & \WX11027_reg/NET0131  ;
  assign n8098 = RESET_pad & \WX11139_reg/NET0131  ;
  assign n8099 = RESET_pad & \WX4652_reg/NET0131  ;
  assign n8100 = RESET_pad & \WX729_reg/NET0131  ;
  assign n8101 = RESET_pad & \WX5957_reg/NET0131  ;
  assign n8102 = RESET_pad & \WX3287_reg/NET0131  ;
  assign n8103 = RESET_pad & \WX801_reg/NET0131  ;
  assign n8104 = RESET_pad & \WX805_reg/NET0131  ;
  assign n8105 = RESET_pad & \WX11149_reg/NET0131  ;
  assign n8106 = RESET_pad & \WX691_reg/NET0131  ;
  assign n8107 = RESET_pad & \WX8557_reg/NET0131  ;
  assign n8108 = RESET_pad & \WX9722_reg/NET0131  ;
  assign n8109 = RESET_pad & \WX9840_reg/NET0131  ;
  assign n8110 = RESET_pad & \WX9764_reg/NET0131  ;
  assign n8111 = RESET_pad & \WX2076_reg/NET0131  ;
  assign n8112 = RESET_pad & \WX7116_reg/NET0131  ;
  assign n8113 = RESET_pad & \WX9796_reg/NET0131  ;
  assign n8114 = RESET_pad & \WX9776_reg/NET0131  ;
  assign n8115 = RESET_pad & \WX11071_reg/NET0131  ;
  assign n8116 = RESET_pad & \WX9760_reg/NET0131  ;
  assign n8117 = RESET_pad & \WX4576_reg/NET0131  ;
  assign n8118 = RESET_pad & \WX803_reg/NET0131  ;
  assign n8119 = RESET_pad & \WX3395_reg/NET0131  ;
  assign n8120 = RESET_pad & \WX4526_reg/NET0131  ;
  assign n8121 = RESET_pad & \WX9790_reg/NET0131  ;
  assign n8122 = RESET_pad & \WX9768_reg/NET0131  ;
  assign n8123 = RESET_pad & \WX653_reg/NET0131  ;
  assign n8124 = RESET_pad & \WX4662_reg/NET0131  ;
  assign n8125 = RESET_pad & \WX4580_reg/NET0131  ;
  assign n8126 = RESET_pad & \WX9728_reg/NET0131  ;
  assign n8127 = RESET_pad & \WX9718_reg/NET0131  ;
  assign n8128 = RESET_pad & \WX3405_reg/NET0131  ;
  assign n8129 = RESET_pad & \WX3245_reg/NET0131  ;
  assign n8130 = RESET_pad & \WX2010_reg/NET0131  ;
  assign n8131 = RESET_pad & \WX4682_reg/NET0131  ;
  assign n8132 = RESET_pad & \WX8589_reg/NET0131  ;
  assign n8133 = RESET_pad & \WX4688_reg/NET0131  ;
  assign n8134 = RESET_pad & \WX9706_reg/NET0131  ;
  assign n8135 = RESET_pad & \WX4690_reg/NET0131  ;
  assign n8136 = RESET_pad & \WX3243_reg/NET0131  ;
  assign n8137 = RESET_pad & \WX3241_reg/NET0131  ;
  assign n8138 = RESET_pad & \WX4698_reg/NET0131  ;
  assign n8139 = RESET_pad & \WX8591_reg/NET0131  ;
  assign n8140 = RESET_pad & \WX3239_reg/NET0131  ;
  assign n8141 = RESET_pad & \WX4704_reg/NET0131  ;
  assign n8142 = RESET_pad & \WX8583_reg/NET0131  ;
  assign n8143 = RESET_pad & \WX11029_reg/NET0131  ;
  assign n8144 = RESET_pad & \WX4712_reg/NET0131  ;
  assign n8145 = RESET_pad & \WX743_reg/NET0131  ;
  assign n8146 = RESET_pad & \WX8565_reg/NET0131  ;
  assign n8147 = RESET_pad & \WX8579_reg/NET0131  ;
  assign n8148 = RESET_pad & \WX3383_reg/NET0131  ;
  assign n8149 = RESET_pad & \WX8559_reg/NET0131  ;
  assign n8150 = RESET_pad & \WX2104_reg/NET0131  ;
  assign n8151 = RESET_pad & \WX4678_reg/NET0131  ;
  assign n8152 = RESET_pad & \WX689_reg/NET0131  ;
  assign n8153 = RESET_pad & \WX3233_reg/NET0131  ;
  assign n8154 = RESET_pad & \WX3393_reg/NET0131  ;
  assign n8155 = RESET_pad & \WX8455_reg/NET0131  ;
  assign n8156 = RESET_pad & \WX3235_reg/NET0131  ;
  assign n8157 = RESET_pad & \WX739_reg/NET0131  ;
  assign n8158 = RESET_pad & \WX8567_reg/NET0131  ;
  assign n8159 = RESET_pad & \WX8573_reg/NET0131  ;
  assign n8160 = RESET_pad & \WX3391_reg/NET0131  ;
  assign n8161 = RESET_pad & \WX10995_reg/NET0131  ;
  assign n8162 = RESET_pad & \WX8571_reg/NET0131  ;
  assign n8163 = RESET_pad & \WX2108_reg/NET0131  ;
  assign n8164 = RESET_pad & \WX2008_reg/NET0131  ;
  assign n8165 = RESET_pad & \WX7242_reg/NET0131  ;
  assign n8166 = RESET_pad & \WX11015_reg/NET0131  ;
  assign n8167 = RESET_pad & \WX9864_reg/NET0131  ;
  assign n8168 = RESET_pad & \WX3385_reg/NET0131  ;
  assign n8169 = RESET_pad & \WX4710_reg/NET0131  ;
  assign n8170 = RESET_pad & \WX779_reg/NET0131  ;
  assign n8171 = RESET_pad & \WX753_reg/NET0131  ;
  assign n8172 = RESET_pad & \WX733_reg/NET0131  ;
  assign n8173 = RESET_pad & \WX2012_reg/NET0131  ;
  assign n8174 = RESET_pad & \WX2086_reg/NET0131  ;
  assign n8175 = RESET_pad & \WX4680_reg/NET0131  ;
  assign n8176 = RESET_pad & \WX4696_reg/NET0131  ;
  assign n8177 = RESET_pad & \WX8561_reg/NET0131  ;
  assign n8178 = RESET_pad & \WX11077_reg/NET0131  ;
  assign n8179 = RESET_pad & \WX2106_reg/NET0131  ;
  assign n8180 = RESET_pad & \WX4686_reg/NET0131  ;
  assign n8181 = RESET_pad & \WX3335_reg/NET0131  ;
  assign n8182 = RESET_pad & \WX4666_reg/NET0131  ;
  assign n8183 = RESET_pad & \WX9830_reg/NET0131  ;
  assign n8184 = RESET_pad & \WX9788_reg/NET0131  ;
  assign n8185 = RESET_pad & \WX4674_reg/NET0131  ;
  assign n8186 = RESET_pad & \WX9838_reg/NET0131  ;
  assign n8187 = RESET_pad & \WX4670_reg/NET0131  ;
  assign n8188 = RESET_pad & \WX3253_reg/NET0131  ;
  assign n8189 = RESET_pad & \WX4664_reg/NET0131  ;
  assign n8190 = RESET_pad & \WX7296_reg/NET0131  ;
  assign n8191 = RESET_pad & \WX4660_reg/NET0131  ;
  assign n8192 = RESET_pad & \WX9696_reg/NET0131  ;
  assign n8193 = RESET_pad & \WX4566_reg/NET0131  ;
  assign n8194 = RESET_pad & \WX11001_reg/NET0131  ;
  assign n8195 = RESET_pad & \WX9812_reg/NET0131  ;
  assign n8196 = RESET_pad & \WX4620_reg/NET0131  ;
  assign n8197 = RESET_pad & \WX3407_reg/NET0131  ;
  assign n8198 = RESET_pad & \WX821_reg/NET0131  ;
  assign n8199 = RESET_pad & \WX8531_reg/NET0131  ;
  assign n8200 = RESET_pad & \WX2102_reg/NET0131  ;
  assign n8201 = RESET_pad & \WX649_reg/NET0131  ;
  assign n8202 = RESET_pad & \WX829_reg/NET0131  ;
  assign n8203 = RESET_pad & \WX8555_reg/NET0131  ;
  assign n8204 = RESET_pad & \WX3295_reg/NET0131  ;
  assign n8205 = RESET_pad & \WX2100_reg/NET0131  ;
  assign n8206 = RESET_pad & \WX825_reg/NET0131  ;
  assign n8207 = RESET_pad & \WX11017_reg/NET0131  ;
  assign n8208 = RESET_pad & \WX5951_reg/NET0131  ;
  assign n8209 = RESET_pad & \WX2098_reg/NET0131  ;
  assign n8210 = RESET_pad & \WX3297_reg/NET0131  ;
  assign n8211 = RESET_pad & \WX5849_reg/NET0131  ;
  assign n8212 = RESET_pad & \WX8553_reg/NET0131  ;
  assign n8213 = RESET_pad & \WX2016_reg/NET0131  ;
  assign n8214 = RESET_pad & \WX11063_reg/NET0131  ;
  assign n8215 = RESET_pad & \WX9700_reg/NET0131  ;
  assign n8216 = RESET_pad & \WX8463_reg/NET0131  ;
  assign n8217 = RESET_pad & \WX2096_reg/NET0131  ;
  assign n8218 = RESET_pad & \WX3331_reg/NET0131  ;
  assign n8219 = RESET_pad & \WX3299_reg/NET0131  ;
  assign n8220 = RESET_pad & \WX8549_reg/NET0131  ;
  assign n8221 = RESET_pad & \WX795_reg/NET0131  ;
  assign n8222 = RESET_pad & \WX3375_reg/NET0131  ;
  assign n8223 = RESET_pad & \WX5859_reg/NET0131  ;
  assign n8224 = RESET_pad & \WX4548_reg/NET0131  ;
  assign n8225 = RESET_pad & \WX3419_reg/NET0131  ;
  assign n8226 = RESET_pad & \WX8545_reg/NET0131  ;
  assign n8227 = RESET_pad & \WX4622_reg/NET0131  ;
  assign n8228 = RESET_pad & \WX8539_reg/NET0131  ;
  assign n8229 = RESET_pad & \WX2094_reg/NET0131  ;
  assign n8230 = RESET_pad & \WX2048_reg/NET0131  ;
  assign n8231 = RESET_pad & \WX723_reg/NET0131  ;
  assign n8232 = RESET_pad & \WX4600_reg/NET0131  ;
  assign n8233 = RESET_pad & \WX4602_reg/NET0131  ;
  assign n8234 = RESET_pad & \WX8405_reg/NET0131  ;
  assign n8235 = RESET_pad & \WX4650_reg/NET0131  ;
  assign n8236 = RESET_pad & \WX8543_reg/NET0131  ;
  assign n8237 = RESET_pad & \WX10997_reg/NET0131  ;
  assign n8238 = RESET_pad & \WX7282_reg/NET0131  ;
  assign n8239 = RESET_pad & \WX9884_reg/NET0131  ;
  assign n8240 = RESET_pad & \WX5899_reg/NET0131  ;
  assign n8241 = RESET_pad & \WX3369_reg/NET0131  ;
  assign n8242 = RESET_pad & \WX4616_reg/NET0131  ;
  assign n8243 = RESET_pad & \WX8457_reg/NET0131  ;
  assign n8244 = RESET_pad & \WX5855_reg/NET0131  ;
  assign n8245 = RESET_pad & \WX8435_reg/NET0131  ;
  assign n8246 = RESET_pad & \WX759_reg/NET0131  ;
  assign n8247 = RESET_pad & \WX8537_reg/NET0131  ;
  assign n8248 = RESET_pad & \WX9854_reg/NET0131  ;
  assign n8249 = RESET_pad & \WX10999_reg/NET0131  ;
  assign n8250 = RESET_pad & \WX7250_reg/NET0131  ;
  assign n8251 = RESET_pad & \WX1978_reg/NET0131  ;
  assign n8252 = RESET_pad & \WX651_reg/NET0131  ;
  assign n8253 = RESET_pad & \WX3387_reg/NET0131  ;
  assign n8254 = RESET_pad & \WX681_reg/NET0131  ;
  assign n8255 = RESET_pad & \WX8535_reg/NET0131  ;
  assign n8256 = RESET_pad & \WX7212_reg/NET0131  ;
  assign n8257 = RESET_pad & \WX5981_reg/NET0131  ;
  assign n8258 = RESET_pad & \WX4586_reg/NET0131  ;
  assign n8259 = RESET_pad & \WX4656_reg/NET0131  ;
  assign n8260 = RESET_pad & \WX3333_reg/NET0131  ;
  assign n8261 = RESET_pad & \WX9826_reg/NET0131  ;
  assign n8262 = RESET_pad & \WX2092_reg/NET0131  ;
  assign n8263 = RESET_pad & \WX4624_reg/NET0131  ;
  assign n8264 = RESET_pad & \WX7136_reg/NET0131  ;
  assign n8265 = RESET_pad & \WX7268_reg/NET0131  ;
  assign n8266 = RESET_pad & \WX4642_reg/NET0131  ;
  assign n8267 = RESET_pad & \WX8409_reg/NET0131  ;
  assign n8268 = RESET_pad & \WX4618_reg/NET0131  ;
  assign n8269 = RESET_pad & \WX4612_reg/NET0131  ;
  assign n8270 = RESET_pad & \WX7292_reg/NET0131  ;
  assign n8271 = RESET_pad & \WX3231_reg/NET0131  ;
  assign n8272 = RESET_pad & \WX8489_reg/NET0131  ;
  assign n8273 = RESET_pad & \WX3305_reg/NET0131  ;
  assign n8274 = RESET_pad & \WX8525_reg/NET0131  ;
  assign n8275 = RESET_pad & \WX11159_reg/NET0131  ;
  assign n8276 = RESET_pad & \WX3367_reg/NET0131  ;
  assign n8277 = RESET_pad & \WX11061_reg/NET0131  ;
  assign n8278 = RESET_pad & \WX8569_reg/NET0131  ;
  assign n8279 = RESET_pad & \WX11125_reg/NET0131  ;
  assign n8280 = RESET_pad & \WX809_reg/NET0131  ;
  assign n8281 = RESET_pad & \WX683_reg/NET0131  ;
  assign n8282 = RESET_pad & \WX8413_reg/NET0131  ;
  assign n8283 = RESET_pad & \WX2062_reg/NET0131  ;
  assign n8284 = RESET_pad & \WX9758_reg/NET0131  ;
  assign n8285 = RESET_pad & \WX3397_reg/NET0131  ;
  assign n8286 = RESET_pad & \WX7300_reg/NET0131  ;
  assign n8287 = RESET_pad & \WX6003_reg/NET0131  ;
  assign n8288 = RESET_pad & \WX4646_reg/NET0131  ;
  assign n8289 = RESET_pad & \WX9880_reg/NET0131  ;
  assign n8290 = RESET_pad & \WX7258_reg/NET0131  ;
  assign n8291 = RESET_pad & \WX8593_reg/NET0131  ;
  assign n8292 = RESET_pad & \WX11057_reg/NET0131  ;
  assign n8293 = RESET_pad & \WX675_reg/NET0131  ;
  assign n8294 = RESET_pad & \WX3371_reg/NET0131  ;
  assign n8295 = RESET_pad & \WX783_reg/NET0131  ;
  assign n8296 = RESET_pad & \WX8411_reg/NET0131  ;
  assign n8297 = RESET_pad & \WX9836_reg/NET0131  ;
  assign n8298 = RESET_pad & \WX11055_reg/NET0131  ;
  assign n8299 = RESET_pad & \WX8467_reg/NET0131  ;
  assign n8300 = RESET_pad & \WX817_reg/NET0131  ;
  assign n8301 = RESET_pad & \WX9870_reg/NET0131  ;
  assign n8302 = RESET_pad & \WX7262_reg/NET0131  ;
  assign n8303 = RESET_pad & \WX7264_reg/NET0131  ;
  assign n8304 = RESET_pad & \WX4604_reg/NET0131  ;
  assign n8305 = RESET_pad & \WX9804_reg/NET0131  ;
  assign n8306 = RESET_pad & \WX8429_reg/NET0131  ;
  assign n8307 = RESET_pad & \WX815_reg/NET0131  ;
  assign n8308 = RESET_pad & \WX5877_reg/NET0131  ;
  assign n8309 = RESET_pad & \WX6001_reg/NET0131  ;
  assign n8310 = RESET_pad & \WX8521_reg/NET0131  ;
  assign n8311 = RESET_pad & \WX7270_reg/NET0131  ;
  assign n8312 = RESET_pad & \WX677_reg/NET0131  ;
  assign n8313 = RESET_pad & \WX5989_reg/NET0131  ;
  assign n8314 = RESET_pad & \WX5993_reg/NET0131  ;
  assign n8315 = RESET_pad & \WX3303_reg/NET0131  ;
  assign n8316 = RESET_pad & \WX7142_reg/NET0131  ;
  assign n8317 = RESET_pad & \WX793_reg/NET0131  ;
  assign n8318 = RESET_pad & \WX9756_reg/NET0131  ;
  assign n8319 = RESET_pad & \WX7260_reg/NET0131  ;
  assign n8320 = RESET_pad & \WX5903_reg/NET0131  ;
  assign n8321 = RESET_pad & \WX11065_reg/NET0131  ;
  assign n8322 = RESET_pad & \WX4534_reg/NET0131  ;
  assign n8323 = RESET_pad & \WX4546_reg/NET0131  ;
  assign n8324 = RESET_pad & \WX2074_reg/NET0131  ;
  assign n8325 = RESET_pad & \WX8483_reg/NET0131  ;
  assign n8326 = RESET_pad & \WX3307_reg/NET0131  ;
  assign n8327 = RESET_pad & \WX9866_reg/NET0131  ;
  assign n8328 = RESET_pad & \WX4610_reg/NET0131  ;
  assign n8329 = RESET_pad & \WX4582_reg/NET0131  ;
  assign n8330 = RESET_pad & \WX5987_reg/NET0131  ;
  assign n8331 = RESET_pad & \WX11051_reg/NET0131  ;
  assign n8332 = RESET_pad & \WX4640_reg/NET0131  ;
  assign n8333 = RESET_pad & \WX655_reg/NET0131  ;
  assign n8334 = RESET_pad & \WX4596_reg/NET0131  ;
  assign n8335 = RESET_pad & \WX673_reg/NET0131  ;
  assign n8336 = RESET_pad & \WX4592_reg/NET0131  ;
  assign n8337 = RESET_pad & \WX7298_reg/NET0131  ;
  assign n8338 = RESET_pad & \WX2078_reg/NET0131  ;
  assign n8339 = RESET_pad & \WX2038_reg/NET0131  ;
  assign n8340 = RESET_pad & \WX11003_reg/NET0131  ;
  assign n8341 = RESET_pad & \WX5881_reg/NET0131  ;
  assign n8342 = RESET_pad & \WX4644_reg/NET0131  ;
  assign n8343 = RESET_pad & \WX2120_reg/NET0131  ;
  assign n8344 = RESET_pad & \WX4654_reg/NET0131  ;
  assign n8345 = RESET_pad & \WX3353_reg/NET0131  ;
  assign n8346 = RESET_pad & \WX5983_reg/NET0131  ;
  assign n8347 = RESET_pad & \WX4572_reg/NET0131  ;
  assign n8348 = RESET_pad & \WX8427_reg/NET0131  ;
  assign n8349 = RESET_pad & \WX4684_reg/NET0131  ;
  assign n8350 = RESET_pad & \WX4694_reg/NET0131  ;
  assign n8351 = RESET_pad & \WX833_reg/NET0131  ;
  assign n8352 = RESET_pad & \WX9886_reg/NET0131  ;
  assign n8353 = RESET_pad & \WX4552_reg/NET0131  ;
  assign n8354 = RESET_pad & \WX4606_reg/NET0131  ;
  assign n8355 = RESET_pad & \WX4536_reg/NET0131  ;
  assign n8356 = RESET_pad & \WX7140_reg/NET0131  ;
  assign n8357 = RESET_pad & \WX5975_reg/NET0131  ;
  assign n8358 = RESET_pad & \WX2110_reg/NET0131  ;
  assign n8359 = RESET_pad & \WX7274_reg/NET0131  ;
  assign n8360 = RESET_pad & \WX5977_reg/NET0131  ;
  assign n8361 = RESET_pad & \WX3417_reg/NET0131  ;
  assign n8362 = RESET_pad & \WX8507_reg/NET0131  ;
  assign n8363 = RESET_pad & \WX9720_reg/NET0131  ;
  assign n8364 = RESET_pad & \WX5971_reg/NET0131  ;
  assign n8365 = RESET_pad & \WX5967_reg/NET0131  ;
  assign n8366 = RESET_pad & \WX7146_reg/NET0131  ;
  assign n8367 = RESET_pad & \WX8541_reg/NET0131  ;
  assign n8368 = RESET_pad & \WX5969_reg/NET0131  ;
  assign n8369 = RESET_pad & \WX3373_reg/NET0131  ;
  assign n8370 = RESET_pad & \WX5963_reg/NET0131  ;
  assign n8371 = RESET_pad & \WX8513_reg/NET0131  ;
  assign n8372 = RESET_pad & \WX8509_reg/NET0131  ;
  assign n8373 = RESET_pad & \WX8433_reg/NET0131  ;
  assign n8374 = RESET_pad & \WX11047_reg/NET0131  ;
  assign n8375 = RESET_pad & \WX1942_reg/NET0131  ;
  assign n8376 = RESET_pad & \WX5961_reg/NET0131  ;
  assign n8377 = RESET_pad & \WX8511_reg/NET0131  ;
  assign n8378 = RESET_pad & \WX8431_reg/NET0131  ;
  assign n8379 = RESET_pad & \WX7286_reg/NET0131  ;
  assign n8380 = RESET_pad & \WX7288_reg/NET0131  ;
  assign n8381 = RESET_pad & \WX3343_reg/NET0131  ;
  assign n8382 = RESET_pad & \WX7112_reg/NET0131  ;
  assign n8383 = RESET_pad & \WX9766_reg/NET0131  ;
  assign n8384 = RESET_pad & \WX3315_reg/NET0131  ;
  assign n8385 = RESET_pad & \WX2070_reg/NET0131  ;
  assign n8386 = RESET_pad & \WX11091_reg/NET0131  ;
  assign n8387 = RESET_pad & \WX3377_reg/NET0131  ;
  assign n8388 = RESET_pad & \WX5943_reg/NET0131  ;
  assign n8389 = RESET_pad & \WX8479_reg/NET0131  ;
  assign n8390 = RESET_pad & \WX1948_reg/NET0131  ;
  assign n8391 = RESET_pad & \WX747_reg/NET0131  ;
  assign n8392 = RESET_pad & \WX8439_reg/NET0131  ;
  assign n8393 = RESET_pad & \WX9738_reg/NET0131  ;
  assign n8394 = RESET_pad & \WX9858_reg/NET0131  ;
  assign n8395 = RESET_pad & \WX7216_reg/NET0131  ;
  assign n8396 = RESET_pad & \WX2022_reg/NET0131  ;
  assign n8397 = RESET_pad & \WX4702_reg/NET0131  ;
  assign n8398 = RESET_pad & \WX4524_reg/NET0131  ;
  assign n8399 = RESET_pad & \WX5853_reg/NET0131  ;
  assign n8400 = RESET_pad & \WX5889_reg/NET0131  ;
  assign n8401 = RESET_pad & \WX8477_reg/NET0131  ;
  assign n8402 = RESET_pad & \WX4608_reg/NET0131  ;
  assign n8403 = RESET_pad & \WX5915_reg/NET0131  ;
  assign n8404 = RESET_pad & \WX8495_reg/NET0131  ;
  assign n8405 = RESET_pad & \WX3313_reg/NET0131  ;
  assign n8406 = RESET_pad & \WX8437_reg/NET0131  ;
  assign n8407 = RESET_pad & \WX5935_reg/NET0131  ;
  assign n8408 = RESET_pad & \WX715_reg/NET0131  ;
  assign n8409 = RESET_pad & \WX8501_reg/NET0131  ;
  assign n8410 = RESET_pad & \WX11009_reg/NET0131  ;
  assign n8411 = RESET_pad & \WX5931_reg/NET0131  ;
  assign n8412 = RESET_pad & \WX4590_reg/NET0131  ;
  assign n8413 = RESET_pad & \WX2124_reg/NET0131  ;
  assign n8414 = RESET_pad & \WX775_reg/NET0131  ;
  assign n8415 = RESET_pad & \WX9792_reg/NET0131  ;
  assign n8416 = RESET_pad & \WX811_reg/NET0131  ;
  assign n8417 = RESET_pad & \WX8499_reg/NET0131  ;
  assign n8418 = RESET_pad & \WX10991_reg/NET0131  ;
  assign n8419 = RESET_pad & \WX7162_reg/NET0131  ;
  assign n8420 = RESET_pad & \WX3411_reg/NET0131  ;
  assign n8421 = RESET_pad & \WX8497_reg/NET0131  ;
  assign n8422 = RESET_pad & \WX703_reg/NET0131  ;
  assign n8423 = RESET_pad & \WX5917_reg/NET0131  ;
  assign n8424 = RESET_pad & \WX11157_reg/NET0131  ;
  assign n8425 = RESET_pad & \WX1970_reg/NET0131  ;
  assign n8426 = RESET_pad & \WX1974_reg/NET0131  ;
  assign n8427 = RESET_pad & \WX8493_reg/NET0131  ;
  assign n8428 = RESET_pad & \WX9828_reg/NET0131  ;
  assign n8429 = RESET_pad & \WX5911_reg/NET0131  ;
  assign n8430 = RESET_pad & \WX797_reg/NET0131  ;
  assign n8431 = RESET_pad & \WX1962_reg/NET0131  ;
  assign n8432 = RESET_pad & \WX2040_reg/NET0131  ;
  assign n8433 = RESET_pad & \WX827_reg/NET0131  ;
  assign n8434 = RESET_pad & \WX8487_reg/NET0131  ;
  assign n8435 = RESET_pad & \WX5913_reg/NET0131  ;
  assign n8436 = RESET_pad & \WX1952_reg/NET0131  ;
  assign n8437 = RESET_pad & \WX5905_reg/NET0131  ;
  assign n8438 = RESET_pad & \WX3345_reg/NET0131  ;
  assign n8439 = RESET_pad & \WX9748_reg/NET0131  ;
  assign n8440 = RESET_pad & \WX2058_reg/NET0131  ;
  assign n8441 = RESET_pad & \WX5907_reg/NET0131  ;
  assign n8442 = RESET_pad & \WX3249_reg/NET0131  ;
  assign n8443 = RESET_pad & \WX1944_reg/NET0131  ;
  assign n8444 = RESET_pad & \WX4630_reg/NET0131  ;
  assign n8445 = RESET_pad & \WX5895_reg/NET0131  ;
  assign n8446 = RESET_pad & \WX5887_reg/NET0131  ;
  assign n8447 = RESET_pad & \WX1938_reg/NET0131  ;
  assign n8448 = RESET_pad & \WX1940_reg/NET0131  ;
  assign n8449 = RESET_pad & \WX8403_reg/NET0131  ;
  assign n8450 = RESET_pad & \WX725_reg/NET0131  ;
  assign n8451 = RESET_pad & \WX5897_reg/NET0131  ;
  assign n8452 = RESET_pad & \WX11173_reg/NET0131  ;
  assign n8453 = RESET_pad & \WX8425_reg/NET0131  ;
  assign n8454 = RESET_pad & \WX7170_reg/NET0131  ;
  assign n8455 = RESET_pad & \WX8465_reg/NET0131  ;
  assign n8456 = RESET_pad & \WX4530_reg/NET0131  ;
  assign n8457 = RESET_pad & \WX7172_reg/NET0131  ;
  assign n8458 = RESET_pad & \WX5893_reg/NET0131  ;
  assign n8459 = RESET_pad & \WX785_reg/NET0131  ;
  assign n8460 = RESET_pad & \WX2050_reg/NET0131  ;
  assign n8461 = RESET_pad & \WX8585_reg/NET0131  ;
  assign n8462 = RESET_pad & \WX8587_reg/NET0131  ;
  assign n8463 = RESET_pad & \WX5891_reg/NET0131  ;
  assign n8464 = RESET_pad & \WX671_reg/NET0131  ;
  assign n8465 = RESET_pad & \WX2028_reg/NET0131  ;
  assign n8466 = RESET_pad & \WX11097_reg/NET0131  ;
  assign n8467 = RESET_pad & \WX2116_reg/NET0131  ;
  assign n8468 = RESET_pad & \WX11151_reg/NET0131  ;
  assign n8469 = RESET_pad & \WX679_reg/NET0131  ;
  assign n8470 = RESET_pad & \WX2024_reg/NET0131  ;
  assign n8471 = RESET_pad & \WX4706_reg/NET0131  ;
  assign n8472 = RESET_pad & \WX7168_reg/NET0131  ;
  assign n8473 = RESET_pad & \WX4554_reg/NET0131  ;
  assign n8474 = RESET_pad & \WX8421_reg/NET0131  ;
  assign n8475 = RESET_pad & \WX2090_reg/NET0131  ;
  assign n8476 = RESET_pad & \WX9784_reg/NET0131  ;
  assign n8477 = RESET_pad & \WX4714_reg/NET0131  ;
  assign n8478 = RESET_pad & \WX11013_reg/NET0131  ;
  assign n8479 = RESET_pad & \WX2052_reg/NET0131  ;
  assign n8480 = RESET_pad & \WX8417_reg/NET0131  ;
  assign n8481 = RESET_pad & \WX3341_reg/NET0131  ;
  assign n8482 = RESET_pad & \WX5883_reg/NET0131  ;
  assign n8483 = RESET_pad & \WX3323_reg/NET0131  ;
  assign n8484 = RESET_pad & \WX9868_reg/NET0131  ;
  assign n8485 = RESET_pad & \WX8461_reg/NET0131  ;
  assign n8486 = RESET_pad & \WX3329_reg/NET0131  ;
  assign n8487 = RESET_pad & \WX11171_reg/NET0131  ;
  assign n8488 = RESET_pad & \WX9734_reg/NET0131  ;
  assign n8489 = RESET_pad & \WX7176_reg/NET0131  ;
  assign n8490 = RESET_pad & \WX2018_reg/NET0131  ;
  assign n8491 = RESET_pad & \WX9834_reg/NET0131  ;
  assign n8492 = RESET_pad & \WX3401_reg/NET0131  ;
  assign n8493 = RESET_pad & \WX2006_reg/NET0131  ;
  assign n8494 = RESET_pad & \WX3337_reg/NET0131  ;
  assign n8495 = RESET_pad & \WX8503_reg/NET0131  ;
  assign n8496 = RESET_pad & \WX5867_reg/NET0131  ;
  assign n8497 = RESET_pad & \WX6005_reg/NET0131  ;
  assign n8498 = RESET_pad & \WX11025_reg/NET0131  ;
  assign n8499 = RESET_pad & \WX1990_reg/NET0131  ;
  assign n8500 = RESET_pad & \WX5831_reg/NET0131  ;
  assign n8501 = RESET_pad & \WX5955_reg/NET0131  ;
  assign n8502 = RESET_pad & \WX8523_reg/NET0131  ;
  assign n8503 = RESET_pad & \WX2084_reg/NET0131  ;
  assign n8504 = RESET_pad & \WX789_reg/NET0131  ;
  assign n8505 = RESET_pad & \WX3381_reg/NET0131  ;
  assign n8506 = RESET_pad & \WX5865_reg/NET0131  ;
  assign n8507 = RESET_pad & \WX5885_reg/NET0131  ;
  assign n8508 = RESET_pad & \WX9794_reg/NET0131  ;
  assign n8509 = RESET_pad & \WX5819_reg/NET0131  ;
  assign n8510 = RESET_pad & \WX5863_reg/NET0131  ;
  assign n8511 = RESET_pad & \WX2042_reg/NET0131  ;
  assign n8512 = RESET_pad & \WX7178_reg/NET0131  ;
  assign n8513 = RESET_pad & \WX813_reg/NET0131  ;
  assign n8514 = RESET_pad & \WX5821_reg/NET0131  ;
  assign n8515 = RESET_pad & \WX5851_reg/NET0131  ;
  assign n8516 = RESET_pad & \WX8473_reg/NET0131  ;
  assign n8517 = RESET_pad & \WX4578_reg/NET0131  ;
  assign n8518 = RESET_pad & \WX3421_reg/NET0131  ;
  assign n8519 = RESET_pad & \WX9732_reg/NET0131  ;
  assign n8520 = RESET_pad & \WX11127_reg/NET0131  ;
  assign n8521 = RESET_pad & \WX5847_reg/NET0131  ;
  assign n8522 = RESET_pad & \WX8469_reg/NET0131  ;
  assign n8523 = RESET_pad & \WX763_reg/NET0131  ;
  assign n8524 = RESET_pad & \WX2036_reg/NET0131  ;
  assign n8525 = RESET_pad & \WX8475_reg/NET0131  ;
  assign n8526 = RESET_pad & \WX11021_reg/NET0131  ;
  assign n8527 = RESET_pad & \WX5901_reg/NET0131  ;
  assign n8528 = RESET_pad & \WX11005_reg/NET0131  ;
  assign n8529 = RESET_pad & \WX3275_reg/NET0131  ;
  assign n8530 = RESET_pad & \WX4632_reg/NET0131  ;
  assign n8531 = RESET_pad & \WX5841_reg/NET0131  ;
  assign n8532 = RESET_pad & \WX5973_reg/NET0131  ;
  assign n8533 = RESET_pad & \WX11019_reg/NET0131  ;
  assign n8534 = RESET_pad & \WX5829_reg/NET0131  ;
  assign n8535 = RESET_pad & \WX647_reg/NET0131  ;
  assign n8536 = RESET_pad & \WX5833_reg/NET0131  ;
  assign n8537 = RESET_pad & \WX5995_reg/NET0131  ;
  assign n8538 = RESET_pad & \WX3261_reg/NET0131  ;
  assign n8539 = RESET_pad & \WX7184_reg/NET0131  ;
  assign n8540 = RESET_pad & \WX11165_reg/NET0131  ;
  assign n8541 = RESET_pad & \WX8419_reg/NET0131  ;
  assign n8542 = RESET_pad & \WX697_reg/NET0131  ;
  assign n8543 = RESET_pad & \WX5823_reg/NET0131  ;
  assign n8544 = RESET_pad & \WX5857_reg/NET0131  ;
  assign n8545 = RESET_pad & \WX717_reg/NET0131  ;
  assign n8546 = RESET_pad & \WX4528_reg/NET0131  ;
  assign n8547 = RESET_pad & \WX5843_reg/NET0131  ;
  assign n8548 = RESET_pad & \WX5827_reg/NET0131  ;
  assign n8549 = RESET_pad & \WX7254_reg/NET0131  ;
  assign n8550 = RESET_pad & \WX5835_reg/NET0131  ;
  assign n8551 = RESET_pad & \WX737_reg/NET0131  ;
  assign n8552 = RESET_pad & \WX3293_reg/NET0131  ;
  assign n8553 = RESET_pad & \WX9846_reg/NET0131  ;
  assign n8554 = RESET_pad & \WX1964_reg/NET0131  ;
  assign n8555 = RESET_pad & \WX9814_reg/NET0131  ;
  assign n8556 = RESET_pad & \WX8505_reg/NET0131  ;
  assign n8557 = RESET_pad & \WX4658_reg/NET0131  ;
  assign n8558 = RESET_pad & \WX5825_reg/NET0131  ;
  assign n8559 = RESET_pad & \WX7188_reg/NET0131  ;
  assign n8560 = RESET_pad & \WX3399_reg/NET0131  ;
  assign n8561 = RESET_pad & \WX2034_reg/NET0131  ;
  assign n8562 = RESET_pad & \WX8471_reg/NET0131  ;
  assign n8563 = RESET_pad & \WX1968_reg/NET0131  ;
  assign n8564 = RESET_pad & \WX7290_reg/NET0131  ;
  assign n8565 = RESET_pad & \WX11101_reg/NET0131  ;
  assign n8566 = RESET_pad & \WX5837_reg/NET0131  ;
  assign n8567 = RESET_pad & \WX8459_reg/NET0131  ;
  assign n8568 = RESET_pad & \WX5817_reg/NET0131  ;
  assign n8569 = RESET_pad & \WX4668_reg/NET0131  ;
  assign n8570 = RESET_pad & \WX4614_reg/NET0131  ;
  assign n8571 = RESET_pad & \WX4672_reg/NET0131  ;
  assign n8572 = RESET_pad & \WX9844_reg/NET0131  ;
  assign n8573 = RESET_pad & \WX4648_reg/NET0131  ;
  assign n8574 = RESET_pad & \WX3325_reg/NET0131  ;
  assign n8575 = RESET_pad & \WX713_reg/NET0131  ;
  assign n8576 = RESET_pad & \WX11069_reg/NET0131  ;
  assign n8577 = RESET_pad & \WX9746_reg/NET0131  ;
  assign n8578 = RESET_pad & \WX9874_reg/NET0131  ;
  assign n8579 = RESET_pad & \WX8451_reg/NET0131  ;
  assign n8580 = RESET_pad & \WX1950_reg/NET0131  ;
  assign n8581 = RESET_pad & \WX5909_reg/NET0131  ;
  assign n8582 = RESET_pad & \WX8515_reg/NET0131  ;
  assign n8583 = RESET_pad & \WX1960_reg/NET0131  ;
  assign n8584 = RESET_pad & \WX7236_reg/NET0131  ;
  assign n8585 = RESET_pad & \WX4700_reg/NET0131  ;
  assign n8586 = RESET_pad & \WX4692_reg/NET0131  ;
  assign n8587 = RESET_pad & \WX1976_reg/NET0131  ;
  assign n8588 = RESET_pad & \WX1980_reg/NET0131  ;
  assign n8589 = RESET_pad & \WX8443_reg/NET0131  ;
  assign n8590 = RESET_pad & \WX1996_reg/NET0131  ;
  assign n8591 = RESET_pad & \WX2032_reg/NET0131  ;
  assign n8592 = RESET_pad & \WX9848_reg/NET0131  ;
  assign n8593 = RESET_pad & \WX11023_reg/NET0131  ;
  assign n8594 = RESET_pad & \WX3317_reg/NET0131  ;
  assign n8595 = RESET_pad & \WX9740_reg/NET0131  ;
  assign n8596 = RESET_pad & \WX2014_reg/NET0131  ;
  assign n8597 = RESET_pad & \WX11155_reg/NET0131  ;
  assign n8598 = RESET_pad & \WX2020_reg/NET0131  ;
  assign n8599 = RESET_pad & \WX6007_reg/NET0131  ;
  assign n8600 = RESET_pad & \WX4708_reg/NET0131  ;
  assign n8601 = RESET_pad & \WX2044_reg/NET0131  ;
  assign n8602 = RESET_pad & \WX2046_reg/NET0131  ;
  assign n8603 = RESET_pad & \WX3359_reg/NET0131  ;
  assign n8604 = RESET_pad & \WX2054_reg/NET0131  ;
  assign n8605 = RESET_pad & \WX5869_reg/NET0131  ;
  assign n8606 = RESET_pad & \WX11179_reg/NET0131  ;
  assign n8607 = RESET_pad & \WX11129_reg/NET0131  ;
  assign n8608 = RESET_pad & \WX11145_reg/NET0131  ;
  assign n8609 = RESET_pad & \WX699_reg/NET0131  ;
  assign n8610 = RESET_pad & \WX2080_reg/NET0131  ;
  assign n8611 = RESET_pad & \WX2082_reg/NET0131  ;
  assign n8612 = RESET_pad & \WX2030_reg/NET0131  ;
  assign n8613 = RESET_pad & \WX11075_reg/NET0131  ;
  assign n8614 = RESET_pad & \WX3311_reg/NET0131  ;
  assign n8615 = RESET_pad & \WX9818_reg/NET0131  ;
  assign n8616 = RESET_pad & \WX701_reg/NET0131  ;
  assign n8617 = RESET_pad & \WX2026_reg/NET0131  ;
  assign n8618 = RESET_pad & \WX5839_reg/NET0131  ;
  assign n8619 = RESET_pad & \WX11007_reg/NET0131  ;
  assign n8620 = RESET_pad & \WX8563_reg/NET0131  ;
  assign n8621 = RESET_pad & \WX3309_reg/NET0131  ;
  assign n8622 = RESET_pad & \WX9710_reg/NET0131  ;
  assign n8623 = RESET_pad & \WX4574_reg/NET0131  ;
  assign n8624 = RESET_pad & \WX7202_reg/NET0131  ;
  assign n8625 = RESET_pad & \WX8415_reg/NET0131  ;
  assign n8626 = RESET_pad & \WX9810_reg/NET0131  ;
  assign n8627 = RESET_pad & \WX3269_reg/NET0131  ;
  assign n8628 = RESET_pad & \WX7200_reg/NET0131  ;
  assign n8629 = RESET_pad & \WX9752_reg/NET0131  ;
  assign n8630 = RESET_pad & \WX7174_reg/NET0131  ;
  assign n8631 = RESET_pad & \WX3389_reg/NET0131  ;
  assign n8632 = RESET_pad & \WX8581_reg/NET0131  ;
  assign n8633 = RESET_pad & \WX5845_reg/NET0131  ;
  assign n8634 = RESET_pad & \WX5873_reg/NET0131  ;
  assign n8635 = RESET_pad & \WX9782_reg/NET0131  ;
  assign n8636 = RESET_pad & \WX7208_reg/NET0131  ;
  assign n8637 = RESET_pad & \WX8485_reg/NET0131  ;
  assign n8638 = RESET_pad & \WX8575_reg/NET0131  ;
  assign n8639 = RESET_pad & \WX8481_reg/NET0131  ;
  assign n8640 = RESET_pad & \WX4532_reg/NET0131  ;
  assign n8641 = RESET_pad & \WX11031_reg/NET0131  ;
  assign n8642 = RESET_pad & \WX7210_reg/NET0131  ;
  assign n8643 = RESET_pad & \WX7206_reg/NET0131  ;
  assign n8644 = RESET_pad & \WX10989_reg/NET0131  ;
  assign n8645 = RESET_pad & \WX765_reg/NET0131  ;
  assign n8646 = RESET_pad & \WX799_reg/NET0131  ;
  assign n8647 = RESET_pad & \WX711_reg/NET0131  ;
  assign n8648 = RESET_pad & \WX751_reg/NET0131  ;
  assign n8649 = RESET_pad & \WX10993_reg/NET0131  ;
  assign n8650 = RESET_pad & \WX3413_reg/NET0131  ;
  assign n8651 = RESET_pad & \WX8577_reg/NET0131  ;
  assign n8652 = RESET_pad & \WX3291_reg/NET0131  ;
  assign n8653 = RESET_pad & \WX741_reg/NET0131  ;
  assign n8654 = RESET_pad & \WX749_reg/NET0131  ;
  assign n8655 = RESET_pad & \WX7266_reg/NET0131  ;
  assign n8656 = RESET_pad & \WX4568_reg/NET0131  ;
  assign n8657 = RESET_pad & \WX8527_reg/NET0131  ;
  assign n8658 = RESET_pad & \WX1982_reg/NET0131  ;
  assign n8659 = RESET_pad & \WX11035_reg/NET0131  ;
  assign n8660 = RESET_pad & \WX11039_reg/NET0131  ;
  assign n8661 = RESET_pad & \WX3251_reg/NET0131  ;
  assign n8662 = RESET_pad & \WX745_reg/NET0131  ;
  assign n8663 = ~\TM0_pad  & ~n1543 ;
  assign n8664 = n2846 & ~n8663 ;
  assign n8665 = \TM0_pad  & ~\_2088__reg/NET0131  ;
  assign n8666 = n1976 & ~n8665 ;
  assign n8667 = ~n5074 & n8666 ;
  assign n8668 = ~n8664 & ~n8667 ;
  assign n8669 = ~\TM0_pad  & ~n1955 ;
  assign n8670 = n2023 & ~n8669 ;
  assign n8671 = \TM0_pad  & ~\_2085__reg/NET0131  ;
  assign n8672 = n1976 & ~n8671 ;
  assign n8673 = ~n5455 & n8672 ;
  assign n8674 = ~n8670 & ~n8673 ;
  assign n8675 = ~\TM0_pad  & ~n1903 ;
  assign n8676 = n3953 & ~n8675 ;
  assign n8677 = \TM0_pad  & ~\_2081__reg/NET0131  ;
  assign n8678 = n1976 & ~n8677 ;
  assign n8679 = ~n5995 & n8678 ;
  assign n8680 = ~n8676 & ~n8679 ;
  assign n8681 = ~\TM0_pad  & ~n1582 ;
  assign n8682 = n2341 & ~n8681 ;
  assign n8683 = \TM0_pad  & ~\_2091__reg/NET0131  ;
  assign n8684 = n1976 & ~n8683 ;
  assign n8685 = ~n4687 & n8684 ;
  assign n8686 = ~n8682 & ~n8685 ;
  assign n8687 = ~\TM0_pad  & ~n1968 ;
  assign n8688 = n3172 & ~n8687 ;
  assign n8689 = \TM0_pad  & ~\_2086__reg/NET0131  ;
  assign n8690 = n1976 & ~n8689 ;
  assign n8691 = ~n5332 & n8690 ;
  assign n8692 = ~n8688 & ~n8691 ;
  assign n8693 = ~\TM0_pad  & ~n1942 ;
  assign n8694 = n3483 & ~n8693 ;
  assign n8695 = \TM0_pad  & ~\_2084__reg/NET0131  ;
  assign n8696 = n1976 & ~n8695 ;
  assign n8697 = ~n5575 & n8696 ;
  assign n8698 = ~n8694 & ~n8697 ;
  assign n8699 = ~\TM0_pad  & ~n1672 ;
  assign n8700 = n4382 & ~n8699 ;
  assign n8701 = \TM0_pad  & ~\_2078__reg/NET0131  ;
  assign n8702 = n1976 & ~n8701 ;
  assign n8703 = ~n6508 & n8702 ;
  assign n8704 = ~n8700 & ~n8703 ;
  assign n8705 = n1974 & ~n3082 ;
  assign n8707 = \TM0_pad  & ~\_2348__reg/NET0131  ;
  assign n8706 = ~\DATA_0_15_pad  & ~\TM0_pad  ;
  assign n8708 = n1976 & ~n8706 ;
  assign n8709 = ~n8707 & n8708 ;
  assign n8710 = ~n8705 & ~n8709 ;
  assign \DATA_9_0_pad  = n1520 ;
  assign \DATA_9_10_pad  = n1533 ;
  assign \DATA_9_11_pad  = n1546 ;
  assign \DATA_9_12_pad  = n1559 ;
  assign \DATA_9_13_pad  = n1572 ;
  assign \DATA_9_14_pad  = n1585 ;
  assign \DATA_9_15_pad  = n1598 ;
  assign \DATA_9_16_pad  = ~n1614 ;
  assign \DATA_9_17_pad  = ~n1630 ;
  assign \DATA_9_18_pad  = ~n1646 ;
  assign \DATA_9_19_pad  = ~n1662 ;
  assign \DATA_9_1_pad  = n1675 ;
  assign \DATA_9_20_pad  = ~n1691 ;
  assign \DATA_9_21_pad  = ~n1707 ;
  assign \DATA_9_22_pad  = ~n1723 ;
  assign \DATA_9_23_pad  = ~n1739 ;
  assign \DATA_9_24_pad  = ~n1755 ;
  assign \DATA_9_25_pad  = ~n1771 ;
  assign \DATA_9_26_pad  = ~n1787 ;
  assign \DATA_9_27_pad  = ~n1803 ;
  assign \DATA_9_28_pad  = ~n1819 ;
  assign \DATA_9_29_pad  = ~n1835 ;
  assign \DATA_9_2_pad  = n1848 ;
  assign \DATA_9_30_pad  = ~n1864 ;
  assign \DATA_9_31_pad  = ~n1880 ;
  assign \DATA_9_3_pad  = n1893 ;
  assign \DATA_9_4_pad  = n1906 ;
  assign \DATA_9_5_pad  = n1919 ;
  assign \DATA_9_6_pad  = n1932 ;
  assign \DATA_9_7_pad  = n1945 ;
  assign \DATA_9_8_pad  = n1958 ;
  assign \DATA_9_9_pad  = n1971 ;
  assign \_al_n0  = 1'b0 ;
  assign \_al_n1  = ~1'b0 ;
  assign \g19/_0_  = ~n1990 ;
  assign \g35/_0_  = ~n2022 ;
  assign \g36/_0_  = ~n2039 ;
  assign \g40/_0_  = ~n2056 ;
  assign \g55780/_0_  = ~n2076 ;
  assign \g55783/_0_  = ~n2096 ;
  assign \g55795/_0_  = ~n2121 ;
  assign \g55796/_0_  = ~n2140 ;
  assign \g55797/_0_  = ~n2172 ;
  assign \g55798/_0_  = ~n2204 ;
  assign \g55799/_0_  = ~n2236 ;
  assign \g55800/_0_  = ~n2268 ;
  assign \g55801/_0_  = ~n2300 ;
  assign \g55802/_0_  = ~n2320 ;
  assign \g55803/_0_  = ~n2340 ;
  assign \g55834/_0_  = ~n2366 ;
  assign \g55835/_0_  = ~n2385 ;
  assign \g55836/_0_  = ~n2404 ;
  assign \g55837/_0_  = ~n2423 ;
  assign \g55838/_0_  = ~n2438 ;
  assign \g55839/_0_  = ~n2457 ;
  assign \g55840/_0_  = ~n2476 ;
  assign \g55841/_0_  = ~n2496 ;
  assign \g55842/_0_  = ~n2516 ;
  assign \g55856/_0_  = n2517 ;
  assign \g55894/_0_  = ~n2542 ;
  assign \g55895/_0_  = ~n2561 ;
  assign \g55896/_0_  = ~n2580 ;
  assign \g55897/_0_  = ~n2599 ;
  assign \g55898/_0_  = ~n2614 ;
  assign \g55899/_0_  = ~n2629 ;
  assign \g55900/_0_  = ~n2648 ;
  assign \g55901/_0_  = ~n2668 ;
  assign \g55902/_0_  = ~n2675 ;
  assign \g55916/_0_  = n2676 ;
  assign \g55953/_0_  = ~n2702 ;
  assign \g55954/_0_  = ~n2721 ;
  assign \g55955/_0_  = ~n2740 ;
  assign \g55956/_0_  = ~n2759 ;
  assign \g55957/_0_  = ~n2774 ;
  assign \g55958/_0_  = ~n2789 ;
  assign \g55959/_0_  = ~n2804 ;
  assign \g55960/_0_  = ~n2824 ;
  assign \g55961/_0_  = ~n2844 ;
  assign \g55975/_0_  = n2845 ;
  assign \g56012/_0_  = ~n2871 ;
  assign \g56013/_0_  = ~n2886 ;
  assign \g56014/_0_  = ~n2905 ;
  assign \g56015/_0_  = ~n2924 ;
  assign \g56016/_0_  = ~n2939 ;
  assign \g56017/_0_  = ~n2954 ;
  assign \g56018/_0_  = ~n2969 ;
  assign \g56019/_0_  = ~n2989 ;
  assign \g56020/_0_  = ~n3009 ;
  assign \g56034/_0_  = n3010 ;
  assign \g56071/_0_  = ~n3036 ;
  assign \g56072/_0_  = ~n3051 ;
  assign \g56073/_0_  = ~n3070 ;
  assign \g56074/_0_  = ~n3085 ;
  assign \g56075/_0_  = ~n3100 ;
  assign \g56076/_0_  = ~n3115 ;
  assign \g56077/_0_  = ~n3130 ;
  assign \g56078/_0_  = ~n3150 ;
  assign \g56079/_0_  = ~n3170 ;
  assign \g56093/_0_  = n3171 ;
  assign \g56130/_0_  = ~n3197 ;
  assign \g56131/_0_  = ~n3212 ;
  assign \g56132/_0_  = ~n3227 ;
  assign \g56133/_0_  = ~n3246 ;
  assign \g56134/_0_  = ~n3261 ;
  assign \g56135/_0_  = ~n3276 ;
  assign \g56136/_0_  = ~n3291 ;
  assign \g56137/_0_  = ~n3311 ;
  assign \g56138/_0_  = ~n3331 ;
  assign \g56152/_0_  = n3332 ;
  assign \g56189/_0_  = ~n3357 ;
  assign \g56190/_0_  = ~n3372 ;
  assign \g56191/_0_  = ~n3377 ;
  assign \g56192/_0_  = ~n3396 ;
  assign \g56193/_0_  = ~n3411 ;
  assign \g56194/_0_  = ~n3426 ;
  assign \g56195/_0_  = ~n3441 ;
  assign \g56196/_0_  = ~n3461 ;
  assign \g56197/_0_  = ~n3481 ;
  assign \g56211/_0_  = n3482 ;
  assign \g56248/_0_  = ~n3508 ;
  assign \g56249/_0_  = ~n3523 ;
  assign \g56250/_0_  = ~n3538 ;
  assign \g56251/_0_  = ~n3557 ;
  assign \g56252/_0_  = ~n3572 ;
  assign \g56253/_0_  = ~n3587 ;
  assign \g56254/_0_  = ~n3602 ;
  assign \g56255/_0_  = ~n3622 ;
  assign \g56256/_0_  = ~n3642 ;
  assign \g56270/_0_  = n3643 ;
  assign \g56307/_0_  = ~n3669 ;
  assign \g56308/_0_  = ~n3684 ;
  assign \g56309/_0_  = ~n3699 ;
  assign \g56310/_0_  = ~n3718 ;
  assign \g56311/_0_  = ~n3733 ;
  assign \g56312/_0_  = ~n3748 ;
  assign \g56313/_0_  = ~n3763 ;
  assign \g56314/_0_  = ~n3783 ;
  assign \g56315/_0_  = ~n3803 ;
  assign \g56329/_0_  = n3804 ;
  assign \g56366/_0_  = ~n3830 ;
  assign \g56367/_0_  = ~n3845 ;
  assign \g56368/_0_  = ~n3860 ;
  assign \g56369/_0_  = ~n3879 ;
  assign \g56370/_0_  = ~n3894 ;
  assign \g56371/_0_  = ~n3909 ;
  assign \g56372/_0_  = ~n3924 ;
  assign \g56373/_0_  = ~n3944 ;
  assign \g56374/_0_  = ~n3951 ;
  assign \g56388/_0_  = n3952 ;
  assign \g56425/_0_  = ~n3978 ;
  assign \g56426/_0_  = ~n3993 ;
  assign \g56427/_0_  = ~n4008 ;
  assign \g56428/_0_  = ~n4027 ;
  assign \g56429/_0_  = ~n4042 ;
  assign \g56430/_0_  = ~n4057 ;
  assign \g56431/_0_  = ~n4072 ;
  assign \g56432/_0_  = ~n4092 ;
  assign \g56433/_0_  = ~n4099 ;
  assign \g56447/_0_  = n4100 ;
  assign \g56484/_0_  = ~n4126 ;
  assign \g56485/_0_  = ~n4141 ;
  assign \g56486/_0_  = ~n4146 ;
  assign \g56487/_0_  = ~n4165 ;
  assign \g56488/_0_  = ~n4180 ;
  assign \g56489/_0_  = ~n4195 ;
  assign \g56490/_0_  = ~n4210 ;
  assign \g56491/_0_  = ~n4230 ;
  assign \g56492/_0_  = ~n4237 ;
  assign \g56507/_0_  = n4238 ;
  assign \g56543/_0_  = ~n4264 ;
  assign \g56544/_0_  = ~n4279 ;
  assign \g56545/_0_  = ~n4294 ;
  assign \g56546/_0_  = ~n4309 ;
  assign \g56547/_0_  = ~n4328 ;
  assign \g56548/_0_  = ~n4343 ;
  assign \g56549/_0_  = ~n4358 ;
  assign \g56551/_0_  = ~n4365 ;
  assign \g56567/_0_  = n4366 ;
  assign \g56602/_0_  = ~n4381 ;
  assign \g56603/_0_  = ~n4407 ;
  assign \g56604/_0_  = ~n4422 ;
  assign \g56605/_0_  = ~n4437 ;
  assign \g56606/_0_  = ~n4452 ;
  assign \g56607/_0_  = ~n4471 ;
  assign \g56608/_0_  = ~n4486 ;
  assign \g56610/_0_  = ~n4493 ;
  assign \g56627/_0_  = n4494 ;
  assign \g56661/_0_  = ~n4509 ;
  assign \g56662/_0_  = ~n4535 ;
  assign \g56663/_0_  = ~n4550 ;
  assign \g56664/_0_  = ~n4565 ;
  assign \g56665/_0_  = ~n4580 ;
  assign \g56666/_0_  = ~n4585 ;
  assign \g56667/_0_  = ~n4600 ;
  assign \g56668/_0_  = ~n4616 ;
  assign \g56686/_0_  = n4617 ;
  assign \g56720/_0_  = ~n4632 ;
  assign \g56721/_0_  = ~n4647 ;
  assign \g56722/_0_  = ~n4662 ;
  assign \g56723/_0_  = ~n4677 ;
  assign \g56724/_0_  = ~n4692 ;
  assign \g56725/_0_  = ~n4707 ;
  assign \g56726/_0_  = ~n4739 ;
  assign \g56727/_0_  = ~n4755 ;
  assign \g56728/_0_  = ~n4761 ;
  assign \g56745/_0_  = n4762 ;
  assign \g56779/_0_  = ~n4777 ;
  assign \g56780/_0_  = ~n4792 ;
  assign \g56781/_0_  = ~n4811 ;
  assign \g56782/_0_  = ~n4826 ;
  assign \g56783/_0_  = ~n4831 ;
  assign \g56784/_0_  = ~n4846 ;
  assign \g56785/_0_  = ~n4865 ;
  assign \g56804/_0_  = n4866 ;
  assign \g56838/_0_  = ~n4881 ;
  assign \g56839/_0_  = ~n4896 ;
  assign \g56840/_0_  = ~n4915 ;
  assign \g56841/_0_  = ~n4930 ;
  assign \g56842/_0_  = ~n4949 ;
  assign \g56843/_0_  = ~n4954 ;
  assign \g56844/_0_  = ~n4973 ;
  assign \g56845/_0_  = ~n4989 ;
  assign \g56846/_0_  = ~n4995 ;
  assign \g56863/_0_  = n4996 ;
  assign \g56897/_0_  = ~n5011 ;
  assign \g56898/_0_  = ~n5030 ;
  assign \g56899/_0_  = ~n5045 ;
  assign \g56900/_0_  = ~n5064 ;
  assign \g56901/_0_  = ~n5079 ;
  assign \g56902/_0_  = ~n5098 ;
  assign \g56903/_0_  = ~n5117 ;
  assign \g56905/_0_  = ~n5123 ;
  assign \g56921/_0_  = n5124 ;
  assign \g56956/_0_  = ~n5143 ;
  assign \g56957/_0_  = ~n5162 ;
  assign \g56958/_0_  = ~n5177 ;
  assign \g56959/_0_  = ~n5196 ;
  assign \g56960/_0_  = ~n5201 ;
  assign \g56961/_0_  = ~n5220 ;
  assign \g56962/_0_  = ~n5239 ;
  assign \g56964/_0_  = ~n5245 ;
  assign \g56980/_0_  = n5246 ;
  assign \g57015/_0_  = ~n5265 ;
  assign \g57016/_0_  = ~n5284 ;
  assign \g57017/_0_  = ~n5303 ;
  assign \g57018/_0_  = ~n5322 ;
  assign \g57019/_0_  = ~n5337 ;
  assign \g57020/_0_  = ~n5356 ;
  assign \g57021/_0_  = ~n5375 ;
  assign \g57023/_0_  = ~n5381 ;
  assign \g57040/_0_  = n5382 ;
  assign \g57074/_0_  = ~n5401 ;
  assign \g57075/_0_  = ~n5407 ;
  assign \g57076/_0_  = ~n5426 ;
  assign \g57077/_0_  = ~n5445 ;
  assign \g57078/_0_  = ~n5460 ;
  assign \g57079/_0_  = ~n5479 ;
  assign \g57080/_0_  = ~n5498 ;
  assign \g57081/_0_  = ~n5514 ;
  assign \g57099/_0_  = n5515 ;
  assign \g57133/_0_  = ~n5521 ;
  assign \g57134/_0_  = ~n5527 ;
  assign \g57135/_0_  = ~n5546 ;
  assign \g57136/_0_  = ~n5565 ;
  assign \g57137/_0_  = ~n5580 ;
  assign \g57138/_0_  = ~n5599 ;
  assign \g57139/_0_  = ~n5618 ;
  assign \g57140/_0_  = ~n5634 ;
  assign \g57141/_0_  = ~n5640 ;
  assign \g57159/_0_  = n5641 ;
  assign \g57193/_0_  = ~n5660 ;
  assign \g57195/_0_  = ~n5679 ;
  assign \g57196/_0_  = ~n5698 ;
  assign \g57197/_0_  = ~n5703 ;
  assign \g57198/_0_  = ~n5722 ;
  assign \g57199/_0_  = ~n5741 ;
  assign \g57200/_0_  = ~n5761 ;
  assign \g57202/_0_  = ~n5767 ;
  assign \g57219/_0_  = n5768 ;
  assign \g57254/_0_  = ~n5787 ;
  assign \g57255/_0_  = ~n5806 ;
  assign \g57256/_0_  = ~n5812 ;
  assign \g57257/_0_  = ~n5831 ;
  assign \g57258/_0_  = ~n5850 ;
  assign \g57259/_0_  = ~n5855 ;
  assign \g57260/_0_  = ~n5874 ;
  assign \g57262/_0_  = ~n5890 ;
  assign \g57263/_0_  = ~n5896 ;
  assign \g57285/_0_  = n5897 ;
  assign \g57318/_0_  = ~n5916 ;
  assign \g57319/_0_  = ~n5935 ;
  assign \g57320/_0_  = ~n5941 ;
  assign \g57321/_0_  = ~n5947 ;
  assign \g57322/_0_  = ~n5966 ;
  assign \g57323/_0_  = ~n5985 ;
  assign \g57324/_0_  = ~n6000 ;
  assign \g57325/_0_  = ~n6019 ;
  assign \g57326/_0_  = ~n6035 ;
  assign \g57328/_0_  = ~n6051 ;
  assign \g57329/_0_  = ~n6058 ;
  assign \g57330/_0_  = ~n6064 ;
  assign \g57350/_0_  = n6065 ;
  assign \g57387/_0_  = ~n6084 ;
  assign \g57388/_0_  = ~n6103 ;
  assign \g57390/_0_  = ~n6109 ;
  assign \g57391/_0_  = ~n6128 ;
  assign \g57392/_0_  = ~n6147 ;
  assign \g57393/_0_  = ~n6152 ;
  assign \g57395/_0_  = ~n6171 ;
  assign \g57396/_0_  = ~n6177 ;
  assign \g57439/_0_  = n6178 ;
  assign \g57476/_0_  = ~n6197 ;
  assign \g57477/_0_  = ~n6216 ;
  assign \g57478/_0_  = ~n6235 ;
  assign \g57479/_0_  = ~n6241 ;
  assign \g57480/_0_  = ~n6260 ;
  assign \g57481/_0_  = ~n6292 ;
  assign \g57482/_0_  = ~n6324 ;
  assign \g57483/_0_  = ~n6343 ;
  assign \g57484/_0_  = ~n6349 ;
  assign \g57485/_0_  = ~n6355 ;
  assign \g57486/_0_  = ~n6361 ;
  assign \g57487/_0_  = ~n6367 ;
  assign \g57488/_0_  = ~n6386 ;
  assign \g57489/_0_  = ~n6405 ;
  assign \g57490/_0_  = ~n6424 ;
  assign \g57491/_0_  = ~n6430 ;
  assign \g57492/_0_  = ~n6449 ;
  assign \g57493/_0_  = ~n6468 ;
  assign \g57494/_0_  = ~n6487 ;
  assign \g57495/_0_  = ~n6493 ;
  assign \g57496/_0_  = ~n6498 ;
  assign \g57497/_0_  = ~n6513 ;
  assign \g57498/_0_  = ~n6518 ;
  assign \g57499/_0_  = ~n6524 ;
  assign \g57500/_0_  = ~n6530 ;
  assign \g57501/_0_  = ~n6536 ;
  assign \g57502/_0_  = ~n6542 ;
  assign \g57503/_0_  = ~n6548 ;
  assign \g57504/_0_  = ~n6554 ;
  assign \g57505/_0_  = ~n6560 ;
  assign \g57524/_0_  = n6561 ;
  assign \g57537/_0_  = n6565 ;
  assign \g57541/_0_  = n6569 ;
  assign \g57543/_0_  = n6573 ;
  assign \g58163/_0_  = n6574 ;
  assign \g58572/_0_  = n6581 ;
  assign \g58573/_0_  = n6588 ;
  assign \g58574/_0_  = n6595 ;
  assign \g58575/_0_  = n6602 ;
  assign \g58576/_0_  = n6609 ;
  assign \g58577/_0_  = n6616 ;
  assign \g58578/_0_  = n6623 ;
  assign \g58579/_0_  = n6630 ;
  assign \g58580/_0_  = n6637 ;
  assign \g58581/_0_  = n6644 ;
  assign \g58582/_0_  = n6651 ;
  assign \g58583/_0_  = n6658 ;
  assign \g58584/_0_  = n6665 ;
  assign \g58585/_0_  = n6672 ;
  assign \g58586/_0_  = n6679 ;
  assign \g58587/_0_  = n6686 ;
  assign \g58588/_0_  = n6693 ;
  assign \g58589/_0_  = n6700 ;
  assign \g58590/_0_  = n6707 ;
  assign \g58591/_0_  = n6714 ;
  assign \g58592/_0_  = n6721 ;
  assign \g58593/_0_  = n6728 ;
  assign \g58594/_0_  = n6735 ;
  assign \g58595/_0_  = n6742 ;
  assign \g58596/_0_  = n6749 ;
  assign \g58597/_0_  = n6756 ;
  assign \g58598/_0_  = n6763 ;
  assign \g58600/_0_  = n6764 ;
  assign \g58602/_0_  = n6765 ;
  assign \g58604/_0_  = n6766 ;
  assign \g58615/_0_  = n6767 ;
  assign \g59240/_0_  = n6771 ;
  assign \g59241/_0_  = n6775 ;
  assign \g59242/_0_  = n6779 ;
  assign \g59243/_0_  = n6783 ;
  assign \g59244/_0_  = n6787 ;
  assign \g59245/_0_  = n6791 ;
  assign \g59246/_0_  = n6795 ;
  assign \g59247/_0_  = n6799 ;
  assign \g59248/_0_  = n6803 ;
  assign \g59249/_0_  = n6807 ;
  assign \g59250/_0_  = n6811 ;
  assign \g59251/_0_  = n6815 ;
  assign \g59252/_0_  = n6819 ;
  assign \g59253/_0_  = n6823 ;
  assign \g59254/_0_  = n6827 ;
  assign \g59255/_0_  = n6831 ;
  assign \g59256/_0_  = n6835 ;
  assign \g59257/_0_  = n6839 ;
  assign \g59258/_0_  = n6843 ;
  assign \g59259/_0_  = n6847 ;
  assign \g59260/_0_  = n6851 ;
  assign \g59261/_0_  = n6855 ;
  assign \g59262/_0_  = n6859 ;
  assign \g59263/_0_  = n6863 ;
  assign \g59264/_0_  = n6867 ;
  assign \g59265/_0_  = n6871 ;
  assign \g59266/_0_  = n6875 ;
  assign \g59267/_0_  = n6879 ;
  assign \g59268/_0_  = n6883 ;
  assign \g59269/_0_  = n6887 ;
  assign \g59270/_0_  = n6891 ;
  assign \g59271/_0_  = n6895 ;
  assign \g59272/_0_  = n6899 ;
  assign \g59273/_0_  = n6903 ;
  assign \g59274/_0_  = n6907 ;
  assign \g59275/_0_  = n6911 ;
  assign \g59276/_0_  = n6915 ;
  assign \g59277/_0_  = n6919 ;
  assign \g59278/_0_  = n6923 ;
  assign \g59279/_0_  = n6927 ;
  assign \g59280/_0_  = n6931 ;
  assign \g59281/_0_  = n6935 ;
  assign \g59282/_0_  = n6939 ;
  assign \g59283/_0_  = n6943 ;
  assign \g59284/_0_  = n6947 ;
  assign \g59285/_0_  = n6951 ;
  assign \g59286/_0_  = n6955 ;
  assign \g59287/_0_  = n6959 ;
  assign \g59288/_0_  = n6963 ;
  assign \g59289/_0_  = n6967 ;
  assign \g59290/_0_  = n6971 ;
  assign \g59291/_0_  = n6975 ;
  assign \g59292/_0_  = n6979 ;
  assign \g59293/_0_  = n6983 ;
  assign \g59294/_0_  = n6987 ;
  assign \g59295/_0_  = n6991 ;
  assign \g59296/_0_  = n6995 ;
  assign \g59297/_0_  = n6999 ;
  assign \g59298/_0_  = n7003 ;
  assign \g59299/_0_  = n7007 ;
  assign \g59300/_0_  = n7011 ;
  assign \g59301/_0_  = n7015 ;
  assign \g59302/_0_  = n7019 ;
  assign \g59303/_0_  = n7023 ;
  assign \g59304/_0_  = n7027 ;
  assign \g59305/_0_  = n7031 ;
  assign \g59306/_0_  = n7035 ;
  assign \g59307/_0_  = n7039 ;
  assign \g59308/_0_  = n7043 ;
  assign \g59309/_0_  = n7047 ;
  assign \g59310/_0_  = n7051 ;
  assign \g59311/_0_  = n7055 ;
  assign \g59312/_0_  = n7059 ;
  assign \g59313/_0_  = n7063 ;
  assign \g59314/_0_  = n7067 ;
  assign \g59315/_0_  = n7071 ;
  assign \g59316/_0_  = n7075 ;
  assign \g59317/_0_  = n7079 ;
  assign \g59318/_0_  = n7083 ;
  assign \g59319/_0_  = n7087 ;
  assign \g59320/_0_  = n7091 ;
  assign \g59321/_0_  = n7095 ;
  assign \g59322/_0_  = n7099 ;
  assign \g59323/_0_  = n7103 ;
  assign \g59324/_0_  = n7107 ;
  assign \g59325/_0_  = n7111 ;
  assign \g59326/_0_  = n7115 ;
  assign \g59327/_0_  = n7119 ;
  assign \g59328/_0_  = n7123 ;
  assign \g59329/_0_  = n7127 ;
  assign \g59330/_0_  = n7131 ;
  assign \g59331/_0_  = n7135 ;
  assign \g59332/_0_  = n7139 ;
  assign \g59333/_0_  = n7143 ;
  assign \g59334/_0_  = n7147 ;
  assign \g59335/_0_  = n7151 ;
  assign \g59336/_0_  = n7155 ;
  assign \g59337/_0_  = n7159 ;
  assign \g59338/_0_  = n7163 ;
  assign \g59339/_0_  = n7167 ;
  assign \g59340/_0_  = n7171 ;
  assign \g59341/_0_  = n7175 ;
  assign \g59342/_0_  = n7179 ;
  assign \g59343/_0_  = n7183 ;
  assign \g59344/_0_  = n7187 ;
  assign \g59345/_0_  = n7191 ;
  assign \g59346/_0_  = n7195 ;
  assign \g59347/_0_  = n7199 ;
  assign \g59348/_0_  = n7203 ;
  assign \g59349/_0_  = n7207 ;
  assign \g59350/_0_  = n7211 ;
  assign \g59351/_0_  = n7215 ;
  assign \g59352/_0_  = n7219 ;
  assign \g59353/_0_  = n7223 ;
  assign \g59354/_0_  = n7227 ;
  assign \g59355/_0_  = n7231 ;
  assign \g59356/_0_  = n7235 ;
  assign \g59357/_0_  = n7239 ;
  assign \g59358/_0_  = n7243 ;
  assign \g59359/_0_  = n7247 ;
  assign \g59360/_0_  = n7251 ;
  assign \g59361/_0_  = n7255 ;
  assign \g59362/_0_  = n7259 ;
  assign \g59363/_0_  = n7263 ;
  assign \g59364/_0_  = n7267 ;
  assign \g59365/_0_  = n7271 ;
  assign \g59366/_0_  = n7275 ;
  assign \g59367/_0_  = n7279 ;
  assign \g59368/_0_  = n7283 ;
  assign \g59369/_0_  = n7287 ;
  assign \g59370/_0_  = n7291 ;
  assign \g59371/_0_  = n7295 ;
  assign \g59372/_0_  = n7299 ;
  assign \g59373/_0_  = n7303 ;
  assign \g59374/_0_  = n7307 ;
  assign \g59375/_0_  = n7311 ;
  assign \g59376/_0_  = n7315 ;
  assign \g59377/_0_  = n7319 ;
  assign \g59378/_0_  = n7323 ;
  assign \g59379/_0_  = n7327 ;
  assign \g59380/_0_  = n7331 ;
  assign \g59381/_0_  = n7335 ;
  assign \g59382/_0_  = n7339 ;
  assign \g59383/_0_  = n7343 ;
  assign \g59384/_0_  = n7347 ;
  assign \g59385/_0_  = n7351 ;
  assign \g59386/_0_  = n7355 ;
  assign \g59387/_0_  = n7359 ;
  assign \g59388/_0_  = n7363 ;
  assign \g59389/_0_  = n7367 ;
  assign \g59390/_0_  = n7371 ;
  assign \g59391/_0_  = n7375 ;
  assign \g59392/_0_  = n7379 ;
  assign \g59393/_0_  = n7383 ;
  assign \g59394/_0_  = n7387 ;
  assign \g59395/_0_  = n7391 ;
  assign \g59396/_0_  = n7395 ;
  assign \g59397/_0_  = n7399 ;
  assign \g59398/_0_  = n7403 ;
  assign \g59399/_0_  = n7407 ;
  assign \g59400/_0_  = n7411 ;
  assign \g59401/_0_  = n7415 ;
  assign \g59402/_0_  = n7419 ;
  assign \g59403/_0_  = n7423 ;
  assign \g59404/_0_  = n7427 ;
  assign \g59405/_0_  = n7431 ;
  assign \g59406/_0_  = n7435 ;
  assign \g59407/_0_  = n7439 ;
  assign \g59408/_0_  = n7443 ;
  assign \g59409/_0_  = n7447 ;
  assign \g59410/_0_  = n7451 ;
  assign \g59411/_0_  = n7455 ;
  assign \g59412/_0_  = n7459 ;
  assign \g59413/_0_  = n7463 ;
  assign \g59414/_0_  = n7467 ;
  assign \g59415/_0_  = n7471 ;
  assign \g59416/_0_  = n7475 ;
  assign \g59417/_0_  = n7479 ;
  assign \g59418/_0_  = n7483 ;
  assign \g59419/_0_  = n7487 ;
  assign \g59420/_0_  = n7491 ;
  assign \g59421/_0_  = n7495 ;
  assign \g59422/_0_  = n7499 ;
  assign \g59423/_0_  = n7503 ;
  assign \g59424/_0_  = n7507 ;
  assign \g59425/_0_  = n7511 ;
  assign \g59426/_0_  = n7515 ;
  assign \g59427/_0_  = n7519 ;
  assign \g59428/_0_  = n7523 ;
  assign \g59429/_0_  = n7527 ;
  assign \g59430/_0_  = n7531 ;
  assign \g59431/_0_  = n7535 ;
  assign \g59432/_0_  = n7539 ;
  assign \g59433/_0_  = n7543 ;
  assign \g59434/_0_  = n7547 ;
  assign \g59435/_0_  = n7551 ;
  assign \g59436/_0_  = n7555 ;
  assign \g59437/_0_  = n7559 ;
  assign \g59438/_0_  = n7563 ;
  assign \g59439/_0_  = n7567 ;
  assign \g59440/_0_  = n7571 ;
  assign \g59441/_0_  = n7575 ;
  assign \g59442/_0_  = n7579 ;
  assign \g59443/_0_  = n7583 ;
  assign \g59444/_0_  = n7587 ;
  assign \g59445/_0_  = n7591 ;
  assign \g59446/_0_  = n7595 ;
  assign \g59447/_0_  = n7599 ;
  assign \g59448/_0_  = n7603 ;
  assign \g59449/_0_  = n7607 ;
  assign \g59450/_0_  = n7611 ;
  assign \g59451/_0_  = n7615 ;
  assign \g59452/_0_  = n7619 ;
  assign \g59453/_0_  = n7623 ;
  assign \g59454/_0_  = n7627 ;
  assign \g59455/_0_  = n7631 ;
  assign \g59456/_0_  = n7635 ;
  assign \g59457/_0_  = n7639 ;
  assign \g59458/_0_  = n7643 ;
  assign \g59459/_0_  = n7647 ;
  assign \g59460/_0_  = n7651 ;
  assign \g59461/_0_  = n7655 ;
  assign \g59462/_0_  = n7659 ;
  assign \g59463/_0_  = n7663 ;
  assign \g59464/_0_  = n7667 ;
  assign \g59465/_0_  = n7671 ;
  assign \g59466/_0_  = n7675 ;
  assign \g59467/_0_  = n7679 ;
  assign \g59468/_0_  = n7683 ;
  assign \g59469/_0_  = n7687 ;
  assign \g59470/_0_  = n7691 ;
  assign \g59471/_0_  = n7695 ;
  assign \g59472/_0_  = n7699 ;
  assign \g59473/_0_  = n7703 ;
  assign \g59474/_0_  = n7707 ;
  assign \g59475/_0_  = n7711 ;
  assign \g59476/_0_  = n7715 ;
  assign \g59477/_0_  = n7719 ;
  assign \g59478/_0_  = n7723 ;
  assign \g59479/_0_  = n7727 ;
  assign \g59480/_0_  = n7731 ;
  assign \g59481/_0_  = n7735 ;
  assign \g59482/_0_  = n7739 ;
  assign \g59483/_0_  = n7743 ;
  assign \g59484/_0_  = n7747 ;
  assign \g59485/_0_  = n7751 ;
  assign \g59486/_0_  = n7755 ;
  assign \g59487/_0_  = n7759 ;
  assign \g59488/_0_  = n7763 ;
  assign \g59489/_0_  = n7767 ;
  assign \g59490/_0_  = n7771 ;
  assign \g59491/_0_  = n7775 ;
  assign \g59492/_0_  = n7779 ;
  assign \g59493/_0_  = n7783 ;
  assign \g59494/_0_  = n7787 ;
  assign \g59495/_0_  = n7791 ;
  assign \g59496/_0_  = n7795 ;
  assign \g59497/_0_  = n7799 ;
  assign \g59498/_0_  = n7800 ;
  assign \g59500/_0_  = n7801 ;
  assign \g59503/_0_  = n7802 ;
  assign \g59512/_0_  = n7803 ;
  assign \g61336/_0_  = n7804 ;
  assign \g61521/_0_  = n7805 ;
  assign \g61523/_0_  = n7806 ;
  assign \g61524/_0_  = n7807 ;
  assign \g61526/_0_  = n7808 ;
  assign \g61527/_0_  = n7809 ;
  assign \g61528/_0_  = n7810 ;
  assign \g61529/_0_  = n7811 ;
  assign \g61530/_0_  = n7812 ;
  assign \g61531/_0_  = n7813 ;
  assign \g61532/_0_  = n7814 ;
  assign \g61533/_0_  = n7815 ;
  assign \g61535/_0_  = n7816 ;
  assign \g61537/_0_  = n7817 ;
  assign \g61539/_0_  = n7818 ;
  assign \g61540/_0_  = n7819 ;
  assign \g61541/_0_  = n7820 ;
  assign \g61542/_0_  = n7821 ;
  assign \g61546/_0_  = n7822 ;
  assign \g61550/_0_  = n7823 ;
  assign \g61551/_0_  = n7824 ;
  assign \g61552/_0_  = n7825 ;
  assign \g61554/_0_  = n7826 ;
  assign \g61555/_0_  = n7827 ;
  assign \g61556/_0_  = n7828 ;
  assign \g61558/_0_  = n7829 ;
  assign \g61559/_0_  = n7830 ;
  assign \g61561/_0_  = n7831 ;
  assign \g61562/_0_  = n7832 ;
  assign \g61563/_0_  = n7833 ;
  assign \g61564/_0_  = n7834 ;
  assign \g61565/_0_  = n7835 ;
  assign \g61566/_0_  = n7836 ;
  assign \g61568/_0_  = n7837 ;
  assign \g61570/_0_  = n7838 ;
  assign \g61571/_0_  = n7839 ;
  assign \g61572/_0_  = n7840 ;
  assign \g61573/_0_  = n7841 ;
  assign \g61577/_0_  = n7842 ;
  assign \g61578/_0_  = n7843 ;
  assign \g61579/_0_  = n7844 ;
  assign \g61580/_0_  = n7845 ;
  assign \g61581/_0_  = n7846 ;
  assign \g61582/_0_  = n7847 ;
  assign \g61583/_0_  = n7848 ;
  assign \g61584/_0_  = n7849 ;
  assign \g61585/_0_  = n7850 ;
  assign \g61586/_0_  = n7851 ;
  assign \g61587/_0_  = n7852 ;
  assign \g61588/_0_  = n7853 ;
  assign \g61589/_0_  = n7854 ;
  assign \g61591/_0_  = n7855 ;
  assign \g61592/_0_  = n7856 ;
  assign \g61594/_0_  = n7857 ;
  assign \g61595/_0_  = n7858 ;
  assign \g61596/_0_  = n7859 ;
  assign \g61597/_0_  = n7860 ;
  assign \g61598/_0_  = n7861 ;
  assign \g61599/_0_  = n7862 ;
  assign \g61600/_0_  = n7863 ;
  assign \g61601/_0_  = n7864 ;
  assign \g61605/_0_  = n7865 ;
  assign \g61606/_0_  = n7866 ;
  assign \g61607/_0_  = n7867 ;
  assign \g61608/_0_  = n7868 ;
  assign \g61609/_0_  = n7869 ;
  assign \g61610/_0_  = n7870 ;
  assign \g61611/_0_  = n7871 ;
  assign \g61612/_0_  = n7872 ;
  assign \g61613/_0_  = n7873 ;
  assign \g61615/_0_  = n7874 ;
  assign \g61616/_0_  = n7875 ;
  assign \g61617/_0_  = n7876 ;
  assign \g61618/_0_  = n7877 ;
  assign \g61619/_0_  = n7878 ;
  assign \g61620/_0_  = n7879 ;
  assign \g61621/_0_  = n7880 ;
  assign \g61623/_0_  = n7881 ;
  assign \g61624/_0_  = n7882 ;
  assign \g61625/_0_  = n7883 ;
  assign \g61626/_0_  = n7884 ;
  assign \g61627/_0_  = n7885 ;
  assign \g61629/_0_  = n7886 ;
  assign \g61630/_0_  = n7887 ;
  assign \g61631/_0_  = n7888 ;
  assign \g61632/_0_  = n7889 ;
  assign \g61633/_0_  = n7890 ;
  assign \g61634/_0_  = n7891 ;
  assign \g61636/_0_  = n7892 ;
  assign \g61638/_0_  = n7893 ;
  assign \g61639/_0_  = n7894 ;
  assign \g61640/_0_  = n7895 ;
  assign \g61641/_0_  = n7896 ;
  assign \g61642/_0_  = n7897 ;
  assign \g61644/_0_  = n7898 ;
  assign \g61647/_0_  = n7899 ;
  assign \g61648/_0_  = n7900 ;
  assign \g61649/_0_  = n7901 ;
  assign \g61650/_0_  = n7902 ;
  assign \g61653/_0_  = n7903 ;
  assign \g61654/_0_  = n7904 ;
  assign \g61655/_0_  = n7905 ;
  assign \g61656/_0_  = n7906 ;
  assign \g61658/_0_  = n7907 ;
  assign \g61661/_0_  = n7908 ;
  assign \g61662/_0_  = n7909 ;
  assign \g61663/_0_  = n7910 ;
  assign \g61664/_0_  = n7911 ;
  assign \g61666/_0_  = n7912 ;
  assign \g61667/_0_  = n7913 ;
  assign \g61668/_0_  = n7914 ;
  assign \g61670/_0_  = n7915 ;
  assign \g61671/_0_  = n7916 ;
  assign \g61672/_0_  = n7917 ;
  assign \g61673/_0_  = n7918 ;
  assign \g61675/_0_  = n7919 ;
  assign \g61676/_0_  = n7920 ;
  assign \g61680/_0_  = n7921 ;
  assign \g61681/_0_  = n7922 ;
  assign \g61682/_0_  = n7923 ;
  assign \g61683/_0_  = n7924 ;
  assign \g61684/_0_  = n7925 ;
  assign \g61686/_0_  = n7926 ;
  assign \g61687/_0_  = n7927 ;
  assign \g61688/_0_  = n7928 ;
  assign \g61689/_0_  = n7929 ;
  assign \g61690/_0_  = n7930 ;
  assign \g61691/_0_  = n7931 ;
  assign \g61693/_0_  = n7932 ;
  assign \g61694/_0_  = n7933 ;
  assign \g61696/_0_  = n7934 ;
  assign \g61697/_0_  = n7935 ;
  assign \g61698/_0_  = n7936 ;
  assign \g61699/_0_  = n7937 ;
  assign \g61700/_0_  = n7938 ;
  assign \g61701/_0_  = n7939 ;
  assign \g61702/_0_  = n7940 ;
  assign \g61703/_0_  = n7941 ;
  assign \g61704/_0_  = n7942 ;
  assign \g61705/_0_  = n7943 ;
  assign \g61706/_0_  = n7944 ;
  assign \g61707/_0_  = n7945 ;
  assign \g61708/_0_  = n7946 ;
  assign \g61711/_0_  = n7947 ;
  assign \g61712/_0_  = n7948 ;
  assign \g61714/_0_  = n7949 ;
  assign \g61716/_0_  = n7950 ;
  assign \g61717/_0_  = n7951 ;
  assign \g61719/_0_  = n7952 ;
  assign \g61720/_0_  = n7953 ;
  assign \g61721/_0_  = n7954 ;
  assign \g61724/_0_  = n7955 ;
  assign \g61725/_0_  = n7956 ;
  assign \g61728/_0_  = n7957 ;
  assign \g61729/_0_  = n7958 ;
  assign \g61731/_0_  = n7959 ;
  assign \g61732/_0_  = n7960 ;
  assign \g61733/_0_  = n7961 ;
  assign \g61736/_0_  = n7962 ;
  assign \g61737/_0_  = n7963 ;
  assign \g61739/_0_  = n7964 ;
  assign \g61740/_0_  = n7965 ;
  assign \g61741/_0_  = n7966 ;
  assign \g61743/_0_  = n7967 ;
  assign \g61744/_0_  = n7968 ;
  assign \g61745/_0_  = n7969 ;
  assign \g61746/_0_  = n7970 ;
  assign \g61747/_0_  = n7971 ;
  assign \g61748/_0_  = n7972 ;
  assign \g61749/_0_  = n7973 ;
  assign \g61750/_0_  = n7974 ;
  assign \g61751/_0_  = n7975 ;
  assign \g61752/_0_  = n7976 ;
  assign \g61753/_0_  = n7977 ;
  assign \g61754/_0_  = n7978 ;
  assign \g61755/_0_  = n7979 ;
  assign \g61757/_0_  = n7980 ;
  assign \g61758/_0_  = n7981 ;
  assign \g61759/_0_  = n7982 ;
  assign \g61760/_0_  = n7983 ;
  assign \g61761/_0_  = n7984 ;
  assign \g61762/_0_  = n7985 ;
  assign \g61763/_0_  = n7986 ;
  assign \g61764/_0_  = n7987 ;
  assign \g61765/_0_  = n7988 ;
  assign \g61766/_0_  = n7989 ;
  assign \g61767/_0_  = n7990 ;
  assign \g61768/_0_  = n7991 ;
  assign \g61769/_0_  = n7992 ;
  assign \g61770/_0_  = n7993 ;
  assign \g61771/_0_  = n7994 ;
  assign \g61772/_0_  = n7995 ;
  assign \g61773/_0_  = n7996 ;
  assign \g61774/_0_  = n7997 ;
  assign \g61775/_0_  = n7998 ;
  assign \g61776/_0_  = n7999 ;
  assign \g61777/_0_  = n8000 ;
  assign \g61778/_0_  = n8001 ;
  assign \g61780/_0_  = n8002 ;
  assign \g61781/_0_  = n8003 ;
  assign \g61783/_0_  = n8004 ;
  assign \g61784/_0_  = n8005 ;
  assign \g61786/_0_  = n8006 ;
  assign \g61787/_0_  = n8007 ;
  assign \g61790/_0_  = n8008 ;
  assign \g61791/_0_  = n8009 ;
  assign \g61794/_0_  = n8010 ;
  assign \g61795/_0_  = n8011 ;
  assign \g61796/_0_  = n8012 ;
  assign \g61797/_0_  = n8013 ;
  assign \g61798/_0_  = n8014 ;
  assign \g61799/_0_  = n8015 ;
  assign \g61800/_0_  = n8016 ;
  assign \g61801/_0_  = n8017 ;
  assign \g61802/_0_  = n8018 ;
  assign \g61803/_0_  = n8019 ;
  assign \g61805/_0_  = n8020 ;
  assign \g61806/_0_  = n8021 ;
  assign \g61807/_0_  = n8022 ;
  assign \g61808/_0_  = n8023 ;
  assign \g61809/_0_  = n8024 ;
  assign \g61810/_0_  = n8025 ;
  assign \g61811/_0_  = n8026 ;
  assign \g61812/_0_  = n8027 ;
  assign \g61813/_0_  = n8028 ;
  assign \g61816/_0_  = n8029 ;
  assign \g61817/_0_  = n8030 ;
  assign \g61818/_0_  = n8031 ;
  assign \g61820/_0_  = n8032 ;
  assign \g61822/_0_  = n8033 ;
  assign \g61823/_0_  = n8034 ;
  assign \g61825/_0_  = n8035 ;
  assign \g61826/_0_  = n8036 ;
  assign \g61827/_0_  = n8037 ;
  assign \g61828/_0_  = n8038 ;
  assign \g61829/_0_  = n8039 ;
  assign \g61832/_0_  = n8040 ;
  assign \g61834/_0_  = n8041 ;
  assign \g61835/_0_  = n8042 ;
  assign \g61837/_0_  = n8043 ;
  assign \g61838/_0_  = n8044 ;
  assign \g61839/_0_  = n8045 ;
  assign \g61840/_0_  = n8046 ;
  assign \g61844/_0_  = n8047 ;
  assign \g61847/_0_  = n8048 ;
  assign \g61848/_0_  = n8049 ;
  assign \g61849/_0_  = n8050 ;
  assign \g61850/_0_  = n8051 ;
  assign \g61851/_0_  = n8052 ;
  assign \g61853/_0_  = n8053 ;
  assign \g61854/_0_  = n8054 ;
  assign \g61855/_0_  = n8055 ;
  assign \g61856/_0_  = n8056 ;
  assign \g61858/_0_  = n8057 ;
  assign \g61859/_0_  = n8058 ;
  assign \g61861/_0_  = n8059 ;
  assign \g61862/_0_  = n8060 ;
  assign \g61863/_0_  = n8061 ;
  assign \g61864/_0_  = n8062 ;
  assign \g61865/_0_  = n8063 ;
  assign \g61866/_0_  = n8064 ;
  assign \g61867/_0_  = n8065 ;
  assign \g61868/_0_  = n8066 ;
  assign \g61869/_0_  = n8067 ;
  assign \g61870/_0_  = n8068 ;
  assign \g61871/_0_  = n8069 ;
  assign \g61873/_0_  = n8070 ;
  assign \g61874/_0_  = n8071 ;
  assign \g61875/_0_  = n8072 ;
  assign \g61877/_0_  = n8073 ;
  assign \g61878/_0_  = n8074 ;
  assign \g61879/_0_  = n8075 ;
  assign \g61880/_0_  = n8076 ;
  assign \g61881/_0_  = n8077 ;
  assign \g61883/_0_  = n8078 ;
  assign \g61884/_0_  = n8079 ;
  assign \g61886/_0_  = n8080 ;
  assign \g61887/_0_  = n8081 ;
  assign \g61890/_0_  = n8082 ;
  assign \g61891/_0_  = n8083 ;
  assign \g61892/_0_  = n8084 ;
  assign \g61893/_0_  = n8085 ;
  assign \g61894/_0_  = n8086 ;
  assign \g61895/_0_  = n8087 ;
  assign \g61900/_0_  = n8088 ;
  assign \g61901/_0_  = n8089 ;
  assign \g61902/_0_  = n8090 ;
  assign \g61904/_0_  = n8091 ;
  assign \g61905/_0_  = n8092 ;
  assign \g61906/_0_  = n8093 ;
  assign \g61907/_0_  = n8094 ;
  assign \g61914/_0_  = n8095 ;
  assign \g61915/_0_  = n8096 ;
  assign \g61917/_0_  = n8097 ;
  assign \g61919/_0_  = n8098 ;
  assign \g61921/_0_  = n8099 ;
  assign \g61924/_0_  = n8100 ;
  assign \g61925/_0_  = n8101 ;
  assign \g61926/_0_  = n8102 ;
  assign \g61927/_0_  = n8103 ;
  assign \g61928/_0_  = n8104 ;
  assign \g61929/_0_  = n8105 ;
  assign \g61930/_0_  = n8106 ;
  assign \g61931/_0_  = n8107 ;
  assign \g61932/_0_  = n8108 ;
  assign \g61933/_0_  = n8109 ;
  assign \g61934/_0_  = n8110 ;
  assign \g61935/_0_  = n8111 ;
  assign \g61936/_0_  = n8112 ;
  assign \g61937/_0_  = n8113 ;
  assign \g61938/_0_  = n8114 ;
  assign \g61939/_0_  = n8115 ;
  assign \g61943/_0_  = n8116 ;
  assign \g61944/_0_  = n8117 ;
  assign \g61945/_0_  = n8118 ;
  assign \g61947/_0_  = n8119 ;
  assign \g61948/_0_  = n8120 ;
  assign \g61949/_0_  = n8121 ;
  assign \g61950/_0_  = n8122 ;
  assign \g61951/_0_  = n8123 ;
  assign \g61952/_0_  = n8124 ;
  assign \g61953/_0_  = n8125 ;
  assign \g61955/_0_  = n8126 ;
  assign \g61956/_0_  = n8127 ;
  assign \g61957/_0_  = n8128 ;
  assign \g61958/_0_  = n8129 ;
  assign \g61959/_0_  = n8130 ;
  assign \g61960/_0_  = n8131 ;
  assign \g61961/_0_  = n8132 ;
  assign \g61962/_0_  = n8133 ;
  assign \g61963/_0_  = n8134 ;
  assign \g61964/_0_  = n8135 ;
  assign \g61965/_0_  = n8136 ;
  assign \g61966/_0_  = n8137 ;
  assign \g61967/_0_  = n8138 ;
  assign \g61968/_0_  = n8139 ;
  assign \g61969/_0_  = n8140 ;
  assign \g61970/_0_  = n8141 ;
  assign \g61971/_0_  = n8142 ;
  assign \g61972/_0_  = n8143 ;
  assign \g61973/_0_  = n8144 ;
  assign \g61974/_0_  = n8145 ;
  assign \g61976/_0_  = n8146 ;
  assign \g61978/_0_  = n8147 ;
  assign \g61980/_0_  = n8148 ;
  assign \g61981/_0_  = n8149 ;
  assign \g61982/_0_  = n8150 ;
  assign \g61983/_0_  = n8151 ;
  assign \g61984/_0_  = n8152 ;
  assign \g61985/_0_  = n8153 ;
  assign \g61986/_0_  = n8154 ;
  assign \g61987/_0_  = n8155 ;
  assign \g61988/_0_  = n8156 ;
  assign \g61989/_0_  = n8157 ;
  assign \g61990/_0_  = n8158 ;
  assign \g61992/_0_  = n8159 ;
  assign \g61994/_0_  = n8160 ;
  assign \g61995/_0_  = n8161 ;
  assign \g61996/_0_  = n8162 ;
  assign \g61997/_0_  = n8163 ;
  assign \g61998/_0_  = n8164 ;
  assign \g62000/_0_  = n8165 ;
  assign \g62001/_0_  = n8166 ;
  assign \g62002/_0_  = n8167 ;
  assign \g62003/_0_  = n8168 ;
  assign \g62004/_0_  = n8169 ;
  assign \g62005/_0_  = n8170 ;
  assign \g62007/_0_  = n8171 ;
  assign \g62008/_0_  = n8172 ;
  assign \g62009/_0_  = n8173 ;
  assign \g62010/_0_  = n8174 ;
  assign \g62011/_0_  = n8175 ;
  assign \g62012/_0_  = n8176 ;
  assign \g62013/_0_  = n8177 ;
  assign \g62014/_0_  = n8178 ;
  assign \g62015/_0_  = n8179 ;
  assign \g62016/_0_  = n8180 ;
  assign \g62017/_0_  = n8181 ;
  assign \g62018/_0_  = n8182 ;
  assign \g62019/_0_  = n8183 ;
  assign \g62020/_0_  = n8184 ;
  assign \g62021/_0_  = n8185 ;
  assign \g62022/_0_  = n8186 ;
  assign \g62023/_0_  = n8187 ;
  assign \g62024/_0_  = n8188 ;
  assign \g62025/_0_  = n8189 ;
  assign \g62026/_0_  = n8190 ;
  assign \g62027/_0_  = n8191 ;
  assign \g62030/_0_  = n8192 ;
  assign \g62033/_0_  = n8193 ;
  assign \g62034/_0_  = n8194 ;
  assign \g62036/_0_  = n8195 ;
  assign \g62038/_0_  = n8196 ;
  assign \g62041/_0_  = n8197 ;
  assign \g62042/_0_  = n8198 ;
  assign \g62043/_0_  = n8199 ;
  assign \g62044/_0_  = n8200 ;
  assign \g62045/_0_  = n8201 ;
  assign \g62046/_0_  = n8202 ;
  assign \g62047/_0_  = n8203 ;
  assign \g62048/_0_  = n8204 ;
  assign \g62050/_0_  = n8205 ;
  assign \g62051/_0_  = n8206 ;
  assign \g62052/_0_  = n8207 ;
  assign \g62055/_0_  = n8208 ;
  assign \g62057/_0_  = n8209 ;
  assign \g62058/_0_  = n8210 ;
  assign \g62059/_0_  = n8211 ;
  assign \g62060/_0_  = n8212 ;
  assign \g62061/_0_  = n8213 ;
  assign \g62062/_0_  = n8214 ;
  assign \g62064/_0_  = n8215 ;
  assign \g62065/_0_  = n8216 ;
  assign \g62066/_0_  = n8217 ;
  assign \g62067/_0_  = n8218 ;
  assign \g62068/_0_  = n8219 ;
  assign \g62072/_0_  = n8220 ;
  assign \g62073/_0_  = n8221 ;
  assign \g62074/_0_  = n8222 ;
  assign \g62075/_0_  = n8223 ;
  assign \g62076/_0_  = n8224 ;
  assign \g62077/_0_  = n8225 ;
  assign \g62078/_0_  = n8226 ;
  assign \g62080/_0_  = n8227 ;
  assign \g62081/_0_  = n8228 ;
  assign \g62082/_0_  = n8229 ;
  assign \g62084/_0_  = n8230 ;
  assign \g62085/_0_  = n8231 ;
  assign \g62086/_0_  = n8232 ;
  assign \g62087/_0_  = n8233 ;
  assign \g62088/_0_  = n8234 ;
  assign \g62089/_0_  = n8235 ;
  assign \g62090/_0_  = n8236 ;
  assign \g62091/_0_  = n8237 ;
  assign \g62092/_0_  = n8238 ;
  assign \g62094/_0_  = n8239 ;
  assign \g62096/_0_  = n8240 ;
  assign \g62097/_0_  = n8241 ;
  assign \g62098/_0_  = n8242 ;
  assign \g62099/_0_  = n8243 ;
  assign \g62100/_0_  = n8244 ;
  assign \g62101/_0_  = n8245 ;
  assign \g62102/_0_  = n8246 ;
  assign \g62104/_0_  = n8247 ;
  assign \g62106/_0_  = n8248 ;
  assign \g62107/_0_  = n8249 ;
  assign \g62108/_0_  = n8250 ;
  assign \g62110/_0_  = n8251 ;
  assign \g62112/_0_  = n8252 ;
  assign \g62113/_0_  = n8253 ;
  assign \g62114/_0_  = n8254 ;
  assign \g62116/_0_  = n8255 ;
  assign \g62117/_0_  = n8256 ;
  assign \g62118/_0_  = n8257 ;
  assign \g62119/_0_  = n8258 ;
  assign \g62120/_0_  = n8259 ;
  assign \g62121/_0_  = n8260 ;
  assign \g62122/_0_  = n8261 ;
  assign \g62124/_0_  = n8262 ;
  assign \g62126/_0_  = n8263 ;
  assign \g62127/_0_  = n8264 ;
  assign \g62128/_0_  = n8265 ;
  assign \g62129/_0_  = n8266 ;
  assign \g62130/_0_  = n8267 ;
  assign \g62131/_0_  = n8268 ;
  assign \g62132/_0_  = n8269 ;
  assign \g62133/_0_  = n8270 ;
  assign \g62135/_0_  = n8271 ;
  assign \g62136/_0_  = n8272 ;
  assign \g62137/_0_  = n8273 ;
  assign \g62138/_0_  = n8274 ;
  assign \g62140/_0_  = n8275 ;
  assign \g62143/_0_  = n8276 ;
  assign \g62144/_0_  = n8277 ;
  assign \g62149/_0_  = n8278 ;
  assign \g62150/_0_  = n8279 ;
  assign \g62151/_0_  = n8280 ;
  assign \g62153/_0_  = n8281 ;
  assign \g62155/_0_  = n8282 ;
  assign \g62156/_0_  = n8283 ;
  assign \g62158/_0_  = n8284 ;
  assign \g62160/_0_  = n8285 ;
  assign \g62161/_0_  = n8286 ;
  assign \g62162/_0_  = n8287 ;
  assign \g62164/_0_  = n8288 ;
  assign \g62165/_0_  = n8289 ;
  assign \g62166/_0_  = n8290 ;
  assign \g62167/_0_  = n8291 ;
  assign \g62168/_0_  = n8292 ;
  assign \g62169/_0_  = n8293 ;
  assign \g62172/_0_  = n8294 ;
  assign \g62173/_0_  = n8295 ;
  assign \g62175/_0_  = n8296 ;
  assign \g62176/_0_  = n8297 ;
  assign \g62177/_0_  = n8298 ;
  assign \g62178/_0_  = n8299 ;
  assign \g62179/_0_  = n8300 ;
  assign \g62180/_0_  = n8301 ;
  assign \g62181/_0_  = n8302 ;
  assign \g62182/_0_  = n8303 ;
  assign \g62183/_0_  = n8304 ;
  assign \g62184/_0_  = n8305 ;
  assign \g62185/_0_  = n8306 ;
  assign \g62186/_0_  = n8307 ;
  assign \g62188/_0_  = n8308 ;
  assign \g62189/_0_  = n8309 ;
  assign \g62190/_0_  = n8310 ;
  assign \g62191/_0_  = n8311 ;
  assign \g62193/_0_  = n8312 ;
  assign \g62194/_0_  = n8313 ;
  assign \g62195/_0_  = n8314 ;
  assign \g62196/_0_  = n8315 ;
  assign \g62197/_0_  = n8316 ;
  assign \g62200/_0_  = n8317 ;
  assign \g62201/_0_  = n8318 ;
  assign \g62202/_0_  = n8319 ;
  assign \g62203/_0_  = n8320 ;
  assign \g62205/_0_  = n8321 ;
  assign \g62206/_0_  = n8322 ;
  assign \g62207/_0_  = n8323 ;
  assign \g62208/_0_  = n8324 ;
  assign \g62209/_0_  = n8325 ;
  assign \g62210/_0_  = n8326 ;
  assign \g62211/_0_  = n8327 ;
  assign \g62215/_0_  = n8328 ;
  assign \g62218/_0_  = n8329 ;
  assign \g62219/_0_  = n8330 ;
  assign \g62221/_0_  = n8331 ;
  assign \g62222/_0_  = n8332 ;
  assign \g62223/_0_  = n8333 ;
  assign \g62224/_0_  = n8334 ;
  assign \g62225/_0_  = n8335 ;
  assign \g62226/_0_  = n8336 ;
  assign \g62229/_0_  = n8337 ;
  assign \g62230/_0_  = n8338 ;
  assign \g62231/_0_  = n8339 ;
  assign \g62233/_0_  = n8340 ;
  assign \g62236/_0_  = n8341 ;
  assign \g62237/_0_  = n8342 ;
  assign \g62238/_0_  = n8343 ;
  assign \g62240/_0_  = n8344 ;
  assign \g62241/_0_  = n8345 ;
  assign \g62243/_0_  = n8346 ;
  assign \g62244/_0_  = n8347 ;
  assign \g62245/_0_  = n8348 ;
  assign \g62247/_0_  = n8349 ;
  assign \g62248/_0_  = n8350 ;
  assign \g62250/_0_  = n8351 ;
  assign \g62252/_0_  = n8352 ;
  assign \g62253/_0_  = n8353 ;
  assign \g62255/_0_  = n8354 ;
  assign \g62256/_0_  = n8355 ;
  assign \g62257/_0_  = n8356 ;
  assign \g62258/_0_  = n8357 ;
  assign \g62259/_0_  = n8358 ;
  assign \g62260/_0_  = n8359 ;
  assign \g62261/_0_  = n8360 ;
  assign \g62262/_0_  = n8361 ;
  assign \g62263/_0_  = n8362 ;
  assign \g62264/_0_  = n8363 ;
  assign \g62265/_0_  = n8364 ;
  assign \g62267/_0_  = n8365 ;
  assign \g62269/_0_  = n8366 ;
  assign \g62270/_0_  = n8367 ;
  assign \g62272/_0_  = n8368 ;
  assign \g62274/_0_  = n8369 ;
  assign \g62277/_0_  = n8370 ;
  assign \g62279/_0_  = n8371 ;
  assign \g62280/_0_  = n8372 ;
  assign \g62281/_0_  = n8373 ;
  assign \g62283/_0_  = n8374 ;
  assign \g62284/_0_  = n8375 ;
  assign \g62285/_0_  = n8376 ;
  assign \g62286/_0_  = n8377 ;
  assign \g62288/_0_  = n8378 ;
  assign \g62289/_0_  = n8379 ;
  assign \g62290/_0_  = n8380 ;
  assign \g62294/_0_  = n8381 ;
  assign \g62295/_0_  = n8382 ;
  assign \g62296/_0_  = n8383 ;
  assign \g62297/_0_  = n8384 ;
  assign \g62298/_0_  = n8385 ;
  assign \g62299/_0_  = n8386 ;
  assign \g62303/_0_  = n8387 ;
  assign \g62305/_0_  = n8388 ;
  assign \g62306/_0_  = n8389 ;
  assign \g62307/_0_  = n8390 ;
  assign \g62309/_0_  = n8391 ;
  assign \g62311/_0_  = n8392 ;
  assign \g62312/_0_  = n8393 ;
  assign \g62313/_0_  = n8394 ;
  assign \g62314/_0_  = n8395 ;
  assign \g62315/_0_  = n8396 ;
  assign \g62316/_0_  = n8397 ;
  assign \g62317/_0_  = n8398 ;
  assign \g62318/_0_  = n8399 ;
  assign \g62319/_0_  = n8400 ;
  assign \g62320/_0_  = n8401 ;
  assign \g62322/_0_  = n8402 ;
  assign \g62324/_0_  = n8403 ;
  assign \g62325/_0_  = n8404 ;
  assign \g62326/_0_  = n8405 ;
  assign \g62327/_0_  = n8406 ;
  assign \g62329/_0_  = n8407 ;
  assign \g62330/_0_  = n8408 ;
  assign \g62331/_0_  = n8409 ;
  assign \g62332/_0_  = n8410 ;
  assign \g62333/_0_  = n8411 ;
  assign \g62335/_0_  = n8412 ;
  assign \g62336/_0_  = n8413 ;
  assign \g62338/_0_  = n8414 ;
  assign \g62341/_0_  = n8415 ;
  assign \g62342/_0_  = n8416 ;
  assign \g62344/_0_  = n8417 ;
  assign \g62345/_0_  = n8418 ;
  assign \g62348/_0_  = n8419 ;
  assign \g62349/_0_  = n8420 ;
  assign \g62350/_0_  = n8421 ;
  assign \g62353/_0_  = n8422 ;
  assign \g62354/_0_  = n8423 ;
  assign \g62355/_0_  = n8424 ;
  assign \g62356/_0_  = n8425 ;
  assign \g62359/_0_  = n8426 ;
  assign \g62362/_0_  = n8427 ;
  assign \g62363/_0_  = n8428 ;
  assign \g62364/_0_  = n8429 ;
  assign \g62365/_0_  = n8430 ;
  assign \g62366/_0_  = n8431 ;
  assign \g62367/_0_  = n8432 ;
  assign \g62368/_0_  = n8433 ;
  assign \g62369/_0_  = n8434 ;
  assign \g62370/_0_  = n8435 ;
  assign \g62371/_0_  = n8436 ;
  assign \g62372/_0_  = n8437 ;
  assign \g62373/_0_  = n8438 ;
  assign \g62374/_0_  = n8439 ;
  assign \g62376/_0_  = n8440 ;
  assign \g62467/_0_  = n8441 ;
  assign \g62468/_0_  = n8442 ;
  assign \g62469/_0_  = n8443 ;
  assign \g62470/_0_  = n8444 ;
  assign \g62471/_0_  = n8445 ;
  assign \g62472/_0_  = n8446 ;
  assign \g62473/_0_  = n8447 ;
  assign \g62474/_0_  = n8448 ;
  assign \g62475/_0_  = n8449 ;
  assign \g62478/_0_  = n8450 ;
  assign \g62480/_0_  = n8451 ;
  assign \g62481/_0_  = n8452 ;
  assign \g62482/_0_  = n8453 ;
  assign \g62483/_0_  = n8454 ;
  assign \g62484/_0_  = n8455 ;
  assign \g62485/_0_  = n8456 ;
  assign \g62486/_0_  = n8457 ;
  assign \g62487/_0_  = n8458 ;
  assign \g62488/_0_  = n8459 ;
  assign \g62489/_0_  = n8460 ;
  assign \g62490/_0_  = n8461 ;
  assign \g62491/_0_  = n8462 ;
  assign \g62492/_0_  = n8463 ;
  assign \g62493/_0_  = n8464 ;
  assign \g62494/_0_  = n8465 ;
  assign \g62495/_0_  = n8466 ;
  assign \g62496/_0_  = n8467 ;
  assign \g62497/_0_  = n8468 ;
  assign \g62498/_0_  = n8469 ;
  assign \g62499/_0_  = n8470 ;
  assign \g62500/_0_  = n8471 ;
  assign \g62501/_0_  = n8472 ;
  assign \g62502/_0_  = n8473 ;
  assign \g62503/_0_  = n8474 ;
  assign \g62504/_0_  = n8475 ;
  assign \g62509/_0_  = n8476 ;
  assign \g62510/_0_  = n8477 ;
  assign \g62511/_0_  = n8478 ;
  assign \g62512/_0_  = n8479 ;
  assign \g62513/_0_  = n8480 ;
  assign \g62514/_0_  = n8481 ;
  assign \g62515/_0_  = n8482 ;
  assign \g62516/_0_  = n8483 ;
  assign \g62517/_0_  = n8484 ;
  assign \g62518/_0_  = n8485 ;
  assign \g62519/_0_  = n8486 ;
  assign \g62520/_0_  = n8487 ;
  assign \g62521/_0_  = n8488 ;
  assign \g62523/_0_  = n8489 ;
  assign \g62526/_0_  = n8490 ;
  assign \g62528/_0_  = n8491 ;
  assign \g62529/_0_  = n8492 ;
  assign \g62531/_0_  = n8493 ;
  assign \g62532/_0_  = n8494 ;
  assign \g62533/_0_  = n8495 ;
  assign \g62534/_0_  = n8496 ;
  assign \g62535/_0_  = n8497 ;
  assign \g62536/_0_  = n8498 ;
  assign \g62537/_0_  = n8499 ;
  assign \g62539/_0_  = n8500 ;
  assign \g62540/_0_  = n8501 ;
  assign \g62541/_0_  = n8502 ;
  assign \g62542/_0_  = n8503 ;
  assign \g62543/_0_  = n8504 ;
  assign \g62544/_0_  = n8505 ;
  assign \g62545/_0_  = n8506 ;
  assign \g62547/_0_  = n8507 ;
  assign \g62548/_0_  = n8508 ;
  assign \g62549/_0_  = n8509 ;
  assign \g62550/_0_  = n8510 ;
  assign \g62551/_0_  = n8511 ;
  assign \g62552/_0_  = n8512 ;
  assign \g62553/_0_  = n8513 ;
  assign \g62554/_0_  = n8514 ;
  assign \g62555/_0_  = n8515 ;
  assign \g62556/_0_  = n8516 ;
  assign \g62557/_0_  = n8517 ;
  assign \g62560/_0_  = n8518 ;
  assign \g62562/_0_  = n8519 ;
  assign \g62563/_0_  = n8520 ;
  assign \g62564/_0_  = n8521 ;
  assign \g62565/_0_  = n8522 ;
  assign \g62566/_0_  = n8523 ;
  assign \g62567/_0_  = n8524 ;
  assign \g62569/_0_  = n8525 ;
  assign \g62570/_0_  = n8526 ;
  assign \g62571/_0_  = n8527 ;
  assign \g62572/_0_  = n8528 ;
  assign \g62573/_0_  = n8529 ;
  assign \g62574/_0_  = n8530 ;
  assign \g62576/_0_  = n8531 ;
  assign \g62577/_0_  = n8532 ;
  assign \g62581/_0_  = n8533 ;
  assign \g62582/_0_  = n8534 ;
  assign \g62584/_0_  = n8535 ;
  assign \g62585/_0_  = n8536 ;
  assign \g62586/_0_  = n8537 ;
  assign \g62588/_0_  = n8538 ;
  assign \g62589/_0_  = n8539 ;
  assign \g62593/_0_  = n8540 ;
  assign \g62594/_0_  = n8541 ;
  assign \g62595/_0_  = n8542 ;
  assign \g62596/_0_  = n8543 ;
  assign \g62597/_0_  = n8544 ;
  assign \g62598/_0_  = n8545 ;
  assign \g62599/_0_  = n8546 ;
  assign \g62600/_0_  = n8547 ;
  assign \g62601/_0_  = n8548 ;
  assign \g62602/_0_  = n8549 ;
  assign \g62603/_0_  = n8550 ;
  assign \g62604/_0_  = n8551 ;
  assign \g62605/_0_  = n8552 ;
  assign \g62606/_0_  = n8553 ;
  assign \g62607/_0_  = n8554 ;
  assign \g62608/_0_  = n8555 ;
  assign \g62609/_0_  = n8556 ;
  assign \g62610/_0_  = n8557 ;
  assign \g62612/_0_  = n8558 ;
  assign \g62613/_0_  = n8559 ;
  assign \g62614/_0_  = n8560 ;
  assign \g62615/_0_  = n8561 ;
  assign \g62617/_0_  = n8562 ;
  assign \g62618/_0_  = n8563 ;
  assign \g62620/_0_  = n8564 ;
  assign \g62621/_0_  = n8565 ;
  assign \g62622/_0_  = n8566 ;
  assign \g62624/_0_  = n8567 ;
  assign \g62625/_0_  = n8568 ;
  assign \g62626/_0_  = n8569 ;
  assign \g62627/_0_  = n8570 ;
  assign \g62629/_0_  = n8571 ;
  assign \g62630/_0_  = n8572 ;
  assign \g62632/_0_  = n8573 ;
  assign \g62633/_0_  = n8574 ;
  assign \g62635/_0_  = n8575 ;
  assign \g62636/_0_  = n8576 ;
  assign \g62637/_0_  = n8577 ;
  assign \g62638/_0_  = n8578 ;
  assign \g62640/_0_  = n8579 ;
  assign \g62641/_0_  = n8580 ;
  assign \g62642/_0_  = n8581 ;
  assign \g62643/_0_  = n8582 ;
  assign \g62644/_0_  = n8583 ;
  assign \g62646/_0_  = n8584 ;
  assign \g62647/_0_  = n8585 ;
  assign \g62649/_0_  = n8586 ;
  assign \g62650/_0_  = n8587 ;
  assign \g62651/_0_  = n8588 ;
  assign \g62653/_0_  = n8589 ;
  assign \g62655/_0_  = n8590 ;
  assign \g62656/_0_  = n8591 ;
  assign \g62657/_0_  = n8592 ;
  assign \g62658/_0_  = n8593 ;
  assign \g62660/_0_  = n8594 ;
  assign \g62661/_0_  = n8595 ;
  assign \g62662/_0_  = n8596 ;
  assign \g62663/_0_  = n8597 ;
  assign \g62664/_0_  = n8598 ;
  assign \g62665/_0_  = n8599 ;
  assign \g62667/_0_  = n8600 ;
  assign \g62669/_0_  = n8601 ;
  assign \g62670/_0_  = n8602 ;
  assign \g62671/_0_  = n8603 ;
  assign \g62672/_0_  = n8604 ;
  assign \g62674/_0_  = n8605 ;
  assign \g62675/_0_  = n8606 ;
  assign \g62676/_0_  = n8607 ;
  assign \g62677/_0_  = n8608 ;
  assign \g62678/_0_  = n8609 ;
  assign \g62679/_0_  = n8610 ;
  assign \g62680/_0_  = n8611 ;
  assign \g62681/_0_  = n8612 ;
  assign \g62682/_0_  = n8613 ;
  assign \g62684/_0_  = n8614 ;
  assign \g62685/_0_  = n8615 ;
  assign \g62686/_0_  = n8616 ;
  assign \g62687/_0_  = n8617 ;
  assign \g62690/_0_  = n8618 ;
  assign \g62693/_0_  = n8619 ;
  assign \g62698/_0_  = n8620 ;
  assign \g62699/_0_  = n8621 ;
  assign \g62700/_0_  = n8622 ;
  assign \g62701/_0_  = n8623 ;
  assign \g62702/_0_  = n8624 ;
  assign \g62703/_0_  = n8625 ;
  assign \g62704/_0_  = n8626 ;
  assign \g62709/_0_  = n8627 ;
  assign \g62710/_0_  = n8628 ;
  assign \g62711/_0_  = n8629 ;
  assign \g62714/_0_  = n8630 ;
  assign \g62715/_0_  = n8631 ;
  assign \g62717/_0_  = n8632 ;
  assign \g62718/_0_  = n8633 ;
  assign \g62719/_0_  = n8634 ;
  assign \g62720/_0_  = n8635 ;
  assign \g62721/_0_  = n8636 ;
  assign \g62723/_0_  = n8637 ;
  assign \g62725/_0_  = n8638 ;
  assign \g62726/_0_  = n8639 ;
  assign \g62729/_0_  = n8640 ;
  assign \g62731/_0_  = n8641 ;
  assign \g62733/_0_  = n8642 ;
  assign \g62738/_0_  = n8643 ;
  assign \g62741/_0_  = n8644 ;
  assign \g62742/_0_  = n8645 ;
  assign \g62744/_0_  = n8646 ;
  assign \g62745/_0_  = n8647 ;
  assign \g62746/_0_  = n8648 ;
  assign \g62747/_0_  = n8649 ;
  assign \g62748/_0_  = n8650 ;
  assign \g62749/_0_  = n8651 ;
  assign \g62753/_0_  = n8652 ;
  assign \g62755/_0_  = n8653 ;
  assign \g62756/_0_  = n8654 ;
  assign \g62758/_0_  = n8655 ;
  assign \g62759/_0_  = n8656 ;
  assign \g62760/_0_  = n8657 ;
  assign \g62761/_0_  = n8658 ;
  assign \g62763/_0_  = n8659 ;
  assign \g62766/_0_  = n8660 ;
  assign \g62767/_0_  = n8661 ;
  assign \g62768/_0_  = n8662 ;
  assign \g65554/_0_  = ~n8668 ;
  assign \g65561/_0_  = ~n8674 ;
  assign \g65569/_0_  = ~n8680 ;
  assign \g65580/_0_  = ~n8686 ;
  assign \g65599/_0_  = ~n8692 ;
  assign \g65606/_0_  = ~n8698 ;
  assign \g65636/_0_  = ~n8704 ;
  assign \g65864/_0_  = ~n8710 ;
endmodule
