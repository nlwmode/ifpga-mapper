module top( \G0_pad  , \G10_pad  , \G11_pad  , \G12_pad  , \G13_pad  , \G14_pad  , \G15_pad  , \G16_pad  , \G18_pad  , \G1_pad  , \G2_pad  , \G38_reg/NET0131  , \G39_reg/NET0131  , \G3_pad  , \G40_reg/NET0131  , \G41_reg/NET0131  , \G42_reg/NET0131  , \G4_pad  , \G5_pad  , \G6_pad  , \G7_pad  , \G8_pad  , \G9_pad  , \G288_pad  , \G290_pad  , \G296_pad  , \G302_pad  , \G310_pad  , \G312_pad  , \G315_pad  , \G327_pad  , \G45_pad  , \G47_pad  , \G49_pad  , \G53_pad  , \G55_pad  , \_al_n0  , \_al_n1  , \g1452/_0_  , \g1456/_1_  , \g1462/_0_  , \g1463/_0_  , \g1504/_3_  , \g1524/_1_  , \g1524/_2_  , \g1527/_3_  , \g31/_0_  , \g45/_1_  );
  input \G0_pad  ;
  input \G10_pad  ;
  input \G11_pad  ;
  input \G12_pad  ;
  input \G13_pad  ;
  input \G14_pad  ;
  input \G15_pad  ;
  input \G16_pad  ;
  input \G18_pad  ;
  input \G1_pad  ;
  input \G2_pad  ;
  input \G38_reg/NET0131  ;
  input \G39_reg/NET0131  ;
  input \G3_pad  ;
  input \G40_reg/NET0131  ;
  input \G41_reg/NET0131  ;
  input \G42_reg/NET0131  ;
  input \G4_pad  ;
  input \G5_pad  ;
  input \G6_pad  ;
  input \G7_pad  ;
  input \G8_pad  ;
  input \G9_pad  ;
  output \G288_pad  ;
  output \G290_pad  ;
  output \G296_pad  ;
  output \G302_pad  ;
  output \G310_pad  ;
  output \G312_pad  ;
  output \G315_pad  ;
  output \G327_pad  ;
  output \G45_pad  ;
  output \G47_pad  ;
  output \G49_pad  ;
  output \G53_pad  ;
  output \G55_pad  ;
  output \_al_n0  ;
  output \_al_n1  ;
  output \g1452/_0_  ;
  output \g1456/_1_  ;
  output \g1462/_0_  ;
  output \g1463/_0_  ;
  output \g1504/_3_  ;
  output \g1524/_1_  ;
  output \g1524/_2_  ;
  output \g1527/_3_  ;
  output \g31/_0_  ;
  output \g45/_1_  ;
  wire n24 , n25 , n26 , n27 , n28 , n29 , n30 , n31 , n32 , n33 , n34 , n35 , n36 , n37 , n38 , n39 , n40 , n41 , n42 , n43 , n44 , n45 , n46 , n47 , n48 , n49 , n50 , n51 , n52 , n53 , n54 , n55 , n56 , n57 , n58 , n59 , n60 , n61 , n62 , n63 , n64 , n65 , n66 , n67 , n68 , n69 , n70 , n71 , n72 , n73 , n74 , n75 , n76 , n77 , n78 , n79 , n80 , n81 , n82 , n83 , n84 , n85 , n86 , n87 , n88 , n89 , n90 , n91 , n92 , n93 , n94 , n95 , n96 , n97 , n98 , n99 , n100 , n101 , n102 , n103 , n104 , n105 , n106 , n107 , n108 , n109 , n110 , n111 , n112 , n113 , n114 , n115 , n116 , n117 , n118 , n119 , n120 , n121 , n122 , n123 , n124 , n125 , n126 , n127 , n128 , n129 , n130 , n131 , n132 , n133 , n134 , n135 , n136 , n137 , n138 , n139 , n140 , n141 , n142 , n143 , n144 , n145 , n146 , n147 , n148 , n149 , n150 , n151 , n152 , n153 , n154 , n155 , n156 , n157 , n158 , n159 , n160 , n161 , n162 , n163 , n164 , n165 , n166 , n167 , n168 , n169 , n170 , n171 , n172 , n173 , n174 , n175 , n176 , n177 , n178 , n179 , n180 , n181 , n182 , n183 , n184 , n185 , n186 , n187 , n188 , n189 , n190 , n191 , n192 , n193 , n194 , n195 , n196 , n197 , n198 , n199 , n200 , n201 , n202 , n203 , n204 , n205 , n206 , n207 , n208 , n209 , n210 , n211 , n212 , n213 , n214 , n215 , n216 , n217 , n218 , n219 , n220 , n221 , n222 , n223 , n224 , n225 , n226 , n227 , n228 , n229 , n230 , n231 , n232 , n233 , n234 , n235 , n236 , n237 , n238 , n239 , n240 , n241 , n242 , n243 , n244 , n245 , n246 , n247 , n248 , n249 , n250 , n251 , n252 , n253 , n254 , n255 , n256 , n257 , n258 , n259 , n260 , n261 , n262 , n263 , n264 , n265 , n266 , n267 , n268 , n269 , n270 , n271 , n272 , n273 , n274 , n275 , n276 , n277 ;
  assign n24 = ~\G41_reg/NET0131  & ~\G42_reg/NET0131  ;
  assign n25 = ~\G38_reg/NET0131  & \G39_reg/NET0131  ;
  assign n26 = \G40_reg/NET0131  & n25 ;
  assign n27 = n24 & n26 ;
  assign n28 = \G15_pad  & ~\G42_reg/NET0131  ;
  assign n29 = ~\G40_reg/NET0131  & ~\G41_reg/NET0131  ;
  assign n30 = \G39_reg/NET0131  & n29 ;
  assign n31 = n28 & n30 ;
  assign n32 = \G40_reg/NET0131  & \G41_reg/NET0131  ;
  assign n33 = ~\G42_reg/NET0131  & n32 ;
  assign n34 = n25 & n33 ;
  assign n39 = ~\G38_reg/NET0131  & ~\G39_reg/NET0131  ;
  assign n40 = \G16_pad  & ~\G4_pad  ;
  assign n41 = \G40_reg/NET0131  & ~n40 ;
  assign n42 = \G16_pad  & ~\G40_reg/NET0131  ;
  assign n43 = ~\G1_pad  & n24 ;
  assign n44 = n42 & n43 ;
  assign n45 = ~n41 & ~n44 ;
  assign n46 = n39 & ~n45 ;
  assign n52 = \G38_reg/NET0131  & n24 ;
  assign n53 = \G40_reg/NET0131  & ~n52 ;
  assign n54 = \G39_reg/NET0131  & \G4_pad  ;
  assign n55 = ~n53 & n54 ;
  assign n35 = \G39_reg/NET0131  & ~\G40_reg/NET0131  ;
  assign n36 = \G41_reg/NET0131  & \G42_reg/NET0131  ;
  assign n37 = ~\G16_pad  & ~n36 ;
  assign n38 = n35 & n37 ;
  assign n48 = ~\G39_reg/NET0131  & \G41_reg/NET0131  ;
  assign n47 = \G38_reg/NET0131  & ~\G40_reg/NET0131  ;
  assign n49 = \G42_reg/NET0131  & ~n47 ;
  assign n50 = n48 & n49 ;
  assign n51 = ~n40 & n50 ;
  assign n56 = ~n38 & ~n51 ;
  assign n57 = ~n55 & n56 ;
  assign n58 = ~n46 & n57 ;
  assign n59 = ~\G41_reg/NET0131  & \G42_reg/NET0131  ;
  assign n60 = n26 & n59 ;
  assign n62 = ~\G38_reg/NET0131  & n36 ;
  assign n61 = \G39_reg/NET0131  & \G40_reg/NET0131  ;
  assign n63 = \G16_pad  & n61 ;
  assign n64 = n62 & n63 ;
  assign n65 = ~\G39_reg/NET0131  & ~\G40_reg/NET0131  ;
  assign n66 = n24 & n65 ;
  assign n67 = \G40_reg/NET0131  & n36 ;
  assign n68 = \G39_reg/NET0131  & n67 ;
  assign n69 = ~n66 & ~n68 ;
  assign n70 = ~\G38_reg/NET0131  & ~n69 ;
  assign n71 = \G15_pad  & \G42_reg/NET0131  ;
  assign n72 = n30 & n71 ;
  assign n75 = n33 & n40 ;
  assign n73 = \G10_pad  & \G11_pad  ;
  assign n74 = ~\G12_pad  & ~n73 ;
  assign n76 = ~\G10_pad  & ~\G11_pad  ;
  assign n77 = \G15_pad  & n39 ;
  assign n78 = ~n76 & n77 ;
  assign n79 = ~n74 & n78 ;
  assign n80 = n75 & n79 ;
  assign n81 = ~\G5_pad  & n27 ;
  assign n82 = \G38_reg/NET0131  & ~\G39_reg/NET0131  ;
  assign n83 = ~n61 & ~n65 ;
  assign n84 = ~n52 & ~n83 ;
  assign n85 = ~n82 & ~n84 ;
  assign n86 = ~n50 & ~n85 ;
  assign n87 = ~\G40_reg/NET0131  & ~\G42_reg/NET0131  ;
  assign n88 = \G41_reg/NET0131  & n87 ;
  assign n89 = n39 & n88 ;
  assign n90 = \G5_pad  & n27 ;
  assign n91 = \G13_pad  & \G15_pad  ;
  assign n92 = \G42_reg/NET0131  & ~n91 ;
  assign n93 = ~\G38_reg/NET0131  & n28 ;
  assign n94 = ~n92 & ~n93 ;
  assign n95 = \G40_reg/NET0131  & ~n94 ;
  assign n96 = ~\G39_reg/NET0131  & ~n95 ;
  assign n97 = \G6_pad  & \G7_pad  ;
  assign n98 = \G8_pad  & \G9_pad  ;
  assign n99 = n97 & n98 ;
  assign n100 = ~\G40_reg/NET0131  & ~n99 ;
  assign n101 = \G38_reg/NET0131  & \G39_reg/NET0131  ;
  assign n102 = ~n100 & n101 ;
  assign n103 = ~\G15_pad  & ~\G40_reg/NET0131  ;
  assign n104 = \G41_reg/NET0131  & ~n103 ;
  assign n105 = ~n102 & n104 ;
  assign n106 = ~n96 & n105 ;
  assign n111 = ~\G7_pad  & ~\G8_pad  ;
  assign n112 = \G9_pad  & n111 ;
  assign n109 = \G15_pad  & \G40_reg/NET0131  ;
  assign n110 = ~\G42_reg/NET0131  & \G6_pad  ;
  assign n113 = n109 & n110 ;
  assign n114 = n112 & n113 ;
  assign n107 = ~\G1_pad  & n29 ;
  assign n108 = ~\G15_pad  & \G42_reg/NET0131  ;
  assign n115 = ~n107 & ~n108 ;
  assign n116 = ~n114 & n115 ;
  assign n117 = n39 & ~n116 ;
  assign n118 = ~n28 & ~n108 ;
  assign n119 = \G39_reg/NET0131  & ~n118 ;
  assign n120 = ~\G39_reg/NET0131  & ~\G41_reg/NET0131  ;
  assign n121 = \G42_reg/NET0131  & n120 ;
  assign n122 = ~n119 & ~n121 ;
  assign n123 = ~\G40_reg/NET0131  & ~n122 ;
  assign n124 = ~n117 & ~n123 ;
  assign n125 = ~n106 & n124 ;
  assign n126 = \G16_pad  & ~n125 ;
  assign n127 = ~\G41_reg/NET0131  & \G5_pad  ;
  assign n128 = ~\G42_reg/NET0131  & ~n127 ;
  assign n129 = ~\G1_pad  & ~\G3_pad  ;
  assign n130 = n59 & n129 ;
  assign n131 = ~\G2_pad  & n130 ;
  assign n132 = ~n128 & ~n131 ;
  assign n133 = n61 & ~n132 ;
  assign n134 = ~\G40_reg/NET0131  & ~n36 ;
  assign n135 = \G4_pad  & ~n134 ;
  assign n136 = \G14_pad  & \G15_pad  ;
  assign n137 = n88 & n136 ;
  assign n138 = ~n135 & ~n137 ;
  assign n139 = ~\G39_reg/NET0131  & ~n138 ;
  assign n140 = ~n133 & ~n139 ;
  assign n141 = ~\G38_reg/NET0131  & ~n140 ;
  assign n142 = ~\G39_reg/NET0131  & \G4_pad  ;
  assign n143 = ~\G0_pad  & \G38_reg/NET0131  ;
  assign n144 = \G39_reg/NET0131  & n143 ;
  assign n145 = ~n142 & ~n144 ;
  assign n146 = n67 & ~n145 ;
  assign n147 = ~n55 & ~n146 ;
  assign n148 = ~n141 & n147 ;
  assign n149 = ~n126 & n148 ;
  assign n150 = ~\G18_pad  & ~n149 ;
  assign n172 = ~\G38_reg/NET0131  & ~n128 ;
  assign n173 = ~n130 & n172 ;
  assign n169 = ~\G4_pad  & n24 ;
  assign n168 = ~\G0_pad  & n36 ;
  assign n170 = \G38_reg/NET0131  & ~n168 ;
  assign n171 = ~n169 & n170 ;
  assign n174 = n61 & ~n171 ;
  assign n175 = ~n173 & n174 ;
  assign n176 = \G2_pad  & n129 ;
  assign n177 = ~\G16_pad  & n176 ;
  assign n178 = ~\G41_reg/NET0131  & ~n177 ;
  assign n179 = ~\G14_pad  & \G15_pad  ;
  assign n180 = \G41_reg/NET0131  & ~n179 ;
  assign n181 = n87 & ~n180 ;
  assign n182 = n39 & n181 ;
  assign n183 = ~n178 & n182 ;
  assign n152 = \G38_reg/NET0131  & ~n36 ;
  assign n153 = ~\G39_reg/NET0131  & ~\G4_pad  ;
  assign n157 = \G16_pad  & ~n103 ;
  assign n158 = n153 & n157 ;
  assign n159 = ~n152 & n158 ;
  assign n151 = ~\G40_reg/NET0131  & ~n62 ;
  assign n154 = ~\G42_reg/NET0131  & ~n76 ;
  assign n155 = \G15_pad  & n32 ;
  assign n156 = ~n154 & n155 ;
  assign n160 = ~n151 & ~n156 ;
  assign n161 = n159 & n160 ;
  assign n162 = \G15_pad  & \G38_reg/NET0131  ;
  assign n163 = n99 & n162 ;
  assign n164 = \G16_pad  & ~n163 ;
  assign n165 = ~\G4_pad  & n35 ;
  assign n166 = n36 & n165 ;
  assign n167 = ~n164 & n166 ;
  assign n184 = ~n161 & ~n167 ;
  assign n185 = ~n183 & n184 ;
  assign n186 = ~n175 & n185 ;
  assign n187 = ~\G18_pad  & ~n186 ;
  assign n195 = ~\G38_reg/NET0131  & n66 ;
  assign n196 = n177 & n195 ;
  assign n188 = ~n37 & n165 ;
  assign n189 = n74 & n154 ;
  assign n191 = n40 & n48 ;
  assign n190 = \G38_reg/NET0131  & ~\G42_reg/NET0131  ;
  assign n192 = n109 & ~n190 ;
  assign n193 = n191 & n192 ;
  assign n194 = ~n189 & n193 ;
  assign n197 = ~n188 & ~n194 ;
  assign n198 = ~n196 & n197 ;
  assign n199 = ~n175 & n198 ;
  assign n200 = ~\G18_pad  & ~n199 ;
  assign n201 = ~\G16_pad  & ~\G1_pad  ;
  assign n202 = ~\G38_reg/NET0131  & n201 ;
  assign n206 = n29 & ~n202 ;
  assign n203 = \G0_pad  & n190 ;
  assign n204 = \G16_pad  & \G38_reg/NET0131  ;
  assign n205 = \G42_reg/NET0131  & ~n204 ;
  assign n207 = ~n203 & ~n205 ;
  assign n208 = n206 & n207 ;
  assign n209 = \G10_pad  & \G12_pad  ;
  assign n210 = ~\G11_pad  & ~n209 ;
  assign n211 = \G15_pad  & ~\G38_reg/NET0131  ;
  assign n212 = ~n210 & n211 ;
  assign n213 = n75 & n212 ;
  assign n214 = ~n208 & ~n213 ;
  assign n215 = ~\G39_reg/NET0131  & ~n214 ;
  assign n219 = \G41_reg/NET0131  & ~n143 ;
  assign n216 = \G1_pad  & ~\G38_reg/NET0131  ;
  assign n217 = ~\G41_reg/NET0131  & ~n216 ;
  assign n218 = \G42_reg/NET0131  & n61 ;
  assign n220 = ~n217 & n218 ;
  assign n221 = ~n219 & n220 ;
  assign n222 = ~\G4_pad  & ~n65 ;
  assign n223 = ~n120 & n204 ;
  assign n224 = n222 & n223 ;
  assign n225 = ~n33 & ~n218 ;
  assign n226 = n224 & n225 ;
  assign n227 = ~n221 & ~n226 ;
  assign n228 = ~n215 & n227 ;
  assign n229 = ~\G18_pad  & ~n228 ;
  assign n231 = \G39_reg/NET0131  & ~\G42_reg/NET0131  ;
  assign n232 = ~\G41_reg/NET0131  & ~n231 ;
  assign n230 = ~n61 & ~n87 ;
  assign n233 = n216 & ~n230 ;
  assign n234 = n232 & n233 ;
  assign n235 = \G15_pad  & n89 ;
  assign n236 = n39 & n137 ;
  assign n237 = \G3_pad  & n66 ;
  assign n238 = n202 & n237 ;
  assign n252 = ~\G39_reg/NET0131  & ~n135 ;
  assign n249 = n59 & n109 ;
  assign n250 = \G16_pad  & ~n87 ;
  assign n251 = ~n249 & n250 ;
  assign n253 = ~n181 & ~n251 ;
  assign n254 = n252 & n253 ;
  assign n239 = ~\G41_reg/NET0131  & ~\G5_pad  ;
  assign n242 = \G40_reg/NET0131  & ~n142 ;
  assign n243 = ~n239 & n242 ;
  assign n240 = ~\G16_pad  & \G39_reg/NET0131  ;
  assign n241 = \G42_reg/NET0131  & ~n240 ;
  assign n244 = ~n232 & ~n241 ;
  assign n245 = n243 & n244 ;
  assign n246 = ~n42 & ~n83 ;
  assign n247 = n176 & n232 ;
  assign n248 = n246 & n247 ;
  assign n255 = ~n245 & ~n248 ;
  assign n256 = ~n254 & n255 ;
  assign n257 = ~\G38_reg/NET0131  & ~n256 ;
  assign n266 = \G39_reg/NET0131  & n71 ;
  assign n267 = ~n99 & n266 ;
  assign n268 = \G15_pad  & ~n25 ;
  assign n269 = \G41_reg/NET0131  & ~n82 ;
  assign n270 = ~n268 & n269 ;
  assign n271 = ~n267 & ~n270 ;
  assign n272 = ~\G40_reg/NET0131  & n40 ;
  assign n273 = ~n271 & n272 ;
  assign n258 = \G16_pad  & n91 ;
  assign n259 = n153 & ~n258 ;
  assign n260 = ~n144 & ~n259 ;
  assign n261 = n67 & ~n260 ;
  assign n262 = \G16_pad  & ~\G41_reg/NET0131  ;
  assign n263 = ~n71 & n262 ;
  assign n264 = ~n36 & n165 ;
  assign n265 = ~n263 & n264 ;
  assign n274 = ~n261 & ~n265 ;
  assign n275 = ~n273 & n274 ;
  assign n276 = ~n257 & n275 ;
  assign n277 = ~\G18_pad  & ~n276 ;
  assign \G288_pad  = n27 ;
  assign \G290_pad  = n31 ;
  assign \G296_pad  = n34 ;
  assign \G302_pad  = ~n58 ;
  assign \G310_pad  = n60 ;
  assign \G312_pad  = n64 ;
  assign \G315_pad  = n70 ;
  assign \G327_pad  = n72 ;
  assign \G45_pad  = n80 ;
  assign \G47_pad  = n81 ;
  assign \G49_pad  = ~n86 ;
  assign \G53_pad  = n89 ;
  assign \G55_pad  = n90 ;
  assign \_al_n0  = 1'b0 ;
  assign \_al_n1  = ~1'b0 ;
  assign \g1452/_0_  = n150 ;
  assign \g1456/_1_  = n187 ;
  assign \g1462/_0_  = n200 ;
  assign \g1463/_0_  = n229 ;
  assign \g1504/_3_  = n234 ;
  assign \g1524/_1_  = n235 ;
  assign \g1524/_2_  = n236 ;
  assign \g1527/_3_  = n238 ;
  assign \g31/_0_  = n277 ;
  assign \g45/_1_  = n167 ;
endmodule
