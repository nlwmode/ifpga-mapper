module top (\A[0] , \A[1] , \A[2] , \A[3] , \A[4] , \A[5] , \A[6] , \A[7] , \A[8] , \A[9] , \A[10] , \A[11] , \A[12] , \A[13] , \A[14] , \A[15] , \A[16] , \A[17] , \A[18] , \A[19] , \A[20] , \A[21] , \A[22] , \A[23] , \A[24] , \A[25] , \A[26] , \A[27] , \A[28] , \A[29] , \A[30] , \A[31] , \A[32] , \A[33] , \A[34] , \A[35] , \A[36] , \A[37] , \A[38] , \A[39] , \A[40] , \A[41] , \A[42] , \A[43] , \A[44] , \A[45] , \A[46] , \A[47] , \A[48] , \A[49] , \A[50] , \A[51] , \A[52] , \A[53] , \A[54] , \A[55] , \A[56] , \A[57] , \A[58] , \A[59] , \A[60] , \A[61] , \A[62] , \A[63] , \A[64] , \A[65] , \A[66] , \A[67] , \A[68] , \A[69] , \A[70] , \A[71] , \A[72] , \A[73] , \A[74] , \A[75] , \A[76] , \A[77] , \A[78] , \A[79] , \A[80] , \A[81] , \A[82] , \A[83] , \A[84] , \A[85] , \A[86] , \A[87] , \A[88] , \A[89] , \A[90] , \A[91] , \A[92] , \A[93] , \A[94] , \A[95] , \A[96] , \A[97] , \A[98] , \A[99] , \A[100] , \A[101] , \A[102] , \A[103] , \A[104] , \A[105] , \A[106] , \A[107] , \A[108] , \A[109] , \A[110] , \A[111] , \A[112] , \A[113] , \A[114] , \A[115] , \A[116] , \A[117] , \A[118] , \A[119] , \A[120] , \A[121] , \A[122] , \A[123] , \A[124] , \A[125] , \A[126] , \A[127] , \P[0] , \P[1] , \P[2] , \P[3] , \P[4] , \P[5] , \P[6] , F);
	input \A[0]  ;
	input \A[1]  ;
	input \A[2]  ;
	input \A[3]  ;
	input \A[4]  ;
	input \A[5]  ;
	input \A[6]  ;
	input \A[7]  ;
	input \A[8]  ;
	input \A[9]  ;
	input \A[10]  ;
	input \A[11]  ;
	input \A[12]  ;
	input \A[13]  ;
	input \A[14]  ;
	input \A[15]  ;
	input \A[16]  ;
	input \A[17]  ;
	input \A[18]  ;
	input \A[19]  ;
	input \A[20]  ;
	input \A[21]  ;
	input \A[22]  ;
	input \A[23]  ;
	input \A[24]  ;
	input \A[25]  ;
	input \A[26]  ;
	input \A[27]  ;
	input \A[28]  ;
	input \A[29]  ;
	input \A[30]  ;
	input \A[31]  ;
	input \A[32]  ;
	input \A[33]  ;
	input \A[34]  ;
	input \A[35]  ;
	input \A[36]  ;
	input \A[37]  ;
	input \A[38]  ;
	input \A[39]  ;
	input \A[40]  ;
	input \A[41]  ;
	input \A[42]  ;
	input \A[43]  ;
	input \A[44]  ;
	input \A[45]  ;
	input \A[46]  ;
	input \A[47]  ;
	input \A[48]  ;
	input \A[49]  ;
	input \A[50]  ;
	input \A[51]  ;
	input \A[52]  ;
	input \A[53]  ;
	input \A[54]  ;
	input \A[55]  ;
	input \A[56]  ;
	input \A[57]  ;
	input \A[58]  ;
	input \A[59]  ;
	input \A[60]  ;
	input \A[61]  ;
	input \A[62]  ;
	input \A[63]  ;
	input \A[64]  ;
	input \A[65]  ;
	input \A[66]  ;
	input \A[67]  ;
	input \A[68]  ;
	input \A[69]  ;
	input \A[70]  ;
	input \A[71]  ;
	input \A[72]  ;
	input \A[73]  ;
	input \A[74]  ;
	input \A[75]  ;
	input \A[76]  ;
	input \A[77]  ;
	input \A[78]  ;
	input \A[79]  ;
	input \A[80]  ;
	input \A[81]  ;
	input \A[82]  ;
	input \A[83]  ;
	input \A[84]  ;
	input \A[85]  ;
	input \A[86]  ;
	input \A[87]  ;
	input \A[88]  ;
	input \A[89]  ;
	input \A[90]  ;
	input \A[91]  ;
	input \A[92]  ;
	input \A[93]  ;
	input \A[94]  ;
	input \A[95]  ;
	input \A[96]  ;
	input \A[97]  ;
	input \A[98]  ;
	input \A[99]  ;
	input \A[100]  ;
	input \A[101]  ;
	input \A[102]  ;
	input \A[103]  ;
	input \A[104]  ;
	input \A[105]  ;
	input \A[106]  ;
	input \A[107]  ;
	input \A[108]  ;
	input \A[109]  ;
	input \A[110]  ;
	input \A[111]  ;
	input \A[112]  ;
	input \A[113]  ;
	input \A[114]  ;
	input \A[115]  ;
	input \A[116]  ;
	input \A[117]  ;
	input \A[118]  ;
	input \A[119]  ;
	input \A[120]  ;
	input \A[121]  ;
	input \A[122]  ;
	input \A[123]  ;
	input \A[124]  ;
	input \A[125]  ;
	input \A[126]  ;
	input \A[127]  ;
	output \P[0]  ;
	output \P[1]  ;
	output \P[2]  ;
	output \P[3]  ;
	output \P[4]  ;
	output \P[5]  ;
	output \P[6]  ;
	output F ;
	wire _w400_ ;
	wire _w399_ ;
	wire _w398_ ;
	wire _w397_ ;
	wire _w396_ ;
	wire _w395_ ;
	wire _w394_ ;
	wire _w393_ ;
	wire _w392_ ;
	wire _w391_ ;
	wire _w390_ ;
	wire _w389_ ;
	wire _w388_ ;
	wire _w387_ ;
	wire _w256_ ;
	wire _w255_ ;
	wire _w254_ ;
	wire _w253_ ;
	wire _w252_ ;
	wire _w251_ ;
	wire _w250_ ;
	wire _w249_ ;
	wire _w248_ ;
	wire _w247_ ;
	wire _w246_ ;
	wire _w245_ ;
	wire _w244_ ;
	wire _w243_ ;
	wire _w242_ ;
	wire _w241_ ;
	wire _w240_ ;
	wire _w239_ ;
	wire _w238_ ;
	wire _w237_ ;
	wire _w236_ ;
	wire _w235_ ;
	wire _w234_ ;
	wire _w233_ ;
	wire _w232_ ;
	wire _w231_ ;
	wire _w230_ ;
	wire _w229_ ;
	wire _w228_ ;
	wire _w227_ ;
	wire _w226_ ;
	wire _w225_ ;
	wire _w224_ ;
	wire _w223_ ;
	wire _w222_ ;
	wire _w221_ ;
	wire _w220_ ;
	wire _w219_ ;
	wire _w218_ ;
	wire _w217_ ;
	wire _w216_ ;
	wire _w215_ ;
	wire _w214_ ;
	wire _w213_ ;
	wire _w212_ ;
	wire _w211_ ;
	wire _w210_ ;
	wire _w209_ ;
	wire _w208_ ;
	wire _w207_ ;
	wire _w206_ ;
	wire _w205_ ;
	wire _w204_ ;
	wire _w203_ ;
	wire _w202_ ;
	wire _w201_ ;
	wire _w200_ ;
	wire _w199_ ;
	wire _w198_ ;
	wire _w197_ ;
	wire _w196_ ;
	wire _w195_ ;
	wire _w194_ ;
	wire _w193_ ;
	wire _w192_ ;
	wire _w191_ ;
	wire _w190_ ;
	wire _w189_ ;
	wire _w158_ ;
	wire _w157_ ;
	wire _w156_ ;
	wire _w155_ ;
	wire _w154_ ;
	wire _w153_ ;
	wire _w152_ ;
	wire _w151_ ;
	wire _w150_ ;
	wire _w149_ ;
	wire _w148_ ;
	wire _w147_ ;
	wire _w146_ ;
	wire _w145_ ;
	wire _w144_ ;
	wire _w143_ ;
	wire _w130_ ;
	wire _w131_ ;
	wire _w132_ ;
	wire _w133_ ;
	wire _w134_ ;
	wire _w135_ ;
	wire _w136_ ;
	wire _w137_ ;
	wire _w138_ ;
	wire _w139_ ;
	wire _w140_ ;
	wire _w141_ ;
	wire _w142_ ;
	wire _w159_ ;
	wire _w160_ ;
	wire _w161_ ;
	wire _w162_ ;
	wire _w163_ ;
	wire _w164_ ;
	wire _w165_ ;
	wire _w166_ ;
	wire _w167_ ;
	wire _w168_ ;
	wire _w169_ ;
	wire _w170_ ;
	wire _w171_ ;
	wire _w172_ ;
	wire _w173_ ;
	wire _w174_ ;
	wire _w175_ ;
	wire _w176_ ;
	wire _w177_ ;
	wire _w178_ ;
	wire _w179_ ;
	wire _w180_ ;
	wire _w181_ ;
	wire _w182_ ;
	wire _w183_ ;
	wire _w184_ ;
	wire _w185_ ;
	wire _w186_ ;
	wire _w187_ ;
	wire _w188_ ;
	wire _w257_ ;
	wire _w258_ ;
	wire _w259_ ;
	wire _w260_ ;
	wire _w261_ ;
	wire _w262_ ;
	wire _w263_ ;
	wire _w264_ ;
	wire _w265_ ;
	wire _w266_ ;
	wire _w267_ ;
	wire _w268_ ;
	wire _w269_ ;
	wire _w270_ ;
	wire _w271_ ;
	wire _w272_ ;
	wire _w273_ ;
	wire _w274_ ;
	wire _w275_ ;
	wire _w276_ ;
	wire _w277_ ;
	wire _w278_ ;
	wire _w279_ ;
	wire _w280_ ;
	wire _w281_ ;
	wire _w282_ ;
	wire _w283_ ;
	wire _w284_ ;
	wire _w285_ ;
	wire _w286_ ;
	wire _w287_ ;
	wire _w288_ ;
	wire _w289_ ;
	wire _w290_ ;
	wire _w291_ ;
	wire _w292_ ;
	wire _w293_ ;
	wire _w294_ ;
	wire _w295_ ;
	wire _w296_ ;
	wire _w297_ ;
	wire _w298_ ;
	wire _w299_ ;
	wire _w300_ ;
	wire _w301_ ;
	wire _w302_ ;
	wire _w303_ ;
	wire _w304_ ;
	wire _w305_ ;
	wire _w306_ ;
	wire _w307_ ;
	wire _w308_ ;
	wire _w309_ ;
	wire _w310_ ;
	wire _w311_ ;
	wire _w312_ ;
	wire _w313_ ;
	wire _w314_ ;
	wire _w315_ ;
	wire _w316_ ;
	wire _w317_ ;
	wire _w318_ ;
	wire _w319_ ;
	wire _w320_ ;
	wire _w321_ ;
	wire _w322_ ;
	wire _w323_ ;
	wire _w324_ ;
	wire _w325_ ;
	wire _w326_ ;
	wire _w327_ ;
	wire _w328_ ;
	wire _w329_ ;
	wire _w330_ ;
	wire _w331_ ;
	wire _w332_ ;
	wire _w333_ ;
	wire _w334_ ;
	wire _w335_ ;
	wire _w336_ ;
	wire _w337_ ;
	wire _w338_ ;
	wire _w339_ ;
	wire _w340_ ;
	wire _w341_ ;
	wire _w342_ ;
	wire _w343_ ;
	wire _w344_ ;
	wire _w345_ ;
	wire _w346_ ;
	wire _w347_ ;
	wire _w348_ ;
	wire _w349_ ;
	wire _w350_ ;
	wire _w351_ ;
	wire _w352_ ;
	wire _w353_ ;
	wire _w354_ ;
	wire _w355_ ;
	wire _w356_ ;
	wire _w357_ ;
	wire _w358_ ;
	wire _w359_ ;
	wire _w360_ ;
	wire _w361_ ;
	wire _w362_ ;
	wire _w363_ ;
	wire _w364_ ;
	wire _w365_ ;
	wire _w366_ ;
	wire _w367_ ;
	wire _w368_ ;
	wire _w369_ ;
	wire _w370_ ;
	wire _w371_ ;
	wire _w372_ ;
	wire _w373_ ;
	wire _w374_ ;
	wire _w375_ ;
	wire _w376_ ;
	wire _w377_ ;
	wire _w378_ ;
	wire _w379_ ;
	wire _w380_ ;
	wire _w381_ ;
	wire _w382_ ;
	wire _w383_ ;
	wire _w384_ ;
	wire _w385_ ;
	wire _w386_ ;
	LUT2 #(
		.INIT('h2)
	) name0 (
		\A[76] ,
		\A[77] ,
		_w130_
	);
	LUT4 #(
		.INIT('h000d)
	) name1 (
		\A[73] ,
		\A[74] ,
		\A[75] ,
		\A[77] ,
		_w131_
	);
	LUT2 #(
		.INIT('h1)
	) name2 (
		_w130_,
		_w131_,
		_w132_
	);
	LUT4 #(
		.INIT('h000d)
	) name3 (
		\A[64] ,
		\A[65] ,
		\A[66] ,
		\A[68] ,
		_w133_
	);
	LUT4 #(
		.INIT('h000d)
	) name4 (
		\A[67] ,
		\A[68] ,
		\A[69] ,
		\A[71] ,
		_w134_
	);
	LUT2 #(
		.INIT('h4)
	) name5 (
		_w133_,
		_w134_,
		_w135_
	);
	LUT4 #(
		.INIT('h000d)
	) name6 (
		\A[55] ,
		\A[56] ,
		\A[57] ,
		\A[59] ,
		_w136_
	);
	LUT4 #(
		.INIT('h000d)
	) name7 (
		\A[58] ,
		\A[59] ,
		\A[60] ,
		\A[62] ,
		_w137_
	);
	LUT2 #(
		.INIT('h4)
	) name8 (
		_w136_,
		_w137_,
		_w138_
	);
	LUT4 #(
		.INIT('h000d)
	) name9 (
		\A[46] ,
		\A[47] ,
		\A[48] ,
		\A[50] ,
		_w139_
	);
	LUT4 #(
		.INIT('h000d)
	) name10 (
		\A[49] ,
		\A[50] ,
		\A[51] ,
		\A[53] ,
		_w140_
	);
	LUT2 #(
		.INIT('h4)
	) name11 (
		_w139_,
		_w140_,
		_w141_
	);
	LUT4 #(
		.INIT('h000d)
	) name12 (
		\A[37] ,
		\A[38] ,
		\A[39] ,
		\A[41] ,
		_w142_
	);
	LUT4 #(
		.INIT('h000d)
	) name13 (
		\A[40] ,
		\A[41] ,
		\A[42] ,
		\A[44] ,
		_w143_
	);
	LUT2 #(
		.INIT('h4)
	) name14 (
		_w142_,
		_w143_,
		_w144_
	);
	LUT4 #(
		.INIT('h000d)
	) name15 (
		\A[28] ,
		\A[29] ,
		\A[30] ,
		\A[32] ,
		_w145_
	);
	LUT4 #(
		.INIT('h000d)
	) name16 (
		\A[31] ,
		\A[32] ,
		\A[33] ,
		\A[35] ,
		_w146_
	);
	LUT2 #(
		.INIT('h4)
	) name17 (
		_w145_,
		_w146_,
		_w147_
	);
	LUT4 #(
		.INIT('h000d)
	) name18 (
		\A[19] ,
		\A[20] ,
		\A[21] ,
		\A[23] ,
		_w148_
	);
	LUT4 #(
		.INIT('h000d)
	) name19 (
		\A[22] ,
		\A[23] ,
		\A[24] ,
		\A[26] ,
		_w149_
	);
	LUT2 #(
		.INIT('h4)
	) name20 (
		_w148_,
		_w149_,
		_w150_
	);
	LUT4 #(
		.INIT('h000d)
	) name21 (
		\A[10] ,
		\A[11] ,
		\A[12] ,
		\A[14] ,
		_w151_
	);
	LUT4 #(
		.INIT('h000d)
	) name22 (
		\A[13] ,
		\A[14] ,
		\A[15] ,
		\A[17] ,
		_w152_
	);
	LUT2 #(
		.INIT('h4)
	) name23 (
		_w151_,
		_w152_,
		_w153_
	);
	LUT4 #(
		.INIT('h000d)
	) name24 (
		\A[1] ,
		\A[2] ,
		\A[3] ,
		\A[5] ,
		_w154_
	);
	LUT4 #(
		.INIT('h000d)
	) name25 (
		\A[4] ,
		\A[5] ,
		\A[6] ,
		\A[8] ,
		_w155_
	);
	LUT4 #(
		.INIT('h000d)
	) name26 (
		\A[7] ,
		\A[8] ,
		\A[9] ,
		\A[11] ,
		_w156_
	);
	LUT4 #(
		.INIT('h8a00)
	) name27 (
		_w152_,
		_w154_,
		_w155_,
		_w156_,
		_w157_
	);
	LUT4 #(
		.INIT('h000d)
	) name28 (
		\A[16] ,
		\A[17] ,
		\A[18] ,
		\A[20] ,
		_w158_
	);
	LUT2 #(
		.INIT('h8)
	) name29 (
		_w149_,
		_w158_,
		_w159_
	);
	LUT4 #(
		.INIT('h5455)
	) name30 (
		_w150_,
		_w153_,
		_w157_,
		_w159_,
		_w160_
	);
	LUT4 #(
		.INIT('h000d)
	) name31 (
		\A[25] ,
		\A[26] ,
		\A[27] ,
		\A[29] ,
		_w161_
	);
	LUT2 #(
		.INIT('h8)
	) name32 (
		_w146_,
		_w161_,
		_w162_
	);
	LUT4 #(
		.INIT('h000d)
	) name33 (
		\A[34] ,
		\A[35] ,
		\A[36] ,
		\A[38] ,
		_w163_
	);
	LUT2 #(
		.INIT('h8)
	) name34 (
		_w143_,
		_w163_,
		_w164_
	);
	LUT4 #(
		.INIT('h1500)
	) name35 (
		_w147_,
		_w160_,
		_w162_,
		_w164_,
		_w165_
	);
	LUT4 #(
		.INIT('h000d)
	) name36 (
		\A[43] ,
		\A[44] ,
		\A[45] ,
		\A[47] ,
		_w166_
	);
	LUT2 #(
		.INIT('h8)
	) name37 (
		_w140_,
		_w166_,
		_w167_
	);
	LUT4 #(
		.INIT('h5455)
	) name38 (
		_w141_,
		_w144_,
		_w165_,
		_w167_,
		_w168_
	);
	LUT4 #(
		.INIT('h000d)
	) name39 (
		\A[52] ,
		\A[53] ,
		\A[54] ,
		\A[56] ,
		_w169_
	);
	LUT2 #(
		.INIT('h8)
	) name40 (
		_w137_,
		_w169_,
		_w170_
	);
	LUT4 #(
		.INIT('h000d)
	) name41 (
		\A[61] ,
		\A[62] ,
		\A[63] ,
		\A[65] ,
		_w171_
	);
	LUT2 #(
		.INIT('h8)
	) name42 (
		_w134_,
		_w171_,
		_w172_
	);
	LUT4 #(
		.INIT('h1500)
	) name43 (
		_w138_,
		_w168_,
		_w170_,
		_w172_,
		_w173_
	);
	LUT4 #(
		.INIT('h000d)
	) name44 (
		\A[70] ,
		\A[71] ,
		\A[72] ,
		\A[74] ,
		_w174_
	);
	LUT2 #(
		.INIT('h4)
	) name45 (
		_w130_,
		_w174_,
		_w175_
	);
	LUT4 #(
		.INIT('h5455)
	) name46 (
		_w132_,
		_w135_,
		_w173_,
		_w175_,
		_w176_
	);
	LUT2 #(
		.INIT('h1)
	) name47 (
		\A[78] ,
		\A[80] ,
		_w177_
	);
	LUT4 #(
		.INIT('h000d)
	) name48 (
		\A[79] ,
		\A[80] ,
		\A[81] ,
		\A[83] ,
		_w178_
	);
	LUT3 #(
		.INIT('h0d)
	) name49 (
		\A[82] ,
		\A[83] ,
		\A[84] ,
		_w179_
	);
	LUT4 #(
		.INIT('h4f00)
	) name50 (
		_w176_,
		_w177_,
		_w178_,
		_w179_,
		_w180_
	);
	LUT2 #(
		.INIT('h2)
	) name51 (
		\A[126] ,
		\A[127] ,
		_w181_
	);
	LUT4 #(
		.INIT('h000d)
	) name52 (
		\A[120] ,
		\A[121] ,
		\A[122] ,
		\A[124] ,
		_w182_
	);
	LUT4 #(
		.INIT('h000d)
	) name53 (
		\A[123] ,
		\A[124] ,
		\A[125] ,
		\A[127] ,
		_w183_
	);
	LUT2 #(
		.INIT('h4)
	) name54 (
		_w182_,
		_w183_,
		_w184_
	);
	LUT4 #(
		.INIT('h000d)
	) name55 (
		\A[111] ,
		\A[112] ,
		\A[113] ,
		\A[115] ,
		_w185_
	);
	LUT4 #(
		.INIT('h000d)
	) name56 (
		\A[114] ,
		\A[115] ,
		\A[116] ,
		\A[118] ,
		_w186_
	);
	LUT2 #(
		.INIT('h4)
	) name57 (
		_w185_,
		_w186_,
		_w187_
	);
	LUT4 #(
		.INIT('h000d)
	) name58 (
		\A[102] ,
		\A[103] ,
		\A[104] ,
		\A[106] ,
		_w188_
	);
	LUT4 #(
		.INIT('h000d)
	) name59 (
		\A[105] ,
		\A[106] ,
		\A[107] ,
		\A[109] ,
		_w189_
	);
	LUT2 #(
		.INIT('h4)
	) name60 (
		_w188_,
		_w189_,
		_w190_
	);
	LUT4 #(
		.INIT('h000d)
	) name61 (
		\A[93] ,
		\A[94] ,
		\A[95] ,
		\A[97] ,
		_w191_
	);
	LUT4 #(
		.INIT('h000d)
	) name62 (
		\A[96] ,
		\A[97] ,
		\A[98] ,
		\A[100] ,
		_w192_
	);
	LUT2 #(
		.INIT('h4)
	) name63 (
		_w191_,
		_w192_,
		_w193_
	);
	LUT4 #(
		.INIT('h00fb)
	) name64 (
		\A[85] ,
		\A[87] ,
		\A[88] ,
		\A[89] ,
		_w194_
	);
	LUT4 #(
		.INIT('h00a2)
	) name65 (
		\A[85] ,
		\A[86] ,
		\A[87] ,
		\A[88] ,
		_w195_
	);
	LUT3 #(
		.INIT('h04)
	) name66 (
		\A[91] ,
		_w194_,
		_w195_,
		_w196_
	);
	LUT4 #(
		.INIT('h000d)
	) name67 (
		\A[90] ,
		\A[91] ,
		\A[92] ,
		\A[94] ,
		_w197_
	);
	LUT2 #(
		.INIT('h8)
	) name68 (
		_w192_,
		_w197_,
		_w198_
	);
	LUT4 #(
		.INIT('h000d)
	) name69 (
		\A[99] ,
		\A[100] ,
		\A[101] ,
		\A[103] ,
		_w199_
	);
	LUT2 #(
		.INIT('h8)
	) name70 (
		_w189_,
		_w199_,
		_w200_
	);
	LUT4 #(
		.INIT('h4500)
	) name71 (
		_w193_,
		_w196_,
		_w198_,
		_w200_,
		_w201_
	);
	LUT4 #(
		.INIT('h000d)
	) name72 (
		\A[108] ,
		\A[109] ,
		\A[110] ,
		\A[112] ,
		_w202_
	);
	LUT2 #(
		.INIT('h8)
	) name73 (
		_w186_,
		_w202_,
		_w203_
	);
	LUT4 #(
		.INIT('h5455)
	) name74 (
		_w187_,
		_w190_,
		_w201_,
		_w203_,
		_w204_
	);
	LUT4 #(
		.INIT('h000d)
	) name75 (
		\A[117] ,
		\A[118] ,
		\A[119] ,
		\A[121] ,
		_w205_
	);
	LUT2 #(
		.INIT('h8)
	) name76 (
		_w183_,
		_w205_,
		_w206_
	);
	LUT4 #(
		.INIT('h0111)
	) name77 (
		_w181_,
		_w184_,
		_w204_,
		_w206_,
		_w207_
	);
	LUT4 #(
		.INIT('h000d)
	) name78 (
		\A[116] ,
		\A[117] ,
		\A[118] ,
		\A[120] ,
		_w208_
	);
	LUT4 #(
		.INIT('h000d)
	) name79 (
		\A[119] ,
		\A[120] ,
		\A[121] ,
		\A[123] ,
		_w209_
	);
	LUT2 #(
		.INIT('h4)
	) name80 (
		_w208_,
		_w209_,
		_w210_
	);
	LUT4 #(
		.INIT('h000d)
	) name81 (
		\A[107] ,
		\A[108] ,
		\A[109] ,
		\A[111] ,
		_w211_
	);
	LUT4 #(
		.INIT('h000d)
	) name82 (
		\A[110] ,
		\A[111] ,
		\A[112] ,
		\A[114] ,
		_w212_
	);
	LUT2 #(
		.INIT('h4)
	) name83 (
		_w211_,
		_w212_,
		_w213_
	);
	LUT2 #(
		.INIT('h2)
	) name84 (
		\A[98] ,
		\A[99] ,
		_w214_
	);
	LUT4 #(
		.INIT('h000d)
	) name85 (
		\A[95] ,
		\A[96] ,
		\A[97] ,
		\A[99] ,
		_w215_
	);
	LUT2 #(
		.INIT('h1)
	) name86 (
		\A[100] ,
		\A[102] ,
		_w216_
	);
	LUT2 #(
		.INIT('h4)
	) name87 (
		_w215_,
		_w216_,
		_w217_
	);
	LUT4 #(
		.INIT('h000d)
	) name88 (
		\A[86] ,
		\A[87] ,
		\A[88] ,
		\A[90] ,
		_w218_
	);
	LUT4 #(
		.INIT('h000d)
	) name89 (
		\A[89] ,
		\A[90] ,
		\A[91] ,
		\A[93] ,
		_w219_
	);
	LUT4 #(
		.INIT('h000d)
	) name90 (
		\A[92] ,
		\A[93] ,
		\A[94] ,
		\A[96] ,
		_w220_
	);
	LUT4 #(
		.INIT('h8a00)
	) name91 (
		_w216_,
		_w218_,
		_w219_,
		_w220_,
		_w221_
	);
	LUT4 #(
		.INIT('h000d)
	) name92 (
		\A[101] ,
		\A[102] ,
		\A[103] ,
		\A[105] ,
		_w222_
	);
	LUT4 #(
		.INIT('hab00)
	) name93 (
		_w214_,
		_w217_,
		_w221_,
		_w222_,
		_w223_
	);
	LUT4 #(
		.INIT('h000d)
	) name94 (
		\A[104] ,
		\A[105] ,
		\A[106] ,
		\A[108] ,
		_w224_
	);
	LUT2 #(
		.INIT('h8)
	) name95 (
		_w212_,
		_w224_,
		_w225_
	);
	LUT4 #(
		.INIT('h000d)
	) name96 (
		\A[113] ,
		\A[114] ,
		\A[115] ,
		\A[117] ,
		_w226_
	);
	LUT2 #(
		.INIT('h8)
	) name97 (
		_w209_,
		_w226_,
		_w227_
	);
	LUT4 #(
		.INIT('h4500)
	) name98 (
		_w213_,
		_w223_,
		_w225_,
		_w227_,
		_w228_
	);
	LUT4 #(
		.INIT('h000d)
	) name99 (
		\A[122] ,
		\A[123] ,
		\A[124] ,
		\A[126] ,
		_w229_
	);
	LUT3 #(
		.INIT('h0d)
	) name100 (
		\A[125] ,
		\A[126] ,
		\A[127] ,
		_w230_
	);
	LUT4 #(
		.INIT('hef00)
	) name101 (
		_w210_,
		_w228_,
		_w229_,
		_w230_,
		_w231_
	);
	LUT2 #(
		.INIT('h2)
	) name102 (
		_w179_,
		_w231_,
		_w232_
	);
	LUT4 #(
		.INIT('h4f00)
	) name103 (
		_w176_,
		_w177_,
		_w178_,
		_w232_,
		_w233_
	);
	LUT3 #(
		.INIT('hf4)
	) name104 (
		_w180_,
		_w207_,
		_w233_,
		_w234_
	);
	LUT2 #(
		.INIT('h1)
	) name105 (
		\A[124] ,
		\A[125] ,
		_w235_
	);
	LUT4 #(
		.INIT('h000e)
	) name106 (
		\A[118] ,
		\A[119] ,
		\A[120] ,
		\A[121] ,
		_w236_
	);
	LUT4 #(
		.INIT('h000e)
	) name107 (
		\A[112] ,
		\A[113] ,
		\A[114] ,
		\A[115] ,
		_w237_
	);
	LUT4 #(
		.INIT('h000e)
	) name108 (
		\A[106] ,
		\A[107] ,
		\A[108] ,
		\A[109] ,
		_w238_
	);
	LUT2 #(
		.INIT('h1)
	) name109 (
		\A[100] ,
		\A[101] ,
		_w239_
	);
	LUT4 #(
		.INIT('h000e)
	) name110 (
		\A[94] ,
		\A[95] ,
		\A[96] ,
		\A[97] ,
		_w240_
	);
	LUT2 #(
		.INIT('h1)
	) name111 (
		\A[84] ,
		\A[85] ,
		_w241_
	);
	LUT4 #(
		.INIT('h000e)
	) name112 (
		\A[82] ,
		\A[83] ,
		\A[88] ,
		\A[89] ,
		_w242_
	);
	LUT4 #(
		.INIT('h000e)
	) name113 (
		\A[76] ,
		\A[77] ,
		\A[78] ,
		\A[79] ,
		_w243_
	);
	LUT4 #(
		.INIT('h000e)
	) name114 (
		\A[70] ,
		\A[71] ,
		\A[72] ,
		\A[73] ,
		_w244_
	);
	LUT4 #(
		.INIT('h000e)
	) name115 (
		\A[64] ,
		\A[65] ,
		\A[66] ,
		\A[67] ,
		_w245_
	);
	LUT4 #(
		.INIT('h000e)
	) name116 (
		\A[58] ,
		\A[59] ,
		\A[60] ,
		\A[61] ,
		_w246_
	);
	LUT4 #(
		.INIT('h000e)
	) name117 (
		\A[52] ,
		\A[53] ,
		\A[54] ,
		\A[55] ,
		_w247_
	);
	LUT4 #(
		.INIT('h000e)
	) name118 (
		\A[26] ,
		\A[27] ,
		\A[28] ,
		\A[29] ,
		_w248_
	);
	LUT4 #(
		.INIT('h000e)
	) name119 (
		\A[20] ,
		\A[21] ,
		\A[22] ,
		\A[23] ,
		_w249_
	);
	LUT4 #(
		.INIT('h000e)
	) name120 (
		\A[14] ,
		\A[15] ,
		\A[16] ,
		\A[17] ,
		_w250_
	);
	LUT4 #(
		.INIT('h000e)
	) name121 (
		\A[8] ,
		\A[9] ,
		\A[10] ,
		\A[11] ,
		_w251_
	);
	LUT4 #(
		.INIT('h000e)
	) name122 (
		\A[2] ,
		\A[3] ,
		\A[4] ,
		\A[5] ,
		_w252_
	);
	LUT4 #(
		.INIT('h0001)
	) name123 (
		\A[6] ,
		\A[7] ,
		\A[10] ,
		\A[11] ,
		_w253_
	);
	LUT4 #(
		.INIT('h0001)
	) name124 (
		\A[12] ,
		\A[13] ,
		\A[16] ,
		\A[17] ,
		_w254_
	);
	LUT4 #(
		.INIT('h4500)
	) name125 (
		_w251_,
		_w252_,
		_w253_,
		_w254_,
		_w255_
	);
	LUT4 #(
		.INIT('h0001)
	) name126 (
		\A[18] ,
		\A[19] ,
		\A[22] ,
		\A[23] ,
		_w256_
	);
	LUT4 #(
		.INIT('h5455)
	) name127 (
		_w249_,
		_w250_,
		_w255_,
		_w256_,
		_w257_
	);
	LUT4 #(
		.INIT('h0001)
	) name128 (
		\A[24] ,
		\A[25] ,
		\A[28] ,
		\A[29] ,
		_w258_
	);
	LUT4 #(
		.INIT('h000e)
	) name129 (
		\A[34] ,
		\A[35] ,
		\A[36] ,
		\A[37] ,
		_w259_
	);
	LUT4 #(
		.INIT('h0001)
	) name130 (
		\A[38] ,
		\A[39] ,
		\A[42] ,
		\A[43] ,
		_w260_
	);
	LUT2 #(
		.INIT('h1)
	) name131 (
		\A[44] ,
		\A[45] ,
		_w261_
	);
	LUT4 #(
		.INIT('h000e)
	) name132 (
		\A[40] ,
		\A[41] ,
		\A[42] ,
		\A[43] ,
		_w262_
	);
	LUT4 #(
		.INIT('h00b0)
	) name133 (
		_w259_,
		_w260_,
		_w261_,
		_w262_,
		_w263_
	);
	LUT2 #(
		.INIT('h1)
	) name134 (
		\A[30] ,
		\A[31] ,
		_w264_
	);
	LUT4 #(
		.INIT('h0001)
	) name135 (
		\A[30] ,
		\A[31] ,
		\A[46] ,
		\A[47] ,
		_w265_
	);
	LUT2 #(
		.INIT('h4)
	) name136 (
		_w263_,
		_w265_,
		_w266_
	);
	LUT4 #(
		.INIT('h1500)
	) name137 (
		_w248_,
		_w257_,
		_w258_,
		_w266_,
		_w267_
	);
	LUT2 #(
		.INIT('h1)
	) name138 (
		\A[48] ,
		\A[49] ,
		_w268_
	);
	LUT4 #(
		.INIT('h000e)
	) name139 (
		\A[32] ,
		\A[33] ,
		\A[46] ,
		\A[47] ,
		_w269_
	);
	LUT3 #(
		.INIT('h8c)
	) name140 (
		_w263_,
		_w268_,
		_w269_,
		_w270_
	);
	LUT4 #(
		.INIT('h1500)
	) name141 (
		_w248_,
		_w257_,
		_w258_,
		_w264_,
		_w271_
	);
	LUT4 #(
		.INIT('h000e)
	) name142 (
		\A[36] ,
		\A[37] ,
		\A[38] ,
		\A[39] ,
		_w272_
	);
	LUT4 #(
		.INIT('h0001)
	) name143 (
		\A[40] ,
		\A[41] ,
		\A[44] ,
		\A[45] ,
		_w273_
	);
	LUT4 #(
		.INIT('h000e)
	) name144 (
		\A[42] ,
		\A[43] ,
		\A[44] ,
		\A[45] ,
		_w274_
	);
	LUT4 #(
		.INIT('h0001)
	) name145 (
		\A[32] ,
		\A[33] ,
		\A[46] ,
		\A[47] ,
		_w275_
	);
	LUT4 #(
		.INIT('h0b00)
	) name146 (
		_w272_,
		_w273_,
		_w274_,
		_w275_,
		_w276_
	);
	LUT4 #(
		.INIT('h4044)
	) name147 (
		_w267_,
		_w270_,
		_w271_,
		_w276_,
		_w277_
	);
	LUT4 #(
		.INIT('h0001)
	) name148 (
		\A[50] ,
		\A[51] ,
		\A[54] ,
		\A[55] ,
		_w278_
	);
	LUT4 #(
		.INIT('h0001)
	) name149 (
		\A[56] ,
		\A[57] ,
		\A[60] ,
		\A[61] ,
		_w279_
	);
	LUT4 #(
		.INIT('h4500)
	) name150 (
		_w247_,
		_w277_,
		_w278_,
		_w279_,
		_w280_
	);
	LUT4 #(
		.INIT('h0001)
	) name151 (
		\A[62] ,
		\A[63] ,
		\A[66] ,
		\A[67] ,
		_w281_
	);
	LUT4 #(
		.INIT('h5455)
	) name152 (
		_w245_,
		_w246_,
		_w280_,
		_w281_,
		_w282_
	);
	LUT4 #(
		.INIT('h0001)
	) name153 (
		\A[68] ,
		\A[69] ,
		\A[72] ,
		\A[73] ,
		_w283_
	);
	LUT4 #(
		.INIT('h0001)
	) name154 (
		\A[74] ,
		\A[75] ,
		\A[78] ,
		\A[79] ,
		_w284_
	);
	LUT4 #(
		.INIT('h1500)
	) name155 (
		_w244_,
		_w282_,
		_w283_,
		_w284_,
		_w285_
	);
	LUT4 #(
		.INIT('h0001)
	) name156 (
		\A[80] ,
		\A[81] ,
		\A[88] ,
		\A[89] ,
		_w286_
	);
	LUT4 #(
		.INIT('h5455)
	) name157 (
		_w242_,
		_w243_,
		_w285_,
		_w286_,
		_w287_
	);
	LUT4 #(
		.INIT('h000e)
	) name158 (
		\A[86] ,
		\A[87] ,
		\A[88] ,
		\A[89] ,
		_w288_
	);
	LUT2 #(
		.INIT('h1)
	) name159 (
		\A[90] ,
		\A[91] ,
		_w289_
	);
	LUT2 #(
		.INIT('h4)
	) name160 (
		_w288_,
		_w289_,
		_w290_
	);
	LUT4 #(
		.INIT('h0001)
	) name161 (
		\A[92] ,
		\A[93] ,
		\A[96] ,
		\A[97] ,
		_w291_
	);
	LUT4 #(
		.INIT('h2f00)
	) name162 (
		_w241_,
		_w287_,
		_w290_,
		_w291_,
		_w292_
	);
	LUT4 #(
		.INIT('h000e)
	) name163 (
		\A[98] ,
		\A[99] ,
		\A[100] ,
		\A[101] ,
		_w293_
	);
	LUT2 #(
		.INIT('h1)
	) name164 (
		\A[102] ,
		\A[103] ,
		_w294_
	);
	LUT2 #(
		.INIT('h4)
	) name165 (
		_w293_,
		_w294_,
		_w295_
	);
	LUT4 #(
		.INIT('h5700)
	) name166 (
		_w239_,
		_w240_,
		_w292_,
		_w295_,
		_w296_
	);
	LUT4 #(
		.INIT('h0001)
	) name167 (
		\A[104] ,
		\A[105] ,
		\A[108] ,
		\A[109] ,
		_w297_
	);
	LUT4 #(
		.INIT('h0001)
	) name168 (
		\A[110] ,
		\A[111] ,
		\A[114] ,
		\A[115] ,
		_w298_
	);
	LUT4 #(
		.INIT('h4500)
	) name169 (
		_w238_,
		_w296_,
		_w297_,
		_w298_,
		_w299_
	);
	LUT4 #(
		.INIT('h0001)
	) name170 (
		\A[116] ,
		\A[117] ,
		\A[120] ,
		\A[121] ,
		_w300_
	);
	LUT4 #(
		.INIT('h5455)
	) name171 (
		_w236_,
		_w237_,
		_w299_,
		_w300_,
		_w301_
	);
	LUT2 #(
		.INIT('h1)
	) name172 (
		\A[126] ,
		\A[127] ,
		_w302_
	);
	LUT4 #(
		.INIT('h000e)
	) name173 (
		\A[122] ,
		\A[123] ,
		\A[124] ,
		\A[125] ,
		_w303_
	);
	LUT2 #(
		.INIT('h2)
	) name174 (
		_w302_,
		_w303_,
		_w304_
	);
	LUT3 #(
		.INIT('h2f)
	) name175 (
		_w235_,
		_w301_,
		_w304_,
		_w305_
	);
	LUT4 #(
		.INIT('h0001)
	) name176 (
		\A[68] ,
		\A[69] ,
		\A[70] ,
		\A[71] ,
		_w306_
	);
	LUT4 #(
		.INIT('h0001)
	) name177 (
		\A[64] ,
		\A[65] ,
		\A[66] ,
		\A[67] ,
		_w307_
	);
	LUT2 #(
		.INIT('h2)
	) name178 (
		_w306_,
		_w307_,
		_w308_
	);
	LUT4 #(
		.INIT('h0001)
	) name179 (
		\A[56] ,
		\A[57] ,
		\A[58] ,
		\A[59] ,
		_w309_
	);
	LUT4 #(
		.INIT('h0001)
	) name180 (
		\A[52] ,
		\A[53] ,
		\A[54] ,
		\A[55] ,
		_w310_
	);
	LUT2 #(
		.INIT('h2)
	) name181 (
		_w309_,
		_w310_,
		_w311_
	);
	LUT4 #(
		.INIT('h0001)
	) name182 (
		\A[44] ,
		\A[45] ,
		\A[46] ,
		\A[47] ,
		_w312_
	);
	LUT4 #(
		.INIT('h0001)
	) name183 (
		\A[40] ,
		\A[41] ,
		\A[42] ,
		\A[43] ,
		_w313_
	);
	LUT2 #(
		.INIT('h2)
	) name184 (
		_w312_,
		_w313_,
		_w314_
	);
	LUT4 #(
		.INIT('h0001)
	) name185 (
		\A[32] ,
		\A[33] ,
		\A[34] ,
		\A[35] ,
		_w315_
	);
	LUT4 #(
		.INIT('h0001)
	) name186 (
		\A[28] ,
		\A[29] ,
		\A[30] ,
		\A[31] ,
		_w316_
	);
	LUT2 #(
		.INIT('h2)
	) name187 (
		_w315_,
		_w316_,
		_w317_
	);
	LUT4 #(
		.INIT('h0001)
	) name188 (
		\A[20] ,
		\A[21] ,
		\A[22] ,
		\A[23] ,
		_w318_
	);
	LUT4 #(
		.INIT('h0001)
	) name189 (
		\A[16] ,
		\A[17] ,
		\A[18] ,
		\A[19] ,
		_w319_
	);
	LUT2 #(
		.INIT('h2)
	) name190 (
		_w318_,
		_w319_,
		_w320_
	);
	LUT4 #(
		.INIT('h0001)
	) name191 (
		\A[8] ,
		\A[9] ,
		\A[10] ,
		\A[11] ,
		_w321_
	);
	LUT4 #(
		.INIT('h0001)
	) name192 (
		\A[4] ,
		\A[5] ,
		\A[6] ,
		\A[7] ,
		_w322_
	);
	LUT4 #(
		.INIT('h0001)
	) name193 (
		\A[12] ,
		\A[13] ,
		\A[14] ,
		\A[15] ,
		_w323_
	);
	LUT4 #(
		.INIT('ha200)
	) name194 (
		_w318_,
		_w321_,
		_w322_,
		_w323_,
		_w324_
	);
	LUT4 #(
		.INIT('h0001)
	) name195 (
		\A[24] ,
		\A[25] ,
		\A[26] ,
		\A[27] ,
		_w325_
	);
	LUT2 #(
		.INIT('h8)
	) name196 (
		_w315_,
		_w325_,
		_w326_
	);
	LUT4 #(
		.INIT('h5455)
	) name197 (
		_w317_,
		_w320_,
		_w324_,
		_w326_,
		_w327_
	);
	LUT4 #(
		.INIT('h0001)
	) name198 (
		\A[36] ,
		\A[37] ,
		\A[38] ,
		\A[39] ,
		_w328_
	);
	LUT2 #(
		.INIT('h8)
	) name199 (
		_w312_,
		_w328_,
		_w329_
	);
	LUT4 #(
		.INIT('h0001)
	) name200 (
		\A[48] ,
		\A[49] ,
		\A[50] ,
		\A[51] ,
		_w330_
	);
	LUT2 #(
		.INIT('h8)
	) name201 (
		_w309_,
		_w330_,
		_w331_
	);
	LUT4 #(
		.INIT('h1500)
	) name202 (
		_w314_,
		_w327_,
		_w329_,
		_w331_,
		_w332_
	);
	LUT4 #(
		.INIT('h0001)
	) name203 (
		\A[60] ,
		\A[61] ,
		\A[62] ,
		\A[63] ,
		_w333_
	);
	LUT2 #(
		.INIT('h8)
	) name204 (
		_w306_,
		_w333_,
		_w334_
	);
	LUT4 #(
		.INIT('h5455)
	) name205 (
		_w308_,
		_w311_,
		_w332_,
		_w334_,
		_w335_
	);
	LUT4 #(
		.INIT('h0001)
	) name206 (
		\A[72] ,
		\A[73] ,
		\A[74] ,
		\A[75] ,
		_w336_
	);
	LUT4 #(
		.INIT('h0001)
	) name207 (
		\A[84] ,
		\A[85] ,
		\A[86] ,
		\A[87] ,
		_w337_
	);
	LUT4 #(
		.INIT('h0001)
	) name208 (
		\A[88] ,
		\A[89] ,
		\A[90] ,
		\A[91] ,
		_w338_
	);
	LUT4 #(
		.INIT('h0001)
	) name209 (
		\A[92] ,
		\A[93] ,
		\A[94] ,
		\A[95] ,
		_w339_
	);
	LUT4 #(
		.INIT('h0001)
	) name210 (
		\A[100] ,
		\A[101] ,
		\A[102] ,
		\A[103] ,
		_w340_
	);
	LUT4 #(
		.INIT('hb000)
	) name211 (
		_w337_,
		_w338_,
		_w339_,
		_w340_,
		_w341_
	);
	LUT4 #(
		.INIT('h0001)
	) name212 (
		\A[104] ,
		\A[105] ,
		\A[106] ,
		\A[107] ,
		_w342_
	);
	LUT4 #(
		.INIT('h0001)
	) name213 (
		\A[112] ,
		\A[113] ,
		\A[114] ,
		\A[115] ,
		_w343_
	);
	LUT4 #(
		.INIT('h0001)
	) name214 (
		\A[96] ,
		\A[97] ,
		\A[98] ,
		\A[99] ,
		_w344_
	);
	LUT4 #(
		.INIT('hc040)
	) name215 (
		_w340_,
		_w342_,
		_w343_,
		_w344_,
		_w345_
	);
	LUT4 #(
		.INIT('h0001)
	) name216 (
		\A[76] ,
		\A[77] ,
		\A[78] ,
		\A[79] ,
		_w346_
	);
	LUT4 #(
		.INIT('h0001)
	) name217 (
		\A[116] ,
		\A[117] ,
		\A[118] ,
		\A[119] ,
		_w347_
	);
	LUT4 #(
		.INIT('h0001)
	) name218 (
		\A[108] ,
		\A[109] ,
		\A[110] ,
		\A[111] ,
		_w348_
	);
	LUT4 #(
		.INIT('hc040)
	) name219 (
		_w343_,
		_w346_,
		_w347_,
		_w348_,
		_w349_
	);
	LUT3 #(
		.INIT('hb0)
	) name220 (
		_w341_,
		_w345_,
		_w349_,
		_w350_
	);
	LUT3 #(
		.INIT('h70)
	) name221 (
		_w335_,
		_w336_,
		_w350_,
		_w351_
	);
	LUT2 #(
		.INIT('h4)
	) name222 (
		_w342_,
		_w348_,
		_w352_
	);
	LUT2 #(
		.INIT('h4)
	) name223 (
		_w339_,
		_w344_,
		_w353_
	);
	LUT4 #(
		.INIT('h0001)
	) name224 (
		\A[80] ,
		\A[81] ,
		\A[82] ,
		\A[83] ,
		_w354_
	);
	LUT4 #(
		.INIT('hc040)
	) name225 (
		_w337_,
		_w338_,
		_w344_,
		_w354_,
		_w355_
	);
	LUT2 #(
		.INIT('h8)
	) name226 (
		_w340_,
		_w348_,
		_w356_
	);
	LUT4 #(
		.INIT('h5455)
	) name227 (
		_w352_,
		_w353_,
		_w355_,
		_w356_,
		_w357_
	);
	LUT2 #(
		.INIT('h8)
	) name228 (
		_w336_,
		_w347_,
		_w358_
	);
	LUT3 #(
		.INIT('h70)
	) name229 (
		_w343_,
		_w357_,
		_w358_,
		_w359_
	);
	LUT4 #(
		.INIT('h0001)
	) name230 (
		\A[120] ,
		\A[121] ,
		\A[122] ,
		\A[123] ,
		_w360_
	);
	LUT2 #(
		.INIT('h4)
	) name231 (
		_w346_,
		_w347_,
		_w361_
	);
	LUT4 #(
		.INIT('h80f0)
	) name232 (
		_w343_,
		_w357_,
		_w360_,
		_w361_,
		_w362_
	);
	LUT3 #(
		.INIT('h70)
	) name233 (
		_w335_,
		_w359_,
		_w362_,
		_w363_
	);
	LUT4 #(
		.INIT('h0001)
	) name234 (
		\A[124] ,
		\A[125] ,
		\A[126] ,
		\A[127] ,
		_w364_
	);
	LUT3 #(
		.INIT('h4f)
	) name235 (
		_w351_,
		_w363_,
		_w364_,
		_w365_
	);
	LUT4 #(
		.INIT('h40c0)
	) name236 (
		_w337_,
		_w338_,
		_w339_,
		_w354_,
		_w366_
	);
	LUT4 #(
		.INIT('h0888)
	) name237 (
		_w306_,
		_w307_,
		_w309_,
		_w333_,
		_w367_
	);
	LUT4 #(
		.INIT('h0888)
	) name238 (
		_w312_,
		_w313_,
		_w315_,
		_w328_,
		_w368_
	);
	LUT4 #(
		.INIT('h0888)
	) name239 (
		_w318_,
		_w319_,
		_w321_,
		_w323_,
		_w369_
	);
	LUT4 #(
		.INIT('h8000)
	) name240 (
		_w312_,
		_w313_,
		_w316_,
		_w325_,
		_w370_
	);
	LUT4 #(
		.INIT('h8000)
	) name241 (
		_w306_,
		_w307_,
		_w310_,
		_w330_,
		_w371_
	);
	LUT4 #(
		.INIT('h4500)
	) name242 (
		_w368_,
		_w369_,
		_w370_,
		_w371_,
		_w372_
	);
	LUT4 #(
		.INIT('h8000)
	) name243 (
		_w336_,
		_w338_,
		_w339_,
		_w346_,
		_w373_
	);
	LUT4 #(
		.INIT('h5455)
	) name244 (
		_w366_,
		_w367_,
		_w372_,
		_w373_,
		_w374_
	);
	LUT2 #(
		.INIT('h8)
	) name245 (
		_w360_,
		_w364_,
		_w375_
	);
	LUT2 #(
		.INIT('h8)
	) name246 (
		_w343_,
		_w347_,
		_w376_
	);
	LUT4 #(
		.INIT('h4c00)
	) name247 (
		_w340_,
		_w342_,
		_w344_,
		_w348_,
		_w377_
	);
	LUT3 #(
		.INIT('ha2)
	) name248 (
		_w375_,
		_w376_,
		_w377_,
		_w378_
	);
	LUT4 #(
		.INIT('h40c0)
	) name249 (
		_w342_,
		_w343_,
		_w347_,
		_w348_,
		_w379_
	);
	LUT2 #(
		.INIT('h2)
	) name250 (
		_w375_,
		_w379_,
		_w380_
	);
	LUT3 #(
		.INIT('h27)
	) name251 (
		_w374_,
		_w378_,
		_w380_,
		_w381_
	);
	LUT4 #(
		.INIT('h8000)
	) name252 (
		_w343_,
		_w347_,
		_w360_,
		_w364_,
		_w382_
	);
	LUT4 #(
		.INIT('h8000)
	) name253 (
		_w337_,
		_w338_,
		_w339_,
		_w354_,
		_w383_
	);
	LUT4 #(
		.INIT('h8000)
	) name254 (
		_w306_,
		_w307_,
		_w336_,
		_w346_,
		_w384_
	);
	LUT2 #(
		.INIT('h2)
	) name255 (
		_w383_,
		_w384_,
		_w385_
	);
	LUT4 #(
		.INIT('h8000)
	) name256 (
		_w312_,
		_w313_,
		_w315_,
		_w328_,
		_w386_
	);
	LUT4 #(
		.INIT('h8000)
	) name257 (
		_w316_,
		_w318_,
		_w319_,
		_w325_,
		_w387_
	);
	LUT4 #(
		.INIT('h8000)
	) name258 (
		_w309_,
		_w310_,
		_w330_,
		_w333_,
		_w388_
	);
	LUT4 #(
		.INIT('ha200)
	) name259 (
		_w383_,
		_w386_,
		_w387_,
		_w388_,
		_w389_
	);
	LUT4 #(
		.INIT('h8000)
	) name260 (
		_w340_,
		_w342_,
		_w344_,
		_w348_,
		_w390_
	);
	LUT4 #(
		.INIT('h5755)
	) name261 (
		_w382_,
		_w385_,
		_w389_,
		_w390_,
		_w391_
	);
	LUT2 #(
		.INIT('h8)
	) name262 (
		_w382_,
		_w390_,
		_w392_
	);
	LUT4 #(
		.INIT('h0888)
	) name263 (
		_w383_,
		_w384_,
		_w386_,
		_w388_,
		_w393_
	);
	LUT2 #(
		.INIT('hd)
	) name264 (
		_w392_,
		_w393_,
		_w394_
	);
	LUT4 #(
		.INIT('h8000)
	) name265 (
		_w382_,
		_w383_,
		_w384_,
		_w390_,
		_w395_
	);
	LUT4 #(
		.INIT('h7fff)
	) name266 (
		_w382_,
		_w383_,
		_w384_,
		_w390_,
		_w396_
	);
	LUT4 #(
		.INIT('h0001)
	) name267 (
		\A[0] ,
		\A[1] ,
		\A[2] ,
		\A[3] ,
		_w397_
	);
	LUT4 #(
		.INIT('h8000)
	) name268 (
		_w321_,
		_w322_,
		_w323_,
		_w397_,
		_w398_
	);
	LUT4 #(
		.INIT('h8000)
	) name269 (
		_w386_,
		_w387_,
		_w388_,
		_w398_,
		_w399_
	);
	LUT2 #(
		.INIT('h7)
	) name270 (
		_w395_,
		_w399_,
		_w400_
	);
	assign \P[0]  = _w234_ ;
	assign \P[1]  = _w305_ ;
	assign \P[2]  = _w365_ ;
	assign \P[3]  = _w381_ ;
	assign \P[4]  = _w391_ ;
	assign \P[5]  = _w394_ ;
	assign \P[6]  = _w396_ ;
	assign F = _w400_ ;
endmodule;