module top (\IN_R_reg[0]/NET0131 , \IN_R_reg[1]/NET0131 , \IN_R_reg[2]/NET0131 , \IN_R_reg[3]/NET0131 , \IN_R_reg[4]/NET0131 , \IN_R_reg[5]/NET0131 , \IN_R_reg[6]/NET0131 , \IN_R_reg[7]/NET0131 , \I[0]_pad , \I[1]_pad , \I[2]_pad , \I[3]_pad , \I[4]_pad , \I[5]_pad , \I[6]_pad , \I[7]_pad , \MAR_reg[0]/NET0131 , \MAR_reg[1]/NET0131 , \MAR_reg[2]/NET0131 , \OUT_R_reg[0]/NET0131 , \OUT_R_reg[1]/NET0131 , \OUT_R_reg[2]/NET0131 , \OUT_R_reg[3]/NET0131 , \O[0]_pad , \O[1]_pad , \O[2]_pad , \O[3]_pad , START_pad, \STATO_reg[0]/NET0131 , \STATO_reg[1]/NET0131 , \_al_n0 , \_al_n1 , \g1016/_0_ , \g1017/_0_ , \g1018/_0_ , \g1019/_0_ , \g1041/_0_ , \g1052/_0_ , \g1053/_0_ , \g1054/_0_ , \g1058/_0_ , \g1059/_0_ , \g1060/_0_ , \g1061/_0_ , \g1063/_0_ , \g1090/_0_ , \g1093/_0_ , \g1095/_0_ , \g1098/_0_ , \g1099/_0_ , \g1100/_0_ , \g1101/_0_ , \g1102/_0_ );
	input \IN_R_reg[0]/NET0131  ;
	input \IN_R_reg[1]/NET0131  ;
	input \IN_R_reg[2]/NET0131  ;
	input \IN_R_reg[3]/NET0131  ;
	input \IN_R_reg[4]/NET0131  ;
	input \IN_R_reg[5]/NET0131  ;
	input \IN_R_reg[6]/NET0131  ;
	input \IN_R_reg[7]/NET0131  ;
	input \I[0]_pad  ;
	input \I[1]_pad  ;
	input \I[2]_pad  ;
	input \I[3]_pad  ;
	input \I[4]_pad  ;
	input \I[5]_pad  ;
	input \I[6]_pad  ;
	input \I[7]_pad  ;
	input \MAR_reg[0]/NET0131  ;
	input \MAR_reg[1]/NET0131  ;
	input \MAR_reg[2]/NET0131  ;
	input \OUT_R_reg[0]/NET0131  ;
	input \OUT_R_reg[1]/NET0131  ;
	input \OUT_R_reg[2]/NET0131  ;
	input \OUT_R_reg[3]/NET0131  ;
	input \O[0]_pad  ;
	input \O[1]_pad  ;
	input \O[2]_pad  ;
	input \O[3]_pad  ;
	input START_pad ;
	input \STATO_reg[0]/NET0131  ;
	input \STATO_reg[1]/NET0131  ;
	output \_al_n0  ;
	output \_al_n1  ;
	output \g1016/_0_  ;
	output \g1017/_0_  ;
	output \g1018/_0_  ;
	output \g1019/_0_  ;
	output \g1041/_0_  ;
	output \g1052/_0_  ;
	output \g1053/_0_  ;
	output \g1054/_0_  ;
	output \g1058/_0_  ;
	output \g1059/_0_  ;
	output \g1060/_0_  ;
	output \g1061/_0_  ;
	output \g1063/_0_  ;
	output \g1090/_0_  ;
	output \g1093/_0_  ;
	output \g1095/_0_  ;
	output \g1098/_0_  ;
	output \g1099/_0_  ;
	output \g1100/_0_  ;
	output \g1101/_0_  ;
	output \g1102/_0_  ;
	wire _w167_ ;
	wire _w166_ ;
	wire _w165_ ;
	wire _w164_ ;
	wire _w163_ ;
	wire _w162_ ;
	wire _w161_ ;
	wire _w160_ ;
	wire _w159_ ;
	wire _w158_ ;
	wire _w89_ ;
	wire _w88_ ;
	wire _w87_ ;
	wire _w86_ ;
	wire _w85_ ;
	wire _w84_ ;
	wire _w83_ ;
	wire _w82_ ;
	wire _w81_ ;
	wire _w80_ ;
	wire _w79_ ;
	wire _w78_ ;
	wire _w77_ ;
	wire _w76_ ;
	wire _w75_ ;
	wire _w74_ ;
	wire _w73_ ;
	wire _w72_ ;
	wire _w71_ ;
	wire _w70_ ;
	wire _w69_ ;
	wire _w68_ ;
	wire _w67_ ;
	wire _w66_ ;
	wire _w65_ ;
	wire _w64_ ;
	wire _w63_ ;
	wire _w62_ ;
	wire _w61_ ;
	wire _w60_ ;
	wire _w43_ ;
	wire _w42_ ;
	wire _w41_ ;
	wire _w40_ ;
	wire _w39_ ;
	wire _w38_ ;
	wire _w37_ ;
	wire _w36_ ;
	wire _w35_ ;
	wire _w34_ ;
	wire _w33_ ;
	wire _w32_ ;
	wire _w31_ ;
	wire _w44_ ;
	wire _w45_ ;
	wire _w46_ ;
	wire _w47_ ;
	wire _w48_ ;
	wire _w49_ ;
	wire _w50_ ;
	wire _w51_ ;
	wire _w52_ ;
	wire _w53_ ;
	wire _w54_ ;
	wire _w55_ ;
	wire _w56_ ;
	wire _w57_ ;
	wire _w58_ ;
	wire _w59_ ;
	wire _w90_ ;
	wire _w91_ ;
	wire _w92_ ;
	wire _w93_ ;
	wire _w94_ ;
	wire _w95_ ;
	wire _w96_ ;
	wire _w97_ ;
	wire _w98_ ;
	wire _w99_ ;
	wire _w100_ ;
	wire _w101_ ;
	wire _w102_ ;
	wire _w103_ ;
	wire _w104_ ;
	wire _w105_ ;
	wire _w106_ ;
	wire _w107_ ;
	wire _w108_ ;
	wire _w109_ ;
	wire _w110_ ;
	wire _w111_ ;
	wire _w112_ ;
	wire _w113_ ;
	wire _w114_ ;
	wire _w115_ ;
	wire _w116_ ;
	wire _w117_ ;
	wire _w118_ ;
	wire _w119_ ;
	wire _w120_ ;
	wire _w121_ ;
	wire _w122_ ;
	wire _w123_ ;
	wire _w124_ ;
	wire _w125_ ;
	wire _w126_ ;
	wire _w127_ ;
	wire _w128_ ;
	wire _w129_ ;
	wire _w130_ ;
	wire _w131_ ;
	wire _w132_ ;
	wire _w133_ ;
	wire _w134_ ;
	wire _w135_ ;
	wire _w136_ ;
	wire _w137_ ;
	wire _w138_ ;
	wire _w139_ ;
	wire _w140_ ;
	wire _w141_ ;
	wire _w142_ ;
	wire _w143_ ;
	wire _w144_ ;
	wire _w145_ ;
	wire _w146_ ;
	wire _w147_ ;
	wire _w148_ ;
	wire _w149_ ;
	wire _w150_ ;
	wire _w151_ ;
	wire _w152_ ;
	wire _w153_ ;
	wire _w154_ ;
	wire _w155_ ;
	wire _w156_ ;
	wire _w157_ ;
	LUT2 #(
		.INIT('h4)
	) name0 (
		\STATO_reg[0]/NET0131 ,
		\STATO_reg[1]/NET0131 ,
		_w31_
	);
	LUT2 #(
		.INIT('h2)
	) name1 (
		\STATO_reg[0]/NET0131 ,
		\STATO_reg[1]/NET0131 ,
		_w32_
	);
	LUT2 #(
		.INIT('h1)
	) name2 (
		_w31_,
		_w32_,
		_w33_
	);
	LUT2 #(
		.INIT('h4)
	) name3 (
		\MAR_reg[0]/NET0131 ,
		\MAR_reg[2]/NET0131 ,
		_w34_
	);
	LUT2 #(
		.INIT('h2)
	) name4 (
		\MAR_reg[0]/NET0131 ,
		\MAR_reg[2]/NET0131 ,
		_w35_
	);
	LUT2 #(
		.INIT('h1)
	) name5 (
		\MAR_reg[1]/NET0131 ,
		_w35_,
		_w36_
	);
	LUT2 #(
		.INIT('h4)
	) name6 (
		\IN_R_reg[6]/NET0131 ,
		_w36_,
		_w37_
	);
	LUT2 #(
		.INIT('h2)
	) name7 (
		\MAR_reg[1]/NET0131 ,
		\MAR_reg[2]/NET0131 ,
		_w38_
	);
	LUT2 #(
		.INIT('h4)
	) name8 (
		\MAR_reg[1]/NET0131 ,
		\MAR_reg[2]/NET0131 ,
		_w39_
	);
	LUT2 #(
		.INIT('h1)
	) name9 (
		_w38_,
		_w39_,
		_w40_
	);
	LUT2 #(
		.INIT('h8)
	) name10 (
		\IN_R_reg[7]/NET0131 ,
		_w40_,
		_w41_
	);
	LUT2 #(
		.INIT('h8)
	) name11 (
		\MAR_reg[0]/NET0131 ,
		_w38_,
		_w42_
	);
	LUT2 #(
		.INIT('h2)
	) name12 (
		\IN_R_reg[6]/NET0131 ,
		_w36_,
		_w43_
	);
	LUT2 #(
		.INIT('h4)
	) name13 (
		_w42_,
		_w43_,
		_w44_
	);
	LUT2 #(
		.INIT('h1)
	) name14 (
		_w37_,
		_w41_,
		_w45_
	);
	LUT2 #(
		.INIT('h4)
	) name15 (
		_w44_,
		_w45_,
		_w46_
	);
	LUT2 #(
		.INIT('h1)
	) name16 (
		_w34_,
		_w46_,
		_w47_
	);
	LUT2 #(
		.INIT('h8)
	) name17 (
		\IN_R_reg[5]/NET0131 ,
		\MAR_reg[2]/NET0131 ,
		_w48_
	);
	LUT2 #(
		.INIT('h1)
	) name18 (
		\IN_R_reg[0]/NET0131 ,
		_w48_,
		_w49_
	);
	LUT2 #(
		.INIT('h1)
	) name19 (
		\MAR_reg[0]/NET0131 ,
		_w49_,
		_w50_
	);
	LUT2 #(
		.INIT('h2)
	) name20 (
		\IN_R_reg[4]/NET0131 ,
		_w35_,
		_w51_
	);
	LUT2 #(
		.INIT('h4)
	) name21 (
		\IN_R_reg[4]/NET0131 ,
		_w35_,
		_w52_
	);
	LUT2 #(
		.INIT('h1)
	) name22 (
		_w51_,
		_w52_,
		_w53_
	);
	LUT2 #(
		.INIT('h4)
	) name23 (
		_w50_,
		_w53_,
		_w54_
	);
	LUT2 #(
		.INIT('h2)
	) name24 (
		\MAR_reg[1]/NET0131 ,
		_w54_,
		_w55_
	);
	LUT2 #(
		.INIT('h4)
	) name25 (
		\IN_R_reg[2]/NET0131 ,
		\MAR_reg[0]/NET0131 ,
		_w56_
	);
	LUT2 #(
		.INIT('h4)
	) name26 (
		_w40_,
		_w56_,
		_w57_
	);
	LUT2 #(
		.INIT('h8)
	) name27 (
		\MAR_reg[0]/NET0131 ,
		\MAR_reg[1]/NET0131 ,
		_w58_
	);
	LUT2 #(
		.INIT('h1)
	) name28 (
		\MAR_reg[0]/NET0131 ,
		\MAR_reg[1]/NET0131 ,
		_w59_
	);
	LUT2 #(
		.INIT('h1)
	) name29 (
		_w58_,
		_w59_,
		_w60_
	);
	LUT2 #(
		.INIT('h8)
	) name30 (
		\MAR_reg[0]/NET0131 ,
		\MAR_reg[2]/NET0131 ,
		_w61_
	);
	LUT2 #(
		.INIT('h2)
	) name31 (
		\IN_R_reg[2]/NET0131 ,
		_w61_,
		_w62_
	);
	LUT2 #(
		.INIT('h8)
	) name32 (
		_w60_,
		_w62_,
		_w63_
	);
	LUT2 #(
		.INIT('h8)
	) name33 (
		\IN_R_reg[1]/NET0131 ,
		\MAR_reg[2]/NET0131 ,
		_w64_
	);
	LUT2 #(
		.INIT('h8)
	) name34 (
		\MAR_reg[1]/NET0131 ,
		\MAR_reg[2]/NET0131 ,
		_w65_
	);
	LUT2 #(
		.INIT('h1)
	) name35 (
		\IN_R_reg[1]/NET0131 ,
		_w65_,
		_w66_
	);
	LUT2 #(
		.INIT('h2)
	) name36 (
		_w60_,
		_w64_,
		_w67_
	);
	LUT2 #(
		.INIT('h4)
	) name37 (
		_w66_,
		_w67_,
		_w68_
	);
	LUT2 #(
		.INIT('h1)
	) name38 (
		\IN_R_reg[3]/NET0131 ,
		_w38_,
		_w69_
	);
	LUT2 #(
		.INIT('h1)
	) name39 (
		\MAR_reg[0]/NET0131 ,
		\MAR_reg[2]/NET0131 ,
		_w70_
	);
	LUT2 #(
		.INIT('h4)
	) name40 (
		\IN_R_reg[7]/NET0131 ,
		\MAR_reg[1]/NET0131 ,
		_w71_
	);
	LUT2 #(
		.INIT('h4)
	) name41 (
		_w70_,
		_w71_,
		_w72_
	);
	LUT2 #(
		.INIT('h1)
	) name42 (
		_w69_,
		_w72_,
		_w73_
	);
	LUT2 #(
		.INIT('h1)
	) name43 (
		_w61_,
		_w73_,
		_w74_
	);
	LUT2 #(
		.INIT('h1)
	) name44 (
		\IN_R_reg[5]/NET0131 ,
		\MAR_reg[2]/NET0131 ,
		_w75_
	);
	LUT2 #(
		.INIT('h1)
	) name45 (
		\IN_R_reg[0]/NET0131 ,
		_w70_,
		_w76_
	);
	LUT2 #(
		.INIT('h1)
	) name46 (
		_w75_,
		_w76_,
		_w77_
	);
	LUT2 #(
		.INIT('h1)
	) name47 (
		\MAR_reg[1]/NET0131 ,
		_w77_,
		_w78_
	);
	LUT2 #(
		.INIT('h1)
	) name48 (
		_w57_,
		_w63_,
		_w79_
	);
	LUT2 #(
		.INIT('h4)
	) name49 (
		_w68_,
		_w79_,
		_w80_
	);
	LUT2 #(
		.INIT('h1)
	) name50 (
		_w74_,
		_w78_,
		_w81_
	);
	LUT2 #(
		.INIT('h8)
	) name51 (
		_w80_,
		_w81_,
		_w82_
	);
	LUT2 #(
		.INIT('h4)
	) name52 (
		_w55_,
		_w82_,
		_w83_
	);
	LUT2 #(
		.INIT('h4)
	) name53 (
		_w47_,
		_w83_,
		_w84_
	);
	LUT2 #(
		.INIT('h2)
	) name54 (
		\STATO_reg[1]/NET0131 ,
		_w84_,
		_w85_
	);
	LUT2 #(
		.INIT('h1)
	) name55 (
		_w33_,
		_w85_,
		_w86_
	);
	LUT2 #(
		.INIT('h2)
	) name56 (
		\OUT_R_reg[3]/NET0131 ,
		_w86_,
		_w87_
	);
	LUT2 #(
		.INIT('h2)
	) name57 (
		\MAR_reg[0]/NET0131 ,
		\OUT_R_reg[3]/NET0131 ,
		_w88_
	);
	LUT2 #(
		.INIT('h8)
	) name58 (
		_w40_,
		_w88_,
		_w89_
	);
	LUT2 #(
		.INIT('h2)
	) name59 (
		_w31_,
		_w89_,
		_w90_
	);
	LUT2 #(
		.INIT('h8)
	) name60 (
		_w84_,
		_w90_,
		_w91_
	);
	LUT2 #(
		.INIT('h1)
	) name61 (
		_w87_,
		_w91_,
		_w92_
	);
	LUT2 #(
		.INIT('h2)
	) name62 (
		\OUT_R_reg[1]/NET0131 ,
		_w86_,
		_w93_
	);
	LUT2 #(
		.INIT('h4)
	) name63 (
		\OUT_R_reg[1]/NET0131 ,
		_w61_,
		_w94_
	);
	LUT2 #(
		.INIT('h2)
	) name64 (
		_w31_,
		_w94_,
		_w95_
	);
	LUT2 #(
		.INIT('h8)
	) name65 (
		_w84_,
		_w95_,
		_w96_
	);
	LUT2 #(
		.INIT('h1)
	) name66 (
		_w93_,
		_w96_,
		_w97_
	);
	LUT2 #(
		.INIT('h2)
	) name67 (
		\OUT_R_reg[0]/NET0131 ,
		_w86_,
		_w98_
	);
	LUT2 #(
		.INIT('h4)
	) name68 (
		\MAR_reg[0]/NET0131 ,
		\MAR_reg[1]/NET0131 ,
		_w99_
	);
	LUT2 #(
		.INIT('h1)
	) name69 (
		\OUT_R_reg[0]/NET0131 ,
		_w99_,
		_w100_
	);
	LUT2 #(
		.INIT('h2)
	) name70 (
		_w31_,
		_w100_,
		_w101_
	);
	LUT2 #(
		.INIT('h8)
	) name71 (
		_w84_,
		_w101_,
		_w102_
	);
	LUT2 #(
		.INIT('h1)
	) name72 (
		_w98_,
		_w102_,
		_w103_
	);
	LUT2 #(
		.INIT('h2)
	) name73 (
		\OUT_R_reg[2]/NET0131 ,
		_w86_,
		_w104_
	);
	LUT2 #(
		.INIT('h8)
	) name74 (
		\MAR_reg[1]/NET0131 ,
		_w61_,
		_w105_
	);
	LUT2 #(
		.INIT('h1)
	) name75 (
		\MAR_reg[0]/NET0131 ,
		_w40_,
		_w106_
	);
	LUT2 #(
		.INIT('h1)
	) name76 (
		\OUT_R_reg[2]/NET0131 ,
		_w105_,
		_w107_
	);
	LUT2 #(
		.INIT('h4)
	) name77 (
		_w106_,
		_w107_,
		_w108_
	);
	LUT2 #(
		.INIT('h2)
	) name78 (
		_w31_,
		_w108_,
		_w109_
	);
	LUT2 #(
		.INIT('h8)
	) name79 (
		_w84_,
		_w109_,
		_w110_
	);
	LUT2 #(
		.INIT('h1)
	) name80 (
		_w104_,
		_w110_,
		_w111_
	);
	LUT2 #(
		.INIT('h8)
	) name81 (
		\STATO_reg[0]/NET0131 ,
		_w58_,
		_w112_
	);
	LUT2 #(
		.INIT('h1)
	) name82 (
		\MAR_reg[2]/NET0131 ,
		_w112_,
		_w113_
	);
	LUT2 #(
		.INIT('h1)
	) name83 (
		_w32_,
		_w113_,
		_w114_
	);
	LUT2 #(
		.INIT('h2)
	) name84 (
		\MAR_reg[1]/NET0131 ,
		\STATO_reg[0]/NET0131 ,
		_w115_
	);
	LUT2 #(
		.INIT('h8)
	) name85 (
		\STATO_reg[0]/NET0131 ,
		\STATO_reg[1]/NET0131 ,
		_w116_
	);
	LUT2 #(
		.INIT('h4)
	) name86 (
		_w59_,
		_w116_,
		_w117_
	);
	LUT2 #(
		.INIT('h4)
	) name87 (
		_w42_,
		_w117_,
		_w118_
	);
	LUT2 #(
		.INIT('h1)
	) name88 (
		_w115_,
		_w118_,
		_w119_
	);
	LUT2 #(
		.INIT('h8)
	) name89 (
		\STATO_reg[1]/NET0131 ,
		_w105_,
		_w120_
	);
	LUT2 #(
		.INIT('h2)
	) name90 (
		\STATO_reg[0]/NET0131 ,
		_w120_,
		_w121_
	);
	LUT2 #(
		.INIT('h1)
	) name91 (
		START_pad,
		_w31_,
		_w122_
	);
	LUT2 #(
		.INIT('h1)
	) name92 (
		_w121_,
		_w122_,
		_w123_
	);
	LUT2 #(
		.INIT('h4)
	) name93 (
		START_pad,
		_w105_,
		_w124_
	);
	LUT2 #(
		.INIT('h2)
	) name94 (
		_w116_,
		_w124_,
		_w125_
	);
	LUT2 #(
		.INIT('h2)
	) name95 (
		_w33_,
		_w125_,
		_w126_
	);
	LUT2 #(
		.INIT('h8)
	) name96 (
		_w116_,
		_w124_,
		_w127_
	);
	LUT2 #(
		.INIT('h2)
	) name97 (
		\O[0]_pad ,
		_w127_,
		_w128_
	);
	LUT2 #(
		.INIT('h8)
	) name98 (
		\OUT_R_reg[0]/NET0131 ,
		_w127_,
		_w129_
	);
	LUT2 #(
		.INIT('h1)
	) name99 (
		_w128_,
		_w129_,
		_w130_
	);
	LUT2 #(
		.INIT('h2)
	) name100 (
		\O[1]_pad ,
		_w127_,
		_w131_
	);
	LUT2 #(
		.INIT('h8)
	) name101 (
		\OUT_R_reg[1]/NET0131 ,
		_w127_,
		_w132_
	);
	LUT2 #(
		.INIT('h1)
	) name102 (
		_w131_,
		_w132_,
		_w133_
	);
	LUT2 #(
		.INIT('h2)
	) name103 (
		\O[2]_pad ,
		_w127_,
		_w134_
	);
	LUT2 #(
		.INIT('h8)
	) name104 (
		\OUT_R_reg[2]/NET0131 ,
		_w127_,
		_w135_
	);
	LUT2 #(
		.INIT('h1)
	) name105 (
		_w134_,
		_w135_,
		_w136_
	);
	LUT2 #(
		.INIT('h2)
	) name106 (
		\O[3]_pad ,
		_w127_,
		_w137_
	);
	LUT2 #(
		.INIT('h8)
	) name107 (
		\OUT_R_reg[3]/NET0131 ,
		_w127_,
		_w138_
	);
	LUT2 #(
		.INIT('h1)
	) name108 (
		_w137_,
		_w138_,
		_w139_
	);
	LUT2 #(
		.INIT('h2)
	) name109 (
		\MAR_reg[0]/NET0131 ,
		\STATO_reg[0]/NET0131 ,
		_w140_
	);
	LUT2 #(
		.INIT('h2)
	) name110 (
		\MAR_reg[0]/NET0131 ,
		_w65_,
		_w141_
	);
	LUT2 #(
		.INIT('h2)
	) name111 (
		_w116_,
		_w141_,
		_w142_
	);
	LUT2 #(
		.INIT('h1)
	) name112 (
		_w140_,
		_w142_,
		_w143_
	);
	LUT2 #(
		.INIT('h2)
	) name113 (
		\IN_R_reg[2]/NET0131 ,
		_w32_,
		_w144_
	);
	LUT2 #(
		.INIT('h8)
	) name114 (
		\I[2]_pad ,
		_w32_,
		_w145_
	);
	LUT2 #(
		.INIT('h1)
	) name115 (
		_w144_,
		_w145_,
		_w146_
	);
	LUT2 #(
		.INIT('h2)
	) name116 (
		\IN_R_reg[6]/NET0131 ,
		_w32_,
		_w147_
	);
	LUT2 #(
		.INIT('h8)
	) name117 (
		\I[6]_pad ,
		_w32_,
		_w148_
	);
	LUT2 #(
		.INIT('h1)
	) name118 (
		_w147_,
		_w148_,
		_w149_
	);
	LUT2 #(
		.INIT('h2)
	) name119 (
		\IN_R_reg[7]/NET0131 ,
		_w32_,
		_w150_
	);
	LUT2 #(
		.INIT('h8)
	) name120 (
		\I[7]_pad ,
		_w32_,
		_w151_
	);
	LUT2 #(
		.INIT('h1)
	) name121 (
		_w150_,
		_w151_,
		_w152_
	);
	LUT2 #(
		.INIT('h2)
	) name122 (
		\IN_R_reg[3]/NET0131 ,
		_w32_,
		_w153_
	);
	LUT2 #(
		.INIT('h8)
	) name123 (
		\I[3]_pad ,
		_w32_,
		_w154_
	);
	LUT2 #(
		.INIT('h1)
	) name124 (
		_w153_,
		_w154_,
		_w155_
	);
	LUT2 #(
		.INIT('h2)
	) name125 (
		\IN_R_reg[0]/NET0131 ,
		_w32_,
		_w156_
	);
	LUT2 #(
		.INIT('h8)
	) name126 (
		\I[0]_pad ,
		_w32_,
		_w157_
	);
	LUT2 #(
		.INIT('h1)
	) name127 (
		_w156_,
		_w157_,
		_w158_
	);
	LUT2 #(
		.INIT('h2)
	) name128 (
		\IN_R_reg[4]/NET0131 ,
		_w32_,
		_w159_
	);
	LUT2 #(
		.INIT('h8)
	) name129 (
		\I[4]_pad ,
		_w32_,
		_w160_
	);
	LUT2 #(
		.INIT('h1)
	) name130 (
		_w159_,
		_w160_,
		_w161_
	);
	LUT2 #(
		.INIT('h2)
	) name131 (
		\IN_R_reg[5]/NET0131 ,
		_w32_,
		_w162_
	);
	LUT2 #(
		.INIT('h8)
	) name132 (
		\I[5]_pad ,
		_w32_,
		_w163_
	);
	LUT2 #(
		.INIT('h1)
	) name133 (
		_w162_,
		_w163_,
		_w164_
	);
	LUT2 #(
		.INIT('h2)
	) name134 (
		\IN_R_reg[1]/NET0131 ,
		_w32_,
		_w165_
	);
	LUT2 #(
		.INIT('h8)
	) name135 (
		\I[1]_pad ,
		_w32_,
		_w166_
	);
	LUT2 #(
		.INIT('h1)
	) name136 (
		_w165_,
		_w166_,
		_w167_
	);
	assign \_al_n0  = 1'b0;
	assign \_al_n1  = 1'b0;
	assign \g1016/_0_  = _w92_ ;
	assign \g1017/_0_  = _w97_ ;
	assign \g1018/_0_  = _w103_ ;
	assign \g1019/_0_  = _w111_ ;
	assign \g1041/_0_  = _w114_ ;
	assign \g1052/_0_  = _w119_ ;
	assign \g1053/_0_  = _w123_ ;
	assign \g1054/_0_  = _w126_ ;
	assign \g1058/_0_  = _w130_ ;
	assign \g1059/_0_  = _w133_ ;
	assign \g1060/_0_  = _w136_ ;
	assign \g1061/_0_  = _w139_ ;
	assign \g1063/_0_  = _w143_ ;
	assign \g1090/_0_  = _w146_ ;
	assign \g1093/_0_  = _w149_ ;
	assign \g1095/_0_  = _w152_ ;
	assign \g1098/_0_  = _w155_ ;
	assign \g1099/_0_  = _w158_ ;
	assign \g1100/_0_  = _w161_ ;
	assign \g1101/_0_  = _w164_ ;
	assign \g1102/_0_  = _w167_ ;
endmodule;