module top( \101GAT(25)_pad  , \106GAT(26)_pad  , \111GAT(27)_pad  , \116GAT(28)_pad  , \121GAT(29)_pad  , \126GAT(30)_pad  , \130GAT(31)_pad  , \135GAT(32)_pad  , \138GAT(33)_pad  , \13GAT(2)_pad  , \143GAT(34)_pad  , \146GAT(35)_pad  , \149GAT(36)_pad  , \152GAT(37)_pad  , \153GAT(38)_pad  , \156GAT(39)_pad  , \159GAT(40)_pad  , \165GAT(41)_pad  , \171GAT(42)_pad  , \177GAT(43)_pad  , \17GAT(3)_pad  , \183GAT(44)_pad  , \189GAT(45)_pad  , \195GAT(46)_pad  , \1GAT(0)_pad  , \201GAT(47)_pad  , \207GAT(48)_pad  , \210GAT(49)_pad  , \219GAT(50)_pad  , \228GAT(51)_pad  , \237GAT(52)_pad  , \246GAT(53)_pad  , \255GAT(54)_pad  , \259GAT(55)_pad  , \260GAT(56)_pad  , \261GAT(57)_pad  , \267GAT(58)_pad  , \268GAT(59)_pad  , \26GAT(4)_pad  , \29GAT(5)_pad  , \36GAT(6)_pad  , \42GAT(7)_pad  , \51GAT(8)_pad  , \55GAT(9)_pad  , \59GAT(10)_pad  , \68GAT(11)_pad  , \72GAT(12)_pad  , \73GAT(13)_pad  , \74GAT(14)_pad  , \75GAT(15)_pad  , \80GAT(16)_pad  , \85GAT(17)_pad  , \86GAT(18)_pad  , \87GAT(19)_pad  , \88GAT(20)_pad  , \89GAT(21)_pad  , \8GAT(1)_pad  , \90GAT(22)_pad  , \91GAT(23)_pad  , \96GAT(24)_pad  , \273GAT(103)  , \388GAT(133)_pad  , \389GAT(132)_pad  , \391GAT(124)_pad  , \393GAT(165)  , \418GAT(168)_pad  , \419GAT(164)_pad  , \420GAT(158)_pad  , \421GAT(162)_pad  , \422GAT(161)_pad  , \423GAT(155)_pad  , \446GAT(183)_pad  , \448GAT(179)_pad  , \449GAT(176)_pad  , \450GAT(173)_pad  , \767GAT(349)_pad  , \768GAT(334)_pad  , \811GAT(378)  , \837GAT(396)  , \838GAT(395)  , \839GAT(394)  , \854GAT(419)  , \866GAT(426)_pad  , \867GAT(432)  , \868GAT(431)  , \869GAT(430)  );
  input \101GAT(25)_pad  ;
  input \106GAT(26)_pad  ;
  input \111GAT(27)_pad  ;
  input \116GAT(28)_pad  ;
  input \121GAT(29)_pad  ;
  input \126GAT(30)_pad  ;
  input \130GAT(31)_pad  ;
  input \135GAT(32)_pad  ;
  input \138GAT(33)_pad  ;
  input \13GAT(2)_pad  ;
  input \143GAT(34)_pad  ;
  input \146GAT(35)_pad  ;
  input \149GAT(36)_pad  ;
  input \152GAT(37)_pad  ;
  input \153GAT(38)_pad  ;
  input \156GAT(39)_pad  ;
  input \159GAT(40)_pad  ;
  input \165GAT(41)_pad  ;
  input \171GAT(42)_pad  ;
  input \177GAT(43)_pad  ;
  input \17GAT(3)_pad  ;
  input \183GAT(44)_pad  ;
  input \189GAT(45)_pad  ;
  input \195GAT(46)_pad  ;
  input \1GAT(0)_pad  ;
  input \201GAT(47)_pad  ;
  input \207GAT(48)_pad  ;
  input \210GAT(49)_pad  ;
  input \219GAT(50)_pad  ;
  input \228GAT(51)_pad  ;
  input \237GAT(52)_pad  ;
  input \246GAT(53)_pad  ;
  input \255GAT(54)_pad  ;
  input \259GAT(55)_pad  ;
  input \260GAT(56)_pad  ;
  input \261GAT(57)_pad  ;
  input \267GAT(58)_pad  ;
  input \268GAT(59)_pad  ;
  input \26GAT(4)_pad  ;
  input \29GAT(5)_pad  ;
  input \36GAT(6)_pad  ;
  input \42GAT(7)_pad  ;
  input \51GAT(8)_pad  ;
  input \55GAT(9)_pad  ;
  input \59GAT(10)_pad  ;
  input \68GAT(11)_pad  ;
  input \72GAT(12)_pad  ;
  input \73GAT(13)_pad  ;
  input \74GAT(14)_pad  ;
  input \75GAT(15)_pad  ;
  input \80GAT(16)_pad  ;
  input \85GAT(17)_pad  ;
  input \86GAT(18)_pad  ;
  input \87GAT(19)_pad  ;
  input \88GAT(20)_pad  ;
  input \89GAT(21)_pad  ;
  input \8GAT(1)_pad  ;
  input \90GAT(22)_pad  ;
  input \91GAT(23)_pad  ;
  input \96GAT(24)_pad  ;
  output \273GAT(103)  ;
  output \388GAT(133)_pad  ;
  output \389GAT(132)_pad  ;
  output \391GAT(124)_pad  ;
  output \393GAT(165)  ;
  output \418GAT(168)_pad  ;
  output \419GAT(164)_pad  ;
  output \420GAT(158)_pad  ;
  output \421GAT(162)_pad  ;
  output \422GAT(161)_pad  ;
  output \423GAT(155)_pad  ;
  output \446GAT(183)_pad  ;
  output \448GAT(179)_pad  ;
  output \449GAT(176)_pad  ;
  output \450GAT(173)_pad  ;
  output \767GAT(349)_pad  ;
  output \768GAT(334)_pad  ;
  output \811GAT(378)  ;
  output \837GAT(396)  ;
  output \838GAT(395)  ;
  output \839GAT(394)  ;
  output \854GAT(419)  ;
  output \866GAT(426)_pad  ;
  output \867GAT(432)  ;
  output \868GAT(431)  ;
  output \869GAT(430)  ;
  wire n61 , n62 , n63 , n64 , n65 , n66 , n67 , n68 , n69 , n70 , n71 , n72 , n73 , n74 , n75 , n76 , n77 , n78 , n79 , n80 , n81 , n82 , n83 , n84 , n85 , n86 , n87 , n88 , n89 , n90 , n91 , n92 , n93 , n94 , n95 , n96 , n97 , n98 , n99 , n100 , n101 , n102 , n103 , n104 , n105 , n106 , n107 , n108 , n109 , n110 , n111 , n112 , n113 , n114 , n115 , n116 , n117 , n118 , n119 , n120 , n121 , n122 , n123 , n124 , n125 , n126 , n127 , n128 , n129 , n130 , n131 , n132 , n133 , n134 , n135 , n136 , n137 , n138 , n139 , n140 , n141 , n142 , n143 , n144 , n145 , n146 , n147 , n148 , n149 , n150 , n151 , n152 , n153 , n154 , n155 , n156 , n157 , n158 , n159 , n160 , n161 , n162 , n163 , n164 , n165 , n166 , n167 , n168 , n169 , n170 , n171 , n172 , n173 , n174 , n175 , n176 , n177 , n178 , n179 , n180 , n181 , n182 , n183 , n184 , n185 , n186 , n187 , n188 , n189 , n190 , n191 , n192 , n193 , n194 , n195 , n196 , n197 , n198 , n199 , n200 , n201 , n202 , n203 , n204 , n205 , n206 , n207 , n208 , n209 , n210 , n211 , n212 , n213 , n214 , n215 , n216 , n217 , n218 , n219 , n220 , n221 , n222 , n223 , n224 , n225 , n226 , n227 , n228 , n229 , n230 , n231 , n232 , n233 , n234 , n235 , n236 , n237 , n238 , n239 , n240 , n241 , n242 , n243 , n244 , n245 , n246 , n247 , n248 , n249 , n250 , n251 , n252 , n253 , n254 , n255 , n256 , n257 , n258 , n259 , n260 , n261 , n262 , n263 , n264 , n265 , n266 , n267 , n268 , n269 , n270 , n271 , n272 , n273 , n274 , n275 , n276 , n277 , n278 , n279 , n280 , n281 , n282 , n283 , n284 , n285 , n286 , n287 , n288 , n289 , n290 , n291 , n292 , n293 , n294 , n295 , n296 , n297 , n298 , n299 , n300 , n301 , n302 , n303 , n304 , n305 , n306 , n307 , n308 , n309 , n310 , n311 , n312 , n313 , n314 , n315 , n316 , n317 , n318 , n319 , n320 , n321 , n322 , n323 , n324 , n325 , n326 , n327 , n328 , n329 , n330 , n331 , n332 , n333 , n334 , n335 , n336 , n337 , n338 , n339 , n340 , n341 , n342 , n343 , n344 , n345 , n346 , n347 , n348 , n349 , n350 , n351 , n352 , n353 , n354 , n355 , n356 , n357 , n358 , n359 , n360 , n361 , n362 , n363 , n364 , n365 , n366 , n367 ;
  assign n61 = \29GAT(5)_pad  & \36GAT(6)_pad  ;
  assign n62 = \42GAT(7)_pad  & n61 ;
  assign n63 = \29GAT(5)_pad  & \75GAT(15)_pad  ;
  assign n64 = \42GAT(7)_pad  & n63 ;
  assign n65 = \80GAT(16)_pad  & n61 ;
  assign n66 = \85GAT(17)_pad  & \86GAT(18)_pad  ;
  assign n67 = \1GAT(0)_pad  & \26GAT(4)_pad  ;
  assign n68 = \51GAT(8)_pad  & n67 ;
  assign n69 = \13GAT(2)_pad  & \17GAT(3)_pad  ;
  assign n70 = \1GAT(0)_pad  & \8GAT(1)_pad  ;
  assign n71 = n69 & n70 ;
  assign n72 = n67 & n69 ;
  assign n73 = ~n62 & n72 ;
  assign n74 = \59GAT(10)_pad  & \75GAT(15)_pad  ;
  assign n75 = \80GAT(16)_pad  & n74 ;
  assign n76 = \36GAT(6)_pad  & \59GAT(10)_pad  ;
  assign n77 = \80GAT(16)_pad  & n76 ;
  assign n78 = \42GAT(7)_pad  & n76 ;
  assign n79 = ~\87GAT(19)_pad  & ~\88GAT(20)_pad  ;
  assign n80 = \90GAT(22)_pad  & ~n79 ;
  assign n81 = n62 & n72 ;
  assign n82 = \13GAT(2)_pad  & \55GAT(9)_pad  ;
  assign n83 = n70 & n82 ;
  assign n84 = \29GAT(5)_pad  & \68GAT(11)_pad  ;
  assign n85 = n83 & n84 ;
  assign n86 = \59GAT(10)_pad  & \68GAT(11)_pad  ;
  assign n87 = n83 & n86 ;
  assign n88 = \74GAT(14)_pad  & n87 ;
  assign n89 = \89GAT(21)_pad  & ~n79 ;
  assign n90 = \111GAT(27)_pad  & ~\91GAT(23)_pad  ;
  assign n91 = ~\111GAT(27)_pad  & \91GAT(23)_pad  ;
  assign n92 = ~n90 & ~n91 ;
  assign n93 = ~\126GAT(30)_pad  & ~\96GAT(24)_pad  ;
  assign n94 = \126GAT(30)_pad  & \96GAT(24)_pad  ;
  assign n95 = ~n93 & ~n94 ;
  assign n96 = n92 & ~n95 ;
  assign n97 = ~n92 & n95 ;
  assign n98 = ~n96 & ~n97 ;
  assign n99 = ~\101GAT(25)_pad  & ~\121GAT(29)_pad  ;
  assign n100 = \101GAT(25)_pad  & \121GAT(29)_pad  ;
  assign n101 = ~n99 & ~n100 ;
  assign n102 = \116GAT(28)_pad  & ~\135GAT(32)_pad  ;
  assign n103 = ~\116GAT(28)_pad  & \135GAT(32)_pad  ;
  assign n104 = ~n102 & ~n103 ;
  assign n105 = n101 & n104 ;
  assign n106 = ~n101 & ~n104 ;
  assign n107 = ~n105 & ~n106 ;
  assign n108 = \106GAT(26)_pad  & ~\130GAT(31)_pad  ;
  assign n109 = ~\106GAT(26)_pad  & \130GAT(31)_pad  ;
  assign n110 = ~n108 & ~n109 ;
  assign n111 = n107 & ~n110 ;
  assign n112 = ~n107 & n110 ;
  assign n113 = ~n111 & ~n112 ;
  assign n114 = n98 & n113 ;
  assign n115 = ~n98 & ~n113 ;
  assign n116 = ~n114 & ~n115 ;
  assign n117 = \171GAT(42)_pad  & ~\177GAT(43)_pad  ;
  assign n118 = ~\171GAT(42)_pad  & \177GAT(43)_pad  ;
  assign n119 = ~n117 & ~n118 ;
  assign n120 = ~\130GAT(31)_pad  & ~\183GAT(44)_pad  ;
  assign n121 = \130GAT(31)_pad  & \183GAT(44)_pad  ;
  assign n122 = ~n120 & ~n121 ;
  assign n123 = n119 & ~n122 ;
  assign n124 = ~n119 & n122 ;
  assign n125 = ~n123 & ~n124 ;
  assign n126 = ~\159GAT(40)_pad  & ~\195GAT(46)_pad  ;
  assign n127 = \159GAT(40)_pad  & \195GAT(46)_pad  ;
  assign n128 = ~n126 & ~n127 ;
  assign n129 = \189GAT(45)_pad  & ~\207GAT(48)_pad  ;
  assign n130 = ~\189GAT(45)_pad  & \207GAT(48)_pad  ;
  assign n131 = ~n129 & ~n130 ;
  assign n132 = n128 & n131 ;
  assign n133 = ~n128 & ~n131 ;
  assign n134 = ~n132 & ~n133 ;
  assign n135 = \165GAT(41)_pad  & ~\201GAT(47)_pad  ;
  assign n136 = ~\165GAT(41)_pad  & \201GAT(47)_pad  ;
  assign n137 = ~n135 & ~n136 ;
  assign n138 = n134 & ~n137 ;
  assign n139 = ~n134 & n137 ;
  assign n140 = ~n138 & ~n139 ;
  assign n141 = n125 & n140 ;
  assign n142 = ~n125 & ~n140 ;
  assign n143 = ~n141 & ~n142 ;
  assign n149 = \42GAT(7)_pad  & n74 ;
  assign n148 = \17GAT(3)_pad  & \51GAT(8)_pad  ;
  assign n150 = n70 & n148 ;
  assign n151 = ~n149 & n150 ;
  assign n153 = \17GAT(3)_pad  & ~\42GAT(7)_pad  ;
  assign n154 = ~\17GAT(3)_pad  & \42GAT(7)_pad  ;
  assign n155 = ~n153 & ~n154 ;
  assign n152 = \156GAT(39)_pad  & \59GAT(10)_pad  ;
  assign n156 = n68 & n152 ;
  assign n157 = ~n155 & n156 ;
  assign n158 = ~n151 & ~n157 ;
  assign n159 = \126GAT(30)_pad  & ~n158 ;
  assign n160 = \55GAT(9)_pad  & n68 ;
  assign n161 = ~\268GAT(59)_pad  & \80GAT(16)_pad  ;
  assign n162 = n63 & n161 ;
  assign n163 = n160 & n162 ;
  assign n164 = n67 & n148 ;
  assign n165 = ~n152 & n164 ;
  assign n166 = \1GAT(0)_pad  & ~n165 ;
  assign n167 = \153GAT(38)_pad  & ~n166 ;
  assign n168 = ~n163 & ~n167 ;
  assign n169 = ~n159 & n168 ;
  assign n170 = \201GAT(47)_pad  & ~n169 ;
  assign n171 = ~\201GAT(47)_pad  & n169 ;
  assign n174 = \261GAT(57)_pad  & ~n171 ;
  assign n175 = ~n170 & n174 ;
  assign n172 = ~n170 & ~n171 ;
  assign n173 = ~\261GAT(57)_pad  & ~n172 ;
  assign n176 = \219GAT(50)_pad  & ~n173 ;
  assign n177 = ~n175 & n176 ;
  assign n178 = \228GAT(51)_pad  & n172 ;
  assign n179 = \201GAT(47)_pad  & \237GAT(52)_pad  ;
  assign n180 = ~\246GAT(53)_pad  & ~n179 ;
  assign n181 = ~n169 & ~n180 ;
  assign n144 = \42GAT(7)_pad  & \72GAT(12)_pad  ;
  assign n145 = \73GAT(13)_pad  & n144 ;
  assign n146 = n87 & n145 ;
  assign n147 = \201GAT(47)_pad  & n146 ;
  assign n182 = \121GAT(29)_pad  & \210GAT(49)_pad  ;
  assign n183 = \255GAT(54)_pad  & \267GAT(58)_pad  ;
  assign n184 = ~n182 & ~n183 ;
  assign n185 = ~n147 & n184 ;
  assign n186 = ~n181 & n185 ;
  assign n187 = ~n178 & n186 ;
  assign n188 = ~n177 & n187 ;
  assign n190 = \111GAT(27)_pad  & ~n158 ;
  assign n191 = \143GAT(34)_pad  & ~n166 ;
  assign n192 = ~n163 & ~n191 ;
  assign n193 = ~n190 & n192 ;
  assign n194 = \183GAT(44)_pad  & ~n193 ;
  assign n195 = ~\183GAT(44)_pad  & n193 ;
  assign n196 = ~n194 & ~n195 ;
  assign n197 = \121GAT(29)_pad  & ~n158 ;
  assign n198 = \149GAT(36)_pad  & ~n166 ;
  assign n199 = ~n163 & ~n198 ;
  assign n200 = ~n197 & n199 ;
  assign n201 = \195GAT(46)_pad  & ~n200 ;
  assign n202 = ~n170 & ~n174 ;
  assign n203 = ~n201 & n202 ;
  assign n204 = ~\195GAT(46)_pad  & n200 ;
  assign n205 = \116GAT(28)_pad  & ~n158 ;
  assign n206 = \146GAT(35)_pad  & ~n166 ;
  assign n207 = ~n163 & ~n206 ;
  assign n208 = ~n205 & n207 ;
  assign n209 = ~\189GAT(45)_pad  & n208 ;
  assign n210 = ~n204 & ~n209 ;
  assign n211 = ~n203 & n210 ;
  assign n212 = \189GAT(45)_pad  & ~n208 ;
  assign n213 = ~n211 & ~n212 ;
  assign n215 = n196 & ~n213 ;
  assign n214 = ~n196 & n213 ;
  assign n216 = \219GAT(50)_pad  & ~n214 ;
  assign n217 = ~n215 & n216 ;
  assign n222 = \228GAT(51)_pad  & n196 ;
  assign n218 = \183GAT(44)_pad  & \237GAT(52)_pad  ;
  assign n219 = ~\246GAT(53)_pad  & ~n218 ;
  assign n220 = ~n193 & ~n219 ;
  assign n189 = \183GAT(44)_pad  & n146 ;
  assign n221 = \106GAT(26)_pad  & \210GAT(49)_pad  ;
  assign n223 = ~n189 & ~n221 ;
  assign n224 = ~n220 & n223 ;
  assign n225 = ~n222 & n224 ;
  assign n226 = ~n217 & n225 ;
  assign n227 = ~n209 & ~n212 ;
  assign n229 = ~n202 & ~n204 ;
  assign n230 = ~n201 & ~n229 ;
  assign n232 = n227 & ~n230 ;
  assign n231 = ~n227 & n230 ;
  assign n233 = \219GAT(50)_pad  & ~n231 ;
  assign n234 = ~n232 & n233 ;
  assign n228 = \228GAT(51)_pad  & n227 ;
  assign n235 = \189GAT(45)_pad  & \237GAT(52)_pad  ;
  assign n236 = ~\246GAT(53)_pad  & ~n235 ;
  assign n237 = ~n208 & ~n236 ;
  assign n239 = \189GAT(45)_pad  & n146 ;
  assign n238 = \111GAT(27)_pad  & \210GAT(49)_pad  ;
  assign n240 = \255GAT(54)_pad  & \259GAT(55)_pad  ;
  assign n241 = ~n238 & ~n240 ;
  assign n242 = ~n239 & n241 ;
  assign n243 = ~n237 & n242 ;
  assign n244 = ~n228 & n243 ;
  assign n245 = ~n234 & n244 ;
  assign n246 = ~n201 & ~n204 ;
  assign n249 = ~n202 & n246 ;
  assign n248 = n202 & ~n246 ;
  assign n250 = \219GAT(50)_pad  & ~n248 ;
  assign n251 = ~n249 & n250 ;
  assign n247 = \228GAT(51)_pad  & n246 ;
  assign n254 = \195GAT(46)_pad  & \237GAT(52)_pad  ;
  assign n255 = ~\246GAT(53)_pad  & ~n254 ;
  assign n256 = ~n200 & ~n255 ;
  assign n253 = \195GAT(46)_pad  & n146 ;
  assign n252 = \116GAT(28)_pad  & \210GAT(49)_pad  ;
  assign n257 = \255GAT(54)_pad  & \260GAT(56)_pad  ;
  assign n258 = ~n252 & ~n257 ;
  assign n259 = ~n253 & n258 ;
  assign n260 = ~n256 & n259 ;
  assign n261 = ~n247 & n260 ;
  assign n262 = ~n251 & n261 ;
  assign n263 = \106GAT(26)_pad  & ~n158 ;
  assign n264 = ~n152 & n160 ;
  assign n265 = \153GAT(38)_pad  & n264 ;
  assign n266 = \138GAT(33)_pad  & \152GAT(37)_pad  ;
  assign n267 = n162 & n164 ;
  assign n268 = ~n266 & ~n267 ;
  assign n269 = ~n265 & n268 ;
  assign n270 = ~n263 & n269 ;
  assign n271 = \177GAT(43)_pad  & ~n270 ;
  assign n272 = ~\177GAT(43)_pad  & n270 ;
  assign n273 = ~n271 & ~n272 ;
  assign n275 = ~n194 & ~n215 ;
  assign n277 = n273 & ~n275 ;
  assign n276 = ~n273 & n275 ;
  assign n278 = \219GAT(50)_pad  & ~n276 ;
  assign n279 = ~n277 & n278 ;
  assign n274 = \228GAT(51)_pad  & n273 ;
  assign n280 = \177GAT(43)_pad  & \237GAT(52)_pad  ;
  assign n281 = ~\246GAT(53)_pad  & ~n280 ;
  assign n282 = ~n270 & ~n281 ;
  assign n283 = \177GAT(43)_pad  & n146 ;
  assign n284 = \101GAT(25)_pad  & \210GAT(49)_pad  ;
  assign n285 = ~n283 & ~n284 ;
  assign n286 = ~n282 & n285 ;
  assign n287 = ~n274 & n286 ;
  assign n288 = ~n279 & n287 ;
  assign n289 = \91GAT(23)_pad  & ~n158 ;
  assign n291 = \143GAT(34)_pad  & n264 ;
  assign n290 = \138GAT(33)_pad  & \8GAT(1)_pad  ;
  assign n292 = ~n267 & ~n290 ;
  assign n293 = ~n291 & n292 ;
  assign n294 = ~n289 & n293 ;
  assign n295 = \159GAT(40)_pad  & ~n294 ;
  assign n296 = ~\159GAT(40)_pad  & n294 ;
  assign n297 = \101GAT(25)_pad  & ~n158 ;
  assign n299 = \149GAT(36)_pad  & n264 ;
  assign n298 = \138GAT(33)_pad  & \17GAT(3)_pad  ;
  assign n300 = ~n267 & ~n298 ;
  assign n301 = ~n299 & n300 ;
  assign n302 = ~n297 & n301 ;
  assign n303 = \171GAT(42)_pad  & ~n302 ;
  assign n304 = ~n272 & ~n275 ;
  assign n305 = ~n271 & ~n304 ;
  assign n306 = ~n303 & n305 ;
  assign n307 = ~\171GAT(42)_pad  & n302 ;
  assign n308 = \96GAT(24)_pad  & ~n158 ;
  assign n310 = \146GAT(35)_pad  & n264 ;
  assign n309 = \138GAT(33)_pad  & \51GAT(8)_pad  ;
  assign n311 = ~n267 & ~n309 ;
  assign n312 = ~n310 & n311 ;
  assign n313 = ~n308 & n312 ;
  assign n314 = ~\165GAT(41)_pad  & n313 ;
  assign n315 = ~n307 & ~n314 ;
  assign n316 = ~n306 & n315 ;
  assign n317 = \165GAT(41)_pad  & ~n313 ;
  assign n318 = ~n316 & ~n317 ;
  assign n319 = ~n296 & ~n318 ;
  assign n320 = ~n295 & ~n319 ;
  assign n321 = ~n295 & ~n296 ;
  assign n323 = n318 & ~n321 ;
  assign n322 = ~n318 & n321 ;
  assign n324 = \219GAT(50)_pad  & ~n322 ;
  assign n325 = ~n323 & n324 ;
  assign n326 = \228GAT(51)_pad  & n321 ;
  assign n327 = \159GAT(40)_pad  & \237GAT(52)_pad  ;
  assign n328 = ~\246GAT(53)_pad  & ~n327 ;
  assign n329 = ~n294 & ~n328 ;
  assign n330 = \159GAT(40)_pad  & n146 ;
  assign n331 = \210GAT(49)_pad  & \268GAT(59)_pad  ;
  assign n332 = ~n330 & ~n331 ;
  assign n333 = ~n329 & n332 ;
  assign n334 = ~n326 & n333 ;
  assign n335 = ~n325 & n334 ;
  assign n337 = ~n314 & ~n317 ;
  assign n338 = ~n305 & ~n307 ;
  assign n339 = ~n303 & ~n338 ;
  assign n341 = n337 & ~n339 ;
  assign n340 = ~n337 & n339 ;
  assign n342 = \219GAT(50)_pad  & ~n340 ;
  assign n343 = ~n341 & n342 ;
  assign n348 = \228GAT(51)_pad  & n337 ;
  assign n344 = \165GAT(41)_pad  & \237GAT(52)_pad  ;
  assign n345 = ~\246GAT(53)_pad  & ~n344 ;
  assign n346 = ~n313 & ~n345 ;
  assign n336 = \165GAT(41)_pad  & n146 ;
  assign n347 = \210GAT(49)_pad  & \91GAT(23)_pad  ;
  assign n349 = ~n336 & ~n347 ;
  assign n350 = ~n346 & n349 ;
  assign n351 = ~n348 & n350 ;
  assign n352 = ~n343 & n351 ;
  assign n353 = ~n303 & ~n307 ;
  assign n356 = n305 & ~n353 ;
  assign n355 = ~n305 & n353 ;
  assign n357 = \219GAT(50)_pad  & ~n355 ;
  assign n358 = ~n356 & n357 ;
  assign n354 = \228GAT(51)_pad  & n353 ;
  assign n359 = \171GAT(42)_pad  & \237GAT(52)_pad  ;
  assign n360 = ~\246GAT(53)_pad  & ~n359 ;
  assign n361 = ~n302 & ~n360 ;
  assign n362 = \171GAT(42)_pad  & n146 ;
  assign n363 = \210GAT(49)_pad  & \96GAT(24)_pad  ;
  assign n364 = ~n362 & ~n363 ;
  assign n365 = ~n361 & n364 ;
  assign n366 = ~n354 & n365 ;
  assign n367 = ~n358 & n366 ;
  assign \273GAT(103)  = n62 ;
  assign \388GAT(133)_pad  = n64 ;
  assign \389GAT(132)_pad  = n65 ;
  assign \391GAT(124)_pad  = n66 ;
  assign \393GAT(165)  = n68 ;
  assign \418GAT(168)_pad  = n71 ;
  assign \419GAT(164)_pad  = ~n73 ;
  assign \420GAT(158)_pad  = ~n75 ;
  assign \421GAT(162)_pad  = ~n77 ;
  assign \422GAT(161)_pad  = ~n78 ;
  assign \423GAT(155)_pad  = n80 ;
  assign \446GAT(183)_pad  = ~n81 ;
  assign \448GAT(179)_pad  = n85 ;
  assign \449GAT(176)_pad  = n88 ;
  assign \450GAT(173)_pad  = n89 ;
  assign \767GAT(349)_pad  = ~n116 ;
  assign \768GAT(334)_pad  = ~n143 ;
  assign \811GAT(378)  = ~n188 ;
  assign \837GAT(396)  = ~n226 ;
  assign \838GAT(395)  = ~n245 ;
  assign \839GAT(394)  = ~n262 ;
  assign \854GAT(419)  = ~n288 ;
  assign \866GAT(426)_pad  = ~n320 ;
  assign \867GAT(432)  = ~n335 ;
  assign \868GAT(431)  = ~n352 ;
  assign \869GAT(430)  = ~n367 ;
endmodule
