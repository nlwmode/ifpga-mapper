module top (a_pad, \b0_pad , b_pad, \c0_pad , c_pad, \d0_pad , d_pad, \e0_pad , e_pad, f_pad, g_pad, \h0_pad , h_pad, i_pad, j_pad, k_pad, l_pad, m_pad, o_pad, t_pad, v_pad, \a0_pad , \f0_pad , \g0_pad , \i0_pad , \j0_pad , \k0_pad , \l0_pad , \m0_pad , \n0_pad , \o0_pad , \p0_pad , w_pad, x_pad, y_pad, z_pad);
	input a_pad ;
	input \b0_pad  ;
	input b_pad ;
	input \c0_pad  ;
	input c_pad ;
	input \d0_pad  ;
	input d_pad ;
	input \e0_pad  ;
	input e_pad ;
	input f_pad ;
	input g_pad ;
	input \h0_pad  ;
	input h_pad ;
	input i_pad ;
	input j_pad ;
	input k_pad ;
	input l_pad ;
	input m_pad ;
	input o_pad ;
	input t_pad ;
	input v_pad ;
	output \a0_pad  ;
	output \f0_pad  ;
	output \g0_pad  ;
	output \i0_pad  ;
	output \j0_pad  ;
	output \k0_pad  ;
	output \l0_pad  ;
	output \m0_pad  ;
	output \n0_pad  ;
	output \o0_pad  ;
	output \p0_pad  ;
	output w_pad ;
	output x_pad ;
	output y_pad ;
	output z_pad ;
	wire _w55_ ;
	wire _w54_ ;
	wire _w53_ ;
	wire _w52_ ;
	wire _w34_ ;
	wire _w33_ ;
	wire _w32_ ;
	wire _w31_ ;
	wire _w30_ ;
	wire _w29_ ;
	wire _w28_ ;
	wire _w27_ ;
	wire _w26_ ;
	wire _w25_ ;
	wire _w24_ ;
	wire _w35_ ;
	wire _w22_ ;
	wire _w51_ ;
	wire _w36_ ;
	wire _w37_ ;
	wire _w38_ ;
	wire _w39_ ;
	wire _w40_ ;
	wire _w41_ ;
	wire _w42_ ;
	wire _w43_ ;
	wire _w44_ ;
	wire _w45_ ;
	wire _w46_ ;
	wire _w47_ ;
	wire _w48_ ;
	wire _w49_ ;
	wire _w50_ ;
	LUT1 #(
		.INIT('h1)
	) name0 (
		t_pad,
		_w22_
	);
	LUT2 #(
		.INIT('h8)
	) name1 (
		i_pad,
		j_pad,
		_w24_
	);
	LUT2 #(
		.INIT('h7)
	) name2 (
		i_pad,
		j_pad,
		_w25_
	);
	LUT3 #(
		.INIT('h40)
	) name3 (
		\c0_pad ,
		i_pad,
		k_pad,
		_w26_
	);
	LUT4 #(
		.INIT('h1000)
	) name4 (
		a_pad,
		\c0_pad ,
		i_pad,
		k_pad,
		_w27_
	);
	LUT4 #(
		.INIT('h00bf)
	) name5 (
		\c0_pad ,
		i_pad,
		k_pad,
		o_pad,
		_w28_
	);
	LUT3 #(
		.INIT('h02)
	) name6 (
		m_pad,
		_w28_,
		_w27_,
		_w29_
	);
	LUT4 #(
		.INIT('h2000)
	) name7 (
		b_pad,
		\c0_pad ,
		i_pad,
		k_pad,
		_w30_
	);
	LUT4 #(
		.INIT('h1333)
	) name8 (
		\c0_pad ,
		\h0_pad ,
		i_pad,
		k_pad,
		_w31_
	);
	LUT3 #(
		.INIT('h02)
	) name9 (
		m_pad,
		_w31_,
		_w30_,
		_w32_
	);
	LUT4 #(
		.INIT('h1555)
	) name10 (
		\c0_pad ,
		c_pad,
		i_pad,
		k_pad,
		_w33_
	);
	LUT4 #(
		.INIT('h7f00)
	) name11 (
		\c0_pad ,
		i_pad,
		k_pad,
		m_pad,
		_w34_
	);
	LUT2 #(
		.INIT('h4)
	) name12 (
		_w33_,
		_w34_,
		_w35_
	);
	LUT2 #(
		.INIT('h2)
	) name13 (
		\e0_pad ,
		\h0_pad ,
		_w36_
	);
	LUT4 #(
		.INIT('h8c80)
	) name14 (
		d_pad,
		m_pad,
		_w26_,
		_w36_,
		_w37_
	);
	LUT4 #(
		.INIT('h1000)
	) name15 (
		\c0_pad ,
		e_pad,
		i_pad,
		k_pad,
		_w38_
	);
	LUT4 #(
		.INIT('h2333)
	) name16 (
		\c0_pad ,
		\d0_pad ,
		i_pad,
		k_pad,
		_w39_
	);
	LUT3 #(
		.INIT('h02)
	) name17 (
		m_pad,
		_w39_,
		_w38_,
		_w40_
	);
	LUT4 #(
		.INIT('h1000)
	) name18 (
		\c0_pad ,
		f_pad,
		i_pad,
		k_pad,
		_w41_
	);
	LUT4 #(
		.INIT('h00bf)
	) name19 (
		\c0_pad ,
		i_pad,
		k_pad,
		t_pad,
		_w42_
	);
	LUT3 #(
		.INIT('h02)
	) name20 (
		m_pad,
		_w42_,
		_w41_,
		_w43_
	);
	LUT4 #(
		.INIT('h1000)
	) name21 (
		\c0_pad ,
		g_pad,
		i_pad,
		k_pad,
		_w44_
	);
	LUT4 #(
		.INIT('h4555)
	) name22 (
		\b0_pad ,
		\c0_pad ,
		i_pad,
		k_pad,
		_w45_
	);
	LUT3 #(
		.INIT('h02)
	) name23 (
		m_pad,
		_w45_,
		_w44_,
		_w46_
	);
	LUT4 #(
		.INIT('h1000)
	) name24 (
		\c0_pad ,
		h_pad,
		i_pad,
		k_pad,
		_w47_
	);
	LUT4 #(
		.INIT('h00bf)
	) name25 (
		\c0_pad ,
		i_pad,
		k_pad,
		v_pad,
		_w48_
	);
	LUT3 #(
		.INIT('h02)
	) name26 (
		m_pad,
		_w48_,
		_w47_,
		_w49_
	);
	LUT2 #(
		.INIT('h8)
	) name27 (
		l_pad,
		v_pad,
		_w50_
	);
	LUT4 #(
		.INIT('h2000)
	) name28 (
		\c0_pad ,
		\h0_pad ,
		i_pad,
		k_pad,
		_w51_
	);
	LUT4 #(
		.INIT('h2333)
	) name29 (
		\c0_pad ,
		\h0_pad ,
		i_pad,
		k_pad,
		_w52_
	);
	LUT2 #(
		.INIT('h4)
	) name30 (
		l_pad,
		m_pad,
		_w53_
	);
	LUT2 #(
		.INIT('h4)
	) name31 (
		_w52_,
		_w53_,
		_w54_
	);
	LUT2 #(
		.INIT('h8)
	) name32 (
		m_pad,
		_w51_,
		_w55_
	);
	assign \a0_pad  = _w22_ ;
	assign \f0_pad  = _w24_ ;
	assign \g0_pad  = _w25_ ;
	assign \i0_pad  = _w29_ ;
	assign \j0_pad  = _w32_ ;
	assign \k0_pad  = _w35_ ;
	assign \l0_pad  = _w37_ ;
	assign \m0_pad  = _w40_ ;
	assign \n0_pad  = _w43_ ;
	assign \o0_pad  = _w46_ ;
	assign \p0_pad  = _w49_ ;
	assign w_pad = _w50_ ;
	assign x_pad = _w51_ ;
	assign y_pad = _w54_ ;
	assign z_pad = _w55_ ;
endmodule;