module top( \a0_pad  , a_pad , \b0_pad  , b_pad , \c0_pad  , c_pad , \d0_pad  , d_pad , \e0_pad  , e_pad , \f0_pad  , f_pad , \g0_pad  , g_pad , \h0_pad  , h_pad , \i0_pad  , i_pad , \j0_pad  , j_pad , \k0_pad  , k_pad , \l0_pad  , l_pad , \m0_pad  , m_pad , \n0_pad  , n_pad , \o0_pad  , o_pad , p_pad , q_pad , r_pad , s_pad , t_pad , u_pad , v_pad , w_pad , x_pad , y_pad , z_pad , \a1_pad  , \b1_pad  , \c1_pad  , \d1_pad  , \e1_pad  , \f1_pad  , \g1_pad  , \h1_pad  , \i1_pad  , \j1_pad  , \j4  , \p0_pad  , \q0_pad  , \r0_pad  , \s0_pad  , \t0_pad  , \u277_syn_3  , \v0_pad  , \w0_pad  , \y0_pad  , \z0_pad  );
  input \a0_pad  ;
  input a_pad ;
  input \b0_pad  ;
  input b_pad ;
  input \c0_pad  ;
  input c_pad ;
  input \d0_pad  ;
  input d_pad ;
  input \e0_pad  ;
  input e_pad ;
  input \f0_pad  ;
  input f_pad ;
  input \g0_pad  ;
  input g_pad ;
  input \h0_pad  ;
  input h_pad ;
  input \i0_pad  ;
  input i_pad ;
  input \j0_pad  ;
  input j_pad ;
  input \k0_pad  ;
  input k_pad ;
  input \l0_pad  ;
  input l_pad ;
  input \m0_pad  ;
  input m_pad ;
  input \n0_pad  ;
  input n_pad ;
  input \o0_pad  ;
  input o_pad ;
  input p_pad ;
  input q_pad ;
  input r_pad ;
  input s_pad ;
  input t_pad ;
  input u_pad ;
  input v_pad ;
  input w_pad ;
  input x_pad ;
  input y_pad ;
  input z_pad ;
  output \a1_pad  ;
  output \b1_pad  ;
  output \c1_pad  ;
  output \d1_pad  ;
  output \e1_pad  ;
  output \f1_pad  ;
  output \g1_pad  ;
  output \h1_pad  ;
  output \i1_pad  ;
  output \j1_pad  ;
  output \j4  ;
  output \p0_pad  ;
  output \q0_pad  ;
  output \r0_pad  ;
  output \s0_pad  ;
  output \t0_pad  ;
  output \u277_syn_3  ;
  output \v0_pad  ;
  output \w0_pad  ;
  output \y0_pad  ;
  output \z0_pad  ;
  wire n42 , n43 , n44 , n45 , n46 , n47 , n48 , n49 , n50 , n51 , n52 , n53 , n54 , n55 , n56 , n57 , n58 , n59 , n60 , n61 , n62 , n63 , n64 , n65 , n66 , n67 , n68 , n69 , n70 , n71 , n72 , n73 , n74 , n75 , n76 , n77 , n78 , n79 , n80 , n81 , n82 , n83 , n84 , n85 , n86 , n87 , n88 , n89 , n90 , n91 , n92 , n93 , n94 , n95 , n96 , n97 , n98 , n99 , n100 , n101 , n102 , n103 , n104 , n105 , n106 , n107 , n108 , n109 , n110 , n111 , n112 , n113 , n114 , n115 , n116 , n117 , n118 , n119 , n120 , n121 ;
  assign n42 = ~\c0_pad  & \j0_pad  ;
  assign n43 = ~\b0_pad  & ~i_pad ;
  assign n44 = n42 & ~n43 ;
  assign n45 = \b0_pad  & e_pad ;
  assign n46 = n44 & ~n45 ;
  assign n47 = \d0_pad  & i_pad ;
  assign n48 = \n0_pad  & \o0_pad  ;
  assign n49 = n47 & n48 ;
  assign n50 = ~\e0_pad  & ~j_pad ;
  assign n51 = ~n49 & n50 ;
  assign n52 = ~n46 & n51 ;
  assign n53 = ~\k0_pad  & ~n42 ;
  assign n54 = \b0_pad  & ~e_pad ;
  assign n55 = ~n53 & n54 ;
  assign n56 = ~e_pad & k_pad ;
  assign n57 = ~n55 & ~n56 ;
  assign n58 = n48 & ~n57 ;
  assign n59 = \c0_pad  & \j0_pad  ;
  assign n60 = ~\l0_pad  & ~n59 ;
  assign n61 = \b0_pad  & ~n60 ;
  assign n62 = ~n58 & ~n61 ;
  assign n63 = ~s_pad & ~t_pad ;
  assign n64 = u_pad & n63 ;
  assign n65 = n61 & n64 ;
  assign n66 = ~\e0_pad  & ~\g0_pad  ;
  assign n67 = \j0_pad  & \k0_pad  ;
  assign n68 = \c0_pad  & ~n67 ;
  assign n69 = \b0_pad  & ~n68 ;
  assign n70 = n66 & ~n69 ;
  assign n71 = ~e_pad & ~n_pad ;
  assign n72 = n48 & n71 ;
  assign n73 = ~n70 & n72 ;
  assign n74 = ~n65 & ~n73 ;
  assign n75 = \a0_pad  & \b0_pad  ;
  assign n76 = \i0_pad  & n75 ;
  assign n77 = m_pad & n76 ;
  assign n78 = b_pad & w_pad ;
  assign n79 = ~x_pad & n78 ;
  assign n80 = x_pad & ~y_pad ;
  assign n81 = n78 & n80 ;
  assign n82 = ~\c0_pad  & i_pad ;
  assign n83 = ~\b0_pad  & ~n82 ;
  assign n84 = \j0_pad  & ~n83 ;
  assign n85 = n51 & ~n84 ;
  assign n86 = \b0_pad  & \c0_pad  ;
  assign n87 = ~\l0_pad  & ~n86 ;
  assign n88 = ~p_pad & ~n62 ;
  assign n89 = q_pad & ~n88 ;
  assign n90 = \b0_pad  & ~n53 ;
  assign n91 = n66 & ~n90 ;
  assign n92 = e_pad & ~n91 ;
  assign n94 = e_pad & ~n44 ;
  assign n93 = ~c_pad & ~n47 ;
  assign n95 = n48 & ~n93 ;
  assign n96 = ~n94 & n95 ;
  assign n97 = ~\b0_pad  & \l0_pad  ;
  assign n98 = \j0_pad  & n86 ;
  assign n99 = ~n97 & ~n98 ;
  assign n100 = v_pad & ~n99 ;
  assign n101 = ~v_pad & ~n99 ;
  assign n107 = a_pad & ~z_pad ;
  assign n106 = ~o_pad & z_pad ;
  assign n108 = \m0_pad  & ~n106 ;
  assign n109 = ~n107 & n108 ;
  assign n102 = ~p_pad & r_pad ;
  assign n103 = ~\f0_pad  & ~\h0_pad  ;
  assign n104 = ~n102 & n103 ;
  assign n105 = o_pad & ~n104 ;
  assign n110 = d_pad & ~n105 ;
  assign n111 = ~n109 & n110 ;
  assign n112 = l_pad & n76 ;
  assign n117 = ~e_pad & f_pad ;
  assign n118 = n48 & n117 ;
  assign n119 = ~n91 & n118 ;
  assign n113 = \b0_pad  & g_pad ;
  assign n114 = \l0_pad  & n113 ;
  assign n115 = h_pad & ~n48 ;
  assign n116 = n55 & n115 ;
  assign n120 = ~n114 & ~n116 ;
  assign n121 = ~n119 & n120 ;
  assign \a1_pad  = n52 ;
  assign \b1_pad  = n62 ;
  assign \c1_pad  = ~n74 ;
  assign \d1_pad  = n74 ;
  assign \e1_pad  = n77 ;
  assign \f1_pad  = n79 ;
  assign \g1_pad  = n81 ;
  assign \h1_pad  = ~n52 ;
  assign \i1_pad  = n52 ;
  assign \j1_pad  = n85 ;
  assign \j4  = ~n87 ;
  assign \p0_pad  = ~n89 ;
  assign \q0_pad  = ~n92 ;
  assign \r0_pad  = ~n96 ;
  assign \s0_pad  = ~n100 ;
  assign \t0_pad  = ~n101 ;
  assign \u277_syn_3  = n48 ;
  assign \v0_pad  = n87 ;
  assign \w0_pad  = n111 ;
  assign \y0_pad  = n112 ;
  assign \z0_pad  = ~n121 ;
endmodule
