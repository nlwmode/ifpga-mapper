module top (\103GAT(6)_pad , \120GAT(7)_pad , \137GAT(8)_pad , \154GAT(9)_pad , \171GAT(10)_pad , \188GAT(11)_pad , \18GAT(1)_pad , \1GAT(0)_pad , \205GAT(12)_pad , \222GAT(13)_pad , \239GAT(14)_pad , \256GAT(15)_pad , \273GAT(16)_pad , \290GAT(17)_pad , \307GAT(18)_pad , \324GAT(19)_pad , \341GAT(20)_pad , \358GAT(21)_pad , \35GAT(2)_pad , \375GAT(22)_pad , \392GAT(23)_pad , \409GAT(24)_pad , \426GAT(25)_pad , \443GAT(26)_pad , \460GAT(27)_pad , \477GAT(28)_pad , \494GAT(29)_pad , \511GAT(30)_pad , \528GAT(31)_pad , \52GAT(3)_pad , \69GAT(4)_pad , \86GAT(5)_pad , \1581GAT(423)_pad , \1901GAT(561)_pad , \2223GAT(700)_pad , \2548GAT(840)_pad , \2877GAT(983)_pad , \3211GAT(1128)_pad , \3552GAT(1275)_pad , \3895GAT(1423)_pad , \4241GAT(1572)_pad , \4591GAT(1722)_pad , \4946GAT(1876)_pad , \5308GAT(2031)_pad , \545GAT(287)_pad , \5672GAT(2187)_pad , \5971GAT(2309)_pad , \6123GAT(2368)_pad , \6150GAT(2378)_pad , \6160GAT(2383)_pad , \6170GAT(2388)_pad , \6180GAT(2393)_pad , \6190GAT(2398)_pad , \6200GAT(2403)_pad , \6210GAT(2408)_pad , \6220GAT(2413)_pad , \6230GAT(2418)_pad , \6240GAT(2423)_pad , \6250GAT(2428)_pad , \6260GAT(2433)_pad , \6270GAT(2438)_pad , \6280GAT(2443)_pad , \6287GAT(2444)_pad , \6288GAT(2447)_pad );
	input \103GAT(6)_pad  ;
	input \120GAT(7)_pad  ;
	input \137GAT(8)_pad  ;
	input \154GAT(9)_pad  ;
	input \171GAT(10)_pad  ;
	input \188GAT(11)_pad  ;
	input \18GAT(1)_pad  ;
	input \1GAT(0)_pad  ;
	input \205GAT(12)_pad  ;
	input \222GAT(13)_pad  ;
	input \239GAT(14)_pad  ;
	input \256GAT(15)_pad  ;
	input \273GAT(16)_pad  ;
	input \290GAT(17)_pad  ;
	input \307GAT(18)_pad  ;
	input \324GAT(19)_pad  ;
	input \341GAT(20)_pad  ;
	input \358GAT(21)_pad  ;
	input \35GAT(2)_pad  ;
	input \375GAT(22)_pad  ;
	input \392GAT(23)_pad  ;
	input \409GAT(24)_pad  ;
	input \426GAT(25)_pad  ;
	input \443GAT(26)_pad  ;
	input \460GAT(27)_pad  ;
	input \477GAT(28)_pad  ;
	input \494GAT(29)_pad  ;
	input \511GAT(30)_pad  ;
	input \528GAT(31)_pad  ;
	input \52GAT(3)_pad  ;
	input \69GAT(4)_pad  ;
	input \86GAT(5)_pad  ;
	output \1581GAT(423)_pad  ;
	output \1901GAT(561)_pad  ;
	output \2223GAT(700)_pad  ;
	output \2548GAT(840)_pad  ;
	output \2877GAT(983)_pad  ;
	output \3211GAT(1128)_pad  ;
	output \3552GAT(1275)_pad  ;
	output \3895GAT(1423)_pad  ;
	output \4241GAT(1572)_pad  ;
	output \4591GAT(1722)_pad  ;
	output \4946GAT(1876)_pad  ;
	output \5308GAT(2031)_pad  ;
	output \545GAT(287)_pad  ;
	output \5672GAT(2187)_pad  ;
	output \5971GAT(2309)_pad  ;
	output \6123GAT(2368)_pad  ;
	output \6150GAT(2378)_pad  ;
	output \6160GAT(2383)_pad  ;
	output \6170GAT(2388)_pad  ;
	output \6180GAT(2393)_pad  ;
	output \6190GAT(2398)_pad  ;
	output \6200GAT(2403)_pad  ;
	output \6210GAT(2408)_pad  ;
	output \6220GAT(2413)_pad  ;
	output \6230GAT(2418)_pad  ;
	output \6240GAT(2423)_pad  ;
	output \6250GAT(2428)_pad  ;
	output \6260GAT(2433)_pad  ;
	output \6270GAT(2438)_pad  ;
	output \6280GAT(2443)_pad  ;
	output \6287GAT(2444)_pad  ;
	output \6288GAT(2447)_pad  ;
	wire _w875_ ;
	wire _w874_ ;
	wire _w873_ ;
	wire _w872_ ;
	wire _w871_ ;
	wire _w870_ ;
	wire _w869_ ;
	wire _w868_ ;
	wire _w867_ ;
	wire _w866_ ;
	wire _w865_ ;
	wire _w864_ ;
	wire _w863_ ;
	wire _w862_ ;
	wire _w861_ ;
	wire _w860_ ;
	wire _w859_ ;
	wire _w858_ ;
	wire _w857_ ;
	wire _w856_ ;
	wire _w855_ ;
	wire _w854_ ;
	wire _w853_ ;
	wire _w852_ ;
	wire _w851_ ;
	wire _w850_ ;
	wire _w849_ ;
	wire _w848_ ;
	wire _w847_ ;
	wire _w846_ ;
	wire _w845_ ;
	wire _w844_ ;
	wire _w843_ ;
	wire _w842_ ;
	wire _w841_ ;
	wire _w840_ ;
	wire _w839_ ;
	wire _w838_ ;
	wire _w837_ ;
	wire _w836_ ;
	wire _w835_ ;
	wire _w834_ ;
	wire _w833_ ;
	wire _w832_ ;
	wire _w831_ ;
	wire _w830_ ;
	wire _w829_ ;
	wire _w828_ ;
	wire _w827_ ;
	wire _w826_ ;
	wire _w825_ ;
	wire _w824_ ;
	wire _w823_ ;
	wire _w822_ ;
	wire _w821_ ;
	wire _w820_ ;
	wire _w819_ ;
	wire _w818_ ;
	wire _w817_ ;
	wire _w816_ ;
	wire _w815_ ;
	wire _w814_ ;
	wire _w813_ ;
	wire _w812_ ;
	wire _w811_ ;
	wire _w810_ ;
	wire _w809_ ;
	wire _w808_ ;
	wire _w807_ ;
	wire _w806_ ;
	wire _w805_ ;
	wire _w804_ ;
	wire _w803_ ;
	wire _w802_ ;
	wire _w801_ ;
	wire _w800_ ;
	wire _w799_ ;
	wire _w798_ ;
	wire _w797_ ;
	wire _w796_ ;
	wire _w795_ ;
	wire _w794_ ;
	wire _w793_ ;
	wire _w792_ ;
	wire _w791_ ;
	wire _w790_ ;
	wire _w789_ ;
	wire _w788_ ;
	wire _w787_ ;
	wire _w786_ ;
	wire _w785_ ;
	wire _w784_ ;
	wire _w783_ ;
	wire _w782_ ;
	wire _w781_ ;
	wire _w780_ ;
	wire _w779_ ;
	wire _w778_ ;
	wire _w777_ ;
	wire _w776_ ;
	wire _w775_ ;
	wire _w774_ ;
	wire _w773_ ;
	wire _w772_ ;
	wire _w771_ ;
	wire _w770_ ;
	wire _w769_ ;
	wire _w768_ ;
	wire _w767_ ;
	wire _w766_ ;
	wire _w765_ ;
	wire _w764_ ;
	wire _w763_ ;
	wire _w762_ ;
	wire _w761_ ;
	wire _w760_ ;
	wire _w759_ ;
	wire _w758_ ;
	wire _w757_ ;
	wire _w756_ ;
	wire _w755_ ;
	wire _w754_ ;
	wire _w753_ ;
	wire _w752_ ;
	wire _w751_ ;
	wire _w750_ ;
	wire _w749_ ;
	wire _w748_ ;
	wire _w747_ ;
	wire _w746_ ;
	wire _w745_ ;
	wire _w744_ ;
	wire _w743_ ;
	wire _w742_ ;
	wire _w741_ ;
	wire _w740_ ;
	wire _w739_ ;
	wire _w738_ ;
	wire _w737_ ;
	wire _w736_ ;
	wire _w735_ ;
	wire _w734_ ;
	wire _w733_ ;
	wire _w732_ ;
	wire _w731_ ;
	wire _w730_ ;
	wire _w729_ ;
	wire _w728_ ;
	wire _w727_ ;
	wire _w726_ ;
	wire _w725_ ;
	wire _w724_ ;
	wire _w723_ ;
	wire _w722_ ;
	wire _w721_ ;
	wire _w720_ ;
	wire _w719_ ;
	wire _w718_ ;
	wire _w717_ ;
	wire _w716_ ;
	wire _w715_ ;
	wire _w714_ ;
	wire _w713_ ;
	wire _w712_ ;
	wire _w711_ ;
	wire _w710_ ;
	wire _w709_ ;
	wire _w708_ ;
	wire _w707_ ;
	wire _w706_ ;
	wire _w705_ ;
	wire _w704_ ;
	wire _w703_ ;
	wire _w702_ ;
	wire _w701_ ;
	wire _w700_ ;
	wire _w699_ ;
	wire _w698_ ;
	wire _w697_ ;
	wire _w696_ ;
	wire _w695_ ;
	wire _w694_ ;
	wire _w693_ ;
	wire _w692_ ;
	wire _w691_ ;
	wire _w690_ ;
	wire _w689_ ;
	wire _w688_ ;
	wire _w687_ ;
	wire _w686_ ;
	wire _w685_ ;
	wire _w684_ ;
	wire _w683_ ;
	wire _w682_ ;
	wire _w681_ ;
	wire _w680_ ;
	wire _w679_ ;
	wire _w678_ ;
	wire _w677_ ;
	wire _w676_ ;
	wire _w675_ ;
	wire _w674_ ;
	wire _w673_ ;
	wire _w672_ ;
	wire _w671_ ;
	wire _w670_ ;
	wire _w669_ ;
	wire _w668_ ;
	wire _w667_ ;
	wire _w666_ ;
	wire _w665_ ;
	wire _w664_ ;
	wire _w663_ ;
	wire _w662_ ;
	wire _w661_ ;
	wire _w660_ ;
	wire _w659_ ;
	wire _w658_ ;
	wire _w657_ ;
	wire _w656_ ;
	wire _w655_ ;
	wire _w654_ ;
	wire _w653_ ;
	wire _w652_ ;
	wire _w651_ ;
	wire _w650_ ;
	wire _w649_ ;
	wire _w648_ ;
	wire _w647_ ;
	wire _w646_ ;
	wire _w645_ ;
	wire _w644_ ;
	wire _w643_ ;
	wire _w642_ ;
	wire _w641_ ;
	wire _w640_ ;
	wire _w639_ ;
	wire _w638_ ;
	wire _w637_ ;
	wire _w636_ ;
	wire _w635_ ;
	wire _w634_ ;
	wire _w633_ ;
	wire _w632_ ;
	wire _w631_ ;
	wire _w630_ ;
	wire _w629_ ;
	wire _w628_ ;
	wire _w627_ ;
	wire _w626_ ;
	wire _w625_ ;
	wire _w624_ ;
	wire _w623_ ;
	wire _w622_ ;
	wire _w621_ ;
	wire _w620_ ;
	wire _w619_ ;
	wire _w618_ ;
	wire _w617_ ;
	wire _w616_ ;
	wire _w615_ ;
	wire _w614_ ;
	wire _w613_ ;
	wire _w612_ ;
	wire _w611_ ;
	wire _w610_ ;
	wire _w609_ ;
	wire _w608_ ;
	wire _w607_ ;
	wire _w606_ ;
	wire _w605_ ;
	wire _w604_ ;
	wire _w603_ ;
	wire _w602_ ;
	wire _w601_ ;
	wire _w600_ ;
	wire _w599_ ;
	wire _w598_ ;
	wire _w597_ ;
	wire _w596_ ;
	wire _w595_ ;
	wire _w594_ ;
	wire _w593_ ;
	wire _w592_ ;
	wire _w591_ ;
	wire _w590_ ;
	wire _w589_ ;
	wire _w588_ ;
	wire _w587_ ;
	wire _w586_ ;
	wire _w585_ ;
	wire _w584_ ;
	wire _w583_ ;
	wire _w582_ ;
	wire _w581_ ;
	wire _w580_ ;
	wire _w579_ ;
	wire _w578_ ;
	wire _w577_ ;
	wire _w576_ ;
	wire _w575_ ;
	wire _w290_ ;
	wire _w289_ ;
	wire _w288_ ;
	wire _w287_ ;
	wire _w286_ ;
	wire _w285_ ;
	wire _w284_ ;
	wire _w283_ ;
	wire _w282_ ;
	wire _w281_ ;
	wire _w280_ ;
	wire _w279_ ;
	wire _w278_ ;
	wire _w277_ ;
	wire _w276_ ;
	wire _w275_ ;
	wire _w274_ ;
	wire _w273_ ;
	wire _w272_ ;
	wire _w271_ ;
	wire _w270_ ;
	wire _w269_ ;
	wire _w268_ ;
	wire _w267_ ;
	wire _w266_ ;
	wire _w265_ ;
	wire _w264_ ;
	wire _w263_ ;
	wire _w262_ ;
	wire _w261_ ;
	wire _w260_ ;
	wire _w259_ ;
	wire _w258_ ;
	wire _w257_ ;
	wire _w256_ ;
	wire _w255_ ;
	wire _w254_ ;
	wire _w253_ ;
	wire _w252_ ;
	wire _w251_ ;
	wire _w250_ ;
	wire _w249_ ;
	wire _w248_ ;
	wire _w247_ ;
	wire _w246_ ;
	wire _w245_ ;
	wire _w244_ ;
	wire _w243_ ;
	wire _w242_ ;
	wire _w241_ ;
	wire _w240_ ;
	wire _w239_ ;
	wire _w238_ ;
	wire _w237_ ;
	wire _w236_ ;
	wire _w235_ ;
	wire _w234_ ;
	wire _w233_ ;
	wire _w232_ ;
	wire _w231_ ;
	wire _w230_ ;
	wire _w229_ ;
	wire _w228_ ;
	wire _w227_ ;
	wire _w226_ ;
	wire _w225_ ;
	wire _w224_ ;
	wire _w223_ ;
	wire _w222_ ;
	wire _w221_ ;
	wire _w220_ ;
	wire _w219_ ;
	wire _w218_ ;
	wire _w217_ ;
	wire _w216_ ;
	wire _w215_ ;
	wire _w214_ ;
	wire _w213_ ;
	wire _w212_ ;
	wire _w211_ ;
	wire _w210_ ;
	wire _w209_ ;
	wire _w208_ ;
	wire _w207_ ;
	wire _w206_ ;
	wire _w205_ ;
	wire _w204_ ;
	wire _w203_ ;
	wire _w202_ ;
	wire _w201_ ;
	wire _w200_ ;
	wire _w199_ ;
	wire _w198_ ;
	wire _w197_ ;
	wire _w196_ ;
	wire _w195_ ;
	wire _w194_ ;
	wire _w193_ ;
	wire _w192_ ;
	wire _w191_ ;
	wire _w190_ ;
	wire _w189_ ;
	wire _w188_ ;
	wire _w187_ ;
	wire _w186_ ;
	wire _w185_ ;
	wire _w184_ ;
	wire _w183_ ;
	wire _w182_ ;
	wire _w181_ ;
	wire _w180_ ;
	wire _w179_ ;
	wire _w178_ ;
	wire _w177_ ;
	wire _w176_ ;
	wire _w175_ ;
	wire _w174_ ;
	wire _w173_ ;
	wire _w172_ ;
	wire _w171_ ;
	wire _w170_ ;
	wire _w169_ ;
	wire _w168_ ;
	wire _w167_ ;
	wire _w166_ ;
	wire _w165_ ;
	wire _w164_ ;
	wire _w163_ ;
	wire _w162_ ;
	wire _w161_ ;
	wire _w92_ ;
	wire _w91_ ;
	wire _w90_ ;
	wire _w89_ ;
	wire _w88_ ;
	wire _w87_ ;
	wire _w86_ ;
	wire _w85_ ;
	wire _w84_ ;
	wire _w83_ ;
	wire _w82_ ;
	wire _w81_ ;
	wire _w80_ ;
	wire _w79_ ;
	wire _w78_ ;
	wire _w77_ ;
	wire _w76_ ;
	wire _w75_ ;
	wire _w74_ ;
	wire _w73_ ;
	wire _w72_ ;
	wire _w71_ ;
	wire _w70_ ;
	wire _w69_ ;
	wire _w68_ ;
	wire _w67_ ;
	wire _w66_ ;
	wire _w65_ ;
	wire _w64_ ;
	wire _w63_ ;
	wire _w46_ ;
	wire _w45_ ;
	wire _w44_ ;
	wire _w43_ ;
	wire _w42_ ;
	wire _w41_ ;
	wire _w40_ ;
	wire _w39_ ;
	wire _w38_ ;
	wire _w37_ ;
	wire _w36_ ;
	wire _w35_ ;
	wire _w34_ ;
	wire _w47_ ;
	wire _w48_ ;
	wire _w49_ ;
	wire _w50_ ;
	wire _w51_ ;
	wire _w52_ ;
	wire _w53_ ;
	wire _w54_ ;
	wire _w55_ ;
	wire _w56_ ;
	wire _w57_ ;
	wire _w58_ ;
	wire _w59_ ;
	wire _w60_ ;
	wire _w61_ ;
	wire _w62_ ;
	wire _w93_ ;
	wire _w94_ ;
	wire _w95_ ;
	wire _w96_ ;
	wire _w97_ ;
	wire _w98_ ;
	wire _w99_ ;
	wire _w100_ ;
	wire _w101_ ;
	wire _w102_ ;
	wire _w103_ ;
	wire _w104_ ;
	wire _w105_ ;
	wire _w106_ ;
	wire _w107_ ;
	wire _w108_ ;
	wire _w109_ ;
	wire _w110_ ;
	wire _w111_ ;
	wire _w112_ ;
	wire _w113_ ;
	wire _w114_ ;
	wire _w115_ ;
	wire _w116_ ;
	wire _w117_ ;
	wire _w118_ ;
	wire _w119_ ;
	wire _w120_ ;
	wire _w121_ ;
	wire _w122_ ;
	wire _w123_ ;
	wire _w124_ ;
	wire _w125_ ;
	wire _w126_ ;
	wire _w127_ ;
	wire _w128_ ;
	wire _w129_ ;
	wire _w130_ ;
	wire _w131_ ;
	wire _w132_ ;
	wire _w133_ ;
	wire _w134_ ;
	wire _w135_ ;
	wire _w136_ ;
	wire _w137_ ;
	wire _w138_ ;
	wire _w139_ ;
	wire _w140_ ;
	wire _w141_ ;
	wire _w142_ ;
	wire _w143_ ;
	wire _w144_ ;
	wire _w145_ ;
	wire _w146_ ;
	wire _w147_ ;
	wire _w148_ ;
	wire _w149_ ;
	wire _w150_ ;
	wire _w151_ ;
	wire _w152_ ;
	wire _w153_ ;
	wire _w154_ ;
	wire _w155_ ;
	wire _w156_ ;
	wire _w157_ ;
	wire _w158_ ;
	wire _w159_ ;
	wire _w160_ ;
	wire _w291_ ;
	wire _w292_ ;
	wire _w293_ ;
	wire _w294_ ;
	wire _w295_ ;
	wire _w296_ ;
	wire _w297_ ;
	wire _w298_ ;
	wire _w299_ ;
	wire _w300_ ;
	wire _w301_ ;
	wire _w302_ ;
	wire _w303_ ;
	wire _w304_ ;
	wire _w305_ ;
	wire _w306_ ;
	wire _w307_ ;
	wire _w308_ ;
	wire _w309_ ;
	wire _w310_ ;
	wire _w311_ ;
	wire _w312_ ;
	wire _w313_ ;
	wire _w314_ ;
	wire _w315_ ;
	wire _w316_ ;
	wire _w317_ ;
	wire _w318_ ;
	wire _w319_ ;
	wire _w320_ ;
	wire _w321_ ;
	wire _w322_ ;
	wire _w323_ ;
	wire _w324_ ;
	wire _w325_ ;
	wire _w326_ ;
	wire _w327_ ;
	wire _w328_ ;
	wire _w329_ ;
	wire _w330_ ;
	wire _w331_ ;
	wire _w332_ ;
	wire _w333_ ;
	wire _w334_ ;
	wire _w335_ ;
	wire _w336_ ;
	wire _w337_ ;
	wire _w338_ ;
	wire _w339_ ;
	wire _w340_ ;
	wire _w341_ ;
	wire _w342_ ;
	wire _w343_ ;
	wire _w344_ ;
	wire _w345_ ;
	wire _w346_ ;
	wire _w347_ ;
	wire _w348_ ;
	wire _w349_ ;
	wire _w350_ ;
	wire _w351_ ;
	wire _w352_ ;
	wire _w353_ ;
	wire _w354_ ;
	wire _w355_ ;
	wire _w356_ ;
	wire _w357_ ;
	wire _w358_ ;
	wire _w359_ ;
	wire _w360_ ;
	wire _w361_ ;
	wire _w362_ ;
	wire _w363_ ;
	wire _w364_ ;
	wire _w365_ ;
	wire _w366_ ;
	wire _w367_ ;
	wire _w368_ ;
	wire _w369_ ;
	wire _w370_ ;
	wire _w371_ ;
	wire _w372_ ;
	wire _w373_ ;
	wire _w374_ ;
	wire _w375_ ;
	wire _w376_ ;
	wire _w377_ ;
	wire _w378_ ;
	wire _w379_ ;
	wire _w380_ ;
	wire _w381_ ;
	wire _w382_ ;
	wire _w383_ ;
	wire _w384_ ;
	wire _w385_ ;
	wire _w386_ ;
	wire _w387_ ;
	wire _w388_ ;
	wire _w389_ ;
	wire _w390_ ;
	wire _w391_ ;
	wire _w392_ ;
	wire _w393_ ;
	wire _w394_ ;
	wire _w395_ ;
	wire _w396_ ;
	wire _w397_ ;
	wire _w398_ ;
	wire _w399_ ;
	wire _w400_ ;
	wire _w401_ ;
	wire _w402_ ;
	wire _w403_ ;
	wire _w404_ ;
	wire _w405_ ;
	wire _w406_ ;
	wire _w407_ ;
	wire _w408_ ;
	wire _w409_ ;
	wire _w410_ ;
	wire _w411_ ;
	wire _w412_ ;
	wire _w413_ ;
	wire _w414_ ;
	wire _w415_ ;
	wire _w416_ ;
	wire _w417_ ;
	wire _w418_ ;
	wire _w419_ ;
	wire _w420_ ;
	wire _w421_ ;
	wire _w422_ ;
	wire _w423_ ;
	wire _w424_ ;
	wire _w425_ ;
	wire _w426_ ;
	wire _w427_ ;
	wire _w428_ ;
	wire _w429_ ;
	wire _w430_ ;
	wire _w431_ ;
	wire _w432_ ;
	wire _w433_ ;
	wire _w434_ ;
	wire _w435_ ;
	wire _w436_ ;
	wire _w437_ ;
	wire _w438_ ;
	wire _w439_ ;
	wire _w440_ ;
	wire _w441_ ;
	wire _w442_ ;
	wire _w443_ ;
	wire _w444_ ;
	wire _w445_ ;
	wire _w446_ ;
	wire _w447_ ;
	wire _w448_ ;
	wire _w449_ ;
	wire _w450_ ;
	wire _w451_ ;
	wire _w452_ ;
	wire _w453_ ;
	wire _w454_ ;
	wire _w455_ ;
	wire _w456_ ;
	wire _w457_ ;
	wire _w458_ ;
	wire _w459_ ;
	wire _w460_ ;
	wire _w461_ ;
	wire _w462_ ;
	wire _w463_ ;
	wire _w464_ ;
	wire _w465_ ;
	wire _w466_ ;
	wire _w467_ ;
	wire _w468_ ;
	wire _w469_ ;
	wire _w470_ ;
	wire _w471_ ;
	wire _w472_ ;
	wire _w473_ ;
	wire _w474_ ;
	wire _w475_ ;
	wire _w476_ ;
	wire _w477_ ;
	wire _w478_ ;
	wire _w479_ ;
	wire _w480_ ;
	wire _w481_ ;
	wire _w482_ ;
	wire _w483_ ;
	wire _w484_ ;
	wire _w485_ ;
	wire _w486_ ;
	wire _w487_ ;
	wire _w488_ ;
	wire _w489_ ;
	wire _w490_ ;
	wire _w491_ ;
	wire _w492_ ;
	wire _w493_ ;
	wire _w494_ ;
	wire _w495_ ;
	wire _w496_ ;
	wire _w497_ ;
	wire _w498_ ;
	wire _w499_ ;
	wire _w500_ ;
	wire _w501_ ;
	wire _w502_ ;
	wire _w503_ ;
	wire _w504_ ;
	wire _w505_ ;
	wire _w506_ ;
	wire _w507_ ;
	wire _w508_ ;
	wire _w509_ ;
	wire _w510_ ;
	wire _w511_ ;
	wire _w512_ ;
	wire _w513_ ;
	wire _w514_ ;
	wire _w515_ ;
	wire _w516_ ;
	wire _w517_ ;
	wire _w518_ ;
	wire _w519_ ;
	wire _w520_ ;
	wire _w521_ ;
	wire _w522_ ;
	wire _w523_ ;
	wire _w524_ ;
	wire _w525_ ;
	wire _w526_ ;
	wire _w527_ ;
	wire _w528_ ;
	wire _w529_ ;
	wire _w530_ ;
	wire _w531_ ;
	wire _w532_ ;
	wire _w533_ ;
	wire _w534_ ;
	wire _w535_ ;
	wire _w536_ ;
	wire _w537_ ;
	wire _w538_ ;
	wire _w539_ ;
	wire _w540_ ;
	wire _w541_ ;
	wire _w542_ ;
	wire _w543_ ;
	wire _w544_ ;
	wire _w545_ ;
	wire _w546_ ;
	wire _w547_ ;
	wire _w548_ ;
	wire _w549_ ;
	wire _w550_ ;
	wire _w551_ ;
	wire _w552_ ;
	wire _w553_ ;
	wire _w554_ ;
	wire _w555_ ;
	wire _w556_ ;
	wire _w557_ ;
	wire _w558_ ;
	wire _w559_ ;
	wire _w560_ ;
	wire _w561_ ;
	wire _w562_ ;
	wire _w563_ ;
	wire _w564_ ;
	wire _w565_ ;
	wire _w566_ ;
	wire _w567_ ;
	wire _w568_ ;
	wire _w569_ ;
	wire _w570_ ;
	wire _w571_ ;
	wire _w572_ ;
	wire _w573_ ;
	wire _w574_ ;
	LUT4 #(
		.INIT('h8000)
	) name0 (
		\18GAT(1)_pad ,
		\1GAT(0)_pad ,
		\273GAT(16)_pad ,
		\290GAT(17)_pad ,
		_w34_
	);
	LUT4 #(
		.INIT('h6ca0)
	) name1 (
		\18GAT(1)_pad ,
		\1GAT(0)_pad ,
		\273GAT(16)_pad ,
		\290GAT(17)_pad ,
		_w35_
	);
	LUT2 #(
		.INIT('h8)
	) name2 (
		\1GAT(0)_pad ,
		\307GAT(18)_pad ,
		_w36_
	);
	LUT2 #(
		.INIT('h4)
	) name3 (
		\35GAT(2)_pad ,
		_w34_,
		_w37_
	);
	LUT2 #(
		.INIT('h8)
	) name4 (
		\18GAT(1)_pad ,
		\290GAT(17)_pad ,
		_w38_
	);
	LUT2 #(
		.INIT('h8)
	) name5 (
		\273GAT(16)_pad ,
		\35GAT(2)_pad ,
		_w39_
	);
	LUT3 #(
		.INIT('h43)
	) name6 (
		\1GAT(0)_pad ,
		_w38_,
		_w39_,
		_w40_
	);
	LUT3 #(
		.INIT('ha9)
	) name7 (
		_w36_,
		_w37_,
		_w40_,
		_w41_
	);
	LUT2 #(
		.INIT('h8)
	) name8 (
		\1GAT(0)_pad ,
		\324GAT(19)_pad ,
		_w42_
	);
	LUT3 #(
		.INIT('h0e)
	) name9 (
		_w36_,
		_w37_,
		_w40_,
		_w43_
	);
	LUT2 #(
		.INIT('h8)
	) name10 (
		\18GAT(1)_pad ,
		\307GAT(18)_pad ,
		_w44_
	);
	LUT3 #(
		.INIT('h08)
	) name11 (
		\18GAT(1)_pad ,
		\273GAT(16)_pad ,
		\52GAT(3)_pad ,
		_w45_
	);
	LUT2 #(
		.INIT('h8)
	) name12 (
		\273GAT(16)_pad ,
		\52GAT(3)_pad ,
		_w46_
	);
	LUT2 #(
		.INIT('h8)
	) name13 (
		\290GAT(17)_pad ,
		\35GAT(2)_pad ,
		_w47_
	);
	LUT3 #(
		.INIT('hbc)
	) name14 (
		\18GAT(1)_pad ,
		_w46_,
		_w47_,
		_w48_
	);
	LUT4 #(
		.INIT('hb7c0)
	) name15 (
		\18GAT(1)_pad ,
		\273GAT(16)_pad ,
		\52GAT(3)_pad ,
		_w47_,
		_w49_
	);
	LUT2 #(
		.INIT('h9)
	) name16 (
		_w44_,
		_w49_,
		_w50_
	);
	LUT3 #(
		.INIT('h69)
	) name17 (
		_w42_,
		_w43_,
		_w50_,
		_w51_
	);
	LUT2 #(
		.INIT('h8)
	) name18 (
		\1GAT(0)_pad ,
		\341GAT(20)_pad ,
		_w52_
	);
	LUT3 #(
		.INIT('h8e)
	) name19 (
		_w42_,
		_w43_,
		_w50_,
		_w53_
	);
	LUT2 #(
		.INIT('h8)
	) name20 (
		\18GAT(1)_pad ,
		\324GAT(19)_pad ,
		_w54_
	);
	LUT3 #(
		.INIT('he0)
	) name21 (
		_w44_,
		_w45_,
		_w48_,
		_w55_
	);
	LUT2 #(
		.INIT('h8)
	) name22 (
		\307GAT(18)_pad ,
		\35GAT(2)_pad ,
		_w56_
	);
	LUT3 #(
		.INIT('h08)
	) name23 (
		\273GAT(16)_pad ,
		\35GAT(2)_pad ,
		\69GAT(4)_pad ,
		_w57_
	);
	LUT2 #(
		.INIT('h8)
	) name24 (
		\273GAT(16)_pad ,
		\69GAT(4)_pad ,
		_w58_
	);
	LUT2 #(
		.INIT('h8)
	) name25 (
		\290GAT(17)_pad ,
		\52GAT(3)_pad ,
		_w59_
	);
	LUT3 #(
		.INIT('hbc)
	) name26 (
		\35GAT(2)_pad ,
		_w58_,
		_w59_,
		_w60_
	);
	LUT4 #(
		.INIT('hd7a0)
	) name27 (
		\273GAT(16)_pad ,
		\35GAT(2)_pad ,
		\69GAT(4)_pad ,
		_w59_,
		_w61_
	);
	LUT2 #(
		.INIT('h9)
	) name28 (
		_w56_,
		_w61_,
		_w62_
	);
	LUT3 #(
		.INIT('h96)
	) name29 (
		_w54_,
		_w55_,
		_w62_,
		_w63_
	);
	LUT3 #(
		.INIT('h69)
	) name30 (
		_w52_,
		_w53_,
		_w63_,
		_w64_
	);
	LUT2 #(
		.INIT('h8)
	) name31 (
		\1GAT(0)_pad ,
		\358GAT(21)_pad ,
		_w65_
	);
	LUT3 #(
		.INIT('h8e)
	) name32 (
		_w52_,
		_w53_,
		_w63_,
		_w66_
	);
	LUT2 #(
		.INIT('h8)
	) name33 (
		\18GAT(1)_pad ,
		\341GAT(20)_pad ,
		_w67_
	);
	LUT3 #(
		.INIT('h8e)
	) name34 (
		_w54_,
		_w55_,
		_w62_,
		_w68_
	);
	LUT2 #(
		.INIT('h8)
	) name35 (
		\324GAT(19)_pad ,
		\35GAT(2)_pad ,
		_w69_
	);
	LUT3 #(
		.INIT('he0)
	) name36 (
		_w56_,
		_w57_,
		_w60_,
		_w70_
	);
	LUT2 #(
		.INIT('h8)
	) name37 (
		\307GAT(18)_pad ,
		\52GAT(3)_pad ,
		_w71_
	);
	LUT3 #(
		.INIT('h08)
	) name38 (
		\273GAT(16)_pad ,
		\52GAT(3)_pad ,
		\86GAT(5)_pad ,
		_w72_
	);
	LUT4 #(
		.INIT('h153f)
	) name39 (
		\273GAT(16)_pad ,
		\290GAT(17)_pad ,
		\69GAT(4)_pad ,
		\86GAT(5)_pad ,
		_w73_
	);
	LUT4 #(
		.INIT('h8000)
	) name40 (
		\273GAT(16)_pad ,
		\290GAT(17)_pad ,
		\69GAT(4)_pad ,
		\86GAT(5)_pad ,
		_w74_
	);
	LUT3 #(
		.INIT('h23)
	) name41 (
		\52GAT(3)_pad ,
		_w73_,
		_w74_,
		_w75_
	);
	LUT4 #(
		.INIT('h0203)
	) name42 (
		\52GAT(3)_pad ,
		_w72_,
		_w73_,
		_w74_,
		_w76_
	);
	LUT2 #(
		.INIT('h9)
	) name43 (
		_w71_,
		_w76_,
		_w77_
	);
	LUT3 #(
		.INIT('h96)
	) name44 (
		_w69_,
		_w70_,
		_w77_,
		_w78_
	);
	LUT3 #(
		.INIT('h96)
	) name45 (
		_w67_,
		_w68_,
		_w78_,
		_w79_
	);
	LUT3 #(
		.INIT('h69)
	) name46 (
		_w65_,
		_w66_,
		_w79_,
		_w80_
	);
	LUT2 #(
		.INIT('h8)
	) name47 (
		\1GAT(0)_pad ,
		\375GAT(22)_pad ,
		_w81_
	);
	LUT3 #(
		.INIT('h8e)
	) name48 (
		_w65_,
		_w66_,
		_w79_,
		_w82_
	);
	LUT2 #(
		.INIT('h8)
	) name49 (
		\18GAT(1)_pad ,
		\358GAT(21)_pad ,
		_w83_
	);
	LUT3 #(
		.INIT('h8e)
	) name50 (
		_w67_,
		_w68_,
		_w78_,
		_w84_
	);
	LUT2 #(
		.INIT('h8)
	) name51 (
		\341GAT(20)_pad ,
		\35GAT(2)_pad ,
		_w85_
	);
	LUT3 #(
		.INIT('h8e)
	) name52 (
		_w69_,
		_w70_,
		_w77_,
		_w86_
	);
	LUT2 #(
		.INIT('h8)
	) name53 (
		\324GAT(19)_pad ,
		\52GAT(3)_pad ,
		_w87_
	);
	LUT2 #(
		.INIT('h8)
	) name54 (
		\307GAT(18)_pad ,
		\69GAT(4)_pad ,
		_w88_
	);
	LUT4 #(
		.INIT('h8000)
	) name55 (
		\103GAT(6)_pad ,
		\273GAT(16)_pad ,
		\290GAT(17)_pad ,
		\86GAT(5)_pad ,
		_w89_
	);
	LUT4 #(
		.INIT('h7888)
	) name56 (
		\103GAT(6)_pad ,
		\273GAT(16)_pad ,
		\290GAT(17)_pad ,
		\86GAT(5)_pad ,
		_w90_
	);
	LUT3 #(
		.INIT('h69)
	) name57 (
		_w74_,
		_w88_,
		_w90_,
		_w91_
	);
	LUT4 #(
		.INIT('h7300)
	) name58 (
		_w71_,
		_w75_,
		_w76_,
		_w91_,
		_w92_
	);
	LUT4 #(
		.INIT('h008c)
	) name59 (
		_w71_,
		_w75_,
		_w76_,
		_w91_,
		_w93_
	);
	LUT4 #(
		.INIT('he01f)
	) name60 (
		_w71_,
		_w72_,
		_w75_,
		_w91_,
		_w94_
	);
	LUT2 #(
		.INIT('h9)
	) name61 (
		_w87_,
		_w94_,
		_w95_
	);
	LUT3 #(
		.INIT('h96)
	) name62 (
		_w85_,
		_w86_,
		_w95_,
		_w96_
	);
	LUT3 #(
		.INIT('h96)
	) name63 (
		_w83_,
		_w84_,
		_w96_,
		_w97_
	);
	LUT3 #(
		.INIT('h69)
	) name64 (
		_w81_,
		_w82_,
		_w97_,
		_w98_
	);
	LUT2 #(
		.INIT('h8)
	) name65 (
		\1GAT(0)_pad ,
		\392GAT(23)_pad ,
		_w99_
	);
	LUT3 #(
		.INIT('h8e)
	) name66 (
		_w81_,
		_w82_,
		_w97_,
		_w100_
	);
	LUT2 #(
		.INIT('h8)
	) name67 (
		\18GAT(1)_pad ,
		\375GAT(22)_pad ,
		_w101_
	);
	LUT3 #(
		.INIT('h8e)
	) name68 (
		_w83_,
		_w84_,
		_w96_,
		_w102_
	);
	LUT2 #(
		.INIT('h8)
	) name69 (
		\358GAT(21)_pad ,
		\35GAT(2)_pad ,
		_w103_
	);
	LUT3 #(
		.INIT('h8e)
	) name70 (
		_w85_,
		_w86_,
		_w95_,
		_w104_
	);
	LUT2 #(
		.INIT('h8)
	) name71 (
		\341GAT(20)_pad ,
		\52GAT(3)_pad ,
		_w105_
	);
	LUT3 #(
		.INIT('h32)
	) name72 (
		_w87_,
		_w92_,
		_w93_,
		_w106_
	);
	LUT2 #(
		.INIT('h8)
	) name73 (
		\324GAT(19)_pad ,
		\69GAT(4)_pad ,
		_w107_
	);
	LUT3 #(
		.INIT('he8)
	) name74 (
		_w74_,
		_w88_,
		_w90_,
		_w108_
	);
	LUT2 #(
		.INIT('h8)
	) name75 (
		\307GAT(18)_pad ,
		\86GAT(5)_pad ,
		_w109_
	);
	LUT2 #(
		.INIT('h4)
	) name76 (
		\120GAT(7)_pad ,
		_w89_,
		_w110_
	);
	LUT2 #(
		.INIT('h8)
	) name77 (
		\103GAT(6)_pad ,
		\290GAT(17)_pad ,
		_w111_
	);
	LUT2 #(
		.INIT('h8)
	) name78 (
		\120GAT(7)_pad ,
		\273GAT(16)_pad ,
		_w112_
	);
	LUT3 #(
		.INIT('h43)
	) name79 (
		\86GAT(5)_pad ,
		_w111_,
		_w112_,
		_w113_
	);
	LUT4 #(
		.INIT('h1114)
	) name80 (
		_w108_,
		_w109_,
		_w110_,
		_w113_,
		_w114_
	);
	LUT4 #(
		.INIT('h8882)
	) name81 (
		_w108_,
		_w109_,
		_w110_,
		_w113_,
		_w115_
	);
	LUT4 #(
		.INIT('h6669)
	) name82 (
		_w108_,
		_w109_,
		_w110_,
		_w113_,
		_w116_
	);
	LUT2 #(
		.INIT('h9)
	) name83 (
		_w107_,
		_w116_,
		_w117_
	);
	LUT3 #(
		.INIT('h96)
	) name84 (
		_w105_,
		_w106_,
		_w117_,
		_w118_
	);
	LUT3 #(
		.INIT('h96)
	) name85 (
		_w103_,
		_w104_,
		_w118_,
		_w119_
	);
	LUT3 #(
		.INIT('h96)
	) name86 (
		_w101_,
		_w102_,
		_w119_,
		_w120_
	);
	LUT3 #(
		.INIT('h69)
	) name87 (
		_w99_,
		_w100_,
		_w120_,
		_w121_
	);
	LUT2 #(
		.INIT('h8)
	) name88 (
		\1GAT(0)_pad ,
		\409GAT(24)_pad ,
		_w122_
	);
	LUT3 #(
		.INIT('h8e)
	) name89 (
		_w99_,
		_w100_,
		_w120_,
		_w123_
	);
	LUT2 #(
		.INIT('h8)
	) name90 (
		\18GAT(1)_pad ,
		\392GAT(23)_pad ,
		_w124_
	);
	LUT3 #(
		.INIT('h8e)
	) name91 (
		_w101_,
		_w102_,
		_w119_,
		_w125_
	);
	LUT2 #(
		.INIT('h8)
	) name92 (
		\35GAT(2)_pad ,
		\375GAT(22)_pad ,
		_w126_
	);
	LUT3 #(
		.INIT('h8e)
	) name93 (
		_w103_,
		_w104_,
		_w118_,
		_w127_
	);
	LUT2 #(
		.INIT('h8)
	) name94 (
		\358GAT(21)_pad ,
		\52GAT(3)_pad ,
		_w128_
	);
	LUT3 #(
		.INIT('h8e)
	) name95 (
		_w105_,
		_w106_,
		_w117_,
		_w129_
	);
	LUT2 #(
		.INIT('h8)
	) name96 (
		\341GAT(20)_pad ,
		\69GAT(4)_pad ,
		_w130_
	);
	LUT3 #(
		.INIT('h32)
	) name97 (
		_w107_,
		_w114_,
		_w115_,
		_w131_
	);
	LUT2 #(
		.INIT('h8)
	) name98 (
		\324GAT(19)_pad ,
		\86GAT(5)_pad ,
		_w132_
	);
	LUT3 #(
		.INIT('h0e)
	) name99 (
		_w109_,
		_w110_,
		_w113_,
		_w133_
	);
	LUT2 #(
		.INIT('h8)
	) name100 (
		\103GAT(6)_pad ,
		\307GAT(18)_pad ,
		_w134_
	);
	LUT3 #(
		.INIT('h20)
	) name101 (
		\103GAT(6)_pad ,
		\137GAT(8)_pad ,
		\273GAT(16)_pad ,
		_w135_
	);
	LUT2 #(
		.INIT('h8)
	) name102 (
		\137GAT(8)_pad ,
		\273GAT(16)_pad ,
		_w136_
	);
	LUT2 #(
		.INIT('h8)
	) name103 (
		\120GAT(7)_pad ,
		\290GAT(17)_pad ,
		_w137_
	);
	LUT3 #(
		.INIT('hbc)
	) name104 (
		\103GAT(6)_pad ,
		_w136_,
		_w137_,
		_w138_
	);
	LUT4 #(
		.INIT('h9fc0)
	) name105 (
		\103GAT(6)_pad ,
		\137GAT(8)_pad ,
		\273GAT(16)_pad ,
		_w137_,
		_w139_
	);
	LUT2 #(
		.INIT('h9)
	) name106 (
		_w134_,
		_w139_,
		_w140_
	);
	LUT3 #(
		.INIT('h96)
	) name107 (
		_w132_,
		_w133_,
		_w140_,
		_w141_
	);
	LUT3 #(
		.INIT('h96)
	) name108 (
		_w130_,
		_w131_,
		_w141_,
		_w142_
	);
	LUT3 #(
		.INIT('h96)
	) name109 (
		_w128_,
		_w129_,
		_w142_,
		_w143_
	);
	LUT3 #(
		.INIT('h96)
	) name110 (
		_w126_,
		_w127_,
		_w143_,
		_w144_
	);
	LUT3 #(
		.INIT('h96)
	) name111 (
		_w124_,
		_w125_,
		_w144_,
		_w145_
	);
	LUT3 #(
		.INIT('h69)
	) name112 (
		_w122_,
		_w123_,
		_w145_,
		_w146_
	);
	LUT2 #(
		.INIT('h8)
	) name113 (
		\1GAT(0)_pad ,
		\426GAT(25)_pad ,
		_w147_
	);
	LUT3 #(
		.INIT('h8e)
	) name114 (
		_w122_,
		_w123_,
		_w145_,
		_w148_
	);
	LUT2 #(
		.INIT('h8)
	) name115 (
		\18GAT(1)_pad ,
		\409GAT(24)_pad ,
		_w149_
	);
	LUT3 #(
		.INIT('h8e)
	) name116 (
		_w124_,
		_w125_,
		_w144_,
		_w150_
	);
	LUT2 #(
		.INIT('h8)
	) name117 (
		\35GAT(2)_pad ,
		\392GAT(23)_pad ,
		_w151_
	);
	LUT3 #(
		.INIT('h8e)
	) name118 (
		_w126_,
		_w127_,
		_w143_,
		_w152_
	);
	LUT2 #(
		.INIT('h8)
	) name119 (
		\375GAT(22)_pad ,
		\52GAT(3)_pad ,
		_w153_
	);
	LUT3 #(
		.INIT('h8e)
	) name120 (
		_w128_,
		_w129_,
		_w142_,
		_w154_
	);
	LUT2 #(
		.INIT('h8)
	) name121 (
		\358GAT(21)_pad ,
		\69GAT(4)_pad ,
		_w155_
	);
	LUT3 #(
		.INIT('h8e)
	) name122 (
		_w130_,
		_w131_,
		_w141_,
		_w156_
	);
	LUT2 #(
		.INIT('h8)
	) name123 (
		\341GAT(20)_pad ,
		\86GAT(5)_pad ,
		_w157_
	);
	LUT3 #(
		.INIT('h8e)
	) name124 (
		_w132_,
		_w133_,
		_w140_,
		_w158_
	);
	LUT2 #(
		.INIT('h8)
	) name125 (
		\103GAT(6)_pad ,
		\324GAT(19)_pad ,
		_w159_
	);
	LUT3 #(
		.INIT('he0)
	) name126 (
		_w134_,
		_w135_,
		_w138_,
		_w160_
	);
	LUT2 #(
		.INIT('h8)
	) name127 (
		\120GAT(7)_pad ,
		\307GAT(18)_pad ,
		_w161_
	);
	LUT3 #(
		.INIT('h20)
	) name128 (
		\120GAT(7)_pad ,
		\154GAT(9)_pad ,
		\273GAT(16)_pad ,
		_w162_
	);
	LUT2 #(
		.INIT('h8)
	) name129 (
		\154GAT(9)_pad ,
		\273GAT(16)_pad ,
		_w163_
	);
	LUT2 #(
		.INIT('h8)
	) name130 (
		\137GAT(8)_pad ,
		\290GAT(17)_pad ,
		_w164_
	);
	LUT3 #(
		.INIT('hbc)
	) name131 (
		\120GAT(7)_pad ,
		_w163_,
		_w164_,
		_w165_
	);
	LUT4 #(
		.INIT('h9fc0)
	) name132 (
		\120GAT(7)_pad ,
		\154GAT(9)_pad ,
		\273GAT(16)_pad ,
		_w164_,
		_w166_
	);
	LUT2 #(
		.INIT('h9)
	) name133 (
		_w161_,
		_w166_,
		_w167_
	);
	LUT3 #(
		.INIT('h96)
	) name134 (
		_w159_,
		_w160_,
		_w167_,
		_w168_
	);
	LUT3 #(
		.INIT('h96)
	) name135 (
		_w157_,
		_w158_,
		_w168_,
		_w169_
	);
	LUT3 #(
		.INIT('h96)
	) name136 (
		_w155_,
		_w156_,
		_w169_,
		_w170_
	);
	LUT3 #(
		.INIT('h96)
	) name137 (
		_w153_,
		_w154_,
		_w170_,
		_w171_
	);
	LUT3 #(
		.INIT('h96)
	) name138 (
		_w151_,
		_w152_,
		_w171_,
		_w172_
	);
	LUT3 #(
		.INIT('h96)
	) name139 (
		_w149_,
		_w150_,
		_w172_,
		_w173_
	);
	LUT3 #(
		.INIT('h69)
	) name140 (
		_w147_,
		_w148_,
		_w173_,
		_w174_
	);
	LUT2 #(
		.INIT('h8)
	) name141 (
		\1GAT(0)_pad ,
		\443GAT(26)_pad ,
		_w175_
	);
	LUT3 #(
		.INIT('h8e)
	) name142 (
		_w147_,
		_w148_,
		_w173_,
		_w176_
	);
	LUT2 #(
		.INIT('h8)
	) name143 (
		\18GAT(1)_pad ,
		\426GAT(25)_pad ,
		_w177_
	);
	LUT3 #(
		.INIT('h8e)
	) name144 (
		_w149_,
		_w150_,
		_w172_,
		_w178_
	);
	LUT2 #(
		.INIT('h8)
	) name145 (
		\35GAT(2)_pad ,
		\409GAT(24)_pad ,
		_w179_
	);
	LUT3 #(
		.INIT('h8e)
	) name146 (
		_w151_,
		_w152_,
		_w171_,
		_w180_
	);
	LUT2 #(
		.INIT('h8)
	) name147 (
		\392GAT(23)_pad ,
		\52GAT(3)_pad ,
		_w181_
	);
	LUT3 #(
		.INIT('h8e)
	) name148 (
		_w153_,
		_w154_,
		_w170_,
		_w182_
	);
	LUT2 #(
		.INIT('h8)
	) name149 (
		\375GAT(22)_pad ,
		\69GAT(4)_pad ,
		_w183_
	);
	LUT3 #(
		.INIT('h8e)
	) name150 (
		_w155_,
		_w156_,
		_w169_,
		_w184_
	);
	LUT2 #(
		.INIT('h8)
	) name151 (
		\358GAT(21)_pad ,
		\86GAT(5)_pad ,
		_w185_
	);
	LUT3 #(
		.INIT('h8e)
	) name152 (
		_w157_,
		_w158_,
		_w168_,
		_w186_
	);
	LUT2 #(
		.INIT('h8)
	) name153 (
		\103GAT(6)_pad ,
		\341GAT(20)_pad ,
		_w187_
	);
	LUT3 #(
		.INIT('h8e)
	) name154 (
		_w159_,
		_w160_,
		_w167_,
		_w188_
	);
	LUT2 #(
		.INIT('h8)
	) name155 (
		\120GAT(7)_pad ,
		\324GAT(19)_pad ,
		_w189_
	);
	LUT3 #(
		.INIT('he0)
	) name156 (
		_w161_,
		_w162_,
		_w165_,
		_w190_
	);
	LUT2 #(
		.INIT('h8)
	) name157 (
		\137GAT(8)_pad ,
		\307GAT(18)_pad ,
		_w191_
	);
	LUT3 #(
		.INIT('h20)
	) name158 (
		\137GAT(8)_pad ,
		\171GAT(10)_pad ,
		\273GAT(16)_pad ,
		_w192_
	);
	LUT2 #(
		.INIT('h8)
	) name159 (
		\171GAT(10)_pad ,
		\273GAT(16)_pad ,
		_w193_
	);
	LUT2 #(
		.INIT('h8)
	) name160 (
		\154GAT(9)_pad ,
		\290GAT(17)_pad ,
		_w194_
	);
	LUT3 #(
		.INIT('hbc)
	) name161 (
		\137GAT(8)_pad ,
		_w193_,
		_w194_,
		_w195_
	);
	LUT4 #(
		.INIT('h9fc0)
	) name162 (
		\137GAT(8)_pad ,
		\171GAT(10)_pad ,
		\273GAT(16)_pad ,
		_w194_,
		_w196_
	);
	LUT2 #(
		.INIT('h9)
	) name163 (
		_w191_,
		_w196_,
		_w197_
	);
	LUT3 #(
		.INIT('h96)
	) name164 (
		_w189_,
		_w190_,
		_w197_,
		_w198_
	);
	LUT3 #(
		.INIT('h96)
	) name165 (
		_w187_,
		_w188_,
		_w198_,
		_w199_
	);
	LUT3 #(
		.INIT('h96)
	) name166 (
		_w185_,
		_w186_,
		_w199_,
		_w200_
	);
	LUT3 #(
		.INIT('h96)
	) name167 (
		_w183_,
		_w184_,
		_w200_,
		_w201_
	);
	LUT3 #(
		.INIT('h96)
	) name168 (
		_w181_,
		_w182_,
		_w201_,
		_w202_
	);
	LUT3 #(
		.INIT('h96)
	) name169 (
		_w179_,
		_w180_,
		_w202_,
		_w203_
	);
	LUT3 #(
		.INIT('h96)
	) name170 (
		_w177_,
		_w178_,
		_w203_,
		_w204_
	);
	LUT3 #(
		.INIT('h69)
	) name171 (
		_w175_,
		_w176_,
		_w204_,
		_w205_
	);
	LUT2 #(
		.INIT('h8)
	) name172 (
		\1GAT(0)_pad ,
		\460GAT(27)_pad ,
		_w206_
	);
	LUT3 #(
		.INIT('h8e)
	) name173 (
		_w175_,
		_w176_,
		_w204_,
		_w207_
	);
	LUT2 #(
		.INIT('h8)
	) name174 (
		\18GAT(1)_pad ,
		\443GAT(26)_pad ,
		_w208_
	);
	LUT3 #(
		.INIT('h8e)
	) name175 (
		_w177_,
		_w178_,
		_w203_,
		_w209_
	);
	LUT2 #(
		.INIT('h8)
	) name176 (
		\35GAT(2)_pad ,
		\426GAT(25)_pad ,
		_w210_
	);
	LUT3 #(
		.INIT('h8e)
	) name177 (
		_w179_,
		_w180_,
		_w202_,
		_w211_
	);
	LUT2 #(
		.INIT('h8)
	) name178 (
		\409GAT(24)_pad ,
		\52GAT(3)_pad ,
		_w212_
	);
	LUT3 #(
		.INIT('h8e)
	) name179 (
		_w181_,
		_w182_,
		_w201_,
		_w213_
	);
	LUT2 #(
		.INIT('h8)
	) name180 (
		\392GAT(23)_pad ,
		\69GAT(4)_pad ,
		_w214_
	);
	LUT3 #(
		.INIT('h8e)
	) name181 (
		_w183_,
		_w184_,
		_w200_,
		_w215_
	);
	LUT2 #(
		.INIT('h8)
	) name182 (
		\375GAT(22)_pad ,
		\86GAT(5)_pad ,
		_w216_
	);
	LUT3 #(
		.INIT('h8e)
	) name183 (
		_w185_,
		_w186_,
		_w199_,
		_w217_
	);
	LUT2 #(
		.INIT('h8)
	) name184 (
		\103GAT(6)_pad ,
		\358GAT(21)_pad ,
		_w218_
	);
	LUT3 #(
		.INIT('h8e)
	) name185 (
		_w187_,
		_w188_,
		_w198_,
		_w219_
	);
	LUT2 #(
		.INIT('h8)
	) name186 (
		\120GAT(7)_pad ,
		\341GAT(20)_pad ,
		_w220_
	);
	LUT3 #(
		.INIT('h8e)
	) name187 (
		_w189_,
		_w190_,
		_w197_,
		_w221_
	);
	LUT2 #(
		.INIT('h8)
	) name188 (
		\137GAT(8)_pad ,
		\324GAT(19)_pad ,
		_w222_
	);
	LUT3 #(
		.INIT('he0)
	) name189 (
		_w191_,
		_w192_,
		_w195_,
		_w223_
	);
	LUT2 #(
		.INIT('h8)
	) name190 (
		\154GAT(9)_pad ,
		\307GAT(18)_pad ,
		_w224_
	);
	LUT3 #(
		.INIT('h20)
	) name191 (
		\154GAT(9)_pad ,
		\188GAT(11)_pad ,
		\273GAT(16)_pad ,
		_w225_
	);
	LUT2 #(
		.INIT('h8)
	) name192 (
		\188GAT(11)_pad ,
		\273GAT(16)_pad ,
		_w226_
	);
	LUT2 #(
		.INIT('h8)
	) name193 (
		\171GAT(10)_pad ,
		\290GAT(17)_pad ,
		_w227_
	);
	LUT3 #(
		.INIT('hbc)
	) name194 (
		\154GAT(9)_pad ,
		_w226_,
		_w227_,
		_w228_
	);
	LUT4 #(
		.INIT('h9fc0)
	) name195 (
		\154GAT(9)_pad ,
		\188GAT(11)_pad ,
		\273GAT(16)_pad ,
		_w227_,
		_w229_
	);
	LUT2 #(
		.INIT('h9)
	) name196 (
		_w224_,
		_w229_,
		_w230_
	);
	LUT3 #(
		.INIT('h96)
	) name197 (
		_w222_,
		_w223_,
		_w230_,
		_w231_
	);
	LUT3 #(
		.INIT('h96)
	) name198 (
		_w220_,
		_w221_,
		_w231_,
		_w232_
	);
	LUT3 #(
		.INIT('h96)
	) name199 (
		_w218_,
		_w219_,
		_w232_,
		_w233_
	);
	LUT3 #(
		.INIT('h96)
	) name200 (
		_w216_,
		_w217_,
		_w233_,
		_w234_
	);
	LUT3 #(
		.INIT('h96)
	) name201 (
		_w214_,
		_w215_,
		_w234_,
		_w235_
	);
	LUT3 #(
		.INIT('h96)
	) name202 (
		_w212_,
		_w213_,
		_w235_,
		_w236_
	);
	LUT3 #(
		.INIT('h96)
	) name203 (
		_w210_,
		_w211_,
		_w236_,
		_w237_
	);
	LUT3 #(
		.INIT('h96)
	) name204 (
		_w208_,
		_w209_,
		_w237_,
		_w238_
	);
	LUT3 #(
		.INIT('h69)
	) name205 (
		_w206_,
		_w207_,
		_w238_,
		_w239_
	);
	LUT2 #(
		.INIT('h8)
	) name206 (
		\1GAT(0)_pad ,
		\477GAT(28)_pad ,
		_w240_
	);
	LUT3 #(
		.INIT('h8e)
	) name207 (
		_w206_,
		_w207_,
		_w238_,
		_w241_
	);
	LUT2 #(
		.INIT('h8)
	) name208 (
		\18GAT(1)_pad ,
		\460GAT(27)_pad ,
		_w242_
	);
	LUT3 #(
		.INIT('h8e)
	) name209 (
		_w208_,
		_w209_,
		_w237_,
		_w243_
	);
	LUT2 #(
		.INIT('h8)
	) name210 (
		\35GAT(2)_pad ,
		\443GAT(26)_pad ,
		_w244_
	);
	LUT3 #(
		.INIT('h8e)
	) name211 (
		_w210_,
		_w211_,
		_w236_,
		_w245_
	);
	LUT2 #(
		.INIT('h8)
	) name212 (
		\426GAT(25)_pad ,
		\52GAT(3)_pad ,
		_w246_
	);
	LUT3 #(
		.INIT('h8e)
	) name213 (
		_w212_,
		_w213_,
		_w235_,
		_w247_
	);
	LUT2 #(
		.INIT('h8)
	) name214 (
		\409GAT(24)_pad ,
		\69GAT(4)_pad ,
		_w248_
	);
	LUT3 #(
		.INIT('h8e)
	) name215 (
		_w214_,
		_w215_,
		_w234_,
		_w249_
	);
	LUT2 #(
		.INIT('h8)
	) name216 (
		\392GAT(23)_pad ,
		\86GAT(5)_pad ,
		_w250_
	);
	LUT3 #(
		.INIT('h8e)
	) name217 (
		_w216_,
		_w217_,
		_w233_,
		_w251_
	);
	LUT2 #(
		.INIT('h8)
	) name218 (
		\103GAT(6)_pad ,
		\375GAT(22)_pad ,
		_w252_
	);
	LUT3 #(
		.INIT('h8e)
	) name219 (
		_w218_,
		_w219_,
		_w232_,
		_w253_
	);
	LUT2 #(
		.INIT('h8)
	) name220 (
		\120GAT(7)_pad ,
		\358GAT(21)_pad ,
		_w254_
	);
	LUT3 #(
		.INIT('h8e)
	) name221 (
		_w220_,
		_w221_,
		_w231_,
		_w255_
	);
	LUT2 #(
		.INIT('h8)
	) name222 (
		\137GAT(8)_pad ,
		\341GAT(20)_pad ,
		_w256_
	);
	LUT3 #(
		.INIT('h8e)
	) name223 (
		_w222_,
		_w223_,
		_w230_,
		_w257_
	);
	LUT2 #(
		.INIT('h8)
	) name224 (
		\154GAT(9)_pad ,
		\324GAT(19)_pad ,
		_w258_
	);
	LUT3 #(
		.INIT('he0)
	) name225 (
		_w224_,
		_w225_,
		_w228_,
		_w259_
	);
	LUT2 #(
		.INIT('h8)
	) name226 (
		\171GAT(10)_pad ,
		\307GAT(18)_pad ,
		_w260_
	);
	LUT3 #(
		.INIT('h20)
	) name227 (
		\171GAT(10)_pad ,
		\205GAT(12)_pad ,
		\273GAT(16)_pad ,
		_w261_
	);
	LUT2 #(
		.INIT('h8)
	) name228 (
		\205GAT(12)_pad ,
		\273GAT(16)_pad ,
		_w262_
	);
	LUT2 #(
		.INIT('h8)
	) name229 (
		\188GAT(11)_pad ,
		\290GAT(17)_pad ,
		_w263_
	);
	LUT3 #(
		.INIT('hbc)
	) name230 (
		\171GAT(10)_pad ,
		_w262_,
		_w263_,
		_w264_
	);
	LUT4 #(
		.INIT('h9fc0)
	) name231 (
		\171GAT(10)_pad ,
		\205GAT(12)_pad ,
		\273GAT(16)_pad ,
		_w263_,
		_w265_
	);
	LUT2 #(
		.INIT('h9)
	) name232 (
		_w260_,
		_w265_,
		_w266_
	);
	LUT3 #(
		.INIT('h96)
	) name233 (
		_w258_,
		_w259_,
		_w266_,
		_w267_
	);
	LUT3 #(
		.INIT('h96)
	) name234 (
		_w256_,
		_w257_,
		_w267_,
		_w268_
	);
	LUT3 #(
		.INIT('h96)
	) name235 (
		_w254_,
		_w255_,
		_w268_,
		_w269_
	);
	LUT3 #(
		.INIT('h96)
	) name236 (
		_w252_,
		_w253_,
		_w269_,
		_w270_
	);
	LUT3 #(
		.INIT('h96)
	) name237 (
		_w250_,
		_w251_,
		_w270_,
		_w271_
	);
	LUT3 #(
		.INIT('h96)
	) name238 (
		_w248_,
		_w249_,
		_w271_,
		_w272_
	);
	LUT3 #(
		.INIT('h96)
	) name239 (
		_w246_,
		_w247_,
		_w272_,
		_w273_
	);
	LUT3 #(
		.INIT('h96)
	) name240 (
		_w244_,
		_w245_,
		_w273_,
		_w274_
	);
	LUT3 #(
		.INIT('h96)
	) name241 (
		_w242_,
		_w243_,
		_w274_,
		_w275_
	);
	LUT3 #(
		.INIT('h69)
	) name242 (
		_w240_,
		_w241_,
		_w275_,
		_w276_
	);
	LUT2 #(
		.INIT('h8)
	) name243 (
		\1GAT(0)_pad ,
		\273GAT(16)_pad ,
		_w277_
	);
	LUT2 #(
		.INIT('h8)
	) name244 (
		\1GAT(0)_pad ,
		\494GAT(29)_pad ,
		_w278_
	);
	LUT3 #(
		.INIT('h8e)
	) name245 (
		_w240_,
		_w241_,
		_w275_,
		_w279_
	);
	LUT2 #(
		.INIT('h8)
	) name246 (
		\18GAT(1)_pad ,
		\477GAT(28)_pad ,
		_w280_
	);
	LUT3 #(
		.INIT('h8e)
	) name247 (
		_w242_,
		_w243_,
		_w274_,
		_w281_
	);
	LUT2 #(
		.INIT('h8)
	) name248 (
		\35GAT(2)_pad ,
		\460GAT(27)_pad ,
		_w282_
	);
	LUT3 #(
		.INIT('h8e)
	) name249 (
		_w244_,
		_w245_,
		_w273_,
		_w283_
	);
	LUT2 #(
		.INIT('h8)
	) name250 (
		\443GAT(26)_pad ,
		\52GAT(3)_pad ,
		_w284_
	);
	LUT3 #(
		.INIT('h8e)
	) name251 (
		_w246_,
		_w247_,
		_w272_,
		_w285_
	);
	LUT2 #(
		.INIT('h8)
	) name252 (
		\426GAT(25)_pad ,
		\69GAT(4)_pad ,
		_w286_
	);
	LUT3 #(
		.INIT('h8e)
	) name253 (
		_w248_,
		_w249_,
		_w271_,
		_w287_
	);
	LUT2 #(
		.INIT('h8)
	) name254 (
		\409GAT(24)_pad ,
		\86GAT(5)_pad ,
		_w288_
	);
	LUT3 #(
		.INIT('h8e)
	) name255 (
		_w250_,
		_w251_,
		_w270_,
		_w289_
	);
	LUT2 #(
		.INIT('h8)
	) name256 (
		\103GAT(6)_pad ,
		\392GAT(23)_pad ,
		_w290_
	);
	LUT3 #(
		.INIT('h8e)
	) name257 (
		_w252_,
		_w253_,
		_w269_,
		_w291_
	);
	LUT2 #(
		.INIT('h8)
	) name258 (
		\120GAT(7)_pad ,
		\375GAT(22)_pad ,
		_w292_
	);
	LUT3 #(
		.INIT('h8e)
	) name259 (
		_w254_,
		_w255_,
		_w268_,
		_w293_
	);
	LUT2 #(
		.INIT('h8)
	) name260 (
		\137GAT(8)_pad ,
		\358GAT(21)_pad ,
		_w294_
	);
	LUT3 #(
		.INIT('h8e)
	) name261 (
		_w256_,
		_w257_,
		_w267_,
		_w295_
	);
	LUT2 #(
		.INIT('h8)
	) name262 (
		\154GAT(9)_pad ,
		\341GAT(20)_pad ,
		_w296_
	);
	LUT3 #(
		.INIT('h8e)
	) name263 (
		_w258_,
		_w259_,
		_w266_,
		_w297_
	);
	LUT2 #(
		.INIT('h8)
	) name264 (
		\171GAT(10)_pad ,
		\324GAT(19)_pad ,
		_w298_
	);
	LUT3 #(
		.INIT('he0)
	) name265 (
		_w260_,
		_w261_,
		_w264_,
		_w299_
	);
	LUT2 #(
		.INIT('h8)
	) name266 (
		\188GAT(11)_pad ,
		\307GAT(18)_pad ,
		_w300_
	);
	LUT3 #(
		.INIT('h20)
	) name267 (
		\188GAT(11)_pad ,
		\222GAT(13)_pad ,
		\273GAT(16)_pad ,
		_w301_
	);
	LUT2 #(
		.INIT('h8)
	) name268 (
		\222GAT(13)_pad ,
		\273GAT(16)_pad ,
		_w302_
	);
	LUT2 #(
		.INIT('h8)
	) name269 (
		\205GAT(12)_pad ,
		\290GAT(17)_pad ,
		_w303_
	);
	LUT3 #(
		.INIT('hbc)
	) name270 (
		\188GAT(11)_pad ,
		_w302_,
		_w303_,
		_w304_
	);
	LUT4 #(
		.INIT('h9fc0)
	) name271 (
		\188GAT(11)_pad ,
		\222GAT(13)_pad ,
		\273GAT(16)_pad ,
		_w303_,
		_w305_
	);
	LUT2 #(
		.INIT('h9)
	) name272 (
		_w300_,
		_w305_,
		_w306_
	);
	LUT3 #(
		.INIT('h96)
	) name273 (
		_w298_,
		_w299_,
		_w306_,
		_w307_
	);
	LUT3 #(
		.INIT('h96)
	) name274 (
		_w296_,
		_w297_,
		_w307_,
		_w308_
	);
	LUT3 #(
		.INIT('h96)
	) name275 (
		_w294_,
		_w295_,
		_w308_,
		_w309_
	);
	LUT3 #(
		.INIT('h96)
	) name276 (
		_w292_,
		_w293_,
		_w309_,
		_w310_
	);
	LUT3 #(
		.INIT('h96)
	) name277 (
		_w290_,
		_w291_,
		_w310_,
		_w311_
	);
	LUT3 #(
		.INIT('h96)
	) name278 (
		_w288_,
		_w289_,
		_w311_,
		_w312_
	);
	LUT3 #(
		.INIT('h96)
	) name279 (
		_w286_,
		_w287_,
		_w312_,
		_w313_
	);
	LUT3 #(
		.INIT('h96)
	) name280 (
		_w284_,
		_w285_,
		_w313_,
		_w314_
	);
	LUT3 #(
		.INIT('h96)
	) name281 (
		_w282_,
		_w283_,
		_w314_,
		_w315_
	);
	LUT3 #(
		.INIT('h96)
	) name282 (
		_w280_,
		_w281_,
		_w315_,
		_w316_
	);
	LUT3 #(
		.INIT('h69)
	) name283 (
		_w278_,
		_w279_,
		_w316_,
		_w317_
	);
	LUT2 #(
		.INIT('h8)
	) name284 (
		\1GAT(0)_pad ,
		\511GAT(30)_pad ,
		_w318_
	);
	LUT3 #(
		.INIT('h8e)
	) name285 (
		_w278_,
		_w279_,
		_w316_,
		_w319_
	);
	LUT2 #(
		.INIT('h8)
	) name286 (
		\18GAT(1)_pad ,
		\494GAT(29)_pad ,
		_w320_
	);
	LUT3 #(
		.INIT('h8e)
	) name287 (
		_w280_,
		_w281_,
		_w315_,
		_w321_
	);
	LUT2 #(
		.INIT('h8)
	) name288 (
		\35GAT(2)_pad ,
		\477GAT(28)_pad ,
		_w322_
	);
	LUT3 #(
		.INIT('h8e)
	) name289 (
		_w282_,
		_w283_,
		_w314_,
		_w323_
	);
	LUT2 #(
		.INIT('h8)
	) name290 (
		\460GAT(27)_pad ,
		\52GAT(3)_pad ,
		_w324_
	);
	LUT3 #(
		.INIT('h8e)
	) name291 (
		_w284_,
		_w285_,
		_w313_,
		_w325_
	);
	LUT2 #(
		.INIT('h8)
	) name292 (
		\443GAT(26)_pad ,
		\69GAT(4)_pad ,
		_w326_
	);
	LUT3 #(
		.INIT('h8e)
	) name293 (
		_w286_,
		_w287_,
		_w312_,
		_w327_
	);
	LUT2 #(
		.INIT('h8)
	) name294 (
		\426GAT(25)_pad ,
		\86GAT(5)_pad ,
		_w328_
	);
	LUT3 #(
		.INIT('h8e)
	) name295 (
		_w288_,
		_w289_,
		_w311_,
		_w329_
	);
	LUT2 #(
		.INIT('h8)
	) name296 (
		\103GAT(6)_pad ,
		\409GAT(24)_pad ,
		_w330_
	);
	LUT3 #(
		.INIT('h8e)
	) name297 (
		_w290_,
		_w291_,
		_w310_,
		_w331_
	);
	LUT2 #(
		.INIT('h8)
	) name298 (
		\120GAT(7)_pad ,
		\392GAT(23)_pad ,
		_w332_
	);
	LUT3 #(
		.INIT('h8e)
	) name299 (
		_w292_,
		_w293_,
		_w309_,
		_w333_
	);
	LUT2 #(
		.INIT('h8)
	) name300 (
		\137GAT(8)_pad ,
		\375GAT(22)_pad ,
		_w334_
	);
	LUT3 #(
		.INIT('h8e)
	) name301 (
		_w294_,
		_w295_,
		_w308_,
		_w335_
	);
	LUT2 #(
		.INIT('h8)
	) name302 (
		\154GAT(9)_pad ,
		\358GAT(21)_pad ,
		_w336_
	);
	LUT3 #(
		.INIT('h8e)
	) name303 (
		_w296_,
		_w297_,
		_w307_,
		_w337_
	);
	LUT2 #(
		.INIT('h8)
	) name304 (
		\171GAT(10)_pad ,
		\341GAT(20)_pad ,
		_w338_
	);
	LUT3 #(
		.INIT('h8e)
	) name305 (
		_w298_,
		_w299_,
		_w306_,
		_w339_
	);
	LUT2 #(
		.INIT('h8)
	) name306 (
		\188GAT(11)_pad ,
		\324GAT(19)_pad ,
		_w340_
	);
	LUT3 #(
		.INIT('he0)
	) name307 (
		_w300_,
		_w301_,
		_w304_,
		_w341_
	);
	LUT2 #(
		.INIT('h8)
	) name308 (
		\205GAT(12)_pad ,
		\307GAT(18)_pad ,
		_w342_
	);
	LUT3 #(
		.INIT('h20)
	) name309 (
		\205GAT(12)_pad ,
		\239GAT(14)_pad ,
		\273GAT(16)_pad ,
		_w343_
	);
	LUT2 #(
		.INIT('h8)
	) name310 (
		\239GAT(14)_pad ,
		\273GAT(16)_pad ,
		_w344_
	);
	LUT2 #(
		.INIT('h8)
	) name311 (
		\222GAT(13)_pad ,
		\290GAT(17)_pad ,
		_w345_
	);
	LUT3 #(
		.INIT('hbc)
	) name312 (
		\205GAT(12)_pad ,
		_w344_,
		_w345_,
		_w346_
	);
	LUT4 #(
		.INIT('h9fc0)
	) name313 (
		\205GAT(12)_pad ,
		\239GAT(14)_pad ,
		\273GAT(16)_pad ,
		_w345_,
		_w347_
	);
	LUT2 #(
		.INIT('h9)
	) name314 (
		_w342_,
		_w347_,
		_w348_
	);
	LUT3 #(
		.INIT('h96)
	) name315 (
		_w340_,
		_w341_,
		_w348_,
		_w349_
	);
	LUT3 #(
		.INIT('h96)
	) name316 (
		_w338_,
		_w339_,
		_w349_,
		_w350_
	);
	LUT3 #(
		.INIT('h96)
	) name317 (
		_w336_,
		_w337_,
		_w350_,
		_w351_
	);
	LUT3 #(
		.INIT('h96)
	) name318 (
		_w334_,
		_w335_,
		_w351_,
		_w352_
	);
	LUT3 #(
		.INIT('h96)
	) name319 (
		_w332_,
		_w333_,
		_w352_,
		_w353_
	);
	LUT3 #(
		.INIT('h96)
	) name320 (
		_w330_,
		_w331_,
		_w353_,
		_w354_
	);
	LUT3 #(
		.INIT('h96)
	) name321 (
		_w328_,
		_w329_,
		_w354_,
		_w355_
	);
	LUT3 #(
		.INIT('h96)
	) name322 (
		_w326_,
		_w327_,
		_w355_,
		_w356_
	);
	LUT3 #(
		.INIT('h96)
	) name323 (
		_w324_,
		_w325_,
		_w356_,
		_w357_
	);
	LUT3 #(
		.INIT('h96)
	) name324 (
		_w322_,
		_w323_,
		_w357_,
		_w358_
	);
	LUT3 #(
		.INIT('h96)
	) name325 (
		_w320_,
		_w321_,
		_w358_,
		_w359_
	);
	LUT3 #(
		.INIT('h69)
	) name326 (
		_w318_,
		_w319_,
		_w359_,
		_w360_
	);
	LUT2 #(
		.INIT('h8)
	) name327 (
		\1GAT(0)_pad ,
		\528GAT(31)_pad ,
		_w361_
	);
	LUT3 #(
		.INIT('h8e)
	) name328 (
		_w318_,
		_w319_,
		_w359_,
		_w362_
	);
	LUT2 #(
		.INIT('h8)
	) name329 (
		\18GAT(1)_pad ,
		\511GAT(30)_pad ,
		_w363_
	);
	LUT3 #(
		.INIT('h8e)
	) name330 (
		_w320_,
		_w321_,
		_w358_,
		_w364_
	);
	LUT2 #(
		.INIT('h8)
	) name331 (
		\35GAT(2)_pad ,
		\494GAT(29)_pad ,
		_w365_
	);
	LUT3 #(
		.INIT('h8e)
	) name332 (
		_w322_,
		_w323_,
		_w357_,
		_w366_
	);
	LUT2 #(
		.INIT('h8)
	) name333 (
		\477GAT(28)_pad ,
		\52GAT(3)_pad ,
		_w367_
	);
	LUT3 #(
		.INIT('h8e)
	) name334 (
		_w324_,
		_w325_,
		_w356_,
		_w368_
	);
	LUT2 #(
		.INIT('h8)
	) name335 (
		\460GAT(27)_pad ,
		\69GAT(4)_pad ,
		_w369_
	);
	LUT3 #(
		.INIT('h8e)
	) name336 (
		_w326_,
		_w327_,
		_w355_,
		_w370_
	);
	LUT2 #(
		.INIT('h8)
	) name337 (
		\443GAT(26)_pad ,
		\86GAT(5)_pad ,
		_w371_
	);
	LUT3 #(
		.INIT('h8e)
	) name338 (
		_w328_,
		_w329_,
		_w354_,
		_w372_
	);
	LUT2 #(
		.INIT('h8)
	) name339 (
		\103GAT(6)_pad ,
		\426GAT(25)_pad ,
		_w373_
	);
	LUT3 #(
		.INIT('h8e)
	) name340 (
		_w330_,
		_w331_,
		_w353_,
		_w374_
	);
	LUT2 #(
		.INIT('h8)
	) name341 (
		\120GAT(7)_pad ,
		\409GAT(24)_pad ,
		_w375_
	);
	LUT3 #(
		.INIT('h8e)
	) name342 (
		_w332_,
		_w333_,
		_w352_,
		_w376_
	);
	LUT2 #(
		.INIT('h8)
	) name343 (
		\137GAT(8)_pad ,
		\392GAT(23)_pad ,
		_w377_
	);
	LUT3 #(
		.INIT('h8e)
	) name344 (
		_w334_,
		_w335_,
		_w351_,
		_w378_
	);
	LUT2 #(
		.INIT('h8)
	) name345 (
		\154GAT(9)_pad ,
		\375GAT(22)_pad ,
		_w379_
	);
	LUT3 #(
		.INIT('h8e)
	) name346 (
		_w336_,
		_w337_,
		_w350_,
		_w380_
	);
	LUT2 #(
		.INIT('h8)
	) name347 (
		\171GAT(10)_pad ,
		\358GAT(21)_pad ,
		_w381_
	);
	LUT3 #(
		.INIT('h8e)
	) name348 (
		_w338_,
		_w339_,
		_w349_,
		_w382_
	);
	LUT2 #(
		.INIT('h8)
	) name349 (
		\188GAT(11)_pad ,
		\341GAT(20)_pad ,
		_w383_
	);
	LUT3 #(
		.INIT('h8e)
	) name350 (
		_w340_,
		_w341_,
		_w348_,
		_w384_
	);
	LUT2 #(
		.INIT('h8)
	) name351 (
		\205GAT(12)_pad ,
		\324GAT(19)_pad ,
		_w385_
	);
	LUT3 #(
		.INIT('he0)
	) name352 (
		_w342_,
		_w343_,
		_w346_,
		_w386_
	);
	LUT2 #(
		.INIT('h8)
	) name353 (
		\222GAT(13)_pad ,
		\307GAT(18)_pad ,
		_w387_
	);
	LUT3 #(
		.INIT('h20)
	) name354 (
		\222GAT(13)_pad ,
		\256GAT(15)_pad ,
		\273GAT(16)_pad ,
		_w388_
	);
	LUT2 #(
		.INIT('h8)
	) name355 (
		\256GAT(15)_pad ,
		\273GAT(16)_pad ,
		_w389_
	);
	LUT2 #(
		.INIT('h8)
	) name356 (
		\239GAT(14)_pad ,
		\290GAT(17)_pad ,
		_w390_
	);
	LUT3 #(
		.INIT('hbc)
	) name357 (
		\222GAT(13)_pad ,
		_w389_,
		_w390_,
		_w391_
	);
	LUT4 #(
		.INIT('h9fc0)
	) name358 (
		\222GAT(13)_pad ,
		\256GAT(15)_pad ,
		\273GAT(16)_pad ,
		_w390_,
		_w392_
	);
	LUT2 #(
		.INIT('h9)
	) name359 (
		_w387_,
		_w392_,
		_w393_
	);
	LUT3 #(
		.INIT('h96)
	) name360 (
		_w385_,
		_w386_,
		_w393_,
		_w394_
	);
	LUT3 #(
		.INIT('h96)
	) name361 (
		_w383_,
		_w384_,
		_w394_,
		_w395_
	);
	LUT3 #(
		.INIT('h96)
	) name362 (
		_w381_,
		_w382_,
		_w395_,
		_w396_
	);
	LUT3 #(
		.INIT('h96)
	) name363 (
		_w379_,
		_w380_,
		_w396_,
		_w397_
	);
	LUT3 #(
		.INIT('h96)
	) name364 (
		_w377_,
		_w378_,
		_w397_,
		_w398_
	);
	LUT3 #(
		.INIT('h96)
	) name365 (
		_w375_,
		_w376_,
		_w398_,
		_w399_
	);
	LUT3 #(
		.INIT('h96)
	) name366 (
		_w373_,
		_w374_,
		_w399_,
		_w400_
	);
	LUT3 #(
		.INIT('h96)
	) name367 (
		_w371_,
		_w372_,
		_w400_,
		_w401_
	);
	LUT3 #(
		.INIT('h96)
	) name368 (
		_w369_,
		_w370_,
		_w401_,
		_w402_
	);
	LUT3 #(
		.INIT('h96)
	) name369 (
		_w367_,
		_w368_,
		_w402_,
		_w403_
	);
	LUT3 #(
		.INIT('h96)
	) name370 (
		_w365_,
		_w366_,
		_w403_,
		_w404_
	);
	LUT3 #(
		.INIT('h96)
	) name371 (
		_w363_,
		_w364_,
		_w404_,
		_w405_
	);
	LUT3 #(
		.INIT('h69)
	) name372 (
		_w361_,
		_w362_,
		_w405_,
		_w406_
	);
	LUT3 #(
		.INIT('h8e)
	) name373 (
		_w361_,
		_w362_,
		_w405_,
		_w407_
	);
	LUT2 #(
		.INIT('h8)
	) name374 (
		\18GAT(1)_pad ,
		\528GAT(31)_pad ,
		_w408_
	);
	LUT3 #(
		.INIT('h8e)
	) name375 (
		_w363_,
		_w364_,
		_w404_,
		_w409_
	);
	LUT2 #(
		.INIT('h8)
	) name376 (
		\35GAT(2)_pad ,
		\511GAT(30)_pad ,
		_w410_
	);
	LUT3 #(
		.INIT('h8e)
	) name377 (
		_w365_,
		_w366_,
		_w403_,
		_w411_
	);
	LUT2 #(
		.INIT('h8)
	) name378 (
		\494GAT(29)_pad ,
		\52GAT(3)_pad ,
		_w412_
	);
	LUT3 #(
		.INIT('h8e)
	) name379 (
		_w367_,
		_w368_,
		_w402_,
		_w413_
	);
	LUT2 #(
		.INIT('h8)
	) name380 (
		\477GAT(28)_pad ,
		\69GAT(4)_pad ,
		_w414_
	);
	LUT3 #(
		.INIT('h8e)
	) name381 (
		_w369_,
		_w370_,
		_w401_,
		_w415_
	);
	LUT2 #(
		.INIT('h8)
	) name382 (
		\460GAT(27)_pad ,
		\86GAT(5)_pad ,
		_w416_
	);
	LUT3 #(
		.INIT('h8e)
	) name383 (
		_w371_,
		_w372_,
		_w400_,
		_w417_
	);
	LUT2 #(
		.INIT('h8)
	) name384 (
		\103GAT(6)_pad ,
		\443GAT(26)_pad ,
		_w418_
	);
	LUT3 #(
		.INIT('h8e)
	) name385 (
		_w373_,
		_w374_,
		_w399_,
		_w419_
	);
	LUT2 #(
		.INIT('h8)
	) name386 (
		\120GAT(7)_pad ,
		\426GAT(25)_pad ,
		_w420_
	);
	LUT3 #(
		.INIT('h8e)
	) name387 (
		_w375_,
		_w376_,
		_w398_,
		_w421_
	);
	LUT2 #(
		.INIT('h8)
	) name388 (
		\137GAT(8)_pad ,
		\409GAT(24)_pad ,
		_w422_
	);
	LUT3 #(
		.INIT('h8e)
	) name389 (
		_w377_,
		_w378_,
		_w397_,
		_w423_
	);
	LUT2 #(
		.INIT('h8)
	) name390 (
		\154GAT(9)_pad ,
		\392GAT(23)_pad ,
		_w424_
	);
	LUT3 #(
		.INIT('h8e)
	) name391 (
		_w379_,
		_w380_,
		_w396_,
		_w425_
	);
	LUT2 #(
		.INIT('h8)
	) name392 (
		\171GAT(10)_pad ,
		\375GAT(22)_pad ,
		_w426_
	);
	LUT3 #(
		.INIT('h8e)
	) name393 (
		_w381_,
		_w382_,
		_w395_,
		_w427_
	);
	LUT2 #(
		.INIT('h8)
	) name394 (
		\188GAT(11)_pad ,
		\358GAT(21)_pad ,
		_w428_
	);
	LUT3 #(
		.INIT('h8e)
	) name395 (
		_w383_,
		_w384_,
		_w394_,
		_w429_
	);
	LUT2 #(
		.INIT('h8)
	) name396 (
		\205GAT(12)_pad ,
		\341GAT(20)_pad ,
		_w430_
	);
	LUT3 #(
		.INIT('h8e)
	) name397 (
		_w385_,
		_w386_,
		_w393_,
		_w431_
	);
	LUT2 #(
		.INIT('h8)
	) name398 (
		\222GAT(13)_pad ,
		\324GAT(19)_pad ,
		_w432_
	);
	LUT3 #(
		.INIT('he0)
	) name399 (
		_w387_,
		_w388_,
		_w391_,
		_w433_
	);
	LUT2 #(
		.INIT('h8)
	) name400 (
		\239GAT(14)_pad ,
		\307GAT(18)_pad ,
		_w434_
	);
	LUT4 #(
		.INIT('h4c00)
	) name401 (
		\239GAT(14)_pad ,
		\256GAT(15)_pad ,
		\273GAT(16)_pad ,
		\290GAT(17)_pad ,
		_w435_
	);
	LUT2 #(
		.INIT('h9)
	) name402 (
		_w434_,
		_w435_,
		_w436_
	);
	LUT4 #(
		.INIT('h7300)
	) name403 (
		_w387_,
		_w391_,
		_w392_,
		_w436_,
		_w437_
	);
	LUT4 #(
		.INIT('h008c)
	) name404 (
		_w387_,
		_w391_,
		_w392_,
		_w436_,
		_w438_
	);
	LUT4 #(
		.INIT('he01f)
	) name405 (
		_w387_,
		_w388_,
		_w391_,
		_w436_,
		_w439_
	);
	LUT2 #(
		.INIT('h9)
	) name406 (
		_w432_,
		_w439_,
		_w440_
	);
	LUT3 #(
		.INIT('h96)
	) name407 (
		_w430_,
		_w431_,
		_w440_,
		_w441_
	);
	LUT3 #(
		.INIT('h96)
	) name408 (
		_w428_,
		_w429_,
		_w441_,
		_w442_
	);
	LUT3 #(
		.INIT('h96)
	) name409 (
		_w426_,
		_w427_,
		_w442_,
		_w443_
	);
	LUT3 #(
		.INIT('h96)
	) name410 (
		_w424_,
		_w425_,
		_w443_,
		_w444_
	);
	LUT3 #(
		.INIT('h96)
	) name411 (
		_w422_,
		_w423_,
		_w444_,
		_w445_
	);
	LUT3 #(
		.INIT('h96)
	) name412 (
		_w420_,
		_w421_,
		_w445_,
		_w446_
	);
	LUT3 #(
		.INIT('h96)
	) name413 (
		_w418_,
		_w419_,
		_w446_,
		_w447_
	);
	LUT3 #(
		.INIT('h96)
	) name414 (
		_w416_,
		_w417_,
		_w447_,
		_w448_
	);
	LUT3 #(
		.INIT('h96)
	) name415 (
		_w414_,
		_w415_,
		_w448_,
		_w449_
	);
	LUT3 #(
		.INIT('h96)
	) name416 (
		_w412_,
		_w413_,
		_w449_,
		_w450_
	);
	LUT3 #(
		.INIT('h96)
	) name417 (
		_w410_,
		_w411_,
		_w450_,
		_w451_
	);
	LUT3 #(
		.INIT('h96)
	) name418 (
		_w408_,
		_w409_,
		_w451_,
		_w452_
	);
	LUT2 #(
		.INIT('h9)
	) name419 (
		_w407_,
		_w452_,
		_w453_
	);
	LUT3 #(
		.INIT('h8e)
	) name420 (
		_w408_,
		_w409_,
		_w451_,
		_w454_
	);
	LUT2 #(
		.INIT('h8)
	) name421 (
		\35GAT(2)_pad ,
		\528GAT(31)_pad ,
		_w455_
	);
	LUT3 #(
		.INIT('h8e)
	) name422 (
		_w410_,
		_w411_,
		_w450_,
		_w456_
	);
	LUT2 #(
		.INIT('h8)
	) name423 (
		\511GAT(30)_pad ,
		\52GAT(3)_pad ,
		_w457_
	);
	LUT3 #(
		.INIT('h8e)
	) name424 (
		_w412_,
		_w413_,
		_w449_,
		_w458_
	);
	LUT2 #(
		.INIT('h8)
	) name425 (
		\494GAT(29)_pad ,
		\69GAT(4)_pad ,
		_w459_
	);
	LUT3 #(
		.INIT('h8e)
	) name426 (
		_w414_,
		_w415_,
		_w448_,
		_w460_
	);
	LUT2 #(
		.INIT('h8)
	) name427 (
		\477GAT(28)_pad ,
		\86GAT(5)_pad ,
		_w461_
	);
	LUT3 #(
		.INIT('h8e)
	) name428 (
		_w416_,
		_w417_,
		_w447_,
		_w462_
	);
	LUT2 #(
		.INIT('h8)
	) name429 (
		\103GAT(6)_pad ,
		\460GAT(27)_pad ,
		_w463_
	);
	LUT3 #(
		.INIT('h8e)
	) name430 (
		_w418_,
		_w419_,
		_w446_,
		_w464_
	);
	LUT2 #(
		.INIT('h8)
	) name431 (
		\120GAT(7)_pad ,
		\443GAT(26)_pad ,
		_w465_
	);
	LUT3 #(
		.INIT('h8e)
	) name432 (
		_w420_,
		_w421_,
		_w445_,
		_w466_
	);
	LUT2 #(
		.INIT('h8)
	) name433 (
		\137GAT(8)_pad ,
		\426GAT(25)_pad ,
		_w467_
	);
	LUT3 #(
		.INIT('h8e)
	) name434 (
		_w422_,
		_w423_,
		_w444_,
		_w468_
	);
	LUT2 #(
		.INIT('h8)
	) name435 (
		\154GAT(9)_pad ,
		\409GAT(24)_pad ,
		_w469_
	);
	LUT3 #(
		.INIT('h8e)
	) name436 (
		_w424_,
		_w425_,
		_w443_,
		_w470_
	);
	LUT2 #(
		.INIT('h8)
	) name437 (
		\171GAT(10)_pad ,
		\392GAT(23)_pad ,
		_w471_
	);
	LUT3 #(
		.INIT('h8e)
	) name438 (
		_w426_,
		_w427_,
		_w442_,
		_w472_
	);
	LUT2 #(
		.INIT('h8)
	) name439 (
		\188GAT(11)_pad ,
		\375GAT(22)_pad ,
		_w473_
	);
	LUT3 #(
		.INIT('h8e)
	) name440 (
		_w428_,
		_w429_,
		_w441_,
		_w474_
	);
	LUT2 #(
		.INIT('h8)
	) name441 (
		\205GAT(12)_pad ,
		\358GAT(21)_pad ,
		_w475_
	);
	LUT3 #(
		.INIT('h8e)
	) name442 (
		_w430_,
		_w431_,
		_w440_,
		_w476_
	);
	LUT2 #(
		.INIT('h8)
	) name443 (
		\222GAT(13)_pad ,
		\341GAT(20)_pad ,
		_w477_
	);
	LUT3 #(
		.INIT('h32)
	) name444 (
		_w432_,
		_w437_,
		_w438_,
		_w478_
	);
	LUT2 #(
		.INIT('h8)
	) name445 (
		\239GAT(14)_pad ,
		\324GAT(19)_pad ,
		_w479_
	);
	LUT4 #(
		.INIT('h007f)
	) name446 (
		\239GAT(14)_pad ,
		\273GAT(16)_pad ,
		\290GAT(17)_pad ,
		\307GAT(18)_pad ,
		_w480_
	);
	LUT3 #(
		.INIT('h80)
	) name447 (
		\239GAT(14)_pad ,
		\290GAT(17)_pad ,
		\307GAT(18)_pad ,
		_w481_
	);
	LUT4 #(
		.INIT('h3339)
	) name448 (
		\256GAT(15)_pad ,
		_w479_,
		_w480_,
		_w481_,
		_w482_
	);
	LUT4 #(
		.INIT('h7100)
	) name449 (
		_w432_,
		_w433_,
		_w436_,
		_w482_,
		_w483_
	);
	LUT4 #(
		.INIT('h008e)
	) name450 (
		_w432_,
		_w433_,
		_w436_,
		_w482_,
		_w484_
	);
	LUT4 #(
		.INIT('h32cd)
	) name451 (
		_w432_,
		_w437_,
		_w438_,
		_w482_,
		_w485_
	);
	LUT2 #(
		.INIT('h9)
	) name452 (
		_w477_,
		_w485_,
		_w486_
	);
	LUT3 #(
		.INIT('h96)
	) name453 (
		_w475_,
		_w476_,
		_w486_,
		_w487_
	);
	LUT3 #(
		.INIT('h96)
	) name454 (
		_w473_,
		_w474_,
		_w487_,
		_w488_
	);
	LUT3 #(
		.INIT('h96)
	) name455 (
		_w471_,
		_w472_,
		_w488_,
		_w489_
	);
	LUT3 #(
		.INIT('h96)
	) name456 (
		_w469_,
		_w470_,
		_w489_,
		_w490_
	);
	LUT3 #(
		.INIT('h96)
	) name457 (
		_w467_,
		_w468_,
		_w490_,
		_w491_
	);
	LUT3 #(
		.INIT('h96)
	) name458 (
		_w465_,
		_w466_,
		_w491_,
		_w492_
	);
	LUT3 #(
		.INIT('h96)
	) name459 (
		_w463_,
		_w464_,
		_w492_,
		_w493_
	);
	LUT3 #(
		.INIT('h96)
	) name460 (
		_w461_,
		_w462_,
		_w493_,
		_w494_
	);
	LUT3 #(
		.INIT('h96)
	) name461 (
		_w459_,
		_w460_,
		_w494_,
		_w495_
	);
	LUT3 #(
		.INIT('h96)
	) name462 (
		_w457_,
		_w458_,
		_w495_,
		_w496_
	);
	LUT3 #(
		.INIT('h96)
	) name463 (
		_w455_,
		_w456_,
		_w496_,
		_w497_
	);
	LUT4 #(
		.INIT('hd22d)
	) name464 (
		_w407_,
		_w452_,
		_w454_,
		_w497_,
		_w498_
	);
	LUT4 #(
		.INIT('h20f2)
	) name465 (
		_w407_,
		_w452_,
		_w454_,
		_w497_,
		_w499_
	);
	LUT3 #(
		.INIT('h8e)
	) name466 (
		_w455_,
		_w456_,
		_w496_,
		_w500_
	);
	LUT2 #(
		.INIT('h8)
	) name467 (
		\528GAT(31)_pad ,
		\52GAT(3)_pad ,
		_w501_
	);
	LUT3 #(
		.INIT('h8e)
	) name468 (
		_w457_,
		_w458_,
		_w495_,
		_w502_
	);
	LUT2 #(
		.INIT('h8)
	) name469 (
		\511GAT(30)_pad ,
		\69GAT(4)_pad ,
		_w503_
	);
	LUT3 #(
		.INIT('h8e)
	) name470 (
		_w459_,
		_w460_,
		_w494_,
		_w504_
	);
	LUT2 #(
		.INIT('h8)
	) name471 (
		\494GAT(29)_pad ,
		\86GAT(5)_pad ,
		_w505_
	);
	LUT3 #(
		.INIT('h8e)
	) name472 (
		_w461_,
		_w462_,
		_w493_,
		_w506_
	);
	LUT2 #(
		.INIT('h8)
	) name473 (
		\103GAT(6)_pad ,
		\477GAT(28)_pad ,
		_w507_
	);
	LUT3 #(
		.INIT('h8e)
	) name474 (
		_w463_,
		_w464_,
		_w492_,
		_w508_
	);
	LUT2 #(
		.INIT('h8)
	) name475 (
		\120GAT(7)_pad ,
		\460GAT(27)_pad ,
		_w509_
	);
	LUT3 #(
		.INIT('h8e)
	) name476 (
		_w465_,
		_w466_,
		_w491_,
		_w510_
	);
	LUT2 #(
		.INIT('h8)
	) name477 (
		\137GAT(8)_pad ,
		\443GAT(26)_pad ,
		_w511_
	);
	LUT3 #(
		.INIT('h8e)
	) name478 (
		_w467_,
		_w468_,
		_w490_,
		_w512_
	);
	LUT2 #(
		.INIT('h8)
	) name479 (
		\154GAT(9)_pad ,
		\426GAT(25)_pad ,
		_w513_
	);
	LUT3 #(
		.INIT('h8e)
	) name480 (
		_w469_,
		_w470_,
		_w489_,
		_w514_
	);
	LUT2 #(
		.INIT('h8)
	) name481 (
		\171GAT(10)_pad ,
		\409GAT(24)_pad ,
		_w515_
	);
	LUT3 #(
		.INIT('h8e)
	) name482 (
		_w471_,
		_w472_,
		_w488_,
		_w516_
	);
	LUT2 #(
		.INIT('h8)
	) name483 (
		\188GAT(11)_pad ,
		\392GAT(23)_pad ,
		_w517_
	);
	LUT3 #(
		.INIT('h8e)
	) name484 (
		_w473_,
		_w474_,
		_w487_,
		_w518_
	);
	LUT2 #(
		.INIT('h8)
	) name485 (
		\205GAT(12)_pad ,
		\375GAT(22)_pad ,
		_w519_
	);
	LUT3 #(
		.INIT('h8e)
	) name486 (
		_w475_,
		_w476_,
		_w486_,
		_w520_
	);
	LUT2 #(
		.INIT('h8)
	) name487 (
		\222GAT(13)_pad ,
		\358GAT(21)_pad ,
		_w521_
	);
	LUT3 #(
		.INIT('h32)
	) name488 (
		_w477_,
		_w483_,
		_w484_,
		_w522_
	);
	LUT2 #(
		.INIT('h8)
	) name489 (
		\239GAT(14)_pad ,
		\341GAT(20)_pad ,
		_w523_
	);
	LUT4 #(
		.INIT('h0a08)
	) name490 (
		\256GAT(15)_pad ,
		_w479_,
		_w480_,
		_w481_,
		_w524_
	);
	LUT4 #(
		.INIT('h3c87)
	) name491 (
		\256GAT(15)_pad ,
		\324GAT(19)_pad ,
		_w523_,
		_w524_,
		_w525_
	);
	LUT4 #(
		.INIT('h7100)
	) name492 (
		_w477_,
		_w478_,
		_w482_,
		_w525_,
		_w526_
	);
	LUT4 #(
		.INIT('h008e)
	) name493 (
		_w477_,
		_w478_,
		_w482_,
		_w525_,
		_w527_
	);
	LUT4 #(
		.INIT('h32cd)
	) name494 (
		_w477_,
		_w483_,
		_w484_,
		_w525_,
		_w528_
	);
	LUT2 #(
		.INIT('h9)
	) name495 (
		_w521_,
		_w528_,
		_w529_
	);
	LUT3 #(
		.INIT('h96)
	) name496 (
		_w519_,
		_w520_,
		_w529_,
		_w530_
	);
	LUT3 #(
		.INIT('h96)
	) name497 (
		_w517_,
		_w518_,
		_w530_,
		_w531_
	);
	LUT3 #(
		.INIT('h96)
	) name498 (
		_w515_,
		_w516_,
		_w531_,
		_w532_
	);
	LUT3 #(
		.INIT('h96)
	) name499 (
		_w513_,
		_w514_,
		_w532_,
		_w533_
	);
	LUT3 #(
		.INIT('h96)
	) name500 (
		_w511_,
		_w512_,
		_w533_,
		_w534_
	);
	LUT3 #(
		.INIT('h96)
	) name501 (
		_w509_,
		_w510_,
		_w534_,
		_w535_
	);
	LUT3 #(
		.INIT('h96)
	) name502 (
		_w507_,
		_w508_,
		_w535_,
		_w536_
	);
	LUT3 #(
		.INIT('h96)
	) name503 (
		_w505_,
		_w506_,
		_w536_,
		_w537_
	);
	LUT3 #(
		.INIT('h96)
	) name504 (
		_w503_,
		_w504_,
		_w537_,
		_w538_
	);
	LUT3 #(
		.INIT('h96)
	) name505 (
		_w501_,
		_w502_,
		_w538_,
		_w539_
	);
	LUT2 #(
		.INIT('h4)
	) name506 (
		_w500_,
		_w539_,
		_w540_
	);
	LUT2 #(
		.INIT('h2)
	) name507 (
		_w500_,
		_w539_,
		_w541_
	);
	LUT2 #(
		.INIT('h9)
	) name508 (
		_w500_,
		_w539_,
		_w542_
	);
	LUT2 #(
		.INIT('h6)
	) name509 (
		_w499_,
		_w542_,
		_w543_
	);
	LUT3 #(
		.INIT('h8e)
	) name510 (
		_w501_,
		_w502_,
		_w538_,
		_w544_
	);
	LUT2 #(
		.INIT('h8)
	) name511 (
		\528GAT(31)_pad ,
		\69GAT(4)_pad ,
		_w545_
	);
	LUT3 #(
		.INIT('h8e)
	) name512 (
		_w503_,
		_w504_,
		_w537_,
		_w546_
	);
	LUT2 #(
		.INIT('h8)
	) name513 (
		\511GAT(30)_pad ,
		\86GAT(5)_pad ,
		_w547_
	);
	LUT3 #(
		.INIT('h8e)
	) name514 (
		_w505_,
		_w506_,
		_w536_,
		_w548_
	);
	LUT2 #(
		.INIT('h8)
	) name515 (
		\103GAT(6)_pad ,
		\494GAT(29)_pad ,
		_w549_
	);
	LUT3 #(
		.INIT('h8e)
	) name516 (
		_w507_,
		_w508_,
		_w535_,
		_w550_
	);
	LUT2 #(
		.INIT('h8)
	) name517 (
		\120GAT(7)_pad ,
		\477GAT(28)_pad ,
		_w551_
	);
	LUT3 #(
		.INIT('h8e)
	) name518 (
		_w509_,
		_w510_,
		_w534_,
		_w552_
	);
	LUT2 #(
		.INIT('h8)
	) name519 (
		\137GAT(8)_pad ,
		\460GAT(27)_pad ,
		_w553_
	);
	LUT3 #(
		.INIT('h8e)
	) name520 (
		_w511_,
		_w512_,
		_w533_,
		_w554_
	);
	LUT2 #(
		.INIT('h8)
	) name521 (
		\154GAT(9)_pad ,
		\443GAT(26)_pad ,
		_w555_
	);
	LUT3 #(
		.INIT('h8e)
	) name522 (
		_w513_,
		_w514_,
		_w532_,
		_w556_
	);
	LUT2 #(
		.INIT('h8)
	) name523 (
		\171GAT(10)_pad ,
		\426GAT(25)_pad ,
		_w557_
	);
	LUT3 #(
		.INIT('h8e)
	) name524 (
		_w515_,
		_w516_,
		_w531_,
		_w558_
	);
	LUT2 #(
		.INIT('h8)
	) name525 (
		\188GAT(11)_pad ,
		\409GAT(24)_pad ,
		_w559_
	);
	LUT3 #(
		.INIT('h8e)
	) name526 (
		_w517_,
		_w518_,
		_w530_,
		_w560_
	);
	LUT2 #(
		.INIT('h8)
	) name527 (
		\205GAT(12)_pad ,
		\392GAT(23)_pad ,
		_w561_
	);
	LUT3 #(
		.INIT('h8e)
	) name528 (
		_w519_,
		_w520_,
		_w529_,
		_w562_
	);
	LUT2 #(
		.INIT('h8)
	) name529 (
		\222GAT(13)_pad ,
		\375GAT(22)_pad ,
		_w563_
	);
	LUT3 #(
		.INIT('h32)
	) name530 (
		_w521_,
		_w526_,
		_w527_,
		_w564_
	);
	LUT2 #(
		.INIT('h8)
	) name531 (
		\239GAT(14)_pad ,
		\358GAT(21)_pad ,
		_w565_
	);
	LUT4 #(
		.INIT('hfc80)
	) name532 (
		\256GAT(15)_pad ,
		\324GAT(19)_pad ,
		_w523_,
		_w524_,
		_w566_
	);
	LUT2 #(
		.INIT('h8)
	) name533 (
		\256GAT(15)_pad ,
		\341GAT(20)_pad ,
		_w567_
	);
	LUT3 #(
		.INIT('h69)
	) name534 (
		_w565_,
		_w566_,
		_w567_,
		_w568_
	);
	LUT4 #(
		.INIT('h7100)
	) name535 (
		_w521_,
		_w522_,
		_w525_,
		_w568_,
		_w569_
	);
	LUT4 #(
		.INIT('h008e)
	) name536 (
		_w521_,
		_w522_,
		_w525_,
		_w568_,
		_w570_
	);
	LUT4 #(
		.INIT('h32cd)
	) name537 (
		_w521_,
		_w526_,
		_w527_,
		_w568_,
		_w571_
	);
	LUT2 #(
		.INIT('h9)
	) name538 (
		_w563_,
		_w571_,
		_w572_
	);
	LUT3 #(
		.INIT('h96)
	) name539 (
		_w561_,
		_w562_,
		_w572_,
		_w573_
	);
	LUT3 #(
		.INIT('h96)
	) name540 (
		_w559_,
		_w560_,
		_w573_,
		_w574_
	);
	LUT3 #(
		.INIT('h96)
	) name541 (
		_w557_,
		_w558_,
		_w574_,
		_w575_
	);
	LUT3 #(
		.INIT('h96)
	) name542 (
		_w555_,
		_w556_,
		_w575_,
		_w576_
	);
	LUT3 #(
		.INIT('h96)
	) name543 (
		_w553_,
		_w554_,
		_w576_,
		_w577_
	);
	LUT3 #(
		.INIT('h96)
	) name544 (
		_w551_,
		_w552_,
		_w577_,
		_w578_
	);
	LUT3 #(
		.INIT('h96)
	) name545 (
		_w549_,
		_w550_,
		_w578_,
		_w579_
	);
	LUT3 #(
		.INIT('h96)
	) name546 (
		_w547_,
		_w548_,
		_w579_,
		_w580_
	);
	LUT3 #(
		.INIT('h96)
	) name547 (
		_w545_,
		_w546_,
		_w580_,
		_w581_
	);
	LUT2 #(
		.INIT('h4)
	) name548 (
		_w544_,
		_w581_,
		_w582_
	);
	LUT2 #(
		.INIT('h9)
	) name549 (
		_w544_,
		_w581_,
		_w583_
	);
	LUT4 #(
		.INIT('h7100)
	) name550 (
		_w499_,
		_w500_,
		_w539_,
		_w583_,
		_w584_
	);
	LUT4 #(
		.INIT('hcd32)
	) name551 (
		_w499_,
		_w540_,
		_w541_,
		_w583_,
		_w585_
	);
	LUT3 #(
		.INIT('h8e)
	) name552 (
		_w545_,
		_w546_,
		_w580_,
		_w586_
	);
	LUT2 #(
		.INIT('h8)
	) name553 (
		\528GAT(31)_pad ,
		\86GAT(5)_pad ,
		_w587_
	);
	LUT3 #(
		.INIT('h8e)
	) name554 (
		_w547_,
		_w548_,
		_w579_,
		_w588_
	);
	LUT2 #(
		.INIT('h8)
	) name555 (
		\103GAT(6)_pad ,
		\511GAT(30)_pad ,
		_w589_
	);
	LUT3 #(
		.INIT('h8e)
	) name556 (
		_w549_,
		_w550_,
		_w578_,
		_w590_
	);
	LUT2 #(
		.INIT('h8)
	) name557 (
		\120GAT(7)_pad ,
		\494GAT(29)_pad ,
		_w591_
	);
	LUT3 #(
		.INIT('h8e)
	) name558 (
		_w551_,
		_w552_,
		_w577_,
		_w592_
	);
	LUT2 #(
		.INIT('h8)
	) name559 (
		\137GAT(8)_pad ,
		\477GAT(28)_pad ,
		_w593_
	);
	LUT3 #(
		.INIT('h8e)
	) name560 (
		_w553_,
		_w554_,
		_w576_,
		_w594_
	);
	LUT2 #(
		.INIT('h8)
	) name561 (
		\154GAT(9)_pad ,
		\460GAT(27)_pad ,
		_w595_
	);
	LUT3 #(
		.INIT('h8e)
	) name562 (
		_w555_,
		_w556_,
		_w575_,
		_w596_
	);
	LUT2 #(
		.INIT('h8)
	) name563 (
		\171GAT(10)_pad ,
		\443GAT(26)_pad ,
		_w597_
	);
	LUT3 #(
		.INIT('h8e)
	) name564 (
		_w557_,
		_w558_,
		_w574_,
		_w598_
	);
	LUT2 #(
		.INIT('h8)
	) name565 (
		\188GAT(11)_pad ,
		\426GAT(25)_pad ,
		_w599_
	);
	LUT3 #(
		.INIT('h8e)
	) name566 (
		_w559_,
		_w560_,
		_w573_,
		_w600_
	);
	LUT2 #(
		.INIT('h8)
	) name567 (
		\205GAT(12)_pad ,
		\409GAT(24)_pad ,
		_w601_
	);
	LUT3 #(
		.INIT('h8e)
	) name568 (
		_w561_,
		_w562_,
		_w572_,
		_w602_
	);
	LUT2 #(
		.INIT('h8)
	) name569 (
		\222GAT(13)_pad ,
		\392GAT(23)_pad ,
		_w603_
	);
	LUT3 #(
		.INIT('h32)
	) name570 (
		_w563_,
		_w569_,
		_w570_,
		_w604_
	);
	LUT2 #(
		.INIT('h8)
	) name571 (
		\239GAT(14)_pad ,
		\375GAT(22)_pad ,
		_w605_
	);
	LUT3 #(
		.INIT('he8)
	) name572 (
		_w565_,
		_w566_,
		_w567_,
		_w606_
	);
	LUT2 #(
		.INIT('h8)
	) name573 (
		\256GAT(15)_pad ,
		\358GAT(21)_pad ,
		_w607_
	);
	LUT4 #(
		.INIT('h0017)
	) name574 (
		_w565_,
		_w566_,
		_w567_,
		_w607_,
		_w608_
	);
	LUT4 #(
		.INIT('he800)
	) name575 (
		_w565_,
		_w566_,
		_w567_,
		_w607_,
		_w609_
	);
	LUT4 #(
		.INIT('h17e8)
	) name576 (
		_w565_,
		_w566_,
		_w567_,
		_w607_,
		_w610_
	);
	LUT2 #(
		.INIT('h9)
	) name577 (
		_w605_,
		_w610_,
		_w611_
	);
	LUT4 #(
		.INIT('h7100)
	) name578 (
		_w563_,
		_w564_,
		_w568_,
		_w611_,
		_w612_
	);
	LUT4 #(
		.INIT('h008e)
	) name579 (
		_w563_,
		_w564_,
		_w568_,
		_w611_,
		_w613_
	);
	LUT4 #(
		.INIT('h32cd)
	) name580 (
		_w563_,
		_w569_,
		_w570_,
		_w611_,
		_w614_
	);
	LUT2 #(
		.INIT('h9)
	) name581 (
		_w603_,
		_w614_,
		_w615_
	);
	LUT3 #(
		.INIT('h96)
	) name582 (
		_w601_,
		_w602_,
		_w615_,
		_w616_
	);
	LUT3 #(
		.INIT('h96)
	) name583 (
		_w599_,
		_w600_,
		_w616_,
		_w617_
	);
	LUT3 #(
		.INIT('h96)
	) name584 (
		_w597_,
		_w598_,
		_w617_,
		_w618_
	);
	LUT3 #(
		.INIT('h96)
	) name585 (
		_w595_,
		_w596_,
		_w618_,
		_w619_
	);
	LUT3 #(
		.INIT('h96)
	) name586 (
		_w593_,
		_w594_,
		_w619_,
		_w620_
	);
	LUT3 #(
		.INIT('h96)
	) name587 (
		_w591_,
		_w592_,
		_w620_,
		_w621_
	);
	LUT3 #(
		.INIT('h96)
	) name588 (
		_w589_,
		_w590_,
		_w621_,
		_w622_
	);
	LUT3 #(
		.INIT('h96)
	) name589 (
		_w587_,
		_w588_,
		_w622_,
		_w623_
	);
	LUT2 #(
		.INIT('h4)
	) name590 (
		_w586_,
		_w623_,
		_w624_
	);
	LUT2 #(
		.INIT('h2)
	) name591 (
		_w586_,
		_w623_,
		_w625_
	);
	LUT2 #(
		.INIT('h9)
	) name592 (
		_w586_,
		_w623_,
		_w626_
	);
	LUT3 #(
		.INIT('he1)
	) name593 (
		_w582_,
		_w584_,
		_w626_,
		_w627_
	);
	LUT4 #(
		.INIT('h0f01)
	) name594 (
		_w582_,
		_w584_,
		_w624_,
		_w625_,
		_w628_
	);
	LUT3 #(
		.INIT('h8e)
	) name595 (
		_w587_,
		_w588_,
		_w622_,
		_w629_
	);
	LUT2 #(
		.INIT('h8)
	) name596 (
		\103GAT(6)_pad ,
		\528GAT(31)_pad ,
		_w630_
	);
	LUT3 #(
		.INIT('h8e)
	) name597 (
		_w589_,
		_w590_,
		_w621_,
		_w631_
	);
	LUT2 #(
		.INIT('h8)
	) name598 (
		\120GAT(7)_pad ,
		\511GAT(30)_pad ,
		_w632_
	);
	LUT3 #(
		.INIT('h8e)
	) name599 (
		_w591_,
		_w592_,
		_w620_,
		_w633_
	);
	LUT2 #(
		.INIT('h8)
	) name600 (
		\137GAT(8)_pad ,
		\494GAT(29)_pad ,
		_w634_
	);
	LUT3 #(
		.INIT('h8e)
	) name601 (
		_w593_,
		_w594_,
		_w619_,
		_w635_
	);
	LUT2 #(
		.INIT('h8)
	) name602 (
		\154GAT(9)_pad ,
		\477GAT(28)_pad ,
		_w636_
	);
	LUT3 #(
		.INIT('h8e)
	) name603 (
		_w595_,
		_w596_,
		_w618_,
		_w637_
	);
	LUT2 #(
		.INIT('h8)
	) name604 (
		\171GAT(10)_pad ,
		\460GAT(27)_pad ,
		_w638_
	);
	LUT3 #(
		.INIT('h8e)
	) name605 (
		_w597_,
		_w598_,
		_w617_,
		_w639_
	);
	LUT2 #(
		.INIT('h8)
	) name606 (
		\188GAT(11)_pad ,
		\443GAT(26)_pad ,
		_w640_
	);
	LUT3 #(
		.INIT('h8e)
	) name607 (
		_w599_,
		_w600_,
		_w616_,
		_w641_
	);
	LUT2 #(
		.INIT('h8)
	) name608 (
		\205GAT(12)_pad ,
		\426GAT(25)_pad ,
		_w642_
	);
	LUT3 #(
		.INIT('h8e)
	) name609 (
		_w601_,
		_w602_,
		_w615_,
		_w643_
	);
	LUT2 #(
		.INIT('h8)
	) name610 (
		\222GAT(13)_pad ,
		\409GAT(24)_pad ,
		_w644_
	);
	LUT3 #(
		.INIT('h32)
	) name611 (
		_w603_,
		_w612_,
		_w613_,
		_w645_
	);
	LUT2 #(
		.INIT('h8)
	) name612 (
		\239GAT(14)_pad ,
		\392GAT(23)_pad ,
		_w646_
	);
	LUT3 #(
		.INIT('h32)
	) name613 (
		_w605_,
		_w608_,
		_w609_,
		_w647_
	);
	LUT2 #(
		.INIT('h8)
	) name614 (
		\256GAT(15)_pad ,
		\375GAT(22)_pad ,
		_w648_
	);
	LUT4 #(
		.INIT('h0017)
	) name615 (
		_w605_,
		_w606_,
		_w607_,
		_w648_,
		_w649_
	);
	LUT4 #(
		.INIT('he800)
	) name616 (
		_w605_,
		_w606_,
		_w607_,
		_w648_,
		_w650_
	);
	LUT4 #(
		.INIT('hcd32)
	) name617 (
		_w605_,
		_w608_,
		_w609_,
		_w648_,
		_w651_
	);
	LUT2 #(
		.INIT('h9)
	) name618 (
		_w646_,
		_w651_,
		_w652_
	);
	LUT4 #(
		.INIT('h7100)
	) name619 (
		_w603_,
		_w604_,
		_w611_,
		_w652_,
		_w653_
	);
	LUT4 #(
		.INIT('h008e)
	) name620 (
		_w603_,
		_w604_,
		_w611_,
		_w652_,
		_w654_
	);
	LUT4 #(
		.INIT('h32cd)
	) name621 (
		_w603_,
		_w612_,
		_w613_,
		_w652_,
		_w655_
	);
	LUT2 #(
		.INIT('h9)
	) name622 (
		_w644_,
		_w655_,
		_w656_
	);
	LUT3 #(
		.INIT('h96)
	) name623 (
		_w642_,
		_w643_,
		_w656_,
		_w657_
	);
	LUT3 #(
		.INIT('h96)
	) name624 (
		_w640_,
		_w641_,
		_w657_,
		_w658_
	);
	LUT3 #(
		.INIT('h96)
	) name625 (
		_w638_,
		_w639_,
		_w658_,
		_w659_
	);
	LUT3 #(
		.INIT('h96)
	) name626 (
		_w636_,
		_w637_,
		_w659_,
		_w660_
	);
	LUT3 #(
		.INIT('h96)
	) name627 (
		_w634_,
		_w635_,
		_w660_,
		_w661_
	);
	LUT3 #(
		.INIT('h96)
	) name628 (
		_w632_,
		_w633_,
		_w661_,
		_w662_
	);
	LUT3 #(
		.INIT('h96)
	) name629 (
		_w630_,
		_w631_,
		_w662_,
		_w663_
	);
	LUT2 #(
		.INIT('h4)
	) name630 (
		_w629_,
		_w663_,
		_w664_
	);
	LUT2 #(
		.INIT('h2)
	) name631 (
		_w629_,
		_w663_,
		_w665_
	);
	LUT2 #(
		.INIT('h9)
	) name632 (
		_w629_,
		_w663_,
		_w666_
	);
	LUT2 #(
		.INIT('h6)
	) name633 (
		_w628_,
		_w666_,
		_w667_
	);
	LUT3 #(
		.INIT('h8e)
	) name634 (
		_w630_,
		_w631_,
		_w662_,
		_w668_
	);
	LUT2 #(
		.INIT('h8)
	) name635 (
		\120GAT(7)_pad ,
		\528GAT(31)_pad ,
		_w669_
	);
	LUT3 #(
		.INIT('h8e)
	) name636 (
		_w632_,
		_w633_,
		_w661_,
		_w670_
	);
	LUT2 #(
		.INIT('h8)
	) name637 (
		\137GAT(8)_pad ,
		\511GAT(30)_pad ,
		_w671_
	);
	LUT3 #(
		.INIT('h8e)
	) name638 (
		_w634_,
		_w635_,
		_w660_,
		_w672_
	);
	LUT2 #(
		.INIT('h8)
	) name639 (
		\154GAT(9)_pad ,
		\494GAT(29)_pad ,
		_w673_
	);
	LUT3 #(
		.INIT('h8e)
	) name640 (
		_w636_,
		_w637_,
		_w659_,
		_w674_
	);
	LUT2 #(
		.INIT('h8)
	) name641 (
		\171GAT(10)_pad ,
		\477GAT(28)_pad ,
		_w675_
	);
	LUT3 #(
		.INIT('h8e)
	) name642 (
		_w638_,
		_w639_,
		_w658_,
		_w676_
	);
	LUT2 #(
		.INIT('h8)
	) name643 (
		\188GAT(11)_pad ,
		\460GAT(27)_pad ,
		_w677_
	);
	LUT3 #(
		.INIT('h8e)
	) name644 (
		_w640_,
		_w641_,
		_w657_,
		_w678_
	);
	LUT2 #(
		.INIT('h8)
	) name645 (
		\205GAT(12)_pad ,
		\443GAT(26)_pad ,
		_w679_
	);
	LUT3 #(
		.INIT('h8e)
	) name646 (
		_w642_,
		_w643_,
		_w656_,
		_w680_
	);
	LUT2 #(
		.INIT('h8)
	) name647 (
		\222GAT(13)_pad ,
		\426GAT(25)_pad ,
		_w681_
	);
	LUT3 #(
		.INIT('h32)
	) name648 (
		_w644_,
		_w653_,
		_w654_,
		_w682_
	);
	LUT2 #(
		.INIT('h8)
	) name649 (
		\239GAT(14)_pad ,
		\409GAT(24)_pad ,
		_w683_
	);
	LUT3 #(
		.INIT('h32)
	) name650 (
		_w646_,
		_w649_,
		_w650_,
		_w684_
	);
	LUT2 #(
		.INIT('h8)
	) name651 (
		\256GAT(15)_pad ,
		\392GAT(23)_pad ,
		_w685_
	);
	LUT4 #(
		.INIT('h0017)
	) name652 (
		_w646_,
		_w647_,
		_w648_,
		_w685_,
		_w686_
	);
	LUT4 #(
		.INIT('he800)
	) name653 (
		_w646_,
		_w647_,
		_w648_,
		_w685_,
		_w687_
	);
	LUT4 #(
		.INIT('hcd32)
	) name654 (
		_w646_,
		_w649_,
		_w650_,
		_w685_,
		_w688_
	);
	LUT2 #(
		.INIT('h9)
	) name655 (
		_w683_,
		_w688_,
		_w689_
	);
	LUT4 #(
		.INIT('h7100)
	) name656 (
		_w644_,
		_w645_,
		_w652_,
		_w689_,
		_w690_
	);
	LUT4 #(
		.INIT('h008e)
	) name657 (
		_w644_,
		_w645_,
		_w652_,
		_w689_,
		_w691_
	);
	LUT4 #(
		.INIT('h32cd)
	) name658 (
		_w644_,
		_w653_,
		_w654_,
		_w689_,
		_w692_
	);
	LUT2 #(
		.INIT('h9)
	) name659 (
		_w681_,
		_w692_,
		_w693_
	);
	LUT3 #(
		.INIT('h96)
	) name660 (
		_w679_,
		_w680_,
		_w693_,
		_w694_
	);
	LUT3 #(
		.INIT('h96)
	) name661 (
		_w677_,
		_w678_,
		_w694_,
		_w695_
	);
	LUT3 #(
		.INIT('h96)
	) name662 (
		_w675_,
		_w676_,
		_w695_,
		_w696_
	);
	LUT3 #(
		.INIT('h96)
	) name663 (
		_w673_,
		_w674_,
		_w696_,
		_w697_
	);
	LUT3 #(
		.INIT('h96)
	) name664 (
		_w671_,
		_w672_,
		_w697_,
		_w698_
	);
	LUT3 #(
		.INIT('h96)
	) name665 (
		_w669_,
		_w670_,
		_w698_,
		_w699_
	);
	LUT2 #(
		.INIT('h4)
	) name666 (
		_w668_,
		_w699_,
		_w700_
	);
	LUT2 #(
		.INIT('h9)
	) name667 (
		_w668_,
		_w699_,
		_w701_
	);
	LUT4 #(
		.INIT('h7100)
	) name668 (
		_w628_,
		_w629_,
		_w663_,
		_w701_,
		_w702_
	);
	LUT4 #(
		.INIT('hcd32)
	) name669 (
		_w628_,
		_w664_,
		_w665_,
		_w701_,
		_w703_
	);
	LUT3 #(
		.INIT('h8e)
	) name670 (
		_w669_,
		_w670_,
		_w698_,
		_w704_
	);
	LUT2 #(
		.INIT('h8)
	) name671 (
		\137GAT(8)_pad ,
		\528GAT(31)_pad ,
		_w705_
	);
	LUT3 #(
		.INIT('h8e)
	) name672 (
		_w671_,
		_w672_,
		_w697_,
		_w706_
	);
	LUT2 #(
		.INIT('h8)
	) name673 (
		\154GAT(9)_pad ,
		\511GAT(30)_pad ,
		_w707_
	);
	LUT3 #(
		.INIT('h8e)
	) name674 (
		_w673_,
		_w674_,
		_w696_,
		_w708_
	);
	LUT2 #(
		.INIT('h8)
	) name675 (
		\171GAT(10)_pad ,
		\494GAT(29)_pad ,
		_w709_
	);
	LUT3 #(
		.INIT('h8e)
	) name676 (
		_w675_,
		_w676_,
		_w695_,
		_w710_
	);
	LUT2 #(
		.INIT('h8)
	) name677 (
		\188GAT(11)_pad ,
		\477GAT(28)_pad ,
		_w711_
	);
	LUT3 #(
		.INIT('h8e)
	) name678 (
		_w677_,
		_w678_,
		_w694_,
		_w712_
	);
	LUT2 #(
		.INIT('h8)
	) name679 (
		\205GAT(12)_pad ,
		\460GAT(27)_pad ,
		_w713_
	);
	LUT3 #(
		.INIT('h8e)
	) name680 (
		_w679_,
		_w680_,
		_w693_,
		_w714_
	);
	LUT2 #(
		.INIT('h8)
	) name681 (
		\222GAT(13)_pad ,
		\443GAT(26)_pad ,
		_w715_
	);
	LUT3 #(
		.INIT('h32)
	) name682 (
		_w681_,
		_w690_,
		_w691_,
		_w716_
	);
	LUT2 #(
		.INIT('h8)
	) name683 (
		\239GAT(14)_pad ,
		\426GAT(25)_pad ,
		_w717_
	);
	LUT3 #(
		.INIT('h32)
	) name684 (
		_w683_,
		_w686_,
		_w687_,
		_w718_
	);
	LUT2 #(
		.INIT('h8)
	) name685 (
		\256GAT(15)_pad ,
		\409GAT(24)_pad ,
		_w719_
	);
	LUT4 #(
		.INIT('h0017)
	) name686 (
		_w683_,
		_w684_,
		_w685_,
		_w719_,
		_w720_
	);
	LUT4 #(
		.INIT('he800)
	) name687 (
		_w683_,
		_w684_,
		_w685_,
		_w719_,
		_w721_
	);
	LUT4 #(
		.INIT('hcd32)
	) name688 (
		_w683_,
		_w686_,
		_w687_,
		_w719_,
		_w722_
	);
	LUT2 #(
		.INIT('h9)
	) name689 (
		_w717_,
		_w722_,
		_w723_
	);
	LUT4 #(
		.INIT('h7100)
	) name690 (
		_w681_,
		_w682_,
		_w689_,
		_w723_,
		_w724_
	);
	LUT4 #(
		.INIT('h008e)
	) name691 (
		_w681_,
		_w682_,
		_w689_,
		_w723_,
		_w725_
	);
	LUT4 #(
		.INIT('h32cd)
	) name692 (
		_w681_,
		_w690_,
		_w691_,
		_w723_,
		_w726_
	);
	LUT2 #(
		.INIT('h9)
	) name693 (
		_w715_,
		_w726_,
		_w727_
	);
	LUT3 #(
		.INIT('h96)
	) name694 (
		_w713_,
		_w714_,
		_w727_,
		_w728_
	);
	LUT3 #(
		.INIT('h96)
	) name695 (
		_w711_,
		_w712_,
		_w728_,
		_w729_
	);
	LUT3 #(
		.INIT('h96)
	) name696 (
		_w709_,
		_w710_,
		_w729_,
		_w730_
	);
	LUT3 #(
		.INIT('h96)
	) name697 (
		_w707_,
		_w708_,
		_w730_,
		_w731_
	);
	LUT3 #(
		.INIT('h96)
	) name698 (
		_w705_,
		_w706_,
		_w731_,
		_w732_
	);
	LUT2 #(
		.INIT('h4)
	) name699 (
		_w704_,
		_w732_,
		_w733_
	);
	LUT2 #(
		.INIT('h2)
	) name700 (
		_w704_,
		_w732_,
		_w734_
	);
	LUT2 #(
		.INIT('h9)
	) name701 (
		_w704_,
		_w732_,
		_w735_
	);
	LUT3 #(
		.INIT('he1)
	) name702 (
		_w700_,
		_w702_,
		_w735_,
		_w736_
	);
	LUT4 #(
		.INIT('h0f01)
	) name703 (
		_w700_,
		_w702_,
		_w733_,
		_w734_,
		_w737_
	);
	LUT3 #(
		.INIT('h8e)
	) name704 (
		_w705_,
		_w706_,
		_w731_,
		_w738_
	);
	LUT2 #(
		.INIT('h8)
	) name705 (
		\154GAT(9)_pad ,
		\528GAT(31)_pad ,
		_w739_
	);
	LUT3 #(
		.INIT('h8e)
	) name706 (
		_w707_,
		_w708_,
		_w730_,
		_w740_
	);
	LUT2 #(
		.INIT('h8)
	) name707 (
		\171GAT(10)_pad ,
		\511GAT(30)_pad ,
		_w741_
	);
	LUT3 #(
		.INIT('h8e)
	) name708 (
		_w709_,
		_w710_,
		_w729_,
		_w742_
	);
	LUT2 #(
		.INIT('h8)
	) name709 (
		\188GAT(11)_pad ,
		\494GAT(29)_pad ,
		_w743_
	);
	LUT3 #(
		.INIT('h8e)
	) name710 (
		_w711_,
		_w712_,
		_w728_,
		_w744_
	);
	LUT2 #(
		.INIT('h8)
	) name711 (
		\205GAT(12)_pad ,
		\477GAT(28)_pad ,
		_w745_
	);
	LUT3 #(
		.INIT('h8e)
	) name712 (
		_w713_,
		_w714_,
		_w727_,
		_w746_
	);
	LUT2 #(
		.INIT('h8)
	) name713 (
		\222GAT(13)_pad ,
		\460GAT(27)_pad ,
		_w747_
	);
	LUT3 #(
		.INIT('h32)
	) name714 (
		_w715_,
		_w724_,
		_w725_,
		_w748_
	);
	LUT2 #(
		.INIT('h8)
	) name715 (
		\239GAT(14)_pad ,
		\443GAT(26)_pad ,
		_w749_
	);
	LUT3 #(
		.INIT('h32)
	) name716 (
		_w717_,
		_w720_,
		_w721_,
		_w750_
	);
	LUT2 #(
		.INIT('h8)
	) name717 (
		\256GAT(15)_pad ,
		\426GAT(25)_pad ,
		_w751_
	);
	LUT4 #(
		.INIT('h0017)
	) name718 (
		_w717_,
		_w718_,
		_w719_,
		_w751_,
		_w752_
	);
	LUT4 #(
		.INIT('he800)
	) name719 (
		_w717_,
		_w718_,
		_w719_,
		_w751_,
		_w753_
	);
	LUT4 #(
		.INIT('hcd32)
	) name720 (
		_w717_,
		_w720_,
		_w721_,
		_w751_,
		_w754_
	);
	LUT2 #(
		.INIT('h9)
	) name721 (
		_w749_,
		_w754_,
		_w755_
	);
	LUT4 #(
		.INIT('h7100)
	) name722 (
		_w715_,
		_w716_,
		_w723_,
		_w755_,
		_w756_
	);
	LUT4 #(
		.INIT('h008e)
	) name723 (
		_w715_,
		_w716_,
		_w723_,
		_w755_,
		_w757_
	);
	LUT4 #(
		.INIT('h32cd)
	) name724 (
		_w715_,
		_w724_,
		_w725_,
		_w755_,
		_w758_
	);
	LUT2 #(
		.INIT('h9)
	) name725 (
		_w747_,
		_w758_,
		_w759_
	);
	LUT3 #(
		.INIT('h96)
	) name726 (
		_w745_,
		_w746_,
		_w759_,
		_w760_
	);
	LUT3 #(
		.INIT('h96)
	) name727 (
		_w743_,
		_w744_,
		_w760_,
		_w761_
	);
	LUT3 #(
		.INIT('h96)
	) name728 (
		_w741_,
		_w742_,
		_w761_,
		_w762_
	);
	LUT3 #(
		.INIT('h96)
	) name729 (
		_w739_,
		_w740_,
		_w762_,
		_w763_
	);
	LUT2 #(
		.INIT('h4)
	) name730 (
		_w738_,
		_w763_,
		_w764_
	);
	LUT2 #(
		.INIT('h2)
	) name731 (
		_w738_,
		_w763_,
		_w765_
	);
	LUT2 #(
		.INIT('h9)
	) name732 (
		_w738_,
		_w763_,
		_w766_
	);
	LUT2 #(
		.INIT('h6)
	) name733 (
		_w737_,
		_w766_,
		_w767_
	);
	LUT3 #(
		.INIT('h8e)
	) name734 (
		_w739_,
		_w740_,
		_w762_,
		_w768_
	);
	LUT2 #(
		.INIT('h8)
	) name735 (
		\171GAT(10)_pad ,
		\528GAT(31)_pad ,
		_w769_
	);
	LUT3 #(
		.INIT('h8e)
	) name736 (
		_w741_,
		_w742_,
		_w761_,
		_w770_
	);
	LUT2 #(
		.INIT('h8)
	) name737 (
		\188GAT(11)_pad ,
		\511GAT(30)_pad ,
		_w771_
	);
	LUT3 #(
		.INIT('h8e)
	) name738 (
		_w743_,
		_w744_,
		_w760_,
		_w772_
	);
	LUT2 #(
		.INIT('h8)
	) name739 (
		\205GAT(12)_pad ,
		\494GAT(29)_pad ,
		_w773_
	);
	LUT3 #(
		.INIT('h8e)
	) name740 (
		_w745_,
		_w746_,
		_w759_,
		_w774_
	);
	LUT2 #(
		.INIT('h8)
	) name741 (
		\222GAT(13)_pad ,
		\477GAT(28)_pad ,
		_w775_
	);
	LUT3 #(
		.INIT('h32)
	) name742 (
		_w747_,
		_w756_,
		_w757_,
		_w776_
	);
	LUT2 #(
		.INIT('h8)
	) name743 (
		\239GAT(14)_pad ,
		\460GAT(27)_pad ,
		_w777_
	);
	LUT3 #(
		.INIT('h32)
	) name744 (
		_w749_,
		_w752_,
		_w753_,
		_w778_
	);
	LUT2 #(
		.INIT('h8)
	) name745 (
		\256GAT(15)_pad ,
		\443GAT(26)_pad ,
		_w779_
	);
	LUT4 #(
		.INIT('h0017)
	) name746 (
		_w749_,
		_w750_,
		_w751_,
		_w779_,
		_w780_
	);
	LUT4 #(
		.INIT('he800)
	) name747 (
		_w749_,
		_w750_,
		_w751_,
		_w779_,
		_w781_
	);
	LUT4 #(
		.INIT('hcd32)
	) name748 (
		_w749_,
		_w752_,
		_w753_,
		_w779_,
		_w782_
	);
	LUT2 #(
		.INIT('h9)
	) name749 (
		_w777_,
		_w782_,
		_w783_
	);
	LUT4 #(
		.INIT('h7100)
	) name750 (
		_w747_,
		_w748_,
		_w755_,
		_w783_,
		_w784_
	);
	LUT4 #(
		.INIT('h008e)
	) name751 (
		_w747_,
		_w748_,
		_w755_,
		_w783_,
		_w785_
	);
	LUT4 #(
		.INIT('h32cd)
	) name752 (
		_w747_,
		_w756_,
		_w757_,
		_w783_,
		_w786_
	);
	LUT2 #(
		.INIT('h9)
	) name753 (
		_w775_,
		_w786_,
		_w787_
	);
	LUT3 #(
		.INIT('h96)
	) name754 (
		_w773_,
		_w774_,
		_w787_,
		_w788_
	);
	LUT3 #(
		.INIT('h96)
	) name755 (
		_w771_,
		_w772_,
		_w788_,
		_w789_
	);
	LUT3 #(
		.INIT('h96)
	) name756 (
		_w769_,
		_w770_,
		_w789_,
		_w790_
	);
	LUT2 #(
		.INIT('h4)
	) name757 (
		_w768_,
		_w790_,
		_w791_
	);
	LUT2 #(
		.INIT('h9)
	) name758 (
		_w768_,
		_w790_,
		_w792_
	);
	LUT4 #(
		.INIT('h7100)
	) name759 (
		_w737_,
		_w738_,
		_w763_,
		_w792_,
		_w793_
	);
	LUT4 #(
		.INIT('hcd32)
	) name760 (
		_w737_,
		_w764_,
		_w765_,
		_w792_,
		_w794_
	);
	LUT3 #(
		.INIT('h8e)
	) name761 (
		_w769_,
		_w770_,
		_w789_,
		_w795_
	);
	LUT2 #(
		.INIT('h8)
	) name762 (
		\188GAT(11)_pad ,
		\528GAT(31)_pad ,
		_w796_
	);
	LUT3 #(
		.INIT('h8e)
	) name763 (
		_w771_,
		_w772_,
		_w788_,
		_w797_
	);
	LUT2 #(
		.INIT('h8)
	) name764 (
		\205GAT(12)_pad ,
		\511GAT(30)_pad ,
		_w798_
	);
	LUT3 #(
		.INIT('h8e)
	) name765 (
		_w773_,
		_w774_,
		_w787_,
		_w799_
	);
	LUT2 #(
		.INIT('h8)
	) name766 (
		\222GAT(13)_pad ,
		\494GAT(29)_pad ,
		_w800_
	);
	LUT3 #(
		.INIT('h32)
	) name767 (
		_w775_,
		_w784_,
		_w785_,
		_w801_
	);
	LUT2 #(
		.INIT('h8)
	) name768 (
		\239GAT(14)_pad ,
		\477GAT(28)_pad ,
		_w802_
	);
	LUT3 #(
		.INIT('h32)
	) name769 (
		_w777_,
		_w780_,
		_w781_,
		_w803_
	);
	LUT2 #(
		.INIT('h8)
	) name770 (
		\256GAT(15)_pad ,
		\460GAT(27)_pad ,
		_w804_
	);
	LUT4 #(
		.INIT('h0017)
	) name771 (
		_w777_,
		_w778_,
		_w779_,
		_w804_,
		_w805_
	);
	LUT4 #(
		.INIT('he800)
	) name772 (
		_w777_,
		_w778_,
		_w779_,
		_w804_,
		_w806_
	);
	LUT4 #(
		.INIT('hcd32)
	) name773 (
		_w777_,
		_w780_,
		_w781_,
		_w804_,
		_w807_
	);
	LUT2 #(
		.INIT('h9)
	) name774 (
		_w802_,
		_w807_,
		_w808_
	);
	LUT4 #(
		.INIT('h7100)
	) name775 (
		_w775_,
		_w776_,
		_w783_,
		_w808_,
		_w809_
	);
	LUT4 #(
		.INIT('h008e)
	) name776 (
		_w775_,
		_w776_,
		_w783_,
		_w808_,
		_w810_
	);
	LUT4 #(
		.INIT('h32cd)
	) name777 (
		_w775_,
		_w784_,
		_w785_,
		_w808_,
		_w811_
	);
	LUT2 #(
		.INIT('h9)
	) name778 (
		_w800_,
		_w811_,
		_w812_
	);
	LUT3 #(
		.INIT('h96)
	) name779 (
		_w798_,
		_w799_,
		_w812_,
		_w813_
	);
	LUT3 #(
		.INIT('h96)
	) name780 (
		_w796_,
		_w797_,
		_w813_,
		_w814_
	);
	LUT2 #(
		.INIT('h4)
	) name781 (
		_w795_,
		_w814_,
		_w815_
	);
	LUT2 #(
		.INIT('h2)
	) name782 (
		_w795_,
		_w814_,
		_w816_
	);
	LUT2 #(
		.INIT('h9)
	) name783 (
		_w795_,
		_w814_,
		_w817_
	);
	LUT3 #(
		.INIT('he1)
	) name784 (
		_w791_,
		_w793_,
		_w817_,
		_w818_
	);
	LUT4 #(
		.INIT('h0f01)
	) name785 (
		_w791_,
		_w793_,
		_w815_,
		_w816_,
		_w819_
	);
	LUT3 #(
		.INIT('h8e)
	) name786 (
		_w796_,
		_w797_,
		_w813_,
		_w820_
	);
	LUT2 #(
		.INIT('h8)
	) name787 (
		\205GAT(12)_pad ,
		\528GAT(31)_pad ,
		_w821_
	);
	LUT3 #(
		.INIT('h8e)
	) name788 (
		_w798_,
		_w799_,
		_w812_,
		_w822_
	);
	LUT2 #(
		.INIT('h8)
	) name789 (
		\222GAT(13)_pad ,
		\511GAT(30)_pad ,
		_w823_
	);
	LUT3 #(
		.INIT('h32)
	) name790 (
		_w800_,
		_w809_,
		_w810_,
		_w824_
	);
	LUT2 #(
		.INIT('h8)
	) name791 (
		\239GAT(14)_pad ,
		\494GAT(29)_pad ,
		_w825_
	);
	LUT3 #(
		.INIT('h32)
	) name792 (
		_w802_,
		_w805_,
		_w806_,
		_w826_
	);
	LUT2 #(
		.INIT('h8)
	) name793 (
		\256GAT(15)_pad ,
		\477GAT(28)_pad ,
		_w827_
	);
	LUT4 #(
		.INIT('h0017)
	) name794 (
		_w802_,
		_w803_,
		_w804_,
		_w827_,
		_w828_
	);
	LUT4 #(
		.INIT('he800)
	) name795 (
		_w802_,
		_w803_,
		_w804_,
		_w827_,
		_w829_
	);
	LUT4 #(
		.INIT('hcd32)
	) name796 (
		_w802_,
		_w805_,
		_w806_,
		_w827_,
		_w830_
	);
	LUT2 #(
		.INIT('h9)
	) name797 (
		_w825_,
		_w830_,
		_w831_
	);
	LUT4 #(
		.INIT('h7100)
	) name798 (
		_w800_,
		_w801_,
		_w808_,
		_w831_,
		_w832_
	);
	LUT4 #(
		.INIT('h008e)
	) name799 (
		_w800_,
		_w801_,
		_w808_,
		_w831_,
		_w833_
	);
	LUT4 #(
		.INIT('h32cd)
	) name800 (
		_w800_,
		_w809_,
		_w810_,
		_w831_,
		_w834_
	);
	LUT2 #(
		.INIT('h9)
	) name801 (
		_w823_,
		_w834_,
		_w835_
	);
	LUT3 #(
		.INIT('h96)
	) name802 (
		_w821_,
		_w822_,
		_w835_,
		_w836_
	);
	LUT2 #(
		.INIT('h4)
	) name803 (
		_w820_,
		_w836_,
		_w837_
	);
	LUT2 #(
		.INIT('h2)
	) name804 (
		_w820_,
		_w836_,
		_w838_
	);
	LUT2 #(
		.INIT('h9)
	) name805 (
		_w820_,
		_w836_,
		_w839_
	);
	LUT2 #(
		.INIT('h6)
	) name806 (
		_w819_,
		_w839_,
		_w840_
	);
	LUT3 #(
		.INIT('h8e)
	) name807 (
		_w821_,
		_w822_,
		_w835_,
		_w841_
	);
	LUT2 #(
		.INIT('h8)
	) name808 (
		\222GAT(13)_pad ,
		\528GAT(31)_pad ,
		_w842_
	);
	LUT3 #(
		.INIT('h32)
	) name809 (
		_w823_,
		_w832_,
		_w833_,
		_w843_
	);
	LUT2 #(
		.INIT('h8)
	) name810 (
		\239GAT(14)_pad ,
		\511GAT(30)_pad ,
		_w844_
	);
	LUT3 #(
		.INIT('h32)
	) name811 (
		_w825_,
		_w828_,
		_w829_,
		_w845_
	);
	LUT2 #(
		.INIT('h8)
	) name812 (
		\256GAT(15)_pad ,
		\494GAT(29)_pad ,
		_w846_
	);
	LUT4 #(
		.INIT('h0017)
	) name813 (
		_w825_,
		_w826_,
		_w827_,
		_w846_,
		_w847_
	);
	LUT4 #(
		.INIT('he800)
	) name814 (
		_w825_,
		_w826_,
		_w827_,
		_w846_,
		_w848_
	);
	LUT4 #(
		.INIT('hcd32)
	) name815 (
		_w825_,
		_w828_,
		_w829_,
		_w846_,
		_w849_
	);
	LUT2 #(
		.INIT('h9)
	) name816 (
		_w844_,
		_w849_,
		_w850_
	);
	LUT4 #(
		.INIT('h7100)
	) name817 (
		_w823_,
		_w824_,
		_w831_,
		_w850_,
		_w851_
	);
	LUT4 #(
		.INIT('h008e)
	) name818 (
		_w823_,
		_w824_,
		_w831_,
		_w850_,
		_w852_
	);
	LUT4 #(
		.INIT('h32cd)
	) name819 (
		_w823_,
		_w832_,
		_w833_,
		_w850_,
		_w853_
	);
	LUT2 #(
		.INIT('h9)
	) name820 (
		_w842_,
		_w853_,
		_w854_
	);
	LUT2 #(
		.INIT('h4)
	) name821 (
		_w841_,
		_w854_,
		_w855_
	);
	LUT2 #(
		.INIT('h9)
	) name822 (
		_w841_,
		_w854_,
		_w856_
	);
	LUT4 #(
		.INIT('h7100)
	) name823 (
		_w819_,
		_w820_,
		_w836_,
		_w856_,
		_w857_
	);
	LUT4 #(
		.INIT('hcd32)
	) name824 (
		_w819_,
		_w837_,
		_w838_,
		_w856_,
		_w858_
	);
	LUT2 #(
		.INIT('h8)
	) name825 (
		\239GAT(14)_pad ,
		\528GAT(31)_pad ,
		_w859_
	);
	LUT3 #(
		.INIT('h32)
	) name826 (
		_w844_,
		_w847_,
		_w848_,
		_w860_
	);
	LUT2 #(
		.INIT('h8)
	) name827 (
		\256GAT(15)_pad ,
		\511GAT(30)_pad ,
		_w861_
	);
	LUT4 #(
		.INIT('h0017)
	) name828 (
		_w844_,
		_w845_,
		_w846_,
		_w861_,
		_w862_
	);
	LUT4 #(
		.INIT('he800)
	) name829 (
		_w844_,
		_w845_,
		_w846_,
		_w861_,
		_w863_
	);
	LUT4 #(
		.INIT('hcd32)
	) name830 (
		_w844_,
		_w847_,
		_w848_,
		_w861_,
		_w864_
	);
	LUT2 #(
		.INIT('h9)
	) name831 (
		_w859_,
		_w864_,
		_w865_
	);
	LUT4 #(
		.INIT('h7100)
	) name832 (
		_w842_,
		_w843_,
		_w850_,
		_w865_,
		_w866_
	);
	LUT4 #(
		.INIT('h32cd)
	) name833 (
		_w842_,
		_w851_,
		_w852_,
		_w865_,
		_w867_
	);
	LUT3 #(
		.INIT('he1)
	) name834 (
		_w855_,
		_w857_,
		_w867_,
		_w868_
	);
	LUT2 #(
		.INIT('h8)
	) name835 (
		\256GAT(15)_pad ,
		\528GAT(31)_pad ,
		_w869_
	);
	LUT4 #(
		.INIT('h0017)
	) name836 (
		_w859_,
		_w860_,
		_w861_,
		_w869_,
		_w870_
	);
	LUT4 #(
		.INIT('h010f)
	) name837 (
		_w855_,
		_w857_,
		_w866_,
		_w867_,
		_w871_
	);
	LUT4 #(
		.INIT('he800)
	) name838 (
		_w859_,
		_w860_,
		_w861_,
		_w869_,
		_w872_
	);
	LUT4 #(
		.INIT('hcd32)
	) name839 (
		_w859_,
		_w862_,
		_w863_,
		_w869_,
		_w873_
	);
	LUT3 #(
		.INIT('h54)
	) name840 (
		_w870_,
		_w871_,
		_w872_,
		_w874_
	);
	LUT2 #(
		.INIT('h6)
	) name841 (
		_w871_,
		_w873_,
		_w875_
	);
	assign \1581GAT(423)_pad  = _w35_ ;
	assign \1901GAT(561)_pad  = _w41_ ;
	assign \2223GAT(700)_pad  = _w51_ ;
	assign \2548GAT(840)_pad  = _w64_ ;
	assign \2877GAT(983)_pad  = _w80_ ;
	assign \3211GAT(1128)_pad  = _w98_ ;
	assign \3552GAT(1275)_pad  = _w121_ ;
	assign \3895GAT(1423)_pad  = _w146_ ;
	assign \4241GAT(1572)_pad  = _w174_ ;
	assign \4591GAT(1722)_pad  = _w205_ ;
	assign \4946GAT(1876)_pad  = _w239_ ;
	assign \5308GAT(2031)_pad  = _w276_ ;
	assign \545GAT(287)_pad  = _w277_ ;
	assign \5672GAT(2187)_pad  = _w317_ ;
	assign \5971GAT(2309)_pad  = _w360_ ;
	assign \6123GAT(2368)_pad  = _w406_ ;
	assign \6150GAT(2378)_pad  = _w453_ ;
	assign \6160GAT(2383)_pad  = _w498_ ;
	assign \6170GAT(2388)_pad  = _w543_ ;
	assign \6180GAT(2393)_pad  = _w585_ ;
	assign \6190GAT(2398)_pad  = _w627_ ;
	assign \6200GAT(2403)_pad  = _w667_ ;
	assign \6210GAT(2408)_pad  = _w703_ ;
	assign \6220GAT(2413)_pad  = _w736_ ;
	assign \6230GAT(2418)_pad  = _w767_ ;
	assign \6240GAT(2423)_pad  = _w794_ ;
	assign \6250GAT(2428)_pad  = _w818_ ;
	assign \6260GAT(2433)_pad  = _w840_ ;
	assign \6270GAT(2438)_pad  = _w858_ ;
	assign \6280GAT(2443)_pad  = _w868_ ;
	assign \6287GAT(2444)_pad  = _w874_ ;
	assign \6288GAT(2447)_pad  = _w875_ ;
endmodule;