module top( \1_pad  , \2_pad  , \3_pad  , \4_pad  , \5_pad  , \6_pad  , \7_pad  , \24_pad  , \25_pad  , \26_pad  , \27_pad  );
  input \1_pad  ;
  input \2_pad  ;
  input \3_pad  ;
  input \4_pad  ;
  input \5_pad  ;
  input \6_pad  ;
  input \7_pad  ;
  output \24_pad  ;
  output \25_pad  ;
  output \26_pad  ;
  output \27_pad  ;
  wire n8 , n9 , n10 , n11 , n12 , n13 , n14 , n15 , n16 , n17 , n18 , n19 , n20 , n21 , n22 , n23 , n24 , n25 , n26 , n27 , n28 , n29 , n30 , n31 ;
  assign n8 = \2_pad  & \5_pad  ;
  assign n9 = ~\2_pad  & ~\5_pad  ;
  assign n10 = \3_pad  & \6_pad  ;
  assign n11 = ~\3_pad  & ~\6_pad  ;
  assign n12 = \1_pad  & \4_pad  ;
  assign n13 = ~\1_pad  & ~\4_pad  ;
  assign n14 = \7_pad  & ~n13 ;
  assign n15 = ~n12 & ~n14 ;
  assign n16 = ~n11 & ~n15 ;
  assign n17 = ~n10 & ~n16 ;
  assign n18 = ~n9 & ~n17 ;
  assign n19 = ~n8 & ~n18 ;
  assign n20 = ~n8 & ~n9 ;
  assign n21 = ~n17 & n20 ;
  assign n22 = n17 & ~n20 ;
  assign n23 = ~n21 & ~n22 ;
  assign n24 = ~n10 & ~n11 ;
  assign n25 = ~n15 & n24 ;
  assign n26 = n15 & ~n24 ;
  assign n27 = ~n25 & ~n26 ;
  assign n28 = ~n12 & ~n13 ;
  assign n29 = ~\7_pad  & n28 ;
  assign n30 = \7_pad  & ~n28 ;
  assign n31 = ~n29 & ~n30 ;
  assign \24_pad  = ~n19 ;
  assign \25_pad  = n23 ;
  assign \26_pad  = n27 ;
  assign \27_pad  = ~n31 ;
endmodule
