module top (\FP_R_reg[10]/P0001 , \FP_R_reg[11]/P0001 , \FP_R_reg[12]/P0001 , \FP_R_reg[13]/P0001 , \FP_R_reg[14]/P0001 , \FP_R_reg[15]/P0001 , \FP_R_reg[16]/P0001 , \FP_R_reg[17]/P0001 , \FP_R_reg[18]/P0001 , \FP_R_reg[19]/P0001 , \FP_R_reg[1]/P0001 , \FP_R_reg[20]/P0001 , \FP_R_reg[21]/P0001 , \FP_R_reg[22]/P0001 , \FP_R_reg[23]/P0001 , \FP_R_reg[24]/P0001 , \FP_R_reg[25]/P0001 , \FP_R_reg[26]/P0001 , \FP_R_reg[27]/P0001 , \FP_R_reg[28]/P0001 , \FP_R_reg[29]/P0001 , \FP_R_reg[2]/P0001 , \FP_R_reg[30]/P0001 , \FP_R_reg[31]/P0001 , \FP_R_reg[32]/P0001 , \FP_R_reg[33]/NET0131 , \FP_R_reg[34]/NET0131 , \FP_R_reg[35]/NET0131 , \FP_R_reg[36]/NET0131 , \FP_R_reg[37]/NET0131 , \FP_R_reg[38]/NET0131 , \FP_R_reg[39]/NET0131 , \FP_R_reg[3]/P0001 , \FP_R_reg[40]/NET0131 , \FP_R_reg[41]/NET0131 , \FP_R_reg[42]/NET0131 , \FP_R_reg[43]/NET0131 , \FP_R_reg[44]/NET0131 , \FP_R_reg[45]/NET0131 , \FP_R_reg[46]/NET0131 , \FP_R_reg[47]/NET0131 , \FP_R_reg[48]/NET0131 , \FP_R_reg[49]/NET0131 , \FP_R_reg[4]/P0001 , \FP_R_reg[50]/NET0131 , \FP_R_reg[51]/NET0131 , \FP_R_reg[52]/NET0131 , \FP_R_reg[53]/NET0131 , \FP_R_reg[54]/NET0131 , \FP_R_reg[55]/NET0131 , \FP_R_reg[56]/NET0131 , \FP_R_reg[57]/NET0131 , \FP_R_reg[58]/NET0131 , \FP_R_reg[59]/NET0131 , \FP_R_reg[5]/P0001 , \FP_R_reg[60]/NET0131 , \FP_R_reg[61]/NET0131 , \FP_R_reg[62]/NET0131 , \FP_R_reg[63]/NET0131 , \FP_R_reg[64]/NET0131 , \FP_R_reg[6]/P0001 , \FP_R_reg[7]/P0001 , \FP_R_reg[8]/P0001 , \FP_R_reg[9]/P0001 , decrypt_pad, \desIn[0]_pad , \desIn[10]_pad , \desIn[11]_pad , \desIn[12]_pad , \desIn[13]_pad , \desIn[14]_pad , \desIn[15]_pad , \desIn[16]_pad , \desIn[17]_pad , \desIn[18]_pad , \desIn[19]_pad , \desIn[1]_pad , \desIn[20]_pad , \desIn[21]_pad , \desIn[22]_pad , \desIn[23]_pad , \desIn[24]_pad , \desIn[25]_pad , \desIn[26]_pad , \desIn[27]_pad , \desIn[28]_pad , \desIn[29]_pad , \desIn[2]_pad , \desIn[30]_pad , \desIn[31]_pad , \desIn[32]_pad , \desIn[33]_pad , \desIn[34]_pad , \desIn[35]_pad , \desIn[36]_pad , \desIn[37]_pad , \desIn[38]_pad , \desIn[39]_pad , \desIn[3]_pad , \desIn[40]_pad , \desIn[41]_pad , \desIn[42]_pad , \desIn[43]_pad , \desIn[44]_pad , \desIn[45]_pad , \desIn[46]_pad , \desIn[47]_pad , \desIn[48]_pad , \desIn[49]_pad , \desIn[4]_pad , \desIn[50]_pad , \desIn[51]_pad , \desIn[52]_pad , \desIn[53]_pad , \desIn[54]_pad , \desIn[55]_pad , \desIn[56]_pad , \desIn[57]_pad , \desIn[58]_pad , \desIn[59]_pad , \desIn[5]_pad , \desIn[60]_pad , \desIn[61]_pad , \desIn[62]_pad , \desIn[63]_pad , \desIn[6]_pad , \desIn[7]_pad , \desIn[8]_pad , \desIn[9]_pad , \key1[0]_pad , \key1[10]_pad , \key1[11]_pad , \key1[12]_pad , \key1[13]_pad , \key1[14]_pad , \key1[15]_pad , \key1[16]_pad , \key1[17]_pad , \key1[18]_pad , \key1[19]_pad , \key1[1]_pad , \key1[20]_pad , \key1[21]_pad , \key1[22]_pad , \key1[23]_pad , \key1[24]_pad , \key1[25]_pad , \key1[26]_pad , \key1[27]_pad , \key1[28]_pad , \key1[29]_pad , \key1[2]_pad , \key1[30]_pad , \key1[31]_pad , \key1[32]_pad , \key1[33]_pad , \key1[34]_pad , \key1[35]_pad , \key1[36]_pad , \key1[37]_pad , \key1[38]_pad , \key1[39]_pad , \key1[3]_pad , \key1[40]_pad , \key1[41]_pad , \key1[42]_pad , \key1[43]_pad , \key1[44]_pad , \key1[45]_pad , \key1[46]_pad , \key1[47]_pad , \key1[48]_pad , \key1[49]_pad , \key1[4]_pad , \key1[50]_pad , \key1[51]_pad , \key1[52]_pad , \key1[53]_pad , \key1[54]_pad , \key1[55]_pad , \key1[5]_pad , \key1[6]_pad , \key1[7]_pad , \key1[8]_pad , \key1[9]_pad , \key2[0]_pad , \key2[10]_pad , \key2[11]_pad , \key2[12]_pad , \key2[13]_pad , \key2[14]_pad , \key2[15]_pad , \key2[16]_pad , \key2[17]_pad , \key2[18]_pad , \key2[19]_pad , \key2[1]_pad , \key2[20]_pad , \key2[21]_pad , \key2[22]_pad , \key2[23]_pad , \key2[24]_pad , \key2[25]_pad , \key2[26]_pad , \key2[27]_pad , \key2[28]_pad , \key2[29]_pad , \key2[2]_pad , \key2[30]_pad , \key2[31]_pad , \key2[32]_pad , \key2[33]_pad , \key2[34]_pad , \key2[35]_pad , \key2[36]_pad , \key2[37]_pad , \key2[38]_pad , \key2[39]_pad , \key2[3]_pad , \key2[40]_pad , \key2[41]_pad , \key2[42]_pad , \key2[43]_pad , \key2[44]_pad , \key2[45]_pad , \key2[46]_pad , \key2[47]_pad , \key2[48]_pad , \key2[49]_pad , \key2[4]_pad , \key2[50]_pad , \key2[51]_pad , \key2[52]_pad , \key2[53]_pad , \key2[54]_pad , \key2[55]_pad , \key2[5]_pad , \key2[6]_pad , \key2[7]_pad , \key2[8]_pad , \key2[9]_pad , \key3[0]_pad , \key3[10]_pad , \key3[11]_pad , \key3[12]_pad , \key3[13]_pad , \key3[14]_pad , \key3[15]_pad , \key3[16]_pad , \key3[17]_pad , \key3[18]_pad , \key3[19]_pad , \key3[1]_pad , \key3[20]_pad , \key3[21]_pad , \key3[22]_pad , \key3[23]_pad , \key3[24]_pad , \key3[25]_pad , \key3[26]_pad , \key3[27]_pad , \key3[28]_pad , \key3[29]_pad , \key3[2]_pad , \key3[30]_pad , \key3[31]_pad , \key3[32]_pad , \key3[33]_pad , \key3[34]_pad , \key3[35]_pad , \key3[36]_pad , \key3[37]_pad , \key3[38]_pad , \key3[39]_pad , \key3[3]_pad , \key3[40]_pad , \key3[41]_pad , \key3[42]_pad , \key3[43]_pad , \key3[44]_pad , \key3[45]_pad , \key3[46]_pad , \key3[47]_pad , \key3[48]_pad , \key3[49]_pad , \key3[4]_pad , \key3[50]_pad , \key3[51]_pad , \key3[52]_pad , \key3[53]_pad , \key3[54]_pad , \key3[55]_pad , \key3[5]_pad , \key3[6]_pad , \key3[7]_pad , \key3[8]_pad , \key3[9]_pad , \roundSel[0]_pad , \roundSel[1]_pad , \roundSel[2]_pad , \roundSel[3]_pad , \roundSel[4]_pad , \roundSel[5]_pad , \_al_n0 , \_al_n1 , \desOut[0]_pad , \desOut[11]_pad , \desOut[12]_pad , \desOut[13]_pad , \desOut[14]_pad , \desOut[15]_pad , \desOut[18]_pad , \desOut[1]_pad , \desOut[22]_pad , \desOut[23]_pad , \desOut[24]_pad , \desOut[25]_pad , \desOut[26]_pad , \desOut[28]_pad , \desOut[2]_pad , \desOut[30]_pad , \desOut[32]_pad , \desOut[34]_pad , \desOut[35]_pad , \desOut[37]_pad , \desOut[38]_pad , \desOut[39]_pad , \desOut[3]_pad , \desOut[40]_pad , \desOut[42]_pad , \desOut[44]_pad , \desOut[45]_pad , \desOut[46]_pad , \desOut[48]_pad , \desOut[4]_pad , \desOut[50]_pad , \desOut[52]_pad , \desOut[54]_pad , \desOut[56]_pad , \desOut[57]_pad , \desOut[59]_pad , \desOut[5]_pad , \desOut[60]_pad , \desOut[61]_pad , \desOut[63]_pad , \desOut[6]_pad , \desOut[8]_pad , \desOut[9]_pad , \g13525_dup/_0_ , \g13583_dup/_0_ , \g17813/_3_ , \g17816/_3_ , \g17819/_3_ , \g17822/_3_ , \g17836/_3_ , \g17871/_3_ , \g17878/_1_ , \g17881/_3_ , \g17966/_2_ , \g17969/_3_ , \g17996/_2_ , \g19574_dup/_3_ , \g19619_dup/_3_ , \g19756_dup/_3_ , \g20263/_3_ , \g20541/_2_ , \g20691/_1_ , \g20740_dup/_3_ , \g67/_2_ );
	input \FP_R_reg[10]/P0001  ;
	input \FP_R_reg[11]/P0001  ;
	input \FP_R_reg[12]/P0001  ;
	input \FP_R_reg[13]/P0001  ;
	input \FP_R_reg[14]/P0001  ;
	input \FP_R_reg[15]/P0001  ;
	input \FP_R_reg[16]/P0001  ;
	input \FP_R_reg[17]/P0001  ;
	input \FP_R_reg[18]/P0001  ;
	input \FP_R_reg[19]/P0001  ;
	input \FP_R_reg[1]/P0001  ;
	input \FP_R_reg[20]/P0001  ;
	input \FP_R_reg[21]/P0001  ;
	input \FP_R_reg[22]/P0001  ;
	input \FP_R_reg[23]/P0001  ;
	input \FP_R_reg[24]/P0001  ;
	input \FP_R_reg[25]/P0001  ;
	input \FP_R_reg[26]/P0001  ;
	input \FP_R_reg[27]/P0001  ;
	input \FP_R_reg[28]/P0001  ;
	input \FP_R_reg[29]/P0001  ;
	input \FP_R_reg[2]/P0001  ;
	input \FP_R_reg[30]/P0001  ;
	input \FP_R_reg[31]/P0001  ;
	input \FP_R_reg[32]/P0001  ;
	input \FP_R_reg[33]/NET0131  ;
	input \FP_R_reg[34]/NET0131  ;
	input \FP_R_reg[35]/NET0131  ;
	input \FP_R_reg[36]/NET0131  ;
	input \FP_R_reg[37]/NET0131  ;
	input \FP_R_reg[38]/NET0131  ;
	input \FP_R_reg[39]/NET0131  ;
	input \FP_R_reg[3]/P0001  ;
	input \FP_R_reg[40]/NET0131  ;
	input \FP_R_reg[41]/NET0131  ;
	input \FP_R_reg[42]/NET0131  ;
	input \FP_R_reg[43]/NET0131  ;
	input \FP_R_reg[44]/NET0131  ;
	input \FP_R_reg[45]/NET0131  ;
	input \FP_R_reg[46]/NET0131  ;
	input \FP_R_reg[47]/NET0131  ;
	input \FP_R_reg[48]/NET0131  ;
	input \FP_R_reg[49]/NET0131  ;
	input \FP_R_reg[4]/P0001  ;
	input \FP_R_reg[50]/NET0131  ;
	input \FP_R_reg[51]/NET0131  ;
	input \FP_R_reg[52]/NET0131  ;
	input \FP_R_reg[53]/NET0131  ;
	input \FP_R_reg[54]/NET0131  ;
	input \FP_R_reg[55]/NET0131  ;
	input \FP_R_reg[56]/NET0131  ;
	input \FP_R_reg[57]/NET0131  ;
	input \FP_R_reg[58]/NET0131  ;
	input \FP_R_reg[59]/NET0131  ;
	input \FP_R_reg[5]/P0001  ;
	input \FP_R_reg[60]/NET0131  ;
	input \FP_R_reg[61]/NET0131  ;
	input \FP_R_reg[62]/NET0131  ;
	input \FP_R_reg[63]/NET0131  ;
	input \FP_R_reg[64]/NET0131  ;
	input \FP_R_reg[6]/P0001  ;
	input \FP_R_reg[7]/P0001  ;
	input \FP_R_reg[8]/P0001  ;
	input \FP_R_reg[9]/P0001  ;
	input decrypt_pad ;
	input \desIn[0]_pad  ;
	input \desIn[10]_pad  ;
	input \desIn[11]_pad  ;
	input \desIn[12]_pad  ;
	input \desIn[13]_pad  ;
	input \desIn[14]_pad  ;
	input \desIn[15]_pad  ;
	input \desIn[16]_pad  ;
	input \desIn[17]_pad  ;
	input \desIn[18]_pad  ;
	input \desIn[19]_pad  ;
	input \desIn[1]_pad  ;
	input \desIn[20]_pad  ;
	input \desIn[21]_pad  ;
	input \desIn[22]_pad  ;
	input \desIn[23]_pad  ;
	input \desIn[24]_pad  ;
	input \desIn[25]_pad  ;
	input \desIn[26]_pad  ;
	input \desIn[27]_pad  ;
	input \desIn[28]_pad  ;
	input \desIn[29]_pad  ;
	input \desIn[2]_pad  ;
	input \desIn[30]_pad  ;
	input \desIn[31]_pad  ;
	input \desIn[32]_pad  ;
	input \desIn[33]_pad  ;
	input \desIn[34]_pad  ;
	input \desIn[35]_pad  ;
	input \desIn[36]_pad  ;
	input \desIn[37]_pad  ;
	input \desIn[38]_pad  ;
	input \desIn[39]_pad  ;
	input \desIn[3]_pad  ;
	input \desIn[40]_pad  ;
	input \desIn[41]_pad  ;
	input \desIn[42]_pad  ;
	input \desIn[43]_pad  ;
	input \desIn[44]_pad  ;
	input \desIn[45]_pad  ;
	input \desIn[46]_pad  ;
	input \desIn[47]_pad  ;
	input \desIn[48]_pad  ;
	input \desIn[49]_pad  ;
	input \desIn[4]_pad  ;
	input \desIn[50]_pad  ;
	input \desIn[51]_pad  ;
	input \desIn[52]_pad  ;
	input \desIn[53]_pad  ;
	input \desIn[54]_pad  ;
	input \desIn[55]_pad  ;
	input \desIn[56]_pad  ;
	input \desIn[57]_pad  ;
	input \desIn[58]_pad  ;
	input \desIn[59]_pad  ;
	input \desIn[5]_pad  ;
	input \desIn[60]_pad  ;
	input \desIn[61]_pad  ;
	input \desIn[62]_pad  ;
	input \desIn[63]_pad  ;
	input \desIn[6]_pad  ;
	input \desIn[7]_pad  ;
	input \desIn[8]_pad  ;
	input \desIn[9]_pad  ;
	input \key1[0]_pad  ;
	input \key1[10]_pad  ;
	input \key1[11]_pad  ;
	input \key1[12]_pad  ;
	input \key1[13]_pad  ;
	input \key1[14]_pad  ;
	input \key1[15]_pad  ;
	input \key1[16]_pad  ;
	input \key1[17]_pad  ;
	input \key1[18]_pad  ;
	input \key1[19]_pad  ;
	input \key1[1]_pad  ;
	input \key1[20]_pad  ;
	input \key1[21]_pad  ;
	input \key1[22]_pad  ;
	input \key1[23]_pad  ;
	input \key1[24]_pad  ;
	input \key1[25]_pad  ;
	input \key1[26]_pad  ;
	input \key1[27]_pad  ;
	input \key1[28]_pad  ;
	input \key1[29]_pad  ;
	input \key1[2]_pad  ;
	input \key1[30]_pad  ;
	input \key1[31]_pad  ;
	input \key1[32]_pad  ;
	input \key1[33]_pad  ;
	input \key1[34]_pad  ;
	input \key1[35]_pad  ;
	input \key1[36]_pad  ;
	input \key1[37]_pad  ;
	input \key1[38]_pad  ;
	input \key1[39]_pad  ;
	input \key1[3]_pad  ;
	input \key1[40]_pad  ;
	input \key1[41]_pad  ;
	input \key1[42]_pad  ;
	input \key1[43]_pad  ;
	input \key1[44]_pad  ;
	input \key1[45]_pad  ;
	input \key1[46]_pad  ;
	input \key1[47]_pad  ;
	input \key1[48]_pad  ;
	input \key1[49]_pad  ;
	input \key1[4]_pad  ;
	input \key1[50]_pad  ;
	input \key1[51]_pad  ;
	input \key1[52]_pad  ;
	input \key1[53]_pad  ;
	input \key1[54]_pad  ;
	input \key1[55]_pad  ;
	input \key1[5]_pad  ;
	input \key1[6]_pad  ;
	input \key1[7]_pad  ;
	input \key1[8]_pad  ;
	input \key1[9]_pad  ;
	input \key2[0]_pad  ;
	input \key2[10]_pad  ;
	input \key2[11]_pad  ;
	input \key2[12]_pad  ;
	input \key2[13]_pad  ;
	input \key2[14]_pad  ;
	input \key2[15]_pad  ;
	input \key2[16]_pad  ;
	input \key2[17]_pad  ;
	input \key2[18]_pad  ;
	input \key2[19]_pad  ;
	input \key2[1]_pad  ;
	input \key2[20]_pad  ;
	input \key2[21]_pad  ;
	input \key2[22]_pad  ;
	input \key2[23]_pad  ;
	input \key2[24]_pad  ;
	input \key2[25]_pad  ;
	input \key2[26]_pad  ;
	input \key2[27]_pad  ;
	input \key2[28]_pad  ;
	input \key2[29]_pad  ;
	input \key2[2]_pad  ;
	input \key2[30]_pad  ;
	input \key2[31]_pad  ;
	input \key2[32]_pad  ;
	input \key2[33]_pad  ;
	input \key2[34]_pad  ;
	input \key2[35]_pad  ;
	input \key2[36]_pad  ;
	input \key2[37]_pad  ;
	input \key2[38]_pad  ;
	input \key2[39]_pad  ;
	input \key2[3]_pad  ;
	input \key2[40]_pad  ;
	input \key2[41]_pad  ;
	input \key2[42]_pad  ;
	input \key2[43]_pad  ;
	input \key2[44]_pad  ;
	input \key2[45]_pad  ;
	input \key2[46]_pad  ;
	input \key2[47]_pad  ;
	input \key2[48]_pad  ;
	input \key2[49]_pad  ;
	input \key2[4]_pad  ;
	input \key2[50]_pad  ;
	input \key2[51]_pad  ;
	input \key2[52]_pad  ;
	input \key2[53]_pad  ;
	input \key2[54]_pad  ;
	input \key2[55]_pad  ;
	input \key2[5]_pad  ;
	input \key2[6]_pad  ;
	input \key2[7]_pad  ;
	input \key2[8]_pad  ;
	input \key2[9]_pad  ;
	input \key3[0]_pad  ;
	input \key3[10]_pad  ;
	input \key3[11]_pad  ;
	input \key3[12]_pad  ;
	input \key3[13]_pad  ;
	input \key3[14]_pad  ;
	input \key3[15]_pad  ;
	input \key3[16]_pad  ;
	input \key3[17]_pad  ;
	input \key3[18]_pad  ;
	input \key3[19]_pad  ;
	input \key3[1]_pad  ;
	input \key3[20]_pad  ;
	input \key3[21]_pad  ;
	input \key3[22]_pad  ;
	input \key3[23]_pad  ;
	input \key3[24]_pad  ;
	input \key3[25]_pad  ;
	input \key3[26]_pad  ;
	input \key3[27]_pad  ;
	input \key3[28]_pad  ;
	input \key3[29]_pad  ;
	input \key3[2]_pad  ;
	input \key3[30]_pad  ;
	input \key3[31]_pad  ;
	input \key3[32]_pad  ;
	input \key3[33]_pad  ;
	input \key3[34]_pad  ;
	input \key3[35]_pad  ;
	input \key3[36]_pad  ;
	input \key3[37]_pad  ;
	input \key3[38]_pad  ;
	input \key3[39]_pad  ;
	input \key3[3]_pad  ;
	input \key3[40]_pad  ;
	input \key3[41]_pad  ;
	input \key3[42]_pad  ;
	input \key3[43]_pad  ;
	input \key3[44]_pad  ;
	input \key3[45]_pad  ;
	input \key3[46]_pad  ;
	input \key3[47]_pad  ;
	input \key3[48]_pad  ;
	input \key3[49]_pad  ;
	input \key3[4]_pad  ;
	input \key3[50]_pad  ;
	input \key3[51]_pad  ;
	input \key3[52]_pad  ;
	input \key3[53]_pad  ;
	input \key3[54]_pad  ;
	input \key3[55]_pad  ;
	input \key3[5]_pad  ;
	input \key3[6]_pad  ;
	input \key3[7]_pad  ;
	input \key3[8]_pad  ;
	input \key3[9]_pad  ;
	input \roundSel[0]_pad  ;
	input \roundSel[1]_pad  ;
	input \roundSel[2]_pad  ;
	input \roundSel[3]_pad  ;
	input \roundSel[4]_pad  ;
	input \roundSel[5]_pad  ;
	output \_al_n0  ;
	output \_al_n1  ;
	output \desOut[0]_pad  ;
	output \desOut[11]_pad  ;
	output \desOut[12]_pad  ;
	output \desOut[13]_pad  ;
	output \desOut[14]_pad  ;
	output \desOut[15]_pad  ;
	output \desOut[18]_pad  ;
	output \desOut[1]_pad  ;
	output \desOut[22]_pad  ;
	output \desOut[23]_pad  ;
	output \desOut[24]_pad  ;
	output \desOut[25]_pad  ;
	output \desOut[26]_pad  ;
	output \desOut[28]_pad  ;
	output \desOut[2]_pad  ;
	output \desOut[30]_pad  ;
	output \desOut[32]_pad  ;
	output \desOut[34]_pad  ;
	output \desOut[35]_pad  ;
	output \desOut[37]_pad  ;
	output \desOut[38]_pad  ;
	output \desOut[39]_pad  ;
	output \desOut[3]_pad  ;
	output \desOut[40]_pad  ;
	output \desOut[42]_pad  ;
	output \desOut[44]_pad  ;
	output \desOut[45]_pad  ;
	output \desOut[46]_pad  ;
	output \desOut[48]_pad  ;
	output \desOut[4]_pad  ;
	output \desOut[50]_pad  ;
	output \desOut[52]_pad  ;
	output \desOut[54]_pad  ;
	output \desOut[56]_pad  ;
	output \desOut[57]_pad  ;
	output \desOut[59]_pad  ;
	output \desOut[5]_pad  ;
	output \desOut[60]_pad  ;
	output \desOut[61]_pad  ;
	output \desOut[63]_pad  ;
	output \desOut[6]_pad  ;
	output \desOut[8]_pad  ;
	output \desOut[9]_pad  ;
	output \g13525_dup/_0_  ;
	output \g13583_dup/_0_  ;
	output \g17813/_3_  ;
	output \g17816/_3_  ;
	output \g17819/_3_  ;
	output \g17822/_3_  ;
	output \g17836/_3_  ;
	output \g17871/_3_  ;
	output \g17878/_1_  ;
	output \g17881/_3_  ;
	output \g17966/_2_  ;
	output \g17969/_3_  ;
	output \g17996/_2_  ;
	output \g19574_dup/_3_  ;
	output \g19619_dup/_3_  ;
	output \g19756_dup/_3_  ;
	output \g20263/_3_  ;
	output \g20541/_2_  ;
	output \g20691/_1_  ;
	output \g20740_dup/_3_  ;
	output \g67/_2_  ;
	wire _w2604_ ;
	wire _w2603_ ;
	wire _w2602_ ;
	wire _w2601_ ;
	wire _w2600_ ;
	wire _w2599_ ;
	wire _w2598_ ;
	wire _w2597_ ;
	wire _w2596_ ;
	wire _w2595_ ;
	wire _w2594_ ;
	wire _w2593_ ;
	wire _w2592_ ;
	wire _w2591_ ;
	wire _w2590_ ;
	wire _w2589_ ;
	wire _w2588_ ;
	wire _w2587_ ;
	wire _w2586_ ;
	wire _w2585_ ;
	wire _w2584_ ;
	wire _w2583_ ;
	wire _w2582_ ;
	wire _w2581_ ;
	wire _w2580_ ;
	wire _w2579_ ;
	wire _w2578_ ;
	wire _w2577_ ;
	wire _w2576_ ;
	wire _w2575_ ;
	wire _w2574_ ;
	wire _w2573_ ;
	wire _w2572_ ;
	wire _w2571_ ;
	wire _w2570_ ;
	wire _w2569_ ;
	wire _w2568_ ;
	wire _w2567_ ;
	wire _w2566_ ;
	wire _w2565_ ;
	wire _w2564_ ;
	wire _w2563_ ;
	wire _w2562_ ;
	wire _w2561_ ;
	wire _w2560_ ;
	wire _w2559_ ;
	wire _w2558_ ;
	wire _w2557_ ;
	wire _w2556_ ;
	wire _w2555_ ;
	wire _w2554_ ;
	wire _w2553_ ;
	wire _w2552_ ;
	wire _w2551_ ;
	wire _w2550_ ;
	wire _w2549_ ;
	wire _w2548_ ;
	wire _w2547_ ;
	wire _w2546_ ;
	wire _w2545_ ;
	wire _w2544_ ;
	wire _w2543_ ;
	wire _w2542_ ;
	wire _w2541_ ;
	wire _w2540_ ;
	wire _w2539_ ;
	wire _w2538_ ;
	wire _w2537_ ;
	wire _w2536_ ;
	wire _w2535_ ;
	wire _w2534_ ;
	wire _w2533_ ;
	wire _w2532_ ;
	wire _w2531_ ;
	wire _w2530_ ;
	wire _w2529_ ;
	wire _w2528_ ;
	wire _w2527_ ;
	wire _w2526_ ;
	wire _w2525_ ;
	wire _w2524_ ;
	wire _w2523_ ;
	wire _w2522_ ;
	wire _w2521_ ;
	wire _w2520_ ;
	wire _w2519_ ;
	wire _w2518_ ;
	wire _w2517_ ;
	wire _w2516_ ;
	wire _w2515_ ;
	wire _w2514_ ;
	wire _w2513_ ;
	wire _w2512_ ;
	wire _w2511_ ;
	wire _w2510_ ;
	wire _w2509_ ;
	wire _w2508_ ;
	wire _w2507_ ;
	wire _w2506_ ;
	wire _w2505_ ;
	wire _w2504_ ;
	wire _w2503_ ;
	wire _w2502_ ;
	wire _w2501_ ;
	wire _w2500_ ;
	wire _w2499_ ;
	wire _w2498_ ;
	wire _w2497_ ;
	wire _w2496_ ;
	wire _w2495_ ;
	wire _w2494_ ;
	wire _w2493_ ;
	wire _w2492_ ;
	wire _w2491_ ;
	wire _w2490_ ;
	wire _w2489_ ;
	wire _w2488_ ;
	wire _w2487_ ;
	wire _w2486_ ;
	wire _w2485_ ;
	wire _w2484_ ;
	wire _w2483_ ;
	wire _w2482_ ;
	wire _w2481_ ;
	wire _w2480_ ;
	wire _w2479_ ;
	wire _w2478_ ;
	wire _w2477_ ;
	wire _w2476_ ;
	wire _w2475_ ;
	wire _w2474_ ;
	wire _w2473_ ;
	wire _w2472_ ;
	wire _w2471_ ;
	wire _w2470_ ;
	wire _w2469_ ;
	wire _w2468_ ;
	wire _w2467_ ;
	wire _w2466_ ;
	wire _w2465_ ;
	wire _w2464_ ;
	wire _w2463_ ;
	wire _w2462_ ;
	wire _w2461_ ;
	wire _w2460_ ;
	wire _w2459_ ;
	wire _w2458_ ;
	wire _w2457_ ;
	wire _w2456_ ;
	wire _w2455_ ;
	wire _w2454_ ;
	wire _w2453_ ;
	wire _w2452_ ;
	wire _w2451_ ;
	wire _w2450_ ;
	wire _w2449_ ;
	wire _w2448_ ;
	wire _w2447_ ;
	wire _w2446_ ;
	wire _w2445_ ;
	wire _w2444_ ;
	wire _w2443_ ;
	wire _w2442_ ;
	wire _w2441_ ;
	wire _w2440_ ;
	wire _w2439_ ;
	wire _w2438_ ;
	wire _w2437_ ;
	wire _w2436_ ;
	wire _w2435_ ;
	wire _w2434_ ;
	wire _w2433_ ;
	wire _w2432_ ;
	wire _w2431_ ;
	wire _w2430_ ;
	wire _w2429_ ;
	wire _w2428_ ;
	wire _w2427_ ;
	wire _w2426_ ;
	wire _w2425_ ;
	wire _w2424_ ;
	wire _w2423_ ;
	wire _w2422_ ;
	wire _w2421_ ;
	wire _w2420_ ;
	wire _w2419_ ;
	wire _w2418_ ;
	wire _w2417_ ;
	wire _w2416_ ;
	wire _w2415_ ;
	wire _w2414_ ;
	wire _w2413_ ;
	wire _w2412_ ;
	wire _w2411_ ;
	wire _w2410_ ;
	wire _w2409_ ;
	wire _w2408_ ;
	wire _w2407_ ;
	wire _w2406_ ;
	wire _w2405_ ;
	wire _w2404_ ;
	wire _w2403_ ;
	wire _w2402_ ;
	wire _w2401_ ;
	wire _w2400_ ;
	wire _w2399_ ;
	wire _w2398_ ;
	wire _w2397_ ;
	wire _w2396_ ;
	wire _w2395_ ;
	wire _w2394_ ;
	wire _w2393_ ;
	wire _w2392_ ;
	wire _w2391_ ;
	wire _w2390_ ;
	wire _w2389_ ;
	wire _w2388_ ;
	wire _w2387_ ;
	wire _w2386_ ;
	wire _w2385_ ;
	wire _w2384_ ;
	wire _w2383_ ;
	wire _w2382_ ;
	wire _w2381_ ;
	wire _w2380_ ;
	wire _w2379_ ;
	wire _w2378_ ;
	wire _w2377_ ;
	wire _w2376_ ;
	wire _w2375_ ;
	wire _w2374_ ;
	wire _w2373_ ;
	wire _w2372_ ;
	wire _w2371_ ;
	wire _w2370_ ;
	wire _w2369_ ;
	wire _w2368_ ;
	wire _w2367_ ;
	wire _w2366_ ;
	wire _w2365_ ;
	wire _w2364_ ;
	wire _w2363_ ;
	wire _w2362_ ;
	wire _w2361_ ;
	wire _w2360_ ;
	wire _w2359_ ;
	wire _w2358_ ;
	wire _w2357_ ;
	wire _w2356_ ;
	wire _w2355_ ;
	wire _w2354_ ;
	wire _w2353_ ;
	wire _w2352_ ;
	wire _w2351_ ;
	wire _w2350_ ;
	wire _w2349_ ;
	wire _w2348_ ;
	wire _w2347_ ;
	wire _w2346_ ;
	wire _w2345_ ;
	wire _w2344_ ;
	wire _w2343_ ;
	wire _w2342_ ;
	wire _w2341_ ;
	wire _w2340_ ;
	wire _w2339_ ;
	wire _w2338_ ;
	wire _w2337_ ;
	wire _w2336_ ;
	wire _w2335_ ;
	wire _w2334_ ;
	wire _w2333_ ;
	wire _w2332_ ;
	wire _w2331_ ;
	wire _w2330_ ;
	wire _w2329_ ;
	wire _w2328_ ;
	wire _w2327_ ;
	wire _w2326_ ;
	wire _w2325_ ;
	wire _w2324_ ;
	wire _w2323_ ;
	wire _w2322_ ;
	wire _w2321_ ;
	wire _w2320_ ;
	wire _w2319_ ;
	wire _w2318_ ;
	wire _w2317_ ;
	wire _w2316_ ;
	wire _w2315_ ;
	wire _w2314_ ;
	wire _w2313_ ;
	wire _w2312_ ;
	wire _w2311_ ;
	wire _w2310_ ;
	wire _w2309_ ;
	wire _w2308_ ;
	wire _w2307_ ;
	wire _w2306_ ;
	wire _w2305_ ;
	wire _w2304_ ;
	wire _w2303_ ;
	wire _w2302_ ;
	wire _w2301_ ;
	wire _w2300_ ;
	wire _w2299_ ;
	wire _w2298_ ;
	wire _w2297_ ;
	wire _w2296_ ;
	wire _w2295_ ;
	wire _w2294_ ;
	wire _w2293_ ;
	wire _w2292_ ;
	wire _w2291_ ;
	wire _w2290_ ;
	wire _w2289_ ;
	wire _w2288_ ;
	wire _w2287_ ;
	wire _w2286_ ;
	wire _w2285_ ;
	wire _w2284_ ;
	wire _w2283_ ;
	wire _w2282_ ;
	wire _w2281_ ;
	wire _w2280_ ;
	wire _w2279_ ;
	wire _w2278_ ;
	wire _w2277_ ;
	wire _w2276_ ;
	wire _w2275_ ;
	wire _w2274_ ;
	wire _w2273_ ;
	wire _w2272_ ;
	wire _w2271_ ;
	wire _w2270_ ;
	wire _w2269_ ;
	wire _w2268_ ;
	wire _w2267_ ;
	wire _w2266_ ;
	wire _w2265_ ;
	wire _w2264_ ;
	wire _w2263_ ;
	wire _w2262_ ;
	wire _w2261_ ;
	wire _w2260_ ;
	wire _w2259_ ;
	wire _w2258_ ;
	wire _w2257_ ;
	wire _w2256_ ;
	wire _w2255_ ;
	wire _w2254_ ;
	wire _w2253_ ;
	wire _w2252_ ;
	wire _w2251_ ;
	wire _w2250_ ;
	wire _w2249_ ;
	wire _w2248_ ;
	wire _w2247_ ;
	wire _w2246_ ;
	wire _w2245_ ;
	wire _w2244_ ;
	wire _w2243_ ;
	wire _w2242_ ;
	wire _w2241_ ;
	wire _w2240_ ;
	wire _w2239_ ;
	wire _w2238_ ;
	wire _w2237_ ;
	wire _w2236_ ;
	wire _w2235_ ;
	wire _w2234_ ;
	wire _w2233_ ;
	wire _w2232_ ;
	wire _w2231_ ;
	wire _w2230_ ;
	wire _w2229_ ;
	wire _w2228_ ;
	wire _w2227_ ;
	wire _w2226_ ;
	wire _w2225_ ;
	wire _w2224_ ;
	wire _w2223_ ;
	wire _w2222_ ;
	wire _w2221_ ;
	wire _w2220_ ;
	wire _w2219_ ;
	wire _w2218_ ;
	wire _w2217_ ;
	wire _w2216_ ;
	wire _w2215_ ;
	wire _w2214_ ;
	wire _w2213_ ;
	wire _w2212_ ;
	wire _w2211_ ;
	wire _w2210_ ;
	wire _w2209_ ;
	wire _w2208_ ;
	wire _w2207_ ;
	wire _w2206_ ;
	wire _w2205_ ;
	wire _w2204_ ;
	wire _w2203_ ;
	wire _w2202_ ;
	wire _w2201_ ;
	wire _w2200_ ;
	wire _w2199_ ;
	wire _w2198_ ;
	wire _w2197_ ;
	wire _w2196_ ;
	wire _w2195_ ;
	wire _w2194_ ;
	wire _w2193_ ;
	wire _w2192_ ;
	wire _w2191_ ;
	wire _w2190_ ;
	wire _w2189_ ;
	wire _w2188_ ;
	wire _w2187_ ;
	wire _w2186_ ;
	wire _w2185_ ;
	wire _w2184_ ;
	wire _w2183_ ;
	wire _w2182_ ;
	wire _w2181_ ;
	wire _w2180_ ;
	wire _w2179_ ;
	wire _w2178_ ;
	wire _w2177_ ;
	wire _w2176_ ;
	wire _w2175_ ;
	wire _w2174_ ;
	wire _w2173_ ;
	wire _w2172_ ;
	wire _w2171_ ;
	wire _w2170_ ;
	wire _w2169_ ;
	wire _w2168_ ;
	wire _w2167_ ;
	wire _w2166_ ;
	wire _w2165_ ;
	wire _w2164_ ;
	wire _w2163_ ;
	wire _w2162_ ;
	wire _w2161_ ;
	wire _w2160_ ;
	wire _w2159_ ;
	wire _w2158_ ;
	wire _w2157_ ;
	wire _w2156_ ;
	wire _w2155_ ;
	wire _w2154_ ;
	wire _w2153_ ;
	wire _w2152_ ;
	wire _w2151_ ;
	wire _w2150_ ;
	wire _w2149_ ;
	wire _w2148_ ;
	wire _w2147_ ;
	wire _w2146_ ;
	wire _w2145_ ;
	wire _w2144_ ;
	wire _w2143_ ;
	wire _w2142_ ;
	wire _w2141_ ;
	wire _w2140_ ;
	wire _w2139_ ;
	wire _w2138_ ;
	wire _w2137_ ;
	wire _w2136_ ;
	wire _w2135_ ;
	wire _w2134_ ;
	wire _w2133_ ;
	wire _w2132_ ;
	wire _w2131_ ;
	wire _w2130_ ;
	wire _w2129_ ;
	wire _w2128_ ;
	wire _w2127_ ;
	wire _w2126_ ;
	wire _w2125_ ;
	wire _w2124_ ;
	wire _w2123_ ;
	wire _w2122_ ;
	wire _w2121_ ;
	wire _w2120_ ;
	wire _w2119_ ;
	wire _w2118_ ;
	wire _w2117_ ;
	wire _w2116_ ;
	wire _w2115_ ;
	wire _w2114_ ;
	wire _w2113_ ;
	wire _w2112_ ;
	wire _w2111_ ;
	wire _w2110_ ;
	wire _w2109_ ;
	wire _w2108_ ;
	wire _w2107_ ;
	wire _w2106_ ;
	wire _w2105_ ;
	wire _w2104_ ;
	wire _w2103_ ;
	wire _w2102_ ;
	wire _w2101_ ;
	wire _w2100_ ;
	wire _w2099_ ;
	wire _w2098_ ;
	wire _w2097_ ;
	wire _w2096_ ;
	wire _w2095_ ;
	wire _w2094_ ;
	wire _w2093_ ;
	wire _w2092_ ;
	wire _w2091_ ;
	wire _w2090_ ;
	wire _w2089_ ;
	wire _w2088_ ;
	wire _w2087_ ;
	wire _w2086_ ;
	wire _w2085_ ;
	wire _w2084_ ;
	wire _w2083_ ;
	wire _w2082_ ;
	wire _w2081_ ;
	wire _w2080_ ;
	wire _w2079_ ;
	wire _w2078_ ;
	wire _w2077_ ;
	wire _w2076_ ;
	wire _w2075_ ;
	wire _w2074_ ;
	wire _w2073_ ;
	wire _w2072_ ;
	wire _w2071_ ;
	wire _w2070_ ;
	wire _w2069_ ;
	wire _w2068_ ;
	wire _w2067_ ;
	wire _w2066_ ;
	wire _w2065_ ;
	wire _w2064_ ;
	wire _w2063_ ;
	wire _w2062_ ;
	wire _w2061_ ;
	wire _w2060_ ;
	wire _w2059_ ;
	wire _w2058_ ;
	wire _w2057_ ;
	wire _w2056_ ;
	wire _w2055_ ;
	wire _w2054_ ;
	wire _w2053_ ;
	wire _w2052_ ;
	wire _w2051_ ;
	wire _w2050_ ;
	wire _w2049_ ;
	wire _w2048_ ;
	wire _w2047_ ;
	wire _w2046_ ;
	wire _w2045_ ;
	wire _w2044_ ;
	wire _w2043_ ;
	wire _w2042_ ;
	wire _w2041_ ;
	wire _w2040_ ;
	wire _w2039_ ;
	wire _w2038_ ;
	wire _w2037_ ;
	wire _w2036_ ;
	wire _w2035_ ;
	wire _w2034_ ;
	wire _w2033_ ;
	wire _w2032_ ;
	wire _w2031_ ;
	wire _w2030_ ;
	wire _w2029_ ;
	wire _w2028_ ;
	wire _w2027_ ;
	wire _w2026_ ;
	wire _w2025_ ;
	wire _w2024_ ;
	wire _w2023_ ;
	wire _w2022_ ;
	wire _w2021_ ;
	wire _w2020_ ;
	wire _w2019_ ;
	wire _w2018_ ;
	wire _w2017_ ;
	wire _w2016_ ;
	wire _w2015_ ;
	wire _w2014_ ;
	wire _w2013_ ;
	wire _w2012_ ;
	wire _w2011_ ;
	wire _w2010_ ;
	wire _w2009_ ;
	wire _w2008_ ;
	wire _w2007_ ;
	wire _w2006_ ;
	wire _w2005_ ;
	wire _w2004_ ;
	wire _w2003_ ;
	wire _w2002_ ;
	wire _w2001_ ;
	wire _w2000_ ;
	wire _w1999_ ;
	wire _w1998_ ;
	wire _w1997_ ;
	wire _w1996_ ;
	wire _w1995_ ;
	wire _w1994_ ;
	wire _w1993_ ;
	wire _w1992_ ;
	wire _w1991_ ;
	wire _w1990_ ;
	wire _w1989_ ;
	wire _w1988_ ;
	wire _w1987_ ;
	wire _w1986_ ;
	wire _w1985_ ;
	wire _w1984_ ;
	wire _w1983_ ;
	wire _w1982_ ;
	wire _w1981_ ;
	wire _w1980_ ;
	wire _w1979_ ;
	wire _w1978_ ;
	wire _w1977_ ;
	wire _w1976_ ;
	wire _w1975_ ;
	wire _w1974_ ;
	wire _w1973_ ;
	wire _w1972_ ;
	wire _w1971_ ;
	wire _w1970_ ;
	wire _w1969_ ;
	wire _w1968_ ;
	wire _w1967_ ;
	wire _w1966_ ;
	wire _w1965_ ;
	wire _w1964_ ;
	wire _w1963_ ;
	wire _w1962_ ;
	wire _w1961_ ;
	wire _w1960_ ;
	wire _w1959_ ;
	wire _w1958_ ;
	wire _w1957_ ;
	wire _w1956_ ;
	wire _w1955_ ;
	wire _w1954_ ;
	wire _w1953_ ;
	wire _w1952_ ;
	wire _w1951_ ;
	wire _w1950_ ;
	wire _w1949_ ;
	wire _w1948_ ;
	wire _w1947_ ;
	wire _w1946_ ;
	wire _w1945_ ;
	wire _w1944_ ;
	wire _w1943_ ;
	wire _w1942_ ;
	wire _w1941_ ;
	wire _w1940_ ;
	wire _w1939_ ;
	wire _w1938_ ;
	wire _w1937_ ;
	wire _w1936_ ;
	wire _w1935_ ;
	wire _w1934_ ;
	wire _w1933_ ;
	wire _w1932_ ;
	wire _w1931_ ;
	wire _w1930_ ;
	wire _w1929_ ;
	wire _w1928_ ;
	wire _w1927_ ;
	wire _w1926_ ;
	wire _w1925_ ;
	wire _w1924_ ;
	wire _w1923_ ;
	wire _w1922_ ;
	wire _w1921_ ;
	wire _w1920_ ;
	wire _w1919_ ;
	wire _w1918_ ;
	wire _w1917_ ;
	wire _w1916_ ;
	wire _w1915_ ;
	wire _w1914_ ;
	wire _w1913_ ;
	wire _w1912_ ;
	wire _w1911_ ;
	wire _w1910_ ;
	wire _w1909_ ;
	wire _w1908_ ;
	wire _w1907_ ;
	wire _w1906_ ;
	wire _w1905_ ;
	wire _w1904_ ;
	wire _w1903_ ;
	wire _w1902_ ;
	wire _w1901_ ;
	wire _w1900_ ;
	wire _w1899_ ;
	wire _w1898_ ;
	wire _w1897_ ;
	wire _w1896_ ;
	wire _w1895_ ;
	wire _w1894_ ;
	wire _w1893_ ;
	wire _w1892_ ;
	wire _w1891_ ;
	wire _w1890_ ;
	wire _w1889_ ;
	wire _w1888_ ;
	wire _w1887_ ;
	wire _w1886_ ;
	wire _w1885_ ;
	wire _w1884_ ;
	wire _w1883_ ;
	wire _w1882_ ;
	wire _w1881_ ;
	wire _w1880_ ;
	wire _w1879_ ;
	wire _w1878_ ;
	wire _w1877_ ;
	wire _w1876_ ;
	wire _w1875_ ;
	wire _w1874_ ;
	wire _w1873_ ;
	wire _w1872_ ;
	wire _w1871_ ;
	wire _w1870_ ;
	wire _w1869_ ;
	wire _w1868_ ;
	wire _w1867_ ;
	wire _w1866_ ;
	wire _w1865_ ;
	wire _w1864_ ;
	wire _w1863_ ;
	wire _w1862_ ;
	wire _w1861_ ;
	wire _w1860_ ;
	wire _w1859_ ;
	wire _w1858_ ;
	wire _w1857_ ;
	wire _w1856_ ;
	wire _w1855_ ;
	wire _w1854_ ;
	wire _w1853_ ;
	wire _w1852_ ;
	wire _w1851_ ;
	wire _w1850_ ;
	wire _w1849_ ;
	wire _w1848_ ;
	wire _w1847_ ;
	wire _w1846_ ;
	wire _w1845_ ;
	wire _w1844_ ;
	wire _w1843_ ;
	wire _w1842_ ;
	wire _w1841_ ;
	wire _w1840_ ;
	wire _w1839_ ;
	wire _w1838_ ;
	wire _w1837_ ;
	wire _w1836_ ;
	wire _w1835_ ;
	wire _w1834_ ;
	wire _w1833_ ;
	wire _w1832_ ;
	wire _w1831_ ;
	wire _w1830_ ;
	wire _w1829_ ;
	wire _w1828_ ;
	wire _w1827_ ;
	wire _w1826_ ;
	wire _w1825_ ;
	wire _w1824_ ;
	wire _w1823_ ;
	wire _w1822_ ;
	wire _w1821_ ;
	wire _w1820_ ;
	wire _w1819_ ;
	wire _w1818_ ;
	wire _w1817_ ;
	wire _w1816_ ;
	wire _w1815_ ;
	wire _w1814_ ;
	wire _w1813_ ;
	wire _w1812_ ;
	wire _w1811_ ;
	wire _w1810_ ;
	wire _w1809_ ;
	wire _w1808_ ;
	wire _w1807_ ;
	wire _w1806_ ;
	wire _w1805_ ;
	wire _w1804_ ;
	wire _w1803_ ;
	wire _w1802_ ;
	wire _w1801_ ;
	wire _w1800_ ;
	wire _w1799_ ;
	wire _w1798_ ;
	wire _w1797_ ;
	wire _w1796_ ;
	wire _w1795_ ;
	wire _w1794_ ;
	wire _w1793_ ;
	wire _w1792_ ;
	wire _w1791_ ;
	wire _w1790_ ;
	wire _w1789_ ;
	wire _w1788_ ;
	wire _w1787_ ;
	wire _w1786_ ;
	wire _w1785_ ;
	wire _w1784_ ;
	wire _w1783_ ;
	wire _w1782_ ;
	wire _w1781_ ;
	wire _w1780_ ;
	wire _w1779_ ;
	wire _w1778_ ;
	wire _w1777_ ;
	wire _w1776_ ;
	wire _w1775_ ;
	wire _w1774_ ;
	wire _w1773_ ;
	wire _w1772_ ;
	wire _w1771_ ;
	wire _w1770_ ;
	wire _w1769_ ;
	wire _w1768_ ;
	wire _w1767_ ;
	wire _w1766_ ;
	wire _w1765_ ;
	wire _w1764_ ;
	wire _w1763_ ;
	wire _w1762_ ;
	wire _w1761_ ;
	wire _w1760_ ;
	wire _w1759_ ;
	wire _w1758_ ;
	wire _w1757_ ;
	wire _w1756_ ;
	wire _w1755_ ;
	wire _w1754_ ;
	wire _w1753_ ;
	wire _w1752_ ;
	wire _w1751_ ;
	wire _w1750_ ;
	wire _w1749_ ;
	wire _w1748_ ;
	wire _w1747_ ;
	wire _w1746_ ;
	wire _w1745_ ;
	wire _w1744_ ;
	wire _w1743_ ;
	wire _w1742_ ;
	wire _w1741_ ;
	wire _w1740_ ;
	wire _w1739_ ;
	wire _w1738_ ;
	wire _w1737_ ;
	wire _w1736_ ;
	wire _w1735_ ;
	wire _w1734_ ;
	wire _w1733_ ;
	wire _w1732_ ;
	wire _w1731_ ;
	wire _w1730_ ;
	wire _w1729_ ;
	wire _w1728_ ;
	wire _w1727_ ;
	wire _w1726_ ;
	wire _w1725_ ;
	wire _w1724_ ;
	wire _w1723_ ;
	wire _w1722_ ;
	wire _w1721_ ;
	wire _w1720_ ;
	wire _w1719_ ;
	wire _w1718_ ;
	wire _w1717_ ;
	wire _w1716_ ;
	wire _w1715_ ;
	wire _w1714_ ;
	wire _w1713_ ;
	wire _w1712_ ;
	wire _w1711_ ;
	wire _w1710_ ;
	wire _w1709_ ;
	wire _w1708_ ;
	wire _w1707_ ;
	wire _w1706_ ;
	wire _w1705_ ;
	wire _w1704_ ;
	wire _w1703_ ;
	wire _w1702_ ;
	wire _w1701_ ;
	wire _w1700_ ;
	wire _w1699_ ;
	wire _w1698_ ;
	wire _w1697_ ;
	wire _w1696_ ;
	wire _w1695_ ;
	wire _w1694_ ;
	wire _w1693_ ;
	wire _w1692_ ;
	wire _w1691_ ;
	wire _w1690_ ;
	wire _w1689_ ;
	wire _w1688_ ;
	wire _w1687_ ;
	wire _w1686_ ;
	wire _w1685_ ;
	wire _w1684_ ;
	wire _w1683_ ;
	wire _w1682_ ;
	wire _w1681_ ;
	wire _w1680_ ;
	wire _w1679_ ;
	wire _w1678_ ;
	wire _w1677_ ;
	wire _w1676_ ;
	wire _w1675_ ;
	wire _w1674_ ;
	wire _w1673_ ;
	wire _w1672_ ;
	wire _w1671_ ;
	wire _w1670_ ;
	wire _w1669_ ;
	wire _w1668_ ;
	wire _w1667_ ;
	wire _w1666_ ;
	wire _w1665_ ;
	wire _w1664_ ;
	wire _w1663_ ;
	wire _w1662_ ;
	wire _w1661_ ;
	wire _w1660_ ;
	wire _w1659_ ;
	wire _w1658_ ;
	wire _w1657_ ;
	wire _w1656_ ;
	wire _w1655_ ;
	wire _w1654_ ;
	wire _w1653_ ;
	wire _w1652_ ;
	wire _w1651_ ;
	wire _w1650_ ;
	wire _w1649_ ;
	wire _w1648_ ;
	wire _w1647_ ;
	wire _w1646_ ;
	wire _w1645_ ;
	wire _w1644_ ;
	wire _w1643_ ;
	wire _w1642_ ;
	wire _w1641_ ;
	wire _w1640_ ;
	wire _w1639_ ;
	wire _w1638_ ;
	wire _w1637_ ;
	wire _w1636_ ;
	wire _w1635_ ;
	wire _w1634_ ;
	wire _w1633_ ;
	wire _w1632_ ;
	wire _w1631_ ;
	wire _w1630_ ;
	wire _w1629_ ;
	wire _w1628_ ;
	wire _w1627_ ;
	wire _w1626_ ;
	wire _w1625_ ;
	wire _w1624_ ;
	wire _w1623_ ;
	wire _w1622_ ;
	wire _w1621_ ;
	wire _w1620_ ;
	wire _w1619_ ;
	wire _w1618_ ;
	wire _w1617_ ;
	wire _w1616_ ;
	wire _w1615_ ;
	wire _w1614_ ;
	wire _w1613_ ;
	wire _w1612_ ;
	wire _w1611_ ;
	wire _w1610_ ;
	wire _w1609_ ;
	wire _w1608_ ;
	wire _w1607_ ;
	wire _w1606_ ;
	wire _w1605_ ;
	wire _w1604_ ;
	wire _w1603_ ;
	wire _w1602_ ;
	wire _w1601_ ;
	wire _w1600_ ;
	wire _w1599_ ;
	wire _w1598_ ;
	wire _w1597_ ;
	wire _w1596_ ;
	wire _w1595_ ;
	wire _w1594_ ;
	wire _w1593_ ;
	wire _w1592_ ;
	wire _w1591_ ;
	wire _w1590_ ;
	wire _w1589_ ;
	wire _w1588_ ;
	wire _w1587_ ;
	wire _w1586_ ;
	wire _w1585_ ;
	wire _w1584_ ;
	wire _w1583_ ;
	wire _w1582_ ;
	wire _w1581_ ;
	wire _w1580_ ;
	wire _w1579_ ;
	wire _w1578_ ;
	wire _w1577_ ;
	wire _w1576_ ;
	wire _w1575_ ;
	wire _w1574_ ;
	wire _w1573_ ;
	wire _w1572_ ;
	wire _w1571_ ;
	wire _w1570_ ;
	wire _w1569_ ;
	wire _w1568_ ;
	wire _w1567_ ;
	wire _w1566_ ;
	wire _w1565_ ;
	wire _w1564_ ;
	wire _w1563_ ;
	wire _w1562_ ;
	wire _w1561_ ;
	wire _w1560_ ;
	wire _w1559_ ;
	wire _w1558_ ;
	wire _w1557_ ;
	wire _w1556_ ;
	wire _w1555_ ;
	wire _w1554_ ;
	wire _w1553_ ;
	wire _w1552_ ;
	wire _w1551_ ;
	wire _w1550_ ;
	wire _w1549_ ;
	wire _w1548_ ;
	wire _w1547_ ;
	wire _w1546_ ;
	wire _w1545_ ;
	wire _w1544_ ;
	wire _w1543_ ;
	wire _w1542_ ;
	wire _w1541_ ;
	wire _w1540_ ;
	wire _w1539_ ;
	wire _w1538_ ;
	wire _w1537_ ;
	wire _w1536_ ;
	wire _w1535_ ;
	wire _w1534_ ;
	wire _w1533_ ;
	wire _w1532_ ;
	wire _w1531_ ;
	wire _w1530_ ;
	wire _w1529_ ;
	wire _w1528_ ;
	wire _w1527_ ;
	wire _w1526_ ;
	wire _w1525_ ;
	wire _w1524_ ;
	wire _w1523_ ;
	wire _w1522_ ;
	wire _w1521_ ;
	wire _w1520_ ;
	wire _w1519_ ;
	wire _w1518_ ;
	wire _w1517_ ;
	wire _w1516_ ;
	wire _w1515_ ;
	wire _w1514_ ;
	wire _w1513_ ;
	wire _w1512_ ;
	wire _w1511_ ;
	wire _w1510_ ;
	wire _w1509_ ;
	wire _w1508_ ;
	wire _w1507_ ;
	wire _w1506_ ;
	wire _w1505_ ;
	wire _w1504_ ;
	wire _w1503_ ;
	wire _w1502_ ;
	wire _w1501_ ;
	wire _w1500_ ;
	wire _w1499_ ;
	wire _w1498_ ;
	wire _w1497_ ;
	wire _w1496_ ;
	wire _w1495_ ;
	wire _w1494_ ;
	wire _w1493_ ;
	wire _w1492_ ;
	wire _w1491_ ;
	wire _w1490_ ;
	wire _w1489_ ;
	wire _w1488_ ;
	wire _w1487_ ;
	wire _w1486_ ;
	wire _w1485_ ;
	wire _w1484_ ;
	wire _w1483_ ;
	wire _w1482_ ;
	wire _w1481_ ;
	wire _w1480_ ;
	wire _w1479_ ;
	wire _w1478_ ;
	wire _w1477_ ;
	wire _w1476_ ;
	wire _w1475_ ;
	wire _w1474_ ;
	wire _w1473_ ;
	wire _w1472_ ;
	wire _w1471_ ;
	wire _w1470_ ;
	wire _w1469_ ;
	wire _w1468_ ;
	wire _w1467_ ;
	wire _w1466_ ;
	wire _w1465_ ;
	wire _w1464_ ;
	wire _w1463_ ;
	wire _w1462_ ;
	wire _w1461_ ;
	wire _w1460_ ;
	wire _w1459_ ;
	wire _w1458_ ;
	wire _w1457_ ;
	wire _w1456_ ;
	wire _w1455_ ;
	wire _w1454_ ;
	wire _w1453_ ;
	wire _w1452_ ;
	wire _w1451_ ;
	wire _w1450_ ;
	wire _w1449_ ;
	wire _w1448_ ;
	wire _w1447_ ;
	wire _w1446_ ;
	wire _w1445_ ;
	wire _w1444_ ;
	wire _w1443_ ;
	wire _w1442_ ;
	wire _w1441_ ;
	wire _w1440_ ;
	wire _w1439_ ;
	wire _w1438_ ;
	wire _w1437_ ;
	wire _w1436_ ;
	wire _w1435_ ;
	wire _w1434_ ;
	wire _w1433_ ;
	wire _w1432_ ;
	wire _w1431_ ;
	wire _w1430_ ;
	wire _w1429_ ;
	wire _w1428_ ;
	wire _w1427_ ;
	wire _w1426_ ;
	wire _w1425_ ;
	wire _w1424_ ;
	wire _w1423_ ;
	wire _w1422_ ;
	wire _w1421_ ;
	wire _w1420_ ;
	wire _w1419_ ;
	wire _w1418_ ;
	wire _w1417_ ;
	wire _w1416_ ;
	wire _w1415_ ;
	wire _w1414_ ;
	wire _w845_ ;
	wire _w844_ ;
	wire _w843_ ;
	wire _w842_ ;
	wire _w841_ ;
	wire _w840_ ;
	wire _w839_ ;
	wire _w838_ ;
	wire _w837_ ;
	wire _w836_ ;
	wire _w835_ ;
	wire _w834_ ;
	wire _w833_ ;
	wire _w832_ ;
	wire _w831_ ;
	wire _w830_ ;
	wire _w829_ ;
	wire _w828_ ;
	wire _w827_ ;
	wire _w826_ ;
	wire _w825_ ;
	wire _w824_ ;
	wire _w823_ ;
	wire _w822_ ;
	wire _w821_ ;
	wire _w820_ ;
	wire _w819_ ;
	wire _w818_ ;
	wire _w817_ ;
	wire _w816_ ;
	wire _w815_ ;
	wire _w814_ ;
	wire _w813_ ;
	wire _w812_ ;
	wire _w811_ ;
	wire _w810_ ;
	wire _w809_ ;
	wire _w808_ ;
	wire _w807_ ;
	wire _w806_ ;
	wire _w805_ ;
	wire _w804_ ;
	wire _w803_ ;
	wire _w802_ ;
	wire _w801_ ;
	wire _w800_ ;
	wire _w799_ ;
	wire _w798_ ;
	wire _w797_ ;
	wire _w796_ ;
	wire _w795_ ;
	wire _w794_ ;
	wire _w793_ ;
	wire _w792_ ;
	wire _w791_ ;
	wire _w790_ ;
	wire _w789_ ;
	wire _w788_ ;
	wire _w787_ ;
	wire _w786_ ;
	wire _w785_ ;
	wire _w784_ ;
	wire _w783_ ;
	wire _w782_ ;
	wire _w781_ ;
	wire _w780_ ;
	wire _w779_ ;
	wire _w778_ ;
	wire _w777_ ;
	wire _w776_ ;
	wire _w775_ ;
	wire _w774_ ;
	wire _w773_ ;
	wire _w772_ ;
	wire _w771_ ;
	wire _w770_ ;
	wire _w769_ ;
	wire _w768_ ;
	wire _w767_ ;
	wire _w766_ ;
	wire _w765_ ;
	wire _w764_ ;
	wire _w763_ ;
	wire _w762_ ;
	wire _w761_ ;
	wire _w760_ ;
	wire _w759_ ;
	wire _w758_ ;
	wire _w757_ ;
	wire _w756_ ;
	wire _w755_ ;
	wire _w754_ ;
	wire _w753_ ;
	wire _w752_ ;
	wire _w751_ ;
	wire _w750_ ;
	wire _w749_ ;
	wire _w748_ ;
	wire _w747_ ;
	wire _w746_ ;
	wire _w745_ ;
	wire _w744_ ;
	wire _w743_ ;
	wire _w742_ ;
	wire _w741_ ;
	wire _w740_ ;
	wire _w739_ ;
	wire _w738_ ;
	wire _w737_ ;
	wire _w736_ ;
	wire _w735_ ;
	wire _w734_ ;
	wire _w733_ ;
	wire _w732_ ;
	wire _w731_ ;
	wire _w730_ ;
	wire _w729_ ;
	wire _w728_ ;
	wire _w727_ ;
	wire _w726_ ;
	wire _w725_ ;
	wire _w724_ ;
	wire _w723_ ;
	wire _w722_ ;
	wire _w721_ ;
	wire _w720_ ;
	wire _w719_ ;
	wire _w718_ ;
	wire _w717_ ;
	wire _w716_ ;
	wire _w715_ ;
	wire _w714_ ;
	wire _w713_ ;
	wire _w712_ ;
	wire _w711_ ;
	wire _w710_ ;
	wire _w709_ ;
	wire _w708_ ;
	wire _w707_ ;
	wire _w706_ ;
	wire _w705_ ;
	wire _w704_ ;
	wire _w703_ ;
	wire _w702_ ;
	wire _w701_ ;
	wire _w700_ ;
	wire _w699_ ;
	wire _w698_ ;
	wire _w697_ ;
	wire _w696_ ;
	wire _w695_ ;
	wire _w694_ ;
	wire _w693_ ;
	wire _w692_ ;
	wire _w691_ ;
	wire _w690_ ;
	wire _w689_ ;
	wire _w688_ ;
	wire _w687_ ;
	wire _w686_ ;
	wire _w685_ ;
	wire _w684_ ;
	wire _w683_ ;
	wire _w682_ ;
	wire _w681_ ;
	wire _w680_ ;
	wire _w679_ ;
	wire _w678_ ;
	wire _w677_ ;
	wire _w676_ ;
	wire _w675_ ;
	wire _w674_ ;
	wire _w673_ ;
	wire _w672_ ;
	wire _w671_ ;
	wire _w670_ ;
	wire _w669_ ;
	wire _w668_ ;
	wire _w667_ ;
	wire _w666_ ;
	wire _w665_ ;
	wire _w664_ ;
	wire _w663_ ;
	wire _w662_ ;
	wire _w661_ ;
	wire _w660_ ;
	wire _w659_ ;
	wire _w658_ ;
	wire _w657_ ;
	wire _w656_ ;
	wire _w655_ ;
	wire _w654_ ;
	wire _w653_ ;
	wire _w652_ ;
	wire _w651_ ;
	wire _w650_ ;
	wire _w649_ ;
	wire _w648_ ;
	wire _w647_ ;
	wire _w646_ ;
	wire _w645_ ;
	wire _w644_ ;
	wire _w643_ ;
	wire _w642_ ;
	wire _w641_ ;
	wire _w640_ ;
	wire _w639_ ;
	wire _w638_ ;
	wire _w637_ ;
	wire _w636_ ;
	wire _w635_ ;
	wire _w634_ ;
	wire _w633_ ;
	wire _w632_ ;
	wire _w631_ ;
	wire _w630_ ;
	wire _w629_ ;
	wire _w628_ ;
	wire _w627_ ;
	wire _w626_ ;
	wire _w625_ ;
	wire _w624_ ;
	wire _w623_ ;
	wire _w622_ ;
	wire _w621_ ;
	wire _w620_ ;
	wire _w619_ ;
	wire _w618_ ;
	wire _w617_ ;
	wire _w616_ ;
	wire _w615_ ;
	wire _w614_ ;
	wire _w613_ ;
	wire _w612_ ;
	wire _w611_ ;
	wire _w610_ ;
	wire _w609_ ;
	wire _w608_ ;
	wire _w607_ ;
	wire _w606_ ;
	wire _w605_ ;
	wire _w604_ ;
	wire _w603_ ;
	wire _w602_ ;
	wire _w601_ ;
	wire _w600_ ;
	wire _w599_ ;
	wire _w598_ ;
	wire _w597_ ;
	wire _w596_ ;
	wire _w595_ ;
	wire _w594_ ;
	wire _w593_ ;
	wire _w592_ ;
	wire _w591_ ;
	wire _w590_ ;
	wire _w589_ ;
	wire _w588_ ;
	wire _w587_ ;
	wire _w586_ ;
	wire _w585_ ;
	wire _w584_ ;
	wire _w583_ ;
	wire _w582_ ;
	wire _w581_ ;
	wire _w580_ ;
	wire _w579_ ;
	wire _w578_ ;
	wire _w577_ ;
	wire _w576_ ;
	wire _w575_ ;
	wire _w574_ ;
	wire _w573_ ;
	wire _w572_ ;
	wire _w571_ ;
	wire _w570_ ;
	wire _w569_ ;
	wire _w568_ ;
	wire _w567_ ;
	wire _w566_ ;
	wire _w565_ ;
	wire _w564_ ;
	wire _w563_ ;
	wire _w562_ ;
	wire _w431_ ;
	wire _w430_ ;
	wire _w429_ ;
	wire _w428_ ;
	wire _w427_ ;
	wire _w426_ ;
	wire _w425_ ;
	wire _w424_ ;
	wire _w423_ ;
	wire _w422_ ;
	wire _w421_ ;
	wire _w420_ ;
	wire _w419_ ;
	wire _w418_ ;
	wire _w417_ ;
	wire _w416_ ;
	wire _w415_ ;
	wire _w414_ ;
	wire _w413_ ;
	wire _w412_ ;
	wire _w411_ ;
	wire _w410_ ;
	wire _w409_ ;
	wire _w408_ ;
	wire _w407_ ;
	wire _w406_ ;
	wire _w405_ ;
	wire _w404_ ;
	wire _w403_ ;
	wire _w402_ ;
	wire _w401_ ;
	wire _w400_ ;
	wire _w399_ ;
	wire _w398_ ;
	wire _w397_ ;
	wire _w396_ ;
	wire _w395_ ;
	wire _w394_ ;
	wire _w393_ ;
	wire _w392_ ;
	wire _w391_ ;
	wire _w390_ ;
	wire _w389_ ;
	wire _w388_ ;
	wire _w387_ ;
	wire _w386_ ;
	wire _w385_ ;
	wire _w384_ ;
	wire _w383_ ;
	wire _w382_ ;
	wire _w381_ ;
	wire _w380_ ;
	wire _w379_ ;
	wire _w378_ ;
	wire _w377_ ;
	wire _w376_ ;
	wire _w375_ ;
	wire _w374_ ;
	wire _w373_ ;
	wire _w372_ ;
	wire _w371_ ;
	wire _w370_ ;
	wire _w369_ ;
	wire _w368_ ;
	wire _w367_ ;
	wire _w366_ ;
	wire _w365_ ;
	wire _w364_ ;
	wire _w333_ ;
	wire _w332_ ;
	wire _w331_ ;
	wire _w330_ ;
	wire _w329_ ;
	wire _w328_ ;
	wire _w327_ ;
	wire _w326_ ;
	wire _w325_ ;
	wire _w324_ ;
	wire _w323_ ;
	wire _w322_ ;
	wire _w321_ ;
	wire _w320_ ;
	wire _w319_ ;
	wire _w318_ ;
	wire _w305_ ;
	wire _w306_ ;
	wire _w307_ ;
	wire _w308_ ;
	wire _w309_ ;
	wire _w310_ ;
	wire _w311_ ;
	wire _w312_ ;
	wire _w313_ ;
	wire _w314_ ;
	wire _w315_ ;
	wire _w316_ ;
	wire _w317_ ;
	wire _w334_ ;
	wire _w335_ ;
	wire _w336_ ;
	wire _w337_ ;
	wire _w338_ ;
	wire _w339_ ;
	wire _w340_ ;
	wire _w341_ ;
	wire _w342_ ;
	wire _w343_ ;
	wire _w344_ ;
	wire _w345_ ;
	wire _w346_ ;
	wire _w347_ ;
	wire _w348_ ;
	wire _w349_ ;
	wire _w350_ ;
	wire _w351_ ;
	wire _w352_ ;
	wire _w353_ ;
	wire _w354_ ;
	wire _w355_ ;
	wire _w356_ ;
	wire _w357_ ;
	wire _w358_ ;
	wire _w359_ ;
	wire _w360_ ;
	wire _w361_ ;
	wire _w362_ ;
	wire _w363_ ;
	wire _w432_ ;
	wire _w433_ ;
	wire _w434_ ;
	wire _w435_ ;
	wire _w436_ ;
	wire _w437_ ;
	wire _w438_ ;
	wire _w439_ ;
	wire _w440_ ;
	wire _w441_ ;
	wire _w442_ ;
	wire _w443_ ;
	wire _w444_ ;
	wire _w445_ ;
	wire _w446_ ;
	wire _w447_ ;
	wire _w448_ ;
	wire _w449_ ;
	wire _w450_ ;
	wire _w451_ ;
	wire _w452_ ;
	wire _w453_ ;
	wire _w454_ ;
	wire _w455_ ;
	wire _w456_ ;
	wire _w457_ ;
	wire _w458_ ;
	wire _w459_ ;
	wire _w460_ ;
	wire _w461_ ;
	wire _w462_ ;
	wire _w463_ ;
	wire _w464_ ;
	wire _w465_ ;
	wire _w466_ ;
	wire _w467_ ;
	wire _w468_ ;
	wire _w469_ ;
	wire _w470_ ;
	wire _w471_ ;
	wire _w472_ ;
	wire _w473_ ;
	wire _w474_ ;
	wire _w475_ ;
	wire _w476_ ;
	wire _w477_ ;
	wire _w478_ ;
	wire _w479_ ;
	wire _w480_ ;
	wire _w481_ ;
	wire _w482_ ;
	wire _w483_ ;
	wire _w484_ ;
	wire _w485_ ;
	wire _w486_ ;
	wire _w487_ ;
	wire _w488_ ;
	wire _w489_ ;
	wire _w490_ ;
	wire _w491_ ;
	wire _w492_ ;
	wire _w493_ ;
	wire _w494_ ;
	wire _w495_ ;
	wire _w496_ ;
	wire _w497_ ;
	wire _w498_ ;
	wire _w499_ ;
	wire _w500_ ;
	wire _w501_ ;
	wire _w502_ ;
	wire _w503_ ;
	wire _w504_ ;
	wire _w505_ ;
	wire _w506_ ;
	wire _w507_ ;
	wire _w508_ ;
	wire _w509_ ;
	wire _w510_ ;
	wire _w511_ ;
	wire _w512_ ;
	wire _w513_ ;
	wire _w514_ ;
	wire _w515_ ;
	wire _w516_ ;
	wire _w517_ ;
	wire _w518_ ;
	wire _w519_ ;
	wire _w520_ ;
	wire _w521_ ;
	wire _w522_ ;
	wire _w523_ ;
	wire _w524_ ;
	wire _w525_ ;
	wire _w526_ ;
	wire _w527_ ;
	wire _w528_ ;
	wire _w529_ ;
	wire _w530_ ;
	wire _w531_ ;
	wire _w532_ ;
	wire _w533_ ;
	wire _w534_ ;
	wire _w535_ ;
	wire _w536_ ;
	wire _w537_ ;
	wire _w538_ ;
	wire _w539_ ;
	wire _w540_ ;
	wire _w541_ ;
	wire _w542_ ;
	wire _w543_ ;
	wire _w544_ ;
	wire _w545_ ;
	wire _w546_ ;
	wire _w547_ ;
	wire _w548_ ;
	wire _w549_ ;
	wire _w550_ ;
	wire _w551_ ;
	wire _w552_ ;
	wire _w553_ ;
	wire _w554_ ;
	wire _w555_ ;
	wire _w556_ ;
	wire _w557_ ;
	wire _w558_ ;
	wire _w559_ ;
	wire _w560_ ;
	wire _w561_ ;
	wire _w846_ ;
	wire _w847_ ;
	wire _w848_ ;
	wire _w849_ ;
	wire _w850_ ;
	wire _w851_ ;
	wire _w852_ ;
	wire _w853_ ;
	wire _w854_ ;
	wire _w855_ ;
	wire _w856_ ;
	wire _w857_ ;
	wire _w858_ ;
	wire _w859_ ;
	wire _w860_ ;
	wire _w861_ ;
	wire _w862_ ;
	wire _w863_ ;
	wire _w864_ ;
	wire _w865_ ;
	wire _w866_ ;
	wire _w867_ ;
	wire _w868_ ;
	wire _w869_ ;
	wire _w870_ ;
	wire _w871_ ;
	wire _w872_ ;
	wire _w873_ ;
	wire _w874_ ;
	wire _w875_ ;
	wire _w876_ ;
	wire _w877_ ;
	wire _w878_ ;
	wire _w879_ ;
	wire _w880_ ;
	wire _w881_ ;
	wire _w882_ ;
	wire _w883_ ;
	wire _w884_ ;
	wire _w885_ ;
	wire _w886_ ;
	wire _w887_ ;
	wire _w888_ ;
	wire _w889_ ;
	wire _w890_ ;
	wire _w891_ ;
	wire _w892_ ;
	wire _w893_ ;
	wire _w894_ ;
	wire _w895_ ;
	wire _w896_ ;
	wire _w897_ ;
	wire _w898_ ;
	wire _w899_ ;
	wire _w900_ ;
	wire _w901_ ;
	wire _w902_ ;
	wire _w903_ ;
	wire _w904_ ;
	wire _w905_ ;
	wire _w906_ ;
	wire _w907_ ;
	wire _w908_ ;
	wire _w909_ ;
	wire _w910_ ;
	wire _w911_ ;
	wire _w912_ ;
	wire _w913_ ;
	wire _w914_ ;
	wire _w915_ ;
	wire _w916_ ;
	wire _w917_ ;
	wire _w918_ ;
	wire _w919_ ;
	wire _w920_ ;
	wire _w921_ ;
	wire _w922_ ;
	wire _w923_ ;
	wire _w924_ ;
	wire _w925_ ;
	wire _w926_ ;
	wire _w927_ ;
	wire _w928_ ;
	wire _w929_ ;
	wire _w930_ ;
	wire _w931_ ;
	wire _w932_ ;
	wire _w933_ ;
	wire _w934_ ;
	wire _w935_ ;
	wire _w936_ ;
	wire _w937_ ;
	wire _w938_ ;
	wire _w939_ ;
	wire _w940_ ;
	wire _w941_ ;
	wire _w942_ ;
	wire _w943_ ;
	wire _w944_ ;
	wire _w945_ ;
	wire _w946_ ;
	wire _w947_ ;
	wire _w948_ ;
	wire _w949_ ;
	wire _w950_ ;
	wire _w951_ ;
	wire _w952_ ;
	wire _w953_ ;
	wire _w954_ ;
	wire _w955_ ;
	wire _w956_ ;
	wire _w957_ ;
	wire _w958_ ;
	wire _w959_ ;
	wire _w960_ ;
	wire _w961_ ;
	wire _w962_ ;
	wire _w963_ ;
	wire _w964_ ;
	wire _w965_ ;
	wire _w966_ ;
	wire _w967_ ;
	wire _w968_ ;
	wire _w969_ ;
	wire _w970_ ;
	wire _w971_ ;
	wire _w972_ ;
	wire _w973_ ;
	wire _w974_ ;
	wire _w975_ ;
	wire _w976_ ;
	wire _w977_ ;
	wire _w978_ ;
	wire _w979_ ;
	wire _w980_ ;
	wire _w981_ ;
	wire _w982_ ;
	wire _w983_ ;
	wire _w984_ ;
	wire _w985_ ;
	wire _w986_ ;
	wire _w987_ ;
	wire _w988_ ;
	wire _w989_ ;
	wire _w990_ ;
	wire _w991_ ;
	wire _w992_ ;
	wire _w993_ ;
	wire _w994_ ;
	wire _w995_ ;
	wire _w996_ ;
	wire _w997_ ;
	wire _w998_ ;
	wire _w999_ ;
	wire _w1000_ ;
	wire _w1001_ ;
	wire _w1002_ ;
	wire _w1003_ ;
	wire _w1004_ ;
	wire _w1005_ ;
	wire _w1006_ ;
	wire _w1007_ ;
	wire _w1008_ ;
	wire _w1009_ ;
	wire _w1010_ ;
	wire _w1011_ ;
	wire _w1012_ ;
	wire _w1013_ ;
	wire _w1014_ ;
	wire _w1015_ ;
	wire _w1016_ ;
	wire _w1017_ ;
	wire _w1018_ ;
	wire _w1019_ ;
	wire _w1020_ ;
	wire _w1021_ ;
	wire _w1022_ ;
	wire _w1023_ ;
	wire _w1024_ ;
	wire _w1025_ ;
	wire _w1026_ ;
	wire _w1027_ ;
	wire _w1028_ ;
	wire _w1029_ ;
	wire _w1030_ ;
	wire _w1031_ ;
	wire _w1032_ ;
	wire _w1033_ ;
	wire _w1034_ ;
	wire _w1035_ ;
	wire _w1036_ ;
	wire _w1037_ ;
	wire _w1038_ ;
	wire _w1039_ ;
	wire _w1040_ ;
	wire _w1041_ ;
	wire _w1042_ ;
	wire _w1043_ ;
	wire _w1044_ ;
	wire _w1045_ ;
	wire _w1046_ ;
	wire _w1047_ ;
	wire _w1048_ ;
	wire _w1049_ ;
	wire _w1050_ ;
	wire _w1051_ ;
	wire _w1052_ ;
	wire _w1053_ ;
	wire _w1054_ ;
	wire _w1055_ ;
	wire _w1056_ ;
	wire _w1057_ ;
	wire _w1058_ ;
	wire _w1059_ ;
	wire _w1060_ ;
	wire _w1061_ ;
	wire _w1062_ ;
	wire _w1063_ ;
	wire _w1064_ ;
	wire _w1065_ ;
	wire _w1066_ ;
	wire _w1067_ ;
	wire _w1068_ ;
	wire _w1069_ ;
	wire _w1070_ ;
	wire _w1071_ ;
	wire _w1072_ ;
	wire _w1073_ ;
	wire _w1074_ ;
	wire _w1075_ ;
	wire _w1076_ ;
	wire _w1077_ ;
	wire _w1078_ ;
	wire _w1079_ ;
	wire _w1080_ ;
	wire _w1081_ ;
	wire _w1082_ ;
	wire _w1083_ ;
	wire _w1084_ ;
	wire _w1085_ ;
	wire _w1086_ ;
	wire _w1087_ ;
	wire _w1088_ ;
	wire _w1089_ ;
	wire _w1090_ ;
	wire _w1091_ ;
	wire _w1092_ ;
	wire _w1093_ ;
	wire _w1094_ ;
	wire _w1095_ ;
	wire _w1096_ ;
	wire _w1097_ ;
	wire _w1098_ ;
	wire _w1099_ ;
	wire _w1100_ ;
	wire _w1101_ ;
	wire _w1102_ ;
	wire _w1103_ ;
	wire _w1104_ ;
	wire _w1105_ ;
	wire _w1106_ ;
	wire _w1107_ ;
	wire _w1108_ ;
	wire _w1109_ ;
	wire _w1110_ ;
	wire _w1111_ ;
	wire _w1112_ ;
	wire _w1113_ ;
	wire _w1114_ ;
	wire _w1115_ ;
	wire _w1116_ ;
	wire _w1117_ ;
	wire _w1118_ ;
	wire _w1119_ ;
	wire _w1120_ ;
	wire _w1121_ ;
	wire _w1122_ ;
	wire _w1123_ ;
	wire _w1124_ ;
	wire _w1125_ ;
	wire _w1126_ ;
	wire _w1127_ ;
	wire _w1128_ ;
	wire _w1129_ ;
	wire _w1130_ ;
	wire _w1131_ ;
	wire _w1132_ ;
	wire _w1133_ ;
	wire _w1134_ ;
	wire _w1135_ ;
	wire _w1136_ ;
	wire _w1137_ ;
	wire _w1138_ ;
	wire _w1139_ ;
	wire _w1140_ ;
	wire _w1141_ ;
	wire _w1142_ ;
	wire _w1143_ ;
	wire _w1144_ ;
	wire _w1145_ ;
	wire _w1146_ ;
	wire _w1147_ ;
	wire _w1148_ ;
	wire _w1149_ ;
	wire _w1150_ ;
	wire _w1151_ ;
	wire _w1152_ ;
	wire _w1153_ ;
	wire _w1154_ ;
	wire _w1155_ ;
	wire _w1156_ ;
	wire _w1157_ ;
	wire _w1158_ ;
	wire _w1159_ ;
	wire _w1160_ ;
	wire _w1161_ ;
	wire _w1162_ ;
	wire _w1163_ ;
	wire _w1164_ ;
	wire _w1165_ ;
	wire _w1166_ ;
	wire _w1167_ ;
	wire _w1168_ ;
	wire _w1169_ ;
	wire _w1170_ ;
	wire _w1171_ ;
	wire _w1172_ ;
	wire _w1173_ ;
	wire _w1174_ ;
	wire _w1175_ ;
	wire _w1176_ ;
	wire _w1177_ ;
	wire _w1178_ ;
	wire _w1179_ ;
	wire _w1180_ ;
	wire _w1181_ ;
	wire _w1182_ ;
	wire _w1183_ ;
	wire _w1184_ ;
	wire _w1185_ ;
	wire _w1186_ ;
	wire _w1187_ ;
	wire _w1188_ ;
	wire _w1189_ ;
	wire _w1190_ ;
	wire _w1191_ ;
	wire _w1192_ ;
	wire _w1193_ ;
	wire _w1194_ ;
	wire _w1195_ ;
	wire _w1196_ ;
	wire _w1197_ ;
	wire _w1198_ ;
	wire _w1199_ ;
	wire _w1200_ ;
	wire _w1201_ ;
	wire _w1202_ ;
	wire _w1203_ ;
	wire _w1204_ ;
	wire _w1205_ ;
	wire _w1206_ ;
	wire _w1207_ ;
	wire _w1208_ ;
	wire _w1209_ ;
	wire _w1210_ ;
	wire _w1211_ ;
	wire _w1212_ ;
	wire _w1213_ ;
	wire _w1214_ ;
	wire _w1215_ ;
	wire _w1216_ ;
	wire _w1217_ ;
	wire _w1218_ ;
	wire _w1219_ ;
	wire _w1220_ ;
	wire _w1221_ ;
	wire _w1222_ ;
	wire _w1223_ ;
	wire _w1224_ ;
	wire _w1225_ ;
	wire _w1226_ ;
	wire _w1227_ ;
	wire _w1228_ ;
	wire _w1229_ ;
	wire _w1230_ ;
	wire _w1231_ ;
	wire _w1232_ ;
	wire _w1233_ ;
	wire _w1234_ ;
	wire _w1235_ ;
	wire _w1236_ ;
	wire _w1237_ ;
	wire _w1238_ ;
	wire _w1239_ ;
	wire _w1240_ ;
	wire _w1241_ ;
	wire _w1242_ ;
	wire _w1243_ ;
	wire _w1244_ ;
	wire _w1245_ ;
	wire _w1246_ ;
	wire _w1247_ ;
	wire _w1248_ ;
	wire _w1249_ ;
	wire _w1250_ ;
	wire _w1251_ ;
	wire _w1252_ ;
	wire _w1253_ ;
	wire _w1254_ ;
	wire _w1255_ ;
	wire _w1256_ ;
	wire _w1257_ ;
	wire _w1258_ ;
	wire _w1259_ ;
	wire _w1260_ ;
	wire _w1261_ ;
	wire _w1262_ ;
	wire _w1263_ ;
	wire _w1264_ ;
	wire _w1265_ ;
	wire _w1266_ ;
	wire _w1267_ ;
	wire _w1268_ ;
	wire _w1269_ ;
	wire _w1270_ ;
	wire _w1271_ ;
	wire _w1272_ ;
	wire _w1273_ ;
	wire _w1274_ ;
	wire _w1275_ ;
	wire _w1276_ ;
	wire _w1277_ ;
	wire _w1278_ ;
	wire _w1279_ ;
	wire _w1280_ ;
	wire _w1281_ ;
	wire _w1282_ ;
	wire _w1283_ ;
	wire _w1284_ ;
	wire _w1285_ ;
	wire _w1286_ ;
	wire _w1287_ ;
	wire _w1288_ ;
	wire _w1289_ ;
	wire _w1290_ ;
	wire _w1291_ ;
	wire _w1292_ ;
	wire _w1293_ ;
	wire _w1294_ ;
	wire _w1295_ ;
	wire _w1296_ ;
	wire _w1297_ ;
	wire _w1298_ ;
	wire _w1299_ ;
	wire _w1300_ ;
	wire _w1301_ ;
	wire _w1302_ ;
	wire _w1303_ ;
	wire _w1304_ ;
	wire _w1305_ ;
	wire _w1306_ ;
	wire _w1307_ ;
	wire _w1308_ ;
	wire _w1309_ ;
	wire _w1310_ ;
	wire _w1311_ ;
	wire _w1312_ ;
	wire _w1313_ ;
	wire _w1314_ ;
	wire _w1315_ ;
	wire _w1316_ ;
	wire _w1317_ ;
	wire _w1318_ ;
	wire _w1319_ ;
	wire _w1320_ ;
	wire _w1321_ ;
	wire _w1322_ ;
	wire _w1323_ ;
	wire _w1324_ ;
	wire _w1325_ ;
	wire _w1326_ ;
	wire _w1327_ ;
	wire _w1328_ ;
	wire _w1329_ ;
	wire _w1330_ ;
	wire _w1331_ ;
	wire _w1332_ ;
	wire _w1333_ ;
	wire _w1334_ ;
	wire _w1335_ ;
	wire _w1336_ ;
	wire _w1337_ ;
	wire _w1338_ ;
	wire _w1339_ ;
	wire _w1340_ ;
	wire _w1341_ ;
	wire _w1342_ ;
	wire _w1343_ ;
	wire _w1344_ ;
	wire _w1345_ ;
	wire _w1346_ ;
	wire _w1347_ ;
	wire _w1348_ ;
	wire _w1349_ ;
	wire _w1350_ ;
	wire _w1351_ ;
	wire _w1352_ ;
	wire _w1353_ ;
	wire _w1354_ ;
	wire _w1355_ ;
	wire _w1356_ ;
	wire _w1357_ ;
	wire _w1358_ ;
	wire _w1359_ ;
	wire _w1360_ ;
	wire _w1361_ ;
	wire _w1362_ ;
	wire _w1363_ ;
	wire _w1364_ ;
	wire _w1365_ ;
	wire _w1366_ ;
	wire _w1367_ ;
	wire _w1368_ ;
	wire _w1369_ ;
	wire _w1370_ ;
	wire _w1371_ ;
	wire _w1372_ ;
	wire _w1373_ ;
	wire _w1374_ ;
	wire _w1375_ ;
	wire _w1376_ ;
	wire _w1377_ ;
	wire _w1378_ ;
	wire _w1379_ ;
	wire _w1380_ ;
	wire _w1381_ ;
	wire _w1382_ ;
	wire _w1383_ ;
	wire _w1384_ ;
	wire _w1385_ ;
	wire _w1386_ ;
	wire _w1387_ ;
	wire _w1388_ ;
	wire _w1389_ ;
	wire _w1390_ ;
	wire _w1391_ ;
	wire _w1392_ ;
	wire _w1393_ ;
	wire _w1394_ ;
	wire _w1395_ ;
	wire _w1396_ ;
	wire _w1397_ ;
	wire _w1398_ ;
	wire _w1399_ ;
	wire _w1400_ ;
	wire _w1401_ ;
	wire _w1402_ ;
	wire _w1403_ ;
	wire _w1404_ ;
	wire _w1405_ ;
	wire _w1406_ ;
	wire _w1407_ ;
	wire _w1408_ ;
	wire _w1409_ ;
	wire _w1410_ ;
	wire _w1411_ ;
	wire _w1412_ ;
	wire _w1413_ ;
	LUT4 #(
		.INIT('h0001)
	) name0 (
		\roundSel[0]_pad ,
		\roundSel[1]_pad ,
		\roundSel[2]_pad ,
		\roundSel[3]_pad ,
		_w305_
	);
	LUT4 #(
		.INIT('h0200)
	) name1 (
		\desIn[27]_pad ,
		\roundSel[4]_pad ,
		\roundSel[5]_pad ,
		_w305_,
		_w306_
	);
	LUT2 #(
		.INIT('h4)
	) name2 (
		\roundSel[4]_pad ,
		\roundSel[5]_pad ,
		_w307_
	);
	LUT4 #(
		.INIT('h4155)
	) name3 (
		\FP_R_reg[20]/P0001 ,
		\roundSel[4]_pad ,
		\roundSel[5]_pad ,
		_w305_,
		_w308_
	);
	LUT4 #(
		.INIT('he8ff)
	) name4 (
		\FP_R_reg[52]/NET0131 ,
		\roundSel[4]_pad ,
		\roundSel[5]_pad ,
		_w305_,
		_w309_
	);
	LUT3 #(
		.INIT('h45)
	) name5 (
		_w306_,
		_w308_,
		_w309_,
		_w310_
	);
	LUT3 #(
		.INIT('hba)
	) name6 (
		_w306_,
		_w308_,
		_w309_,
		_w311_
	);
	LUT4 #(
		.INIT('h0002)
	) name7 (
		\roundSel[0]_pad ,
		\roundSel[1]_pad ,
		\roundSel[2]_pad ,
		\roundSel[3]_pad ,
		_w312_
	);
	LUT3 #(
		.INIT('h59)
	) name8 (
		decrypt_pad,
		\roundSel[4]_pad ,
		\roundSel[5]_pad ,
		_w313_
	);
	LUT4 #(
		.INIT('h0408)
	) name9 (
		decrypt_pad,
		\key3[30]_pad ,
		\roundSel[4]_pad ,
		\roundSel[5]_pad ,
		_w314_
	);
	LUT3 #(
		.INIT('h08)
	) name10 (
		\key2[30]_pad ,
		\roundSel[4]_pad ,
		\roundSel[5]_pad ,
		_w315_
	);
	LUT4 #(
		.INIT('h0804)
	) name11 (
		decrypt_pad,
		\key1[30]_pad ,
		\roundSel[4]_pad ,
		\roundSel[5]_pad ,
		_w316_
	);
	LUT4 #(
		.INIT('haaa8)
	) name12 (
		_w313_,
		_w315_,
		_w316_,
		_w314_,
		_w317_
	);
	LUT4 #(
		.INIT('h0408)
	) name13 (
		decrypt_pad,
		\key3[9]_pad ,
		\roundSel[4]_pad ,
		\roundSel[5]_pad ,
		_w318_
	);
	LUT3 #(
		.INIT('h08)
	) name14 (
		\key2[9]_pad ,
		\roundSel[4]_pad ,
		\roundSel[5]_pad ,
		_w319_
	);
	LUT4 #(
		.INIT('h0804)
	) name15 (
		decrypt_pad,
		\key1[9]_pad ,
		\roundSel[4]_pad ,
		\roundSel[5]_pad ,
		_w320_
	);
	LUT4 #(
		.INIT('h5554)
	) name16 (
		_w313_,
		_w319_,
		_w320_,
		_w318_,
		_w321_
	);
	LUT3 #(
		.INIT('ha8)
	) name17 (
		_w312_,
		_w317_,
		_w321_,
		_w322_
	);
	LUT4 #(
		.INIT('h0040)
	) name18 (
		\roundSel[0]_pad ,
		\roundSel[1]_pad ,
		\roundSel[2]_pad ,
		\roundSel[3]_pad ,
		_w323_
	);
	LUT4 #(
		.INIT('h0408)
	) name19 (
		decrypt_pad,
		\key3[49]_pad ,
		\roundSel[4]_pad ,
		\roundSel[5]_pad ,
		_w324_
	);
	LUT3 #(
		.INIT('h08)
	) name20 (
		\key2[49]_pad ,
		\roundSel[4]_pad ,
		\roundSel[5]_pad ,
		_w325_
	);
	LUT4 #(
		.INIT('h0804)
	) name21 (
		decrypt_pad,
		\key1[49]_pad ,
		\roundSel[4]_pad ,
		\roundSel[5]_pad ,
		_w326_
	);
	LUT4 #(
		.INIT('h5554)
	) name22 (
		_w313_,
		_w325_,
		_w326_,
		_w324_,
		_w327_
	);
	LUT4 #(
		.INIT('h0408)
	) name23 (
		decrypt_pad,
		\key3[14]_pad ,
		\roundSel[4]_pad ,
		\roundSel[5]_pad ,
		_w328_
	);
	LUT3 #(
		.INIT('h08)
	) name24 (
		\key2[14]_pad ,
		\roundSel[4]_pad ,
		\roundSel[5]_pad ,
		_w329_
	);
	LUT4 #(
		.INIT('h0804)
	) name25 (
		decrypt_pad,
		\key1[14]_pad ,
		\roundSel[4]_pad ,
		\roundSel[5]_pad ,
		_w330_
	);
	LUT4 #(
		.INIT('haaa8)
	) name26 (
		_w313_,
		_w329_,
		_w330_,
		_w328_,
		_w331_
	);
	LUT3 #(
		.INIT('ha8)
	) name27 (
		_w323_,
		_w327_,
		_w331_,
		_w332_
	);
	LUT4 #(
		.INIT('h0020)
	) name28 (
		\roundSel[0]_pad ,
		\roundSel[1]_pad ,
		\roundSel[2]_pad ,
		\roundSel[3]_pad ,
		_w333_
	);
	LUT4 #(
		.INIT('h0408)
	) name29 (
		decrypt_pad,
		\key3[8]_pad ,
		\roundSel[4]_pad ,
		\roundSel[5]_pad ,
		_w334_
	);
	LUT3 #(
		.INIT('h08)
	) name30 (
		\key2[8]_pad ,
		\roundSel[4]_pad ,
		\roundSel[5]_pad ,
		_w335_
	);
	LUT4 #(
		.INIT('h0804)
	) name31 (
		decrypt_pad,
		\key1[8]_pad ,
		\roundSel[4]_pad ,
		\roundSel[5]_pad ,
		_w336_
	);
	LUT4 #(
		.INIT('h5554)
	) name32 (
		_w313_,
		_w335_,
		_w336_,
		_w334_,
		_w337_
	);
	LUT4 #(
		.INIT('h0408)
	) name33 (
		decrypt_pad,
		\key3[0]_pad ,
		\roundSel[4]_pad ,
		\roundSel[5]_pad ,
		_w338_
	);
	LUT3 #(
		.INIT('h08)
	) name34 (
		\key2[0]_pad ,
		\roundSel[4]_pad ,
		\roundSel[5]_pad ,
		_w339_
	);
	LUT4 #(
		.INIT('h0804)
	) name35 (
		decrypt_pad,
		\key1[0]_pad ,
		\roundSel[4]_pad ,
		\roundSel[5]_pad ,
		_w340_
	);
	LUT4 #(
		.INIT('haaa8)
	) name36 (
		_w313_,
		_w339_,
		_w340_,
		_w338_,
		_w341_
	);
	LUT3 #(
		.INIT('ha8)
	) name37 (
		_w333_,
		_w337_,
		_w341_,
		_w342_
	);
	LUT4 #(
		.INIT('h0010)
	) name38 (
		\roundSel[0]_pad ,
		\roundSel[1]_pad ,
		\roundSel[2]_pad ,
		\roundSel[3]_pad ,
		_w343_
	);
	LUT4 #(
		.INIT('h0408)
	) name39 (
		decrypt_pad,
		\key3[45]_pad ,
		\roundSel[4]_pad ,
		\roundSel[5]_pad ,
		_w344_
	);
	LUT3 #(
		.INIT('h08)
	) name40 (
		\key2[45]_pad ,
		\roundSel[4]_pad ,
		\roundSel[5]_pad ,
		_w345_
	);
	LUT4 #(
		.INIT('h0804)
	) name41 (
		decrypt_pad,
		\key1[45]_pad ,
		\roundSel[4]_pad ,
		\roundSel[5]_pad ,
		_w346_
	);
	LUT4 #(
		.INIT('haaa8)
	) name42 (
		_w313_,
		_w345_,
		_w346_,
		_w344_,
		_w347_
	);
	LUT4 #(
		.INIT('h0408)
	) name43 (
		decrypt_pad,
		\key3[22]_pad ,
		\roundSel[4]_pad ,
		\roundSel[5]_pad ,
		_w348_
	);
	LUT3 #(
		.INIT('h08)
	) name44 (
		\key2[22]_pad ,
		\roundSel[4]_pad ,
		\roundSel[5]_pad ,
		_w349_
	);
	LUT4 #(
		.INIT('h0804)
	) name45 (
		decrypt_pad,
		\key1[22]_pad ,
		\roundSel[4]_pad ,
		\roundSel[5]_pad ,
		_w350_
	);
	LUT4 #(
		.INIT('h5554)
	) name46 (
		_w313_,
		_w349_,
		_w350_,
		_w348_,
		_w351_
	);
	LUT3 #(
		.INIT('ha8)
	) name47 (
		_w343_,
		_w347_,
		_w351_,
		_w352_
	);
	LUT4 #(
		.INIT('h0001)
	) name48 (
		_w322_,
		_w332_,
		_w342_,
		_w352_,
		_w353_
	);
	LUT4 #(
		.INIT('h0408)
	) name49 (
		decrypt_pad,
		\key3[16]_pad ,
		\roundSel[4]_pad ,
		\roundSel[5]_pad ,
		_w354_
	);
	LUT3 #(
		.INIT('h08)
	) name50 (
		\key2[16]_pad ,
		\roundSel[4]_pad ,
		\roundSel[5]_pad ,
		_w355_
	);
	LUT4 #(
		.INIT('h0804)
	) name51 (
		decrypt_pad,
		\key1[16]_pad ,
		\roundSel[4]_pad ,
		\roundSel[5]_pad ,
		_w356_
	);
	LUT4 #(
		.INIT('h5554)
	) name52 (
		_w313_,
		_w355_,
		_w356_,
		_w354_,
		_w357_
	);
	LUT4 #(
		.INIT('h0408)
	) name53 (
		decrypt_pad,
		\key3[23]_pad ,
		\roundSel[4]_pad ,
		\roundSel[5]_pad ,
		_w358_
	);
	LUT3 #(
		.INIT('h08)
	) name54 (
		\key2[23]_pad ,
		\roundSel[4]_pad ,
		\roundSel[5]_pad ,
		_w359_
	);
	LUT4 #(
		.INIT('h0804)
	) name55 (
		decrypt_pad,
		\key1[23]_pad ,
		\roundSel[4]_pad ,
		\roundSel[5]_pad ,
		_w360_
	);
	LUT4 #(
		.INIT('haaa8)
	) name56 (
		_w313_,
		_w359_,
		_w360_,
		_w358_,
		_w361_
	);
	LUT3 #(
		.INIT('ha8)
	) name57 (
		_w305_,
		_w357_,
		_w361_,
		_w362_
	);
	LUT4 #(
		.INIT('h2000)
	) name58 (
		\roundSel[0]_pad ,
		\roundSel[1]_pad ,
		\roundSel[2]_pad ,
		\roundSel[3]_pad ,
		_w363_
	);
	LUT4 #(
		.INIT('h0408)
	) name59 (
		decrypt_pad,
		\key3[44]_pad ,
		\roundSel[4]_pad ,
		\roundSel[5]_pad ,
		_w364_
	);
	LUT3 #(
		.INIT('h08)
	) name60 (
		\key2[44]_pad ,
		\roundSel[4]_pad ,
		\roundSel[5]_pad ,
		_w365_
	);
	LUT4 #(
		.INIT('h0804)
	) name61 (
		decrypt_pad,
		\key1[44]_pad ,
		\roundSel[4]_pad ,
		\roundSel[5]_pad ,
		_w366_
	);
	LUT4 #(
		.INIT('h5554)
	) name62 (
		_w313_,
		_w365_,
		_w366_,
		_w364_,
		_w367_
	);
	LUT4 #(
		.INIT('h0408)
	) name63 (
		decrypt_pad,
		\key3[50]_pad ,
		\roundSel[4]_pad ,
		\roundSel[5]_pad ,
		_w368_
	);
	LUT3 #(
		.INIT('h08)
	) name64 (
		\key2[50]_pad ,
		\roundSel[4]_pad ,
		\roundSel[5]_pad ,
		_w369_
	);
	LUT4 #(
		.INIT('h0804)
	) name65 (
		decrypt_pad,
		\key1[50]_pad ,
		\roundSel[4]_pad ,
		\roundSel[5]_pad ,
		_w370_
	);
	LUT4 #(
		.INIT('haaa8)
	) name66 (
		_w313_,
		_w369_,
		_w370_,
		_w368_,
		_w371_
	);
	LUT3 #(
		.INIT('ha8)
	) name67 (
		_w363_,
		_w367_,
		_w371_,
		_w372_
	);
	LUT4 #(
		.INIT('h0800)
	) name68 (
		\roundSel[0]_pad ,
		\roundSel[1]_pad ,
		\roundSel[2]_pad ,
		\roundSel[3]_pad ,
		_w373_
	);
	LUT4 #(
		.INIT('haaa8)
	) name69 (
		_w313_,
		_w349_,
		_w350_,
		_w348_,
		_w374_
	);
	LUT4 #(
		.INIT('h5554)
	) name70 (
		_w313_,
		_w345_,
		_w346_,
		_w344_,
		_w375_
	);
	LUT3 #(
		.INIT('ha8)
	) name71 (
		_w373_,
		_w374_,
		_w375_,
		_w376_
	);
	LUT4 #(
		.INIT('h0080)
	) name72 (
		\roundSel[0]_pad ,
		\roundSel[1]_pad ,
		\roundSel[2]_pad ,
		\roundSel[3]_pad ,
		_w377_
	);
	LUT4 #(
		.INIT('h0408)
	) name73 (
		decrypt_pad,
		\key3[35]_pad ,
		\roundSel[4]_pad ,
		\roundSel[5]_pad ,
		_w378_
	);
	LUT3 #(
		.INIT('h08)
	) name74 (
		\key2[35]_pad ,
		\roundSel[4]_pad ,
		\roundSel[5]_pad ,
		_w379_
	);
	LUT4 #(
		.INIT('h0804)
	) name75 (
		decrypt_pad,
		\key1[35]_pad ,
		\roundSel[4]_pad ,
		\roundSel[5]_pad ,
		_w380_
	);
	LUT4 #(
		.INIT('h5554)
	) name76 (
		_w313_,
		_w379_,
		_w380_,
		_w378_,
		_w381_
	);
	LUT4 #(
		.INIT('h0408)
	) name77 (
		decrypt_pad,
		\key3[28]_pad ,
		\roundSel[4]_pad ,
		\roundSel[5]_pad ,
		_w382_
	);
	LUT3 #(
		.INIT('h08)
	) name78 (
		\key2[28]_pad ,
		\roundSel[4]_pad ,
		\roundSel[5]_pad ,
		_w383_
	);
	LUT4 #(
		.INIT('h0804)
	) name79 (
		decrypt_pad,
		\key1[28]_pad ,
		\roundSel[4]_pad ,
		\roundSel[5]_pad ,
		_w384_
	);
	LUT4 #(
		.INIT('haaa8)
	) name80 (
		_w313_,
		_w383_,
		_w384_,
		_w382_,
		_w385_
	);
	LUT3 #(
		.INIT('ha8)
	) name81 (
		_w377_,
		_w381_,
		_w385_,
		_w386_
	);
	LUT4 #(
		.INIT('h0001)
	) name82 (
		_w362_,
		_w372_,
		_w376_,
		_w386_,
		_w387_
	);
	LUT4 #(
		.INIT('h1000)
	) name83 (
		\roundSel[0]_pad ,
		\roundSel[1]_pad ,
		\roundSel[2]_pad ,
		\roundSel[3]_pad ,
		_w388_
	);
	LUT4 #(
		.INIT('h0408)
	) name84 (
		decrypt_pad,
		\key3[36]_pad ,
		\roundSel[4]_pad ,
		\roundSel[5]_pad ,
		_w389_
	);
	LUT3 #(
		.INIT('h08)
	) name85 (
		\key2[36]_pad ,
		\roundSel[4]_pad ,
		\roundSel[5]_pad ,
		_w390_
	);
	LUT4 #(
		.INIT('h0804)
	) name86 (
		decrypt_pad,
		\key1[36]_pad ,
		\roundSel[4]_pad ,
		\roundSel[5]_pad ,
		_w391_
	);
	LUT4 #(
		.INIT('haaa8)
	) name87 (
		_w313_,
		_w390_,
		_w391_,
		_w389_,
		_w392_
	);
	LUT4 #(
		.INIT('h0408)
	) name88 (
		decrypt_pad,
		\key3[31]_pad ,
		\roundSel[4]_pad ,
		\roundSel[5]_pad ,
		_w393_
	);
	LUT3 #(
		.INIT('h08)
	) name89 (
		\key2[31]_pad ,
		\roundSel[4]_pad ,
		\roundSel[5]_pad ,
		_w394_
	);
	LUT4 #(
		.INIT('h0804)
	) name90 (
		decrypt_pad,
		\key1[31]_pad ,
		\roundSel[4]_pad ,
		\roundSel[5]_pad ,
		_w395_
	);
	LUT4 #(
		.INIT('h5554)
	) name91 (
		_w313_,
		_w394_,
		_w395_,
		_w393_,
		_w396_
	);
	LUT3 #(
		.INIT('ha8)
	) name92 (
		_w388_,
		_w392_,
		_w396_,
		_w397_
	);
	LUT4 #(
		.INIT('h4000)
	) name93 (
		\roundSel[0]_pad ,
		\roundSel[1]_pad ,
		\roundSel[2]_pad ,
		\roundSel[3]_pad ,
		_w398_
	);
	LUT4 #(
		.INIT('h5554)
	) name94 (
		_w313_,
		_w315_,
		_w316_,
		_w314_,
		_w399_
	);
	LUT4 #(
		.INIT('haaa8)
	) name95 (
		_w313_,
		_w319_,
		_w320_,
		_w318_,
		_w400_
	);
	LUT3 #(
		.INIT('ha8)
	) name96 (
		_w398_,
		_w399_,
		_w400_,
		_w401_
	);
	LUT4 #(
		.INIT('h8000)
	) name97 (
		\roundSel[0]_pad ,
		\roundSel[1]_pad ,
		\roundSel[2]_pad ,
		\roundSel[3]_pad ,
		_w402_
	);
	LUT4 #(
		.INIT('haaa8)
	) name98 (
		_w313_,
		_w355_,
		_w356_,
		_w354_,
		_w403_
	);
	LUT4 #(
		.INIT('h5554)
	) name99 (
		_w313_,
		_w359_,
		_w360_,
		_w358_,
		_w404_
	);
	LUT3 #(
		.INIT('ha8)
	) name100 (
		_w402_,
		_w403_,
		_w404_,
		_w405_
	);
	LUT4 #(
		.INIT('h0008)
	) name101 (
		\roundSel[0]_pad ,
		\roundSel[1]_pad ,
		\roundSel[2]_pad ,
		\roundSel[3]_pad ,
		_w406_
	);
	LUT4 #(
		.INIT('haaa8)
	) name102 (
		_w313_,
		_w394_,
		_w395_,
		_w393_,
		_w407_
	);
	LUT4 #(
		.INIT('h5554)
	) name103 (
		_w313_,
		_w390_,
		_w391_,
		_w389_,
		_w408_
	);
	LUT3 #(
		.INIT('ha8)
	) name104 (
		_w406_,
		_w407_,
		_w408_,
		_w409_
	);
	LUT4 #(
		.INIT('h0001)
	) name105 (
		_w397_,
		_w401_,
		_w405_,
		_w409_,
		_w410_
	);
	LUT4 #(
		.INIT('h0200)
	) name106 (
		\roundSel[0]_pad ,
		\roundSel[1]_pad ,
		\roundSel[2]_pad ,
		\roundSel[3]_pad ,
		_w411_
	);
	LUT4 #(
		.INIT('haaa8)
	) name107 (
		_w313_,
		_w325_,
		_w326_,
		_w324_,
		_w412_
	);
	LUT4 #(
		.INIT('h5554)
	) name108 (
		_w313_,
		_w329_,
		_w330_,
		_w328_,
		_w413_
	);
	LUT3 #(
		.INIT('ha8)
	) name109 (
		_w411_,
		_w412_,
		_w413_,
		_w414_
	);
	LUT4 #(
		.INIT('h0004)
	) name110 (
		\roundSel[0]_pad ,
		\roundSel[1]_pad ,
		\roundSel[2]_pad ,
		\roundSel[3]_pad ,
		_w415_
	);
	LUT4 #(
		.INIT('haaa8)
	) name111 (
		_w313_,
		_w365_,
		_w366_,
		_w364_,
		_w416_
	);
	LUT4 #(
		.INIT('h5554)
	) name112 (
		_w313_,
		_w369_,
		_w370_,
		_w368_,
		_w417_
	);
	LUT3 #(
		.INIT('ha8)
	) name113 (
		_w415_,
		_w416_,
		_w417_,
		_w418_
	);
	LUT4 #(
		.INIT('h0100)
	) name114 (
		\roundSel[0]_pad ,
		\roundSel[1]_pad ,
		\roundSel[2]_pad ,
		\roundSel[3]_pad ,
		_w419_
	);
	LUT4 #(
		.INIT('haaa8)
	) name115 (
		_w313_,
		_w379_,
		_w380_,
		_w378_,
		_w420_
	);
	LUT4 #(
		.INIT('h5554)
	) name116 (
		_w313_,
		_w383_,
		_w384_,
		_w382_,
		_w421_
	);
	LUT3 #(
		.INIT('ha8)
	) name117 (
		_w419_,
		_w420_,
		_w421_,
		_w422_
	);
	LUT4 #(
		.INIT('h0400)
	) name118 (
		\roundSel[0]_pad ,
		\roundSel[1]_pad ,
		\roundSel[2]_pad ,
		\roundSel[3]_pad ,
		_w423_
	);
	LUT4 #(
		.INIT('haaa8)
	) name119 (
		_w313_,
		_w335_,
		_w336_,
		_w334_,
		_w424_
	);
	LUT4 #(
		.INIT('h5554)
	) name120 (
		_w313_,
		_w339_,
		_w340_,
		_w338_,
		_w425_
	);
	LUT3 #(
		.INIT('ha8)
	) name121 (
		_w423_,
		_w424_,
		_w425_,
		_w426_
	);
	LUT4 #(
		.INIT('h0001)
	) name122 (
		_w414_,
		_w418_,
		_w422_,
		_w426_,
		_w427_
	);
	LUT4 #(
		.INIT('h8000)
	) name123 (
		_w410_,
		_w427_,
		_w353_,
		_w387_,
		_w428_
	);
	LUT2 #(
		.INIT('h9)
	) name124 (
		_w310_,
		_w428_,
		_w429_
	);
	LUT4 #(
		.INIT('h0408)
	) name125 (
		decrypt_pad,
		\key3[51]_pad ,
		\roundSel[4]_pad ,
		\roundSel[5]_pad ,
		_w430_
	);
	LUT3 #(
		.INIT('h08)
	) name126 (
		\key2[51]_pad ,
		\roundSel[4]_pad ,
		\roundSel[5]_pad ,
		_w431_
	);
	LUT4 #(
		.INIT('h0804)
	) name127 (
		decrypt_pad,
		\key1[51]_pad ,
		\roundSel[4]_pad ,
		\roundSel[5]_pad ,
		_w432_
	);
	LUT4 #(
		.INIT('haaa8)
	) name128 (
		_w313_,
		_w431_,
		_w432_,
		_w430_,
		_w433_
	);
	LUT3 #(
		.INIT('hc8)
	) name129 (
		_w396_,
		_w402_,
		_w433_,
		_w434_
	);
	LUT4 #(
		.INIT('h5554)
	) name130 (
		_w313_,
		_w431_,
		_w432_,
		_w430_,
		_w435_
	);
	LUT3 #(
		.INIT('ha8)
	) name131 (
		_w305_,
		_w407_,
		_w435_,
		_w436_
	);
	LUT4 #(
		.INIT('h0408)
	) name132 (
		decrypt_pad,
		\key3[21]_pad ,
		\roundSel[4]_pad ,
		\roundSel[5]_pad ,
		_w437_
	);
	LUT3 #(
		.INIT('h08)
	) name133 (
		\key2[21]_pad ,
		\roundSel[4]_pad ,
		\roundSel[5]_pad ,
		_w438_
	);
	LUT4 #(
		.INIT('h0804)
	) name134 (
		decrypt_pad,
		\key1[21]_pad ,
		\roundSel[4]_pad ,
		\roundSel[5]_pad ,
		_w439_
	);
	LUT4 #(
		.INIT('haaa8)
	) name135 (
		_w313_,
		_w438_,
		_w439_,
		_w437_,
		_w440_
	);
	LUT4 #(
		.INIT('h0408)
	) name136 (
		decrypt_pad,
		\key3[2]_pad ,
		\roundSel[4]_pad ,
		\roundSel[5]_pad ,
		_w441_
	);
	LUT3 #(
		.INIT('h08)
	) name137 (
		\key2[2]_pad ,
		\roundSel[4]_pad ,
		\roundSel[5]_pad ,
		_w442_
	);
	LUT4 #(
		.INIT('h0804)
	) name138 (
		decrypt_pad,
		\key1[2]_pad ,
		\roundSel[4]_pad ,
		\roundSel[5]_pad ,
		_w443_
	);
	LUT4 #(
		.INIT('h5554)
	) name139 (
		_w313_,
		_w442_,
		_w443_,
		_w441_,
		_w444_
	);
	LUT3 #(
		.INIT('ha8)
	) name140 (
		_w343_,
		_w440_,
		_w444_,
		_w445_
	);
	LUT4 #(
		.INIT('h0408)
	) name141 (
		decrypt_pad,
		\key3[15]_pad ,
		\roundSel[4]_pad ,
		\roundSel[5]_pad ,
		_w446_
	);
	LUT3 #(
		.INIT('h08)
	) name142 (
		\key2[15]_pad ,
		\roundSel[4]_pad ,
		\roundSel[5]_pad ,
		_w447_
	);
	LUT4 #(
		.INIT('h0804)
	) name143 (
		decrypt_pad,
		\key1[15]_pad ,
		\roundSel[4]_pad ,
		\roundSel[5]_pad ,
		_w448_
	);
	LUT4 #(
		.INIT('h5554)
	) name144 (
		_w313_,
		_w447_,
		_w448_,
		_w446_,
		_w449_
	);
	LUT3 #(
		.INIT('ha8)
	) name145 (
		_w377_,
		_w424_,
		_w449_,
		_w450_
	);
	LUT4 #(
		.INIT('h0001)
	) name146 (
		_w434_,
		_w436_,
		_w445_,
		_w450_,
		_w451_
	);
	LUT4 #(
		.INIT('h0408)
	) name147 (
		decrypt_pad,
		\key3[29]_pad ,
		\roundSel[4]_pad ,
		\roundSel[5]_pad ,
		_w452_
	);
	LUT3 #(
		.INIT('h08)
	) name148 (
		\key2[29]_pad ,
		\roundSel[4]_pad ,
		\roundSel[5]_pad ,
		_w453_
	);
	LUT4 #(
		.INIT('h0804)
	) name149 (
		decrypt_pad,
		\key1[29]_pad ,
		\roundSel[4]_pad ,
		\roundSel[5]_pad ,
		_w454_
	);
	LUT4 #(
		.INIT('h5554)
	) name150 (
		_w313_,
		_w453_,
		_w454_,
		_w452_,
		_w455_
	);
	LUT3 #(
		.INIT('ha8)
	) name151 (
		_w323_,
		_w412_,
		_w455_,
		_w456_
	);
	LUT4 #(
		.INIT('haaa8)
	) name152 (
		_w313_,
		_w453_,
		_w454_,
		_w452_,
		_w457_
	);
	LUT3 #(
		.INIT('hc8)
	) name153 (
		_w327_,
		_w411_,
		_w457_,
		_w458_
	);
	LUT4 #(
		.INIT('haaa8)
	) name154 (
		_w313_,
		_w442_,
		_w443_,
		_w441_,
		_w459_
	);
	LUT4 #(
		.INIT('h5554)
	) name155 (
		_w313_,
		_w438_,
		_w439_,
		_w437_,
		_w460_
	);
	LUT3 #(
		.INIT('ha8)
	) name156 (
		_w373_,
		_w459_,
		_w460_,
		_w461_
	);
	LUT4 #(
		.INIT('h0408)
	) name157 (
		decrypt_pad,
		\key3[7]_pad ,
		\roundSel[4]_pad ,
		\roundSel[5]_pad ,
		_w462_
	);
	LUT3 #(
		.INIT('h08)
	) name158 (
		\key2[7]_pad ,
		\roundSel[4]_pad ,
		\roundSel[5]_pad ,
		_w463_
	);
	LUT4 #(
		.INIT('h0804)
	) name159 (
		decrypt_pad,
		\key1[7]_pad ,
		\roundSel[4]_pad ,
		\roundSel[5]_pad ,
		_w464_
	);
	LUT4 #(
		.INIT('h5554)
	) name160 (
		_w313_,
		_w463_,
		_w464_,
		_w462_,
		_w465_
	);
	LUT3 #(
		.INIT('ha8)
	) name161 (
		_w388_,
		_w403_,
		_w465_,
		_w466_
	);
	LUT4 #(
		.INIT('h0001)
	) name162 (
		_w456_,
		_w458_,
		_w461_,
		_w466_,
		_w467_
	);
	LUT4 #(
		.INIT('h0408)
	) name163 (
		decrypt_pad,
		\key3[38]_pad ,
		\roundSel[4]_pad ,
		\roundSel[5]_pad ,
		_w468_
	);
	LUT3 #(
		.INIT('h08)
	) name164 (
		\key2[38]_pad ,
		\roundSel[4]_pad ,
		\roundSel[5]_pad ,
		_w469_
	);
	LUT4 #(
		.INIT('h0804)
	) name165 (
		decrypt_pad,
		\key1[38]_pad ,
		\roundSel[4]_pad ,
		\roundSel[5]_pad ,
		_w470_
	);
	LUT4 #(
		.INIT('h5554)
	) name166 (
		_w313_,
		_w469_,
		_w470_,
		_w468_,
		_w471_
	);
	LUT3 #(
		.INIT('hc8)
	) name167 (
		_w416_,
		_w398_,
		_w471_,
		_w472_
	);
	LUT4 #(
		.INIT('haaa8)
	) name168 (
		_w313_,
		_w469_,
		_w470_,
		_w468_,
		_w473_
	);
	LUT3 #(
		.INIT('hc8)
	) name169 (
		_w367_,
		_w312_,
		_w473_,
		_w474_
	);
	LUT4 #(
		.INIT('h0408)
	) name170 (
		decrypt_pad,
		\key3[43]_pad ,
		\roundSel[4]_pad ,
		\roundSel[5]_pad ,
		_w475_
	);
	LUT3 #(
		.INIT('h08)
	) name171 (
		\key2[43]_pad ,
		\roundSel[4]_pad ,
		\roundSel[5]_pad ,
		_w476_
	);
	LUT4 #(
		.INIT('h0804)
	) name172 (
		decrypt_pad,
		\key1[43]_pad ,
		\roundSel[4]_pad ,
		\roundSel[5]_pad ,
		_w477_
	);
	LUT4 #(
		.INIT('h5554)
	) name173 (
		_w313_,
		_w476_,
		_w477_,
		_w475_,
		_w478_
	);
	LUT3 #(
		.INIT('ha8)
	) name174 (
		_w333_,
		_w420_,
		_w478_,
		_w479_
	);
	LUT4 #(
		.INIT('haaa8)
	) name175 (
		_w313_,
		_w447_,
		_w448_,
		_w446_,
		_w480_
	);
	LUT3 #(
		.INIT('hc8)
	) name176 (
		_w337_,
		_w419_,
		_w480_,
		_w481_
	);
	LUT4 #(
		.INIT('h0001)
	) name177 (
		_w472_,
		_w474_,
		_w479_,
		_w481_,
		_w482_
	);
	LUT4 #(
		.INIT('haaa8)
	) name178 (
		_w313_,
		_w463_,
		_w464_,
		_w462_,
		_w483_
	);
	LUT3 #(
		.INIT('hc8)
	) name179 (
		_w357_,
		_w406_,
		_w483_,
		_w484_
	);
	LUT4 #(
		.INIT('h0408)
	) name180 (
		decrypt_pad,
		\key3[52]_pad ,
		\roundSel[4]_pad ,
		\roundSel[5]_pad ,
		_w485_
	);
	LUT3 #(
		.INIT('h08)
	) name181 (
		\key2[52]_pad ,
		\roundSel[4]_pad ,
		\roundSel[5]_pad ,
		_w486_
	);
	LUT4 #(
		.INIT('h0804)
	) name182 (
		decrypt_pad,
		\key1[52]_pad ,
		\roundSel[4]_pad ,
		\roundSel[5]_pad ,
		_w487_
	);
	LUT4 #(
		.INIT('haaa8)
	) name183 (
		_w313_,
		_w486_,
		_w487_,
		_w485_,
		_w488_
	);
	LUT3 #(
		.INIT('ha8)
	) name184 (
		_w415_,
		_w399_,
		_w488_,
		_w489_
	);
	LUT4 #(
		.INIT('h5554)
	) name185 (
		_w313_,
		_w486_,
		_w487_,
		_w485_,
		_w490_
	);
	LUT3 #(
		.INIT('ha8)
	) name186 (
		_w363_,
		_w317_,
		_w490_,
		_w491_
	);
	LUT4 #(
		.INIT('haaa8)
	) name187 (
		_w313_,
		_w476_,
		_w477_,
		_w475_,
		_w492_
	);
	LUT3 #(
		.INIT('hc8)
	) name188 (
		_w381_,
		_w423_,
		_w492_,
		_w493_
	);
	LUT4 #(
		.INIT('h0001)
	) name189 (
		_w484_,
		_w489_,
		_w491_,
		_w493_,
		_w494_
	);
	LUT4 #(
		.INIT('h8000)
	) name190 (
		_w482_,
		_w494_,
		_w451_,
		_w467_,
		_w495_
	);
	LUT4 #(
		.INIT('h0200)
	) name191 (
		\desIn[3]_pad ,
		\roundSel[4]_pad ,
		\roundSel[5]_pad ,
		_w305_,
		_w496_
	);
	LUT4 #(
		.INIT('h4155)
	) name192 (
		\FP_R_reg[17]/P0001 ,
		\roundSel[4]_pad ,
		\roundSel[5]_pad ,
		_w305_,
		_w497_
	);
	LUT4 #(
		.INIT('he8ff)
	) name193 (
		\FP_R_reg[49]/NET0131 ,
		\roundSel[4]_pad ,
		\roundSel[5]_pad ,
		_w305_,
		_w498_
	);
	LUT3 #(
		.INIT('h45)
	) name194 (
		_w496_,
		_w497_,
		_w498_,
		_w499_
	);
	LUT3 #(
		.INIT('hba)
	) name195 (
		_w496_,
		_w497_,
		_w498_,
		_w500_
	);
	LUT2 #(
		.INIT('h9)
	) name196 (
		_w495_,
		_w499_,
		_w501_
	);
	LUT3 #(
		.INIT('hc8)
	) name197 (
		_w337_,
		_w415_,
		_w459_,
		_w502_
	);
	LUT3 #(
		.INIT('hc8)
	) name198 (
		_w375_,
		_w419_,
		_w488_,
		_w503_
	);
	LUT3 #(
		.INIT('ha8)
	) name199 (
		_w312_,
		_w351_,
		_w492_,
		_w504_
	);
	LUT3 #(
		.INIT('ha8)
	) name200 (
		_w373_,
		_w420_,
		_w399_,
		_w505_
	);
	LUT4 #(
		.INIT('h0001)
	) name201 (
		_w502_,
		_w503_,
		_w504_,
		_w505_,
		_w506_
	);
	LUT3 #(
		.INIT('he0)
	) name202 (
		_w357_,
		_w412_,
		_w388_,
		_w507_
	);
	LUT3 #(
		.INIT('ha8)
	) name203 (
		_w377_,
		_w347_,
		_w490_,
		_w508_
	);
	LUT3 #(
		.INIT('hc8)
	) name204 (
		_w374_,
		_w398_,
		_w478_,
		_w509_
	);
	LUT3 #(
		.INIT('ha8)
	) name205 (
		_w323_,
		_w407_,
		_w465_,
		_w510_
	);
	LUT4 #(
		.INIT('h0001)
	) name206 (
		_w507_,
		_w508_,
		_w509_,
		_w510_,
		_w511_
	);
	LUT3 #(
		.INIT('ha8)
	) name207 (
		_w411_,
		_w396_,
		_w483_,
		_w512_
	);
	LUT3 #(
		.INIT('ha8)
	) name208 (
		_w402_,
		_w408_,
		_w457_,
		_w513_
	);
	LUT3 #(
		.INIT('hc8)
	) name209 (
		_w367_,
		_w423_,
		_w440_,
		_w514_
	);
	LUT3 #(
		.INIT('he0)
	) name210 (
		_w381_,
		_w317_,
		_w343_,
		_w515_
	);
	LUT4 #(
		.INIT('h0001)
	) name211 (
		_w512_,
		_w513_,
		_w514_,
		_w515_,
		_w516_
	);
	LUT3 #(
		.INIT('he0)
	) name212 (
		_w327_,
		_w403_,
		_w406_,
		_w517_
	);
	LUT3 #(
		.INIT('ha8)
	) name213 (
		_w305_,
		_w392_,
		_w455_,
		_w518_
	);
	LUT3 #(
		.INIT('ha8)
	) name214 (
		_w363_,
		_w424_,
		_w444_,
		_w519_
	);
	LUT3 #(
		.INIT('ha8)
	) name215 (
		_w333_,
		_w416_,
		_w460_,
		_w520_
	);
	LUT4 #(
		.INIT('h0001)
	) name216 (
		_w517_,
		_w518_,
		_w519_,
		_w520_,
		_w521_
	);
	LUT4 #(
		.INIT('h8000)
	) name217 (
		_w516_,
		_w521_,
		_w506_,
		_w511_,
		_w522_
	);
	LUT4 #(
		.INIT('h0200)
	) name218 (
		\desIn[61]_pad ,
		\roundSel[4]_pad ,
		\roundSel[5]_pad ,
		_w305_,
		_w523_
	);
	LUT4 #(
		.INIT('h4155)
	) name219 (
		\FP_R_reg[16]/P0001 ,
		\roundSel[4]_pad ,
		\roundSel[5]_pad ,
		_w305_,
		_w524_
	);
	LUT4 #(
		.INIT('he8ff)
	) name220 (
		\FP_R_reg[48]/NET0131 ,
		\roundSel[4]_pad ,
		\roundSel[5]_pad ,
		_w305_,
		_w525_
	);
	LUT3 #(
		.INIT('h45)
	) name221 (
		_w523_,
		_w524_,
		_w525_,
		_w526_
	);
	LUT3 #(
		.INIT('hba)
	) name222 (
		_w523_,
		_w524_,
		_w525_,
		_w527_
	);
	LUT2 #(
		.INIT('h9)
	) name223 (
		_w522_,
		_w526_,
		_w528_
	);
	LUT3 #(
		.INIT('ha8)
	) name224 (
		_w363_,
		_w413_,
		_w433_,
		_w529_
	);
	LUT3 #(
		.INIT('ha8)
	) name225 (
		_w305_,
		_w375_,
		_w488_,
		_w530_
	);
	LUT3 #(
		.INIT('ha8)
	) name226 (
		_w323_,
		_w417_,
		_w480_,
		_w531_
	);
	LUT3 #(
		.INIT('hc8)
	) name227 (
		_w371_,
		_w411_,
		_w449_,
		_w532_
	);
	LUT4 #(
		.INIT('h0001)
	) name228 (
		_w529_,
		_w530_,
		_w531_,
		_w532_,
		_w533_
	);
	LUT3 #(
		.INIT('hc8)
	) name229 (
		_w425_,
		_w398_,
		_w473_,
		_w534_
	);
	LUT3 #(
		.INIT('ha8)
	) name230 (
		_w419_,
		_w392_,
		_w455_,
		_w535_
	);
	LUT4 #(
		.INIT('h0408)
	) name231 (
		decrypt_pad,
		\key3[42]_pad ,
		\roundSel[4]_pad ,
		\roundSel[5]_pad ,
		_w536_
	);
	LUT3 #(
		.INIT('h08)
	) name232 (
		\key2[42]_pad ,
		\roundSel[4]_pad ,
		\roundSel[5]_pad ,
		_w537_
	);
	LUT4 #(
		.INIT('h0804)
	) name233 (
		decrypt_pad,
		\key1[42]_pad ,
		\roundSel[4]_pad ,
		\roundSel[5]_pad ,
		_w538_
	);
	LUT4 #(
		.INIT('h5554)
	) name234 (
		_w313_,
		_w537_,
		_w538_,
		_w536_,
		_w539_
	);
	LUT3 #(
		.INIT('hc8)
	) name235 (
		_w361_,
		_w373_,
		_w539_,
		_w540_
	);
	LUT3 #(
		.INIT('hc8)
	) name236 (
		_w331_,
		_w415_,
		_w435_,
		_w541_
	);
	LUT4 #(
		.INIT('h0001)
	) name237 (
		_w534_,
		_w535_,
		_w540_,
		_w541_,
		_w542_
	);
	LUT3 #(
		.INIT('ha8)
	) name238 (
		_w312_,
		_w341_,
		_w471_,
		_w543_
	);
	LUT3 #(
		.INIT('ha8)
	) name239 (
		_w377_,
		_w408_,
		_w457_,
		_w544_
	);
	LUT4 #(
		.INIT('h0408)
	) name240 (
		decrypt_pad,
		\key3[37]_pad ,
		\roundSel[4]_pad ,
		\roundSel[5]_pad ,
		_w545_
	);
	LUT3 #(
		.INIT('h08)
	) name241 (
		\key2[37]_pad ,
		\roundSel[4]_pad ,
		\roundSel[5]_pad ,
		_w546_
	);
	LUT4 #(
		.INIT('h0804)
	) name242 (
		decrypt_pad,
		\key1[37]_pad ,
		\roundSel[4]_pad ,
		\roundSel[5]_pad ,
		_w547_
	);
	LUT4 #(
		.INIT('h5554)
	) name243 (
		_w313_,
		_w546_,
		_w547_,
		_w545_,
		_w548_
	);
	LUT3 #(
		.INIT('hc8)
	) name244 (
		_w385_,
		_w406_,
		_w548_,
		_w549_
	);
	LUT4 #(
		.INIT('h0408)
	) name245 (
		decrypt_pad,
		\key3[1]_pad ,
		\roundSel[4]_pad ,
		\roundSel[5]_pad ,
		_w550_
	);
	LUT3 #(
		.INIT('h08)
	) name246 (
		\key2[1]_pad ,
		\roundSel[4]_pad ,
		\roundSel[5]_pad ,
		_w551_
	);
	LUT4 #(
		.INIT('h0804)
	) name247 (
		decrypt_pad,
		\key1[1]_pad ,
		\roundSel[4]_pad ,
		\roundSel[5]_pad ,
		_w552_
	);
	LUT4 #(
		.INIT('haaa8)
	) name248 (
		_w313_,
		_w551_,
		_w552_,
		_w550_,
		_w553_
	);
	LUT3 #(
		.INIT('hc8)
	) name249 (
		_w321_,
		_w333_,
		_w553_,
		_w554_
	);
	LUT4 #(
		.INIT('h0001)
	) name250 (
		_w543_,
		_w544_,
		_w549_,
		_w554_,
		_w555_
	);
	LUT4 #(
		.INIT('haaa8)
	) name251 (
		_w313_,
		_w546_,
		_w547_,
		_w545_,
		_w556_
	);
	LUT3 #(
		.INIT('hc8)
	) name252 (
		_w421_,
		_w388_,
		_w556_,
		_w557_
	);
	LUT3 #(
		.INIT('hc8)
	) name253 (
		_w347_,
		_w402_,
		_w490_,
		_w558_
	);
	LUT4 #(
		.INIT('haaa8)
	) name254 (
		_w313_,
		_w537_,
		_w538_,
		_w536_,
		_w559_
	);
	LUT3 #(
		.INIT('ha8)
	) name255 (
		_w343_,
		_w404_,
		_w559_,
		_w560_
	);
	LUT4 #(
		.INIT('h5554)
	) name256 (
		_w313_,
		_w551_,
		_w552_,
		_w550_,
		_w561_
	);
	LUT3 #(
		.INIT('ha8)
	) name257 (
		_w423_,
		_w400_,
		_w561_,
		_w562_
	);
	LUT4 #(
		.INIT('h0001)
	) name258 (
		_w557_,
		_w558_,
		_w560_,
		_w562_,
		_w563_
	);
	LUT4 #(
		.INIT('h8000)
	) name259 (
		_w555_,
		_w563_,
		_w533_,
		_w542_,
		_w564_
	);
	LUT4 #(
		.INIT('h0200)
	) name260 (
		\desIn[35]_pad ,
		\roundSel[4]_pad ,
		\roundSel[5]_pad ,
		_w305_,
		_w565_
	);
	LUT4 #(
		.INIT('h4155)
	) name261 (
		\FP_R_reg[21]/P0001 ,
		\roundSel[4]_pad ,
		\roundSel[5]_pad ,
		_w305_,
		_w566_
	);
	LUT4 #(
		.INIT('he8ff)
	) name262 (
		\FP_R_reg[53]/NET0131 ,
		\roundSel[4]_pad ,
		\roundSel[5]_pad ,
		_w305_,
		_w567_
	);
	LUT3 #(
		.INIT('h45)
	) name263 (
		_w565_,
		_w566_,
		_w567_,
		_w568_
	);
	LUT3 #(
		.INIT('hba)
	) name264 (
		_w565_,
		_w566_,
		_w567_,
		_w569_
	);
	LUT2 #(
		.INIT('h9)
	) name265 (
		_w564_,
		_w568_,
		_w570_
	);
	LUT4 #(
		.INIT('h9009)
	) name266 (
		_w522_,
		_w526_,
		_w564_,
		_w568_,
		_w571_
	);
	LUT3 #(
		.INIT('ha8)
	) name267 (
		_w343_,
		_w459_,
		_w465_,
		_w572_
	);
	LUT3 #(
		.INIT('hc8)
	) name268 (
		_w367_,
		_w419_,
		_w433_,
		_w573_
	);
	LUT3 #(
		.INIT('hc8)
	) name269 (
		_w337_,
		_w402_,
		_w553_,
		_w574_
	);
	LUT3 #(
		.INIT('ha8)
	) name270 (
		_w312_,
		_w327_,
		_w480_,
		_w575_
	);
	LUT4 #(
		.INIT('h0001)
	) name271 (
		_w572_,
		_w573_,
		_w574_,
		_w575_,
		_w576_
	);
	LUT3 #(
		.INIT('ha8)
	) name272 (
		_w388_,
		_w440_,
		_w478_,
		_w577_
	);
	LUT3 #(
		.INIT('ha8)
	) name273 (
		_w305_,
		_w424_,
		_w561_,
		_w578_
	);
	LUT3 #(
		.INIT('hc8)
	) name274 (
		_w381_,
		_w415_,
		_w457_,
		_w579_
	);
	LUT3 #(
		.INIT('hc8)
	) name275 (
		_w317_,
		_w323_,
		_w471_,
		_w580_
	);
	LUT4 #(
		.INIT('h0001)
	) name276 (
		_w577_,
		_w578_,
		_w579_,
		_w580_,
		_w581_
	);
	LUT3 #(
		.INIT('hc8)
	) name277 (
		_w357_,
		_w423_,
		_w488_,
		_w582_
	);
	LUT3 #(
		.INIT('ha8)
	) name278 (
		_w377_,
		_w416_,
		_w435_,
		_w583_
	);
	LUT3 #(
		.INIT('ha8)
	) name279 (
		_w363_,
		_w420_,
		_w455_,
		_w584_
	);
	LUT3 #(
		.INIT('ha8)
	) name280 (
		_w406_,
		_w460_,
		_w492_,
		_w585_
	);
	LUT4 #(
		.INIT('h0001)
	) name281 (
		_w582_,
		_w583_,
		_w584_,
		_w585_,
		_w586_
	);
	LUT3 #(
		.INIT('ha8)
	) name282 (
		_w411_,
		_w399_,
		_w473_,
		_w587_
	);
	LUT3 #(
		.INIT('hc8)
	) name283 (
		_w412_,
		_w398_,
		_w449_,
		_w588_
	);
	LUT3 #(
		.INIT('ha8)
	) name284 (
		_w333_,
		_w403_,
		_w490_,
		_w589_
	);
	LUT3 #(
		.INIT('ha8)
	) name285 (
		_w373_,
		_w444_,
		_w483_,
		_w590_
	);
	LUT4 #(
		.INIT('h0001)
	) name286 (
		_w587_,
		_w588_,
		_w589_,
		_w590_,
		_w591_
	);
	LUT4 #(
		.INIT('h8000)
	) name287 (
		_w586_,
		_w591_,
		_w576_,
		_w581_,
		_w592_
	);
	LUT4 #(
		.INIT('h0100)
	) name288 (
		\desIn[19]_pad ,
		\roundSel[4]_pad ,
		\roundSel[5]_pad ,
		_w305_,
		_w593_
	);
	LUT4 #(
		.INIT('h2800)
	) name289 (
		\FP_R_reg[51]/NET0131 ,
		\roundSel[4]_pad ,
		\roundSel[5]_pad ,
		_w305_,
		_w594_
	);
	LUT4 #(
		.INIT('h7c55)
	) name290 (
		\FP_R_reg[19]/P0001 ,
		\roundSel[4]_pad ,
		\roundSel[5]_pad ,
		_w305_,
		_w595_
	);
	LUT3 #(
		.INIT('h45)
	) name291 (
		_w593_,
		_w594_,
		_w595_,
		_w596_
	);
	LUT2 #(
		.INIT('h9)
	) name292 (
		_w592_,
		_w596_,
		_w597_
	);
	LUT4 #(
		.INIT('h0660)
	) name293 (
		_w495_,
		_w499_,
		_w522_,
		_w526_,
		_w598_
	);
	LUT4 #(
		.INIT('h006e)
	) name294 (
		_w501_,
		_w528_,
		_w570_,
		_w597_,
		_w599_
	);
	LUT3 #(
		.INIT('hc8)
	) name295 (
		_w361_,
		_w411_,
		_w478_,
		_w600_
	);
	LUT3 #(
		.INIT('hc8)
	) name296 (
		_w331_,
		_w402_,
		_w460_,
		_w601_
	);
	LUT3 #(
		.INIT('ha8)
	) name297 (
		_w305_,
		_w413_,
		_w440_,
		_w602_
	);
	LUT3 #(
		.INIT('ha8)
	) name298 (
		_w323_,
		_w404_,
		_w492_,
		_w603_
	);
	LUT4 #(
		.INIT('h0001)
	) name299 (
		_w600_,
		_w601_,
		_w602_,
		_w603_,
		_w604_
	);
	LUT3 #(
		.INIT('ha8)
	) name300 (
		_w333_,
		_w457_,
		_w548_,
		_w605_
	);
	LUT3 #(
		.INIT('ha8)
	) name301 (
		_w419_,
		_w400_,
		_w444_,
		_w606_
	);
	LUT3 #(
		.INIT('ha8)
	) name302 (
		_w388_,
		_w473_,
		_w561_,
		_w607_
	);
	LUT3 #(
		.INIT('hc8)
	) name303 (
		_w421_,
		_w398_,
		_w483_,
		_w608_
	);
	LUT4 #(
		.INIT('h0001)
	) name304 (
		_w605_,
		_w606_,
		_w607_,
		_w608_,
		_w609_
	);
	LUT3 #(
		.INIT('ha8)
	) name305 (
		_w423_,
		_w455_,
		_w556_,
		_w610_
	);
	LUT3 #(
		.INIT('ha8)
	) name306 (
		_w377_,
		_w321_,
		_w459_,
		_w611_
	);
	LUT3 #(
		.INIT('ha8)
	) name307 (
		_w406_,
		_w471_,
		_w553_,
		_w612_
	);
	LUT3 #(
		.INIT('ha8)
	) name308 (
		_w373_,
		_w433_,
		_w449_,
		_w613_
	);
	LUT4 #(
		.INIT('h0001)
	) name309 (
		_w610_,
		_w611_,
		_w612_,
		_w613_,
		_w614_
	);
	LUT3 #(
		.INIT('ha8)
	) name310 (
		_w415_,
		_w490_,
		_w559_,
		_w615_
	);
	LUT3 #(
		.INIT('hc8)
	) name311 (
		_w385_,
		_w312_,
		_w465_,
		_w616_
	);
	LUT3 #(
		.INIT('ha8)
	) name312 (
		_w363_,
		_w488_,
		_w539_,
		_w617_
	);
	LUT3 #(
		.INIT('ha8)
	) name313 (
		_w343_,
		_w435_,
		_w480_,
		_w618_
	);
	LUT4 #(
		.INIT('h0001)
	) name314 (
		_w615_,
		_w616_,
		_w617_,
		_w618_,
		_w619_
	);
	LUT4 #(
		.INIT('h8000)
	) name315 (
		_w614_,
		_w619_,
		_w604_,
		_w609_,
		_w620_
	);
	LUT4 #(
		.INIT('h0200)
	) name316 (
		\desIn[11]_pad ,
		\roundSel[4]_pad ,
		\roundSel[5]_pad ,
		_w305_,
		_w621_
	);
	LUT4 #(
		.INIT('h4155)
	) name317 (
		\FP_R_reg[18]/P0001 ,
		\roundSel[4]_pad ,
		\roundSel[5]_pad ,
		_w305_,
		_w622_
	);
	LUT4 #(
		.INIT('he8ff)
	) name318 (
		\FP_R_reg[50]/NET0131 ,
		\roundSel[4]_pad ,
		\roundSel[5]_pad ,
		_w305_,
		_w623_
	);
	LUT3 #(
		.INIT('h45)
	) name319 (
		_w621_,
		_w622_,
		_w623_,
		_w624_
	);
	LUT3 #(
		.INIT('hba)
	) name320 (
		_w621_,
		_w622_,
		_w623_,
		_w625_
	);
	LUT2 #(
		.INIT('h9)
	) name321 (
		_w620_,
		_w624_,
		_w626_
	);
	LUT4 #(
		.INIT('h0660)
	) name322 (
		_w522_,
		_w526_,
		_w564_,
		_w568_,
		_w627_
	);
	LUT4 #(
		.INIT('h0660)
	) name323 (
		_w495_,
		_w499_,
		_w564_,
		_w568_,
		_w628_
	);
	LUT3 #(
		.INIT('h27)
	) name324 (
		_w626_,
		_w627_,
		_w628_,
		_w629_
	);
	LUT2 #(
		.INIT('h4)
	) name325 (
		_w501_,
		_w571_,
		_w630_
	);
	LUT4 #(
		.INIT('h0990)
	) name326 (
		_w495_,
		_w499_,
		_w620_,
		_w624_,
		_w631_
	);
	LUT2 #(
		.INIT('h4)
	) name327 (
		_w528_,
		_w631_,
		_w632_
	);
	LUT3 #(
		.INIT('h8c)
	) name328 (
		_w528_,
		_w597_,
		_w631_,
		_w633_
	);
	LUT4 #(
		.INIT('h7077)
	) name329 (
		_w599_,
		_w629_,
		_w630_,
		_w633_,
		_w634_
	);
	LUT4 #(
		.INIT('h0990)
	) name330 (
		_w522_,
		_w526_,
		_w564_,
		_w568_,
		_w635_
	);
	LUT4 #(
		.INIT('hf75f)
	) name331 (
		_w501_,
		_w528_,
		_w570_,
		_w626_,
		_w636_
	);
	LUT3 #(
		.INIT('h8a)
	) name332 (
		_w429_,
		_w634_,
		_w636_,
		_w637_
	);
	LUT3 #(
		.INIT('h40)
	) name333 (
		_w501_,
		_w626_,
		_w627_,
		_w638_
	);
	LUT4 #(
		.INIT('hf6ff)
	) name334 (
		_w501_,
		_w528_,
		_w570_,
		_w626_,
		_w639_
	);
	LUT4 #(
		.INIT('hf6ef)
	) name335 (
		_w501_,
		_w528_,
		_w570_,
		_w626_,
		_w640_
	);
	LUT2 #(
		.INIT('h1)
	) name336 (
		_w597_,
		_w640_,
		_w641_
	);
	LUT2 #(
		.INIT('h2)
	) name337 (
		_w528_,
		_w628_,
		_w642_
	);
	LUT4 #(
		.INIT('h0004)
	) name338 (
		_w429_,
		_w597_,
		_w598_,
		_w631_,
		_w643_
	);
	LUT2 #(
		.INIT('h4)
	) name339 (
		_w642_,
		_w643_,
		_w644_
	);
	LUT4 #(
		.INIT('h0990)
	) name340 (
		_w495_,
		_w499_,
		_w564_,
		_w568_,
		_w645_
	);
	LUT4 #(
		.INIT('h0660)
	) name341 (
		_w310_,
		_w428_,
		_w620_,
		_w624_,
		_w646_
	);
	LUT4 #(
		.INIT('hd800)
	) name342 (
		_w597_,
		_w598_,
		_w645_,
		_w646_,
		_w647_
	);
	LUT4 #(
		.INIT('h6006)
	) name343 (
		_w522_,
		_w526_,
		_w564_,
		_w568_,
		_w648_
	);
	LUT2 #(
		.INIT('h8)
	) name344 (
		_w501_,
		_w648_,
		_w649_
	);
	LUT4 #(
		.INIT('h6006)
	) name345 (
		_w310_,
		_w428_,
		_w620_,
		_w624_,
		_w650_
	);
	LUT3 #(
		.INIT('h80)
	) name346 (
		_w501_,
		_w648_,
		_w650_,
		_w651_
	);
	LUT4 #(
		.INIT('h6006)
	) name347 (
		_w495_,
		_w499_,
		_w620_,
		_w624_,
		_w652_
	);
	LUT4 #(
		.INIT('h9009)
	) name348 (
		_w522_,
		_w526_,
		_w592_,
		_w596_,
		_w653_
	);
	LUT4 #(
		.INIT('ha7f7)
	) name349 (
		_w501_,
		_w571_,
		_w626_,
		_w653_,
		_w654_
	);
	LUT3 #(
		.INIT('h10)
	) name350 (
		_w651_,
		_w647_,
		_w654_,
		_w655_
	);
	LUT3 #(
		.INIT('h10)
	) name351 (
		_w641_,
		_w644_,
		_w655_,
		_w656_
	);
	LUT4 #(
		.INIT('h0100)
	) name352 (
		\desIn[0]_pad ,
		\roundSel[4]_pad ,
		\roundSel[5]_pad ,
		_w305_,
		_w657_
	);
	LUT4 #(
		.INIT('h2800)
	) name353 (
		\FP_R_reg[25]/P0001 ,
		\roundSel[4]_pad ,
		\roundSel[5]_pad ,
		_w305_,
		_w658_
	);
	LUT4 #(
		.INIT('h7c55)
	) name354 (
		\FP_R_reg[57]/NET0131 ,
		\roundSel[4]_pad ,
		\roundSel[5]_pad ,
		_w305_,
		_w659_
	);
	LUT3 #(
		.INIT('h45)
	) name355 (
		_w657_,
		_w658_,
		_w659_,
		_w660_
	);
	LUT3 #(
		.INIT('h4b)
	) name356 (
		_w637_,
		_w656_,
		_w660_,
		_w661_
	);
	LUT4 #(
		.INIT('h0408)
	) name357 (
		decrypt_pad,
		\key3[4]_pad ,
		\roundSel[4]_pad ,
		\roundSel[5]_pad ,
		_w662_
	);
	LUT3 #(
		.INIT('h08)
	) name358 (
		\key2[4]_pad ,
		\roundSel[4]_pad ,
		\roundSel[5]_pad ,
		_w663_
	);
	LUT4 #(
		.INIT('h0804)
	) name359 (
		decrypt_pad,
		\key1[4]_pad ,
		\roundSel[4]_pad ,
		\roundSel[5]_pad ,
		_w664_
	);
	LUT4 #(
		.INIT('haaa8)
	) name360 (
		_w313_,
		_w663_,
		_w664_,
		_w662_,
		_w665_
	);
	LUT4 #(
		.INIT('h0408)
	) name361 (
		decrypt_pad,
		\key3[12]_pad ,
		\roundSel[4]_pad ,
		\roundSel[5]_pad ,
		_w666_
	);
	LUT3 #(
		.INIT('h08)
	) name362 (
		\key2[12]_pad ,
		\roundSel[4]_pad ,
		\roundSel[5]_pad ,
		_w667_
	);
	LUT4 #(
		.INIT('h0804)
	) name363 (
		decrypt_pad,
		\key1[12]_pad ,
		\roundSel[4]_pad ,
		\roundSel[5]_pad ,
		_w668_
	);
	LUT4 #(
		.INIT('h5554)
	) name364 (
		_w313_,
		_w667_,
		_w668_,
		_w666_,
		_w669_
	);
	LUT3 #(
		.INIT('ha8)
	) name365 (
		_w415_,
		_w665_,
		_w669_,
		_w670_
	);
	LUT4 #(
		.INIT('h5554)
	) name366 (
		_w313_,
		_w663_,
		_w664_,
		_w662_,
		_w671_
	);
	LUT4 #(
		.INIT('haaa8)
	) name367 (
		_w313_,
		_w667_,
		_w668_,
		_w666_,
		_w672_
	);
	LUT3 #(
		.INIT('ha8)
	) name368 (
		_w363_,
		_w671_,
		_w672_,
		_w673_
	);
	LUT4 #(
		.INIT('h0408)
	) name369 (
		decrypt_pad,
		\key3[27]_pad ,
		\roundSel[4]_pad ,
		\roundSel[5]_pad ,
		_w674_
	);
	LUT3 #(
		.INIT('h08)
	) name370 (
		\key2[27]_pad ,
		\roundSel[4]_pad ,
		\roundSel[5]_pad ,
		_w675_
	);
	LUT4 #(
		.INIT('h0804)
	) name371 (
		decrypt_pad,
		\key1[27]_pad ,
		\roundSel[4]_pad ,
		\roundSel[5]_pad ,
		_w676_
	);
	LUT4 #(
		.INIT('h5554)
	) name372 (
		_w313_,
		_w675_,
		_w676_,
		_w674_,
		_w677_
	);
	LUT4 #(
		.INIT('h0408)
	) name373 (
		decrypt_pad,
		\key3[46]_pad ,
		\roundSel[4]_pad ,
		\roundSel[5]_pad ,
		_w678_
	);
	LUT3 #(
		.INIT('h08)
	) name374 (
		\key2[46]_pad ,
		\roundSel[4]_pad ,
		\roundSel[5]_pad ,
		_w679_
	);
	LUT4 #(
		.INIT('h0804)
	) name375 (
		decrypt_pad,
		\key1[46]_pad ,
		\roundSel[4]_pad ,
		\roundSel[5]_pad ,
		_w680_
	);
	LUT4 #(
		.INIT('haaa8)
	) name376 (
		_w313_,
		_w679_,
		_w680_,
		_w678_,
		_w681_
	);
	LUT3 #(
		.INIT('ha8)
	) name377 (
		_w333_,
		_w677_,
		_w681_,
		_w682_
	);
	LUT4 #(
		.INIT('h0408)
	) name378 (
		decrypt_pad,
		\key3[33]_pad ,
		\roundSel[4]_pad ,
		\roundSel[5]_pad ,
		_w683_
	);
	LUT3 #(
		.INIT('h08)
	) name379 (
		\key2[33]_pad ,
		\roundSel[4]_pad ,
		\roundSel[5]_pad ,
		_w684_
	);
	LUT4 #(
		.INIT('h0804)
	) name380 (
		decrypt_pad,
		\key1[33]_pad ,
		\roundSel[4]_pad ,
		\roundSel[5]_pad ,
		_w685_
	);
	LUT4 #(
		.INIT('haaa8)
	) name381 (
		_w313_,
		_w684_,
		_w685_,
		_w683_,
		_w686_
	);
	LUT4 #(
		.INIT('h0408)
	) name382 (
		decrypt_pad,
		\key3[40]_pad ,
		\roundSel[4]_pad ,
		\roundSel[5]_pad ,
		_w687_
	);
	LUT3 #(
		.INIT('h08)
	) name383 (
		\key2[40]_pad ,
		\roundSel[4]_pad ,
		\roundSel[5]_pad ,
		_w688_
	);
	LUT4 #(
		.INIT('h0804)
	) name384 (
		decrypt_pad,
		\key1[40]_pad ,
		\roundSel[4]_pad ,
		\roundSel[5]_pad ,
		_w689_
	);
	LUT4 #(
		.INIT('h5554)
	) name385 (
		_w313_,
		_w688_,
		_w689_,
		_w687_,
		_w690_
	);
	LUT3 #(
		.INIT('ha8)
	) name386 (
		_w402_,
		_w686_,
		_w690_,
		_w691_
	);
	LUT4 #(
		.INIT('h0001)
	) name387 (
		_w670_,
		_w673_,
		_w682_,
		_w691_,
		_w692_
	);
	LUT4 #(
		.INIT('h0408)
	) name388 (
		decrypt_pad,
		\key3[24]_pad ,
		\roundSel[4]_pad ,
		\roundSel[5]_pad ,
		_w693_
	);
	LUT3 #(
		.INIT('h08)
	) name389 (
		\key2[24]_pad ,
		\roundSel[4]_pad ,
		\roundSel[5]_pad ,
		_w694_
	);
	LUT4 #(
		.INIT('h0804)
	) name390 (
		decrypt_pad,
		\key1[24]_pad ,
		\roundSel[4]_pad ,
		\roundSel[5]_pad ,
		_w695_
	);
	LUT4 #(
		.INIT('haaa8)
	) name391 (
		_w313_,
		_w694_,
		_w695_,
		_w693_,
		_w696_
	);
	LUT4 #(
		.INIT('h0408)
	) name392 (
		decrypt_pad,
		\key3[17]_pad ,
		\roundSel[4]_pad ,
		\roundSel[5]_pad ,
		_w697_
	);
	LUT3 #(
		.INIT('h08)
	) name393 (
		\key2[17]_pad ,
		\roundSel[4]_pad ,
		\roundSel[5]_pad ,
		_w698_
	);
	LUT4 #(
		.INIT('h0804)
	) name394 (
		decrypt_pad,
		\key1[17]_pad ,
		\roundSel[4]_pad ,
		\roundSel[5]_pad ,
		_w699_
	);
	LUT4 #(
		.INIT('h5554)
	) name395 (
		_w313_,
		_w698_,
		_w699_,
		_w697_,
		_w700_
	);
	LUT3 #(
		.INIT('ha8)
	) name396 (
		_w419_,
		_w696_,
		_w700_,
		_w701_
	);
	LUT4 #(
		.INIT('haaa8)
	) name397 (
		_w313_,
		_w675_,
		_w676_,
		_w674_,
		_w702_
	);
	LUT4 #(
		.INIT('h5554)
	) name398 (
		_w313_,
		_w679_,
		_w680_,
		_w678_,
		_w703_
	);
	LUT3 #(
		.INIT('ha8)
	) name399 (
		_w423_,
		_w702_,
		_w703_,
		_w704_
	);
	LUT4 #(
		.INIT('h0408)
	) name400 (
		decrypt_pad,
		\key3[47]_pad ,
		\roundSel[4]_pad ,
		\roundSel[5]_pad ,
		_w705_
	);
	LUT3 #(
		.INIT('h08)
	) name401 (
		\key2[47]_pad ,
		\roundSel[4]_pad ,
		\roundSel[5]_pad ,
		_w706_
	);
	LUT4 #(
		.INIT('h0804)
	) name402 (
		decrypt_pad,
		\key1[47]_pad ,
		\roundSel[4]_pad ,
		\roundSel[5]_pad ,
		_w707_
	);
	LUT4 #(
		.INIT('h5554)
	) name403 (
		_w313_,
		_w706_,
		_w707_,
		_w705_,
		_w708_
	);
	LUT4 #(
		.INIT('h0408)
	) name404 (
		decrypt_pad,
		\key3[26]_pad ,
		\roundSel[4]_pad ,
		\roundSel[5]_pad ,
		_w709_
	);
	LUT3 #(
		.INIT('h08)
	) name405 (
		\key2[26]_pad ,
		\roundSel[4]_pad ,
		\roundSel[5]_pad ,
		_w710_
	);
	LUT4 #(
		.INIT('h0804)
	) name406 (
		decrypt_pad,
		\key1[26]_pad ,
		\roundSel[4]_pad ,
		\roundSel[5]_pad ,
		_w711_
	);
	LUT4 #(
		.INIT('haaa8)
	) name407 (
		_w313_,
		_w710_,
		_w711_,
		_w709_,
		_w712_
	);
	LUT3 #(
		.INIT('ha8)
	) name408 (
		_w398_,
		_w708_,
		_w712_,
		_w713_
	);
	LUT4 #(
		.INIT('h0408)
	) name409 (
		decrypt_pad,
		\key3[32]_pad ,
		\roundSel[4]_pad ,
		\roundSel[5]_pad ,
		_w714_
	);
	LUT3 #(
		.INIT('h08)
	) name410 (
		\key2[32]_pad ,
		\roundSel[4]_pad ,
		\roundSel[5]_pad ,
		_w715_
	);
	LUT4 #(
		.INIT('h0804)
	) name411 (
		decrypt_pad,
		\key1[32]_pad ,
		\roundSel[4]_pad ,
		\roundSel[5]_pad ,
		_w716_
	);
	LUT4 #(
		.INIT('h5554)
	) name412 (
		_w313_,
		_w715_,
		_w716_,
		_w714_,
		_w717_
	);
	LUT4 #(
		.INIT('h0408)
	) name413 (
		decrypt_pad,
		\key3[41]_pad ,
		\roundSel[4]_pad ,
		\roundSel[5]_pad ,
		_w718_
	);
	LUT3 #(
		.INIT('h08)
	) name414 (
		\key2[41]_pad ,
		\roundSel[4]_pad ,
		\roundSel[5]_pad ,
		_w719_
	);
	LUT4 #(
		.INIT('h0804)
	) name415 (
		decrypt_pad,
		\key1[41]_pad ,
		\roundSel[4]_pad ,
		\roundSel[5]_pad ,
		_w720_
	);
	LUT4 #(
		.INIT('haaa8)
	) name416 (
		_w313_,
		_w719_,
		_w720_,
		_w718_,
		_w721_
	);
	LUT3 #(
		.INIT('ha8)
	) name417 (
		_w373_,
		_w717_,
		_w721_,
		_w722_
	);
	LUT4 #(
		.INIT('h0001)
	) name418 (
		_w701_,
		_w704_,
		_w713_,
		_w722_,
		_w723_
	);
	LUT4 #(
		.INIT('h5554)
	) name419 (
		_w313_,
		_w694_,
		_w695_,
		_w693_,
		_w724_
	);
	LUT4 #(
		.INIT('haaa8)
	) name420 (
		_w313_,
		_w698_,
		_w699_,
		_w697_,
		_w725_
	);
	LUT3 #(
		.INIT('ha8)
	) name421 (
		_w377_,
		_w724_,
		_w725_,
		_w726_
	);
	LUT4 #(
		.INIT('h0408)
	) name422 (
		decrypt_pad,
		\key3[13]_pad ,
		\roundSel[4]_pad ,
		\roundSel[5]_pad ,
		_w727_
	);
	LUT3 #(
		.INIT('h08)
	) name423 (
		\key2[13]_pad ,
		\roundSel[4]_pad ,
		\roundSel[5]_pad ,
		_w728_
	);
	LUT4 #(
		.INIT('h0804)
	) name424 (
		decrypt_pad,
		\key1[13]_pad ,
		\roundSel[4]_pad ,
		\roundSel[5]_pad ,
		_w729_
	);
	LUT4 #(
		.INIT('haaa8)
	) name425 (
		_w313_,
		_w728_,
		_w729_,
		_w727_,
		_w730_
	);
	LUT4 #(
		.INIT('h0408)
	) name426 (
		decrypt_pad,
		\key3[3]_pad ,
		\roundSel[4]_pad ,
		\roundSel[5]_pad ,
		_w731_
	);
	LUT3 #(
		.INIT('h08)
	) name427 (
		\key2[3]_pad ,
		\roundSel[4]_pad ,
		\roundSel[5]_pad ,
		_w732_
	);
	LUT4 #(
		.INIT('h0804)
	) name428 (
		decrypt_pad,
		\key1[3]_pad ,
		\roundSel[4]_pad ,
		\roundSel[5]_pad ,
		_w733_
	);
	LUT4 #(
		.INIT('h5554)
	) name429 (
		_w313_,
		_w732_,
		_w733_,
		_w731_,
		_w734_
	);
	LUT3 #(
		.INIT('ha8)
	) name430 (
		_w411_,
		_w730_,
		_w734_,
		_w735_
	);
	LUT4 #(
		.INIT('h5554)
	) name431 (
		_w313_,
		_w684_,
		_w685_,
		_w683_,
		_w736_
	);
	LUT4 #(
		.INIT('haaa8)
	) name432 (
		_w313_,
		_w688_,
		_w689_,
		_w687_,
		_w737_
	);
	LUT3 #(
		.INIT('ha8)
	) name433 (
		_w305_,
		_w736_,
		_w737_,
		_w738_
	);
	LUT4 #(
		.INIT('haaa8)
	) name434 (
		_w313_,
		_w706_,
		_w707_,
		_w705_,
		_w739_
	);
	LUT4 #(
		.INIT('h5554)
	) name435 (
		_w313_,
		_w710_,
		_w711_,
		_w709_,
		_w740_
	);
	LUT3 #(
		.INIT('ha8)
	) name436 (
		_w312_,
		_w739_,
		_w740_,
		_w741_
	);
	LUT4 #(
		.INIT('h0001)
	) name437 (
		_w726_,
		_w735_,
		_w738_,
		_w741_,
		_w742_
	);
	LUT4 #(
		.INIT('h0408)
	) name438 (
		decrypt_pad,
		\key3[18]_pad ,
		\roundSel[4]_pad ,
		\roundSel[5]_pad ,
		_w743_
	);
	LUT3 #(
		.INIT('h08)
	) name439 (
		\key2[18]_pad ,
		\roundSel[4]_pad ,
		\roundSel[5]_pad ,
		_w744_
	);
	LUT4 #(
		.INIT('h0804)
	) name440 (
		decrypt_pad,
		\key1[18]_pad ,
		\roundSel[4]_pad ,
		\roundSel[5]_pad ,
		_w745_
	);
	LUT4 #(
		.INIT('h5554)
	) name441 (
		_w313_,
		_w744_,
		_w745_,
		_w743_,
		_w746_
	);
	LUT4 #(
		.INIT('h0408)
	) name442 (
		decrypt_pad,
		\key3[55]_pad ,
		\roundSel[4]_pad ,
		\roundSel[5]_pad ,
		_w747_
	);
	LUT3 #(
		.INIT('h08)
	) name443 (
		\key2[55]_pad ,
		\roundSel[4]_pad ,
		\roundSel[5]_pad ,
		_w748_
	);
	LUT4 #(
		.INIT('h0804)
	) name444 (
		decrypt_pad,
		\key1[55]_pad ,
		\roundSel[4]_pad ,
		\roundSel[5]_pad ,
		_w749_
	);
	LUT4 #(
		.INIT('haaa8)
	) name445 (
		_w313_,
		_w748_,
		_w749_,
		_w747_,
		_w750_
	);
	LUT3 #(
		.INIT('ha8)
	) name446 (
		_w388_,
		_w746_,
		_w750_,
		_w751_
	);
	LUT4 #(
		.INIT('h5554)
	) name447 (
		_w313_,
		_w728_,
		_w729_,
		_w727_,
		_w752_
	);
	LUT4 #(
		.INIT('haaa8)
	) name448 (
		_w313_,
		_w732_,
		_w733_,
		_w731_,
		_w753_
	);
	LUT3 #(
		.INIT('ha8)
	) name449 (
		_w323_,
		_w752_,
		_w753_,
		_w754_
	);
	LUT4 #(
		.INIT('haaa8)
	) name450 (
		_w313_,
		_w744_,
		_w745_,
		_w743_,
		_w755_
	);
	LUT4 #(
		.INIT('h5554)
	) name451 (
		_w313_,
		_w748_,
		_w749_,
		_w747_,
		_w756_
	);
	LUT3 #(
		.INIT('ha8)
	) name452 (
		_w406_,
		_w755_,
		_w756_,
		_w757_
	);
	LUT4 #(
		.INIT('haaa8)
	) name453 (
		_w313_,
		_w715_,
		_w716_,
		_w714_,
		_w758_
	);
	LUT4 #(
		.INIT('h5554)
	) name454 (
		_w313_,
		_w719_,
		_w720_,
		_w718_,
		_w759_
	);
	LUT3 #(
		.INIT('ha8)
	) name455 (
		_w343_,
		_w758_,
		_w759_,
		_w760_
	);
	LUT4 #(
		.INIT('h0001)
	) name456 (
		_w751_,
		_w754_,
		_w757_,
		_w760_,
		_w761_
	);
	LUT4 #(
		.INIT('h8000)
	) name457 (
		_w742_,
		_w761_,
		_w692_,
		_w723_,
		_w762_
	);
	LUT2 #(
		.INIT('h9)
	) name458 (
		_w526_,
		_w762_,
		_w763_
	);
	LUT4 #(
		.INIT('h0408)
	) name459 (
		decrypt_pad,
		\key3[53]_pad ,
		\roundSel[4]_pad ,
		\roundSel[5]_pad ,
		_w764_
	);
	LUT3 #(
		.INIT('h08)
	) name460 (
		\key2[53]_pad ,
		\roundSel[4]_pad ,
		\roundSel[5]_pad ,
		_w765_
	);
	LUT4 #(
		.INIT('h0804)
	) name461 (
		decrypt_pad,
		\key1[53]_pad ,
		\roundSel[4]_pad ,
		\roundSel[5]_pad ,
		_w766_
	);
	LUT4 #(
		.INIT('haaa8)
	) name462 (
		_w313_,
		_w765_,
		_w766_,
		_w764_,
		_w767_
	);
	LUT3 #(
		.INIT('ha8)
	) name463 (
		_w411_,
		_w746_,
		_w767_,
		_w768_
	);
	LUT4 #(
		.INIT('h0408)
	) name464 (
		decrypt_pad,
		\key3[39]_pad ,
		\roundSel[4]_pad ,
		\roundSel[5]_pad ,
		_w769_
	);
	LUT3 #(
		.INIT('h08)
	) name465 (
		\key2[39]_pad ,
		\roundSel[4]_pad ,
		\roundSel[5]_pad ,
		_w770_
	);
	LUT4 #(
		.INIT('h0804)
	) name466 (
		decrypt_pad,
		\key1[39]_pad ,
		\roundSel[4]_pad ,
		\roundSel[5]_pad ,
		_w771_
	);
	LUT4 #(
		.INIT('h5554)
	) name467 (
		_w313_,
		_w770_,
		_w771_,
		_w769_,
		_w772_
	);
	LUT3 #(
		.INIT('ha8)
	) name468 (
		_w377_,
		_w758_,
		_w772_,
		_w773_
	);
	LUT4 #(
		.INIT('h5554)
	) name469 (
		_w313_,
		_w765_,
		_w766_,
		_w764_,
		_w774_
	);
	LUT3 #(
		.INIT('ha8)
	) name470 (
		_w323_,
		_w755_,
		_w774_,
		_w775_
	);
	LUT4 #(
		.INIT('h0408)
	) name471 (
		decrypt_pad,
		\key3[19]_pad ,
		\roundSel[4]_pad ,
		\roundSel[5]_pad ,
		_w776_
	);
	LUT3 #(
		.INIT('h08)
	) name472 (
		\key2[19]_pad ,
		\roundSel[4]_pad ,
		\roundSel[5]_pad ,
		_w777_
	);
	LUT4 #(
		.INIT('h0804)
	) name473 (
		decrypt_pad,
		\key1[19]_pad ,
		\roundSel[4]_pad ,
		\roundSel[5]_pad ,
		_w778_
	);
	LUT4 #(
		.INIT('h5554)
	) name474 (
		_w313_,
		_w777_,
		_w778_,
		_w776_,
		_w779_
	);
	LUT3 #(
		.INIT('ha8)
	) name475 (
		_w363_,
		_w702_,
		_w779_,
		_w780_
	);
	LUT4 #(
		.INIT('h0001)
	) name476 (
		_w768_,
		_w773_,
		_w775_,
		_w780_,
		_w781_
	);
	LUT3 #(
		.INIT('ha8)
	) name477 (
		_w343_,
		_w724_,
		_w739_,
		_w782_
	);
	LUT4 #(
		.INIT('h0408)
	) name478 (
		decrypt_pad,
		\key3[48]_pad ,
		\roundSel[4]_pad ,
		\roundSel[5]_pad ,
		_w783_
	);
	LUT3 #(
		.INIT('h08)
	) name479 (
		\key2[48]_pad ,
		\roundSel[4]_pad ,
		\roundSel[5]_pad ,
		_w784_
	);
	LUT4 #(
		.INIT('h0804)
	) name480 (
		decrypt_pad,
		\key1[48]_pad ,
		\roundSel[4]_pad ,
		\roundSel[5]_pad ,
		_w785_
	);
	LUT4 #(
		.INIT('h5554)
	) name481 (
		_w313_,
		_w784_,
		_w785_,
		_w783_,
		_w786_
	);
	LUT3 #(
		.INIT('ha8)
	) name482 (
		_w305_,
		_w750_,
		_w786_,
		_w787_
	);
	LUT4 #(
		.INIT('haaa8)
	) name483 (
		_w313_,
		_w784_,
		_w785_,
		_w783_,
		_w788_
	);
	LUT3 #(
		.INIT('ha8)
	) name484 (
		_w402_,
		_w756_,
		_w788_,
		_w789_
	);
	LUT4 #(
		.INIT('h0408)
	) name485 (
		decrypt_pad,
		\key3[10]_pad ,
		\roundSel[4]_pad ,
		\roundSel[5]_pad ,
		_w790_
	);
	LUT3 #(
		.INIT('h08)
	) name486 (
		\key2[10]_pad ,
		\roundSel[4]_pad ,
		\roundSel[5]_pad ,
		_w791_
	);
	LUT4 #(
		.INIT('h0804)
	) name487 (
		decrypt_pad,
		\key1[10]_pad ,
		\roundSel[4]_pad ,
		\roundSel[5]_pad ,
		_w792_
	);
	LUT4 #(
		.INIT('haaa8)
	) name488 (
		_w313_,
		_w791_,
		_w792_,
		_w790_,
		_w793_
	);
	LUT3 #(
		.INIT('ha8)
	) name489 (
		_w423_,
		_w671_,
		_w793_,
		_w794_
	);
	LUT4 #(
		.INIT('h0001)
	) name490 (
		_w782_,
		_w787_,
		_w789_,
		_w794_,
		_w795_
	);
	LUT3 #(
		.INIT('ha8)
	) name491 (
		_w406_,
		_w686_,
		_w752_,
		_w796_
	);
	LUT4 #(
		.INIT('haaa8)
	) name492 (
		_w313_,
		_w770_,
		_w771_,
		_w769_,
		_w797_
	);
	LUT3 #(
		.INIT('ha8)
	) name493 (
		_w419_,
		_w717_,
		_w797_,
		_w798_
	);
	LUT4 #(
		.INIT('h0408)
	) name494 (
		decrypt_pad,
		\key3[5]_pad ,
		\roundSel[4]_pad ,
		\roundSel[5]_pad ,
		_w799_
	);
	LUT3 #(
		.INIT('h08)
	) name495 (
		\key2[5]_pad ,
		\roundSel[4]_pad ,
		\roundSel[5]_pad ,
		_w800_
	);
	LUT4 #(
		.INIT('h0804)
	) name496 (
		decrypt_pad,
		\key1[5]_pad ,
		\roundSel[4]_pad ,
		\roundSel[5]_pad ,
		_w801_
	);
	LUT4 #(
		.INIT('h5554)
	) name497 (
		_w313_,
		_w800_,
		_w801_,
		_w799_,
		_w802_
	);
	LUT3 #(
		.INIT('ha8)
	) name498 (
		_w398_,
		_w721_,
		_w802_,
		_w803_
	);
	LUT3 #(
		.INIT('ha8)
	) name499 (
		_w388_,
		_w730_,
		_w736_,
		_w804_
	);
	LUT4 #(
		.INIT('h0001)
	) name500 (
		_w796_,
		_w798_,
		_w803_,
		_w804_,
		_w805_
	);
	LUT4 #(
		.INIT('haaa8)
	) name501 (
		_w313_,
		_w800_,
		_w801_,
		_w799_,
		_w806_
	);
	LUT3 #(
		.INIT('ha8)
	) name502 (
		_w312_,
		_w759_,
		_w806_,
		_w807_
	);
	LUT3 #(
		.INIT('ha8)
	) name503 (
		_w373_,
		_w696_,
		_w708_,
		_w808_
	);
	LUT4 #(
		.INIT('h5554)
	) name504 (
		_w313_,
		_w791_,
		_w792_,
		_w790_,
		_w809_
	);
	LUT3 #(
		.INIT('ha8)
	) name505 (
		_w333_,
		_w665_,
		_w809_,
		_w810_
	);
	LUT4 #(
		.INIT('haaa8)
	) name506 (
		_w313_,
		_w777_,
		_w778_,
		_w776_,
		_w811_
	);
	LUT3 #(
		.INIT('ha8)
	) name507 (
		_w415_,
		_w677_,
		_w811_,
		_w812_
	);
	LUT4 #(
		.INIT('h0001)
	) name508 (
		_w807_,
		_w808_,
		_w810_,
		_w812_,
		_w813_
	);
	LUT4 #(
		.INIT('h8000)
	) name509 (
		_w805_,
		_w813_,
		_w781_,
		_w795_,
		_w814_
	);
	LUT4 #(
		.INIT('h0200)
	) name510 (
		\desIn[37]_pad ,
		\roundSel[4]_pad ,
		\roundSel[5]_pad ,
		_w305_,
		_w815_
	);
	LUT4 #(
		.INIT('h4155)
	) name511 (
		\FP_R_reg[13]/P0001 ,
		\roundSel[4]_pad ,
		\roundSel[5]_pad ,
		_w305_,
		_w816_
	);
	LUT4 #(
		.INIT('he8ff)
	) name512 (
		\FP_R_reg[45]/NET0131 ,
		\roundSel[4]_pad ,
		\roundSel[5]_pad ,
		_w305_,
		_w817_
	);
	LUT3 #(
		.INIT('h45)
	) name513 (
		_w815_,
		_w816_,
		_w817_,
		_w818_
	);
	LUT3 #(
		.INIT('hba)
	) name514 (
		_w815_,
		_w816_,
		_w817_,
		_w819_
	);
	LUT2 #(
		.INIT('h9)
	) name515 (
		_w814_,
		_w818_,
		_w820_
	);
	LUT4 #(
		.INIT('h0408)
	) name516 (
		decrypt_pad,
		\key3[20]_pad ,
		\roundSel[4]_pad ,
		\roundSel[5]_pad ,
		_w821_
	);
	LUT3 #(
		.INIT('h08)
	) name517 (
		\key2[20]_pad ,
		\roundSel[4]_pad ,
		\roundSel[5]_pad ,
		_w822_
	);
	LUT4 #(
		.INIT('h0804)
	) name518 (
		decrypt_pad,
		\key1[20]_pad ,
		\roundSel[4]_pad ,
		\roundSel[5]_pad ,
		_w823_
	);
	LUT4 #(
		.INIT('h5554)
	) name519 (
		_w313_,
		_w822_,
		_w823_,
		_w821_,
		_w824_
	);
	LUT3 #(
		.INIT('ha8)
	) name520 (
		_w363_,
		_w824_,
		_w767_,
		_w825_
	);
	LUT3 #(
		.INIT('ha8)
	) name521 (
		_w377_,
		_w686_,
		_w690_,
		_w826_
	);
	LUT3 #(
		.INIT('ha8)
	) name522 (
		_w402_,
		_w724_,
		_w725_,
		_w827_
	);
	LUT4 #(
		.INIT('h0408)
	) name523 (
		decrypt_pad,
		\key3[6]_pad ,
		\roundSel[4]_pad ,
		\roundSel[5]_pad ,
		_w828_
	);
	LUT3 #(
		.INIT('h08)
	) name524 (
		\key2[6]_pad ,
		\roundSel[4]_pad ,
		\roundSel[5]_pad ,
		_w829_
	);
	LUT4 #(
		.INIT('h0804)
	) name525 (
		decrypt_pad,
		\key1[6]_pad ,
		\roundSel[4]_pad ,
		\roundSel[5]_pad ,
		_w830_
	);
	LUT4 #(
		.INIT('h5554)
	) name526 (
		_w313_,
		_w829_,
		_w830_,
		_w828_,
		_w831_
	);
	LUT3 #(
		.INIT('ha8)
	) name527 (
		_w398_,
		_w793_,
		_w831_,
		_w832_
	);
	LUT4 #(
		.INIT('h0001)
	) name528 (
		_w825_,
		_w826_,
		_w827_,
		_w832_,
		_w833_
	);
	LUT4 #(
		.INIT('h0408)
	) name529 (
		decrypt_pad,
		\key3[11]_pad ,
		\roundSel[4]_pad ,
		\roundSel[5]_pad ,
		_w834_
	);
	LUT3 #(
		.INIT('h08)
	) name530 (
		\key2[11]_pad ,
		\roundSel[4]_pad ,
		\roundSel[5]_pad ,
		_w835_
	);
	LUT4 #(
		.INIT('h0804)
	) name531 (
		decrypt_pad,
		\key1[11]_pad ,
		\roundSel[4]_pad ,
		\roundSel[5]_pad ,
		_w836_
	);
	LUT4 #(
		.INIT('h5554)
	) name532 (
		_w313_,
		_w835_,
		_w836_,
		_w834_,
		_w837_
	);
	LUT3 #(
		.INIT('ha8)
	) name533 (
		_w333_,
		_w837_,
		_w806_,
		_w838_
	);
	LUT4 #(
		.INIT('h0408)
	) name534 (
		decrypt_pad,
		\key3[34]_pad ,
		\roundSel[4]_pad ,
		\roundSel[5]_pad ,
		_w839_
	);
	LUT3 #(
		.INIT('h08)
	) name535 (
		\key2[34]_pad ,
		\roundSel[4]_pad ,
		\roundSel[5]_pad ,
		_w840_
	);
	LUT4 #(
		.INIT('h0804)
	) name536 (
		decrypt_pad,
		\key1[34]_pad ,
		\roundSel[4]_pad ,
		\roundSel[5]_pad ,
		_w841_
	);
	LUT4 #(
		.INIT('haaa8)
	) name537 (
		_w313_,
		_w840_,
		_w841_,
		_w839_,
		_w842_
	);
	LUT3 #(
		.INIT('ha8)
	) name538 (
		_w406_,
		_w842_,
		_w772_,
		_w843_
	);
	LUT4 #(
		.INIT('h0408)
	) name539 (
		decrypt_pad,
		\key3[25]_pad ,
		\roundSel[4]_pad ,
		\roundSel[5]_pad ,
		_w844_
	);
	LUT3 #(
		.INIT('h08)
	) name540 (
		\key2[25]_pad ,
		\roundSel[4]_pad ,
		\roundSel[5]_pad ,
		_w845_
	);
	LUT4 #(
		.INIT('h0804)
	) name541 (
		decrypt_pad,
		\key1[25]_pad ,
		\roundSel[4]_pad ,
		\roundSel[5]_pad ,
		_w846_
	);
	LUT4 #(
		.INIT('haaa8)
	) name542 (
		_w313_,
		_w845_,
		_w846_,
		_w844_,
		_w847_
	);
	LUT3 #(
		.INIT('ha8)
	) name543 (
		_w373_,
		_w847_,
		_w786_,
		_w848_
	);
	LUT4 #(
		.INIT('haaa8)
	) name544 (
		_w313_,
		_w829_,
		_w830_,
		_w828_,
		_w849_
	);
	LUT3 #(
		.INIT('ha8)
	) name545 (
		_w312_,
		_w809_,
		_w849_,
		_w850_
	);
	LUT4 #(
		.INIT('h0001)
	) name546 (
		_w838_,
		_w843_,
		_w848_,
		_w850_,
		_w851_
	);
	LUT3 #(
		.INIT('ha8)
	) name547 (
		_w419_,
		_w736_,
		_w737_,
		_w852_
	);
	LUT4 #(
		.INIT('h0408)
	) name548 (
		decrypt_pad,
		\key3[54]_pad ,
		\roundSel[4]_pad ,
		\roundSel[5]_pad ,
		_w853_
	);
	LUT3 #(
		.INIT('h08)
	) name549 (
		\key2[54]_pad ,
		\roundSel[4]_pad ,
		\roundSel[5]_pad ,
		_w854_
	);
	LUT4 #(
		.INIT('h0804)
	) name550 (
		decrypt_pad,
		\key1[54]_pad ,
		\roundSel[4]_pad ,
		\roundSel[5]_pad ,
		_w855_
	);
	LUT4 #(
		.INIT('h5554)
	) name551 (
		_w313_,
		_w854_,
		_w855_,
		_w853_,
		_w856_
	);
	LUT3 #(
		.INIT('ha8)
	) name552 (
		_w323_,
		_w856_,
		_w811_,
		_w857_
	);
	LUT4 #(
		.INIT('haaa8)
	) name553 (
		_w313_,
		_w835_,
		_w836_,
		_w834_,
		_w858_
	);
	LUT3 #(
		.INIT('ha8)
	) name554 (
		_w423_,
		_w802_,
		_w858_,
		_w859_
	);
	LUT4 #(
		.INIT('haaa8)
	) name555 (
		_w313_,
		_w822_,
		_w823_,
		_w821_,
		_w860_
	);
	LUT3 #(
		.INIT('ha8)
	) name556 (
		_w415_,
		_w860_,
		_w774_,
		_w861_
	);
	LUT4 #(
		.INIT('h0001)
	) name557 (
		_w852_,
		_w857_,
		_w859_,
		_w861_,
		_w862_
	);
	LUT4 #(
		.INIT('h5554)
	) name558 (
		_w313_,
		_w840_,
		_w841_,
		_w839_,
		_w863_
	);
	LUT3 #(
		.INIT('ha8)
	) name559 (
		_w388_,
		_w863_,
		_w797_,
		_w864_
	);
	LUT4 #(
		.INIT('haaa8)
	) name560 (
		_w313_,
		_w854_,
		_w855_,
		_w853_,
		_w865_
	);
	LUT3 #(
		.INIT('ha8)
	) name561 (
		_w411_,
		_w865_,
		_w779_,
		_w866_
	);
	LUT3 #(
		.INIT('ha8)
	) name562 (
		_w305_,
		_w696_,
		_w700_,
		_w867_
	);
	LUT4 #(
		.INIT('h5554)
	) name563 (
		_w313_,
		_w845_,
		_w846_,
		_w844_,
		_w868_
	);
	LUT3 #(
		.INIT('ha8)
	) name564 (
		_w343_,
		_w868_,
		_w788_,
		_w869_
	);
	LUT4 #(
		.INIT('h0001)
	) name565 (
		_w864_,
		_w866_,
		_w867_,
		_w869_,
		_w870_
	);
	LUT4 #(
		.INIT('h8000)
	) name566 (
		_w862_,
		_w870_,
		_w833_,
		_w851_,
		_w871_
	);
	LUT4 #(
		.INIT('h0200)
	) name567 (
		\desIn[45]_pad ,
		\roundSel[4]_pad ,
		\roundSel[5]_pad ,
		_w305_,
		_w872_
	);
	LUT4 #(
		.INIT('h4155)
	) name568 (
		\FP_R_reg[14]/P0001 ,
		\roundSel[4]_pad ,
		\roundSel[5]_pad ,
		_w305_,
		_w873_
	);
	LUT4 #(
		.INIT('he8ff)
	) name569 (
		\FP_R_reg[46]/NET0131 ,
		\roundSel[4]_pad ,
		\roundSel[5]_pad ,
		_w305_,
		_w874_
	);
	LUT3 #(
		.INIT('h45)
	) name570 (
		_w872_,
		_w873_,
		_w874_,
		_w875_
	);
	LUT3 #(
		.INIT('hba)
	) name571 (
		_w872_,
		_w873_,
		_w874_,
		_w876_
	);
	LUT2 #(
		.INIT('h6)
	) name572 (
		_w871_,
		_w875_,
		_w877_
	);
	LUT4 #(
		.INIT('h0990)
	) name573 (
		_w814_,
		_w818_,
		_w871_,
		_w875_,
		_w878_
	);
	LUT3 #(
		.INIT('ha8)
	) name574 (
		_w343_,
		_w767_,
		_w802_,
		_w879_
	);
	LUT3 #(
		.INIT('ha8)
	) name575 (
		_w402_,
		_w671_,
		_w865_,
		_w880_
	);
	LUT3 #(
		.INIT('ha8)
	) name576 (
		_w411_,
		_w724_,
		_w842_,
		_w881_
	);
	LUT3 #(
		.INIT('ha8)
	) name577 (
		_w323_,
		_w696_,
		_w863_,
		_w882_
	);
	LUT4 #(
		.INIT('h0001)
	) name578 (
		_w879_,
		_w880_,
		_w881_,
		_w882_,
		_w883_
	);
	LUT3 #(
		.INIT('ha8)
	) name579 (
		_w305_,
		_w665_,
		_w856_,
		_w884_
	);
	LUT3 #(
		.INIT('ha8)
	) name580 (
		_w377_,
		_w730_,
		_w824_,
		_w885_
	);
	LUT3 #(
		.INIT('ha8)
	) name581 (
		_w419_,
		_w752_,
		_w860_,
		_w886_
	);
	LUT3 #(
		.INIT('ha8)
	) name582 (
		_w363_,
		_w686_,
		_w868_,
		_w887_
	);
	LUT4 #(
		.INIT('h0001)
	) name583 (
		_w884_,
		_w885_,
		_w886_,
		_w887_,
		_w888_
	);
	LUT3 #(
		.INIT('ha8)
	) name584 (
		_w423_,
		_w788_,
		_w809_,
		_w889_
	);
	LUT3 #(
		.INIT('ha8)
	) name585 (
		_w398_,
		_w739_,
		_w837_,
		_w890_
	);
	LUT3 #(
		.INIT('ha8)
	) name586 (
		_w373_,
		_w774_,
		_w806_,
		_w891_
	);
	LUT3 #(
		.INIT('ha8)
	) name587 (
		_w388_,
		_w772_,
		_w811_,
		_w892_
	);
	LUT4 #(
		.INIT('h0001)
	) name588 (
		_w889_,
		_w890_,
		_w891_,
		_w892_,
		_w893_
	);
	LUT3 #(
		.INIT('ha8)
	) name589 (
		_w415_,
		_w736_,
		_w847_,
		_w894_
	);
	LUT3 #(
		.INIT('ha8)
	) name590 (
		_w333_,
		_w786_,
		_w793_,
		_w895_
	);
	LUT3 #(
		.INIT('ha8)
	) name591 (
		_w312_,
		_w708_,
		_w858_,
		_w896_
	);
	LUT3 #(
		.INIT('ha8)
	) name592 (
		_w406_,
		_w779_,
		_w797_,
		_w897_
	);
	LUT4 #(
		.INIT('h0001)
	) name593 (
		_w894_,
		_w895_,
		_w896_,
		_w897_,
		_w898_
	);
	LUT4 #(
		.INIT('h8000)
	) name594 (
		_w893_,
		_w898_,
		_w883_,
		_w888_,
		_w899_
	);
	LUT3 #(
		.INIT('h40)
	) name595 (
		\FP_R_reg[44]/NET0131 ,
		_w305_,
		_w307_,
		_w900_
	);
	LUT4 #(
		.INIT('hb0aa)
	) name596 (
		\FP_R_reg[12]/P0001 ,
		\roundSel[4]_pad ,
		\roundSel[5]_pad ,
		_w305_,
		_w901_
	);
	LUT4 #(
		.INIT('h0800)
	) name597 (
		\FP_R_reg[44]/NET0131 ,
		\roundSel[4]_pad ,
		\roundSel[5]_pad ,
		_w305_,
		_w902_
	);
	LUT4 #(
		.INIT('h0200)
	) name598 (
		\desIn[29]_pad ,
		\roundSel[4]_pad ,
		\roundSel[5]_pad ,
		_w305_,
		_w903_
	);
	LUT4 #(
		.INIT('h1011)
	) name599 (
		_w902_,
		_w903_,
		_w900_,
		_w901_,
		_w904_
	);
	LUT4 #(
		.INIT('hefee)
	) name600 (
		_w902_,
		_w903_,
		_w900_,
		_w901_,
		_w905_
	);
	LUT2 #(
		.INIT('h9)
	) name601 (
		_w899_,
		_w904_,
		_w906_
	);
	LUT3 #(
		.INIT('ha8)
	) name602 (
		_w388_,
		_w753_,
		_w756_,
		_w907_
	);
	LUT3 #(
		.INIT('ha8)
	) name603 (
		_w419_,
		_w665_,
		_w856_,
		_w908_
	);
	LUT3 #(
		.INIT('ha8)
	) name604 (
		_w333_,
		_w712_,
		_w717_,
		_w909_
	);
	LUT3 #(
		.INIT('ha8)
	) name605 (
		_w373_,
		_w669_,
		_w681_,
		_w910_
	);
	LUT4 #(
		.INIT('h0001)
	) name606 (
		_w907_,
		_w908_,
		_w909_,
		_w910_,
		_w911_
	);
	LUT3 #(
		.INIT('ha8)
	) name607 (
		_w323_,
		_w746_,
		_w737_,
		_w912_
	);
	LUT3 #(
		.INIT('ha8)
	) name608 (
		_w377_,
		_w671_,
		_w865_,
		_w913_
	);
	LUT3 #(
		.INIT('ha8)
	) name609 (
		_w305_,
		_w752_,
		_w860_,
		_w914_
	);
	LUT3 #(
		.INIT('ha8)
	) name610 (
		_w411_,
		_w690_,
		_w755_,
		_w915_
	);
	LUT4 #(
		.INIT('h0001)
	) name611 (
		_w912_,
		_w913_,
		_w914_,
		_w915_,
		_w916_
	);
	LUT3 #(
		.INIT('ha8)
	) name612 (
		_w398_,
		_w677_,
		_w849_,
		_w917_
	);
	LUT3 #(
		.INIT('ha8)
	) name613 (
		_w402_,
		_w730_,
		_w824_,
		_w918_
	);
	LUT3 #(
		.INIT('ha8)
	) name614 (
		_w415_,
		_w700_,
		_w721_,
		_w919_
	);
	LUT3 #(
		.INIT('ha8)
	) name615 (
		_w312_,
		_w702_,
		_w831_,
		_w920_
	);
	LUT4 #(
		.INIT('h0001)
	) name616 (
		_w917_,
		_w918_,
		_w919_,
		_w920_,
		_w921_
	);
	LUT3 #(
		.INIT('ha8)
	) name617 (
		_w406_,
		_w750_,
		_w734_,
		_w922_
	);
	LUT3 #(
		.INIT('ha8)
	) name618 (
		_w343_,
		_w703_,
		_w672_,
		_w923_
	);
	LUT3 #(
		.INIT('ha8)
	) name619 (
		_w363_,
		_w759_,
		_w725_,
		_w924_
	);
	LUT3 #(
		.INIT('ha8)
	) name620 (
		_w423_,
		_w758_,
		_w740_,
		_w925_
	);
	LUT4 #(
		.INIT('h0001)
	) name621 (
		_w922_,
		_w923_,
		_w924_,
		_w925_,
		_w926_
	);
	LUT4 #(
		.INIT('h8000)
	) name622 (
		_w921_,
		_w926_,
		_w911_,
		_w916_,
		_w927_
	);
	LUT2 #(
		.INIT('h9)
	) name623 (
		_w499_,
		_w927_,
		_w928_
	);
	LUT4 #(
		.INIT('h4182)
	) name624 (
		_w499_,
		_w899_,
		_w904_,
		_w927_,
		_w929_
	);
	LUT3 #(
		.INIT('ha8)
	) name625 (
		_w323_,
		_w702_,
		_w802_,
		_w930_
	);
	LUT3 #(
		.INIT('ha8)
	) name626 (
		_w419_,
		_w759_,
		_w788_,
		_w931_
	);
	LUT3 #(
		.INIT('ha8)
	) name627 (
		_w305_,
		_w758_,
		_w868_,
		_w932_
	);
	LUT3 #(
		.INIT('ha8)
	) name628 (
		_w373_,
		_w686_,
		_w724_,
		_w933_
	);
	LUT4 #(
		.INIT('h0001)
	) name629 (
		_w930_,
		_w931_,
		_w932_,
		_w933_,
		_w934_
	);
	LUT3 #(
		.INIT('ha8)
	) name630 (
		_w406_,
		_w708_,
		_w793_,
		_w935_
	);
	LUT3 #(
		.INIT('ha8)
	) name631 (
		_w398_,
		_w755_,
		_w772_,
		_w936_
	);
	LUT3 #(
		.INIT('ha8)
	) name632 (
		_w388_,
		_w739_,
		_w809_,
		_w937_
	);
	LUT3 #(
		.INIT('ha8)
	) name633 (
		_w363_,
		_w665_,
		_w774_,
		_w938_
	);
	LUT4 #(
		.INIT('h0001)
	) name634 (
		_w935_,
		_w936_,
		_w937_,
		_w938_,
		_w939_
	);
	LUT3 #(
		.INIT('ha8)
	) name635 (
		_w377_,
		_w721_,
		_w786_,
		_w940_
	);
	LUT3 #(
		.INIT('ha8)
	) name636 (
		_w333_,
		_w730_,
		_w779_,
		_w941_
	);
	LUT3 #(
		.INIT('ha8)
	) name637 (
		_w312_,
		_w746_,
		_w797_,
		_w942_
	);
	LUT3 #(
		.INIT('ha8)
	) name638 (
		_w423_,
		_w752_,
		_w811_,
		_w943_
	);
	LUT4 #(
		.INIT('h0001)
	) name639 (
		_w940_,
		_w941_,
		_w942_,
		_w943_,
		_w944_
	);
	LUT3 #(
		.INIT('ha8)
	) name640 (
		_w343_,
		_w696_,
		_w736_,
		_w945_
	);
	LUT3 #(
		.INIT('ha8)
	) name641 (
		_w415_,
		_w671_,
		_w767_,
		_w946_
	);
	LUT3 #(
		.INIT('ha8)
	) name642 (
		_w402_,
		_w717_,
		_w847_,
		_w947_
	);
	LUT3 #(
		.INIT('ha8)
	) name643 (
		_w411_,
		_w677_,
		_w806_,
		_w948_
	);
	LUT4 #(
		.INIT('h0001)
	) name644 (
		_w945_,
		_w946_,
		_w947_,
		_w948_,
		_w949_
	);
	LUT4 #(
		.INIT('h8000)
	) name645 (
		_w944_,
		_w949_,
		_w934_,
		_w939_,
		_w950_
	);
	LUT4 #(
		.INIT('h0200)
	) name646 (
		\desIn[53]_pad ,
		\roundSel[4]_pad ,
		\roundSel[5]_pad ,
		_w305_,
		_w951_
	);
	LUT4 #(
		.INIT('h4155)
	) name647 (
		\FP_R_reg[15]/P0001 ,
		\roundSel[4]_pad ,
		\roundSel[5]_pad ,
		_w305_,
		_w952_
	);
	LUT4 #(
		.INIT('he8ff)
	) name648 (
		\FP_R_reg[47]/NET0131 ,
		\roundSel[4]_pad ,
		\roundSel[5]_pad ,
		_w305_,
		_w953_
	);
	LUT3 #(
		.INIT('h45)
	) name649 (
		_w951_,
		_w952_,
		_w953_,
		_w954_
	);
	LUT3 #(
		.INIT('hba)
	) name650 (
		_w951_,
		_w952_,
		_w953_,
		_w955_
	);
	LUT2 #(
		.INIT('h9)
	) name651 (
		_w950_,
		_w954_,
		_w956_
	);
	LUT4 #(
		.INIT('h2814)
	) name652 (
		_w499_,
		_w899_,
		_w904_,
		_w927_,
		_w957_
	);
	LUT4 #(
		.INIT('h0042)
	) name653 (
		_w906_,
		_w878_,
		_w928_,
		_w956_,
		_w958_
	);
	LUT4 #(
		.INIT('h8241)
	) name654 (
		_w499_,
		_w899_,
		_w904_,
		_w927_,
		_w959_
	);
	LUT4 #(
		.INIT('h6006)
	) name655 (
		_w814_,
		_w818_,
		_w871_,
		_w875_,
		_w960_
	);
	LUT4 #(
		.INIT('hcdef)
	) name656 (
		_w820_,
		_w877_,
		_w957_,
		_w959_,
		_w961_
	);
	LUT4 #(
		.INIT('h1428)
	) name657 (
		_w499_,
		_w899_,
		_w904_,
		_w927_,
		_w962_
	);
	LUT4 #(
		.INIT('h9009)
	) name658 (
		_w814_,
		_w818_,
		_w950_,
		_w954_,
		_w963_
	);
	LUT2 #(
		.INIT('h8)
	) name659 (
		_w962_,
		_w963_,
		_w964_
	);
	LUT4 #(
		.INIT('h0660)
	) name660 (
		_w814_,
		_w818_,
		_w871_,
		_w875_,
		_w965_
	);
	LUT4 #(
		.INIT('h9009)
	) name661 (
		_w899_,
		_w904_,
		_w950_,
		_w954_,
		_w966_
	);
	LUT3 #(
		.INIT('h80)
	) name662 (
		_w928_,
		_w966_,
		_w965_,
		_w967_
	);
	LUT4 #(
		.INIT('h0002)
	) name663 (
		_w961_,
		_w964_,
		_w967_,
		_w958_,
		_w968_
	);
	LUT2 #(
		.INIT('h2)
	) name664 (
		_w763_,
		_w968_,
		_w969_
	);
	LUT3 #(
		.INIT('h80)
	) name665 (
		_w877_,
		_w956_,
		_w957_,
		_w970_
	);
	LUT4 #(
		.INIT('h1428)
	) name666 (
		_w499_,
		_w814_,
		_w818_,
		_w927_,
		_w971_
	);
	LUT3 #(
		.INIT('ha8)
	) name667 (
		_w966_,
		_w960_,
		_w971_,
		_w972_
	);
	LUT4 #(
		.INIT('h0660)
	) name668 (
		_w814_,
		_w818_,
		_w950_,
		_w954_,
		_w973_
	);
	LUT2 #(
		.INIT('h8)
	) name669 (
		_w962_,
		_w973_,
		_w974_
	);
	LUT3 #(
		.INIT('h01)
	) name670 (
		_w972_,
		_w970_,
		_w974_,
		_w975_
	);
	LUT4 #(
		.INIT('h0660)
	) name671 (
		_w871_,
		_w875_,
		_w950_,
		_w954_,
		_w976_
	);
	LUT4 #(
		.INIT('ha888)
	) name672 (
		_w906_,
		_w878_,
		_w928_,
		_w976_,
		_w977_
	);
	LUT4 #(
		.INIT('h6006)
	) name673 (
		_w899_,
		_w904_,
		_w814_,
		_w818_,
		_w978_
	);
	LUT3 #(
		.INIT('h10)
	) name674 (
		_w877_,
		_w928_,
		_w978_,
		_w979_
	);
	LUT3 #(
		.INIT('h40)
	) name675 (
		_w820_,
		_w877_,
		_w962_,
		_w980_
	);
	LUT4 #(
		.INIT('hffeb)
	) name676 (
		_w906_,
		_w820_,
		_w877_,
		_w928_,
		_w981_
	);
	LUT2 #(
		.INIT('h4)
	) name677 (
		_w977_,
		_w981_,
		_w982_
	);
	LUT3 #(
		.INIT('h15)
	) name678 (
		_w763_,
		_w975_,
		_w982_,
		_w983_
	);
	LUT3 #(
		.INIT('h45)
	) name679 (
		_w956_,
		_w980_,
		_w961_,
		_w984_
	);
	LUT3 #(
		.INIT('h40)
	) name680 (
		_w877_,
		_w956_,
		_w978_,
		_w985_
	);
	LUT3 #(
		.INIT('h80)
	) name681 (
		_w877_,
		_w963_,
		_w929_,
		_w986_
	);
	LUT2 #(
		.INIT('h1)
	) name682 (
		_w985_,
		_w986_,
		_w987_
	);
	LUT2 #(
		.INIT('h4)
	) name683 (
		_w984_,
		_w987_,
		_w988_
	);
	LUT4 #(
		.INIT('h0100)
	) name684 (
		\desIn[12]_pad ,
		\roundSel[4]_pad ,
		\roundSel[5]_pad ,
		_w305_,
		_w989_
	);
	LUT4 #(
		.INIT('h2800)
	) name685 (
		\FP_R_reg[10]/P0001 ,
		\roundSel[4]_pad ,
		\roundSel[5]_pad ,
		_w305_,
		_w990_
	);
	LUT4 #(
		.INIT('h7c55)
	) name686 (
		\FP_R_reg[42]/NET0131 ,
		\roundSel[4]_pad ,
		\roundSel[5]_pad ,
		_w305_,
		_w991_
	);
	LUT3 #(
		.INIT('h45)
	) name687 (
		_w989_,
		_w990_,
		_w991_,
		_w992_
	);
	LUT4 #(
		.INIT('h10ef)
	) name688 (
		_w983_,
		_w969_,
		_w988_,
		_w992_,
		_w993_
	);
	LUT4 #(
		.INIT('h0200)
	) name689 (
		\desIn[13]_pad ,
		\roundSel[4]_pad ,
		\roundSel[5]_pad ,
		_w305_,
		_w994_
	);
	LUT4 #(
		.INIT('h4155)
	) name690 (
		\FP_R_reg[10]/P0001 ,
		\roundSel[4]_pad ,
		\roundSel[5]_pad ,
		_w305_,
		_w995_
	);
	LUT4 #(
		.INIT('he8ff)
	) name691 (
		\FP_R_reg[42]/NET0131 ,
		\roundSel[4]_pad ,
		\roundSel[5]_pad ,
		_w305_,
		_w996_
	);
	LUT3 #(
		.INIT('h45)
	) name692 (
		_w994_,
		_w995_,
		_w996_,
		_w997_
	);
	LUT3 #(
		.INIT('hba)
	) name693 (
		_w994_,
		_w995_,
		_w996_,
		_w998_
	);
	LUT4 #(
		.INIT('h0200)
	) name694 (
		\desIn[63]_pad ,
		\roundSel[4]_pad ,
		\roundSel[5]_pad ,
		_w305_,
		_w999_
	);
	LUT4 #(
		.INIT('h4155)
	) name695 (
		\FP_R_reg[8]/P0001 ,
		\roundSel[4]_pad ,
		\roundSel[5]_pad ,
		_w305_,
		_w1000_
	);
	LUT4 #(
		.INIT('he8ff)
	) name696 (
		\FP_R_reg[40]/NET0131 ,
		\roundSel[4]_pad ,
		\roundSel[5]_pad ,
		_w305_,
		_w1001_
	);
	LUT3 #(
		.INIT('h45)
	) name697 (
		_w999_,
		_w1000_,
		_w1001_,
		_w1002_
	);
	LUT3 #(
		.INIT('hba)
	) name698 (
		_w999_,
		_w1000_,
		_w1001_,
		_w1003_
	);
	LUT3 #(
		.INIT('ha8)
	) name699 (
		_w411_,
		_w672_,
		_w863_,
		_w1004_
	);
	LUT3 #(
		.INIT('ha8)
	) name700 (
		_w415_,
		_w753_,
		_w837_,
		_w1005_
	);
	LUT3 #(
		.INIT('ha8)
	) name701 (
		_w406_,
		_w725_,
		_w856_,
		_w1006_
	);
	LUT3 #(
		.INIT('ha8)
	) name702 (
		_w377_,
		_w756_,
		_w788_,
		_w1007_
	);
	LUT4 #(
		.INIT('h0001)
	) name703 (
		_w1004_,
		_w1005_,
		_w1006_,
		_w1007_,
		_w1008_
	);
	LUT3 #(
		.INIT('ha8)
	) name704 (
		_w305_,
		_w717_,
		_w797_,
		_w1009_
	);
	LUT3 #(
		.INIT('ha8)
	) name705 (
		_w388_,
		_w700_,
		_w865_,
		_w1010_
	);
	LUT3 #(
		.INIT('ha8)
	) name706 (
		_w373_,
		_w737_,
		_w831_,
		_w1011_
	);
	LUT3 #(
		.INIT('ha8)
	) name707 (
		_w343_,
		_w690_,
		_w849_,
		_w1012_
	);
	LUT4 #(
		.INIT('h0001)
	) name708 (
		_w1009_,
		_w1010_,
		_w1011_,
		_w1012_,
		_w1013_
	);
	LUT3 #(
		.INIT('ha8)
	) name709 (
		_w419_,
		_w750_,
		_w786_,
		_w1014_
	);
	LUT3 #(
		.INIT('ha8)
	) name710 (
		_w312_,
		_w681_,
		_w868_,
		_w1015_
	);
	LUT3 #(
		.INIT('ha8)
	) name711 (
		_w402_,
		_w758_,
		_w772_,
		_w1016_
	);
	LUT3 #(
		.INIT('ha8)
	) name712 (
		_w423_,
		_w712_,
		_w824_,
		_w1017_
	);
	LUT4 #(
		.INIT('h0001)
	) name713 (
		_w1014_,
		_w1015_,
		_w1016_,
		_w1017_,
		_w1018_
	);
	LUT3 #(
		.INIT('ha8)
	) name714 (
		_w363_,
		_w734_,
		_w858_,
		_w1019_
	);
	LUT3 #(
		.INIT('ha8)
	) name715 (
		_w333_,
		_w740_,
		_w860_,
		_w1020_
	);
	LUT3 #(
		.INIT('ha8)
	) name716 (
		_w398_,
		_w703_,
		_w847_,
		_w1021_
	);
	LUT3 #(
		.INIT('ha8)
	) name717 (
		_w323_,
		_w669_,
		_w842_,
		_w1022_
	);
	LUT4 #(
		.INIT('h0001)
	) name718 (
		_w1019_,
		_w1020_,
		_w1021_,
		_w1022_,
		_w1023_
	);
	LUT4 #(
		.INIT('h8000)
	) name719 (
		_w1018_,
		_w1023_,
		_w1008_,
		_w1013_,
		_w1024_
	);
	LUT2 #(
		.INIT('h6)
	) name720 (
		_w1002_,
		_w1024_,
		_w1025_
	);
	LUT3 #(
		.INIT('ha8)
	) name721 (
		_w419_,
		_w758_,
		_w868_,
		_w1026_
	);
	LUT3 #(
		.INIT('ha8)
	) name722 (
		_w363_,
		_w669_,
		_w860_,
		_w1027_
	);
	LUT3 #(
		.INIT('ha8)
	) name723 (
		_w398_,
		_w756_,
		_w842_,
		_w1028_
	);
	LUT3 #(
		.INIT('ha8)
	) name724 (
		_w343_,
		_w700_,
		_w737_,
		_w1029_
	);
	LUT4 #(
		.INIT('h0001)
	) name725 (
		_w1026_,
		_w1027_,
		_w1028_,
		_w1029_,
		_w1030_
	);
	LUT3 #(
		.INIT('ha8)
	) name726 (
		_w305_,
		_w759_,
		_w788_,
		_w1031_
	);
	LUT3 #(
		.INIT('ha8)
	) name727 (
		_w411_,
		_w681_,
		_w837_,
		_w1032_
	);
	LUT3 #(
		.INIT('ha8)
	) name728 (
		_w388_,
		_w740_,
		_w849_,
		_w1033_
	);
	LUT3 #(
		.INIT('ha8)
	) name729 (
		_w373_,
		_w690_,
		_w725_,
		_w1034_
	);
	LUT4 #(
		.INIT('h0001)
	) name730 (
		_w1031_,
		_w1032_,
		_w1033_,
		_w1034_,
		_w1035_
	);
	LUT3 #(
		.INIT('ha8)
	) name731 (
		_w333_,
		_w734_,
		_w865_,
		_w1036_
	);
	LUT3 #(
		.INIT('ha8)
	) name732 (
		_w402_,
		_w721_,
		_w786_,
		_w1037_
	);
	LUT3 #(
		.INIT('ha8)
	) name733 (
		_w415_,
		_w672_,
		_w824_,
		_w1038_
	);
	LUT3 #(
		.INIT('ha8)
	) name734 (
		_w312_,
		_w750_,
		_w863_,
		_w1039_
	);
	LUT4 #(
		.INIT('h0001)
	) name735 (
		_w1036_,
		_w1037_,
		_w1038_,
		_w1039_,
		_w1040_
	);
	LUT3 #(
		.INIT('ha8)
	) name736 (
		_w406_,
		_w712_,
		_w831_,
		_w1041_
	);
	LUT3 #(
		.INIT('ha8)
	) name737 (
		_w323_,
		_w703_,
		_w858_,
		_w1042_
	);
	LUT3 #(
		.INIT('ha8)
	) name738 (
		_w377_,
		_w717_,
		_w847_,
		_w1043_
	);
	LUT3 #(
		.INIT('ha8)
	) name739 (
		_w423_,
		_w753_,
		_w856_,
		_w1044_
	);
	LUT4 #(
		.INIT('h0001)
	) name740 (
		_w1041_,
		_w1042_,
		_w1043_,
		_w1044_,
		_w1045_
	);
	LUT4 #(
		.INIT('h8000)
	) name741 (
		_w1040_,
		_w1045_,
		_w1030_,
		_w1035_,
		_w1046_
	);
	LUT3 #(
		.INIT('h40)
	) name742 (
		\FP_R_reg[39]/NET0131 ,
		_w305_,
		_w307_,
		_w1047_
	);
	LUT4 #(
		.INIT('hb0aa)
	) name743 (
		\FP_R_reg[7]/P0001 ,
		\roundSel[4]_pad ,
		\roundSel[5]_pad ,
		_w305_,
		_w1048_
	);
	LUT4 #(
		.INIT('h0800)
	) name744 (
		\FP_R_reg[39]/NET0131 ,
		\roundSel[4]_pad ,
		\roundSel[5]_pad ,
		_w305_,
		_w1049_
	);
	LUT4 #(
		.INIT('h0200)
	) name745 (
		\desIn[55]_pad ,
		\roundSel[4]_pad ,
		\roundSel[5]_pad ,
		_w305_,
		_w1050_
	);
	LUT4 #(
		.INIT('h1011)
	) name746 (
		_w1049_,
		_w1050_,
		_w1047_,
		_w1048_,
		_w1051_
	);
	LUT4 #(
		.INIT('hefee)
	) name747 (
		_w1049_,
		_w1050_,
		_w1047_,
		_w1048_,
		_w1052_
	);
	LUT2 #(
		.INIT('h9)
	) name748 (
		_w1046_,
		_w1051_,
		_w1053_
	);
	LUT4 #(
		.INIT('h0200)
	) name749 (
		\desIn[39]_pad ,
		\roundSel[4]_pad ,
		\roundSel[5]_pad ,
		_w305_,
		_w1054_
	);
	LUT4 #(
		.INIT('h4155)
	) name750 (
		\FP_R_reg[5]/P0001 ,
		\roundSel[4]_pad ,
		\roundSel[5]_pad ,
		_w305_,
		_w1055_
	);
	LUT4 #(
		.INIT('he8ff)
	) name751 (
		\FP_R_reg[37]/NET0131 ,
		\roundSel[4]_pad ,
		\roundSel[5]_pad ,
		_w305_,
		_w1056_
	);
	LUT3 #(
		.INIT('h45)
	) name752 (
		_w1054_,
		_w1055_,
		_w1056_,
		_w1057_
	);
	LUT3 #(
		.INIT('hba)
	) name753 (
		_w1054_,
		_w1055_,
		_w1056_,
		_w1058_
	);
	LUT3 #(
		.INIT('ha8)
	) name754 (
		_w419_,
		_w690_,
		_w739_,
		_w1059_
	);
	LUT3 #(
		.INIT('ha8)
	) name755 (
		_w406_,
		_w703_,
		_w721_,
		_w1060_
	);
	LUT3 #(
		.INIT('ha8)
	) name756 (
		_w415_,
		_w702_,
		_w734_,
		_w1061_
	);
	LUT3 #(
		.INIT('ha8)
	) name757 (
		_w312_,
		_w700_,
		_w730_,
		_w1062_
	);
	LUT4 #(
		.INIT('h0001)
	) name758 (
		_w1059_,
		_w1060_,
		_w1061_,
		_w1062_,
		_w1063_
	);
	LUT3 #(
		.INIT('ha8)
	) name759 (
		_w377_,
		_w708_,
		_w737_,
		_w1064_
	);
	LUT3 #(
		.INIT('ha8)
	) name760 (
		_w323_,
		_w712_,
		_w671_,
		_w1065_
	);
	LUT3 #(
		.INIT('ha8)
	) name761 (
		_w398_,
		_w752_,
		_w725_,
		_w1066_
	);
	LUT3 #(
		.INIT('ha8)
	) name762 (
		_w373_,
		_w756_,
		_w758_,
		_w1067_
	);
	LUT4 #(
		.INIT('h0001)
	) name763 (
		_w1064_,
		_w1065_,
		_w1066_,
		_w1067_,
		_w1068_
	);
	LUT3 #(
		.INIT('ha8)
	) name764 (
		_w343_,
		_w717_,
		_w750_,
		_w1069_
	);
	LUT3 #(
		.INIT('ha8)
	) name765 (
		_w402_,
		_w696_,
		_w831_,
		_w1070_
	);
	LUT3 #(
		.INIT('ha8)
	) name766 (
		_w388_,
		_w681_,
		_w759_,
		_w1071_
	);
	LUT3 #(
		.INIT('ha8)
	) name767 (
		_w423_,
		_w669_,
		_w755_,
		_w1072_
	);
	LUT4 #(
		.INIT('h0001)
	) name768 (
		_w1069_,
		_w1070_,
		_w1071_,
		_w1072_,
		_w1073_
	);
	LUT3 #(
		.INIT('ha8)
	) name769 (
		_w333_,
		_w672_,
		_w746_,
		_w1074_
	);
	LUT3 #(
		.INIT('ha8)
	) name770 (
		_w411_,
		_w665_,
		_w740_,
		_w1075_
	);
	LUT3 #(
		.INIT('ha8)
	) name771 (
		_w305_,
		_w724_,
		_w849_,
		_w1076_
	);
	LUT3 #(
		.INIT('ha8)
	) name772 (
		_w363_,
		_w677_,
		_w753_,
		_w1077_
	);
	LUT4 #(
		.INIT('h0001)
	) name773 (
		_w1074_,
		_w1075_,
		_w1076_,
		_w1077_,
		_w1078_
	);
	LUT4 #(
		.INIT('h8000)
	) name774 (
		_w1073_,
		_w1078_,
		_w1063_,
		_w1068_,
		_w1079_
	);
	LUT2 #(
		.INIT('h6)
	) name775 (
		_w1057_,
		_w1079_,
		_w1080_
	);
	LUT4 #(
		.INIT('h0200)
	) name776 (
		\desIn[5]_pad ,
		\roundSel[4]_pad ,
		\roundSel[5]_pad ,
		_w305_,
		_w1081_
	);
	LUT4 #(
		.INIT('h4155)
	) name777 (
		\FP_R_reg[9]/P0001 ,
		\roundSel[4]_pad ,
		\roundSel[5]_pad ,
		_w305_,
		_w1082_
	);
	LUT4 #(
		.INIT('he8ff)
	) name778 (
		\FP_R_reg[41]/NET0131 ,
		\roundSel[4]_pad ,
		\roundSel[5]_pad ,
		_w305_,
		_w1083_
	);
	LUT3 #(
		.INIT('h45)
	) name779 (
		_w1081_,
		_w1082_,
		_w1083_,
		_w1084_
	);
	LUT3 #(
		.INIT('hba)
	) name780 (
		_w1081_,
		_w1082_,
		_w1083_,
		_w1085_
	);
	LUT3 #(
		.INIT('ha8)
	) name781 (
		_w377_,
		_w734_,
		_w767_,
		_w1086_
	);
	LUT3 #(
		.INIT('ha8)
	) name782 (
		_w312_,
		_w712_,
		_w802_,
		_w1087_
	);
	LUT3 #(
		.INIT('ha8)
	) name783 (
		_w323_,
		_w700_,
		_w797_,
		_w1088_
	);
	LUT3 #(
		.INIT('ha8)
	) name784 (
		_w333_,
		_w847_,
		_w831_,
		_w1089_
	);
	LUT4 #(
		.INIT('h0001)
	) name785 (
		_w1086_,
		_w1087_,
		_w1088_,
		_w1089_,
		_w1090_
	);
	LUT3 #(
		.INIT('ha8)
	) name786 (
		_w305_,
		_w669_,
		_w811_,
		_w1091_
	);
	LUT3 #(
		.INIT('ha8)
	) name787 (
		_w343_,
		_w824_,
		_w858_,
		_w1092_
	);
	LUT3 #(
		.INIT('ha8)
	) name788 (
		_w388_,
		_w856_,
		_w842_,
		_w1093_
	);
	LUT3 #(
		.INIT('ha8)
	) name789 (
		_w415_,
		_w737_,
		_w786_,
		_w1094_
	);
	LUT4 #(
		.INIT('h0001)
	) name790 (
		_w1091_,
		_w1092_,
		_w1093_,
		_w1094_,
		_w1095_
	);
	LUT3 #(
		.INIT('ha8)
	) name791 (
		_w423_,
		_w868_,
		_w849_,
		_w1096_
	);
	LUT3 #(
		.INIT('ha8)
	) name792 (
		_w419_,
		_w753_,
		_w774_,
		_w1097_
	);
	LUT3 #(
		.INIT('ha8)
	) name793 (
		_w373_,
		_w860_,
		_w837_,
		_w1098_
	);
	LUT3 #(
		.INIT('ha8)
	) name794 (
		_w398_,
		_w740_,
		_w806_,
		_w1099_
	);
	LUT4 #(
		.INIT('h0001)
	) name795 (
		_w1096_,
		_w1097_,
		_w1098_,
		_w1099_,
		_w1100_
	);
	LUT3 #(
		.INIT('ha8)
	) name796 (
		_w411_,
		_w725_,
		_w772_,
		_w1101_
	);
	LUT3 #(
		.INIT('ha8)
	) name797 (
		_w406_,
		_w865_,
		_w863_,
		_w1102_
	);
	LUT3 #(
		.INIT('ha8)
	) name798 (
		_w402_,
		_w672_,
		_w779_,
		_w1103_
	);
	LUT3 #(
		.INIT('ha8)
	) name799 (
		_w363_,
		_w690_,
		_w788_,
		_w1104_
	);
	LUT4 #(
		.INIT('h0001)
	) name800 (
		_w1101_,
		_w1102_,
		_w1103_,
		_w1104_,
		_w1105_
	);
	LUT4 #(
		.INIT('h8000)
	) name801 (
		_w1100_,
		_w1105_,
		_w1090_,
		_w1095_,
		_w1106_
	);
	LUT2 #(
		.INIT('h6)
	) name802 (
		_w1084_,
		_w1106_,
		_w1107_
	);
	LUT4 #(
		.INIT('h0200)
	) name803 (
		\desIn[31]_pad ,
		\roundSel[4]_pad ,
		\roundSel[5]_pad ,
		_w305_,
		_w1108_
	);
	LUT4 #(
		.INIT('h4155)
	) name804 (
		\FP_R_reg[4]/P0001 ,
		\roundSel[4]_pad ,
		\roundSel[5]_pad ,
		_w305_,
		_w1109_
	);
	LUT4 #(
		.INIT('he8ff)
	) name805 (
		\FP_R_reg[36]/NET0131 ,
		\roundSel[4]_pad ,
		\roundSel[5]_pad ,
		_w305_,
		_w1110_
	);
	LUT3 #(
		.INIT('h45)
	) name806 (
		_w1108_,
		_w1109_,
		_w1110_,
		_w1111_
	);
	LUT3 #(
		.INIT('hba)
	) name807 (
		_w1108_,
		_w1109_,
		_w1110_,
		_w1112_
	);
	LUT3 #(
		.INIT('ha8)
	) name808 (
		_w377_,
		_w665_,
		_w837_,
		_w1113_
	);
	LUT3 #(
		.INIT('ha8)
	) name809 (
		_w343_,
		_w774_,
		_w811_,
		_w1114_
	);
	LUT3 #(
		.INIT('ha8)
	) name810 (
		_w415_,
		_w724_,
		_w788_,
		_w1115_
	);
	LUT3 #(
		.INIT('ha8)
	) name811 (
		_w398_,
		_w730_,
		_w863_,
		_w1116_
	);
	LUT4 #(
		.INIT('h0001)
	) name812 (
		_w1113_,
		_w1114_,
		_w1115_,
		_w1116_,
		_w1117_
	);
	LUT3 #(
		.INIT('ha8)
	) name813 (
		_w305_,
		_w702_,
		_w824_,
		_w1118_
	);
	LUT3 #(
		.INIT('ha8)
	) name814 (
		_w333_,
		_w686_,
		_w772_,
		_w1119_
	);
	LUT3 #(
		.INIT('ha8)
	) name815 (
		_w373_,
		_w767_,
		_w779_,
		_w1120_
	);
	LUT3 #(
		.INIT('ha8)
	) name816 (
		_w388_,
		_w802_,
		_w793_,
		_w1121_
	);
	LUT4 #(
		.INIT('h0001)
	) name817 (
		_w1118_,
		_w1119_,
		_w1120_,
		_w1121_,
		_w1122_
	);
	LUT3 #(
		.INIT('ha8)
	) name818 (
		_w423_,
		_w736_,
		_w797_,
		_w1123_
	);
	LUT3 #(
		.INIT('ha8)
	) name819 (
		_w402_,
		_w677_,
		_w860_,
		_w1124_
	);
	LUT3 #(
		.INIT('ha8)
	) name820 (
		_w411_,
		_w708_,
		_w847_,
		_w1125_
	);
	LUT3 #(
		.INIT('ha8)
	) name821 (
		_w323_,
		_w739_,
		_w868_,
		_w1126_
	);
	LUT4 #(
		.INIT('h0001)
	) name822 (
		_w1123_,
		_w1124_,
		_w1125_,
		_w1126_,
		_w1127_
	);
	LUT3 #(
		.INIT('ha8)
	) name823 (
		_w406_,
		_w809_,
		_w806_,
		_w1128_
	);
	LUT3 #(
		.INIT('ha8)
	) name824 (
		_w363_,
		_w696_,
		_w786_,
		_w1129_
	);
	LUT3 #(
		.INIT('ha8)
	) name825 (
		_w419_,
		_w671_,
		_w858_,
		_w1130_
	);
	LUT3 #(
		.INIT('ha8)
	) name826 (
		_w312_,
		_w752_,
		_w842_,
		_w1131_
	);
	LUT4 #(
		.INIT('h0001)
	) name827 (
		_w1128_,
		_w1129_,
		_w1130_,
		_w1131_,
		_w1132_
	);
	LUT4 #(
		.INIT('h8000)
	) name828 (
		_w1127_,
		_w1132_,
		_w1117_,
		_w1122_,
		_w1133_
	);
	LUT2 #(
		.INIT('h9)
	) name829 (
		_w1111_,
		_w1133_,
		_w1134_
	);
	LUT4 #(
		.INIT('h0990)
	) name830 (
		_w1084_,
		_w1106_,
		_w1111_,
		_w1133_,
		_w1135_
	);
	LUT4 #(
		.INIT('h0200)
	) name831 (
		\desIn[47]_pad ,
		\roundSel[4]_pad ,
		\roundSel[5]_pad ,
		_w305_,
		_w1136_
	);
	LUT4 #(
		.INIT('h4155)
	) name832 (
		\FP_R_reg[6]/P0001 ,
		\roundSel[4]_pad ,
		\roundSel[5]_pad ,
		_w305_,
		_w1137_
	);
	LUT4 #(
		.INIT('he8ff)
	) name833 (
		\FP_R_reg[38]/NET0131 ,
		\roundSel[4]_pad ,
		\roundSel[5]_pad ,
		_w305_,
		_w1138_
	);
	LUT3 #(
		.INIT('h45)
	) name834 (
		_w1136_,
		_w1137_,
		_w1138_,
		_w1139_
	);
	LUT3 #(
		.INIT('hba)
	) name835 (
		_w1136_,
		_w1137_,
		_w1138_,
		_w1140_
	);
	LUT3 #(
		.INIT('ha8)
	) name836 (
		_w419_,
		_w730_,
		_w831_,
		_w1141_
	);
	LUT3 #(
		.INIT('ha8)
	) name837 (
		_w423_,
		_w721_,
		_w734_,
		_w1142_
	);
	LUT3 #(
		.INIT('ha8)
	) name838 (
		_w398_,
		_w671_,
		_w737_,
		_w1143_
	);
	LUT3 #(
		.INIT('ha8)
	) name839 (
		_w363_,
		_w712_,
		_w746_,
		_w1144_
	);
	LUT4 #(
		.INIT('h0001)
	) name840 (
		_w1141_,
		_w1142_,
		_w1143_,
		_w1144_,
		_w1145_
	);
	LUT3 #(
		.INIT('ha8)
	) name841 (
		_w305_,
		_w708_,
		_w865_,
		_w1146_
	);
	LUT3 #(
		.INIT('ha8)
	) name842 (
		_w323_,
		_w677_,
		_w725_,
		_w1147_
	);
	LUT3 #(
		.INIT('ha8)
	) name843 (
		_w333_,
		_w753_,
		_w759_,
		_w1148_
	);
	LUT3 #(
		.INIT('ha8)
	) name844 (
		_w312_,
		_w665_,
		_w690_,
		_w1149_
	);
	LUT4 #(
		.INIT('h0001)
	) name845 (
		_w1146_,
		_w1147_,
		_w1148_,
		_w1149_,
		_w1150_
	);
	LUT3 #(
		.INIT('ha8)
	) name846 (
		_w388_,
		_w717_,
		_w672_,
		_w1151_
	);
	LUT3 #(
		.INIT('ha8)
	) name847 (
		_w377_,
		_w752_,
		_w849_,
		_w1152_
	);
	LUT3 #(
		.INIT('ha8)
	) name848 (
		_w415_,
		_w755_,
		_w740_,
		_w1153_
	);
	LUT3 #(
		.INIT('ha8)
	) name849 (
		_w373_,
		_w703_,
		_w750_,
		_w1154_
	);
	LUT4 #(
		.INIT('h0001)
	) name850 (
		_w1151_,
		_w1152_,
		_w1153_,
		_w1154_,
		_w1155_
	);
	LUT3 #(
		.INIT('ha8)
	) name851 (
		_w406_,
		_w669_,
		_w758_,
		_w1156_
	);
	LUT3 #(
		.INIT('ha8)
	) name852 (
		_w411_,
		_w700_,
		_w702_,
		_w1157_
	);
	LUT3 #(
		.INIT('ha8)
	) name853 (
		_w402_,
		_w739_,
		_w856_,
		_w1158_
	);
	LUT3 #(
		.INIT('ha8)
	) name854 (
		_w343_,
		_w681_,
		_w756_,
		_w1159_
	);
	LUT4 #(
		.INIT('h0001)
	) name855 (
		_w1156_,
		_w1157_,
		_w1158_,
		_w1159_,
		_w1160_
	);
	LUT4 #(
		.INIT('h8000)
	) name856 (
		_w1155_,
		_w1160_,
		_w1145_,
		_w1150_,
		_w1161_
	);
	LUT2 #(
		.INIT('h9)
	) name857 (
		_w1139_,
		_w1161_,
		_w1162_
	);
	LUT4 #(
		.INIT('h9009)
	) name858 (
		_w1139_,
		_w1161_,
		_w1111_,
		_w1133_,
		_w1163_
	);
	LUT4 #(
		.INIT('h20fd)
	) name859 (
		_w1080_,
		_w1107_,
		_w1134_,
		_w1163_,
		_w1164_
	);
	LUT2 #(
		.INIT('h1)
	) name860 (
		_w1053_,
		_w1164_,
		_w1165_
	);
	LUT4 #(
		.INIT('h0990)
	) name861 (
		_w1057_,
		_w1079_,
		_w1084_,
		_w1106_,
		_w1166_
	);
	LUT4 #(
		.INIT('h5410)
	) name862 (
		_w1162_,
		_w1080_,
		_w1107_,
		_w1135_,
		_w1167_
	);
	LUT4 #(
		.INIT('h0990)
	) name863 (
		_w1139_,
		_w1161_,
		_w1057_,
		_w1079_,
		_w1168_
	);
	LUT4 #(
		.INIT('h9009)
	) name864 (
		_w1084_,
		_w1106_,
		_w1111_,
		_w1133_,
		_w1169_
	);
	LUT3 #(
		.INIT('h80)
	) name865 (
		_w1053_,
		_w1168_,
		_w1169_,
		_w1170_
	);
	LUT4 #(
		.INIT('h0660)
	) name866 (
		_w1139_,
		_w1161_,
		_w1057_,
		_w1079_,
		_w1171_
	);
	LUT4 #(
		.INIT('h0990)
	) name867 (
		_w1084_,
		_w1106_,
		_w1046_,
		_w1051_,
		_w1172_
	);
	LUT4 #(
		.INIT('h9bdf)
	) name868 (
		_w1162_,
		_w1080_,
		_w1135_,
		_w1172_,
		_w1173_
	);
	LUT3 #(
		.INIT('h10)
	) name869 (
		_w1167_,
		_w1170_,
		_w1173_,
		_w1174_
	);
	LUT3 #(
		.INIT('h8a)
	) name870 (
		_w1025_,
		_w1165_,
		_w1174_,
		_w1175_
	);
	LUT4 #(
		.INIT('h9009)
	) name871 (
		_w1057_,
		_w1079_,
		_w1111_,
		_w1133_,
		_w1176_
	);
	LUT4 #(
		.INIT('h6006)
	) name872 (
		_w1139_,
		_w1161_,
		_w1057_,
		_w1079_,
		_w1177_
	);
	LUT3 #(
		.INIT('ha8)
	) name873 (
		_w1053_,
		_w1176_,
		_w1177_,
		_w1178_
	);
	LUT4 #(
		.INIT('h6006)
	) name874 (
		_w1084_,
		_w1106_,
		_w1111_,
		_w1133_,
		_w1179_
	);
	LUT4 #(
		.INIT('h9009)
	) name875 (
		_w1057_,
		_w1079_,
		_w1084_,
		_w1106_,
		_w1180_
	);
	LUT4 #(
		.INIT('h4100)
	) name876 (
		_w1162_,
		_w1080_,
		_w1107_,
		_w1134_,
		_w1181_
	);
	LUT3 #(
		.INIT('h54)
	) name877 (
		_w1025_,
		_w1178_,
		_w1181_,
		_w1182_
	);
	LUT3 #(
		.INIT('h20)
	) name878 (
		_w1107_,
		_w1134_,
		_w1168_,
		_w1183_
	);
	LUT3 #(
		.INIT('h8c)
	) name879 (
		_w1162_,
		_w1053_,
		_w1176_,
		_w1184_
	);
	LUT4 #(
		.INIT('h009f)
	) name880 (
		_w1162_,
		_w1080_,
		_w1135_,
		_w1053_,
		_w1185_
	);
	LUT3 #(
		.INIT('h0b)
	) name881 (
		_w1183_,
		_w1184_,
		_w1185_,
		_w1186_
	);
	LUT4 #(
		.INIT('h0660)
	) name882 (
		_w1084_,
		_w1106_,
		_w1111_,
		_w1133_,
		_w1187_
	);
	LUT3 #(
		.INIT('h9d)
	) name883 (
		_w1107_,
		_w1134_,
		_w1168_,
		_w1188_
	);
	LUT4 #(
		.INIT('h0990)
	) name884 (
		_w1002_,
		_w1024_,
		_w1046_,
		_w1051_,
		_w1189_
	);
	LUT2 #(
		.INIT('h4)
	) name885 (
		_w1177_,
		_w1189_,
		_w1190_
	);
	LUT2 #(
		.INIT('h4)
	) name886 (
		_w1188_,
		_w1190_,
		_w1191_
	);
	LUT3 #(
		.INIT('h01)
	) name887 (
		_w1182_,
		_w1186_,
		_w1191_,
		_w1192_
	);
	LUT4 #(
		.INIT('h0100)
	) name888 (
		\desIn[14]_pad ,
		\roundSel[4]_pad ,
		\roundSel[5]_pad ,
		_w305_,
		_w1193_
	);
	LUT4 #(
		.INIT('h2800)
	) name889 (
		\FP_R_reg[2]/P0001 ,
		\roundSel[4]_pad ,
		\roundSel[5]_pad ,
		_w305_,
		_w1194_
	);
	LUT4 #(
		.INIT('h7c55)
	) name890 (
		\FP_R_reg[34]/NET0131 ,
		\roundSel[4]_pad ,
		\roundSel[5]_pad ,
		_w305_,
		_w1195_
	);
	LUT3 #(
		.INIT('h45)
	) name891 (
		_w1193_,
		_w1194_,
		_w1195_,
		_w1196_
	);
	LUT3 #(
		.INIT('h4b)
	) name892 (
		_w1175_,
		_w1192_,
		_w1196_,
		_w1197_
	);
	LUT3 #(
		.INIT('h40)
	) name893 (
		\FP_R_reg[34]/NET0131 ,
		_w305_,
		_w307_,
		_w1198_
	);
	LUT4 #(
		.INIT('hb0aa)
	) name894 (
		\FP_R_reg[2]/P0001 ,
		\roundSel[4]_pad ,
		\roundSel[5]_pad ,
		_w305_,
		_w1199_
	);
	LUT4 #(
		.INIT('h0800)
	) name895 (
		\FP_R_reg[34]/NET0131 ,
		\roundSel[4]_pad ,
		\roundSel[5]_pad ,
		_w305_,
		_w1200_
	);
	LUT4 #(
		.INIT('h0200)
	) name896 (
		\desIn[15]_pad ,
		\roundSel[4]_pad ,
		\roundSel[5]_pad ,
		_w305_,
		_w1201_
	);
	LUT4 #(
		.INIT('h1011)
	) name897 (
		_w1200_,
		_w1201_,
		_w1198_,
		_w1199_,
		_w1202_
	);
	LUT4 #(
		.INIT('hefee)
	) name898 (
		_w1200_,
		_w1201_,
		_w1198_,
		_w1199_,
		_w1203_
	);
	LUT4 #(
		.INIT('h0200)
	) name899 (
		\desIn[51]_pad ,
		\roundSel[4]_pad ,
		\roundSel[5]_pad ,
		_w305_,
		_w1204_
	);
	LUT4 #(
		.INIT('h4155)
	) name900 (
		\FP_R_reg[23]/P0001 ,
		\roundSel[4]_pad ,
		\roundSel[5]_pad ,
		_w305_,
		_w1205_
	);
	LUT4 #(
		.INIT('he8ff)
	) name901 (
		\FP_R_reg[55]/NET0131 ,
		\roundSel[4]_pad ,
		\roundSel[5]_pad ,
		_w305_,
		_w1206_
	);
	LUT3 #(
		.INIT('h45)
	) name902 (
		_w1204_,
		_w1205_,
		_w1206_,
		_w1207_
	);
	LUT3 #(
		.INIT('hba)
	) name903 (
		_w1204_,
		_w1205_,
		_w1206_,
		_w1208_
	);
	LUT3 #(
		.INIT('hc8)
	) name904 (
		_w327_,
		_w333_,
		_w347_,
		_w1209_
	);
	LUT3 #(
		.INIT('ha8)
	) name905 (
		_w363_,
		_w392_,
		_w399_,
		_w1210_
	);
	LUT3 #(
		.INIT('ha8)
	) name906 (
		_w411_,
		_w420_,
		_w425_,
		_w1211_
	);
	LUT3 #(
		.INIT('he0)
	) name907 (
		_w357_,
		_w371_,
		_w398_,
		_w1212_
	);
	LUT4 #(
		.INIT('h0001)
	) name908 (
		_w1209_,
		_w1210_,
		_w1211_,
		_w1212_,
		_w1213_
	);
	LUT3 #(
		.INIT('hc8)
	) name909 (
		_w413_,
		_w419_,
		_w440_,
		_w1214_
	);
	LUT3 #(
		.INIT('he0)
	) name910 (
		_w351_,
		_w416_,
		_w406_,
		_w1215_
	);
	LUT3 #(
		.INIT('hc8)
	) name911 (
		_w317_,
		_w415_,
		_w408_,
		_w1216_
	);
	LUT3 #(
		.INIT('hc8)
	) name912 (
		_w321_,
		_w402_,
		_w459_,
		_w1217_
	);
	LUT4 #(
		.INIT('h0001)
	) name913 (
		_w1214_,
		_w1215_,
		_w1216_,
		_w1217_,
		_w1218_
	);
	LUT3 #(
		.INIT('he0)
	) name914 (
		_w375_,
		_w412_,
		_w423_,
		_w1219_
	);
	LUT3 #(
		.INIT('hc8)
	) name915 (
		_w381_,
		_w323_,
		_w341_,
		_w1220_
	);
	LUT3 #(
		.INIT('ha8)
	) name916 (
		_w377_,
		_w331_,
		_w460_,
		_w1221_
	);
	LUT3 #(
		.INIT('he0)
	) name917 (
		_w367_,
		_w374_,
		_w388_,
		_w1222_
	);
	LUT4 #(
		.INIT('h0001)
	) name918 (
		_w1219_,
		_w1220_,
		_w1221_,
		_w1222_,
		_w1223_
	);
	LUT3 #(
		.INIT('ha8)
	) name919 (
		_w312_,
		_w417_,
		_w403_,
		_w1224_
	);
	LUT3 #(
		.INIT('ha8)
	) name920 (
		_w305_,
		_w400_,
		_w444_,
		_w1225_
	);
	LUT3 #(
		.INIT('hc8)
	) name921 (
		_w337_,
		_w343_,
		_w407_,
		_w1226_
	);
	LUT3 #(
		.INIT('ha8)
	) name922 (
		_w373_,
		_w424_,
		_w396_,
		_w1227_
	);
	LUT4 #(
		.INIT('h0001)
	) name923 (
		_w1224_,
		_w1225_,
		_w1226_,
		_w1227_,
		_w1228_
	);
	LUT4 #(
		.INIT('h8000)
	) name924 (
		_w1223_,
		_w1228_,
		_w1213_,
		_w1218_,
		_w1229_
	);
	LUT2 #(
		.INIT('h9)
	) name925 (
		_w1207_,
		_w1229_,
		_w1230_
	);
	LUT3 #(
		.INIT('ha8)
	) name926 (
		_w377_,
		_w420_,
		_w539_,
		_w1231_
	);
	LUT3 #(
		.INIT('ha8)
	) name927 (
		_w333_,
		_w449_,
		_w483_,
		_w1232_
	);
	LUT3 #(
		.INIT('ha8)
	) name928 (
		_w323_,
		_w440_,
		_w561_,
		_w1233_
	);
	LUT3 #(
		.INIT('ha8)
	) name929 (
		_w363_,
		_w459_,
		_w435_,
		_w1234_
	);
	LUT4 #(
		.INIT('h0001)
	) name930 (
		_w1231_,
		_w1232_,
		_w1233_,
		_w1234_,
		_w1235_
	);
	LUT3 #(
		.INIT('ha8)
	) name931 (
		_w305_,
		_w317_,
		_w404_,
		_w1236_
	);
	LUT3 #(
		.INIT('ha8)
	) name932 (
		_w388_,
		_w492_,
		_w471_,
		_w1237_
	);
	LUT3 #(
		.INIT('ha8)
	) name933 (
		_w411_,
		_w460_,
		_w553_,
		_w1238_
	);
	LUT3 #(
		.INIT('he0)
	) name934 (
		_w361_,
		_w399_,
		_w402_,
		_w1239_
	);
	LUT4 #(
		.INIT('h0001)
	) name935 (
		_w1236_,
		_w1237_,
		_w1238_,
		_w1239_,
		_w1240_
	);
	LUT3 #(
		.INIT('hc8)
	) name936 (
		_w381_,
		_w419_,
		_w559_,
		_w1241_
	);
	LUT3 #(
		.INIT('ha8)
	) name937 (
		_w373_,
		_w457_,
		_w490_,
		_w1242_
	);
	LUT3 #(
		.INIT('ha8)
	) name938 (
		_w343_,
		_w455_,
		_w488_,
		_w1243_
	);
	LUT3 #(
		.INIT('ha8)
	) name939 (
		_w423_,
		_w465_,
		_w480_,
		_w1244_
	);
	LUT4 #(
		.INIT('h0001)
	) name940 (
		_w1241_,
		_w1242_,
		_w1243_,
		_w1244_,
		_w1245_
	);
	LUT3 #(
		.INIT('ha8)
	) name941 (
		_w406_,
		_w473_,
		_w478_,
		_w1246_
	);
	LUT3 #(
		.INIT('hc8)
	) name942 (
		_w357_,
		_w312_,
		_w556_,
		_w1247_
	);
	LUT3 #(
		.INIT('ha8)
	) name943 (
		_w415_,
		_w433_,
		_w444_,
		_w1248_
	);
	LUT3 #(
		.INIT('ha8)
	) name944 (
		_w398_,
		_w403_,
		_w548_,
		_w1249_
	);
	LUT4 #(
		.INIT('h0001)
	) name945 (
		_w1246_,
		_w1247_,
		_w1248_,
		_w1249_,
		_w1250_
	);
	LUT4 #(
		.INIT('h8000)
	) name946 (
		_w1245_,
		_w1250_,
		_w1235_,
		_w1240_,
		_w1251_
	);
	LUT4 #(
		.INIT('h0200)
	) name947 (
		\desIn[1]_pad ,
		\roundSel[4]_pad ,
		\roundSel[5]_pad ,
		_w305_,
		_w1252_
	);
	LUT4 #(
		.INIT('h4155)
	) name948 (
		\FP_R_reg[25]/P0001 ,
		\roundSel[4]_pad ,
		\roundSel[5]_pad ,
		_w305_,
		_w1253_
	);
	LUT4 #(
		.INIT('he8ff)
	) name949 (
		\FP_R_reg[57]/NET0131 ,
		\roundSel[4]_pad ,
		\roundSel[5]_pad ,
		_w305_,
		_w1254_
	);
	LUT3 #(
		.INIT('h45)
	) name950 (
		_w1252_,
		_w1253_,
		_w1254_,
		_w1255_
	);
	LUT3 #(
		.INIT('hba)
	) name951 (
		_w1252_,
		_w1253_,
		_w1254_,
		_w1256_
	);
	LUT2 #(
		.INIT('h9)
	) name952 (
		_w1251_,
		_w1255_,
		_w1257_
	);
	LUT3 #(
		.INIT('hc8)
	) name953 (
		_w371_,
		_w377_,
		_w444_,
		_w1258_
	);
	LUT3 #(
		.INIT('hc8)
	) name954 (
		_w367_,
		_w343_,
		_w424_,
		_w1259_
	);
	LUT3 #(
		.INIT('hc8)
	) name955 (
		_w413_,
		_w402_,
		_w483_,
		_w1260_
	);
	LUT3 #(
		.INIT('ha8)
	) name956 (
		_w305_,
		_w331_,
		_w465_,
		_w1261_
	);
	LUT4 #(
		.INIT('h0001)
	) name957 (
		_w1258_,
		_w1259_,
		_w1260_,
		_w1261_,
		_w1262_
	);
	LUT3 #(
		.INIT('hc8)
	) name958 (
		_w357_,
		_w323_,
		_w392_,
		_w1263_
	);
	LUT3 #(
		.INIT('ha8)
	) name959 (
		_w363_,
		_w381_,
		_w347_,
		_w1264_
	);
	LUT3 #(
		.INIT('ha8)
	) name960 (
		_w411_,
		_w403_,
		_w408_,
		_w1265_
	);
	LUT3 #(
		.INIT('he0)
	) name961 (
		_w317_,
		_w351_,
		_w423_,
		_w1266_
	);
	LUT4 #(
		.INIT('h0001)
	) name962 (
		_w1263_,
		_w1264_,
		_w1265_,
		_w1266_,
		_w1267_
	);
	LUT3 #(
		.INIT('hc8)
	) name963 (
		_w327_,
		_w388_,
		_w407_,
		_w1268_
	);
	LUT3 #(
		.INIT('hc8)
	) name964 (
		_w374_,
		_w333_,
		_w399_,
		_w1269_
	);
	LUT3 #(
		.INIT('hc8)
	) name965 (
		_w417_,
		_w419_,
		_w459_,
		_w1270_
	);
	LUT3 #(
		.INIT('hc8)
	) name966 (
		_w341_,
		_w398_,
		_w460_,
		_w1271_
	);
	LUT4 #(
		.INIT('h0001)
	) name967 (
		_w1268_,
		_w1269_,
		_w1270_,
		_w1271_,
		_w1272_
	);
	LUT3 #(
		.INIT('ha8)
	) name968 (
		_w312_,
		_w425_,
		_w440_,
		_w1273_
	);
	LUT3 #(
		.INIT('ha8)
	) name969 (
		_w373_,
		_w337_,
		_w416_,
		_w1274_
	);
	LUT3 #(
		.INIT('he0)
	) name970 (
		_w412_,
		_w396_,
		_w406_,
		_w1275_
	);
	LUT3 #(
		.INIT('hc8)
	) name971 (
		_w375_,
		_w415_,
		_w420_,
		_w1276_
	);
	LUT4 #(
		.INIT('h0001)
	) name972 (
		_w1273_,
		_w1274_,
		_w1275_,
		_w1276_,
		_w1277_
	);
	LUT4 #(
		.INIT('h8000)
	) name973 (
		_w1272_,
		_w1277_,
		_w1262_,
		_w1267_,
		_w1278_
	);
	LUT2 #(
		.INIT('h9)
	) name974 (
		_w310_,
		_w1278_,
		_w1279_
	);
	LUT3 #(
		.INIT('hc8)
	) name975 (
		_w361_,
		_w343_,
		_w421_,
		_w1280_
	);
	LUT3 #(
		.INIT('hc8)
	) name976 (
		_w331_,
		_w423_,
		_w548_,
		_w1281_
	);
	LUT3 #(
		.INIT('ha8)
	) name977 (
		_w363_,
		_w417_,
		_w553_,
		_w1282_
	);
	LUT3 #(
		.INIT('ha8)
	) name978 (
		_w305_,
		_w351_,
		_w457_,
		_w1283_
	);
	LUT4 #(
		.INIT('h0001)
	) name979 (
		_w1280_,
		_w1281_,
		_w1282_,
		_w1283_,
		_w1284_
	);
	LUT3 #(
		.INIT('hc8)
	) name980 (
		_w375_,
		_w377_,
		_w473_,
		_w1285_
	);
	LUT3 #(
		.INIT('hc8)
	) name981 (
		_w374_,
		_w402_,
		_w455_,
		_w1286_
	);
	LUT3 #(
		.INIT('ha8)
	) name982 (
		_w373_,
		_w385_,
		_w404_,
		_w1287_
	);
	LUT3 #(
		.INIT('ha8)
	) name983 (
		_w333_,
		_w413_,
		_w556_,
		_w1288_
	);
	LUT4 #(
		.INIT('h0001)
	) name984 (
		_w1285_,
		_w1286_,
		_w1287_,
		_w1288_,
		_w1289_
	);
	LUT3 #(
		.INIT('hc8)
	) name985 (
		_w371_,
		_w415_,
		_w561_,
		_w1290_
	);
	LUT3 #(
		.INIT('hc8)
	) name986 (
		_w400_,
		_w406_,
		_w539_,
		_w1291_
	);
	LUT3 #(
		.INIT('hc8)
	) name987 (
		_w321_,
		_w388_,
		_w559_,
		_w1292_
	);
	LUT3 #(
		.INIT('ha8)
	) name988 (
		_w312_,
		_w392_,
		_w449_,
		_w1293_
	);
	LUT4 #(
		.INIT('h0001)
	) name989 (
		_w1290_,
		_w1291_,
		_w1292_,
		_w1293_,
		_w1294_
	);
	LUT3 #(
		.INIT('hc8)
	) name990 (
		_w347_,
		_w419_,
		_w471_,
		_w1295_
	);
	LUT3 #(
		.INIT('ha8)
	) name991 (
		_w398_,
		_w408_,
		_w480_,
		_w1296_
	);
	LUT3 #(
		.INIT('hc8)
	) name992 (
		_w341_,
		_w411_,
		_w435_,
		_w1297_
	);
	LUT3 #(
		.INIT('ha8)
	) name993 (
		_w323_,
		_w425_,
		_w433_,
		_w1298_
	);
	LUT4 #(
		.INIT('h0001)
	) name994 (
		_w1295_,
		_w1296_,
		_w1297_,
		_w1298_,
		_w1299_
	);
	LUT4 #(
		.INIT('h8000)
	) name995 (
		_w1294_,
		_w1299_,
		_w1284_,
		_w1289_,
		_w1300_
	);
	LUT2 #(
		.INIT('h9)
	) name996 (
		_w568_,
		_w1300_,
		_w1301_
	);
	LUT4 #(
		.INIT('h4812)
	) name997 (
		_w310_,
		_w568_,
		_w1278_,
		_w1300_,
		_w1302_
	);
	LUT4 #(
		.INIT('h0660)
	) name998 (
		_w310_,
		_w1278_,
		_w1251_,
		_w1255_,
		_w1303_
	);
	LUT4 #(
		.INIT('h0041)
	) name999 (
		_w1279_,
		_w1301_,
		_w1257_,
		_w1230_,
		_w1304_
	);
	LUT3 #(
		.INIT('hc8)
	) name1000 (
		_w385_,
		_w333_,
		_w408_,
		_w1305_
	);
	LUT3 #(
		.INIT('ha8)
	) name1001 (
		_w419_,
		_w424_,
		_w561_,
		_w1306_
	);
	LUT3 #(
		.INIT('hc8)
	) name1002 (
		_w347_,
		_w415_,
		_w404_,
		_w1307_
	);
	LUT3 #(
		.INIT('hc8)
	) name1003 (
		_w371_,
		_w373_,
		_w413_,
		_w1308_
	);
	LUT4 #(
		.INIT('h0001)
	) name1004 (
		_w1305_,
		_w1306_,
		_w1307_,
		_w1308_,
		_w1309_
	);
	LUT3 #(
		.INIT('hc8)
	) name1005 (
		_w421_,
		_w423_,
		_w392_,
		_w1310_
	);
	LUT3 #(
		.INIT('hc8)
	) name1006 (
		_w416_,
		_w402_,
		_w435_,
		_w1311_
	);
	LUT3 #(
		.INIT('hc8)
	) name1007 (
		_w425_,
		_w388_,
		_w400_,
		_w1312_
	);
	LUT3 #(
		.INIT('hc8)
	) name1008 (
		_w396_,
		_w398_,
		_w556_,
		_w1313_
	);
	LUT4 #(
		.INIT('h0001)
	) name1009 (
		_w1310_,
		_w1311_,
		_w1312_,
		_w1313_,
		_w1314_
	);
	LUT3 #(
		.INIT('hc8)
	) name1010 (
		_w361_,
		_w363_,
		_w375_,
		_w1315_
	);
	LUT3 #(
		.INIT('ha8)
	) name1011 (
		_w377_,
		_w337_,
		_w553_,
		_w1316_
	);
	LUT3 #(
		.INIT('hc8)
	) name1012 (
		_w331_,
		_w343_,
		_w417_,
		_w1317_
	);
	LUT3 #(
		.INIT('he0)
	) name1013 (
		_w321_,
		_w341_,
		_w406_,
		_w1318_
	);
	LUT4 #(
		.INIT('h0001)
	) name1014 (
		_w1315_,
		_w1316_,
		_w1317_,
		_w1318_,
		_w1319_
	);
	LUT3 #(
		.INIT('ha8)
	) name1015 (
		_w312_,
		_w407_,
		_w548_,
		_w1320_
	);
	LUT3 #(
		.INIT('ha8)
	) name1016 (
		_w305_,
		_w367_,
		_w433_,
		_w1321_
	);
	LUT3 #(
		.INIT('hc8)
	) name1017 (
		_w374_,
		_w411_,
		_w539_,
		_w1322_
	);
	LUT3 #(
		.INIT('ha8)
	) name1018 (
		_w323_,
		_w351_,
		_w559_,
		_w1323_
	);
	LUT4 #(
		.INIT('h0001)
	) name1019 (
		_w1320_,
		_w1321_,
		_w1322_,
		_w1323_,
		_w1324_
	);
	LUT4 #(
		.INIT('h8000)
	) name1020 (
		_w1319_,
		_w1324_,
		_w1309_,
		_w1314_,
		_w1325_
	);
	LUT4 #(
		.INIT('h0200)
	) name1021 (
		\desIn[43]_pad ,
		\roundSel[4]_pad ,
		\roundSel[5]_pad ,
		_w305_,
		_w1326_
	);
	LUT4 #(
		.INIT('h4155)
	) name1022 (
		\FP_R_reg[22]/P0001 ,
		\roundSel[4]_pad ,
		\roundSel[5]_pad ,
		_w305_,
		_w1327_
	);
	LUT4 #(
		.INIT('he8ff)
	) name1023 (
		\FP_R_reg[54]/NET0131 ,
		\roundSel[4]_pad ,
		\roundSel[5]_pad ,
		_w305_,
		_w1328_
	);
	LUT3 #(
		.INIT('h45)
	) name1024 (
		_w1326_,
		_w1327_,
		_w1328_,
		_w1329_
	);
	LUT3 #(
		.INIT('hba)
	) name1025 (
		_w1326_,
		_w1327_,
		_w1328_,
		_w1330_
	);
	LUT2 #(
		.INIT('h9)
	) name1026 (
		_w1325_,
		_w1329_,
		_w1331_
	);
	LUT4 #(
		.INIT('h2814)
	) name1027 (
		_w568_,
		_w1325_,
		_w1329_,
		_w1300_,
		_w1332_
	);
	LUT4 #(
		.INIT('h7525)
	) name1028 (
		_w1279_,
		_w1331_,
		_w1301_,
		_w1257_,
		_w1333_
	);
	LUT4 #(
		.INIT('h9009)
	) name1029 (
		_w568_,
		_w1300_,
		_w1251_,
		_w1255_,
		_w1334_
	);
	LUT4 #(
		.INIT('h0200)
	) name1030 (
		\desIn[59]_pad ,
		\roundSel[4]_pad ,
		\roundSel[5]_pad ,
		_w305_,
		_w1335_
	);
	LUT4 #(
		.INIT('h4155)
	) name1031 (
		\FP_R_reg[24]/P0001 ,
		\roundSel[4]_pad ,
		\roundSel[5]_pad ,
		_w305_,
		_w1336_
	);
	LUT4 #(
		.INIT('he8ff)
	) name1032 (
		\FP_R_reg[56]/NET0131 ,
		\roundSel[4]_pad ,
		\roundSel[5]_pad ,
		_w305_,
		_w1337_
	);
	LUT3 #(
		.INIT('h45)
	) name1033 (
		_w1335_,
		_w1336_,
		_w1337_,
		_w1338_
	);
	LUT3 #(
		.INIT('hba)
	) name1034 (
		_w1335_,
		_w1336_,
		_w1337_,
		_w1339_
	);
	LUT3 #(
		.INIT('ha8)
	) name1035 (
		_w377_,
		_w403_,
		_w404_,
		_w1340_
	);
	LUT3 #(
		.INIT('ha8)
	) name1036 (
		_w415_,
		_w465_,
		_w553_,
		_w1341_
	);
	LUT3 #(
		.INIT('ha8)
	) name1037 (
		_w411_,
		_w444_,
		_w556_,
		_w1342_
	);
	LUT3 #(
		.INIT('he0)
	) name1038 (
		_w357_,
		_w361_,
		_w419_,
		_w1343_
	);
	LUT4 #(
		.INIT('h0001)
	) name1039 (
		_w1340_,
		_w1341_,
		_w1342_,
		_w1343_,
		_w1344_
	);
	LUT3 #(
		.INIT('ha8)
	) name1040 (
		_w305_,
		_w420_,
		_w421_,
		_w1345_
	);
	LUT3 #(
		.INIT('ha8)
	) name1041 (
		_w423_,
		_w433_,
		_w478_,
		_w1346_
	);
	LUT3 #(
		.INIT('ha8)
	) name1042 (
		_w406_,
		_w490_,
		_w480_,
		_w1347_
	);
	LUT3 #(
		.INIT('ha8)
	) name1043 (
		_w398_,
		_w440_,
		_w539_,
		_w1348_
	);
	LUT4 #(
		.INIT('h0001)
	) name1044 (
		_w1345_,
		_w1346_,
		_w1347_,
		_w1348_,
		_w1349_
	);
	LUT3 #(
		.INIT('he0)
	) name1045 (
		_w381_,
		_w385_,
		_w402_,
		_w1350_
	);
	LUT3 #(
		.INIT('ha8)
	) name1046 (
		_w323_,
		_w459_,
		_w548_,
		_w1351_
	);
	LUT3 #(
		.INIT('ha8)
	) name1047 (
		_w333_,
		_w435_,
		_w492_,
		_w1352_
	);
	LUT3 #(
		.INIT('ha8)
	) name1048 (
		_w343_,
		_w457_,
		_w471_,
		_w1353_
	);
	LUT4 #(
		.INIT('h0001)
	) name1049 (
		_w1350_,
		_w1351_,
		_w1352_,
		_w1353_,
		_w1354_
	);
	LUT3 #(
		.INIT('ha8)
	) name1050 (
		_w373_,
		_w455_,
		_w473_,
		_w1355_
	);
	LUT3 #(
		.INIT('ha8)
	) name1051 (
		_w363_,
		_w483_,
		_w561_,
		_w1356_
	);
	LUT3 #(
		.INIT('ha8)
	) name1052 (
		_w388_,
		_w449_,
		_w488_,
		_w1357_
	);
	LUT3 #(
		.INIT('ha8)
	) name1053 (
		_w312_,
		_w460_,
		_w559_,
		_w1358_
	);
	LUT4 #(
		.INIT('h0001)
	) name1054 (
		_w1355_,
		_w1356_,
		_w1357_,
		_w1358_,
		_w1359_
	);
	LUT4 #(
		.INIT('h8000)
	) name1055 (
		_w1354_,
		_w1359_,
		_w1344_,
		_w1349_,
		_w1360_
	);
	LUT2 #(
		.INIT('h9)
	) name1056 (
		_w1338_,
		_w1360_,
		_w1361_
	);
	LUT4 #(
		.INIT('h007f)
	) name1057 (
		_w1279_,
		_w1331_,
		_w1334_,
		_w1361_,
		_w1362_
	);
	LUT4 #(
		.INIT('h0d00)
	) name1058 (
		_w1230_,
		_w1333_,
		_w1304_,
		_w1362_,
		_w1363_
	);
	LUT4 #(
		.INIT('h1248)
	) name1059 (
		_w310_,
		_w568_,
		_w1278_,
		_w1300_,
		_w1364_
	);
	LUT4 #(
		.INIT('hdadf)
	) name1060 (
		_w1279_,
		_w1331_,
		_w1301_,
		_w1257_,
		_w1365_
	);
	LUT2 #(
		.INIT('h2)
	) name1061 (
		_w1230_,
		_w1365_,
		_w1366_
	);
	LUT2 #(
		.INIT('h4)
	) name1062 (
		_w1257_,
		_w1332_,
		_w1367_
	);
	LUT4 #(
		.INIT('h2184)
	) name1063 (
		_w310_,
		_w568_,
		_w1278_,
		_w1300_,
		_w1368_
	);
	LUT3 #(
		.INIT('h8c)
	) name1064 (
		_w1230_,
		_w1361_,
		_w1368_,
		_w1369_
	);
	LUT4 #(
		.INIT('h0990)
	) name1065 (
		_w1325_,
		_w1329_,
		_w1251_,
		_w1255_,
		_w1370_
	);
	LUT4 #(
		.INIT('h9669)
	) name1066 (
		_w1325_,
		_w1329_,
		_w1251_,
		_w1255_,
		_w1371_
	);
	LUT2 #(
		.INIT('h2)
	) name1067 (
		_w1364_,
		_w1371_,
		_w1372_
	);
	LUT4 #(
		.INIT('h197f)
	) name1068 (
		_w1331_,
		_w1257_,
		_w1302_,
		_w1364_,
		_w1373_
	);
	LUT3 #(
		.INIT('h40)
	) name1069 (
		_w1367_,
		_w1369_,
		_w1373_,
		_w1374_
	);
	LUT4 #(
		.INIT('h6006)
	) name1070 (
		_w1325_,
		_w1329_,
		_w1207_,
		_w1229_,
		_w1375_
	);
	LUT3 #(
		.INIT('h80)
	) name1071 (
		_w1257_,
		_w1364_,
		_w1375_,
		_w1376_
	);
	LUT4 #(
		.INIT('h0660)
	) name1072 (
		_w1325_,
		_w1329_,
		_w1207_,
		_w1229_,
		_w1377_
	);
	LUT4 #(
		.INIT('h0990)
	) name1073 (
		_w310_,
		_w1278_,
		_w1251_,
		_w1255_,
		_w1378_
	);
	LUT4 #(
		.INIT('h9009)
	) name1074 (
		_w310_,
		_w1278_,
		_w1251_,
		_w1255_,
		_w1379_
	);
	LUT4 #(
		.INIT('hc480)
	) name1075 (
		_w1301_,
		_w1377_,
		_w1378_,
		_w1379_,
		_w1380_
	);
	LUT2 #(
		.INIT('h1)
	) name1076 (
		_w1376_,
		_w1380_,
		_w1381_
	);
	LUT4 #(
		.INIT('hba00)
	) name1077 (
		_w1363_,
		_w1366_,
		_w1374_,
		_w1381_,
		_w1382_
	);
	LUT4 #(
		.INIT('h0100)
	) name1078 (
		\desIn[18]_pad ,
		\roundSel[4]_pad ,
		\roundSel[5]_pad ,
		_w305_,
		_w1383_
	);
	LUT4 #(
		.INIT('h2800)
	) name1079 (
		\FP_R_reg[19]/P0001 ,
		\roundSel[4]_pad ,
		\roundSel[5]_pad ,
		_w305_,
		_w1384_
	);
	LUT4 #(
		.INIT('h7c55)
	) name1080 (
		\FP_R_reg[51]/NET0131 ,
		\roundSel[4]_pad ,
		\roundSel[5]_pad ,
		_w305_,
		_w1385_
	);
	LUT3 #(
		.INIT('h45)
	) name1081 (
		_w1383_,
		_w1384_,
		_w1385_,
		_w1386_
	);
	LUT2 #(
		.INIT('h9)
	) name1082 (
		_w1382_,
		_w1386_,
		_w1387_
	);
	LUT4 #(
		.INIT('hf7c7)
	) name1083 (
		_w501_,
		_w528_,
		_w570_,
		_w626_,
		_w1388_
	);
	LUT4 #(
		.INIT('h0cbc)
	) name1084 (
		_w501_,
		_w528_,
		_w570_,
		_w626_,
		_w1389_
	);
	LUT4 #(
		.INIT('hfa10)
	) name1085 (
		_w597_,
		_w652_,
		_w1388_,
		_w1389_,
		_w1390_
	);
	LUT3 #(
		.INIT('h20)
	) name1086 (
		_w528_,
		_w626_,
		_w628_,
		_w1391_
	);
	LUT4 #(
		.INIT('h0200)
	) name1087 (
		_w528_,
		_w597_,
		_w626_,
		_w628_,
		_w1392_
	);
	LUT4 #(
		.INIT('h6006)
	) name1088 (
		_w592_,
		_w596_,
		_w620_,
		_w624_,
		_w1393_
	);
	LUT3 #(
		.INIT('h80)
	) name1089 (
		_w570_,
		_w598_,
		_w1393_,
		_w1394_
	);
	LUT2 #(
		.INIT('h1)
	) name1090 (
		_w1392_,
		_w1394_,
		_w1395_
	);
	LUT3 #(
		.INIT('he0)
	) name1091 (
		_w429_,
		_w1390_,
		_w1395_,
		_w1396_
	);
	LUT4 #(
		.INIT('hfd3d)
	) name1092 (
		_w501_,
		_w528_,
		_w570_,
		_w626_,
		_w1397_
	);
	LUT2 #(
		.INIT('h8)
	) name1093 (
		_w635_,
		_w652_,
		_w1398_
	);
	LUT4 #(
		.INIT('h5d7f)
	) name1094 (
		_w528_,
		_w570_,
		_w631_,
		_w652_,
		_w1399_
	);
	LUT4 #(
		.INIT('h7200)
	) name1095 (
		_w597_,
		_w649_,
		_w1397_,
		_w1399_,
		_w1400_
	);
	LUT3 #(
		.INIT('h20)
	) name1096 (
		_w501_,
		_w626_,
		_w635_,
		_w1401_
	);
	LUT4 #(
		.INIT('hbff6)
	) name1097 (
		_w501_,
		_w528_,
		_w570_,
		_w626_,
		_w1402_
	);
	LUT2 #(
		.INIT('h2)
	) name1098 (
		_w597_,
		_w1402_,
		_w1403_
	);
	LUT3 #(
		.INIT('h0d)
	) name1099 (
		_w429_,
		_w1400_,
		_w1403_,
		_w1404_
	);
	LUT4 #(
		.INIT('h0100)
	) name1100 (
		\desIn[22]_pad ,
		\roundSel[4]_pad ,
		\roundSel[5]_pad ,
		_w305_,
		_w1405_
	);
	LUT4 #(
		.INIT('h2800)
	) name1101 (
		\FP_R_reg[3]/P0001 ,
		\roundSel[4]_pad ,
		\roundSel[5]_pad ,
		_w305_,
		_w1406_
	);
	LUT4 #(
		.INIT('h7c55)
	) name1102 (
		\FP_R_reg[35]/NET0131 ,
		\roundSel[4]_pad ,
		\roundSel[5]_pad ,
		_w305_,
		_w1407_
	);
	LUT3 #(
		.INIT('h45)
	) name1103 (
		_w1405_,
		_w1406_,
		_w1407_,
		_w1408_
	);
	LUT3 #(
		.INIT('h87)
	) name1104 (
		_w1396_,
		_w1404_,
		_w1408_,
		_w1409_
	);
	LUT4 #(
		.INIT('h0200)
	) name1105 (
		\desIn[23]_pad ,
		\roundSel[4]_pad ,
		\roundSel[5]_pad ,
		_w305_,
		_w1410_
	);
	LUT4 #(
		.INIT('h4155)
	) name1106 (
		\FP_R_reg[3]/P0001 ,
		\roundSel[4]_pad ,
		\roundSel[5]_pad ,
		_w305_,
		_w1411_
	);
	LUT4 #(
		.INIT('he8ff)
	) name1107 (
		\FP_R_reg[35]/NET0131 ,
		\roundSel[4]_pad ,
		\roundSel[5]_pad ,
		_w305_,
		_w1412_
	);
	LUT3 #(
		.INIT('h45)
	) name1108 (
		_w1410_,
		_w1411_,
		_w1412_,
		_w1413_
	);
	LUT3 #(
		.INIT('hba)
	) name1109 (
		_w1410_,
		_w1411_,
		_w1412_,
		_w1414_
	);
	LUT4 #(
		.INIT('h3cdf)
	) name1110 (
		_w1162_,
		_w1080_,
		_w1107_,
		_w1134_,
		_w1415_
	);
	LUT2 #(
		.INIT('h2)
	) name1111 (
		_w1053_,
		_w1415_,
		_w1416_
	);
	LUT4 #(
		.INIT('h0660)
	) name1112 (
		_w1139_,
		_w1161_,
		_w1084_,
		_w1106_,
		_w1417_
	);
	LUT4 #(
		.INIT('h0660)
	) name1113 (
		_w1111_,
		_w1133_,
		_w1046_,
		_w1051_,
		_w1418_
	);
	LUT3 #(
		.INIT('he0)
	) name1114 (
		_w1180_,
		_w1417_,
		_w1418_,
		_w1419_
	);
	LUT3 #(
		.INIT('h40)
	) name1115 (
		_w1162_,
		_w1080_,
		_w1169_,
		_w1420_
	);
	LUT4 #(
		.INIT('h6006)
	) name1116 (
		_w1139_,
		_w1161_,
		_w1046_,
		_w1051_,
		_w1421_
	);
	LUT4 #(
		.INIT('h23ef)
	) name1117 (
		_w1107_,
		_w1134_,
		_w1168_,
		_w1421_,
		_w1422_
	);
	LUT3 #(
		.INIT('h10)
	) name1118 (
		_w1420_,
		_w1419_,
		_w1422_,
		_w1423_
	);
	LUT3 #(
		.INIT('h45)
	) name1119 (
		_w1025_,
		_w1416_,
		_w1423_,
		_w1424_
	);
	LUT3 #(
		.INIT('h02)
	) name1120 (
		_w1080_,
		_w1135_,
		_w1179_,
		_w1425_
	);
	LUT4 #(
		.INIT('hddf7)
	) name1121 (
		_w1162_,
		_w1080_,
		_w1135_,
		_w1179_,
		_w1426_
	);
	LUT2 #(
		.INIT('h2)
	) name1122 (
		_w1025_,
		_w1426_,
		_w1427_
	);
	LUT4 #(
		.INIT('h8cf3)
	) name1123 (
		_w1162_,
		_w1080_,
		_w1107_,
		_w1134_,
		_w1428_
	);
	LUT4 #(
		.INIT('h0660)
	) name1124 (
		_w1002_,
		_w1024_,
		_w1046_,
		_w1051_,
		_w1429_
	);
	LUT2 #(
		.INIT('h4)
	) name1125 (
		_w1428_,
		_w1429_,
		_w1430_
	);
	LUT4 #(
		.INIT('hd5f7)
	) name1126 (
		_w1162_,
		_w1080_,
		_w1134_,
		_w1179_,
		_w1431_
	);
	LUT4 #(
		.INIT('h0660)
	) name1127 (
		_w1002_,
		_w1024_,
		_w1111_,
		_w1133_,
		_w1432_
	);
	LUT4 #(
		.INIT('ha800)
	) name1128 (
		_w1053_,
		_w1180_,
		_w1417_,
		_w1432_,
		_w1433_
	);
	LUT3 #(
		.INIT('h0e)
	) name1129 (
		_w1053_,
		_w1431_,
		_w1433_,
		_w1434_
	);
	LUT3 #(
		.INIT('h10)
	) name1130 (
		_w1427_,
		_w1430_,
		_w1434_,
		_w1435_
	);
	LUT4 #(
		.INIT('h0100)
	) name1131 (
		\desIn[24]_pad ,
		\roundSel[4]_pad ,
		\roundSel[5]_pad ,
		_w305_,
		_w1436_
	);
	LUT4 #(
		.INIT('h2800)
	) name1132 (
		\FP_R_reg[28]/P0001 ,
		\roundSel[4]_pad ,
		\roundSel[5]_pad ,
		_w305_,
		_w1437_
	);
	LUT4 #(
		.INIT('h7c55)
	) name1133 (
		\FP_R_reg[60]/NET0131 ,
		\roundSel[4]_pad ,
		\roundSel[5]_pad ,
		_w305_,
		_w1438_
	);
	LUT3 #(
		.INIT('h45)
	) name1134 (
		_w1436_,
		_w1437_,
		_w1438_,
		_w1439_
	);
	LUT3 #(
		.INIT('h4b)
	) name1135 (
		_w1424_,
		_w1435_,
		_w1439_,
		_w1440_
	);
	LUT4 #(
		.INIT('h0200)
	) name1136 (
		\desIn[25]_pad ,
		\roundSel[4]_pad ,
		\roundSel[5]_pad ,
		_w305_,
		_w1441_
	);
	LUT4 #(
		.INIT('h4155)
	) name1137 (
		\FP_R_reg[28]/P0001 ,
		\roundSel[4]_pad ,
		\roundSel[5]_pad ,
		_w305_,
		_w1442_
	);
	LUT4 #(
		.INIT('he8ff)
	) name1138 (
		\FP_R_reg[60]/NET0131 ,
		\roundSel[4]_pad ,
		\roundSel[5]_pad ,
		_w305_,
		_w1443_
	);
	LUT3 #(
		.INIT('h45)
	) name1139 (
		_w1441_,
		_w1442_,
		_w1443_,
		_w1444_
	);
	LUT3 #(
		.INIT('hba)
	) name1140 (
		_w1441_,
		_w1442_,
		_w1443_,
		_w1445_
	);
	LUT4 #(
		.INIT('h5d7f)
	) name1141 (
		_w820_,
		_w877_,
		_w957_,
		_w959_,
		_w1446_
	);
	LUT4 #(
		.INIT('h37bf)
	) name1142 (
		_w820_,
		_w956_,
		_w957_,
		_w929_,
		_w1447_
	);
	LUT3 #(
		.INIT('h40)
	) name1143 (
		_w877_,
		_w962_,
		_w973_,
		_w1448_
	);
	LUT4 #(
		.INIT('h0990)
	) name1144 (
		_w899_,
		_w904_,
		_w814_,
		_w818_,
		_w1449_
	);
	LUT4 #(
		.INIT('h9669)
	) name1145 (
		_w899_,
		_w904_,
		_w814_,
		_w818_,
		_w1450_
	);
	LUT2 #(
		.INIT('h2)
	) name1146 (
		_w976_,
		_w1450_,
		_w1451_
	);
	LUT4 #(
		.INIT('h0200)
	) name1147 (
		_w1446_,
		_w1448_,
		_w1451_,
		_w1447_,
		_w1452_
	);
	LUT2 #(
		.INIT('h2)
	) name1148 (
		_w763_,
		_w1452_,
		_w1453_
	);
	LUT3 #(
		.INIT('ha8)
	) name1149 (
		_w959_,
		_w963_,
		_w965_,
		_w1454_
	);
	LUT4 #(
		.INIT('h6006)
	) name1150 (
		_w814_,
		_w818_,
		_w950_,
		_w954_,
		_w1455_
	);
	LUT2 #(
		.INIT('h8)
	) name1151 (
		_w962_,
		_w1455_,
		_w1456_
	);
	LUT3 #(
		.INIT('h01)
	) name1152 (
		_w985_,
		_w1456_,
		_w1454_,
		_w1457_
	);
	LUT4 #(
		.INIT('h2814)
	) name1153 (
		_w499_,
		_w814_,
		_w818_,
		_w927_,
		_w1458_
	);
	LUT4 #(
		.INIT('h3310)
	) name1154 (
		_w877_,
		_w956_,
		_w929_,
		_w1458_,
		_w1459_
	);
	LUT2 #(
		.INIT('h2)
	) name1155 (
		_w981_,
		_w1459_,
		_w1460_
	);
	LUT2 #(
		.INIT('h8)
	) name1156 (
		_w960_,
		_w929_,
		_w1461_
	);
	LUT4 #(
		.INIT('haebf)
	) name1157 (
		_w820_,
		_w877_,
		_w962_,
		_w929_,
		_w1462_
	);
	LUT3 #(
		.INIT('h80)
	) name1158 (
		_w928_,
		_w976_,
		_w978_,
		_w1463_
	);
	LUT4 #(
		.INIT('h0031)
	) name1159 (
		_w956_,
		_w986_,
		_w1462_,
		_w1463_,
		_w1464_
	);
	LUT4 #(
		.INIT('hea00)
	) name1160 (
		_w763_,
		_w1457_,
		_w1460_,
		_w1464_,
		_w1465_
	);
	LUT4 #(
		.INIT('h0100)
	) name1161 (
		\desIn[26]_pad ,
		\roundSel[4]_pad ,
		\roundSel[5]_pad ,
		_w305_,
		_w1466_
	);
	LUT4 #(
		.INIT('h2800)
	) name1162 (
		\FP_R_reg[20]/P0001 ,
		\roundSel[4]_pad ,
		\roundSel[5]_pad ,
		_w305_,
		_w1467_
	);
	LUT4 #(
		.INIT('h7c55)
	) name1163 (
		\FP_R_reg[52]/NET0131 ,
		\roundSel[4]_pad ,
		\roundSel[5]_pad ,
		_w305_,
		_w1468_
	);
	LUT3 #(
		.INIT('h45)
	) name1164 (
		_w1466_,
		_w1467_,
		_w1468_,
		_w1469_
	);
	LUT3 #(
		.INIT('h4b)
	) name1165 (
		_w1453_,
		_w1465_,
		_w1469_,
		_w1470_
	);
	LUT4 #(
		.INIT('h0200)
	) name1166 (
		\desIn[28]_pad ,
		\roundSel[4]_pad ,
		\roundSel[5]_pad ,
		_w305_,
		_w1471_
	);
	LUT4 #(
		.INIT('h4155)
	) name1167 (
		\FP_R_reg[44]/NET0131 ,
		\roundSel[4]_pad ,
		\roundSel[5]_pad ,
		_w305_,
		_w1472_
	);
	LUT4 #(
		.INIT('he8ff)
	) name1168 (
		\FP_R_reg[12]/P0001 ,
		\roundSel[4]_pad ,
		\roundSel[5]_pad ,
		_w305_,
		_w1473_
	);
	LUT3 #(
		.INIT('h45)
	) name1169 (
		_w1471_,
		_w1472_,
		_w1473_,
		_w1474_
	);
	LUT3 #(
		.INIT('hc8)
	) name1170 (
		_w374_,
		_w323_,
		_w444_,
		_w1475_
	);
	LUT3 #(
		.INIT('ha8)
	) name1171 (
		_w419_,
		_w408_,
		_w492_,
		_w1476_
	);
	LUT3 #(
		.INIT('ha8)
	) name1172 (
		_w377_,
		_w392_,
		_w478_,
		_w1477_
	);
	LUT3 #(
		.INIT('hc8)
	) name1173 (
		_w375_,
		_w312_,
		_w483_,
		_w1478_
	);
	LUT4 #(
		.INIT('h0001)
	) name1174 (
		_w1475_,
		_w1476_,
		_w1477_,
		_w1478_,
		_w1479_
	);
	LUT3 #(
		.INIT('ha8)
	) name1175 (
		_w363_,
		_w407_,
		_w460_,
		_w1480_
	);
	LUT3 #(
		.INIT('ha8)
	) name1176 (
		_w305_,
		_w341_,
		_w490_,
		_w1481_
	);
	LUT3 #(
		.INIT('ha8)
	) name1177 (
		_w343_,
		_w412_,
		_w399_,
		_w1482_
	);
	LUT3 #(
		.INIT('ha8)
	) name1178 (
		_w373_,
		_w317_,
		_w327_,
		_w1483_
	);
	LUT4 #(
		.INIT('h0001)
	) name1179 (
		_w1480_,
		_w1481_,
		_w1482_,
		_w1483_,
		_w1484_
	);
	LUT3 #(
		.INIT('hc8)
	) name1180 (
		_w337_,
		_w423_,
		_w403_,
		_w1485_
	);
	LUT3 #(
		.INIT('hc8)
	) name1181 (
		_w425_,
		_w402_,
		_w488_,
		_w1486_
	);
	LUT3 #(
		.INIT('hc8)
	) name1182 (
		_w351_,
		_w411_,
		_w459_,
		_w1487_
	);
	LUT3 #(
		.INIT('he0)
	) name1183 (
		_w367_,
		_w420_,
		_w406_,
		_w1488_
	);
	LUT4 #(
		.INIT('h0001)
	) name1184 (
		_w1485_,
		_w1486_,
		_w1487_,
		_w1488_,
		_w1489_
	);
	LUT3 #(
		.INIT('hc8)
	) name1185 (
		_w357_,
		_w333_,
		_w424_,
		_w1490_
	);
	LUT3 #(
		.INIT('hc8)
	) name1186 (
		_w347_,
		_w398_,
		_w465_,
		_w1491_
	);
	LUT3 #(
		.INIT('ha8)
	) name1187 (
		_w415_,
		_w396_,
		_w440_,
		_w1492_
	);
	LUT3 #(
		.INIT('he0)
	) name1188 (
		_w381_,
		_w416_,
		_w388_,
		_w1493_
	);
	LUT4 #(
		.INIT('h0001)
	) name1189 (
		_w1490_,
		_w1491_,
		_w1492_,
		_w1493_,
		_w1494_
	);
	LUT4 #(
		.INIT('h8000)
	) name1190 (
		_w1489_,
		_w1494_,
		_w1479_,
		_w1484_,
		_w1495_
	);
	LUT4 #(
		.INIT('h0200)
	) name1191 (
		\desIn[17]_pad ,
		\roundSel[4]_pad ,
		\roundSel[5]_pad ,
		_w305_,
		_w1496_
	);
	LUT4 #(
		.INIT('h4155)
	) name1192 (
		\FP_R_reg[27]/P0001 ,
		\roundSel[4]_pad ,
		\roundSel[5]_pad ,
		_w305_,
		_w1497_
	);
	LUT4 #(
		.INIT('he8ff)
	) name1193 (
		\FP_R_reg[59]/NET0131 ,
		\roundSel[4]_pad ,
		\roundSel[5]_pad ,
		_w305_,
		_w1498_
	);
	LUT3 #(
		.INIT('h45)
	) name1194 (
		_w1496_,
		_w1497_,
		_w1498_,
		_w1499_
	);
	LUT3 #(
		.INIT('hba)
	) name1195 (
		_w1496_,
		_w1497_,
		_w1498_,
		_w1500_
	);
	LUT2 #(
		.INIT('h9)
	) name1196 (
		_w1495_,
		_w1499_,
		_w1501_
	);
	LUT3 #(
		.INIT('he0)
	) name1197 (
		_w374_,
		_w413_,
		_w423_,
		_w1502_
	);
	LUT3 #(
		.INIT('hc8)
	) name1198 (
		_w317_,
		_w402_,
		_w548_,
		_w1503_
	);
	LUT3 #(
		.INIT('ha8)
	) name1199 (
		_w411_,
		_w421_,
		_w424_,
		_w1504_
	);
	LUT3 #(
		.INIT('ha8)
	) name1200 (
		_w363_,
		_w396_,
		_w400_,
		_w1505_
	);
	LUT4 #(
		.INIT('h0001)
	) name1201 (
		_w1502_,
		_w1503_,
		_w1504_,
		_w1505_,
		_w1506_
	);
	LUT3 #(
		.INIT('ha8)
	) name1202 (
		_w377_,
		_w327_,
		_w559_,
		_w1507_
	);
	LUT3 #(
		.INIT('hc8)
	) name1203 (
		_w385_,
		_w323_,
		_w337_,
		_w1508_
	);
	LUT3 #(
		.INIT('hc8)
	) name1204 (
		_w341_,
		_w343_,
		_w408_,
		_w1509_
	);
	LUT3 #(
		.INIT('ha8)
	) name1205 (
		_w305_,
		_w399_,
		_w556_,
		_w1510_
	);
	LUT4 #(
		.INIT('h0001)
	) name1206 (
		_w1507_,
		_w1508_,
		_w1509_,
		_w1510_,
		_w1511_
	);
	LUT3 #(
		.INIT('ha8)
	) name1207 (
		_w373_,
		_w425_,
		_w392_,
		_w1512_
	);
	LUT3 #(
		.INIT('hc8)
	) name1208 (
		_w321_,
		_w415_,
		_w407_,
		_w1513_
	);
	LUT3 #(
		.INIT('he0)
	) name1209 (
		_w371_,
		_w375_,
		_w388_,
		_w1514_
	);
	LUT3 #(
		.INIT('ha8)
	) name1210 (
		_w312_,
		_w416_,
		_w404_,
		_w1515_
	);
	LUT4 #(
		.INIT('h0001)
	) name1211 (
		_w1512_,
		_w1513_,
		_w1514_,
		_w1515_,
		_w1516_
	);
	LUT3 #(
		.INIT('he0)
	) name1212 (
		_w361_,
		_w367_,
		_w398_,
		_w1517_
	);
	LUT3 #(
		.INIT('hc8)
	) name1213 (
		_w331_,
		_w333_,
		_w351_,
		_w1518_
	);
	LUT3 #(
		.INIT('he0)
	) name1214 (
		_w347_,
		_w417_,
		_w406_,
		_w1519_
	);
	LUT3 #(
		.INIT('hc8)
	) name1215 (
		_w412_,
		_w419_,
		_w539_,
		_w1520_
	);
	LUT4 #(
		.INIT('h0001)
	) name1216 (
		_w1517_,
		_w1518_,
		_w1519_,
		_w1520_,
		_w1521_
	);
	LUT4 #(
		.INIT('h8000)
	) name1217 (
		_w1516_,
		_w1521_,
		_w1506_,
		_w1511_,
		_w1522_
	);
	LUT2 #(
		.INIT('h9)
	) name1218 (
		_w1255_,
		_w1522_,
		_w1523_
	);
	LUT3 #(
		.INIT('ha8)
	) name1219 (
		_w373_,
		_w435_,
		_w553_,
		_w1524_
	);
	LUT3 #(
		.INIT('hc8)
	) name1220 (
		_w331_,
		_w419_,
		_w465_,
		_w1525_
	);
	LUT3 #(
		.INIT('hc8)
	) name1221 (
		_w321_,
		_w398_,
		_w492_,
		_w1526_
	);
	LUT3 #(
		.INIT('ha8)
	) name1222 (
		_w388_,
		_w480_,
		_w548_,
		_w1527_
	);
	LUT4 #(
		.INIT('h0001)
	) name1223 (
		_w1524_,
		_w1525_,
		_w1526_,
		_w1527_,
		_w1528_
	);
	LUT3 #(
		.INIT('hc8)
	) name1224 (
		_w385_,
		_w411_,
		_w490_,
		_w1529_
	);
	LUT3 #(
		.INIT('ha8)
	) name1225 (
		_w377_,
		_w413_,
		_w483_,
		_w1530_
	);
	LUT3 #(
		.INIT('hc8)
	) name1226 (
		_w371_,
		_w402_,
		_w444_,
		_w1531_
	);
	LUT3 #(
		.INIT('ha8)
	) name1227 (
		_w312_,
		_w400_,
		_w478_,
		_w1532_
	);
	LUT4 #(
		.INIT('h0001)
	) name1228 (
		_w1529_,
		_w1530_,
		_w1531_,
		_w1532_,
		_w1533_
	);
	LUT3 #(
		.INIT('ha8)
	) name1229 (
		_w406_,
		_w449_,
		_w556_,
		_w1534_
	);
	LUT3 #(
		.INIT('ha8)
	) name1230 (
		_w305_,
		_w417_,
		_w459_,
		_w1535_
	);
	LUT3 #(
		.INIT('ha8)
	) name1231 (
		_w363_,
		_w404_,
		_w457_,
		_w1536_
	);
	LUT3 #(
		.INIT('ha8)
	) name1232 (
		_w333_,
		_w473_,
		_w539_,
		_w1537_
	);
	LUT4 #(
		.INIT('h0001)
	) name1233 (
		_w1534_,
		_w1535_,
		_w1536_,
		_w1537_,
		_w1538_
	);
	LUT3 #(
		.INIT('ha8)
	) name1234 (
		_w423_,
		_w471_,
		_w559_,
		_w1539_
	);
	LUT3 #(
		.INIT('hc8)
	) name1235 (
		_w361_,
		_w415_,
		_w455_,
		_w1540_
	);
	LUT3 #(
		.INIT('ha8)
	) name1236 (
		_w323_,
		_w421_,
		_w488_,
		_w1541_
	);
	LUT3 #(
		.INIT('ha8)
	) name1237 (
		_w343_,
		_w433_,
		_w561_,
		_w1542_
	);
	LUT4 #(
		.INIT('h0001)
	) name1238 (
		_w1539_,
		_w1540_,
		_w1541_,
		_w1542_,
		_w1543_
	);
	LUT4 #(
		.INIT('h8000)
	) name1239 (
		_w1538_,
		_w1543_,
		_w1528_,
		_w1533_,
		_w1544_
	);
	LUT2 #(
		.INIT('h6)
	) name1240 (
		_w1338_,
		_w1544_,
		_w1545_
	);
	LUT4 #(
		.INIT('h8421)
	) name1241 (
		_w1255_,
		_w1338_,
		_w1522_,
		_w1544_,
		_w1546_
	);
	LUT3 #(
		.INIT('hc8)
	) name1242 (
		_w357_,
		_w373_,
		_w440_,
		_w1547_
	);
	LUT3 #(
		.INIT('ha8)
	) name1243 (
		_w419_,
		_w396_,
		_w473_,
		_w1548_
	);
	LUT3 #(
		.INIT('hc8)
	) name1244 (
		_w327_,
		_w415_,
		_w492_,
		_w1549_
	);
	LUT3 #(
		.INIT('ha8)
	) name1245 (
		_w312_,
		_w337_,
		_w457_,
		_w1550_
	);
	LUT4 #(
		.INIT('h0001)
	) name1246 (
		_w1547_,
		_w1548_,
		_w1549_,
		_w1550_,
		_w1551_
	);
	LUT3 #(
		.INIT('ha8)
	) name1247 (
		_w343_,
		_w403_,
		_w460_,
		_w1552_
	);
	LUT3 #(
		.INIT('hc8)
	) name1248 (
		_w351_,
		_w402_,
		_w480_,
		_w1553_
	);
	LUT3 #(
		.INIT('ha8)
	) name1249 (
		_w363_,
		_w412_,
		_w478_,
		_w1554_
	);
	LUT3 #(
		.INIT('ha8)
	) name1250 (
		_w423_,
		_w399_,
		_w483_,
		_w1555_
	);
	LUT4 #(
		.INIT('h0001)
	) name1251 (
		_w1552_,
		_w1553_,
		_w1554_,
		_w1555_,
		_w1556_
	);
	LUT3 #(
		.INIT('hc8)
	) name1252 (
		_w420_,
		_w388_,
		_w444_,
		_w1557_
	);
	LUT3 #(
		.INIT('ha8)
	) name1253 (
		_w305_,
		_w374_,
		_w449_,
		_w1558_
	);
	LUT3 #(
		.INIT('hc8)
	) name1254 (
		_w424_,
		_w398_,
		_w455_,
		_w1559_
	);
	LUT3 #(
		.INIT('hc8)
	) name1255 (
		_w381_,
		_w406_,
		_w459_,
		_w1560_
	);
	LUT4 #(
		.INIT('h0001)
	) name1256 (
		_w1557_,
		_w1558_,
		_w1559_,
		_w1560_,
		_w1561_
	);
	LUT3 #(
		.INIT('hc8)
	) name1257 (
		_w317_,
		_w333_,
		_w465_,
		_w1562_
	);
	LUT3 #(
		.INIT('ha8)
	) name1258 (
		_w377_,
		_w407_,
		_w471_,
		_w1563_
	);
	LUT3 #(
		.INIT('hc8)
	) name1259 (
		_w367_,
		_w411_,
		_w488_,
		_w1564_
	);
	LUT3 #(
		.INIT('ha8)
	) name1260 (
		_w323_,
		_w416_,
		_w490_,
		_w1565_
	);
	LUT4 #(
		.INIT('h0001)
	) name1261 (
		_w1562_,
		_w1563_,
		_w1564_,
		_w1565_,
		_w1566_
	);
	LUT4 #(
		.INIT('h8000)
	) name1262 (
		_w1561_,
		_w1566_,
		_w1551_,
		_w1556_,
		_w1567_
	);
	LUT4 #(
		.INIT('h0200)
	) name1263 (
		\desIn[9]_pad ,
		\roundSel[4]_pad ,
		\roundSel[5]_pad ,
		_w305_,
		_w1568_
	);
	LUT4 #(
		.INIT('h4155)
	) name1264 (
		\FP_R_reg[26]/P0001 ,
		\roundSel[4]_pad ,
		\roundSel[5]_pad ,
		_w305_,
		_w1569_
	);
	LUT4 #(
		.INIT('he8ff)
	) name1265 (
		\FP_R_reg[58]/NET0131 ,
		\roundSel[4]_pad ,
		\roundSel[5]_pad ,
		_w305_,
		_w1570_
	);
	LUT3 #(
		.INIT('h45)
	) name1266 (
		_w1568_,
		_w1569_,
		_w1570_,
		_w1571_
	);
	LUT3 #(
		.INIT('hba)
	) name1267 (
		_w1568_,
		_w1569_,
		_w1570_,
		_w1572_
	);
	LUT2 #(
		.INIT('h6)
	) name1268 (
		_w1567_,
		_w1571_,
		_w1573_
	);
	LUT4 #(
		.INIT('h0660)
	) name1269 (
		_w1255_,
		_w1522_,
		_w1567_,
		_w1571_,
		_w1574_
	);
	LUT3 #(
		.INIT('ha8)
	) name1270 (
		_w363_,
		_w425_,
		_w556_,
		_w1575_
	);
	LUT3 #(
		.INIT('ha8)
	) name1271 (
		_w377_,
		_w351_,
		_w480_,
		_w1576_
	);
	LUT3 #(
		.INIT('hc8)
	) name1272 (
		_w371_,
		_w423_,
		_w539_,
		_w1577_
	);
	LUT3 #(
		.INIT('ha8)
	) name1273 (
		_w411_,
		_w392_,
		_w561_,
		_w1578_
	);
	LUT4 #(
		.INIT('h0001)
	) name1274 (
		_w1575_,
		_w1576_,
		_w1577_,
		_w1578_,
		_w1579_
	);
	LUT3 #(
		.INIT('ha8)
	) name1275 (
		_w333_,
		_w417_,
		_w559_,
		_w1580_
	);
	LUT3 #(
		.INIT('ha8)
	) name1276 (
		_w305_,
		_w396_,
		_w473_,
		_w1581_
	);
	LUT3 #(
		.INIT('ha8)
	) name1277 (
		_w402_,
		_w407_,
		_w471_,
		_w1582_
	);
	LUT3 #(
		.INIT('ha8)
	) name1278 (
		_w373_,
		_w421_,
		_w400_,
		_w1583_
	);
	LUT4 #(
		.INIT('h0001)
	) name1279 (
		_w1580_,
		_w1581_,
		_w1582_,
		_w1583_,
		_w1584_
	);
	LUT3 #(
		.INIT('hc8)
	) name1280 (
		_w341_,
		_w415_,
		_w548_,
		_w1585_
	);
	LUT3 #(
		.INIT('hc8)
	) name1281 (
		_w374_,
		_w419_,
		_w449_,
		_w1586_
	);
	LUT3 #(
		.INIT('ha8)
	) name1282 (
		_w312_,
		_w347_,
		_w435_,
		_w1587_
	);
	LUT3 #(
		.INIT('he0)
	) name1283 (
		_w385_,
		_w321_,
		_w343_,
		_w1588_
	);
	LUT4 #(
		.INIT('h0001)
	) name1284 (
		_w1585_,
		_w1586_,
		_w1587_,
		_w1588_,
		_w1589_
	);
	LUT3 #(
		.INIT('ha8)
	) name1285 (
		_w323_,
		_w408_,
		_w553_,
		_w1590_
	);
	LUT3 #(
		.INIT('hc8)
	) name1286 (
		_w375_,
		_w398_,
		_w433_,
		_w1591_
	);
	LUT3 #(
		.INIT('he0)
	) name1287 (
		_w361_,
		_w413_,
		_w388_,
		_w1592_
	);
	LUT3 #(
		.INIT('he0)
	) name1288 (
		_w331_,
		_w404_,
		_w406_,
		_w1593_
	);
	LUT4 #(
		.INIT('h0001)
	) name1289 (
		_w1590_,
		_w1591_,
		_w1592_,
		_w1593_,
		_w1594_
	);
	LUT4 #(
		.INIT('h8000)
	) name1290 (
		_w1589_,
		_w1594_,
		_w1579_,
		_w1584_,
		_w1595_
	);
	LUT4 #(
		.INIT('h0200)
	) name1291 (
		\desIn[33]_pad ,
		\roundSel[4]_pad ,
		\roundSel[5]_pad ,
		_w305_,
		_w1596_
	);
	LUT4 #(
		.INIT('h4155)
	) name1292 (
		\FP_R_reg[29]/P0001 ,
		\roundSel[4]_pad ,
		\roundSel[5]_pad ,
		_w305_,
		_w1597_
	);
	LUT4 #(
		.INIT('he8ff)
	) name1293 (
		\FP_R_reg[61]/NET0131 ,
		\roundSel[4]_pad ,
		\roundSel[5]_pad ,
		_w305_,
		_w1598_
	);
	LUT3 #(
		.INIT('h45)
	) name1294 (
		_w1596_,
		_w1597_,
		_w1598_,
		_w1599_
	);
	LUT3 #(
		.INIT('hba)
	) name1295 (
		_w1596_,
		_w1597_,
		_w1598_,
		_w1600_
	);
	LUT2 #(
		.INIT('h6)
	) name1296 (
		_w1595_,
		_w1599_,
		_w1601_
	);
	LUT4 #(
		.INIT('h0660)
	) name1297 (
		_w1338_,
		_w1544_,
		_w1595_,
		_w1599_,
		_w1602_
	);
	LUT4 #(
		.INIT('ha888)
	) name1298 (
		_w1501_,
		_w1546_,
		_w1574_,
		_w1602_,
		_w1603_
	);
	LUT4 #(
		.INIT('h0990)
	) name1299 (
		_w1338_,
		_w1544_,
		_w1595_,
		_w1599_,
		_w1604_
	);
	LUT4 #(
		.INIT('h6006)
	) name1300 (
		_w1255_,
		_w1522_,
		_w1567_,
		_w1571_,
		_w1605_
	);
	LUT2 #(
		.INIT('h8)
	) name1301 (
		_w1604_,
		_w1605_,
		_w1606_
	);
	LUT4 #(
		.INIT('h9009)
	) name1302 (
		_w1255_,
		_w1522_,
		_w1567_,
		_w1571_,
		_w1607_
	);
	LUT3 #(
		.INIT('hc8)
	) name1303 (
		_w321_,
		_w411_,
		_w416_,
		_w1608_
	);
	LUT3 #(
		.INIT('he0)
	) name1304 (
		_w374_,
		_w425_,
		_w406_,
		_w1609_
	);
	LUT3 #(
		.INIT('hc8)
	) name1305 (
		_w413_,
		_w415_,
		_w424_,
		_w1610_
	);
	LUT3 #(
		.INIT('ha8)
	) name1306 (
		_w363_,
		_w331_,
		_w337_,
		_w1611_
	);
	LUT4 #(
		.INIT('h0001)
	) name1307 (
		_w1608_,
		_w1609_,
		_w1610_,
		_w1611_,
		_w1612_
	);
	LUT3 #(
		.INIT('hc8)
	) name1308 (
		_w361_,
		_w377_,
		_w399_,
		_w1613_
	);
	LUT3 #(
		.INIT('he0)
	) name1309 (
		_w341_,
		_w351_,
		_w388_,
		_w1614_
	);
	LUT3 #(
		.INIT('hc8)
	) name1310 (
		_w417_,
		_w423_,
		_w407_,
		_w1615_
	);
	LUT3 #(
		.INIT('hc8)
	) name1311 (
		_w317_,
		_w419_,
		_w404_,
		_w1616_
	);
	LUT4 #(
		.INIT('h0001)
	) name1312 (
		_w1613_,
		_w1614_,
		_w1615_,
		_w1616_,
		_w1617_
	);
	LUT3 #(
		.INIT('he0)
	) name1313 (
		_w385_,
		_w327_,
		_w398_,
		_w1618_
	);
	LUT3 #(
		.INIT('hc8)
	) name1314 (
		_w375_,
		_w343_,
		_w392_,
		_w1619_
	);
	LUT3 #(
		.INIT('hc8)
	) name1315 (
		_w420_,
		_w402_,
		_w539_,
		_w1620_
	);
	LUT3 #(
		.INIT('ha8)
	) name1316 (
		_w373_,
		_w347_,
		_w408_,
		_w1621_
	);
	LUT4 #(
		.INIT('h0001)
	) name1317 (
		_w1618_,
		_w1619_,
		_w1620_,
		_w1621_,
		_w1622_
	);
	LUT3 #(
		.INIT('hc8)
	) name1318 (
		_w367_,
		_w323_,
		_w400_,
		_w1623_
	);
	LUT3 #(
		.INIT('hc8)
	) name1319 (
		_w371_,
		_w333_,
		_w396_,
		_w1624_
	);
	LUT3 #(
		.INIT('ha8)
	) name1320 (
		_w305_,
		_w381_,
		_w559_,
		_w1625_
	);
	LUT3 #(
		.INIT('ha8)
	) name1321 (
		_w312_,
		_w412_,
		_w421_,
		_w1626_
	);
	LUT4 #(
		.INIT('h0001)
	) name1322 (
		_w1623_,
		_w1624_,
		_w1625_,
		_w1626_,
		_w1627_
	);
	LUT4 #(
		.INIT('h8000)
	) name1323 (
		_w1622_,
		_w1627_,
		_w1612_,
		_w1617_,
		_w1628_
	);
	LUT2 #(
		.INIT('h9)
	) name1324 (
		_w1444_,
		_w1628_,
		_w1629_
	);
	LUT3 #(
		.INIT('h70)
	) name1325 (
		_w1602_,
		_w1607_,
		_w1629_,
		_w1630_
	);
	LUT4 #(
		.INIT('h9009)
	) name1326 (
		_w1338_,
		_w1544_,
		_w1595_,
		_w1599_,
		_w1631_
	);
	LUT3 #(
		.INIT('h40)
	) name1327 (
		_w1523_,
		_w1573_,
		_w1631_,
		_w1632_
	);
	LUT4 #(
		.INIT('h4182)
	) name1328 (
		_w1255_,
		_w1495_,
		_w1499_,
		_w1522_,
		_w1633_
	);
	LUT4 #(
		.INIT('h6006)
	) name1329 (
		_w1338_,
		_w1544_,
		_w1595_,
		_w1599_,
		_w1634_
	);
	LUT4 #(
		.INIT('hc100)
	) name1330 (
		_w1501_,
		_w1523_,
		_w1573_,
		_w1634_,
		_w1635_
	);
	LUT4 #(
		.INIT('h0100)
	) name1331 (
		_w1606_,
		_w1632_,
		_w1635_,
		_w1630_,
		_w1636_
	);
	LUT4 #(
		.INIT('h6996)
	) name1332 (
		_w1255_,
		_w1522_,
		_w1567_,
		_w1571_,
		_w1637_
	);
	LUT4 #(
		.INIT('h9669)
	) name1333 (
		_w1338_,
		_w1544_,
		_w1595_,
		_w1599_,
		_w1638_
	);
	LUT3 #(
		.INIT('h40)
	) name1334 (
		_w1546_,
		_w1638_,
		_w1637_,
		_w1639_
	);
	LUT4 #(
		.INIT('h0660)
	) name1335 (
		_w1255_,
		_w1522_,
		_w1595_,
		_w1599_,
		_w1640_
	);
	LUT4 #(
		.INIT('h3101)
	) name1336 (
		_w1501_,
		_w1545_,
		_w1573_,
		_w1640_,
		_w1641_
	);
	LUT3 #(
		.INIT('he0)
	) name1337 (
		_w1607_,
		_w1633_,
		_w1634_,
		_w1642_
	);
	LUT4 #(
		.INIT('h9009)
	) name1338 (
		_w1255_,
		_w1522_,
		_w1595_,
		_w1599_,
		_w1643_
	);
	LUT4 #(
		.INIT('h6996)
	) name1339 (
		_w1255_,
		_w1522_,
		_w1595_,
		_w1599_,
		_w1644_
	);
	LUT2 #(
		.INIT('h1)
	) name1340 (
		_w1501_,
		_w1644_,
		_w1645_
	);
	LUT4 #(
		.INIT('h0001)
	) name1341 (
		_w1629_,
		_w1641_,
		_w1642_,
		_w1645_,
		_w1646_
	);
	LUT4 #(
		.INIT('hb0bb)
	) name1342 (
		_w1603_,
		_w1636_,
		_w1639_,
		_w1646_,
		_w1647_
	);
	LUT2 #(
		.INIT('h9)
	) name1343 (
		_w1474_,
		_w1647_,
		_w1648_
	);
	LUT3 #(
		.INIT('ha8)
	) name1344 (
		_w402_,
		_w752_,
		_w849_,
		_w1649_
	);
	LUT3 #(
		.INIT('ha8)
	) name1345 (
		_w398_,
		_w696_,
		_w824_,
		_w1650_
	);
	LUT3 #(
		.INIT('ha8)
	) name1346 (
		_w388_,
		_w767_,
		_w786_,
		_w1651_
	);
	LUT3 #(
		.INIT('ha8)
	) name1347 (
		_w377_,
		_w739_,
		_w856_,
		_w1652_
	);
	LUT4 #(
		.INIT('h0001)
	) name1348 (
		_w1649_,
		_w1650_,
		_w1651_,
		_w1652_,
		_w1653_
	);
	LUT3 #(
		.INIT('ha8)
	) name1349 (
		_w419_,
		_w708_,
		_w865_,
		_w1654_
	);
	LUT3 #(
		.INIT('ha8)
	) name1350 (
		_w411_,
		_w736_,
		_w858_,
		_w1655_
	);
	LUT3 #(
		.INIT('ha8)
	) name1351 (
		_w343_,
		_w806_,
		_w772_,
		_w1656_
	);
	LUT3 #(
		.INIT('ha8)
	) name1352 (
		_w312_,
		_w724_,
		_w860_,
		_w1657_
	);
	LUT4 #(
		.INIT('h0001)
	) name1353 (
		_w1654_,
		_w1655_,
		_w1656_,
		_w1657_,
		_w1658_
	);
	LUT3 #(
		.INIT('ha8)
	) name1354 (
		_w305_,
		_w730_,
		_w831_,
		_w1659_
	);
	LUT3 #(
		.INIT('ha8)
	) name1355 (
		_w415_,
		_w842_,
		_w809_,
		_w1660_
	);
	LUT3 #(
		.INIT('ha8)
	) name1356 (
		_w333_,
		_w868_,
		_w811_,
		_w1661_
	);
	LUT3 #(
		.INIT('ha8)
	) name1357 (
		_w363_,
		_w863_,
		_w793_,
		_w1662_
	);
	LUT4 #(
		.INIT('h0001)
	) name1358 (
		_w1659_,
		_w1660_,
		_w1661_,
		_w1662_,
		_w1663_
	);
	LUT3 #(
		.INIT('ha8)
	) name1359 (
		_w323_,
		_w686_,
		_w837_,
		_w1664_
	);
	LUT3 #(
		.INIT('ha8)
	) name1360 (
		_w373_,
		_w802_,
		_w797_,
		_w1665_
	);
	LUT3 #(
		.INIT('ha8)
	) name1361 (
		_w406_,
		_w788_,
		_w774_,
		_w1666_
	);
	LUT3 #(
		.INIT('ha8)
	) name1362 (
		_w423_,
		_w847_,
		_w779_,
		_w1667_
	);
	LUT4 #(
		.INIT('h0001)
	) name1363 (
		_w1664_,
		_w1665_,
		_w1666_,
		_w1667_,
		_w1668_
	);
	LUT4 #(
		.INIT('h8000)
	) name1364 (
		_w1663_,
		_w1668_,
		_w1653_,
		_w1658_,
		_w1669_
	);
	LUT2 #(
		.INIT('h6)
	) name1365 (
		_w1111_,
		_w1669_,
		_w1670_
	);
	LUT3 #(
		.INIT('ha8)
	) name1366 (
		_w305_,
		_w753_,
		_w774_,
		_w1671_
	);
	LUT3 #(
		.INIT('ha8)
	) name1367 (
		_w343_,
		_w702_,
		_w671_,
		_w1672_
	);
	LUT3 #(
		.INIT('ha8)
	) name1368 (
		_w398_,
		_w681_,
		_w809_,
		_w1673_
	);
	LUT3 #(
		.INIT('ha8)
	) name1369 (
		_w312_,
		_w703_,
		_w793_,
		_w1674_
	);
	LUT4 #(
		.INIT('h0001)
	) name1370 (
		_w1671_,
		_w1672_,
		_w1673_,
		_w1674_,
		_w1675_
	);
	LUT3 #(
		.INIT('ha8)
	) name1371 (
		_w419_,
		_w669_,
		_w811_,
		_w1676_
	);
	LUT3 #(
		.INIT('ha8)
	) name1372 (
		_w363_,
		_w758_,
		_w724_,
		_w1677_
	);
	LUT3 #(
		.INIT('ha8)
	) name1373 (
		_w423_,
		_w759_,
		_w739_,
		_w1678_
	);
	LUT3 #(
		.INIT('ha8)
	) name1374 (
		_w415_,
		_w696_,
		_w717_,
		_w1679_
	);
	LUT4 #(
		.INIT('h0001)
	) name1375 (
		_w1676_,
		_w1677_,
		_w1678_,
		_w1679_,
		_w1680_
	);
	LUT3 #(
		.INIT('ha8)
	) name1376 (
		_w333_,
		_w708_,
		_w721_,
		_w1681_
	);
	LUT3 #(
		.INIT('ha8)
	) name1377 (
		_w402_,
		_w734_,
		_w767_,
		_w1682_
	);
	LUT3 #(
		.INIT('ha8)
	) name1378 (
		_w373_,
		_w665_,
		_w677_,
		_w1683_
	);
	LUT3 #(
		.INIT('ha8)
	) name1379 (
		_w388_,
		_w752_,
		_w755_,
		_w1684_
	);
	LUT4 #(
		.INIT('h0001)
	) name1380 (
		_w1681_,
		_w1682_,
		_w1683_,
		_w1684_,
		_w1685_
	);
	LUT3 #(
		.INIT('ha8)
	) name1381 (
		_w406_,
		_w746_,
		_w730_,
		_w1686_
	);
	LUT3 #(
		.INIT('ha8)
	) name1382 (
		_w323_,
		_w750_,
		_w736_,
		_w1687_
	);
	LUT3 #(
		.INIT('ha8)
	) name1383 (
		_w377_,
		_w672_,
		_w779_,
		_w1688_
	);
	LUT3 #(
		.INIT('ha8)
	) name1384 (
		_w411_,
		_w686_,
		_w756_,
		_w1689_
	);
	LUT4 #(
		.INIT('h0001)
	) name1385 (
		_w1686_,
		_w1687_,
		_w1688_,
		_w1689_,
		_w1690_
	);
	LUT4 #(
		.INIT('h8000)
	) name1386 (
		_w1685_,
		_w1690_,
		_w1675_,
		_w1680_,
		_w1691_
	);
	LUT2 #(
		.INIT('h9)
	) name1387 (
		_w1413_,
		_w1691_,
		_w1692_
	);
	LUT3 #(
		.INIT('ha8)
	) name1388 (
		_w363_,
		_w837_,
		_w811_,
		_w1693_
	);
	LUT3 #(
		.INIT('ha8)
	) name1389 (
		_w377_,
		_w696_,
		_w831_,
		_w1694_
	);
	LUT3 #(
		.INIT('ha8)
	) name1390 (
		_w343_,
		_w786_,
		_w797_,
		_w1695_
	);
	LUT3 #(
		.INIT('ha8)
	) name1391 (
		_w423_,
		_w842_,
		_w774_,
		_w1696_
	);
	LUT4 #(
		.INIT('h0001)
	) name1392 (
		_w1693_,
		_w1694_,
		_w1695_,
		_w1696_,
		_w1697_
	);
	LUT3 #(
		.INIT('ha8)
	) name1393 (
		_w411_,
		_w860_,
		_w809_,
		_w1698_
	);
	LUT3 #(
		.INIT('ha8)
	) name1394 (
		_w305_,
		_w690_,
		_w739_,
		_w1699_
	);
	LUT3 #(
		.INIT('ha8)
	) name1395 (
		_w402_,
		_w708_,
		_w737_,
		_w1700_
	);
	LUT3 #(
		.INIT('ha8)
	) name1396 (
		_w323_,
		_w824_,
		_w793_,
		_w1701_
	);
	LUT4 #(
		.INIT('h0001)
	) name1397 (
		_w1698_,
		_w1699_,
		_w1700_,
		_w1701_,
		_w1702_
	);
	LUT3 #(
		.INIT('ha8)
	) name1398 (
		_w398_,
		_w686_,
		_w856_,
		_w1703_
	);
	LUT3 #(
		.INIT('ha8)
	) name1399 (
		_w419_,
		_w724_,
		_w849_,
		_w1704_
	);
	LUT3 #(
		.INIT('ha8)
	) name1400 (
		_w415_,
		_w858_,
		_w779_,
		_w1705_
	);
	LUT3 #(
		.INIT('ha8)
	) name1401 (
		_w312_,
		_w736_,
		_w865_,
		_w1706_
	);
	LUT4 #(
		.INIT('h0001)
	) name1402 (
		_w1703_,
		_w1704_,
		_w1705_,
		_w1706_,
		_w1707_
	);
	LUT3 #(
		.INIT('ha8)
	) name1403 (
		_w406_,
		_w802_,
		_w847_,
		_w1708_
	);
	LUT3 #(
		.INIT('ha8)
	) name1404 (
		_w373_,
		_w788_,
		_w772_,
		_w1709_
	);
	LUT3 #(
		.INIT('ha8)
	) name1405 (
		_w333_,
		_w767_,
		_w863_,
		_w1710_
	);
	LUT3 #(
		.INIT('ha8)
	) name1406 (
		_w388_,
		_w868_,
		_w806_,
		_w1711_
	);
	LUT4 #(
		.INIT('h0001)
	) name1407 (
		_w1708_,
		_w1709_,
		_w1710_,
		_w1711_,
		_w1712_
	);
	LUT4 #(
		.INIT('h8000)
	) name1408 (
		_w1707_,
		_w1712_,
		_w1697_,
		_w1702_,
		_w1713_
	);
	LUT4 #(
		.INIT('h0200)
	) name1409 (
		\desIn[57]_pad ,
		\roundSel[4]_pad ,
		\roundSel[5]_pad ,
		_w305_,
		_w1714_
	);
	LUT4 #(
		.INIT('h4155)
	) name1410 (
		\FP_R_reg[32]/P0001 ,
		\roundSel[4]_pad ,
		\roundSel[5]_pad ,
		_w305_,
		_w1715_
	);
	LUT4 #(
		.INIT('he8ff)
	) name1411 (
		\FP_R_reg[64]/NET0131 ,
		\roundSel[4]_pad ,
		\roundSel[5]_pad ,
		_w305_,
		_w1716_
	);
	LUT3 #(
		.INIT('h45)
	) name1412 (
		_w1714_,
		_w1715_,
		_w1716_,
		_w1717_
	);
	LUT3 #(
		.INIT('hba)
	) name1413 (
		_w1714_,
		_w1715_,
		_w1716_,
		_w1718_
	);
	LUT2 #(
		.INIT('h9)
	) name1414 (
		_w1713_,
		_w1717_,
		_w1719_
	);
	LUT3 #(
		.INIT('ha8)
	) name1415 (
		_w343_,
		_w669_,
		_w753_,
		_w1720_
	);
	LUT3 #(
		.INIT('ha8)
	) name1416 (
		_w377_,
		_w677_,
		_w860_,
		_w1721_
	);
	LUT3 #(
		.INIT('ha8)
	) name1417 (
		_w402_,
		_w665_,
		_w837_,
		_w1722_
	);
	LUT3 #(
		.INIT('ha8)
	) name1418 (
		_w323_,
		_w759_,
		_w849_,
		_w1723_
	);
	LUT4 #(
		.INIT('h0001)
	) name1419 (
		_w1720_,
		_w1721_,
		_w1722_,
		_w1723_,
		_w1724_
	);
	LUT3 #(
		.INIT('ha8)
	) name1420 (
		_w312_,
		_w755_,
		_w856_,
		_w1725_
	);
	LUT3 #(
		.INIT('ha8)
	) name1421 (
		_w419_,
		_w702_,
		_w824_,
		_w1726_
	);
	LUT3 #(
		.INIT('ha8)
	) name1422 (
		_w333_,
		_w756_,
		_w725_,
		_w1727_
	);
	LUT3 #(
		.INIT('ha8)
	) name1423 (
		_w388_,
		_w703_,
		_w712_,
		_w1728_
	);
	LUT4 #(
		.INIT('h0001)
	) name1424 (
		_w1725_,
		_w1726_,
		_w1727_,
		_w1728_,
		_w1729_
	);
	LUT3 #(
		.INIT('ha8)
	) name1425 (
		_w363_,
		_w717_,
		_w737_,
		_w1730_
	);
	LUT3 #(
		.INIT('ha8)
	) name1426 (
		_w305_,
		_w671_,
		_w858_,
		_w1731_
	);
	LUT3 #(
		.INIT('ha8)
	) name1427 (
		_w411_,
		_w721_,
		_w831_,
		_w1732_
	);
	LUT3 #(
		.INIT('ha8)
	) name1428 (
		_w423_,
		_w700_,
		_w750_,
		_w1733_
	);
	LUT4 #(
		.INIT('h0001)
	) name1429 (
		_w1730_,
		_w1731_,
		_w1732_,
		_w1733_,
		_w1734_
	);
	LUT3 #(
		.INIT('ha8)
	) name1430 (
		_w398_,
		_w746_,
		_w865_,
		_w1735_
	);
	LUT3 #(
		.INIT('ha8)
	) name1431 (
		_w406_,
		_w681_,
		_w740_,
		_w1736_
	);
	LUT3 #(
		.INIT('ha8)
	) name1432 (
		_w415_,
		_w690_,
		_w758_,
		_w1737_
	);
	LUT3 #(
		.INIT('ha8)
	) name1433 (
		_w373_,
		_w672_,
		_w734_,
		_w1738_
	);
	LUT4 #(
		.INIT('h0001)
	) name1434 (
		_w1735_,
		_w1736_,
		_w1737_,
		_w1738_,
		_w1739_
	);
	LUT4 #(
		.INIT('h8000)
	) name1435 (
		_w1734_,
		_w1739_,
		_w1724_,
		_w1729_,
		_w1740_
	);
	LUT3 #(
		.INIT('h40)
	) name1436 (
		\FP_R_reg[33]/NET0131 ,
		_w305_,
		_w307_,
		_w1741_
	);
	LUT4 #(
		.INIT('hb0aa)
	) name1437 (
		\FP_R_reg[1]/P0001 ,
		\roundSel[4]_pad ,
		\roundSel[5]_pad ,
		_w305_,
		_w1742_
	);
	LUT4 #(
		.INIT('h0800)
	) name1438 (
		\FP_R_reg[33]/NET0131 ,
		\roundSel[4]_pad ,
		\roundSel[5]_pad ,
		_w305_,
		_w1743_
	);
	LUT4 #(
		.INIT('h0200)
	) name1439 (
		\desIn[7]_pad ,
		\roundSel[4]_pad ,
		\roundSel[5]_pad ,
		_w305_,
		_w1744_
	);
	LUT4 #(
		.INIT('h1011)
	) name1440 (
		_w1743_,
		_w1744_,
		_w1741_,
		_w1742_,
		_w1745_
	);
	LUT4 #(
		.INIT('hefee)
	) name1441 (
		_w1743_,
		_w1744_,
		_w1741_,
		_w1742_,
		_w1746_
	);
	LUT2 #(
		.INIT('h9)
	) name1442 (
		_w1740_,
		_w1745_,
		_w1747_
	);
	LUT3 #(
		.INIT('ha8)
	) name1443 (
		_w323_,
		_w681_,
		_w724_,
		_w1748_
	);
	LUT3 #(
		.INIT('ha8)
	) name1444 (
		_w402_,
		_w740_,
		_w811_,
		_w1749_
	);
	LUT3 #(
		.INIT('ha8)
	) name1445 (
		_w343_,
		_w677_,
		_w755_,
		_w1750_
	);
	LUT3 #(
		.INIT('ha8)
	) name1446 (
		_w363_,
		_w708_,
		_w750_,
		_w1751_
	);
	LUT4 #(
		.INIT('h0001)
	) name1447 (
		_w1748_,
		_w1749_,
		_w1750_,
		_w1751_,
		_w1752_
	);
	LUT3 #(
		.INIT('ha8)
	) name1448 (
		_w373_,
		_w702_,
		_w746_,
		_w1753_
	);
	LUT3 #(
		.INIT('ha8)
	) name1449 (
		_w312_,
		_w669_,
		_w686_,
		_w1754_
	);
	LUT3 #(
		.INIT('ha8)
	) name1450 (
		_w406_,
		_w665_,
		_w759_,
		_w1755_
	);
	LUT3 #(
		.INIT('ha8)
	) name1451 (
		_w415_,
		_w756_,
		_w739_,
		_w1756_
	);
	LUT4 #(
		.INIT('h0001)
	) name1452 (
		_w1753_,
		_w1754_,
		_w1755_,
		_w1756_,
		_w1757_
	);
	LUT3 #(
		.INIT('ha8)
	) name1453 (
		_w305_,
		_w712_,
		_w779_,
		_w1758_
	);
	LUT3 #(
		.INIT('ha8)
	) name1454 (
		_w423_,
		_w717_,
		_w730_,
		_w1759_
	);
	LUT3 #(
		.INIT('ha8)
	) name1455 (
		_w411_,
		_w696_,
		_w703_,
		_w1760_
	);
	LUT3 #(
		.INIT('ha8)
	) name1456 (
		_w377_,
		_w753_,
		_w809_,
		_w1761_
	);
	LUT4 #(
		.INIT('h0001)
	) name1457 (
		_w1758_,
		_w1759_,
		_w1760_,
		_w1761_,
		_w1762_
	);
	LUT3 #(
		.INIT('ha8)
	) name1458 (
		_w388_,
		_w721_,
		_w671_,
		_w1763_
	);
	LUT3 #(
		.INIT('ha8)
	) name1459 (
		_w398_,
		_w672_,
		_w736_,
		_w1764_
	);
	LUT3 #(
		.INIT('ha8)
	) name1460 (
		_w333_,
		_w752_,
		_w758_,
		_w1765_
	);
	LUT3 #(
		.INIT('ha8)
	) name1461 (
		_w419_,
		_w734_,
		_w793_,
		_w1766_
	);
	LUT4 #(
		.INIT('h0001)
	) name1462 (
		_w1763_,
		_w1764_,
		_w1765_,
		_w1766_,
		_w1767_
	);
	LUT4 #(
		.INIT('h8000)
	) name1463 (
		_w1762_,
		_w1767_,
		_w1752_,
		_w1757_,
		_w1768_
	);
	LUT2 #(
		.INIT('h6)
	) name1464 (
		_w1202_,
		_w1768_,
		_w1769_
	);
	LUT4 #(
		.INIT('h1428)
	) name1465 (
		_w1202_,
		_w1740_,
		_w1745_,
		_w1768_,
		_w1770_
	);
	LUT3 #(
		.INIT('ha8)
	) name1466 (
		_w411_,
		_w671_,
		_w797_,
		_w1771_
	);
	LUT3 #(
		.INIT('ha8)
	) name1467 (
		_w377_,
		_w755_,
		_w868_,
		_w1772_
	);
	LUT3 #(
		.INIT('ha8)
	) name1468 (
		_w343_,
		_w686_,
		_w809_,
		_w1773_
	);
	LUT3 #(
		.INIT('ha8)
	) name1469 (
		_w323_,
		_w665_,
		_w772_,
		_w1774_
	);
	LUT4 #(
		.INIT('h0001)
	) name1470 (
		_w1771_,
		_w1772_,
		_w1773_,
		_w1774_,
		_w1775_
	);
	LUT3 #(
		.INIT('ha8)
	) name1471 (
		_w423_,
		_w708_,
		_w767_,
		_w1776_
	);
	LUT3 #(
		.INIT('ha8)
	) name1472 (
		_w402_,
		_w759_,
		_w842_,
		_w1777_
	);
	LUT3 #(
		.INIT('ha8)
	) name1473 (
		_w305_,
		_w721_,
		_w863_,
		_w1778_
	);
	LUT3 #(
		.INIT('ha8)
	) name1474 (
		_w363_,
		_w730_,
		_w802_,
		_w1779_
	);
	LUT4 #(
		.INIT('h0001)
	) name1475 (
		_w1776_,
		_w1777_,
		_w1778_,
		_w1779_,
		_w1780_
	);
	LUT3 #(
		.INIT('ha8)
	) name1476 (
		_w388_,
		_w696_,
		_w779_,
		_w1781_
	);
	LUT3 #(
		.INIT('ha8)
	) name1477 (
		_w419_,
		_w746_,
		_w847_,
		_w1782_
	);
	LUT3 #(
		.INIT('ha8)
	) name1478 (
		_w398_,
		_w702_,
		_w786_,
		_w1783_
	);
	LUT3 #(
		.INIT('ha8)
	) name1479 (
		_w312_,
		_w677_,
		_w788_,
		_w1784_
	);
	LUT4 #(
		.INIT('h0001)
	) name1480 (
		_w1781_,
		_w1782_,
		_w1783_,
		_w1784_,
		_w1785_
	);
	LUT3 #(
		.INIT('ha8)
	) name1481 (
		_w373_,
		_w736_,
		_w793_,
		_w1786_
	);
	LUT3 #(
		.INIT('ha8)
	) name1482 (
		_w415_,
		_w752_,
		_w806_,
		_w1787_
	);
	LUT3 #(
		.INIT('ha8)
	) name1483 (
		_w406_,
		_w724_,
		_w811_,
		_w1788_
	);
	LUT3 #(
		.INIT('ha8)
	) name1484 (
		_w333_,
		_w739_,
		_w774_,
		_w1789_
	);
	LUT4 #(
		.INIT('h0001)
	) name1485 (
		_w1786_,
		_w1787_,
		_w1788_,
		_w1789_,
		_w1790_
	);
	LUT4 #(
		.INIT('h8000)
	) name1486 (
		_w1785_,
		_w1790_,
		_w1775_,
		_w1780_,
		_w1791_
	);
	LUT2 #(
		.INIT('h9)
	) name1487 (
		_w1057_,
		_w1791_,
		_w1792_
	);
	LUT4 #(
		.INIT('h8241)
	) name1488 (
		_w1057_,
		_w1713_,
		_w1717_,
		_w1791_,
		_w1793_
	);
	LUT2 #(
		.INIT('h8)
	) name1489 (
		_w1793_,
		_w1770_,
		_w1794_
	);
	LUT4 #(
		.INIT('ha022)
	) name1490 (
		_w1692_,
		_w1719_,
		_w1793_,
		_w1770_,
		_w1795_
	);
	LUT4 #(
		.INIT('h0144)
	) name1491 (
		_w1692_,
		_w1719_,
		_w1747_,
		_w1769_,
		_w1796_
	);
	LUT4 #(
		.INIT('h8241)
	) name1492 (
		_w1202_,
		_w1740_,
		_w1745_,
		_w1768_,
		_w1797_
	);
	LUT4 #(
		.INIT('h9009)
	) name1493 (
		_w1713_,
		_w1717_,
		_w1740_,
		_w1745_,
		_w1798_
	);
	LUT3 #(
		.INIT('h40)
	) name1494 (
		_w1792_,
		_w1769_,
		_w1798_,
		_w1799_
	);
	LUT4 #(
		.INIT('hf73f)
	) name1495 (
		_w1719_,
		_w1747_,
		_w1792_,
		_w1769_,
		_w1800_
	);
	LUT4 #(
		.INIT('h5455)
	) name1496 (
		_w1670_,
		_w1795_,
		_w1796_,
		_w1800_,
		_w1801_
	);
	LUT4 #(
		.INIT('h1428)
	) name1497 (
		_w1057_,
		_w1740_,
		_w1745_,
		_w1791_,
		_w1802_
	);
	LUT4 #(
		.INIT('h8008)
	) name1498 (
		_w1692_,
		_w1719_,
		_w1747_,
		_w1792_,
		_w1803_
	);
	LUT4 #(
		.INIT('h2814)
	) name1499 (
		_w1057_,
		_w1713_,
		_w1717_,
		_w1791_,
		_w1804_
	);
	LUT4 #(
		.INIT('h0018)
	) name1500 (
		_w1719_,
		_w1747_,
		_w1792_,
		_w1769_,
		_w1805_
	);
	LUT3 #(
		.INIT('ha8)
	) name1501 (
		_w1670_,
		_w1803_,
		_w1805_,
		_w1806_
	);
	LUT4 #(
		.INIT('h1248)
	) name1502 (
		_w1111_,
		_w1413_,
		_w1669_,
		_w1691_,
		_w1807_
	);
	LUT4 #(
		.INIT('h1428)
	) name1503 (
		_w1057_,
		_w1713_,
		_w1717_,
		_w1791_,
		_w1808_
	);
	LUT4 #(
		.INIT('hdade)
	) name1504 (
		_w1719_,
		_w1747_,
		_w1792_,
		_w1769_,
		_w1809_
	);
	LUT4 #(
		.INIT('h4182)
	) name1505 (
		_w1202_,
		_w1740_,
		_w1745_,
		_w1768_,
		_w1810_
	);
	LUT4 #(
		.INIT('h0990)
	) name1506 (
		_w1413_,
		_w1691_,
		_w1713_,
		_w1717_,
		_w1811_
	);
	LUT4 #(
		.INIT('he400)
	) name1507 (
		_w1792_,
		_w1797_,
		_w1810_,
		_w1811_,
		_w1812_
	);
	LUT3 #(
		.INIT('h0d)
	) name1508 (
		_w1807_,
		_w1809_,
		_w1812_,
		_w1813_
	);
	LUT4 #(
		.INIT('h0100)
	) name1509 (
		\desIn[2]_pad ,
		\roundSel[4]_pad ,
		\roundSel[5]_pad ,
		_w305_,
		_w1814_
	);
	LUT4 #(
		.INIT('h2800)
	) name1510 (
		\FP_R_reg[17]/P0001 ,
		\roundSel[4]_pad ,
		\roundSel[5]_pad ,
		_w305_,
		_w1815_
	);
	LUT4 #(
		.INIT('h7c55)
	) name1511 (
		\FP_R_reg[49]/NET0131 ,
		\roundSel[4]_pad ,
		\roundSel[5]_pad ,
		_w305_,
		_w1816_
	);
	LUT3 #(
		.INIT('h45)
	) name1512 (
		_w1814_,
		_w1815_,
		_w1816_,
		_w1817_
	);
	LUT4 #(
		.INIT('h10ef)
	) name1513 (
		_w1806_,
		_w1801_,
		_w1813_,
		_w1817_,
		_w1818_
	);
	LUT3 #(
		.INIT('h20)
	) name1514 (
		_w1331_,
		_w1301_,
		_w1379_,
		_w1819_
	);
	LUT4 #(
		.INIT('he65f)
	) name1515 (
		_w1279_,
		_w1331_,
		_w1301_,
		_w1257_,
		_w1820_
	);
	LUT3 #(
		.INIT('h80)
	) name1516 (
		_w1331_,
		_w1257_,
		_w1364_,
		_w1821_
	);
	LUT4 #(
		.INIT('hfbaf)
	) name1517 (
		_w1279_,
		_w1331_,
		_w1301_,
		_w1257_,
		_w1822_
	);
	LUT4 #(
		.INIT('h1428)
	) name1518 (
		_w568_,
		_w1325_,
		_w1329_,
		_w1300_,
		_w1823_
	);
	LUT4 #(
		.INIT('h5d7f)
	) name1519 (
		_w1279_,
		_w1257_,
		_w1377_,
		_w1823_,
		_w1824_
	);
	LUT4 #(
		.INIT('he400)
	) name1520 (
		_w1230_,
		_w1822_,
		_w1820_,
		_w1824_,
		_w1825_
	);
	LUT4 #(
		.INIT('h0660)
	) name1521 (
		_w310_,
		_w1278_,
		_w1325_,
		_w1329_,
		_w1826_
	);
	LUT4 #(
		.INIT('h3310)
	) name1522 (
		_w1257_,
		_w1230_,
		_w1332_,
		_w1826_,
		_w1827_
	);
	LUT3 #(
		.INIT('h10)
	) name1523 (
		_w1279_,
		_w1257_,
		_w1332_,
		_w1828_
	);
	LUT4 #(
		.INIT('h2777)
	) name1524 (
		_w1331_,
		_w1334_,
		_w1230_,
		_w1379_,
		_w1829_
	);
	LUT3 #(
		.INIT('h10)
	) name1525 (
		_w1828_,
		_w1827_,
		_w1829_,
		_w1830_
	);
	LUT4 #(
		.INIT('h9009)
	) name1526 (
		_w1325_,
		_w1329_,
		_w1207_,
		_w1229_,
		_w1831_
	);
	LUT4 #(
		.INIT('h4900)
	) name1527 (
		_w1279_,
		_w1301_,
		_w1257_,
		_w1831_,
		_w1832_
	);
	LUT2 #(
		.INIT('h8)
	) name1528 (
		_w1301_,
		_w1379_,
		_w1833_
	);
	LUT4 #(
		.INIT('h028a)
	) name1529 (
		_w1331_,
		_w1301_,
		_w1378_,
		_w1379_,
		_w1834_
	);
	LUT3 #(
		.INIT('h32)
	) name1530 (
		_w1331_,
		_w1230_,
		_w1303_,
		_w1835_
	);
	LUT3 #(
		.INIT('h45)
	) name1531 (
		_w1832_,
		_w1834_,
		_w1835_,
		_w1836_
	);
	LUT4 #(
		.INIT('he400)
	) name1532 (
		_w1361_,
		_w1825_,
		_w1830_,
		_w1836_,
		_w1837_
	);
	LUT4 #(
		.INIT('h0100)
	) name1533 (
		\desIn[30]_pad ,
		\roundSel[4]_pad ,
		\roundSel[5]_pad ,
		_w305_,
		_w1838_
	);
	LUT4 #(
		.INIT('h2800)
	) name1534 (
		\FP_R_reg[4]/P0001 ,
		\roundSel[4]_pad ,
		\roundSel[5]_pad ,
		_w305_,
		_w1839_
	);
	LUT4 #(
		.INIT('h7c55)
	) name1535 (
		\FP_R_reg[36]/NET0131 ,
		\roundSel[4]_pad ,
		\roundSel[5]_pad ,
		_w305_,
		_w1840_
	);
	LUT3 #(
		.INIT('h45)
	) name1536 (
		_w1838_,
		_w1839_,
		_w1840_,
		_w1841_
	);
	LUT2 #(
		.INIT('h9)
	) name1537 (
		_w1837_,
		_w1841_,
		_w1842_
	);
	LUT3 #(
		.INIT('h80)
	) name1538 (
		_w1331_,
		_w1301_,
		_w1378_,
		_w1843_
	);
	LUT2 #(
		.INIT('h2)
	) name1539 (
		_w1302_,
		_w1370_,
		_w1844_
	);
	LUT3 #(
		.INIT('ha8)
	) name1540 (
		_w1230_,
		_w1843_,
		_w1844_,
		_w1845_
	);
	LUT4 #(
		.INIT('h7f7a)
	) name1541 (
		_w1279_,
		_w1331_,
		_w1257_,
		_w1332_,
		_w1846_
	);
	LUT2 #(
		.INIT('h1)
	) name1542 (
		_w1230_,
		_w1846_,
		_w1847_
	);
	LUT2 #(
		.INIT('h8)
	) name1543 (
		_w1377_,
		_w1378_,
		_w1848_
	);
	LUT3 #(
		.INIT('h01)
	) name1544 (
		_w1372_,
		_w1819_,
		_w1848_,
		_w1849_
	);
	LUT4 #(
		.INIT('ha8aa)
	) name1545 (
		_w1361_,
		_w1845_,
		_w1847_,
		_w1849_,
		_w1850_
	);
	LUT4 #(
		.INIT('h5fb4)
	) name1546 (
		_w1279_,
		_w1331_,
		_w1301_,
		_w1257_,
		_w1851_
	);
	LUT4 #(
		.INIT('hcd6f)
	) name1547 (
		_w1279_,
		_w1331_,
		_w1301_,
		_w1257_,
		_w1852_
	);
	LUT4 #(
		.INIT('h3120)
	) name1548 (
		_w1230_,
		_w1821_,
		_w1851_,
		_w1852_,
		_w1853_
	);
	LUT4 #(
		.INIT('h0777)
	) name1549 (
		_w1334_,
		_w1375_,
		_w1378_,
		_w1823_,
		_w1854_
	);
	LUT3 #(
		.INIT('he0)
	) name1550 (
		_w1361_,
		_w1853_,
		_w1854_,
		_w1855_
	);
	LUT4 #(
		.INIT('h0100)
	) name1551 (
		\desIn[32]_pad ,
		\roundSel[4]_pad ,
		\roundSel[5]_pad ,
		_w305_,
		_w1856_
	);
	LUT4 #(
		.INIT('h2800)
	) name1552 (
		\FP_R_reg[29]/P0001 ,
		\roundSel[4]_pad ,
		\roundSel[5]_pad ,
		_w305_,
		_w1857_
	);
	LUT4 #(
		.INIT('h7c55)
	) name1553 (
		\FP_R_reg[61]/NET0131 ,
		\roundSel[4]_pad ,
		\roundSel[5]_pad ,
		_w305_,
		_w1858_
	);
	LUT3 #(
		.INIT('h45)
	) name1554 (
		_w1856_,
		_w1857_,
		_w1858_,
		_w1859_
	);
	LUT3 #(
		.INIT('hb4)
	) name1555 (
		_w1850_,
		_w1855_,
		_w1859_,
		_w1860_
	);
	LUT3 #(
		.INIT('hc8)
	) name1556 (
		_w371_,
		_w419_,
		_w478_,
		_w1861_
	);
	LUT3 #(
		.INIT('ha8)
	) name1557 (
		_w377_,
		_w417_,
		_w492_,
		_w1862_
	);
	LUT3 #(
		.INIT('ha8)
	) name1558 (
		_w333_,
		_w404_,
		_w480_,
		_w1863_
	);
	LUT3 #(
		.INIT('ha8)
	) name1559 (
		_w411_,
		_w400_,
		_w455_,
		_w1864_
	);
	LUT4 #(
		.INIT('h0001)
	) name1560 (
		_w1861_,
		_w1862_,
		_w1863_,
		_w1864_,
		_w1865_
	);
	LUT3 #(
		.INIT('hc8)
	) name1561 (
		_w321_,
		_w323_,
		_w457_,
		_w1866_
	);
	LUT3 #(
		.INIT('ha8)
	) name1562 (
		_w363_,
		_w421_,
		_w473_,
		_w1867_
	);
	LUT3 #(
		.INIT('hc8)
	) name1563 (
		_w413_,
		_w398_,
		_w488_,
		_w1868_
	);
	LUT3 #(
		.INIT('hc8)
	) name1564 (
		_w361_,
		_w423_,
		_w449_,
		_w1869_
	);
	LUT4 #(
		.INIT('h0001)
	) name1565 (
		_w1866_,
		_w1867_,
		_w1868_,
		_w1869_,
		_w1870_
	);
	LUT3 #(
		.INIT('hc8)
	) name1566 (
		_w385_,
		_w415_,
		_w471_,
		_w1871_
	);
	LUT3 #(
		.INIT('ha8)
	) name1567 (
		_w343_,
		_w548_,
		_w553_,
		_w1872_
	);
	LUT3 #(
		.INIT('ha8)
	) name1568 (
		_w373_,
		_w556_,
		_w561_,
		_w1873_
	);
	LUT3 #(
		.INIT('ha8)
	) name1569 (
		_w388_,
		_w433_,
		_w539_,
		_w1874_
	);
	LUT4 #(
		.INIT('h0001)
	) name1570 (
		_w1871_,
		_w1872_,
		_w1873_,
		_w1874_,
		_w1875_
	);
	LUT3 #(
		.INIT('ha8)
	) name1571 (
		_w305_,
		_w425_,
		_w483_,
		_w1876_
	);
	LUT3 #(
		.INIT('hc8)
	) name1572 (
		_w341_,
		_w402_,
		_w465_,
		_w1877_
	);
	LUT3 #(
		.INIT('ha8)
	) name1573 (
		_w406_,
		_w435_,
		_w559_,
		_w1878_
	);
	LUT3 #(
		.INIT('ha8)
	) name1574 (
		_w312_,
		_w331_,
		_w490_,
		_w1879_
	);
	LUT4 #(
		.INIT('h0001)
	) name1575 (
		_w1876_,
		_w1877_,
		_w1878_,
		_w1879_,
		_w1880_
	);
	LUT4 #(
		.INIT('h8000)
	) name1576 (
		_w1875_,
		_w1880_,
		_w1865_,
		_w1870_,
		_w1881_
	);
	LUT2 #(
		.INIT('h9)
	) name1577 (
		_w1717_,
		_w1881_,
		_w1882_
	);
	LUT3 #(
		.INIT('hc8)
	) name1578 (
		_w371_,
		_w343_,
		_w425_,
		_w1883_
	);
	LUT3 #(
		.INIT('ha8)
	) name1579 (
		_w305_,
		_w327_,
		_w553_,
		_w1884_
	);
	LUT3 #(
		.INIT('hc8)
	) name1580 (
		_w361_,
		_w323_,
		_w396_,
		_w1885_
	);
	LUT3 #(
		.INIT('ha8)
	) name1581 (
		_w411_,
		_w404_,
		_w407_,
		_w1886_
	);
	LUT4 #(
		.INIT('h0001)
	) name1582 (
		_w1883_,
		_w1884_,
		_w1885_,
		_w1886_,
		_w1887_
	);
	LUT3 #(
		.INIT('ha8)
	) name1583 (
		_w363_,
		_w385_,
		_w351_,
		_w1888_
	);
	LUT3 #(
		.INIT('hc8)
	) name1584 (
		_w367_,
		_w377_,
		_w556_,
		_w1889_
	);
	LUT3 #(
		.INIT('hc8)
	) name1585 (
		_w412_,
		_w402_,
		_w561_,
		_w1890_
	);
	LUT3 #(
		.INIT('he0)
	) name1586 (
		_w321_,
		_w347_,
		_w423_,
		_w1891_
	);
	LUT4 #(
		.INIT('h0001)
	) name1587 (
		_w1888_,
		_w1889_,
		_w1890_,
		_w1891_,
		_w1892_
	);
	LUT3 #(
		.INIT('hc8)
	) name1588 (
		_w337_,
		_w398_,
		_w559_,
		_w1893_
	);
	LUT3 #(
		.INIT('hc8)
	) name1589 (
		_w416_,
		_w419_,
		_w548_,
		_w1894_
	);
	LUT3 #(
		.INIT('he0)
	) name1590 (
		_w413_,
		_w392_,
		_w406_,
		_w1895_
	);
	LUT3 #(
		.INIT('hc8)
	) name1591 (
		_w331_,
		_w388_,
		_w408_,
		_w1896_
	);
	LUT4 #(
		.INIT('h0001)
	) name1592 (
		_w1893_,
		_w1894_,
		_w1895_,
		_w1896_,
		_w1897_
	);
	LUT3 #(
		.INIT('ha8)
	) name1593 (
		_w373_,
		_w341_,
		_w417_,
		_w1898_
	);
	LUT3 #(
		.INIT('ha8)
	) name1594 (
		_w312_,
		_w424_,
		_w539_,
		_w1899_
	);
	LUT3 #(
		.INIT('hc8)
	) name1595 (
		_w375_,
		_w333_,
		_w400_,
		_w1900_
	);
	LUT3 #(
		.INIT('hc8)
	) name1596 (
		_w374_,
		_w415_,
		_w421_,
		_w1901_
	);
	LUT4 #(
		.INIT('h0001)
	) name1597 (
		_w1898_,
		_w1899_,
		_w1900_,
		_w1901_,
		_w1902_
	);
	LUT4 #(
		.INIT('h8000)
	) name1598 (
		_w1897_,
		_w1902_,
		_w1887_,
		_w1892_,
		_w1903_
	);
	LUT4 #(
		.INIT('h0200)
	) name1599 (
		\desIn[49]_pad ,
		\roundSel[4]_pad ,
		\roundSel[5]_pad ,
		_w305_,
		_w1904_
	);
	LUT4 #(
		.INIT('h4155)
	) name1600 (
		\FP_R_reg[31]/P0001 ,
		\roundSel[4]_pad ,
		\roundSel[5]_pad ,
		_w305_,
		_w1905_
	);
	LUT4 #(
		.INIT('he8ff)
	) name1601 (
		\FP_R_reg[63]/NET0131 ,
		\roundSel[4]_pad ,
		\roundSel[5]_pad ,
		_w305_,
		_w1906_
	);
	LUT3 #(
		.INIT('h45)
	) name1602 (
		_w1904_,
		_w1905_,
		_w1906_,
		_w1907_
	);
	LUT3 #(
		.INIT('hba)
	) name1603 (
		_w1904_,
		_w1905_,
		_w1906_,
		_w1908_
	);
	LUT2 #(
		.INIT('h9)
	) name1604 (
		_w1903_,
		_w1907_,
		_w1909_
	);
	LUT3 #(
		.INIT('he0)
	) name1605 (
		_w381_,
		_w331_,
		_w398_,
		_w1910_
	);
	LUT3 #(
		.INIT('ha8)
	) name1606 (
		_w305_,
		_w385_,
		_w460_,
		_w1911_
	);
	LUT3 #(
		.INIT('ha8)
	) name1607 (
		_w312_,
		_w413_,
		_w420_,
		_w1912_
	);
	LUT3 #(
		.INIT('hc8)
	) name1608 (
		_w416_,
		_w423_,
		_w408_,
		_w1913_
	);
	LUT4 #(
		.INIT('h0001)
	) name1609 (
		_w1910_,
		_w1911_,
		_w1912_,
		_w1913_,
		_w1914_
	);
	LUT3 #(
		.INIT('hc8)
	) name1610 (
		_w371_,
		_w323_,
		_w399_,
		_w1915_
	);
	LUT3 #(
		.INIT('hc8)
	) name1611 (
		_w421_,
		_w402_,
		_w440_,
		_w1916_
	);
	LUT3 #(
		.INIT('hc8)
	) name1612 (
		_w321_,
		_w419_,
		_w403_,
		_w1917_
	);
	LUT3 #(
		.INIT('ha8)
	) name1613 (
		_w373_,
		_w351_,
		_w407_,
		_w1918_
	);
	LUT4 #(
		.INIT('h0001)
	) name1614 (
		_w1915_,
		_w1916_,
		_w1917_,
		_w1918_,
		_w1919_
	);
	LUT3 #(
		.INIT('ha8)
	) name1615 (
		_w363_,
		_w327_,
		_w341_,
		_w1920_
	);
	LUT3 #(
		.INIT('hc8)
	) name1616 (
		_w357_,
		_w377_,
		_w400_,
		_w1921_
	);
	LUT3 #(
		.INIT('hc8)
	) name1617 (
		_w412_,
		_w415_,
		_w425_,
		_w1922_
	);
	LUT3 #(
		.INIT('hc8)
	) name1618 (
		_w367_,
		_w333_,
		_w392_,
		_w1923_
	);
	LUT4 #(
		.INIT('h0001)
	) name1619 (
		_w1920_,
		_w1921_,
		_w1922_,
		_w1923_,
		_w1924_
	);
	LUT3 #(
		.INIT('hc8)
	) name1620 (
		_w374_,
		_w343_,
		_w396_,
		_w1925_
	);
	LUT3 #(
		.INIT('he0)
	) name1621 (
		_w337_,
		_w347_,
		_w388_,
		_w1926_
	);
	LUT3 #(
		.INIT('he0)
	) name1622 (
		_w375_,
		_w424_,
		_w406_,
		_w1927_
	);
	LUT3 #(
		.INIT('hc8)
	) name1623 (
		_w317_,
		_w411_,
		_w417_,
		_w1928_
	);
	LUT4 #(
		.INIT('h0001)
	) name1624 (
		_w1925_,
		_w1926_,
		_w1927_,
		_w1928_,
		_w1929_
	);
	LUT4 #(
		.INIT('h8000)
	) name1625 (
		_w1924_,
		_w1929_,
		_w1914_,
		_w1919_,
		_w1930_
	);
	LUT2 #(
		.INIT('h6)
	) name1626 (
		_w1745_,
		_w1930_,
		_w1931_
	);
	LUT3 #(
		.INIT('ha8)
	) name1627 (
		_w323_,
		_w420_,
		_w449_,
		_w1932_
	);
	LUT3 #(
		.INIT('ha8)
	) name1628 (
		_w377_,
		_w412_,
		_w561_,
		_w1933_
	);
	LUT3 #(
		.INIT('ha8)
	) name1629 (
		_w343_,
		_w483_,
		_w478_,
		_w1934_
	);
	LUT3 #(
		.INIT('ha8)
	) name1630 (
		_w423_,
		_w457_,
		_w460_,
		_w1935_
	);
	LUT4 #(
		.INIT('h0001)
	) name1631 (
		_w1932_,
		_w1933_,
		_w1934_,
		_w1935_,
		_w1936_
	);
	LUT3 #(
		.INIT('hc8)
	) name1632 (
		_w381_,
		_w411_,
		_w480_,
		_w1937_
	);
	LUT3 #(
		.INIT('ha8)
	) name1633 (
		_w305_,
		_w416_,
		_w548_,
		_w1938_
	);
	LUT3 #(
		.INIT('hc8)
	) name1634 (
		_w367_,
		_w402_,
		_w556_,
		_w1939_
	);
	LUT3 #(
		.INIT('ha8)
	) name1635 (
		_w363_,
		_w403_,
		_w471_,
		_w1940_
	);
	LUT4 #(
		.INIT('h0001)
	) name1636 (
		_w1937_,
		_w1938_,
		_w1939_,
		_w1940_,
		_w1941_
	);
	LUT3 #(
		.INIT('ha8)
	) name1637 (
		_w333_,
		_w455_,
		_w440_,
		_w1942_
	);
	LUT3 #(
		.INIT('hc8)
	) name1638 (
		_w327_,
		_w419_,
		_w553_,
		_w1943_
	);
	LUT3 #(
		.INIT('ha8)
	) name1639 (
		_w388_,
		_w459_,
		_w490_,
		_w1944_
	);
	LUT3 #(
		.INIT('hc8)
	) name1640 (
		_w317_,
		_w398_,
		_w435_,
		_w1945_
	);
	LUT4 #(
		.INIT('h0001)
	) name1641 (
		_w1942_,
		_w1943_,
		_w1944_,
		_w1945_,
		_w1946_
	);
	LUT3 #(
		.INIT('ha8)
	) name1642 (
		_w373_,
		_w465_,
		_w492_,
		_w1947_
	);
	LUT3 #(
		.INIT('ha8)
	) name1643 (
		_w312_,
		_w399_,
		_w433_,
		_w1948_
	);
	LUT3 #(
		.INIT('ha8)
	) name1644 (
		_w406_,
		_w444_,
		_w488_,
		_w1949_
	);
	LUT3 #(
		.INIT('hc8)
	) name1645 (
		_w357_,
		_w415_,
		_w473_,
		_w1950_
	);
	LUT4 #(
		.INIT('h0001)
	) name1646 (
		_w1947_,
		_w1948_,
		_w1949_,
		_w1950_,
		_w1951_
	);
	LUT4 #(
		.INIT('h8000)
	) name1647 (
		_w1946_,
		_w1951_,
		_w1936_,
		_w1941_,
		_w1952_
	);
	LUT4 #(
		.INIT('h0200)
	) name1648 (
		\desIn[41]_pad ,
		\roundSel[4]_pad ,
		\roundSel[5]_pad ,
		_w305_,
		_w1953_
	);
	LUT4 #(
		.INIT('h4155)
	) name1649 (
		\FP_R_reg[30]/P0001 ,
		\roundSel[4]_pad ,
		\roundSel[5]_pad ,
		_w305_,
		_w1954_
	);
	LUT4 #(
		.INIT('he8ff)
	) name1650 (
		\FP_R_reg[62]/NET0131 ,
		\roundSel[4]_pad ,
		\roundSel[5]_pad ,
		_w305_,
		_w1955_
	);
	LUT3 #(
		.INIT('h45)
	) name1651 (
		_w1953_,
		_w1954_,
		_w1955_,
		_w1956_
	);
	LUT3 #(
		.INIT('hba)
	) name1652 (
		_w1953_,
		_w1954_,
		_w1955_,
		_w1957_
	);
	LUT2 #(
		.INIT('h9)
	) name1653 (
		_w1952_,
		_w1956_,
		_w1958_
	);
	LUT3 #(
		.INIT('ha8)
	) name1654 (
		_w333_,
		_w421_,
		_w433_,
		_w1959_
	);
	LUT3 #(
		.INIT('hc8)
	) name1655 (
		_w341_,
		_w419_,
		_w490_,
		_w1960_
	);
	LUT3 #(
		.INIT('ha8)
	) name1656 (
		_w373_,
		_w559_,
		_w548_,
		_w1961_
	);
	LUT3 #(
		.INIT('hc8)
	) name1657 (
		_w417_,
		_w398_,
		_w457_,
		_w1962_
	);
	LUT4 #(
		.INIT('h0001)
	) name1658 (
		_w1959_,
		_w1960_,
		_w1961_,
		_w1962_,
		_w1963_
	);
	LUT3 #(
		.INIT('hc8)
	) name1659 (
		_w371_,
		_w312_,
		_w455_,
		_w1964_
	);
	LUT3 #(
		.INIT('ha8)
	) name1660 (
		_w305_,
		_w408_,
		_w492_,
		_w1965_
	);
	LUT3 #(
		.INIT('ha8)
	) name1661 (
		_w363_,
		_w321_,
		_w480_,
		_w1966_
	);
	LUT3 #(
		.INIT('hc8)
	) name1662 (
		_w361_,
		_w406_,
		_w561_,
		_w1967_
	);
	LUT4 #(
		.INIT('h0001)
	) name1663 (
		_w1964_,
		_w1965_,
		_w1966_,
		_w1967_,
		_w1968_
	);
	LUT3 #(
		.INIT('ha8)
	) name1664 (
		_w415_,
		_w400_,
		_w449_,
		_w1969_
	);
	LUT3 #(
		.INIT('hc8)
	) name1665 (
		_w392_,
		_w402_,
		_w478_,
		_w1970_
	);
	LUT3 #(
		.INIT('hc8)
	) name1666 (
		_w385_,
		_w423_,
		_w435_,
		_w1971_
	);
	LUT3 #(
		.INIT('ha8)
	) name1667 (
		_w323_,
		_w413_,
		_w473_,
		_w1972_
	);
	LUT4 #(
		.INIT('h0001)
	) name1668 (
		_w1969_,
		_w1970_,
		_w1971_,
		_w1972_,
		_w1973_
	);
	LUT3 #(
		.INIT('hc8)
	) name1669 (
		_w331_,
		_w411_,
		_w471_,
		_w1974_
	);
	LUT3 #(
		.INIT('ha8)
	) name1670 (
		_w377_,
		_w425_,
		_w488_,
		_w1975_
	);
	LUT3 #(
		.INIT('ha8)
	) name1671 (
		_w343_,
		_w539_,
		_w556_,
		_w1976_
	);
	LUT3 #(
		.INIT('ha8)
	) name1672 (
		_w388_,
		_w404_,
		_w553_,
		_w1977_
	);
	LUT4 #(
		.INIT('h0001)
	) name1673 (
		_w1974_,
		_w1975_,
		_w1976_,
		_w1977_,
		_w1978_
	);
	LUT4 #(
		.INIT('h8000)
	) name1674 (
		_w1973_,
		_w1978_,
		_w1963_,
		_w1968_,
		_w1979_
	);
	LUT2 #(
		.INIT('h9)
	) name1675 (
		_w1599_,
		_w1979_,
		_w1980_
	);
	LUT4 #(
		.INIT('h1428)
	) name1676 (
		_w1599_,
		_w1952_,
		_w1956_,
		_w1979_,
		_w1981_
	);
	LUT3 #(
		.INIT('ha8)
	) name1677 (
		_w373_,
		_w471_,
		_w480_,
		_w1982_
	);
	LUT3 #(
		.INIT('hc8)
	) name1678 (
		_w385_,
		_w419_,
		_w460_,
		_w1983_
	);
	LUT3 #(
		.INIT('ha8)
	) name1679 (
		_w398_,
		_w404_,
		_w459_,
		_w1984_
	);
	LUT3 #(
		.INIT('hc8)
	) name1680 (
		_w361_,
		_w312_,
		_w444_,
		_w1985_
	);
	LUT4 #(
		.INIT('h0001)
	) name1681 (
		_w1982_,
		_w1983_,
		_w1984_,
		_w1985_,
		_w1986_
	);
	LUT3 #(
		.INIT('ha8)
	) name1682 (
		_w343_,
		_w449_,
		_w473_,
		_w1987_
	);
	LUT3 #(
		.INIT('he0)
	) name1683 (
		_w357_,
		_w400_,
		_w402_,
		_w1988_
	);
	LUT3 #(
		.INIT('ha8)
	) name1684 (
		_w406_,
		_w455_,
		_w433_,
		_w1989_
	);
	LUT3 #(
		.INIT('ha8)
	) name1685 (
		_w333_,
		_w488_,
		_w561_,
		_w1990_
	);
	LUT4 #(
		.INIT('h0001)
	) name1686 (
		_w1987_,
		_w1988_,
		_w1989_,
		_w1990_,
		_w1991_
	);
	LUT3 #(
		.INIT('ha8)
	) name1687 (
		_w363_,
		_w492_,
		_w548_,
		_w1992_
	);
	LUT3 #(
		.INIT('ha8)
	) name1688 (
		_w377_,
		_w421_,
		_w440_,
		_w1993_
	);
	LUT3 #(
		.INIT('ha8)
	) name1689 (
		_w411_,
		_w465_,
		_w559_,
		_w1994_
	);
	LUT3 #(
		.INIT('ha8)
	) name1690 (
		_w423_,
		_w490_,
		_w553_,
		_w1995_
	);
	LUT4 #(
		.INIT('h0001)
	) name1691 (
		_w1992_,
		_w1993_,
		_w1994_,
		_w1995_,
		_w1996_
	);
	LUT3 #(
		.INIT('ha8)
	) name1692 (
		_w323_,
		_w483_,
		_w539_,
		_w1997_
	);
	LUT3 #(
		.INIT('ha8)
	) name1693 (
		_w305_,
		_w321_,
		_w403_,
		_w1998_
	);
	LUT3 #(
		.INIT('ha8)
	) name1694 (
		_w388_,
		_w457_,
		_w435_,
		_w1999_
	);
	LUT3 #(
		.INIT('ha8)
	) name1695 (
		_w415_,
		_w478_,
		_w556_,
		_w2000_
	);
	LUT4 #(
		.INIT('h0001)
	) name1696 (
		_w1997_,
		_w1998_,
		_w1999_,
		_w2000_,
		_w2001_
	);
	LUT4 #(
		.INIT('h8000)
	) name1697 (
		_w1996_,
		_w2001_,
		_w1986_,
		_w1991_,
		_w2002_
	);
	LUT2 #(
		.INIT('h9)
	) name1698 (
		_w1444_,
		_w2002_,
		_w2003_
	);
	LUT4 #(
		.INIT('h1428)
	) name1699 (
		_w1444_,
		_w1745_,
		_w1930_,
		_w2002_,
		_w2004_
	);
	LUT4 #(
		.INIT('h2814)
	) name1700 (
		_w1444_,
		_w1952_,
		_w1956_,
		_w2002_,
		_w2005_
	);
	LUT4 #(
		.INIT('h76f2)
	) name1701 (
		_w1958_,
		_w1980_,
		_w1931_,
		_w2003_,
		_w2006_
	);
	LUT2 #(
		.INIT('h2)
	) name1702 (
		_w1909_,
		_w2006_,
		_w2007_
	);
	LUT4 #(
		.INIT('h2814)
	) name1703 (
		_w1444_,
		_w1745_,
		_w1930_,
		_w2002_,
		_w2008_
	);
	LUT4 #(
		.INIT('ha820)
	) name1704 (
		_w1958_,
		_w1980_,
		_w2004_,
		_w2008_,
		_w2009_
	);
	LUT4 #(
		.INIT('h4182)
	) name1705 (
		_w1599_,
		_w1952_,
		_w1956_,
		_w1979_,
		_w2010_
	);
	LUT4 #(
		.INIT('h8241)
	) name1706 (
		_w1444_,
		_w1745_,
		_w1930_,
		_w2002_,
		_w2011_
	);
	LUT4 #(
		.INIT('ha3ff)
	) name1707 (
		_w1958_,
		_w2010_,
		_w1931_,
		_w2003_,
		_w2012_
	);
	LUT3 #(
		.INIT('h10)
	) name1708 (
		_w1931_,
		_w2003_,
		_w1981_,
		_w2013_
	);
	LUT4 #(
		.INIT('h000e)
	) name1709 (
		_w1909_,
		_w2012_,
		_w2009_,
		_w2013_,
		_w2014_
	);
	LUT3 #(
		.INIT('h8a)
	) name1710 (
		_w1882_,
		_w2007_,
		_w2014_,
		_w2015_
	);
	LUT4 #(
		.INIT('h1dff)
	) name1711 (
		_w1958_,
		_w1980_,
		_w1931_,
		_w2003_,
		_w2016_
	);
	LUT2 #(
		.INIT('h2)
	) name1712 (
		_w1909_,
		_w2016_,
		_w2017_
	);
	LUT4 #(
		.INIT('h4182)
	) name1713 (
		_w1444_,
		_w1952_,
		_w1956_,
		_w2002_,
		_w2018_
	);
	LUT4 #(
		.INIT('h2184)
	) name1714 (
		_w1599_,
		_w1745_,
		_w1979_,
		_w1930_,
		_w2019_
	);
	LUT4 #(
		.INIT('h1428)
	) name1715 (
		_w1444_,
		_w1903_,
		_w1907_,
		_w2002_,
		_w2020_
	);
	LUT4 #(
		.INIT('h575f)
	) name1716 (
		_w1980_,
		_w1931_,
		_w2018_,
		_w2020_,
		_w2021_
	);
	LUT4 #(
		.INIT('h4182)
	) name1717 (
		_w1444_,
		_w1745_,
		_w1930_,
		_w2002_,
		_w2022_
	);
	LUT4 #(
		.INIT('h6006)
	) name1718 (
		_w1903_,
		_w1907_,
		_w1952_,
		_w1956_,
		_w2023_
	);
	LUT4 #(
		.INIT('hcedf)
	) name1719 (
		_w1931_,
		_w2003_,
		_w1981_,
		_w2023_,
		_w2024_
	);
	LUT3 #(
		.INIT('h80)
	) name1720 (
		_w2010_,
		_w1931_,
		_w2003_,
		_w2025_
	);
	LUT4 #(
		.INIT('h0660)
	) name1721 (
		_w1903_,
		_w1907_,
		_w1952_,
		_w1956_,
		_w2026_
	);
	LUT4 #(
		.INIT('h2814)
	) name1722 (
		_w1599_,
		_w1952_,
		_w1956_,
		_w1979_,
		_w2027_
	);
	LUT3 #(
		.INIT('ha8)
	) name1723 (
		_w2011_,
		_w2026_,
		_w2027_,
		_w2028_
	);
	LUT4 #(
		.INIT('h1000)
	) name1724 (
		_w2025_,
		_w2028_,
		_w2021_,
		_w2024_,
		_w2029_
	);
	LUT3 #(
		.INIT('h20)
	) name1725 (
		_w1909_,
		_w2003_,
		_w1981_,
		_w2030_
	);
	LUT3 #(
		.INIT('h80)
	) name1726 (
		_w1980_,
		_w2011_,
		_w2026_,
		_w2031_
	);
	LUT2 #(
		.INIT('h1)
	) name1727 (
		_w2030_,
		_w2031_,
		_w2032_
	);
	LUT4 #(
		.INIT('hba00)
	) name1728 (
		_w1882_,
		_w2017_,
		_w2029_,
		_w2032_,
		_w2033_
	);
	LUT4 #(
		.INIT('h0100)
	) name1729 (
		\desIn[34]_pad ,
		\roundSel[4]_pad ,
		\roundSel[5]_pad ,
		_w305_,
		_w2034_
	);
	LUT4 #(
		.INIT('h2800)
	) name1730 (
		\FP_R_reg[21]/P0001 ,
		\roundSel[4]_pad ,
		\roundSel[5]_pad ,
		_w305_,
		_w2035_
	);
	LUT4 #(
		.INIT('h7c55)
	) name1731 (
		\FP_R_reg[53]/NET0131 ,
		\roundSel[4]_pad ,
		\roundSel[5]_pad ,
		_w305_,
		_w2036_
	);
	LUT3 #(
		.INIT('h45)
	) name1732 (
		_w2034_,
		_w2035_,
		_w2036_,
		_w2037_
	);
	LUT3 #(
		.INIT('h4b)
	) name1733 (
		_w2015_,
		_w2033_,
		_w2037_,
		_w2038_
	);
	LUT4 #(
		.INIT('h802a)
	) name1734 (
		_w1909_,
		_w1980_,
		_w1931_,
		_w2005_,
		_w2039_
	);
	LUT3 #(
		.INIT('h15)
	) name1735 (
		_w1909_,
		_w2010_,
		_w2003_,
		_w2040_
	);
	LUT4 #(
		.INIT('h5154)
	) name1736 (
		_w1909_,
		_w1958_,
		_w1980_,
		_w2003_,
		_w2041_
	);
	LUT3 #(
		.INIT('h80)
	) name1737 (
		_w1958_,
		_w1980_,
		_w2022_,
		_w2042_
	);
	LUT4 #(
		.INIT('haa02)
	) name1738 (
		_w1882_,
		_w2039_,
		_w2041_,
		_w2042_,
		_w2043_
	);
	LUT4 #(
		.INIT('h4812)
	) name1739 (
		_w1599_,
		_w1745_,
		_w1979_,
		_w1930_,
		_w2044_
	);
	LUT4 #(
		.INIT('hdffc)
	) name1740 (
		_w1958_,
		_w1980_,
		_w1931_,
		_w2003_,
		_w2045_
	);
	LUT4 #(
		.INIT('h0032)
	) name1741 (
		_w2005_,
		_w2008_,
		_w2019_,
		_w2027_,
		_w2046_
	);
	LUT4 #(
		.INIT('h0777)
	) name1742 (
		_w1981_,
		_w2004_,
		_w2018_,
		_w2044_,
		_w2047_
	);
	LUT4 #(
		.INIT('h0e00)
	) name1743 (
		_w1882_,
		_w2045_,
		_w2046_,
		_w2047_,
		_w2048_
	);
	LUT4 #(
		.INIT('h5404)
	) name1744 (
		_w1909_,
		_w1980_,
		_w1931_,
		_w2018_,
		_w2049_
	);
	LUT3 #(
		.INIT('hc4)
	) name1745 (
		_w1909_,
		_w2005_,
		_w2019_,
		_w2050_
	);
	LUT3 #(
		.INIT('h80)
	) name1746 (
		_w1958_,
		_w1980_,
		_w2011_,
		_w2051_
	);
	LUT4 #(
		.INIT('h5554)
	) name1747 (
		_w1882_,
		_w2050_,
		_w2051_,
		_w2049_,
		_w2052_
	);
	LUT3 #(
		.INIT('h80)
	) name1748 (
		_w1980_,
		_w2008_,
		_w2026_,
		_w2053_
	);
	LUT4 #(
		.INIT('h000d)
	) name1749 (
		_w1909_,
		_w2048_,
		_w2052_,
		_w2053_,
		_w2054_
	);
	LUT4 #(
		.INIT('h0100)
	) name1750 (
		\desIn[38]_pad ,
		\roundSel[4]_pad ,
		\roundSel[5]_pad ,
		_w305_,
		_w2055_
	);
	LUT4 #(
		.INIT('h2800)
	) name1751 (
		\FP_R_reg[5]/P0001 ,
		\roundSel[4]_pad ,
		\roundSel[5]_pad ,
		_w305_,
		_w2056_
	);
	LUT4 #(
		.INIT('h7c55)
	) name1752 (
		\FP_R_reg[37]/NET0131 ,
		\roundSel[4]_pad ,
		\roundSel[5]_pad ,
		_w305_,
		_w2057_
	);
	LUT3 #(
		.INIT('h45)
	) name1753 (
		_w2055_,
		_w2056_,
		_w2057_,
		_w2058_
	);
	LUT3 #(
		.INIT('hb4)
	) name1754 (
		_w2043_,
		_w2054_,
		_w2058_,
		_w2059_
	);
	LUT3 #(
		.INIT('ha8)
	) name1755 (
		_w363_,
		_w703_,
		_w865_,
		_w2060_
	);
	LUT3 #(
		.INIT('ha8)
	) name1756 (
		_w419_,
		_w721_,
		_w863_,
		_w2061_
	);
	LUT3 #(
		.INIT('ha8)
	) name1757 (
		_w402_,
		_w755_,
		_w868_,
		_w2062_
	);
	LUT3 #(
		.INIT('ha8)
	) name1758 (
		_w343_,
		_w725_,
		_w740_,
		_w2063_
	);
	LUT4 #(
		.INIT('h0001)
	) name1759 (
		_w2060_,
		_w2061_,
		_w2062_,
		_w2063_,
		_w2064_
	);
	LUT3 #(
		.INIT('ha8)
	) name1760 (
		_w323_,
		_w756_,
		_w860_,
		_w2065_
	);
	LUT3 #(
		.INIT('ha8)
	) name1761 (
		_w305_,
		_w746_,
		_w847_,
		_w2066_
	);
	LUT3 #(
		.INIT('ha8)
	) name1762 (
		_w398_,
		_w717_,
		_w858_,
		_w2067_
	);
	LUT3 #(
		.INIT('ha8)
	) name1763 (
		_w411_,
		_w750_,
		_w824_,
		_w2068_
	);
	LUT4 #(
		.INIT('h0001)
	) name1764 (
		_w2065_,
		_w2066_,
		_w2067_,
		_w2068_,
		_w2069_
	);
	LUT3 #(
		.INIT('ha8)
	) name1765 (
		_w406_,
		_w690_,
		_w753_,
		_w2070_
	);
	LUT3 #(
		.INIT('ha8)
	) name1766 (
		_w377_,
		_w759_,
		_w842_,
		_w2071_
	);
	LUT3 #(
		.INIT('ha8)
	) name1767 (
		_w312_,
		_w758_,
		_w837_,
		_w2072_
	);
	LUT3 #(
		.INIT('ha8)
	) name1768 (
		_w415_,
		_w681_,
		_w856_,
		_w2073_
	);
	LUT4 #(
		.INIT('h0001)
	) name1769 (
		_w2070_,
		_w2071_,
		_w2072_,
		_w2073_,
		_w2074_
	);
	LUT3 #(
		.INIT('ha8)
	) name1770 (
		_w423_,
		_w672_,
		_w831_,
		_w2075_
	);
	LUT3 #(
		.INIT('ha8)
	) name1771 (
		_w373_,
		_w700_,
		_w712_,
		_w2076_
	);
	LUT3 #(
		.INIT('ha8)
	) name1772 (
		_w388_,
		_w734_,
		_w737_,
		_w2077_
	);
	LUT3 #(
		.INIT('ha8)
	) name1773 (
		_w333_,
		_w669_,
		_w849_,
		_w2078_
	);
	LUT4 #(
		.INIT('h0001)
	) name1774 (
		_w2075_,
		_w2076_,
		_w2077_,
		_w2078_,
		_w2079_
	);
	LUT4 #(
		.INIT('h8000)
	) name1775 (
		_w2074_,
		_w2079_,
		_w2064_,
		_w2069_,
		_w2080_
	);
	LUT2 #(
		.INIT('h6)
	) name1776 (
		_w1084_,
		_w2080_,
		_w2081_
	);
	LUT3 #(
		.INIT('ha8)
	) name1777 (
		_w305_,
		_w756_,
		_w806_,
		_w2082_
	);
	LUT3 #(
		.INIT('ha8)
	) name1778 (
		_w343_,
		_w865_,
		_w831_,
		_w2083_
	);
	LUT3 #(
		.INIT('ha8)
	) name1779 (
		_w402_,
		_w750_,
		_w802_,
		_w2084_
	);
	LUT3 #(
		.INIT('ha8)
	) name1780 (
		_w411_,
		_w753_,
		_w868_,
		_w2085_
	);
	LUT4 #(
		.INIT('h0001)
	) name1781 (
		_w2082_,
		_w2083_,
		_w2084_,
		_w2085_,
		_w2086_
	);
	LUT3 #(
		.INIT('ha8)
	) name1782 (
		_w377_,
		_w703_,
		_w797_,
		_w2087_
	);
	LUT3 #(
		.INIT('ha8)
	) name1783 (
		_w323_,
		_w734_,
		_w847_,
		_w2088_
	);
	LUT3 #(
		.INIT('ha8)
	) name1784 (
		_w363_,
		_w740_,
		_w842_,
		_w2089_
	);
	LUT3 #(
		.INIT('ha8)
	) name1785 (
		_w423_,
		_w725_,
		_w837_,
		_w2090_
	);
	LUT4 #(
		.INIT('h0001)
	) name1786 (
		_w2087_,
		_w2088_,
		_w2089_,
		_w2090_,
		_w2091_
	);
	LUT3 #(
		.INIT('ha8)
	) name1787 (
		_w406_,
		_w737_,
		_w824_,
		_w2092_
	);
	LUT3 #(
		.INIT('ha8)
	) name1788 (
		_w419_,
		_w681_,
		_w772_,
		_w2093_
	);
	LUT3 #(
		.INIT('ha8)
	) name1789 (
		_w415_,
		_w712_,
		_w863_,
		_w2094_
	);
	LUT3 #(
		.INIT('ha8)
	) name1790 (
		_w333_,
		_w700_,
		_w858_,
		_w2095_
	);
	LUT4 #(
		.INIT('h0001)
	) name1791 (
		_w2092_,
		_w2093_,
		_w2094_,
		_w2095_,
		_w2096_
	);
	LUT3 #(
		.INIT('ha8)
	) name1792 (
		_w398_,
		_w669_,
		_w788_,
		_w2097_
	);
	LUT3 #(
		.INIT('ha8)
	) name1793 (
		_w388_,
		_w690_,
		_w860_,
		_w2098_
	);
	LUT3 #(
		.INIT('ha8)
	) name1794 (
		_w373_,
		_w856_,
		_w849_,
		_w2099_
	);
	LUT3 #(
		.INIT('ha8)
	) name1795 (
		_w312_,
		_w672_,
		_w786_,
		_w2100_
	);
	LUT4 #(
		.INIT('h0001)
	) name1796 (
		_w2097_,
		_w2098_,
		_w2099_,
		_w2100_,
		_w2101_
	);
	LUT4 #(
		.INIT('h8000)
	) name1797 (
		_w2096_,
		_w2101_,
		_w2086_,
		_w2091_,
		_w2102_
	);
	LUT2 #(
		.INIT('h6)
	) name1798 (
		_w818_,
		_w2102_,
		_w2103_
	);
	LUT4 #(
		.INIT('h4182)
	) name1799 (
		_w818_,
		_w1084_,
		_w2080_,
		_w2102_,
		_w2104_
	);
	LUT3 #(
		.INIT('ha8)
	) name1800 (
		_w363_,
		_w856_,
		_w806_,
		_w2105_
	);
	LUT3 #(
		.INIT('ha8)
	) name1801 (
		_w402_,
		_w712_,
		_w736_,
		_w2106_
	);
	LUT3 #(
		.INIT('ha8)
	) name1802 (
		_w323_,
		_w767_,
		_w831_,
		_w2107_
	);
	LUT3 #(
		.INIT('ha8)
	) name1803 (
		_w423_,
		_w860_,
		_w772_,
		_w2108_
	);
	LUT4 #(
		.INIT('h0001)
	) name1804 (
		_w2105_,
		_w2106_,
		_w2107_,
		_w2108_,
		_w2109_
	);
	LUT3 #(
		.INIT('ha8)
	) name1805 (
		_w415_,
		_w802_,
		_w865_,
		_w2110_
	);
	LUT3 #(
		.INIT('ha8)
	) name1806 (
		_w377_,
		_w700_,
		_w793_,
		_w2111_
	);
	LUT3 #(
		.INIT('ha8)
	) name1807 (
		_w305_,
		_w686_,
		_w740_,
		_w2112_
	);
	LUT3 #(
		.INIT('ha8)
	) name1808 (
		_w398_,
		_w690_,
		_w811_,
		_w2113_
	);
	LUT4 #(
		.INIT('h0001)
	) name1809 (
		_w2110_,
		_w2111_,
		_w2112_,
		_w2113_,
		_w2114_
	);
	LUT3 #(
		.INIT('ha8)
	) name1810 (
		_w411_,
		_w774_,
		_w849_,
		_w2115_
	);
	LUT3 #(
		.INIT('ha8)
	) name1811 (
		_w419_,
		_w725_,
		_w809_,
		_w2116_
	);
	LUT3 #(
		.INIT('ha8)
	) name1812 (
		_w373_,
		_w868_,
		_w842_,
		_w2117_
	);
	LUT3 #(
		.INIT('ha8)
	) name1813 (
		_w312_,
		_w737_,
		_w779_,
		_w2118_
	);
	LUT4 #(
		.INIT('h0001)
	) name1814 (
		_w2115_,
		_w2116_,
		_w2117_,
		_w2118_,
		_w2119_
	);
	LUT3 #(
		.INIT('ha8)
	) name1815 (
		_w406_,
		_w786_,
		_w858_,
		_w2120_
	);
	LUT3 #(
		.INIT('ha8)
	) name1816 (
		_w333_,
		_w824_,
		_w797_,
		_w2121_
	);
	LUT3 #(
		.INIT('ha8)
	) name1817 (
		_w388_,
		_w788_,
		_w837_,
		_w2122_
	);
	LUT3 #(
		.INIT('ha8)
	) name1818 (
		_w343_,
		_w863_,
		_w847_,
		_w2123_
	);
	LUT4 #(
		.INIT('h0001)
	) name1819 (
		_w2120_,
		_w2121_,
		_w2122_,
		_w2123_,
		_w2124_
	);
	LUT4 #(
		.INIT('h8000)
	) name1820 (
		_w2119_,
		_w2124_,
		_w2109_,
		_w2114_,
		_w2125_
	);
	LUT2 #(
		.INIT('h9)
	) name1821 (
		_w997_,
		_w2125_,
		_w2126_
	);
	LUT3 #(
		.INIT('ha8)
	) name1822 (
		_w343_,
		_w856_,
		_w860_,
		_w2127_
	);
	LUT3 #(
		.INIT('ha8)
	) name1823 (
		_w305_,
		_w703_,
		_w767_,
		_w2128_
	);
	LUT3 #(
		.INIT('ha8)
	) name1824 (
		_w402_,
		_w681_,
		_w774_,
		_w2129_
	);
	LUT3 #(
		.INIT('ha8)
	) name1825 (
		_w323_,
		_w740_,
		_w788_,
		_w2130_
	);
	LUT4 #(
		.INIT('h0001)
	) name1826 (
		_w2127_,
		_w2128_,
		_w2129_,
		_w2130_,
		_w2131_
	);
	LUT3 #(
		.INIT('ha8)
	) name1827 (
		_w406_,
		_w837_,
		_w849_,
		_w2132_
	);
	LUT3 #(
		.INIT('ha8)
	) name1828 (
		_w419_,
		_w672_,
		_w802_,
		_w2133_
	);
	LUT3 #(
		.INIT('ha8)
	) name1829 (
		_w388_,
		_w858_,
		_w831_,
		_w2134_
	);
	LUT3 #(
		.INIT('ha8)
	) name1830 (
		_w415_,
		_w725_,
		_w868_,
		_w2135_
	);
	LUT4 #(
		.INIT('h0001)
	) name1831 (
		_w2132_,
		_w2133_,
		_w2134_,
		_w2135_,
		_w2136_
	);
	LUT3 #(
		.INIT('ha8)
	) name1832 (
		_w373_,
		_w824_,
		_w865_,
		_w2137_
	);
	LUT3 #(
		.INIT('ha8)
	) name1833 (
		_w312_,
		_w753_,
		_w772_,
		_w2138_
	);
	LUT3 #(
		.INIT('ha8)
	) name1834 (
		_w333_,
		_w690_,
		_w842_,
		_w2139_
	);
	LUT3 #(
		.INIT('ha8)
	) name1835 (
		_w398_,
		_w734_,
		_w797_,
		_w2140_
	);
	LUT4 #(
		.INIT('h0001)
	) name1836 (
		_w2137_,
		_w2138_,
		_w2139_,
		_w2140_,
		_w2141_
	);
	LUT3 #(
		.INIT('ha8)
	) name1837 (
		_w363_,
		_w700_,
		_w847_,
		_w2142_
	);
	LUT3 #(
		.INIT('ha8)
	) name1838 (
		_w411_,
		_w712_,
		_w786_,
		_w2143_
	);
	LUT3 #(
		.INIT('ha8)
	) name1839 (
		_w423_,
		_w737_,
		_w863_,
		_w2144_
	);
	LUT3 #(
		.INIT('ha8)
	) name1840 (
		_w377_,
		_w669_,
		_w806_,
		_w2145_
	);
	LUT4 #(
		.INIT('h0001)
	) name1841 (
		_w2142_,
		_w2143_,
		_w2144_,
		_w2145_,
		_w2146_
	);
	LUT4 #(
		.INIT('h8000)
	) name1842 (
		_w2141_,
		_w2146_,
		_w2131_,
		_w2136_,
		_w2147_
	);
	LUT2 #(
		.INIT('h6)
	) name1843 (
		_w1002_,
		_w2147_,
		_w2148_
	);
	LUT4 #(
		.INIT('h8421)
	) name1844 (
		_w997_,
		_w1002_,
		_w2125_,
		_w2147_,
		_w2149_
	);
	LUT3 #(
		.INIT('ha8)
	) name1845 (
		_w406_,
		_w700_,
		_w672_,
		_w2150_
	);
	LUT3 #(
		.INIT('ha8)
	) name1846 (
		_w388_,
		_w669_,
		_w725_,
		_w2151_
	);
	LUT3 #(
		.INIT('ha8)
	) name1847 (
		_w343_,
		_w712_,
		_w734_,
		_w2152_
	);
	LUT3 #(
		.INIT('ha8)
	) name1848 (
		_w415_,
		_w750_,
		_w831_,
		_w2153_
	);
	LUT4 #(
		.INIT('h0001)
	) name1849 (
		_w2150_,
		_w2151_,
		_w2152_,
		_w2153_,
		_w2154_
	);
	LUT3 #(
		.INIT('ha8)
	) name1850 (
		_w402_,
		_w702_,
		_w863_,
		_w2155_
	);
	LUT3 #(
		.INIT('ha8)
	) name1851 (
		_w398_,
		_w759_,
		_w860_,
		_w2156_
	);
	LUT3 #(
		.INIT('ha8)
	) name1852 (
		_w333_,
		_w703_,
		_w737_,
		_w2157_
	);
	LUT3 #(
		.INIT('ha8)
	) name1853 (
		_w411_,
		_w758_,
		_w856_,
		_w2158_
	);
	LUT4 #(
		.INIT('h0001)
	) name1854 (
		_w2155_,
		_w2156_,
		_w2157_,
		_w2158_,
		_w2159_
	);
	LUT3 #(
		.INIT('ha8)
	) name1855 (
		_w377_,
		_w746_,
		_w858_,
		_w2160_
	);
	LUT3 #(
		.INIT('ha8)
	) name1856 (
		_w373_,
		_w753_,
		_w740_,
		_w2161_
	);
	LUT3 #(
		.INIT('ha8)
	) name1857 (
		_w363_,
		_w756_,
		_w849_,
		_w2162_
	);
	LUT3 #(
		.INIT('ha8)
	) name1858 (
		_w323_,
		_w717_,
		_w865_,
		_w2163_
	);
	LUT4 #(
		.INIT('h0001)
	) name1859 (
		_w2160_,
		_w2161_,
		_w2162_,
		_w2163_,
		_w2164_
	);
	LUT3 #(
		.INIT('ha8)
	) name1860 (
		_w419_,
		_w755_,
		_w837_,
		_w2165_
	);
	LUT3 #(
		.INIT('ha8)
	) name1861 (
		_w423_,
		_w681_,
		_w690_,
		_w2166_
	);
	LUT3 #(
		.INIT('ha8)
	) name1862 (
		_w312_,
		_w721_,
		_w824_,
		_w2167_
	);
	LUT3 #(
		.INIT('ha8)
	) name1863 (
		_w305_,
		_w677_,
		_w842_,
		_w2168_
	);
	LUT4 #(
		.INIT('h0001)
	) name1864 (
		_w2165_,
		_w2166_,
		_w2167_,
		_w2168_,
		_w2169_
	);
	LUT4 #(
		.INIT('h8000)
	) name1865 (
		_w2164_,
		_w2169_,
		_w2154_,
		_w2159_,
		_w2170_
	);
	LUT4 #(
		.INIT('h0200)
	) name1866 (
		\desIn[21]_pad ,
		\roundSel[4]_pad ,
		\roundSel[5]_pad ,
		_w305_,
		_w2171_
	);
	LUT4 #(
		.INIT('h4155)
	) name1867 (
		\FP_R_reg[11]/P0001 ,
		\roundSel[4]_pad ,
		\roundSel[5]_pad ,
		_w305_,
		_w2172_
	);
	LUT4 #(
		.INIT('he8ff)
	) name1868 (
		\FP_R_reg[43]/NET0131 ,
		\roundSel[4]_pad ,
		\roundSel[5]_pad ,
		_w305_,
		_w2173_
	);
	LUT3 #(
		.INIT('h45)
	) name1869 (
		_w2171_,
		_w2172_,
		_w2173_,
		_w2174_
	);
	LUT3 #(
		.INIT('hba)
	) name1870 (
		_w2171_,
		_w2172_,
		_w2173_,
		_w2175_
	);
	LUT2 #(
		.INIT('h9)
	) name1871 (
		_w2170_,
		_w2174_,
		_w2176_
	);
	LUT4 #(
		.INIT('h2600)
	) name1872 (
		_w2104_,
		_w2126_,
		_w2148_,
		_w2176_,
		_w2177_
	);
	LUT4 #(
		.INIT('h1428)
	) name1873 (
		_w1002_,
		_w1084_,
		_w2080_,
		_w2147_,
		_w2178_
	);
	LUT4 #(
		.INIT('h0001)
	) name1874 (
		_w2104_,
		_w2149_,
		_w2176_,
		_w2178_,
		_w2179_
	);
	LUT3 #(
		.INIT('ha8)
	) name1875 (
		_w406_,
		_w702_,
		_w717_,
		_w2180_
	);
	LUT3 #(
		.INIT('ha8)
	) name1876 (
		_w363_,
		_w681_,
		_w752_,
		_w2181_
	);
	LUT3 #(
		.INIT('ha8)
	) name1877 (
		_w323_,
		_w708_,
		_w672_,
		_w2182_
	);
	LUT3 #(
		.INIT('ha8)
	) name1878 (
		_w415_,
		_w703_,
		_w730_,
		_w2183_
	);
	LUT4 #(
		.INIT('h0001)
	) name1879 (
		_w2180_,
		_w2181_,
		_w2182_,
		_w2183_,
		_w2184_
	);
	LUT3 #(
		.INIT('ha8)
	) name1880 (
		_w419_,
		_w686_,
		_w740_,
		_w2185_
	);
	LUT3 #(
		.INIT('ha8)
	) name1881 (
		_w388_,
		_w677_,
		_w758_,
		_w2186_
	);
	LUT3 #(
		.INIT('ha8)
	) name1882 (
		_w411_,
		_w669_,
		_w739_,
		_w2187_
	);
	LUT3 #(
		.INIT('ha8)
	) name1883 (
		_w402_,
		_w700_,
		_w793_,
		_w2188_
	);
	LUT4 #(
		.INIT('h0001)
	) name1884 (
		_w2185_,
		_w2186_,
		_w2187_,
		_w2188_,
		_w2189_
	);
	LUT3 #(
		.INIT('ha8)
	) name1885 (
		_w343_,
		_w721_,
		_w746_,
		_w2190_
	);
	LUT3 #(
		.INIT('ha8)
	) name1886 (
		_w373_,
		_w755_,
		_w759_,
		_w2191_
	);
	LUT3 #(
		.INIT('ha8)
	) name1887 (
		_w377_,
		_w712_,
		_w736_,
		_w2192_
	);
	LUT3 #(
		.INIT('ha8)
	) name1888 (
		_w423_,
		_w665_,
		_w756_,
		_w2193_
	);
	LUT4 #(
		.INIT('h0001)
	) name1889 (
		_w2190_,
		_w2191_,
		_w2192_,
		_w2193_,
		_w2194_
	);
	LUT3 #(
		.INIT('ha8)
	) name1890 (
		_w312_,
		_w696_,
		_w734_,
		_w2195_
	);
	LUT3 #(
		.INIT('ha8)
	) name1891 (
		_w398_,
		_w753_,
		_w724_,
		_w2196_
	);
	LUT3 #(
		.INIT('ha8)
	) name1892 (
		_w305_,
		_w725_,
		_w809_,
		_w2197_
	);
	LUT3 #(
		.INIT('ha8)
	) name1893 (
		_w333_,
		_w671_,
		_w750_,
		_w2198_
	);
	LUT4 #(
		.INIT('h0001)
	) name1894 (
		_w2195_,
		_w2196_,
		_w2197_,
		_w2198_,
		_w2199_
	);
	LUT4 #(
		.INIT('h8000)
	) name1895 (
		_w2194_,
		_w2199_,
		_w2184_,
		_w2189_,
		_w2200_
	);
	LUT2 #(
		.INIT('h9)
	) name1896 (
		_w904_,
		_w2200_,
		_w2201_
	);
	LUT4 #(
		.INIT('h1428)
	) name1897 (
		_w997_,
		_w1084_,
		_w2080_,
		_w2125_,
		_w2202_
	);
	LUT4 #(
		.INIT('h1248)
	) name1898 (
		_w818_,
		_w1002_,
		_w2102_,
		_w2147_,
		_w2203_
	);
	LUT4 #(
		.INIT('h8421)
	) name1899 (
		_w818_,
		_w1002_,
		_w2102_,
		_w2147_,
		_w2204_
	);
	LUT4 #(
		.INIT('h6996)
	) name1900 (
		_w818_,
		_w1002_,
		_w2102_,
		_w2147_,
		_w2205_
	);
	LUT2 #(
		.INIT('h2)
	) name1901 (
		_w2202_,
		_w2205_,
		_w2206_
	);
	LUT4 #(
		.INIT('h2814)
	) name1902 (
		_w818_,
		_w1084_,
		_w2080_,
		_w2102_,
		_w2207_
	);
	LUT3 #(
		.INIT('h80)
	) name1903 (
		_w2126_,
		_w2148_,
		_w2207_,
		_w2208_
	);
	LUT4 #(
		.INIT('h0001)
	) name1904 (
		_w2179_,
		_w2206_,
		_w2201_,
		_w2208_,
		_w2209_
	);
	LUT4 #(
		.INIT('h2184)
	) name1905 (
		_w818_,
		_w1002_,
		_w2102_,
		_w2147_,
		_w2210_
	);
	LUT4 #(
		.INIT('h084c)
	) name1906 (
		_w2126_,
		_w2176_,
		_w2203_,
		_w2210_,
		_w2211_
	);
	LUT4 #(
		.INIT('h0203)
	) name1907 (
		_w2081_,
		_w2149_,
		_w2176_,
		_w2203_,
		_w2212_
	);
	LUT4 #(
		.INIT('h6006)
	) name1908 (
		_w997_,
		_w2125_,
		_w2170_,
		_w2174_,
		_w2213_
	);
	LUT4 #(
		.INIT('h4812)
	) name1909 (
		_w818_,
		_w1002_,
		_w2102_,
		_w2147_,
		_w2214_
	);
	LUT3 #(
		.INIT('h80)
	) name1910 (
		_w2081_,
		_w2213_,
		_w2214_,
		_w2215_
	);
	LUT4 #(
		.INIT('h8241)
	) name1911 (
		_w997_,
		_w1084_,
		_w2080_,
		_w2125_,
		_w2216_
	);
	LUT3 #(
		.INIT('h8c)
	) name1912 (
		_w2204_,
		_w2201_,
		_w2216_,
		_w2217_
	);
	LUT4 #(
		.INIT('h0e00)
	) name1913 (
		_w2211_,
		_w2212_,
		_w2215_,
		_w2217_,
		_w2218_
	);
	LUT3 #(
		.INIT('h08)
	) name1914 (
		_w2104_,
		_w2126_,
		_w2176_,
		_w2219_
	);
	LUT4 #(
		.INIT('h9009)
	) name1915 (
		_w1002_,
		_w2147_,
		_w2170_,
		_w2174_,
		_w2220_
	);
	LUT3 #(
		.INIT('h80)
	) name1916 (
		_w2126_,
		_w2207_,
		_w2220_,
		_w2221_
	);
	LUT2 #(
		.INIT('h1)
	) name1917 (
		_w2219_,
		_w2221_,
		_w2222_
	);
	LUT4 #(
		.INIT('hf400)
	) name1918 (
		_w2177_,
		_w2209_,
		_w2218_,
		_w2222_,
		_w2223_
	);
	LUT4 #(
		.INIT('h0100)
	) name1919 (
		\desIn[40]_pad ,
		\roundSel[4]_pad ,
		\roundSel[5]_pad ,
		_w305_,
		_w2224_
	);
	LUT4 #(
		.INIT('h2800)
	) name1920 (
		\FP_R_reg[30]/P0001 ,
		\roundSel[4]_pad ,
		\roundSel[5]_pad ,
		_w305_,
		_w2225_
	);
	LUT4 #(
		.INIT('h7c55)
	) name1921 (
		\FP_R_reg[62]/NET0131 ,
		\roundSel[4]_pad ,
		\roundSel[5]_pad ,
		_w305_,
		_w2226_
	);
	LUT3 #(
		.INIT('h45)
	) name1922 (
		_w2224_,
		_w2225_,
		_w2226_,
		_w2227_
	);
	LUT2 #(
		.INIT('h6)
	) name1923 (
		_w2223_,
		_w2227_,
		_w2228_
	);
	LUT4 #(
		.INIT('hff67)
	) name1924 (
		_w1523_,
		_w1545_,
		_w1573_,
		_w1601_,
		_w2229_
	);
	LUT4 #(
		.INIT('h8241)
	) name1925 (
		_w1338_,
		_w1495_,
		_w1499_,
		_w1544_,
		_w2230_
	);
	LUT4 #(
		.INIT('hd100)
	) name1926 (
		_w1523_,
		_w1573_,
		_w1643_,
		_w2230_,
		_w2231_
	);
	LUT4 #(
		.INIT('haebf)
	) name1927 (
		_w1523_,
		_w1573_,
		_w1602_,
		_w1634_,
		_w2232_
	);
	LUT4 #(
		.INIT('h0e00)
	) name1928 (
		_w1501_,
		_w2229_,
		_w2231_,
		_w2232_,
		_w2233_
	);
	LUT2 #(
		.INIT('h2)
	) name1929 (
		_w1629_,
		_w2233_,
		_w2234_
	);
	LUT2 #(
		.INIT('h8)
	) name1930 (
		_w1546_,
		_w1601_,
		_w2235_
	);
	LUT4 #(
		.INIT('h5efe)
	) name1931 (
		_w1545_,
		_w1573_,
		_w1601_,
		_w1605_,
		_w2236_
	);
	LUT3 #(
		.INIT('h45)
	) name1932 (
		_w1501_,
		_w2235_,
		_w2236_,
		_w2237_
	);
	LUT3 #(
		.INIT('h20)
	) name1933 (
		_w1573_,
		_w1633_,
		_w1634_,
		_w2238_
	);
	LUT3 #(
		.INIT('ha8)
	) name1934 (
		_w1574_,
		_w1604_,
		_w2230_,
		_w2239_
	);
	LUT3 #(
		.INIT('h10)
	) name1935 (
		_w1545_,
		_w1601_,
		_w1607_,
		_w2240_
	);
	LUT3 #(
		.INIT('h01)
	) name1936 (
		_w2239_,
		_w2240_,
		_w2238_,
		_w2241_
	);
	LUT3 #(
		.INIT('h45)
	) name1937 (
		_w1629_,
		_w2237_,
		_w2241_,
		_w2242_
	);
	LUT4 #(
		.INIT('h5d7f)
	) name1938 (
		_w1545_,
		_w1601_,
		_w1607_,
		_w1605_,
		_w2243_
	);
	LUT2 #(
		.INIT('h4)
	) name1939 (
		_w1523_,
		_w1604_,
		_w2244_
	);
	LUT3 #(
		.INIT('ha2)
	) name1940 (
		_w1501_,
		_w2243_,
		_w2244_,
		_w2245_
	);
	LUT3 #(
		.INIT('h10)
	) name1941 (
		_w1501_,
		_w1545_,
		_w1607_,
		_w2246_
	);
	LUT4 #(
		.INIT('h2184)
	) name1942 (
		_w1255_,
		_w1338_,
		_w1522_,
		_w1544_,
		_w2247_
	);
	LUT4 #(
		.INIT('hc480)
	) name1943 (
		_w1501_,
		_w1573_,
		_w1640_,
		_w2247_,
		_w2248_
	);
	LUT2 #(
		.INIT('h1)
	) name1944 (
		_w2246_,
		_w2248_,
		_w2249_
	);
	LUT2 #(
		.INIT('h4)
	) name1945 (
		_w2245_,
		_w2249_,
		_w2250_
	);
	LUT4 #(
		.INIT('h0100)
	) name1946 (
		\desIn[42]_pad ,
		\roundSel[4]_pad ,
		\roundSel[5]_pad ,
		_w305_,
		_w2251_
	);
	LUT4 #(
		.INIT('h2800)
	) name1947 (
		\FP_R_reg[22]/P0001 ,
		\roundSel[4]_pad ,
		\roundSel[5]_pad ,
		_w305_,
		_w2252_
	);
	LUT4 #(
		.INIT('h7c55)
	) name1948 (
		\FP_R_reg[54]/NET0131 ,
		\roundSel[4]_pad ,
		\roundSel[5]_pad ,
		_w305_,
		_w2253_
	);
	LUT3 #(
		.INIT('h45)
	) name1949 (
		_w2251_,
		_w2252_,
		_w2253_,
		_w2254_
	);
	LUT4 #(
		.INIT('h10ef)
	) name1950 (
		_w2242_,
		_w2234_,
		_w2250_,
		_w2254_,
		_w2255_
	);
	LUT2 #(
		.INIT('h8)
	) name1951 (
		_w626_,
		_w645_,
		_w2256_
	);
	LUT4 #(
		.INIT('h2fef)
	) name1952 (
		_w501_,
		_w528_,
		_w570_,
		_w631_,
		_w2257_
	);
	LUT4 #(
		.INIT('ha8aa)
	) name1953 (
		_w597_,
		_w1391_,
		_w2256_,
		_w2257_,
		_w2258_
	);
	LUT4 #(
		.INIT('h3edc)
	) name1954 (
		_w501_,
		_w528_,
		_w570_,
		_w626_,
		_w2259_
	);
	LUT4 #(
		.INIT('hbffd)
	) name1955 (
		_w501_,
		_w528_,
		_w570_,
		_w626_,
		_w2260_
	);
	LUT3 #(
		.INIT('he0)
	) name1956 (
		_w597_,
		_w2259_,
		_w2260_,
		_w2261_
	);
	LUT3 #(
		.INIT('h45)
	) name1957 (
		_w429_,
		_w2258_,
		_w2261_,
		_w2262_
	);
	LUT2 #(
		.INIT('h4)
	) name1958 (
		_w631_,
		_w648_,
		_w2263_
	);
	LUT4 #(
		.INIT('hf737)
	) name1959 (
		_w501_,
		_w528_,
		_w570_,
		_w626_,
		_w2264_
	);
	LUT3 #(
		.INIT('h45)
	) name1960 (
		_w597_,
		_w2263_,
		_w2264_,
		_w2265_
	);
	LUT4 #(
		.INIT('h0990)
	) name1961 (
		_w592_,
		_w596_,
		_w620_,
		_w624_,
		_w2266_
	);
	LUT4 #(
		.INIT('h2100)
	) name1962 (
		_w501_,
		_w528_,
		_w570_,
		_w2266_,
		_w2267_
	);
	LUT4 #(
		.INIT('h9669)
	) name1963 (
		_w495_,
		_w499_,
		_w620_,
		_w624_,
		_w2268_
	);
	LUT4 #(
		.INIT('hf7dd)
	) name1964 (
		_w528_,
		_w570_,
		_w1393_,
		_w2268_,
		_w2269_
	);
	LUT2 #(
		.INIT('h4)
	) name1965 (
		_w2267_,
		_w2269_,
		_w2270_
	);
	LUT4 #(
		.INIT('h1200)
	) name1966 (
		_w501_,
		_w528_,
		_w570_,
		_w626_,
		_w2271_
	);
	LUT4 #(
		.INIT('hfe54)
	) name1967 (
		_w597_,
		_w638_,
		_w1401_,
		_w2271_,
		_w2272_
	);
	LUT4 #(
		.INIT('h0075)
	) name1968 (
		_w429_,
		_w2265_,
		_w2270_,
		_w2272_,
		_w2273_
	);
	LUT4 #(
		.INIT('h0100)
	) name1969 (
		\desIn[44]_pad ,
		\roundSel[4]_pad ,
		\roundSel[5]_pad ,
		_w305_,
		_w2274_
	);
	LUT4 #(
		.INIT('h2800)
	) name1970 (
		\FP_R_reg[14]/P0001 ,
		\roundSel[4]_pad ,
		\roundSel[5]_pad ,
		_w305_,
		_w2275_
	);
	LUT4 #(
		.INIT('h7c55)
	) name1971 (
		\FP_R_reg[46]/NET0131 ,
		\roundSel[4]_pad ,
		\roundSel[5]_pad ,
		_w305_,
		_w2276_
	);
	LUT3 #(
		.INIT('h45)
	) name1972 (
		_w2274_,
		_w2275_,
		_w2276_,
		_w2277_
	);
	LUT3 #(
		.INIT('h4b)
	) name1973 (
		_w2262_,
		_w2273_,
		_w2277_,
		_w2278_
	);
	LUT4 #(
		.INIT('h6006)
	) name1974 (
		_w1002_,
		_w2147_,
		_w2170_,
		_w2174_,
		_w2279_
	);
	LUT4 #(
		.INIT('h4182)
	) name1975 (
		_w997_,
		_w1084_,
		_w2080_,
		_w2125_,
		_w2280_
	);
	LUT4 #(
		.INIT('he696)
	) name1976 (
		_w2081_,
		_w2126_,
		_w2205_,
		_w2279_,
		_w2281_
	);
	LUT2 #(
		.INIT('h1)
	) name1977 (
		_w2201_,
		_w2281_,
		_w2282_
	);
	LUT4 #(
		.INIT('hcfbb)
	) name1978 (
		_w2081_,
		_w2103_,
		_w2126_,
		_w2148_,
		_w2283_
	);
	LUT4 #(
		.INIT('hcd99)
	) name1979 (
		_w2081_,
		_w2103_,
		_w2126_,
		_w2148_,
		_w2284_
	);
	LUT2 #(
		.INIT('h8)
	) name1980 (
		_w2202_,
		_w2203_,
		_w2285_
	);
	LUT4 #(
		.INIT('hd5df)
	) name1981 (
		_w2081_,
		_w2103_,
		_w2126_,
		_w2203_,
		_w2286_
	);
	LUT4 #(
		.INIT('h08aa)
	) name1982 (
		_w2176_,
		_w2201_,
		_w2284_,
		_w2286_,
		_w2287_
	);
	LUT2 #(
		.INIT('h2)
	) name1983 (
		_w2148_,
		_w2280_,
		_w2288_
	);
	LUT4 #(
		.INIT('h2814)
	) name1984 (
		_w904_,
		_w2170_,
		_w2174_,
		_w2200_,
		_w2289_
	);
	LUT3 #(
		.INIT('h10)
	) name1985 (
		_w2104_,
		_w2207_,
		_w2289_,
		_w2290_
	);
	LUT4 #(
		.INIT('h8241)
	) name1986 (
		_w904_,
		_w1084_,
		_w2080_,
		_w2200_,
		_w2291_
	);
	LUT3 #(
		.INIT('h80)
	) name1987 (
		_w2126_,
		_w2203_,
		_w2291_,
		_w2292_
	);
	LUT3 #(
		.INIT('h0b)
	) name1988 (
		_w2288_,
		_w2290_,
		_w2292_,
		_w2293_
	);
	LUT4 #(
		.INIT('h0100)
	) name1989 (
		\desIn[46]_pad ,
		\roundSel[4]_pad ,
		\roundSel[5]_pad ,
		_w305_,
		_w2294_
	);
	LUT4 #(
		.INIT('h2800)
	) name1990 (
		\FP_R_reg[6]/P0001 ,
		\roundSel[4]_pad ,
		\roundSel[5]_pad ,
		_w305_,
		_w2295_
	);
	LUT4 #(
		.INIT('h7c55)
	) name1991 (
		\FP_R_reg[38]/NET0131 ,
		\roundSel[4]_pad ,
		\roundSel[5]_pad ,
		_w305_,
		_w2296_
	);
	LUT3 #(
		.INIT('h45)
	) name1992 (
		_w2294_,
		_w2295_,
		_w2296_,
		_w2297_
	);
	LUT4 #(
		.INIT('h10ef)
	) name1993 (
		_w2287_,
		_w2282_,
		_w2293_,
		_w2297_,
		_w2298_
	);
	LUT4 #(
		.INIT('h2814)
	) name1994 (
		_w1057_,
		_w1740_,
		_w1745_,
		_w1791_,
		_w2299_
	);
	LUT4 #(
		.INIT('haa20)
	) name1995 (
		_w1692_,
		_w1769_,
		_w1808_,
		_w2299_,
		_w2300_
	);
	LUT4 #(
		.INIT('h4182)
	) name1996 (
		_w1202_,
		_w1413_,
		_w1691_,
		_w1768_,
		_w2301_
	);
	LUT2 #(
		.INIT('h8)
	) name1997 (
		_w1804_,
		_w2301_,
		_w2302_
	);
	LUT4 #(
		.INIT('h0660)
	) name1998 (
		_w1713_,
		_w1717_,
		_w1740_,
		_w1745_,
		_w2303_
	);
	LUT4 #(
		.INIT('hbfbc)
	) name1999 (
		_w1692_,
		_w1719_,
		_w1747_,
		_w1769_,
		_w2304_
	);
	LUT3 #(
		.INIT('h80)
	) name2000 (
		_w1719_,
		_w1802_,
		_w1769_,
		_w2305_
	);
	LUT3 #(
		.INIT('h45)
	) name2001 (
		_w1670_,
		_w1747_,
		_w1804_,
		_w2306_
	);
	LUT4 #(
		.INIT('h1000)
	) name2002 (
		_w2302_,
		_w2305_,
		_w2306_,
		_w2304_,
		_w2307_
	);
	LUT4 #(
		.INIT('h8241)
	) name2003 (
		_w1202_,
		_w1413_,
		_w1691_,
		_w1768_,
		_w2308_
	);
	LUT3 #(
		.INIT('h40)
	) name2004 (
		_w1792_,
		_w1798_,
		_w2308_,
		_w2309_
	);
	LUT2 #(
		.INIT('h1)
	) name2005 (
		_w1794_,
		_w2309_,
		_w2310_
	);
	LUT2 #(
		.INIT('h8)
	) name2006 (
		_w1747_,
		_w1808_,
		_w2311_
	);
	LUT4 #(
		.INIT('h77cf)
	) name2007 (
		_w1692_,
		_w1719_,
		_w1747_,
		_w1792_,
		_w2312_
	);
	LUT4 #(
		.INIT('h2aaa)
	) name2008 (
		_w1670_,
		_w1747_,
		_w1804_,
		_w2308_,
		_w2313_
	);
	LUT3 #(
		.INIT('hd0)
	) name2009 (
		_w1769_,
		_w2312_,
		_w2313_,
		_w2314_
	);
	LUT4 #(
		.INIT('h0bbb)
	) name2010 (
		_w2300_,
		_w2307_,
		_w2310_,
		_w2314_,
		_w2315_
	);
	LUT3 #(
		.INIT('h20)
	) name2011 (
		_w1792_,
		_w1769_,
		_w2303_,
		_w2316_
	);
	LUT4 #(
		.INIT('hdd5f)
	) name2012 (
		_w1747_,
		_w1792_,
		_w1793_,
		_w1769_,
		_w2317_
	);
	LUT3 #(
		.INIT('h45)
	) name2013 (
		_w1692_,
		_w2316_,
		_w2317_,
		_w2318_
	);
	LUT4 #(
		.INIT('hf7a7)
	) name2014 (
		_w1719_,
		_w1802_,
		_w1769_,
		_w2299_,
		_w2319_
	);
	LUT3 #(
		.INIT('h40)
	) name2015 (
		_w1792_,
		_w2303_,
		_w2308_,
		_w2320_
	);
	LUT4 #(
		.INIT('h9009)
	) name2016 (
		_w1413_,
		_w1691_,
		_w1713_,
		_w1717_,
		_w2321_
	);
	LUT2 #(
		.INIT('h8)
	) name2017 (
		_w1770_,
		_w2321_,
		_w2322_
	);
	LUT4 #(
		.INIT('h000d)
	) name2018 (
		_w1807_,
		_w2319_,
		_w2320_,
		_w2322_,
		_w2323_
	);
	LUT2 #(
		.INIT('h4)
	) name2019 (
		_w2318_,
		_w2323_,
		_w2324_
	);
	LUT4 #(
		.INIT('h0100)
	) name2020 (
		\desIn[48]_pad ,
		\roundSel[4]_pad ,
		\roundSel[5]_pad ,
		_w305_,
		_w2325_
	);
	LUT4 #(
		.INIT('h2800)
	) name2021 (
		\FP_R_reg[31]/P0001 ,
		\roundSel[4]_pad ,
		\roundSel[5]_pad ,
		_w305_,
		_w2326_
	);
	LUT4 #(
		.INIT('h7c55)
	) name2022 (
		\FP_R_reg[63]/NET0131 ,
		\roundSel[4]_pad ,
		\roundSel[5]_pad ,
		_w305_,
		_w2327_
	);
	LUT3 #(
		.INIT('h45)
	) name2023 (
		_w2325_,
		_w2326_,
		_w2327_,
		_w2328_
	);
	LUT3 #(
		.INIT('h4b)
	) name2024 (
		_w2315_,
		_w2324_,
		_w2328_,
		_w2329_
	);
	LUT4 #(
		.INIT('h0096)
	) name2025 (
		_w1719_,
		_w1747_,
		_w1792_,
		_w1769_,
		_w2330_
	);
	LUT4 #(
		.INIT('hb100)
	) name2026 (
		_w1747_,
		_w1792_,
		_w1804_,
		_w2301_,
		_w2331_
	);
	LUT4 #(
		.INIT('h5554)
	) name2027 (
		_w1670_,
		_w1799_,
		_w2331_,
		_w2330_,
		_w2332_
	);
	LUT4 #(
		.INIT('h1054)
	) name2028 (
		_w1692_,
		_w1747_,
		_w1792_,
		_w1804_,
		_w2333_
	);
	LUT4 #(
		.INIT('h8a82)
	) name2029 (
		_w1692_,
		_w1747_,
		_w1792_,
		_w1769_,
		_w2334_
	);
	LUT4 #(
		.INIT('h7fde)
	) name2030 (
		_w1719_,
		_w1747_,
		_w1792_,
		_w1769_,
		_w2335_
	);
	LUT4 #(
		.INIT('hdc00)
	) name2031 (
		_w2311_,
		_w2333_,
		_w2334_,
		_w2335_,
		_w2336_
	);
	LUT4 #(
		.INIT('h7fbf)
	) name2032 (
		_w1719_,
		_w1747_,
		_w1792_,
		_w1769_,
		_w2337_
	);
	LUT2 #(
		.INIT('h1)
	) name2033 (
		_w1692_,
		_w2337_,
		_w2338_
	);
	LUT4 #(
		.INIT('h000d)
	) name2034 (
		_w1670_,
		_w2336_,
		_w2338_,
		_w2332_,
		_w2339_
	);
	LUT4 #(
		.INIT('h0100)
	) name2035 (
		\desIn[4]_pad ,
		\roundSel[4]_pad ,
		\roundSel[5]_pad ,
		_w305_,
		_w2340_
	);
	LUT4 #(
		.INIT('h2800)
	) name2036 (
		\FP_R_reg[9]/P0001 ,
		\roundSel[4]_pad ,
		\roundSel[5]_pad ,
		_w305_,
		_w2341_
	);
	LUT4 #(
		.INIT('h7c55)
	) name2037 (
		\FP_R_reg[41]/NET0131 ,
		\roundSel[4]_pad ,
		\roundSel[5]_pad ,
		_w305_,
		_w2342_
	);
	LUT3 #(
		.INIT('h45)
	) name2038 (
		_w2340_,
		_w2341_,
		_w2342_,
		_w2343_
	);
	LUT2 #(
		.INIT('h9)
	) name2039 (
		_w2339_,
		_w2343_,
		_w2344_
	);
	LUT4 #(
		.INIT('h5504)
	) name2040 (
		_w1692_,
		_w1793_,
		_w1769_,
		_w1798_,
		_w2345_
	);
	LUT3 #(
		.INIT('h80)
	) name2041 (
		_w1692_,
		_w1747_,
		_w1808_,
		_w2346_
	);
	LUT2 #(
		.INIT('h8)
	) name2042 (
		_w1804_,
		_w2308_,
		_w2347_
	);
	LUT3 #(
		.INIT('he7)
	) name2043 (
		_w1747_,
		_w1792_,
		_w1769_,
		_w2348_
	);
	LUT4 #(
		.INIT('h0100)
	) name2044 (
		_w2345_,
		_w2346_,
		_w2347_,
		_w2348_,
		_w2349_
	);
	LUT2 #(
		.INIT('h2)
	) name2045 (
		_w1670_,
		_w2349_,
		_w2350_
	);
	LUT3 #(
		.INIT('h80)
	) name2046 (
		_w1692_,
		_w1747_,
		_w1804_,
		_w2351_
	);
	LUT4 #(
		.INIT('h0001)
	) name2047 (
		_w1794_,
		_w2309_,
		_w2320_,
		_w2351_,
		_w2352_
	);
	LUT4 #(
		.INIT('hebe9)
	) name2048 (
		_w1719_,
		_w1747_,
		_w1792_,
		_w1769_,
		_w2353_
	);
	LUT4 #(
		.INIT('h2184)
	) name2049 (
		_w1111_,
		_w1413_,
		_w1669_,
		_w1691_,
		_w2354_
	);
	LUT2 #(
		.INIT('h4)
	) name2050 (
		_w2353_,
		_w2354_,
		_w2355_
	);
	LUT4 #(
		.INIT('h8000)
	) name2051 (
		_w1692_,
		_w1747_,
		_w1769_,
		_w1808_,
		_w2356_
	);
	LUT4 #(
		.INIT('h1428)
	) name2052 (
		_w1202_,
		_w1413_,
		_w1691_,
		_w1768_,
		_w2357_
	);
	LUT4 #(
		.INIT('h1800)
	) name2053 (
		_w1719_,
		_w1747_,
		_w1792_,
		_w2357_,
		_w2358_
	);
	LUT3 #(
		.INIT('h40)
	) name2054 (
		_w1692_,
		_w1793_,
		_w1797_,
		_w2359_
	);
	LUT4 #(
		.INIT('h0001)
	) name2055 (
		_w2322_,
		_w2358_,
		_w2359_,
		_w2356_,
		_w2360_
	);
	LUT4 #(
		.INIT('h0e00)
	) name2056 (
		_w1670_,
		_w2352_,
		_w2355_,
		_w2360_,
		_w2361_
	);
	LUT4 #(
		.INIT('h0100)
	) name2057 (
		\desIn[50]_pad ,
		\roundSel[4]_pad ,
		\roundSel[5]_pad ,
		_w305_,
		_w2362_
	);
	LUT4 #(
		.INIT('h2800)
	) name2058 (
		\FP_R_reg[23]/P0001 ,
		\roundSel[4]_pad ,
		\roundSel[5]_pad ,
		_w305_,
		_w2363_
	);
	LUT4 #(
		.INIT('h7c55)
	) name2059 (
		\FP_R_reg[55]/NET0131 ,
		\roundSel[4]_pad ,
		\roundSel[5]_pad ,
		_w305_,
		_w2364_
	);
	LUT3 #(
		.INIT('h45)
	) name2060 (
		_w2362_,
		_w2363_,
		_w2364_,
		_w2365_
	);
	LUT3 #(
		.INIT('hb4)
	) name2061 (
		_w2350_,
		_w2361_,
		_w2365_,
		_w2366_
	);
	LUT4 #(
		.INIT('h33bc)
	) name2062 (
		_w1958_,
		_w1980_,
		_w1931_,
		_w2003_,
		_w2367_
	);
	LUT2 #(
		.INIT('h8)
	) name2063 (
		_w1981_,
		_w2008_,
		_w2368_
	);
	LUT4 #(
		.INIT('h5504)
	) name2064 (
		_w1882_,
		_w1909_,
		_w2367_,
		_w2368_,
		_w2369_
	);
	LUT2 #(
		.INIT('h8)
	) name2065 (
		_w2023_,
		_w2044_,
		_w2370_
	);
	LUT4 #(
		.INIT('h9dbf)
	) name2066 (
		_w1958_,
		_w1980_,
		_w2003_,
		_w2011_,
		_w2371_
	);
	LUT3 #(
		.INIT('h20)
	) name2067 (
		_w1909_,
		_w1980_,
		_w2004_,
		_w2372_
	);
	LUT3 #(
		.INIT('h80)
	) name2068 (
		_w1980_,
		_w1931_,
		_w2018_,
		_w2373_
	);
	LUT4 #(
		.INIT('h0100)
	) name2069 (
		_w2372_,
		_w2370_,
		_w2373_,
		_w2371_,
		_w2374_
	);
	LUT4 #(
		.INIT('h1428)
	) name2070 (
		_w1599_,
		_w1717_,
		_w1881_,
		_w1979_,
		_w2375_
	);
	LUT4 #(
		.INIT('h13df)
	) name2071 (
		_w1931_,
		_w2003_,
		_w1981_,
		_w2375_,
		_w2376_
	);
	LUT4 #(
		.INIT('hff7b)
	) name2072 (
		_w1958_,
		_w1980_,
		_w1931_,
		_w2003_,
		_w2377_
	);
	LUT3 #(
		.INIT('h80)
	) name2073 (
		_w2040_,
		_w2376_,
		_w2377_,
		_w2378_
	);
	LUT4 #(
		.INIT('ha8aa)
	) name2074 (
		_w1909_,
		_w1931_,
		_w2003_,
		_w1981_,
		_w2379_
	);
	LUT2 #(
		.INIT('h4)
	) name2075 (
		_w2042_,
		_w2379_,
		_w2380_
	);
	LUT4 #(
		.INIT('hddd0)
	) name2076 (
		_w1882_,
		_w2374_,
		_w2378_,
		_w2380_,
		_w2381_
	);
	LUT4 #(
		.INIT('h0100)
	) name2077 (
		\desIn[52]_pad ,
		\roundSel[4]_pad ,
		\roundSel[5]_pad ,
		_w305_,
		_w2382_
	);
	LUT4 #(
		.INIT('h2800)
	) name2078 (
		\FP_R_reg[15]/P0001 ,
		\roundSel[4]_pad ,
		\roundSel[5]_pad ,
		_w305_,
		_w2383_
	);
	LUT4 #(
		.INIT('h7c55)
	) name2079 (
		\FP_R_reg[47]/NET0131 ,
		\roundSel[4]_pad ,
		\roundSel[5]_pad ,
		_w305_,
		_w2384_
	);
	LUT3 #(
		.INIT('h45)
	) name2080 (
		_w2382_,
		_w2383_,
		_w2384_,
		_w2385_
	);
	LUT3 #(
		.INIT('h4b)
	) name2081 (
		_w2369_,
		_w2381_,
		_w2385_,
		_w2386_
	);
	LUT4 #(
		.INIT('h0100)
	) name2082 (
		\desIn[54]_pad ,
		\roundSel[4]_pad ,
		\roundSel[5]_pad ,
		_w305_,
		_w2387_
	);
	LUT4 #(
		.INIT('h2800)
	) name2083 (
		\FP_R_reg[7]/P0001 ,
		\roundSel[4]_pad ,
		\roundSel[5]_pad ,
		_w305_,
		_w2388_
	);
	LUT4 #(
		.INIT('h7c55)
	) name2084 (
		\FP_R_reg[39]/NET0131 ,
		\roundSel[4]_pad ,
		\roundSel[5]_pad ,
		_w305_,
		_w2389_
	);
	LUT3 #(
		.INIT('h45)
	) name2085 (
		_w2387_,
		_w2388_,
		_w2389_,
		_w2390_
	);
	LUT2 #(
		.INIT('h8)
	) name2086 (
		_w1605_,
		_w1631_,
		_w2391_
	);
	LUT2 #(
		.INIT('h1)
	) name2087 (
		_w1607_,
		_w1638_,
		_w2392_
	);
	LUT4 #(
		.INIT('h8c22)
	) name2088 (
		_w1523_,
		_w1573_,
		_w1601_,
		_w1638_,
		_w2393_
	);
	LUT4 #(
		.INIT('h2814)
	) name2089 (
		_w1444_,
		_w1495_,
		_w1499_,
		_w1628_,
		_w2394_
	);
	LUT4 #(
		.INIT('h4182)
	) name2090 (
		_w1444_,
		_w1495_,
		_w1499_,
		_w1628_,
		_w2395_
	);
	LUT4 #(
		.INIT('h9669)
	) name2091 (
		_w1444_,
		_w1495_,
		_w1499_,
		_w1628_,
		_w2396_
	);
	LUT3 #(
		.INIT('h70)
	) name2092 (
		_w1602_,
		_w1605_,
		_w2396_,
		_w2397_
	);
	LUT2 #(
		.INIT('h4)
	) name2093 (
		_w2393_,
		_w2397_,
		_w2398_
	);
	LUT2 #(
		.INIT('h2)
	) name2094 (
		_w1545_,
		_w1637_,
		_w2399_
	);
	LUT2 #(
		.INIT('h2)
	) name2095 (
		_w1523_,
		_w1638_,
		_w2400_
	);
	LUT3 #(
		.INIT('hb0)
	) name2096 (
		_w1573_,
		_w1604_,
		_w2394_,
		_w2401_
	);
	LUT3 #(
		.INIT('h10)
	) name2097 (
		_w2400_,
		_w2399_,
		_w2401_,
		_w2402_
	);
	LUT3 #(
		.INIT('hb0)
	) name2098 (
		_w1573_,
		_w1602_,
		_w2395_,
		_w2403_
	);
	LUT3 #(
		.INIT('h10)
	) name2099 (
		_w2240_,
		_w2392_,
		_w2403_,
		_w2404_
	);
	LUT4 #(
		.INIT('h00ab)
	) name2100 (
		_w2391_,
		_w2398_,
		_w2402_,
		_w2404_,
		_w2405_
	);
	LUT2 #(
		.INIT('h6)
	) name2101 (
		_w2390_,
		_w2405_,
		_w2406_
	);
	LUT4 #(
		.INIT('hb85f)
	) name2102 (
		_w1523_,
		_w1545_,
		_w1573_,
		_w1601_,
		_w2407_
	);
	LUT2 #(
		.INIT('h2)
	) name2103 (
		_w1501_,
		_w2407_,
		_w2408_
	);
	LUT3 #(
		.INIT('h40)
	) name2104 (
		_w1545_,
		_w1601_,
		_w1607_,
		_w2409_
	);
	LUT2 #(
		.INIT('h2)
	) name2105 (
		_w1574_,
		_w1638_,
		_w2410_
	);
	LUT4 #(
		.INIT('h4e5f)
	) name2106 (
		_w1523_,
		_w1573_,
		_w1602_,
		_w1631_,
		_w2411_
	);
	LUT4 #(
		.INIT('h2322)
	) name2107 (
		_w1501_,
		_w2409_,
		_w2410_,
		_w2411_,
		_w2412_
	);
	LUT3 #(
		.INIT('h8a)
	) name2108 (
		_w1629_,
		_w2408_,
		_w2412_,
		_w2413_
	);
	LUT3 #(
		.INIT('h80)
	) name2109 (
		_w1523_,
		_w1573_,
		_w1604_,
		_w2414_
	);
	LUT4 #(
		.INIT('h4d6f)
	) name2110 (
		_w1545_,
		_w1601_,
		_w1607_,
		_w1605_,
		_w2415_
	);
	LUT2 #(
		.INIT('h4)
	) name2111 (
		_w2414_,
		_w2415_,
		_w2416_
	);
	LUT4 #(
		.INIT('hcfee)
	) name2112 (
		_w1523_,
		_w1545_,
		_w1573_,
		_w1601_,
		_w2417_
	);
	LUT4 #(
		.INIT('h0015)
	) name2113 (
		_w1501_,
		_w1573_,
		_w1604_,
		_w1644_,
		_w2418_
	);
	LUT3 #(
		.INIT('h0d)
	) name2114 (
		_w1501_,
		_w2417_,
		_w2418_,
		_w2419_
	);
	LUT3 #(
		.INIT('h80)
	) name2115 (
		_w1501_,
		_w1605_,
		_w1634_,
		_w2420_
	);
	LUT4 #(
		.INIT('hf7d7)
	) name2116 (
		_w1523_,
		_w1545_,
		_w1573_,
		_w1601_,
		_w2421_
	);
	LUT3 #(
		.INIT('h32)
	) name2117 (
		_w1501_,
		_w2420_,
		_w2421_,
		_w2422_
	);
	LUT4 #(
		.INIT('hea00)
	) name2118 (
		_w1629_,
		_w2416_,
		_w2419_,
		_w2422_,
		_w2423_
	);
	LUT4 #(
		.INIT('h0100)
	) name2119 (
		\desIn[56]_pad ,
		\roundSel[4]_pad ,
		\roundSel[5]_pad ,
		_w305_,
		_w2424_
	);
	LUT4 #(
		.INIT('h2800)
	) name2120 (
		\FP_R_reg[32]/P0001 ,
		\roundSel[4]_pad ,
		\roundSel[5]_pad ,
		_w305_,
		_w2425_
	);
	LUT4 #(
		.INIT('h7c55)
	) name2121 (
		\FP_R_reg[64]/NET0131 ,
		\roundSel[4]_pad ,
		\roundSel[5]_pad ,
		_w305_,
		_w2426_
	);
	LUT3 #(
		.INIT('h45)
	) name2122 (
		_w2424_,
		_w2425_,
		_w2426_,
		_w2427_
	);
	LUT3 #(
		.INIT('h4b)
	) name2123 (
		_w2413_,
		_w2423_,
		_w2427_,
		_w2428_
	);
	LUT4 #(
		.INIT('hd1ee)
	) name2124 (
		_w2081_,
		_w2103_,
		_w2126_,
		_w2148_,
		_w2429_
	);
	LUT2 #(
		.INIT('h8)
	) name2125 (
		_w2081_,
		_w2149_,
		_w2430_
	);
	LUT3 #(
		.INIT('h7d)
	) name2126 (
		_w2103_,
		_w2126_,
		_w2148_,
		_w2431_
	);
	LUT4 #(
		.INIT('h0e04)
	) name2127 (
		_w2201_,
		_w2429_,
		_w2430_,
		_w2431_,
		_w2432_
	);
	LUT4 #(
		.INIT('h92d6)
	) name2128 (
		_w2081_,
		_w2103_,
		_w2148_,
		_w2279_,
		_w2433_
	);
	LUT3 #(
		.INIT('h40)
	) name2129 (
		_w2081_,
		_w2126_,
		_w2210_,
		_w2434_
	);
	LUT4 #(
		.INIT('hcc04)
	) name2130 (
		_w2126_,
		_w2201_,
		_w2433_,
		_w2434_,
		_w2435_
	);
	LUT4 #(
		.INIT('h1600)
	) name2131 (
		_w2081_,
		_w2103_,
		_w2148_,
		_w2176_,
		_w2436_
	);
	LUT4 #(
		.INIT('h9009)
	) name2132 (
		_w997_,
		_w2125_,
		_w2170_,
		_w2174_,
		_w2437_
	);
	LUT4 #(
		.INIT('h8400)
	) name2133 (
		_w2081_,
		_w2103_,
		_w2148_,
		_w2437_,
		_w2438_
	);
	LUT4 #(
		.INIT('h00ab)
	) name2134 (
		_w2201_,
		_w2285_,
		_w2436_,
		_w2438_,
		_w2439_
	);
	LUT4 #(
		.INIT('h3200)
	) name2135 (
		_w2176_,
		_w2435_,
		_w2432_,
		_w2439_,
		_w2440_
	);
	LUT4 #(
		.INIT('h0100)
	) name2136 (
		\desIn[60]_pad ,
		\roundSel[4]_pad ,
		\roundSel[5]_pad ,
		_w305_,
		_w2441_
	);
	LUT4 #(
		.INIT('h2800)
	) name2137 (
		\FP_R_reg[16]/P0001 ,
		\roundSel[4]_pad ,
		\roundSel[5]_pad ,
		_w305_,
		_w2442_
	);
	LUT4 #(
		.INIT('h7c55)
	) name2138 (
		\FP_R_reg[48]/NET0131 ,
		\roundSel[4]_pad ,
		\roundSel[5]_pad ,
		_w305_,
		_w2443_
	);
	LUT3 #(
		.INIT('h45)
	) name2139 (
		_w2441_,
		_w2442_,
		_w2443_,
		_w2444_
	);
	LUT2 #(
		.INIT('h9)
	) name2140 (
		_w2440_,
		_w2444_,
		_w2445_
	);
	LUT3 #(
		.INIT('h4c)
	) name2141 (
		_w877_,
		_w956_,
		_w962_,
		_w2446_
	);
	LUT2 #(
		.INIT('h8)
	) name2142 (
		_w928_,
		_w1449_,
		_w2447_
	);
	LUT3 #(
		.INIT('h13)
	) name2143 (
		_w877_,
		_w956_,
		_w929_,
		_w2448_
	);
	LUT4 #(
		.INIT('hb0bb)
	) name2144 (
		_w1461_,
		_w2446_,
		_w2447_,
		_w2448_,
		_w2449_
	);
	LUT3 #(
		.INIT('h80)
	) name2145 (
		_w820_,
		_w877_,
		_w929_,
		_w2450_
	);
	LUT2 #(
		.INIT('h2)
	) name2146 (
		_w1446_,
		_w2450_,
		_w2451_
	);
	LUT3 #(
		.INIT('h45)
	) name2147 (
		_w763_,
		_w2449_,
		_w2451_,
		_w2452_
	);
	LUT2 #(
		.INIT('h1)
	) name2148 (
		_w877_,
		_w957_,
		_w2453_
	);
	LUT3 #(
		.INIT('h02)
	) name2149 (
		_w820_,
		_w956_,
		_w929_,
		_w2454_
	);
	LUT3 #(
		.INIT('h20)
	) name2150 (
		_w820_,
		_w877_,
		_w929_,
		_w2455_
	);
	LUT4 #(
		.INIT('hfef6)
	) name2151 (
		_w906_,
		_w820_,
		_w877_,
		_w928_,
		_w2456_
	);
	LUT4 #(
		.INIT('h20aa)
	) name2152 (
		_w763_,
		_w2453_,
		_w2454_,
		_w2456_,
		_w2457_
	);
	LUT3 #(
		.INIT('h8a)
	) name2153 (
		_w956_,
		_w979_,
		_w961_,
		_w2458_
	);
	LUT2 #(
		.INIT('h8)
	) name2154 (
		_w877_,
		_w1449_,
		_w2459_
	);
	LUT4 #(
		.INIT('h9009)
	) name2155 (
		_w526_,
		_w762_,
		_w950_,
		_w954_,
		_w2460_
	);
	LUT4 #(
		.INIT('hec00)
	) name2156 (
		_w877_,
		_w1458_,
		_w1449_,
		_w2460_,
		_w2461_
	);
	LUT4 #(
		.INIT('h0200)
	) name2157 (
		_w820_,
		_w877_,
		_w956_,
		_w929_,
		_w2462_
	);
	LUT3 #(
		.INIT('h01)
	) name2158 (
		_w1448_,
		_w2462_,
		_w2461_,
		_w2463_
	);
	LUT3 #(
		.INIT('h10)
	) name2159 (
		_w2458_,
		_w2457_,
		_w2463_,
		_w2464_
	);
	LUT4 #(
		.INIT('h0100)
	) name2160 (
		\desIn[6]_pad ,
		\roundSel[4]_pad ,
		\roundSel[5]_pad ,
		_w305_,
		_w2465_
	);
	LUT4 #(
		.INIT('h2800)
	) name2161 (
		\FP_R_reg[1]/P0001 ,
		\roundSel[4]_pad ,
		\roundSel[5]_pad ,
		_w305_,
		_w2466_
	);
	LUT4 #(
		.INIT('h7c55)
	) name2162 (
		\FP_R_reg[33]/NET0131 ,
		\roundSel[4]_pad ,
		\roundSel[5]_pad ,
		_w305_,
		_w2467_
	);
	LUT3 #(
		.INIT('h45)
	) name2163 (
		_w2465_,
		_w2466_,
		_w2467_,
		_w2468_
	);
	LUT3 #(
		.INIT('h4b)
	) name2164 (
		_w2452_,
		_w2464_,
		_w2468_,
		_w2469_
	);
	LUT4 #(
		.INIT('h0100)
	) name2165 (
		\desIn[8]_pad ,
		\roundSel[4]_pad ,
		\roundSel[5]_pad ,
		_w305_,
		_w2470_
	);
	LUT4 #(
		.INIT('h2800)
	) name2166 (
		\FP_R_reg[26]/P0001 ,
		\roundSel[4]_pad ,
		\roundSel[5]_pad ,
		_w305_,
		_w2471_
	);
	LUT4 #(
		.INIT('h7c55)
	) name2167 (
		\FP_R_reg[58]/NET0131 ,
		\roundSel[4]_pad ,
		\roundSel[5]_pad ,
		_w305_,
		_w2472_
	);
	LUT3 #(
		.INIT('h45)
	) name2168 (
		_w2470_,
		_w2471_,
		_w2472_,
		_w2473_
	);
	LUT4 #(
		.INIT('h8fdf)
	) name2169 (
		_w906_,
		_w877_,
		_w928_,
		_w965_,
		_w2474_
	);
	LUT2 #(
		.INIT('h1)
	) name2170 (
		_w956_,
		_w2474_,
		_w2475_
	);
	LUT3 #(
		.INIT('hc8)
	) name2171 (
		_w878_,
		_w962_,
		_w1455_,
		_w2476_
	);
	LUT3 #(
		.INIT('h04)
	) name2172 (
		_w877_,
		_w957_,
		_w973_,
		_w2477_
	);
	LUT3 #(
		.INIT('h01)
	) name2173 (
		_w2455_,
		_w2477_,
		_w2476_,
		_w2478_
	);
	LUT3 #(
		.INIT('h8a)
	) name2174 (
		_w763_,
		_w2475_,
		_w2478_,
		_w2479_
	);
	LUT3 #(
		.INIT('h10)
	) name2175 (
		_w877_,
		_w957_,
		_w963_,
		_w2480_
	);
	LUT4 #(
		.INIT('hb5bf)
	) name2176 (
		_w906_,
		_w878_,
		_w928_,
		_w963_,
		_w2481_
	);
	LUT4 #(
		.INIT('h5455)
	) name2177 (
		_w763_,
		_w2459_,
		_w2480_,
		_w2481_,
		_w2482_
	);
	LUT4 #(
		.INIT('h0660)
	) name2178 (
		_w526_,
		_w762_,
		_w950_,
		_w954_,
		_w2483_
	);
	LUT4 #(
		.INIT('hf400)
	) name2179 (
		_w906_,
		_w960_,
		_w971_,
		_w2483_,
		_w2484_
	);
	LUT3 #(
		.INIT('h80)
	) name2180 (
		_w878_,
		_w956_,
		_w957_,
		_w2485_
	);
	LUT3 #(
		.INIT('h80)
	) name2181 (
		_w877_,
		_w973_,
		_w929_,
		_w2486_
	);
	LUT4 #(
		.INIT('h0084)
	) name2182 (
		_w906_,
		_w878_,
		_w928_,
		_w956_,
		_w2487_
	);
	LUT4 #(
		.INIT('h0001)
	) name2183 (
		_w967_,
		_w2485_,
		_w2486_,
		_w2487_,
		_w2488_
	);
	LUT3 #(
		.INIT('h10)
	) name2184 (
		_w2482_,
		_w2484_,
		_w2488_,
		_w2489_
	);
	LUT3 #(
		.INIT('h65)
	) name2185 (
		_w2473_,
		_w2479_,
		_w2489_,
		_w2490_
	);
	LUT4 #(
		.INIT('hcdef)
	) name2186 (
		_w1162_,
		_w1080_,
		_w1169_,
		_w1179_,
		_w2491_
	);
	LUT3 #(
		.INIT('h23)
	) name2187 (
		_w1080_,
		_w1053_,
		_w1187_,
		_w2492_
	);
	LUT4 #(
		.INIT('h67ef)
	) name2188 (
		_w1107_,
		_w1134_,
		_w1168_,
		_w1171_,
		_w2493_
	);
	LUT3 #(
		.INIT('h80)
	) name2189 (
		_w2491_,
		_w2492_,
		_w2493_,
		_w2494_
	);
	LUT3 #(
		.INIT('h8c)
	) name2190 (
		_w1166_,
		_w1053_,
		_w1163_,
		_w2495_
	);
	LUT2 #(
		.INIT('h4)
	) name2191 (
		_w1425_,
		_w2495_,
		_w2496_
	);
	LUT3 #(
		.INIT('ha8)
	) name2192 (
		_w1135_,
		_w1177_,
		_w1421_,
		_w2497_
	);
	LUT4 #(
		.INIT('h2aaa)
	) name2193 (
		_w1025_,
		_w1166_,
		_w1134_,
		_w1421_,
		_w2498_
	);
	LUT2 #(
		.INIT('h4)
	) name2194 (
		_w2497_,
		_w2498_,
		_w2499_
	);
	LUT3 #(
		.INIT('he0)
	) name2195 (
		_w2494_,
		_w2496_,
		_w2499_,
		_w2500_
	);
	LUT4 #(
		.INIT('h0f0d)
	) name2196 (
		_w1080_,
		_w1135_,
		_w1053_,
		_w1417_,
		_w2501_
	);
	LUT2 #(
		.INIT('h8)
	) name2197 (
		_w1162_,
		_w1135_,
		_w2502_
	);
	LUT3 #(
		.INIT('h4c)
	) name2198 (
		_w1107_,
		_w1053_,
		_w1171_,
		_w2503_
	);
	LUT3 #(
		.INIT('h45)
	) name2199 (
		_w2501_,
		_w2502_,
		_w2503_,
		_w2504_
	);
	LUT3 #(
		.INIT('h10)
	) name2200 (
		_w1162_,
		_w1080_,
		_w1187_,
		_w2505_
	);
	LUT4 #(
		.INIT('h0040)
	) name2201 (
		_w1025_,
		_w1173_,
		_w2491_,
		_w2505_,
		_w2506_
	);
	LUT2 #(
		.INIT('h4)
	) name2202 (
		_w2504_,
		_w2506_,
		_w2507_
	);
	LUT4 #(
		.INIT('h0100)
	) name2203 (
		\desIn[36]_pad ,
		\roundSel[4]_pad ,
		\roundSel[5]_pad ,
		_w305_,
		_w2508_
	);
	LUT4 #(
		.INIT('h2800)
	) name2204 (
		\FP_R_reg[13]/P0001 ,
		\roundSel[4]_pad ,
		\roundSel[5]_pad ,
		_w305_,
		_w2509_
	);
	LUT4 #(
		.INIT('h7c55)
	) name2205 (
		\FP_R_reg[45]/NET0131 ,
		\roundSel[4]_pad ,
		\roundSel[5]_pad ,
		_w305_,
		_w2510_
	);
	LUT3 #(
		.INIT('h45)
	) name2206 (
		_w2508_,
		_w2509_,
		_w2510_,
		_w2511_
	);
	LUT3 #(
		.INIT('h1e)
	) name2207 (
		_w2500_,
		_w2507_,
		_w2511_,
		_w2512_
	);
	LUT4 #(
		.INIT('he400)
	) name2208 (
		_w1080_,
		_w1107_,
		_w1135_,
		_w1053_,
		_w2513_
	);
	LUT4 #(
		.INIT('h3aff)
	) name2209 (
		_w1162_,
		_w1080_,
		_w1107_,
		_w1134_,
		_w2514_
	);
	LUT4 #(
		.INIT('h0032)
	) name2210 (
		_w1053_,
		_w1183_,
		_w2514_,
		_w2513_,
		_w2515_
	);
	LUT3 #(
		.INIT('h80)
	) name2211 (
		_w1134_,
		_w1053_,
		_w1180_,
		_w2516_
	);
	LUT4 #(
		.INIT('h5d7f)
	) name2212 (
		_w1162_,
		_w1080_,
		_w1169_,
		_w1179_,
		_w2517_
	);
	LUT4 #(
		.INIT('hd9fb)
	) name2213 (
		_w1162_,
		_w1080_,
		_w1169_,
		_w1418_,
		_w2518_
	);
	LUT3 #(
		.INIT('h40)
	) name2214 (
		_w2516_,
		_w2517_,
		_w2518_,
		_w2519_
	);
	LUT4 #(
		.INIT('hf5ef)
	) name2215 (
		_w1162_,
		_w1080_,
		_w1107_,
		_w1134_,
		_w2520_
	);
	LUT2 #(
		.INIT('h8)
	) name2216 (
		_w1180_,
		_w1418_,
		_w2521_
	);
	LUT3 #(
		.INIT('h0d)
	) name2217 (
		_w1053_,
		_w2520_,
		_w2521_,
		_w2522_
	);
	LUT4 #(
		.INIT('hd800)
	) name2218 (
		_w1025_,
		_w2519_,
		_w2515_,
		_w2522_,
		_w2523_
	);
	LUT4 #(
		.INIT('h0100)
	) name2219 (
		\desIn[10]_pad ,
		\roundSel[4]_pad ,
		\roundSel[5]_pad ,
		_w305_,
		_w2524_
	);
	LUT4 #(
		.INIT('h2800)
	) name2220 (
		\FP_R_reg[18]/P0001 ,
		\roundSel[4]_pad ,
		\roundSel[5]_pad ,
		_w305_,
		_w2525_
	);
	LUT4 #(
		.INIT('h7c55)
	) name2221 (
		\FP_R_reg[50]/NET0131 ,
		\roundSel[4]_pad ,
		\roundSel[5]_pad ,
		_w305_,
		_w2526_
	);
	LUT3 #(
		.INIT('h45)
	) name2222 (
		_w2524_,
		_w2525_,
		_w2526_,
		_w2527_
	);
	LUT2 #(
		.INIT('h9)
	) name2223 (
		_w2523_,
		_w2527_,
		_w2528_
	);
	LUT4 #(
		.INIT('hd9fb)
	) name2224 (
		_w1331_,
		_w1301_,
		_w1257_,
		_w1230_,
		_w2529_
	);
	LUT4 #(
		.INIT('h0301)
	) name2225 (
		_w1279_,
		_w1819_,
		_w1848_,
		_w2529_,
		_w2530_
	);
	LUT4 #(
		.INIT('h0060)
	) name2226 (
		_w1279_,
		_w1331_,
		_w1301_,
		_w1230_,
		_w2531_
	);
	LUT4 #(
		.INIT('hcc80)
	) name2227 (
		_w1257_,
		_w1230_,
		_w1364_,
		_w1826_,
		_w2532_
	);
	LUT2 #(
		.INIT('h1)
	) name2228 (
		_w2531_,
		_w2532_,
		_w2533_
	);
	LUT3 #(
		.INIT('h15)
	) name2229 (
		_w1361_,
		_w2530_,
		_w2533_,
		_w2534_
	);
	LUT4 #(
		.INIT('h2133)
	) name2230 (
		_w1279_,
		_w1331_,
		_w1301_,
		_w1257_,
		_w2535_
	);
	LUT4 #(
		.INIT('h1113)
	) name2231 (
		_w1331_,
		_w1230_,
		_w1302_,
		_w1379_,
		_w2536_
	);
	LUT2 #(
		.INIT('h4)
	) name2232 (
		_w2535_,
		_w2536_,
		_w2537_
	);
	LUT4 #(
		.INIT('hbcbf)
	) name2233 (
		_w1279_,
		_w1331_,
		_w1301_,
		_w1378_,
		_w2538_
	);
	LUT3 #(
		.INIT('h8a)
	) name2234 (
		_w1230_,
		_w1833_,
		_w2538_,
		_w2539_
	);
	LUT4 #(
		.INIT('h77ef)
	) name2235 (
		_w1279_,
		_w1331_,
		_w1301_,
		_w1257_,
		_w2540_
	);
	LUT4 #(
		.INIT('he040)
	) name2236 (
		_w1301_,
		_w1303_,
		_w1377_,
		_w1378_,
		_w2541_
	);
	LUT4 #(
		.INIT('h0301)
	) name2237 (
		_w1230_,
		_w1376_,
		_w2541_,
		_w2540_,
		_w2542_
	);
	LUT4 #(
		.INIT('h5700)
	) name2238 (
		_w1361_,
		_w2537_,
		_w2539_,
		_w2542_,
		_w2543_
	);
	LUT4 #(
		.INIT('h0100)
	) name2239 (
		\desIn[20]_pad ,
		\roundSel[4]_pad ,
		\roundSel[5]_pad ,
		_w305_,
		_w2544_
	);
	LUT4 #(
		.INIT('h2800)
	) name2240 (
		\FP_R_reg[11]/P0001 ,
		\roundSel[4]_pad ,
		\roundSel[5]_pad ,
		_w305_,
		_w2545_
	);
	LUT4 #(
		.INIT('h7c55)
	) name2241 (
		\FP_R_reg[43]/NET0131 ,
		\roundSel[4]_pad ,
		\roundSel[5]_pad ,
		_w305_,
		_w2546_
	);
	LUT3 #(
		.INIT('h45)
	) name2242 (
		_w2544_,
		_w2545_,
		_w2546_,
		_w2547_
	);
	LUT3 #(
		.INIT('hb4)
	) name2243 (
		_w2534_,
		_w2543_,
		_w2547_,
		_w2548_
	);
	LUT4 #(
		.INIT('h707d)
	) name2244 (
		_w1980_,
		_w1931_,
		_w2003_,
		_w1981_,
		_w2549_
	);
	LUT4 #(
		.INIT('hf3bf)
	) name2245 (
		_w1958_,
		_w1980_,
		_w1931_,
		_w2003_,
		_w2550_
	);
	LUT4 #(
		.INIT('hdef6)
	) name2246 (
		_w1958_,
		_w1980_,
		_w1931_,
		_w2003_,
		_w2551_
	);
	LUT4 #(
		.INIT('hd800)
	) name2247 (
		_w1909_,
		_w2550_,
		_w2549_,
		_w2551_,
		_w2552_
	);
	LUT3 #(
		.INIT('h2a)
	) name2248 (
		_w1909_,
		_w1980_,
		_w2018_,
		_w2553_
	);
	LUT3 #(
		.INIT('hb4)
	) name2249 (
		_w1958_,
		_w1980_,
		_w1931_,
		_w2554_
	);
	LUT2 #(
		.INIT('h8)
	) name2250 (
		_w2011_,
		_w2023_,
		_w2555_
	);
	LUT4 #(
		.INIT('h67ef)
	) name2251 (
		_w1980_,
		_w1931_,
		_w2018_,
		_w2020_,
		_w2556_
	);
	LUT4 #(
		.INIT('h0700)
	) name2252 (
		_w2553_,
		_w2554_,
		_w2555_,
		_w2556_,
		_w2557_
	);
	LUT4 #(
		.INIT('h4182)
	) name2253 (
		_w1745_,
		_w1903_,
		_w1907_,
		_w1930_,
		_w2558_
	);
	LUT2 #(
		.INIT('h8)
	) name2254 (
		_w2010_,
		_w2558_,
		_w2559_
	);
	LUT4 #(
		.INIT('h000b)
	) name2255 (
		_w1909_,
		_w2046_,
		_w2053_,
		_w2559_,
		_w2560_
	);
	LUT4 #(
		.INIT('hd800)
	) name2256 (
		_w1882_,
		_w2552_,
		_w2557_,
		_w2560_,
		_w2561_
	);
	LUT4 #(
		.INIT('h0100)
	) name2257 (
		\desIn[16]_pad ,
		\roundSel[4]_pad ,
		\roundSel[5]_pad ,
		_w305_,
		_w2562_
	);
	LUT4 #(
		.INIT('h2800)
	) name2258 (
		\FP_R_reg[27]/P0001 ,
		\roundSel[4]_pad ,
		\roundSel[5]_pad ,
		_w305_,
		_w2563_
	);
	LUT4 #(
		.INIT('h7c55)
	) name2259 (
		\FP_R_reg[59]/NET0131 ,
		\roundSel[4]_pad ,
		\roundSel[5]_pad ,
		_w305_,
		_w2564_
	);
	LUT3 #(
		.INIT('h45)
	) name2260 (
		_w2562_,
		_w2563_,
		_w2564_,
		_w2565_
	);
	LUT2 #(
		.INIT('h9)
	) name2261 (
		_w2561_,
		_w2565_,
		_w2566_
	);
	LUT4 #(
		.INIT('hbfbe)
	) name2262 (
		_w501_,
		_w528_,
		_w570_,
		_w626_,
		_w2567_
	);
	LUT2 #(
		.INIT('h8)
	) name2263 (
		_w528_,
		_w2266_,
		_w2568_
	);
	LUT4 #(
		.INIT('h0032)
	) name2264 (
		_w597_,
		_w2271_,
		_w2567_,
		_w2568_,
		_w2569_
	);
	LUT2 #(
		.INIT('h2)
	) name2265 (
		_w429_,
		_w2569_,
		_w2570_
	);
	LUT3 #(
		.INIT('h08)
	) name2266 (
		_w501_,
		_w571_,
		_w597_,
		_w2571_
	);
	LUT3 #(
		.INIT('h04)
	) name2267 (
		_w632_,
		_w639_,
		_w2571_,
		_w2572_
	);
	LUT4 #(
		.INIT('hbf8f)
	) name2268 (
		_w501_,
		_w528_,
		_w570_,
		_w652_,
		_w2573_
	);
	LUT3 #(
		.INIT('h31)
	) name2269 (
		_w597_,
		_w1392_,
		_w2573_,
		_w2574_
	);
	LUT4 #(
		.INIT('hf5df)
	) name2270 (
		_w501_,
		_w528_,
		_w570_,
		_w626_,
		_w2575_
	);
	LUT4 #(
		.INIT('h0702)
	) name2271 (
		_w597_,
		_w1398_,
		_w1394_,
		_w2575_,
		_w2576_
	);
	LUT4 #(
		.INIT('hea00)
	) name2272 (
		_w429_,
		_w2572_,
		_w2574_,
		_w2576_,
		_w2577_
	);
	LUT4 #(
		.INIT('h0100)
	) name2273 (
		\desIn[62]_pad ,
		\roundSel[4]_pad ,
		\roundSel[5]_pad ,
		_w305_,
		_w2578_
	);
	LUT4 #(
		.INIT('h2800)
	) name2274 (
		\FP_R_reg[8]/P0001 ,
		\roundSel[4]_pad ,
		\roundSel[5]_pad ,
		_w305_,
		_w2579_
	);
	LUT4 #(
		.INIT('h7c55)
	) name2275 (
		\FP_R_reg[40]/NET0131 ,
		\roundSel[4]_pad ,
		\roundSel[5]_pad ,
		_w305_,
		_w2580_
	);
	LUT3 #(
		.INIT('h45)
	) name2276 (
		_w2578_,
		_w2579_,
		_w2580_,
		_w2581_
	);
	LUT3 #(
		.INIT('h4b)
	) name2277 (
		_w2570_,
		_w2577_,
		_w2581_,
		_w2582_
	);
	LUT4 #(
		.INIT('h385f)
	) name2278 (
		_w2081_,
		_w2103_,
		_w2126_,
		_w2148_,
		_w2583_
	);
	LUT3 #(
		.INIT('h80)
	) name2279 (
		_w2081_,
		_w2103_,
		_w2149_,
		_w2584_
	);
	LUT4 #(
		.INIT('h3302)
	) name2280 (
		_w2176_,
		_w2201_,
		_w2583_,
		_w2584_,
		_w2585_
	);
	LUT3 #(
		.INIT('h01)
	) name2281 (
		_w2176_,
		_w2202_,
		_w2205_,
		_w2586_
	);
	LUT3 #(
		.INIT('h20)
	) name2282 (
		_w2081_,
		_w2210_,
		_w2213_,
		_w2587_
	);
	LUT2 #(
		.INIT('h1)
	) name2283 (
		_w2586_,
		_w2587_,
		_w2588_
	);
	LUT4 #(
		.INIT('hcfaf)
	) name2284 (
		_w2081_,
		_w2103_,
		_w2126_,
		_w2148_,
		_w2589_
	);
	LUT3 #(
		.INIT('h08)
	) name2285 (
		_w2202_,
		_w2205_,
		_w2279_,
		_w2590_
	);
	LUT3 #(
		.INIT('h0d)
	) name2286 (
		_w2176_,
		_w2589_,
		_w2590_,
		_w2591_
	);
	LUT3 #(
		.INIT('h2a)
	) name2287 (
		_w2201_,
		_w2588_,
		_w2591_,
		_w2592_
	);
	LUT4 #(
		.INIT('h1428)
	) name2288 (
		_w904_,
		_w2170_,
		_w2174_,
		_w2200_,
		_w2593_
	);
	LUT3 #(
		.INIT('hb0)
	) name2289 (
		_w2206_,
		_w2283_,
		_w2593_,
		_w2594_
	);
	LUT4 #(
		.INIT('h0990)
	) name2290 (
		_w997_,
		_w2125_,
		_w2170_,
		_w2174_,
		_w2595_
	);
	LUT3 #(
		.INIT('h40)
	) name2291 (
		_w2081_,
		_w2204_,
		_w2595_,
		_w2596_
	);
	LUT3 #(
		.INIT('h40)
	) name2292 (
		_w2103_,
		_w2280_,
		_w2279_,
		_w2597_
	);
	LUT3 #(
		.INIT('h01)
	) name2293 (
		_w2215_,
		_w2597_,
		_w2596_,
		_w2598_
	);
	LUT2 #(
		.INIT('h4)
	) name2294 (
		_w2594_,
		_w2598_,
		_w2599_
	);
	LUT4 #(
		.INIT('h0100)
	) name2295 (
		\desIn[58]_pad ,
		\roundSel[4]_pad ,
		\roundSel[5]_pad ,
		_w305_,
		_w2600_
	);
	LUT4 #(
		.INIT('h2800)
	) name2296 (
		\FP_R_reg[24]/P0001 ,
		\roundSel[4]_pad ,
		\roundSel[5]_pad ,
		_w305_,
		_w2601_
	);
	LUT4 #(
		.INIT('h7c55)
	) name2297 (
		\FP_R_reg[56]/NET0131 ,
		\roundSel[4]_pad ,
		\roundSel[5]_pad ,
		_w305_,
		_w2602_
	);
	LUT3 #(
		.INIT('h45)
	) name2298 (
		_w2600_,
		_w2601_,
		_w2602_,
		_w2603_
	);
	LUT4 #(
		.INIT('h10ef)
	) name2299 (
		_w2592_,
		_w2585_,
		_w2599_,
		_w2603_,
		_w2604_
	);
	assign \_al_n0  = 1'b0;
	assign \_al_n1  = 1'b1;
	assign \desOut[0]_pad  = _w661_ ;
	assign \desOut[11]_pad  = _w625_ ;
	assign \desOut[12]_pad  = _w993_ ;
	assign \desOut[13]_pad  = _w998_ ;
	assign \desOut[14]_pad  = _w1197_ ;
	assign \desOut[15]_pad  = _w1203_ ;
	assign \desOut[18]_pad  = _w1387_ ;
	assign \desOut[1]_pad  = _w1256_ ;
	assign \desOut[22]_pad  = _w1409_ ;
	assign \desOut[23]_pad  = _w1414_ ;
	assign \desOut[24]_pad  = _w1440_ ;
	assign \desOut[25]_pad  = _w1445_ ;
	assign \desOut[26]_pad  = _w1470_ ;
	assign \desOut[28]_pad  = _w1648_ ;
	assign \desOut[2]_pad  = _w1818_ ;
	assign \desOut[30]_pad  = _w1842_ ;
	assign \desOut[32]_pad  = _w1860_ ;
	assign \desOut[34]_pad  = _w2038_ ;
	assign \desOut[35]_pad  = _w569_ ;
	assign \desOut[37]_pad  = _w819_ ;
	assign \desOut[38]_pad  = _w2059_ ;
	assign \desOut[39]_pad  = _w1058_ ;
	assign \desOut[3]_pad  = _w500_ ;
	assign \desOut[40]_pad  = _w2228_ ;
	assign \desOut[42]_pad  = _w2255_ ;
	assign \desOut[44]_pad  = _w2278_ ;
	assign \desOut[45]_pad  = _w876_ ;
	assign \desOut[46]_pad  = _w2298_ ;
	assign \desOut[48]_pad  = _w2329_ ;
	assign \desOut[4]_pad  = _w2344_ ;
	assign \desOut[50]_pad  = _w2366_ ;
	assign \desOut[52]_pad  = _w2386_ ;
	assign \desOut[54]_pad  = _w2406_ ;
	assign \desOut[56]_pad  = _w2428_ ;
	assign \desOut[57]_pad  = _w1718_ ;
	assign \desOut[59]_pad  = _w1339_ ;
	assign \desOut[5]_pad  = _w1085_ ;
	assign \desOut[60]_pad  = _w2445_ ;
	assign \desOut[61]_pad  = _w527_ ;
	assign \desOut[63]_pad  = _w1003_ ;
	assign \desOut[6]_pad  = _w2469_ ;
	assign \desOut[8]_pad  = _w2490_ ;
	assign \desOut[9]_pad  = _w1572_ ;
	assign \g13525_dup/_0_  = _w2512_ ;
	assign \g13583_dup/_0_  = _w2528_ ;
	assign \g17813/_3_  = _w1112_ ;
	assign \g17816/_3_  = _w1957_ ;
	assign \g17819/_3_  = _w955_ ;
	assign \g17822/_3_  = _w1208_ ;
	assign \g17836/_3_  = _w1500_ ;
	assign \g17871/_3_  = _w1140_ ;
	assign \g17878/_1_  = _w311_ ;
	assign \g17881/_3_  = _w2175_ ;
	assign \g17966/_2_  = _w1908_ ;
	assign \g17969/_3_  = _w1330_ ;
	assign \g17996/_2_  = _w905_ ;
	assign \g19574_dup/_3_  = _w2548_ ;
	assign \g19619_dup/_3_  = _w2566_ ;
	assign \g19756_dup/_3_  = _w2582_ ;
	assign \g20263/_3_  = _w1600_ ;
	assign \g20541/_2_  = _w1746_ ;
	assign \g20691/_1_  = _w596_ ;
	assign \g20740_dup/_3_  = _w2604_ ;
	assign \g67/_2_  = _w1052_ ;
endmodule;