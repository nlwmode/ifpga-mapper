module top( CLR_pad , \v0_pad  , \v10_reg/NET0131  , \v11_reg/NET0131  , \v12_reg/NET0131  , \v1_pad  , \v2_pad  , \v3_pad  , \v4_pad  , \v5_pad  , \v6_pad  , \v7_reg/NET0131  , \v8_reg/NET0131  , \v9_reg/NET0131  , \_al_n0  , \_al_n1  , \g1757/_0_  , \g1763/_1_  , \g1787/_3_  , \g1800/_3_  , \g1821/_2_  , \g1940/_1_  , \g25/_0_  , \g2783/_3_  , \g2823/_0_  , \g38/_1_  , \g40/_1_  , \v13_D_11_pad  , \v13_D_12_pad  , \v13_D_13_pad  , \v13_D_14_pad  , \v13_D_16_pad  , \v13_D_18_pad  , \v13_D_19_pad  , \v13_D_21_pad  , \v13_D_22_pad  , \v13_D_23_pad  , \v13_D_24_pad  , \v13_D_7_pad  , \v13_D_8_pad  , \v13_D_9_pad  );
  input CLR_pad ;
  input \v0_pad  ;
  input \v10_reg/NET0131  ;
  input \v11_reg/NET0131  ;
  input \v12_reg/NET0131  ;
  input \v1_pad  ;
  input \v2_pad  ;
  input \v3_pad  ;
  input \v4_pad  ;
  input \v5_pad  ;
  input \v6_pad  ;
  input \v7_reg/NET0131  ;
  input \v8_reg/NET0131  ;
  input \v9_reg/NET0131  ;
  output \_al_n0  ;
  output \_al_n1  ;
  output \g1757/_0_  ;
  output \g1763/_1_  ;
  output \g1787/_3_  ;
  output \g1800/_3_  ;
  output \g1821/_2_  ;
  output \g1940/_1_  ;
  output \g25/_0_  ;
  output \g2783/_3_  ;
  output \g2823/_0_  ;
  output \g38/_1_  ;
  output \g40/_1_  ;
  output \v13_D_11_pad  ;
  output \v13_D_12_pad  ;
  output \v13_D_13_pad  ;
  output \v13_D_14_pad  ;
  output \v13_D_16_pad  ;
  output \v13_D_18_pad  ;
  output \v13_D_19_pad  ;
  output \v13_D_21_pad  ;
  output \v13_D_22_pad  ;
  output \v13_D_23_pad  ;
  output \v13_D_24_pad  ;
  output \v13_D_7_pad  ;
  output \v13_D_8_pad  ;
  output \v13_D_9_pad  ;
  wire n15 , n16 , n17 , n18 , n19 , n20 , n21 , n22 , n23 , n24 , n25 , n26 , n27 , n28 , n29 , n30 , n31 , n32 , n33 , n34 , n35 , n36 , n37 , n38 , n39 , n40 , n41 , n42 , n43 , n44 , n45 , n46 , n47 , n48 , n49 , n50 , n51 , n52 , n53 , n54 , n55 , n56 , n57 , n58 , n59 , n60 , n61 , n62 , n63 , n64 , n65 , n66 , n67 , n68 , n69 , n70 , n71 , n72 , n73 , n74 , n75 , n76 , n77 , n78 , n79 , n80 , n81 , n82 , n83 , n84 , n85 , n86 , n87 , n88 , n89 , n90 , n91 , n92 , n93 , n94 , n95 , n96 , n97 , n98 , n99 , n100 , n101 , n102 , n103 , n104 , n105 , n106 , n107 , n108 , n109 , n110 , n111 , n112 , n113 , n114 , n115 , n116 , n117 , n118 , n119 , n120 , n121 , n122 , n123 , n124 , n125 , n126 , n127 , n128 , n129 , n130 , n131 , n132 , n133 , n134 , n135 , n136 , n137 , n138 , n139 , n140 , n141 , n142 , n143 , n144 , n145 , n146 , n147 , n148 , n149 , n150 , n151 , n152 , n153 , n154 , n155 , n156 , n157 , n158 , n159 , n160 , n161 , n162 , n163 , n164 , n165 , n166 , n167 , n168 , n169 , n170 , n171 , n172 , n173 , n174 , n175 , n176 , n177 , n178 , n179 , n180 , n181 , n182 , n183 , n184 , n185 , n186 , n187 , n188 , n189 , n190 , n191 , n192 , n193 , n194 , n195 , n196 , n197 , n198 , n199 , n200 , n201 , n202 , n203 , n204 , n205 , n206 , n207 , n208 , n209 , n210 , n211 , n212 , n213 , n214 , n215 , n216 , n217 , n218 , n219 , n220 , n221 , n222 , n223 , n224 , n225 , n226 , n227 , n228 , n229 , n230 , n231 , n232 , n233 , n234 , n235 , n236 , n237 , n238 , n239 , n240 , n241 , n242 , n243 , n244 , n245 , n246 , n247 , n248 , n249 , n250 , n251 , n252 , n253 , n254 , n255 , n256 , n257 , n258 , n259 , n260 , n261 , n262 , n263 , n264 , n265 , n266 , n267 , n268 , n269 , n270 , n271 , n272 , n273 , n274 , n275 , n276 , n277 , n278 , n279 , n280 , n281 , n282 , n283 , n284 , n285 , n286 , n287 , n288 , n289 , n290 , n291 , n292 , n293 , n294 , n295 , n296 , n297 , n298 , n299 , n300 , n301 , n302 , n303 , n304 , n305 , n306 , n307 , n308 , n309 , n310 , n311 , n312 , n313 , n314 , n315 , n316 , n317 , n318 , n319 , n320 , n321 , n322 , n323 , n324 , n325 , n326 , n327 , n328 , n329 , n330 , n331 , n332 , n333 , n334 , n335 , n336 , n337 , n338 , n339 , n340 , n341 , n342 , n343 , n344 , n345 , n346 , n347 , n348 , n349 , n350 , n351 , n352 , n353 , n354 , n355 , n356 , n357 , n358 , n359 , n360 , n361 , n362 , n363 , n364 , n365 , n366 , n367 , n368 , n369 , n370 , n371 , n372 , n373 , n374 , n375 , n376 , n377 , n378 , n379 , n380 , n381 , n382 , n383 , n384 , n385 , n386 , n387 , n388 , n389 , n390 , n391 , n392 , n393 , n394 , n395 , n396 , n397 , n398 , n399 , n400 , n401 , n402 , n403 , n404 , n405 , n406 , n407 , n408 , n409 , n410 , n411 , n412 , n413 , n414 , n415 , n416 , n417 , n418 , n419 , n420 , n421 , n422 , n423 , n424 , n425 , n426 , n427 , n428 , n429 , n430 , n431 , n432 , n433 , n434 , n435 , n436 , n437 , n438 , n439 , n440 , n441 , n442 , n443 , n444 , n445 , n446 , n447 , n448 , n449 , n450 , n451 , n452 , n453 , n454 , n455 , n456 , n457 , n458 , n459 , n460 , n461 , n462 , n463 , n464 , n465 , n466 , n467 , n468 , n469 , n470 , n471 , n472 , n473 , n474 , n475 , n476 , n477 , n478 , n479 , n480 , n481 , n482 , n483 , n484 , n485 , n486 , n487 , n488 , n489 , n490 , n491 , n492 , n493 , n494 , n495 , n496 , n497 , n498 , n499 , n500 , n501 , n502 , n503 , n504 , n505 , n506 , n507 , n508 , n509 , n510 , n511 , n512 , n513 , n514 , n515 , n516 , n517 , n518 , n519 , n520 , n521 , n522 , n523 , n524 , n525 , n526 , n527 , n528 , n529 , n530 , n531 , n532 , n533 , n534 , n535 , n536 , n537 , n538 , n539 , n540 , n541 , n542 , n543 , n544 , n545 , n546 , n547 , n548 , n549 , n550 , n551 , n552 , n553 , n554 , n555 , n556 , n557 , n558 , n559 , n560 , n561 , n562 , n563 , n564 , n565 , n566 , n567 , n568 , n569 , n570 , n571 , n572 , n573 , n574 , n575 , n576 , n577 , n578 , n579 ;
  assign n25 = ~\v10_reg/NET0131  & \v11_reg/NET0131  ;
  assign n26 = \v10_reg/NET0131  & ~\v11_reg/NET0131  ;
  assign n27 = ~n25 & ~n26 ;
  assign n28 = ~\v10_reg/NET0131  & ~\v3_pad  ;
  assign n29 = ~\v6_pad  & n28 ;
  assign n30 = n27 & ~n29 ;
  assign n31 = \v12_reg/NET0131  & ~n30 ;
  assign n15 = \v10_reg/NET0131  & ~\v12_reg/NET0131  ;
  assign n16 = ~\v11_reg/NET0131  & n15 ;
  assign n17 = \v9_reg/NET0131  & ~n16 ;
  assign n18 = \v10_reg/NET0131  & \v11_reg/NET0131  ;
  assign n19 = ~\v0_pad  & n18 ;
  assign n20 = ~\v10_reg/NET0131  & ~\v11_reg/NET0131  ;
  assign n21 = ~n19 & ~n20 ;
  assign n22 = \v4_pad  & \v5_pad  ;
  assign n23 = ~\v12_reg/NET0131  & n22 ;
  assign n24 = ~n21 & n23 ;
  assign n32 = ~n17 & ~n24 ;
  assign n33 = ~n31 & n32 ;
  assign n34 = ~\v8_reg/NET0131  & ~n33 ;
  assign n39 = \v11_reg/NET0131  & \v12_reg/NET0131  ;
  assign n40 = ~\v10_reg/NET0131  & ~\v1_pad  ;
  assign n41 = n39 & n40 ;
  assign n35 = \v12_reg/NET0131  & ~\v3_pad  ;
  assign n36 = \v10_reg/NET0131  & ~\v8_reg/NET0131  ;
  assign n37 = n35 & n36 ;
  assign n38 = ~\v8_reg/NET0131  & \v9_reg/NET0131  ;
  assign n42 = ~n37 & ~n38 ;
  assign n43 = ~n41 & n42 ;
  assign n44 = \v2_pad  & ~n43 ;
  assign n45 = \v9_reg/NET0131  & n39 ;
  assign n46 = ~\v10_reg/NET0131  & \v8_reg/NET0131  ;
  assign n47 = ~\v12_reg/NET0131  & ~\v9_reg/NET0131  ;
  assign n48 = n46 & n47 ;
  assign n49 = ~n45 & ~n48 ;
  assign n50 = ~n44 & n49 ;
  assign n51 = ~n34 & n50 ;
  assign n52 = ~\v7_reg/NET0131  & ~n51 ;
  assign n75 = \v11_reg/NET0131  & ~n46 ;
  assign n76 = ~\v12_reg/NET0131  & ~n36 ;
  assign n77 = n75 & n76 ;
  assign n71 = ~\v12_reg/NET0131  & \v9_reg/NET0131  ;
  assign n72 = n18 & n71 ;
  assign n54 = \v12_reg/NET0131  & ~\v9_reg/NET0131  ;
  assign n73 = \v11_reg/NET0131  & ~n54 ;
  assign n74 = n46 & ~n73 ;
  assign n78 = ~n72 & ~n74 ;
  assign n79 = ~n77 & n78 ;
  assign n80 = \v7_reg/NET0131  & ~n79 ;
  assign n64 = \v12_reg/NET0131  & \v1_pad  ;
  assign n65 = ~\v10_reg/NET0131  & n64 ;
  assign n66 = \v8_reg/NET0131  & n23 ;
  assign n67 = ~n65 & ~n66 ;
  assign n68 = \v11_reg/NET0131  & ~\v2_pad  ;
  assign n69 = ~\v7_reg/NET0131  & n68 ;
  assign n70 = ~n67 & n69 ;
  assign n53 = ~\v2_pad  & \v8_reg/NET0131  ;
  assign n55 = \v7_reg/NET0131  & n54 ;
  assign n56 = \v11_reg/NET0131  & n15 ;
  assign n57 = ~n55 & ~n56 ;
  assign n58 = n53 & ~n57 ;
  assign n59 = ~\v10_reg/NET0131  & ~\v12_reg/NET0131  ;
  assign n60 = \v3_pad  & n59 ;
  assign n61 = ~n54 & ~n60 ;
  assign n62 = ~\v11_reg/NET0131  & \v8_reg/NET0131  ;
  assign n63 = ~n61 & n62 ;
  assign n81 = ~n58 & ~n63 ;
  assign n82 = ~n70 & n81 ;
  assign n83 = ~n80 & n82 ;
  assign n84 = ~n52 & n83 ;
  assign n85 = CLR_pad & ~n84 ;
  assign n118 = ~\v8_reg/NET0131  & ~\v9_reg/NET0131  ;
  assign n119 = \v12_reg/NET0131  & n25 ;
  assign n120 = ~\v0_pad  & \v11_reg/NET0131  ;
  assign n121 = n15 & ~n120 ;
  assign n122 = ~n119 & ~n121 ;
  assign n123 = n118 & ~n122 ;
  assign n112 = ~\v10_reg/NET0131  & ~\v9_reg/NET0131  ;
  assign n113 = n23 & n112 ;
  assign n114 = ~\v11_reg/NET0131  & n113 ;
  assign n89 = ~\v11_reg/NET0131  & ~\v8_reg/NET0131  ;
  assign n90 = n71 & n89 ;
  assign n115 = n39 & n53 ;
  assign n116 = ~n90 & ~n115 ;
  assign n117 = n40 & ~n116 ;
  assign n129 = ~n114 & ~n117 ;
  assign n130 = ~n123 & n129 ;
  assign n86 = ~\v9_reg/NET0131  & ~n64 ;
  assign n87 = \v11_reg/NET0131  & n46 ;
  assign n88 = ~n86 & n87 ;
  assign n91 = ~\v10_reg/NET0131  & n90 ;
  assign n92 = ~n88 & ~n91 ;
  assign n93 = \v2_pad  & ~n92 ;
  assign n109 = \v8_reg/NET0131  & \v9_reg/NET0131  ;
  assign n110 = \v12_reg/NET0131  & ~n18 ;
  assign n111 = n109 & n110 ;
  assign n103 = ~\v11_reg/NET0131  & ~\v6_pad  ;
  assign n104 = ~\v10_reg/NET0131  & ~\v8_reg/NET0131  ;
  assign n105 = n71 & n104 ;
  assign n106 = n103 & n105 ;
  assign n107 = \v9_reg/NET0131  & ~n22 ;
  assign n108 = n87 & n107 ;
  assign n126 = ~n106 & ~n108 ;
  assign n127 = ~n111 & n126 ;
  assign n94 = \v2_pad  & n26 ;
  assign n95 = ~n22 & n36 ;
  assign n96 = ~n94 & ~n95 ;
  assign n97 = n47 & ~n96 ;
  assign n100 = ~\v11_reg/NET0131  & \v3_pad  ;
  assign n101 = ~\v12_reg/NET0131  & n46 ;
  assign n102 = n100 & n101 ;
  assign n98 = \v12_reg/NET0131  & \v9_reg/NET0131  ;
  assign n99 = n26 & n98 ;
  assign n124 = ~\v7_reg/NET0131  & ~n99 ;
  assign n125 = ~n102 & n124 ;
  assign n128 = ~n97 & n125 ;
  assign n131 = n127 & n128 ;
  assign n132 = ~n93 & n131 ;
  assign n133 = n130 & n132 ;
  assign n139 = ~\v12_reg/NET0131  & ~n20 ;
  assign n140 = \v9_reg/NET0131  & ~n139 ;
  assign n137 = \v12_reg/NET0131  & ~n68 ;
  assign n138 = n27 & n137 ;
  assign n141 = \v8_reg/NET0131  & ~n138 ;
  assign n142 = ~n140 & n141 ;
  assign n134 = \v11_reg/NET0131  & ~\v12_reg/NET0131  ;
  assign n135 = \v10_reg/NET0131  & ~\v9_reg/NET0131  ;
  assign n136 = n134 & ~n135 ;
  assign n143 = \v7_reg/NET0131  & ~n136 ;
  assign n144 = ~n142 & n143 ;
  assign n145 = ~n133 & ~n144 ;
  assign n146 = \v11_reg/NET0131  & \v3_pad  ;
  assign n147 = n48 & ~n146 ;
  assign n148 = ~\v6_pad  & n104 ;
  assign n149 = ~\v7_reg/NET0131  & ~\v9_reg/NET0131  ;
  assign n150 = n35 & n149 ;
  assign n151 = n148 & n150 ;
  assign n152 = ~n147 & ~n151 ;
  assign n153 = ~n145 & n152 ;
  assign n154 = CLR_pad & ~n153 ;
  assign n155 = ~\v7_reg/NET0131  & ~\v8_reg/NET0131  ;
  assign n156 = n114 & n155 ;
  assign n157 = \v11_reg/NET0131  & \v9_reg/NET0131  ;
  assign n158 = \v0_pad  & \v11_reg/NET0131  ;
  assign n159 = n149 & ~n158 ;
  assign n160 = ~n157 & ~n159 ;
  assign n161 = \v10_reg/NET0131  & ~n160 ;
  assign n162 = \v8_reg/NET0131  & ~n112 ;
  assign n163 = \v11_reg/NET0131  & n162 ;
  assign n164 = ~n161 & ~n163 ;
  assign n165 = ~\v12_reg/NET0131  & ~n164 ;
  assign n166 = ~\v8_reg/NET0131  & ~n25 ;
  assign n167 = ~\v12_reg/NET0131  & ~n166 ;
  assign n168 = \v11_reg/NET0131  & n135 ;
  assign n169 = \v8_reg/NET0131  & n168 ;
  assign n170 = ~n167 & ~n169 ;
  assign n171 = \v7_reg/NET0131  & ~n170 ;
  assign n172 = ~n165 & ~n171 ;
  assign n173 = \v2_pad  & ~n172 ;
  assign n174 = ~n156 & ~n173 ;
  assign n175 = ~\v2_pad  & \v9_reg/NET0131  ;
  assign n176 = \v11_reg/NET0131  & n175 ;
  assign n177 = ~n94 & ~n176 ;
  assign n178 = ~\v12_reg/NET0131  & ~n177 ;
  assign n179 = \v8_reg/NET0131  & ~n178 ;
  assign n180 = \v11_reg/NET0131  & ~n104 ;
  assign n181 = ~\v4_pad  & \v5_pad  ;
  assign n182 = ~\v10_reg/NET0131  & ~n181 ;
  assign n183 = ~\v9_reg/NET0131  & ~n182 ;
  assign n184 = ~n180 & ~n183 ;
  assign n185 = ~\v12_reg/NET0131  & ~n184 ;
  assign n186 = \v11_reg/NET0131  & n112 ;
  assign n187 = ~n185 & ~n186 ;
  assign n188 = ~n179 & ~n187 ;
  assign n189 = ~\v7_reg/NET0131  & ~n188 ;
  assign n194 = \v7_reg/NET0131  & n112 ;
  assign n195 = ~\v12_reg/NET0131  & ~n194 ;
  assign n190 = ~\v10_reg/NET0131  & n54 ;
  assign n191 = ~\v11_reg/NET0131  & n190 ;
  assign n192 = \v9_reg/NET0131  & ~n20 ;
  assign n193 = \v8_reg/NET0131  & ~n192 ;
  assign n196 = ~n191 & n193 ;
  assign n197 = ~n195 & n196 ;
  assign n198 = ~n189 & ~n197 ;
  assign n199 = ~n21 & n118 ;
  assign n200 = \v11_reg/NET0131  & \v8_reg/NET0131  ;
  assign n201 = n175 & n200 ;
  assign n202 = ~n199 & ~n201 ;
  assign n203 = ~\v12_reg/NET0131  & ~\v7_reg/NET0131  ;
  assign n204 = \v4_pad  & ~\v5_pad  ;
  assign n205 = n203 & n204 ;
  assign n206 = ~n202 & n205 ;
  assign n207 = ~\v1_pad  & \v6_pad  ;
  assign n208 = \v8_reg/NET0131  & ~n207 ;
  assign n209 = \v10_reg/NET0131  & ~\v7_reg/NET0131  ;
  assign n210 = n98 & n146 ;
  assign n211 = n209 & n210 ;
  assign n212 = n208 & n211 ;
  assign n213 = \v10_reg/NET0131  & ~\v2_pad  ;
  assign n214 = ~n22 & n213 ;
  assign n215 = n134 & ~n214 ;
  assign n216 = \v9_reg/NET0131  & ~n215 ;
  assign n217 = n162 & ~n216 ;
  assign n232 = \v6_pad  & n20 ;
  assign n233 = \v12_reg/NET0131  & n232 ;
  assign n234 = n118 & n233 ;
  assign n236 = n200 & n207 ;
  assign n218 = \v12_reg/NET0131  & \v3_pad  ;
  assign n235 = ~\v0_pad  & \v10_reg/NET0131  ;
  assign n237 = n218 & n235 ;
  assign n238 = n236 & n237 ;
  assign n239 = ~n234 & ~n238 ;
  assign n240 = ~n217 & n239 ;
  assign n219 = n20 & n118 ;
  assign n220 = \v10_reg/NET0131  & n158 ;
  assign n221 = n208 & n220 ;
  assign n222 = ~n219 & ~n221 ;
  assign n223 = n218 & ~n222 ;
  assign n224 = ~\v11_reg/NET0131  & ~n47 ;
  assign n225 = \v11_reg/NET0131  & ~n38 ;
  assign n226 = ~n224 & ~n225 ;
  assign n227 = ~\v9_reg/NET0131  & n22 ;
  assign n228 = ~\v0_pad  & ~\v12_reg/NET0131  ;
  assign n229 = n227 & n228 ;
  assign n230 = ~n226 & ~n229 ;
  assign n231 = \v10_reg/NET0131  & ~n230 ;
  assign n241 = ~n223 & ~n231 ;
  assign n242 = n240 & n241 ;
  assign n243 = ~\v7_reg/NET0131  & ~n242 ;
  assign n246 = ~\v12_reg/NET0131  & ~\v8_reg/NET0131  ;
  assign n247 = ~n224 & ~n246 ;
  assign n248 = ~\v10_reg/NET0131  & ~n89 ;
  assign n249 = ~n247 & n248 ;
  assign n250 = ~n72 & ~n249 ;
  assign n251 = \v7_reg/NET0131  & ~n250 ;
  assign n244 = \v8_reg/NET0131  & n135 ;
  assign n245 = ~n137 & n244 ;
  assign n252 = ~\v12_reg/NET0131  & ~\v2_pad  ;
  assign n253 = \v1_pad  & ~\v7_reg/NET0131  ;
  assign n254 = n38 & n253 ;
  assign n255 = n252 & n254 ;
  assign n256 = n232 & n255 ;
  assign n257 = ~n245 & ~n256 ;
  assign n258 = ~n251 & n257 ;
  assign n259 = ~n243 & n258 ;
  assign n260 = CLR_pad & ~n259 ;
  assign n261 = ~\v8_reg/NET0131  & n158 ;
  assign n262 = n26 & ~n53 ;
  assign n263 = ~n261 & ~n262 ;
  assign n264 = n149 & ~n263 ;
  assign n265 = \v11_reg/NET0131  & ~n135 ;
  assign n266 = ~\v10_reg/NET0131  & \v9_reg/NET0131  ;
  assign n267 = ~\v8_reg/NET0131  & ~n266 ;
  assign n268 = n265 & n267 ;
  assign n270 = ~n149 & ~n200 ;
  assign n269 = \v8_reg/NET0131  & ~\v9_reg/NET0131  ;
  assign n271 = n22 & ~n269 ;
  assign n272 = ~n270 & n271 ;
  assign n273 = ~n268 & ~n272 ;
  assign n274 = ~n264 & n273 ;
  assign n275 = ~\v12_reg/NET0131  & ~n274 ;
  assign n276 = \v11_reg/NET0131  & ~n252 ;
  assign n277 = ~\v7_reg/NET0131  & ~n276 ;
  assign n278 = n26 & ~n47 ;
  assign n279 = \v8_reg/NET0131  & ~n98 ;
  assign n280 = ~n186 & n279 ;
  assign n281 = ~n278 & n280 ;
  assign n282 = ~n277 & n281 ;
  assign n283 = ~n275 & ~n282 ;
  assign n290 = ~\v12_reg/NET0131  & \v1_pad  ;
  assign n291 = n18 & ~n207 ;
  assign n292 = ~n290 & ~n291 ;
  assign n293 = \v3_pad  & ~n292 ;
  assign n295 = \v12_reg/NET0131  & ~\v8_reg/NET0131  ;
  assign n296 = n26 & n295 ;
  assign n294 = ~\v12_reg/NET0131  & ~n89 ;
  assign n297 = \v9_reg/NET0131  & ~n294 ;
  assign n298 = ~n296 & n297 ;
  assign n299 = ~n293 & n298 ;
  assign n286 = n26 & n71 ;
  assign n284 = n71 & n103 ;
  assign n285 = ~n15 & n157 ;
  assign n287 = ~n284 & ~n285 ;
  assign n288 = ~n286 & n287 ;
  assign n289 = ~\v8_reg/NET0131  & ~n288 ;
  assign n300 = n118 & n235 ;
  assign n301 = n22 & n134 ;
  assign n302 = n300 & n301 ;
  assign n303 = ~n289 & ~n302 ;
  assign n304 = ~n299 & n303 ;
  assign n305 = ~\v7_reg/NET0131  & ~n304 ;
  assign n306 = n22 & n200 ;
  assign n307 = ~n89 & ~n306 ;
  assign n308 = ~\v7_reg/NET0131  & n71 ;
  assign n309 = ~n307 & n308 ;
  assign n310 = \v7_reg/NET0131  & \v8_reg/NET0131  ;
  assign n311 = n54 & n310 ;
  assign n312 = ~n309 & ~n311 ;
  assign n313 = ~\v2_pad  & ~n312 ;
  assign n314 = \v7_reg/NET0131  & ~n18 ;
  assign n315 = ~n47 & n314 ;
  assign n316 = n193 & n315 ;
  assign n317 = ~n313 & ~n316 ;
  assign n318 = ~n305 & n317 ;
  assign n319 = CLR_pad & ~n318 ;
  assign n326 = ~\v12_reg/NET0131  & ~n112 ;
  assign n327 = ~\v2_pad  & ~n107 ;
  assign n328 = n326 & n327 ;
  assign n323 = ~\v3_pad  & ~\v9_reg/NET0131  ;
  assign n324 = n134 & ~n323 ;
  assign n325 = ~\v10_reg/NET0131  & ~n324 ;
  assign n320 = \v0_pad  & n207 ;
  assign n321 = \v3_pad  & n98 ;
  assign n322 = ~n320 & n321 ;
  assign n329 = ~n224 & ~n322 ;
  assign n330 = ~n325 & n329 ;
  assign n331 = ~n328 & n330 ;
  assign n332 = \v8_reg/NET0131  & ~n331 ;
  assign n337 = ~\v1_pad  & n266 ;
  assign n338 = ~n168 & ~n337 ;
  assign n339 = n246 & ~n338 ;
  assign n334 = ~\v11_reg/NET0131  & n54 ;
  assign n335 = ~n105 & ~n334 ;
  assign n336 = ~\v6_pad  & ~n335 ;
  assign n333 = ~\v10_reg/NET0131  & n45 ;
  assign n340 = ~n278 & ~n333 ;
  assign n341 = ~n336 & n340 ;
  assign n342 = ~n339 & n341 ;
  assign n343 = ~n332 & n342 ;
  assign n344 = ~\v7_reg/NET0131  & ~n343 ;
  assign n347 = ~\v8_reg/NET0131  & ~n71 ;
  assign n345 = ~\v10_reg/NET0131  & ~n200 ;
  assign n346 = ~\v11_reg/NET0131  & ~\v12_reg/NET0131  ;
  assign n348 = n345 & ~n346 ;
  assign n349 = ~n347 & n348 ;
  assign n354 = ~\v12_reg/NET0131  & \v2_pad  ;
  assign n355 = ~\v7_reg/NET0131  & n266 ;
  assign n356 = n354 & n355 ;
  assign n361 = ~n349 & ~n356 ;
  assign n350 = \v10_reg/NET0131  & \v8_reg/NET0131  ;
  assign n351 = \v11_reg/NET0131  & \v2_pad  ;
  assign n352 = n55 & n351 ;
  assign n353 = n350 & n352 ;
  assign n357 = ~\v11_reg/NET0131  & ~n244 ;
  assign n358 = ~\v12_reg/NET0131  & \v7_reg/NET0131  ;
  assign n359 = ~n180 & n358 ;
  assign n360 = ~n357 & n359 ;
  assign n362 = ~n353 & ~n360 ;
  assign n363 = n361 & n362 ;
  assign n364 = ~n344 & n363 ;
  assign n365 = CLR_pad & ~n364 ;
  assign n380 = \v11_reg/NET0131  & n322 ;
  assign n381 = ~n22 & n59 ;
  assign n382 = ~n119 & ~n284 ;
  assign n383 = ~n381 & n382 ;
  assign n384 = ~n380 & n383 ;
  assign n385 = \v8_reg/NET0131  & ~n384 ;
  assign n377 = ~n168 & ~n266 ;
  assign n378 = ~n232 & n377 ;
  assign n379 = n295 & ~n378 ;
  assign n366 = ~n71 & ~n104 ;
  assign n367 = ~\v3_pad  & ~n246 ;
  assign n368 = ~n366 & n367 ;
  assign n369 = ~n113 & ~n368 ;
  assign n370 = ~\v11_reg/NET0131  & ~n369 ;
  assign n371 = ~\v11_reg/NET0131  & ~n354 ;
  assign n372 = ~n59 & ~n371 ;
  assign n373 = n269 & ~n372 ;
  assign n374 = \v10_reg/NET0131  & ~n38 ;
  assign n375 = ~n104 & n354 ;
  assign n376 = ~n374 & n375 ;
  assign n386 = ~n373 & ~n376 ;
  assign n387 = ~n370 & n386 ;
  assign n388 = ~n379 & n387 ;
  assign n389 = ~n385 & n388 ;
  assign n390 = ~\v7_reg/NET0131  & ~n389 ;
  assign n391 = \v10_reg/NET0131  & ~n54 ;
  assign n392 = n62 & ~n190 ;
  assign n393 = ~n391 & n392 ;
  assign n394 = ~\v11_reg/NET0131  & ~n46 ;
  assign n395 = \v9_reg/NET0131  & n358 ;
  assign n396 = ~n394 & n395 ;
  assign n397 = ~n393 & ~n396 ;
  assign n398 = ~n390 & n397 ;
  assign n399 = CLR_pad & ~n398 ;
  assign n402 = ~\v9_reg/NET0131  & ~n26 ;
  assign n403 = ~n158 & n402 ;
  assign n404 = ~\v8_reg/NET0131  & ~n403 ;
  assign n405 = \v8_reg/NET0131  & ~n68 ;
  assign n406 = \v6_pad  & n100 ;
  assign n407 = n405 & ~n406 ;
  assign n401 = n22 & ~n62 ;
  assign n408 = ~\v12_reg/NET0131  & ~n401 ;
  assign n409 = ~n407 & n408 ;
  assign n410 = ~n404 & n409 ;
  assign n411 = ~\v7_reg/NET0131  & ~n410 ;
  assign n400 = n104 & n134 ;
  assign n412 = ~n193 & ~n400 ;
  assign n413 = ~n411 & n412 ;
  assign n415 = ~\v10_reg/NET0131  & n22 ;
  assign n416 = ~\v12_reg/NET0131  & ~n158 ;
  assign n417 = ~n415 & n416 ;
  assign n414 = \v12_reg/NET0131  & ~n26 ;
  assign n418 = ~\v9_reg/NET0131  & ~n414 ;
  assign n419 = ~n417 & n418 ;
  assign n420 = ~n72 & ~n419 ;
  assign n421 = ~\v7_reg/NET0131  & ~n420 ;
  assign n422 = ~\v12_reg/NET0131  & n186 ;
  assign n423 = ~n421 & ~n422 ;
  assign n424 = ~\v8_reg/NET0131  & ~n423 ;
  assign n425 = ~n98 & ~n112 ;
  assign n426 = n276 & n425 ;
  assign n427 = ~n358 & ~n426 ;
  assign n428 = \v8_reg/NET0131  & ~n427 ;
  assign n429 = ~n424 & ~n428 ;
  assign n430 = \v11_reg/NET0131  & ~n235 ;
  assign n431 = ~\v9_reg/NET0131  & ~n430 ;
  assign n432 = ~\v8_reg/NET0131  & n431 ;
  assign n433 = ~n201 & ~n432 ;
  assign n434 = n22 & ~n433 ;
  assign n435 = n162 & n351 ;
  assign n436 = ~n434 & ~n435 ;
  assign n437 = ~\v12_reg/NET0131  & ~n436 ;
  assign n438 = ~n15 & ~n295 ;
  assign n439 = ~\v9_reg/NET0131  & ~n27 ;
  assign n440 = ~n438 & n439 ;
  assign n441 = ~n437 & ~n440 ;
  assign n442 = ~\v7_reg/NET0131  & ~n441 ;
  assign n443 = ~n39 & n112 ;
  assign n444 = ~n286 & ~n443 ;
  assign n445 = \v8_reg/NET0131  & ~n444 ;
  assign n446 = ~n400 & ~n445 ;
  assign n447 = \v7_reg/NET0131  & ~n446 ;
  assign n448 = ~n200 & ~n203 ;
  assign n449 = ~\v9_reg/NET0131  & ~n448 ;
  assign n450 = ~n290 & ~n449 ;
  assign n451 = ~n157 & n290 ;
  assign n452 = \v10_reg/NET0131  & ~n451 ;
  assign n453 = ~n450 & n452 ;
  assign n454 = ~n447 & ~n453 ;
  assign n455 = ~n442 & n454 ;
  assign n458 = ~\v8_reg/NET0131  & ~n431 ;
  assign n460 = ~\v12_reg/NET0131  & ~n22 ;
  assign n459 = ~\v4_pad  & ~\v5_pad  ;
  assign n461 = ~n26 & ~n459 ;
  assign n462 = n460 & n461 ;
  assign n463 = ~n405 & n462 ;
  assign n464 = ~n458 & n463 ;
  assign n465 = ~\v7_reg/NET0131  & ~n464 ;
  assign n456 = ~\v8_reg/NET0131  & ~n265 ;
  assign n457 = n358 & ~n456 ;
  assign n466 = ~n193 & ~n457 ;
  assign n467 = ~n465 & n466 ;
  assign n468 = n308 & n406 ;
  assign n469 = ~n352 & ~n468 ;
  assign n470 = n350 & ~n469 ;
  assign n471 = n22 & n219 ;
  assign n472 = \v8_reg/NET0131  & n175 ;
  assign n473 = ~n300 & ~n472 ;
  assign n474 = \v11_reg/NET0131  & ~n459 ;
  assign n475 = ~n473 & n474 ;
  assign n476 = ~n471 & ~n475 ;
  assign n477 = n203 & ~n476 ;
  assign n478 = n54 & n148 ;
  assign n479 = \v6_pad  & n15 ;
  assign n480 = n109 & n479 ;
  assign n481 = ~n478 & ~n480 ;
  assign n482 = ~\v7_reg/NET0131  & n100 ;
  assign n483 = ~n481 & n482 ;
  assign n484 = ~n353 & ~n483 ;
  assign n485 = n89 & n227 ;
  assign n486 = \v2_pad  & n109 ;
  assign n487 = ~n485 & ~n486 ;
  assign n488 = ~\v10_reg/NET0131  & n203 ;
  assign n489 = ~n487 & n488 ;
  assign n490 = n286 & n310 ;
  assign n491 = n62 & n252 ;
  assign n492 = \v12_reg/NET0131  & n38 ;
  assign n493 = ~n491 & ~n492 ;
  assign n494 = ~\v10_reg/NET0131  & ~\v7_reg/NET0131  ;
  assign n495 = ~n493 & n494 ;
  assign n496 = ~n490 & ~n495 ;
  assign n497 = \v0_pad  & n56 ;
  assign n498 = ~n233 & ~n497 ;
  assign n499 = ~\v9_reg/NET0131  & ~n498 ;
  assign n500 = \v10_reg/NET0131  & n45 ;
  assign n501 = ~n499 & ~n500 ;
  assign n502 = n155 & ~n501 ;
  assign n511 = ~\v10_reg/NET0131  & n109 ;
  assign n510 = \v10_reg/NET0131  & ~n109 ;
  assign n512 = n358 & ~n510 ;
  assign n513 = ~n511 & n512 ;
  assign n504 = ~\v12_reg/NET0131  & ~\v5_pad  ;
  assign n515 = \v9_reg/NET0131  & n504 ;
  assign n516 = ~n55 & ~n515 ;
  assign n514 = ~\v10_reg/NET0131  & \v7_reg/NET0131  ;
  assign n517 = n53 & ~n514 ;
  assign n518 = ~n516 & n517 ;
  assign n519 = ~n513 & ~n518 ;
  assign n520 = \v11_reg/NET0131  & ~n519 ;
  assign n503 = n100 & n480 ;
  assign n505 = n27 & ~n504 ;
  assign n506 = n118 & ~n139 ;
  assign n507 = ~n505 & n506 ;
  assign n508 = ~n503 & ~n507 ;
  assign n509 = ~\v7_reg/NET0131  & ~n508 ;
  assign n521 = n53 & n514 ;
  assign n522 = ~\v5_pad  & n18 ;
  assign n523 = n155 & n522 ;
  assign n524 = ~n521 & ~n523 ;
  assign n525 = ~\v0_pad  & n47 ;
  assign n526 = ~n524 & n525 ;
  assign n527 = ~n509 & ~n526 ;
  assign n528 = ~n520 & n527 ;
  assign n529 = ~n190 & ~n326 ;
  assign n530 = n62 & ~n529 ;
  assign n531 = n71 & n75 ;
  assign n532 = ~n530 & ~n531 ;
  assign n533 = \v7_reg/NET0131  & ~n532 ;
  assign n534 = ~n16 & ~n119 ;
  assign n535 = ~\v8_reg/NET0131  & ~n534 ;
  assign n536 = ~\v12_reg/NET0131  & n94 ;
  assign n537 = ~n535 & ~n536 ;
  assign n538 = ~\v9_reg/NET0131  & ~n537 ;
  assign n539 = ~n201 & ~n300 ;
  assign n540 = ~\v12_reg/NET0131  & ~n181 ;
  assign n541 = ~n539 & n540 ;
  assign n542 = ~n538 & ~n541 ;
  assign n543 = ~\v7_reg/NET0131  & ~n542 ;
  assign n544 = ~n533 & ~n543 ;
  assign n553 = \v11_reg/NET0131  & ~n228 ;
  assign n554 = ~\v9_reg/NET0131  & ~n16 ;
  assign n555 = ~n553 & n554 ;
  assign n556 = ~\v8_reg/NET0131  & ~n555 ;
  assign n548 = ~\v8_reg/NET0131  & ~n15 ;
  assign n549 = \v10_reg/NET0131  & n252 ;
  assign n550 = ~n548 & ~n549 ;
  assign n551 = ~\v9_reg/NET0131  & ~n550 ;
  assign n552 = ~\v11_reg/NET0131  & ~n551 ;
  assign n545 = \v11_reg/NET0131  & ~\v8_reg/NET0131  ;
  assign n546 = ~n175 & ~n545 ;
  assign n547 = ~n181 & ~n546 ;
  assign n557 = n112 & ~n346 ;
  assign n558 = ~\v7_reg/NET0131  & ~n98 ;
  assign n559 = ~n557 & n558 ;
  assign n560 = ~n547 & n559 ;
  assign n561 = ~n552 & n560 ;
  assign n562 = ~n556 & n561 ;
  assign n563 = \v9_reg/NET0131  & ~n346 ;
  assign n564 = ~n39 & n350 ;
  assign n565 = ~n563 & n564 ;
  assign n566 = \v7_reg/NET0131  & ~n400 ;
  assign n567 = ~n565 & n566 ;
  assign n568 = ~n562 & ~n567 ;
  assign n569 = n46 & ~n47 ;
  assign n570 = ~n157 & n569 ;
  assign n571 = ~n568 & ~n570 ;
  assign n572 = ~\v9_reg/NET0131  & n53 ;
  assign n573 = ~n261 & ~n572 ;
  assign n574 = n209 & ~n573 ;
  assign n575 = ~n310 & ~n545 ;
  assign n576 = \v9_reg/NET0131  & ~n345 ;
  assign n577 = ~n575 & n576 ;
  assign n578 = ~n574 & ~n577 ;
  assign n579 = ~\v12_reg/NET0131  & ~n578 ;
  assign \_al_n0  = 1'b0 ;
  assign \_al_n1  = ~1'b0 ;
  assign \g1757/_0_  = n85 ;
  assign \g1763/_1_  = n154 ;
  assign \g1787/_3_  = ~n174 ;
  assign \g1800/_3_  = ~n198 ;
  assign \g1821/_2_  = n206 ;
  assign \g1940/_1_  = n212 ;
  assign \g25/_0_  = n260 ;
  assign \g2783/_3_  = ~n283 ;
  assign \g2823/_0_  = n319 ;
  assign \g38/_1_  = n365 ;
  assign \g40/_1_  = n399 ;
  assign \v13_D_11_pad  = ~n413 ;
  assign \v13_D_12_pad  = ~n429 ;
  assign \v13_D_13_pad  = ~n455 ;
  assign \v13_D_14_pad  = ~n467 ;
  assign \v13_D_16_pad  = n470 ;
  assign \v13_D_18_pad  = n477 ;
  assign \v13_D_19_pad  = ~n484 ;
  assign \v13_D_21_pad  = n489 ;
  assign \v13_D_22_pad  = ~n496 ;
  assign \v13_D_23_pad  = n502 ;
  assign \v13_D_24_pad  = ~n528 ;
  assign \v13_D_7_pad  = ~n544 ;
  assign \v13_D_8_pad  = ~n571 ;
  assign \v13_D_9_pad  = n579 ;
endmodule
