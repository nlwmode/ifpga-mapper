module top( a_pad , b_pad , c_pad , d_pad , e_pad , f_pad , g_pad , h_pad , i_pad , j_pad , k_pad , l_pad , m_pad , n_pad , o_pad , p_pad , q_pad , r_pad , s_pad , t_pad , u_pad );
  input a_pad ;
  input b_pad ;
  input c_pad ;
  input d_pad ;
  input e_pad ;
  input f_pad ;
  input g_pad ;
  input h_pad ;
  input i_pad ;
  input j_pad ;
  input k_pad ;
  input l_pad ;
  input m_pad ;
  input n_pad ;
  input o_pad ;
  input p_pad ;
  output q_pad ;
  output r_pad ;
  output s_pad ;
  output t_pad ;
  output u_pad ;
  wire n17 , n18 , n19 , n20 , n21 , n22 , n23 , n24 , n25 , n26 , n27 , n28 , n29 , n30 , n31 , n32 , n33 , n34 , n35 , n36 , n37 , n38 , n39 , n40 , n41 , n42 , n43 , n44 , n45 , n46 , n47 , n48 ;
  assign n17 = ~e_pad & f_pad ;
  assign n18 = a_pad & n17 ;
  assign n19 = c_pad & d_pad ;
  assign n21 = j_pad & ~n19 ;
  assign n20 = ~j_pad & n19 ;
  assign n22 = e_pad & f_pad ;
  assign n23 = ~n20 & n22 ;
  assign n24 = ~n21 & n23 ;
  assign n25 = ~n18 & ~n24 ;
  assign n26 = b_pad & n17 ;
  assign n28 = l_pad & ~n20 ;
  assign n27 = ~l_pad & n20 ;
  assign n29 = n22 & ~n27 ;
  assign n30 = ~n28 & n29 ;
  assign n31 = ~n26 & ~n30 ;
  assign n32 = g_pad & n17 ;
  assign n33 = m_pad & ~n27 ;
  assign n34 = ~l_pad & ~m_pad ;
  assign n35 = n20 & n34 ;
  assign n36 = n22 & ~n35 ;
  assign n37 = ~n33 & n36 ;
  assign n38 = ~n32 & ~n37 ;
  assign n39 = h_pad & n17 ;
  assign n41 = ~n_pad & n35 ;
  assign n40 = n_pad & ~n35 ;
  assign n42 = n22 & ~n40 ;
  assign n43 = ~n41 & n42 ;
  assign n44 = ~n39 & ~n43 ;
  assign n45 = d_pad & i_pad ;
  assign n46 = k_pad & o_pad ;
  assign n47 = p_pad & n46 ;
  assign n48 = n45 & n47 ;
  assign q_pad = n25 ;
  assign r_pad = n31 ;
  assign s_pad = n38 ;
  assign t_pad = n44 ;
  assign u_pad = n48 ;
endmodule
