module top (\g102_pad , \g10_reg/NET0131 , \g11_reg/NET0131 , \g1293_pad , \g14_reg/NET0131 , \g15_reg/NET0131 , \g18_reg/NET0131 , \g197_reg/NET0131 , \g19_reg/NET0131 , \g1_reg/NET0131 , \g204_reg/NET0131 , \g205_reg/NET0131 , \g206_reg/NET0131 , \g207_reg/NET0131 , \g208_reg/NET0131 , \g209_reg/NET0131 , \g210_reg/NET0131 , \g211_reg/NET0131 , \g212_reg/NET0131 , \g218_reg/NET0131 , \g224_reg/NET0131 , \g230_reg/NET0131 , \g236_reg/NET0131 , \g242_reg/NET0131 , \g248_reg/NET0131 , \g24_reg/NET0131 , \g254_reg/NET0131 , \g25_reg/NET0131 , \g260_reg/NET0131 , \g266_reg/NET0131 , \g269_reg/NET0131 , \g276_reg/NET0131 , \g277_reg/NET0131 , \g278_reg/NET0131 , \g279_reg/NET0131 , \g280_reg/NET0131 , \g281_reg/NET0131 , \g282_reg/NET0131 , \g283_reg/NET0131 , \g28_reg/NET0131 , \g293_reg/NET0131 , \g297_reg/NET0131 , \g29_reg/NET0131 , \g2_reg/NET0131 , \g33_reg/NET0131 , \g3_reg/NET0131 , \g402_reg/NET0131 , \g406_reg/NET0131 , \g4099_pad , \g4100_pad , \g4101_pad , \g4102_pad , \g4103_pad , \g4104_pad , \g4105_pad , \g4108_pad , \g410_reg/NET0131 , \g4110_pad , \g4112_pad , \g414_reg/NET0131 , \g418_reg/NET0131 , \g422_reg/NET0131 , \g426_reg/NET0131 , \g430_reg/NET0131 , \g434_reg/NET0131 , \g437_reg/NET0131 , \g441_reg/NET0131 , \g4422_pad , \g445_reg/NET0131 , \g449_reg/NET0131 , \g453_reg/NET0131 , \g457_reg/NET0131 , \g461_reg/NET0131 , \g465_reg/NET0131 , \g471_reg/NET0131 , \g478_reg/NET0131 , \g486_reg/NET0131 , \g489_reg/NET0131 , \g48_reg/NET0131 , \g492_reg/NET0131 , \g496_reg/NET0131 , \g500_reg/NET0131 , \g504_reg/NET0131 , \g508_reg/NET0131 , \g512_reg/NET0131 , \g536_reg/NET0131 , \g541_reg/NET0131 , \g545_reg/NET0131 , \g548_reg/NET0131 , \g551_reg/NET0131 , \g554_reg/NET0131 , \g557_pad , \g558_pad , \g559_pad , \g560_pad , \g561_pad , \g562_pad , \g563_pad , \g567_pad , \g571_reg/NET0131 , \g574_reg/NET0131 , \g578_reg/NET0131 , \g582_reg/NET0131 , \g586_reg/NET0131 , \g590_reg/NET0131 , \g594_reg/NET0131 , \g598_reg/NET0131 , \g602_reg/NET0131 , \g606_reg/NET0131 , \g610_reg/NET0131 , \g613_reg/NET0131 , \g616_reg/NET0131 , \g619_reg/NET0131 , \g622_reg/NET0131 , \g625_reg/NET0131 , \g628_reg/NET0131 , \g631_reg/NET0131 , \g634_reg/NET0131 , \g638_reg/NET0131 , \g639_pad , \g642_reg/NET0131 , \g646_reg/NET0131 , \g650_reg/NET0131 , \g654_reg/NET0131 , \g662_reg/NET0131 , \g669_reg/NET0131 , \g672_reg/NET0131 , \g675_reg/NET0131 , \g676_reg/NET0131 , \g677_reg/NET0131 , \g678_reg/NET0131 , \g679_reg/NET0131 , \g680_reg/NET0131 , \g681_reg/NET0131 , \g682_reg/NET0131 , \g683_reg/NET0131 , \g684_reg/NET0131 , \g685_reg/NET0131 , \g687_reg/NET0131 , \g688_reg/NET0131 , \g689_reg/NET0131 , \g698_reg/NET0131 , \g6_reg/NET0131 , \g702_pad , \g7_reg/NET0131 , \g89_pad , \_al_n1 , \g10560/_0_ , \g10562/_1_ , \g10564/_1_ , \g10566/_1_ , \g10567/_0_ , \g10569/_1_ , \g10580/_0_ , \g10616/_2_ , \g10627/_2_ , \g10628/_0_ , \g10629/_2_ , \g10630/_2_ , \g10633/_2_ , \g10635/_2_ , \g10636/_2_ , \g10637/_2_ , \g10641/_0_ , \g10649/_0_ , \g10672/_0_ , \g10673/_0_ , \g10680/_0_ , \g10683/_0_ , \g10686/_0_ , \g10695/_0_ , \g10700/_0_ , \g10703/_0_ , \g10704/_0_ , \g10748/_0_ , \g10750/_2_ , \g10757/_0_ , \g10758/_0_ , \g10782/_0_ , \g10826/_0_ , \g10827/_0_ , \g10828/_1_ , \g10832/_2_ , \g10834/_2_ , \g10836/_0_ , \g10837/_1__syn_2 , \g10868/_0_ , \g10904/_0_ , \g10913/_0_ , \g10915/_0_ , \g10922/_0_ , \g10938/_0_ , \g10939/_0_ , \g10940/_0_ , \g10941/_0_ , \g10942/_0_ , \g10944/_2_ , \g10977/_0_ , \g10980/_0_ , \g11020/_0_ , \g11028/_0_ , \g11051/_0_ , \g11057/_0_ , \g11109/_0_ , \g11113/_2_ , \g11156/_0_ , \g11172/_3_ , \g11193/_0_ , \g11219/_0_ , \g11355/_0_ , \g11384/_0_ , \g11442/_0_ , \g11448/_0_ , \g11558/_0_ , \g11559/_0_ , \g11824/_1_ , \g11853/_0_ , \g11854/_0_ , \g11977/_0_ , \g11981/_0_ , \g2584_pad , \g4121_pad , \g4809_pad , \g5692_pad , \g6282_pad , \g6284_pad , \g6360_pad , \g6362_pad , \g6364_pad , \g6366_pad , \g6368_pad , \g6370_pad , \g6372_pad , \g6374_pad );
	input \g102_pad  ;
	input \g10_reg/NET0131  ;
	input \g11_reg/NET0131  ;
	input \g1293_pad  ;
	input \g14_reg/NET0131  ;
	input \g15_reg/NET0131  ;
	input \g18_reg/NET0131  ;
	input \g197_reg/NET0131  ;
	input \g19_reg/NET0131  ;
	input \g1_reg/NET0131  ;
	input \g204_reg/NET0131  ;
	input \g205_reg/NET0131  ;
	input \g206_reg/NET0131  ;
	input \g207_reg/NET0131  ;
	input \g208_reg/NET0131  ;
	input \g209_reg/NET0131  ;
	input \g210_reg/NET0131  ;
	input \g211_reg/NET0131  ;
	input \g212_reg/NET0131  ;
	input \g218_reg/NET0131  ;
	input \g224_reg/NET0131  ;
	input \g230_reg/NET0131  ;
	input \g236_reg/NET0131  ;
	input \g242_reg/NET0131  ;
	input \g248_reg/NET0131  ;
	input \g24_reg/NET0131  ;
	input \g254_reg/NET0131  ;
	input \g25_reg/NET0131  ;
	input \g260_reg/NET0131  ;
	input \g266_reg/NET0131  ;
	input \g269_reg/NET0131  ;
	input \g276_reg/NET0131  ;
	input \g277_reg/NET0131  ;
	input \g278_reg/NET0131  ;
	input \g279_reg/NET0131  ;
	input \g280_reg/NET0131  ;
	input \g281_reg/NET0131  ;
	input \g282_reg/NET0131  ;
	input \g283_reg/NET0131  ;
	input \g28_reg/NET0131  ;
	input \g293_reg/NET0131  ;
	input \g297_reg/NET0131  ;
	input \g29_reg/NET0131  ;
	input \g2_reg/NET0131  ;
	input \g33_reg/NET0131  ;
	input \g3_reg/NET0131  ;
	input \g402_reg/NET0131  ;
	input \g406_reg/NET0131  ;
	input \g4099_pad  ;
	input \g4100_pad  ;
	input \g4101_pad  ;
	input \g4102_pad  ;
	input \g4103_pad  ;
	input \g4104_pad  ;
	input \g4105_pad  ;
	input \g4108_pad  ;
	input \g410_reg/NET0131  ;
	input \g4110_pad  ;
	input \g4112_pad  ;
	input \g414_reg/NET0131  ;
	input \g418_reg/NET0131  ;
	input \g422_reg/NET0131  ;
	input \g426_reg/NET0131  ;
	input \g430_reg/NET0131  ;
	input \g434_reg/NET0131  ;
	input \g437_reg/NET0131  ;
	input \g441_reg/NET0131  ;
	input \g4422_pad  ;
	input \g445_reg/NET0131  ;
	input \g449_reg/NET0131  ;
	input \g453_reg/NET0131  ;
	input \g457_reg/NET0131  ;
	input \g461_reg/NET0131  ;
	input \g465_reg/NET0131  ;
	input \g471_reg/NET0131  ;
	input \g478_reg/NET0131  ;
	input \g486_reg/NET0131  ;
	input \g489_reg/NET0131  ;
	input \g48_reg/NET0131  ;
	input \g492_reg/NET0131  ;
	input \g496_reg/NET0131  ;
	input \g500_reg/NET0131  ;
	input \g504_reg/NET0131  ;
	input \g508_reg/NET0131  ;
	input \g512_reg/NET0131  ;
	input \g536_reg/NET0131  ;
	input \g541_reg/NET0131  ;
	input \g545_reg/NET0131  ;
	input \g548_reg/NET0131  ;
	input \g551_reg/NET0131  ;
	input \g554_reg/NET0131  ;
	input \g557_pad  ;
	input \g558_pad  ;
	input \g559_pad  ;
	input \g560_pad  ;
	input \g561_pad  ;
	input \g562_pad  ;
	input \g563_pad  ;
	input \g567_pad  ;
	input \g571_reg/NET0131  ;
	input \g574_reg/NET0131  ;
	input \g578_reg/NET0131  ;
	input \g582_reg/NET0131  ;
	input \g586_reg/NET0131  ;
	input \g590_reg/NET0131  ;
	input \g594_reg/NET0131  ;
	input \g598_reg/NET0131  ;
	input \g602_reg/NET0131  ;
	input \g606_reg/NET0131  ;
	input \g610_reg/NET0131  ;
	input \g613_reg/NET0131  ;
	input \g616_reg/NET0131  ;
	input \g619_reg/NET0131  ;
	input \g622_reg/NET0131  ;
	input \g625_reg/NET0131  ;
	input \g628_reg/NET0131  ;
	input \g631_reg/NET0131  ;
	input \g634_reg/NET0131  ;
	input \g638_reg/NET0131  ;
	input \g639_pad  ;
	input \g642_reg/NET0131  ;
	input \g646_reg/NET0131  ;
	input \g650_reg/NET0131  ;
	input \g654_reg/NET0131  ;
	input \g662_reg/NET0131  ;
	input \g669_reg/NET0131  ;
	input \g672_reg/NET0131  ;
	input \g675_reg/NET0131  ;
	input \g676_reg/NET0131  ;
	input \g677_reg/NET0131  ;
	input \g678_reg/NET0131  ;
	input \g679_reg/NET0131  ;
	input \g680_reg/NET0131  ;
	input \g681_reg/NET0131  ;
	input \g682_reg/NET0131  ;
	input \g683_reg/NET0131  ;
	input \g684_reg/NET0131  ;
	input \g685_reg/NET0131  ;
	input \g687_reg/NET0131  ;
	input \g688_reg/NET0131  ;
	input \g689_reg/NET0131  ;
	input \g698_reg/NET0131  ;
	input \g6_reg/NET0131  ;
	input \g702_pad  ;
	input \g7_reg/NET0131  ;
	input \g89_pad  ;
	output \_al_n1  ;
	output \g10560/_0_  ;
	output \g10562/_1_  ;
	output \g10564/_1_  ;
	output \g10566/_1_  ;
	output \g10567/_0_  ;
	output \g10569/_1_  ;
	output \g10580/_0_  ;
	output \g10616/_2_  ;
	output \g10627/_2_  ;
	output \g10628/_0_  ;
	output \g10629/_2_  ;
	output \g10630/_2_  ;
	output \g10633/_2_  ;
	output \g10635/_2_  ;
	output \g10636/_2_  ;
	output \g10637/_2_  ;
	output \g10641/_0_  ;
	output \g10649/_0_  ;
	output \g10672/_0_  ;
	output \g10673/_0_  ;
	output \g10680/_0_  ;
	output \g10683/_0_  ;
	output \g10686/_0_  ;
	output \g10695/_0_  ;
	output \g10700/_0_  ;
	output \g10703/_0_  ;
	output \g10704/_0_  ;
	output \g10748/_0_  ;
	output \g10750/_2_  ;
	output \g10757/_0_  ;
	output \g10758/_0_  ;
	output \g10782/_0_  ;
	output \g10826/_0_  ;
	output \g10827/_0_  ;
	output \g10828/_1_  ;
	output \g10832/_2_  ;
	output \g10834/_2_  ;
	output \g10836/_0_  ;
	output \g10837/_1__syn_2  ;
	output \g10868/_0_  ;
	output \g10904/_0_  ;
	output \g10913/_0_  ;
	output \g10915/_0_  ;
	output \g10922/_0_  ;
	output \g10938/_0_  ;
	output \g10939/_0_  ;
	output \g10940/_0_  ;
	output \g10941/_0_  ;
	output \g10942/_0_  ;
	output \g10944/_2_  ;
	output \g10977/_0_  ;
	output \g10980/_0_  ;
	output \g11020/_0_  ;
	output \g11028/_0_  ;
	output \g11051/_0_  ;
	output \g11057/_0_  ;
	output \g11109/_0_  ;
	output \g11113/_2_  ;
	output \g11156/_0_  ;
	output \g11172/_3_  ;
	output \g11193/_0_  ;
	output \g11219/_0_  ;
	output \g11355/_0_  ;
	output \g11384/_0_  ;
	output \g11442/_0_  ;
	output \g11448/_0_  ;
	output \g11558/_0_  ;
	output \g11559/_0_  ;
	output \g11824/_1_  ;
	output \g11853/_0_  ;
	output \g11854/_0_  ;
	output \g11977/_0_  ;
	output \g11981/_0_  ;
	output \g2584_pad  ;
	output \g4121_pad  ;
	output \g4809_pad  ;
	output \g5692_pad  ;
	output \g6282_pad  ;
	output \g6284_pad  ;
	output \g6360_pad  ;
	output \g6362_pad  ;
	output \g6364_pad  ;
	output \g6366_pad  ;
	output \g6368_pad  ;
	output \g6370_pad  ;
	output \g6372_pad  ;
	output \g6374_pad  ;
	wire _w813_ ;
	wire _w812_ ;
	wire _w811_ ;
	wire _w810_ ;
	wire _w809_ ;
	wire _w808_ ;
	wire _w807_ ;
	wire _w806_ ;
	wire _w805_ ;
	wire _w804_ ;
	wire _w803_ ;
	wire _w802_ ;
	wire _w801_ ;
	wire _w800_ ;
	wire _w799_ ;
	wire _w798_ ;
	wire _w797_ ;
	wire _w796_ ;
	wire _w795_ ;
	wire _w794_ ;
	wire _w793_ ;
	wire _w792_ ;
	wire _w791_ ;
	wire _w790_ ;
	wire _w789_ ;
	wire _w788_ ;
	wire _w787_ ;
	wire _w786_ ;
	wire _w785_ ;
	wire _w784_ ;
	wire _w783_ ;
	wire _w782_ ;
	wire _w781_ ;
	wire _w780_ ;
	wire _w779_ ;
	wire _w778_ ;
	wire _w777_ ;
	wire _w776_ ;
	wire _w775_ ;
	wire _w774_ ;
	wire _w773_ ;
	wire _w772_ ;
	wire _w771_ ;
	wire _w770_ ;
	wire _w769_ ;
	wire _w768_ ;
	wire _w767_ ;
	wire _w766_ ;
	wire _w765_ ;
	wire _w764_ ;
	wire _w763_ ;
	wire _w762_ ;
	wire _w761_ ;
	wire _w760_ ;
	wire _w759_ ;
	wire _w758_ ;
	wire _w757_ ;
	wire _w756_ ;
	wire _w755_ ;
	wire _w754_ ;
	wire _w753_ ;
	wire _w752_ ;
	wire _w751_ ;
	wire _w750_ ;
	wire _w749_ ;
	wire _w748_ ;
	wire _w747_ ;
	wire _w746_ ;
	wire _w745_ ;
	wire _w744_ ;
	wire _w743_ ;
	wire _w742_ ;
	wire _w741_ ;
	wire _w740_ ;
	wire _w739_ ;
	wire _w738_ ;
	wire _w737_ ;
	wire _w736_ ;
	wire _w735_ ;
	wire _w734_ ;
	wire _w733_ ;
	wire _w732_ ;
	wire _w731_ ;
	wire _w730_ ;
	wire _w729_ ;
	wire _w728_ ;
	wire _w727_ ;
	wire _w726_ ;
	wire _w725_ ;
	wire _w724_ ;
	wire _w723_ ;
	wire _w722_ ;
	wire _w721_ ;
	wire _w720_ ;
	wire _w719_ ;
	wire _w718_ ;
	wire _w717_ ;
	wire _w716_ ;
	wire _w715_ ;
	wire _w714_ ;
	wire _w713_ ;
	wire _w712_ ;
	wire _w711_ ;
	wire _w710_ ;
	wire _w709_ ;
	wire _w708_ ;
	wire _w707_ ;
	wire _w706_ ;
	wire _w705_ ;
	wire _w704_ ;
	wire _w703_ ;
	wire _w702_ ;
	wire _w701_ ;
	wire _w700_ ;
	wire _w699_ ;
	wire _w698_ ;
	wire _w697_ ;
	wire _w696_ ;
	wire _w695_ ;
	wire _w694_ ;
	wire _w693_ ;
	wire _w692_ ;
	wire _w691_ ;
	wire _w690_ ;
	wire _w689_ ;
	wire _w688_ ;
	wire _w403_ ;
	wire _w402_ ;
	wire _w401_ ;
	wire _w400_ ;
	wire _w399_ ;
	wire _w398_ ;
	wire _w397_ ;
	wire _w396_ ;
	wire _w395_ ;
	wire _w394_ ;
	wire _w393_ ;
	wire _w392_ ;
	wire _w391_ ;
	wire _w390_ ;
	wire _w389_ ;
	wire _w388_ ;
	wire _w387_ ;
	wire _w386_ ;
	wire _w385_ ;
	wire _w384_ ;
	wire _w383_ ;
	wire _w382_ ;
	wire _w381_ ;
	wire _w380_ ;
	wire _w379_ ;
	wire _w378_ ;
	wire _w377_ ;
	wire _w376_ ;
	wire _w375_ ;
	wire _w374_ ;
	wire _w373_ ;
	wire _w372_ ;
	wire _w371_ ;
	wire _w370_ ;
	wire _w369_ ;
	wire _w368_ ;
	wire _w367_ ;
	wire _w366_ ;
	wire _w365_ ;
	wire _w364_ ;
	wire _w363_ ;
	wire _w362_ ;
	wire _w361_ ;
	wire _w360_ ;
	wire _w359_ ;
	wire _w358_ ;
	wire _w357_ ;
	wire _w356_ ;
	wire _w355_ ;
	wire _w354_ ;
	wire _w353_ ;
	wire _w352_ ;
	wire _w351_ ;
	wire _w350_ ;
	wire _w349_ ;
	wire _w348_ ;
	wire _w347_ ;
	wire _w346_ ;
	wire _w345_ ;
	wire _w344_ ;
	wire _w343_ ;
	wire _w342_ ;
	wire _w341_ ;
	wire _w340_ ;
	wire _w339_ ;
	wire _w338_ ;
	wire _w337_ ;
	wire _w336_ ;
	wire _w335_ ;
	wire _w334_ ;
	wire _w333_ ;
	wire _w332_ ;
	wire _w331_ ;
	wire _w330_ ;
	wire _w329_ ;
	wire _w328_ ;
	wire _w327_ ;
	wire _w326_ ;
	wire _w325_ ;
	wire _w324_ ;
	wire _w323_ ;
	wire _w322_ ;
	wire _w321_ ;
	wire _w320_ ;
	wire _w319_ ;
	wire _w318_ ;
	wire _w317_ ;
	wire _w316_ ;
	wire _w315_ ;
	wire _w314_ ;
	wire _w313_ ;
	wire _w312_ ;
	wire _w311_ ;
	wire _w310_ ;
	wire _w309_ ;
	wire _w308_ ;
	wire _w307_ ;
	wire _w306_ ;
	wire _w305_ ;
	wire _w304_ ;
	wire _w303_ ;
	wire _w302_ ;
	wire _w301_ ;
	wire _w300_ ;
	wire _w299_ ;
	wire _w298_ ;
	wire _w297_ ;
	wire _w296_ ;
	wire _w295_ ;
	wire _w294_ ;
	wire _w293_ ;
	wire _w292_ ;
	wire _w291_ ;
	wire _w290_ ;
	wire _w289_ ;
	wire _w288_ ;
	wire _w287_ ;
	wire _w286_ ;
	wire _w285_ ;
	wire _w284_ ;
	wire _w283_ ;
	wire _w282_ ;
	wire _w281_ ;
	wire _w280_ ;
	wire _w279_ ;
	wire _w278_ ;
	wire _w277_ ;
	wire _w276_ ;
	wire _w275_ ;
	wire _w274_ ;
	wire _w205_ ;
	wire _w204_ ;
	wire _w203_ ;
	wire _w202_ ;
	wire _w201_ ;
	wire _w200_ ;
	wire _w199_ ;
	wire _w198_ ;
	wire _w197_ ;
	wire _w196_ ;
	wire _w195_ ;
	wire _w194_ ;
	wire _w193_ ;
	wire _w192_ ;
	wire _w191_ ;
	wire _w190_ ;
	wire _w189_ ;
	wire _w188_ ;
	wire _w187_ ;
	wire _w186_ ;
	wire _w185_ ;
	wire _w184_ ;
	wire _w183_ ;
	wire _w182_ ;
	wire _w181_ ;
	wire _w180_ ;
	wire _w179_ ;
	wire _w178_ ;
	wire _w177_ ;
	wire _w176_ ;
	wire _w159_ ;
	wire _w158_ ;
	wire _w157_ ;
	wire _w156_ ;
	wire _w155_ ;
	wire _w154_ ;
	wire _w153_ ;
	wire _w152_ ;
	wire _w151_ ;
	wire _w150_ ;
	wire _w149_ ;
	wire _w148_ ;
	wire _w147_ ;
	wire _w160_ ;
	wire _w161_ ;
	wire _w162_ ;
	wire _w163_ ;
	wire _w164_ ;
	wire _w165_ ;
	wire _w166_ ;
	wire _w167_ ;
	wire _w168_ ;
	wire _w169_ ;
	wire _w170_ ;
	wire _w171_ ;
	wire _w172_ ;
	wire _w173_ ;
	wire _w174_ ;
	wire _w175_ ;
	wire _w206_ ;
	wire _w207_ ;
	wire _w208_ ;
	wire _w209_ ;
	wire _w210_ ;
	wire _w211_ ;
	wire _w212_ ;
	wire _w213_ ;
	wire _w214_ ;
	wire _w215_ ;
	wire _w216_ ;
	wire _w217_ ;
	wire _w218_ ;
	wire _w219_ ;
	wire _w220_ ;
	wire _w221_ ;
	wire _w222_ ;
	wire _w223_ ;
	wire _w224_ ;
	wire _w225_ ;
	wire _w226_ ;
	wire _w227_ ;
	wire _w228_ ;
	wire _w229_ ;
	wire _w230_ ;
	wire _w231_ ;
	wire _w232_ ;
	wire _w233_ ;
	wire _w234_ ;
	wire _w235_ ;
	wire _w236_ ;
	wire _w237_ ;
	wire _w238_ ;
	wire _w239_ ;
	wire _w240_ ;
	wire _w241_ ;
	wire _w242_ ;
	wire _w243_ ;
	wire _w244_ ;
	wire _w245_ ;
	wire _w246_ ;
	wire _w247_ ;
	wire _w248_ ;
	wire _w249_ ;
	wire _w250_ ;
	wire _w251_ ;
	wire _w252_ ;
	wire _w253_ ;
	wire _w254_ ;
	wire _w255_ ;
	wire _w256_ ;
	wire _w257_ ;
	wire _w258_ ;
	wire _w259_ ;
	wire _w260_ ;
	wire _w261_ ;
	wire _w262_ ;
	wire _w263_ ;
	wire _w264_ ;
	wire _w265_ ;
	wire _w266_ ;
	wire _w267_ ;
	wire _w268_ ;
	wire _w269_ ;
	wire _w270_ ;
	wire _w271_ ;
	wire _w272_ ;
	wire _w273_ ;
	wire _w404_ ;
	wire _w405_ ;
	wire _w406_ ;
	wire _w407_ ;
	wire _w408_ ;
	wire _w409_ ;
	wire _w410_ ;
	wire _w411_ ;
	wire _w412_ ;
	wire _w413_ ;
	wire _w414_ ;
	wire _w415_ ;
	wire _w416_ ;
	wire _w417_ ;
	wire _w418_ ;
	wire _w419_ ;
	wire _w420_ ;
	wire _w421_ ;
	wire _w422_ ;
	wire _w423_ ;
	wire _w424_ ;
	wire _w425_ ;
	wire _w426_ ;
	wire _w427_ ;
	wire _w428_ ;
	wire _w429_ ;
	wire _w430_ ;
	wire _w431_ ;
	wire _w432_ ;
	wire _w433_ ;
	wire _w434_ ;
	wire _w435_ ;
	wire _w436_ ;
	wire _w437_ ;
	wire _w438_ ;
	wire _w439_ ;
	wire _w440_ ;
	wire _w441_ ;
	wire _w442_ ;
	wire _w443_ ;
	wire _w444_ ;
	wire _w445_ ;
	wire _w446_ ;
	wire _w447_ ;
	wire _w448_ ;
	wire _w449_ ;
	wire _w450_ ;
	wire _w451_ ;
	wire _w452_ ;
	wire _w453_ ;
	wire _w454_ ;
	wire _w455_ ;
	wire _w456_ ;
	wire _w457_ ;
	wire _w458_ ;
	wire _w459_ ;
	wire _w460_ ;
	wire _w461_ ;
	wire _w462_ ;
	wire _w463_ ;
	wire _w464_ ;
	wire _w465_ ;
	wire _w466_ ;
	wire _w467_ ;
	wire _w468_ ;
	wire _w469_ ;
	wire _w470_ ;
	wire _w471_ ;
	wire _w472_ ;
	wire _w473_ ;
	wire _w474_ ;
	wire _w475_ ;
	wire _w476_ ;
	wire _w477_ ;
	wire _w478_ ;
	wire _w479_ ;
	wire _w480_ ;
	wire _w481_ ;
	wire _w482_ ;
	wire _w483_ ;
	wire _w484_ ;
	wire _w485_ ;
	wire _w486_ ;
	wire _w487_ ;
	wire _w488_ ;
	wire _w489_ ;
	wire _w490_ ;
	wire _w491_ ;
	wire _w492_ ;
	wire _w493_ ;
	wire _w494_ ;
	wire _w495_ ;
	wire _w496_ ;
	wire _w497_ ;
	wire _w498_ ;
	wire _w499_ ;
	wire _w500_ ;
	wire _w501_ ;
	wire _w502_ ;
	wire _w503_ ;
	wire _w504_ ;
	wire _w505_ ;
	wire _w506_ ;
	wire _w507_ ;
	wire _w508_ ;
	wire _w509_ ;
	wire _w510_ ;
	wire _w511_ ;
	wire _w512_ ;
	wire _w513_ ;
	wire _w514_ ;
	wire _w515_ ;
	wire _w516_ ;
	wire _w517_ ;
	wire _w518_ ;
	wire _w519_ ;
	wire _w520_ ;
	wire _w521_ ;
	wire _w522_ ;
	wire _w523_ ;
	wire _w524_ ;
	wire _w525_ ;
	wire _w526_ ;
	wire _w527_ ;
	wire _w528_ ;
	wire _w529_ ;
	wire _w530_ ;
	wire _w531_ ;
	wire _w532_ ;
	wire _w533_ ;
	wire _w534_ ;
	wire _w535_ ;
	wire _w536_ ;
	wire _w537_ ;
	wire _w538_ ;
	wire _w539_ ;
	wire _w540_ ;
	wire _w541_ ;
	wire _w542_ ;
	wire _w543_ ;
	wire _w544_ ;
	wire _w545_ ;
	wire _w546_ ;
	wire _w547_ ;
	wire _w548_ ;
	wire _w549_ ;
	wire _w550_ ;
	wire _w551_ ;
	wire _w552_ ;
	wire _w553_ ;
	wire _w554_ ;
	wire _w555_ ;
	wire _w556_ ;
	wire _w557_ ;
	wire _w558_ ;
	wire _w559_ ;
	wire _w560_ ;
	wire _w561_ ;
	wire _w562_ ;
	wire _w563_ ;
	wire _w564_ ;
	wire _w565_ ;
	wire _w566_ ;
	wire _w567_ ;
	wire _w568_ ;
	wire _w569_ ;
	wire _w570_ ;
	wire _w571_ ;
	wire _w572_ ;
	wire _w573_ ;
	wire _w574_ ;
	wire _w575_ ;
	wire _w576_ ;
	wire _w577_ ;
	wire _w578_ ;
	wire _w579_ ;
	wire _w580_ ;
	wire _w581_ ;
	wire _w582_ ;
	wire _w583_ ;
	wire _w584_ ;
	wire _w585_ ;
	wire _w586_ ;
	wire _w587_ ;
	wire _w588_ ;
	wire _w589_ ;
	wire _w590_ ;
	wire _w591_ ;
	wire _w592_ ;
	wire _w593_ ;
	wire _w594_ ;
	wire _w595_ ;
	wire _w596_ ;
	wire _w597_ ;
	wire _w598_ ;
	wire _w599_ ;
	wire _w600_ ;
	wire _w601_ ;
	wire _w602_ ;
	wire _w603_ ;
	wire _w604_ ;
	wire _w605_ ;
	wire _w606_ ;
	wire _w607_ ;
	wire _w608_ ;
	wire _w609_ ;
	wire _w610_ ;
	wire _w611_ ;
	wire _w612_ ;
	wire _w613_ ;
	wire _w614_ ;
	wire _w615_ ;
	wire _w616_ ;
	wire _w617_ ;
	wire _w618_ ;
	wire _w619_ ;
	wire _w620_ ;
	wire _w621_ ;
	wire _w622_ ;
	wire _w623_ ;
	wire _w624_ ;
	wire _w625_ ;
	wire _w626_ ;
	wire _w627_ ;
	wire _w628_ ;
	wire _w629_ ;
	wire _w630_ ;
	wire _w631_ ;
	wire _w632_ ;
	wire _w633_ ;
	wire _w634_ ;
	wire _w635_ ;
	wire _w636_ ;
	wire _w637_ ;
	wire _w638_ ;
	wire _w639_ ;
	wire _w640_ ;
	wire _w641_ ;
	wire _w642_ ;
	wire _w643_ ;
	wire _w644_ ;
	wire _w645_ ;
	wire _w646_ ;
	wire _w647_ ;
	wire _w648_ ;
	wire _w649_ ;
	wire _w650_ ;
	wire _w651_ ;
	wire _w652_ ;
	wire _w653_ ;
	wire _w654_ ;
	wire _w655_ ;
	wire _w656_ ;
	wire _w657_ ;
	wire _w658_ ;
	wire _w659_ ;
	wire _w660_ ;
	wire _w661_ ;
	wire _w662_ ;
	wire _w663_ ;
	wire _w664_ ;
	wire _w665_ ;
	wire _w666_ ;
	wire _w667_ ;
	wire _w668_ ;
	wire _w669_ ;
	wire _w670_ ;
	wire _w671_ ;
	wire _w672_ ;
	wire _w673_ ;
	wire _w674_ ;
	wire _w675_ ;
	wire _w676_ ;
	wire _w677_ ;
	wire _w678_ ;
	wire _w679_ ;
	wire _w680_ ;
	wire _w681_ ;
	wire _w682_ ;
	wire _w683_ ;
	wire _w684_ ;
	wire _w685_ ;
	wire _w686_ ;
	wire _w687_ ;
	LUT2 #(
		.INIT('h8)
	) name0 (
		\g602_reg/NET0131 ,
		\g610_reg/NET0131 ,
		_w147_
	);
	LUT2 #(
		.INIT('h8)
	) name1 (
		\g613_reg/NET0131 ,
		_w147_,
		_w148_
	);
	LUT2 #(
		.INIT('h8)
	) name2 (
		\g616_reg/NET0131 ,
		_w148_,
		_w149_
	);
	LUT2 #(
		.INIT('h8)
	) name3 (
		\g619_reg/NET0131 ,
		_w149_,
		_w150_
	);
	LUT2 #(
		.INIT('h8)
	) name4 (
		\g622_reg/NET0131 ,
		_w150_,
		_w151_
	);
	LUT2 #(
		.INIT('h8)
	) name5 (
		\g625_reg/NET0131 ,
		_w151_,
		_w152_
	);
	LUT2 #(
		.INIT('h8)
	) name6 (
		\g628_reg/NET0131 ,
		_w152_,
		_w153_
	);
	LUT2 #(
		.INIT('h8)
	) name7 (
		\g631_reg/NET0131 ,
		_w153_,
		_w154_
	);
	LUT2 #(
		.INIT('h8)
	) name8 (
		\g578_reg/NET0131 ,
		_w154_,
		_w155_
	);
	LUT2 #(
		.INIT('h8)
	) name9 (
		\g582_reg/NET0131 ,
		_w155_,
		_w156_
	);
	LUT2 #(
		.INIT('h8)
	) name10 (
		\g586_reg/NET0131 ,
		_w156_,
		_w157_
	);
	LUT2 #(
		.INIT('h8)
	) name11 (
		\g574_reg/NET0131 ,
		_w157_,
		_w158_
	);
	LUT2 #(
		.INIT('h1)
	) name12 (
		\g590_reg/NET0131 ,
		_w158_,
		_w159_
	);
	LUT2 #(
		.INIT('h8)
	) name13 (
		\g590_reg/NET0131 ,
		_w158_,
		_w160_
	);
	LUT2 #(
		.INIT('h1)
	) name14 (
		_w159_,
		_w160_,
		_w161_
	);
	LUT2 #(
		.INIT('h8)
	) name15 (
		\g594_reg/NET0131 ,
		_w160_,
		_w162_
	);
	LUT2 #(
		.INIT('h2)
	) name16 (
		\g639_pad ,
		_w162_,
		_w163_
	);
	LUT2 #(
		.INIT('h4)
	) name17 (
		_w161_,
		_w163_,
		_w164_
	);
	LUT2 #(
		.INIT('h1)
	) name18 (
		\g582_reg/NET0131 ,
		_w155_,
		_w165_
	);
	LUT2 #(
		.INIT('h1)
	) name19 (
		_w156_,
		_w165_,
		_w166_
	);
	LUT2 #(
		.INIT('h8)
	) name20 (
		_w163_,
		_w166_,
		_w167_
	);
	LUT2 #(
		.INIT('h1)
	) name21 (
		\g586_reg/NET0131 ,
		_w156_,
		_w168_
	);
	LUT2 #(
		.INIT('h1)
	) name22 (
		_w157_,
		_w168_,
		_w169_
	);
	LUT2 #(
		.INIT('h8)
	) name23 (
		_w163_,
		_w169_,
		_w170_
	);
	LUT2 #(
		.INIT('h1)
	) name24 (
		\g594_reg/NET0131 ,
		_w160_,
		_w171_
	);
	LUT2 #(
		.INIT('h2)
	) name25 (
		_w163_,
		_w171_,
		_w172_
	);
	LUT2 #(
		.INIT('h1)
	) name26 (
		\g574_reg/NET0131 ,
		_w157_,
		_w173_
	);
	LUT2 #(
		.INIT('h1)
	) name27 (
		_w158_,
		_w173_,
		_w174_
	);
	LUT2 #(
		.INIT('h2)
	) name28 (
		_w163_,
		_w174_,
		_w175_
	);
	LUT2 #(
		.INIT('h1)
	) name29 (
		\g578_reg/NET0131 ,
		_w154_,
		_w176_
	);
	LUT2 #(
		.INIT('h1)
	) name30 (
		_w155_,
		_w176_,
		_w177_
	);
	LUT2 #(
		.INIT('h8)
	) name31 (
		_w163_,
		_w177_,
		_w178_
	);
	LUT2 #(
		.INIT('h2)
	) name32 (
		\g19_reg/NET0131 ,
		\g25_reg/NET0131 ,
		_w179_
	);
	LUT2 #(
		.INIT('h4)
	) name33 (
		\g19_reg/NET0131 ,
		\g25_reg/NET0131 ,
		_w180_
	);
	LUT2 #(
		.INIT('h1)
	) name34 (
		_w179_,
		_w180_,
		_w181_
	);
	LUT2 #(
		.INIT('h1)
	) name35 (
		\g3_reg/NET0131 ,
		\g7_reg/NET0131 ,
		_w182_
	);
	LUT2 #(
		.INIT('h8)
	) name36 (
		\g3_reg/NET0131 ,
		\g7_reg/NET0131 ,
		_w183_
	);
	LUT2 #(
		.INIT('h1)
	) name37 (
		_w182_,
		_w183_,
		_w184_
	);
	LUT2 #(
		.INIT('h8)
	) name38 (
		\g33_reg/NET0131 ,
		_w184_,
		_w185_
	);
	LUT2 #(
		.INIT('h1)
	) name39 (
		\g33_reg/NET0131 ,
		_w184_,
		_w186_
	);
	LUT2 #(
		.INIT('h1)
	) name40 (
		_w185_,
		_w186_,
		_w187_
	);
	LUT2 #(
		.INIT('h2)
	) name41 (
		\g11_reg/NET0131 ,
		\g15_reg/NET0131 ,
		_w188_
	);
	LUT2 #(
		.INIT('h4)
	) name42 (
		\g11_reg/NET0131 ,
		\g15_reg/NET0131 ,
		_w189_
	);
	LUT2 #(
		.INIT('h1)
	) name43 (
		_w188_,
		_w189_,
		_w190_
	);
	LUT2 #(
		.INIT('h8)
	) name44 (
		\g29_reg/NET0131 ,
		_w190_,
		_w191_
	);
	LUT2 #(
		.INIT('h1)
	) name45 (
		\g29_reg/NET0131 ,
		_w190_,
		_w192_
	);
	LUT2 #(
		.INIT('h1)
	) name46 (
		_w191_,
		_w192_,
		_w193_
	);
	LUT2 #(
		.INIT('h2)
	) name47 (
		_w187_,
		_w193_,
		_w194_
	);
	LUT2 #(
		.INIT('h4)
	) name48 (
		_w187_,
		_w193_,
		_w195_
	);
	LUT2 #(
		.INIT('h1)
	) name49 (
		_w194_,
		_w195_,
		_w196_
	);
	LUT2 #(
		.INIT('h8)
	) name50 (
		_w181_,
		_w196_,
		_w197_
	);
	LUT2 #(
		.INIT('h1)
	) name51 (
		_w181_,
		_w196_,
		_w198_
	);
	LUT2 #(
		.INIT('h1)
	) name52 (
		_w197_,
		_w198_,
		_w199_
	);
	LUT2 #(
		.INIT('h8)
	) name53 (
		\g1293_pad ,
		\g702_pad ,
		_w200_
	);
	LUT2 #(
		.INIT('h4)
	) name54 (
		\g266_reg/NET0131 ,
		\g4110_pad ,
		_w201_
	);
	LUT2 #(
		.INIT('h8)
	) name55 (
		\g662_reg/NET0131 ,
		_w201_,
		_w202_
	);
	LUT2 #(
		.INIT('h8)
	) name56 (
		_w200_,
		_w202_,
		_w203_
	);
	LUT2 #(
		.INIT('h8)
	) name57 (
		\g676_reg/NET0131 ,
		_w203_,
		_w204_
	);
	LUT2 #(
		.INIT('h4)
	) name58 (
		\g698_reg/NET0131 ,
		_w204_,
		_w205_
	);
	LUT2 #(
		.INIT('h1)
	) name59 (
		\g688_reg/NET0131 ,
		\g689_reg/NET0131 ,
		_w206_
	);
	LUT2 #(
		.INIT('h8)
	) name60 (
		_w205_,
		_w206_,
		_w207_
	);
	LUT2 #(
		.INIT('h4)
	) name61 (
		\g687_reg/NET0131 ,
		_w207_,
		_w208_
	);
	LUT2 #(
		.INIT('h8)
	) name62 (
		\g204_reg/NET0131 ,
		\g205_reg/NET0131 ,
		_w209_
	);
	LUT2 #(
		.INIT('h8)
	) name63 (
		\g206_reg/NET0131 ,
		_w209_,
		_w210_
	);
	LUT2 #(
		.INIT('h8)
	) name64 (
		\g207_reg/NET0131 ,
		_w210_,
		_w211_
	);
	LUT2 #(
		.INIT('h8)
	) name65 (
		\g208_reg/NET0131 ,
		_w211_,
		_w212_
	);
	LUT2 #(
		.INIT('h8)
	) name66 (
		\g209_reg/NET0131 ,
		_w212_,
		_w213_
	);
	LUT2 #(
		.INIT('h2)
	) name67 (
		\g208_reg/NET0131 ,
		\g209_reg/NET0131 ,
		_w214_
	);
	LUT2 #(
		.INIT('h4)
	) name68 (
		\g208_reg/NET0131 ,
		\g209_reg/NET0131 ,
		_w215_
	);
	LUT2 #(
		.INIT('h1)
	) name69 (
		_w214_,
		_w215_,
		_w216_
	);
	LUT2 #(
		.INIT('h8)
	) name70 (
		_w211_,
		_w215_,
		_w217_
	);
	LUT2 #(
		.INIT('h1)
	) name71 (
		_w216_,
		_w217_,
		_w218_
	);
	LUT2 #(
		.INIT('h1)
	) name72 (
		\g471_reg/NET0131 ,
		_w218_,
		_w219_
	);
	LUT2 #(
		.INIT('h2)
	) name73 (
		\g471_reg/NET0131 ,
		_w217_,
		_w220_
	);
	LUT2 #(
		.INIT('h1)
	) name74 (
		_w219_,
		_w220_,
		_w221_
	);
	LUT2 #(
		.INIT('h4)
	) name75 (
		\g204_reg/NET0131 ,
		\g680_reg/NET0131 ,
		_w222_
	);
	LUT2 #(
		.INIT('h8)
	) name76 (
		\g204_reg/NET0131 ,
		\g679_reg/NET0131 ,
		_w223_
	);
	LUT2 #(
		.INIT('h1)
	) name77 (
		\g205_reg/NET0131 ,
		_w222_,
		_w224_
	);
	LUT2 #(
		.INIT('h4)
	) name78 (
		_w223_,
		_w224_,
		_w225_
	);
	LUT2 #(
		.INIT('h8)
	) name79 (
		\g204_reg/NET0131 ,
		\g677_reg/NET0131 ,
		_w226_
	);
	LUT2 #(
		.INIT('h4)
	) name80 (
		\g204_reg/NET0131 ,
		\g678_reg/NET0131 ,
		_w227_
	);
	LUT2 #(
		.INIT('h2)
	) name81 (
		\g205_reg/NET0131 ,
		_w226_,
		_w228_
	);
	LUT2 #(
		.INIT('h4)
	) name82 (
		_w227_,
		_w228_,
		_w229_
	);
	LUT2 #(
		.INIT('h1)
	) name83 (
		_w225_,
		_w229_,
		_w230_
	);
	LUT2 #(
		.INIT('h2)
	) name84 (
		\g206_reg/NET0131 ,
		_w230_,
		_w231_
	);
	LUT2 #(
		.INIT('h4)
	) name85 (
		\g204_reg/NET0131 ,
		\g684_reg/NET0131 ,
		_w232_
	);
	LUT2 #(
		.INIT('h8)
	) name86 (
		\g204_reg/NET0131 ,
		\g683_reg/NET0131 ,
		_w233_
	);
	LUT2 #(
		.INIT('h1)
	) name87 (
		\g205_reg/NET0131 ,
		_w232_,
		_w234_
	);
	LUT2 #(
		.INIT('h4)
	) name88 (
		_w233_,
		_w234_,
		_w235_
	);
	LUT2 #(
		.INIT('h8)
	) name89 (
		\g204_reg/NET0131 ,
		\g681_reg/NET0131 ,
		_w236_
	);
	LUT2 #(
		.INIT('h4)
	) name90 (
		\g204_reg/NET0131 ,
		\g682_reg/NET0131 ,
		_w237_
	);
	LUT2 #(
		.INIT('h2)
	) name91 (
		\g205_reg/NET0131 ,
		_w236_,
		_w238_
	);
	LUT2 #(
		.INIT('h4)
	) name92 (
		_w237_,
		_w238_,
		_w239_
	);
	LUT2 #(
		.INIT('h1)
	) name93 (
		_w235_,
		_w239_,
		_w240_
	);
	LUT2 #(
		.INIT('h1)
	) name94 (
		\g206_reg/NET0131 ,
		_w240_,
		_w241_
	);
	LUT2 #(
		.INIT('h1)
	) name95 (
		_w231_,
		_w241_,
		_w242_
	);
	LUT2 #(
		.INIT('h1)
	) name96 (
		\g471_reg/NET0131 ,
		_w242_,
		_w243_
	);
	LUT2 #(
		.INIT('h8)
	) name97 (
		\g471_reg/NET0131 ,
		_w242_,
		_w244_
	);
	LUT2 #(
		.INIT('h2)
	) name98 (
		_w216_,
		_w243_,
		_w245_
	);
	LUT2 #(
		.INIT('h4)
	) name99 (
		_w244_,
		_w245_,
		_w246_
	);
	LUT2 #(
		.INIT('h1)
	) name100 (
		_w221_,
		_w246_,
		_w247_
	);
	LUT2 #(
		.INIT('h8)
	) name101 (
		\g210_reg/NET0131 ,
		\g211_reg/NET0131 ,
		_w248_
	);
	LUT2 #(
		.INIT('h4)
	) name102 (
		_w247_,
		_w248_,
		_w249_
	);
	LUT2 #(
		.INIT('h8)
	) name103 (
		_w213_,
		_w249_,
		_w250_
	);
	LUT2 #(
		.INIT('h4)
	) name104 (
		\g210_reg/NET0131 ,
		\g211_reg/NET0131 ,
		_w251_
	);
	LUT2 #(
		.INIT('h8)
	) name105 (
		_w213_,
		_w251_,
		_w252_
	);
	LUT2 #(
		.INIT('h2)
	) name106 (
		\g210_reg/NET0131 ,
		\g211_reg/NET0131 ,
		_w253_
	);
	LUT2 #(
		.INIT('h8)
	) name107 (
		_w213_,
		_w253_,
		_w254_
	);
	LUT2 #(
		.INIT('h8)
	) name108 (
		_w246_,
		_w254_,
		_w255_
	);
	LUT2 #(
		.INIT('h1)
	) name109 (
		\g210_reg/NET0131 ,
		\g211_reg/NET0131 ,
		_w256_
	);
	LUT2 #(
		.INIT('h4)
	) name110 (
		\g471_reg/NET0131 ,
		_w256_,
		_w257_
	);
	LUT2 #(
		.INIT('h4)
	) name111 (
		_w218_,
		_w257_,
		_w258_
	);
	LUT2 #(
		.INIT('h1)
	) name112 (
		_w252_,
		_w258_,
		_w259_
	);
	LUT2 #(
		.INIT('h4)
	) name113 (
		_w255_,
		_w259_,
		_w260_
	);
	LUT2 #(
		.INIT('h4)
	) name114 (
		_w250_,
		_w260_,
		_w261_
	);
	LUT2 #(
		.INIT('h8)
	) name115 (
		\g211_reg/NET0131 ,
		_w261_,
		_w262_
	);
	LUT2 #(
		.INIT('h4)
	) name116 (
		_w246_,
		_w254_,
		_w263_
	);
	LUT2 #(
		.INIT('h4)
	) name117 (
		_w213_,
		_w248_,
		_w264_
	);
	LUT2 #(
		.INIT('h4)
	) name118 (
		_w247_,
		_w264_,
		_w265_
	);
	LUT2 #(
		.INIT('h4)
	) name119 (
		_w212_,
		_w253_,
		_w266_
	);
	LUT2 #(
		.INIT('h8)
	) name120 (
		_w246_,
		_w266_,
		_w267_
	);
	LUT2 #(
		.INIT('h1)
	) name121 (
		_w265_,
		_w267_,
		_w268_
	);
	LUT2 #(
		.INIT('h4)
	) name122 (
		_w263_,
		_w268_,
		_w269_
	);
	LUT2 #(
		.INIT('h4)
	) name123 (
		_w262_,
		_w269_,
		_w270_
	);
	LUT2 #(
		.INIT('h2)
	) name124 (
		\g197_reg/NET0131 ,
		_w270_,
		_w271_
	);
	LUT2 #(
		.INIT('h4)
	) name125 (
		\g197_reg/NET0131 ,
		\g684_reg/NET0131 ,
		_w272_
	);
	LUT2 #(
		.INIT('h1)
	) name126 (
		_w271_,
		_w272_,
		_w273_
	);
	LUT2 #(
		.INIT('h2)
	) name127 (
		_w208_,
		_w273_,
		_w274_
	);
	LUT2 #(
		.INIT('h8)
	) name128 (
		\g687_reg/NET0131 ,
		_w207_,
		_w275_
	);
	LUT2 #(
		.INIT('h8)
	) name129 (
		\g276_reg/NET0131 ,
		\g277_reg/NET0131 ,
		_w276_
	);
	LUT2 #(
		.INIT('h8)
	) name130 (
		\g278_reg/NET0131 ,
		_w276_,
		_w277_
	);
	LUT2 #(
		.INIT('h8)
	) name131 (
		\g279_reg/NET0131 ,
		_w277_,
		_w278_
	);
	LUT2 #(
		.INIT('h8)
	) name132 (
		\g280_reg/NET0131 ,
		_w278_,
		_w279_
	);
	LUT2 #(
		.INIT('h8)
	) name133 (
		\g281_reg/NET0131 ,
		_w279_,
		_w280_
	);
	LUT2 #(
		.INIT('h4)
	) name134 (
		\g280_reg/NET0131 ,
		\g281_reg/NET0131 ,
		_w281_
	);
	LUT2 #(
		.INIT('h2)
	) name135 (
		\g280_reg/NET0131 ,
		\g281_reg/NET0131 ,
		_w282_
	);
	LUT2 #(
		.INIT('h1)
	) name136 (
		_w281_,
		_w282_,
		_w283_
	);
	LUT2 #(
		.INIT('h4)
	) name137 (
		\g276_reg/NET0131 ,
		\g680_reg/NET0131 ,
		_w284_
	);
	LUT2 #(
		.INIT('h8)
	) name138 (
		\g276_reg/NET0131 ,
		\g679_reg/NET0131 ,
		_w285_
	);
	LUT2 #(
		.INIT('h1)
	) name139 (
		\g277_reg/NET0131 ,
		_w284_,
		_w286_
	);
	LUT2 #(
		.INIT('h4)
	) name140 (
		_w285_,
		_w286_,
		_w287_
	);
	LUT2 #(
		.INIT('h8)
	) name141 (
		\g276_reg/NET0131 ,
		\g677_reg/NET0131 ,
		_w288_
	);
	LUT2 #(
		.INIT('h4)
	) name142 (
		\g276_reg/NET0131 ,
		\g678_reg/NET0131 ,
		_w289_
	);
	LUT2 #(
		.INIT('h2)
	) name143 (
		\g277_reg/NET0131 ,
		_w288_,
		_w290_
	);
	LUT2 #(
		.INIT('h4)
	) name144 (
		_w289_,
		_w290_,
		_w291_
	);
	LUT2 #(
		.INIT('h1)
	) name145 (
		_w287_,
		_w291_,
		_w292_
	);
	LUT2 #(
		.INIT('h2)
	) name146 (
		\g278_reg/NET0131 ,
		_w292_,
		_w293_
	);
	LUT2 #(
		.INIT('h4)
	) name147 (
		\g276_reg/NET0131 ,
		\g684_reg/NET0131 ,
		_w294_
	);
	LUT2 #(
		.INIT('h8)
	) name148 (
		\g276_reg/NET0131 ,
		\g683_reg/NET0131 ,
		_w295_
	);
	LUT2 #(
		.INIT('h1)
	) name149 (
		\g277_reg/NET0131 ,
		_w294_,
		_w296_
	);
	LUT2 #(
		.INIT('h4)
	) name150 (
		_w295_,
		_w296_,
		_w297_
	);
	LUT2 #(
		.INIT('h4)
	) name151 (
		\g276_reg/NET0131 ,
		\g682_reg/NET0131 ,
		_w298_
	);
	LUT2 #(
		.INIT('h8)
	) name152 (
		\g276_reg/NET0131 ,
		\g681_reg/NET0131 ,
		_w299_
	);
	LUT2 #(
		.INIT('h2)
	) name153 (
		\g277_reg/NET0131 ,
		_w298_,
		_w300_
	);
	LUT2 #(
		.INIT('h4)
	) name154 (
		_w299_,
		_w300_,
		_w301_
	);
	LUT2 #(
		.INIT('h1)
	) name155 (
		_w297_,
		_w301_,
		_w302_
	);
	LUT2 #(
		.INIT('h1)
	) name156 (
		\g278_reg/NET0131 ,
		_w302_,
		_w303_
	);
	LUT2 #(
		.INIT('h1)
	) name157 (
		_w293_,
		_w303_,
		_w304_
	);
	LUT2 #(
		.INIT('h2)
	) name158 (
		\g478_reg/NET0131 ,
		_w304_,
		_w305_
	);
	LUT2 #(
		.INIT('h4)
	) name159 (
		\g478_reg/NET0131 ,
		_w304_,
		_w306_
	);
	LUT2 #(
		.INIT('h1)
	) name160 (
		_w305_,
		_w306_,
		_w307_
	);
	LUT2 #(
		.INIT('h8)
	) name161 (
		_w283_,
		_w307_,
		_w308_
	);
	LUT2 #(
		.INIT('h8)
	) name162 (
		_w278_,
		_w281_,
		_w309_
	);
	LUT2 #(
		.INIT('h1)
	) name163 (
		_w283_,
		_w309_,
		_w310_
	);
	LUT2 #(
		.INIT('h2)
	) name164 (
		\g478_reg/NET0131 ,
		_w310_,
		_w311_
	);
	LUT2 #(
		.INIT('h4)
	) name165 (
		\g478_reg/NET0131 ,
		_w310_,
		_w312_
	);
	LUT2 #(
		.INIT('h1)
	) name166 (
		_w311_,
		_w312_,
		_w313_
	);
	LUT2 #(
		.INIT('h4)
	) name167 (
		_w283_,
		_w313_,
		_w314_
	);
	LUT2 #(
		.INIT('h8)
	) name168 (
		\g282_reg/NET0131 ,
		\g283_reg/NET0131 ,
		_w315_
	);
	LUT2 #(
		.INIT('h4)
	) name169 (
		_w314_,
		_w315_,
		_w316_
	);
	LUT2 #(
		.INIT('h4)
	) name170 (
		_w308_,
		_w316_,
		_w317_
	);
	LUT2 #(
		.INIT('h2)
	) name171 (
		\g282_reg/NET0131 ,
		_w317_,
		_w318_
	);
	LUT2 #(
		.INIT('h2)
	) name172 (
		_w280_,
		_w318_,
		_w319_
	);
	LUT2 #(
		.INIT('h2)
	) name173 (
		\g283_reg/NET0131 ,
		_w319_,
		_w320_
	);
	LUT2 #(
		.INIT('h2)
	) name174 (
		_w283_,
		_w307_,
		_w321_
	);
	LUT2 #(
		.INIT('h2)
	) name175 (
		\g282_reg/NET0131 ,
		\g283_reg/NET0131 ,
		_w322_
	);
	LUT2 #(
		.INIT('h8)
	) name176 (
		_w321_,
		_w322_,
		_w323_
	);
	LUT2 #(
		.INIT('h1)
	) name177 (
		_w317_,
		_w323_,
		_w324_
	);
	LUT2 #(
		.INIT('h1)
	) name178 (
		_w280_,
		_w324_,
		_w325_
	);
	LUT2 #(
		.INIT('h8)
	) name179 (
		_w280_,
		_w322_,
		_w326_
	);
	LUT2 #(
		.INIT('h4)
	) name180 (
		_w321_,
		_w326_,
		_w327_
	);
	LUT2 #(
		.INIT('h1)
	) name181 (
		_w325_,
		_w327_,
		_w328_
	);
	LUT2 #(
		.INIT('h4)
	) name182 (
		_w320_,
		_w328_,
		_w329_
	);
	LUT2 #(
		.INIT('h2)
	) name183 (
		\g269_reg/NET0131 ,
		_w329_,
		_w330_
	);
	LUT2 #(
		.INIT('h4)
	) name184 (
		\g269_reg/NET0131 ,
		\g684_reg/NET0131 ,
		_w331_
	);
	LUT2 #(
		.INIT('h1)
	) name185 (
		_w330_,
		_w331_,
		_w332_
	);
	LUT2 #(
		.INIT('h2)
	) name186 (
		_w275_,
		_w332_,
		_w333_
	);
	LUT2 #(
		.INIT('h8)
	) name187 (
		\g689_reg/NET0131 ,
		_w205_,
		_w334_
	);
	LUT2 #(
		.INIT('h8)
	) name188 (
		\g689_reg/NET0131 ,
		\g698_reg/NET0131 ,
		_w335_
	);
	LUT2 #(
		.INIT('h4)
	) name189 (
		\g688_reg/NET0131 ,
		_w335_,
		_w336_
	);
	LUT2 #(
		.INIT('h4)
	) name190 (
		\g685_reg/NET0131 ,
		_w336_,
		_w337_
	);
	LUT2 #(
		.INIT('h8)
	) name191 (
		_w204_,
		_w337_,
		_w338_
	);
	LUT2 #(
		.INIT('h1)
	) name192 (
		_w334_,
		_w338_,
		_w339_
	);
	LUT2 #(
		.INIT('h2)
	) name193 (
		\g684_reg/NET0131 ,
		_w339_,
		_w340_
	);
	LUT2 #(
		.INIT('h8)
	) name194 (
		\g685_reg/NET0131 ,
		_w336_,
		_w341_
	);
	LUT2 #(
		.INIT('h4)
	) name195 (
		\g682_reg/NET0131 ,
		_w341_,
		_w342_
	);
	LUT2 #(
		.INIT('h8)
	) name196 (
		\g683_reg/NET0131 ,
		\g684_reg/NET0131 ,
		_w343_
	);
	LUT2 #(
		.INIT('h4)
	) name197 (
		\g681_reg/NET0131 ,
		_w343_,
		_w344_
	);
	LUT2 #(
		.INIT('h8)
	) name198 (
		_w342_,
		_w344_,
		_w345_
	);
	LUT2 #(
		.INIT('h8)
	) name199 (
		_w203_,
		_w345_,
		_w346_
	);
	LUT2 #(
		.INIT('h8)
	) name200 (
		\g677_reg/NET0131 ,
		_w346_,
		_w347_
	);
	LUT2 #(
		.INIT('h8)
	) name201 (
		\g500_reg/NET0131 ,
		_w347_,
		_w348_
	);
	LUT2 #(
		.INIT('h1)
	) name202 (
		\g678_reg/NET0131 ,
		\g679_reg/NET0131 ,
		_w349_
	);
	LUT2 #(
		.INIT('h8)
	) name203 (
		\g688_reg/NET0131 ,
		_w335_,
		_w350_
	);
	LUT2 #(
		.INIT('h8)
	) name204 (
		_w203_,
		_w350_,
		_w351_
	);
	LUT2 #(
		.INIT('h8)
	) name205 (
		\g680_reg/NET0131 ,
		_w349_,
		_w352_
	);
	LUT2 #(
		.INIT('h8)
	) name206 (
		_w351_,
		_w352_,
		_w353_
	);
	LUT2 #(
		.INIT('h8)
	) name207 (
		\g684_reg/NET0131 ,
		_w341_,
		_w354_
	);
	LUT2 #(
		.INIT('h8)
	) name208 (
		_w203_,
		_w354_,
		_w355_
	);
	LUT2 #(
		.INIT('h4)
	) name209 (
		\g680_reg/NET0131 ,
		_w351_,
		_w356_
	);
	LUT2 #(
		.INIT('h4)
	) name210 (
		\g679_reg/NET0131 ,
		_w356_,
		_w357_
	);
	LUT2 #(
		.INIT('h8)
	) name211 (
		\g678_reg/NET0131 ,
		_w356_,
		_w358_
	);
	LUT2 #(
		.INIT('h8)
	) name212 (
		\g679_reg/NET0131 ,
		_w358_,
		_w359_
	);
	LUT2 #(
		.INIT('h1)
	) name213 (
		_w353_,
		_w355_,
		_w360_
	);
	LUT2 #(
		.INIT('h4)
	) name214 (
		_w207_,
		_w360_,
		_w361_
	);
	LUT2 #(
		.INIT('h4)
	) name215 (
		_w357_,
		_w361_,
		_w362_
	);
	LUT2 #(
		.INIT('h2)
	) name216 (
		_w339_,
		_w359_,
		_w363_
	);
	LUT2 #(
		.INIT('h8)
	) name217 (
		_w362_,
		_w363_,
		_w364_
	);
	LUT2 #(
		.INIT('h1)
	) name218 (
		_w348_,
		_w364_,
		_w365_
	);
	LUT2 #(
		.INIT('h8)
	) name219 (
		_w203_,
		_w343_,
		_w366_
	);
	LUT2 #(
		.INIT('h8)
	) name220 (
		\g682_reg/NET0131 ,
		_w341_,
		_w367_
	);
	LUT2 #(
		.INIT('h8)
	) name221 (
		_w366_,
		_w367_,
		_w368_
	);
	LUT2 #(
		.INIT('h4)
	) name222 (
		\g677_reg/NET0131 ,
		_w368_,
		_w369_
	);
	LUT2 #(
		.INIT('h8)
	) name223 (
		\g434_reg/NET0131 ,
		_w369_,
		_w370_
	);
	LUT2 #(
		.INIT('h8)
	) name224 (
		\g677_reg/NET0131 ,
		_w368_,
		_w371_
	);
	LUT2 #(
		.INIT('h8)
	) name225 (
		\g430_reg/NET0131 ,
		_w371_,
		_w372_
	);
	LUT2 #(
		.INIT('h8)
	) name226 (
		\g557_pad ,
		_w359_,
		_w373_
	);
	LUT2 #(
		.INIT('h1)
	) name227 (
		_w370_,
		_w372_,
		_w374_
	);
	LUT2 #(
		.INIT('h4)
	) name228 (
		_w340_,
		_w374_,
		_w375_
	);
	LUT2 #(
		.INIT('h4)
	) name229 (
		_w373_,
		_w375_,
		_w376_
	);
	LUT2 #(
		.INIT('h8)
	) name230 (
		_w365_,
		_w376_,
		_w377_
	);
	LUT2 #(
		.INIT('h4)
	) name231 (
		_w333_,
		_w377_,
		_w378_
	);
	LUT2 #(
		.INIT('h4)
	) name232 (
		_w274_,
		_w378_,
		_w379_
	);
	LUT2 #(
		.INIT('h4)
	) name233 (
		\g197_reg/NET0131 ,
		\g683_reg/NET0131 ,
		_w380_
	);
	LUT2 #(
		.INIT('h4)
	) name234 (
		\g211_reg/NET0131 ,
		_w221_,
		_w381_
	);
	LUT2 #(
		.INIT('h2)
	) name235 (
		\g210_reg/NET0131 ,
		_w381_,
		_w382_
	);
	LUT2 #(
		.INIT('h8)
	) name236 (
		_w268_,
		_w382_,
		_w383_
	);
	LUT2 #(
		.INIT('h2)
	) name237 (
		_w261_,
		_w383_,
		_w384_
	);
	LUT2 #(
		.INIT('h4)
	) name238 (
		_w263_,
		_w384_,
		_w385_
	);
	LUT2 #(
		.INIT('h2)
	) name239 (
		\g197_reg/NET0131 ,
		_w385_,
		_w386_
	);
	LUT2 #(
		.INIT('h1)
	) name240 (
		_w380_,
		_w386_,
		_w387_
	);
	LUT2 #(
		.INIT('h2)
	) name241 (
		_w208_,
		_w387_,
		_w388_
	);
	LUT2 #(
		.INIT('h1)
	) name242 (
		\g283_reg/NET0131 ,
		_w283_,
		_w389_
	);
	LUT2 #(
		.INIT('h4)
	) name243 (
		_w313_,
		_w389_,
		_w390_
	);
	LUT2 #(
		.INIT('h2)
	) name244 (
		\g282_reg/NET0131 ,
		_w390_,
		_w391_
	);
	LUT2 #(
		.INIT('h2)
	) name245 (
		_w324_,
		_w391_,
		_w392_
	);
	LUT2 #(
		.INIT('h1)
	) name246 (
		_w325_,
		_w392_,
		_w393_
	);
	LUT2 #(
		.INIT('h1)
	) name247 (
		\g282_reg/NET0131 ,
		\g283_reg/NET0131 ,
		_w394_
	);
	LUT2 #(
		.INIT('h4)
	) name248 (
		\g478_reg/NET0131 ,
		_w394_,
		_w395_
	);
	LUT2 #(
		.INIT('h4)
	) name249 (
		_w310_,
		_w395_,
		_w396_
	);
	LUT2 #(
		.INIT('h4)
	) name250 (
		\g282_reg/NET0131 ,
		\g283_reg/NET0131 ,
		_w397_
	);
	LUT2 #(
		.INIT('h8)
	) name251 (
		_w280_,
		_w397_,
		_w398_
	);
	LUT2 #(
		.INIT('h1)
	) name252 (
		_w396_,
		_w398_,
		_w399_
	);
	LUT2 #(
		.INIT('h4)
	) name253 (
		_w393_,
		_w399_,
		_w400_
	);
	LUT2 #(
		.INIT('h2)
	) name254 (
		\g269_reg/NET0131 ,
		_w400_,
		_w401_
	);
	LUT2 #(
		.INIT('h4)
	) name255 (
		\g269_reg/NET0131 ,
		\g683_reg/NET0131 ,
		_w402_
	);
	LUT2 #(
		.INIT('h1)
	) name256 (
		_w401_,
		_w402_,
		_w403_
	);
	LUT2 #(
		.INIT('h2)
	) name257 (
		_w275_,
		_w403_,
		_w404_
	);
	LUT2 #(
		.INIT('h2)
	) name258 (
		\g683_reg/NET0131 ,
		_w339_,
		_w405_
	);
	LUT2 #(
		.INIT('h8)
	) name259 (
		\g426_reg/NET0131 ,
		_w371_,
		_w406_
	);
	LUT2 #(
		.INIT('h8)
	) name260 (
		\g437_reg/NET0131 ,
		_w369_,
		_w407_
	);
	LUT2 #(
		.INIT('h8)
	) name261 (
		\g558_pad ,
		_w359_,
		_w408_
	);
	LUT2 #(
		.INIT('h1)
	) name262 (
		_w406_,
		_w407_,
		_w409_
	);
	LUT2 #(
		.INIT('h4)
	) name263 (
		_w405_,
		_w409_,
		_w410_
	);
	LUT2 #(
		.INIT('h4)
	) name264 (
		_w408_,
		_w410_,
		_w411_
	);
	LUT2 #(
		.INIT('h8)
	) name265 (
		_w365_,
		_w411_,
		_w412_
	);
	LUT2 #(
		.INIT('h4)
	) name266 (
		_w404_,
		_w412_,
		_w413_
	);
	LUT2 #(
		.INIT('h4)
	) name267 (
		_w388_,
		_w413_,
		_w414_
	);
	LUT2 #(
		.INIT('h8)
	) name268 (
		\g567_pad ,
		\g598_reg/NET0131 ,
		_w415_
	);
	LUT2 #(
		.INIT('h8)
	) name269 (
		\g634_reg/NET0131 ,
		_w415_,
		_w416_
	);
	LUT2 #(
		.INIT('h8)
	) name270 (
		\g642_reg/NET0131 ,
		_w416_,
		_w417_
	);
	LUT2 #(
		.INIT('h8)
	) name271 (
		\g606_reg/NET0131 ,
		_w417_,
		_w418_
	);
	LUT2 #(
		.INIT('h8)
	) name272 (
		\g646_reg/NET0131 ,
		_w418_,
		_w419_
	);
	LUT2 #(
		.INIT('h8)
	) name273 (
		\g650_reg/NET0131 ,
		_w419_,
		_w420_
	);
	LUT2 #(
		.INIT('h8)
	) name274 (
		\g654_reg/NET0131 ,
		_w420_,
		_w421_
	);
	LUT2 #(
		.INIT('h1)
	) name275 (
		\g571_reg/NET0131 ,
		_w421_,
		_w422_
	);
	LUT2 #(
		.INIT('h8)
	) name276 (
		\g571_reg/NET0131 ,
		_w421_,
		_w423_
	);
	LUT2 #(
		.INIT('h2)
	) name277 (
		\g638_reg/NET0131 ,
		_w422_,
		_w424_
	);
	LUT2 #(
		.INIT('h4)
	) name278 (
		_w423_,
		_w424_,
		_w425_
	);
	LUT2 #(
		.INIT('h4)
	) name279 (
		\g269_reg/NET0131 ,
		\g679_reg/NET0131 ,
		_w426_
	);
	LUT2 #(
		.INIT('h1)
	) name280 (
		_w280_,
		_w395_,
		_w427_
	);
	LUT2 #(
		.INIT('h8)
	) name281 (
		\g269_reg/NET0131 ,
		_w427_,
		_w428_
	);
	LUT2 #(
		.INIT('h1)
	) name282 (
		\g278_reg/NET0131 ,
		_w276_,
		_w429_
	);
	LUT2 #(
		.INIT('h1)
	) name283 (
		_w277_,
		_w429_,
		_w430_
	);
	LUT2 #(
		.INIT('h8)
	) name284 (
		_w428_,
		_w430_,
		_w431_
	);
	LUT2 #(
		.INIT('h1)
	) name285 (
		_w426_,
		_w431_,
		_w432_
	);
	LUT2 #(
		.INIT('h2)
	) name286 (
		_w275_,
		_w432_,
		_w433_
	);
	LUT2 #(
		.INIT('h8)
	) name287 (
		\g410_reg/NET0131 ,
		_w371_,
		_w434_
	);
	LUT2 #(
		.INIT('h8)
	) name288 (
		\g681_reg/NET0131 ,
		_w342_,
		_w435_
	);
	LUT2 #(
		.INIT('h8)
	) name289 (
		_w366_,
		_w435_,
		_w436_
	);
	LUT2 #(
		.INIT('h8)
	) name290 (
		\g551_reg/NET0131 ,
		_w436_,
		_w437_
	);
	LUT2 #(
		.INIT('h4)
	) name291 (
		\g683_reg/NET0131 ,
		_w354_,
		_w438_
	);
	LUT2 #(
		.INIT('h8)
	) name292 (
		_w203_,
		_w438_,
		_w439_
	);
	LUT2 #(
		.INIT('h8)
	) name293 (
		\g293_reg/NET0131 ,
		_w439_,
		_w440_
	);
	LUT2 #(
		.INIT('h8)
	) name294 (
		\g453_reg/NET0131 ,
		_w369_,
		_w441_
	);
	LUT2 #(
		.INIT('h4)
	) name295 (
		\g677_reg/NET0131 ,
		_w346_,
		_w442_
	);
	LUT2 #(
		.INIT('h8)
	) name296 (
		\g536_reg/NET0131 ,
		_w442_,
		_w443_
	);
	LUT2 #(
		.INIT('h8)
	) name297 (
		\g508_reg/NET0131 ,
		_w347_,
		_w444_
	);
	LUT2 #(
		.INIT('h4)
	) name298 (
		\g197_reg/NET0131 ,
		\g679_reg/NET0131 ,
		_w445_
	);
	LUT2 #(
		.INIT('h2)
	) name299 (
		\g197_reg/NET0131 ,
		_w258_,
		_w446_
	);
	LUT2 #(
		.INIT('h1)
	) name300 (
		_w213_,
		_w257_,
		_w447_
	);
	LUT2 #(
		.INIT('h1)
	) name301 (
		_w213_,
		_w218_,
		_w448_
	);
	LUT2 #(
		.INIT('h1)
	) name302 (
		_w447_,
		_w448_,
		_w449_
	);
	LUT2 #(
		.INIT('h2)
	) name303 (
		_w446_,
		_w449_,
		_w450_
	);
	LUT2 #(
		.INIT('h1)
	) name304 (
		\g206_reg/NET0131 ,
		_w209_,
		_w451_
	);
	LUT2 #(
		.INIT('h1)
	) name305 (
		_w210_,
		_w451_,
		_w452_
	);
	LUT2 #(
		.INIT('h8)
	) name306 (
		_w450_,
		_w452_,
		_w453_
	);
	LUT2 #(
		.INIT('h1)
	) name307 (
		_w445_,
		_w453_,
		_w454_
	);
	LUT2 #(
		.INIT('h2)
	) name308 (
		_w208_,
		_w454_,
		_w455_
	);
	LUT2 #(
		.INIT('h8)
	) name309 (
		\g562_pad ,
		_w358_,
		_w456_
	);
	LUT2 #(
		.INIT('h2)
	) name310 (
		_w339_,
		_w456_,
		_w457_
	);
	LUT2 #(
		.INIT('h2)
	) name311 (
		\g679_reg/NET0131 ,
		_w457_,
		_w458_
	);
	LUT2 #(
		.INIT('h1)
	) name312 (
		_w434_,
		_w437_,
		_w459_
	);
	LUT2 #(
		.INIT('h1)
	) name313 (
		_w440_,
		_w441_,
		_w460_
	);
	LUT2 #(
		.INIT('h8)
	) name314 (
		_w459_,
		_w460_,
		_w461_
	);
	LUT2 #(
		.INIT('h1)
	) name315 (
		_w443_,
		_w444_,
		_w462_
	);
	LUT2 #(
		.INIT('h8)
	) name316 (
		_w461_,
		_w462_,
		_w463_
	);
	LUT2 #(
		.INIT('h1)
	) name317 (
		_w364_,
		_w458_,
		_w464_
	);
	LUT2 #(
		.INIT('h8)
	) name318 (
		_w463_,
		_w464_,
		_w465_
	);
	LUT2 #(
		.INIT('h4)
	) name319 (
		_w433_,
		_w465_,
		_w466_
	);
	LUT2 #(
		.INIT('h4)
	) name320 (
		_w455_,
		_w466_,
		_w467_
	);
	LUT2 #(
		.INIT('h4)
	) name321 (
		\g197_reg/NET0131 ,
		\g680_reg/NET0131 ,
		_w468_
	);
	LUT2 #(
		.INIT('h1)
	) name322 (
		\g207_reg/NET0131 ,
		_w210_,
		_w469_
	);
	LUT2 #(
		.INIT('h1)
	) name323 (
		_w211_,
		_w469_,
		_w470_
	);
	LUT2 #(
		.INIT('h1)
	) name324 (
		_w449_,
		_w470_,
		_w471_
	);
	LUT2 #(
		.INIT('h2)
	) name325 (
		_w446_,
		_w471_,
		_w472_
	);
	LUT2 #(
		.INIT('h1)
	) name326 (
		_w468_,
		_w472_,
		_w473_
	);
	LUT2 #(
		.INIT('h2)
	) name327 (
		_w208_,
		_w473_,
		_w474_
	);
	LUT2 #(
		.INIT('h4)
	) name328 (
		\g269_reg/NET0131 ,
		\g680_reg/NET0131 ,
		_w475_
	);
	LUT2 #(
		.INIT('h1)
	) name329 (
		\g279_reg/NET0131 ,
		_w277_,
		_w476_
	);
	LUT2 #(
		.INIT('h1)
	) name330 (
		_w278_,
		_w476_,
		_w477_
	);
	LUT2 #(
		.INIT('h8)
	) name331 (
		_w310_,
		_w395_,
		_w478_
	);
	LUT2 #(
		.INIT('h1)
	) name332 (
		_w280_,
		_w478_,
		_w479_
	);
	LUT2 #(
		.INIT('h4)
	) name333 (
		_w477_,
		_w479_,
		_w480_
	);
	LUT2 #(
		.INIT('h2)
	) name334 (
		\g269_reg/NET0131 ,
		_w396_,
		_w481_
	);
	LUT2 #(
		.INIT('h4)
	) name335 (
		_w480_,
		_w481_,
		_w482_
	);
	LUT2 #(
		.INIT('h1)
	) name336 (
		_w475_,
		_w482_,
		_w483_
	);
	LUT2 #(
		.INIT('h2)
	) name337 (
		_w275_,
		_w483_,
		_w484_
	);
	LUT2 #(
		.INIT('h8)
	) name338 (
		\g414_reg/NET0131 ,
		_w371_,
		_w485_
	);
	LUT2 #(
		.INIT('h8)
	) name339 (
		\g449_reg/NET0131 ,
		_w369_,
		_w486_
	);
	LUT2 #(
		.INIT('h8)
	) name340 (
		\g512_reg/NET0131 ,
		_w347_,
		_w487_
	);
	LUT2 #(
		.INIT('h2)
	) name341 (
		\g680_reg/NET0131 ,
		_w339_,
		_w488_
	);
	LUT2 #(
		.INIT('h8)
	) name342 (
		\g541_reg/NET0131 ,
		_w442_,
		_w489_
	);
	LUT2 #(
		.INIT('h8)
	) name343 (
		\g554_reg/NET0131 ,
		_w436_,
		_w490_
	);
	LUT2 #(
		.INIT('h8)
	) name344 (
		\g297_reg/NET0131 ,
		_w439_,
		_w491_
	);
	LUT2 #(
		.INIT('h8)
	) name345 (
		\g561_pad ,
		_w359_,
		_w492_
	);
	LUT2 #(
		.INIT('h1)
	) name346 (
		_w485_,
		_w486_,
		_w493_
	);
	LUT2 #(
		.INIT('h1)
	) name347 (
		_w490_,
		_w491_,
		_w494_
	);
	LUT2 #(
		.INIT('h8)
	) name348 (
		_w493_,
		_w494_,
		_w495_
	);
	LUT2 #(
		.INIT('h1)
	) name349 (
		_w487_,
		_w488_,
		_w496_
	);
	LUT2 #(
		.INIT('h1)
	) name350 (
		_w489_,
		_w492_,
		_w497_
	);
	LUT2 #(
		.INIT('h8)
	) name351 (
		_w496_,
		_w497_,
		_w498_
	);
	LUT2 #(
		.INIT('h4)
	) name352 (
		_w364_,
		_w495_,
		_w499_
	);
	LUT2 #(
		.INIT('h8)
	) name353 (
		_w498_,
		_w499_,
		_w500_
	);
	LUT2 #(
		.INIT('h4)
	) name354 (
		_w474_,
		_w500_,
		_w501_
	);
	LUT2 #(
		.INIT('h4)
	) name355 (
		_w484_,
		_w501_,
		_w502_
	);
	LUT2 #(
		.INIT('h4)
	) name356 (
		\g197_reg/NET0131 ,
		\g682_reg/NET0131 ,
		_w503_
	);
	LUT2 #(
		.INIT('h1)
	) name357 (
		\g209_reg/NET0131 ,
		_w212_,
		_w504_
	);
	LUT2 #(
		.INIT('h1)
	) name358 (
		_w213_,
		_w504_,
		_w505_
	);
	LUT2 #(
		.INIT('h1)
	) name359 (
		_w258_,
		_w505_,
		_w506_
	);
	LUT2 #(
		.INIT('h2)
	) name360 (
		\g197_reg/NET0131 ,
		_w449_,
		_w507_
	);
	LUT2 #(
		.INIT('h4)
	) name361 (
		_w506_,
		_w507_,
		_w508_
	);
	LUT2 #(
		.INIT('h1)
	) name362 (
		_w503_,
		_w508_,
		_w509_
	);
	LUT2 #(
		.INIT('h2)
	) name363 (
		_w208_,
		_w509_,
		_w510_
	);
	LUT2 #(
		.INIT('h1)
	) name364 (
		\g281_reg/NET0131 ,
		_w395_,
		_w511_
	);
	LUT2 #(
		.INIT('h4)
	) name365 (
		_w279_,
		_w511_,
		_w512_
	);
	LUT2 #(
		.INIT('h2)
	) name366 (
		_w479_,
		_w512_,
		_w513_
	);
	LUT2 #(
		.INIT('h2)
	) name367 (
		\g269_reg/NET0131 ,
		_w513_,
		_w514_
	);
	LUT2 #(
		.INIT('h1)
	) name368 (
		\g269_reg/NET0131 ,
		\g682_reg/NET0131 ,
		_w515_
	);
	LUT2 #(
		.INIT('h1)
	) name369 (
		_w514_,
		_w515_,
		_w516_
	);
	LUT2 #(
		.INIT('h8)
	) name370 (
		_w275_,
		_w516_,
		_w517_
	);
	LUT2 #(
		.INIT('h2)
	) name371 (
		\g682_reg/NET0131 ,
		_w339_,
		_w518_
	);
	LUT2 #(
		.INIT('h8)
	) name372 (
		\g422_reg/NET0131 ,
		_w371_,
		_w519_
	);
	LUT2 #(
		.INIT('h8)
	) name373 (
		\g441_reg/NET0131 ,
		_w369_,
		_w520_
	);
	LUT2 #(
		.INIT('h8)
	) name374 (
		\g559_pad ,
		_w359_,
		_w521_
	);
	LUT2 #(
		.INIT('h1)
	) name375 (
		_w519_,
		_w520_,
		_w522_
	);
	LUT2 #(
		.INIT('h4)
	) name376 (
		_w518_,
		_w522_,
		_w523_
	);
	LUT2 #(
		.INIT('h4)
	) name377 (
		_w521_,
		_w523_,
		_w524_
	);
	LUT2 #(
		.INIT('h4)
	) name378 (
		_w364_,
		_w524_,
		_w525_
	);
	LUT2 #(
		.INIT('h4)
	) name379 (
		_w510_,
		_w525_,
		_w526_
	);
	LUT2 #(
		.INIT('h4)
	) name380 (
		_w517_,
		_w526_,
		_w527_
	);
	LUT2 #(
		.INIT('h4)
	) name381 (
		\g269_reg/NET0131 ,
		\g678_reg/NET0131 ,
		_w528_
	);
	LUT2 #(
		.INIT('h1)
	) name382 (
		\g276_reg/NET0131 ,
		\g277_reg/NET0131 ,
		_w529_
	);
	LUT2 #(
		.INIT('h1)
	) name383 (
		_w276_,
		_w529_,
		_w530_
	);
	LUT2 #(
		.INIT('h8)
	) name384 (
		_w428_,
		_w530_,
		_w531_
	);
	LUT2 #(
		.INIT('h1)
	) name385 (
		_w528_,
		_w531_,
		_w532_
	);
	LUT2 #(
		.INIT('h2)
	) name386 (
		_w275_,
		_w532_,
		_w533_
	);
	LUT2 #(
		.INIT('h8)
	) name387 (
		\g548_reg/NET0131 ,
		_w436_,
		_w534_
	);
	LUT2 #(
		.INIT('h8)
	) name388 (
		\g457_reg/NET0131 ,
		_w369_,
		_w535_
	);
	LUT2 #(
		.INIT('h8)
	) name389 (
		\g406_reg/NET0131 ,
		_w371_,
		_w536_
	);
	LUT2 #(
		.INIT('h8)
	) name390 (
		\g465_reg/NET0131 ,
		_w442_,
		_w537_
	);
	LUT2 #(
		.INIT('h8)
	) name391 (
		\g563_pad ,
		_w359_,
		_w538_
	);
	LUT2 #(
		.INIT('h8)
	) name392 (
		\g504_reg/NET0131 ,
		_w347_,
		_w539_
	);
	LUT2 #(
		.INIT('h8)
	) name393 (
		\g672_reg/NET0131 ,
		_w353_,
		_w540_
	);
	LUT2 #(
		.INIT('h8)
	) name394 (
		\g269_reg/NET0131 ,
		_w439_,
		_w541_
	);
	LUT2 #(
		.INIT('h8)
	) name395 (
		_w349_,
		_w356_,
		_w542_
	);
	LUT2 #(
		.INIT('h8)
	) name396 (
		\g492_reg/NET0131 ,
		_w542_,
		_w543_
	);
	LUT2 #(
		.INIT('h4)
	) name397 (
		\g197_reg/NET0131 ,
		\g678_reg/NET0131 ,
		_w544_
	);
	LUT2 #(
		.INIT('h1)
	) name398 (
		\g204_reg/NET0131 ,
		\g205_reg/NET0131 ,
		_w545_
	);
	LUT2 #(
		.INIT('h1)
	) name399 (
		_w209_,
		_w545_,
		_w546_
	);
	LUT2 #(
		.INIT('h8)
	) name400 (
		_w450_,
		_w546_,
		_w547_
	);
	LUT2 #(
		.INIT('h1)
	) name401 (
		_w544_,
		_w547_,
		_w548_
	);
	LUT2 #(
		.INIT('h2)
	) name402 (
		_w208_,
		_w548_,
		_w549_
	);
	LUT2 #(
		.INIT('h4)
	) name403 (
		\g489_reg/NET0131 ,
		_w357_,
		_w550_
	);
	LUT2 #(
		.INIT('h2)
	) name404 (
		_w339_,
		_w550_,
		_w551_
	);
	LUT2 #(
		.INIT('h2)
	) name405 (
		\g678_reg/NET0131 ,
		_w551_,
		_w552_
	);
	LUT2 #(
		.INIT('h1)
	) name406 (
		_w534_,
		_w540_,
		_w553_
	);
	LUT2 #(
		.INIT('h1)
	) name407 (
		_w535_,
		_w536_,
		_w554_
	);
	LUT2 #(
		.INIT('h1)
	) name408 (
		_w541_,
		_w543_,
		_w555_
	);
	LUT2 #(
		.INIT('h8)
	) name409 (
		_w554_,
		_w555_,
		_w556_
	);
	LUT2 #(
		.INIT('h4)
	) name410 (
		_w537_,
		_w553_,
		_w557_
	);
	LUT2 #(
		.INIT('h1)
	) name411 (
		_w538_,
		_w539_,
		_w558_
	);
	LUT2 #(
		.INIT('h8)
	) name412 (
		_w557_,
		_w558_,
		_w559_
	);
	LUT2 #(
		.INIT('h4)
	) name413 (
		_w364_,
		_w556_,
		_w560_
	);
	LUT2 #(
		.INIT('h4)
	) name414 (
		_w552_,
		_w560_,
		_w561_
	);
	LUT2 #(
		.INIT('h4)
	) name415 (
		_w533_,
		_w559_,
		_w562_
	);
	LUT2 #(
		.INIT('h8)
	) name416 (
		_w561_,
		_w562_,
		_w563_
	);
	LUT2 #(
		.INIT('h4)
	) name417 (
		_w549_,
		_w563_,
		_w564_
	);
	LUT2 #(
		.INIT('h4)
	) name418 (
		\g269_reg/NET0131 ,
		\g677_reg/NET0131 ,
		_w565_
	);
	LUT2 #(
		.INIT('h4)
	) name419 (
		\g276_reg/NET0131 ,
		_w428_,
		_w566_
	);
	LUT2 #(
		.INIT('h1)
	) name420 (
		_w565_,
		_w566_,
		_w567_
	);
	LUT2 #(
		.INIT('h2)
	) name421 (
		_w275_,
		_w567_,
		_w568_
	);
	LUT2 #(
		.INIT('h4)
	) name422 (
		\g197_reg/NET0131 ,
		\g677_reg/NET0131 ,
		_w569_
	);
	LUT2 #(
		.INIT('h4)
	) name423 (
		\g204_reg/NET0131 ,
		_w450_,
		_w570_
	);
	LUT2 #(
		.INIT('h1)
	) name424 (
		_w569_,
		_w570_,
		_w571_
	);
	LUT2 #(
		.INIT('h2)
	) name425 (
		_w208_,
		_w571_,
		_w572_
	);
	LUT2 #(
		.INIT('h8)
	) name426 (
		\g669_reg/NET0131 ,
		_w353_,
		_w573_
	);
	LUT2 #(
		.INIT('h8)
	) name427 (
		\g545_reg/NET0131 ,
		_w436_,
		_w574_
	);
	LUT2 #(
		.INIT('h8)
	) name428 (
		\g402_reg/NET0131 ,
		_w371_,
		_w575_
	);
	LUT2 #(
		.INIT('h8)
	) name429 (
		\g496_reg/NET0131 ,
		_w542_,
		_w576_
	);
	LUT2 #(
		.INIT('h2)
	) name430 (
		\g677_reg/NET0131 ,
		_w339_,
		_w577_
	);
	LUT2 #(
		.INIT('h8)
	) name431 (
		\g4422_pad ,
		_w359_,
		_w578_
	);
	LUT2 #(
		.INIT('h8)
	) name432 (
		\g197_reg/NET0131 ,
		_w439_,
		_w579_
	);
	LUT2 #(
		.INIT('h1)
	) name433 (
		\g486_reg/NET0131 ,
		\g679_reg/NET0131 ,
		_w580_
	);
	LUT2 #(
		.INIT('h8)
	) name434 (
		_w358_,
		_w580_,
		_w581_
	);
	LUT2 #(
		.INIT('h8)
	) name435 (
		\g461_reg/NET0131 ,
		_w369_,
		_w582_
	);
	LUT2 #(
		.INIT('h1)
	) name436 (
		_w573_,
		_w574_,
		_w583_
	);
	LUT2 #(
		.INIT('h1)
	) name437 (
		_w575_,
		_w576_,
		_w584_
	);
	LUT2 #(
		.INIT('h1)
	) name438 (
		_w579_,
		_w581_,
		_w585_
	);
	LUT2 #(
		.INIT('h4)
	) name439 (
		_w582_,
		_w585_,
		_w586_
	);
	LUT2 #(
		.INIT('h8)
	) name440 (
		_w583_,
		_w584_,
		_w587_
	);
	LUT2 #(
		.INIT('h1)
	) name441 (
		_w348_,
		_w577_,
		_w588_
	);
	LUT2 #(
		.INIT('h4)
	) name442 (
		_w578_,
		_w588_,
		_w589_
	);
	LUT2 #(
		.INIT('h8)
	) name443 (
		_w586_,
		_w587_,
		_w590_
	);
	LUT2 #(
		.INIT('h4)
	) name444 (
		_w364_,
		_w590_,
		_w591_
	);
	LUT2 #(
		.INIT('h4)
	) name445 (
		_w568_,
		_w589_,
		_w592_
	);
	LUT2 #(
		.INIT('h8)
	) name446 (
		_w591_,
		_w592_,
		_w593_
	);
	LUT2 #(
		.INIT('h4)
	) name447 (
		_w572_,
		_w593_,
		_w594_
	);
	LUT2 #(
		.INIT('h4)
	) name448 (
		\g269_reg/NET0131 ,
		\g681_reg/NET0131 ,
		_w595_
	);
	LUT2 #(
		.INIT('h1)
	) name449 (
		\g280_reg/NET0131 ,
		_w278_,
		_w596_
	);
	LUT2 #(
		.INIT('h1)
	) name450 (
		_w279_,
		_w596_,
		_w597_
	);
	LUT2 #(
		.INIT('h2)
	) name451 (
		_w427_,
		_w597_,
		_w598_
	);
	LUT2 #(
		.INIT('h2)
	) name452 (
		\g269_reg/NET0131 ,
		_w598_,
		_w599_
	);
	LUT2 #(
		.INIT('h1)
	) name453 (
		_w595_,
		_w599_,
		_w600_
	);
	LUT2 #(
		.INIT('h2)
	) name454 (
		_w275_,
		_w600_,
		_w601_
	);
	LUT2 #(
		.INIT('h4)
	) name455 (
		\g197_reg/NET0131 ,
		\g681_reg/NET0131 ,
		_w602_
	);
	LUT2 #(
		.INIT('h1)
	) name456 (
		\g208_reg/NET0131 ,
		_w211_,
		_w603_
	);
	LUT2 #(
		.INIT('h1)
	) name457 (
		_w212_,
		_w603_,
		_w604_
	);
	LUT2 #(
		.INIT('h2)
	) name458 (
		_w447_,
		_w604_,
		_w605_
	);
	LUT2 #(
		.INIT('h2)
	) name459 (
		\g197_reg/NET0131 ,
		_w605_,
		_w606_
	);
	LUT2 #(
		.INIT('h1)
	) name460 (
		_w602_,
		_w606_,
		_w607_
	);
	LUT2 #(
		.INIT('h2)
	) name461 (
		_w208_,
		_w607_,
		_w608_
	);
	LUT2 #(
		.INIT('h8)
	) name462 (
		\g560_pad ,
		_w359_,
		_w609_
	);
	LUT2 #(
		.INIT('h8)
	) name463 (
		\g445_reg/NET0131 ,
		_w369_,
		_w610_
	);
	LUT2 #(
		.INIT('h2)
	) name464 (
		\g681_reg/NET0131 ,
		_w339_,
		_w611_
	);
	LUT2 #(
		.INIT('h8)
	) name465 (
		\g418_reg/NET0131 ,
		_w371_,
		_w612_
	);
	LUT2 #(
		.INIT('h1)
	) name466 (
		_w610_,
		_w612_,
		_w613_
	);
	LUT2 #(
		.INIT('h4)
	) name467 (
		_w609_,
		_w613_,
		_w614_
	);
	LUT2 #(
		.INIT('h4)
	) name468 (
		_w611_,
		_w614_,
		_w615_
	);
	LUT2 #(
		.INIT('h4)
	) name469 (
		_w364_,
		_w615_,
		_w616_
	);
	LUT2 #(
		.INIT('h1)
	) name470 (
		_w601_,
		_w608_,
		_w617_
	);
	LUT2 #(
		.INIT('h8)
	) name471 (
		_w616_,
		_w617_,
		_w618_
	);
	LUT2 #(
		.INIT('h1)
	) name472 (
		\g631_reg/NET0131 ,
		_w153_,
		_w619_
	);
	LUT2 #(
		.INIT('h2)
	) name473 (
		\g639_pad ,
		_w154_,
		_w620_
	);
	LUT2 #(
		.INIT('h4)
	) name474 (
		_w619_,
		_w620_,
		_w621_
	);
	LUT2 #(
		.INIT('h1)
	) name475 (
		\g654_reg/NET0131 ,
		_w420_,
		_w622_
	);
	LUT2 #(
		.INIT('h2)
	) name476 (
		\g638_reg/NET0131 ,
		_w421_,
		_w623_
	);
	LUT2 #(
		.INIT('h4)
	) name477 (
		_w622_,
		_w623_,
		_w624_
	);
	LUT2 #(
		.INIT('h1)
	) name478 (
		\g628_reg/NET0131 ,
		_w152_,
		_w625_
	);
	LUT2 #(
		.INIT('h2)
	) name479 (
		\g639_pad ,
		_w153_,
		_w626_
	);
	LUT2 #(
		.INIT('h4)
	) name480 (
		_w625_,
		_w626_,
		_w627_
	);
	LUT2 #(
		.INIT('h1)
	) name481 (
		_w270_,
		_w384_,
		_w628_
	);
	LUT2 #(
		.INIT('h1)
	) name482 (
		_w329_,
		_w400_,
		_w629_
	);
	LUT2 #(
		.INIT('h1)
	) name483 (
		\g650_reg/NET0131 ,
		_w419_,
		_w630_
	);
	LUT2 #(
		.INIT('h2)
	) name484 (
		\g638_reg/NET0131 ,
		_w420_,
		_w631_
	);
	LUT2 #(
		.INIT('h4)
	) name485 (
		_w630_,
		_w631_,
		_w632_
	);
	LUT2 #(
		.INIT('h2)
	) name486 (
		\g18_reg/NET0131 ,
		\g28_reg/NET0131 ,
		_w633_
	);
	LUT2 #(
		.INIT('h4)
	) name487 (
		\g18_reg/NET0131 ,
		\g28_reg/NET0131 ,
		_w634_
	);
	LUT2 #(
		.INIT('h1)
	) name488 (
		_w633_,
		_w634_,
		_w635_
	);
	LUT2 #(
		.INIT('h1)
	) name489 (
		\g10_reg/NET0131 ,
		\g1_reg/NET0131 ,
		_w636_
	);
	LUT2 #(
		.INIT('h8)
	) name490 (
		\g10_reg/NET0131 ,
		\g1_reg/NET0131 ,
		_w637_
	);
	LUT2 #(
		.INIT('h1)
	) name491 (
		_w636_,
		_w637_,
		_w638_
	);
	LUT2 #(
		.INIT('h2)
	) name492 (
		_w635_,
		_w638_,
		_w639_
	);
	LUT2 #(
		.INIT('h4)
	) name493 (
		_w635_,
		_w638_,
		_w640_
	);
	LUT2 #(
		.INIT('h1)
	) name494 (
		_w639_,
		_w640_,
		_w641_
	);
	LUT2 #(
		.INIT('h1)
	) name495 (
		\g14_reg/NET0131 ,
		\g48_reg/NET0131 ,
		_w642_
	);
	LUT2 #(
		.INIT('h8)
	) name496 (
		\g14_reg/NET0131 ,
		\g48_reg/NET0131 ,
		_w643_
	);
	LUT2 #(
		.INIT('h1)
	) name497 (
		_w642_,
		_w643_,
		_w644_
	);
	LUT2 #(
		.INIT('h8)
	) name498 (
		\g2_reg/NET0131 ,
		_w644_,
		_w645_
	);
	LUT2 #(
		.INIT('h1)
	) name499 (
		\g2_reg/NET0131 ,
		_w644_,
		_w646_
	);
	LUT2 #(
		.INIT('h1)
	) name500 (
		_w645_,
		_w646_,
		_w647_
	);
	LUT2 #(
		.INIT('h2)
	) name501 (
		\g24_reg/NET0131 ,
		\g6_reg/NET0131 ,
		_w648_
	);
	LUT2 #(
		.INIT('h4)
	) name502 (
		\g24_reg/NET0131 ,
		\g6_reg/NET0131 ,
		_w649_
	);
	LUT2 #(
		.INIT('h1)
	) name503 (
		_w648_,
		_w649_,
		_w650_
	);
	LUT2 #(
		.INIT('h2)
	) name504 (
		_w647_,
		_w650_,
		_w651_
	);
	LUT2 #(
		.INIT('h4)
	) name505 (
		_w647_,
		_w650_,
		_w652_
	);
	LUT2 #(
		.INIT('h1)
	) name506 (
		_w651_,
		_w652_,
		_w653_
	);
	LUT2 #(
		.INIT('h8)
	) name507 (
		_w641_,
		_w653_,
		_w654_
	);
	LUT2 #(
		.INIT('h1)
	) name508 (
		_w641_,
		_w653_,
		_w655_
	);
	LUT2 #(
		.INIT('h1)
	) name509 (
		_w654_,
		_w655_,
		_w656_
	);
	LUT2 #(
		.INIT('h1)
	) name510 (
		\g4110_pad ,
		_w656_,
		_w657_
	);
	LUT2 #(
		.INIT('h2)
	) name511 (
		\g676_reg/NET0131 ,
		_w657_,
		_w658_
	);
	LUT2 #(
		.INIT('h4)
	) name512 (
		\g4110_pad ,
		_w200_,
		_w659_
	);
	LUT2 #(
		.INIT('h8)
	) name513 (
		_w658_,
		_w659_,
		_w660_
	);
	LUT2 #(
		.INIT('h8)
	) name514 (
		_w345_,
		_w660_,
		_w661_
	);
	LUT2 #(
		.INIT('h4)
	) name515 (
		\g677_reg/NET0131 ,
		_w661_,
		_w662_
	);
	LUT2 #(
		.INIT('h8)
	) name516 (
		\g679_reg/NET0131 ,
		_w662_,
		_w663_
	);
	LUT2 #(
		.INIT('h1)
	) name517 (
		\g218_reg/NET0131 ,
		\g504_reg/NET0131 ,
		_w664_
	);
	LUT2 #(
		.INIT('h8)
	) name518 (
		\g218_reg/NET0131 ,
		\g504_reg/NET0131 ,
		_w665_
	);
	LUT2 #(
		.INIT('h1)
	) name519 (
		_w664_,
		_w665_,
		_w666_
	);
	LUT2 #(
		.INIT('h1)
	) name520 (
		\g230_reg/NET0131 ,
		\g512_reg/NET0131 ,
		_w667_
	);
	LUT2 #(
		.INIT('h8)
	) name521 (
		\g230_reg/NET0131 ,
		\g512_reg/NET0131 ,
		_w668_
	);
	LUT2 #(
		.INIT('h1)
	) name522 (
		_w667_,
		_w668_,
		_w669_
	);
	LUT2 #(
		.INIT('h1)
	) name523 (
		\g224_reg/NET0131 ,
		\g508_reg/NET0131 ,
		_w670_
	);
	LUT2 #(
		.INIT('h8)
	) name524 (
		\g224_reg/NET0131 ,
		\g508_reg/NET0131 ,
		_w671_
	);
	LUT2 #(
		.INIT('h1)
	) name525 (
		_w670_,
		_w671_,
		_w672_
	);
	LUT2 #(
		.INIT('h1)
	) name526 (
		\g212_reg/NET0131 ,
		\g248_reg/NET0131 ,
		_w673_
	);
	LUT2 #(
		.INIT('h1)
	) name527 (
		\g254_reg/NET0131 ,
		\g500_reg/NET0131 ,
		_w674_
	);
	LUT2 #(
		.INIT('h8)
	) name528 (
		_w673_,
		_w674_,
		_w675_
	);
	LUT2 #(
		.INIT('h8)
	) name529 (
		\g212_reg/NET0131 ,
		\g248_reg/NET0131 ,
		_w676_
	);
	LUT2 #(
		.INIT('h8)
	) name530 (
		\g254_reg/NET0131 ,
		\g500_reg/NET0131 ,
		_w677_
	);
	LUT2 #(
		.INIT('h8)
	) name531 (
		_w676_,
		_w677_,
		_w678_
	);
	LUT2 #(
		.INIT('h1)
	) name532 (
		_w675_,
		_w678_,
		_w679_
	);
	LUT2 #(
		.INIT('h1)
	) name533 (
		\g236_reg/NET0131 ,
		\g242_reg/NET0131 ,
		_w680_
	);
	LUT2 #(
		.INIT('h4)
	) name534 (
		\g260_reg/NET0131 ,
		_w680_,
		_w681_
	);
	LUT2 #(
		.INIT('h4)
	) name535 (
		_w666_,
		_w681_,
		_w682_
	);
	LUT2 #(
		.INIT('h1)
	) name536 (
		_w669_,
		_w672_,
		_w683_
	);
	LUT2 #(
		.INIT('h8)
	) name537 (
		_w682_,
		_w683_,
		_w684_
	);
	LUT2 #(
		.INIT('h4)
	) name538 (
		_w679_,
		_w684_,
		_w685_
	);
	LUT2 #(
		.INIT('h1)
	) name539 (
		\g465_reg/NET0131 ,
		_w217_,
		_w686_
	);
	LUT2 #(
		.INIT('h2)
	) name540 (
		\g465_reg/NET0131 ,
		_w309_,
		_w687_
	);
	LUT2 #(
		.INIT('h2)
	) name541 (
		_w685_,
		_w686_,
		_w688_
	);
	LUT2 #(
		.INIT('h4)
	) name542 (
		_w687_,
		_w688_,
		_w689_
	);
	LUT2 #(
		.INIT('h2)
	) name543 (
		\g536_reg/NET0131 ,
		_w689_,
		_w690_
	);
	LUT2 #(
		.INIT('h4)
	) name544 (
		_w662_,
		_w690_,
		_w691_
	);
	LUT2 #(
		.INIT('h1)
	) name545 (
		_w663_,
		_w691_,
		_w692_
	);
	LUT2 #(
		.INIT('h1)
	) name546 (
		\g625_reg/NET0131 ,
		_w151_,
		_w693_
	);
	LUT2 #(
		.INIT('h2)
	) name547 (
		\g639_pad ,
		_w152_,
		_w694_
	);
	LUT2 #(
		.INIT('h4)
	) name548 (
		_w693_,
		_w694_,
		_w695_
	);
	LUT2 #(
		.INIT('h1)
	) name549 (
		\g646_reg/NET0131 ,
		_w418_,
		_w696_
	);
	LUT2 #(
		.INIT('h2)
	) name550 (
		\g638_reg/NET0131 ,
		_w419_,
		_w697_
	);
	LUT2 #(
		.INIT('h4)
	) name551 (
		_w696_,
		_w697_,
		_w698_
	);
	LUT2 #(
		.INIT('h1)
	) name552 (
		\g492_reg/NET0131 ,
		_w317_,
		_w699_
	);
	LUT2 #(
		.INIT('h1)
	) name553 (
		\g496_reg/NET0131 ,
		_w249_,
		_w700_
	);
	LUT2 #(
		.INIT('h8)
	) name554 (
		\g677_reg/NET0131 ,
		_w661_,
		_w701_
	);
	LUT2 #(
		.INIT('h1)
	) name555 (
		\g622_reg/NET0131 ,
		_w150_,
		_w702_
	);
	LUT2 #(
		.INIT('h2)
	) name556 (
		\g639_pad ,
		_w151_,
		_w703_
	);
	LUT2 #(
		.INIT('h4)
	) name557 (
		_w702_,
		_w703_,
		_w704_
	);
	LUT2 #(
		.INIT('h8)
	) name558 (
		_w438_,
		_w660_,
		_w705_
	);
	LUT2 #(
		.INIT('h1)
	) name559 (
		\g606_reg/NET0131 ,
		_w417_,
		_w706_
	);
	LUT2 #(
		.INIT('h2)
	) name560 (
		\g638_reg/NET0131 ,
		_w418_,
		_w707_
	);
	LUT2 #(
		.INIT('h4)
	) name561 (
		_w706_,
		_w707_,
		_w708_
	);
	LUT2 #(
		.INIT('h2)
	) name562 (
		\g4101_pad ,
		\g4105_pad ,
		_w709_
	);
	LUT2 #(
		.INIT('h4)
	) name563 (
		\g4101_pad ,
		\g4105_pad ,
		_w710_
	);
	LUT2 #(
		.INIT('h1)
	) name564 (
		_w709_,
		_w710_,
		_w711_
	);
	LUT2 #(
		.INIT('h8)
	) name565 (
		\g4103_pad ,
		_w711_,
		_w712_
	);
	LUT2 #(
		.INIT('h1)
	) name566 (
		\g4103_pad ,
		_w711_,
		_w713_
	);
	LUT2 #(
		.INIT('h1)
	) name567 (
		_w712_,
		_w713_,
		_w714_
	);
	LUT2 #(
		.INIT('h2)
	) name568 (
		\g4099_pad ,
		_w714_,
		_w715_
	);
	LUT2 #(
		.INIT('h4)
	) name569 (
		\g4099_pad ,
		_w714_,
		_w716_
	);
	LUT2 #(
		.INIT('h1)
	) name570 (
		_w715_,
		_w716_,
		_w717_
	);
	LUT2 #(
		.INIT('h1)
	) name571 (
		\g4100_pad ,
		\g4102_pad ,
		_w718_
	);
	LUT2 #(
		.INIT('h8)
	) name572 (
		\g4100_pad ,
		\g4102_pad ,
		_w719_
	);
	LUT2 #(
		.INIT('h1)
	) name573 (
		_w718_,
		_w719_,
		_w720_
	);
	LUT2 #(
		.INIT('h4)
	) name574 (
		_w656_,
		_w720_,
		_w721_
	);
	LUT2 #(
		.INIT('h2)
	) name575 (
		_w656_,
		_w720_,
		_w722_
	);
	LUT2 #(
		.INIT('h1)
	) name576 (
		_w721_,
		_w722_,
		_w723_
	);
	LUT2 #(
		.INIT('h8)
	) name577 (
		_w717_,
		_w723_,
		_w724_
	);
	LUT2 #(
		.INIT('h1)
	) name578 (
		_w717_,
		_w723_,
		_w725_
	);
	LUT2 #(
		.INIT('h1)
	) name579 (
		_w724_,
		_w725_,
		_w726_
	);
	LUT2 #(
		.INIT('h4)
	) name580 (
		\g4104_pad ,
		_w726_,
		_w727_
	);
	LUT2 #(
		.INIT('h1)
	) name581 (
		\g669_reg/NET0131 ,
		_w727_,
		_w728_
	);
	LUT2 #(
		.INIT('h1)
	) name582 (
		\g619_reg/NET0131 ,
		_w149_,
		_w729_
	);
	LUT2 #(
		.INIT('h2)
	) name583 (
		\g639_pad ,
		_w150_,
		_w730_
	);
	LUT2 #(
		.INIT('h4)
	) name584 (
		_w729_,
		_w730_,
		_w731_
	);
	LUT2 #(
		.INIT('h1)
	) name585 (
		\g642_reg/NET0131 ,
		_w416_,
		_w732_
	);
	LUT2 #(
		.INIT('h2)
	) name586 (
		\g638_reg/NET0131 ,
		_w417_,
		_w733_
	);
	LUT2 #(
		.INIT('h4)
	) name587 (
		_w732_,
		_w733_,
		_w734_
	);
	LUT2 #(
		.INIT('h4)
	) name588 (
		\g4104_pad ,
		_w657_,
		_w735_
	);
	LUT2 #(
		.INIT('h1)
	) name589 (
		\g672_reg/NET0131 ,
		_w735_,
		_w736_
	);
	LUT2 #(
		.INIT('h4)
	) name590 (
		\g536_reg/NET0131 ,
		_w685_,
		_w737_
	);
	LUT2 #(
		.INIT('h4)
	) name591 (
		\g541_reg/NET0131 ,
		_w737_,
		_w738_
	);
	LUT2 #(
		.INIT('h4)
	) name592 (
		\g590_reg/NET0131 ,
		\g594_reg/NET0131 ,
		_w739_
	);
	LUT2 #(
		.INIT('h2)
	) name593 (
		\g590_reg/NET0131 ,
		\g594_reg/NET0131 ,
		_w740_
	);
	LUT2 #(
		.INIT('h4)
	) name594 (
		\g578_reg/NET0131 ,
		\g682_reg/NET0131 ,
		_w741_
	);
	LUT2 #(
		.INIT('h8)
	) name595 (
		\g578_reg/NET0131 ,
		\g681_reg/NET0131 ,
		_w742_
	);
	LUT2 #(
		.INIT('h2)
	) name596 (
		\g582_reg/NET0131 ,
		_w741_,
		_w743_
	);
	LUT2 #(
		.INIT('h4)
	) name597 (
		_w742_,
		_w743_,
		_w744_
	);
	LUT2 #(
		.INIT('h4)
	) name598 (
		\g578_reg/NET0131 ,
		\g684_reg/NET0131 ,
		_w745_
	);
	LUT2 #(
		.INIT('h8)
	) name599 (
		\g578_reg/NET0131 ,
		\g683_reg/NET0131 ,
		_w746_
	);
	LUT2 #(
		.INIT('h1)
	) name600 (
		\g582_reg/NET0131 ,
		_w745_,
		_w747_
	);
	LUT2 #(
		.INIT('h4)
	) name601 (
		_w746_,
		_w747_,
		_w748_
	);
	LUT2 #(
		.INIT('h1)
	) name602 (
		_w744_,
		_w748_,
		_w749_
	);
	LUT2 #(
		.INIT('h1)
	) name603 (
		\g586_reg/NET0131 ,
		_w749_,
		_w750_
	);
	LUT2 #(
		.INIT('h4)
	) name604 (
		\g578_reg/NET0131 ,
		\g680_reg/NET0131 ,
		_w751_
	);
	LUT2 #(
		.INIT('h8)
	) name605 (
		\g578_reg/NET0131 ,
		\g679_reg/NET0131 ,
		_w752_
	);
	LUT2 #(
		.INIT('h1)
	) name606 (
		\g582_reg/NET0131 ,
		_w751_,
		_w753_
	);
	LUT2 #(
		.INIT('h4)
	) name607 (
		_w752_,
		_w753_,
		_w754_
	);
	LUT2 #(
		.INIT('h4)
	) name608 (
		\g578_reg/NET0131 ,
		\g678_reg/NET0131 ,
		_w755_
	);
	LUT2 #(
		.INIT('h8)
	) name609 (
		\g578_reg/NET0131 ,
		\g677_reg/NET0131 ,
		_w756_
	);
	LUT2 #(
		.INIT('h2)
	) name610 (
		\g582_reg/NET0131 ,
		_w755_,
		_w757_
	);
	LUT2 #(
		.INIT('h4)
	) name611 (
		_w756_,
		_w757_,
		_w758_
	);
	LUT2 #(
		.INIT('h1)
	) name612 (
		_w754_,
		_w758_,
		_w759_
	);
	LUT2 #(
		.INIT('h2)
	) name613 (
		\g586_reg/NET0131 ,
		_w759_,
		_w760_
	);
	LUT2 #(
		.INIT('h1)
	) name614 (
		_w750_,
		_w760_,
		_w761_
	);
	LUT2 #(
		.INIT('h1)
	) name615 (
		_w739_,
		_w740_,
		_w762_
	);
	LUT2 #(
		.INIT('h4)
	) name616 (
		_w761_,
		_w762_,
		_w763_
	);
	LUT2 #(
		.INIT('h8)
	) name617 (
		\g574_reg/NET0131 ,
		\g578_reg/NET0131 ,
		_w764_
	);
	LUT2 #(
		.INIT('h8)
	) name618 (
		\g582_reg/NET0131 ,
		\g586_reg/NET0131 ,
		_w765_
	);
	LUT2 #(
		.INIT('h8)
	) name619 (
		_w764_,
		_w765_,
		_w766_
	);
	LUT2 #(
		.INIT('h8)
	) name620 (
		_w739_,
		_w766_,
		_w767_
	);
	LUT2 #(
		.INIT('h1)
	) name621 (
		_w763_,
		_w767_,
		_w768_
	);
	LUT2 #(
		.INIT('h1)
	) name622 (
		\g616_reg/NET0131 ,
		_w148_,
		_w769_
	);
	LUT2 #(
		.INIT('h2)
	) name623 (
		\g639_pad ,
		_w149_,
		_w770_
	);
	LUT2 #(
		.INIT('h4)
	) name624 (
		_w769_,
		_w770_,
		_w771_
	);
	LUT2 #(
		.INIT('h1)
	) name625 (
		\g634_reg/NET0131 ,
		_w415_,
		_w772_
	);
	LUT2 #(
		.INIT('h2)
	) name626 (
		\g638_reg/NET0131 ,
		_w416_,
		_w773_
	);
	LUT2 #(
		.INIT('h4)
	) name627 (
		_w772_,
		_w773_,
		_w774_
	);
	LUT2 #(
		.INIT('h1)
	) name628 (
		\g613_reg/NET0131 ,
		_w147_,
		_w775_
	);
	LUT2 #(
		.INIT('h1)
	) name629 (
		_w148_,
		_w775_,
		_w776_
	);
	LUT2 #(
		.INIT('h2)
	) name630 (
		\g639_pad ,
		_w776_,
		_w777_
	);
	LUT2 #(
		.INIT('h8)
	) name631 (
		\g465_reg/NET0131 ,
		\g478_reg/NET0131 ,
		_w778_
	);
	LUT2 #(
		.INIT('h4)
	) name632 (
		\g465_reg/NET0131 ,
		\g471_reg/NET0131 ,
		_w779_
	);
	LUT2 #(
		.INIT('h1)
	) name633 (
		_w778_,
		_w779_,
		_w780_
	);
	LUT2 #(
		.INIT('h1)
	) name634 (
		\g567_pad ,
		\g598_reg/NET0131 ,
		_w781_
	);
	LUT2 #(
		.INIT('h2)
	) name635 (
		\g638_reg/NET0131 ,
		_w415_,
		_w782_
	);
	LUT2 #(
		.INIT('h4)
	) name636 (
		_w781_,
		_w782_,
		_w783_
	);
	LUT2 #(
		.INIT('h1)
	) name637 (
		\g602_reg/NET0131 ,
		\g610_reg/NET0131 ,
		_w784_
	);
	LUT2 #(
		.INIT('h2)
	) name638 (
		\g639_pad ,
		_w147_,
		_w785_
	);
	LUT2 #(
		.INIT('h4)
	) name639 (
		_w784_,
		_w785_,
		_w786_
	);
	LUT2 #(
		.INIT('h4)
	) name640 (
		\g266_reg/NET0131 ,
		\g4108_pad ,
		_w787_
	);
	LUT2 #(
		.INIT('h4)
	) name641 (
		\g602_reg/NET0131 ,
		\g639_pad ,
		_w788_
	);
	LUT2 #(
		.INIT('h4)
	) name642 (
		\g680_reg/NET0131 ,
		_w662_,
		_w789_
	);
	LUT2 #(
		.INIT('h1)
	) name643 (
		\g465_reg/NET0131 ,
		_w213_,
		_w790_
	);
	LUT2 #(
		.INIT('h2)
	) name644 (
		\g465_reg/NET0131 ,
		_w280_,
		_w791_
	);
	LUT2 #(
		.INIT('h2)
	) name645 (
		_w737_,
		_w790_,
		_w792_
	);
	LUT2 #(
		.INIT('h4)
	) name646 (
		_w791_,
		_w792_,
		_w793_
	);
	LUT2 #(
		.INIT('h1)
	) name647 (
		\g541_reg/NET0131 ,
		_w793_,
		_w794_
	);
	LUT2 #(
		.INIT('h4)
	) name648 (
		_w662_,
		_w794_,
		_w795_
	);
	LUT2 #(
		.INIT('h1)
	) name649 (
		_w789_,
		_w795_,
		_w796_
	);
	LUT2 #(
		.INIT('h4)
	) name650 (
		\g102_pad ,
		\g89_pad ,
		_w797_
	);
	LUT2 #(
		.INIT('h8)
	) name651 (
		\g567_pad ,
		\g638_reg/NET0131 ,
		_w798_
	);
	LUT2 #(
		.INIT('h4)
	) name652 (
		\g489_reg/NET0131 ,
		\g492_reg/NET0131 ,
		_w799_
	);
	LUT2 #(
		.INIT('h4)
	) name653 (
		\g486_reg/NET0131 ,
		\g496_reg/NET0131 ,
		_w800_
	);
	LUT2 #(
		.INIT('h1)
	) name654 (
		_w799_,
		_w800_,
		_w801_
	);
	LUT2 #(
		.INIT('h4)
	) name655 (
		\g4104_pad ,
		\g675_reg/NET0131 ,
		_w802_
	);
	LUT2 #(
		.INIT('h8)
	) name656 (
		_w658_,
		_w802_,
		_w803_
	);
	LUT2 #(
		.INIT('h8)
	) name657 (
		\g4110_pad ,
		_w803_,
		_w804_
	);
	LUT2 #(
		.INIT('h4)
	) name658 (
		_w199_,
		_w804_,
		_w805_
	);
	LUT2 #(
		.INIT('h4)
	) name659 (
		\g25_reg/NET0131 ,
		_w804_,
		_w806_
	);
	LUT2 #(
		.INIT('h4)
	) name660 (
		\g29_reg/NET0131 ,
		_w804_,
		_w807_
	);
	LUT2 #(
		.INIT('h4)
	) name661 (
		\g3_reg/NET0131 ,
		_w804_,
		_w808_
	);
	LUT2 #(
		.INIT('h4)
	) name662 (
		\g33_reg/NET0131 ,
		_w804_,
		_w809_
	);
	LUT2 #(
		.INIT('h4)
	) name663 (
		\g7_reg/NET0131 ,
		_w804_,
		_w810_
	);
	LUT2 #(
		.INIT('h4)
	) name664 (
		\g11_reg/NET0131 ,
		_w804_,
		_w811_
	);
	LUT2 #(
		.INIT('h4)
	) name665 (
		\g15_reg/NET0131 ,
		_w804_,
		_w812_
	);
	LUT2 #(
		.INIT('h4)
	) name666 (
		\g19_reg/NET0131 ,
		_w804_,
		_w813_
	);
	assign \_al_n1  = 1'b0;
	assign \g10560/_0_  = _w164_ ;
	assign \g10562/_1_  = _w167_ ;
	assign \g10564/_1_  = _w170_ ;
	assign \g10566/_1_  = _w172_ ;
	assign \g10567/_0_  = _w175_ ;
	assign \g10569/_1_  = _w178_ ;
	assign \g10580/_0_  = _w199_ ;
	assign \g10616/_2_  = _w379_ ;
	assign \g10627/_2_  = _w414_ ;
	assign \g10628/_0_  = _w425_ ;
	assign \g10629/_2_  = _w467_ ;
	assign \g10630/_2_  = _w502_ ;
	assign \g10633/_2_  = _w527_ ;
	assign \g10635/_2_  = _w564_ ;
	assign \g10636/_2_  = _w594_ ;
	assign \g10637/_2_  = _w618_ ;
	assign \g10641/_0_  = _w621_ ;
	assign \g10649/_0_  = _w624_ ;
	assign \g10672/_0_  = _w332_ ;
	assign \g10673/_0_  = _w273_ ;
	assign \g10680/_0_  = _w627_ ;
	assign \g10683/_0_  = _w628_ ;
	assign \g10686/_0_  = _w629_ ;
	assign \g10695/_0_  = _w403_ ;
	assign \g10700/_0_  = _w632_ ;
	assign \g10703/_0_  = _w270_ ;
	assign \g10704/_0_  = _w692_ ;
	assign \g10748/_0_  = _w695_ ;
	assign \g10750/_2_  = _w384_ ;
	assign \g10757/_0_  = _w516_ ;
	assign \g10758/_0_  = _w509_ ;
	assign \g10782/_0_  = _w698_ ;
	assign \g10826/_0_  = _w699_ ;
	assign \g10827/_0_  = _w700_ ;
	assign \g10828/_1_  = _w701_ ;
	assign \g10832/_2_  = _w607_ ;
	assign \g10834/_2_  = _w600_ ;
	assign \g10836/_0_  = _w704_ ;
	assign \g10837/_1__syn_2  = _w705_ ;
	assign \g10868/_0_  = _w708_ ;
	assign \g10904/_0_  = _w728_ ;
	assign \g10913/_0_  = _w483_ ;
	assign \g10915/_0_  = _w473_ ;
	assign \g10922/_0_  = _w731_ ;
	assign \g10938/_0_  = _w567_ ;
	assign \g10939/_0_  = _w532_ ;
	assign \g10940/_0_  = _w571_ ;
	assign \g10941/_0_  = _w548_ ;
	assign \g10942/_0_  = _w432_ ;
	assign \g10944/_2_  = _w454_ ;
	assign \g10977/_0_  = _w734_ ;
	assign \g10980/_0_  = _w736_ ;
	assign \g11020/_0_  = _w726_ ;
	assign \g11028/_0_  = _w738_ ;
	assign \g11051/_0_  = _w768_ ;
	assign \g11057/_0_  = _w771_ ;
	assign \g11109/_0_  = _w774_ ;
	assign \g11113/_2_  = _w685_ ;
	assign \g11156/_0_  = _w777_ ;
	assign \g11172/_3_  = _w780_ ;
	assign \g11193/_0_  = _w783_ ;
	assign \g11219/_0_  = _w786_ ;
	assign \g11355/_0_  = \g678_reg/NET0131 ;
	assign \g11384/_0_  = \g677_reg/NET0131 ;
	assign \g11442/_0_  = _w787_ ;
	assign \g11448/_0_  = _w788_ ;
	assign \g11558/_0_  = \g266_reg/NET0131 ;
	assign \g11559/_0_  = \g4112_pad ;
	assign \g11824/_1_  = _w387_ ;
	assign \g11853/_0_  = _w796_ ;
	assign \g11854/_0_  = _w662_ ;
	assign \g11977/_0_  = _w329_ ;
	assign \g11981/_0_  = _w400_ ;
	assign \g2584_pad  = _w797_ ;
	assign \g4121_pad  = _w798_ ;
	assign \g4809_pad  = _w801_ ;
	assign \g5692_pad  = 1'b0;
	assign \g6282_pad  = _w803_ ;
	assign \g6284_pad  = _w805_ ;
	assign \g6360_pad  = _w806_ ;
	assign \g6362_pad  = _w807_ ;
	assign \g6364_pad  = _w808_ ;
	assign \g6366_pad  = _w809_ ;
	assign \g6368_pad  = _w810_ ;
	assign \g6370_pad  = _w811_ ;
	assign \g6372_pad  = _w812_ ;
	assign \g6374_pad  = _w813_ ;
endmodule;