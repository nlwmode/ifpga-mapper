module top (a_pad, b_pad, c_pad, e_pad, f_pad, g_pad, h_pad, i_pad, j_pad, k_pad, l_pad, m_pad, n_pad, o_pad, p_pad, q_pad, r_pad, s_pad, t_pad, u_pad, v_pad, w_pad, x_pad, y_pad, \a0_pad , \b0_pad , \c0_pad , \d0_pad , \e0_pad , \f0_pad , \g0_pad , \h0_pad , \i0_pad , \j0_pad , \k0_pad , \l0_pad , \m0_pad , \n0_pad , \o0_pad , \p0_pad , \q0_pad , \r0_pad , \s0_pad , \t0_pad , z_pad);
	input a_pad ;
	input b_pad ;
	input c_pad ;
	input e_pad ;
	input f_pad ;
	input g_pad ;
	input h_pad ;
	input i_pad ;
	input j_pad ;
	input k_pad ;
	input l_pad ;
	input m_pad ;
	input n_pad ;
	input o_pad ;
	input p_pad ;
	input q_pad ;
	input r_pad ;
	input s_pad ;
	input t_pad ;
	input u_pad ;
	input v_pad ;
	input w_pad ;
	input x_pad ;
	input y_pad ;
	output \a0_pad  ;
	output \b0_pad  ;
	output \c0_pad  ;
	output \d0_pad  ;
	output \e0_pad  ;
	output \f0_pad  ;
	output \g0_pad  ;
	output \h0_pad  ;
	output \i0_pad  ;
	output \j0_pad  ;
	output \k0_pad  ;
	output \l0_pad  ;
	output \m0_pad  ;
	output \n0_pad  ;
	output \o0_pad  ;
	output \p0_pad  ;
	output \q0_pad  ;
	output \r0_pad  ;
	output \s0_pad  ;
	output \t0_pad  ;
	output z_pad ;
	wire _w98_ ;
	wire _w97_ ;
	wire _w96_ ;
	wire _w95_ ;
	wire _w94_ ;
	wire _w93_ ;
	wire _w92_ ;
	wire _w91_ ;
	wire _w90_ ;
	wire _w89_ ;
	wire _w88_ ;
	wire _w87_ ;
	wire _w86_ ;
	wire _w85_ ;
	wire _w54_ ;
	wire _w53_ ;
	wire _w52_ ;
	wire _w51_ ;
	wire _w50_ ;
	wire _w49_ ;
	wire _w48_ ;
	wire _w47_ ;
	wire _w46_ ;
	wire _w45_ ;
	wire _w44_ ;
	wire _w43_ ;
	wire _w42_ ;
	wire _w41_ ;
	wire _w40_ ;
	wire _w39_ ;
	wire _w26_ ;
	wire _w27_ ;
	wire _w28_ ;
	wire _w29_ ;
	wire _w30_ ;
	wire _w31_ ;
	wire _w32_ ;
	wire _w33_ ;
	wire _w34_ ;
	wire _w35_ ;
	wire _w36_ ;
	wire _w37_ ;
	wire _w38_ ;
	wire _w55_ ;
	wire _w56_ ;
	wire _w57_ ;
	wire _w58_ ;
	wire _w59_ ;
	wire _w60_ ;
	wire _w61_ ;
	wire _w62_ ;
	wire _w63_ ;
	wire _w64_ ;
	wire _w65_ ;
	wire _w66_ ;
	wire _w67_ ;
	wire _w68_ ;
	wire _w69_ ;
	wire _w70_ ;
	wire _w71_ ;
	wire _w72_ ;
	wire _w73_ ;
	wire _w74_ ;
	wire _w75_ ;
	wire _w76_ ;
	wire _w77_ ;
	wire _w78_ ;
	wire _w79_ ;
	wire _w80_ ;
	wire _w81_ ;
	wire _w82_ ;
	wire _w83_ ;
	wire _w84_ ;
	LUT4 #(
		.INIT('ha800)
	) name0 (
		f_pad,
		t_pad,
		u_pad,
		v_pad,
		_w26_
	);
	LUT4 #(
		.INIT('h1110)
	) name1 (
		s_pad,
		t_pad,
		v_pad,
		y_pad,
		_w27_
	);
	LUT2 #(
		.INIT('h2)
	) name2 (
		u_pad,
		v_pad,
		_w28_
	);
	LUT2 #(
		.INIT('h4)
	) name3 (
		u_pad,
		v_pad,
		_w29_
	);
	LUT2 #(
		.INIT('h9)
	) name4 (
		u_pad,
		v_pad,
		_w30_
	);
	LUT4 #(
		.INIT('h0051)
	) name5 (
		w_pad,
		_w27_,
		_w30_,
		_w26_,
		_w31_
	);
	LUT3 #(
		.INIT('ha2)
	) name6 (
		q_pad,
		v_pad,
		w_pad,
		_w32_
	);
	LUT4 #(
		.INIT('h0002)
	) name7 (
		s_pad,
		t_pad,
		v_pad,
		y_pad,
		_w33_
	);
	LUT3 #(
		.INIT('h13)
	) name8 (
		u_pad,
		_w32_,
		_w33_,
		_w34_
	);
	LUT2 #(
		.INIT('h4)
	) name9 (
		_w31_,
		_w34_,
		_w35_
	);
	LUT4 #(
		.INIT('he0f0)
	) name10 (
		s_pad,
		t_pad,
		u_pad,
		y_pad,
		_w36_
	);
	LUT2 #(
		.INIT('h1)
	) name11 (
		v_pad,
		_w36_,
		_w37_
	);
	LUT4 #(
		.INIT('h5700)
	) name12 (
		g_pad,
		t_pad,
		u_pad,
		v_pad,
		_w38_
	);
	LUT3 #(
		.INIT('h0d)
	) name13 (
		w_pad,
		_w33_,
		_w38_,
		_w39_
	);
	LUT2 #(
		.INIT('h4)
	) name14 (
		_w37_,
		_w39_,
		_w40_
	);
	LUT2 #(
		.INIT('h1)
	) name15 (
		u_pad,
		w_pad,
		_w41_
	);
	LUT4 #(
		.INIT('h3320)
	) name16 (
		q_pad,
		v_pad,
		_w27_,
		_w41_,
		_w42_
	);
	LUT3 #(
		.INIT('h51)
	) name17 (
		h_pad,
		u_pad,
		v_pad,
		_w43_
	);
	LUT4 #(
		.INIT('h2aaa)
	) name18 (
		q_pad,
		u_pad,
		_w33_,
		_w43_,
		_w44_
	);
	LUT4 #(
		.INIT('h5404)
	) name19 (
		h_pad,
		t_pad,
		u_pad,
		v_pad,
		_w45_
	);
	LUT3 #(
		.INIT('h02)
	) name20 (
		s_pad,
		t_pad,
		u_pad,
		_w46_
	);
	LUT4 #(
		.INIT('h000d)
	) name21 (
		w_pad,
		_w33_,
		_w45_,
		_w46_,
		_w47_
	);
	LUT4 #(
		.INIT('h3302)
	) name22 (
		w_pad,
		_w42_,
		_w44_,
		_w47_,
		_w48_
	);
	LUT4 #(
		.INIT('h00f7)
	) name23 (
		s_pad,
		t_pad,
		u_pad,
		v_pad,
		_w49_
	);
	LUT4 #(
		.INIT('h5700)
	) name24 (
		i_pad,
		t_pad,
		u_pad,
		v_pad,
		_w50_
	);
	LUT3 #(
		.INIT('h01)
	) name25 (
		w_pad,
		_w50_,
		_w49_,
		_w51_
	);
	LUT4 #(
		.INIT('h0207)
	) name26 (
		s_pad,
		t_pad,
		u_pad,
		v_pad,
		_w52_
	);
	LUT4 #(
		.INIT('ha800)
	) name27 (
		j_pad,
		t_pad,
		u_pad,
		v_pad,
		_w53_
	);
	LUT3 #(
		.INIT('h54)
	) name28 (
		w_pad,
		_w52_,
		_w53_,
		_w54_
	);
	LUT2 #(
		.INIT('h1)
	) name29 (
		a_pad,
		k_pad,
		_w55_
	);
	LUT3 #(
		.INIT('h10)
	) name30 (
		a_pad,
		k_pad,
		l_pad,
		_w56_
	);
	LUT2 #(
		.INIT('h4)
	) name31 (
		m_pad,
		n_pad,
		_w57_
	);
	LUT3 #(
		.INIT('h04)
	) name32 (
		a_pad,
		k_pad,
		l_pad,
		_w58_
	);
	LUT3 #(
		.INIT('hba)
	) name33 (
		_w56_,
		_w57_,
		_w58_,
		_w59_
	);
	LUT3 #(
		.INIT('h80)
	) name34 (
		k_pad,
		l_pad,
		m_pad,
		_w60_
	);
	LUT4 #(
		.INIT('h1540)
	) name35 (
		a_pad,
		k_pad,
		l_pad,
		m_pad,
		_w61_
	);
	LUT4 #(
		.INIT('h5551)
	) name36 (
		a_pad,
		k_pad,
		l_pad,
		m_pad,
		_w62_
	);
	LUT3 #(
		.INIT('h60)
	) name37 (
		n_pad,
		_w60_,
		_w62_,
		_w63_
	);
	LUT4 #(
		.INIT('h0200)
	) name38 (
		k_pad,
		l_pad,
		m_pad,
		n_pad,
		_w64_
	);
	LUT3 #(
		.INIT('ha8)
	) name39 (
		o_pad,
		x_pad,
		_w64_,
		_w65_
	);
	LUT4 #(
		.INIT('h1114)
	) name40 (
		a_pad,
		o_pad,
		x_pad,
		_w64_,
		_w66_
	);
	LUT2 #(
		.INIT('h4)
	) name41 (
		q_pad,
		r_pad,
		_w67_
	);
	LUT4 #(
		.INIT('h8880)
	) name42 (
		o_pad,
		p_pad,
		x_pad,
		_w64_,
		_w68_
	);
	LUT4 #(
		.INIT('h0414)
	) name43 (
		a_pad,
		p_pad,
		_w65_,
		_w67_,
		_w69_
	);
	LUT3 #(
		.INIT('h14)
	) name44 (
		a_pad,
		q_pad,
		_w68_,
		_w70_
	);
	LUT3 #(
		.INIT('h13)
	) name45 (
		q_pad,
		r_pad,
		_w68_,
		_w71_
	);
	LUT3 #(
		.INIT('h6e)
	) name46 (
		p_pad,
		q_pad,
		r_pad,
		_w72_
	);
	LUT4 #(
		.INIT('h00a8)
	) name47 (
		o_pad,
		x_pad,
		_w64_,
		_w72_,
		_w73_
	);
	LUT2 #(
		.INIT('h1)
	) name48 (
		a_pad,
		_w73_,
		_w74_
	);
	LUT2 #(
		.INIT('h4)
	) name49 (
		_w71_,
		_w74_,
		_w75_
	);
	LUT3 #(
		.INIT('h10)
	) name50 (
		p_pad,
		q_pad,
		r_pad,
		_w76_
	);
	LUT4 #(
		.INIT('ha800)
	) name51 (
		o_pad,
		x_pad,
		_w64_,
		_w76_,
		_w77_
	);
	LUT3 #(
		.INIT('h14)
	) name52 (
		a_pad,
		s_pad,
		_w77_,
		_w78_
	);
	LUT4 #(
		.INIT('h3133)
	) name53 (
		s_pad,
		t_pad,
		_w29_,
		_w77_,
		_w79_
	);
	LUT4 #(
		.INIT('h1555)
	) name54 (
		a_pad,
		s_pad,
		t_pad,
		_w77_,
		_w80_
	);
	LUT2 #(
		.INIT('h4)
	) name55 (
		_w79_,
		_w80_,
		_w81_
	);
	LUT4 #(
		.INIT('h870f)
	) name56 (
		s_pad,
		t_pad,
		u_pad,
		_w77_,
		_w82_
	);
	LUT2 #(
		.INIT('h1)
	) name57 (
		a_pad,
		_w82_,
		_w83_
	);
	LUT2 #(
		.INIT('h4)
	) name58 (
		t_pad,
		u_pad,
		_w84_
	);
	LUT2 #(
		.INIT('h9)
	) name59 (
		t_pad,
		u_pad,
		_w85_
	);
	LUT4 #(
		.INIT('h4ccc)
	) name60 (
		s_pad,
		v_pad,
		_w77_,
		_w85_,
		_w86_
	);
	LUT4 #(
		.INIT('h8000)
	) name61 (
		s_pad,
		t_pad,
		_w28_,
		_w77_,
		_w87_
	);
	LUT3 #(
		.INIT('h54)
	) name62 (
		a_pad,
		_w86_,
		_w87_,
		_w88_
	);
	LUT3 #(
		.INIT('h10)
	) name63 (
		s_pad,
		v_pad,
		y_pad,
		_w89_
	);
	LUT3 #(
		.INIT('h15)
	) name64 (
		w_pad,
		_w84_,
		_w89_,
		_w90_
	);
	LUT3 #(
		.INIT('h15)
	) name65 (
		a_pad,
		u_pad,
		_w33_,
		_w91_
	);
	LUT2 #(
		.INIT('h4)
	) name66 (
		_w90_,
		_w91_,
		_w92_
	);
	LUT3 #(
		.INIT('h14)
	) name67 (
		a_pad,
		b_pad,
		x_pad,
		_w93_
	);
	LUT3 #(
		.INIT('h14)
	) name68 (
		a_pad,
		c_pad,
		y_pad,
		_w94_
	);
	LUT3 #(
		.INIT('ha8)
	) name69 (
		e_pad,
		t_pad,
		u_pad,
		_w95_
	);
	LUT4 #(
		.INIT('hfd00)
	) name70 (
		s_pad,
		t_pad,
		u_pad,
		v_pad,
		_w96_
	);
	LUT3 #(
		.INIT('h0d)
	) name71 (
		u_pad,
		v_pad,
		w_pad,
		_w97_
	);
	LUT3 #(
		.INIT('hb0)
	) name72 (
		_w95_,
		_w96_,
		_w97_,
		_w98_
	);
	assign \a0_pad  = _w35_ ;
	assign \b0_pad  = _w40_ ;
	assign \c0_pad  = _w48_ ;
	assign \d0_pad  = _w51_ ;
	assign \e0_pad  = _w54_ ;
	assign \f0_pad  = _w55_ ;
	assign \g0_pad  = _w59_ ;
	assign \h0_pad  = _w61_ ;
	assign \i0_pad  = _w63_ ;
	assign \j0_pad  = _w66_ ;
	assign \k0_pad  = _w69_ ;
	assign \l0_pad  = _w70_ ;
	assign \m0_pad  = _w75_ ;
	assign \n0_pad  = _w78_ ;
	assign \o0_pad  = _w81_ ;
	assign \p0_pad  = _w83_ ;
	assign \q0_pad  = _w88_ ;
	assign \r0_pad  = _w92_ ;
	assign \s0_pad  = _w93_ ;
	assign \t0_pad  = _w94_ ;
	assign z_pad = _w98_ ;
endmodule;