module top (mc_cke_pad_o__pad, mc_vpen_pad_o_pad, \mem_ack_r_reg/P0001 , \poc_o[0]_pad , \poc_o[10]_pad , \poc_o[11]_pad , \poc_o[12]_pad , \poc_o[13]_pad , \poc_o[14]_pad , \poc_o[15]_pad , \poc_o[16]_pad , \poc_o[17]_pad , \poc_o[18]_pad , \poc_o[19]_pad , \poc_o[1]_pad , \poc_o[20]_pad , \poc_o[21]_pad , \poc_o[22]_pad , \poc_o[23]_pad , \poc_o[24]_pad , \poc_o[25]_pad , \poc_o[26]_pad , \poc_o[27]_pad , \poc_o[28]_pad , \poc_o[29]_pad , \poc_o[2]_pad , \poc_o[30]_pad , \poc_o[31]_pad , \poc_o[3]_pad , \poc_o[4]_pad , \poc_o[5]_pad , \poc_o[6]_pad , \poc_o[7]_pad , \poc_o[8]_pad , \poc_o[9]_pad , suspended_o_pad, \u0_cs_reg[0]/NET0131 , \u0_cs_reg[1]/NET0131 , \u0_csc_mask_r_reg[0]/NET0131 , \u0_csc_mask_r_reg[10]/NET0131 , \u0_csc_mask_r_reg[1]/NET0131 , \u0_csc_mask_r_reg[2]/NET0131 , \u0_csc_mask_r_reg[3]/NET0131 , \u0_csc_mask_r_reg[4]/NET0131 , \u0_csc_mask_r_reg[5]/NET0131 , \u0_csc_mask_r_reg[6]/NET0131 , \u0_csc_mask_r_reg[7]/NET0131 , \u0_csc_mask_r_reg[8]/NET0131 , \u0_csc_mask_r_reg[9]/NET0131 , \u0_csc_reg[10]/NET0131 , \u0_csc_reg[11]/NET0131 , \u0_csc_reg[1]/NET0131 , \u0_csc_reg[2]/NET0131 , \u0_csc_reg[3]/NET0131 , \u0_csc_reg[4]/NET0131 , \u0_csc_reg[5]/NET0131 , \u0_csc_reg[6]/NET0131 , \u0_csc_reg[7]/NET0131 , \u0_csc_reg[9]/NET0131 , \u0_csr_r2_reg[0]/NET0131 , \u0_csr_r2_reg[1]/NET0131 , \u0_csr_r2_reg[2]/NET0131 , \u0_csr_r2_reg[3]/NET0131 , \u0_csr_r2_reg[4]/NET0131 , \u0_csr_r2_reg[5]/NET0131 , \u0_csr_r2_reg[6]/NET0131 , \u0_csr_r2_reg[7]/NET0131 , \u0_csr_r_reg[0]/P0001 , \u0_csr_r_reg[10]/NET0131 , \u0_csr_r_reg[2]/NET0131 , \u0_csr_r_reg[3]/NET0131 , \u0_csr_r_reg[4]/NET0131 , \u0_csr_r_reg[5]/NET0131 , \u0_csr_r_reg[6]/NET0131 , \u0_csr_r_reg[7]/NET0131 , \u0_csr_r_reg[8]/NET0131 , \u0_csr_r_reg[9]/NET0131 , \u0_init_ack_r_reg/P0001 , \u0_init_req_reg/NET0131 , \u0_lmr_ack_r_reg/P0001 , \u0_lmr_req_reg/NET0131 , \u0_rf_we_reg/NET0131 , \u0_rst_r2_reg/NET0131 , \u0_sp_csc_reg[10]/NET0131 , \u0_sp_csc_reg[1]/NET0131 , \u0_sp_csc_reg[2]/NET0131 , \u0_sp_csc_reg[3]/NET0131 , \u0_sp_csc_reg[4]/NET0131 , \u0_sp_csc_reg[5]/NET0131 , \u0_sp_csc_reg[6]/NET0131 , \u0_sp_csc_reg[7]/NET0131 , \u0_sp_csc_reg[9]/NET0131 , \u0_sp_tms_reg[0]/NET0131 , \u0_sp_tms_reg[10]/NET0131 , \u0_sp_tms_reg[11]/NET0131 , \u0_sp_tms_reg[12]/NET0131 , \u0_sp_tms_reg[13]/NET0131 , \u0_sp_tms_reg[14]/NET0131 , \u0_sp_tms_reg[15]/NET0131 , \u0_sp_tms_reg[16]/NET0131 , \u0_sp_tms_reg[17]/NET0131 , \u0_sp_tms_reg[18]/NET0131 , \u0_sp_tms_reg[19]/NET0131 , \u0_sp_tms_reg[1]/NET0131 , \u0_sp_tms_reg[20]/NET0131 , \u0_sp_tms_reg[21]/NET0131 , \u0_sp_tms_reg[22]/NET0131 , \u0_sp_tms_reg[23]/NET0131 , \u0_sp_tms_reg[24]/NET0131 , \u0_sp_tms_reg[25]/NET0131 , \u0_sp_tms_reg[26]/NET0131 , \u0_sp_tms_reg[27]/NET0131 , \u0_sp_tms_reg[2]/NET0131 , \u0_sp_tms_reg[3]/NET0131 , \u0_sp_tms_reg[4]/NET0131 , \u0_sp_tms_reg[5]/NET0131 , \u0_sp_tms_reg[6]/NET0131 , \u0_sp_tms_reg[7]/NET0131 , \u0_sp_tms_reg[8]/NET0131 , \u0_sp_tms_reg[9]/NET0131 , \u0_spec_req_cs_reg[0]/NET0131 , \u0_spec_req_cs_reg[1]/NET0131 , \u0_sreq_cs_le_reg/NET0131 , \u0_tms_reg[0]/NET0131 , \u0_tms_reg[10]/NET0131 , \u0_tms_reg[11]/NET0131 , \u0_tms_reg[12]/NET0131 , \u0_tms_reg[13]/NET0131 , \u0_tms_reg[14]/NET0131 , \u0_tms_reg[15]/NET0131 , \u0_tms_reg[16]/NET0131 , \u0_tms_reg[17]/NET0131 , \u0_tms_reg[18]/NET0131 , \u0_tms_reg[19]/NET0131 , \u0_tms_reg[1]/NET0131 , \u0_tms_reg[20]/NET0131 , \u0_tms_reg[21]/NET0131 , \u0_tms_reg[22]/NET0131 , \u0_tms_reg[23]/NET0131 , \u0_tms_reg[24]/NET0131 , \u0_tms_reg[25]/NET0131 , \u0_tms_reg[26]/NET0131 , \u0_tms_reg[27]/NET0131 , \u0_tms_reg[2]/NET0131 , \u0_tms_reg[3]/NET0131 , \u0_tms_reg[4]/NET0131 , \u0_tms_reg[5]/NET0131 , \u0_tms_reg[6]/NET0131 , \u0_tms_reg[7]/NET0131 , \u0_tms_reg[8]/NET0131 , \u0_tms_reg[9]/NET0131 , \u0_u0_addr_r_reg[2]/P0001 , \u0_u0_addr_r_reg[3]/P0001 , \u0_u0_addr_r_reg[4]/P0001 , \u0_u0_addr_r_reg[5]/P0001 , \u0_u0_addr_r_reg[6]/P0001 , \u0_u0_csc_reg[0]/NET0131 , \u0_u0_csc_reg[10]/P0001 , \u0_u0_csc_reg[11]/P0001 , \u0_u0_csc_reg[12]/P0001 , \u0_u0_csc_reg[13]/P0001 , \u0_u0_csc_reg[14]/P0001 , \u0_u0_csc_reg[15]/P0001 , \u0_u0_csc_reg[16]/P0001 , \u0_u0_csc_reg[17]/P0001 , \u0_u0_csc_reg[18]/P0001 , \u0_u0_csc_reg[19]/P0001 , \u0_u0_csc_reg[1]/NET0131 , \u0_u0_csc_reg[20]/P0001 , \u0_u0_csc_reg[21]/P0001 , \u0_u0_csc_reg[22]/P0001 , \u0_u0_csc_reg[23]/P0001 , \u0_u0_csc_reg[24]/P0001 , \u0_u0_csc_reg[25]/P0001 , \u0_u0_csc_reg[26]/P0001 , \u0_u0_csc_reg[27]/P0001 , \u0_u0_csc_reg[28]/P0001 , \u0_u0_csc_reg[29]/P0001 , \u0_u0_csc_reg[2]/NET0131 , \u0_u0_csc_reg[30]/P0001 , \u0_u0_csc_reg[31]/P0001 , \u0_u0_csc_reg[3]/NET0131 , \u0_u0_csc_reg[4]/P0001 , \u0_u0_csc_reg[5]/P0001 , \u0_u0_csc_reg[6]/P0001 , \u0_u0_csc_reg[7]/P0001 , \u0_u0_csc_reg[8]/P0001 , \u0_u0_csc_reg[9]/P0001 , \u0_u0_init_req_reg/NET0131 , \u0_u0_init_req_we_reg/NET0131 , \u0_u0_inited_reg/NET0131 , \u0_u0_lmr_req_reg/NET0131 , \u0_u0_lmr_req_we_reg/NET0131 , \u0_u0_tms_reg[0]/P0001 , \u0_u0_tms_reg[10]/P0001 , \u0_u0_tms_reg[11]/P0001 , \u0_u0_tms_reg[12]/P0001 , \u0_u0_tms_reg[13]/P0001 , \u0_u0_tms_reg[14]/P0001 , \u0_u0_tms_reg[15]/P0001 , \u0_u0_tms_reg[16]/P0001 , \u0_u0_tms_reg[17]/P0001 , \u0_u0_tms_reg[18]/P0001 , \u0_u0_tms_reg[19]/P0001 , \u0_u0_tms_reg[1]/P0001 , \u0_u0_tms_reg[20]/P0001 , \u0_u0_tms_reg[21]/P0001 , \u0_u0_tms_reg[22]/P0001 , \u0_u0_tms_reg[23]/P0001 , \u0_u0_tms_reg[24]/P0001 , \u0_u0_tms_reg[25]/P0001 , \u0_u0_tms_reg[26]/P0001 , \u0_u0_tms_reg[27]/P0001 , \u0_u0_tms_reg[28]/P0001 , \u0_u0_tms_reg[29]/P0001 , \u0_u0_tms_reg[2]/P0001 , \u0_u0_tms_reg[30]/P0001 , \u0_u0_tms_reg[31]/P0001 , \u0_u0_tms_reg[3]/P0001 , \u0_u0_tms_reg[4]/P0001 , \u0_u0_tms_reg[5]/P0001 , \u0_u0_tms_reg[6]/P0001 , \u0_u0_tms_reg[7]/P0001 , \u0_u0_tms_reg[8]/P0001 , \u0_u0_tms_reg[9]/P0001 , \u0_u1_csc_reg[0]/NET0131 , \u0_u1_csc_reg[10]/P0001 , \u0_u1_csc_reg[11]/P0001 , \u0_u1_csc_reg[12]/P0001 , \u0_u1_csc_reg[13]/P0001 , \u0_u1_csc_reg[14]/P0001 , \u0_u1_csc_reg[15]/P0001 , \u0_u1_csc_reg[16]/P0001 , \u0_u1_csc_reg[17]/P0001 , \u0_u1_csc_reg[18]/P0001 , \u0_u1_csc_reg[19]/P0001 , \u0_u1_csc_reg[1]/NET0131 , \u0_u1_csc_reg[20]/P0001 , \u0_u1_csc_reg[21]/P0001 , \u0_u1_csc_reg[22]/P0001 , \u0_u1_csc_reg[23]/P0001 , \u0_u1_csc_reg[24]/P0001 , \u0_u1_csc_reg[25]/P0001 , \u0_u1_csc_reg[26]/P0001 , \u0_u1_csc_reg[27]/P0001 , \u0_u1_csc_reg[28]/P0001 , \u0_u1_csc_reg[29]/P0001 , \u0_u1_csc_reg[2]/NET0131 , \u0_u1_csc_reg[30]/P0001 , \u0_u1_csc_reg[31]/P0001 , \u0_u1_csc_reg[3]/NET0131 , \u0_u1_csc_reg[4]/P0001 , \u0_u1_csc_reg[5]/P0001 , \u0_u1_csc_reg[6]/P0001 , \u0_u1_csc_reg[7]/P0001 , \u0_u1_csc_reg[8]/P0001 , \u0_u1_csc_reg[9]/P0001 , \u0_u1_init_req_reg/NET0131 , \u0_u1_init_req_we_reg/NET0131 , \u0_u1_inited_reg/NET0131 , \u0_u1_lmr_req_reg/NET0131 , \u0_u1_lmr_req_we_reg/NET0131 , \u0_u1_tms_reg[0]/P0001 , \u0_u1_tms_reg[10]/P0001 , \u0_u1_tms_reg[11]/P0001 , \u0_u1_tms_reg[12]/P0001 , \u0_u1_tms_reg[13]/P0001 , \u0_u1_tms_reg[14]/P0001 , \u0_u1_tms_reg[15]/P0001 , \u0_u1_tms_reg[16]/P0001 , \u0_u1_tms_reg[17]/P0001 , \u0_u1_tms_reg[18]/P0001 , \u0_u1_tms_reg[19]/P0001 , \u0_u1_tms_reg[1]/P0001 , \u0_u1_tms_reg[20]/P0001 , \u0_u1_tms_reg[21]/P0001 , \u0_u1_tms_reg[22]/P0001 , \u0_u1_tms_reg[23]/P0001 , \u0_u1_tms_reg[24]/P0001 , \u0_u1_tms_reg[25]/P0001 , \u0_u1_tms_reg[26]/P0001 , \u0_u1_tms_reg[27]/P0001 , \u0_u1_tms_reg[28]/P0001 , \u0_u1_tms_reg[29]/P0001 , \u0_u1_tms_reg[2]/P0001 , \u0_u1_tms_reg[30]/P0001 , \u0_u1_tms_reg[31]/P0001 , \u0_u1_tms_reg[3]/P0001 , \u0_u1_tms_reg[4]/P0001 , \u0_u1_tms_reg[5]/P0001 , \u0_u1_tms_reg[6]/P0001 , \u0_u1_tms_reg[7]/P0001 , \u0_u1_tms_reg[8]/P0001 , \u0_u1_tms_reg[9]/P0001 , \u0_wp_err_reg/NET0131 , \u1_acs_addr_reg[0]/P0001 , \u1_acs_addr_reg[10]/P0001 , \u1_acs_addr_reg[11]/P0001 , \u1_acs_addr_reg[12]/P0001 , \u1_acs_addr_reg[13]/P0001 , \u1_acs_addr_reg[14]/P0001 , \u1_acs_addr_reg[15]/P0001 , \u1_acs_addr_reg[16]/P0001 , \u1_acs_addr_reg[17]/P0001 , \u1_acs_addr_reg[18]/P0001 , \u1_acs_addr_reg[19]/P0001 , \u1_acs_addr_reg[1]/P0001 , \u1_acs_addr_reg[20]/P0001 , \u1_acs_addr_reg[21]/P0001 , \u1_acs_addr_reg[22]/P0001 , \u1_acs_addr_reg[23]/P0001 , \u1_acs_addr_reg[2]/P0001 , \u1_acs_addr_reg[3]/P0001 , \u1_acs_addr_reg[4]/P0001 , \u1_acs_addr_reg[5]/P0001 , \u1_acs_addr_reg[6]/P0001 , \u1_acs_addr_reg[7]/P0001 , \u1_acs_addr_reg[8]/P0001 , \u1_acs_addr_reg[9]/P0001 , \u1_bank_adr_reg[0]/P0001 , \u1_bank_adr_reg[1]/P0001 , \u1_col_adr_reg[0]/P0001 , \u1_col_adr_reg[1]/P0001 , \u1_col_adr_reg[2]/P0001 , \u1_col_adr_reg[3]/P0001 , \u1_col_adr_reg[4]/P0001 , \u1_col_adr_reg[5]/P0001 , \u1_col_adr_reg[6]/P0001 , \u1_col_adr_reg[7]/P0001 , \u1_col_adr_reg[8]/P0001 , \u1_col_adr_reg[9]/P0001 , \u1_row_adr_reg[0]/P0001 , \u1_row_adr_reg[10]/P0001 , \u1_row_adr_reg[11]/P0001 , \u1_row_adr_reg[12]/P0001 , \u1_row_adr_reg[1]/P0001 , \u1_row_adr_reg[2]/P0001 , \u1_row_adr_reg[3]/P0001 , \u1_row_adr_reg[4]/P0001 , \u1_row_adr_reg[5]/P0001 , \u1_row_adr_reg[6]/P0001 , \u1_row_adr_reg[7]/P0001 , \u1_row_adr_reg[8]/P0001 , \u1_row_adr_reg[9]/P0001 , \u1_sram_addr_reg[0]/P0001 , \u1_sram_addr_reg[10]/P0001 , \u1_sram_addr_reg[11]/P0001 , \u1_sram_addr_reg[12]/P0001 , \u1_sram_addr_reg[13]/P0001 , \u1_sram_addr_reg[14]/P0001 , \u1_sram_addr_reg[15]/P0001 , \u1_sram_addr_reg[16]/P0001 , \u1_sram_addr_reg[17]/P0001 , \u1_sram_addr_reg[18]/P0001 , \u1_sram_addr_reg[19]/P0001 , \u1_sram_addr_reg[1]/P0001 , \u1_sram_addr_reg[20]/P0001 , \u1_sram_addr_reg[21]/P0001 , \u1_sram_addr_reg[22]/P0001 , \u1_sram_addr_reg[23]/P0001 , \u1_sram_addr_reg[2]/P0001 , \u1_sram_addr_reg[3]/P0001 , \u1_sram_addr_reg[4]/P0001 , \u1_sram_addr_reg[5]/P0001 , \u1_sram_addr_reg[6]/P0001 , \u1_sram_addr_reg[7]/P0001 , \u1_sram_addr_reg[8]/P0001 , \u1_sram_addr_reg[9]/P0001 , \u1_u0_out_r_reg[0]/P0001 , \u1_u0_out_r_reg[10]/P0001 , \u1_u0_out_r_reg[11]/P0001 , \u1_u0_out_r_reg[12]/P0001 , \u1_u0_out_r_reg[1]/P0001 , \u1_u0_out_r_reg[2]/P0001 , \u1_u0_out_r_reg[3]/P0001 , \u1_u0_out_r_reg[4]/P0001 , \u1_u0_out_r_reg[5]/P0001 , \u1_u0_out_r_reg[6]/P0001 , \u1_u0_out_r_reg[7]/P0001 , \u1_u0_out_r_reg[8]/P0001 , \u1_u0_out_r_reg[9]/P0001 , \u2_bank_open_reg/P0001 , \u2_row_same_reg/P0001 , \u2_u0_b0_last_row_reg[0]/P0001 , \u2_u0_b0_last_row_reg[10]/P0001 , \u2_u0_b0_last_row_reg[11]/P0001 , \u2_u0_b0_last_row_reg[12]/P0001 , \u2_u0_b0_last_row_reg[1]/P0001 , \u2_u0_b0_last_row_reg[2]/P0001 , \u2_u0_b0_last_row_reg[3]/P0001 , \u2_u0_b0_last_row_reg[4]/P0001 , \u2_u0_b0_last_row_reg[5]/P0001 , \u2_u0_b0_last_row_reg[6]/P0001 , \u2_u0_b0_last_row_reg[7]/P0001 , \u2_u0_b0_last_row_reg[8]/P0001 , \u2_u0_b0_last_row_reg[9]/P0001 , \u2_u0_b1_last_row_reg[0]/P0001 , \u2_u0_b1_last_row_reg[10]/P0001 , \u2_u0_b1_last_row_reg[11]/P0001 , \u2_u0_b1_last_row_reg[12]/P0001 , \u2_u0_b1_last_row_reg[1]/P0001 , \u2_u0_b1_last_row_reg[2]/P0001 , \u2_u0_b1_last_row_reg[3]/P0001 , \u2_u0_b1_last_row_reg[4]/P0001 , \u2_u0_b1_last_row_reg[5]/P0001 , \u2_u0_b1_last_row_reg[6]/P0001 , \u2_u0_b1_last_row_reg[7]/P0001 , \u2_u0_b1_last_row_reg[8]/P0001 , \u2_u0_b1_last_row_reg[9]/P0001 , \u2_u0_b2_last_row_reg[0]/P0001 , \u2_u0_b2_last_row_reg[10]/P0001 , \u2_u0_b2_last_row_reg[11]/P0001 , \u2_u0_b2_last_row_reg[12]/P0001 , \u2_u0_b2_last_row_reg[1]/P0001 , \u2_u0_b2_last_row_reg[2]/P0001 , \u2_u0_b2_last_row_reg[3]/P0001 , \u2_u0_b2_last_row_reg[4]/P0001 , \u2_u0_b2_last_row_reg[5]/P0001 , \u2_u0_b2_last_row_reg[6]/P0001 , \u2_u0_b2_last_row_reg[7]/P0001 , \u2_u0_b2_last_row_reg[8]/P0001 , \u2_u0_b2_last_row_reg[9]/P0001 , \u2_u0_b3_last_row_reg[0]/P0001 , \u2_u0_b3_last_row_reg[10]/P0001 , \u2_u0_b3_last_row_reg[11]/P0001 , \u2_u0_b3_last_row_reg[12]/P0001 , \u2_u0_b3_last_row_reg[1]/P0001 , \u2_u0_b3_last_row_reg[2]/P0001 , \u2_u0_b3_last_row_reg[3]/P0001 , \u2_u0_b3_last_row_reg[4]/P0001 , \u2_u0_b3_last_row_reg[5]/P0001 , \u2_u0_b3_last_row_reg[6]/P0001 , \u2_u0_b3_last_row_reg[7]/P0001 , \u2_u0_b3_last_row_reg[8]/P0001 , \u2_u0_b3_last_row_reg[9]/P0001 , \u2_u0_bank0_open_reg/NET0131 , \u2_u0_bank1_open_reg/NET0131 , \u2_u0_bank2_open_reg/NET0131 , \u2_u0_bank3_open_reg/NET0131 , \u2_u1_b0_last_row_reg[0]/P0001 , \u2_u1_b0_last_row_reg[10]/P0001 , \u2_u1_b0_last_row_reg[11]/P0001 , \u2_u1_b0_last_row_reg[12]/P0001 , \u2_u1_b0_last_row_reg[1]/P0001 , \u2_u1_b0_last_row_reg[2]/P0001 , \u2_u1_b0_last_row_reg[3]/P0001 , \u2_u1_b0_last_row_reg[4]/P0001 , \u2_u1_b0_last_row_reg[5]/P0001 , \u2_u1_b0_last_row_reg[6]/P0001 , \u2_u1_b0_last_row_reg[7]/P0001 , \u2_u1_b0_last_row_reg[8]/P0001 , \u2_u1_b0_last_row_reg[9]/P0001 , \u2_u1_b1_last_row_reg[0]/P0001 , \u2_u1_b1_last_row_reg[10]/P0001 , \u2_u1_b1_last_row_reg[11]/P0001 , \u2_u1_b1_last_row_reg[12]/P0001 , \u2_u1_b1_last_row_reg[1]/P0001 , \u2_u1_b1_last_row_reg[2]/P0001 , \u2_u1_b1_last_row_reg[3]/P0001 , \u2_u1_b1_last_row_reg[4]/P0001 , \u2_u1_b1_last_row_reg[5]/P0001 , \u2_u1_b1_last_row_reg[6]/P0001 , \u2_u1_b1_last_row_reg[7]/P0001 , \u2_u1_b1_last_row_reg[8]/P0001 , \u2_u1_b1_last_row_reg[9]/P0001 , \u2_u1_b2_last_row_reg[0]/P0001 , \u2_u1_b2_last_row_reg[10]/P0001 , \u2_u1_b2_last_row_reg[11]/P0001 , \u2_u1_b2_last_row_reg[12]/P0001 , \u2_u1_b2_last_row_reg[1]/P0001 , \u2_u1_b2_last_row_reg[2]/P0001 , \u2_u1_b2_last_row_reg[3]/P0001 , \u2_u1_b2_last_row_reg[4]/P0001 , \u2_u1_b2_last_row_reg[5]/P0001 , \u2_u1_b2_last_row_reg[6]/P0001 , \u2_u1_b2_last_row_reg[7]/P0001 , \u2_u1_b2_last_row_reg[8]/P0001 , \u2_u1_b2_last_row_reg[9]/P0001 , \u2_u1_b3_last_row_reg[0]/P0001 , \u2_u1_b3_last_row_reg[10]/P0001 , \u2_u1_b3_last_row_reg[11]/P0001 , \u2_u1_b3_last_row_reg[12]/P0001 , \u2_u1_b3_last_row_reg[1]/P0001 , \u2_u1_b3_last_row_reg[2]/P0001 , \u2_u1_b3_last_row_reg[3]/P0001 , \u2_u1_b3_last_row_reg[4]/P0001 , \u2_u1_b3_last_row_reg[5]/P0001 , \u2_u1_b3_last_row_reg[6]/P0001 , \u2_u1_b3_last_row_reg[7]/P0001 , \u2_u1_b3_last_row_reg[8]/P0001 , \u2_u1_b3_last_row_reg[9]/P0001 , \u2_u1_bank0_open_reg/NET0131 , \u2_u1_bank1_open_reg/NET0131 , \u2_u1_bank2_open_reg/NET0131 , \u2_u1_bank3_open_reg/NET0131 , \u3_byte0_reg[0]/P0001 , \u3_byte0_reg[1]/P0001 , \u3_byte0_reg[2]/P0001 , \u3_byte0_reg[3]/P0001 , \u3_byte0_reg[4]/P0001 , \u3_byte0_reg[5]/P0001 , \u3_byte0_reg[6]/P0001 , \u3_byte0_reg[7]/P0001 , \u3_byte1_reg[0]/P0001 , \u3_byte1_reg[1]/P0001 , \u3_byte1_reg[2]/P0001 , \u3_byte1_reg[3]/P0001 , \u3_byte1_reg[4]/P0001 , \u3_byte1_reg[5]/P0001 , \u3_byte1_reg[6]/P0001 , \u3_byte1_reg[7]/P0001 , \u3_byte2_reg[0]/P0001 , \u3_byte2_reg[1]/P0001 , \u3_byte2_reg[2]/P0001 , \u3_byte2_reg[3]/P0001 , \u3_byte2_reg[4]/P0001 , \u3_byte2_reg[5]/P0001 , \u3_byte2_reg[6]/P0001 , \u3_byte2_reg[7]/P0001 , \u3_u0_r0_reg[0]/P0001 , \u3_u0_r0_reg[10]/P0001 , \u3_u0_r0_reg[11]/P0001 , \u3_u0_r0_reg[12]/P0001 , \u3_u0_r0_reg[13]/P0001 , \u3_u0_r0_reg[14]/P0001 , \u3_u0_r0_reg[15]/P0001 , \u3_u0_r0_reg[16]/P0001 , \u3_u0_r0_reg[17]/P0001 , \u3_u0_r0_reg[18]/P0001 , \u3_u0_r0_reg[19]/P0001 , \u3_u0_r0_reg[1]/P0001 , \u3_u0_r0_reg[20]/P0001 , \u3_u0_r0_reg[21]/P0001 , \u3_u0_r0_reg[22]/P0001 , \u3_u0_r0_reg[23]/P0001 , \u3_u0_r0_reg[24]/P0001 , \u3_u0_r0_reg[25]/P0001 , \u3_u0_r0_reg[26]/P0001 , \u3_u0_r0_reg[27]/P0001 , \u3_u0_r0_reg[28]/P0001 , \u3_u0_r0_reg[29]/P0001 , \u3_u0_r0_reg[2]/P0001 , \u3_u0_r0_reg[30]/P0001 , \u3_u0_r0_reg[31]/P0001 , \u3_u0_r0_reg[32]/P0001 , \u3_u0_r0_reg[33]/P0001 , \u3_u0_r0_reg[34]/P0001 , \u3_u0_r0_reg[35]/P0001 , \u3_u0_r0_reg[3]/P0001 , \u3_u0_r0_reg[4]/P0001 , \u3_u0_r0_reg[5]/P0001 , \u3_u0_r0_reg[6]/P0001 , \u3_u0_r0_reg[7]/P0001 , \u3_u0_r0_reg[8]/P0001 , \u3_u0_r0_reg[9]/P0001 , \u3_u0_r1_reg[0]/P0001 , \u3_u0_r1_reg[10]/P0001 , \u3_u0_r1_reg[11]/P0001 , \u3_u0_r1_reg[12]/P0001 , \u3_u0_r1_reg[13]/P0001 , \u3_u0_r1_reg[14]/P0001 , \u3_u0_r1_reg[15]/P0001 , \u3_u0_r1_reg[16]/P0001 , \u3_u0_r1_reg[17]/P0001 , \u3_u0_r1_reg[18]/P0001 , \u3_u0_r1_reg[19]/P0001 , \u3_u0_r1_reg[1]/P0001 , \u3_u0_r1_reg[20]/P0001 , \u3_u0_r1_reg[21]/P0001 , \u3_u0_r1_reg[22]/P0001 , \u3_u0_r1_reg[23]/P0001 , \u3_u0_r1_reg[24]/P0001 , \u3_u0_r1_reg[25]/P0001 , \u3_u0_r1_reg[26]/P0001 , \u3_u0_r1_reg[27]/P0001 , \u3_u0_r1_reg[28]/P0001 , \u3_u0_r1_reg[29]/P0001 , \u3_u0_r1_reg[2]/P0001 , \u3_u0_r1_reg[30]/P0001 , \u3_u0_r1_reg[31]/P0001 , \u3_u0_r1_reg[32]/P0001 , \u3_u0_r1_reg[33]/P0001 , \u3_u0_r1_reg[34]/P0001 , \u3_u0_r1_reg[35]/P0001 , \u3_u0_r1_reg[3]/P0001 , \u3_u0_r1_reg[4]/P0001 , \u3_u0_r1_reg[5]/P0001 , \u3_u0_r1_reg[6]/P0001 , \u3_u0_r1_reg[7]/P0001 , \u3_u0_r1_reg[8]/P0001 , \u3_u0_r1_reg[9]/P0001 , \u3_u0_r2_reg[0]/P0001 , \u3_u0_r2_reg[10]/P0001 , \u3_u0_r2_reg[11]/P0001 , \u3_u0_r2_reg[12]/P0001 , \u3_u0_r2_reg[13]/P0001 , \u3_u0_r2_reg[14]/P0001 , \u3_u0_r2_reg[15]/P0001 , \u3_u0_r2_reg[16]/P0001 , \u3_u0_r2_reg[17]/P0001 , \u3_u0_r2_reg[18]/P0001 , \u3_u0_r2_reg[19]/P0001 , \u3_u0_r2_reg[1]/P0001 , \u3_u0_r2_reg[20]/P0001 , \u3_u0_r2_reg[21]/P0001 , \u3_u0_r2_reg[22]/P0001 , \u3_u0_r2_reg[23]/P0001 , \u3_u0_r2_reg[24]/P0001 , \u3_u0_r2_reg[25]/P0001 , \u3_u0_r2_reg[26]/P0001 , \u3_u0_r2_reg[27]/P0001 , \u3_u0_r2_reg[28]/P0001 , \u3_u0_r2_reg[29]/P0001 , \u3_u0_r2_reg[2]/P0001 , \u3_u0_r2_reg[30]/P0001 , \u3_u0_r2_reg[31]/P0001 , \u3_u0_r2_reg[32]/P0001 , \u3_u0_r2_reg[33]/P0001 , \u3_u0_r2_reg[34]/P0001 , \u3_u0_r2_reg[35]/P0001 , \u3_u0_r2_reg[3]/P0001 , \u3_u0_r2_reg[4]/P0001 , \u3_u0_r2_reg[5]/P0001 , \u3_u0_r2_reg[6]/P0001 , \u3_u0_r2_reg[7]/P0001 , \u3_u0_r2_reg[8]/P0001 , \u3_u0_r2_reg[9]/P0001 , \u3_u0_r3_reg[0]/P0001 , \u3_u0_r3_reg[10]/P0001 , \u3_u0_r3_reg[11]/P0001 , \u3_u0_r3_reg[12]/P0001 , \u3_u0_r3_reg[13]/P0001 , \u3_u0_r3_reg[14]/P0001 , \u3_u0_r3_reg[15]/P0001 , \u3_u0_r3_reg[16]/P0001 , \u3_u0_r3_reg[17]/P0001 , \u3_u0_r3_reg[18]/P0001 , \u3_u0_r3_reg[19]/P0001 , \u3_u0_r3_reg[1]/P0001 , \u3_u0_r3_reg[20]/P0001 , \u3_u0_r3_reg[21]/P0001 , \u3_u0_r3_reg[22]/P0001 , \u3_u0_r3_reg[23]/P0001 , \u3_u0_r3_reg[24]/P0001 , \u3_u0_r3_reg[25]/P0001 , \u3_u0_r3_reg[26]/P0001 , \u3_u0_r3_reg[27]/P0001 , \u3_u0_r3_reg[28]/P0001 , \u3_u0_r3_reg[29]/P0001 , \u3_u0_r3_reg[2]/P0001 , \u3_u0_r3_reg[30]/P0001 , \u3_u0_r3_reg[31]/P0001 , \u3_u0_r3_reg[32]/P0001 , \u3_u0_r3_reg[33]/P0001 , \u3_u0_r3_reg[34]/P0001 , \u3_u0_r3_reg[35]/P0001 , \u3_u0_r3_reg[3]/P0001 , \u3_u0_r3_reg[4]/P0001 , \u3_u0_r3_reg[5]/P0001 , \u3_u0_r3_reg[6]/P0001 , \u3_u0_r3_reg[7]/P0001 , \u3_u0_r3_reg[8]/P0001 , \u3_u0_r3_reg[9]/P0001 , \u3_u0_rd_adr_reg[0]/NET0131 , \u3_u0_rd_adr_reg[1]/NET0131 , \u3_u0_rd_adr_reg[2]/NET0131 , \u3_u0_rd_adr_reg[3]/NET0131 , \u3_u0_wr_adr_reg[0]/NET0131 , \u3_u0_wr_adr_reg[1]/NET0131 , \u3_u0_wr_adr_reg[2]/NET0131 , \u3_u0_wr_adr_reg[3]/NET0131 , \u4_ps_cnt_reg[0]/NET0131 , \u4_ps_cnt_reg[1]/NET0131 , \u4_ps_cnt_reg[2]/NET0131 , \u4_ps_cnt_reg[3]/NET0131 , \u4_ps_cnt_reg[4]/NET0131 , \u4_ps_cnt_reg[5]/NET0131 , \u4_ps_cnt_reg[6]/NET0131 , \u4_ps_cnt_reg[7]/NET0131 , \u4_rfr_ce_reg/NET0131 , \u4_rfr_clr_reg/P0001 , \u4_rfr_cnt_reg[0]/NET0131 , \u4_rfr_cnt_reg[1]/NET0131 , \u4_rfr_cnt_reg[2]/NET0131 , \u4_rfr_cnt_reg[3]/NET0131 , \u4_rfr_cnt_reg[4]/NET0131 , \u4_rfr_cnt_reg[5]/NET0131 , \u4_rfr_cnt_reg[6]/NET0131 , \u4_rfr_cnt_reg[7]/NET0131 , \u4_rfr_early_reg/NET0131 , \u4_rfr_en_reg/NET0131 , \u4_rfr_req_reg/NET0131 , \u5_ack_cnt_reg[0]/NET0131 , \u5_ack_cnt_reg[1]/NET0131 , \u5_ack_cnt_reg[2]/NET0131 , \u5_ack_cnt_reg[3]/NET0131 , \u5_ap_en_reg/NET0131 , \u5_burst_act_rd_reg/P0001 , \u5_burst_cnt_reg[0]/NET0131 , \u5_burst_cnt_reg[10]/NET0131 , \u5_burst_cnt_reg[1]/NET0131 , \u5_burst_cnt_reg[2]/NET0131 , \u5_burst_cnt_reg[3]/NET0131 , \u5_burst_cnt_reg[4]/NET0131 , \u5_burst_cnt_reg[5]/NET0131 , \u5_burst_cnt_reg[6]/NET0131 , \u5_burst_cnt_reg[7]/NET0131 , \u5_burst_cnt_reg[8]/NET0131 , \u5_burst_cnt_reg[9]/NET0131 , \u5_cke_o_del_reg/P0001 , \u5_cke_r_reg/NET0131 , \u5_cmd_a10_r_reg/P0001 , \u5_cmd_asserted2_reg/NET0131 , \u5_cmd_asserted_reg/NET0131 , \u5_cmd_del_reg[0]/NET0131 , \u5_cmd_del_reg[1]/NET0131 , \u5_cmd_del_reg[2]/NET0131 , \u5_cmd_del_reg[3]/NET0131 , \u5_cnt_reg/NET0131 , \u5_cs_le_r_reg/P0001 , \u5_cs_le_reg/P0001 , \u5_data_oe_r2_reg/NET0131 , \u5_data_oe_reg/NET0131 , \u5_dv_r_reg/NET0131 , \u5_ir_cnt_done_reg/P0001 , \u5_ir_cnt_reg[0]/P0001 , \u5_ir_cnt_reg[1]/P0001 , \u5_ir_cnt_reg[2]/P0001 , \u5_ir_cnt_reg[3]/P0001 , \u5_lmr_ack_reg/NET0131 , \u5_lookup_ready1_reg/NET0131 , \u5_lookup_ready2_reg/NET0131 , \u5_mc_adv_r1_reg/NET0131 , \u5_mc_adv_r_reg/NET0131 , \u5_mc_c_oe_reg/NET0131 , \u5_mc_le_reg/NET0131 , \u5_mem_ack_r_reg/NET0131 , \u5_no_wb_cycle_reg/NET0131 , \u5_oe__reg/NET0131 , \u5_pack_le0_reg/P0001 , \u5_pack_le1_reg/P0001 , \u5_resume_req_r_reg/NET0131 , \u5_rfr_ack_r_reg/NET0131 , \u5_state_reg[0]/NET0131 , \u5_state_reg[10]/NET0131 , \u5_state_reg[11]/NET0131 , \u5_state_reg[12]/NET0131 , \u5_state_reg[13]/NET0131 , \u5_state_reg[14]/NET0131 , \u5_state_reg[15]/NET0131 , \u5_state_reg[16]/NET0131 , \u5_state_reg[17]/NET0131 , \u5_state_reg[18]/NET0131 , \u5_state_reg[19]/NET0131 , \u5_state_reg[1]/NET0131 , \u5_state_reg[20]/NET0131 , \u5_state_reg[21]/NET0131 , \u5_state_reg[22]/NET0131 , \u5_state_reg[23]/NET0131 , \u5_state_reg[24]/NET0131 , \u5_state_reg[25]/NET0131 , \u5_state_reg[26]/NET0131 , \u5_state_reg[27]/NET0131 , \u5_state_reg[28]/NET0131 , \u5_state_reg[29]/NET0131 , \u5_state_reg[2]/NET0131 , \u5_state_reg[30]/NET0131 , \u5_state_reg[31]/NET0131 , \u5_state_reg[32]/NET0131 , \u5_state_reg[33]/NET0131 , \u5_state_reg[34]/NET0131 , \u5_state_reg[35]/NET0131 , \u5_state_reg[36]/NET0131 , \u5_state_reg[37]/NET0131 , \u5_state_reg[38]/NET0131 , \u5_state_reg[39]/NET0131 , \u5_state_reg[3]/NET0131 , \u5_state_reg[40]/NET0131 , \u5_state_reg[41]/NET0131 , \u5_state_reg[42]/NET0131 , \u5_state_reg[43]/NET0131 , \u5_state_reg[44]/NET0131 , \u5_state_reg[45]/NET0131 , \u5_state_reg[46]/NET0131 , \u5_state_reg[47]/NET0131 , \u5_state_reg[48]/NET0131 , \u5_state_reg[49]/NET0131 , \u5_state_reg[4]/NET0131 , \u5_state_reg[50]/NET0131 , \u5_state_reg[51]/NET0131 , \u5_state_reg[52]/NET0131 , \u5_state_reg[53]/NET0131 , \u5_state_reg[54]/NET0131 , \u5_state_reg[55]/NET0131 , \u5_state_reg[56]/NET0131 , \u5_state_reg[57]/NET0131 , \u5_state_reg[58]/NET0131 , \u5_state_reg[59]/NET0131 , \u5_state_reg[5]/NET0131 , \u5_state_reg[60]/NET0131 , \u5_state_reg[61]/NET0131 , \u5_state_reg[62]/NET0131 , \u5_state_reg[63]/NET0131 , \u5_state_reg[64]/NET0131 , \u5_state_reg[65]/NET0131 , \u5_state_reg[6]/NET0131 , \u5_state_reg[7]/NET0131 , \u5_state_reg[8]/NET0131 , \u5_state_reg[9]/NET0131 , \u5_susp_req_r_reg/NET0131 , \u5_susp_sel_r_reg/NET0131 , \u5_timer2_reg[0]/P0001 , \u5_timer2_reg[1]/P0001 , \u5_timer2_reg[2]/P0001 , \u5_timer2_reg[3]/P0001 , \u5_timer2_reg[4]/P0001 , \u5_timer2_reg[5]/P0001 , \u5_timer2_reg[6]/P0001 , \u5_timer2_reg[7]/P0001 , \u5_timer2_reg[8]/P0001 , \u5_timer_reg[0]/NET0131 , \u5_timer_reg[1]/NET0131 , \u5_timer_reg[2]/NET0131 , \u5_timer_reg[3]/NET0131 , \u5_timer_reg[4]/NET0131 , \u5_timer_reg[5]/NET0131 , \u5_timer_reg[6]/NET0131 , \u5_timer_reg[7]/NET0131 , \u5_tmr2_done_reg/NET0131 , \u5_tmr_done_reg/NET0131 , \u5_wb_cycle_reg/NET0131 , \u5_wb_stb_first_reg/NET0131 , \u5_wb_wait_r_reg/P0001 , \u5_wb_write_go_r_reg/NET0131 , \u5_wr_cycle_reg/NET0131 , \u6_read_go_r1_reg/NET0131 , \u6_read_go_r_reg/NET0131 , \u6_rmw_en_reg/NET0131 , \u6_rmw_r_reg/NET0131 , \u6_wb_first_r_reg/NET0131 , \u6_wr_hold_reg/NET0131 , \u6_write_go_r1_reg/NET0131 , \u6_write_go_r_reg/NET0131 , \u7_mc_ack_r_reg/NET0131 , \u7_mc_br_r_reg/P0001 , \u7_mc_data_ir_reg[0]/P0001 , \u7_mc_data_ir_reg[10]/P0001 , \u7_mc_data_ir_reg[11]/P0001 , \u7_mc_data_ir_reg[12]/P0001 , \u7_mc_data_ir_reg[13]/P0001 , \u7_mc_data_ir_reg[14]/P0001 , \u7_mc_data_ir_reg[15]/P0001 , \u7_mc_data_ir_reg[16]/P0001 , \u7_mc_data_ir_reg[17]/P0001 , \u7_mc_data_ir_reg[18]/P0001 , \u7_mc_data_ir_reg[19]/P0001 , \u7_mc_data_ir_reg[1]/P0001 , \u7_mc_data_ir_reg[20]/P0001 , \u7_mc_data_ir_reg[21]/P0001 , \u7_mc_data_ir_reg[22]/P0001 , \u7_mc_data_ir_reg[23]/P0001 , \u7_mc_data_ir_reg[24]/P0001 , \u7_mc_data_ir_reg[25]/P0001 , \u7_mc_data_ir_reg[26]/P0001 , \u7_mc_data_ir_reg[27]/P0001 , \u7_mc_data_ir_reg[28]/P0001 , \u7_mc_data_ir_reg[29]/P0001 , \u7_mc_data_ir_reg[2]/P0001 , \u7_mc_data_ir_reg[30]/P0001 , \u7_mc_data_ir_reg[31]/P0001 , \u7_mc_data_ir_reg[3]/P0001 , \u7_mc_data_ir_reg[4]/P0001 , \u7_mc_data_ir_reg[5]/P0001 , \u7_mc_data_ir_reg[6]/P0001 , \u7_mc_data_ir_reg[7]/P0001 , \u7_mc_data_ir_reg[8]/P0001 , \u7_mc_data_ir_reg[9]/P0001 , \u7_mc_dqm_r2_reg[0]/P0001 , \u7_mc_dqm_r2_reg[1]/P0001 , \u7_mc_dqm_r2_reg[2]/P0001 , \u7_mc_dqm_r2_reg[3]/P0001 , \u7_mc_dqm_r_reg[0]/P0001 , \u7_mc_dqm_r_reg[1]/P0001 , \u7_mc_dqm_r_reg[2]/P0001 , \u7_mc_dqm_r_reg[3]/P0001 , wb_ack_o_pad, \wb_addr_i[0]_pad , \wb_addr_i[10]_pad , \wb_addr_i[11]_pad , \wb_addr_i[12]_pad , \wb_addr_i[13]_pad , \wb_addr_i[14]_pad , \wb_addr_i[15]_pad , \wb_addr_i[16]_pad , \wb_addr_i[17]_pad , \wb_addr_i[18]_pad , \wb_addr_i[19]_pad , \wb_addr_i[1]_pad , \wb_addr_i[20]_pad , \wb_addr_i[21]_pad , \wb_addr_i[22]_pad , \wb_addr_i[23]_pad , \wb_addr_i[24]_pad , \wb_addr_i[25]_pad , \wb_addr_i[26]_pad , \wb_addr_i[27]_pad , \wb_addr_i[28]_pad , \wb_addr_i[29]_pad , \wb_addr_i[2]_pad , \wb_addr_i[30]_pad , \wb_addr_i[31]_pad , \wb_addr_i[3]_pad , \wb_addr_i[4]_pad , \wb_addr_i[5]_pad , \wb_addr_i[6]_pad , \wb_addr_i[7]_pad , \wb_addr_i[8]_pad , \wb_addr_i[9]_pad , wb_cyc_i_pad, \wb_data_i[0]_pad , \wb_data_i[10]_pad , \wb_data_i[11]_pad , \wb_data_i[12]_pad , \wb_data_i[13]_pad , \wb_data_i[14]_pad , \wb_data_i[15]_pad , \wb_data_i[16]_pad , \wb_data_i[17]_pad , \wb_data_i[18]_pad , \wb_data_i[19]_pad , \wb_data_i[1]_pad , \wb_data_i[20]_pad , \wb_data_i[21]_pad , \wb_data_i[22]_pad , \wb_data_i[23]_pad , \wb_data_i[24]_pad , \wb_data_i[25]_pad , \wb_data_i[26]_pad , \wb_data_i[27]_pad , \wb_data_i[28]_pad , \wb_data_i[29]_pad , \wb_data_i[2]_pad , \wb_data_i[30]_pad , \wb_data_i[31]_pad , \wb_data_i[3]_pad , \wb_data_i[4]_pad , \wb_data_i[5]_pad , \wb_data_i[6]_pad , \wb_data_i[7]_pad , \wb_data_i[8]_pad , \wb_data_i[9]_pad , wb_err_o_pad, \wb_sel_i[0]_pad , \wb_sel_i[1]_pad , \wb_sel_i[2]_pad , \wb_sel_i[3]_pad , wb_stb_i_pad, wb_we_i_pad, \_al_n0 , \_al_n1 , \g22/_0_ , \g23/_0_ , \g25_dup61718/_2_ , \g43466/_0_ , \g43467/_0_ , \g43468/_0_ , \g43469/_0_ , \g43470/_0_ , \g43471/_0_ , \g43472/_0_ , \g43473/_0_ , \g43474/_0_ , \g43475/_0_ , \g43476/_0_ , \g43477/_0_ , \g43478/_0_ , \g43512/_0_ , \g43513/_0_ , \g43544/_3_ , \g43545/_0_ , \g43554/_0_ , \g43555/_0_ , \g43557/_0_ , \g43558/_0_ , \g43571/_2_ , \g43632/_0_ , \g43633/_0_ , \g43635/_0_ , \g43636/_0_ , \g43637/_0_ , \g43638/_0_ , \g43639/_0_ , \g43640/_0_ , \g43642/_0_ , \g43662/_0_ , \g43663/_0_ , \g43664/_0_ , \g43665/_0_ , \g43668/_0_ , \g43670/_0_ , \g43671/_0_ , \g43673/_0_ , \g43674/_0_ , \g43692/_0_ , \g43695/_0_ , \g43696/_0_ , \g43697/_0_ , \g43698/_0_ , \g43700/_0_ , \g43701/_0_ , \g43703/_0_ , \g43705/_0_ , \g43707/_0_ , \g43708/_0_ , \g43710/_0_ , \g43717/_0_ , \g43719/_0_ , \g43720/_0_ , \g43721/_0_ , \g43722/_1_ , \g43723/_0_ , \g43725/_0_ , \g43729/_0_ , \g43731/_0_ , \g43734/_0_ , \g43735/_0_ , \g43737/_0_ , \g43744/_0_ , \g43747/_0_ , \g43760/_2_ , \g43770/_1_ , \g43775/_2_ , \g43780/_2_ , \g43786/_0_ , \g43787/_1_ , \g43847/_0_ , \g43848/_1_ , \g43858/_1_ , \g43891/_3_ , \g43895/_0_ , \g43934/_0_ , \g43936/_3_ , \g43954/_3_ , \g43961/_0_ , \g44016/_1_ , \g44067/_0_ , \g44094/_0_ , \g44096/_0_ , \g44104/_0_ , \g44122/_0_ , \g44172/_0_ , \g44209/_0_ , \g44219/_0_ , \g44220/_0_ , \g44222/_0_ , \g44223/_0_ , \g44241/_2_ , \g44252/_0_ , \g44253/_0_ , \g44255/_2_ , \g44263/_2_ , \g44470/_0_ , \g44538/_0_ , \g44539/_0_ , \g44540/_0_ , \g44541/_0_ , \g44542/_0_ , \g44543/_0_ , \g44544/_0_ , \g44545/_0_ , \g44546/_0_ , \g44547/_0_ , \g44548/_0_ , \g44549/_0_ , \g44550/_0_ , \g44551/_0_ , \g44552/_0_ , \g44553/_0_ , \g44554/_0_ , \g44555/_0_ , \g44556/_0_ , \g44557/_0_ , \g44558/_0_ , \g44559/_0_ , \g44560/_0_ , \g44561/_0_ , \g44562/_0_ , \g44563/_0_ , \g44564/_0_ , \g44565/_0_ , \g44566/_0_ , \g44567/_0_ , \g44568/_0_ , \g44569/_0_ , \g44570/_0_ , \g44571/_0_ , \g44572/_0_ , \g44573/_0_ , \g44574/_0_ , \g44575/_0_ , \g44576/_0_ , \g44577/_0_ , \g44578/_0_ , \g44579/_0_ , \g44580/_0_ , \g44581/_0_ , \g44582/_0_ , \g44583/_0_ , \g44584/_0_ , \g44585/_0_ , \g44586/_0_ , \g44588/_0_ , \g44589/_0_ , \g44590/_0_ , \g44591/_0_ , \g44592/_0_ , \g44593/_0_ , \g44594/_0_ , \g44595/_0_ , \g44596/_0_ , \g44636/_2_ , \g44646/_0_ , \g44647/_0_ , \g44648/_0_ , \g44649/_0_ , \g44650/_0_ , \g44651/_0_ , \g44652/_0_ , \g44653/_0_ , \g44654/_0_ , \g44655/_0_ , \g44656/_0_ , \g44657/_0_ , \g44665/_0_ , \g44666/_0_ , \g44667/_0_ , \g44668/_0_ , \g44752/_0_ , \g44753/_0_ , \g44873/_0_ , \g44939/_0_ , \g44942/_0_ , \g44945/_0_ , \g45023/_2_ , \g45090/_0_ , \g45141/_0_ , \g45147/_3_ , \g45155/_0_ , \g45190/_0_ , \g45195/_2_ , \g45199/_2_ , \g45201/_2_ , \g45324/_0_ , \g45334/_2_ , \g45336/_0_ , \g45388/_0_ , \g45391/_0_ , \g45413/_2_ , \g45530/_0_ , \g45532/_0_ , \g45533/_0_ , \g45534/_0_ , \g45739/_2_ , \g45743/_2_ , \g45767/_0_ , \g45782/_0_ , \g45830/_3_ , \g45834/_3_ , \g45835/_3_ , \g45836/_3_ , \g45837/_3_ , \g45839/_3_ , \g45840/_3_ , \g45841/_3_ , \g45842/_3_ , \g45843/_3_ , \g45844/_3_ , \g45845/_3_ , \g46191/_0_ , \g46193/_3_ , \g46256/_3_ , \g46257/_3_ , \g46258/_3_ , \g46259/_3_ , \g46260/_3_ , \g46261/_3_ , \g46262/_3_ , \g46263/_3_ , \g46278/_0_ , \g46292/_0_ , \g46293/_0_ , \g46312/_0_ , \g46367/_2_ , \g46370/_2_ , \g46380/_2_ , \g46386/_2_ , \g46388/_2_ , \g46392/_2_ , \g46395/_2_ , \g46399/_2_ , \g46420/_0_ , \g46446/_0_ , \g46493/_0_ , \g46510/_0_ , \g46669/_2_ , \g46691/_0_ , \g46708/_0_ , \g46721/_00_ , \g46776/_0_ , \g46777/_0_ , \g46778/_0_ , \g46779/_0_ , \g46780/_0_ , \g46782/_0_ , \g46784/_0_ , \g46932/_0_ , \g47112/_0_ , \g47124/_0_ , \g47265/_0_ , \g47270/_0_ , \g47275/_0_ , \g47300/_1_ , \g47305/_1_ , \g47338/_0_ , \g47339/_0_ , \g47352/_0_ , \g47699/_3_ , \g47711/_0_ , \g47719/_3_ , \g47721/_3_ , \g47723/_3_ , \g47853/_0_ , \g48094/_0_ , \g48095/_0_ , \g48177/_2_ , \g48194/_0_ , \g48369/_2_ , \g48371/_2_ , \g48373/_2_ , \g48375/_2_ , \g48377/_2_ , \g48379/_2_ , \g48381/_2_ , \g48383/_2_ , \g48385/_2_ , \g48535/_0_ , \g48569/_0_ , \g48570/_0_ , \g48571/_0_ , \g48836/_0_ , \g48843/_0_ , \g49187/_3_ , \g49375/_2_ , \g49633/_0_ , \g49788/_1_ , \g49800/_1_ , \g49802/_1_ , \g49806/_1_ , \g49853/_1_ , \g49883/_0_ , \g49884/_0_ , \g49885/_0_ , \g49886/_0_ , \g49976/_1_ , \g50038/_0_ , \g50082/_0_ , \g50083/_0_ , \g50167/_3_ , \g50168/_3_ , \g50169/_3_ , \g50170/_3_ , \g50171/_3_ , \g50177/_0_ , \g50190/_0_ , \g50236/_0_ , \g50251/_3_ , \g50256/_0_ , \g50318/_3_ , \g50319/_3_ , \g50350/_3_ , \g50351/_3_ , \g50352/_3_ , \g50353/_3_ , \g50354/_3_ , \g50355/_3_ , \g50361/_2_ , \g50366/_0_ , \g50393/_0_ , \g50552/_1_ , \g51108/_0_ , \g51160/_0_ , \g51290/_1_ , \g51327/_3_ , \g51328/_3_ , \g51329/_3_ , \g51330/_3_ , \g51331/_3_ , \g51332/_3_ , \g51333/_3_ , \g51334/_3_ , \g51339/_3_ , \g51340/_3_ , \g51341/_3_ , \g51342/_3_ , \g51343/_3_ , \g51346/_0_ , \g51347/_0_ , \g51348/_0_ , \g51381/_3_ , \g51382/_3_ , \g51383/_3_ , \g51386/_3_ , \g51387/_3_ , \g51405/_3_ , \g51410/_3_ , \g51883/_0_ , \g51916/_0_ , \g51947/_0_ , \g51948/_0_ , \g51949/_0_ , \g51950/_0_ , \g51951/_0_ , \g51952/_0_ , \g51953/_0_ , \g51954/_0_ , \g51955/_0_ , \g51956/_0_ , \g51957/_0_ , \g51958/_0_ , \g51959/_0_ , \g51960/_0_ , \g51961/_0_ , \g51962/_0_ , \g51963/_0_ , \g51964/_0_ , \g51965/_0_ , \g51967/_0_ , \g51968/_0_ , \g51969/_0_ , \g51970/_0_ , \g51971/_0_ , \g51972/_0_ , \g51973/_0_ , \g51974/_0_ , \g51975/_0_ , \g51976/_0_ , \g51977/_0_ , \g51978/_0_ , \g51979/_0_ , \g51980/_0_ , \g51981/_0_ , \g51982/_0_ , \g51983/_0_ , \g51984/_0_ , \g51985/_0_ , \g51986/_0_ , \g51987/_0_ , \g51988/_0_ , \g51989/_0_ , \g51990/_0_ , \g51991/_0_ , \g51992/_0_ , \g51993/_0_ , \g51994/_0_ , \g51995/_0_ , \g51996/_0_ , \g51997/_0_ , \g51998/_0_ , \g51999/_0_ , \g52000/_0_ , \g52001/_0_ , \g52002/_0_ , \g52003/_0_ , \g52004/_0_ , \g52005/_0_ , \g52006/_0_ , \g52007/_0_ , \g52008/_0_ , \g52009/_0_ , \g52010/_0_ , \g52011/_0_ , \g52012/_0_ , \g52013/_0_ , \g52014/_0_ , \g52015/_0_ , \g52016/_0_ , \g52017/_0_ , \g52018/_0_ , \g52019/_0_ , \g52020/_0_ , \g52021/_0_ , \g52022/_0_ , \g52023/_0_ , \g52024/_0_ , \g52025/_0_ , \g52026/_0_ , \g52027/_0_ , \g52028/_0_ , \g52029/_0_ , \g52030/_0_ , \g52031/_0_ , \g52032/_0_ , \g52033/_0_ , \g52034/_0_ , \g52035/_0_ , \g52036/_0_ , \g52037/_0_ , \g52038/_0_ , \g52039/_0_ , \g52040/_0_ , \g52041/_0_ , \g52042/_0_ , \g52043/_0_ , \g52044/_0_ , \g52045/_0_ , \g52046/_0_ , \g52047/_0_ , \g52049/_0_ , \g52050/_0_ , \g52051/_0_ , \g52052/_0_ , \g52053/_0_ , \g52054/_0_ , \g52055/_0_ , \g52056/_0_ , \g52057/_0_ , \g52058/_0_ , \g52061/_0_ , \g52065/_0_ , \g52066/_0_ , \g52067/_0_ , \g52068/_0_ , \g52069/_0_ , \g52070/_0_ , \g52071/_0_ , \g52073/_0_ , \g52074/_0_ , \g52075/_0_ , \g52082/_0_ , \g52083/_0_ , \g52158/_0_ , \g52201/_0_ , \g52202/_0_ , \g52346/_0_ , \g52351/_0_ , \g52390/_0_ , \g52847/_0_ , \g52854/_0_ , \g52968/_0_ , \g52969/_0_ , \g52970/_0_ , \g52971/_0_ , \g52984/_0_ , \g52994/_0_ , \g53019/_0_ , \g53030/_0_ , \g53094/_1_ , \g53106/_0_ , \g53150/_0_ , \g53256/_0_ , \g53297/_0_ , \g53345/_0_ , \g53359/_0_ , \g53375/_0_ , \g53474/_1__syn_2 , \g53475/_2_ , \g53593/_0_ , \g53643/_1_ , \g53655/_0_ , \g53710/_0_ , \g53786/_0_ , \g53837/_0_ , \g53888/_1_ , \g53909/_0_ , \g54253/_2_ , \g54394/_3_ , \g54413/_0_ , \g55420/_0_ , \g55587/_0_ , \g55852/_0_ , \g57020/_0_ , \g59450/_0_ , \g59488/_2_ , \g59752/_0_ , \g59786/_0_ , \g59854/_0_ , \g59878/_0_ , \g59902/_0_ , \g59924/_0_ , \g59947/_0_ , \g59972/_0_ , \g59996/_0_ , \g60017/_0_ , \g60040/_0_ , \g60064/_0_ , \g60095/_0_ , \g60119/_0_ , \g60145/_1_ , \g60165/_0_ , \g60407/_2_ , \g60408/_0_ , \g60613/_2_ , \g60649/_0_ , \g60771/_0_ , \g60908/_1_ , \g60911/_0_ , \g60977/_0_ , \g61/_0_ , \g61002/_0_ , \g61308/_0_ , \g61312/_1_ , \g61314/_0_ , \g61319/_1_ , \g61342/_1_ , \g61360/_0_ , \g61377/_0_ , \g61423/_1_ , \g61426/_0_ , \g61479/_1_ , \g61523/_1_ , \g61558/_1_ , \g61652/_0_ , \g61866/_0_ , \g61868/_1_ , \g61887/_0_ , \u7_mc_dqm_r_reg[0]/P0001_reg_syn_3 , \u7_mc_dqm_r_reg[1]/P0001_reg_syn_3 , \u7_mc_dqm_r_reg[2]/P0001_reg_syn_3 , \u7_mc_dqm_r_reg[3]/P0001_reg_syn_3 , \u7_mc_we__reg/_05_ );
	input mc_cke_pad_o__pad ;
	input mc_vpen_pad_o_pad ;
	input \mem_ack_r_reg/P0001  ;
	input \poc_o[0]_pad  ;
	input \poc_o[10]_pad  ;
	input \poc_o[11]_pad  ;
	input \poc_o[12]_pad  ;
	input \poc_o[13]_pad  ;
	input \poc_o[14]_pad  ;
	input \poc_o[15]_pad  ;
	input \poc_o[16]_pad  ;
	input \poc_o[17]_pad  ;
	input \poc_o[18]_pad  ;
	input \poc_o[19]_pad  ;
	input \poc_o[1]_pad  ;
	input \poc_o[20]_pad  ;
	input \poc_o[21]_pad  ;
	input \poc_o[22]_pad  ;
	input \poc_o[23]_pad  ;
	input \poc_o[24]_pad  ;
	input \poc_o[25]_pad  ;
	input \poc_o[26]_pad  ;
	input \poc_o[27]_pad  ;
	input \poc_o[28]_pad  ;
	input \poc_o[29]_pad  ;
	input \poc_o[2]_pad  ;
	input \poc_o[30]_pad  ;
	input \poc_o[31]_pad  ;
	input \poc_o[3]_pad  ;
	input \poc_o[4]_pad  ;
	input \poc_o[5]_pad  ;
	input \poc_o[6]_pad  ;
	input \poc_o[7]_pad  ;
	input \poc_o[8]_pad  ;
	input \poc_o[9]_pad  ;
	input suspended_o_pad ;
	input \u0_cs_reg[0]/NET0131  ;
	input \u0_cs_reg[1]/NET0131  ;
	input \u0_csc_mask_r_reg[0]/NET0131  ;
	input \u0_csc_mask_r_reg[10]/NET0131  ;
	input \u0_csc_mask_r_reg[1]/NET0131  ;
	input \u0_csc_mask_r_reg[2]/NET0131  ;
	input \u0_csc_mask_r_reg[3]/NET0131  ;
	input \u0_csc_mask_r_reg[4]/NET0131  ;
	input \u0_csc_mask_r_reg[5]/NET0131  ;
	input \u0_csc_mask_r_reg[6]/NET0131  ;
	input \u0_csc_mask_r_reg[7]/NET0131  ;
	input \u0_csc_mask_r_reg[8]/NET0131  ;
	input \u0_csc_mask_r_reg[9]/NET0131  ;
	input \u0_csc_reg[10]/NET0131  ;
	input \u0_csc_reg[11]/NET0131  ;
	input \u0_csc_reg[1]/NET0131  ;
	input \u0_csc_reg[2]/NET0131  ;
	input \u0_csc_reg[3]/NET0131  ;
	input \u0_csc_reg[4]/NET0131  ;
	input \u0_csc_reg[5]/NET0131  ;
	input \u0_csc_reg[6]/NET0131  ;
	input \u0_csc_reg[7]/NET0131  ;
	input \u0_csc_reg[9]/NET0131  ;
	input \u0_csr_r2_reg[0]/NET0131  ;
	input \u0_csr_r2_reg[1]/NET0131  ;
	input \u0_csr_r2_reg[2]/NET0131  ;
	input \u0_csr_r2_reg[3]/NET0131  ;
	input \u0_csr_r2_reg[4]/NET0131  ;
	input \u0_csr_r2_reg[5]/NET0131  ;
	input \u0_csr_r2_reg[6]/NET0131  ;
	input \u0_csr_r2_reg[7]/NET0131  ;
	input \u0_csr_r_reg[0]/P0001  ;
	input \u0_csr_r_reg[10]/NET0131  ;
	input \u0_csr_r_reg[2]/NET0131  ;
	input \u0_csr_r_reg[3]/NET0131  ;
	input \u0_csr_r_reg[4]/NET0131  ;
	input \u0_csr_r_reg[5]/NET0131  ;
	input \u0_csr_r_reg[6]/NET0131  ;
	input \u0_csr_r_reg[7]/NET0131  ;
	input \u0_csr_r_reg[8]/NET0131  ;
	input \u0_csr_r_reg[9]/NET0131  ;
	input \u0_init_ack_r_reg/P0001  ;
	input \u0_init_req_reg/NET0131  ;
	input \u0_lmr_ack_r_reg/P0001  ;
	input \u0_lmr_req_reg/NET0131  ;
	input \u0_rf_we_reg/NET0131  ;
	input \u0_rst_r2_reg/NET0131  ;
	input \u0_sp_csc_reg[10]/NET0131  ;
	input \u0_sp_csc_reg[1]/NET0131  ;
	input \u0_sp_csc_reg[2]/NET0131  ;
	input \u0_sp_csc_reg[3]/NET0131  ;
	input \u0_sp_csc_reg[4]/NET0131  ;
	input \u0_sp_csc_reg[5]/NET0131  ;
	input \u0_sp_csc_reg[6]/NET0131  ;
	input \u0_sp_csc_reg[7]/NET0131  ;
	input \u0_sp_csc_reg[9]/NET0131  ;
	input \u0_sp_tms_reg[0]/NET0131  ;
	input \u0_sp_tms_reg[10]/NET0131  ;
	input \u0_sp_tms_reg[11]/NET0131  ;
	input \u0_sp_tms_reg[12]/NET0131  ;
	input \u0_sp_tms_reg[13]/NET0131  ;
	input \u0_sp_tms_reg[14]/NET0131  ;
	input \u0_sp_tms_reg[15]/NET0131  ;
	input \u0_sp_tms_reg[16]/NET0131  ;
	input \u0_sp_tms_reg[17]/NET0131  ;
	input \u0_sp_tms_reg[18]/NET0131  ;
	input \u0_sp_tms_reg[19]/NET0131  ;
	input \u0_sp_tms_reg[1]/NET0131  ;
	input \u0_sp_tms_reg[20]/NET0131  ;
	input \u0_sp_tms_reg[21]/NET0131  ;
	input \u0_sp_tms_reg[22]/NET0131  ;
	input \u0_sp_tms_reg[23]/NET0131  ;
	input \u0_sp_tms_reg[24]/NET0131  ;
	input \u0_sp_tms_reg[25]/NET0131  ;
	input \u0_sp_tms_reg[26]/NET0131  ;
	input \u0_sp_tms_reg[27]/NET0131  ;
	input \u0_sp_tms_reg[2]/NET0131  ;
	input \u0_sp_tms_reg[3]/NET0131  ;
	input \u0_sp_tms_reg[4]/NET0131  ;
	input \u0_sp_tms_reg[5]/NET0131  ;
	input \u0_sp_tms_reg[6]/NET0131  ;
	input \u0_sp_tms_reg[7]/NET0131  ;
	input \u0_sp_tms_reg[8]/NET0131  ;
	input \u0_sp_tms_reg[9]/NET0131  ;
	input \u0_spec_req_cs_reg[0]/NET0131  ;
	input \u0_spec_req_cs_reg[1]/NET0131  ;
	input \u0_sreq_cs_le_reg/NET0131  ;
	input \u0_tms_reg[0]/NET0131  ;
	input \u0_tms_reg[10]/NET0131  ;
	input \u0_tms_reg[11]/NET0131  ;
	input \u0_tms_reg[12]/NET0131  ;
	input \u0_tms_reg[13]/NET0131  ;
	input \u0_tms_reg[14]/NET0131  ;
	input \u0_tms_reg[15]/NET0131  ;
	input \u0_tms_reg[16]/NET0131  ;
	input \u0_tms_reg[17]/NET0131  ;
	input \u0_tms_reg[18]/NET0131  ;
	input \u0_tms_reg[19]/NET0131  ;
	input \u0_tms_reg[1]/NET0131  ;
	input \u0_tms_reg[20]/NET0131  ;
	input \u0_tms_reg[21]/NET0131  ;
	input \u0_tms_reg[22]/NET0131  ;
	input \u0_tms_reg[23]/NET0131  ;
	input \u0_tms_reg[24]/NET0131  ;
	input \u0_tms_reg[25]/NET0131  ;
	input \u0_tms_reg[26]/NET0131  ;
	input \u0_tms_reg[27]/NET0131  ;
	input \u0_tms_reg[2]/NET0131  ;
	input \u0_tms_reg[3]/NET0131  ;
	input \u0_tms_reg[4]/NET0131  ;
	input \u0_tms_reg[5]/NET0131  ;
	input \u0_tms_reg[6]/NET0131  ;
	input \u0_tms_reg[7]/NET0131  ;
	input \u0_tms_reg[8]/NET0131  ;
	input \u0_tms_reg[9]/NET0131  ;
	input \u0_u0_addr_r_reg[2]/P0001  ;
	input \u0_u0_addr_r_reg[3]/P0001  ;
	input \u0_u0_addr_r_reg[4]/P0001  ;
	input \u0_u0_addr_r_reg[5]/P0001  ;
	input \u0_u0_addr_r_reg[6]/P0001  ;
	input \u0_u0_csc_reg[0]/NET0131  ;
	input \u0_u0_csc_reg[10]/P0001  ;
	input \u0_u0_csc_reg[11]/P0001  ;
	input \u0_u0_csc_reg[12]/P0001  ;
	input \u0_u0_csc_reg[13]/P0001  ;
	input \u0_u0_csc_reg[14]/P0001  ;
	input \u0_u0_csc_reg[15]/P0001  ;
	input \u0_u0_csc_reg[16]/P0001  ;
	input \u0_u0_csc_reg[17]/P0001  ;
	input \u0_u0_csc_reg[18]/P0001  ;
	input \u0_u0_csc_reg[19]/P0001  ;
	input \u0_u0_csc_reg[1]/NET0131  ;
	input \u0_u0_csc_reg[20]/P0001  ;
	input \u0_u0_csc_reg[21]/P0001  ;
	input \u0_u0_csc_reg[22]/P0001  ;
	input \u0_u0_csc_reg[23]/P0001  ;
	input \u0_u0_csc_reg[24]/P0001  ;
	input \u0_u0_csc_reg[25]/P0001  ;
	input \u0_u0_csc_reg[26]/P0001  ;
	input \u0_u0_csc_reg[27]/P0001  ;
	input \u0_u0_csc_reg[28]/P0001  ;
	input \u0_u0_csc_reg[29]/P0001  ;
	input \u0_u0_csc_reg[2]/NET0131  ;
	input \u0_u0_csc_reg[30]/P0001  ;
	input \u0_u0_csc_reg[31]/P0001  ;
	input \u0_u0_csc_reg[3]/NET0131  ;
	input \u0_u0_csc_reg[4]/P0001  ;
	input \u0_u0_csc_reg[5]/P0001  ;
	input \u0_u0_csc_reg[6]/P0001  ;
	input \u0_u0_csc_reg[7]/P0001  ;
	input \u0_u0_csc_reg[8]/P0001  ;
	input \u0_u0_csc_reg[9]/P0001  ;
	input \u0_u0_init_req_reg/NET0131  ;
	input \u0_u0_init_req_we_reg/NET0131  ;
	input \u0_u0_inited_reg/NET0131  ;
	input \u0_u0_lmr_req_reg/NET0131  ;
	input \u0_u0_lmr_req_we_reg/NET0131  ;
	input \u0_u0_tms_reg[0]/P0001  ;
	input \u0_u0_tms_reg[10]/P0001  ;
	input \u0_u0_tms_reg[11]/P0001  ;
	input \u0_u0_tms_reg[12]/P0001  ;
	input \u0_u0_tms_reg[13]/P0001  ;
	input \u0_u0_tms_reg[14]/P0001  ;
	input \u0_u0_tms_reg[15]/P0001  ;
	input \u0_u0_tms_reg[16]/P0001  ;
	input \u0_u0_tms_reg[17]/P0001  ;
	input \u0_u0_tms_reg[18]/P0001  ;
	input \u0_u0_tms_reg[19]/P0001  ;
	input \u0_u0_tms_reg[1]/P0001  ;
	input \u0_u0_tms_reg[20]/P0001  ;
	input \u0_u0_tms_reg[21]/P0001  ;
	input \u0_u0_tms_reg[22]/P0001  ;
	input \u0_u0_tms_reg[23]/P0001  ;
	input \u0_u0_tms_reg[24]/P0001  ;
	input \u0_u0_tms_reg[25]/P0001  ;
	input \u0_u0_tms_reg[26]/P0001  ;
	input \u0_u0_tms_reg[27]/P0001  ;
	input \u0_u0_tms_reg[28]/P0001  ;
	input \u0_u0_tms_reg[29]/P0001  ;
	input \u0_u0_tms_reg[2]/P0001  ;
	input \u0_u0_tms_reg[30]/P0001  ;
	input \u0_u0_tms_reg[31]/P0001  ;
	input \u0_u0_tms_reg[3]/P0001  ;
	input \u0_u0_tms_reg[4]/P0001  ;
	input \u0_u0_tms_reg[5]/P0001  ;
	input \u0_u0_tms_reg[6]/P0001  ;
	input \u0_u0_tms_reg[7]/P0001  ;
	input \u0_u0_tms_reg[8]/P0001  ;
	input \u0_u0_tms_reg[9]/P0001  ;
	input \u0_u1_csc_reg[0]/NET0131  ;
	input \u0_u1_csc_reg[10]/P0001  ;
	input \u0_u1_csc_reg[11]/P0001  ;
	input \u0_u1_csc_reg[12]/P0001  ;
	input \u0_u1_csc_reg[13]/P0001  ;
	input \u0_u1_csc_reg[14]/P0001  ;
	input \u0_u1_csc_reg[15]/P0001  ;
	input \u0_u1_csc_reg[16]/P0001  ;
	input \u0_u1_csc_reg[17]/P0001  ;
	input \u0_u1_csc_reg[18]/P0001  ;
	input \u0_u1_csc_reg[19]/P0001  ;
	input \u0_u1_csc_reg[1]/NET0131  ;
	input \u0_u1_csc_reg[20]/P0001  ;
	input \u0_u1_csc_reg[21]/P0001  ;
	input \u0_u1_csc_reg[22]/P0001  ;
	input \u0_u1_csc_reg[23]/P0001  ;
	input \u0_u1_csc_reg[24]/P0001  ;
	input \u0_u1_csc_reg[25]/P0001  ;
	input \u0_u1_csc_reg[26]/P0001  ;
	input \u0_u1_csc_reg[27]/P0001  ;
	input \u0_u1_csc_reg[28]/P0001  ;
	input \u0_u1_csc_reg[29]/P0001  ;
	input \u0_u1_csc_reg[2]/NET0131  ;
	input \u0_u1_csc_reg[30]/P0001  ;
	input \u0_u1_csc_reg[31]/P0001  ;
	input \u0_u1_csc_reg[3]/NET0131  ;
	input \u0_u1_csc_reg[4]/P0001  ;
	input \u0_u1_csc_reg[5]/P0001  ;
	input \u0_u1_csc_reg[6]/P0001  ;
	input \u0_u1_csc_reg[7]/P0001  ;
	input \u0_u1_csc_reg[8]/P0001  ;
	input \u0_u1_csc_reg[9]/P0001  ;
	input \u0_u1_init_req_reg/NET0131  ;
	input \u0_u1_init_req_we_reg/NET0131  ;
	input \u0_u1_inited_reg/NET0131  ;
	input \u0_u1_lmr_req_reg/NET0131  ;
	input \u0_u1_lmr_req_we_reg/NET0131  ;
	input \u0_u1_tms_reg[0]/P0001  ;
	input \u0_u1_tms_reg[10]/P0001  ;
	input \u0_u1_tms_reg[11]/P0001  ;
	input \u0_u1_tms_reg[12]/P0001  ;
	input \u0_u1_tms_reg[13]/P0001  ;
	input \u0_u1_tms_reg[14]/P0001  ;
	input \u0_u1_tms_reg[15]/P0001  ;
	input \u0_u1_tms_reg[16]/P0001  ;
	input \u0_u1_tms_reg[17]/P0001  ;
	input \u0_u1_tms_reg[18]/P0001  ;
	input \u0_u1_tms_reg[19]/P0001  ;
	input \u0_u1_tms_reg[1]/P0001  ;
	input \u0_u1_tms_reg[20]/P0001  ;
	input \u0_u1_tms_reg[21]/P0001  ;
	input \u0_u1_tms_reg[22]/P0001  ;
	input \u0_u1_tms_reg[23]/P0001  ;
	input \u0_u1_tms_reg[24]/P0001  ;
	input \u0_u1_tms_reg[25]/P0001  ;
	input \u0_u1_tms_reg[26]/P0001  ;
	input \u0_u1_tms_reg[27]/P0001  ;
	input \u0_u1_tms_reg[28]/P0001  ;
	input \u0_u1_tms_reg[29]/P0001  ;
	input \u0_u1_tms_reg[2]/P0001  ;
	input \u0_u1_tms_reg[30]/P0001  ;
	input \u0_u1_tms_reg[31]/P0001  ;
	input \u0_u1_tms_reg[3]/P0001  ;
	input \u0_u1_tms_reg[4]/P0001  ;
	input \u0_u1_tms_reg[5]/P0001  ;
	input \u0_u1_tms_reg[6]/P0001  ;
	input \u0_u1_tms_reg[7]/P0001  ;
	input \u0_u1_tms_reg[8]/P0001  ;
	input \u0_u1_tms_reg[9]/P0001  ;
	input \u0_wp_err_reg/NET0131  ;
	input \u1_acs_addr_reg[0]/P0001  ;
	input \u1_acs_addr_reg[10]/P0001  ;
	input \u1_acs_addr_reg[11]/P0001  ;
	input \u1_acs_addr_reg[12]/P0001  ;
	input \u1_acs_addr_reg[13]/P0001  ;
	input \u1_acs_addr_reg[14]/P0001  ;
	input \u1_acs_addr_reg[15]/P0001  ;
	input \u1_acs_addr_reg[16]/P0001  ;
	input \u1_acs_addr_reg[17]/P0001  ;
	input \u1_acs_addr_reg[18]/P0001  ;
	input \u1_acs_addr_reg[19]/P0001  ;
	input \u1_acs_addr_reg[1]/P0001  ;
	input \u1_acs_addr_reg[20]/P0001  ;
	input \u1_acs_addr_reg[21]/P0001  ;
	input \u1_acs_addr_reg[22]/P0001  ;
	input \u1_acs_addr_reg[23]/P0001  ;
	input \u1_acs_addr_reg[2]/P0001  ;
	input \u1_acs_addr_reg[3]/P0001  ;
	input \u1_acs_addr_reg[4]/P0001  ;
	input \u1_acs_addr_reg[5]/P0001  ;
	input \u1_acs_addr_reg[6]/P0001  ;
	input \u1_acs_addr_reg[7]/P0001  ;
	input \u1_acs_addr_reg[8]/P0001  ;
	input \u1_acs_addr_reg[9]/P0001  ;
	input \u1_bank_adr_reg[0]/P0001  ;
	input \u1_bank_adr_reg[1]/P0001  ;
	input \u1_col_adr_reg[0]/P0001  ;
	input \u1_col_adr_reg[1]/P0001  ;
	input \u1_col_adr_reg[2]/P0001  ;
	input \u1_col_adr_reg[3]/P0001  ;
	input \u1_col_adr_reg[4]/P0001  ;
	input \u1_col_adr_reg[5]/P0001  ;
	input \u1_col_adr_reg[6]/P0001  ;
	input \u1_col_adr_reg[7]/P0001  ;
	input \u1_col_adr_reg[8]/P0001  ;
	input \u1_col_adr_reg[9]/P0001  ;
	input \u1_row_adr_reg[0]/P0001  ;
	input \u1_row_adr_reg[10]/P0001  ;
	input \u1_row_adr_reg[11]/P0001  ;
	input \u1_row_adr_reg[12]/P0001  ;
	input \u1_row_adr_reg[1]/P0001  ;
	input \u1_row_adr_reg[2]/P0001  ;
	input \u1_row_adr_reg[3]/P0001  ;
	input \u1_row_adr_reg[4]/P0001  ;
	input \u1_row_adr_reg[5]/P0001  ;
	input \u1_row_adr_reg[6]/P0001  ;
	input \u1_row_adr_reg[7]/P0001  ;
	input \u1_row_adr_reg[8]/P0001  ;
	input \u1_row_adr_reg[9]/P0001  ;
	input \u1_sram_addr_reg[0]/P0001  ;
	input \u1_sram_addr_reg[10]/P0001  ;
	input \u1_sram_addr_reg[11]/P0001  ;
	input \u1_sram_addr_reg[12]/P0001  ;
	input \u1_sram_addr_reg[13]/P0001  ;
	input \u1_sram_addr_reg[14]/P0001  ;
	input \u1_sram_addr_reg[15]/P0001  ;
	input \u1_sram_addr_reg[16]/P0001  ;
	input \u1_sram_addr_reg[17]/P0001  ;
	input \u1_sram_addr_reg[18]/P0001  ;
	input \u1_sram_addr_reg[19]/P0001  ;
	input \u1_sram_addr_reg[1]/P0001  ;
	input \u1_sram_addr_reg[20]/P0001  ;
	input \u1_sram_addr_reg[21]/P0001  ;
	input \u1_sram_addr_reg[22]/P0001  ;
	input \u1_sram_addr_reg[23]/P0001  ;
	input \u1_sram_addr_reg[2]/P0001  ;
	input \u1_sram_addr_reg[3]/P0001  ;
	input \u1_sram_addr_reg[4]/P0001  ;
	input \u1_sram_addr_reg[5]/P0001  ;
	input \u1_sram_addr_reg[6]/P0001  ;
	input \u1_sram_addr_reg[7]/P0001  ;
	input \u1_sram_addr_reg[8]/P0001  ;
	input \u1_sram_addr_reg[9]/P0001  ;
	input \u1_u0_out_r_reg[0]/P0001  ;
	input \u1_u0_out_r_reg[10]/P0001  ;
	input \u1_u0_out_r_reg[11]/P0001  ;
	input \u1_u0_out_r_reg[12]/P0001  ;
	input \u1_u0_out_r_reg[1]/P0001  ;
	input \u1_u0_out_r_reg[2]/P0001  ;
	input \u1_u0_out_r_reg[3]/P0001  ;
	input \u1_u0_out_r_reg[4]/P0001  ;
	input \u1_u0_out_r_reg[5]/P0001  ;
	input \u1_u0_out_r_reg[6]/P0001  ;
	input \u1_u0_out_r_reg[7]/P0001  ;
	input \u1_u0_out_r_reg[8]/P0001  ;
	input \u1_u0_out_r_reg[9]/P0001  ;
	input \u2_bank_open_reg/P0001  ;
	input \u2_row_same_reg/P0001  ;
	input \u2_u0_b0_last_row_reg[0]/P0001  ;
	input \u2_u0_b0_last_row_reg[10]/P0001  ;
	input \u2_u0_b0_last_row_reg[11]/P0001  ;
	input \u2_u0_b0_last_row_reg[12]/P0001  ;
	input \u2_u0_b0_last_row_reg[1]/P0001  ;
	input \u2_u0_b0_last_row_reg[2]/P0001  ;
	input \u2_u0_b0_last_row_reg[3]/P0001  ;
	input \u2_u0_b0_last_row_reg[4]/P0001  ;
	input \u2_u0_b0_last_row_reg[5]/P0001  ;
	input \u2_u0_b0_last_row_reg[6]/P0001  ;
	input \u2_u0_b0_last_row_reg[7]/P0001  ;
	input \u2_u0_b0_last_row_reg[8]/P0001  ;
	input \u2_u0_b0_last_row_reg[9]/P0001  ;
	input \u2_u0_b1_last_row_reg[0]/P0001  ;
	input \u2_u0_b1_last_row_reg[10]/P0001  ;
	input \u2_u0_b1_last_row_reg[11]/P0001  ;
	input \u2_u0_b1_last_row_reg[12]/P0001  ;
	input \u2_u0_b1_last_row_reg[1]/P0001  ;
	input \u2_u0_b1_last_row_reg[2]/P0001  ;
	input \u2_u0_b1_last_row_reg[3]/P0001  ;
	input \u2_u0_b1_last_row_reg[4]/P0001  ;
	input \u2_u0_b1_last_row_reg[5]/P0001  ;
	input \u2_u0_b1_last_row_reg[6]/P0001  ;
	input \u2_u0_b1_last_row_reg[7]/P0001  ;
	input \u2_u0_b1_last_row_reg[8]/P0001  ;
	input \u2_u0_b1_last_row_reg[9]/P0001  ;
	input \u2_u0_b2_last_row_reg[0]/P0001  ;
	input \u2_u0_b2_last_row_reg[10]/P0001  ;
	input \u2_u0_b2_last_row_reg[11]/P0001  ;
	input \u2_u0_b2_last_row_reg[12]/P0001  ;
	input \u2_u0_b2_last_row_reg[1]/P0001  ;
	input \u2_u0_b2_last_row_reg[2]/P0001  ;
	input \u2_u0_b2_last_row_reg[3]/P0001  ;
	input \u2_u0_b2_last_row_reg[4]/P0001  ;
	input \u2_u0_b2_last_row_reg[5]/P0001  ;
	input \u2_u0_b2_last_row_reg[6]/P0001  ;
	input \u2_u0_b2_last_row_reg[7]/P0001  ;
	input \u2_u0_b2_last_row_reg[8]/P0001  ;
	input \u2_u0_b2_last_row_reg[9]/P0001  ;
	input \u2_u0_b3_last_row_reg[0]/P0001  ;
	input \u2_u0_b3_last_row_reg[10]/P0001  ;
	input \u2_u0_b3_last_row_reg[11]/P0001  ;
	input \u2_u0_b3_last_row_reg[12]/P0001  ;
	input \u2_u0_b3_last_row_reg[1]/P0001  ;
	input \u2_u0_b3_last_row_reg[2]/P0001  ;
	input \u2_u0_b3_last_row_reg[3]/P0001  ;
	input \u2_u0_b3_last_row_reg[4]/P0001  ;
	input \u2_u0_b3_last_row_reg[5]/P0001  ;
	input \u2_u0_b3_last_row_reg[6]/P0001  ;
	input \u2_u0_b3_last_row_reg[7]/P0001  ;
	input \u2_u0_b3_last_row_reg[8]/P0001  ;
	input \u2_u0_b3_last_row_reg[9]/P0001  ;
	input \u2_u0_bank0_open_reg/NET0131  ;
	input \u2_u0_bank1_open_reg/NET0131  ;
	input \u2_u0_bank2_open_reg/NET0131  ;
	input \u2_u0_bank3_open_reg/NET0131  ;
	input \u2_u1_b0_last_row_reg[0]/P0001  ;
	input \u2_u1_b0_last_row_reg[10]/P0001  ;
	input \u2_u1_b0_last_row_reg[11]/P0001  ;
	input \u2_u1_b0_last_row_reg[12]/P0001  ;
	input \u2_u1_b0_last_row_reg[1]/P0001  ;
	input \u2_u1_b0_last_row_reg[2]/P0001  ;
	input \u2_u1_b0_last_row_reg[3]/P0001  ;
	input \u2_u1_b0_last_row_reg[4]/P0001  ;
	input \u2_u1_b0_last_row_reg[5]/P0001  ;
	input \u2_u1_b0_last_row_reg[6]/P0001  ;
	input \u2_u1_b0_last_row_reg[7]/P0001  ;
	input \u2_u1_b0_last_row_reg[8]/P0001  ;
	input \u2_u1_b0_last_row_reg[9]/P0001  ;
	input \u2_u1_b1_last_row_reg[0]/P0001  ;
	input \u2_u1_b1_last_row_reg[10]/P0001  ;
	input \u2_u1_b1_last_row_reg[11]/P0001  ;
	input \u2_u1_b1_last_row_reg[12]/P0001  ;
	input \u2_u1_b1_last_row_reg[1]/P0001  ;
	input \u2_u1_b1_last_row_reg[2]/P0001  ;
	input \u2_u1_b1_last_row_reg[3]/P0001  ;
	input \u2_u1_b1_last_row_reg[4]/P0001  ;
	input \u2_u1_b1_last_row_reg[5]/P0001  ;
	input \u2_u1_b1_last_row_reg[6]/P0001  ;
	input \u2_u1_b1_last_row_reg[7]/P0001  ;
	input \u2_u1_b1_last_row_reg[8]/P0001  ;
	input \u2_u1_b1_last_row_reg[9]/P0001  ;
	input \u2_u1_b2_last_row_reg[0]/P0001  ;
	input \u2_u1_b2_last_row_reg[10]/P0001  ;
	input \u2_u1_b2_last_row_reg[11]/P0001  ;
	input \u2_u1_b2_last_row_reg[12]/P0001  ;
	input \u2_u1_b2_last_row_reg[1]/P0001  ;
	input \u2_u1_b2_last_row_reg[2]/P0001  ;
	input \u2_u1_b2_last_row_reg[3]/P0001  ;
	input \u2_u1_b2_last_row_reg[4]/P0001  ;
	input \u2_u1_b2_last_row_reg[5]/P0001  ;
	input \u2_u1_b2_last_row_reg[6]/P0001  ;
	input \u2_u1_b2_last_row_reg[7]/P0001  ;
	input \u2_u1_b2_last_row_reg[8]/P0001  ;
	input \u2_u1_b2_last_row_reg[9]/P0001  ;
	input \u2_u1_b3_last_row_reg[0]/P0001  ;
	input \u2_u1_b3_last_row_reg[10]/P0001  ;
	input \u2_u1_b3_last_row_reg[11]/P0001  ;
	input \u2_u1_b3_last_row_reg[12]/P0001  ;
	input \u2_u1_b3_last_row_reg[1]/P0001  ;
	input \u2_u1_b3_last_row_reg[2]/P0001  ;
	input \u2_u1_b3_last_row_reg[3]/P0001  ;
	input \u2_u1_b3_last_row_reg[4]/P0001  ;
	input \u2_u1_b3_last_row_reg[5]/P0001  ;
	input \u2_u1_b3_last_row_reg[6]/P0001  ;
	input \u2_u1_b3_last_row_reg[7]/P0001  ;
	input \u2_u1_b3_last_row_reg[8]/P0001  ;
	input \u2_u1_b3_last_row_reg[9]/P0001  ;
	input \u2_u1_bank0_open_reg/NET0131  ;
	input \u2_u1_bank1_open_reg/NET0131  ;
	input \u2_u1_bank2_open_reg/NET0131  ;
	input \u2_u1_bank3_open_reg/NET0131  ;
	input \u3_byte0_reg[0]/P0001  ;
	input \u3_byte0_reg[1]/P0001  ;
	input \u3_byte0_reg[2]/P0001  ;
	input \u3_byte0_reg[3]/P0001  ;
	input \u3_byte0_reg[4]/P0001  ;
	input \u3_byte0_reg[5]/P0001  ;
	input \u3_byte0_reg[6]/P0001  ;
	input \u3_byte0_reg[7]/P0001  ;
	input \u3_byte1_reg[0]/P0001  ;
	input \u3_byte1_reg[1]/P0001  ;
	input \u3_byte1_reg[2]/P0001  ;
	input \u3_byte1_reg[3]/P0001  ;
	input \u3_byte1_reg[4]/P0001  ;
	input \u3_byte1_reg[5]/P0001  ;
	input \u3_byte1_reg[6]/P0001  ;
	input \u3_byte1_reg[7]/P0001  ;
	input \u3_byte2_reg[0]/P0001  ;
	input \u3_byte2_reg[1]/P0001  ;
	input \u3_byte2_reg[2]/P0001  ;
	input \u3_byte2_reg[3]/P0001  ;
	input \u3_byte2_reg[4]/P0001  ;
	input \u3_byte2_reg[5]/P0001  ;
	input \u3_byte2_reg[6]/P0001  ;
	input \u3_byte2_reg[7]/P0001  ;
	input \u3_u0_r0_reg[0]/P0001  ;
	input \u3_u0_r0_reg[10]/P0001  ;
	input \u3_u0_r0_reg[11]/P0001  ;
	input \u3_u0_r0_reg[12]/P0001  ;
	input \u3_u0_r0_reg[13]/P0001  ;
	input \u3_u0_r0_reg[14]/P0001  ;
	input \u3_u0_r0_reg[15]/P0001  ;
	input \u3_u0_r0_reg[16]/P0001  ;
	input \u3_u0_r0_reg[17]/P0001  ;
	input \u3_u0_r0_reg[18]/P0001  ;
	input \u3_u0_r0_reg[19]/P0001  ;
	input \u3_u0_r0_reg[1]/P0001  ;
	input \u3_u0_r0_reg[20]/P0001  ;
	input \u3_u0_r0_reg[21]/P0001  ;
	input \u3_u0_r0_reg[22]/P0001  ;
	input \u3_u0_r0_reg[23]/P0001  ;
	input \u3_u0_r0_reg[24]/P0001  ;
	input \u3_u0_r0_reg[25]/P0001  ;
	input \u3_u0_r0_reg[26]/P0001  ;
	input \u3_u0_r0_reg[27]/P0001  ;
	input \u3_u0_r0_reg[28]/P0001  ;
	input \u3_u0_r0_reg[29]/P0001  ;
	input \u3_u0_r0_reg[2]/P0001  ;
	input \u3_u0_r0_reg[30]/P0001  ;
	input \u3_u0_r0_reg[31]/P0001  ;
	input \u3_u0_r0_reg[32]/P0001  ;
	input \u3_u0_r0_reg[33]/P0001  ;
	input \u3_u0_r0_reg[34]/P0001  ;
	input \u3_u0_r0_reg[35]/P0001  ;
	input \u3_u0_r0_reg[3]/P0001  ;
	input \u3_u0_r0_reg[4]/P0001  ;
	input \u3_u0_r0_reg[5]/P0001  ;
	input \u3_u0_r0_reg[6]/P0001  ;
	input \u3_u0_r0_reg[7]/P0001  ;
	input \u3_u0_r0_reg[8]/P0001  ;
	input \u3_u0_r0_reg[9]/P0001  ;
	input \u3_u0_r1_reg[0]/P0001  ;
	input \u3_u0_r1_reg[10]/P0001  ;
	input \u3_u0_r1_reg[11]/P0001  ;
	input \u3_u0_r1_reg[12]/P0001  ;
	input \u3_u0_r1_reg[13]/P0001  ;
	input \u3_u0_r1_reg[14]/P0001  ;
	input \u3_u0_r1_reg[15]/P0001  ;
	input \u3_u0_r1_reg[16]/P0001  ;
	input \u3_u0_r1_reg[17]/P0001  ;
	input \u3_u0_r1_reg[18]/P0001  ;
	input \u3_u0_r1_reg[19]/P0001  ;
	input \u3_u0_r1_reg[1]/P0001  ;
	input \u3_u0_r1_reg[20]/P0001  ;
	input \u3_u0_r1_reg[21]/P0001  ;
	input \u3_u0_r1_reg[22]/P0001  ;
	input \u3_u0_r1_reg[23]/P0001  ;
	input \u3_u0_r1_reg[24]/P0001  ;
	input \u3_u0_r1_reg[25]/P0001  ;
	input \u3_u0_r1_reg[26]/P0001  ;
	input \u3_u0_r1_reg[27]/P0001  ;
	input \u3_u0_r1_reg[28]/P0001  ;
	input \u3_u0_r1_reg[29]/P0001  ;
	input \u3_u0_r1_reg[2]/P0001  ;
	input \u3_u0_r1_reg[30]/P0001  ;
	input \u3_u0_r1_reg[31]/P0001  ;
	input \u3_u0_r1_reg[32]/P0001  ;
	input \u3_u0_r1_reg[33]/P0001  ;
	input \u3_u0_r1_reg[34]/P0001  ;
	input \u3_u0_r1_reg[35]/P0001  ;
	input \u3_u0_r1_reg[3]/P0001  ;
	input \u3_u0_r1_reg[4]/P0001  ;
	input \u3_u0_r1_reg[5]/P0001  ;
	input \u3_u0_r1_reg[6]/P0001  ;
	input \u3_u0_r1_reg[7]/P0001  ;
	input \u3_u0_r1_reg[8]/P0001  ;
	input \u3_u0_r1_reg[9]/P0001  ;
	input \u3_u0_r2_reg[0]/P0001  ;
	input \u3_u0_r2_reg[10]/P0001  ;
	input \u3_u0_r2_reg[11]/P0001  ;
	input \u3_u0_r2_reg[12]/P0001  ;
	input \u3_u0_r2_reg[13]/P0001  ;
	input \u3_u0_r2_reg[14]/P0001  ;
	input \u3_u0_r2_reg[15]/P0001  ;
	input \u3_u0_r2_reg[16]/P0001  ;
	input \u3_u0_r2_reg[17]/P0001  ;
	input \u3_u0_r2_reg[18]/P0001  ;
	input \u3_u0_r2_reg[19]/P0001  ;
	input \u3_u0_r2_reg[1]/P0001  ;
	input \u3_u0_r2_reg[20]/P0001  ;
	input \u3_u0_r2_reg[21]/P0001  ;
	input \u3_u0_r2_reg[22]/P0001  ;
	input \u3_u0_r2_reg[23]/P0001  ;
	input \u3_u0_r2_reg[24]/P0001  ;
	input \u3_u0_r2_reg[25]/P0001  ;
	input \u3_u0_r2_reg[26]/P0001  ;
	input \u3_u0_r2_reg[27]/P0001  ;
	input \u3_u0_r2_reg[28]/P0001  ;
	input \u3_u0_r2_reg[29]/P0001  ;
	input \u3_u0_r2_reg[2]/P0001  ;
	input \u3_u0_r2_reg[30]/P0001  ;
	input \u3_u0_r2_reg[31]/P0001  ;
	input \u3_u0_r2_reg[32]/P0001  ;
	input \u3_u0_r2_reg[33]/P0001  ;
	input \u3_u0_r2_reg[34]/P0001  ;
	input \u3_u0_r2_reg[35]/P0001  ;
	input \u3_u0_r2_reg[3]/P0001  ;
	input \u3_u0_r2_reg[4]/P0001  ;
	input \u3_u0_r2_reg[5]/P0001  ;
	input \u3_u0_r2_reg[6]/P0001  ;
	input \u3_u0_r2_reg[7]/P0001  ;
	input \u3_u0_r2_reg[8]/P0001  ;
	input \u3_u0_r2_reg[9]/P0001  ;
	input \u3_u0_r3_reg[0]/P0001  ;
	input \u3_u0_r3_reg[10]/P0001  ;
	input \u3_u0_r3_reg[11]/P0001  ;
	input \u3_u0_r3_reg[12]/P0001  ;
	input \u3_u0_r3_reg[13]/P0001  ;
	input \u3_u0_r3_reg[14]/P0001  ;
	input \u3_u0_r3_reg[15]/P0001  ;
	input \u3_u0_r3_reg[16]/P0001  ;
	input \u3_u0_r3_reg[17]/P0001  ;
	input \u3_u0_r3_reg[18]/P0001  ;
	input \u3_u0_r3_reg[19]/P0001  ;
	input \u3_u0_r3_reg[1]/P0001  ;
	input \u3_u0_r3_reg[20]/P0001  ;
	input \u3_u0_r3_reg[21]/P0001  ;
	input \u3_u0_r3_reg[22]/P0001  ;
	input \u3_u0_r3_reg[23]/P0001  ;
	input \u3_u0_r3_reg[24]/P0001  ;
	input \u3_u0_r3_reg[25]/P0001  ;
	input \u3_u0_r3_reg[26]/P0001  ;
	input \u3_u0_r3_reg[27]/P0001  ;
	input \u3_u0_r3_reg[28]/P0001  ;
	input \u3_u0_r3_reg[29]/P0001  ;
	input \u3_u0_r3_reg[2]/P0001  ;
	input \u3_u0_r3_reg[30]/P0001  ;
	input \u3_u0_r3_reg[31]/P0001  ;
	input \u3_u0_r3_reg[32]/P0001  ;
	input \u3_u0_r3_reg[33]/P0001  ;
	input \u3_u0_r3_reg[34]/P0001  ;
	input \u3_u0_r3_reg[35]/P0001  ;
	input \u3_u0_r3_reg[3]/P0001  ;
	input \u3_u0_r3_reg[4]/P0001  ;
	input \u3_u0_r3_reg[5]/P0001  ;
	input \u3_u0_r3_reg[6]/P0001  ;
	input \u3_u0_r3_reg[7]/P0001  ;
	input \u3_u0_r3_reg[8]/P0001  ;
	input \u3_u0_r3_reg[9]/P0001  ;
	input \u3_u0_rd_adr_reg[0]/NET0131  ;
	input \u3_u0_rd_adr_reg[1]/NET0131  ;
	input \u3_u0_rd_adr_reg[2]/NET0131  ;
	input \u3_u0_rd_adr_reg[3]/NET0131  ;
	input \u3_u0_wr_adr_reg[0]/NET0131  ;
	input \u3_u0_wr_adr_reg[1]/NET0131  ;
	input \u3_u0_wr_adr_reg[2]/NET0131  ;
	input \u3_u0_wr_adr_reg[3]/NET0131  ;
	input \u4_ps_cnt_reg[0]/NET0131  ;
	input \u4_ps_cnt_reg[1]/NET0131  ;
	input \u4_ps_cnt_reg[2]/NET0131  ;
	input \u4_ps_cnt_reg[3]/NET0131  ;
	input \u4_ps_cnt_reg[4]/NET0131  ;
	input \u4_ps_cnt_reg[5]/NET0131  ;
	input \u4_ps_cnt_reg[6]/NET0131  ;
	input \u4_ps_cnt_reg[7]/NET0131  ;
	input \u4_rfr_ce_reg/NET0131  ;
	input \u4_rfr_clr_reg/P0001  ;
	input \u4_rfr_cnt_reg[0]/NET0131  ;
	input \u4_rfr_cnt_reg[1]/NET0131  ;
	input \u4_rfr_cnt_reg[2]/NET0131  ;
	input \u4_rfr_cnt_reg[3]/NET0131  ;
	input \u4_rfr_cnt_reg[4]/NET0131  ;
	input \u4_rfr_cnt_reg[5]/NET0131  ;
	input \u4_rfr_cnt_reg[6]/NET0131  ;
	input \u4_rfr_cnt_reg[7]/NET0131  ;
	input \u4_rfr_early_reg/NET0131  ;
	input \u4_rfr_en_reg/NET0131  ;
	input \u4_rfr_req_reg/NET0131  ;
	input \u5_ack_cnt_reg[0]/NET0131  ;
	input \u5_ack_cnt_reg[1]/NET0131  ;
	input \u5_ack_cnt_reg[2]/NET0131  ;
	input \u5_ack_cnt_reg[3]/NET0131  ;
	input \u5_ap_en_reg/NET0131  ;
	input \u5_burst_act_rd_reg/P0001  ;
	input \u5_burst_cnt_reg[0]/NET0131  ;
	input \u5_burst_cnt_reg[10]/NET0131  ;
	input \u5_burst_cnt_reg[1]/NET0131  ;
	input \u5_burst_cnt_reg[2]/NET0131  ;
	input \u5_burst_cnt_reg[3]/NET0131  ;
	input \u5_burst_cnt_reg[4]/NET0131  ;
	input \u5_burst_cnt_reg[5]/NET0131  ;
	input \u5_burst_cnt_reg[6]/NET0131  ;
	input \u5_burst_cnt_reg[7]/NET0131  ;
	input \u5_burst_cnt_reg[8]/NET0131  ;
	input \u5_burst_cnt_reg[9]/NET0131  ;
	input \u5_cke_o_del_reg/P0001  ;
	input \u5_cke_r_reg/NET0131  ;
	input \u5_cmd_a10_r_reg/P0001  ;
	input \u5_cmd_asserted2_reg/NET0131  ;
	input \u5_cmd_asserted_reg/NET0131  ;
	input \u5_cmd_del_reg[0]/NET0131  ;
	input \u5_cmd_del_reg[1]/NET0131  ;
	input \u5_cmd_del_reg[2]/NET0131  ;
	input \u5_cmd_del_reg[3]/NET0131  ;
	input \u5_cnt_reg/NET0131  ;
	input \u5_cs_le_r_reg/P0001  ;
	input \u5_cs_le_reg/P0001  ;
	input \u5_data_oe_r2_reg/NET0131  ;
	input \u5_data_oe_reg/NET0131  ;
	input \u5_dv_r_reg/NET0131  ;
	input \u5_ir_cnt_done_reg/P0001  ;
	input \u5_ir_cnt_reg[0]/P0001  ;
	input \u5_ir_cnt_reg[1]/P0001  ;
	input \u5_ir_cnt_reg[2]/P0001  ;
	input \u5_ir_cnt_reg[3]/P0001  ;
	input \u5_lmr_ack_reg/NET0131  ;
	input \u5_lookup_ready1_reg/NET0131  ;
	input \u5_lookup_ready2_reg/NET0131  ;
	input \u5_mc_adv_r1_reg/NET0131  ;
	input \u5_mc_adv_r_reg/NET0131  ;
	input \u5_mc_c_oe_reg/NET0131  ;
	input \u5_mc_le_reg/NET0131  ;
	input \u5_mem_ack_r_reg/NET0131  ;
	input \u5_no_wb_cycle_reg/NET0131  ;
	input \u5_oe__reg/NET0131  ;
	input \u5_pack_le0_reg/P0001  ;
	input \u5_pack_le1_reg/P0001  ;
	input \u5_resume_req_r_reg/NET0131  ;
	input \u5_rfr_ack_r_reg/NET0131  ;
	input \u5_state_reg[0]/NET0131  ;
	input \u5_state_reg[10]/NET0131  ;
	input \u5_state_reg[11]/NET0131  ;
	input \u5_state_reg[12]/NET0131  ;
	input \u5_state_reg[13]/NET0131  ;
	input \u5_state_reg[14]/NET0131  ;
	input \u5_state_reg[15]/NET0131  ;
	input \u5_state_reg[16]/NET0131  ;
	input \u5_state_reg[17]/NET0131  ;
	input \u5_state_reg[18]/NET0131  ;
	input \u5_state_reg[19]/NET0131  ;
	input \u5_state_reg[1]/NET0131  ;
	input \u5_state_reg[20]/NET0131  ;
	input \u5_state_reg[21]/NET0131  ;
	input \u5_state_reg[22]/NET0131  ;
	input \u5_state_reg[23]/NET0131  ;
	input \u5_state_reg[24]/NET0131  ;
	input \u5_state_reg[25]/NET0131  ;
	input \u5_state_reg[26]/NET0131  ;
	input \u5_state_reg[27]/NET0131  ;
	input \u5_state_reg[28]/NET0131  ;
	input \u5_state_reg[29]/NET0131  ;
	input \u5_state_reg[2]/NET0131  ;
	input \u5_state_reg[30]/NET0131  ;
	input \u5_state_reg[31]/NET0131  ;
	input \u5_state_reg[32]/NET0131  ;
	input \u5_state_reg[33]/NET0131  ;
	input \u5_state_reg[34]/NET0131  ;
	input \u5_state_reg[35]/NET0131  ;
	input \u5_state_reg[36]/NET0131  ;
	input \u5_state_reg[37]/NET0131  ;
	input \u5_state_reg[38]/NET0131  ;
	input \u5_state_reg[39]/NET0131  ;
	input \u5_state_reg[3]/NET0131  ;
	input \u5_state_reg[40]/NET0131  ;
	input \u5_state_reg[41]/NET0131  ;
	input \u5_state_reg[42]/NET0131  ;
	input \u5_state_reg[43]/NET0131  ;
	input \u5_state_reg[44]/NET0131  ;
	input \u5_state_reg[45]/NET0131  ;
	input \u5_state_reg[46]/NET0131  ;
	input \u5_state_reg[47]/NET0131  ;
	input \u5_state_reg[48]/NET0131  ;
	input \u5_state_reg[49]/NET0131  ;
	input \u5_state_reg[4]/NET0131  ;
	input \u5_state_reg[50]/NET0131  ;
	input \u5_state_reg[51]/NET0131  ;
	input \u5_state_reg[52]/NET0131  ;
	input \u5_state_reg[53]/NET0131  ;
	input \u5_state_reg[54]/NET0131  ;
	input \u5_state_reg[55]/NET0131  ;
	input \u5_state_reg[56]/NET0131  ;
	input \u5_state_reg[57]/NET0131  ;
	input \u5_state_reg[58]/NET0131  ;
	input \u5_state_reg[59]/NET0131  ;
	input \u5_state_reg[5]/NET0131  ;
	input \u5_state_reg[60]/NET0131  ;
	input \u5_state_reg[61]/NET0131  ;
	input \u5_state_reg[62]/NET0131  ;
	input \u5_state_reg[63]/NET0131  ;
	input \u5_state_reg[64]/NET0131  ;
	input \u5_state_reg[65]/NET0131  ;
	input \u5_state_reg[6]/NET0131  ;
	input \u5_state_reg[7]/NET0131  ;
	input \u5_state_reg[8]/NET0131  ;
	input \u5_state_reg[9]/NET0131  ;
	input \u5_susp_req_r_reg/NET0131  ;
	input \u5_susp_sel_r_reg/NET0131  ;
	input \u5_timer2_reg[0]/P0001  ;
	input \u5_timer2_reg[1]/P0001  ;
	input \u5_timer2_reg[2]/P0001  ;
	input \u5_timer2_reg[3]/P0001  ;
	input \u5_timer2_reg[4]/P0001  ;
	input \u5_timer2_reg[5]/P0001  ;
	input \u5_timer2_reg[6]/P0001  ;
	input \u5_timer2_reg[7]/P0001  ;
	input \u5_timer2_reg[8]/P0001  ;
	input \u5_timer_reg[0]/NET0131  ;
	input \u5_timer_reg[1]/NET0131  ;
	input \u5_timer_reg[2]/NET0131  ;
	input \u5_timer_reg[3]/NET0131  ;
	input \u5_timer_reg[4]/NET0131  ;
	input \u5_timer_reg[5]/NET0131  ;
	input \u5_timer_reg[6]/NET0131  ;
	input \u5_timer_reg[7]/NET0131  ;
	input \u5_tmr2_done_reg/NET0131  ;
	input \u5_tmr_done_reg/NET0131  ;
	input \u5_wb_cycle_reg/NET0131  ;
	input \u5_wb_stb_first_reg/NET0131  ;
	input \u5_wb_wait_r_reg/P0001  ;
	input \u5_wb_write_go_r_reg/NET0131  ;
	input \u5_wr_cycle_reg/NET0131  ;
	input \u6_read_go_r1_reg/NET0131  ;
	input \u6_read_go_r_reg/NET0131  ;
	input \u6_rmw_en_reg/NET0131  ;
	input \u6_rmw_r_reg/NET0131  ;
	input \u6_wb_first_r_reg/NET0131  ;
	input \u6_wr_hold_reg/NET0131  ;
	input \u6_write_go_r1_reg/NET0131  ;
	input \u6_write_go_r_reg/NET0131  ;
	input \u7_mc_ack_r_reg/NET0131  ;
	input \u7_mc_br_r_reg/P0001  ;
	input \u7_mc_data_ir_reg[0]/P0001  ;
	input \u7_mc_data_ir_reg[10]/P0001  ;
	input \u7_mc_data_ir_reg[11]/P0001  ;
	input \u7_mc_data_ir_reg[12]/P0001  ;
	input \u7_mc_data_ir_reg[13]/P0001  ;
	input \u7_mc_data_ir_reg[14]/P0001  ;
	input \u7_mc_data_ir_reg[15]/P0001  ;
	input \u7_mc_data_ir_reg[16]/P0001  ;
	input \u7_mc_data_ir_reg[17]/P0001  ;
	input \u7_mc_data_ir_reg[18]/P0001  ;
	input \u7_mc_data_ir_reg[19]/P0001  ;
	input \u7_mc_data_ir_reg[1]/P0001  ;
	input \u7_mc_data_ir_reg[20]/P0001  ;
	input \u7_mc_data_ir_reg[21]/P0001  ;
	input \u7_mc_data_ir_reg[22]/P0001  ;
	input \u7_mc_data_ir_reg[23]/P0001  ;
	input \u7_mc_data_ir_reg[24]/P0001  ;
	input \u7_mc_data_ir_reg[25]/P0001  ;
	input \u7_mc_data_ir_reg[26]/P0001  ;
	input \u7_mc_data_ir_reg[27]/P0001  ;
	input \u7_mc_data_ir_reg[28]/P0001  ;
	input \u7_mc_data_ir_reg[29]/P0001  ;
	input \u7_mc_data_ir_reg[2]/P0001  ;
	input \u7_mc_data_ir_reg[30]/P0001  ;
	input \u7_mc_data_ir_reg[31]/P0001  ;
	input \u7_mc_data_ir_reg[3]/P0001  ;
	input \u7_mc_data_ir_reg[4]/P0001  ;
	input \u7_mc_data_ir_reg[5]/P0001  ;
	input \u7_mc_data_ir_reg[6]/P0001  ;
	input \u7_mc_data_ir_reg[7]/P0001  ;
	input \u7_mc_data_ir_reg[8]/P0001  ;
	input \u7_mc_data_ir_reg[9]/P0001  ;
	input \u7_mc_dqm_r2_reg[0]/P0001  ;
	input \u7_mc_dqm_r2_reg[1]/P0001  ;
	input \u7_mc_dqm_r2_reg[2]/P0001  ;
	input \u7_mc_dqm_r2_reg[3]/P0001  ;
	input \u7_mc_dqm_r_reg[0]/P0001  ;
	input \u7_mc_dqm_r_reg[1]/P0001  ;
	input \u7_mc_dqm_r_reg[2]/P0001  ;
	input \u7_mc_dqm_r_reg[3]/P0001  ;
	input wb_ack_o_pad ;
	input \wb_addr_i[0]_pad  ;
	input \wb_addr_i[10]_pad  ;
	input \wb_addr_i[11]_pad  ;
	input \wb_addr_i[12]_pad  ;
	input \wb_addr_i[13]_pad  ;
	input \wb_addr_i[14]_pad  ;
	input \wb_addr_i[15]_pad  ;
	input \wb_addr_i[16]_pad  ;
	input \wb_addr_i[17]_pad  ;
	input \wb_addr_i[18]_pad  ;
	input \wb_addr_i[19]_pad  ;
	input \wb_addr_i[1]_pad  ;
	input \wb_addr_i[20]_pad  ;
	input \wb_addr_i[21]_pad  ;
	input \wb_addr_i[22]_pad  ;
	input \wb_addr_i[23]_pad  ;
	input \wb_addr_i[24]_pad  ;
	input \wb_addr_i[25]_pad  ;
	input \wb_addr_i[26]_pad  ;
	input \wb_addr_i[27]_pad  ;
	input \wb_addr_i[28]_pad  ;
	input \wb_addr_i[29]_pad  ;
	input \wb_addr_i[2]_pad  ;
	input \wb_addr_i[30]_pad  ;
	input \wb_addr_i[31]_pad  ;
	input \wb_addr_i[3]_pad  ;
	input \wb_addr_i[4]_pad  ;
	input \wb_addr_i[5]_pad  ;
	input \wb_addr_i[6]_pad  ;
	input \wb_addr_i[7]_pad  ;
	input \wb_addr_i[8]_pad  ;
	input \wb_addr_i[9]_pad  ;
	input wb_cyc_i_pad ;
	input \wb_data_i[0]_pad  ;
	input \wb_data_i[10]_pad  ;
	input \wb_data_i[11]_pad  ;
	input \wb_data_i[12]_pad  ;
	input \wb_data_i[13]_pad  ;
	input \wb_data_i[14]_pad  ;
	input \wb_data_i[15]_pad  ;
	input \wb_data_i[16]_pad  ;
	input \wb_data_i[17]_pad  ;
	input \wb_data_i[18]_pad  ;
	input \wb_data_i[19]_pad  ;
	input \wb_data_i[1]_pad  ;
	input \wb_data_i[20]_pad  ;
	input \wb_data_i[21]_pad  ;
	input \wb_data_i[22]_pad  ;
	input \wb_data_i[23]_pad  ;
	input \wb_data_i[24]_pad  ;
	input \wb_data_i[25]_pad  ;
	input \wb_data_i[26]_pad  ;
	input \wb_data_i[27]_pad  ;
	input \wb_data_i[28]_pad  ;
	input \wb_data_i[29]_pad  ;
	input \wb_data_i[2]_pad  ;
	input \wb_data_i[30]_pad  ;
	input \wb_data_i[31]_pad  ;
	input \wb_data_i[3]_pad  ;
	input \wb_data_i[4]_pad  ;
	input \wb_data_i[5]_pad  ;
	input \wb_data_i[6]_pad  ;
	input \wb_data_i[7]_pad  ;
	input \wb_data_i[8]_pad  ;
	input \wb_data_i[9]_pad  ;
	input wb_err_o_pad ;
	input \wb_sel_i[0]_pad  ;
	input \wb_sel_i[1]_pad  ;
	input \wb_sel_i[2]_pad  ;
	input \wb_sel_i[3]_pad  ;
	input wb_stb_i_pad ;
	input wb_we_i_pad ;
	output \_al_n0  ;
	output \_al_n1  ;
	output \g22/_0_  ;
	output \g23/_0_  ;
	output \g25_dup61718/_2_  ;
	output \g43466/_0_  ;
	output \g43467/_0_  ;
	output \g43468/_0_  ;
	output \g43469/_0_  ;
	output \g43470/_0_  ;
	output \g43471/_0_  ;
	output \g43472/_0_  ;
	output \g43473/_0_  ;
	output \g43474/_0_  ;
	output \g43475/_0_  ;
	output \g43476/_0_  ;
	output \g43477/_0_  ;
	output \g43478/_0_  ;
	output \g43512/_0_  ;
	output \g43513/_0_  ;
	output \g43544/_3_  ;
	output \g43545/_0_  ;
	output \g43554/_0_  ;
	output \g43555/_0_  ;
	output \g43557/_0_  ;
	output \g43558/_0_  ;
	output \g43571/_2_  ;
	output \g43632/_0_  ;
	output \g43633/_0_  ;
	output \g43635/_0_  ;
	output \g43636/_0_  ;
	output \g43637/_0_  ;
	output \g43638/_0_  ;
	output \g43639/_0_  ;
	output \g43640/_0_  ;
	output \g43642/_0_  ;
	output \g43662/_0_  ;
	output \g43663/_0_  ;
	output \g43664/_0_  ;
	output \g43665/_0_  ;
	output \g43668/_0_  ;
	output \g43670/_0_  ;
	output \g43671/_0_  ;
	output \g43673/_0_  ;
	output \g43674/_0_  ;
	output \g43692/_0_  ;
	output \g43695/_0_  ;
	output \g43696/_0_  ;
	output \g43697/_0_  ;
	output \g43698/_0_  ;
	output \g43700/_0_  ;
	output \g43701/_0_  ;
	output \g43703/_0_  ;
	output \g43705/_0_  ;
	output \g43707/_0_  ;
	output \g43708/_0_  ;
	output \g43710/_0_  ;
	output \g43717/_0_  ;
	output \g43719/_0_  ;
	output \g43720/_0_  ;
	output \g43721/_0_  ;
	output \g43722/_1_  ;
	output \g43723/_0_  ;
	output \g43725/_0_  ;
	output \g43729/_0_  ;
	output \g43731/_0_  ;
	output \g43734/_0_  ;
	output \g43735/_0_  ;
	output \g43737/_0_  ;
	output \g43744/_0_  ;
	output \g43747/_0_  ;
	output \g43760/_2_  ;
	output \g43770/_1_  ;
	output \g43775/_2_  ;
	output \g43780/_2_  ;
	output \g43786/_0_  ;
	output \g43787/_1_  ;
	output \g43847/_0_  ;
	output \g43848/_1_  ;
	output \g43858/_1_  ;
	output \g43891/_3_  ;
	output \g43895/_0_  ;
	output \g43934/_0_  ;
	output \g43936/_3_  ;
	output \g43954/_3_  ;
	output \g43961/_0_  ;
	output \g44016/_1_  ;
	output \g44067/_0_  ;
	output \g44094/_0_  ;
	output \g44096/_0_  ;
	output \g44104/_0_  ;
	output \g44122/_0_  ;
	output \g44172/_0_  ;
	output \g44209/_0_  ;
	output \g44219/_0_  ;
	output \g44220/_0_  ;
	output \g44222/_0_  ;
	output \g44223/_0_  ;
	output \g44241/_2_  ;
	output \g44252/_0_  ;
	output \g44253/_0_  ;
	output \g44255/_2_  ;
	output \g44263/_2_  ;
	output \g44470/_0_  ;
	output \g44538/_0_  ;
	output \g44539/_0_  ;
	output \g44540/_0_  ;
	output \g44541/_0_  ;
	output \g44542/_0_  ;
	output \g44543/_0_  ;
	output \g44544/_0_  ;
	output \g44545/_0_  ;
	output \g44546/_0_  ;
	output \g44547/_0_  ;
	output \g44548/_0_  ;
	output \g44549/_0_  ;
	output \g44550/_0_  ;
	output \g44551/_0_  ;
	output \g44552/_0_  ;
	output \g44553/_0_  ;
	output \g44554/_0_  ;
	output \g44555/_0_  ;
	output \g44556/_0_  ;
	output \g44557/_0_  ;
	output \g44558/_0_  ;
	output \g44559/_0_  ;
	output \g44560/_0_  ;
	output \g44561/_0_  ;
	output \g44562/_0_  ;
	output \g44563/_0_  ;
	output \g44564/_0_  ;
	output \g44565/_0_  ;
	output \g44566/_0_  ;
	output \g44567/_0_  ;
	output \g44568/_0_  ;
	output \g44569/_0_  ;
	output \g44570/_0_  ;
	output \g44571/_0_  ;
	output \g44572/_0_  ;
	output \g44573/_0_  ;
	output \g44574/_0_  ;
	output \g44575/_0_  ;
	output \g44576/_0_  ;
	output \g44577/_0_  ;
	output \g44578/_0_  ;
	output \g44579/_0_  ;
	output \g44580/_0_  ;
	output \g44581/_0_  ;
	output \g44582/_0_  ;
	output \g44583/_0_  ;
	output \g44584/_0_  ;
	output \g44585/_0_  ;
	output \g44586/_0_  ;
	output \g44588/_0_  ;
	output \g44589/_0_  ;
	output \g44590/_0_  ;
	output \g44591/_0_  ;
	output \g44592/_0_  ;
	output \g44593/_0_  ;
	output \g44594/_0_  ;
	output \g44595/_0_  ;
	output \g44596/_0_  ;
	output \g44636/_2_  ;
	output \g44646/_0_  ;
	output \g44647/_0_  ;
	output \g44648/_0_  ;
	output \g44649/_0_  ;
	output \g44650/_0_  ;
	output \g44651/_0_  ;
	output \g44652/_0_  ;
	output \g44653/_0_  ;
	output \g44654/_0_  ;
	output \g44655/_0_  ;
	output \g44656/_0_  ;
	output \g44657/_0_  ;
	output \g44665/_0_  ;
	output \g44666/_0_  ;
	output \g44667/_0_  ;
	output \g44668/_0_  ;
	output \g44752/_0_  ;
	output \g44753/_0_  ;
	output \g44873/_0_  ;
	output \g44939/_0_  ;
	output \g44942/_0_  ;
	output \g44945/_0_  ;
	output \g45023/_2_  ;
	output \g45090/_0_  ;
	output \g45141/_0_  ;
	output \g45147/_3_  ;
	output \g45155/_0_  ;
	output \g45190/_0_  ;
	output \g45195/_2_  ;
	output \g45199/_2_  ;
	output \g45201/_2_  ;
	output \g45324/_0_  ;
	output \g45334/_2_  ;
	output \g45336/_0_  ;
	output \g45388/_0_  ;
	output \g45391/_0_  ;
	output \g45413/_2_  ;
	output \g45530/_0_  ;
	output \g45532/_0_  ;
	output \g45533/_0_  ;
	output \g45534/_0_  ;
	output \g45739/_2_  ;
	output \g45743/_2_  ;
	output \g45767/_0_  ;
	output \g45782/_0_  ;
	output \g45830/_3_  ;
	output \g45834/_3_  ;
	output \g45835/_3_  ;
	output \g45836/_3_  ;
	output \g45837/_3_  ;
	output \g45839/_3_  ;
	output \g45840/_3_  ;
	output \g45841/_3_  ;
	output \g45842/_3_  ;
	output \g45843/_3_  ;
	output \g45844/_3_  ;
	output \g45845/_3_  ;
	output \g46191/_0_  ;
	output \g46193/_3_  ;
	output \g46256/_3_  ;
	output \g46257/_3_  ;
	output \g46258/_3_  ;
	output \g46259/_3_  ;
	output \g46260/_3_  ;
	output \g46261/_3_  ;
	output \g46262/_3_  ;
	output \g46263/_3_  ;
	output \g46278/_0_  ;
	output \g46292/_0_  ;
	output \g46293/_0_  ;
	output \g46312/_0_  ;
	output \g46367/_2_  ;
	output \g46370/_2_  ;
	output \g46380/_2_  ;
	output \g46386/_2_  ;
	output \g46388/_2_  ;
	output \g46392/_2_  ;
	output \g46395/_2_  ;
	output \g46399/_2_  ;
	output \g46420/_0_  ;
	output \g46446/_0_  ;
	output \g46493/_0_  ;
	output \g46510/_0_  ;
	output \g46669/_2_  ;
	output \g46691/_0_  ;
	output \g46708/_0_  ;
	output \g46721/_00_  ;
	output \g46776/_0_  ;
	output \g46777/_0_  ;
	output \g46778/_0_  ;
	output \g46779/_0_  ;
	output \g46780/_0_  ;
	output \g46782/_0_  ;
	output \g46784/_0_  ;
	output \g46932/_0_  ;
	output \g47112/_0_  ;
	output \g47124/_0_  ;
	output \g47265/_0_  ;
	output \g47270/_0_  ;
	output \g47275/_0_  ;
	output \g47300/_1_  ;
	output \g47305/_1_  ;
	output \g47338/_0_  ;
	output \g47339/_0_  ;
	output \g47352/_0_  ;
	output \g47699/_3_  ;
	output \g47711/_0_  ;
	output \g47719/_3_  ;
	output \g47721/_3_  ;
	output \g47723/_3_  ;
	output \g47853/_0_  ;
	output \g48094/_0_  ;
	output \g48095/_0_  ;
	output \g48177/_2_  ;
	output \g48194/_0_  ;
	output \g48369/_2_  ;
	output \g48371/_2_  ;
	output \g48373/_2_  ;
	output \g48375/_2_  ;
	output \g48377/_2_  ;
	output \g48379/_2_  ;
	output \g48381/_2_  ;
	output \g48383/_2_  ;
	output \g48385/_2_  ;
	output \g48535/_0_  ;
	output \g48569/_0_  ;
	output \g48570/_0_  ;
	output \g48571/_0_  ;
	output \g48836/_0_  ;
	output \g48843/_0_  ;
	output \g49187/_3_  ;
	output \g49375/_2_  ;
	output \g49633/_0_  ;
	output \g49788/_1_  ;
	output \g49800/_1_  ;
	output \g49802/_1_  ;
	output \g49806/_1_  ;
	output \g49853/_1_  ;
	output \g49883/_0_  ;
	output \g49884/_0_  ;
	output \g49885/_0_  ;
	output \g49886/_0_  ;
	output \g49976/_1_  ;
	output \g50038/_0_  ;
	output \g50082/_0_  ;
	output \g50083/_0_  ;
	output \g50167/_3_  ;
	output \g50168/_3_  ;
	output \g50169/_3_  ;
	output \g50170/_3_  ;
	output \g50171/_3_  ;
	output \g50177/_0_  ;
	output \g50190/_0_  ;
	output \g50236/_0_  ;
	output \g50251/_3_  ;
	output \g50256/_0_  ;
	output \g50318/_3_  ;
	output \g50319/_3_  ;
	output \g50350/_3_  ;
	output \g50351/_3_  ;
	output \g50352/_3_  ;
	output \g50353/_3_  ;
	output \g50354/_3_  ;
	output \g50355/_3_  ;
	output \g50361/_2_  ;
	output \g50366/_0_  ;
	output \g50393/_0_  ;
	output \g50552/_1_  ;
	output \g51108/_0_  ;
	output \g51160/_0_  ;
	output \g51290/_1_  ;
	output \g51327/_3_  ;
	output \g51328/_3_  ;
	output \g51329/_3_  ;
	output \g51330/_3_  ;
	output \g51331/_3_  ;
	output \g51332/_3_  ;
	output \g51333/_3_  ;
	output \g51334/_3_  ;
	output \g51339/_3_  ;
	output \g51340/_3_  ;
	output \g51341/_3_  ;
	output \g51342/_3_  ;
	output \g51343/_3_  ;
	output \g51346/_0_  ;
	output \g51347/_0_  ;
	output \g51348/_0_  ;
	output \g51381/_3_  ;
	output \g51382/_3_  ;
	output \g51383/_3_  ;
	output \g51386/_3_  ;
	output \g51387/_3_  ;
	output \g51405/_3_  ;
	output \g51410/_3_  ;
	output \g51883/_0_  ;
	output \g51916/_0_  ;
	output \g51947/_0_  ;
	output \g51948/_0_  ;
	output \g51949/_0_  ;
	output \g51950/_0_  ;
	output \g51951/_0_  ;
	output \g51952/_0_  ;
	output \g51953/_0_  ;
	output \g51954/_0_  ;
	output \g51955/_0_  ;
	output \g51956/_0_  ;
	output \g51957/_0_  ;
	output \g51958/_0_  ;
	output \g51959/_0_  ;
	output \g51960/_0_  ;
	output \g51961/_0_  ;
	output \g51962/_0_  ;
	output \g51963/_0_  ;
	output \g51964/_0_  ;
	output \g51965/_0_  ;
	output \g51967/_0_  ;
	output \g51968/_0_  ;
	output \g51969/_0_  ;
	output \g51970/_0_  ;
	output \g51971/_0_  ;
	output \g51972/_0_  ;
	output \g51973/_0_  ;
	output \g51974/_0_  ;
	output \g51975/_0_  ;
	output \g51976/_0_  ;
	output \g51977/_0_  ;
	output \g51978/_0_  ;
	output \g51979/_0_  ;
	output \g51980/_0_  ;
	output \g51981/_0_  ;
	output \g51982/_0_  ;
	output \g51983/_0_  ;
	output \g51984/_0_  ;
	output \g51985/_0_  ;
	output \g51986/_0_  ;
	output \g51987/_0_  ;
	output \g51988/_0_  ;
	output \g51989/_0_  ;
	output \g51990/_0_  ;
	output \g51991/_0_  ;
	output \g51992/_0_  ;
	output \g51993/_0_  ;
	output \g51994/_0_  ;
	output \g51995/_0_  ;
	output \g51996/_0_  ;
	output \g51997/_0_  ;
	output \g51998/_0_  ;
	output \g51999/_0_  ;
	output \g52000/_0_  ;
	output \g52001/_0_  ;
	output \g52002/_0_  ;
	output \g52003/_0_  ;
	output \g52004/_0_  ;
	output \g52005/_0_  ;
	output \g52006/_0_  ;
	output \g52007/_0_  ;
	output \g52008/_0_  ;
	output \g52009/_0_  ;
	output \g52010/_0_  ;
	output \g52011/_0_  ;
	output \g52012/_0_  ;
	output \g52013/_0_  ;
	output \g52014/_0_  ;
	output \g52015/_0_  ;
	output \g52016/_0_  ;
	output \g52017/_0_  ;
	output \g52018/_0_  ;
	output \g52019/_0_  ;
	output \g52020/_0_  ;
	output \g52021/_0_  ;
	output \g52022/_0_  ;
	output \g52023/_0_  ;
	output \g52024/_0_  ;
	output \g52025/_0_  ;
	output \g52026/_0_  ;
	output \g52027/_0_  ;
	output \g52028/_0_  ;
	output \g52029/_0_  ;
	output \g52030/_0_  ;
	output \g52031/_0_  ;
	output \g52032/_0_  ;
	output \g52033/_0_  ;
	output \g52034/_0_  ;
	output \g52035/_0_  ;
	output \g52036/_0_  ;
	output \g52037/_0_  ;
	output \g52038/_0_  ;
	output \g52039/_0_  ;
	output \g52040/_0_  ;
	output \g52041/_0_  ;
	output \g52042/_0_  ;
	output \g52043/_0_  ;
	output \g52044/_0_  ;
	output \g52045/_0_  ;
	output \g52046/_0_  ;
	output \g52047/_0_  ;
	output \g52049/_0_  ;
	output \g52050/_0_  ;
	output \g52051/_0_  ;
	output \g52052/_0_  ;
	output \g52053/_0_  ;
	output \g52054/_0_  ;
	output \g52055/_0_  ;
	output \g52056/_0_  ;
	output \g52057/_0_  ;
	output \g52058/_0_  ;
	output \g52061/_0_  ;
	output \g52065/_0_  ;
	output \g52066/_0_  ;
	output \g52067/_0_  ;
	output \g52068/_0_  ;
	output \g52069/_0_  ;
	output \g52070/_0_  ;
	output \g52071/_0_  ;
	output \g52073/_0_  ;
	output \g52074/_0_  ;
	output \g52075/_0_  ;
	output \g52082/_0_  ;
	output \g52083/_0_  ;
	output \g52158/_0_  ;
	output \g52201/_0_  ;
	output \g52202/_0_  ;
	output \g52346/_0_  ;
	output \g52351/_0_  ;
	output \g52390/_0_  ;
	output \g52847/_0_  ;
	output \g52854/_0_  ;
	output \g52968/_0_  ;
	output \g52969/_0_  ;
	output \g52970/_0_  ;
	output \g52971/_0_  ;
	output \g52984/_0_  ;
	output \g52994/_0_  ;
	output \g53019/_0_  ;
	output \g53030/_0_  ;
	output \g53094/_1_  ;
	output \g53106/_0_  ;
	output \g53150/_0_  ;
	output \g53256/_0_  ;
	output \g53297/_0_  ;
	output \g53345/_0_  ;
	output \g53359/_0_  ;
	output \g53375/_0_  ;
	output \g53474/_1__syn_2  ;
	output \g53475/_2_  ;
	output \g53593/_0_  ;
	output \g53643/_1_  ;
	output \g53655/_0_  ;
	output \g53710/_0_  ;
	output \g53786/_0_  ;
	output \g53837/_0_  ;
	output \g53888/_1_  ;
	output \g53909/_0_  ;
	output \g54253/_2_  ;
	output \g54394/_3_  ;
	output \g54413/_0_  ;
	output \g55420/_0_  ;
	output \g55587/_0_  ;
	output \g55852/_0_  ;
	output \g57020/_0_  ;
	output \g59450/_0_  ;
	output \g59488/_2_  ;
	output \g59752/_0_  ;
	output \g59786/_0_  ;
	output \g59854/_0_  ;
	output \g59878/_0_  ;
	output \g59902/_0_  ;
	output \g59924/_0_  ;
	output \g59947/_0_  ;
	output \g59972/_0_  ;
	output \g59996/_0_  ;
	output \g60017/_0_  ;
	output \g60040/_0_  ;
	output \g60064/_0_  ;
	output \g60095/_0_  ;
	output \g60119/_0_  ;
	output \g60145/_1_  ;
	output \g60165/_0_  ;
	output \g60407/_2_  ;
	output \g60408/_0_  ;
	output \g60613/_2_  ;
	output \g60649/_0_  ;
	output \g60771/_0_  ;
	output \g60908/_1_  ;
	output \g60911/_0_  ;
	output \g60977/_0_  ;
	output \g61/_0_  ;
	output \g61002/_0_  ;
	output \g61308/_0_  ;
	output \g61312/_1_  ;
	output \g61314/_0_  ;
	output \g61319/_1_  ;
	output \g61342/_1_  ;
	output \g61360/_0_  ;
	output \g61377/_0_  ;
	output \g61423/_1_  ;
	output \g61426/_0_  ;
	output \g61479/_1_  ;
	output \g61523/_1_  ;
	output \g61558/_1_  ;
	output \g61652/_0_  ;
	output \g61866/_0_  ;
	output \g61868/_1_  ;
	output \g61887/_0_  ;
	output \u7_mc_dqm_r_reg[0]/P0001_reg_syn_3  ;
	output \u7_mc_dqm_r_reg[1]/P0001_reg_syn_3  ;
	output \u7_mc_dqm_r_reg[2]/P0001_reg_syn_3  ;
	output \u7_mc_dqm_r_reg[3]/P0001_reg_syn_3  ;
	output \u7_mc_we__reg/_05_  ;
	wire _w5408_ ;
	wire _w5407_ ;
	wire _w5406_ ;
	wire _w5405_ ;
	wire _w5404_ ;
	wire _w5403_ ;
	wire _w5402_ ;
	wire _w5401_ ;
	wire _w5400_ ;
	wire _w5399_ ;
	wire _w5398_ ;
	wire _w5397_ ;
	wire _w5396_ ;
	wire _w5395_ ;
	wire _w5394_ ;
	wire _w5393_ ;
	wire _w5392_ ;
	wire _w5391_ ;
	wire _w5390_ ;
	wire _w5389_ ;
	wire _w5388_ ;
	wire _w5387_ ;
	wire _w5386_ ;
	wire _w5384_ ;
	wire _w5383_ ;
	wire _w5382_ ;
	wire _w5381_ ;
	wire _w5380_ ;
	wire _w5379_ ;
	wire _w5378_ ;
	wire _w5377_ ;
	wire _w5376_ ;
	wire _w5375_ ;
	wire _w5374_ ;
	wire _w5373_ ;
	wire _w5372_ ;
	wire _w5371_ ;
	wire _w5370_ ;
	wire _w5369_ ;
	wire _w5368_ ;
	wire _w5367_ ;
	wire _w5366_ ;
	wire _w5365_ ;
	wire _w5364_ ;
	wire _w5363_ ;
	wire _w5362_ ;
	wire _w5361_ ;
	wire _w5360_ ;
	wire _w5359_ ;
	wire _w5358_ ;
	wire _w5357_ ;
	wire _w5356_ ;
	wire _w5355_ ;
	wire _w5354_ ;
	wire _w5353_ ;
	wire _w5352_ ;
	wire _w5351_ ;
	wire _w5350_ ;
	wire _w5349_ ;
	wire _w5348_ ;
	wire _w5347_ ;
	wire _w5346_ ;
	wire _w5345_ ;
	wire _w5344_ ;
	wire _w5343_ ;
	wire _w5342_ ;
	wire _w5341_ ;
	wire _w5340_ ;
	wire _w5339_ ;
	wire _w5338_ ;
	wire _w5337_ ;
	wire _w5336_ ;
	wire _w5335_ ;
	wire _w5334_ ;
	wire _w5333_ ;
	wire _w5332_ ;
	wire _w5331_ ;
	wire _w5330_ ;
	wire _w5329_ ;
	wire _w5328_ ;
	wire _w5327_ ;
	wire _w5326_ ;
	wire _w5325_ ;
	wire _w5324_ ;
	wire _w5323_ ;
	wire _w5322_ ;
	wire _w5321_ ;
	wire _w5320_ ;
	wire _w5319_ ;
	wire _w5318_ ;
	wire _w5317_ ;
	wire _w5316_ ;
	wire _w5315_ ;
	wire _w5314_ ;
	wire _w5313_ ;
	wire _w5312_ ;
	wire _w5311_ ;
	wire _w5310_ ;
	wire _w5309_ ;
	wire _w5308_ ;
	wire _w5307_ ;
	wire _w5306_ ;
	wire _w5305_ ;
	wire _w5304_ ;
	wire _w5303_ ;
	wire _w5302_ ;
	wire _w5301_ ;
	wire _w5300_ ;
	wire _w5299_ ;
	wire _w5298_ ;
	wire _w5297_ ;
	wire _w5296_ ;
	wire _w5295_ ;
	wire _w5294_ ;
	wire _w5293_ ;
	wire _w5292_ ;
	wire _w5291_ ;
	wire _w5290_ ;
	wire _w5289_ ;
	wire _w5288_ ;
	wire _w5287_ ;
	wire _w5286_ ;
	wire _w5285_ ;
	wire _w5284_ ;
	wire _w5283_ ;
	wire _w5282_ ;
	wire _w5281_ ;
	wire _w5280_ ;
	wire _w5279_ ;
	wire _w5278_ ;
	wire _w5277_ ;
	wire _w5276_ ;
	wire _w5275_ ;
	wire _w5274_ ;
	wire _w5273_ ;
	wire _w5272_ ;
	wire _w5271_ ;
	wire _w5270_ ;
	wire _w5269_ ;
	wire _w5268_ ;
	wire _w5267_ ;
	wire _w5266_ ;
	wire _w5265_ ;
	wire _w5264_ ;
	wire _w5263_ ;
	wire _w5262_ ;
	wire _w5261_ ;
	wire _w5260_ ;
	wire _w5259_ ;
	wire _w5258_ ;
	wire _w5257_ ;
	wire _w5256_ ;
	wire _w5255_ ;
	wire _w5254_ ;
	wire _w5253_ ;
	wire _w5252_ ;
	wire _w5251_ ;
	wire _w5250_ ;
	wire _w5249_ ;
	wire _w5248_ ;
	wire _w5247_ ;
	wire _w5246_ ;
	wire _w5245_ ;
	wire _w5244_ ;
	wire _w5243_ ;
	wire _w5242_ ;
	wire _w5241_ ;
	wire _w5240_ ;
	wire _w5239_ ;
	wire _w5238_ ;
	wire _w5237_ ;
	wire _w5236_ ;
	wire _w5235_ ;
	wire _w5234_ ;
	wire _w5233_ ;
	wire _w5232_ ;
	wire _w5231_ ;
	wire _w5230_ ;
	wire _w5229_ ;
	wire _w5228_ ;
	wire _w5227_ ;
	wire _w5226_ ;
	wire _w5225_ ;
	wire _w5224_ ;
	wire _w5223_ ;
	wire _w5222_ ;
	wire _w5221_ ;
	wire _w5220_ ;
	wire _w5219_ ;
	wire _w5218_ ;
	wire _w5217_ ;
	wire _w5216_ ;
	wire _w5215_ ;
	wire _w5214_ ;
	wire _w5213_ ;
	wire _w5212_ ;
	wire _w5211_ ;
	wire _w5210_ ;
	wire _w5209_ ;
	wire _w5208_ ;
	wire _w5207_ ;
	wire _w5206_ ;
	wire _w5205_ ;
	wire _w5204_ ;
	wire _w5203_ ;
	wire _w5202_ ;
	wire _w5201_ ;
	wire _w5200_ ;
	wire _w5199_ ;
	wire _w5198_ ;
	wire _w5197_ ;
	wire _w5196_ ;
	wire _w5195_ ;
	wire _w5194_ ;
	wire _w5193_ ;
	wire _w5192_ ;
	wire _w5191_ ;
	wire _w5190_ ;
	wire _w5189_ ;
	wire _w5188_ ;
	wire _w5187_ ;
	wire _w5186_ ;
	wire _w5185_ ;
	wire _w5184_ ;
	wire _w5183_ ;
	wire _w5182_ ;
	wire _w5181_ ;
	wire _w5180_ ;
	wire _w5179_ ;
	wire _w5178_ ;
	wire _w5177_ ;
	wire _w5176_ ;
	wire _w5175_ ;
	wire _w5174_ ;
	wire _w5173_ ;
	wire _w5172_ ;
	wire _w5171_ ;
	wire _w5170_ ;
	wire _w5169_ ;
	wire _w5168_ ;
	wire _w5167_ ;
	wire _w5166_ ;
	wire _w5165_ ;
	wire _w5164_ ;
	wire _w5163_ ;
	wire _w5162_ ;
	wire _w5161_ ;
	wire _w5160_ ;
	wire _w5159_ ;
	wire _w5158_ ;
	wire _w5157_ ;
	wire _w5156_ ;
	wire _w5155_ ;
	wire _w5154_ ;
	wire _w5153_ ;
	wire _w5152_ ;
	wire _w5151_ ;
	wire _w5150_ ;
	wire _w5149_ ;
	wire _w5148_ ;
	wire _w5147_ ;
	wire _w5146_ ;
	wire _w5145_ ;
	wire _w5144_ ;
	wire _w5143_ ;
	wire _w5142_ ;
	wire _w5141_ ;
	wire _w5140_ ;
	wire _w5139_ ;
	wire _w5138_ ;
	wire _w5137_ ;
	wire _w5136_ ;
	wire _w5135_ ;
	wire _w5134_ ;
	wire _w5133_ ;
	wire _w5132_ ;
	wire _w5131_ ;
	wire _w5130_ ;
	wire _w5129_ ;
	wire _w5128_ ;
	wire _w5127_ ;
	wire _w5126_ ;
	wire _w5125_ ;
	wire _w5124_ ;
	wire _w5123_ ;
	wire _w5122_ ;
	wire _w5121_ ;
	wire _w5120_ ;
	wire _w5119_ ;
	wire _w5118_ ;
	wire _w5117_ ;
	wire _w5116_ ;
	wire _w5115_ ;
	wire _w5114_ ;
	wire _w5113_ ;
	wire _w5112_ ;
	wire _w5111_ ;
	wire _w5110_ ;
	wire _w5109_ ;
	wire _w5108_ ;
	wire _w5107_ ;
	wire _w5106_ ;
	wire _w5105_ ;
	wire _w5104_ ;
	wire _w5103_ ;
	wire _w5102_ ;
	wire _w5101_ ;
	wire _w5100_ ;
	wire _w5099_ ;
	wire _w5098_ ;
	wire _w5097_ ;
	wire _w5096_ ;
	wire _w5095_ ;
	wire _w5094_ ;
	wire _w5093_ ;
	wire _w5092_ ;
	wire _w5091_ ;
	wire _w5090_ ;
	wire _w5089_ ;
	wire _w5088_ ;
	wire _w5087_ ;
	wire _w5086_ ;
	wire _w5085_ ;
	wire _w5084_ ;
	wire _w5083_ ;
	wire _w5082_ ;
	wire _w5081_ ;
	wire _w5080_ ;
	wire _w5079_ ;
	wire _w5078_ ;
	wire _w5077_ ;
	wire _w5076_ ;
	wire _w5075_ ;
	wire _w5074_ ;
	wire _w5073_ ;
	wire _w5072_ ;
	wire _w5071_ ;
	wire _w5070_ ;
	wire _w5069_ ;
	wire _w5068_ ;
	wire _w5067_ ;
	wire _w5066_ ;
	wire _w5065_ ;
	wire _w5064_ ;
	wire _w5063_ ;
	wire _w5062_ ;
	wire _w5061_ ;
	wire _w5060_ ;
	wire _w5059_ ;
	wire _w5058_ ;
	wire _w5057_ ;
	wire _w5056_ ;
	wire _w5055_ ;
	wire _w5054_ ;
	wire _w5053_ ;
	wire _w5052_ ;
	wire _w5051_ ;
	wire _w5050_ ;
	wire _w5049_ ;
	wire _w5048_ ;
	wire _w5047_ ;
	wire _w5046_ ;
	wire _w5045_ ;
	wire _w5044_ ;
	wire _w5043_ ;
	wire _w5042_ ;
	wire _w5041_ ;
	wire _w5040_ ;
	wire _w5039_ ;
	wire _w5038_ ;
	wire _w5037_ ;
	wire _w5036_ ;
	wire _w5035_ ;
	wire _w5034_ ;
	wire _w5033_ ;
	wire _w5032_ ;
	wire _w5031_ ;
	wire _w5030_ ;
	wire _w5029_ ;
	wire _w5028_ ;
	wire _w5027_ ;
	wire _w5026_ ;
	wire _w5025_ ;
	wire _w5024_ ;
	wire _w5023_ ;
	wire _w5022_ ;
	wire _w5021_ ;
	wire _w5020_ ;
	wire _w5019_ ;
	wire _w5018_ ;
	wire _w5017_ ;
	wire _w5016_ ;
	wire _w5015_ ;
	wire _w5014_ ;
	wire _w5013_ ;
	wire _w5012_ ;
	wire _w5011_ ;
	wire _w5010_ ;
	wire _w5009_ ;
	wire _w5008_ ;
	wire _w5007_ ;
	wire _w5006_ ;
	wire _w5005_ ;
	wire _w5004_ ;
	wire _w5003_ ;
	wire _w5002_ ;
	wire _w5001_ ;
	wire _w5000_ ;
	wire _w4999_ ;
	wire _w4998_ ;
	wire _w4997_ ;
	wire _w4996_ ;
	wire _w4995_ ;
	wire _w4994_ ;
	wire _w4993_ ;
	wire _w4992_ ;
	wire _w4991_ ;
	wire _w4990_ ;
	wire _w4989_ ;
	wire _w4988_ ;
	wire _w4987_ ;
	wire _w4986_ ;
	wire _w4985_ ;
	wire _w4984_ ;
	wire _w4983_ ;
	wire _w4982_ ;
	wire _w4981_ ;
	wire _w4980_ ;
	wire _w4979_ ;
	wire _w4978_ ;
	wire _w4977_ ;
	wire _w4976_ ;
	wire _w4975_ ;
	wire _w4974_ ;
	wire _w4973_ ;
	wire _w4972_ ;
	wire _w4971_ ;
	wire _w4970_ ;
	wire _w4969_ ;
	wire _w4968_ ;
	wire _w4967_ ;
	wire _w4966_ ;
	wire _w4965_ ;
	wire _w4964_ ;
	wire _w4963_ ;
	wire _w4962_ ;
	wire _w4961_ ;
	wire _w4960_ ;
	wire _w4959_ ;
	wire _w4958_ ;
	wire _w4957_ ;
	wire _w4956_ ;
	wire _w4955_ ;
	wire _w4954_ ;
	wire _w4953_ ;
	wire _w4952_ ;
	wire _w4951_ ;
	wire _w4950_ ;
	wire _w4949_ ;
	wire _w4948_ ;
	wire _w4947_ ;
	wire _w4946_ ;
	wire _w4945_ ;
	wire _w4944_ ;
	wire _w4943_ ;
	wire _w4942_ ;
	wire _w4941_ ;
	wire _w4940_ ;
	wire _w4939_ ;
	wire _w4938_ ;
	wire _w4937_ ;
	wire _w4936_ ;
	wire _w4935_ ;
	wire _w4934_ ;
	wire _w4933_ ;
	wire _w4932_ ;
	wire _w4931_ ;
	wire _w4930_ ;
	wire _w4929_ ;
	wire _w4928_ ;
	wire _w4927_ ;
	wire _w4926_ ;
	wire _w4925_ ;
	wire _w4924_ ;
	wire _w4923_ ;
	wire _w4922_ ;
	wire _w4921_ ;
	wire _w4920_ ;
	wire _w4919_ ;
	wire _w4918_ ;
	wire _w4917_ ;
	wire _w4916_ ;
	wire _w4915_ ;
	wire _w4914_ ;
	wire _w4913_ ;
	wire _w4912_ ;
	wire _w4911_ ;
	wire _w4910_ ;
	wire _w4909_ ;
	wire _w4908_ ;
	wire _w4907_ ;
	wire _w4906_ ;
	wire _w4905_ ;
	wire _w4904_ ;
	wire _w4903_ ;
	wire _w4902_ ;
	wire _w4901_ ;
	wire _w4900_ ;
	wire _w4899_ ;
	wire _w4898_ ;
	wire _w4897_ ;
	wire _w4896_ ;
	wire _w4895_ ;
	wire _w4894_ ;
	wire _w4893_ ;
	wire _w4892_ ;
	wire _w4891_ ;
	wire _w4890_ ;
	wire _w4889_ ;
	wire _w4888_ ;
	wire _w4887_ ;
	wire _w4886_ ;
	wire _w4885_ ;
	wire _w4884_ ;
	wire _w4883_ ;
	wire _w4882_ ;
	wire _w4881_ ;
	wire _w4880_ ;
	wire _w4879_ ;
	wire _w4878_ ;
	wire _w4877_ ;
	wire _w4876_ ;
	wire _w4875_ ;
	wire _w4874_ ;
	wire _w4873_ ;
	wire _w4872_ ;
	wire _w4871_ ;
	wire _w4870_ ;
	wire _w4869_ ;
	wire _w4868_ ;
	wire _w4867_ ;
	wire _w4866_ ;
	wire _w4865_ ;
	wire _w4864_ ;
	wire _w4863_ ;
	wire _w4862_ ;
	wire _w4861_ ;
	wire _w4860_ ;
	wire _w4859_ ;
	wire _w4858_ ;
	wire _w4857_ ;
	wire _w4856_ ;
	wire _w4855_ ;
	wire _w4854_ ;
	wire _w4853_ ;
	wire _w4852_ ;
	wire _w4851_ ;
	wire _w4850_ ;
	wire _w4849_ ;
	wire _w4848_ ;
	wire _w4847_ ;
	wire _w4846_ ;
	wire _w4845_ ;
	wire _w4844_ ;
	wire _w4843_ ;
	wire _w4842_ ;
	wire _w4841_ ;
	wire _w4840_ ;
	wire _w4839_ ;
	wire _w4838_ ;
	wire _w4837_ ;
	wire _w4836_ ;
	wire _w4835_ ;
	wire _w4834_ ;
	wire _w4833_ ;
	wire _w4832_ ;
	wire _w4831_ ;
	wire _w4830_ ;
	wire _w4829_ ;
	wire _w4828_ ;
	wire _w4827_ ;
	wire _w4826_ ;
	wire _w4825_ ;
	wire _w4824_ ;
	wire _w4823_ ;
	wire _w4822_ ;
	wire _w4821_ ;
	wire _w4820_ ;
	wire _w4819_ ;
	wire _w4818_ ;
	wire _w4817_ ;
	wire _w4816_ ;
	wire _w4815_ ;
	wire _w4814_ ;
	wire _w4813_ ;
	wire _w4812_ ;
	wire _w4811_ ;
	wire _w4810_ ;
	wire _w4809_ ;
	wire _w4808_ ;
	wire _w4807_ ;
	wire _w4806_ ;
	wire _w4805_ ;
	wire _w4804_ ;
	wire _w4803_ ;
	wire _w4802_ ;
	wire _w4801_ ;
	wire _w4800_ ;
	wire _w4799_ ;
	wire _w4798_ ;
	wire _w4797_ ;
	wire _w4796_ ;
	wire _w4795_ ;
	wire _w4794_ ;
	wire _w4793_ ;
	wire _w4792_ ;
	wire _w4791_ ;
	wire _w4790_ ;
	wire _w4789_ ;
	wire _w4788_ ;
	wire _w4787_ ;
	wire _w4786_ ;
	wire _w4785_ ;
	wire _w4784_ ;
	wire _w4783_ ;
	wire _w4782_ ;
	wire _w4781_ ;
	wire _w4780_ ;
	wire _w4779_ ;
	wire _w4778_ ;
	wire _w4777_ ;
	wire _w4776_ ;
	wire _w4775_ ;
	wire _w4774_ ;
	wire _w4773_ ;
	wire _w4772_ ;
	wire _w4771_ ;
	wire _w4770_ ;
	wire _w4769_ ;
	wire _w4768_ ;
	wire _w4767_ ;
	wire _w4766_ ;
	wire _w4765_ ;
	wire _w4764_ ;
	wire _w4763_ ;
	wire _w4762_ ;
	wire _w4761_ ;
	wire _w4760_ ;
	wire _w4759_ ;
	wire _w4758_ ;
	wire _w4757_ ;
	wire _w4756_ ;
	wire _w4755_ ;
	wire _w4754_ ;
	wire _w4753_ ;
	wire _w4752_ ;
	wire _w4751_ ;
	wire _w4750_ ;
	wire _w4749_ ;
	wire _w4748_ ;
	wire _w4747_ ;
	wire _w4746_ ;
	wire _w4745_ ;
	wire _w4744_ ;
	wire _w4743_ ;
	wire _w4742_ ;
	wire _w4741_ ;
	wire _w4740_ ;
	wire _w4739_ ;
	wire _w4738_ ;
	wire _w4737_ ;
	wire _w4736_ ;
	wire _w4735_ ;
	wire _w4734_ ;
	wire _w4733_ ;
	wire _w4732_ ;
	wire _w4731_ ;
	wire _w4730_ ;
	wire _w4729_ ;
	wire _w4728_ ;
	wire _w4727_ ;
	wire _w4726_ ;
	wire _w4725_ ;
	wire _w4724_ ;
	wire _w4723_ ;
	wire _w4722_ ;
	wire _w4721_ ;
	wire _w4720_ ;
	wire _w4719_ ;
	wire _w4718_ ;
	wire _w4717_ ;
	wire _w4716_ ;
	wire _w4715_ ;
	wire _w4714_ ;
	wire _w4713_ ;
	wire _w4712_ ;
	wire _w4711_ ;
	wire _w4710_ ;
	wire _w4709_ ;
	wire _w4708_ ;
	wire _w4707_ ;
	wire _w4706_ ;
	wire _w4705_ ;
	wire _w4704_ ;
	wire _w4703_ ;
	wire _w4702_ ;
	wire _w4701_ ;
	wire _w4700_ ;
	wire _w4699_ ;
	wire _w4698_ ;
	wire _w4697_ ;
	wire _w4696_ ;
	wire _w4695_ ;
	wire _w4694_ ;
	wire _w4693_ ;
	wire _w4692_ ;
	wire _w4691_ ;
	wire _w4690_ ;
	wire _w4689_ ;
	wire _w4688_ ;
	wire _w4687_ ;
	wire _w4686_ ;
	wire _w4685_ ;
	wire _w4684_ ;
	wire _w4683_ ;
	wire _w4682_ ;
	wire _w4681_ ;
	wire _w4680_ ;
	wire _w4679_ ;
	wire _w4678_ ;
	wire _w4677_ ;
	wire _w4676_ ;
	wire _w4675_ ;
	wire _w4674_ ;
	wire _w4673_ ;
	wire _w4672_ ;
	wire _w4671_ ;
	wire _w4670_ ;
	wire _w4669_ ;
	wire _w4668_ ;
	wire _w4667_ ;
	wire _w4666_ ;
	wire _w4665_ ;
	wire _w4664_ ;
	wire _w4663_ ;
	wire _w4662_ ;
	wire _w4661_ ;
	wire _w4660_ ;
	wire _w4659_ ;
	wire _w4658_ ;
	wire _w4657_ ;
	wire _w4656_ ;
	wire _w4655_ ;
	wire _w4654_ ;
	wire _w4653_ ;
	wire _w4652_ ;
	wire _w4651_ ;
	wire _w4650_ ;
	wire _w4649_ ;
	wire _w4648_ ;
	wire _w4647_ ;
	wire _w4646_ ;
	wire _w4645_ ;
	wire _w4644_ ;
	wire _w4643_ ;
	wire _w4642_ ;
	wire _w4641_ ;
	wire _w4640_ ;
	wire _w4639_ ;
	wire _w4638_ ;
	wire _w4637_ ;
	wire _w4636_ ;
	wire _w4635_ ;
	wire _w4634_ ;
	wire _w4633_ ;
	wire _w4632_ ;
	wire _w4631_ ;
	wire _w4630_ ;
	wire _w4629_ ;
	wire _w4628_ ;
	wire _w4627_ ;
	wire _w4626_ ;
	wire _w4625_ ;
	wire _w4624_ ;
	wire _w4623_ ;
	wire _w4622_ ;
	wire _w4621_ ;
	wire _w4620_ ;
	wire _w4619_ ;
	wire _w4618_ ;
	wire _w4617_ ;
	wire _w4616_ ;
	wire _w4615_ ;
	wire _w4614_ ;
	wire _w4613_ ;
	wire _w4612_ ;
	wire _w4611_ ;
	wire _w4610_ ;
	wire _w4609_ ;
	wire _w4608_ ;
	wire _w4607_ ;
	wire _w4606_ ;
	wire _w4605_ ;
	wire _w4604_ ;
	wire _w4603_ ;
	wire _w4602_ ;
	wire _w4601_ ;
	wire _w4600_ ;
	wire _w4599_ ;
	wire _w4598_ ;
	wire _w4597_ ;
	wire _w4596_ ;
	wire _w4595_ ;
	wire _w4594_ ;
	wire _w4593_ ;
	wire _w4592_ ;
	wire _w4591_ ;
	wire _w4590_ ;
	wire _w4589_ ;
	wire _w4588_ ;
	wire _w4587_ ;
	wire _w4586_ ;
	wire _w4585_ ;
	wire _w4584_ ;
	wire _w4583_ ;
	wire _w4582_ ;
	wire _w4581_ ;
	wire _w4580_ ;
	wire _w4579_ ;
	wire _w4578_ ;
	wire _w4577_ ;
	wire _w4576_ ;
	wire _w4575_ ;
	wire _w4574_ ;
	wire _w4573_ ;
	wire _w4572_ ;
	wire _w4571_ ;
	wire _w4570_ ;
	wire _w4569_ ;
	wire _w4568_ ;
	wire _w4567_ ;
	wire _w4566_ ;
	wire _w4565_ ;
	wire _w4564_ ;
	wire _w4563_ ;
	wire _w4562_ ;
	wire _w4561_ ;
	wire _w4560_ ;
	wire _w4559_ ;
	wire _w4558_ ;
	wire _w4557_ ;
	wire _w4556_ ;
	wire _w4555_ ;
	wire _w4554_ ;
	wire _w4553_ ;
	wire _w4552_ ;
	wire _w4551_ ;
	wire _w4550_ ;
	wire _w4549_ ;
	wire _w4548_ ;
	wire _w4547_ ;
	wire _w4546_ ;
	wire _w4545_ ;
	wire _w4544_ ;
	wire _w4543_ ;
	wire _w4542_ ;
	wire _w4541_ ;
	wire _w4540_ ;
	wire _w4539_ ;
	wire _w4538_ ;
	wire _w4537_ ;
	wire _w4536_ ;
	wire _w4535_ ;
	wire _w4534_ ;
	wire _w4533_ ;
	wire _w4532_ ;
	wire _w4531_ ;
	wire _w4530_ ;
	wire _w4529_ ;
	wire _w4528_ ;
	wire _w4527_ ;
	wire _w4526_ ;
	wire _w4525_ ;
	wire _w4524_ ;
	wire _w4523_ ;
	wire _w4522_ ;
	wire _w4521_ ;
	wire _w4520_ ;
	wire _w4519_ ;
	wire _w4518_ ;
	wire _w4517_ ;
	wire _w4516_ ;
	wire _w4515_ ;
	wire _w4514_ ;
	wire _w4513_ ;
	wire _w4512_ ;
	wire _w4511_ ;
	wire _w4510_ ;
	wire _w4509_ ;
	wire _w4508_ ;
	wire _w4507_ ;
	wire _w4506_ ;
	wire _w4505_ ;
	wire _w4504_ ;
	wire _w4503_ ;
	wire _w4502_ ;
	wire _w4501_ ;
	wire _w4500_ ;
	wire _w4499_ ;
	wire _w4498_ ;
	wire _w4497_ ;
	wire _w4496_ ;
	wire _w4495_ ;
	wire _w4494_ ;
	wire _w4493_ ;
	wire _w4492_ ;
	wire _w4491_ ;
	wire _w4490_ ;
	wire _w4489_ ;
	wire _w4488_ ;
	wire _w4487_ ;
	wire _w4486_ ;
	wire _w4485_ ;
	wire _w4484_ ;
	wire _w4483_ ;
	wire _w4482_ ;
	wire _w4481_ ;
	wire _w4480_ ;
	wire _w4479_ ;
	wire _w4478_ ;
	wire _w4477_ ;
	wire _w4476_ ;
	wire _w4475_ ;
	wire _w4474_ ;
	wire _w4473_ ;
	wire _w4472_ ;
	wire _w4471_ ;
	wire _w4470_ ;
	wire _w4469_ ;
	wire _w4468_ ;
	wire _w4467_ ;
	wire _w4466_ ;
	wire _w4465_ ;
	wire _w4464_ ;
	wire _w4463_ ;
	wire _w4462_ ;
	wire _w4461_ ;
	wire _w4460_ ;
	wire _w4459_ ;
	wire _w4458_ ;
	wire _w4457_ ;
	wire _w4456_ ;
	wire _w4455_ ;
	wire _w4454_ ;
	wire _w4453_ ;
	wire _w4452_ ;
	wire _w4451_ ;
	wire _w4450_ ;
	wire _w4449_ ;
	wire _w4448_ ;
	wire _w4447_ ;
	wire _w4446_ ;
	wire _w4445_ ;
	wire _w4444_ ;
	wire _w4443_ ;
	wire _w4442_ ;
	wire _w4441_ ;
	wire _w4440_ ;
	wire _w4439_ ;
	wire _w4438_ ;
	wire _w4437_ ;
	wire _w4436_ ;
	wire _w4435_ ;
	wire _w4434_ ;
	wire _w4433_ ;
	wire _w4432_ ;
	wire _w4431_ ;
	wire _w4430_ ;
	wire _w4429_ ;
	wire _w4428_ ;
	wire _w4427_ ;
	wire _w4426_ ;
	wire _w4425_ ;
	wire _w4424_ ;
	wire _w4423_ ;
	wire _w4422_ ;
	wire _w4421_ ;
	wire _w4420_ ;
	wire _w4419_ ;
	wire _w4418_ ;
	wire _w4417_ ;
	wire _w4416_ ;
	wire _w4415_ ;
	wire _w4414_ ;
	wire _w4413_ ;
	wire _w4412_ ;
	wire _w4411_ ;
	wire _w4410_ ;
	wire _w4409_ ;
	wire _w4408_ ;
	wire _w4407_ ;
	wire _w4406_ ;
	wire _w4405_ ;
	wire _w4404_ ;
	wire _w4403_ ;
	wire _w4402_ ;
	wire _w4401_ ;
	wire _w4400_ ;
	wire _w4399_ ;
	wire _w4398_ ;
	wire _w4397_ ;
	wire _w4396_ ;
	wire _w4395_ ;
	wire _w4394_ ;
	wire _w4393_ ;
	wire _w4392_ ;
	wire _w4391_ ;
	wire _w4390_ ;
	wire _w4389_ ;
	wire _w4388_ ;
	wire _w4387_ ;
	wire _w4386_ ;
	wire _w4385_ ;
	wire _w4384_ ;
	wire _w4383_ ;
	wire _w4382_ ;
	wire _w4381_ ;
	wire _w4380_ ;
	wire _w4379_ ;
	wire _w4378_ ;
	wire _w4377_ ;
	wire _w4376_ ;
	wire _w4375_ ;
	wire _w4374_ ;
	wire _w4373_ ;
	wire _w4372_ ;
	wire _w4371_ ;
	wire _w4370_ ;
	wire _w4369_ ;
	wire _w4368_ ;
	wire _w4367_ ;
	wire _w4366_ ;
	wire _w4365_ ;
	wire _w4364_ ;
	wire _w4363_ ;
	wire _w4362_ ;
	wire _w4361_ ;
	wire _w4360_ ;
	wire _w4359_ ;
	wire _w4358_ ;
	wire _w4357_ ;
	wire _w4356_ ;
	wire _w4355_ ;
	wire _w4354_ ;
	wire _w4353_ ;
	wire _w4352_ ;
	wire _w4351_ ;
	wire _w4350_ ;
	wire _w4349_ ;
	wire _w4348_ ;
	wire _w4347_ ;
	wire _w4346_ ;
	wire _w4345_ ;
	wire _w4344_ ;
	wire _w4343_ ;
	wire _w4342_ ;
	wire _w4341_ ;
	wire _w4340_ ;
	wire _w4339_ ;
	wire _w4338_ ;
	wire _w4337_ ;
	wire _w4336_ ;
	wire _w4335_ ;
	wire _w4334_ ;
	wire _w4333_ ;
	wire _w4332_ ;
	wire _w4331_ ;
	wire _w4330_ ;
	wire _w4329_ ;
	wire _w4328_ ;
	wire _w4327_ ;
	wire _w4326_ ;
	wire _w4325_ ;
	wire _w4324_ ;
	wire _w4323_ ;
	wire _w4322_ ;
	wire _w4321_ ;
	wire _w4320_ ;
	wire _w4319_ ;
	wire _w4318_ ;
	wire _w4317_ ;
	wire _w4316_ ;
	wire _w4315_ ;
	wire _w4314_ ;
	wire _w4313_ ;
	wire _w4312_ ;
	wire _w4311_ ;
	wire _w4310_ ;
	wire _w4309_ ;
	wire _w4308_ ;
	wire _w4307_ ;
	wire _w4306_ ;
	wire _w4305_ ;
	wire _w4304_ ;
	wire _w4303_ ;
	wire _w4302_ ;
	wire _w4301_ ;
	wire _w4300_ ;
	wire _w4299_ ;
	wire _w4298_ ;
	wire _w4297_ ;
	wire _w4296_ ;
	wire _w4295_ ;
	wire _w4294_ ;
	wire _w4293_ ;
	wire _w4292_ ;
	wire _w4291_ ;
	wire _w4290_ ;
	wire _w4289_ ;
	wire _w4288_ ;
	wire _w4287_ ;
	wire _w4286_ ;
	wire _w4285_ ;
	wire _w4284_ ;
	wire _w4283_ ;
	wire _w4282_ ;
	wire _w4281_ ;
	wire _w4280_ ;
	wire _w4279_ ;
	wire _w4278_ ;
	wire _w4277_ ;
	wire _w4276_ ;
	wire _w4275_ ;
	wire _w4274_ ;
	wire _w4273_ ;
	wire _w4272_ ;
	wire _w4271_ ;
	wire _w4270_ ;
	wire _w4269_ ;
	wire _w4268_ ;
	wire _w4267_ ;
	wire _w4266_ ;
	wire _w4265_ ;
	wire _w4264_ ;
	wire _w4263_ ;
	wire _w4262_ ;
	wire _w4261_ ;
	wire _w4260_ ;
	wire _w4259_ ;
	wire _w4258_ ;
	wire _w4257_ ;
	wire _w4256_ ;
	wire _w4255_ ;
	wire _w4254_ ;
	wire _w4253_ ;
	wire _w4252_ ;
	wire _w4251_ ;
	wire _w4250_ ;
	wire _w4249_ ;
	wire _w4248_ ;
	wire _w4247_ ;
	wire _w4246_ ;
	wire _w4245_ ;
	wire _w4244_ ;
	wire _w4243_ ;
	wire _w4242_ ;
	wire _w4241_ ;
	wire _w4240_ ;
	wire _w4239_ ;
	wire _w4238_ ;
	wire _w4237_ ;
	wire _w4236_ ;
	wire _w4235_ ;
	wire _w4234_ ;
	wire _w4233_ ;
	wire _w4232_ ;
	wire _w4231_ ;
	wire _w4230_ ;
	wire _w4229_ ;
	wire _w4228_ ;
	wire _w4227_ ;
	wire _w4226_ ;
	wire _w4225_ ;
	wire _w4224_ ;
	wire _w4223_ ;
	wire _w4222_ ;
	wire _w4221_ ;
	wire _w4220_ ;
	wire _w4219_ ;
	wire _w4218_ ;
	wire _w4217_ ;
	wire _w4216_ ;
	wire _w4215_ ;
	wire _w4214_ ;
	wire _w4213_ ;
	wire _w4212_ ;
	wire _w4211_ ;
	wire _w4210_ ;
	wire _w4209_ ;
	wire _w4208_ ;
	wire _w4207_ ;
	wire _w4206_ ;
	wire _w4205_ ;
	wire _w4204_ ;
	wire _w4203_ ;
	wire _w4202_ ;
	wire _w4201_ ;
	wire _w4200_ ;
	wire _w4199_ ;
	wire _w4198_ ;
	wire _w4197_ ;
	wire _w4196_ ;
	wire _w4195_ ;
	wire _w4194_ ;
	wire _w4193_ ;
	wire _w4192_ ;
	wire _w4191_ ;
	wire _w4190_ ;
	wire _w4189_ ;
	wire _w4188_ ;
	wire _w4187_ ;
	wire _w4186_ ;
	wire _w4185_ ;
	wire _w4184_ ;
	wire _w4183_ ;
	wire _w4182_ ;
	wire _w4181_ ;
	wire _w4180_ ;
	wire _w4179_ ;
	wire _w4178_ ;
	wire _w4177_ ;
	wire _w4176_ ;
	wire _w4175_ ;
	wire _w4174_ ;
	wire _w4173_ ;
	wire _w4172_ ;
	wire _w4171_ ;
	wire _w4170_ ;
	wire _w4169_ ;
	wire _w4168_ ;
	wire _w4167_ ;
	wire _w4166_ ;
	wire _w4165_ ;
	wire _w4164_ ;
	wire _w4163_ ;
	wire _w4162_ ;
	wire _w4161_ ;
	wire _w4160_ ;
	wire _w4159_ ;
	wire _w4158_ ;
	wire _w4157_ ;
	wire _w4156_ ;
	wire _w4155_ ;
	wire _w4154_ ;
	wire _w4153_ ;
	wire _w4152_ ;
	wire _w4151_ ;
	wire _w4150_ ;
	wire _w4149_ ;
	wire _w4148_ ;
	wire _w4147_ ;
	wire _w4146_ ;
	wire _w4145_ ;
	wire _w4144_ ;
	wire _w4143_ ;
	wire _w4142_ ;
	wire _w4141_ ;
	wire _w4140_ ;
	wire _w4139_ ;
	wire _w4138_ ;
	wire _w4137_ ;
	wire _w4136_ ;
	wire _w4135_ ;
	wire _w4134_ ;
	wire _w4133_ ;
	wire _w4132_ ;
	wire _w4131_ ;
	wire _w4130_ ;
	wire _w4129_ ;
	wire _w4128_ ;
	wire _w4127_ ;
	wire _w4126_ ;
	wire _w4125_ ;
	wire _w4124_ ;
	wire _w4123_ ;
	wire _w4122_ ;
	wire _w4121_ ;
	wire _w4120_ ;
	wire _w4119_ ;
	wire _w4118_ ;
	wire _w4117_ ;
	wire _w4116_ ;
	wire _w4115_ ;
	wire _w4114_ ;
	wire _w4113_ ;
	wire _w4112_ ;
	wire _w4111_ ;
	wire _w4110_ ;
	wire _w4109_ ;
	wire _w4108_ ;
	wire _w4107_ ;
	wire _w4106_ ;
	wire _w4105_ ;
	wire _w4104_ ;
	wire _w4103_ ;
	wire _w4102_ ;
	wire _w4101_ ;
	wire _w4100_ ;
	wire _w4099_ ;
	wire _w4098_ ;
	wire _w4097_ ;
	wire _w4096_ ;
	wire _w4095_ ;
	wire _w4094_ ;
	wire _w4093_ ;
	wire _w4092_ ;
	wire _w4091_ ;
	wire _w4090_ ;
	wire _w4089_ ;
	wire _w4088_ ;
	wire _w4087_ ;
	wire _w4086_ ;
	wire _w4085_ ;
	wire _w4084_ ;
	wire _w4083_ ;
	wire _w4082_ ;
	wire _w4081_ ;
	wire _w4080_ ;
	wire _w4079_ ;
	wire _w4078_ ;
	wire _w4077_ ;
	wire _w4076_ ;
	wire _w4075_ ;
	wire _w4074_ ;
	wire _w4073_ ;
	wire _w4072_ ;
	wire _w4071_ ;
	wire _w4070_ ;
	wire _w4069_ ;
	wire _w4068_ ;
	wire _w4067_ ;
	wire _w4066_ ;
	wire _w4065_ ;
	wire _w4064_ ;
	wire _w4063_ ;
	wire _w4062_ ;
	wire _w4061_ ;
	wire _w4060_ ;
	wire _w4059_ ;
	wire _w4058_ ;
	wire _w4057_ ;
	wire _w4056_ ;
	wire _w4055_ ;
	wire _w4054_ ;
	wire _w4053_ ;
	wire _w4052_ ;
	wire _w4051_ ;
	wire _w4050_ ;
	wire _w4049_ ;
	wire _w4048_ ;
	wire _w4047_ ;
	wire _w4046_ ;
	wire _w4045_ ;
	wire _w4044_ ;
	wire _w4043_ ;
	wire _w4042_ ;
	wire _w4041_ ;
	wire _w4040_ ;
	wire _w4039_ ;
	wire _w4038_ ;
	wire _w4037_ ;
	wire _w4036_ ;
	wire _w4035_ ;
	wire _w4034_ ;
	wire _w4033_ ;
	wire _w4032_ ;
	wire _w4031_ ;
	wire _w4030_ ;
	wire _w4029_ ;
	wire _w4028_ ;
	wire _w4027_ ;
	wire _w4026_ ;
	wire _w4025_ ;
	wire _w4024_ ;
	wire _w4023_ ;
	wire _w4022_ ;
	wire _w4021_ ;
	wire _w4020_ ;
	wire _w4019_ ;
	wire _w4018_ ;
	wire _w4017_ ;
	wire _w4016_ ;
	wire _w4015_ ;
	wire _w4014_ ;
	wire _w4013_ ;
	wire _w4012_ ;
	wire _w4011_ ;
	wire _w4010_ ;
	wire _w4009_ ;
	wire _w4008_ ;
	wire _w4007_ ;
	wire _w4006_ ;
	wire _w4005_ ;
	wire _w4004_ ;
	wire _w4003_ ;
	wire _w4002_ ;
	wire _w4001_ ;
	wire _w4000_ ;
	wire _w3999_ ;
	wire _w3998_ ;
	wire _w3997_ ;
	wire _w3996_ ;
	wire _w3995_ ;
	wire _w3994_ ;
	wire _w3993_ ;
	wire _w3992_ ;
	wire _w3991_ ;
	wire _w3990_ ;
	wire _w3989_ ;
	wire _w3988_ ;
	wire _w3987_ ;
	wire _w3986_ ;
	wire _w3985_ ;
	wire _w3984_ ;
	wire _w3983_ ;
	wire _w3982_ ;
	wire _w3981_ ;
	wire _w3980_ ;
	wire _w3979_ ;
	wire _w3978_ ;
	wire _w3977_ ;
	wire _w3976_ ;
	wire _w3975_ ;
	wire _w3974_ ;
	wire _w3973_ ;
	wire _w3972_ ;
	wire _w3971_ ;
	wire _w3970_ ;
	wire _w3969_ ;
	wire _w3968_ ;
	wire _w3967_ ;
	wire _w3966_ ;
	wire _w3965_ ;
	wire _w3964_ ;
	wire _w3963_ ;
	wire _w3962_ ;
	wire _w3961_ ;
	wire _w3960_ ;
	wire _w3959_ ;
	wire _w3958_ ;
	wire _w3957_ ;
	wire _w3956_ ;
	wire _w3955_ ;
	wire _w3954_ ;
	wire _w3953_ ;
	wire _w3952_ ;
	wire _w3951_ ;
	wire _w3950_ ;
	wire _w3949_ ;
	wire _w3948_ ;
	wire _w3947_ ;
	wire _w3946_ ;
	wire _w3945_ ;
	wire _w3944_ ;
	wire _w3943_ ;
	wire _w3942_ ;
	wire _w3941_ ;
	wire _w3940_ ;
	wire _w3939_ ;
	wire _w3938_ ;
	wire _w3937_ ;
	wire _w3936_ ;
	wire _w3935_ ;
	wire _w3934_ ;
	wire _w3933_ ;
	wire _w3932_ ;
	wire _w3931_ ;
	wire _w3930_ ;
	wire _w3929_ ;
	wire _w3928_ ;
	wire _w3927_ ;
	wire _w3926_ ;
	wire _w3925_ ;
	wire _w3924_ ;
	wire _w3923_ ;
	wire _w3922_ ;
	wire _w3921_ ;
	wire _w3920_ ;
	wire _w3919_ ;
	wire _w3918_ ;
	wire _w3917_ ;
	wire _w3916_ ;
	wire _w3915_ ;
	wire _w3914_ ;
	wire _w3913_ ;
	wire _w3912_ ;
	wire _w3911_ ;
	wire _w3910_ ;
	wire _w3909_ ;
	wire _w3908_ ;
	wire _w3907_ ;
	wire _w3906_ ;
	wire _w3905_ ;
	wire _w3904_ ;
	wire _w3903_ ;
	wire _w3902_ ;
	wire _w3901_ ;
	wire _w3900_ ;
	wire _w3899_ ;
	wire _w3898_ ;
	wire _w3897_ ;
	wire _w3896_ ;
	wire _w3895_ ;
	wire _w3894_ ;
	wire _w3893_ ;
	wire _w3892_ ;
	wire _w3891_ ;
	wire _w3890_ ;
	wire _w3889_ ;
	wire _w3888_ ;
	wire _w3887_ ;
	wire _w3886_ ;
	wire _w3885_ ;
	wire _w3884_ ;
	wire _w3883_ ;
	wire _w3882_ ;
	wire _w3881_ ;
	wire _w3880_ ;
	wire _w3879_ ;
	wire _w3878_ ;
	wire _w3877_ ;
	wire _w3876_ ;
	wire _w3875_ ;
	wire _w3874_ ;
	wire _w3873_ ;
	wire _w3872_ ;
	wire _w3871_ ;
	wire _w3870_ ;
	wire _w3869_ ;
	wire _w3868_ ;
	wire _w3867_ ;
	wire _w3866_ ;
	wire _w3865_ ;
	wire _w3864_ ;
	wire _w3863_ ;
	wire _w3862_ ;
	wire _w3861_ ;
	wire _w3860_ ;
	wire _w3859_ ;
	wire _w3858_ ;
	wire _w3857_ ;
	wire _w3856_ ;
	wire _w3855_ ;
	wire _w3854_ ;
	wire _w3853_ ;
	wire _w3852_ ;
	wire _w3851_ ;
	wire _w3850_ ;
	wire _w3849_ ;
	wire _w3848_ ;
	wire _w3847_ ;
	wire _w3846_ ;
	wire _w3845_ ;
	wire _w3844_ ;
	wire _w3843_ ;
	wire _w3842_ ;
	wire _w3841_ ;
	wire _w3840_ ;
	wire _w3839_ ;
	wire _w3838_ ;
	wire _w3837_ ;
	wire _w3836_ ;
	wire _w3835_ ;
	wire _w3834_ ;
	wire _w3833_ ;
	wire _w3832_ ;
	wire _w3831_ ;
	wire _w3830_ ;
	wire _w3829_ ;
	wire _w3828_ ;
	wire _w3827_ ;
	wire _w3826_ ;
	wire _w3825_ ;
	wire _w3824_ ;
	wire _w3823_ ;
	wire _w3822_ ;
	wire _w3821_ ;
	wire _w3820_ ;
	wire _w3819_ ;
	wire _w3818_ ;
	wire _w3817_ ;
	wire _w3816_ ;
	wire _w3815_ ;
	wire _w3814_ ;
	wire _w3813_ ;
	wire _w3812_ ;
	wire _w3811_ ;
	wire _w3810_ ;
	wire _w3809_ ;
	wire _w3808_ ;
	wire _w3807_ ;
	wire _w3806_ ;
	wire _w3805_ ;
	wire _w3804_ ;
	wire _w3803_ ;
	wire _w3802_ ;
	wire _w3801_ ;
	wire _w3800_ ;
	wire _w3799_ ;
	wire _w3798_ ;
	wire _w3797_ ;
	wire _w3796_ ;
	wire _w3795_ ;
	wire _w3794_ ;
	wire _w3793_ ;
	wire _w3792_ ;
	wire _w3791_ ;
	wire _w3790_ ;
	wire _w3789_ ;
	wire _w3788_ ;
	wire _w3787_ ;
	wire _w3786_ ;
	wire _w3785_ ;
	wire _w3784_ ;
	wire _w3783_ ;
	wire _w3782_ ;
	wire _w3781_ ;
	wire _w3780_ ;
	wire _w3779_ ;
	wire _w3778_ ;
	wire _w3777_ ;
	wire _w3776_ ;
	wire _w3775_ ;
	wire _w3774_ ;
	wire _w3773_ ;
	wire _w3772_ ;
	wire _w3771_ ;
	wire _w3770_ ;
	wire _w3769_ ;
	wire _w3768_ ;
	wire _w3767_ ;
	wire _w3766_ ;
	wire _w3765_ ;
	wire _w3764_ ;
	wire _w3763_ ;
	wire _w3762_ ;
	wire _w3761_ ;
	wire _w3760_ ;
	wire _w3759_ ;
	wire _w3758_ ;
	wire _w3757_ ;
	wire _w3756_ ;
	wire _w3755_ ;
	wire _w3754_ ;
	wire _w3753_ ;
	wire _w3752_ ;
	wire _w3751_ ;
	wire _w3750_ ;
	wire _w3749_ ;
	wire _w3748_ ;
	wire _w3747_ ;
	wire _w3746_ ;
	wire _w3745_ ;
	wire _w3744_ ;
	wire _w3743_ ;
	wire _w3742_ ;
	wire _w3741_ ;
	wire _w3740_ ;
	wire _w3739_ ;
	wire _w3738_ ;
	wire _w3737_ ;
	wire _w3736_ ;
	wire _w3735_ ;
	wire _w3734_ ;
	wire _w3733_ ;
	wire _w3732_ ;
	wire _w3731_ ;
	wire _w3730_ ;
	wire _w3729_ ;
	wire _w3728_ ;
	wire _w3727_ ;
	wire _w3726_ ;
	wire _w3725_ ;
	wire _w3724_ ;
	wire _w3723_ ;
	wire _w3722_ ;
	wire _w3721_ ;
	wire _w3720_ ;
	wire _w3719_ ;
	wire _w3718_ ;
	wire _w3717_ ;
	wire _w3716_ ;
	wire _w3715_ ;
	wire _w3714_ ;
	wire _w3713_ ;
	wire _w3712_ ;
	wire _w3711_ ;
	wire _w3710_ ;
	wire _w3709_ ;
	wire _w3708_ ;
	wire _w3707_ ;
	wire _w3706_ ;
	wire _w3705_ ;
	wire _w3704_ ;
	wire _w3703_ ;
	wire _w3702_ ;
	wire _w3701_ ;
	wire _w3700_ ;
	wire _w3699_ ;
	wire _w3698_ ;
	wire _w3697_ ;
	wire _w3696_ ;
	wire _w3695_ ;
	wire _w3694_ ;
	wire _w3693_ ;
	wire _w3692_ ;
	wire _w3691_ ;
	wire _w3690_ ;
	wire _w3689_ ;
	wire _w3688_ ;
	wire _w3687_ ;
	wire _w3686_ ;
	wire _w3685_ ;
	wire _w3684_ ;
	wire _w3683_ ;
	wire _w3682_ ;
	wire _w3681_ ;
	wire _w3680_ ;
	wire _w3679_ ;
	wire _w3678_ ;
	wire _w3677_ ;
	wire _w3676_ ;
	wire _w3675_ ;
	wire _w3674_ ;
	wire _w3673_ ;
	wire _w3672_ ;
	wire _w3671_ ;
	wire _w3670_ ;
	wire _w3669_ ;
	wire _w3668_ ;
	wire _w3667_ ;
	wire _w3666_ ;
	wire _w3665_ ;
	wire _w3664_ ;
	wire _w3663_ ;
	wire _w3662_ ;
	wire _w3661_ ;
	wire _w3660_ ;
	wire _w3659_ ;
	wire _w3658_ ;
	wire _w3657_ ;
	wire _w3656_ ;
	wire _w3655_ ;
	wire _w3654_ ;
	wire _w3653_ ;
	wire _w3652_ ;
	wire _w3651_ ;
	wire _w3650_ ;
	wire _w3649_ ;
	wire _w3648_ ;
	wire _w3647_ ;
	wire _w3646_ ;
	wire _w3645_ ;
	wire _w3644_ ;
	wire _w3643_ ;
	wire _w3642_ ;
	wire _w3641_ ;
	wire _w3640_ ;
	wire _w3639_ ;
	wire _w3638_ ;
	wire _w3637_ ;
	wire _w3636_ ;
	wire _w3635_ ;
	wire _w3634_ ;
	wire _w3633_ ;
	wire _w3632_ ;
	wire _w3631_ ;
	wire _w3630_ ;
	wire _w3629_ ;
	wire _w3628_ ;
	wire _w3627_ ;
	wire _w3626_ ;
	wire _w3625_ ;
	wire _w3624_ ;
	wire _w3623_ ;
	wire _w3622_ ;
	wire _w3621_ ;
	wire _w3620_ ;
	wire _w3619_ ;
	wire _w3618_ ;
	wire _w3617_ ;
	wire _w3616_ ;
	wire _w3615_ ;
	wire _w3614_ ;
	wire _w3613_ ;
	wire _w3612_ ;
	wire _w3611_ ;
	wire _w3610_ ;
	wire _w3609_ ;
	wire _w3608_ ;
	wire _w3607_ ;
	wire _w3606_ ;
	wire _w3605_ ;
	wire _w3604_ ;
	wire _w3603_ ;
	wire _w3602_ ;
	wire _w3601_ ;
	wire _w3600_ ;
	wire _w3599_ ;
	wire _w3598_ ;
	wire _w3597_ ;
	wire _w3596_ ;
	wire _w3595_ ;
	wire _w3594_ ;
	wire _w3593_ ;
	wire _w3592_ ;
	wire _w3591_ ;
	wire _w3590_ ;
	wire _w3589_ ;
	wire _w3588_ ;
	wire _w3587_ ;
	wire _w3586_ ;
	wire _w3585_ ;
	wire _w3584_ ;
	wire _w3583_ ;
	wire _w3582_ ;
	wire _w3581_ ;
	wire _w3580_ ;
	wire _w3579_ ;
	wire _w3578_ ;
	wire _w3577_ ;
	wire _w3576_ ;
	wire _w3575_ ;
	wire _w3574_ ;
	wire _w3573_ ;
	wire _w3572_ ;
	wire _w3571_ ;
	wire _w3570_ ;
	wire _w3569_ ;
	wire _w3568_ ;
	wire _w3567_ ;
	wire _w3566_ ;
	wire _w3565_ ;
	wire _w3564_ ;
	wire _w3563_ ;
	wire _w3562_ ;
	wire _w3561_ ;
	wire _w3560_ ;
	wire _w3559_ ;
	wire _w3558_ ;
	wire _w3557_ ;
	wire _w3556_ ;
	wire _w3555_ ;
	wire _w3554_ ;
	wire _w3553_ ;
	wire _w3552_ ;
	wire _w3551_ ;
	wire _w3550_ ;
	wire _w3549_ ;
	wire _w3548_ ;
	wire _w3547_ ;
	wire _w3546_ ;
	wire _w3545_ ;
	wire _w3544_ ;
	wire _w3543_ ;
	wire _w3542_ ;
	wire _w3541_ ;
	wire _w3540_ ;
	wire _w3539_ ;
	wire _w3538_ ;
	wire _w3537_ ;
	wire _w3536_ ;
	wire _w3535_ ;
	wire _w3534_ ;
	wire _w3533_ ;
	wire _w3532_ ;
	wire _w3531_ ;
	wire _w3530_ ;
	wire _w3529_ ;
	wire _w3528_ ;
	wire _w3527_ ;
	wire _w3526_ ;
	wire _w3525_ ;
	wire _w3524_ ;
	wire _w3523_ ;
	wire _w3522_ ;
	wire _w3521_ ;
	wire _w3520_ ;
	wire _w3519_ ;
	wire _w3518_ ;
	wire _w3517_ ;
	wire _w3516_ ;
	wire _w3515_ ;
	wire _w3514_ ;
	wire _w3513_ ;
	wire _w3512_ ;
	wire _w3511_ ;
	wire _w3510_ ;
	wire _w3509_ ;
	wire _w3508_ ;
	wire _w3507_ ;
	wire _w3506_ ;
	wire _w3505_ ;
	wire _w3504_ ;
	wire _w3503_ ;
	wire _w3502_ ;
	wire _w3501_ ;
	wire _w3500_ ;
	wire _w3499_ ;
	wire _w3498_ ;
	wire _w3497_ ;
	wire _w3496_ ;
	wire _w3495_ ;
	wire _w3494_ ;
	wire _w3493_ ;
	wire _w3492_ ;
	wire _w3491_ ;
	wire _w3490_ ;
	wire _w3489_ ;
	wire _w3488_ ;
	wire _w3487_ ;
	wire _w3486_ ;
	wire _w3485_ ;
	wire _w3484_ ;
	wire _w3483_ ;
	wire _w3482_ ;
	wire _w3481_ ;
	wire _w3480_ ;
	wire _w3479_ ;
	wire _w3478_ ;
	wire _w3477_ ;
	wire _w3476_ ;
	wire _w3475_ ;
	wire _w3474_ ;
	wire _w3473_ ;
	wire _w3472_ ;
	wire _w3471_ ;
	wire _w3470_ ;
	wire _w3469_ ;
	wire _w3468_ ;
	wire _w3467_ ;
	wire _w3466_ ;
	wire _w3465_ ;
	wire _w3464_ ;
	wire _w3463_ ;
	wire _w3462_ ;
	wire _w3461_ ;
	wire _w3460_ ;
	wire _w3459_ ;
	wire _w3458_ ;
	wire _w3457_ ;
	wire _w3456_ ;
	wire _w3455_ ;
	wire _w3454_ ;
	wire _w3453_ ;
	wire _w3452_ ;
	wire _w3451_ ;
	wire _w3450_ ;
	wire _w3449_ ;
	wire _w3448_ ;
	wire _w3447_ ;
	wire _w3446_ ;
	wire _w3445_ ;
	wire _w3444_ ;
	wire _w3443_ ;
	wire _w3442_ ;
	wire _w3441_ ;
	wire _w3440_ ;
	wire _w3439_ ;
	wire _w3438_ ;
	wire _w3437_ ;
	wire _w3436_ ;
	wire _w3435_ ;
	wire _w3434_ ;
	wire _w3433_ ;
	wire _w3432_ ;
	wire _w3431_ ;
	wire _w3430_ ;
	wire _w3429_ ;
	wire _w3428_ ;
	wire _w3427_ ;
	wire _w3426_ ;
	wire _w3425_ ;
	wire _w3424_ ;
	wire _w3423_ ;
	wire _w3422_ ;
	wire _w3421_ ;
	wire _w3420_ ;
	wire _w3419_ ;
	wire _w3418_ ;
	wire _w3417_ ;
	wire _w3416_ ;
	wire _w3415_ ;
	wire _w3414_ ;
	wire _w3413_ ;
	wire _w3412_ ;
	wire _w3411_ ;
	wire _w3410_ ;
	wire _w3409_ ;
	wire _w3408_ ;
	wire _w3407_ ;
	wire _w3406_ ;
	wire _w3405_ ;
	wire _w3404_ ;
	wire _w3403_ ;
	wire _w3402_ ;
	wire _w3401_ ;
	wire _w3400_ ;
	wire _w3399_ ;
	wire _w3398_ ;
	wire _w3397_ ;
	wire _w3396_ ;
	wire _w3395_ ;
	wire _w3394_ ;
	wire _w3393_ ;
	wire _w3392_ ;
	wire _w3391_ ;
	wire _w3390_ ;
	wire _w3389_ ;
	wire _w3388_ ;
	wire _w3387_ ;
	wire _w3386_ ;
	wire _w3385_ ;
	wire _w3384_ ;
	wire _w3383_ ;
	wire _w3382_ ;
	wire _w3381_ ;
	wire _w3380_ ;
	wire _w3379_ ;
	wire _w3378_ ;
	wire _w3377_ ;
	wire _w3376_ ;
	wire _w3375_ ;
	wire _w3374_ ;
	wire _w3373_ ;
	wire _w3372_ ;
	wire _w3371_ ;
	wire _w3370_ ;
	wire _w3369_ ;
	wire _w3368_ ;
	wire _w3367_ ;
	wire _w3366_ ;
	wire _w3365_ ;
	wire _w3364_ ;
	wire _w3363_ ;
	wire _w3362_ ;
	wire _w3361_ ;
	wire _w3360_ ;
	wire _w3359_ ;
	wire _w3358_ ;
	wire _w3357_ ;
	wire _w3356_ ;
	wire _w3355_ ;
	wire _w3354_ ;
	wire _w3353_ ;
	wire _w3352_ ;
	wire _w3351_ ;
	wire _w3350_ ;
	wire _w3349_ ;
	wire _w3348_ ;
	wire _w3347_ ;
	wire _w3346_ ;
	wire _w3345_ ;
	wire _w3344_ ;
	wire _w3343_ ;
	wire _w3342_ ;
	wire _w3341_ ;
	wire _w3340_ ;
	wire _w3339_ ;
	wire _w3338_ ;
	wire _w3337_ ;
	wire _w3336_ ;
	wire _w3335_ ;
	wire _w3334_ ;
	wire _w3333_ ;
	wire _w3332_ ;
	wire _w3331_ ;
	wire _w3330_ ;
	wire _w3329_ ;
	wire _w3328_ ;
	wire _w3327_ ;
	wire _w3326_ ;
	wire _w3325_ ;
	wire _w3324_ ;
	wire _w3323_ ;
	wire _w3322_ ;
	wire _w3321_ ;
	wire _w3320_ ;
	wire _w3319_ ;
	wire _w3318_ ;
	wire _w3317_ ;
	wire _w2068_ ;
	wire _w2067_ ;
	wire _w2066_ ;
	wire _w2065_ ;
	wire _w2064_ ;
	wire _w2063_ ;
	wire _w2062_ ;
	wire _w2061_ ;
	wire _w2060_ ;
	wire _w2059_ ;
	wire _w2058_ ;
	wire _w2057_ ;
	wire _w2056_ ;
	wire _w2055_ ;
	wire _w2054_ ;
	wire _w2053_ ;
	wire _w2052_ ;
	wire _w2051_ ;
	wire _w2050_ ;
	wire _w2049_ ;
	wire _w2048_ ;
	wire _w2047_ ;
	wire _w2046_ ;
	wire _w2045_ ;
	wire _w2044_ ;
	wire _w2043_ ;
	wire _w2042_ ;
	wire _w2041_ ;
	wire _w2040_ ;
	wire _w2039_ ;
	wire _w2038_ ;
	wire _w2037_ ;
	wire _w2036_ ;
	wire _w2035_ ;
	wire _w2034_ ;
	wire _w2033_ ;
	wire _w2032_ ;
	wire _w2031_ ;
	wire _w2030_ ;
	wire _w2029_ ;
	wire _w2028_ ;
	wire _w2027_ ;
	wire _w2026_ ;
	wire _w2025_ ;
	wire _w2024_ ;
	wire _w2023_ ;
	wire _w2022_ ;
	wire _w2021_ ;
	wire _w2020_ ;
	wire _w2019_ ;
	wire _w2018_ ;
	wire _w2017_ ;
	wire _w2016_ ;
	wire _w2015_ ;
	wire _w2014_ ;
	wire _w2013_ ;
	wire _w2012_ ;
	wire _w2011_ ;
	wire _w2010_ ;
	wire _w2009_ ;
	wire _w2008_ ;
	wire _w2007_ ;
	wire _w2006_ ;
	wire _w2005_ ;
	wire _w2004_ ;
	wire _w2003_ ;
	wire _w2002_ ;
	wire _w2001_ ;
	wire _w2000_ ;
	wire _w1999_ ;
	wire _w1998_ ;
	wire _w1997_ ;
	wire _w1996_ ;
	wire _w1995_ ;
	wire _w1994_ ;
	wire _w1993_ ;
	wire _w1992_ ;
	wire _w1991_ ;
	wire _w1990_ ;
	wire _w1989_ ;
	wire _w1988_ ;
	wire _w1987_ ;
	wire _w1986_ ;
	wire _w1985_ ;
	wire _w1984_ ;
	wire _w1983_ ;
	wire _w1982_ ;
	wire _w1981_ ;
	wire _w1980_ ;
	wire _w1979_ ;
	wire _w1978_ ;
	wire _w1977_ ;
	wire _w1976_ ;
	wire _w1975_ ;
	wire _w1974_ ;
	wire _w1973_ ;
	wire _w1972_ ;
	wire _w1971_ ;
	wire _w1970_ ;
	wire _w1969_ ;
	wire _w1968_ ;
	wire _w1967_ ;
	wire _w1966_ ;
	wire _w1965_ ;
	wire _w1964_ ;
	wire _w1963_ ;
	wire _w1962_ ;
	wire _w1961_ ;
	wire _w1960_ ;
	wire _w1959_ ;
	wire _w1958_ ;
	wire _w1957_ ;
	wire _w1956_ ;
	wire _w1955_ ;
	wire _w1954_ ;
	wire _w1953_ ;
	wire _w1952_ ;
	wire _w1951_ ;
	wire _w1950_ ;
	wire _w1949_ ;
	wire _w1948_ ;
	wire _w1947_ ;
	wire _w1946_ ;
	wire _w1945_ ;
	wire _w1944_ ;
	wire _w1943_ ;
	wire _w1942_ ;
	wire _w1941_ ;
	wire _w1940_ ;
	wire _w1939_ ;
	wire _w1938_ ;
	wire _w1937_ ;
	wire _w1936_ ;
	wire _w1935_ ;
	wire _w1934_ ;
	wire _w1933_ ;
	wire _w1932_ ;
	wire _w1931_ ;
	wire _w1930_ ;
	wire _w1929_ ;
	wire _w1928_ ;
	wire _w1927_ ;
	wire _w1926_ ;
	wire _w1925_ ;
	wire _w1924_ ;
	wire _w1923_ ;
	wire _w1922_ ;
	wire _w1921_ ;
	wire _w1920_ ;
	wire _w1919_ ;
	wire _w1918_ ;
	wire _w1917_ ;
	wire _w1916_ ;
	wire _w1915_ ;
	wire _w1914_ ;
	wire _w1913_ ;
	wire _w1912_ ;
	wire _w1911_ ;
	wire _w1910_ ;
	wire _w1909_ ;
	wire _w1908_ ;
	wire _w1907_ ;
	wire _w1906_ ;
	wire _w1905_ ;
	wire _w1904_ ;
	wire _w1903_ ;
	wire _w1902_ ;
	wire _w1901_ ;
	wire _w1900_ ;
	wire _w1899_ ;
	wire _w1898_ ;
	wire _w1897_ ;
	wire _w1896_ ;
	wire _w1895_ ;
	wire _w1894_ ;
	wire _w1893_ ;
	wire _w1892_ ;
	wire _w1891_ ;
	wire _w1890_ ;
	wire _w1889_ ;
	wire _w1888_ ;
	wire _w1887_ ;
	wire _w1886_ ;
	wire _w1885_ ;
	wire _w1884_ ;
	wire _w1883_ ;
	wire _w1882_ ;
	wire _w1881_ ;
	wire _w1880_ ;
	wire _w1879_ ;
	wire _w1878_ ;
	wire _w1877_ ;
	wire _w1876_ ;
	wire _w1875_ ;
	wire _w1874_ ;
	wire _w1873_ ;
	wire _w1872_ ;
	wire _w1871_ ;
	wire _w1870_ ;
	wire _w1869_ ;
	wire _w1868_ ;
	wire _w1867_ ;
	wire _w1866_ ;
	wire _w1865_ ;
	wire _w1864_ ;
	wire _w1863_ ;
	wire _w1862_ ;
	wire _w1861_ ;
	wire _w1860_ ;
	wire _w1859_ ;
	wire _w1858_ ;
	wire _w1857_ ;
	wire _w1856_ ;
	wire _w1855_ ;
	wire _w1854_ ;
	wire _w1853_ ;
	wire _w1852_ ;
	wire _w1851_ ;
	wire _w1850_ ;
	wire _w1849_ ;
	wire _w1847_ ;
	wire _w1846_ ;
	wire _w1845_ ;
	wire _w1844_ ;
	wire _w1843_ ;
	wire _w1842_ ;
	wire _w1841_ ;
	wire _w1840_ ;
	wire _w1839_ ;
	wire _w1838_ ;
	wire _w1837_ ;
	wire _w1836_ ;
	wire _w1835_ ;
	wire _w1834_ ;
	wire _w1833_ ;
	wire _w1832_ ;
	wire _w1831_ ;
	wire _w1830_ ;
	wire _w1829_ ;
	wire _w1828_ ;
	wire _w1827_ ;
	wire _w1826_ ;
	wire _w1825_ ;
	wire _w1824_ ;
	wire _w1823_ ;
	wire _w1822_ ;
	wire _w1821_ ;
	wire _w1820_ ;
	wire _w1819_ ;
	wire _w1818_ ;
	wire _w1817_ ;
	wire _w1816_ ;
	wire _w1815_ ;
	wire _w1814_ ;
	wire _w1813_ ;
	wire _w1812_ ;
	wire _w1811_ ;
	wire _w1810_ ;
	wire _w1809_ ;
	wire _w1808_ ;
	wire _w1807_ ;
	wire _w1806_ ;
	wire _w1805_ ;
	wire _w1804_ ;
	wire _w1803_ ;
	wire _w1802_ ;
	wire _w1801_ ;
	wire _w1800_ ;
	wire _w1799_ ;
	wire _w1798_ ;
	wire _w1797_ ;
	wire _w1796_ ;
	wire _w1795_ ;
	wire _w1794_ ;
	wire _w1793_ ;
	wire _w1792_ ;
	wire _w1791_ ;
	wire _w1790_ ;
	wire _w1789_ ;
	wire _w1788_ ;
	wire _w1787_ ;
	wire _w1786_ ;
	wire _w1785_ ;
	wire _w1784_ ;
	wire _w1783_ ;
	wire _w1782_ ;
	wire _w1781_ ;
	wire _w1780_ ;
	wire _w1779_ ;
	wire _w1778_ ;
	wire _w1777_ ;
	wire _w1776_ ;
	wire _w1775_ ;
	wire _w1774_ ;
	wire _w1773_ ;
	wire _w1772_ ;
	wire _w1771_ ;
	wire _w1770_ ;
	wire _w1769_ ;
	wire _w1768_ ;
	wire _w1767_ ;
	wire _w1766_ ;
	wire _w1765_ ;
	wire _w1764_ ;
	wire _w1763_ ;
	wire _w1762_ ;
	wire _w1761_ ;
	wire _w1760_ ;
	wire _w1759_ ;
	wire _w1758_ ;
	wire _w1757_ ;
	wire _w1756_ ;
	wire _w1755_ ;
	wire _w1754_ ;
	wire _w1753_ ;
	wire _w1752_ ;
	wire _w1751_ ;
	wire _w1750_ ;
	wire _w1749_ ;
	wire _w1748_ ;
	wire _w1747_ ;
	wire _w1746_ ;
	wire _w1745_ ;
	wire _w1744_ ;
	wire _w1743_ ;
	wire _w1742_ ;
	wire _w1741_ ;
	wire _w1740_ ;
	wire _w1739_ ;
	wire _w1738_ ;
	wire _w1737_ ;
	wire _w1736_ ;
	wire _w1735_ ;
	wire _w1734_ ;
	wire _w1733_ ;
	wire _w1732_ ;
	wire _w1731_ ;
	wire _w1730_ ;
	wire _w1729_ ;
	wire _w1728_ ;
	wire _w1727_ ;
	wire _w1726_ ;
	wire _w1725_ ;
	wire _w1724_ ;
	wire _w1723_ ;
	wire _w1722_ ;
	wire _w1721_ ;
	wire _w1720_ ;
	wire _w1719_ ;
	wire _w1718_ ;
	wire _w1717_ ;
	wire _w1716_ ;
	wire _w1715_ ;
	wire _w1714_ ;
	wire _w1713_ ;
	wire _w1712_ ;
	wire _w1711_ ;
	wire _w1710_ ;
	wire _w1709_ ;
	wire _w1708_ ;
	wire _w1707_ ;
	wire _w1706_ ;
	wire _w1705_ ;
	wire _w1704_ ;
	wire _w1703_ ;
	wire _w1702_ ;
	wire _w1701_ ;
	wire _w1700_ ;
	wire _w1699_ ;
	wire _w1698_ ;
	wire _w1697_ ;
	wire _w1696_ ;
	wire _w1695_ ;
	wire _w1694_ ;
	wire _w1693_ ;
	wire _w1692_ ;
	wire _w1691_ ;
	wire _w1690_ ;
	wire _w1689_ ;
	wire _w1688_ ;
	wire _w1687_ ;
	wire _w1686_ ;
	wire _w1685_ ;
	wire _w1684_ ;
	wire _w1683_ ;
	wire _w1682_ ;
	wire _w1681_ ;
	wire _w1680_ ;
	wire _w1679_ ;
	wire _w1678_ ;
	wire _w1677_ ;
	wire _w1676_ ;
	wire _w1675_ ;
	wire _w1674_ ;
	wire _w1673_ ;
	wire _w1672_ ;
	wire _w1671_ ;
	wire _w1670_ ;
	wire _w1669_ ;
	wire _w1668_ ;
	wire _w1667_ ;
	wire _w1666_ ;
	wire _w1665_ ;
	wire _w1664_ ;
	wire _w1663_ ;
	wire _w1662_ ;
	wire _w1661_ ;
	wire _w1660_ ;
	wire _w1659_ ;
	wire _w1658_ ;
	wire _w1657_ ;
	wire _w1656_ ;
	wire _w1655_ ;
	wire _w1654_ ;
	wire _w1653_ ;
	wire _w1652_ ;
	wire _w1651_ ;
	wire _w1650_ ;
	wire _w1649_ ;
	wire _w1648_ ;
	wire _w1647_ ;
	wire _w1646_ ;
	wire _w1645_ ;
	wire _w1644_ ;
	wire _w1643_ ;
	wire _w1642_ ;
	wire _w1641_ ;
	wire _w1640_ ;
	wire _w1639_ ;
	wire _w1638_ ;
	wire _w1637_ ;
	wire _w1636_ ;
	wire _w1635_ ;
	wire _w1634_ ;
	wire _w1633_ ;
	wire _w1632_ ;
	wire _w1631_ ;
	wire _w1630_ ;
	wire _w1629_ ;
	wire _w1628_ ;
	wire _w1627_ ;
	wire _w1626_ ;
	wire _w1625_ ;
	wire _w1624_ ;
	wire _w1623_ ;
	wire _w1622_ ;
	wire _w1621_ ;
	wire _w1620_ ;
	wire _w1619_ ;
	wire _w1618_ ;
	wire _w1617_ ;
	wire _w1616_ ;
	wire _w1615_ ;
	wire _w1614_ ;
	wire _w1613_ ;
	wire _w1612_ ;
	wire _w1611_ ;
	wire _w1610_ ;
	wire _w1609_ ;
	wire _w1608_ ;
	wire _w1607_ ;
	wire _w1606_ ;
	wire _w1605_ ;
	wire _w1604_ ;
	wire _w1603_ ;
	wire _w1602_ ;
	wire _w1601_ ;
	wire _w1600_ ;
	wire _w1599_ ;
	wire _w1598_ ;
	wire _w1597_ ;
	wire _w1596_ ;
	wire _w1595_ ;
	wire _w1594_ ;
	wire _w1593_ ;
	wire _w1592_ ;
	wire _w1591_ ;
	wire _w1590_ ;
	wire _w1589_ ;
	wire _w1588_ ;
	wire _w1587_ ;
	wire _w1586_ ;
	wire _w1585_ ;
	wire _w1584_ ;
	wire _w1583_ ;
	wire _w1582_ ;
	wire _w1581_ ;
	wire _w1580_ ;
	wire _w1579_ ;
	wire _w1578_ ;
	wire _w1577_ ;
	wire _w1576_ ;
	wire _w1575_ ;
	wire _w1574_ ;
	wire _w1573_ ;
	wire _w1572_ ;
	wire _w1571_ ;
	wire _w1570_ ;
	wire _w1569_ ;
	wire _w1568_ ;
	wire _w1567_ ;
	wire _w1566_ ;
	wire _w1565_ ;
	wire _w1564_ ;
	wire _w1563_ ;
	wire _w1562_ ;
	wire _w1561_ ;
	wire _w1560_ ;
	wire _w1559_ ;
	wire _w1558_ ;
	wire _w1557_ ;
	wire _w1556_ ;
	wire _w1555_ ;
	wire _w1554_ ;
	wire _w1553_ ;
	wire _w1552_ ;
	wire _w1551_ ;
	wire _w1550_ ;
	wire _w1549_ ;
	wire _w1548_ ;
	wire _w1547_ ;
	wire _w1546_ ;
	wire _w1545_ ;
	wire _w1544_ ;
	wire _w1543_ ;
	wire _w1542_ ;
	wire _w1541_ ;
	wire _w1540_ ;
	wire _w1539_ ;
	wire _w1538_ ;
	wire _w1537_ ;
	wire _w1536_ ;
	wire _w1535_ ;
	wire _w1534_ ;
	wire _w1533_ ;
	wire _w1532_ ;
	wire _w1531_ ;
	wire _w1530_ ;
	wire _w1529_ ;
	wire _w1528_ ;
	wire _w1527_ ;
	wire _w1526_ ;
	wire _w1525_ ;
	wire _w1524_ ;
	wire _w1523_ ;
	wire _w1522_ ;
	wire _w1521_ ;
	wire _w1520_ ;
	wire _w1519_ ;
	wire _w1518_ ;
	wire _w1517_ ;
	wire _w1516_ ;
	wire _w1515_ ;
	wire _w1514_ ;
	wire _w1513_ ;
	wire _w1512_ ;
	wire _w1511_ ;
	wire _w1510_ ;
	wire _w1509_ ;
	wire _w1508_ ;
	wire _w1507_ ;
	wire _w1506_ ;
	wire _w1505_ ;
	wire _w1504_ ;
	wire _w1503_ ;
	wire _w1502_ ;
	wire _w1501_ ;
	wire _w1216_ ;
	wire _w1215_ ;
	wire _w1214_ ;
	wire _w1213_ ;
	wire _w1212_ ;
	wire _w1211_ ;
	wire _w1210_ ;
	wire _w1209_ ;
	wire _w1208_ ;
	wire _w1207_ ;
	wire _w1206_ ;
	wire _w1205_ ;
	wire _w1204_ ;
	wire _w1203_ ;
	wire _w1202_ ;
	wire _w1201_ ;
	wire _w1200_ ;
	wire _w1199_ ;
	wire _w1198_ ;
	wire _w1197_ ;
	wire _w1196_ ;
	wire _w1195_ ;
	wire _w1194_ ;
	wire _w1193_ ;
	wire _w1192_ ;
	wire _w1191_ ;
	wire _w1190_ ;
	wire _w1189_ ;
	wire _w1188_ ;
	wire _w1187_ ;
	wire _w1186_ ;
	wire _w1185_ ;
	wire _w1184_ ;
	wire _w1183_ ;
	wire _w1182_ ;
	wire _w1181_ ;
	wire _w1180_ ;
	wire _w1179_ ;
	wire _w1178_ ;
	wire _w1177_ ;
	wire _w1176_ ;
	wire _w1175_ ;
	wire _w1174_ ;
	wire _w1173_ ;
	wire _w1172_ ;
	wire _w1171_ ;
	wire _w1170_ ;
	wire _w1169_ ;
	wire _w1168_ ;
	wire _w1167_ ;
	wire _w1166_ ;
	wire _w1165_ ;
	wire _w1164_ ;
	wire _w1163_ ;
	wire _w1162_ ;
	wire _w1161_ ;
	wire _w1160_ ;
	wire _w1159_ ;
	wire _w1158_ ;
	wire _w1157_ ;
	wire _w1156_ ;
	wire _w1155_ ;
	wire _w1154_ ;
	wire _w1153_ ;
	wire _w1152_ ;
	wire _w1151_ ;
	wire _w1150_ ;
	wire _w1149_ ;
	wire _w1148_ ;
	wire _w1147_ ;
	wire _w1146_ ;
	wire _w1145_ ;
	wire _w1144_ ;
	wire _w1143_ ;
	wire _w1142_ ;
	wire _w1141_ ;
	wire _w1140_ ;
	wire _w1139_ ;
	wire _w1138_ ;
	wire _w1137_ ;
	wire _w1136_ ;
	wire _w1135_ ;
	wire _w1134_ ;
	wire _w1133_ ;
	wire _w1132_ ;
	wire _w1131_ ;
	wire _w1130_ ;
	wire _w1129_ ;
	wire _w1128_ ;
	wire _w1127_ ;
	wire _w1126_ ;
	wire _w1125_ ;
	wire _w1124_ ;
	wire _w1123_ ;
	wire _w1122_ ;
	wire _w1121_ ;
	wire _w1120_ ;
	wire _w1119_ ;
	wire _w1118_ ;
	wire _w1117_ ;
	wire _w1116_ ;
	wire _w1115_ ;
	wire _w1114_ ;
	wire _w1113_ ;
	wire _w1112_ ;
	wire _w1111_ ;
	wire _w1110_ ;
	wire _w1109_ ;
	wire _w1108_ ;
	wire _w1107_ ;
	wire _w1106_ ;
	wire _w1105_ ;
	wire _w1104_ ;
	wire _w1103_ ;
	wire _w1102_ ;
	wire _w1101_ ;
	wire _w1100_ ;
	wire _w1099_ ;
	wire _w1098_ ;
	wire _w1097_ ;
	wire _w1096_ ;
	wire _w1095_ ;
	wire _w1094_ ;
	wire _w1093_ ;
	wire _w1092_ ;
	wire _w1091_ ;
	wire _w1090_ ;
	wire _w1089_ ;
	wire _w1088_ ;
	wire _w1087_ ;
	wire _w1018_ ;
	wire _w1017_ ;
	wire _w1016_ ;
	wire _w1015_ ;
	wire _w1014_ ;
	wire _w1013_ ;
	wire _w1012_ ;
	wire _w1011_ ;
	wire _w1010_ ;
	wire _w1009_ ;
	wire _w1008_ ;
	wire _w1007_ ;
	wire _w1005_ ;
	wire _w1004_ ;
	wire _w1003_ ;
	wire _w1002_ ;
	wire _w1001_ ;
	wire _w1000_ ;
	wire _w999_ ;
	wire _w998_ ;
	wire _w997_ ;
	wire _w995_ ;
	wire _w994_ ;
	wire _w993_ ;
	wire _w996_ ;
	wire _w1848_ ;
	wire _w739_ ;
	wire _w3096_ ;
	wire _w1280_ ;
	wire _w992_ ;
	wire _w991_ ;
	wire _w990_ ;
	wire _w989_ ;
	wire _w972_ ;
	wire _w971_ ;
	wire _w970_ ;
	wire _w969_ ;
	wire _w968_ ;
	wire _w967_ ;
	wire _w966_ ;
	wire _w965_ ;
	wire _w1006_ ;
	wire _w1060_ ;
	wire _w964_ ;
	wire _w963_ ;
	wire _w962_ ;
	wire _w973_ ;
	wire _w974_ ;
	wire _w975_ ;
	wire _w976_ ;
	wire _w977_ ;
	wire _w978_ ;
	wire _w979_ ;
	wire _w980_ ;
	wire _w981_ ;
	wire _w982_ ;
	wire _w983_ ;
	wire _w984_ ;
	wire _w985_ ;
	wire _w986_ ;
	wire _w987_ ;
	wire _w988_ ;
	wire _w1019_ ;
	wire _w1020_ ;
	wire _w1021_ ;
	wire _w1022_ ;
	wire _w1023_ ;
	wire _w1024_ ;
	wire _w1025_ ;
	wire _w1026_ ;
	wire _w1027_ ;
	wire _w1028_ ;
	wire _w1029_ ;
	wire _w1030_ ;
	wire _w1031_ ;
	wire _w1032_ ;
	wire _w1033_ ;
	wire _w1034_ ;
	wire _w1035_ ;
	wire _w1036_ ;
	wire _w1037_ ;
	wire _w1038_ ;
	wire _w1039_ ;
	wire _w1040_ ;
	wire _w1041_ ;
	wire _w1042_ ;
	wire _w1043_ ;
	wire _w1044_ ;
	wire _w1045_ ;
	wire _w1046_ ;
	wire _w1047_ ;
	wire _w1048_ ;
	wire _w1049_ ;
	wire _w1050_ ;
	wire _w1051_ ;
	wire _w1052_ ;
	wire _w1053_ ;
	wire _w1054_ ;
	wire _w1055_ ;
	wire _w1056_ ;
	wire _w1057_ ;
	wire _w1058_ ;
	wire _w1059_ ;
	wire _w1061_ ;
	wire _w1062_ ;
	wire _w1063_ ;
	wire _w1064_ ;
	wire _w1065_ ;
	wire _w1066_ ;
	wire _w1067_ ;
	wire _w1068_ ;
	wire _w1380_ ;
	wire _w1069_ ;
	wire _w1070_ ;
	wire _w1071_ ;
	wire _w1072_ ;
	wire _w1073_ ;
	wire _w1074_ ;
	wire _w1075_ ;
	wire _w1076_ ;
	wire _w1077_ ;
	wire _w1078_ ;
	wire _w1079_ ;
	wire _w1080_ ;
	wire _w1081_ ;
	wire _w1082_ ;
	wire _w1083_ ;
	wire _w1084_ ;
	wire _w1085_ ;
	wire _w1086_ ;
	wire _w1217_ ;
	wire _w1218_ ;
	wire _w1219_ ;
	wire _w1220_ ;
	wire _w1221_ ;
	wire _w1222_ ;
	wire _w1223_ ;
	wire _w1224_ ;
	wire _w1225_ ;
	wire _w1226_ ;
	wire _w1227_ ;
	wire _w1228_ ;
	wire _w1229_ ;
	wire _w1230_ ;
	wire _w1231_ ;
	wire _w1232_ ;
	wire _w1233_ ;
	wire _w1234_ ;
	wire _w1235_ ;
	wire _w1236_ ;
	wire _w1237_ ;
	wire _w1238_ ;
	wire _w1239_ ;
	wire _w1240_ ;
	wire _w1241_ ;
	wire _w1242_ ;
	wire _w1243_ ;
	wire _w1244_ ;
	wire _w1245_ ;
	wire _w1246_ ;
	wire _w1247_ ;
	wire _w1248_ ;
	wire _w1249_ ;
	wire _w1250_ ;
	wire _w1251_ ;
	wire _w1252_ ;
	wire _w1253_ ;
	wire _w1254_ ;
	wire _w1255_ ;
	wire _w1256_ ;
	wire _w1257_ ;
	wire _w1258_ ;
	wire _w1259_ ;
	wire _w1260_ ;
	wire _w1261_ ;
	wire _w1262_ ;
	wire _w1263_ ;
	wire _w1264_ ;
	wire _w1265_ ;
	wire _w1266_ ;
	wire _w1267_ ;
	wire _w1268_ ;
	wire _w1269_ ;
	wire _w1270_ ;
	wire _w1271_ ;
	wire _w1272_ ;
	wire _w1273_ ;
	wire _w1274_ ;
	wire _w1275_ ;
	wire _w1276_ ;
	wire _w1277_ ;
	wire _w1278_ ;
	wire _w1279_ ;
	wire _w1281_ ;
	wire _w1282_ ;
	wire _w1283_ ;
	wire _w1284_ ;
	wire _w1285_ ;
	wire _w1286_ ;
	wire _w1287_ ;
	wire _w1288_ ;
	wire _w1289_ ;
	wire _w1290_ ;
	wire _w1291_ ;
	wire _w1292_ ;
	wire _w1293_ ;
	wire _w1294_ ;
	wire _w1295_ ;
	wire _w1296_ ;
	wire _w1297_ ;
	wire _w1298_ ;
	wire _w1299_ ;
	wire _w1300_ ;
	wire _w1301_ ;
	wire _w1302_ ;
	wire _w1303_ ;
	wire _w1304_ ;
	wire _w1305_ ;
	wire _w1306_ ;
	wire _w1307_ ;
	wire _w1308_ ;
	wire _w1309_ ;
	wire _w1310_ ;
	wire _w1311_ ;
	wire _w1312_ ;
	wire _w1313_ ;
	wire _w1314_ ;
	wire _w1315_ ;
	wire _w1316_ ;
	wire _w1317_ ;
	wire _w1318_ ;
	wire _w1319_ ;
	wire _w1320_ ;
	wire _w1321_ ;
	wire _w1322_ ;
	wire _w1323_ ;
	wire _w1324_ ;
	wire _w1325_ ;
	wire _w1326_ ;
	wire _w1327_ ;
	wire _w1328_ ;
	wire _w1329_ ;
	wire _w1330_ ;
	wire _w1331_ ;
	wire _w1332_ ;
	wire _w1333_ ;
	wire _w1334_ ;
	wire _w1335_ ;
	wire _w1336_ ;
	wire _w1337_ ;
	wire _w1338_ ;
	wire _w1339_ ;
	wire _w1340_ ;
	wire _w1341_ ;
	wire _w1342_ ;
	wire _w1343_ ;
	wire _w1344_ ;
	wire _w1345_ ;
	wire _w1346_ ;
	wire _w1347_ ;
	wire _w1348_ ;
	wire _w1349_ ;
	wire _w1350_ ;
	wire _w1351_ ;
	wire _w1352_ ;
	wire _w1353_ ;
	wire _w1354_ ;
	wire _w1355_ ;
	wire _w1356_ ;
	wire _w1357_ ;
	wire _w1358_ ;
	wire _w1359_ ;
	wire _w1360_ ;
	wire _w1361_ ;
	wire _w1362_ ;
	wire _w1363_ ;
	wire _w1364_ ;
	wire _w1365_ ;
	wire _w1366_ ;
	wire _w1367_ ;
	wire _w1368_ ;
	wire _w1369_ ;
	wire _w1370_ ;
	wire _w1371_ ;
	wire _w1372_ ;
	wire _w1373_ ;
	wire _w1374_ ;
	wire _w1375_ ;
	wire _w1376_ ;
	wire _w1377_ ;
	wire _w1378_ ;
	wire _w1379_ ;
	wire _w1381_ ;
	wire _w1382_ ;
	wire _w1383_ ;
	wire _w1384_ ;
	wire _w1385_ ;
	wire _w1386_ ;
	wire _w1387_ ;
	wire _w1388_ ;
	wire _w1389_ ;
	wire _w1390_ ;
	wire _w1391_ ;
	wire _w1392_ ;
	wire _w1393_ ;
	wire _w1394_ ;
	wire _w1395_ ;
	wire _w1396_ ;
	wire _w1397_ ;
	wire _w1398_ ;
	wire _w1399_ ;
	wire _w1400_ ;
	wire _w1401_ ;
	wire _w1402_ ;
	wire _w1403_ ;
	wire _w1404_ ;
	wire _w1405_ ;
	wire _w1406_ ;
	wire _w5385_ ;
	wire _w298_ ;
	wire _w2655_ ;
	wire _w1407_ ;
	wire _w1408_ ;
	wire _w1409_ ;
	wire _w1410_ ;
	wire _w1411_ ;
	wire _w1412_ ;
	wire _w1413_ ;
	wire _w1414_ ;
	wire _w1415_ ;
	wire _w1416_ ;
	wire _w1417_ ;
	wire _w1418_ ;
	wire _w1419_ ;
	wire _w1420_ ;
	wire _w1421_ ;
	wire _w1422_ ;
	wire _w1423_ ;
	wire _w1424_ ;
	wire _w1425_ ;
	wire _w1426_ ;
	wire _w1427_ ;
	wire _w1428_ ;
	wire _w1429_ ;
	wire _w1430_ ;
	wire _w1431_ ;
	wire _w1432_ ;
	wire _w1433_ ;
	wire _w1434_ ;
	wire _w1435_ ;
	wire _w1436_ ;
	wire _w1437_ ;
	wire _w1438_ ;
	wire _w1439_ ;
	wire _w1440_ ;
	wire _w1441_ ;
	wire _w1442_ ;
	wire _w1443_ ;
	wire _w1444_ ;
	wire _w1445_ ;
	wire _w1446_ ;
	wire _w1447_ ;
	wire _w1448_ ;
	wire _w1449_ ;
	wire _w1450_ ;
	wire _w1451_ ;
	wire _w1452_ ;
	wire _w1453_ ;
	wire _w1454_ ;
	wire _w1455_ ;
	wire _w1456_ ;
	wire _w1457_ ;
	wire _w1458_ ;
	wire _w1459_ ;
	wire _w1460_ ;
	wire _w1461_ ;
	wire _w1462_ ;
	wire _w1463_ ;
	wire _w1464_ ;
	wire _w1465_ ;
	wire _w1466_ ;
	wire _w1467_ ;
	wire _w1468_ ;
	wire _w1469_ ;
	wire _w1470_ ;
	wire _w1471_ ;
	wire _w1472_ ;
	wire _w1473_ ;
	wire _w1474_ ;
	wire _w1475_ ;
	wire _w1476_ ;
	wire _w1477_ ;
	wire _w1478_ ;
	wire _w1479_ ;
	wire _w1480_ ;
	wire _w1481_ ;
	wire _w1482_ ;
	wire _w1483_ ;
	wire _w1484_ ;
	wire _w1485_ ;
	wire _w1486_ ;
	wire _w1487_ ;
	wire _w1488_ ;
	wire _w1489_ ;
	wire _w1490_ ;
	wire _w1491_ ;
	wire _w1492_ ;
	wire _w1493_ ;
	wire _w1494_ ;
	wire _w1495_ ;
	wire _w1496_ ;
	wire _w1497_ ;
	wire _w1498_ ;
	wire _w1499_ ;
	wire _w1500_ ;
	wire _w2069_ ;
	wire _w2070_ ;
	wire _w2071_ ;
	wire _w2072_ ;
	wire _w2073_ ;
	wire _w2074_ ;
	wire _w2075_ ;
	wire _w2076_ ;
	wire _w2077_ ;
	wire _w2078_ ;
	wire _w2079_ ;
	wire _w2080_ ;
	wire _w2081_ ;
	wire _w2082_ ;
	wire _w2083_ ;
	wire _w2084_ ;
	wire _w2085_ ;
	wire _w2086_ ;
	wire _w2087_ ;
	wire _w2088_ ;
	wire _w2089_ ;
	wire _w2090_ ;
	wire _w2091_ ;
	wire _w2092_ ;
	wire _w2093_ ;
	wire _w2094_ ;
	wire _w2095_ ;
	wire _w2096_ ;
	wire _w2097_ ;
	wire _w2098_ ;
	wire _w2099_ ;
	wire _w2100_ ;
	wire _w2101_ ;
	wire _w2102_ ;
	wire _w2103_ ;
	wire _w2104_ ;
	wire _w2105_ ;
	wire _w2106_ ;
	wire _w2107_ ;
	wire _w2108_ ;
	wire _w2109_ ;
	wire _w2110_ ;
	wire _w2111_ ;
	wire _w2112_ ;
	wire _w2113_ ;
	wire _w2114_ ;
	wire _w2115_ ;
	wire _w2116_ ;
	wire _w2117_ ;
	wire _w2118_ ;
	wire _w2119_ ;
	wire _w2120_ ;
	wire _w2121_ ;
	wire _w2122_ ;
	wire _w2123_ ;
	wire _w2124_ ;
	wire _w2125_ ;
	wire _w2126_ ;
	wire _w2127_ ;
	wire _w2128_ ;
	wire _w2129_ ;
	wire _w2130_ ;
	wire _w2131_ ;
	wire _w2132_ ;
	wire _w2133_ ;
	wire _w2134_ ;
	wire _w2135_ ;
	wire _w2136_ ;
	wire _w2137_ ;
	wire _w2138_ ;
	wire _w2139_ ;
	wire _w2140_ ;
	wire _w2141_ ;
	wire _w2142_ ;
	wire _w2143_ ;
	wire _w2144_ ;
	wire _w2145_ ;
	wire _w2146_ ;
	wire _w2147_ ;
	wire _w2148_ ;
	wire _w2149_ ;
	wire _w2150_ ;
	wire _w2151_ ;
	wire _w2152_ ;
	wire _w2153_ ;
	wire _w2154_ ;
	wire _w2155_ ;
	wire _w2156_ ;
	wire _w2157_ ;
	wire _w2158_ ;
	wire _w2159_ ;
	wire _w2160_ ;
	wire _w2161_ ;
	wire _w2162_ ;
	wire _w2163_ ;
	wire _w2164_ ;
	wire _w2165_ ;
	wire _w2166_ ;
	wire _w2167_ ;
	wire _w2168_ ;
	wire _w2169_ ;
	wire _w2170_ ;
	wire _w2171_ ;
	wire _w2172_ ;
	wire _w2173_ ;
	wire _w2174_ ;
	wire _w2175_ ;
	wire _w2176_ ;
	wire _w2177_ ;
	wire _w2178_ ;
	wire _w2179_ ;
	wire _w2180_ ;
	wire _w2181_ ;
	wire _w2182_ ;
	wire _w2183_ ;
	wire _w2184_ ;
	wire _w2185_ ;
	wire _w2186_ ;
	wire _w2187_ ;
	wire _w2188_ ;
	wire _w2189_ ;
	wire _w2190_ ;
	wire _w2191_ ;
	wire _w2192_ ;
	wire _w2193_ ;
	wire _w2194_ ;
	wire _w2195_ ;
	wire _w2196_ ;
	wire _w2197_ ;
	wire _w2198_ ;
	wire _w2199_ ;
	wire _w2200_ ;
	wire _w2201_ ;
	wire _w2202_ ;
	wire _w2203_ ;
	wire _w2204_ ;
	wire _w2205_ ;
	wire _w2206_ ;
	wire _w2207_ ;
	wire _w2208_ ;
	wire _w2209_ ;
	wire _w2210_ ;
	wire _w2211_ ;
	wire _w2212_ ;
	wire _w2213_ ;
	wire _w2214_ ;
	wire _w2215_ ;
	wire _w2216_ ;
	wire _w2217_ ;
	wire _w2218_ ;
	wire _w2219_ ;
	wire _w2220_ ;
	wire _w2221_ ;
	wire _w2222_ ;
	wire _w2223_ ;
	wire _w2224_ ;
	wire _w2225_ ;
	wire _w2226_ ;
	wire _w2227_ ;
	wire _w2228_ ;
	wire _w2229_ ;
	wire _w2230_ ;
	wire _w2231_ ;
	wire _w2232_ ;
	wire _w2233_ ;
	wire _w2234_ ;
	wire _w2235_ ;
	wire _w2236_ ;
	wire _w2237_ ;
	wire _w2238_ ;
	wire _w2239_ ;
	wire _w2240_ ;
	wire _w2241_ ;
	wire _w2242_ ;
	wire _w2243_ ;
	wire _w2244_ ;
	wire _w2245_ ;
	wire _w2246_ ;
	wire _w2247_ ;
	wire _w2248_ ;
	wire _w2249_ ;
	wire _w2250_ ;
	wire _w2251_ ;
	wire _w2252_ ;
	wire _w2253_ ;
	wire _w2254_ ;
	wire _w2255_ ;
	wire _w2256_ ;
	wire _w2257_ ;
	wire _w2258_ ;
	wire _w2259_ ;
	wire _w2260_ ;
	wire _w2261_ ;
	wire _w2262_ ;
	wire _w2263_ ;
	wire _w2264_ ;
	wire _w2265_ ;
	wire _w2266_ ;
	wire _w2267_ ;
	wire _w2268_ ;
	wire _w2269_ ;
	wire _w2270_ ;
	wire _w2271_ ;
	wire _w2272_ ;
	wire _w2273_ ;
	wire _w2274_ ;
	wire _w2275_ ;
	wire _w2276_ ;
	wire _w2277_ ;
	wire _w2278_ ;
	wire _w2279_ ;
	wire _w2280_ ;
	wire _w2281_ ;
	wire _w2282_ ;
	wire _w2283_ ;
	wire _w2284_ ;
	wire _w2285_ ;
	wire _w2286_ ;
	wire _w2287_ ;
	wire _w2288_ ;
	wire _w2289_ ;
	wire _w2290_ ;
	wire _w2291_ ;
	wire _w2292_ ;
	wire _w2293_ ;
	wire _w2294_ ;
	wire _w2295_ ;
	wire _w2296_ ;
	wire _w2297_ ;
	wire _w2298_ ;
	wire _w2299_ ;
	wire _w2300_ ;
	wire _w2301_ ;
	wire _w2302_ ;
	wire _w2303_ ;
	wire _w2304_ ;
	wire _w2305_ ;
	wire _w2306_ ;
	wire _w2307_ ;
	wire _w2308_ ;
	wire _w2309_ ;
	wire _w2310_ ;
	wire _w2311_ ;
	wire _w2312_ ;
	wire _w2313_ ;
	wire _w2314_ ;
	wire _w2315_ ;
	wire _w2316_ ;
	wire _w2317_ ;
	wire _w2318_ ;
	wire _w2319_ ;
	wire _w2320_ ;
	wire _w2321_ ;
	wire _w2322_ ;
	wire _w2323_ ;
	wire _w2324_ ;
	wire _w2325_ ;
	wire _w2326_ ;
	wire _w2327_ ;
	wire _w2328_ ;
	wire _w2329_ ;
	wire _w2330_ ;
	wire _w2331_ ;
	wire _w2332_ ;
	wire _w2333_ ;
	wire _w2334_ ;
	wire _w2335_ ;
	wire _w2336_ ;
	wire _w2337_ ;
	wire _w2338_ ;
	wire _w2339_ ;
	wire _w2340_ ;
	wire _w2341_ ;
	wire _w2342_ ;
	wire _w2343_ ;
	wire _w2344_ ;
	wire _w2345_ ;
	wire _w2346_ ;
	wire _w2347_ ;
	wire _w2348_ ;
	wire _w2349_ ;
	wire _w2350_ ;
	wire _w2351_ ;
	wire _w2352_ ;
	wire _w2353_ ;
	wire _w2354_ ;
	wire _w2355_ ;
	wire _w2356_ ;
	wire _w2357_ ;
	wire _w2358_ ;
	wire _w2359_ ;
	wire _w2360_ ;
	wire _w2361_ ;
	wire _w2362_ ;
	wire _w2363_ ;
	wire _w2364_ ;
	wire _w2365_ ;
	wire _w2366_ ;
	wire _w2367_ ;
	wire _w2368_ ;
	wire _w2369_ ;
	wire _w2370_ ;
	wire _w2371_ ;
	wire _w2372_ ;
	wire _w2373_ ;
	wire _w2374_ ;
	wire _w2375_ ;
	wire _w2376_ ;
	wire _w2377_ ;
	wire _w2378_ ;
	wire _w2379_ ;
	wire _w2380_ ;
	wire _w2381_ ;
	wire _w2382_ ;
	wire _w2383_ ;
	wire _w2384_ ;
	wire _w2385_ ;
	wire _w2386_ ;
	wire _w2387_ ;
	wire _w2388_ ;
	wire _w2389_ ;
	wire _w2390_ ;
	wire _w2391_ ;
	wire _w2392_ ;
	wire _w2393_ ;
	wire _w2394_ ;
	wire _w2395_ ;
	wire _w2396_ ;
	wire _w2397_ ;
	wire _w2398_ ;
	wire _w2399_ ;
	wire _w2400_ ;
	wire _w2401_ ;
	wire _w2402_ ;
	wire _w2403_ ;
	wire _w2404_ ;
	wire _w2405_ ;
	wire _w2406_ ;
	wire _w2407_ ;
	wire _w2408_ ;
	wire _w2409_ ;
	wire _w2410_ ;
	wire _w2411_ ;
	wire _w2412_ ;
	wire _w2413_ ;
	wire _w2414_ ;
	wire _w2415_ ;
	wire _w2416_ ;
	wire _w2417_ ;
	wire _w2418_ ;
	wire _w2419_ ;
	wire _w2420_ ;
	wire _w2421_ ;
	wire _w2422_ ;
	wire _w2423_ ;
	wire _w2424_ ;
	wire _w2425_ ;
	wire _w2426_ ;
	wire _w2427_ ;
	wire _w2428_ ;
	wire _w2429_ ;
	wire _w2430_ ;
	wire _w2431_ ;
	wire _w2432_ ;
	wire _w2433_ ;
	wire _w2434_ ;
	wire _w2435_ ;
	wire _w2436_ ;
	wire _w2437_ ;
	wire _w2438_ ;
	wire _w2439_ ;
	wire _w2440_ ;
	wire _w2441_ ;
	wire _w2442_ ;
	wire _w2443_ ;
	wire _w2444_ ;
	wire _w2445_ ;
	wire _w2446_ ;
	wire _w2447_ ;
	wire _w2448_ ;
	wire _w2449_ ;
	wire _w2450_ ;
	wire _w2451_ ;
	wire _w2452_ ;
	wire _w2453_ ;
	wire _w2454_ ;
	wire _w2455_ ;
	wire _w2456_ ;
	wire _w2457_ ;
	wire _w2458_ ;
	wire _w2459_ ;
	wire _w2460_ ;
	wire _w2461_ ;
	wire _w2462_ ;
	wire _w2463_ ;
	wire _w2464_ ;
	wire _w2465_ ;
	wire _w2466_ ;
	wire _w2467_ ;
	wire _w2468_ ;
	wire _w2469_ ;
	wire _w2470_ ;
	wire _w2471_ ;
	wire _w2472_ ;
	wire _w2473_ ;
	wire _w2474_ ;
	wire _w2475_ ;
	wire _w2476_ ;
	wire _w2477_ ;
	wire _w2478_ ;
	wire _w2479_ ;
	wire _w2480_ ;
	wire _w2481_ ;
	wire _w2482_ ;
	wire _w2483_ ;
	wire _w2484_ ;
	wire _w2485_ ;
	wire _w2486_ ;
	wire _w2487_ ;
	wire _w2488_ ;
	wire _w2489_ ;
	wire _w2490_ ;
	wire _w2491_ ;
	wire _w2492_ ;
	wire _w2493_ ;
	wire _w2494_ ;
	wire _w2495_ ;
	wire _w2496_ ;
	wire _w2497_ ;
	wire _w2498_ ;
	wire _w2499_ ;
	wire _w2500_ ;
	wire _w2501_ ;
	wire _w2502_ ;
	wire _w2503_ ;
	wire _w2504_ ;
	wire _w2505_ ;
	wire _w2506_ ;
	wire _w2507_ ;
	wire _w2508_ ;
	wire _w2509_ ;
	wire _w2510_ ;
	wire _w2511_ ;
	wire _w2512_ ;
	wire _w2513_ ;
	wire _w2514_ ;
	wire _w2515_ ;
	wire _w2516_ ;
	wire _w2517_ ;
	wire _w2518_ ;
	wire _w2519_ ;
	wire _w2520_ ;
	wire _w2521_ ;
	wire _w2522_ ;
	wire _w2523_ ;
	wire _w2524_ ;
	wire _w2525_ ;
	wire _w2526_ ;
	wire _w2527_ ;
	wire _w2528_ ;
	wire _w2529_ ;
	wire _w2530_ ;
	wire _w2531_ ;
	wire _w2532_ ;
	wire _w2533_ ;
	wire _w2534_ ;
	wire _w2535_ ;
	wire _w2536_ ;
	wire _w2537_ ;
	wire _w2538_ ;
	wire _w2539_ ;
	wire _w2540_ ;
	wire _w2541_ ;
	wire _w2542_ ;
	wire _w2543_ ;
	wire _w2544_ ;
	wire _w2545_ ;
	wire _w2546_ ;
	wire _w2547_ ;
	wire _w2548_ ;
	wire _w2549_ ;
	wire _w2550_ ;
	wire _w2551_ ;
	wire _w2552_ ;
	wire _w2553_ ;
	wire _w2554_ ;
	wire _w2555_ ;
	wire _w2556_ ;
	wire _w2557_ ;
	wire _w2558_ ;
	wire _w2559_ ;
	wire _w2560_ ;
	wire _w2561_ ;
	wire _w2562_ ;
	wire _w2563_ ;
	wire _w2564_ ;
	wire _w2565_ ;
	wire _w2566_ ;
	wire _w2567_ ;
	wire _w2568_ ;
	wire _w2569_ ;
	wire _w2570_ ;
	wire _w2571_ ;
	wire _w2572_ ;
	wire _w2573_ ;
	wire _w2574_ ;
	wire _w2575_ ;
	wire _w2576_ ;
	wire _w2577_ ;
	wire _w2578_ ;
	wire _w2579_ ;
	wire _w2580_ ;
	wire _w2581_ ;
	wire _w2582_ ;
	wire _w2583_ ;
	wire _w2584_ ;
	wire _w2585_ ;
	wire _w2586_ ;
	wire _w2587_ ;
	wire _w2588_ ;
	wire _w2589_ ;
	wire _w2590_ ;
	wire _w2591_ ;
	wire _w2592_ ;
	wire _w2593_ ;
	wire _w2594_ ;
	wire _w2595_ ;
	wire _w2596_ ;
	wire _w2597_ ;
	wire _w2598_ ;
	wire _w2599_ ;
	wire _w2600_ ;
	wire _w2601_ ;
	wire _w2602_ ;
	wire _w2603_ ;
	wire _w2604_ ;
	wire _w2605_ ;
	wire _w2606_ ;
	wire _w2607_ ;
	wire _w2608_ ;
	wire _w2609_ ;
	wire _w2610_ ;
	wire _w2611_ ;
	wire _w2612_ ;
	wire _w2613_ ;
	wire _w2614_ ;
	wire _w2615_ ;
	wire _w2616_ ;
	wire _w2617_ ;
	wire _w2618_ ;
	wire _w2619_ ;
	wire _w2620_ ;
	wire _w2621_ ;
	wire _w2622_ ;
	wire _w2623_ ;
	wire _w2624_ ;
	wire _w2625_ ;
	wire _w2626_ ;
	wire _w2627_ ;
	wire _w2628_ ;
	wire _w2629_ ;
	wire _w2630_ ;
	wire _w2631_ ;
	wire _w2632_ ;
	wire _w2633_ ;
	wire _w2634_ ;
	wire _w2635_ ;
	wire _w2636_ ;
	wire _w2637_ ;
	wire _w2638_ ;
	wire _w2639_ ;
	wire _w2640_ ;
	wire _w2641_ ;
	wire _w2642_ ;
	wire _w2643_ ;
	wire _w2644_ ;
	wire _w2645_ ;
	wire _w2646_ ;
	wire _w2647_ ;
	wire _w2648_ ;
	wire _w2649_ ;
	wire _w2650_ ;
	wire _w2651_ ;
	wire _w2652_ ;
	wire _w2653_ ;
	wire _w2654_ ;
	wire _w2656_ ;
	wire _w2657_ ;
	wire _w2658_ ;
	wire _w2659_ ;
	wire _w2660_ ;
	wire _w2661_ ;
	wire _w2662_ ;
	wire _w2663_ ;
	wire _w2664_ ;
	wire _w2665_ ;
	wire _w2666_ ;
	wire _w2667_ ;
	wire _w2668_ ;
	wire _w2669_ ;
	wire _w2670_ ;
	wire _w2671_ ;
	wire _w2672_ ;
	wire _w2673_ ;
	wire _w2674_ ;
	wire _w2675_ ;
	wire _w2676_ ;
	wire _w2677_ ;
	wire _w2678_ ;
	wire _w2679_ ;
	wire _w2680_ ;
	wire _w2681_ ;
	wire _w2682_ ;
	wire _w2683_ ;
	wire _w2684_ ;
	wire _w2685_ ;
	wire _w2686_ ;
	wire _w2687_ ;
	wire _w2688_ ;
	wire _w2689_ ;
	wire _w2690_ ;
	wire _w2691_ ;
	wire _w2692_ ;
	wire _w2693_ ;
	wire _w2694_ ;
	wire _w2695_ ;
	wire _w2696_ ;
	wire _w2697_ ;
	wire _w2698_ ;
	wire _w2699_ ;
	wire _w2700_ ;
	wire _w2701_ ;
	wire _w2702_ ;
	wire _w2703_ ;
	wire _w2704_ ;
	wire _w2705_ ;
	wire _w2706_ ;
	wire _w2707_ ;
	wire _w2708_ ;
	wire _w2709_ ;
	wire _w2710_ ;
	wire _w2711_ ;
	wire _w2712_ ;
	wire _w2713_ ;
	wire _w2714_ ;
	wire _w2715_ ;
	wire _w2716_ ;
	wire _w2717_ ;
	wire _w2718_ ;
	wire _w2719_ ;
	wire _w2720_ ;
	wire _w2721_ ;
	wire _w2722_ ;
	wire _w2723_ ;
	wire _w2724_ ;
	wire _w2725_ ;
	wire _w2726_ ;
	wire _w2727_ ;
	wire _w2728_ ;
	wire _w2729_ ;
	wire _w2730_ ;
	wire _w2731_ ;
	wire _w2732_ ;
	wire _w2733_ ;
	wire _w2734_ ;
	wire _w2735_ ;
	wire _w2736_ ;
	wire _w2737_ ;
	wire _w2738_ ;
	wire _w2739_ ;
	wire _w2740_ ;
	wire _w2741_ ;
	wire _w2742_ ;
	wire _w2743_ ;
	wire _w2744_ ;
	wire _w2745_ ;
	wire _w2746_ ;
	wire _w2747_ ;
	wire _w2748_ ;
	wire _w2749_ ;
	wire _w2750_ ;
	wire _w2751_ ;
	wire _w2752_ ;
	wire _w2753_ ;
	wire _w2754_ ;
	wire _w2755_ ;
	wire _w2756_ ;
	wire _w2757_ ;
	wire _w2758_ ;
	wire _w2759_ ;
	wire _w2760_ ;
	wire _w2761_ ;
	wire _w2762_ ;
	wire _w2763_ ;
	wire _w2764_ ;
	wire _w2765_ ;
	wire _w2766_ ;
	wire _w2767_ ;
	wire _w2768_ ;
	wire _w2769_ ;
	wire _w2770_ ;
	wire _w2771_ ;
	wire _w2772_ ;
	wire _w2773_ ;
	wire _w2774_ ;
	wire _w2775_ ;
	wire _w2776_ ;
	wire _w2777_ ;
	wire _w2778_ ;
	wire _w2779_ ;
	wire _w2780_ ;
	wire _w2781_ ;
	wire _w2782_ ;
	wire _w2783_ ;
	wire _w2784_ ;
	wire _w2785_ ;
	wire _w2786_ ;
	wire _w2787_ ;
	wire _w2788_ ;
	wire _w2789_ ;
	wire _w2790_ ;
	wire _w2791_ ;
	wire _w2792_ ;
	wire _w2793_ ;
	wire _w2794_ ;
	wire _w2795_ ;
	wire _w2796_ ;
	wire _w2797_ ;
	wire _w2798_ ;
	wire _w2799_ ;
	wire _w2800_ ;
	wire _w2801_ ;
	wire _w2802_ ;
	wire _w2803_ ;
	wire _w2804_ ;
	wire _w2805_ ;
	wire _w2806_ ;
	wire _w2807_ ;
	wire _w2808_ ;
	wire _w2809_ ;
	wire _w2810_ ;
	wire _w2811_ ;
	wire _w2812_ ;
	wire _w2813_ ;
	wire _w2814_ ;
	wire _w2815_ ;
	wire _w2816_ ;
	wire _w2817_ ;
	wire _w2818_ ;
	wire _w2819_ ;
	wire _w2820_ ;
	wire _w2821_ ;
	wire _w2822_ ;
	wire _w2823_ ;
	wire _w2824_ ;
	wire _w2825_ ;
	wire _w2826_ ;
	wire _w2827_ ;
	wire _w2828_ ;
	wire _w2829_ ;
	wire _w2830_ ;
	wire _w2831_ ;
	wire _w2832_ ;
	wire _w2833_ ;
	wire _w2834_ ;
	wire _w2835_ ;
	wire _w2836_ ;
	wire _w2837_ ;
	wire _w2838_ ;
	wire _w2839_ ;
	wire _w2840_ ;
	wire _w2841_ ;
	wire _w2842_ ;
	wire _w2843_ ;
	wire _w2844_ ;
	wire _w2845_ ;
	wire _w2846_ ;
	wire _w2847_ ;
	wire _w2848_ ;
	wire _w2849_ ;
	wire _w2850_ ;
	wire _w2851_ ;
	wire _w2852_ ;
	wire _w2853_ ;
	wire _w2854_ ;
	wire _w2855_ ;
	wire _w2856_ ;
	wire _w2857_ ;
	wire _w2858_ ;
	wire _w2859_ ;
	wire _w2860_ ;
	wire _w2861_ ;
	wire _w2862_ ;
	wire _w2863_ ;
	wire _w2864_ ;
	wire _w2865_ ;
	wire _w2866_ ;
	wire _w2867_ ;
	wire _w2868_ ;
	wire _w2869_ ;
	wire _w2870_ ;
	wire _w2871_ ;
	wire _w2872_ ;
	wire _w2873_ ;
	wire _w2874_ ;
	wire _w2875_ ;
	wire _w2876_ ;
	wire _w2877_ ;
	wire _w2878_ ;
	wire _w2879_ ;
	wire _w2880_ ;
	wire _w2881_ ;
	wire _w2882_ ;
	wire _w2883_ ;
	wire _w2884_ ;
	wire _w2885_ ;
	wire _w2886_ ;
	wire _w2887_ ;
	wire _w2888_ ;
	wire _w2889_ ;
	wire _w2890_ ;
	wire _w2891_ ;
	wire _w2892_ ;
	wire _w2893_ ;
	wire _w2894_ ;
	wire _w2895_ ;
	wire _w2896_ ;
	wire _w2897_ ;
	wire _w2898_ ;
	wire _w2899_ ;
	wire _w2900_ ;
	wire _w2901_ ;
	wire _w2902_ ;
	wire _w2903_ ;
	wire _w2904_ ;
	wire _w2905_ ;
	wire _w2906_ ;
	wire _w2907_ ;
	wire _w2908_ ;
	wire _w2909_ ;
	wire _w2910_ ;
	wire _w2911_ ;
	wire _w2912_ ;
	wire _w2913_ ;
	wire _w2914_ ;
	wire _w2915_ ;
	wire _w2916_ ;
	wire _w2917_ ;
	wire _w2918_ ;
	wire _w2919_ ;
	wire _w2920_ ;
	wire _w2921_ ;
	wire _w2922_ ;
	wire _w2923_ ;
	wire _w2924_ ;
	wire _w2925_ ;
	wire _w2926_ ;
	wire _w2927_ ;
	wire _w2928_ ;
	wire _w2929_ ;
	wire _w2930_ ;
	wire _w2931_ ;
	wire _w2932_ ;
	wire _w2933_ ;
	wire _w2934_ ;
	wire _w2935_ ;
	wire _w2936_ ;
	wire _w2937_ ;
	wire _w2938_ ;
	wire _w2939_ ;
	wire _w2940_ ;
	wire _w2941_ ;
	wire _w2942_ ;
	wire _w2943_ ;
	wire _w2944_ ;
	wire _w2945_ ;
	wire _w2946_ ;
	wire _w2947_ ;
	wire _w2948_ ;
	wire _w2949_ ;
	wire _w2950_ ;
	wire _w2951_ ;
	wire _w2952_ ;
	wire _w2953_ ;
	wire _w2954_ ;
	wire _w2955_ ;
	wire _w2956_ ;
	wire _w2957_ ;
	wire _w2958_ ;
	wire _w2959_ ;
	wire _w2960_ ;
	wire _w2961_ ;
	wire _w2962_ ;
	wire _w2963_ ;
	wire _w2964_ ;
	wire _w2965_ ;
	wire _w2966_ ;
	wire _w2967_ ;
	wire _w2968_ ;
	wire _w2969_ ;
	wire _w2970_ ;
	wire _w2971_ ;
	wire _w2972_ ;
	wire _w2973_ ;
	wire _w2974_ ;
	wire _w2975_ ;
	wire _w2976_ ;
	wire _w2977_ ;
	wire _w2978_ ;
	wire _w2979_ ;
	wire _w2980_ ;
	wire _w2981_ ;
	wire _w2982_ ;
	wire _w2983_ ;
	wire _w2984_ ;
	wire _w2985_ ;
	wire _w2986_ ;
	wire _w2987_ ;
	wire _w2988_ ;
	wire _w2989_ ;
	wire _w2990_ ;
	wire _w2991_ ;
	wire _w2992_ ;
	wire _w2993_ ;
	wire _w2994_ ;
	wire _w2995_ ;
	wire _w2996_ ;
	wire _w2997_ ;
	wire _w2998_ ;
	wire _w2999_ ;
	wire _w3000_ ;
	wire _w3001_ ;
	wire _w3002_ ;
	wire _w3003_ ;
	wire _w3004_ ;
	wire _w3005_ ;
	wire _w3006_ ;
	wire _w3007_ ;
	wire _w3008_ ;
	wire _w3009_ ;
	wire _w3010_ ;
	wire _w3011_ ;
	wire _w3012_ ;
	wire _w3013_ ;
	wire _w3014_ ;
	wire _w3015_ ;
	wire _w3016_ ;
	wire _w3017_ ;
	wire _w3018_ ;
	wire _w3019_ ;
	wire _w3020_ ;
	wire _w3021_ ;
	wire _w3022_ ;
	wire _w3023_ ;
	wire _w3024_ ;
	wire _w3025_ ;
	wire _w3026_ ;
	wire _w3027_ ;
	wire _w3028_ ;
	wire _w3029_ ;
	wire _w3030_ ;
	wire _w3031_ ;
	wire _w3032_ ;
	wire _w3033_ ;
	wire _w3034_ ;
	wire _w3035_ ;
	wire _w3036_ ;
	wire _w3037_ ;
	wire _w3038_ ;
	wire _w3039_ ;
	wire _w3040_ ;
	wire _w3041_ ;
	wire _w3042_ ;
	wire _w3043_ ;
	wire _w3044_ ;
	wire _w3045_ ;
	wire _w3046_ ;
	wire _w3047_ ;
	wire _w3048_ ;
	wire _w3049_ ;
	wire _w3050_ ;
	wire _w3051_ ;
	wire _w3052_ ;
	wire _w3053_ ;
	wire _w3054_ ;
	wire _w3055_ ;
	wire _w3056_ ;
	wire _w3057_ ;
	wire _w3058_ ;
	wire _w3059_ ;
	wire _w3060_ ;
	wire _w3061_ ;
	wire _w3062_ ;
	wire _w3063_ ;
	wire _w3064_ ;
	wire _w3065_ ;
	wire _w3066_ ;
	wire _w3067_ ;
	wire _w3068_ ;
	wire _w3069_ ;
	wire _w3070_ ;
	wire _w3071_ ;
	wire _w3072_ ;
	wire _w3073_ ;
	wire _w3074_ ;
	wire _w3075_ ;
	wire _w3076_ ;
	wire _w3077_ ;
	wire _w3078_ ;
	wire _w3079_ ;
	wire _w3080_ ;
	wire _w3081_ ;
	wire _w3082_ ;
	wire _w3083_ ;
	wire _w3084_ ;
	wire _w3085_ ;
	wire _w3086_ ;
	wire _w3087_ ;
	wire _w3088_ ;
	wire _w3089_ ;
	wire _w3090_ ;
	wire _w3091_ ;
	wire _w3092_ ;
	wire _w3093_ ;
	wire _w3094_ ;
	wire _w3095_ ;
	wire _w3097_ ;
	wire _w3098_ ;
	wire _w3099_ ;
	wire _w3100_ ;
	wire _w3101_ ;
	wire _w3102_ ;
	wire _w3103_ ;
	wire _w3104_ ;
	wire _w3105_ ;
	wire _w3106_ ;
	wire _w3107_ ;
	wire _w3108_ ;
	wire _w3109_ ;
	wire _w3110_ ;
	wire _w3111_ ;
	wire _w3112_ ;
	wire _w3113_ ;
	wire _w3114_ ;
	wire _w3115_ ;
	wire _w3116_ ;
	wire _w3117_ ;
	wire _w3118_ ;
	wire _w3119_ ;
	wire _w3120_ ;
	wire _w3121_ ;
	wire _w3122_ ;
	wire _w3123_ ;
	wire _w3124_ ;
	wire _w3125_ ;
	wire _w3126_ ;
	wire _w3127_ ;
	wire _w3128_ ;
	wire _w3129_ ;
	wire _w3130_ ;
	wire _w3131_ ;
	wire _w3132_ ;
	wire _w3133_ ;
	wire _w3134_ ;
	wire _w3135_ ;
	wire _w3136_ ;
	wire _w3137_ ;
	wire _w3138_ ;
	wire _w3139_ ;
	wire _w3140_ ;
	wire _w3141_ ;
	wire _w3142_ ;
	wire _w3143_ ;
	wire _w3144_ ;
	wire _w3145_ ;
	wire _w3146_ ;
	wire _w3147_ ;
	wire _w3148_ ;
	wire _w3149_ ;
	wire _w3150_ ;
	wire _w3151_ ;
	wire _w3152_ ;
	wire _w3153_ ;
	wire _w3154_ ;
	wire _w3155_ ;
	wire _w3156_ ;
	wire _w3157_ ;
	wire _w3158_ ;
	wire _w3159_ ;
	wire _w3160_ ;
	wire _w3161_ ;
	wire _w3162_ ;
	wire _w3163_ ;
	wire _w3164_ ;
	wire _w3165_ ;
	wire _w3166_ ;
	wire _w3167_ ;
	wire _w3168_ ;
	wire _w3169_ ;
	wire _w3170_ ;
	wire _w3171_ ;
	wire _w3172_ ;
	wire _w3173_ ;
	wire _w3174_ ;
	wire _w3175_ ;
	wire _w3176_ ;
	wire _w3177_ ;
	wire _w3178_ ;
	wire _w3179_ ;
	wire _w3180_ ;
	wire _w3181_ ;
	wire _w3182_ ;
	wire _w3183_ ;
	wire _w3184_ ;
	wire _w3185_ ;
	wire _w3186_ ;
	wire _w3187_ ;
	wire _w3188_ ;
	wire _w3189_ ;
	wire _w3190_ ;
	wire _w3191_ ;
	wire _w3192_ ;
	wire _w3193_ ;
	wire _w3194_ ;
	wire _w3195_ ;
	wire _w3196_ ;
	wire _w3197_ ;
	wire _w3198_ ;
	wire _w3199_ ;
	wire _w3200_ ;
	wire _w3201_ ;
	wire _w3202_ ;
	wire _w3203_ ;
	wire _w3204_ ;
	wire _w3205_ ;
	wire _w3206_ ;
	wire _w3207_ ;
	wire _w3208_ ;
	wire _w3209_ ;
	wire _w3210_ ;
	wire _w3211_ ;
	wire _w3212_ ;
	wire _w3213_ ;
	wire _w3214_ ;
	wire _w3215_ ;
	wire _w3216_ ;
	wire _w3217_ ;
	wire _w3218_ ;
	wire _w3219_ ;
	wire _w3220_ ;
	wire _w3221_ ;
	wire _w3222_ ;
	wire _w3223_ ;
	wire _w3224_ ;
	wire _w3225_ ;
	wire _w3226_ ;
	wire _w3227_ ;
	wire _w3228_ ;
	wire _w3229_ ;
	wire _w3230_ ;
	wire _w3231_ ;
	wire _w3232_ ;
	wire _w3233_ ;
	wire _w3234_ ;
	wire _w3235_ ;
	wire _w3236_ ;
	wire _w3237_ ;
	wire _w3238_ ;
	wire _w3239_ ;
	wire _w3240_ ;
	wire _w3241_ ;
	wire _w3242_ ;
	wire _w3243_ ;
	wire _w3244_ ;
	wire _w3245_ ;
	wire _w3246_ ;
	wire _w3247_ ;
	wire _w3248_ ;
	wire _w3249_ ;
	wire _w3250_ ;
	wire _w3251_ ;
	wire _w3252_ ;
	wire _w3253_ ;
	wire _w3254_ ;
	wire _w3255_ ;
	wire _w3256_ ;
	wire _w3257_ ;
	wire _w3258_ ;
	wire _w3259_ ;
	wire _w3260_ ;
	wire _w3261_ ;
	wire _w3262_ ;
	wire _w3263_ ;
	wire _w3264_ ;
	wire _w3265_ ;
	wire _w3266_ ;
	wire _w3267_ ;
	wire _w3268_ ;
	wire _w3269_ ;
	wire _w3270_ ;
	wire _w3271_ ;
	wire _w3272_ ;
	wire _w3273_ ;
	wire _w3274_ ;
	wire _w3275_ ;
	wire _w3276_ ;
	wire _w3277_ ;
	wire _w3278_ ;
	wire _w3279_ ;
	wire _w3280_ ;
	wire _w3281_ ;
	wire _w3282_ ;
	wire _w3283_ ;
	wire _w3284_ ;
	wire _w3285_ ;
	wire _w3286_ ;
	wire _w3287_ ;
	wire _w3288_ ;
	wire _w3289_ ;
	wire _w3290_ ;
	wire _w3291_ ;
	wire _w3292_ ;
	wire _w3293_ ;
	wire _w3294_ ;
	wire _w3295_ ;
	wire _w3296_ ;
	wire _w3297_ ;
	wire _w3298_ ;
	wire _w3299_ ;
	wire _w3300_ ;
	wire _w3301_ ;
	wire _w3302_ ;
	wire _w3303_ ;
	wire _w3304_ ;
	wire _w3305_ ;
	wire _w3306_ ;
	wire _w3307_ ;
	wire _w3308_ ;
	wire _w3309_ ;
	wire _w3310_ ;
	wire _w3311_ ;
	wire _w3312_ ;
	wire _w3313_ ;
	wire _w3314_ ;
	wire _w3315_ ;
	wire _w3316_ ;
	LUT1 #(
		.INIT('h1)
	) name0 (
		\u1_acs_addr_reg[0]/P0001 ,
		_w298_
	);
	LUT1 #(
		.INIT('h1)
	) name1 (
		\u5_mc_le_reg/NET0131 ,
		_w739_
	);
	LUT2 #(
		.INIT('h1)
	) name2 (
		\u5_state_reg[40]/NET0131 ,
		\u5_state_reg[41]/NET0131 ,
		_w962_
	);
	LUT4 #(
		.INIT('h0001)
	) name3 (
		\u5_state_reg[38]/NET0131 ,
		\u5_state_reg[39]/NET0131 ,
		\u5_state_reg[40]/NET0131 ,
		\u5_state_reg[41]/NET0131 ,
		_w963_
	);
	LUT2 #(
		.INIT('h1)
	) name4 (
		\u5_state_reg[42]/NET0131 ,
		\u5_state_reg[44]/NET0131 ,
		_w964_
	);
	LUT4 #(
		.INIT('h0001)
	) name5 (
		\u5_state_reg[42]/NET0131 ,
		\u5_state_reg[43]/NET0131 ,
		\u5_state_reg[44]/NET0131 ,
		\u5_state_reg[45]/NET0131 ,
		_w965_
	);
	LUT2 #(
		.INIT('h8)
	) name6 (
		_w963_,
		_w965_,
		_w966_
	);
	LUT2 #(
		.INIT('h1)
	) name7 (
		\u5_state_reg[36]/NET0131 ,
		\u5_state_reg[37]/NET0131 ,
		_w967_
	);
	LUT4 #(
		.INIT('h0001)
	) name8 (
		\u5_state_reg[34]/NET0131 ,
		\u5_state_reg[35]/NET0131 ,
		\u5_state_reg[36]/NET0131 ,
		\u5_state_reg[37]/NET0131 ,
		_w968_
	);
	LUT2 #(
		.INIT('h1)
	) name9 (
		\u5_state_reg[46]/NET0131 ,
		\u5_state_reg[49]/NET0131 ,
		_w969_
	);
	LUT4 #(
		.INIT('h0001)
	) name10 (
		\u5_state_reg[46]/NET0131 ,
		\u5_state_reg[47]/NET0131 ,
		\u5_state_reg[48]/NET0131 ,
		\u5_state_reg[49]/NET0131 ,
		_w970_
	);
	LUT4 #(
		.INIT('h8000)
	) name11 (
		_w963_,
		_w965_,
		_w968_,
		_w970_,
		_w971_
	);
	LUT2 #(
		.INIT('h1)
	) name12 (
		\u5_state_reg[28]/NET0131 ,
		\u5_state_reg[29]/NET0131 ,
		_w972_
	);
	LUT4 #(
		.INIT('h0001)
	) name13 (
		\u5_state_reg[26]/NET0131 ,
		\u5_state_reg[27]/NET0131 ,
		\u5_state_reg[28]/NET0131 ,
		\u5_state_reg[29]/NET0131 ,
		_w973_
	);
	LUT4 #(
		.INIT('h0001)
	) name14 (
		\u5_state_reg[18]/NET0131 ,
		\u5_state_reg[19]/NET0131 ,
		\u5_state_reg[20]/NET0131 ,
		\u5_state_reg[21]/NET0131 ,
		_w974_
	);
	LUT2 #(
		.INIT('h1)
	) name15 (
		\u5_state_reg[22]/NET0131 ,
		\u5_state_reg[24]/NET0131 ,
		_w975_
	);
	LUT4 #(
		.INIT('h0001)
	) name16 (
		\u5_state_reg[22]/NET0131 ,
		\u5_state_reg[23]/NET0131 ,
		\u5_state_reg[24]/NET0131 ,
		\u5_state_reg[25]/NET0131 ,
		_w976_
	);
	LUT4 #(
		.INIT('h0001)
	) name17 (
		\u5_state_reg[30]/NET0131 ,
		\u5_state_reg[31]/NET0131 ,
		\u5_state_reg[32]/NET0131 ,
		\u5_state_reg[33]/NET0131 ,
		_w977_
	);
	LUT2 #(
		.INIT('h8)
	) name18 (
		_w976_,
		_w977_,
		_w978_
	);
	LUT4 #(
		.INIT('h8000)
	) name19 (
		_w973_,
		_w974_,
		_w976_,
		_w977_,
		_w979_
	);
	LUT4 #(
		.INIT('h0001)
	) name20 (
		\u5_state_reg[14]/NET0131 ,
		\u5_state_reg[15]/NET0131 ,
		\u5_state_reg[16]/NET0131 ,
		\u5_state_reg[17]/NET0131 ,
		_w980_
	);
	LUT4 #(
		.INIT('h0001)
	) name21 (
		\u5_state_reg[6]/NET0131 ,
		\u5_state_reg[7]/NET0131 ,
		\u5_state_reg[8]/NET0131 ,
		\u5_state_reg[9]/NET0131 ,
		_w981_
	);
	LUT4 #(
		.INIT('h0001)
	) name22 (
		\u5_state_reg[10]/NET0131 ,
		\u5_state_reg[11]/NET0131 ,
		\u5_state_reg[12]/NET0131 ,
		\u5_state_reg[13]/NET0131 ,
		_w982_
	);
	LUT4 #(
		.INIT('h0001)
	) name23 (
		\u5_state_reg[2]/NET0131 ,
		\u5_state_reg[3]/NET0131 ,
		\u5_state_reg[4]/NET0131 ,
		\u5_state_reg[5]/NET0131 ,
		_w983_
	);
	LUT4 #(
		.INIT('h8000)
	) name24 (
		_w980_,
		_w981_,
		_w982_,
		_w983_,
		_w984_
	);
	LUT4 #(
		.INIT('h0001)
	) name25 (
		\u5_state_reg[62]/NET0131 ,
		\u5_state_reg[63]/NET0131 ,
		\u5_state_reg[64]/NET0131 ,
		\u5_state_reg[65]/NET0131 ,
		_w985_
	);
	LUT2 #(
		.INIT('h1)
	) name26 (
		\u5_state_reg[60]/NET0131 ,
		\u5_state_reg[61]/NET0131 ,
		_w986_
	);
	LUT2 #(
		.INIT('h1)
	) name27 (
		\u5_state_reg[58]/NET0131 ,
		\u5_state_reg[59]/NET0131 ,
		_w987_
	);
	LUT4 #(
		.INIT('h0001)
	) name28 (
		\u5_state_reg[58]/NET0131 ,
		\u5_state_reg[59]/NET0131 ,
		\u5_state_reg[60]/NET0131 ,
		\u5_state_reg[61]/NET0131 ,
		_w988_
	);
	LUT2 #(
		.INIT('h1)
	) name29 (
		\u5_state_reg[0]/NET0131 ,
		\u5_state_reg[1]/NET0131 ,
		_w989_
	);
	LUT3 #(
		.INIT('h80)
	) name30 (
		_w985_,
		_w988_,
		_w989_,
		_w990_
	);
	LUT4 #(
		.INIT('h8000)
	) name31 (
		_w971_,
		_w979_,
		_w984_,
		_w990_,
		_w991_
	);
	LUT2 #(
		.INIT('h1)
	) name32 (
		\u5_state_reg[50]/NET0131 ,
		\u5_state_reg[51]/NET0131 ,
		_w992_
	);
	LUT4 #(
		.INIT('h0001)
	) name33 (
		\u5_state_reg[50]/NET0131 ,
		\u5_state_reg[51]/NET0131 ,
		\u5_state_reg[52]/NET0131 ,
		\u5_state_reg[53]/NET0131 ,
		_w993_
	);
	LUT3 #(
		.INIT('h02)
	) name34 (
		\u5_state_reg[54]/NET0131 ,
		\u5_state_reg[55]/NET0131 ,
		\u5_state_reg[57]/NET0131 ,
		_w994_
	);
	LUT3 #(
		.INIT('h40)
	) name35 (
		\u5_state_reg[56]/NET0131 ,
		_w993_,
		_w994_,
		_w995_
	);
	LUT2 #(
		.INIT('h8)
	) name36 (
		_w991_,
		_w995_,
		_w996_
	);
	LUT2 #(
		.INIT('h4)
	) name37 (
		\u5_dv_r_reg/NET0131 ,
		\u5_mc_adv_r_reg/NET0131 ,
		_w997_
	);
	LUT3 #(
		.INIT('h80)
	) name38 (
		_w991_,
		_w995_,
		_w997_,
		_w998_
	);
	LUT4 #(
		.INIT('h0001)
	) name39 (
		\u5_state_reg[54]/NET0131 ,
		\u5_state_reg[55]/NET0131 ,
		\u5_state_reg[56]/NET0131 ,
		\u5_state_reg[57]/NET0131 ,
		_w999_
	);
	LUT2 #(
		.INIT('h8)
	) name40 (
		_w993_,
		_w999_,
		_w1000_
	);
	LUT4 #(
		.INIT('h8000)
	) name41 (
		_w980_,
		_w981_,
		_w993_,
		_w999_,
		_w1001_
	);
	LUT4 #(
		.INIT('h8000)
	) name42 (
		_w971_,
		_w979_,
		_w990_,
		_w1001_,
		_w1002_
	);
	LUT3 #(
		.INIT('h01)
	) name43 (
		\u5_state_reg[2]/NET0131 ,
		\u5_state_reg[3]/NET0131 ,
		\u5_state_reg[4]/NET0131 ,
		_w1003_
	);
	LUT3 #(
		.INIT('h01)
	) name44 (
		\u5_state_reg[12]/NET0131 ,
		\u5_state_reg[13]/NET0131 ,
		\u5_state_reg[5]/NET0131 ,
		_w1004_
	);
	LUT2 #(
		.INIT('h8)
	) name45 (
		_w1003_,
		_w1004_,
		_w1005_
	);
	LUT2 #(
		.INIT('h4)
	) name46 (
		\u5_state_reg[10]/NET0131 ,
		\u5_state_reg[11]/NET0131 ,
		_w1006_
	);
	LUT2 #(
		.INIT('h4)
	) name47 (
		\u5_cnt_reg/NET0131 ,
		\u5_wb_cycle_reg/NET0131 ,
		_w1007_
	);
	LUT4 #(
		.INIT('h0800)
	) name48 (
		\u5_burst_act_rd_reg/P0001 ,
		\u5_cke_o_del_reg/P0001 ,
		\u5_cnt_reg/NET0131 ,
		\u5_wb_cycle_reg/NET0131 ,
		_w1008_
	);
	LUT2 #(
		.INIT('h8)
	) name49 (
		_w1006_,
		_w1008_,
		_w1009_
	);
	LUT3 #(
		.INIT('h80)
	) name50 (
		_w1002_,
		_w1005_,
		_w1009_,
		_w1010_
	);
	LUT2 #(
		.INIT('he)
	) name51 (
		_w998_,
		_w1010_,
		_w1011_
	);
	LUT3 #(
		.INIT('ha8)
	) name52 (
		\u3_u0_wr_adr_reg[3]/NET0131 ,
		_w998_,
		_w1010_,
		_w1012_
	);
	LUT2 #(
		.INIT('h8)
	) name53 (
		wb_cyc_i_pad,
		wb_stb_i_pad,
		_w1013_
	);
	LUT3 #(
		.INIT('h80)
	) name54 (
		wb_cyc_i_pad,
		wb_stb_i_pad,
		wb_we_i_pad,
		_w1014_
	);
	LUT2 #(
		.INIT('h2)
	) name55 (
		\u6_rmw_en_reg/NET0131 ,
		\u6_wr_hold_reg/NET0131 ,
		_w1015_
	);
	LUT2 #(
		.INIT('h8)
	) name56 (
		_w1014_,
		_w1015_,
		_w1016_
	);
	LUT2 #(
		.INIT('h2)
	) name57 (
		\u5_state_reg[6]/NET0131 ,
		\u5_wb_wait_r_reg/P0001 ,
		_w1017_
	);
	LUT4 #(
		.INIT('h8000)
	) name58 (
		_w970_,
		_w988_,
		_w993_,
		_w999_,
		_w1018_
	);
	LUT2 #(
		.INIT('h8)
	) name59 (
		_w966_,
		_w1018_,
		_w1019_
	);
	LUT4 #(
		.INIT('h0001)
	) name60 (
		\u5_state_reg[10]/NET0131 ,
		\u5_state_reg[11]/NET0131 ,
		\u5_state_reg[8]/NET0131 ,
		\u5_state_reg[9]/NET0131 ,
		_w1020_
	);
	LUT4 #(
		.INIT('h0001)
	) name61 (
		\u5_state_reg[12]/NET0131 ,
		\u5_state_reg[13]/NET0131 ,
		\u5_state_reg[15]/NET0131 ,
		\u5_state_reg[16]/NET0131 ,
		_w1021_
	);
	LUT2 #(
		.INIT('h8)
	) name62 (
		_w1020_,
		_w1021_,
		_w1022_
	);
	LUT2 #(
		.INIT('h1)
	) name63 (
		\u5_state_reg[5]/NET0131 ,
		\u5_state_reg[6]/NET0131 ,
		_w1023_
	);
	LUT3 #(
		.INIT('h10)
	) name64 (
		\u5_state_reg[14]/NET0131 ,
		\u5_state_reg[17]/NET0131 ,
		\u5_state_reg[7]/NET0131 ,
		_w1024_
	);
	LUT4 #(
		.INIT('h8000)
	) name65 (
		_w973_,
		_w974_,
		_w1023_,
		_w1024_,
		_w1025_
	);
	LUT3 #(
		.INIT('h01)
	) name66 (
		\u5_state_reg[30]/NET0131 ,
		\u5_state_reg[31]/NET0131 ,
		\u5_state_reg[32]/NET0131 ,
		_w1026_
	);
	LUT3 #(
		.INIT('hfe)
	) name67 (
		\u5_state_reg[30]/NET0131 ,
		\u5_state_reg[31]/NET0131 ,
		\u5_state_reg[32]/NET0131 ,
		_w1027_
	);
	LUT4 #(
		.INIT('h0001)
	) name68 (
		\u5_state_reg[1]/NET0131 ,
		\u5_state_reg[2]/NET0131 ,
		\u5_state_reg[3]/NET0131 ,
		\u5_state_reg[4]/NET0131 ,
		_w1028_
	);
	LUT2 #(
		.INIT('h8)
	) name69 (
		_w1026_,
		_w1028_,
		_w1029_
	);
	LUT3 #(
		.INIT('h01)
	) name70 (
		\u5_state_reg[33]/NET0131 ,
		\u5_state_reg[34]/NET0131 ,
		\u5_state_reg[35]/NET0131 ,
		_w1030_
	);
	LUT3 #(
		.INIT('h01)
	) name71 (
		\u5_state_reg[0]/NET0131 ,
		\u5_state_reg[36]/NET0131 ,
		\u5_state_reg[37]/NET0131 ,
		_w1031_
	);
	LUT4 #(
		.INIT('h8000)
	) name72 (
		_w976_,
		_w985_,
		_w1030_,
		_w1031_,
		_w1032_
	);
	LUT4 #(
		.INIT('h8000)
	) name73 (
		_w1022_,
		_w1025_,
		_w1029_,
		_w1032_,
		_w1033_
	);
	LUT3 #(
		.INIT('h15)
	) name74 (
		_w1017_,
		_w1019_,
		_w1033_,
		_w1034_
	);
	LUT4 #(
		.INIT('h8000)
	) name75 (
		_w971_,
		_w973_,
		_w990_,
		_w1000_,
		_w1035_
	);
	LUT2 #(
		.INIT('h8)
	) name76 (
		_w974_,
		_w976_,
		_w1036_
	);
	LUT4 #(
		.INIT('h0100)
	) name77 (
		\u5_state_reg[30]/NET0131 ,
		\u5_state_reg[31]/NET0131 ,
		\u5_state_reg[32]/NET0131 ,
		\u5_state_reg[33]/NET0131 ,
		_w1037_
	);
	LUT3 #(
		.INIT('h80)
	) name78 (
		_w984_,
		_w1036_,
		_w1037_,
		_w1038_
	);
	LUT2 #(
		.INIT('h8)
	) name79 (
		_w1035_,
		_w1038_,
		_w1039_
	);
	LUT4 #(
		.INIT('h8000)
	) name80 (
		_w963_,
		_w965_,
		_w993_,
		_w999_,
		_w1040_
	);
	LUT4 #(
		.INIT('h8000)
	) name81 (
		_w979_,
		_w984_,
		_w990_,
		_w1040_,
		_w1041_
	);
	LUT4 #(
		.INIT('h0002)
	) name82 (
		\u5_state_reg[34]/NET0131 ,
		\u5_state_reg[35]/NET0131 ,
		\u5_state_reg[36]/NET0131 ,
		\u5_state_reg[37]/NET0131 ,
		_w1042_
	);
	LUT2 #(
		.INIT('h8)
	) name83 (
		_w970_,
		_w1042_,
		_w1043_
	);
	LUT4 #(
		.INIT('h0777)
	) name84 (
		_w1035_,
		_w1038_,
		_w1041_,
		_w1043_,
		_w1044_
	);
	LUT3 #(
		.INIT('h80)
	) name85 (
		_w1002_,
		_w1005_,
		_w1006_,
		_w1045_
	);
	LUT2 #(
		.INIT('h8)
	) name86 (
		_w974_,
		_w977_,
		_w1046_
	);
	LUT4 #(
		.INIT('h0004)
	) name87 (
		\u5_state_reg[22]/NET0131 ,
		\u5_state_reg[23]/NET0131 ,
		\u5_state_reg[24]/NET0131 ,
		\u5_state_reg[25]/NET0131 ,
		_w1047_
	);
	LUT3 #(
		.INIT('h80)
	) name88 (
		_w984_,
		_w1046_,
		_w1047_,
		_w1048_
	);
	LUT4 #(
		.INIT('h0002)
	) name89 (
		\u5_state_reg[30]/NET0131 ,
		\u5_state_reg[31]/NET0131 ,
		\u5_state_reg[32]/NET0131 ,
		\u5_state_reg[33]/NET0131 ,
		_w1049_
	);
	LUT3 #(
		.INIT('h80)
	) name90 (
		_w984_,
		_w1036_,
		_w1049_,
		_w1050_
	);
	LUT2 #(
		.INIT('h8)
	) name91 (
		_w1035_,
		_w1050_,
		_w1051_
	);
	LUT3 #(
		.INIT('h57)
	) name92 (
		_w1035_,
		_w1048_,
		_w1050_,
		_w1052_
	);
	LUT3 #(
		.INIT('h20)
	) name93 (
		_w1044_,
		_w1045_,
		_w1052_,
		_w1053_
	);
	LUT2 #(
		.INIT('h4)
	) name94 (
		\u5_state_reg[52]/NET0131 ,
		\u5_state_reg[53]/NET0131 ,
		_w1054_
	);
	LUT3 #(
		.INIT('h80)
	) name95 (
		_w992_,
		_w999_,
		_w1054_,
		_w1055_
	);
	LUT2 #(
		.INIT('h8)
	) name96 (
		_w991_,
		_w1055_,
		_w1056_
	);
	LUT3 #(
		.INIT('h57)
	) name97 (
		_w991_,
		_w995_,
		_w1055_,
		_w1057_
	);
	LUT3 #(
		.INIT('h80)
	) name98 (
		_w989_,
		_w993_,
		_w999_,
		_w1058_
	);
	LUT4 #(
		.INIT('h8000)
	) name99 (
		_w971_,
		_w979_,
		_w984_,
		_w1058_,
		_w1059_
	);
	LUT4 #(
		.INIT('h0100)
	) name100 (
		\u5_state_reg[62]/NET0131 ,
		\u5_state_reg[63]/NET0131 ,
		\u5_state_reg[64]/NET0131 ,
		\u5_state_reg[65]/NET0131 ,
		_w1060_
	);
	LUT2 #(
		.INIT('h8)
	) name101 (
		_w988_,
		_w1060_,
		_w1061_
	);
	LUT4 #(
		.INIT('h8000)
	) name102 (
		_w968_,
		_w970_,
		_w993_,
		_w999_,
		_w1062_
	);
	LUT4 #(
		.INIT('h8000)
	) name103 (
		_w979_,
		_w984_,
		_w990_,
		_w1062_,
		_w1063_
	);
	LUT4 #(
		.INIT('h0010)
	) name104 (
		\u5_state_reg[38]/NET0131 ,
		\u5_state_reg[39]/NET0131 ,
		\u5_state_reg[40]/NET0131 ,
		\u5_state_reg[41]/NET0131 ,
		_w1064_
	);
	LUT2 #(
		.INIT('h8)
	) name105 (
		_w965_,
		_w1064_,
		_w1065_
	);
	LUT4 #(
		.INIT('h0777)
	) name106 (
		_w1059_,
		_w1061_,
		_w1063_,
		_w1065_,
		_w1066_
	);
	LUT2 #(
		.INIT('h8)
	) name107 (
		_w1057_,
		_w1066_,
		_w1067_
	);
	LUT4 #(
		.INIT('h8000)
	) name108 (
		_w971_,
		_w974_,
		_w990_,
		_w1000_,
		_w1068_
	);
	LUT4 #(
		.INIT('h0100)
	) name109 (
		\u5_state_reg[26]/NET0131 ,
		\u5_state_reg[27]/NET0131 ,
		\u5_state_reg[28]/NET0131 ,
		\u5_state_reg[29]/NET0131 ,
		_w1069_
	);
	LUT3 #(
		.INIT('h80)
	) name110 (
		_w978_,
		_w984_,
		_w1069_,
		_w1070_
	);
	LUT2 #(
		.INIT('h8)
	) name111 (
		_w1068_,
		_w1070_,
		_w1071_
	);
	LUT3 #(
		.INIT('h08)
	) name112 (
		_w1057_,
		_w1066_,
		_w1071_,
		_w1072_
	);
	LUT2 #(
		.INIT('h8)
	) name113 (
		_w1053_,
		_w1072_,
		_w1073_
	);
	LUT2 #(
		.INIT('h2)
	) name114 (
		\u5_state_reg[10]/NET0131 ,
		\u5_state_reg[11]/NET0131 ,
		_w1074_
	);
	LUT3 #(
		.INIT('h80)
	) name115 (
		_w1002_,
		_w1005_,
		_w1074_,
		_w1075_
	);
	LUT4 #(
		.INIT('h0010)
	) name116 (
		\u5_state_reg[54]/NET0131 ,
		\u5_state_reg[55]/NET0131 ,
		\u5_state_reg[56]/NET0131 ,
		\u5_state_reg[57]/NET0131 ,
		_w1076_
	);
	LUT2 #(
		.INIT('h8)
	) name117 (
		_w993_,
		_w1076_,
		_w1077_
	);
	LUT4 #(
		.INIT('h0010)
	) name118 (
		\u5_state_reg[34]/NET0131 ,
		\u5_state_reg[35]/NET0131 ,
		\u5_state_reg[36]/NET0131 ,
		\u5_state_reg[37]/NET0131 ,
		_w1078_
	);
	LUT2 #(
		.INIT('h8)
	) name119 (
		_w970_,
		_w1078_,
		_w1079_
	);
	LUT4 #(
		.INIT('h135f)
	) name120 (
		_w991_,
		_w1041_,
		_w1077_,
		_w1079_,
		_w1080_
	);
	LUT2 #(
		.INIT('h4)
	) name121 (
		_w1075_,
		_w1080_,
		_w1081_
	);
	LUT2 #(
		.INIT('h2)
	) name122 (
		\u5_state_reg[60]/NET0131 ,
		\u5_state_reg[61]/NET0131 ,
		_w1082_
	);
	LUT3 #(
		.INIT('h80)
	) name123 (
		_w985_,
		_w987_,
		_w1082_,
		_w1083_
	);
	LUT2 #(
		.INIT('h8)
	) name124 (
		_w1059_,
		_w1083_,
		_w1084_
	);
	LUT4 #(
		.INIT('h0010)
	) name125 (
		\u5_state_reg[62]/NET0131 ,
		\u5_state_reg[63]/NET0131 ,
		\u5_state_reg[64]/NET0131 ,
		\u5_state_reg[65]/NET0131 ,
		_w1085_
	);
	LUT2 #(
		.INIT('h8)
	) name126 (
		_w988_,
		_w1085_,
		_w1086_
	);
	LUT2 #(
		.INIT('h8)
	) name127 (
		_w1059_,
		_w1086_,
		_w1087_
	);
	LUT3 #(
		.INIT('h57)
	) name128 (
		_w1059_,
		_w1083_,
		_w1086_,
		_w1088_
	);
	LUT3 #(
		.INIT('h40)
	) name129 (
		_w1075_,
		_w1080_,
		_w1088_,
		_w1089_
	);
	LUT4 #(
		.INIT('h0010)
	) name130 (
		\u5_state_reg[46]/NET0131 ,
		\u5_state_reg[47]/NET0131 ,
		\u5_state_reg[48]/NET0131 ,
		\u5_state_reg[49]/NET0131 ,
		_w1090_
	);
	LUT2 #(
		.INIT('h8)
	) name131 (
		_w968_,
		_w1090_,
		_w1091_
	);
	LUT2 #(
		.INIT('h8)
	) name132 (
		_w1041_,
		_w1091_,
		_w1092_
	);
	LUT4 #(
		.INIT('h0100)
	) name133 (
		\u5_state_reg[54]/NET0131 ,
		\u5_state_reg[55]/NET0131 ,
		\u5_state_reg[56]/NET0131 ,
		\u5_state_reg[57]/NET0131 ,
		_w1093_
	);
	LUT2 #(
		.INIT('h8)
	) name134 (
		_w993_,
		_w1093_,
		_w1094_
	);
	LUT2 #(
		.INIT('h8)
	) name135 (
		_w991_,
		_w1094_,
		_w1095_
	);
	LUT4 #(
		.INIT('h0100)
	) name136 (
		\u5_state_reg[18]/NET0131 ,
		\u5_state_reg[19]/NET0131 ,
		\u5_state_reg[20]/NET0131 ,
		\u5_state_reg[21]/NET0131 ,
		_w1096_
	);
	LUT3 #(
		.INIT('h80)
	) name137 (
		_w978_,
		_w984_,
		_w1096_,
		_w1097_
	);
	LUT4 #(
		.INIT('h135f)
	) name138 (
		_w991_,
		_w1035_,
		_w1094_,
		_w1097_,
		_w1098_
	);
	LUT4 #(
		.INIT('h8000)
	) name139 (
		_w982_,
		_w983_,
		_w993_,
		_w999_,
		_w1099_
	);
	LUT4 #(
		.INIT('h8000)
	) name140 (
		_w971_,
		_w979_,
		_w990_,
		_w1099_,
		_w1100_
	);
	LUT4 #(
		.INIT('h0100)
	) name141 (
		\u5_state_reg[14]/NET0131 ,
		\u5_state_reg[15]/NET0131 ,
		\u5_state_reg[16]/NET0131 ,
		\u5_state_reg[17]/NET0131 ,
		_w1101_
	);
	LUT2 #(
		.INIT('h8)
	) name142 (
		_w981_,
		_w1101_,
		_w1102_
	);
	LUT4 #(
		.INIT('h0100)
	) name143 (
		\u5_state_reg[6]/NET0131 ,
		\u5_state_reg[7]/NET0131 ,
		\u5_state_reg[8]/NET0131 ,
		\u5_state_reg[9]/NET0131 ,
		_w1103_
	);
	LUT2 #(
		.INIT('h8)
	) name144 (
		_w980_,
		_w1103_,
		_w1104_
	);
	LUT2 #(
		.INIT('h8)
	) name145 (
		_w1100_,
		_w1104_,
		_w1105_
	);
	LUT3 #(
		.INIT('h57)
	) name146 (
		_w1100_,
		_w1102_,
		_w1104_,
		_w1106_
	);
	LUT4 #(
		.INIT('h0010)
	) name147 (
		\u5_state_reg[6]/NET0131 ,
		\u5_state_reg[7]/NET0131 ,
		\u5_state_reg[8]/NET0131 ,
		\u5_state_reg[9]/NET0131 ,
		_w1107_
	);
	LUT2 #(
		.INIT('h8)
	) name148 (
		_w980_,
		_w1107_,
		_w1108_
	);
	LUT4 #(
		.INIT('h0004)
	) name149 (
		\u5_state_reg[6]/NET0131 ,
		\u5_state_reg[7]/NET0131 ,
		\u5_state_reg[8]/NET0131 ,
		\u5_state_reg[9]/NET0131 ,
		_w1109_
	);
	LUT2 #(
		.INIT('h8)
	) name150 (
		_w980_,
		_w1109_,
		_w1110_
	);
	LUT3 #(
		.INIT('h57)
	) name151 (
		_w1100_,
		_w1108_,
		_w1110_,
		_w1111_
	);
	LUT4 #(
		.INIT('h4000)
	) name152 (
		_w1092_,
		_w1098_,
		_w1106_,
		_w1111_,
		_w1112_
	);
	LUT4 #(
		.INIT('h8000)
	) name153 (
		_w1053_,
		_w1072_,
		_w1089_,
		_w1112_,
		_w1113_
	);
	LUT2 #(
		.INIT('h1)
	) name154 (
		\u5_lmr_ack_reg/NET0131 ,
		\u5_state_reg[26]/NET0131 ,
		_w1114_
	);
	LUT3 #(
		.INIT('h02)
	) name155 (
		\u0_tms_reg[9]/NET0131 ,
		\u5_lmr_ack_reg/NET0131 ,
		\u5_state_reg[26]/NET0131 ,
		_w1115_
	);
	LUT4 #(
		.INIT('h11d5)
	) name156 (
		\u0_sp_tms_reg[9]/NET0131 ,
		_w976_,
		_w1114_,
		_w1115_,
		_w1116_
	);
	LUT3 #(
		.INIT('h2a)
	) name157 (
		\u0_sp_csc_reg[10]/NET0131 ,
		_w976_,
		_w1114_,
		_w1117_
	);
	LUT3 #(
		.INIT('h02)
	) name158 (
		\u0_csc_reg[10]/NET0131 ,
		\u5_lmr_ack_reg/NET0131 ,
		\u5_state_reg[26]/NET0131 ,
		_w1118_
	);
	LUT4 #(
		.INIT('h11d5)
	) name159 (
		\u0_sp_csc_reg[10]/NET0131 ,
		_w976_,
		_w1114_,
		_w1118_,
		_w1119_
	);
	LUT2 #(
		.INIT('h4)
	) name160 (
		_w1116_,
		_w1119_,
		_w1120_
	);
	LUT3 #(
		.INIT('h02)
	) name161 (
		\u0_tms_reg[1]/NET0131 ,
		\u5_lmr_ack_reg/NET0131 ,
		\u5_state_reg[26]/NET0131 ,
		_w1121_
	);
	LUT4 #(
		.INIT('h11d5)
	) name162 (
		\u0_sp_tms_reg[1]/NET0131 ,
		_w976_,
		_w1114_,
		_w1121_,
		_w1122_
	);
	LUT3 #(
		.INIT('h02)
	) name163 (
		\u0_tms_reg[2]/NET0131 ,
		\u5_lmr_ack_reg/NET0131 ,
		\u5_state_reg[26]/NET0131 ,
		_w1123_
	);
	LUT4 #(
		.INIT('h11d5)
	) name164 (
		\u0_sp_tms_reg[2]/NET0131 ,
		_w976_,
		_w1114_,
		_w1123_,
		_w1124_
	);
	LUT2 #(
		.INIT('h8)
	) name165 (
		_w1122_,
		_w1124_,
		_w1125_
	);
	LUT3 #(
		.INIT('h02)
	) name166 (
		\u0_tms_reg[0]/NET0131 ,
		\u5_lmr_ack_reg/NET0131 ,
		\u5_state_reg[26]/NET0131 ,
		_w1126_
	);
	LUT4 #(
		.INIT('h11d5)
	) name167 (
		\u0_sp_tms_reg[0]/NET0131 ,
		_w976_,
		_w1114_,
		_w1126_,
		_w1127_
	);
	LUT4 #(
		.INIT('h8000)
	) name168 (
		_w1119_,
		_w1122_,
		_w1124_,
		_w1127_,
		_w1128_
	);
	LUT2 #(
		.INIT('h1)
	) name169 (
		_w1120_,
		_w1128_,
		_w1129_
	);
	LUT2 #(
		.INIT('h2)
	) name170 (
		wb_stb_i_pad,
		wb_we_i_pad,
		_w1130_
	);
	LUT3 #(
		.INIT('ha2)
	) name171 (
		\u6_write_go_r1_reg/NET0131 ,
		wb_stb_i_pad,
		wb_we_i_pad,
		_w1131_
	);
	LUT2 #(
		.INIT('h2)
	) name172 (
		wb_cyc_i_pad,
		wb_stb_i_pad,
		_w1132_
	);
	LUT2 #(
		.INIT('h4)
	) name173 (
		\u6_rmw_r_reg/NET0131 ,
		wb_cyc_i_pad,
		_w1133_
	);
	LUT3 #(
		.INIT('h40)
	) name174 (
		\u6_rmw_r_reg/NET0131 ,
		wb_cyc_i_pad,
		wb_stb_i_pad,
		_w1134_
	);
	LUT4 #(
		.INIT('h7000)
	) name175 (
		_w1014_,
		_w1015_,
		_w1131_,
		_w1134_,
		_w1135_
	);
	LUT3 #(
		.INIT('h80)
	) name176 (
		_w1100_,
		_w1108_,
		_w1135_,
		_w1136_
	);
	LUT2 #(
		.INIT('h4)
	) name177 (
		_w1129_,
		_w1136_,
		_w1137_
	);
	LUT3 #(
		.INIT('h45)
	) name178 (
		\u5_ap_en_reg/NET0131 ,
		_w1113_,
		_w1137_,
		_w1138_
	);
	LUT4 #(
		.INIT('h0002)
	) name179 (
		\u5_state_reg[14]/NET0131 ,
		\u5_state_reg[15]/NET0131 ,
		\u5_state_reg[16]/NET0131 ,
		\u5_state_reg[17]/NET0131 ,
		_w1139_
	);
	LUT2 #(
		.INIT('h8)
	) name180 (
		_w981_,
		_w1139_,
		_w1140_
	);
	LUT2 #(
		.INIT('h8)
	) name181 (
		_w1100_,
		_w1140_,
		_w1141_
	);
	LUT3 #(
		.INIT('h01)
	) name182 (
		\u5_state_reg[10]/NET0131 ,
		\u5_state_reg[11]/NET0131 ,
		\u5_state_reg[5]/NET0131 ,
		_w1142_
	);
	LUT2 #(
		.INIT('h8)
	) name183 (
		_w1003_,
		_w1142_,
		_w1143_
	);
	LUT2 #(
		.INIT('h4)
	) name184 (
		\u5_state_reg[12]/NET0131 ,
		\u5_state_reg[13]/NET0131 ,
		_w1144_
	);
	LUT3 #(
		.INIT('h80)
	) name185 (
		_w1002_,
		_w1143_,
		_w1144_,
		_w1145_
	);
	LUT2 #(
		.INIT('h1)
	) name186 (
		_w1141_,
		_w1145_,
		_w1146_
	);
	LUT2 #(
		.INIT('h1)
	) name187 (
		\u5_state_reg[18]/NET0131 ,
		\u5_state_reg[21]/NET0131 ,
		_w1147_
	);
	LUT3 #(
		.INIT('h80)
	) name188 (
		_w978_,
		_w984_,
		_w1147_,
		_w1148_
	);
	LUT2 #(
		.INIT('h2)
	) name189 (
		\u5_state_reg[19]/NET0131 ,
		\u5_state_reg[20]/NET0131 ,
		_w1149_
	);
	LUT3 #(
		.INIT('h80)
	) name190 (
		_w1035_,
		_w1148_,
		_w1149_,
		_w1150_
	);
	LUT4 #(
		.INIT('h0100)
	) name191 (
		\u5_state_reg[46]/NET0131 ,
		\u5_state_reg[47]/NET0131 ,
		\u5_state_reg[48]/NET0131 ,
		\u5_state_reg[49]/NET0131 ,
		_w1151_
	);
	LUT2 #(
		.INIT('h8)
	) name192 (
		_w968_,
		_w1151_,
		_w1152_
	);
	LUT2 #(
		.INIT('h8)
	) name193 (
		_w1041_,
		_w1152_,
		_w1153_
	);
	LUT4 #(
		.INIT('h0002)
	) name194 (
		\u5_state_reg[26]/NET0131 ,
		\u5_state_reg[27]/NET0131 ,
		\u5_state_reg[28]/NET0131 ,
		\u5_state_reg[29]/NET0131 ,
		_w1154_
	);
	LUT3 #(
		.INIT('h80)
	) name195 (
		_w978_,
		_w984_,
		_w1154_,
		_w1155_
	);
	LUT2 #(
		.INIT('h8)
	) name196 (
		_w1068_,
		_w1155_,
		_w1156_
	);
	LUT4 #(
		.INIT('h0004)
	) name197 (
		\u5_state_reg[14]/NET0131 ,
		\u5_state_reg[15]/NET0131 ,
		\u5_state_reg[16]/NET0131 ,
		\u5_state_reg[17]/NET0131 ,
		_w1157_
	);
	LUT2 #(
		.INIT('h8)
	) name198 (
		_w981_,
		_w1157_,
		_w1158_
	);
	LUT2 #(
		.INIT('h8)
	) name199 (
		_w1100_,
		_w1158_,
		_w1159_
	);
	LUT4 #(
		.INIT('h0002)
	) name200 (
		\u5_state_reg[6]/NET0131 ,
		\u5_state_reg[7]/NET0131 ,
		\u5_state_reg[8]/NET0131 ,
		\u5_state_reg[9]/NET0131 ,
		_w1160_
	);
	LUT2 #(
		.INIT('h8)
	) name201 (
		_w980_,
		_w1160_,
		_w1161_
	);
	LUT3 #(
		.INIT('h57)
	) name202 (
		_w1100_,
		_w1158_,
		_w1161_,
		_w1162_
	);
	LUT4 #(
		.INIT('h0100)
	) name203 (
		_w1150_,
		_w1153_,
		_w1156_,
		_w1162_,
		_w1163_
	);
	LUT2 #(
		.INIT('h8)
	) name204 (
		_w1146_,
		_w1163_,
		_w1164_
	);
	LUT3 #(
		.INIT('h04)
	) name205 (
		\u5_state_reg[2]/NET0131 ,
		\u5_state_reg[3]/NET0131 ,
		\u5_state_reg[4]/NET0131 ,
		_w1165_
	);
	LUT3 #(
		.INIT('h40)
	) name206 (
		\u5_state_reg[5]/NET0131 ,
		_w982_,
		_w1165_,
		_w1166_
	);
	LUT4 #(
		.INIT('h0010)
	) name207 (
		\u5_state_reg[30]/NET0131 ,
		\u5_state_reg[31]/NET0131 ,
		\u5_state_reg[32]/NET0131 ,
		\u5_state_reg[33]/NET0131 ,
		_w1167_
	);
	LUT3 #(
		.INIT('h80)
	) name208 (
		_w984_,
		_w1036_,
		_w1167_,
		_w1168_
	);
	LUT2 #(
		.INIT('h8)
	) name209 (
		_w1035_,
		_w1168_,
		_w1169_
	);
	LUT4 #(
		.INIT('h135f)
	) name210 (
		_w1002_,
		_w1035_,
		_w1166_,
		_w1168_,
		_w1170_
	);
	LUT4 #(
		.INIT('h0004)
	) name211 (
		\u5_state_reg[62]/NET0131 ,
		\u5_state_reg[63]/NET0131 ,
		\u5_state_reg[64]/NET0131 ,
		\u5_state_reg[65]/NET0131 ,
		_w1171_
	);
	LUT2 #(
		.INIT('h8)
	) name212 (
		_w988_,
		_w1171_,
		_w1172_
	);
	LUT2 #(
		.INIT('h8)
	) name213 (
		_w1059_,
		_w1172_,
		_w1173_
	);
	LUT4 #(
		.INIT('h8000)
	) name214 (
		_w971_,
		_w979_,
		_w984_,
		_w989_,
		_w1174_
	);
	LUT4 #(
		.INIT('h0001)
	) name215 (
		\u5_state_reg[52]/NET0131 ,
		\u5_state_reg[53]/NET0131 ,
		\u5_state_reg[58]/NET0131 ,
		\u5_state_reg[59]/NET0131 ,
		_w1175_
	);
	LUT4 #(
		.INIT('h8000)
	) name216 (
		_w985_,
		_w986_,
		_w999_,
		_w1175_,
		_w1176_
	);
	LUT2 #(
		.INIT('h2)
	) name217 (
		\u5_state_reg[50]/NET0131 ,
		\u5_state_reg[51]/NET0131 ,
		_w1177_
	);
	LUT2 #(
		.INIT('h8)
	) name218 (
		_w1176_,
		_w1177_,
		_w1178_
	);
	LUT4 #(
		.INIT('h0777)
	) name219 (
		_w1059_,
		_w1172_,
		_w1174_,
		_w1178_,
		_w1179_
	);
	LUT2 #(
		.INIT('h8)
	) name220 (
		_w1170_,
		_w1179_,
		_w1180_
	);
	LUT4 #(
		.INIT('h0100)
	) name221 (
		\u5_state_reg[2]/NET0131 ,
		\u5_state_reg[3]/NET0131 ,
		\u5_state_reg[4]/NET0131 ,
		\u5_state_reg[5]/NET0131 ,
		_w1181_
	);
	LUT2 #(
		.INIT('h8)
	) name222 (
		_w982_,
		_w1181_,
		_w1182_
	);
	LUT4 #(
		.INIT('h8000)
	) name223 (
		_w985_,
		_w988_,
		_w993_,
		_w999_,
		_w1183_
	);
	LUT4 #(
		.INIT('h8000)
	) name224 (
		_w971_,
		_w979_,
		_w984_,
		_w1183_,
		_w1184_
	);
	LUT2 #(
		.INIT('h4)
	) name225 (
		\u5_state_reg[0]/NET0131 ,
		\u5_state_reg[1]/NET0131 ,
		_w1185_
	);
	LUT2 #(
		.INIT('h8)
	) name226 (
		_w1184_,
		_w1185_,
		_w1186_
	);
	LUT4 #(
		.INIT('h0777)
	) name227 (
		_w1002_,
		_w1182_,
		_w1184_,
		_w1185_,
		_w1187_
	);
	LUT2 #(
		.INIT('h4)
	) name228 (
		\u5_state_reg[58]/NET0131 ,
		\u5_state_reg[59]/NET0131 ,
		_w1188_
	);
	LUT3 #(
		.INIT('h80)
	) name229 (
		_w985_,
		_w986_,
		_w1188_,
		_w1189_
	);
	LUT2 #(
		.INIT('h8)
	) name230 (
		_w1059_,
		_w1189_,
		_w1190_
	);
	LUT2 #(
		.INIT('h4)
	) name231 (
		\u5_state_reg[19]/NET0131 ,
		\u5_state_reg[20]/NET0131 ,
		_w1191_
	);
	LUT3 #(
		.INIT('h80)
	) name232 (
		_w1035_,
		_w1148_,
		_w1191_,
		_w1192_
	);
	LUT3 #(
		.INIT('h02)
	) name233 (
		_w1187_,
		_w1190_,
		_w1192_,
		_w1193_
	);
	LUT4 #(
		.INIT('h0100)
	) name234 (
		\u5_state_reg[34]/NET0131 ,
		\u5_state_reg[35]/NET0131 ,
		\u5_state_reg[36]/NET0131 ,
		\u5_state_reg[37]/NET0131 ,
		_w1194_
	);
	LUT2 #(
		.INIT('h8)
	) name235 (
		_w970_,
		_w1194_,
		_w1195_
	);
	LUT2 #(
		.INIT('h8)
	) name236 (
		_w1041_,
		_w1195_,
		_w1196_
	);
	LUT4 #(
		.INIT('h0004)
	) name237 (
		\u5_state_reg[30]/NET0131 ,
		\u5_state_reg[31]/NET0131 ,
		\u5_state_reg[32]/NET0131 ,
		\u5_state_reg[33]/NET0131 ,
		_w1197_
	);
	LUT3 #(
		.INIT('h80)
	) name238 (
		_w984_,
		_w1036_,
		_w1197_,
		_w1198_
	);
	LUT2 #(
		.INIT('h8)
	) name239 (
		_w1035_,
		_w1198_,
		_w1199_
	);
	LUT4 #(
		.INIT('h0010)
	) name240 (
		\u5_state_reg[26]/NET0131 ,
		\u5_state_reg[27]/NET0131 ,
		\u5_state_reg[28]/NET0131 ,
		\u5_state_reg[29]/NET0131 ,
		_w1200_
	);
	LUT3 #(
		.INIT('h80)
	) name241 (
		_w978_,
		_w984_,
		_w1200_,
		_w1201_
	);
	LUT4 #(
		.INIT('h135f)
	) name242 (
		_w1035_,
		_w1068_,
		_w1198_,
		_w1201_,
		_w1202_
	);
	LUT4 #(
		.INIT('h0004)
	) name243 (
		\u5_state_reg[38]/NET0131 ,
		\u5_state_reg[39]/NET0131 ,
		\u5_state_reg[40]/NET0131 ,
		\u5_state_reg[41]/NET0131 ,
		_w1203_
	);
	LUT2 #(
		.INIT('h8)
	) name244 (
		_w965_,
		_w1203_,
		_w1204_
	);
	LUT2 #(
		.INIT('h8)
	) name245 (
		_w1063_,
		_w1204_,
		_w1205_
	);
	LUT2 #(
		.INIT('h2)
	) name246 (
		\u5_state_reg[0]/NET0131 ,
		\u5_state_reg[1]/NET0131 ,
		_w1206_
	);
	LUT2 #(
		.INIT('h8)
	) name247 (
		_w1184_,
		_w1206_,
		_w1207_
	);
	LUT4 #(
		.INIT('h135f)
	) name248 (
		_w1063_,
		_w1184_,
		_w1204_,
		_w1206_,
		_w1208_
	);
	LUT3 #(
		.INIT('h40)
	) name249 (
		_w1196_,
		_w1202_,
		_w1208_,
		_w1209_
	);
	LUT2 #(
		.INIT('h2)
	) name250 (
		\u5_state_reg[58]/NET0131 ,
		\u5_state_reg[59]/NET0131 ,
		_w1210_
	);
	LUT3 #(
		.INIT('h80)
	) name251 (
		_w985_,
		_w986_,
		_w1210_,
		_w1211_
	);
	LUT2 #(
		.INIT('h2)
	) name252 (
		\u5_state_reg[52]/NET0131 ,
		\u5_state_reg[53]/NET0131 ,
		_w1212_
	);
	LUT3 #(
		.INIT('h80)
	) name253 (
		_w992_,
		_w999_,
		_w1212_,
		_w1213_
	);
	LUT2 #(
		.INIT('h8)
	) name254 (
		_w991_,
		_w1213_,
		_w1214_
	);
	LUT4 #(
		.INIT('h153f)
	) name255 (
		_w991_,
		_w1059_,
		_w1211_,
		_w1213_,
		_w1215_
	);
	LUT4 #(
		.INIT('h0004)
	) name256 (
		\u5_state_reg[46]/NET0131 ,
		\u5_state_reg[47]/NET0131 ,
		\u5_state_reg[48]/NET0131 ,
		\u5_state_reg[49]/NET0131 ,
		_w1216_
	);
	LUT2 #(
		.INIT('h8)
	) name257 (
		_w968_,
		_w1216_,
		_w1217_
	);
	LUT2 #(
		.INIT('h8)
	) name258 (
		_w1041_,
		_w1217_,
		_w1218_
	);
	LUT4 #(
		.INIT('h0100)
	) name259 (
		\u5_state_reg[38]/NET0131 ,
		\u5_state_reg[39]/NET0131 ,
		\u5_state_reg[40]/NET0131 ,
		\u5_state_reg[41]/NET0131 ,
		_w1219_
	);
	LUT4 #(
		.INIT('hfefd)
	) name260 (
		\u5_state_reg[38]/NET0131 ,
		\u5_state_reg[39]/NET0131 ,
		\u5_state_reg[40]/NET0131 ,
		\u5_state_reg[41]/NET0131 ,
		_w1220_
	);
	LUT2 #(
		.INIT('h2)
	) name261 (
		_w965_,
		_w1220_,
		_w1221_
	);
	LUT2 #(
		.INIT('h4)
	) name262 (
		\u5_state_reg[60]/NET0131 ,
		\u5_state_reg[61]/NET0131 ,
		_w1222_
	);
	LUT3 #(
		.INIT('h80)
	) name263 (
		_w985_,
		_w987_,
		_w1222_,
		_w1223_
	);
	LUT4 #(
		.INIT('h153f)
	) name264 (
		_w1059_,
		_w1063_,
		_w1221_,
		_w1223_,
		_w1224_
	);
	LUT3 #(
		.INIT('h20)
	) name265 (
		_w1215_,
		_w1218_,
		_w1224_,
		_w1225_
	);
	LUT4 #(
		.INIT('h8000)
	) name266 (
		_w1180_,
		_w1193_,
		_w1209_,
		_w1225_,
		_w1226_
	);
	LUT4 #(
		.INIT('h0100)
	) name267 (
		\u5_state_reg[22]/NET0131 ,
		\u5_state_reg[23]/NET0131 ,
		\u5_state_reg[24]/NET0131 ,
		\u5_state_reg[25]/NET0131 ,
		_w1227_
	);
	LUT3 #(
		.INIT('h80)
	) name268 (
		_w984_,
		_w1046_,
		_w1227_,
		_w1228_
	);
	LUT2 #(
		.INIT('h4)
	) name269 (
		\u5_state_reg[50]/NET0131 ,
		\u5_state_reg[51]/NET0131 ,
		_w1229_
	);
	LUT2 #(
		.INIT('h8)
	) name270 (
		_w1176_,
		_w1229_,
		_w1230_
	);
	LUT2 #(
		.INIT('h8)
	) name271 (
		_w1174_,
		_w1230_,
		_w1231_
	);
	LUT4 #(
		.INIT('h135f)
	) name272 (
		_w1035_,
		_w1174_,
		_w1228_,
		_w1230_,
		_w1232_
	);
	LUT2 #(
		.INIT('h2)
	) name273 (
		\u5_state_reg[44]/NET0131 ,
		\u5_state_reg[45]/NET0131 ,
		_w1233_
	);
	LUT2 #(
		.INIT('h1)
	) name274 (
		\u5_state_reg[42]/NET0131 ,
		\u5_state_reg[43]/NET0131 ,
		_w1234_
	);
	LUT2 #(
		.INIT('h8)
	) name275 (
		_w963_,
		_w1234_,
		_w1235_
	);
	LUT3 #(
		.INIT('h80)
	) name276 (
		_w963_,
		_w1233_,
		_w1234_,
		_w1236_
	);
	LUT2 #(
		.INIT('h8)
	) name277 (
		_w1063_,
		_w1236_,
		_w1237_
	);
	LUT2 #(
		.INIT('h1)
	) name278 (
		\u5_state_reg[44]/NET0131 ,
		\u5_state_reg[45]/NET0131 ,
		_w1238_
	);
	LUT2 #(
		.INIT('h2)
	) name279 (
		\u5_state_reg[42]/NET0131 ,
		\u5_state_reg[43]/NET0131 ,
		_w1239_
	);
	LUT3 #(
		.INIT('h80)
	) name280 (
		_w963_,
		_w1238_,
		_w1239_,
		_w1240_
	);
	LUT3 #(
		.INIT('h57)
	) name281 (
		_w1063_,
		_w1236_,
		_w1240_,
		_w1241_
	);
	LUT2 #(
		.INIT('h4)
	) name282 (
		\u5_state_reg[44]/NET0131 ,
		\u5_state_reg[45]/NET0131 ,
		_w1242_
	);
	LUT3 #(
		.INIT('h80)
	) name283 (
		_w963_,
		_w1234_,
		_w1242_,
		_w1243_
	);
	LUT2 #(
		.INIT('h8)
	) name284 (
		_w1063_,
		_w1243_,
		_w1244_
	);
	LUT2 #(
		.INIT('h4)
	) name285 (
		\u5_state_reg[42]/NET0131 ,
		\u5_state_reg[43]/NET0131 ,
		_w1245_
	);
	LUT3 #(
		.INIT('h80)
	) name286 (
		_w963_,
		_w1238_,
		_w1245_,
		_w1246_
	);
	LUT2 #(
		.INIT('h8)
	) name287 (
		_w1063_,
		_w1246_,
		_w1247_
	);
	LUT3 #(
		.INIT('h57)
	) name288 (
		_w1063_,
		_w1243_,
		_w1246_,
		_w1248_
	);
	LUT3 #(
		.INIT('h04)
	) name289 (
		\u5_state_reg[54]/NET0131 ,
		\u5_state_reg[55]/NET0131 ,
		\u5_state_reg[57]/NET0131 ,
		_w1249_
	);
	LUT3 #(
		.INIT('h40)
	) name290 (
		\u5_state_reg[56]/NET0131 ,
		_w993_,
		_w1249_,
		_w1250_
	);
	LUT4 #(
		.INIT('h0002)
	) name291 (
		\u5_state_reg[62]/NET0131 ,
		\u5_state_reg[63]/NET0131 ,
		\u5_state_reg[64]/NET0131 ,
		\u5_state_reg[65]/NET0131 ,
		_w1251_
	);
	LUT2 #(
		.INIT('h8)
	) name292 (
		_w988_,
		_w1251_,
		_w1252_
	);
	LUT4 #(
		.INIT('h135f)
	) name293 (
		_w991_,
		_w1059_,
		_w1250_,
		_w1252_,
		_w1253_
	);
	LUT4 #(
		.INIT('h8000)
	) name294 (
		_w1232_,
		_w1241_,
		_w1248_,
		_w1253_,
		_w1254_
	);
	LUT4 #(
		.INIT('h0004)
	) name295 (
		\u5_state_reg[34]/NET0131 ,
		\u5_state_reg[35]/NET0131 ,
		\u5_state_reg[36]/NET0131 ,
		\u5_state_reg[37]/NET0131 ,
		_w1255_
	);
	LUT2 #(
		.INIT('h8)
	) name296 (
		_w970_,
		_w1255_,
		_w1256_
	);
	LUT2 #(
		.INIT('h8)
	) name297 (
		_w1041_,
		_w1256_,
		_w1257_
	);
	LUT2 #(
		.INIT('h2)
	) name298 (
		\u5_state_reg[12]/NET0131 ,
		\u5_state_reg[13]/NET0131 ,
		_w1258_
	);
	LUT3 #(
		.INIT('h80)
	) name299 (
		_w1002_,
		_w1143_,
		_w1258_,
		_w1259_
	);
	LUT4 #(
		.INIT('h0002)
	) name300 (
		\u5_state_reg[46]/NET0131 ,
		\u5_state_reg[47]/NET0131 ,
		\u5_state_reg[48]/NET0131 ,
		\u5_state_reg[49]/NET0131 ,
		_w1260_
	);
	LUT2 #(
		.INIT('h8)
	) name301 (
		_w968_,
		_w1260_,
		_w1261_
	);
	LUT2 #(
		.INIT('h8)
	) name302 (
		_w1041_,
		_w1261_,
		_w1262_
	);
	LUT4 #(
		.INIT('h0010)
	) name303 (
		\u5_state_reg[22]/NET0131 ,
		\u5_state_reg[23]/NET0131 ,
		\u5_state_reg[24]/NET0131 ,
		\u5_state_reg[25]/NET0131 ,
		_w1263_
	);
	LUT3 #(
		.INIT('h80)
	) name304 (
		_w984_,
		_w1046_,
		_w1263_,
		_w1264_
	);
	LUT4 #(
		.INIT('h153f)
	) name305 (
		_w1035_,
		_w1041_,
		_w1261_,
		_w1264_,
		_w1265_
	);
	LUT3 #(
		.INIT('h10)
	) name306 (
		_w1257_,
		_w1259_,
		_w1265_,
		_w1266_
	);
	LUT2 #(
		.INIT('h8)
	) name307 (
		_w1254_,
		_w1266_,
		_w1267_
	);
	LUT4 #(
		.INIT('h8000)
	) name308 (
		_w1113_,
		_w1164_,
		_w1226_,
		_w1267_,
		_w1268_
	);
	LUT3 #(
		.INIT('h20)
	) name309 (
		\u5_tmr_done_reg/NET0131 ,
		\u6_rmw_r_reg/NET0131 ,
		wb_cyc_i_pad,
		_w1269_
	);
	LUT4 #(
		.INIT('h7000)
	) name310 (
		_w1014_,
		_w1015_,
		_w1131_,
		_w1269_,
		_w1270_
	);
	LUT3 #(
		.INIT('h80)
	) name311 (
		_w1100_,
		_w1110_,
		_w1270_,
		_w1271_
	);
	LUT4 #(
		.INIT('h5554)
	) name312 (
		_w1129_,
		_w1141_,
		_w1145_,
		_w1271_,
		_w1272_
	);
	LUT4 #(
		.INIT('h0002)
	) name313 (
		\u5_state_reg[2]/NET0131 ,
		\u5_state_reg[3]/NET0131 ,
		\u5_state_reg[4]/NET0131 ,
		\u5_state_reg[5]/NET0131 ,
		_w1273_
	);
	LUT2 #(
		.INIT('h8)
	) name314 (
		_w982_,
		_w1273_,
		_w1274_
	);
	LUT3 #(
		.INIT('h80)
	) name315 (
		\u5_cmd_a10_r_reg/P0001 ,
		_w1002_,
		_w1274_,
		_w1275_
	);
	LUT4 #(
		.INIT('h0010)
	) name316 (
		\u5_state_reg[14]/NET0131 ,
		\u5_state_reg[15]/NET0131 ,
		\u5_state_reg[16]/NET0131 ,
		\u5_state_reg[17]/NET0131 ,
		_w1276_
	);
	LUT2 #(
		.INIT('h8)
	) name317 (
		_w981_,
		_w1276_,
		_w1277_
	);
	LUT3 #(
		.INIT('h2a)
	) name318 (
		\u5_tmr_done_reg/NET0131 ,
		_w976_,
		_w1118_,
		_w1278_
	);
	LUT2 #(
		.INIT('h4)
	) name319 (
		_w1117_,
		_w1278_,
		_w1279_
	);
	LUT3 #(
		.INIT('h8a)
	) name320 (
		\u5_cmd_a10_r_reg/P0001 ,
		_w1117_,
		_w1278_,
		_w1280_
	);
	LUT3 #(
		.INIT('h80)
	) name321 (
		_w1100_,
		_w1277_,
		_w1280_,
		_w1281_
	);
	LUT4 #(
		.INIT('h0002)
	) name322 (
		\u5_state_reg[18]/NET0131 ,
		\u5_state_reg[19]/NET0131 ,
		\u5_state_reg[20]/NET0131 ,
		\u5_state_reg[21]/NET0131 ,
		_w1282_
	);
	LUT3 #(
		.INIT('h80)
	) name323 (
		_w978_,
		_w984_,
		_w1282_,
		_w1283_
	);
	LUT4 #(
		.INIT('h0002)
	) name324 (
		\u5_state_reg[22]/NET0131 ,
		\u5_state_reg[23]/NET0131 ,
		\u5_state_reg[24]/NET0131 ,
		\u5_state_reg[25]/NET0131 ,
		_w1284_
	);
	LUT3 #(
		.INIT('h80)
	) name325 (
		_w984_,
		_w1046_,
		_w1284_,
		_w1285_
	);
	LUT3 #(
		.INIT('h57)
	) name326 (
		_w1035_,
		_w1283_,
		_w1285_,
		_w1286_
	);
	LUT4 #(
		.INIT('h0004)
	) name327 (
		\u5_state_reg[26]/NET0131 ,
		\u5_state_reg[27]/NET0131 ,
		\u5_state_reg[28]/NET0131 ,
		\u5_state_reg[29]/NET0131 ,
		_w1287_
	);
	LUT3 #(
		.INIT('h80)
	) name328 (
		_w978_,
		_w984_,
		_w1287_,
		_w1288_
	);
	LUT4 #(
		.INIT('h0010)
	) name329 (
		\u5_state_reg[2]/NET0131 ,
		\u5_state_reg[3]/NET0131 ,
		\u5_state_reg[4]/NET0131 ,
		\u5_state_reg[5]/NET0131 ,
		_w1289_
	);
	LUT2 #(
		.INIT('h8)
	) name330 (
		_w982_,
		_w1289_,
		_w1290_
	);
	LUT3 #(
		.INIT('h80)
	) name331 (
		\u5_rfr_ack_r_reg/NET0131 ,
		_w982_,
		_w1289_,
		_w1291_
	);
	LUT2 #(
		.INIT('h8)
	) name332 (
		_w1002_,
		_w1291_,
		_w1292_
	);
	LUT4 #(
		.INIT('h153f)
	) name333 (
		_w1002_,
		_w1068_,
		_w1288_,
		_w1291_,
		_w1293_
	);
	LUT4 #(
		.INIT('h1000)
	) name334 (
		_w1275_,
		_w1281_,
		_w1286_,
		_w1293_,
		_w1294_
	);
	LUT2 #(
		.INIT('h4)
	) name335 (
		_w1272_,
		_w1294_,
		_w1295_
	);
	LUT3 #(
		.INIT('h1f)
	) name336 (
		_w1138_,
		_w1268_,
		_w1295_,
		_w1296_
	);
	LUT4 #(
		.INIT('h02aa)
	) name337 (
		_w1034_,
		_w1138_,
		_w1268_,
		_w1295_,
		_w1297_
	);
	LUT4 #(
		.INIT('h0200)
	) name338 (
		_w1187_,
		_w1190_,
		_w1196_,
		_w1202_,
		_w1298_
	);
	LUT3 #(
		.INIT('h57)
	) name339 (
		_w1100_,
		_w1161_,
		_w1277_,
		_w1299_
	);
	LUT2 #(
		.INIT('h8)
	) name340 (
		_w1298_,
		_w1299_,
		_w1300_
	);
	LUT2 #(
		.INIT('h2)
	) name341 (
		\u5_wb_cycle_reg/NET0131 ,
		_w1116_,
		_w1301_
	);
	LUT4 #(
		.INIT('h8000)
	) name342 (
		\u5_wb_cycle_reg/NET0131 ,
		_w1122_,
		_w1124_,
		_w1127_,
		_w1302_
	);
	LUT2 #(
		.INIT('h1)
	) name343 (
		_w1301_,
		_w1302_,
		_w1303_
	);
	LUT4 #(
		.INIT('h0008)
	) name344 (
		_w1100_,
		_w1140_,
		_w1301_,
		_w1302_,
		_w1304_
	);
	LUT2 #(
		.INIT('h8)
	) name345 (
		_w1002_,
		_w1290_,
		_w1305_
	);
	LUT4 #(
		.INIT('h153f)
	) name346 (
		_w1002_,
		_w1068_,
		_w1288_,
		_w1290_,
		_w1306_
	);
	LUT3 #(
		.INIT('h10)
	) name347 (
		_w1169_,
		_w1304_,
		_w1306_,
		_w1307_
	);
	LUT4 #(
		.INIT('h153f)
	) name348 (
		_w1041_,
		_w1100_,
		_w1158_,
		_w1217_,
		_w1308_
	);
	LUT3 #(
		.INIT('h10)
	) name349 (
		_w1259_,
		_w1262_,
		_w1308_,
		_w1309_
	);
	LUT2 #(
		.INIT('h8)
	) name350 (
		_w1208_,
		_w1215_,
		_w1310_
	);
	LUT4 #(
		.INIT('h8000)
	) name351 (
		_w1053_,
		_w1307_,
		_w1309_,
		_w1310_,
		_w1311_
	);
	LUT4 #(
		.INIT('h153f)
	) name352 (
		_w1041_,
		_w1100_,
		_w1108_,
		_w1152_,
		_w1312_
	);
	LUT2 #(
		.INIT('h4)
	) name353 (
		_w1150_,
		_w1312_,
		_w1313_
	);
	LUT4 #(
		.INIT('h135f)
	) name354 (
		_w1041_,
		_w1059_,
		_w1091_,
		_w1172_,
		_w1314_
	);
	LUT4 #(
		.INIT('h135f)
	) name355 (
		_w991_,
		_w1002_,
		_w1094_,
		_w1166_,
		_w1315_
	);
	LUT4 #(
		.INIT('h4000)
	) name356 (
		_w1150_,
		_w1312_,
		_w1314_,
		_w1315_,
		_w1316_
	);
	LUT3 #(
		.INIT('h80)
	) name357 (
		_w1057_,
		_w1066_,
		_w1286_,
		_w1317_
	);
	LUT2 #(
		.INIT('h8)
	) name358 (
		_w1316_,
		_w1317_,
		_w1318_
	);
	LUT4 #(
		.INIT('h153f)
	) name359 (
		_w1063_,
		_w1100_,
		_w1110_,
		_w1221_,
		_w1319_
	);
	LUT4 #(
		.INIT('h153f)
	) name360 (
		_w1002_,
		_w1059_,
		_w1223_,
		_w1274_,
		_w1320_
	);
	LUT4 #(
		.INIT('h0777)
	) name361 (
		_w1035_,
		_w1097_,
		_w1174_,
		_w1178_,
		_w1321_
	);
	LUT3 #(
		.INIT('h80)
	) name362 (
		_w1319_,
		_w1320_,
		_w1321_,
		_w1322_
	);
	LUT4 #(
		.INIT('h0800)
	) name363 (
		_w1089_,
		_w1254_,
		_w1257_,
		_w1322_,
		_w1323_
	);
	LUT4 #(
		.INIT('h8000)
	) name364 (
		_w1300_,
		_w1311_,
		_w1318_,
		_w1323_,
		_w1324_
	);
	LUT4 #(
		.INIT('h7fff)
	) name365 (
		_w1300_,
		_w1311_,
		_w1318_,
		_w1323_,
		_w1325_
	);
	LUT2 #(
		.INIT('h8)
	) name366 (
		\u5_cmd_del_reg[1]/NET0131 ,
		\u5_wr_cycle_reg/NET0131 ,
		_w1326_
	);
	LUT3 #(
		.INIT('h07)
	) name367 (
		_w976_,
		_w1114_,
		_w1326_,
		_w1327_
	);
	LUT3 #(
		.INIT('h08)
	) name368 (
		\u1_row_adr_reg[10]/P0001 ,
		\u5_state_reg[6]/NET0131 ,
		\u5_wb_wait_r_reg/P0001 ,
		_w1328_
	);
	LUT3 #(
		.INIT('h80)
	) name369 (
		\u1_row_adr_reg[10]/P0001 ,
		_w966_,
		_w1018_,
		_w1329_
	);
	LUT3 #(
		.INIT('h13)
	) name370 (
		_w1033_,
		_w1328_,
		_w1329_,
		_w1330_
	);
	LUT4 #(
		.INIT('h1f00)
	) name371 (
		\u5_wr_cycle_reg/NET0131 ,
		_w1324_,
		_w1327_,
		_w1330_,
		_w1331_
	);
	LUT3 #(
		.INIT('h02)
	) name372 (
		\u0_csc_reg[1]/NET0131 ,
		\u5_lmr_ack_reg/NET0131 ,
		\u5_state_reg[26]/NET0131 ,
		_w1332_
	);
	LUT4 #(
		.INIT('h11d5)
	) name373 (
		\u0_sp_csc_reg[1]/NET0131 ,
		_w976_,
		_w1114_,
		_w1332_,
		_w1333_
	);
	LUT3 #(
		.INIT('h02)
	) name374 (
		\u0_csc_reg[3]/NET0131 ,
		\u5_lmr_ack_reg/NET0131 ,
		\u5_state_reg[26]/NET0131 ,
		_w1334_
	);
	LUT4 #(
		.INIT('h11d5)
	) name375 (
		\u0_sp_csc_reg[3]/NET0131 ,
		_w976_,
		_w1114_,
		_w1334_,
		_w1335_
	);
	LUT2 #(
		.INIT('h8)
	) name376 (
		_w1333_,
		_w1335_,
		_w1336_
	);
	LUT3 #(
		.INIT('h02)
	) name377 (
		\u0_csc_reg[2]/NET0131 ,
		\u5_lmr_ack_reg/NET0131 ,
		\u5_state_reg[26]/NET0131 ,
		_w1337_
	);
	LUT4 #(
		.INIT('h11d5)
	) name378 (
		\u0_sp_csc_reg[2]/NET0131 ,
		_w976_,
		_w1114_,
		_w1337_,
		_w1338_
	);
	LUT3 #(
		.INIT('h80)
	) name379 (
		_w1333_,
		_w1335_,
		_w1338_,
		_w1339_
	);
	LUT3 #(
		.INIT('h15)
	) name380 (
		\u0_sp_tms_reg[10]/NET0131 ,
		\u5_cmd_del_reg[1]/NET0131 ,
		\u5_wr_cycle_reg/NET0131 ,
		_w1340_
	);
	LUT3 #(
		.INIT('h70)
	) name381 (
		_w976_,
		_w1114_,
		_w1340_,
		_w1341_
	);
	LUT4 #(
		.INIT('h10f0)
	) name382 (
		\u5_wr_cycle_reg/NET0131 ,
		_w1324_,
		_w1339_,
		_w1341_,
		_w1342_
	);
	LUT2 #(
		.INIT('h4)
	) name383 (
		_w1333_,
		_w1335_,
		_w1343_
	);
	LUT4 #(
		.INIT('h2000)
	) name384 (
		\u6_wr_hold_reg/NET0131 ,
		_w1333_,
		_w1335_,
		_w1338_,
		_w1344_
	);
	LUT2 #(
		.INIT('h4)
	) name385 (
		\u1_sram_addr_reg[10]/P0001 ,
		\u6_wr_hold_reg/NET0131 ,
		_w1345_
	);
	LUT4 #(
		.INIT('h3777)
	) name386 (
		_w1333_,
		_w1335_,
		_w1338_,
		_w1345_,
		_w1346_
	);
	LUT3 #(
		.INIT('he0)
	) name387 (
		\wb_addr_i[12]_pad ,
		_w1344_,
		_w1346_,
		_w1347_
	);
	LUT4 #(
		.INIT('h0080)
	) name388 (
		\u1_acs_addr_reg[10]/P0001 ,
		_w1333_,
		_w1335_,
		_w1338_,
		_w1348_
	);
	LUT2 #(
		.INIT('h1)
	) name389 (
		\u5_rfr_ack_r_reg/NET0131 ,
		_w1348_,
		_w1349_
	);
	LUT2 #(
		.INIT('h4)
	) name390 (
		_w1347_,
		_w1349_,
		_w1350_
	);
	LUT4 #(
		.INIT('hb0ff)
	) name391 (
		_w1297_,
		_w1331_,
		_w1342_,
		_w1350_,
		_w1351_
	);
	LUT3 #(
		.INIT('h51)
	) name392 (
		\u1_col_adr_reg[0]/P0001 ,
		\u5_state_reg[6]/NET0131 ,
		\u5_wb_wait_r_reg/P0001 ,
		_w1352_
	);
	LUT3 #(
		.INIT('h70)
	) name393 (
		_w1019_,
		_w1033_,
		_w1352_,
		_w1353_
	);
	LUT3 #(
		.INIT('h04)
	) name394 (
		\u1_row_adr_reg[0]/P0001 ,
		\u5_state_reg[6]/NET0131 ,
		\u5_wb_wait_r_reg/P0001 ,
		_w1354_
	);
	LUT3 #(
		.INIT('h40)
	) name395 (
		\u1_row_adr_reg[0]/P0001 ,
		_w966_,
		_w1018_,
		_w1355_
	);
	LUT3 #(
		.INIT('h13)
	) name396 (
		_w1033_,
		_w1354_,
		_w1355_,
		_w1356_
	);
	LUT2 #(
		.INIT('h4)
	) name397 (
		_w1353_,
		_w1356_,
		_w1357_
	);
	LUT4 #(
		.INIT('h001f)
	) name398 (
		\u5_wr_cycle_reg/NET0131 ,
		_w1324_,
		_w1327_,
		_w1357_,
		_w1358_
	);
	LUT3 #(
		.INIT('h15)
	) name399 (
		\u0_sp_tms_reg[0]/NET0131 ,
		\u5_cmd_del_reg[1]/NET0131 ,
		\u5_wr_cycle_reg/NET0131 ,
		_w1359_
	);
	LUT3 #(
		.INIT('h70)
	) name400 (
		_w976_,
		_w1114_,
		_w1359_,
		_w1360_
	);
	LUT4 #(
		.INIT('h10f0)
	) name401 (
		\u5_wr_cycle_reg/NET0131 ,
		_w1324_,
		_w1339_,
		_w1360_,
		_w1361_
	);
	LUT4 #(
		.INIT('h0080)
	) name402 (
		\u1_acs_addr_reg[0]/P0001 ,
		_w1333_,
		_w1335_,
		_w1338_,
		_w1362_
	);
	LUT2 #(
		.INIT('h4)
	) name403 (
		\u1_sram_addr_reg[0]/P0001 ,
		\u6_wr_hold_reg/NET0131 ,
		_w1363_
	);
	LUT4 #(
		.INIT('h3777)
	) name404 (
		_w1333_,
		_w1335_,
		_w1338_,
		_w1363_,
		_w1364_
	);
	LUT4 #(
		.INIT('h010f)
	) name405 (
		\wb_addr_i[2]_pad ,
		_w1344_,
		_w1362_,
		_w1364_,
		_w1365_
	);
	LUT3 #(
		.INIT('h4f)
	) name406 (
		_w1358_,
		_w1361_,
		_w1365_,
		_w1366_
	);
	LUT3 #(
		.INIT('h08)
	) name407 (
		\u1_row_adr_reg[11]/P0001 ,
		\u5_state_reg[6]/NET0131 ,
		\u5_wb_wait_r_reg/P0001 ,
		_w1367_
	);
	LUT3 #(
		.INIT('h80)
	) name408 (
		\u1_row_adr_reg[11]/P0001 ,
		_w966_,
		_w1018_,
		_w1368_
	);
	LUT3 #(
		.INIT('h13)
	) name409 (
		_w1033_,
		_w1367_,
		_w1368_,
		_w1369_
	);
	LUT4 #(
		.INIT('h1f00)
	) name410 (
		\u5_wr_cycle_reg/NET0131 ,
		_w1324_,
		_w1327_,
		_w1369_,
		_w1370_
	);
	LUT3 #(
		.INIT('h15)
	) name411 (
		\u0_sp_tms_reg[11]/NET0131 ,
		\u5_cmd_del_reg[1]/NET0131 ,
		\u5_wr_cycle_reg/NET0131 ,
		_w1371_
	);
	LUT3 #(
		.INIT('h70)
	) name412 (
		_w976_,
		_w1114_,
		_w1371_,
		_w1372_
	);
	LUT4 #(
		.INIT('h10f0)
	) name413 (
		\u5_wr_cycle_reg/NET0131 ,
		_w1324_,
		_w1339_,
		_w1372_,
		_w1373_
	);
	LUT4 #(
		.INIT('h0080)
	) name414 (
		\u1_acs_addr_reg[11]/P0001 ,
		_w1333_,
		_w1335_,
		_w1338_,
		_w1374_
	);
	LUT2 #(
		.INIT('h4)
	) name415 (
		\u1_sram_addr_reg[11]/P0001 ,
		\u6_wr_hold_reg/NET0131 ,
		_w1375_
	);
	LUT4 #(
		.INIT('h3777)
	) name416 (
		_w1333_,
		_w1335_,
		_w1338_,
		_w1375_,
		_w1376_
	);
	LUT4 #(
		.INIT('h010f)
	) name417 (
		\wb_addr_i[13]_pad ,
		_w1344_,
		_w1374_,
		_w1376_,
		_w1377_
	);
	LUT3 #(
		.INIT('h4f)
	) name418 (
		_w1370_,
		_w1373_,
		_w1377_,
		_w1378_
	);
	LUT3 #(
		.INIT('h08)
	) name419 (
		\u1_row_adr_reg[12]/P0001 ,
		\u5_state_reg[6]/NET0131 ,
		\u5_wb_wait_r_reg/P0001 ,
		_w1379_
	);
	LUT3 #(
		.INIT('h80)
	) name420 (
		\u1_row_adr_reg[12]/P0001 ,
		_w966_,
		_w1018_,
		_w1380_
	);
	LUT3 #(
		.INIT('h13)
	) name421 (
		_w1033_,
		_w1379_,
		_w1380_,
		_w1381_
	);
	LUT4 #(
		.INIT('h1f00)
	) name422 (
		\u5_wr_cycle_reg/NET0131 ,
		_w1324_,
		_w1327_,
		_w1381_,
		_w1382_
	);
	LUT3 #(
		.INIT('h15)
	) name423 (
		\u0_sp_tms_reg[12]/NET0131 ,
		\u5_cmd_del_reg[1]/NET0131 ,
		\u5_wr_cycle_reg/NET0131 ,
		_w1383_
	);
	LUT3 #(
		.INIT('h70)
	) name424 (
		_w976_,
		_w1114_,
		_w1383_,
		_w1384_
	);
	LUT4 #(
		.INIT('h10f0)
	) name425 (
		\u5_wr_cycle_reg/NET0131 ,
		_w1324_,
		_w1339_,
		_w1384_,
		_w1385_
	);
	LUT4 #(
		.INIT('h0080)
	) name426 (
		\u1_acs_addr_reg[12]/P0001 ,
		_w1333_,
		_w1335_,
		_w1338_,
		_w1386_
	);
	LUT2 #(
		.INIT('h4)
	) name427 (
		\u1_sram_addr_reg[12]/P0001 ,
		\u6_wr_hold_reg/NET0131 ,
		_w1387_
	);
	LUT4 #(
		.INIT('h3777)
	) name428 (
		_w1333_,
		_w1335_,
		_w1338_,
		_w1387_,
		_w1388_
	);
	LUT4 #(
		.INIT('h010f)
	) name429 (
		\wb_addr_i[14]_pad ,
		_w1344_,
		_w1386_,
		_w1388_,
		_w1389_
	);
	LUT3 #(
		.INIT('h4f)
	) name430 (
		_w1382_,
		_w1385_,
		_w1389_,
		_w1390_
	);
	LUT3 #(
		.INIT('h51)
	) name431 (
		\u1_col_adr_reg[1]/P0001 ,
		\u5_state_reg[6]/NET0131 ,
		\u5_wb_wait_r_reg/P0001 ,
		_w1391_
	);
	LUT3 #(
		.INIT('h70)
	) name432 (
		_w1019_,
		_w1033_,
		_w1391_,
		_w1392_
	);
	LUT3 #(
		.INIT('h04)
	) name433 (
		\u1_row_adr_reg[1]/P0001 ,
		\u5_state_reg[6]/NET0131 ,
		\u5_wb_wait_r_reg/P0001 ,
		_w1393_
	);
	LUT3 #(
		.INIT('h40)
	) name434 (
		\u1_row_adr_reg[1]/P0001 ,
		_w966_,
		_w1018_,
		_w1394_
	);
	LUT3 #(
		.INIT('h13)
	) name435 (
		_w1033_,
		_w1393_,
		_w1394_,
		_w1395_
	);
	LUT2 #(
		.INIT('h4)
	) name436 (
		_w1392_,
		_w1395_,
		_w1396_
	);
	LUT4 #(
		.INIT('h001f)
	) name437 (
		\u5_wr_cycle_reg/NET0131 ,
		_w1324_,
		_w1327_,
		_w1396_,
		_w1397_
	);
	LUT3 #(
		.INIT('h15)
	) name438 (
		\u0_sp_tms_reg[1]/NET0131 ,
		\u5_cmd_del_reg[1]/NET0131 ,
		\u5_wr_cycle_reg/NET0131 ,
		_w1398_
	);
	LUT3 #(
		.INIT('h70)
	) name439 (
		_w976_,
		_w1114_,
		_w1398_,
		_w1399_
	);
	LUT4 #(
		.INIT('h10f0)
	) name440 (
		\u5_wr_cycle_reg/NET0131 ,
		_w1324_,
		_w1339_,
		_w1399_,
		_w1400_
	);
	LUT4 #(
		.INIT('h0080)
	) name441 (
		\u1_acs_addr_reg[1]/P0001 ,
		_w1333_,
		_w1335_,
		_w1338_,
		_w1401_
	);
	LUT2 #(
		.INIT('h4)
	) name442 (
		\u1_sram_addr_reg[1]/P0001 ,
		\u6_wr_hold_reg/NET0131 ,
		_w1402_
	);
	LUT4 #(
		.INIT('h3777)
	) name443 (
		_w1333_,
		_w1335_,
		_w1338_,
		_w1402_,
		_w1403_
	);
	LUT4 #(
		.INIT('h010f)
	) name444 (
		\wb_addr_i[3]_pad ,
		_w1344_,
		_w1401_,
		_w1403_,
		_w1404_
	);
	LUT3 #(
		.INIT('h4f)
	) name445 (
		_w1397_,
		_w1400_,
		_w1404_,
		_w1405_
	);
	LUT3 #(
		.INIT('h51)
	) name446 (
		\u1_col_adr_reg[2]/P0001 ,
		\u5_state_reg[6]/NET0131 ,
		\u5_wb_wait_r_reg/P0001 ,
		_w1406_
	);
	LUT3 #(
		.INIT('h70)
	) name447 (
		_w1019_,
		_w1033_,
		_w1406_,
		_w1407_
	);
	LUT3 #(
		.INIT('h04)
	) name448 (
		\u1_row_adr_reg[2]/P0001 ,
		\u5_state_reg[6]/NET0131 ,
		\u5_wb_wait_r_reg/P0001 ,
		_w1408_
	);
	LUT3 #(
		.INIT('h40)
	) name449 (
		\u1_row_adr_reg[2]/P0001 ,
		_w966_,
		_w1018_,
		_w1409_
	);
	LUT3 #(
		.INIT('h13)
	) name450 (
		_w1033_,
		_w1408_,
		_w1409_,
		_w1410_
	);
	LUT2 #(
		.INIT('h4)
	) name451 (
		_w1407_,
		_w1410_,
		_w1411_
	);
	LUT4 #(
		.INIT('h001f)
	) name452 (
		\u5_wr_cycle_reg/NET0131 ,
		_w1324_,
		_w1327_,
		_w1411_,
		_w1412_
	);
	LUT3 #(
		.INIT('h15)
	) name453 (
		\u0_sp_tms_reg[2]/NET0131 ,
		\u5_cmd_del_reg[1]/NET0131 ,
		\u5_wr_cycle_reg/NET0131 ,
		_w1413_
	);
	LUT3 #(
		.INIT('h70)
	) name454 (
		_w976_,
		_w1114_,
		_w1413_,
		_w1414_
	);
	LUT4 #(
		.INIT('h10f0)
	) name455 (
		\u5_wr_cycle_reg/NET0131 ,
		_w1324_,
		_w1339_,
		_w1414_,
		_w1415_
	);
	LUT4 #(
		.INIT('h0080)
	) name456 (
		\u1_acs_addr_reg[2]/P0001 ,
		_w1333_,
		_w1335_,
		_w1338_,
		_w1416_
	);
	LUT2 #(
		.INIT('h4)
	) name457 (
		\u1_sram_addr_reg[2]/P0001 ,
		\u6_wr_hold_reg/NET0131 ,
		_w1417_
	);
	LUT4 #(
		.INIT('h3777)
	) name458 (
		_w1333_,
		_w1335_,
		_w1338_,
		_w1417_,
		_w1418_
	);
	LUT4 #(
		.INIT('h010f)
	) name459 (
		\wb_addr_i[4]_pad ,
		_w1344_,
		_w1416_,
		_w1418_,
		_w1419_
	);
	LUT3 #(
		.INIT('h4f)
	) name460 (
		_w1412_,
		_w1415_,
		_w1419_,
		_w1420_
	);
	LUT3 #(
		.INIT('h51)
	) name461 (
		\u1_col_adr_reg[3]/P0001 ,
		\u5_state_reg[6]/NET0131 ,
		\u5_wb_wait_r_reg/P0001 ,
		_w1421_
	);
	LUT3 #(
		.INIT('h70)
	) name462 (
		_w1019_,
		_w1033_,
		_w1421_,
		_w1422_
	);
	LUT3 #(
		.INIT('h04)
	) name463 (
		\u1_row_adr_reg[3]/P0001 ,
		\u5_state_reg[6]/NET0131 ,
		\u5_wb_wait_r_reg/P0001 ,
		_w1423_
	);
	LUT3 #(
		.INIT('h40)
	) name464 (
		\u1_row_adr_reg[3]/P0001 ,
		_w966_,
		_w1018_,
		_w1424_
	);
	LUT3 #(
		.INIT('h13)
	) name465 (
		_w1033_,
		_w1423_,
		_w1424_,
		_w1425_
	);
	LUT2 #(
		.INIT('h4)
	) name466 (
		_w1422_,
		_w1425_,
		_w1426_
	);
	LUT4 #(
		.INIT('h001f)
	) name467 (
		\u5_wr_cycle_reg/NET0131 ,
		_w1324_,
		_w1327_,
		_w1426_,
		_w1427_
	);
	LUT3 #(
		.INIT('h15)
	) name468 (
		\u0_sp_tms_reg[3]/NET0131 ,
		\u5_cmd_del_reg[1]/NET0131 ,
		\u5_wr_cycle_reg/NET0131 ,
		_w1428_
	);
	LUT3 #(
		.INIT('h70)
	) name469 (
		_w976_,
		_w1114_,
		_w1428_,
		_w1429_
	);
	LUT4 #(
		.INIT('h10f0)
	) name470 (
		\u5_wr_cycle_reg/NET0131 ,
		_w1324_,
		_w1339_,
		_w1429_,
		_w1430_
	);
	LUT4 #(
		.INIT('h0080)
	) name471 (
		\u1_acs_addr_reg[3]/P0001 ,
		_w1333_,
		_w1335_,
		_w1338_,
		_w1431_
	);
	LUT2 #(
		.INIT('h4)
	) name472 (
		\u1_sram_addr_reg[3]/P0001 ,
		\u6_wr_hold_reg/NET0131 ,
		_w1432_
	);
	LUT4 #(
		.INIT('h3777)
	) name473 (
		_w1333_,
		_w1335_,
		_w1338_,
		_w1432_,
		_w1433_
	);
	LUT4 #(
		.INIT('h010f)
	) name474 (
		\wb_addr_i[5]_pad ,
		_w1344_,
		_w1431_,
		_w1433_,
		_w1434_
	);
	LUT3 #(
		.INIT('h4f)
	) name475 (
		_w1427_,
		_w1430_,
		_w1434_,
		_w1435_
	);
	LUT3 #(
		.INIT('h51)
	) name476 (
		\u1_col_adr_reg[4]/P0001 ,
		\u5_state_reg[6]/NET0131 ,
		\u5_wb_wait_r_reg/P0001 ,
		_w1436_
	);
	LUT3 #(
		.INIT('h70)
	) name477 (
		_w1019_,
		_w1033_,
		_w1436_,
		_w1437_
	);
	LUT3 #(
		.INIT('h04)
	) name478 (
		\u1_row_adr_reg[4]/P0001 ,
		\u5_state_reg[6]/NET0131 ,
		\u5_wb_wait_r_reg/P0001 ,
		_w1438_
	);
	LUT3 #(
		.INIT('h40)
	) name479 (
		\u1_row_adr_reg[4]/P0001 ,
		_w966_,
		_w1018_,
		_w1439_
	);
	LUT3 #(
		.INIT('h13)
	) name480 (
		_w1033_,
		_w1438_,
		_w1439_,
		_w1440_
	);
	LUT2 #(
		.INIT('h4)
	) name481 (
		_w1437_,
		_w1440_,
		_w1441_
	);
	LUT4 #(
		.INIT('h001f)
	) name482 (
		\u5_wr_cycle_reg/NET0131 ,
		_w1324_,
		_w1327_,
		_w1441_,
		_w1442_
	);
	LUT3 #(
		.INIT('h15)
	) name483 (
		\u0_sp_tms_reg[4]/NET0131 ,
		\u5_cmd_del_reg[1]/NET0131 ,
		\u5_wr_cycle_reg/NET0131 ,
		_w1443_
	);
	LUT3 #(
		.INIT('h70)
	) name484 (
		_w976_,
		_w1114_,
		_w1443_,
		_w1444_
	);
	LUT4 #(
		.INIT('h10f0)
	) name485 (
		\u5_wr_cycle_reg/NET0131 ,
		_w1324_,
		_w1339_,
		_w1444_,
		_w1445_
	);
	LUT4 #(
		.INIT('h0080)
	) name486 (
		\u1_acs_addr_reg[4]/P0001 ,
		_w1333_,
		_w1335_,
		_w1338_,
		_w1446_
	);
	LUT2 #(
		.INIT('h4)
	) name487 (
		\u1_sram_addr_reg[4]/P0001 ,
		\u6_wr_hold_reg/NET0131 ,
		_w1447_
	);
	LUT4 #(
		.INIT('h3777)
	) name488 (
		_w1333_,
		_w1335_,
		_w1338_,
		_w1447_,
		_w1448_
	);
	LUT4 #(
		.INIT('h010f)
	) name489 (
		\wb_addr_i[6]_pad ,
		_w1344_,
		_w1446_,
		_w1448_,
		_w1449_
	);
	LUT3 #(
		.INIT('h4f)
	) name490 (
		_w1442_,
		_w1445_,
		_w1449_,
		_w1450_
	);
	LUT3 #(
		.INIT('h51)
	) name491 (
		\u1_col_adr_reg[5]/P0001 ,
		\u5_state_reg[6]/NET0131 ,
		\u5_wb_wait_r_reg/P0001 ,
		_w1451_
	);
	LUT3 #(
		.INIT('h70)
	) name492 (
		_w1019_,
		_w1033_,
		_w1451_,
		_w1452_
	);
	LUT3 #(
		.INIT('h04)
	) name493 (
		\u1_row_adr_reg[5]/P0001 ,
		\u5_state_reg[6]/NET0131 ,
		\u5_wb_wait_r_reg/P0001 ,
		_w1453_
	);
	LUT3 #(
		.INIT('h40)
	) name494 (
		\u1_row_adr_reg[5]/P0001 ,
		_w966_,
		_w1018_,
		_w1454_
	);
	LUT3 #(
		.INIT('h13)
	) name495 (
		_w1033_,
		_w1453_,
		_w1454_,
		_w1455_
	);
	LUT2 #(
		.INIT('h4)
	) name496 (
		_w1452_,
		_w1455_,
		_w1456_
	);
	LUT4 #(
		.INIT('h001f)
	) name497 (
		\u5_wr_cycle_reg/NET0131 ,
		_w1324_,
		_w1327_,
		_w1456_,
		_w1457_
	);
	LUT3 #(
		.INIT('h15)
	) name498 (
		\u0_sp_tms_reg[5]/NET0131 ,
		\u5_cmd_del_reg[1]/NET0131 ,
		\u5_wr_cycle_reg/NET0131 ,
		_w1458_
	);
	LUT3 #(
		.INIT('h70)
	) name499 (
		_w976_,
		_w1114_,
		_w1458_,
		_w1459_
	);
	LUT4 #(
		.INIT('h10f0)
	) name500 (
		\u5_wr_cycle_reg/NET0131 ,
		_w1324_,
		_w1339_,
		_w1459_,
		_w1460_
	);
	LUT4 #(
		.INIT('h0080)
	) name501 (
		\u1_acs_addr_reg[5]/P0001 ,
		_w1333_,
		_w1335_,
		_w1338_,
		_w1461_
	);
	LUT2 #(
		.INIT('h4)
	) name502 (
		\u1_sram_addr_reg[5]/P0001 ,
		\u6_wr_hold_reg/NET0131 ,
		_w1462_
	);
	LUT4 #(
		.INIT('h3777)
	) name503 (
		_w1333_,
		_w1335_,
		_w1338_,
		_w1462_,
		_w1463_
	);
	LUT4 #(
		.INIT('h010f)
	) name504 (
		\wb_addr_i[7]_pad ,
		_w1344_,
		_w1461_,
		_w1463_,
		_w1464_
	);
	LUT3 #(
		.INIT('h4f)
	) name505 (
		_w1457_,
		_w1460_,
		_w1464_,
		_w1465_
	);
	LUT3 #(
		.INIT('h51)
	) name506 (
		\u1_col_adr_reg[6]/P0001 ,
		\u5_state_reg[6]/NET0131 ,
		\u5_wb_wait_r_reg/P0001 ,
		_w1466_
	);
	LUT3 #(
		.INIT('h70)
	) name507 (
		_w1019_,
		_w1033_,
		_w1466_,
		_w1467_
	);
	LUT3 #(
		.INIT('h04)
	) name508 (
		\u1_row_adr_reg[6]/P0001 ,
		\u5_state_reg[6]/NET0131 ,
		\u5_wb_wait_r_reg/P0001 ,
		_w1468_
	);
	LUT3 #(
		.INIT('h40)
	) name509 (
		\u1_row_adr_reg[6]/P0001 ,
		_w966_,
		_w1018_,
		_w1469_
	);
	LUT3 #(
		.INIT('h13)
	) name510 (
		_w1033_,
		_w1468_,
		_w1469_,
		_w1470_
	);
	LUT2 #(
		.INIT('h4)
	) name511 (
		_w1467_,
		_w1470_,
		_w1471_
	);
	LUT4 #(
		.INIT('h001f)
	) name512 (
		\u5_wr_cycle_reg/NET0131 ,
		_w1324_,
		_w1327_,
		_w1471_,
		_w1472_
	);
	LUT3 #(
		.INIT('h15)
	) name513 (
		\u0_sp_tms_reg[6]/NET0131 ,
		\u5_cmd_del_reg[1]/NET0131 ,
		\u5_wr_cycle_reg/NET0131 ,
		_w1473_
	);
	LUT3 #(
		.INIT('h70)
	) name514 (
		_w976_,
		_w1114_,
		_w1473_,
		_w1474_
	);
	LUT4 #(
		.INIT('h10f0)
	) name515 (
		\u5_wr_cycle_reg/NET0131 ,
		_w1324_,
		_w1339_,
		_w1474_,
		_w1475_
	);
	LUT4 #(
		.INIT('h0080)
	) name516 (
		\u1_acs_addr_reg[6]/P0001 ,
		_w1333_,
		_w1335_,
		_w1338_,
		_w1476_
	);
	LUT2 #(
		.INIT('h4)
	) name517 (
		\u1_sram_addr_reg[6]/P0001 ,
		\u6_wr_hold_reg/NET0131 ,
		_w1477_
	);
	LUT4 #(
		.INIT('h3777)
	) name518 (
		_w1333_,
		_w1335_,
		_w1338_,
		_w1477_,
		_w1478_
	);
	LUT4 #(
		.INIT('h010f)
	) name519 (
		\wb_addr_i[8]_pad ,
		_w1344_,
		_w1476_,
		_w1478_,
		_w1479_
	);
	LUT3 #(
		.INIT('h4f)
	) name520 (
		_w1472_,
		_w1475_,
		_w1479_,
		_w1480_
	);
	LUT3 #(
		.INIT('h51)
	) name521 (
		\u1_col_adr_reg[7]/P0001 ,
		\u5_state_reg[6]/NET0131 ,
		\u5_wb_wait_r_reg/P0001 ,
		_w1481_
	);
	LUT3 #(
		.INIT('h70)
	) name522 (
		_w1019_,
		_w1033_,
		_w1481_,
		_w1482_
	);
	LUT3 #(
		.INIT('h04)
	) name523 (
		\u1_row_adr_reg[7]/P0001 ,
		\u5_state_reg[6]/NET0131 ,
		\u5_wb_wait_r_reg/P0001 ,
		_w1483_
	);
	LUT3 #(
		.INIT('h40)
	) name524 (
		\u1_row_adr_reg[7]/P0001 ,
		_w966_,
		_w1018_,
		_w1484_
	);
	LUT3 #(
		.INIT('h13)
	) name525 (
		_w1033_,
		_w1483_,
		_w1484_,
		_w1485_
	);
	LUT2 #(
		.INIT('h4)
	) name526 (
		_w1482_,
		_w1485_,
		_w1486_
	);
	LUT4 #(
		.INIT('h001f)
	) name527 (
		\u5_wr_cycle_reg/NET0131 ,
		_w1324_,
		_w1327_,
		_w1486_,
		_w1487_
	);
	LUT3 #(
		.INIT('h15)
	) name528 (
		\u0_sp_tms_reg[7]/NET0131 ,
		\u5_cmd_del_reg[1]/NET0131 ,
		\u5_wr_cycle_reg/NET0131 ,
		_w1488_
	);
	LUT3 #(
		.INIT('h70)
	) name529 (
		_w976_,
		_w1114_,
		_w1488_,
		_w1489_
	);
	LUT4 #(
		.INIT('h10f0)
	) name530 (
		\u5_wr_cycle_reg/NET0131 ,
		_w1324_,
		_w1339_,
		_w1489_,
		_w1490_
	);
	LUT4 #(
		.INIT('h0080)
	) name531 (
		\u1_acs_addr_reg[7]/P0001 ,
		_w1333_,
		_w1335_,
		_w1338_,
		_w1491_
	);
	LUT2 #(
		.INIT('h4)
	) name532 (
		\u1_sram_addr_reg[7]/P0001 ,
		\u6_wr_hold_reg/NET0131 ,
		_w1492_
	);
	LUT4 #(
		.INIT('h3777)
	) name533 (
		_w1333_,
		_w1335_,
		_w1338_,
		_w1492_,
		_w1493_
	);
	LUT4 #(
		.INIT('h010f)
	) name534 (
		\wb_addr_i[9]_pad ,
		_w1344_,
		_w1491_,
		_w1493_,
		_w1494_
	);
	LUT3 #(
		.INIT('h4f)
	) name535 (
		_w1487_,
		_w1490_,
		_w1494_,
		_w1495_
	);
	LUT3 #(
		.INIT('h51)
	) name536 (
		\u1_col_adr_reg[8]/P0001 ,
		\u5_state_reg[6]/NET0131 ,
		\u5_wb_wait_r_reg/P0001 ,
		_w1496_
	);
	LUT3 #(
		.INIT('h70)
	) name537 (
		_w1019_,
		_w1033_,
		_w1496_,
		_w1497_
	);
	LUT3 #(
		.INIT('h04)
	) name538 (
		\u1_row_adr_reg[8]/P0001 ,
		\u5_state_reg[6]/NET0131 ,
		\u5_wb_wait_r_reg/P0001 ,
		_w1498_
	);
	LUT3 #(
		.INIT('h40)
	) name539 (
		\u1_row_adr_reg[8]/P0001 ,
		_w966_,
		_w1018_,
		_w1499_
	);
	LUT3 #(
		.INIT('h13)
	) name540 (
		_w1033_,
		_w1498_,
		_w1499_,
		_w1500_
	);
	LUT2 #(
		.INIT('h4)
	) name541 (
		_w1497_,
		_w1500_,
		_w1501_
	);
	LUT4 #(
		.INIT('h001f)
	) name542 (
		\u5_wr_cycle_reg/NET0131 ,
		_w1324_,
		_w1327_,
		_w1501_,
		_w1502_
	);
	LUT3 #(
		.INIT('h15)
	) name543 (
		\u0_sp_tms_reg[8]/NET0131 ,
		\u5_cmd_del_reg[1]/NET0131 ,
		\u5_wr_cycle_reg/NET0131 ,
		_w1503_
	);
	LUT3 #(
		.INIT('h70)
	) name544 (
		_w976_,
		_w1114_,
		_w1503_,
		_w1504_
	);
	LUT4 #(
		.INIT('h10f0)
	) name545 (
		\u5_wr_cycle_reg/NET0131 ,
		_w1324_,
		_w1339_,
		_w1504_,
		_w1505_
	);
	LUT4 #(
		.INIT('h0080)
	) name546 (
		\u1_acs_addr_reg[8]/P0001 ,
		_w1333_,
		_w1335_,
		_w1338_,
		_w1506_
	);
	LUT2 #(
		.INIT('h4)
	) name547 (
		\u1_sram_addr_reg[8]/P0001 ,
		\u6_wr_hold_reg/NET0131 ,
		_w1507_
	);
	LUT4 #(
		.INIT('h3777)
	) name548 (
		_w1333_,
		_w1335_,
		_w1338_,
		_w1507_,
		_w1508_
	);
	LUT4 #(
		.INIT('h010f)
	) name549 (
		\wb_addr_i[10]_pad ,
		_w1344_,
		_w1506_,
		_w1508_,
		_w1509_
	);
	LUT3 #(
		.INIT('h4f)
	) name550 (
		_w1502_,
		_w1505_,
		_w1509_,
		_w1510_
	);
	LUT3 #(
		.INIT('h51)
	) name551 (
		\u1_col_adr_reg[9]/P0001 ,
		\u5_state_reg[6]/NET0131 ,
		\u5_wb_wait_r_reg/P0001 ,
		_w1511_
	);
	LUT3 #(
		.INIT('h70)
	) name552 (
		_w1019_,
		_w1033_,
		_w1511_,
		_w1512_
	);
	LUT3 #(
		.INIT('h04)
	) name553 (
		\u1_row_adr_reg[9]/P0001 ,
		\u5_state_reg[6]/NET0131 ,
		\u5_wb_wait_r_reg/P0001 ,
		_w1513_
	);
	LUT3 #(
		.INIT('h40)
	) name554 (
		\u1_row_adr_reg[9]/P0001 ,
		_w966_,
		_w1018_,
		_w1514_
	);
	LUT3 #(
		.INIT('h13)
	) name555 (
		_w1033_,
		_w1513_,
		_w1514_,
		_w1515_
	);
	LUT2 #(
		.INIT('h4)
	) name556 (
		_w1512_,
		_w1515_,
		_w1516_
	);
	LUT4 #(
		.INIT('h001f)
	) name557 (
		\u5_wr_cycle_reg/NET0131 ,
		_w1324_,
		_w1327_,
		_w1516_,
		_w1517_
	);
	LUT3 #(
		.INIT('h15)
	) name558 (
		\u0_sp_tms_reg[9]/NET0131 ,
		\u5_cmd_del_reg[1]/NET0131 ,
		\u5_wr_cycle_reg/NET0131 ,
		_w1518_
	);
	LUT3 #(
		.INIT('h70)
	) name559 (
		_w976_,
		_w1114_,
		_w1518_,
		_w1519_
	);
	LUT4 #(
		.INIT('h10f0)
	) name560 (
		\u5_wr_cycle_reg/NET0131 ,
		_w1324_,
		_w1339_,
		_w1519_,
		_w1520_
	);
	LUT4 #(
		.INIT('h0080)
	) name561 (
		\u1_acs_addr_reg[9]/P0001 ,
		_w1333_,
		_w1335_,
		_w1338_,
		_w1521_
	);
	LUT2 #(
		.INIT('h4)
	) name562 (
		\u1_sram_addr_reg[9]/P0001 ,
		\u6_wr_hold_reg/NET0131 ,
		_w1522_
	);
	LUT4 #(
		.INIT('h3777)
	) name563 (
		_w1333_,
		_w1335_,
		_w1338_,
		_w1522_,
		_w1523_
	);
	LUT4 #(
		.INIT('h010f)
	) name564 (
		\wb_addr_i[11]_pad ,
		_w1344_,
		_w1521_,
		_w1523_,
		_w1524_
	);
	LUT3 #(
		.INIT('h4f)
	) name565 (
		_w1517_,
		_w1520_,
		_w1524_,
		_w1525_
	);
	LUT2 #(
		.INIT('h1)
	) name566 (
		\u5_rfr_ack_r_reg/NET0131 ,
		\u5_susp_sel_r_reg/NET0131 ,
		_w1526_
	);
	LUT3 #(
		.INIT('h01)
	) name567 (
		\u0_cs_reg[0]/NET0131 ,
		\u5_lmr_ack_reg/NET0131 ,
		\u5_state_reg[26]/NET0131 ,
		_w1527_
	);
	LUT3 #(
		.INIT('h80)
	) name568 (
		_w976_,
		_w1526_,
		_w1527_,
		_w1528_
	);
	LUT3 #(
		.INIT('h01)
	) name569 (
		\u0_spec_req_cs_reg[0]/NET0131 ,
		\u5_rfr_ack_r_reg/NET0131 ,
		\u5_susp_sel_r_reg/NET0131 ,
		_w1529_
	);
	LUT3 #(
		.INIT('h70)
	) name570 (
		_w976_,
		_w1114_,
		_w1529_,
		_w1530_
	);
	LUT4 #(
		.INIT('h0002)
	) name571 (
		\u0_u0_csc_reg[0]/NET0131 ,
		\u0_u0_csc_reg[1]/NET0131 ,
		\u0_u0_csc_reg[2]/NET0131 ,
		\u0_u0_csc_reg[3]/NET0131 ,
		_w1531_
	);
	LUT2 #(
		.INIT('h1)
	) name572 (
		_w1526_,
		_w1531_,
		_w1532_
	);
	LUT3 #(
		.INIT('h01)
	) name573 (
		_w1528_,
		_w1530_,
		_w1532_,
		_w1533_
	);
	LUT2 #(
		.INIT('h8)
	) name574 (
		\u5_cmd_del_reg[3]/NET0131 ,
		\u5_wr_cycle_reg/NET0131 ,
		_w1534_
	);
	LUT2 #(
		.INIT('h4)
	) name575 (
		\u5_cmd_del_reg[3]/NET0131 ,
		\u5_wr_cycle_reg/NET0131 ,
		_w1535_
	);
	LUT3 #(
		.INIT('h57)
	) name576 (
		_w982_,
		_w1181_,
		_w1289_,
		_w1536_
	);
	LUT3 #(
		.INIT('h51)
	) name577 (
		\u4_rfr_req_reg/NET0131 ,
		_w1002_,
		_w1536_,
		_w1537_
	);
	LUT3 #(
		.INIT('h04)
	) name578 (
		\u5_rfr_ack_r_reg/NET0131 ,
		_w1002_,
		_w1536_,
		_w1538_
	);
	LUT3 #(
		.INIT('h01)
	) name579 (
		_w1187_,
		_w1537_,
		_w1538_,
		_w1539_
	);
	LUT4 #(
		.INIT('h0777)
	) name580 (
		_w1068_,
		_w1070_,
		_w1100_,
		_w1102_,
		_w1540_
	);
	LUT3 #(
		.INIT('h02)
	) name581 (
		\u5_mc_c_oe_reg/NET0131 ,
		\u5_rfr_ack_r_reg/NET0131 ,
		\u5_susp_sel_r_reg/NET0131 ,
		_w1541_
	);
	LUT2 #(
		.INIT('h8)
	) name582 (
		_w1540_,
		_w1541_,
		_w1542_
	);
	LUT3 #(
		.INIT('h02)
	) name583 (
		\u0_tms_reg[19]/NET0131 ,
		\u5_lmr_ack_reg/NET0131 ,
		\u5_state_reg[26]/NET0131 ,
		_w1543_
	);
	LUT4 #(
		.INIT('h11d5)
	) name584 (
		\u0_sp_tms_reg[19]/NET0131 ,
		_w976_,
		_w1114_,
		_w1543_,
		_w1544_
	);
	LUT3 #(
		.INIT('h02)
	) name585 (
		\u0_tms_reg[18]/NET0131 ,
		\u5_lmr_ack_reg/NET0131 ,
		\u5_state_reg[26]/NET0131 ,
		_w1545_
	);
	LUT4 #(
		.INIT('h11d5)
	) name586 (
		\u0_sp_tms_reg[18]/NET0131 ,
		_w976_,
		_w1114_,
		_w1545_,
		_w1546_
	);
	LUT2 #(
		.INIT('h8)
	) name587 (
		_w1544_,
		_w1546_,
		_w1547_
	);
	LUT3 #(
		.INIT('h80)
	) name588 (
		_w1540_,
		_w1541_,
		_w1547_,
		_w1548_
	);
	LUT3 #(
		.INIT('h02)
	) name589 (
		\u0_tms_reg[17]/NET0131 ,
		\u5_lmr_ack_reg/NET0131 ,
		\u5_state_reg[26]/NET0131 ,
		_w1549_
	);
	LUT4 #(
		.INIT('h11d5)
	) name590 (
		\u0_sp_tms_reg[17]/NET0131 ,
		_w976_,
		_w1114_,
		_w1549_,
		_w1550_
	);
	LUT3 #(
		.INIT('h01)
	) name591 (
		\u0_tms_reg[16]/NET0131 ,
		\u5_lmr_ack_reg/NET0131 ,
		\u5_state_reg[26]/NET0131 ,
		_w1551_
	);
	LUT4 #(
		.INIT('h22ea)
	) name592 (
		\u0_sp_tms_reg[16]/NET0131 ,
		_w976_,
		_w1114_,
		_w1551_,
		_w1552_
	);
	LUT2 #(
		.INIT('h2)
	) name593 (
		_w1550_,
		_w1552_,
		_w1553_
	);
	LUT3 #(
		.INIT('h80)
	) name594 (
		_w1540_,
		_w1541_,
		_w1553_,
		_w1554_
	);
	LUT4 #(
		.INIT('h8aaa)
	) name595 (
		_w1153_,
		_w1539_,
		_w1548_,
		_w1554_,
		_w1555_
	);
	LUT4 #(
		.INIT('h5557)
	) name596 (
		_w1063_,
		_w1204_,
		_w1243_,
		_w1246_,
		_w1556_
	);
	LUT4 #(
		.INIT('h153f)
	) name597 (
		_w1041_,
		_w1063_,
		_w1236_,
		_w1261_,
		_w1557_
	);
	LUT3 #(
		.INIT('h40)
	) name598 (
		_w1145_,
		_w1556_,
		_w1557_,
		_w1558_
	);
	LUT4 #(
		.INIT('h153f)
	) name599 (
		_w1035_,
		_w1063_,
		_w1240_,
		_w1264_,
		_w1559_
	);
	LUT3 #(
		.INIT('h02)
	) name600 (
		\u5_state_reg[50]/NET0131 ,
		\u5_state_reg[51]/NET0131 ,
		\u5_tmr2_done_reg/NET0131 ,
		_w1560_
	);
	LUT2 #(
		.INIT('h8)
	) name601 (
		_w1176_,
		_w1560_,
		_w1561_
	);
	LUT4 #(
		.INIT('h0777)
	) name602 (
		_w1068_,
		_w1070_,
		_w1174_,
		_w1561_,
		_w1562_
	);
	LUT4 #(
		.INIT('h4000)
	) name603 (
		_w1084_,
		_w1106_,
		_w1559_,
		_w1562_,
		_w1563_
	);
	LUT4 #(
		.INIT('h7000)
	) name604 (
		_w1014_,
		_w1015_,
		_w1131_,
		_w1133_,
		_w1564_
	);
	LUT3 #(
		.INIT('h20)
	) name605 (
		\u6_read_go_r1_reg/NET0131 ,
		\u6_rmw_r_reg/NET0131 ,
		wb_cyc_i_pad,
		_w1565_
	);
	LUT3 #(
		.INIT('h70)
	) name606 (
		_w1014_,
		_w1015_,
		_w1565_,
		_w1566_
	);
	LUT2 #(
		.INIT('h1)
	) name607 (
		_w1564_,
		_w1566_,
		_w1567_
	);
	LUT3 #(
		.INIT('ha8)
	) name608 (
		_w1132_,
		_w1564_,
		_w1566_,
		_w1568_
	);
	LUT3 #(
		.INIT('h04)
	) name609 (
		_w1333_,
		_w1335_,
		_w1338_,
		_w1569_
	);
	LUT2 #(
		.INIT('h4)
	) name610 (
		_w1568_,
		_w1569_,
		_w1570_
	);
	LUT3 #(
		.INIT('hec)
	) name611 (
		_w1132_,
		_w1564_,
		_w1566_,
		_w1571_
	);
	LUT3 #(
		.INIT('h08)
	) name612 (
		_w1338_,
		_w1343_,
		_w1571_,
		_w1572_
	);
	LUT3 #(
		.INIT('h02)
	) name613 (
		\u0_cs_reg[1]/NET0131 ,
		\u5_lmr_ack_reg/NET0131 ,
		\u5_state_reg[26]/NET0131 ,
		_w1573_
	);
	LUT3 #(
		.INIT('h80)
	) name614 (
		_w976_,
		_w1526_,
		_w1573_,
		_w1574_
	);
	LUT3 #(
		.INIT('h02)
	) name615 (
		\u0_spec_req_cs_reg[1]/NET0131 ,
		\u5_rfr_ack_r_reg/NET0131 ,
		\u5_susp_sel_r_reg/NET0131 ,
		_w1575_
	);
	LUT3 #(
		.INIT('h70)
	) name616 (
		_w976_,
		_w1114_,
		_w1575_,
		_w1576_
	);
	LUT4 #(
		.INIT('h0002)
	) name617 (
		\u0_u1_csc_reg[0]/NET0131 ,
		\u0_u1_csc_reg[1]/NET0131 ,
		\u0_u1_csc_reg[2]/NET0131 ,
		\u0_u1_csc_reg[3]/NET0131 ,
		_w1577_
	);
	LUT2 #(
		.INIT('h4)
	) name618 (
		_w1526_,
		_w1577_,
		_w1578_
	);
	LUT3 #(
		.INIT('h01)
	) name619 (
		_w1574_,
		_w1576_,
		_w1578_,
		_w1579_
	);
	LUT3 #(
		.INIT('ha8)
	) name620 (
		\u5_lookup_ready2_reg/NET0131 ,
		_w1564_,
		_w1566_,
		_w1580_
	);
	LUT3 #(
		.INIT('hb0)
	) name621 (
		_w1533_,
		_w1579_,
		_w1580_,
		_w1581_
	);
	LUT3 #(
		.INIT('h15)
	) name622 (
		\u0_init_req_reg/NET0131 ,
		\u0_lmr_req_reg/NET0131 ,
		\u5_lookup_ready2_reg/NET0131 ,
		_w1582_
	);
	LUT2 #(
		.INIT('h2)
	) name623 (
		\u5_susp_req_r_reg/NET0131 ,
		\u5_wb_cycle_reg/NET0131 ,
		_w1583_
	);
	LUT3 #(
		.INIT('h51)
	) name624 (
		\u4_rfr_req_reg/NET0131 ,
		\u5_susp_req_r_reg/NET0131 ,
		\u5_wb_cycle_reg/NET0131 ,
		_w1584_
	);
	LUT3 #(
		.INIT('h80)
	) name625 (
		_w1185_,
		_w1582_,
		_w1584_,
		_w1585_
	);
	LUT2 #(
		.INIT('h8)
	) name626 (
		_w1184_,
		_w1585_,
		_w1586_
	);
	LUT4 #(
		.INIT('he000)
	) name627 (
		_w1570_,
		_w1572_,
		_w1581_,
		_w1586_,
		_w1587_
	);
	LUT4 #(
		.INIT('h0080)
	) name628 (
		_w1225_,
		_w1558_,
		_w1563_,
		_w1587_,
		_w1588_
	);
	LUT3 #(
		.INIT('h40)
	) name629 (
		\u5_wb_wait_r_reg/P0001 ,
		_w1100_,
		_w1161_,
		_w1589_
	);
	LUT3 #(
		.INIT('h80)
	) name630 (
		_w1100_,
		_w1277_,
		_w1279_,
		_w1590_
	);
	LUT4 #(
		.INIT('h0040)
	) name631 (
		_w1159_,
		_w1286_,
		_w1306_,
		_w1590_,
		_w1591_
	);
	LUT3 #(
		.INIT('h57)
	) name632 (
		_w1041_,
		_w1079_,
		_w1195_,
		_w1592_
	);
	LUT3 #(
		.INIT('h40)
	) name633 (
		\u5_tmr_done_reg/NET0131 ,
		_w1059_,
		_w1086_,
		_w1593_
	);
	LUT4 #(
		.INIT('h0010)
	) name634 (
		_w1156_,
		_w1192_,
		_w1592_,
		_w1593_,
		_w1594_
	);
	LUT3 #(
		.INIT('h40)
	) name635 (
		_w1589_,
		_w1591_,
		_w1594_,
		_w1595_
	);
	LUT4 #(
		.INIT('h2000)
	) name636 (
		_w1314_,
		_w1555_,
		_w1588_,
		_w1595_,
		_w1596_
	);
	LUT4 #(
		.INIT('h8880)
	) name637 (
		_w1100_,
		_w1140_,
		_w1301_,
		_w1302_,
		_w1597_
	);
	LUT4 #(
		.INIT('h8000)
	) name638 (
		_w1122_,
		_w1124_,
		_w1127_,
		_w1541_,
		_w1598_
	);
	LUT4 #(
		.INIT('h7000)
	) name639 (
		_w1187_,
		_w1292_,
		_w1540_,
		_w1598_,
		_w1599_
	);
	LUT3 #(
		.INIT('h80)
	) name640 (
		_w1122_,
		_w1124_,
		_w1127_,
		_w1600_
	);
	LUT4 #(
		.INIT('h2aaa)
	) name641 (
		_w1116_,
		_w1122_,
		_w1124_,
		_w1127_,
		_w1601_
	);
	LUT2 #(
		.INIT('h1)
	) name642 (
		\u5_burst_cnt_reg[0]/NET0131 ,
		\u5_burst_cnt_reg[1]/NET0131 ,
		_w1602_
	);
	LUT3 #(
		.INIT('h01)
	) name643 (
		\u5_burst_cnt_reg[0]/NET0131 ,
		\u5_burst_cnt_reg[1]/NET0131 ,
		\u5_burst_cnt_reg[2]/NET0131 ,
		_w1603_
	);
	LUT4 #(
		.INIT('h0001)
	) name644 (
		\u5_burst_cnt_reg[3]/NET0131 ,
		\u5_burst_cnt_reg[4]/NET0131 ,
		\u5_burst_cnt_reg[5]/NET0131 ,
		\u5_burst_cnt_reg[6]/NET0131 ,
		_w1604_
	);
	LUT2 #(
		.INIT('h8)
	) name645 (
		_w1603_,
		_w1604_,
		_w1605_
	);
	LUT2 #(
		.INIT('h1)
	) name646 (
		\u5_burst_cnt_reg[7]/NET0131 ,
		\u5_burst_cnt_reg[8]/NET0131 ,
		_w1606_
	);
	LUT4 #(
		.INIT('h0001)
	) name647 (
		\u5_burst_cnt_reg[10]/NET0131 ,
		\u5_burst_cnt_reg[7]/NET0131 ,
		\u5_burst_cnt_reg[8]/NET0131 ,
		\u5_burst_cnt_reg[9]/NET0131 ,
		_w1607_
	);
	LUT3 #(
		.INIT('h80)
	) name648 (
		_w1603_,
		_w1604_,
		_w1607_,
		_w1608_
	);
	LUT3 #(
		.INIT('h7f)
	) name649 (
		_w1603_,
		_w1604_,
		_w1607_,
		_w1609_
	);
	LUT4 #(
		.INIT('h1555)
	) name650 (
		\u5_wb_write_go_r_reg/NET0131 ,
		_w1603_,
		_w1604_,
		_w1607_,
		_w1610_
	);
	LUT2 #(
		.INIT('h8)
	) name651 (
		_w1601_,
		_w1610_,
		_w1611_
	);
	LUT2 #(
		.INIT('h4)
	) name652 (
		\u5_cnt_reg/NET0131 ,
		_w1116_,
		_w1612_
	);
	LUT3 #(
		.INIT('h8a)
	) name653 (
		\u5_cke_r_reg/NET0131 ,
		_w1600_,
		_w1612_,
		_w1613_
	);
	LUT3 #(
		.INIT('h10)
	) name654 (
		_w1568_,
		_w1600_,
		_w1612_,
		_w1614_
	);
	LUT4 #(
		.INIT('h5c55)
	) name655 (
		\u5_cke_r_reg/NET0131 ,
		_w1568_,
		_w1600_,
		_w1612_,
		_w1615_
	);
	LUT2 #(
		.INIT('h2)
	) name656 (
		_w1141_,
		_w1615_,
		_w1616_
	);
	LUT4 #(
		.INIT('hb000)
	) name657 (
		_w1539_,
		_w1599_,
		_w1611_,
		_w1616_,
		_w1617_
	);
	LUT2 #(
		.INIT('h1)
	) name658 (
		_w1597_,
		_w1617_,
		_w1618_
	);
	LUT3 #(
		.INIT('h01)
	) name659 (
		_w1534_,
		_w1597_,
		_w1617_,
		_w1619_
	);
	LUT4 #(
		.INIT('hfddd)
	) name660 (
		_w1533_,
		_w1535_,
		_w1596_,
		_w1619_,
		_w1620_
	);
	LUT4 #(
		.INIT('hfeee)
	) name661 (
		_w1535_,
		_w1579_,
		_w1596_,
		_w1619_,
		_w1621_
	);
	LUT2 #(
		.INIT('h2)
	) name662 (
		_w1304_,
		_w1615_,
		_w1622_
	);
	LUT4 #(
		.INIT('h4f00)
	) name663 (
		_w1539_,
		_w1599_,
		_w1611_,
		_w1622_,
		_w1623_
	);
	LUT3 #(
		.INIT('h08)
	) name664 (
		_w1100_,
		_w1277_,
		_w1279_,
		_w1624_
	);
	LUT4 #(
		.INIT('h135f)
	) name665 (
		_w1002_,
		_w1059_,
		_w1182_,
		_w1189_,
		_w1625_
	);
	LUT4 #(
		.INIT('h0800)
	) name666 (
		_w1315_,
		_w1319_,
		_w1624_,
		_w1625_,
		_w1626_
	);
	LUT4 #(
		.INIT('h8000)
	) name667 (
		_w1081_,
		_w1209_,
		_w1313_,
		_w1626_,
		_w1627_
	);
	LUT2 #(
		.INIT('h2)
	) name668 (
		_w1582_,
		_w1583_,
		_w1628_
	);
	LUT3 #(
		.INIT('h08)
	) name669 (
		\u5_lookup_ready2_reg/NET0131 ,
		_w1582_,
		_w1583_,
		_w1629_
	);
	LUT3 #(
		.INIT('he0)
	) name670 (
		_w1564_,
		_w1566_,
		_w1629_,
		_w1630_
	);
	LUT3 #(
		.INIT('hb0)
	) name671 (
		_w1533_,
		_w1579_,
		_w1630_,
		_w1631_
	);
	LUT4 #(
		.INIT('hf0d0)
	) name672 (
		_w1135_,
		_w1333_,
		_w1335_,
		_w1338_,
		_w1632_
	);
	LUT4 #(
		.INIT('h00b0)
	) name673 (
		_w1533_,
		_w1579_,
		_w1630_,
		_w1632_,
		_w1633_
	);
	LUT2 #(
		.INIT('h2)
	) name674 (
		_w1186_,
		_w1633_,
		_w1634_
	);
	LUT3 #(
		.INIT('h20)
	) name675 (
		\u4_rfr_req_reg/NET0131 ,
		\u5_state_reg[0]/NET0131 ,
		\u5_state_reg[1]/NET0131 ,
		_w1635_
	);
	LUT4 #(
		.INIT('h0777)
	) name676 (
		_w1035_,
		_w1168_,
		_w1184_,
		_w1635_,
		_w1636_
	);
	LUT4 #(
		.INIT('h153f)
	) name677 (
		_w991_,
		_w1100_,
		_w1161_,
		_w1213_,
		_w1637_
	);
	LUT4 #(
		.INIT('h8000)
	) name678 (
		_w1320_,
		_w1321_,
		_w1636_,
		_w1637_,
		_w1638_
	);
	LUT3 #(
		.INIT('h80)
	) name679 (
		\u5_tmr_done_reg/NET0131 ,
		_w1059_,
		_w1086_,
		_w1639_
	);
	LUT3 #(
		.INIT('h04)
	) name680 (
		_w1084_,
		_w1106_,
		_w1639_,
		_w1640_
	);
	LUT3 #(
		.INIT('h40)
	) name681 (
		_w1634_,
		_w1638_,
		_w1640_,
		_w1641_
	);
	LUT4 #(
		.INIT('h0008)
	) name682 (
		_w1141_,
		_w1303_,
		_w1613_,
		_w1614_,
		_w1642_
	);
	LUT3 #(
		.INIT('h08)
	) name683 (
		_w1254_,
		_w1266_,
		_w1642_,
		_w1643_
	);
	LUT4 #(
		.INIT('h8000)
	) name684 (
		_w1073_,
		_w1627_,
		_w1641_,
		_w1643_,
		_w1644_
	);
	LUT2 #(
		.INIT('hb)
	) name685 (
		_w1623_,
		_w1644_,
		_w1645_
	);
	LUT2 #(
		.INIT('h8)
	) name686 (
		\u5_cmd_asserted_reg/NET0131 ,
		\u5_mc_le_reg/NET0131 ,
		_w1646_
	);
	LUT2 #(
		.INIT('h4)
	) name687 (
		\u5_cmd_asserted_reg/NET0131 ,
		\u5_mc_le_reg/NET0131 ,
		_w1647_
	);
	LUT3 #(
		.INIT('h01)
	) name688 (
		_w1597_,
		_w1617_,
		_w1646_,
		_w1648_
	);
	LUT3 #(
		.INIT('h13)
	) name689 (
		_w1596_,
		_w1647_,
		_w1648_,
		_w1649_
	);
	LUT4 #(
		.INIT('h0020)
	) name690 (
		_w1135_,
		_w1333_,
		_w1335_,
		_w1338_,
		_w1650_
	);
	LUT3 #(
		.INIT('h80)
	) name691 (
		_w1184_,
		_w1585_,
		_w1650_,
		_w1651_
	);
	LUT3 #(
		.INIT('h15)
	) name692 (
		_w1173_,
		_w1581_,
		_w1651_,
		_w1652_
	);
	LUT3 #(
		.INIT('h0b)
	) name693 (
		_w1539_,
		_w1542_,
		_w1652_,
		_w1653_
	);
	LUT3 #(
		.INIT('h02)
	) name694 (
		\u0_tms_reg[14]/NET0131 ,
		\u5_lmr_ack_reg/NET0131 ,
		\u5_state_reg[26]/NET0131 ,
		_w1654_
	);
	LUT4 #(
		.INIT('h11d5)
	) name695 (
		\u0_sp_tms_reg[14]/NET0131 ,
		_w976_,
		_w1114_,
		_w1654_,
		_w1655_
	);
	LUT4 #(
		.INIT('hea00)
	) name696 (
		_w1173_,
		_w1581_,
		_w1651_,
		_w1655_,
		_w1656_
	);
	LUT4 #(
		.INIT('hf400)
	) name697 (
		_w1539_,
		_w1542_,
		_w1652_,
		_w1656_,
		_w1657_
	);
	LUT3 #(
		.INIT('h20)
	) name698 (
		_w1059_,
		_w1223_,
		_w1252_,
		_w1658_
	);
	LUT3 #(
		.INIT('h10)
	) name699 (
		\u5_state_reg[58]/NET0131 ,
		\u5_state_reg[59]/NET0131 ,
		\u5_tmr_done_reg/NET0131 ,
		_w1659_
	);
	LUT3 #(
		.INIT('h80)
	) name700 (
		_w985_,
		_w1222_,
		_w1659_,
		_w1660_
	);
	LUT2 #(
		.INIT('h8)
	) name701 (
		_w1059_,
		_w1660_,
		_w1661_
	);
	LUT4 #(
		.INIT('h55df)
	) name702 (
		_w1059_,
		_w1223_,
		_w1252_,
		_w1660_,
		_w1662_
	);
	LUT3 #(
		.INIT('h02)
	) name703 (
		\u0_tms_reg[10]/NET0131 ,
		\u5_lmr_ack_reg/NET0131 ,
		\u5_state_reg[26]/NET0131 ,
		_w1663_
	);
	LUT4 #(
		.INIT('h11d5)
	) name704 (
		\u0_sp_tms_reg[10]/NET0131 ,
		_w976_,
		_w1114_,
		_w1663_,
		_w1664_
	);
	LUT2 #(
		.INIT('h4)
	) name705 (
		_w1662_,
		_w1664_,
		_w1665_
	);
	LUT3 #(
		.INIT('h04)
	) name706 (
		_w1338_,
		_w1343_,
		_w1571_,
		_w1666_
	);
	LUT4 #(
		.INIT('h1555)
	) name707 (
		_w1084_,
		_w1581_,
		_w1586_,
		_w1666_,
		_w1667_
	);
	LUT3 #(
		.INIT('h80)
	) name708 (
		_w1124_,
		_w1540_,
		_w1541_,
		_w1668_
	);
	LUT4 #(
		.INIT('hc4c0)
	) name709 (
		_w1539_,
		_w1662_,
		_w1667_,
		_w1668_,
		_w1669_
	);
	LUT2 #(
		.INIT('h1)
	) name710 (
		_w1665_,
		_w1669_,
		_w1670_
	);
	LUT4 #(
		.INIT('h4555)
	) name711 (
		\u5_state_reg[9]/NET0131 ,
		\u5_wb_wait_r_reg/P0001 ,
		_w1100_,
		_w1161_,
		_w1671_
	);
	LUT2 #(
		.INIT('h8)
	) name712 (
		_w1591_,
		_w1671_,
		_w1672_
	);
	LUT4 #(
		.INIT('h0001)
	) name713 (
		\u5_state_reg[17]/NET0131 ,
		\u5_state_reg[20]/NET0131 ,
		\u5_state_reg[24]/NET0131 ,
		\u5_state_reg[26]/NET0131 ,
		_w1673_
	);
	LUT2 #(
		.INIT('h1)
	) name714 (
		\u5_timer_reg[2]/NET0131 ,
		\u5_timer_reg[3]/NET0131 ,
		_w1674_
	);
	LUT4 #(
		.INIT('h0001)
	) name715 (
		\u5_timer_reg[2]/NET0131 ,
		\u5_timer_reg[3]/NET0131 ,
		\u5_timer_reg[4]/NET0131 ,
		\u5_timer_reg[5]/NET0131 ,
		_w1675_
	);
	LUT4 #(
		.INIT('h0001)
	) name716 (
		\u5_timer_reg[0]/NET0131 ,
		\u5_timer_reg[1]/NET0131 ,
		\u5_timer_reg[6]/NET0131 ,
		\u5_timer_reg[7]/NET0131 ,
		_w1676_
	);
	LUT2 #(
		.INIT('h8)
	) name717 (
		_w1675_,
		_w1676_,
		_w1677_
	);
	LUT3 #(
		.INIT('h01)
	) name718 (
		\u5_mc_le_reg/NET0131 ,
		\u5_timer_reg[0]/NET0131 ,
		\u5_timer_reg[1]/NET0131 ,
		_w1678_
	);
	LUT3 #(
		.INIT('h70)
	) name719 (
		_w1675_,
		_w1676_,
		_w1678_,
		_w1679_
	);
	LUT3 #(
		.INIT('h01)
	) name720 (
		\u5_state_reg[30]/NET0131 ,
		\u5_state_reg[31]/NET0131 ,
		\u5_timer_reg[2]/NET0131 ,
		_w1680_
	);
	LUT4 #(
		.INIT('h8f00)
	) name721 (
		_w1675_,
		_w1676_,
		_w1678_,
		_w1680_,
		_w1681_
	);
	LUT3 #(
		.INIT('h10)
	) name722 (
		\u5_state_reg[30]/NET0131 ,
		\u5_state_reg[31]/NET0131 ,
		\u5_timer_reg[2]/NET0131 ,
		_w1682_
	);
	LUT4 #(
		.INIT('h7000)
	) name723 (
		_w1675_,
		_w1676_,
		_w1678_,
		_w1682_,
		_w1683_
	);
	LUT4 #(
		.INIT('hccc8)
	) name724 (
		\u5_state_reg[35]/NET0131 ,
		_w1673_,
		_w1681_,
		_w1683_,
		_w1684_
	);
	LUT3 #(
		.INIT('h2a)
	) name725 (
		\u0_sp_tms_reg[26]/NET0131 ,
		_w976_,
		_w1114_,
		_w1685_
	);
	LUT3 #(
		.INIT('h02)
	) name726 (
		\u0_tms_reg[26]/NET0131 ,
		\u5_lmr_ack_reg/NET0131 ,
		\u5_state_reg[26]/NET0131 ,
		_w1686_
	);
	LUT3 #(
		.INIT('h13)
	) name727 (
		_w976_,
		_w1673_,
		_w1686_,
		_w1687_
	);
	LUT2 #(
		.INIT('h4)
	) name728 (
		_w1685_,
		_w1687_,
		_w1688_
	);
	LUT3 #(
		.INIT('h80)
	) name729 (
		_w1540_,
		_w1541_,
		_w1688_,
		_w1689_
	);
	LUT3 #(
		.INIT('h23)
	) name730 (
		_w1539_,
		_w1684_,
		_w1689_,
		_w1690_
	);
	LUT2 #(
		.INIT('h8)
	) name731 (
		_w1672_,
		_w1690_,
		_w1691_
	);
	LUT3 #(
		.INIT('h02)
	) name732 (
		\u0_tms_reg[22]/NET0131 ,
		\u5_lmr_ack_reg/NET0131 ,
		\u5_state_reg[26]/NET0131 ,
		_w1692_
	);
	LUT4 #(
		.INIT('h11d5)
	) name733 (
		\u0_sp_tms_reg[22]/NET0131 ,
		_w976_,
		_w1114_,
		_w1692_,
		_w1693_
	);
	LUT3 #(
		.INIT('h80)
	) name734 (
		_w1540_,
		_w1541_,
		_w1693_,
		_w1694_
	);
	LUT3 #(
		.INIT('h23)
	) name735 (
		_w1539_,
		_w1591_,
		_w1694_,
		_w1695_
	);
	LUT2 #(
		.INIT('h1)
	) name736 (
		\u5_state_reg[13]/NET0131 ,
		\u5_state_reg[14]/NET0131 ,
		_w1696_
	);
	LUT3 #(
		.INIT('h80)
	) name737 (
		_w1540_,
		_w1541_,
		_w1544_,
		_w1697_
	);
	LUT4 #(
		.INIT('h80c0)
	) name738 (
		_w1539_,
		_w1589_,
		_w1591_,
		_w1697_,
		_w1698_
	);
	LUT3 #(
		.INIT('h04)
	) name739 (
		_w1695_,
		_w1696_,
		_w1698_,
		_w1699_
	);
	LUT3 #(
		.INIT('h01)
	) name740 (
		\u0_tms_reg[21]/NET0131 ,
		\u5_lmr_ack_reg/NET0131 ,
		\u5_state_reg[26]/NET0131 ,
		_w1700_
	);
	LUT4 #(
		.INIT('h22ea)
	) name741 (
		\u0_sp_tms_reg[21]/NET0131 ,
		_w976_,
		_w1114_,
		_w1700_,
		_w1701_
	);
	LUT2 #(
		.INIT('h8)
	) name742 (
		_w1552_,
		_w1701_,
		_w1702_
	);
	LUT3 #(
		.INIT('h08)
	) name743 (
		_w1540_,
		_w1541_,
		_w1702_,
		_w1703_
	);
	LUT2 #(
		.INIT('h1)
	) name744 (
		_w1552_,
		_w1701_,
		_w1704_
	);
	LUT3 #(
		.INIT('h80)
	) name745 (
		_w1540_,
		_w1541_,
		_w1704_,
		_w1705_
	);
	LUT3 #(
		.INIT('h02)
	) name746 (
		\u0_tms_reg[15]/NET0131 ,
		\u5_lmr_ack_reg/NET0131 ,
		\u5_state_reg[26]/NET0131 ,
		_w1706_
	);
	LUT4 #(
		.INIT('h11d5)
	) name747 (
		\u0_sp_tms_reg[15]/NET0131 ,
		_w976_,
		_w1114_,
		_w1706_,
		_w1707_
	);
	LUT3 #(
		.INIT('h02)
	) name748 (
		\u0_tms_reg[20]/NET0131 ,
		\u5_lmr_ack_reg/NET0131 ,
		\u5_state_reg[26]/NET0131 ,
		_w1708_
	);
	LUT4 #(
		.INIT('h11d5)
	) name749 (
		\u0_sp_tms_reg[20]/NET0131 ,
		_w976_,
		_w1114_,
		_w1708_,
		_w1709_
	);
	LUT2 #(
		.INIT('h1)
	) name750 (
		_w1707_,
		_w1709_,
		_w1710_
	);
	LUT3 #(
		.INIT('h08)
	) name751 (
		_w1540_,
		_w1541_,
		_w1710_,
		_w1711_
	);
	LUT3 #(
		.INIT('hab)
	) name752 (
		_w1539_,
		_w1705_,
		_w1711_,
		_w1712_
	);
	LUT4 #(
		.INIT('h4440)
	) name753 (
		_w1539_,
		_w1703_,
		_w1705_,
		_w1711_,
		_w1713_
	);
	LUT3 #(
		.INIT('h0b)
	) name754 (
		_w1539_,
		_w1694_,
		_w1696_,
		_w1714_
	);
	LUT3 #(
		.INIT('h04)
	) name755 (
		_w1539_,
		_w1694_,
		_w1696_,
		_w1715_
	);
	LUT4 #(
		.INIT('h0145)
	) name756 (
		_w1665_,
		_w1713_,
		_w1714_,
		_w1715_,
		_w1716_
	);
	LUT4 #(
		.INIT('h8a00)
	) name757 (
		_w1667_,
		_w1691_,
		_w1699_,
		_w1716_,
		_w1717_
	);
	LUT4 #(
		.INIT('hf040)
	) name758 (
		_w1539_,
		_w1542_,
		_w1652_,
		_w1662_,
		_w1718_
	);
	LUT4 #(
		.INIT('h5455)
	) name759 (
		_w1657_,
		_w1670_,
		_w1717_,
		_w1718_,
		_w1719_
	);
	LUT3 #(
		.INIT('h20)
	) name760 (
		\u5_cmd_asserted_reg/NET0131 ,
		\u5_state_reg[12]/NET0131 ,
		\u5_state_reg[13]/NET0131 ,
		_w1720_
	);
	LUT2 #(
		.INIT('h4)
	) name761 (
		\u5_mem_ack_r_reg/NET0131 ,
		\u5_wb_cycle_reg/NET0131 ,
		_w1721_
	);
	LUT3 #(
		.INIT('h80)
	) name762 (
		_w1135_,
		_w1720_,
		_w1721_,
		_w1722_
	);
	LUT4 #(
		.INIT('h0800)
	) name763 (
		_w1002_,
		_w1143_,
		_w1608_,
		_w1722_,
		_w1723_
	);
	LUT3 #(
		.INIT('hb0)
	) name764 (
		_w1539_,
		_w1599_,
		_w1723_,
		_w1724_
	);
	LUT2 #(
		.INIT('h4)
	) name765 (
		\u5_mem_ack_r_reg/NET0131 ,
		\u5_wr_cycle_reg/NET0131 ,
		_w1725_
	);
	LUT2 #(
		.INIT('h8)
	) name766 (
		_w1135_,
		_w1725_,
		_w1726_
	);
	LUT4 #(
		.INIT('h0800)
	) name767 (
		_w1100_,
		_w1140_,
		_w1608_,
		_w1726_,
		_w1727_
	);
	LUT3 #(
		.INIT('hb0)
	) name768 (
		_w1539_,
		_w1599_,
		_w1727_,
		_w1728_
	);
	LUT4 #(
		.INIT('h8880)
	) name769 (
		\u5_tmr_done_reg/NET0131 ,
		_w1059_,
		_w1086_,
		_w1223_,
		_w1729_
	);
	LUT2 #(
		.INIT('h4)
	) name770 (
		\u5_mem_ack_r_reg/NET0131 ,
		_w1135_,
		_w1730_
	);
	LUT3 #(
		.INIT('h80)
	) name771 (
		_w1100_,
		_w1108_,
		_w1730_,
		_w1731_
	);
	LUT4 #(
		.INIT('h0002)
	) name772 (
		_w1066_,
		_w1231_,
		_w1729_,
		_w1731_,
		_w1732_
	);
	LUT2 #(
		.INIT('h8)
	) name773 (
		wb_stb_i_pad,
		wb_we_i_pad,
		_w1733_
	);
	LUT2 #(
		.INIT('h1)
	) name774 (
		\u5_ack_cnt_reg[0]/NET0131 ,
		\u5_ack_cnt_reg[1]/NET0131 ,
		_w1734_
	);
	LUT4 #(
		.INIT('h0001)
	) name775 (
		\u5_ack_cnt_reg[0]/NET0131 ,
		\u5_ack_cnt_reg[1]/NET0131 ,
		\u5_ack_cnt_reg[2]/NET0131 ,
		\u5_ack_cnt_reg[3]/NET0131 ,
		_w1735_
	);
	LUT4 #(
		.INIT('h0070)
	) name776 (
		_w1014_,
		_w1015_,
		_w1565_,
		_w1735_,
		_w1736_
	);
	LUT3 #(
		.INIT('h10)
	) name777 (
		\u5_mem_ack_r_reg/NET0131 ,
		_w1733_,
		_w1736_,
		_w1737_
	);
	LUT2 #(
		.INIT('h4)
	) name778 (
		_w1568_,
		_w1737_,
		_w1738_
	);
	LUT4 #(
		.INIT('h2000)
	) name779 (
		_w1135_,
		_w1333_,
		_w1335_,
		_w1338_,
		_w1739_
	);
	LUT3 #(
		.INIT('h80)
	) name780 (
		_w1184_,
		_w1585_,
		_w1739_,
		_w1740_
	);
	LUT3 #(
		.INIT('h08)
	) name781 (
		\u5_cmd_asserted_reg/NET0131 ,
		\u5_state_reg[58]/NET0131 ,
		\u5_state_reg[59]/NET0131 ,
		_w1741_
	);
	LUT3 #(
		.INIT('h80)
	) name782 (
		_w985_,
		_w986_,
		_w1741_,
		_w1742_
	);
	LUT3 #(
		.INIT('h80)
	) name783 (
		_w1059_,
		_w1730_,
		_w1742_,
		_w1743_
	);
	LUT2 #(
		.INIT('h4)
	) name784 (
		\u5_mem_ack_r_reg/NET0131 ,
		_w1270_,
		_w1744_
	);
	LUT3 #(
		.INIT('h80)
	) name785 (
		_w1100_,
		_w1110_,
		_w1744_,
		_w1745_
	);
	LUT4 #(
		.INIT('h0007)
	) name786 (
		_w1581_,
		_w1740_,
		_w1743_,
		_w1745_,
		_w1746_
	);
	LUT3 #(
		.INIT('h20)
	) name787 (
		_w1732_,
		_w1738_,
		_w1746_,
		_w1747_
	);
	LUT3 #(
		.INIT('h01)
	) name788 (
		\wb_addr_i[29]_pad ,
		\wb_addr_i[30]_pad ,
		\wb_addr_i[31]_pad ,
		_w1748_
	);
	LUT3 #(
		.INIT('he0)
	) name789 (
		_w1564_,
		_w1566_,
		_w1748_,
		_w1749_
	);
	LUT4 #(
		.INIT('hef00)
	) name790 (
		_w1724_,
		_w1728_,
		_w1747_,
		_w1749_,
		_w1750_
	);
	LUT2 #(
		.INIT('h4)
	) name791 (
		_w1013_,
		_w1750_,
		_w1751_
	);
	LUT4 #(
		.INIT('h0002)
	) name792 (
		\u3_u0_rd_adr_reg[0]/NET0131 ,
		\u3_u0_rd_adr_reg[1]/NET0131 ,
		\u3_u0_rd_adr_reg[2]/NET0131 ,
		\u3_u0_rd_adr_reg[3]/NET0131 ,
		_w1752_
	);
	LUT4 #(
		.INIT('h0004)
	) name793 (
		\u3_u0_rd_adr_reg[0]/NET0131 ,
		\u3_u0_rd_adr_reg[1]/NET0131 ,
		\u3_u0_rd_adr_reg[2]/NET0131 ,
		\u3_u0_rd_adr_reg[3]/NET0131 ,
		_w1753_
	);
	LUT4 #(
		.INIT('h135f)
	) name794 (
		\u3_u0_r0_reg[13]/P0001 ,
		\u3_u0_r1_reg[13]/P0001 ,
		_w1752_,
		_w1753_,
		_w1754_
	);
	LUT4 #(
		.INIT('h0100)
	) name795 (
		\u3_u0_rd_adr_reg[0]/NET0131 ,
		\u3_u0_rd_adr_reg[1]/NET0131 ,
		\u3_u0_rd_adr_reg[2]/NET0131 ,
		\u3_u0_rd_adr_reg[3]/NET0131 ,
		_w1755_
	);
	LUT4 #(
		.INIT('h0010)
	) name796 (
		\u3_u0_rd_adr_reg[0]/NET0131 ,
		\u3_u0_rd_adr_reg[1]/NET0131 ,
		\u3_u0_rd_adr_reg[2]/NET0131 ,
		\u3_u0_rd_adr_reg[3]/NET0131 ,
		_w1756_
	);
	LUT4 #(
		.INIT('h153f)
	) name797 (
		\u3_u0_r2_reg[13]/P0001 ,
		\u3_u0_r3_reg[13]/P0001 ,
		_w1755_,
		_w1756_,
		_w1757_
	);
	LUT4 #(
		.INIT('h135f)
	) name798 (
		\u3_u0_r0_reg[9]/P0001 ,
		\u3_u0_r1_reg[9]/P0001 ,
		_w1752_,
		_w1753_,
		_w1758_
	);
	LUT4 #(
		.INIT('h153f)
	) name799 (
		\u3_u0_r2_reg[9]/P0001 ,
		\u3_u0_r3_reg[9]/P0001 ,
		_w1755_,
		_w1756_,
		_w1759_
	);
	LUT4 #(
		.INIT('h8777)
	) name800 (
		_w1754_,
		_w1757_,
		_w1758_,
		_w1759_,
		_w1760_
	);
	LUT4 #(
		.INIT('h135f)
	) name801 (
		\u3_u0_r0_reg[14]/P0001 ,
		\u3_u0_r1_reg[14]/P0001 ,
		_w1752_,
		_w1753_,
		_w1761_
	);
	LUT4 #(
		.INIT('h153f)
	) name802 (
		\u3_u0_r2_reg[14]/P0001 ,
		\u3_u0_r3_reg[14]/P0001 ,
		_w1755_,
		_w1756_,
		_w1762_
	);
	LUT2 #(
		.INIT('h8)
	) name803 (
		_w1761_,
		_w1762_,
		_w1763_
	);
	LUT4 #(
		.INIT('h135f)
	) name804 (
		\u3_u0_r0_reg[11]/P0001 ,
		\u3_u0_r1_reg[11]/P0001 ,
		_w1752_,
		_w1753_,
		_w1764_
	);
	LUT4 #(
		.INIT('h153f)
	) name805 (
		\u3_u0_r2_reg[11]/P0001 ,
		\u3_u0_r3_reg[11]/P0001 ,
		_w1755_,
		_w1756_,
		_w1765_
	);
	LUT4 #(
		.INIT('h135f)
	) name806 (
		\u3_u0_r0_reg[12]/P0001 ,
		\u3_u0_r1_reg[12]/P0001 ,
		_w1752_,
		_w1753_,
		_w1766_
	);
	LUT4 #(
		.INIT('h153f)
	) name807 (
		\u3_u0_r2_reg[12]/P0001 ,
		\u3_u0_r3_reg[12]/P0001 ,
		_w1755_,
		_w1756_,
		_w1767_
	);
	LUT4 #(
		.INIT('h7888)
	) name808 (
		_w1764_,
		_w1765_,
		_w1766_,
		_w1767_,
		_w1768_
	);
	LUT3 #(
		.INIT('h69)
	) name809 (
		_w1760_,
		_w1763_,
		_w1768_,
		_w1769_
	);
	LUT4 #(
		.INIT('h135f)
	) name810 (
		\u3_u0_r0_reg[8]/P0001 ,
		\u3_u0_r1_reg[8]/P0001 ,
		_w1752_,
		_w1753_,
		_w1770_
	);
	LUT4 #(
		.INIT('h153f)
	) name811 (
		\u3_u0_r2_reg[8]/P0001 ,
		\u3_u0_r3_reg[8]/P0001 ,
		_w1755_,
		_w1756_,
		_w1771_
	);
	LUT4 #(
		.INIT('h135f)
	) name812 (
		\u3_u0_r0_reg[15]/P0001 ,
		\u3_u0_r1_reg[15]/P0001 ,
		_w1752_,
		_w1753_,
		_w1772_
	);
	LUT4 #(
		.INIT('h153f)
	) name813 (
		\u3_u0_r2_reg[15]/P0001 ,
		\u3_u0_r3_reg[15]/P0001 ,
		_w1755_,
		_w1756_,
		_w1773_
	);
	LUT4 #(
		.INIT('h8777)
	) name814 (
		_w1770_,
		_w1771_,
		_w1772_,
		_w1773_,
		_w1774_
	);
	LUT4 #(
		.INIT('h135f)
	) name815 (
		\u3_u0_r0_reg[33]/P0001 ,
		\u3_u0_r1_reg[33]/P0001 ,
		_w1752_,
		_w1753_,
		_w1775_
	);
	LUT4 #(
		.INIT('h153f)
	) name816 (
		\u3_u0_r2_reg[33]/P0001 ,
		\u3_u0_r3_reg[33]/P0001 ,
		_w1755_,
		_w1756_,
		_w1776_
	);
	LUT4 #(
		.INIT('h135f)
	) name817 (
		\u3_u0_r0_reg[10]/P0001 ,
		\u3_u0_r1_reg[10]/P0001 ,
		_w1752_,
		_w1753_,
		_w1777_
	);
	LUT4 #(
		.INIT('h153f)
	) name818 (
		\u3_u0_r2_reg[10]/P0001 ,
		\u3_u0_r3_reg[10]/P0001 ,
		_w1755_,
		_w1756_,
		_w1778_
	);
	LUT4 #(
		.INIT('h8777)
	) name819 (
		_w1775_,
		_w1776_,
		_w1777_,
		_w1778_,
		_w1779_
	);
	LUT2 #(
		.INIT('h6)
	) name820 (
		_w1774_,
		_w1779_,
		_w1780_
	);
	LUT2 #(
		.INIT('h2)
	) name821 (
		_w1769_,
		_w1780_,
		_w1781_
	);
	LUT4 #(
		.INIT('h2002)
	) name822 (
		\wb_sel_i[1]_pad ,
		_w1760_,
		_w1763_,
		_w1768_,
		_w1782_
	);
	LUT3 #(
		.INIT('h82)
	) name823 (
		\wb_sel_i[1]_pad ,
		_w1774_,
		_w1779_,
		_w1783_
	);
	LUT4 #(
		.INIT('h0880)
	) name824 (
		\wb_sel_i[1]_pad ,
		_w1760_,
		_w1763_,
		_w1768_,
		_w1784_
	);
	LUT3 #(
		.INIT('h01)
	) name825 (
		_w1782_,
		_w1783_,
		_w1784_,
		_w1785_
	);
	LUT4 #(
		.INIT('h135f)
	) name826 (
		\u3_u0_r0_reg[30]/P0001 ,
		\u3_u0_r1_reg[30]/P0001 ,
		_w1752_,
		_w1753_,
		_w1786_
	);
	LUT4 #(
		.INIT('h153f)
	) name827 (
		\u3_u0_r2_reg[30]/P0001 ,
		\u3_u0_r3_reg[30]/P0001 ,
		_w1755_,
		_w1756_,
		_w1787_
	);
	LUT4 #(
		.INIT('h153f)
	) name828 (
		\u3_u0_r2_reg[29]/P0001 ,
		\u3_u0_r3_reg[29]/P0001 ,
		_w1755_,
		_w1756_,
		_w1788_
	);
	LUT4 #(
		.INIT('h135f)
	) name829 (
		\u3_u0_r0_reg[29]/P0001 ,
		\u3_u0_r1_reg[29]/P0001 ,
		_w1752_,
		_w1753_,
		_w1789_
	);
	LUT4 #(
		.INIT('h8777)
	) name830 (
		_w1786_,
		_w1787_,
		_w1788_,
		_w1789_,
		_w1790_
	);
	LUT4 #(
		.INIT('h135f)
	) name831 (
		\u3_u0_r0_reg[27]/P0001 ,
		\u3_u0_r3_reg[27]/P0001 ,
		_w1752_,
		_w1755_,
		_w1791_
	);
	LUT4 #(
		.INIT('h135f)
	) name832 (
		\u3_u0_r1_reg[27]/P0001 ,
		\u3_u0_r2_reg[27]/P0001 ,
		_w1753_,
		_w1756_,
		_w1792_
	);
	LUT2 #(
		.INIT('h8)
	) name833 (
		_w1791_,
		_w1792_,
		_w1793_
	);
	LUT4 #(
		.INIT('h135f)
	) name834 (
		\u3_u0_r0_reg[25]/P0001 ,
		\u3_u0_r1_reg[25]/P0001 ,
		_w1752_,
		_w1753_,
		_w1794_
	);
	LUT4 #(
		.INIT('h153f)
	) name835 (
		\u3_u0_r2_reg[25]/P0001 ,
		\u3_u0_r3_reg[25]/P0001 ,
		_w1755_,
		_w1756_,
		_w1795_
	);
	LUT4 #(
		.INIT('h135f)
	) name836 (
		\u3_u0_r0_reg[28]/P0001 ,
		\u3_u0_r1_reg[28]/P0001 ,
		_w1752_,
		_w1753_,
		_w1796_
	);
	LUT4 #(
		.INIT('h153f)
	) name837 (
		\u3_u0_r2_reg[28]/P0001 ,
		\u3_u0_r3_reg[28]/P0001 ,
		_w1755_,
		_w1756_,
		_w1797_
	);
	LUT4 #(
		.INIT('h7888)
	) name838 (
		_w1794_,
		_w1795_,
		_w1796_,
		_w1797_,
		_w1798_
	);
	LUT3 #(
		.INIT('h69)
	) name839 (
		_w1790_,
		_w1793_,
		_w1798_,
		_w1799_
	);
	LUT4 #(
		.INIT('h135f)
	) name840 (
		\u3_u0_r0_reg[24]/P0001 ,
		\u3_u0_r2_reg[24]/P0001 ,
		_w1752_,
		_w1756_,
		_w1800_
	);
	LUT4 #(
		.INIT('h135f)
	) name841 (
		\u3_u0_r1_reg[24]/P0001 ,
		\u3_u0_r3_reg[24]/P0001 ,
		_w1753_,
		_w1755_,
		_w1801_
	);
	LUT4 #(
		.INIT('h135f)
	) name842 (
		\u3_u0_r0_reg[31]/P0001 ,
		\u3_u0_r1_reg[31]/P0001 ,
		_w1752_,
		_w1753_,
		_w1802_
	);
	LUT4 #(
		.INIT('h153f)
	) name843 (
		\u3_u0_r2_reg[31]/P0001 ,
		\u3_u0_r3_reg[31]/P0001 ,
		_w1755_,
		_w1756_,
		_w1803_
	);
	LUT4 #(
		.INIT('h8777)
	) name844 (
		_w1800_,
		_w1801_,
		_w1802_,
		_w1803_,
		_w1804_
	);
	LUT4 #(
		.INIT('h135f)
	) name845 (
		\u3_u0_r1_reg[35]/P0001 ,
		\u3_u0_r3_reg[35]/P0001 ,
		_w1753_,
		_w1755_,
		_w1805_
	);
	LUT4 #(
		.INIT('h135f)
	) name846 (
		\u3_u0_r0_reg[35]/P0001 ,
		\u3_u0_r2_reg[35]/P0001 ,
		_w1752_,
		_w1756_,
		_w1806_
	);
	LUT4 #(
		.INIT('h135f)
	) name847 (
		\u3_u0_r0_reg[26]/P0001 ,
		\u3_u0_r1_reg[26]/P0001 ,
		_w1752_,
		_w1753_,
		_w1807_
	);
	LUT4 #(
		.INIT('h153f)
	) name848 (
		\u3_u0_r2_reg[26]/P0001 ,
		\u3_u0_r3_reg[26]/P0001 ,
		_w1755_,
		_w1756_,
		_w1808_
	);
	LUT4 #(
		.INIT('h8777)
	) name849 (
		_w1805_,
		_w1806_,
		_w1807_,
		_w1808_,
		_w1809_
	);
	LUT2 #(
		.INIT('h6)
	) name850 (
		_w1804_,
		_w1809_,
		_w1810_
	);
	LUT2 #(
		.INIT('h2)
	) name851 (
		_w1799_,
		_w1810_,
		_w1811_
	);
	LUT4 #(
		.INIT('h2002)
	) name852 (
		\wb_sel_i[3]_pad ,
		_w1790_,
		_w1793_,
		_w1798_,
		_w1812_
	);
	LUT3 #(
		.INIT('h82)
	) name853 (
		\wb_sel_i[3]_pad ,
		_w1804_,
		_w1809_,
		_w1813_
	);
	LUT4 #(
		.INIT('h0880)
	) name854 (
		\wb_sel_i[3]_pad ,
		_w1790_,
		_w1793_,
		_w1798_,
		_w1814_
	);
	LUT3 #(
		.INIT('h01)
	) name855 (
		_w1812_,
		_w1813_,
		_w1814_,
		_w1815_
	);
	LUT4 #(
		.INIT('heee0)
	) name856 (
		_w1781_,
		_w1785_,
		_w1811_,
		_w1815_,
		_w1816_
	);
	LUT4 #(
		.INIT('h135f)
	) name857 (
		\u3_u0_r0_reg[21]/P0001 ,
		\u3_u0_r1_reg[21]/P0001 ,
		_w1752_,
		_w1753_,
		_w1817_
	);
	LUT4 #(
		.INIT('h153f)
	) name858 (
		\u3_u0_r2_reg[21]/P0001 ,
		\u3_u0_r3_reg[21]/P0001 ,
		_w1755_,
		_w1756_,
		_w1818_
	);
	LUT4 #(
		.INIT('h135f)
	) name859 (
		\u3_u0_r0_reg[17]/P0001 ,
		\u3_u0_r1_reg[17]/P0001 ,
		_w1752_,
		_w1753_,
		_w1819_
	);
	LUT4 #(
		.INIT('h153f)
	) name860 (
		\u3_u0_r2_reg[17]/P0001 ,
		\u3_u0_r3_reg[17]/P0001 ,
		_w1755_,
		_w1756_,
		_w1820_
	);
	LUT4 #(
		.INIT('h8777)
	) name861 (
		_w1817_,
		_w1818_,
		_w1819_,
		_w1820_,
		_w1821_
	);
	LUT4 #(
		.INIT('h135f)
	) name862 (
		\u3_u0_r0_reg[22]/P0001 ,
		\u3_u0_r1_reg[22]/P0001 ,
		_w1752_,
		_w1753_,
		_w1822_
	);
	LUT4 #(
		.INIT('h153f)
	) name863 (
		\u3_u0_r2_reg[22]/P0001 ,
		\u3_u0_r3_reg[22]/P0001 ,
		_w1755_,
		_w1756_,
		_w1823_
	);
	LUT2 #(
		.INIT('h8)
	) name864 (
		_w1822_,
		_w1823_,
		_w1824_
	);
	LUT4 #(
		.INIT('h135f)
	) name865 (
		\u3_u0_r0_reg[19]/P0001 ,
		\u3_u0_r2_reg[19]/P0001 ,
		_w1752_,
		_w1756_,
		_w1825_
	);
	LUT4 #(
		.INIT('h135f)
	) name866 (
		\u3_u0_r1_reg[19]/P0001 ,
		\u3_u0_r3_reg[19]/P0001 ,
		_w1753_,
		_w1755_,
		_w1826_
	);
	LUT4 #(
		.INIT('h135f)
	) name867 (
		\u3_u0_r0_reg[20]/P0001 ,
		\u3_u0_r3_reg[20]/P0001 ,
		_w1752_,
		_w1755_,
		_w1827_
	);
	LUT4 #(
		.INIT('h135f)
	) name868 (
		\u3_u0_r1_reg[20]/P0001 ,
		\u3_u0_r2_reg[20]/P0001 ,
		_w1753_,
		_w1756_,
		_w1828_
	);
	LUT4 #(
		.INIT('h7888)
	) name869 (
		_w1825_,
		_w1826_,
		_w1827_,
		_w1828_,
		_w1829_
	);
	LUT3 #(
		.INIT('h69)
	) name870 (
		_w1821_,
		_w1824_,
		_w1829_,
		_w1830_
	);
	LUT4 #(
		.INIT('h135f)
	) name871 (
		\u3_u0_r0_reg[16]/P0001 ,
		\u3_u0_r1_reg[16]/P0001 ,
		_w1752_,
		_w1753_,
		_w1831_
	);
	LUT4 #(
		.INIT('h153f)
	) name872 (
		\u3_u0_r2_reg[16]/P0001 ,
		\u3_u0_r3_reg[16]/P0001 ,
		_w1755_,
		_w1756_,
		_w1832_
	);
	LUT4 #(
		.INIT('h135f)
	) name873 (
		\u3_u0_r0_reg[23]/P0001 ,
		\u3_u0_r1_reg[23]/P0001 ,
		_w1752_,
		_w1753_,
		_w1833_
	);
	LUT4 #(
		.INIT('h153f)
	) name874 (
		\u3_u0_r2_reg[23]/P0001 ,
		\u3_u0_r3_reg[23]/P0001 ,
		_w1755_,
		_w1756_,
		_w1834_
	);
	LUT4 #(
		.INIT('h8777)
	) name875 (
		_w1831_,
		_w1832_,
		_w1833_,
		_w1834_,
		_w1835_
	);
	LUT4 #(
		.INIT('h135f)
	) name876 (
		\u3_u0_r0_reg[34]/P0001 ,
		\u3_u0_r1_reg[34]/P0001 ,
		_w1752_,
		_w1753_,
		_w1836_
	);
	LUT4 #(
		.INIT('h153f)
	) name877 (
		\u3_u0_r2_reg[34]/P0001 ,
		\u3_u0_r3_reg[34]/P0001 ,
		_w1755_,
		_w1756_,
		_w1837_
	);
	LUT4 #(
		.INIT('h135f)
	) name878 (
		\u3_u0_r0_reg[18]/P0001 ,
		\u3_u0_r1_reg[18]/P0001 ,
		_w1752_,
		_w1753_,
		_w1838_
	);
	LUT4 #(
		.INIT('h153f)
	) name879 (
		\u3_u0_r2_reg[18]/P0001 ,
		\u3_u0_r3_reg[18]/P0001 ,
		_w1755_,
		_w1756_,
		_w1839_
	);
	LUT4 #(
		.INIT('h8777)
	) name880 (
		_w1836_,
		_w1837_,
		_w1838_,
		_w1839_,
		_w1840_
	);
	LUT2 #(
		.INIT('h6)
	) name881 (
		_w1835_,
		_w1840_,
		_w1841_
	);
	LUT2 #(
		.INIT('h2)
	) name882 (
		_w1830_,
		_w1841_,
		_w1842_
	);
	LUT4 #(
		.INIT('h2002)
	) name883 (
		\wb_sel_i[2]_pad ,
		_w1821_,
		_w1824_,
		_w1829_,
		_w1843_
	);
	LUT3 #(
		.INIT('h82)
	) name884 (
		\wb_sel_i[2]_pad ,
		_w1835_,
		_w1840_,
		_w1844_
	);
	LUT4 #(
		.INIT('h0880)
	) name885 (
		\wb_sel_i[2]_pad ,
		_w1821_,
		_w1824_,
		_w1829_,
		_w1845_
	);
	LUT3 #(
		.INIT('h01)
	) name886 (
		_w1843_,
		_w1844_,
		_w1845_,
		_w1846_
	);
	LUT4 #(
		.INIT('h135f)
	) name887 (
		\u3_u0_r0_reg[0]/P0001 ,
		\u3_u0_r2_reg[0]/P0001 ,
		_w1752_,
		_w1756_,
		_w1847_
	);
	LUT4 #(
		.INIT('h135f)
	) name888 (
		\u3_u0_r1_reg[0]/P0001 ,
		\u3_u0_r3_reg[0]/P0001 ,
		_w1753_,
		_w1755_,
		_w1848_
	);
	LUT4 #(
		.INIT('h135f)
	) name889 (
		\u3_u0_r0_reg[2]/P0001 ,
		\u3_u0_r1_reg[2]/P0001 ,
		_w1752_,
		_w1753_,
		_w1849_
	);
	LUT4 #(
		.INIT('h153f)
	) name890 (
		\u3_u0_r2_reg[2]/P0001 ,
		\u3_u0_r3_reg[2]/P0001 ,
		_w1755_,
		_w1756_,
		_w1850_
	);
	LUT4 #(
		.INIT('h8777)
	) name891 (
		_w1847_,
		_w1848_,
		_w1849_,
		_w1850_,
		_w1851_
	);
	LUT4 #(
		.INIT('h135f)
	) name892 (
		\u3_u0_r0_reg[4]/P0001 ,
		\u3_u0_r1_reg[4]/P0001 ,
		_w1752_,
		_w1753_,
		_w1852_
	);
	LUT4 #(
		.INIT('h153f)
	) name893 (
		\u3_u0_r2_reg[4]/P0001 ,
		\u3_u0_r3_reg[4]/P0001 ,
		_w1755_,
		_w1756_,
		_w1853_
	);
	LUT2 #(
		.INIT('h8)
	) name894 (
		_w1852_,
		_w1853_,
		_w1854_
	);
	LUT4 #(
		.INIT('h153f)
	) name895 (
		\u3_u0_r2_reg[7]/P0001 ,
		\u3_u0_r3_reg[7]/P0001 ,
		_w1755_,
		_w1756_,
		_w1855_
	);
	LUT4 #(
		.INIT('h135f)
	) name896 (
		\u3_u0_r0_reg[7]/P0001 ,
		\u3_u0_r1_reg[7]/P0001 ,
		_w1752_,
		_w1753_,
		_w1856_
	);
	LUT4 #(
		.INIT('h135f)
	) name897 (
		\u3_u0_r1_reg[6]/P0001 ,
		\u3_u0_r2_reg[6]/P0001 ,
		_w1753_,
		_w1756_,
		_w1857_
	);
	LUT4 #(
		.INIT('h135f)
	) name898 (
		\u3_u0_r0_reg[6]/P0001 ,
		\u3_u0_r3_reg[6]/P0001 ,
		_w1752_,
		_w1755_,
		_w1858_
	);
	LUT4 #(
		.INIT('h7888)
	) name899 (
		_w1855_,
		_w1856_,
		_w1857_,
		_w1858_,
		_w1859_
	);
	LUT3 #(
		.INIT('h69)
	) name900 (
		_w1851_,
		_w1854_,
		_w1859_,
		_w1860_
	);
	LUT4 #(
		.INIT('h153f)
	) name901 (
		\u3_u0_r2_reg[5]/P0001 ,
		\u3_u0_r3_reg[5]/P0001 ,
		_w1755_,
		_w1756_,
		_w1861_
	);
	LUT4 #(
		.INIT('h135f)
	) name902 (
		\u3_u0_r0_reg[5]/P0001 ,
		\u3_u0_r1_reg[5]/P0001 ,
		_w1752_,
		_w1753_,
		_w1862_
	);
	LUT4 #(
		.INIT('h135f)
	) name903 (
		\u3_u0_r0_reg[3]/P0001 ,
		\u3_u0_r2_reg[3]/P0001 ,
		_w1752_,
		_w1756_,
		_w1863_
	);
	LUT4 #(
		.INIT('h135f)
	) name904 (
		\u3_u0_r1_reg[3]/P0001 ,
		\u3_u0_r3_reg[3]/P0001 ,
		_w1753_,
		_w1755_,
		_w1864_
	);
	LUT4 #(
		.INIT('h8777)
	) name905 (
		_w1861_,
		_w1862_,
		_w1863_,
		_w1864_,
		_w1865_
	);
	LUT4 #(
		.INIT('h153f)
	) name906 (
		\u3_u0_r2_reg[32]/P0001 ,
		\u3_u0_r3_reg[32]/P0001 ,
		_w1755_,
		_w1756_,
		_w1866_
	);
	LUT4 #(
		.INIT('h135f)
	) name907 (
		\u3_u0_r0_reg[32]/P0001 ,
		\u3_u0_r1_reg[32]/P0001 ,
		_w1752_,
		_w1753_,
		_w1867_
	);
	LUT4 #(
		.INIT('h135f)
	) name908 (
		\u3_u0_r0_reg[1]/P0001 ,
		\u3_u0_r1_reg[1]/P0001 ,
		_w1752_,
		_w1753_,
		_w1868_
	);
	LUT4 #(
		.INIT('h153f)
	) name909 (
		\u3_u0_r2_reg[1]/P0001 ,
		\u3_u0_r3_reg[1]/P0001 ,
		_w1755_,
		_w1756_,
		_w1869_
	);
	LUT4 #(
		.INIT('h8777)
	) name910 (
		_w1866_,
		_w1867_,
		_w1868_,
		_w1869_,
		_w1870_
	);
	LUT2 #(
		.INIT('h6)
	) name911 (
		_w1865_,
		_w1870_,
		_w1871_
	);
	LUT2 #(
		.INIT('h2)
	) name912 (
		_w1860_,
		_w1871_,
		_w1872_
	);
	LUT4 #(
		.INIT('h2002)
	) name913 (
		\wb_sel_i[0]_pad ,
		_w1851_,
		_w1854_,
		_w1859_,
		_w1873_
	);
	LUT3 #(
		.INIT('h82)
	) name914 (
		\wb_sel_i[0]_pad ,
		_w1865_,
		_w1870_,
		_w1874_
	);
	LUT4 #(
		.INIT('h0880)
	) name915 (
		\wb_sel_i[0]_pad ,
		_w1851_,
		_w1854_,
		_w1859_,
		_w1875_
	);
	LUT3 #(
		.INIT('h01)
	) name916 (
		_w1873_,
		_w1874_,
		_w1875_,
		_w1876_
	);
	LUT4 #(
		.INIT('heee0)
	) name917 (
		_w1842_,
		_w1846_,
		_w1872_,
		_w1876_,
		_w1877_
	);
	LUT2 #(
		.INIT('h8)
	) name918 (
		_w1816_,
		_w1877_,
		_w1878_
	);
	LUT2 #(
		.INIT('h2)
	) name919 (
		\u0_csc_reg[11]/NET0131 ,
		wb_we_i_pad,
		_w1879_
	);
	LUT3 #(
		.INIT('he0)
	) name920 (
		_w1564_,
		_w1566_,
		_w1879_,
		_w1880_
	);
	LUT4 #(
		.INIT('hef00)
	) name921 (
		_w1724_,
		_w1728_,
		_w1747_,
		_w1880_,
		_w1881_
	);
	LUT2 #(
		.INIT('h1)
	) name922 (
		\u0_wp_err_reg/NET0131 ,
		\u5_state_reg[65]/NET0131 ,
		_w1882_
	);
	LUT4 #(
		.INIT('h8a00)
	) name923 (
		_w1750_,
		_w1878_,
		_w1881_,
		_w1882_,
		_w1883_
	);
	LUT3 #(
		.INIT('h08)
	) name924 (
		\wb_addr_i[29]_pad ,
		\wb_addr_i[30]_pad ,
		\wb_addr_i[31]_pad ,
		_w1884_
	);
	LUT3 #(
		.INIT('h40)
	) name925 (
		wb_ack_o_pad,
		wb_cyc_i_pad,
		wb_stb_i_pad,
		_w1885_
	);
	LUT2 #(
		.INIT('h8)
	) name926 (
		_w1884_,
		_w1885_,
		_w1886_
	);
	LUT3 #(
		.INIT('hfe)
	) name927 (
		_w1751_,
		_w1883_,
		_w1886_,
		_w1887_
	);
	LUT2 #(
		.INIT('h7)
	) name928 (
		_w1596_,
		_w1618_,
		_w1888_
	);
	LUT3 #(
		.INIT('h80)
	) name929 (
		_w1540_,
		_w1541_,
		_w1707_,
		_w1889_
	);
	LUT3 #(
		.INIT('h23)
	) name930 (
		_w1539_,
		_w1652_,
		_w1889_,
		_w1890_
	);
	LUT3 #(
		.INIT('h02)
	) name931 (
		\u0_tms_reg[11]/NET0131 ,
		\u5_lmr_ack_reg/NET0131 ,
		\u5_state_reg[26]/NET0131 ,
		_w1891_
	);
	LUT4 #(
		.INIT('h11d5)
	) name932 (
		\u0_sp_tms_reg[11]/NET0131 ,
		_w976_,
		_w1114_,
		_w1891_,
		_w1892_
	);
	LUT3 #(
		.INIT('h80)
	) name933 (
		_w1540_,
		_w1541_,
		_w1892_,
		_w1893_
	);
	LUT4 #(
		.INIT('hc8cc)
	) name934 (
		_w1539_,
		_w1652_,
		_w1662_,
		_w1893_,
		_w1894_
	);
	LUT2 #(
		.INIT('h1)
	) name935 (
		_w1890_,
		_w1894_,
		_w1895_
	);
	LUT3 #(
		.INIT('h02)
	) name936 (
		\u0_tms_reg[23]/NET0131 ,
		\u5_lmr_ack_reg/NET0131 ,
		\u5_state_reg[26]/NET0131 ,
		_w1896_
	);
	LUT4 #(
		.INIT('h11d5)
	) name937 (
		\u0_sp_tms_reg[23]/NET0131 ,
		_w976_,
		_w1114_,
		_w1896_,
		_w1897_
	);
	LUT3 #(
		.INIT('h80)
	) name938 (
		_w1540_,
		_w1541_,
		_w1897_,
		_w1898_
	);
	LUT3 #(
		.INIT('h23)
	) name939 (
		_w1539_,
		_w1591_,
		_w1898_,
		_w1899_
	);
	LUT3 #(
		.INIT('h01)
	) name940 (
		\u5_state_reg[30]/NET0131 ,
		\u5_state_reg[31]/NET0131 ,
		\u5_state_reg[35]/NET0131 ,
		_w1900_
	);
	LUT2 #(
		.INIT('h8)
	) name941 (
		_w1673_,
		_w1900_,
		_w1901_
	);
	LUT4 #(
		.INIT('h63ff)
	) name942 (
		\u5_timer_reg[2]/NET0131 ,
		\u5_timer_reg[3]/NET0131 ,
		_w1679_,
		_w1901_,
		_w1902_
	);
	LUT3 #(
		.INIT('h02)
	) name943 (
		\u0_tms_reg[27]/NET0131 ,
		\u5_lmr_ack_reg/NET0131 ,
		\u5_state_reg[26]/NET0131 ,
		_w1903_
	);
	LUT4 #(
		.INIT('h11d5)
	) name944 (
		\u0_sp_tms_reg[27]/NET0131 ,
		_w976_,
		_w1114_,
		_w1903_,
		_w1904_
	);
	LUT3 #(
		.INIT('h80)
	) name945 (
		_w1540_,
		_w1541_,
		_w1904_,
		_w1905_
	);
	LUT4 #(
		.INIT('hd0c0)
	) name946 (
		_w1539_,
		_w1673_,
		_w1902_,
		_w1905_,
		_w1906_
	);
	LUT3 #(
		.INIT('h01)
	) name947 (
		\u5_state_reg[13]/NET0131 ,
		\u5_state_reg[14]/NET0131 ,
		\u5_state_reg[9]/NET0131 ,
		_w1907_
	);
	LUT4 #(
		.INIT('hbf00)
	) name948 (
		\u5_wb_wait_r_reg/P0001 ,
		_w1100_,
		_w1161_,
		_w1907_,
		_w1908_
	);
	LUT2 #(
		.INIT('h8)
	) name949 (
		_w1591_,
		_w1908_,
		_w1909_
	);
	LUT4 #(
		.INIT('h8a88)
	) name950 (
		_w1667_,
		_w1899_,
		_w1906_,
		_w1909_,
		_w1910_
	);
	LUT3 #(
		.INIT('hab)
	) name951 (
		_w1539_,
		_w1694_,
		_w1898_,
		_w1911_
	);
	LUT3 #(
		.INIT('h45)
	) name952 (
		_w1696_,
		_w1713_,
		_w1911_,
		_w1912_
	);
	LUT3 #(
		.INIT('h40)
	) name953 (
		_w1539_,
		_w1694_,
		_w1898_,
		_w1913_
	);
	LUT3 #(
		.INIT('h40)
	) name954 (
		_w1539_,
		_w1703_,
		_w1898_,
		_w1914_
	);
	LUT4 #(
		.INIT('h080a)
	) name955 (
		_w1667_,
		_w1712_,
		_w1913_,
		_w1914_,
		_w1915_
	);
	LUT3 #(
		.INIT('h02)
	) name956 (
		\u0_tms_reg[3]/NET0131 ,
		\u5_lmr_ack_reg/NET0131 ,
		\u5_state_reg[26]/NET0131 ,
		_w1916_
	);
	LUT4 #(
		.INIT('h11d5)
	) name957 (
		\u0_sp_tms_reg[3]/NET0131 ,
		_w976_,
		_w1114_,
		_w1916_,
		_w1917_
	);
	LUT3 #(
		.INIT('h80)
	) name958 (
		_w1540_,
		_w1541_,
		_w1917_,
		_w1918_
	);
	LUT4 #(
		.INIT('hc4c0)
	) name959 (
		_w1539_,
		_w1662_,
		_w1667_,
		_w1918_,
		_w1919_
	);
	LUT2 #(
		.INIT('h4)
	) name960 (
		_w1890_,
		_w1919_,
		_w1920_
	);
	LUT4 #(
		.INIT('h1500)
	) name961 (
		_w1910_,
		_w1912_,
		_w1915_,
		_w1920_,
		_w1921_
	);
	LUT2 #(
		.INIT('h1)
	) name962 (
		_w1895_,
		_w1921_,
		_w1922_
	);
	LUT4 #(
		.INIT('ha8aa)
	) name963 (
		\u5_state_reg[16]/NET0131 ,
		_w1568_,
		_w1600_,
		_w1612_,
		_w1923_
	);
	LUT3 #(
		.INIT('h20)
	) name964 (
		_w1141_,
		_w1613_,
		_w1923_,
		_w1924_
	);
	LUT2 #(
		.INIT('h1)
	) name965 (
		\u5_wb_cycle_reg/NET0131 ,
		_w1116_,
		_w1925_
	);
	LUT4 #(
		.INIT('h4000)
	) name966 (
		\u5_wb_cycle_reg/NET0131 ,
		_w1122_,
		_w1124_,
		_w1127_,
		_w1926_
	);
	LUT2 #(
		.INIT('h1)
	) name967 (
		_w1925_,
		_w1926_,
		_w1927_
	);
	LUT4 #(
		.INIT('h0400)
	) name968 (
		\u5_wb_write_go_r_reg/NET0131 ,
		\u6_read_go_r1_reg/NET0131 ,
		\u6_rmw_r_reg/NET0131 ,
		wb_cyc_i_pad,
		_w1928_
	);
	LUT3 #(
		.INIT('h70)
	) name969 (
		_w1014_,
		_w1015_,
		_w1928_,
		_w1929_
	);
	LUT4 #(
		.INIT('h80aa)
	) name970 (
		\u5_state_reg[16]/NET0131 ,
		_w1014_,
		_w1015_,
		_w1928_,
		_w1930_
	);
	LUT2 #(
		.INIT('h4)
	) name971 (
		_w1608_,
		_w1930_,
		_w1931_
	);
	LUT4 #(
		.INIT('hb000)
	) name972 (
		_w1539_,
		_w1599_,
		_w1927_,
		_w1931_,
		_w1932_
	);
	LUT3 #(
		.INIT('h01)
	) name973 (
		\u5_ap_en_reg/NET0131 ,
		_w1925_,
		_w1926_,
		_w1933_
	);
	LUT4 #(
		.INIT('hf400)
	) name974 (
		_w1539_,
		_w1599_,
		_w1608_,
		_w1933_,
		_w1934_
	);
	LUT4 #(
		.INIT('h004f)
	) name975 (
		_w1539_,
		_w1599_,
		_w1611_,
		_w1615_,
		_w1935_
	);
	LUT4 #(
		.INIT('ha800)
	) name976 (
		_w1141_,
		_w1932_,
		_w1934_,
		_w1935_,
		_w1936_
	);
	LUT2 #(
		.INIT('h2)
	) name977 (
		_w1601_,
		_w1608_,
		_w1937_
	);
	LUT4 #(
		.INIT('h1033)
	) name978 (
		_w1539_,
		_w1564_,
		_w1599_,
		_w1937_,
		_w1938_
	);
	LUT4 #(
		.INIT('h0400)
	) name979 (
		\u5_ap_en_reg/NET0131 ,
		\u5_cmd_asserted_reg/NET0131 ,
		\u5_state_reg[12]/NET0131 ,
		\u5_state_reg[13]/NET0131 ,
		_w1939_
	);
	LUT4 #(
		.INIT('h4000)
	) name980 (
		\u5_wb_cycle_reg/NET0131 ,
		_w1002_,
		_w1143_,
		_w1939_,
		_w1940_
	);
	LUT4 #(
		.INIT('h0800)
	) name981 (
		_w1002_,
		_w1143_,
		_w1608_,
		_w1939_,
		_w1941_
	);
	LUT4 #(
		.INIT('h040f)
	) name982 (
		_w1539_,
		_w1599_,
		_w1940_,
		_w1941_,
		_w1942_
	);
	LUT2 #(
		.INIT('h8)
	) name983 (
		\u5_mem_ack_r_reg/NET0131 ,
		\u5_state_reg[16]/NET0131 ,
		_w1943_
	);
	LUT3 #(
		.INIT('h08)
	) name984 (
		\u5_state_reg[16]/NET0131 ,
		wb_cyc_i_pad,
		wb_stb_i_pad,
		_w1944_
	);
	LUT4 #(
		.INIT('h010f)
	) name985 (
		_w1564_,
		_w1566_,
		_w1943_,
		_w1944_,
		_w1945_
	);
	LUT3 #(
		.INIT('h15)
	) name986 (
		\u5_ap_en_reg/NET0131 ,
		_w976_,
		_w1118_,
		_w1946_
	);
	LUT2 #(
		.INIT('h4)
	) name987 (
		_w1117_,
		_w1946_,
		_w1947_
	);
	LUT2 #(
		.INIT('h2)
	) name988 (
		_w1945_,
		_w1947_,
		_w1948_
	);
	LUT2 #(
		.INIT('h1)
	) name989 (
		_w1564_,
		_w1735_,
		_w1949_
	);
	LUT3 #(
		.INIT('ha8)
	) name990 (
		_w1258_,
		_w1564_,
		_w1735_,
		_w1950_
	);
	LUT3 #(
		.INIT('h80)
	) name991 (
		_w1002_,
		_w1143_,
		_w1950_,
		_w1951_
	);
	LUT3 #(
		.INIT('h80)
	) name992 (
		\u5_cmd_asserted_reg/NET0131 ,
		_w1100_,
		_w1158_,
		_w1952_
	);
	LUT3 #(
		.INIT('h80)
	) name993 (
		\u5_tmr_done_reg/NET0131 ,
		_w976_,
		_w1118_,
		_w1953_
	);
	LUT2 #(
		.INIT('h8)
	) name994 (
		\u0_sp_csc_reg[10]/NET0131 ,
		\u5_tmr_done_reg/NET0131 ,
		_w1954_
	);
	LUT3 #(
		.INIT('h70)
	) name995 (
		_w976_,
		_w1114_,
		_w1954_,
		_w1955_
	);
	LUT2 #(
		.INIT('h1)
	) name996 (
		_w1953_,
		_w1955_,
		_w1956_
	);
	LUT2 #(
		.INIT('h8)
	) name997 (
		\u5_cmd_asserted_reg/NET0131 ,
		\u5_tmr_done_reg/NET0131 ,
		_w1957_
	);
	LUT3 #(
		.INIT('h70)
	) name998 (
		_w976_,
		_w1118_,
		_w1957_,
		_w1958_
	);
	LUT3 #(
		.INIT('h8a)
	) name999 (
		\u5_state_reg[16]/NET0131 ,
		_w1117_,
		_w1958_,
		_w1959_
	);
	LUT4 #(
		.INIT('h8000)
	) name1000 (
		_w1100_,
		_w1277_,
		_w1956_,
		_w1959_,
		_w1960_
	);
	LUT4 #(
		.INIT('h000b)
	) name1001 (
		_w1948_,
		_w1951_,
		_w1952_,
		_w1960_,
		_w1961_
	);
	LUT3 #(
		.INIT('hd0)
	) name1002 (
		_w1938_,
		_w1942_,
		_w1961_,
		_w1962_
	);
	LUT3 #(
		.INIT('hef)
	) name1003 (
		_w1924_,
		_w1936_,
		_w1962_,
		_w1963_
	);
	LUT3 #(
		.INIT('h2a)
	) name1004 (
		\u0_sp_csc_reg[7]/NET0131 ,
		_w976_,
		_w1114_,
		_w1964_
	);
	LUT3 #(
		.INIT('h02)
	) name1005 (
		\u0_csc_reg[7]/NET0131 ,
		\u5_lmr_ack_reg/NET0131 ,
		\u5_state_reg[26]/NET0131 ,
		_w1965_
	);
	LUT4 #(
		.INIT('h11d5)
	) name1006 (
		\u0_sp_csc_reg[7]/NET0131 ,
		_w976_,
		_w1114_,
		_w1965_,
		_w1966_
	);
	LUT3 #(
		.INIT('h02)
	) name1007 (
		\u0_csc_reg[6]/NET0131 ,
		\u5_lmr_ack_reg/NET0131 ,
		\u5_state_reg[26]/NET0131 ,
		_w1967_
	);
	LUT4 #(
		.INIT('h11d5)
	) name1008 (
		\u0_sp_csc_reg[6]/NET0131 ,
		_w976_,
		_w1114_,
		_w1967_,
		_w1968_
	);
	LUT2 #(
		.INIT('h8)
	) name1009 (
		_w1966_,
		_w1968_,
		_w1969_
	);
	LUT3 #(
		.INIT('h2a)
	) name1010 (
		\u0_sp_csc_reg[4]/NET0131 ,
		_w976_,
		_w1114_,
		_w1970_
	);
	LUT3 #(
		.INIT('h02)
	) name1011 (
		\u0_csc_reg[4]/NET0131 ,
		\u5_lmr_ack_reg/NET0131 ,
		\u5_state_reg[26]/NET0131 ,
		_w1971_
	);
	LUT4 #(
		.INIT('h11d5)
	) name1012 (
		\u0_sp_csc_reg[4]/NET0131 ,
		_w976_,
		_w1114_,
		_w1971_,
		_w1972_
	);
	LUT3 #(
		.INIT('h08)
	) name1013 (
		_w1966_,
		_w1968_,
		_w1972_,
		_w1973_
	);
	LUT3 #(
		.INIT('h2a)
	) name1014 (
		\u0_sp_csc_reg[5]/NET0131 ,
		_w976_,
		_w1114_,
		_w1974_
	);
	LUT3 #(
		.INIT('h02)
	) name1015 (
		\u0_csc_reg[5]/NET0131 ,
		\u5_lmr_ack_reg/NET0131 ,
		\u5_state_reg[26]/NET0131 ,
		_w1975_
	);
	LUT4 #(
		.INIT('h11d5)
	) name1016 (
		\u0_sp_csc_reg[5]/NET0131 ,
		_w976_,
		_w1114_,
		_w1975_,
		_w1976_
	);
	LUT4 #(
		.INIT('hf700)
	) name1017 (
		_w1966_,
		_w1968_,
		_w1972_,
		_w1976_,
		_w1977_
	);
	LUT2 #(
		.INIT('h2)
	) name1018 (
		\u5_state_reg[1]/NET0131 ,
		_w1977_,
		_w1978_
	);
	LUT3 #(
		.INIT('hb0)
	) name1019 (
		_w1539_,
		_w1668_,
		_w1978_,
		_w1979_
	);
	LUT3 #(
		.INIT('h80)
	) name1020 (
		\u5_wr_cycle_reg/NET0131 ,
		_w1732_,
		_w1746_,
		_w1980_
	);
	LUT3 #(
		.INIT('h80)
	) name1021 (
		_w1603_,
		_w1604_,
		_w1606_,
		_w1981_
	);
	LUT4 #(
		.INIT('hfe00)
	) name1022 (
		\u5_wr_cycle_reg/NET0131 ,
		_w998_,
		_w1010_,
		_w1981_,
		_w1982_
	);
	LUT4 #(
		.INIT('hef00)
	) name1023 (
		_w1724_,
		_w1728_,
		_w1980_,
		_w1982_,
		_w1983_
	);
	LUT3 #(
		.INIT('h40)
	) name1024 (
		\u5_burst_cnt_reg[7]/NET0131 ,
		_w1603_,
		_w1604_,
		_w1984_
	);
	LUT4 #(
		.INIT('hfe00)
	) name1025 (
		\u5_wr_cycle_reg/NET0131 ,
		_w998_,
		_w1010_,
		_w1984_,
		_w1985_
	);
	LUT4 #(
		.INIT('hef00)
	) name1026 (
		_w1724_,
		_w1728_,
		_w1980_,
		_w1985_,
		_w1986_
	);
	LUT4 #(
		.INIT('hcfcd)
	) name1027 (
		\u5_burst_cnt_reg[8]/NET0131 ,
		\u5_state_reg[1]/NET0131 ,
		_w1983_,
		_w1986_,
		_w1987_
	);
	LUT3 #(
		.INIT('h45)
	) name1028 (
		\u5_state_reg[52]/NET0131 ,
		_w1979_,
		_w1987_,
		_w1988_
	);
	LUT4 #(
		.INIT('hfe00)
	) name1029 (
		\u5_wr_cycle_reg/NET0131 ,
		_w998_,
		_w1010_,
		_w1608_,
		_w1989_
	);
	LUT4 #(
		.INIT('hef00)
	) name1030 (
		_w1724_,
		_w1728_,
		_w1980_,
		_w1989_,
		_w1990_
	);
	LUT4 #(
		.INIT('h4000)
	) name1031 (
		\u5_burst_cnt_reg[9]/NET0131 ,
		_w1603_,
		_w1604_,
		_w1606_,
		_w1991_
	);
	LUT4 #(
		.INIT('hfe00)
	) name1032 (
		\u5_wr_cycle_reg/NET0131 ,
		_w998_,
		_w1010_,
		_w1991_,
		_w1992_
	);
	LUT4 #(
		.INIT('hef00)
	) name1033 (
		_w1724_,
		_w1728_,
		_w1980_,
		_w1992_,
		_w1993_
	);
	LUT4 #(
		.INIT('hcfcd)
	) name1034 (
		\u5_burst_cnt_reg[10]/NET0131 ,
		\u5_state_reg[1]/NET0131 ,
		_w1990_,
		_w1993_,
		_w1994_
	);
	LUT2 #(
		.INIT('h8)
	) name1035 (
		_w1972_,
		_w1976_,
		_w1995_
	);
	LUT4 #(
		.INIT('h7000)
	) name1036 (
		_w1966_,
		_w1968_,
		_w1972_,
		_w1976_,
		_w1996_
	);
	LUT2 #(
		.INIT('h8)
	) name1037 (
		\u5_state_reg[1]/NET0131 ,
		_w1996_,
		_w1997_
	);
	LUT3 #(
		.INIT('hb0)
	) name1038 (
		_w1539_,
		_w1668_,
		_w1997_,
		_w1998_
	);
	LUT3 #(
		.INIT('h51)
	) name1039 (
		\u5_state_reg[52]/NET0131 ,
		_w1994_,
		_w1998_,
		_w1999_
	);
	LUT2 #(
		.INIT('h8)
	) name1040 (
		\u5_state_reg[1]/NET0131 ,
		_w1127_,
		_w2000_
	);
	LUT3 #(
		.INIT('h80)
	) name1041 (
		_w1540_,
		_w1541_,
		_w2000_,
		_w2001_
	);
	LUT4 #(
		.INIT('h0400)
	) name1042 (
		\u5_state_reg[52]/NET0131 ,
		_w1125_,
		_w1539_,
		_w2001_,
		_w2002_
	);
	LUT4 #(
		.INIT('h5554)
	) name1043 (
		\u5_burst_cnt_reg[0]/NET0131 ,
		\u5_wr_cycle_reg/NET0131 ,
		_w998_,
		_w1010_,
		_w2003_
	);
	LUT4 #(
		.INIT('hef00)
	) name1044 (
		_w1724_,
		_w1728_,
		_w1980_,
		_w2003_,
		_w2004_
	);
	LUT4 #(
		.INIT('h0002)
	) name1045 (
		\u5_burst_cnt_reg[0]/NET0131 ,
		\u5_wr_cycle_reg/NET0131 ,
		_w998_,
		_w1010_,
		_w2005_
	);
	LUT4 #(
		.INIT('h20aa)
	) name1046 (
		\u5_burst_cnt_reg[0]/NET0131 ,
		_w1539_,
		_w1599_,
		_w1723_,
		_w2006_
	);
	LUT4 #(
		.INIT('h0b0f)
	) name1047 (
		_w1728_,
		_w1980_,
		_w2005_,
		_w2006_,
		_w2007_
	);
	LUT2 #(
		.INIT('h1)
	) name1048 (
		\u5_state_reg[1]/NET0131 ,
		\u5_state_reg[52]/NET0131 ,
		_w2008_
	);
	LUT4 #(
		.INIT('hefaa)
	) name1049 (
		_w2002_,
		_w2004_,
		_w2007_,
		_w2008_,
		_w2009_
	);
	LUT2 #(
		.INIT('h1)
	) name1050 (
		\u5_state_reg[17]/NET0131 ,
		\u5_tmr_done_reg/NET0131 ,
		_w2010_
	);
	LUT2 #(
		.INIT('h4)
	) name1051 (
		\u5_rfr_ack_r_reg/NET0131 ,
		\u5_tmr_done_reg/NET0131 ,
		_w2011_
	);
	LUT3 #(
		.INIT('h08)
	) name1052 (
		_w982_,
		_w1181_,
		_w2011_,
		_w2012_
	);
	LUT4 #(
		.INIT('h153f)
	) name1053 (
		_w1002_,
		_w1035_,
		_w1168_,
		_w2012_,
		_w2013_
	);
	LUT3 #(
		.INIT('h40)
	) name1054 (
		\u5_cmd_asserted_reg/NET0131 ,
		_w1100_,
		_w1102_,
		_w2014_
	);
	LUT3 #(
		.INIT('hf1)
	) name1055 (
		_w2010_,
		_w2013_,
		_w2014_,
		_w2015_
	);
	LUT4 #(
		.INIT('h0001)
	) name1056 (
		\wb_addr_i[29]_pad ,
		\wb_addr_i[30]_pad ,
		\wb_addr_i[31]_pad ,
		wb_err_o_pad,
		_w2016_
	);
	LUT2 #(
		.INIT('h8)
	) name1057 (
		_w1013_,
		_w2016_,
		_w2017_
	);
	LUT4 #(
		.INIT('h4f00)
	) name1058 (
		_w1878_,
		_w1881_,
		_w1882_,
		_w2017_,
		_w2018_
	);
	LUT4 #(
		.INIT('h222a)
	) name1059 (
		\u5_lookup_ready2_reg/NET0131 ,
		_w1132_,
		_w1564_,
		_w1566_,
		_w2019_
	);
	LUT3 #(
		.INIT('h4c)
	) name1060 (
		_w1333_,
		_w1335_,
		_w1338_,
		_w2020_
	);
	LUT4 #(
		.INIT('h0b3b)
	) name1061 (
		\u5_lookup_ready2_reg/NET0131 ,
		_w1339_,
		_w1568_,
		_w2020_,
		_w2021_
	);
	LUT2 #(
		.INIT('h4)
	) name1062 (
		\u5_cmd_asserted2_reg/NET0131 ,
		\u7_mc_br_r_reg/P0001 ,
		_w2022_
	);
	LUT4 #(
		.INIT('h4f00)
	) name1063 (
		_w1533_,
		_w1579_,
		_w1580_,
		_w2022_,
		_w2023_
	);
	LUT4 #(
		.INIT('h084c)
	) name1064 (
		_w1581_,
		_w1586_,
		_w2021_,
		_w2022_,
		_w2024_
	);
	LUT3 #(
		.INIT('h08)
	) name1065 (
		_w1100_,
		_w1277_,
		_w1956_,
		_w2025_
	);
	LUT2 #(
		.INIT('h1)
	) name1066 (
		\u5_state_reg[1]/NET0131 ,
		\u5_tmr_done_reg/NET0131 ,
		_w2026_
	);
	LUT4 #(
		.INIT('h153f)
	) name1067 (
		_w1002_,
		_w1184_,
		_w1206_,
		_w1274_,
		_w2027_
	);
	LUT3 #(
		.INIT('h08)
	) name1068 (
		\u5_wb_cycle_reg/NET0131 ,
		wb_cyc_i_pad,
		wb_stb_i_pad,
		_w2028_
	);
	LUT4 #(
		.INIT('he0f0)
	) name1069 (
		\u5_cs_le_r_reg/P0001 ,
		\u5_state_reg[1]/NET0131 ,
		\u5_tmr2_done_reg/NET0131 ,
		\u5_wb_cycle_reg/NET0131 ,
		_w2029_
	);
	LUT4 #(
		.INIT('h1f00)
	) name1070 (
		_w1564_,
		_w1566_,
		_w2028_,
		_w2029_,
		_w2030_
	);
	LUT3 #(
		.INIT('h80)
	) name1071 (
		_w1002_,
		_w1166_,
		_w2030_,
		_w2031_
	);
	LUT4 #(
		.INIT('h0054)
	) name1072 (
		_w1095_,
		_w2026_,
		_w2027_,
		_w2031_,
		_w2032_
	);
	LUT3 #(
		.INIT('hef)
	) name1073 (
		_w2024_,
		_w2025_,
		_w2032_,
		_w2033_
	);
	LUT4 #(
		.INIT('hfe00)
	) name1074 (
		\u5_wr_cycle_reg/NET0131 ,
		_w998_,
		_w1010_,
		_w1603_,
		_w2034_
	);
	LUT4 #(
		.INIT('hef00)
	) name1075 (
		_w1724_,
		_w1728_,
		_w1980_,
		_w2034_,
		_w2035_
	);
	LUT4 #(
		.INIT('hfe00)
	) name1076 (
		\u5_wr_cycle_reg/NET0131 ,
		_w998_,
		_w1010_,
		_w1602_,
		_w2036_
	);
	LUT4 #(
		.INIT('hef00)
	) name1077 (
		_w1724_,
		_w1728_,
		_w1980_,
		_w2036_,
		_w2037_
	);
	LUT4 #(
		.INIT('hcfcd)
	) name1078 (
		\u5_burst_cnt_reg[2]/NET0131 ,
		\u5_state_reg[1]/NET0131 ,
		_w2035_,
		_w2037_,
		_w2038_
	);
	LUT2 #(
		.INIT('h4)
	) name1079 (
		_w1122_,
		_w1124_,
		_w2039_
	);
	LUT3 #(
		.INIT('h80)
	) name1080 (
		_w1540_,
		_w1541_,
		_w2039_,
		_w2040_
	);
	LUT4 #(
		.INIT('h4555)
	) name1081 (
		\u5_state_reg[52]/NET0131 ,
		_w1539_,
		_w2001_,
		_w2040_,
		_w2041_
	);
	LUT2 #(
		.INIT('h7)
	) name1082 (
		_w2038_,
		_w2041_,
		_w2042_
	);
	LUT4 #(
		.INIT('h8707)
	) name1083 (
		_w1966_,
		_w1968_,
		_w1972_,
		_w1976_,
		_w2043_
	);
	LUT2 #(
		.INIT('h8)
	) name1084 (
		\u5_state_reg[1]/NET0131 ,
		_w2043_,
		_w2044_
	);
	LUT3 #(
		.INIT('hb0)
	) name1085 (
		_w1539_,
		_w1668_,
		_w2044_,
		_w2045_
	);
	LUT4 #(
		.INIT('h00ed)
	) name1086 (
		\u5_burst_cnt_reg[9]/NET0131 ,
		\u5_state_reg[1]/NET0131 ,
		_w1983_,
		_w2045_,
		_w2046_
	);
	LUT2 #(
		.INIT('h1)
	) name1087 (
		\u5_state_reg[52]/NET0131 ,
		_w2046_,
		_w2047_
	);
	LUT3 #(
		.INIT('h51)
	) name1088 (
		\u5_data_oe_reg/NET0131 ,
		\u5_wb_cycle_reg/NET0131 ,
		\u5_wr_cycle_reg/NET0131 ,
		_w2048_
	);
	LUT3 #(
		.INIT('h31)
	) name1089 (
		\u5_data_oe_reg/NET0131 ,
		\u5_susp_sel_r_reg/NET0131 ,
		\u7_mc_dqm_r2_reg[0]/P0001 ,
		_w2049_
	);
	LUT2 #(
		.INIT('hb)
	) name1090 (
		_w2048_,
		_w2049_,
		_w2050_
	);
	LUT3 #(
		.INIT('h31)
	) name1091 (
		\u5_data_oe_reg/NET0131 ,
		\u5_susp_sel_r_reg/NET0131 ,
		\u7_mc_dqm_r2_reg[1]/P0001 ,
		_w2051_
	);
	LUT2 #(
		.INIT('hb)
	) name1092 (
		_w2048_,
		_w2051_,
		_w2052_
	);
	LUT3 #(
		.INIT('h31)
	) name1093 (
		\u5_data_oe_reg/NET0131 ,
		\u5_susp_sel_r_reg/NET0131 ,
		\u7_mc_dqm_r2_reg[2]/P0001 ,
		_w2053_
	);
	LUT2 #(
		.INIT('hb)
	) name1094 (
		_w2048_,
		_w2053_,
		_w2054_
	);
	LUT3 #(
		.INIT('h31)
	) name1095 (
		\u5_data_oe_reg/NET0131 ,
		\u5_susp_sel_r_reg/NET0131 ,
		\u7_mc_dqm_r2_reg[3]/P0001 ,
		_w2055_
	);
	LUT2 #(
		.INIT('hb)
	) name1096 (
		_w2048_,
		_w2055_,
		_w2056_
	);
	LUT4 #(
		.INIT('hfd01)
	) name1097 (
		\u5_state_reg[2]/NET0131 ,
		_w1613_,
		_w1614_,
		_w1927_,
		_w2057_
	);
	LUT2 #(
		.INIT('h2)
	) name1098 (
		_w1141_,
		_w2057_,
		_w2058_
	);
	LUT4 #(
		.INIT('h5510)
	) name1099 (
		\u5_ap_en_reg/NET0131 ,
		_w1539_,
		_w1599_,
		_w1608_,
		_w2059_
	);
	LUT4 #(
		.INIT('h4055)
	) name1100 (
		\u5_state_reg[2]/NET0131 ,
		_w1014_,
		_w1015_,
		_w1928_,
		_w2060_
	);
	LUT2 #(
		.INIT('h4)
	) name1101 (
		_w1608_,
		_w2060_,
		_w2061_
	);
	LUT3 #(
		.INIT('hb0)
	) name1102 (
		_w1539_,
		_w1599_,
		_w2061_,
		_w2062_
	);
	LUT4 #(
		.INIT('h0008)
	) name1103 (
		_w1141_,
		_w1935_,
		_w2059_,
		_w2062_,
		_w2063_
	);
	LUT3 #(
		.INIT('h80)
	) name1104 (
		_w1002_,
		_w1143_,
		_w1720_,
		_w2064_
	);
	LUT4 #(
		.INIT('haa20)
	) name1105 (
		\u5_wb_cycle_reg/NET0131 ,
		_w1539_,
		_w1599_,
		_w1608_,
		_w2065_
	);
	LUT2 #(
		.INIT('h2)
	) name1106 (
		\u5_ap_en_reg/NET0131 ,
		_w1564_,
		_w2066_
	);
	LUT4 #(
		.INIT('h4f00)
	) name1107 (
		_w1539_,
		_w1599_,
		_w1937_,
		_w2066_,
		_w2067_
	);
	LUT3 #(
		.INIT('ha8)
	) name1108 (
		_w2064_,
		_w2065_,
		_w2067_,
		_w2068_
	);
	LUT2 #(
		.INIT('h2)
	) name1109 (
		\u5_mem_ack_r_reg/NET0131 ,
		\u5_state_reg[2]/NET0131 ,
		_w2069_
	);
	LUT3 #(
		.INIT('h04)
	) name1110 (
		\u5_state_reg[2]/NET0131 ,
		wb_cyc_i_pad,
		wb_stb_i_pad,
		_w2070_
	);
	LUT4 #(
		.INIT('h010f)
	) name1111 (
		_w1564_,
		_w1566_,
		_w2069_,
		_w2070_,
		_w2071_
	);
	LUT2 #(
		.INIT('h4)
	) name1112 (
		_w1947_,
		_w2071_,
		_w2072_
	);
	LUT2 #(
		.INIT('h8)
	) name1113 (
		_w1951_,
		_w2072_,
		_w2073_
	);
	LUT4 #(
		.INIT('h337f)
	) name1114 (
		\u5_tmr_done_reg/NET0131 ,
		_w1059_,
		_w1086_,
		_w1252_,
		_w2074_
	);
	LUT2 #(
		.INIT('h4)
	) name1115 (
		\u5_state_reg[2]/NET0131 ,
		\u7_mc_br_r_reg/P0001 ,
		_w2075_
	);
	LUT3 #(
		.INIT('h08)
	) name1116 (
		_w1041_,
		_w1256_,
		_w2075_,
		_w2076_
	);
	LUT3 #(
		.INIT('h45)
	) name1117 (
		\u5_state_reg[2]/NET0131 ,
		_w1117_,
		_w1958_,
		_w2077_
	);
	LUT4 #(
		.INIT('h0080)
	) name1118 (
		_w1100_,
		_w1277_,
		_w1956_,
		_w2077_,
		_w2078_
	);
	LUT3 #(
		.INIT('h02)
	) name1119 (
		_w2074_,
		_w2076_,
		_w2078_,
		_w2079_
	);
	LUT2 #(
		.INIT('h4)
	) name1120 (
		_w2073_,
		_w2079_,
		_w2080_
	);
	LUT4 #(
		.INIT('h0302)
	) name1121 (
		\u5_tmr_done_reg/NET0131 ,
		_w1156_,
		_w1192_,
		_w1320_,
		_w2081_
	);
	LUT4 #(
		.INIT('h153f)
	) name1122 (
		_w1068_,
		_w1100_,
		_w1102_,
		_w1155_,
		_w2082_
	);
	LUT3 #(
		.INIT('h8a)
	) name1123 (
		\u5_cmd_asserted_reg/NET0131 ,
		_w1192_,
		_w2082_,
		_w2083_
	);
	LUT3 #(
		.INIT('h0d)
	) name1124 (
		\u5_state_reg[2]/NET0131 ,
		_w2081_,
		_w2083_,
		_w2084_
	);
	LUT2 #(
		.INIT('h8)
	) name1125 (
		_w2080_,
		_w2084_,
		_w2085_
	);
	LUT4 #(
		.INIT('hfeff)
	) name1126 (
		_w2058_,
		_w2063_,
		_w2068_,
		_w2085_,
		_w2086_
	);
	LUT3 #(
		.INIT('h08)
	) name1127 (
		_w1059_,
		_w1189_,
		_w1571_,
		_w2087_
	);
	LUT3 #(
		.INIT('h08)
	) name1128 (
		\u5_state_reg[57]/NET0131 ,
		wb_cyc_i_pad,
		wb_stb_i_pad,
		_w2088_
	);
	LUT4 #(
		.INIT('h0070)
	) name1129 (
		_w1014_,
		_w1015_,
		_w1565_,
		_w2088_,
		_w2089_
	);
	LUT2 #(
		.INIT('h2)
	) name1130 (
		_w1077_,
		_w2089_,
		_w2090_
	);
	LUT2 #(
		.INIT('h8)
	) name1131 (
		_w991_,
		_w2090_,
		_w2091_
	);
	LUT3 #(
		.INIT('h10)
	) name1132 (
		\u5_state_reg[57]/NET0131 ,
		\u6_rmw_r_reg/NET0131 ,
		wb_cyc_i_pad,
		_w2092_
	);
	LUT4 #(
		.INIT('h7000)
	) name1133 (
		_w1014_,
		_w1015_,
		_w1131_,
		_w2092_,
		_w2093_
	);
	LUT4 #(
		.INIT('h0057)
	) name1134 (
		_w1132_,
		_w1564_,
		_w1566_,
		_w2093_,
		_w2094_
	);
	LUT3 #(
		.INIT('h80)
	) name1135 (
		_w1059_,
		_w1742_,
		_w2094_,
		_w2095_
	);
	LUT2 #(
		.INIT('h2)
	) name1136 (
		\u5_state_reg[57]/NET0131 ,
		_w1735_,
		_w2096_
	);
	LUT2 #(
		.INIT('h2)
	) name1137 (
		_w1566_,
		_w2096_,
		_w2097_
	);
	LUT3 #(
		.INIT('h08)
	) name1138 (
		_w991_,
		_w1250_,
		_w2097_,
		_w2098_
	);
	LUT4 #(
		.INIT('hfffe)
	) name1139 (
		_w2087_,
		_w2091_,
		_w2095_,
		_w2098_,
		_w2099_
	);
	LUT4 #(
		.INIT('ha080)
	) name1140 (
		_w1059_,
		_w1189_,
		_w1568_,
		_w1742_,
		_w2100_
	);
	LUT3 #(
		.INIT('h20)
	) name1141 (
		\u5_state_reg[59]/NET0131 ,
		\u6_rmw_r_reg/NET0131 ,
		wb_cyc_i_pad,
		_w2101_
	);
	LUT4 #(
		.INIT('h7000)
	) name1142 (
		_w1014_,
		_w1015_,
		_w1131_,
		_w2101_,
		_w2102_
	);
	LUT3 #(
		.INIT('h80)
	) name1143 (
		_w1059_,
		_w1742_,
		_w2102_,
		_w2103_
	);
	LUT2 #(
		.INIT('he)
	) name1144 (
		_w2100_,
		_w2103_,
		_w2104_
	);
	LUT3 #(
		.INIT('h80)
	) name1145 (
		_w1127_,
		_w1540_,
		_w1541_,
		_w2105_
	);
	LUT4 #(
		.INIT('h080c)
	) name1146 (
		_w1539_,
		_w1662_,
		_w1667_,
		_w2105_,
		_w2106_
	);
	LUT3 #(
		.INIT('h01)
	) name1147 (
		\u0_tms_reg[24]/NET0131 ,
		\u5_lmr_ack_reg/NET0131 ,
		\u5_state_reg[26]/NET0131 ,
		_w2107_
	);
	LUT4 #(
		.INIT('h22ea)
	) name1148 (
		\u0_sp_tms_reg[24]/NET0131 ,
		_w976_,
		_w1114_,
		_w2107_,
		_w2108_
	);
	LUT2 #(
		.INIT('h1)
	) name1149 (
		_w1673_,
		_w2108_,
		_w2109_
	);
	LUT3 #(
		.INIT('h80)
	) name1150 (
		_w1540_,
		_w1541_,
		_w2109_,
		_w2110_
	);
	LUT4 #(
		.INIT('hc888)
	) name1151 (
		\u5_mc_le_reg/NET0131 ,
		\u5_timer_reg[0]/NET0131 ,
		_w1675_,
		_w1676_,
		_w2111_
	);
	LUT2 #(
		.INIT('h1)
	) name1152 (
		\u5_mc_le_reg/NET0131 ,
		\u5_timer_reg[0]/NET0131 ,
		_w2112_
	);
	LUT3 #(
		.INIT('h70)
	) name1153 (
		_w1675_,
		_w1676_,
		_w2112_,
		_w2113_
	);
	LUT3 #(
		.INIT('h02)
	) name1154 (
		_w1901_,
		_w2111_,
		_w2113_,
		_w2114_
	);
	LUT4 #(
		.INIT('h5510)
	) name1155 (
		\u5_state_reg[9]/NET0131 ,
		_w1539_,
		_w2110_,
		_w2114_,
		_w2115_
	);
	LUT3 #(
		.INIT('h02)
	) name1156 (
		\u0_tms_reg[4]/NET0131 ,
		\u5_lmr_ack_reg/NET0131 ,
		\u5_state_reg[26]/NET0131 ,
		_w2116_
	);
	LUT4 #(
		.INIT('h11d5)
	) name1157 (
		\u0_sp_tms_reg[4]/NET0131 ,
		_w976_,
		_w1114_,
		_w2116_,
		_w2117_
	);
	LUT2 #(
		.INIT('h8)
	) name1158 (
		\u5_state_reg[9]/NET0131 ,
		_w2117_,
		_w2118_
	);
	LUT3 #(
		.INIT('h80)
	) name1159 (
		_w1540_,
		_w1541_,
		_w2118_,
		_w2119_
	);
	LUT4 #(
		.INIT('h2030)
	) name1160 (
		_w1539_,
		_w1589_,
		_w1591_,
		_w2119_,
		_w2120_
	);
	LUT2 #(
		.INIT('h4)
	) name1161 (
		_w2115_,
		_w2120_,
		_w2121_
	);
	LUT3 #(
		.INIT('h80)
	) name1162 (
		_w1540_,
		_w1541_,
		_w1709_,
		_w2122_
	);
	LUT3 #(
		.INIT('h23)
	) name1163 (
		_w1539_,
		_w1591_,
		_w2122_,
		_w2123_
	);
	LUT3 #(
		.INIT('h80)
	) name1164 (
		_w1540_,
		_w1541_,
		_w1550_,
		_w2124_
	);
	LUT4 #(
		.INIT('h80c0)
	) name1165 (
		_w1539_,
		_w1589_,
		_w1591_,
		_w2124_,
		_w2125_
	);
	LUT3 #(
		.INIT('h02)
	) name1166 (
		_w1696_,
		_w2123_,
		_w2125_,
		_w2126_
	);
	LUT2 #(
		.INIT('h8)
	) name1167 (
		_w1707_,
		_w1709_,
		_w2127_
	);
	LUT3 #(
		.INIT('h80)
	) name1168 (
		_w1540_,
		_w1541_,
		_w2127_,
		_w2128_
	);
	LUT4 #(
		.INIT('h3323)
	) name1169 (
		_w1539_,
		_w1696_,
		_w1711_,
		_w2128_,
		_w2129_
	);
	LUT3 #(
		.INIT('h08)
	) name1170 (
		_w1662_,
		_w1667_,
		_w2129_,
		_w2130_
	);
	LUT4 #(
		.INIT('h1055)
	) name1171 (
		_w2106_,
		_w2121_,
		_w2126_,
		_w2130_,
		_w2131_
	);
	LUT3 #(
		.INIT('h02)
	) name1172 (
		\u0_tms_reg[8]/NET0131 ,
		\u5_lmr_ack_reg/NET0131 ,
		\u5_state_reg[26]/NET0131 ,
		_w2132_
	);
	LUT4 #(
		.INIT('h11d5)
	) name1173 (
		\u0_sp_tms_reg[8]/NET0131 ,
		_w976_,
		_w1114_,
		_w2132_,
		_w2133_
	);
	LUT3 #(
		.INIT('h80)
	) name1174 (
		_w1540_,
		_w1541_,
		_w2133_,
		_w2134_
	);
	LUT3 #(
		.INIT('h23)
	) name1175 (
		_w1539_,
		_w1662_,
		_w2134_,
		_w2135_
	);
	LUT3 #(
		.INIT('h02)
	) name1176 (
		\u0_tms_reg[12]/NET0131 ,
		\u5_lmr_ack_reg/NET0131 ,
		\u5_state_reg[26]/NET0131 ,
		_w2136_
	);
	LUT4 #(
		.INIT('h11d5)
	) name1177 (
		\u0_sp_tms_reg[12]/NET0131 ,
		_w976_,
		_w1114_,
		_w2136_,
		_w2137_
	);
	LUT3 #(
		.INIT('h80)
	) name1178 (
		_w1540_,
		_w1541_,
		_w2137_,
		_w2138_
	);
	LUT3 #(
		.INIT('h23)
	) name1179 (
		_w1539_,
		_w1652_,
		_w2138_,
		_w2139_
	);
	LUT4 #(
		.INIT('hffa2)
	) name1180 (
		_w1652_,
		_w2131_,
		_w2135_,
		_w2139_,
		_w2140_
	);
	LUT3 #(
		.INIT('h02)
	) name1181 (
		\u0_tms_reg[13]/NET0131 ,
		\u5_lmr_ack_reg/NET0131 ,
		\u5_state_reg[26]/NET0131 ,
		_w2141_
	);
	LUT4 #(
		.INIT('h11d5)
	) name1182 (
		\u0_sp_tms_reg[13]/NET0131 ,
		_w976_,
		_w1114_,
		_w2141_,
		_w2142_
	);
	LUT4 #(
		.INIT('hea00)
	) name1183 (
		_w1173_,
		_w1581_,
		_w1651_,
		_w2142_,
		_w2143_
	);
	LUT4 #(
		.INIT('hf400)
	) name1184 (
		_w1539_,
		_w1542_,
		_w1652_,
		_w2143_,
		_w2144_
	);
	LUT3 #(
		.INIT('h80)
	) name1185 (
		_w1122_,
		_w1540_,
		_w1541_,
		_w2145_
	);
	LUT4 #(
		.INIT('hc8cc)
	) name1186 (
		_w1539_,
		_w1662_,
		_w1667_,
		_w2145_,
		_w2146_
	);
	LUT4 #(
		.INIT('h080c)
	) name1187 (
		_w1539_,
		_w1662_,
		_w1667_,
		_w2145_,
		_w2147_
	);
	LUT3 #(
		.INIT('h01)
	) name1188 (
		\u0_tms_reg[25]/NET0131 ,
		\u5_lmr_ack_reg/NET0131 ,
		\u5_state_reg[26]/NET0131 ,
		_w2148_
	);
	LUT4 #(
		.INIT('h22ea)
	) name1189 (
		\u0_sp_tms_reg[25]/NET0131 ,
		_w976_,
		_w1114_,
		_w2148_,
		_w2149_
	);
	LUT2 #(
		.INIT('h1)
	) name1190 (
		_w1673_,
		_w2149_,
		_w2150_
	);
	LUT3 #(
		.INIT('h80)
	) name1191 (
		_w1540_,
		_w1541_,
		_w2150_,
		_w2151_
	);
	LUT4 #(
		.INIT('h80aa)
	) name1192 (
		\u5_timer_reg[1]/NET0131 ,
		_w1675_,
		_w1676_,
		_w2112_,
		_w2152_
	);
	LUT3 #(
		.INIT('h04)
	) name1193 (
		_w1679_,
		_w1901_,
		_w2152_,
		_w2153_
	);
	LUT4 #(
		.INIT('h5510)
	) name1194 (
		\u5_state_reg[9]/NET0131 ,
		_w1539_,
		_w2151_,
		_w2153_,
		_w2154_
	);
	LUT3 #(
		.INIT('h02)
	) name1195 (
		\u0_tms_reg[5]/NET0131 ,
		\u5_lmr_ack_reg/NET0131 ,
		\u5_state_reg[26]/NET0131 ,
		_w2155_
	);
	LUT4 #(
		.INIT('h11d5)
	) name1196 (
		\u0_sp_tms_reg[5]/NET0131 ,
		_w976_,
		_w1114_,
		_w2155_,
		_w2156_
	);
	LUT2 #(
		.INIT('h8)
	) name1197 (
		\u5_state_reg[9]/NET0131 ,
		_w2156_,
		_w2157_
	);
	LUT3 #(
		.INIT('h80)
	) name1198 (
		_w1540_,
		_w1541_,
		_w2157_,
		_w2158_
	);
	LUT4 #(
		.INIT('h2030)
	) name1199 (
		_w1539_,
		_w1589_,
		_w1591_,
		_w2158_,
		_w2159_
	);
	LUT3 #(
		.INIT('h80)
	) name1200 (
		_w1540_,
		_w1541_,
		_w1546_,
		_w2160_
	);
	LUT4 #(
		.INIT('h80c0)
	) name1201 (
		_w1539_,
		_w1589_,
		_w1591_,
		_w2160_,
		_w2161_
	);
	LUT3 #(
		.INIT('h08)
	) name1202 (
		_w1540_,
		_w1541_,
		_w1701_,
		_w2162_
	);
	LUT4 #(
		.INIT('hd0c0)
	) name1203 (
		_w1539_,
		_w1591_,
		_w1696_,
		_w2162_,
		_w2163_
	);
	LUT4 #(
		.INIT('h0b00)
	) name1204 (
		_w2154_,
		_w2159_,
		_w2161_,
		_w2163_,
		_w2164_
	);
	LUT3 #(
		.INIT('h04)
	) name1205 (
		_w1539_,
		_w1703_,
		_w1705_,
		_w2165_
	);
	LUT3 #(
		.INIT('h10)
	) name1206 (
		_w1539_,
		_w1696_,
		_w1711_,
		_w2166_
	);
	LUT3 #(
		.INIT('h23)
	) name1207 (
		_w1539_,
		_w1696_,
		_w1711_,
		_w2167_
	);
	LUT4 #(
		.INIT('h028a)
	) name1208 (
		_w2146_,
		_w2165_,
		_w2166_,
		_w2167_,
		_w2168_
	);
	LUT3 #(
		.INIT('h80)
	) name1209 (
		_w1116_,
		_w1540_,
		_w1541_,
		_w2169_
	);
	LUT4 #(
		.INIT('hc4c0)
	) name1210 (
		_w1539_,
		_w1652_,
		_w1662_,
		_w2169_,
		_w2170_
	);
	LUT2 #(
		.INIT('h4)
	) name1211 (
		_w1653_,
		_w2170_,
		_w2171_
	);
	LUT4 #(
		.INIT('h4500)
	) name1212 (
		_w2147_,
		_w2164_,
		_w2168_,
		_w2171_,
		_w2172_
	);
	LUT2 #(
		.INIT('h1)
	) name1213 (
		_w2144_,
		_w2172_,
		_w2173_
	);
	LUT4 #(
		.INIT('he222)
	) name1214 (
		\u5_state_reg[41]/NET0131 ,
		\u5_tmr2_done_reg/NET0131 ,
		_w1972_,
		_w1976_,
		_w2174_
	);
	LUT3 #(
		.INIT('h80)
	) name1215 (
		_w1041_,
		_w1195_,
		_w2174_,
		_w2175_
	);
	LUT2 #(
		.INIT('h1)
	) name1216 (
		\u5_state_reg[45]/NET0131 ,
		\u5_tmr2_done_reg/NET0131 ,
		_w2176_
	);
	LUT3 #(
		.INIT('h8a)
	) name1217 (
		\u5_tmr2_done_reg/NET0131 ,
		_w1972_,
		_w1976_,
		_w2177_
	);
	LUT3 #(
		.INIT('h08)
	) name1218 (
		_w1041_,
		_w1195_,
		_w2177_,
		_w2178_
	);
	LUT3 #(
		.INIT('h32)
	) name1219 (
		_w1237_,
		_w2176_,
		_w2178_,
		_w2179_
	);
	LUT2 #(
		.INIT('h2)
	) name1220 (
		\u5_state_reg[46]/NET0131 ,
		\u5_tmr2_done_reg/NET0131 ,
		_w2180_
	);
	LUT3 #(
		.INIT('hba)
	) name1221 (
		_w1244_,
		_w1557_,
		_w2180_,
		_w2181_
	);
	LUT4 #(
		.INIT('h0080)
	) name1222 (
		_w1135_,
		_w1333_,
		_w1335_,
		_w1338_,
		_w2182_
	);
	LUT4 #(
		.INIT('hb000)
	) name1223 (
		_w1533_,
		_w1579_,
		_w1580_,
		_w2182_,
		_w2183_
	);
	LUT4 #(
		.INIT('h8a00)
	) name1224 (
		\u5_state_reg[47]/NET0131 ,
		_w1533_,
		_w1579_,
		_w1580_,
		_w2184_
	);
	LUT3 #(
		.INIT('h8c)
	) name1225 (
		\u5_cmd_asserted2_reg/NET0131 ,
		\u5_state_reg[47]/NET0131 ,
		\u7_mc_br_r_reg/P0001 ,
		_w2185_
	);
	LUT4 #(
		.INIT('h4f00)
	) name1226 (
		_w1533_,
		_w1579_,
		_w1580_,
		_w2185_,
		_w2186_
	);
	LUT4 #(
		.INIT('h0023)
	) name1227 (
		_w2021_,
		_w2183_,
		_w2184_,
		_w2186_,
		_w2187_
	);
	LUT2 #(
		.INIT('h2)
	) name1228 (
		_w1586_,
		_w2187_,
		_w2188_
	);
	LUT3 #(
		.INIT('h04)
	) name1229 (
		\u5_cmd_asserted_reg/NET0131 ,
		\u5_state_reg[52]/NET0131 ,
		\u5_state_reg[53]/NET0131 ,
		_w2189_
	);
	LUT3 #(
		.INIT('h80)
	) name1230 (
		_w992_,
		_w999_,
		_w2189_,
		_w2190_
	);
	LUT4 #(
		.INIT('h2000)
	) name1231 (
		\u6_read_go_r1_reg/NET0131 ,
		\u6_rmw_r_reg/NET0131 ,
		wb_cyc_i_pad,
		wb_stb_i_pad,
		_w2191_
	);
	LUT3 #(
		.INIT('h70)
	) name1232 (
		_w1014_,
		_w1015_,
		_w2191_,
		_w2192_
	);
	LUT2 #(
		.INIT('h8)
	) name1233 (
		_w1077_,
		_w2192_,
		_w2193_
	);
	LUT2 #(
		.INIT('h8)
	) name1234 (
		_w991_,
		_w2193_,
		_w2194_
	);
	LUT3 #(
		.INIT('h57)
	) name1235 (
		_w991_,
		_w2190_,
		_w2193_,
		_w2195_
	);
	LUT2 #(
		.INIT('h4)
	) name1236 (
		_w1586_,
		_w2195_,
		_w2196_
	);
	LUT4 #(
		.INIT('h082a)
	) name1237 (
		\u5_state_reg[52]/NET0131 ,
		_w1581_,
		_w2021_,
		_w2022_,
		_w2197_
	);
	LUT3 #(
		.INIT('h70)
	) name1238 (
		_w1572_,
		_w1581_,
		_w2195_,
		_w2198_
	);
	LUT3 #(
		.INIT('h45)
	) name1239 (
		_w2196_,
		_w2197_,
		_w2198_,
		_w2199_
	);
	LUT3 #(
		.INIT('h04)
	) name1240 (
		\u5_cmd_asserted_reg/NET0131 ,
		\u5_state_reg[58]/NET0131 ,
		\u5_state_reg[59]/NET0131 ,
		_w2200_
	);
	LUT3 #(
		.INIT('h80)
	) name1241 (
		_w985_,
		_w986_,
		_w2200_,
		_w2201_
	);
	LUT2 #(
		.INIT('h9)
	) name1242 (
		\u5_state_reg[58]/NET0131 ,
		\u5_state_reg[59]/NET0131 ,
		_w2202_
	);
	LUT3 #(
		.INIT('h08)
	) name1243 (
		_w985_,
		_w986_,
		_w2202_,
		_w2203_
	);
	LUT4 #(
		.INIT('h575f)
	) name1244 (
		_w1059_,
		_w1135_,
		_w2201_,
		_w2203_,
		_w2204_
	);
	LUT2 #(
		.INIT('h4)
	) name1245 (
		_w1586_,
		_w2204_,
		_w2205_
	);
	LUT4 #(
		.INIT('hb000)
	) name1246 (
		_w1533_,
		_w1579_,
		_w1580_,
		_w1739_,
		_w2206_
	);
	LUT4 #(
		.INIT('h8a00)
	) name1247 (
		\u5_state_reg[58]/NET0131 ,
		_w1533_,
		_w1579_,
		_w1580_,
		_w2207_
	);
	LUT3 #(
		.INIT('h23)
	) name1248 (
		_w2021_,
		_w2206_,
		_w2207_,
		_w2208_
	);
	LUT3 #(
		.INIT('h8c)
	) name1249 (
		\u5_cmd_asserted2_reg/NET0131 ,
		\u5_state_reg[58]/NET0131 ,
		\u7_mc_br_r_reg/P0001 ,
		_w2209_
	);
	LUT4 #(
		.INIT('h4f00)
	) name1250 (
		_w1533_,
		_w1579_,
		_w1580_,
		_w2209_,
		_w2210_
	);
	LUT2 #(
		.INIT('h2)
	) name1251 (
		_w2204_,
		_w2210_,
		_w2211_
	);
	LUT3 #(
		.INIT('h15)
	) name1252 (
		_w2205_,
		_w2208_,
		_w2211_,
		_w2212_
	);
	LUT2 #(
		.INIT('h1)
	) name1253 (
		\u5_cmd_asserted_reg/NET0131 ,
		\u5_state_reg[5]/NET0131 ,
		_w2213_
	);
	LUT3 #(
		.INIT('h08)
	) name1254 (
		_w982_,
		_w1289_,
		_w2213_,
		_w2214_
	);
	LUT2 #(
		.INIT('h8)
	) name1255 (
		_w1002_,
		_w2214_,
		_w2215_
	);
	LUT4 #(
		.INIT('h135f)
	) name1256 (
		_w1002_,
		_w1068_,
		_w1182_,
		_w1201_,
		_w2216_
	);
	LUT2 #(
		.INIT('h2)
	) name1257 (
		\u5_state_reg[5]/NET0131 ,
		\u5_tmr_done_reg/NET0131 ,
		_w2217_
	);
	LUT3 #(
		.INIT('hba)
	) name1258 (
		_w2215_,
		_w2216_,
		_w2217_,
		_w2218_
	);
	LUT3 #(
		.INIT('h02)
	) name1259 (
		\u5_state_reg[60]/NET0131 ,
		\u5_tmr2_done_reg/NET0131 ,
		\u7_mc_ack_r_reg/NET0131 ,
		_w2219_
	);
	LUT4 #(
		.INIT('h8000)
	) name1260 (
		_w985_,
		_w987_,
		_w1082_,
		_w2219_,
		_w2220_
	);
	LUT2 #(
		.INIT('h8)
	) name1261 (
		_w1059_,
		_w2220_,
		_w2221_
	);
	LUT4 #(
		.INIT('h153f)
	) name1262 (
		_w1059_,
		_w1184_,
		_w1585_,
		_w2220_,
		_w2222_
	);
	LUT4 #(
		.INIT('h3f37)
	) name1263 (
		\u5_state_reg[60]/NET0131 ,
		_w1581_,
		_w1666_,
		_w2021_,
		_w2223_
	);
	LUT3 #(
		.INIT('h8c)
	) name1264 (
		\u5_cmd_asserted2_reg/NET0131 ,
		\u5_state_reg[60]/NET0131 ,
		\u7_mc_br_r_reg/P0001 ,
		_w2224_
	);
	LUT4 #(
		.INIT('h4f00)
	) name1265 (
		_w1533_,
		_w1579_,
		_w1580_,
		_w2224_,
		_w2225_
	);
	LUT2 #(
		.INIT('h1)
	) name1266 (
		_w2221_,
		_w2225_,
		_w2226_
	);
	LUT3 #(
		.INIT('h15)
	) name1267 (
		_w2222_,
		_w2223_,
		_w2226_,
		_w2227_
	);
	LUT3 #(
		.INIT('h02)
	) name1268 (
		\u5_state_reg[63]/NET0131 ,
		\u5_tmr2_done_reg/NET0131 ,
		\u7_mc_ack_r_reg/NET0131 ,
		_w2228_
	);
	LUT3 #(
		.INIT('h80)
	) name1269 (
		_w1059_,
		_w1172_,
		_w2228_,
		_w2229_
	);
	LUT2 #(
		.INIT('h1)
	) name1270 (
		_w1586_,
		_w2229_,
		_w2230_
	);
	LUT4 #(
		.INIT('hb000)
	) name1271 (
		_w1533_,
		_w1579_,
		_w1580_,
		_w1650_,
		_w2231_
	);
	LUT4 #(
		.INIT('h8a00)
	) name1272 (
		\u5_state_reg[63]/NET0131 ,
		_w1533_,
		_w1579_,
		_w1580_,
		_w2232_
	);
	LUT3 #(
		.INIT('h23)
	) name1273 (
		_w2021_,
		_w2231_,
		_w2232_,
		_w2233_
	);
	LUT3 #(
		.INIT('h8c)
	) name1274 (
		\u5_cmd_asserted2_reg/NET0131 ,
		\u5_state_reg[63]/NET0131 ,
		\u7_mc_br_r_reg/P0001 ,
		_w2234_
	);
	LUT4 #(
		.INIT('h4f00)
	) name1275 (
		_w1533_,
		_w1579_,
		_w1580_,
		_w2234_,
		_w2235_
	);
	LUT2 #(
		.INIT('h1)
	) name1276 (
		_w2229_,
		_w2235_,
		_w2236_
	);
	LUT3 #(
		.INIT('h15)
	) name1277 (
		_w2230_,
		_w2233_,
		_w2236_,
		_w2237_
	);
	LUT2 #(
		.INIT('h1)
	) name1278 (
		\u5_cmd_asserted_reg/NET0131 ,
		\u5_state_reg[7]/NET0131 ,
		_w2238_
	);
	LUT3 #(
		.INIT('h08)
	) name1279 (
		_w1100_,
		_w1161_,
		_w2238_,
		_w2239_
	);
	LUT2 #(
		.INIT('h2)
	) name1280 (
		\u5_tmr_done_reg/NET0131 ,
		\u5_wb_wait_r_reg/P0001 ,
		_w2240_
	);
	LUT3 #(
		.INIT('he2)
	) name1281 (
		\u5_state_reg[7]/NET0131 ,
		\u5_tmr_done_reg/NET0131 ,
		\u5_wb_wait_r_reg/P0001 ,
		_w2241_
	);
	LUT2 #(
		.INIT('h4)
	) name1282 (
		_w1270_,
		_w2241_,
		_w2242_
	);
	LUT3 #(
		.INIT('h80)
	) name1283 (
		_w1100_,
		_w1110_,
		_w2242_,
		_w2243_
	);
	LUT2 #(
		.INIT('he)
	) name1284 (
		_w2239_,
		_w2243_,
		_w2244_
	);
	LUT3 #(
		.INIT('h80)
	) name1285 (
		\u5_wb_wait_r_reg/P0001 ,
		_w976_,
		_w1118_,
		_w2245_
	);
	LUT2 #(
		.INIT('h8)
	) name1286 (
		\u0_sp_csc_reg[10]/NET0131 ,
		\u5_wb_wait_r_reg/P0001 ,
		_w2246_
	);
	LUT3 #(
		.INIT('h70)
	) name1287 (
		_w976_,
		_w1114_,
		_w2246_,
		_w2247_
	);
	LUT2 #(
		.INIT('h1)
	) name1288 (
		_w2245_,
		_w2247_,
		_w2248_
	);
	LUT2 #(
		.INIT('h4)
	) name1289 (
		_w1568_,
		_w2248_,
		_w2249_
	);
	LUT3 #(
		.INIT('h08)
	) name1290 (
		_w1100_,
		_w1108_,
		_w1135_,
		_w2250_
	);
	LUT3 #(
		.INIT('h45)
	) name1291 (
		_w1586_,
		_w2249_,
		_w2250_,
		_w2251_
	);
	LUT3 #(
		.INIT('h80)
	) name1292 (
		\u2_bank_open_reg/P0001 ,
		_w976_,
		_w1118_,
		_w2252_
	);
	LUT2 #(
		.INIT('h8)
	) name1293 (
		\u0_sp_csc_reg[10]/NET0131 ,
		\u2_bank_open_reg/P0001 ,
		_w2253_
	);
	LUT3 #(
		.INIT('h70)
	) name1294 (
		_w976_,
		_w1114_,
		_w2253_,
		_w2254_
	);
	LUT3 #(
		.INIT('ha8)
	) name1295 (
		\u2_row_same_reg/P0001 ,
		_w2252_,
		_w2254_,
		_w2255_
	);
	LUT3 #(
		.INIT('h80)
	) name1296 (
		_w1339_,
		_w2019_,
		_w2255_,
		_w2256_
	);
	LUT4 #(
		.INIT('h33f7)
	) name1297 (
		\u5_state_reg[8]/NET0131 ,
		_w1581_,
		_w2021_,
		_w2256_,
		_w2257_
	);
	LUT3 #(
		.INIT('h8c)
	) name1298 (
		\u5_cmd_asserted2_reg/NET0131 ,
		\u5_state_reg[8]/NET0131 ,
		\u7_mc_br_r_reg/P0001 ,
		_w2258_
	);
	LUT4 #(
		.INIT('h4f00)
	) name1299 (
		_w1533_,
		_w1579_,
		_w1580_,
		_w2258_,
		_w2259_
	);
	LUT3 #(
		.INIT('h0b)
	) name1300 (
		_w2249_,
		_w2250_,
		_w2259_,
		_w2260_
	);
	LUT3 #(
		.INIT('h15)
	) name1301 (
		_w2251_,
		_w2257_,
		_w2260_,
		_w2261_
	);
	LUT4 #(
		.INIT('h0080)
	) name1302 (
		\u5_state_reg[9]/NET0131 ,
		_w1100_,
		_w1108_,
		_w1135_,
		_w2262_
	);
	LUT2 #(
		.INIT('h4)
	) name1303 (
		\u5_cmd_asserted_reg/NET0131 ,
		\u5_state_reg[9]/NET0131 ,
		_w2263_
	);
	LUT4 #(
		.INIT('ha800)
	) name1304 (
		_w1100_,
		_w1102_,
		_w1104_,
		_w2263_,
		_w2264_
	);
	LUT2 #(
		.INIT('h1)
	) name1305 (
		_w2262_,
		_w2264_,
		_w2265_
	);
	LUT3 #(
		.INIT('h80)
	) name1306 (
		_w1100_,
		_w1110_,
		_w2240_,
		_w2266_
	);
	LUT4 #(
		.INIT('h0800)
	) name1307 (
		_w1100_,
		_w1108_,
		_w1568_,
		_w2248_,
		_w2267_
	);
	LUT3 #(
		.INIT('h54)
	) name1308 (
		_w1564_,
		_w2266_,
		_w2267_,
		_w2268_
	);
	LUT2 #(
		.INIT('hd)
	) name1309 (
		_w2265_,
		_w2268_,
		_w2269_
	);
	LUT2 #(
		.INIT('h8)
	) name1310 (
		_w965_,
		_w1219_,
		_w2270_
	);
	LUT3 #(
		.INIT('h02)
	) name1311 (
		\u5_state_reg[42]/NET0131 ,
		\u5_state_reg[43]/NET0131 ,
		\u5_tmr2_done_reg/NET0131 ,
		_w2271_
	);
	LUT3 #(
		.INIT('h80)
	) name1312 (
		_w963_,
		_w1238_,
		_w2271_,
		_w2272_
	);
	LUT3 #(
		.INIT('ha8)
	) name1313 (
		_w1063_,
		_w2270_,
		_w2272_,
		_w2273_
	);
	LUT3 #(
		.INIT('h80)
	) name1314 (
		\u7_mc_ack_r_reg/NET0131 ,
		_w1059_,
		_w1172_,
		_w2274_
	);
	LUT2 #(
		.INIT('he)
	) name1315 (
		_w1593_,
		_w2274_,
		_w2275_
	);
	LUT3 #(
		.INIT('h0e)
	) name1316 (
		\u5_state_reg[65]/NET0131 ,
		\u5_tmr2_done_reg/NET0131 ,
		\u7_mc_ack_r_reg/NET0131 ,
		_w2276_
	);
	LUT4 #(
		.INIT('ha800)
	) name1317 (
		_w1059_,
		_w1083_,
		_w1172_,
		_w2276_,
		_w2277_
	);
	LUT3 #(
		.INIT('h40)
	) name1318 (
		\u5_cmd_asserted_reg/NET0131 ,
		_w1100_,
		_w1161_,
		_w2278_
	);
	LUT3 #(
		.INIT('ha3)
	) name1319 (
		\u5_rfr_ack_r_reg/NET0131 ,
		\u5_state_reg[6]/NET0131 ,
		\u5_tmr_done_reg/NET0131 ,
		_w2279_
	);
	LUT3 #(
		.INIT('h08)
	) name1320 (
		_w982_,
		_w1181_,
		_w2279_,
		_w2280_
	);
	LUT2 #(
		.INIT('h8)
	) name1321 (
		_w1002_,
		_w2280_,
		_w2281_
	);
	LUT3 #(
		.INIT('h01)
	) name1322 (
		_w1586_,
		_w2278_,
		_w2281_,
		_w2282_
	);
	LUT3 #(
		.INIT('h02)
	) name1323 (
		_w1338_,
		_w2252_,
		_w2254_,
		_w2283_
	);
	LUT3 #(
		.INIT('h80)
	) name1324 (
		_w1336_,
		_w2019_,
		_w2283_,
		_w2284_
	);
	LUT4 #(
		.INIT('h33f7)
	) name1325 (
		\u5_state_reg[6]/NET0131 ,
		_w1581_,
		_w2021_,
		_w2284_,
		_w2285_
	);
	LUT3 #(
		.INIT('h8c)
	) name1326 (
		\u5_cmd_asserted2_reg/NET0131 ,
		\u5_state_reg[6]/NET0131 ,
		\u7_mc_br_r_reg/P0001 ,
		_w2286_
	);
	LUT4 #(
		.INIT('h4f00)
	) name1327 (
		_w1533_,
		_w1579_,
		_w1580_,
		_w2286_,
		_w2287_
	);
	LUT3 #(
		.INIT('h01)
	) name1328 (
		_w2278_,
		_w2281_,
		_w2287_,
		_w2288_
	);
	LUT3 #(
		.INIT('h15)
	) name1329 (
		_w2282_,
		_w2285_,
		_w2288_,
		_w2289_
	);
	LUT2 #(
		.INIT('h2)
	) name1330 (
		\u5_wb_cycle_reg/NET0131 ,
		_w1564_,
		_w2290_
	);
	LUT4 #(
		.INIT('h8000)
	) name1331 (
		_w1002_,
		_w1005_,
		_w1006_,
		_w2290_,
		_w2291_
	);
	LUT4 #(
		.INIT('h0b00)
	) name1332 (
		_w1539_,
		_w1599_,
		_w1608_,
		_w2291_,
		_w2292_
	);
	LUT3 #(
		.INIT('h20)
	) name1333 (
		\u5_state_reg[10]/NET0131 ,
		\u5_state_reg[11]/NET0131 ,
		\u5_tmr_done_reg/NET0131 ,
		_w2293_
	);
	LUT3 #(
		.INIT('h80)
	) name1334 (
		_w1002_,
		_w1005_,
		_w2293_,
		_w2294_
	);
	LUT2 #(
		.INIT('he)
	) name1335 (
		_w2292_,
		_w2294_,
		_w2295_
	);
	LUT2 #(
		.INIT('h2)
	) name1336 (
		\u5_state_reg[1]/NET0131 ,
		\u5_state_reg[52]/NET0131 ,
		_w2296_
	);
	LUT3 #(
		.INIT('h80)
	) name1337 (
		_w1125_,
		_w1540_,
		_w1541_,
		_w2297_
	);
	LUT4 #(
		.INIT('h1000)
	) name1338 (
		_w1539_,
		_w2105_,
		_w2296_,
		_w2297_,
		_w2298_
	);
	LUT4 #(
		.INIT('hff60)
	) name1339 (
		\u5_burst_cnt_reg[1]/NET0131 ,
		_w2004_,
		_w2008_,
		_w2298_,
		_w2299_
	);
	LUT4 #(
		.INIT('h0400)
	) name1340 (
		_w1539_,
		_w2040_,
		_w2105_,
		_w2296_,
		_w2300_
	);
	LUT4 #(
		.INIT('hff48)
	) name1341 (
		\u5_burst_cnt_reg[3]/NET0131 ,
		_w2008_,
		_w2035_,
		_w2300_,
		_w2301_
	);
	LUT3 #(
		.INIT('h80)
	) name1342 (
		\u5_resume_req_r_reg/NET0131 ,
		_w1035_,
		_w1050_,
		_w2302_
	);
	LUT3 #(
		.INIT('h08)
	) name1343 (
		\u5_cmd_asserted_reg/NET0131 ,
		\u5_state_reg[52]/NET0131 ,
		\u5_state_reg[53]/NET0131 ,
		_w2303_
	);
	LUT3 #(
		.INIT('h80)
	) name1344 (
		_w992_,
		_w999_,
		_w2303_,
		_w2304_
	);
	LUT3 #(
		.INIT('h04)
	) name1345 (
		\u5_state_reg[52]/NET0131 ,
		\u5_state_reg[53]/NET0131 ,
		\u5_tmr2_done_reg/NET0131 ,
		_w2305_
	);
	LUT3 #(
		.INIT('h80)
	) name1346 (
		_w992_,
		_w999_,
		_w2305_,
		_w2306_
	);
	LUT3 #(
		.INIT('ha8)
	) name1347 (
		_w991_,
		_w2304_,
		_w2306_,
		_w2307_
	);
	LUT4 #(
		.INIT('h0001)
	) name1348 (
		\u5_burst_cnt_reg[0]/NET0131 ,
		\u5_burst_cnt_reg[1]/NET0131 ,
		\u5_burst_cnt_reg[2]/NET0131 ,
		\u5_burst_cnt_reg[3]/NET0131 ,
		_w2308_
	);
	LUT4 #(
		.INIT('hfe00)
	) name1349 (
		\u5_wr_cycle_reg/NET0131 ,
		_w998_,
		_w1010_,
		_w2308_,
		_w2309_
	);
	LUT4 #(
		.INIT('hef00)
	) name1350 (
		_w1724_,
		_w1728_,
		_w1980_,
		_w2309_,
		_w2310_
	);
	LUT4 #(
		.INIT('h90c0)
	) name1351 (
		\u5_burst_cnt_reg[4]/NET0131 ,
		\u5_burst_cnt_reg[5]/NET0131 ,
		_w2008_,
		_w2310_,
		_w2311_
	);
	LUT4 #(
		.INIT('hfe00)
	) name1352 (
		\u5_wr_cycle_reg/NET0131 ,
		_w998_,
		_w1010_,
		_w1605_,
		_w2312_
	);
	LUT4 #(
		.INIT('hef00)
	) name1353 (
		_w1724_,
		_w1728_,
		_w1980_,
		_w2312_,
		_w2313_
	);
	LUT2 #(
		.INIT('h8)
	) name1354 (
		_w2008_,
		_w2313_,
		_w2314_
	);
	LUT2 #(
		.INIT('h1)
	) name1355 (
		\u5_burst_cnt_reg[4]/NET0131 ,
		\u5_burst_cnt_reg[5]/NET0131 ,
		_w2315_
	);
	LUT3 #(
		.INIT('h02)
	) name1356 (
		\u5_burst_cnt_reg[6]/NET0131 ,
		\u5_state_reg[1]/NET0131 ,
		\u5_state_reg[52]/NET0131 ,
		_w2316_
	);
	LUT3 #(
		.INIT('h70)
	) name1357 (
		_w2310_,
		_w2315_,
		_w2316_,
		_w2317_
	);
	LUT2 #(
		.INIT('he)
	) name1358 (
		_w2314_,
		_w2317_,
		_w2318_
	);
	LUT2 #(
		.INIT('he)
	) name1359 (
		\u5_oe__reg/NET0131 ,
		\u5_susp_sel_r_reg/NET0131 ,
		_w2319_
	);
	LUT3 #(
		.INIT('h48)
	) name1360 (
		\u5_burst_cnt_reg[7]/NET0131 ,
		_w2008_,
		_w2313_,
		_w2320_
	);
	LUT3 #(
		.INIT('h48)
	) name1361 (
		\u5_burst_cnt_reg[4]/NET0131 ,
		_w2008_,
		_w2310_,
		_w2321_
	);
	LUT4 #(
		.INIT('h135f)
	) name1362 (
		_w991_,
		_w1041_,
		_w1055_,
		_w1091_,
		_w2322_
	);
	LUT2 #(
		.INIT('h2)
	) name1363 (
		\u5_state_reg[48]/NET0131 ,
		\u5_tmr2_done_reg/NET0131 ,
		_w2323_
	);
	LUT3 #(
		.INIT('hba)
	) name1364 (
		_w1218_,
		_w2322_,
		_w2323_,
		_w2324_
	);
	LUT2 #(
		.INIT('h8)
	) name1365 (
		\u5_wb_cycle_reg/NET0131 ,
		_w1564_,
		_w2325_
	);
	LUT3 #(
		.INIT('h0d)
	) name1366 (
		\u5_wb_cycle_reg/NET0131 ,
		_w1564_,
		_w1608_,
		_w2326_
	);
	LUT4 #(
		.INIT('h040f)
	) name1367 (
		_w1539_,
		_w1599_,
		_w2325_,
		_w2326_,
		_w2327_
	);
	LUT4 #(
		.INIT('h2aaa)
	) name1368 (
		\u5_state_reg[15]/NET0131 ,
		_w1603_,
		_w1604_,
		_w1607_,
		_w2328_
	);
	LUT3 #(
		.INIT('hb0)
	) name1369 (
		_w1539_,
		_w1599_,
		_w2328_,
		_w2329_
	);
	LUT3 #(
		.INIT('ha2)
	) name1370 (
		_w1045_,
		_w2327_,
		_w2329_,
		_w2330_
	);
	LUT3 #(
		.INIT('h40)
	) name1371 (
		\u5_cmd_asserted_reg/NET0131 ,
		_w1100_,
		_w1158_,
		_w2331_
	);
	LUT2 #(
		.INIT('h4)
	) name1372 (
		_w1564_,
		_w1720_,
		_w2332_
	);
	LUT3 #(
		.INIT('h80)
	) name1373 (
		_w1002_,
		_w1143_,
		_w2332_,
		_w2333_
	);
	LUT2 #(
		.INIT('h8)
	) name1374 (
		_w1937_,
		_w2333_,
		_w2334_
	);
	LUT4 #(
		.INIT('h040f)
	) name1375 (
		_w1539_,
		_w1599_,
		_w2331_,
		_w2334_,
		_w2335_
	);
	LUT2 #(
		.INIT('h4)
	) name1376 (
		_w1617_,
		_w2335_,
		_w2336_
	);
	LUT2 #(
		.INIT('hb)
	) name1377 (
		_w2330_,
		_w2336_,
		_w2337_
	);
	LUT3 #(
		.INIT('h80)
	) name1378 (
		_w991_,
		_w1250_,
		_w1736_,
		_w2338_
	);
	LUT2 #(
		.INIT('h2)
	) name1379 (
		_w1566_,
		_w1608_,
		_w2339_
	);
	LUT4 #(
		.INIT('h20aa)
	) name1380 (
		_w996_,
		_w1539_,
		_w1599_,
		_w2339_,
		_w2340_
	);
	LUT2 #(
		.INIT('he)
	) name1381 (
		_w2338_,
		_w2340_,
		_w2341_
	);
	LUT3 #(
		.INIT('h08)
	) name1382 (
		_w1100_,
		_w1140_,
		_w1929_,
		_w2342_
	);
	LUT3 #(
		.INIT('h40)
	) name1383 (
		_w1608_,
		_w1927_,
		_w2342_,
		_w2343_
	);
	LUT3 #(
		.INIT('hb0)
	) name1384 (
		_w1539_,
		_w1599_,
		_w2343_,
		_w2344_
	);
	LUT2 #(
		.INIT('h8)
	) name1385 (
		_w1935_,
		_w2344_,
		_w2345_
	);
	LUT4 #(
		.INIT('h3331)
	) name1386 (
		_w1141_,
		_w1145_,
		_w1613_,
		_w1614_,
		_w2346_
	);
	LUT3 #(
		.INIT('h20)
	) name1387 (
		\u5_cmd_asserted_reg/NET0131 ,
		\u6_rmw_r_reg/NET0131 ,
		wb_cyc_i_pad,
		_w2347_
	);
	LUT4 #(
		.INIT('h7000)
	) name1388 (
		_w1014_,
		_w1015_,
		_w1131_,
		_w2347_,
		_w2348_
	);
	LUT2 #(
		.INIT('h4)
	) name1389 (
		\u5_wb_cycle_reg/NET0131 ,
		_w2348_,
		_w2349_
	);
	LUT2 #(
		.INIT('h4)
	) name1390 (
		_w1608_,
		_w2348_,
		_w2350_
	);
	LUT4 #(
		.INIT('h040f)
	) name1391 (
		_w1539_,
		_w1599_,
		_w2349_,
		_w2350_,
		_w2351_
	);
	LUT2 #(
		.INIT('h4)
	) name1392 (
		\u5_cmd_asserted_reg/NET0131 ,
		\u5_state_reg[14]/NET0131 ,
		_w2352_
	);
	LUT4 #(
		.INIT('h00fd)
	) name1393 (
		_w1141_,
		_w1613_,
		_w1614_,
		_w2352_,
		_w2353_
	);
	LUT3 #(
		.INIT('h15)
	) name1394 (
		_w2346_,
		_w2351_,
		_w2353_,
		_w2354_
	);
	LUT2 #(
		.INIT('he)
	) name1395 (
		_w2345_,
		_w2354_,
		_w2355_
	);
	LUT3 #(
		.INIT('h08)
	) name1396 (
		\u5_data_oe_reg/NET0131 ,
		\u5_mc_c_oe_reg/NET0131 ,
		\u5_susp_sel_r_reg/NET0131 ,
		_w2356_
	);
	LUT2 #(
		.INIT('h1)
	) name1397 (
		\u5_state_reg[24]/NET0131 ,
		\u5_tmr_done_reg/NET0131 ,
		_w2357_
	);
	LUT3 #(
		.INIT('h80)
	) name1398 (
		_w975_,
		_w984_,
		_w1046_,
		_w2358_
	);
	LUT4 #(
		.INIT('h1c3c)
	) name1399 (
		\u5_ir_cnt_done_reg/P0001 ,
		\u5_state_reg[23]/NET0131 ,
		\u5_state_reg[25]/NET0131 ,
		\u5_tmr_done_reg/NET0131 ,
		_w2359_
	);
	LUT4 #(
		.INIT('h2000)
	) name1400 (
		_w1035_,
		_w2357_,
		_w2358_,
		_w2359_,
		_w2360_
	);
	LUT2 #(
		.INIT('h4)
	) name1401 (
		\u5_cmd_asserted_reg/NET0131 ,
		_w1263_,
		_w2361_
	);
	LUT3 #(
		.INIT('h80)
	) name1402 (
		_w984_,
		_w1046_,
		_w2361_,
		_w2362_
	);
	LUT2 #(
		.INIT('h8)
	) name1403 (
		_w1035_,
		_w2362_,
		_w2363_
	);
	LUT2 #(
		.INIT('he)
	) name1404 (
		_w2360_,
		_w2363_,
		_w2364_
	);
	LUT2 #(
		.INIT('h1)
	) name1405 (
		\u5_wb_stb_first_reg/NET0131 ,
		wb_stb_i_pad,
		_w2365_
	);
	LUT4 #(
		.INIT('h1000)
	) name1406 (
		\u6_read_go_r_reg/NET0131 ,
		\u6_write_go_r_reg/NET0131 ,
		wb_cyc_i_pad,
		wb_stb_i_pad,
		_w2366_
	);
	LUT3 #(
		.INIT('h02)
	) name1407 (
		\u6_wb_first_r_reg/NET0131 ,
		wb_ack_o_pad,
		wb_err_o_pad,
		_w2367_
	);
	LUT4 #(
		.INIT('h5551)
	) name1408 (
		\u5_wb_stb_first_reg/NET0131 ,
		\u6_wb_first_r_reg/NET0131 ,
		wb_ack_o_pad,
		wb_err_o_pad,
		_w2368_
	);
	LUT4 #(
		.INIT('h2033)
	) name1409 (
		_w1748_,
		_w2365_,
		_w2366_,
		_w2368_,
		_w2369_
	);
	LUT3 #(
		.INIT('h10)
	) name1410 (
		_w1564_,
		_w1566_,
		_w2369_,
		_w2370_
	);
	LUT4 #(
		.INIT('h4f00)
	) name1411 (
		_w1539_,
		_w1599_,
		_w1723_,
		_w2369_,
		_w2371_
	);
	LUT4 #(
		.INIT('hf4f0)
	) name1412 (
		_w1728_,
		_w1747_,
		_w2370_,
		_w2371_,
		_w2372_
	);
	LUT2 #(
		.INIT('h1)
	) name1413 (
		\u5_cmd_asserted_reg/NET0131 ,
		\u5_state_reg[19]/NET0131 ,
		_w2373_
	);
	LUT3 #(
		.INIT('h08)
	) name1414 (
		_w1035_,
		_w1283_,
		_w2373_,
		_w2374_
	);
	LUT3 #(
		.INIT('h02)
	) name1415 (
		\u5_state_reg[19]/NET0131 ,
		\u5_state_reg[20]/NET0131 ,
		\u5_tmr_done_reg/NET0131 ,
		_w2375_
	);
	LUT3 #(
		.INIT('h80)
	) name1416 (
		_w1035_,
		_w1148_,
		_w2375_,
		_w2376_
	);
	LUT2 #(
		.INIT('he)
	) name1417 (
		_w2374_,
		_w2376_,
		_w2377_
	);
	LUT3 #(
		.INIT('h80)
	) name1418 (
		_w991_,
		_w995_,
		_w2339_,
		_w2378_
	);
	LUT4 #(
		.INIT('h4440)
	) name1419 (
		\u5_state_reg[52]/NET0131 ,
		\u5_state_reg[53]/NET0131 ,
		\u5_state_reg[54]/NET0131 ,
		\u5_tmr2_done_reg/NET0131 ,
		_w2379_
	);
	LUT3 #(
		.INIT('h80)
	) name1420 (
		_w992_,
		_w999_,
		_w2379_,
		_w2380_
	);
	LUT2 #(
		.INIT('h8)
	) name1421 (
		_w991_,
		_w2380_,
		_w2381_
	);
	LUT4 #(
		.INIT('hffb0)
	) name1422 (
		_w1539_,
		_w1599_,
		_w2378_,
		_w2381_,
		_w2382_
	);
	LUT3 #(
		.INIT('h80)
	) name1423 (
		_w1184_,
		_w1185_,
		_w1569_,
		_w2383_
	);
	LUT4 #(
		.INIT('h8000)
	) name1424 (
		_w1184_,
		_w1185_,
		_w1546_,
		_w1569_,
		_w2384_
	);
	LUT3 #(
		.INIT('h80)
	) name1425 (
		_w1540_,
		_w1541_,
		_w2384_,
		_w2385_
	);
	LUT2 #(
		.INIT('h4)
	) name1426 (
		_w1539_,
		_w2385_,
		_w2386_
	);
	LUT2 #(
		.INIT('h8)
	) name1427 (
		_w968_,
		_w969_,
		_w2387_
	);
	LUT3 #(
		.INIT('h1c)
	) name1428 (
		\u5_cmd_asserted_reg/NET0131 ,
		\u5_state_reg[47]/NET0131 ,
		\u5_state_reg[48]/NET0131 ,
		_w2388_
	);
	LUT3 #(
		.INIT('h80)
	) name1429 (
		_w1041_,
		_w2387_,
		_w2388_,
		_w2389_
	);
	LUT4 #(
		.INIT('h8000)
	) name1430 (
		_w1041_,
		_w1655_,
		_w2387_,
		_w2388_,
		_w2390_
	);
	LUT3 #(
		.INIT('h80)
	) name1431 (
		_w1540_,
		_w1541_,
		_w2390_,
		_w2391_
	);
	LUT2 #(
		.INIT('h4)
	) name1432 (
		_w1539_,
		_w2391_,
		_w2392_
	);
	LUT4 #(
		.INIT('h0075)
	) name1433 (
		\u5_state_reg[51]/NET0131 ,
		_w1539_,
		_w1694_,
		_w2389_,
		_w2393_
	);
	LUT2 #(
		.INIT('h1)
	) name1434 (
		_w2392_,
		_w2393_,
		_w2394_
	);
	LUT2 #(
		.INIT('h2)
	) name1435 (
		\u5_state_reg[40]/NET0131 ,
		\u5_state_reg[51]/NET0131 ,
		_w2395_
	);
	LUT3 #(
		.INIT('hb0)
	) name1436 (
		_w1539_,
		_w2169_,
		_w2395_,
		_w2396_
	);
	LUT2 #(
		.INIT('h1)
	) name1437 (
		\u5_state_reg[40]/NET0131 ,
		\u5_state_reg[51]/NET0131 ,
		_w2397_
	);
	LUT4 #(
		.INIT('h0001)
	) name1438 (
		\u5_timer2_reg[0]/P0001 ,
		\u5_timer2_reg[1]/P0001 ,
		\u5_timer2_reg[2]/P0001 ,
		\u5_timer2_reg[3]/P0001 ,
		_w2398_
	);
	LUT3 #(
		.INIT('h01)
	) name1439 (
		\u5_timer2_reg[4]/P0001 ,
		\u5_timer2_reg[5]/P0001 ,
		\u5_timer2_reg[6]/P0001 ,
		_w2399_
	);
	LUT2 #(
		.INIT('h1)
	) name1440 (
		\u5_timer2_reg[7]/P0001 ,
		\u5_timer2_reg[8]/P0001 ,
		_w2400_
	);
	LUT3 #(
		.INIT('h80)
	) name1441 (
		_w2398_,
		_w2399_,
		_w2400_,
		_w2401_
	);
	LUT4 #(
		.INIT('h0001)
	) name1442 (
		\u5_state_reg[36]/NET0131 ,
		\u5_state_reg[41]/NET0131 ,
		\u5_state_reg[43]/NET0131 ,
		\u5_state_reg[45]/NET0131 ,
		_w2402_
	);
	LUT3 #(
		.INIT('h01)
	) name1443 (
		\u5_timer2_reg[0]/P0001 ,
		\u5_timer2_reg[1]/P0001 ,
		\u5_timer2_reg[2]/P0001 ,
		_w2403_
	);
	LUT3 #(
		.INIT('h1e)
	) name1444 (
		\u5_timer2_reg[0]/P0001 ,
		\u5_timer2_reg[1]/P0001 ,
		\u5_timer2_reg[2]/P0001 ,
		_w2404_
	);
	LUT2 #(
		.INIT('h2)
	) name1445 (
		_w2402_,
		_w2404_,
		_w2405_
	);
	LUT3 #(
		.INIT('h20)
	) name1446 (
		_w2397_,
		_w2401_,
		_w2405_,
		_w2406_
	);
	LUT2 #(
		.INIT('h2)
	) name1447 (
		_w2397_,
		_w2402_,
		_w2407_
	);
	LUT4 #(
		.INIT('h040f)
	) name1448 (
		_w1539_,
		_w2145_,
		_w2406_,
		_w2407_,
		_w2408_
	);
	LUT3 #(
		.INIT('h80)
	) name1449 (
		\u5_tmr2_done_reg/NET0131 ,
		_w1041_,
		_w1091_,
		_w2409_
	);
	LUT3 #(
		.INIT('h0b)
	) name1450 (
		_w1539_,
		_w2391_,
		_w2409_,
		_w2410_
	);
	LUT3 #(
		.INIT('hb0)
	) name1451 (
		_w2396_,
		_w2408_,
		_w2410_,
		_w2411_
	);
	LUT2 #(
		.INIT('h4)
	) name1452 (
		_w2389_,
		_w2409_,
		_w2412_
	);
	LUT3 #(
		.INIT('h80)
	) name1453 (
		_w1184_,
		_w1185_,
		_w1343_,
		_w2413_
	);
	LUT2 #(
		.INIT('h1)
	) name1454 (
		_w1214_,
		_w2413_,
		_w2414_
	);
	LUT4 #(
		.INIT('h4f00)
	) name1455 (
		_w1539_,
		_w2124_,
		_w2412_,
		_w2414_,
		_w2415_
	);
	LUT4 #(
		.INIT('h5455)
	) name1456 (
		_w2386_,
		_w2394_,
		_w2411_,
		_w2415_,
		_w2416_
	);
	LUT3 #(
		.INIT('h2a)
	) name1457 (
		\u5_state_reg[37]/NET0131 ,
		_w976_,
		_w1975_,
		_w2417_
	);
	LUT3 #(
		.INIT('h80)
	) name1458 (
		\u1_acs_addr_reg[12]/P0001 ,
		\u1_u0_out_r_reg[12]/P0001 ,
		\u5_tmr2_done_reg/NET0131 ,
		_w2418_
	);
	LUT4 #(
		.INIT('h7500)
	) name1459 (
		_w964_,
		_w1974_,
		_w2417_,
		_w2418_,
		_w2419_
	);
	LUT3 #(
		.INIT('h80)
	) name1460 (
		\u1_acs_addr_reg[13]/P0001 ,
		\u1_acs_addr_reg[14]/P0001 ,
		\u1_acs_addr_reg[15]/P0001 ,
		_w2420_
	);
	LUT3 #(
		.INIT('h80)
	) name1461 (
		\u1_acs_addr_reg[16]/P0001 ,
		\u1_acs_addr_reg[17]/P0001 ,
		\u1_acs_addr_reg[18]/P0001 ,
		_w2421_
	);
	LUT3 #(
		.INIT('h80)
	) name1462 (
		\u1_acs_addr_reg[19]/P0001 ,
		\u1_acs_addr_reg[20]/P0001 ,
		\u1_acs_addr_reg[21]/P0001 ,
		_w2422_
	);
	LUT4 #(
		.INIT('h8000)
	) name1463 (
		_w2419_,
		_w2420_,
		_w2421_,
		_w2422_,
		_w2423_
	);
	LUT2 #(
		.INIT('h1)
	) name1464 (
		\u5_cs_le_reg/P0001 ,
		wb_we_i_pad,
		_w2424_
	);
	LUT4 #(
		.INIT('h9300)
	) name1465 (
		\u1_acs_addr_reg[22]/P0001 ,
		\u1_acs_addr_reg[23]/P0001 ,
		_w2423_,
		_w2424_,
		_w2425_
	);
	LUT3 #(
		.INIT('h2a)
	) name1466 (
		\wb_addr_i[25]_pad ,
		_w976_,
		_w1971_,
		_w2426_
	);
	LUT4 #(
		.INIT('h0e0f)
	) name1467 (
		_w1970_,
		_w1976_,
		_w2424_,
		_w2426_,
		_w2427_
	);
	LUT3 #(
		.INIT('h2a)
	) name1468 (
		\wb_addr_i[24]_pad ,
		_w976_,
		_w1975_,
		_w2428_
	);
	LUT3 #(
		.INIT('h10)
	) name1469 (
		_w1972_,
		_w1974_,
		_w2428_,
		_w2429_
	);
	LUT3 #(
		.INIT('h2a)
	) name1470 (
		\wb_addr_i[23]_pad ,
		_w976_,
		_w1971_,
		_w2430_
	);
	LUT3 #(
		.INIT('h40)
	) name1471 (
		_w1970_,
		_w1976_,
		_w2430_,
		_w2431_
	);
	LUT3 #(
		.INIT('h02)
	) name1472 (
		_w2427_,
		_w2429_,
		_w2431_,
		_w2432_
	);
	LUT2 #(
		.INIT('h1)
	) name1473 (
		_w2425_,
		_w2432_,
		_w2433_
	);
	LUT3 #(
		.INIT('hb0)
	) name1474 (
		_w1539_,
		_w2124_,
		_w2383_,
		_w2434_
	);
	LUT4 #(
		.INIT('h004f)
	) name1475 (
		_w1539_,
		_w2124_,
		_w2383_,
		_w2414_,
		_w2435_
	);
	LUT4 #(
		.INIT('h8000)
	) name1476 (
		_w1041_,
		_w2142_,
		_w2387_,
		_w2388_,
		_w2436_
	);
	LUT3 #(
		.INIT('h80)
	) name1477 (
		_w1540_,
		_w1541_,
		_w2436_,
		_w2437_
	);
	LUT2 #(
		.INIT('h4)
	) name1478 (
		_w1539_,
		_w2437_,
		_w2438_
	);
	LUT4 #(
		.INIT('h0075)
	) name1479 (
		\u5_state_reg[51]/NET0131 ,
		_w1539_,
		_w2162_,
		_w2389_,
		_w2439_
	);
	LUT2 #(
		.INIT('h1)
	) name1480 (
		_w2438_,
		_w2439_,
		_w2440_
	);
	LUT2 #(
		.INIT('h6)
	) name1481 (
		\u5_timer2_reg[0]/P0001 ,
		\u5_timer2_reg[1]/P0001 ,
		_w2441_
	);
	LUT2 #(
		.INIT('h2)
	) name1482 (
		_w2402_,
		_w2441_,
		_w2442_
	);
	LUT3 #(
		.INIT('h20)
	) name1483 (
		_w2397_,
		_w2401_,
		_w2442_,
		_w2443_
	);
	LUT4 #(
		.INIT('h004f)
	) name1484 (
		_w1539_,
		_w2105_,
		_w2407_,
		_w2443_,
		_w2444_
	);
	LUT3 #(
		.INIT('hb0)
	) name1485 (
		_w1539_,
		_w2134_,
		_w2395_,
		_w2445_
	);
	LUT3 #(
		.INIT('h23)
	) name1486 (
		_w1539_,
		_w2409_,
		_w2437_,
		_w2446_
	);
	LUT3 #(
		.INIT('hd0)
	) name1487 (
		_w2444_,
		_w2445_,
		_w2446_,
		_w2447_
	);
	LUT3 #(
		.INIT('h08)
	) name1488 (
		_w1540_,
		_w1541_,
		_w1552_,
		_w2448_
	);
	LUT3 #(
		.INIT('h8c)
	) name1489 (
		_w1539_,
		_w2412_,
		_w2448_,
		_w2449_
	);
	LUT2 #(
		.INIT('h1)
	) name1490 (
		_w2434_,
		_w2449_,
		_w2450_
	);
	LUT4 #(
		.INIT('h5455)
	) name1491 (
		_w2435_,
		_w2440_,
		_w2447_,
		_w2450_,
		_w2451_
	);
	LUT3 #(
		.INIT('hb0)
	) name1492 (
		_w1539_,
		_w1697_,
		_w2383_,
		_w2452_
	);
	LUT3 #(
		.INIT('h80)
	) name1493 (
		_w1540_,
		_w1541_,
		_w1664_,
		_w2453_
	);
	LUT3 #(
		.INIT('h8c)
	) name1494 (
		_w1539_,
		_w2395_,
		_w2453_,
		_w2454_
	);
	LUT2 #(
		.INIT('h2)
	) name1495 (
		_w1124_,
		_w2402_,
		_w2455_
	);
	LUT3 #(
		.INIT('h80)
	) name1496 (
		_w1540_,
		_w1541_,
		_w2455_,
		_w2456_
	);
	LUT4 #(
		.INIT('h7f00)
	) name1497 (
		_w2398_,
		_w2399_,
		_w2400_,
		_w2403_,
		_w2457_
	);
	LUT4 #(
		.INIT('hd500)
	) name1498 (
		_w2398_,
		_w2399_,
		_w2400_,
		_w2402_,
		_w2458_
	);
	LUT4 #(
		.INIT('h08cc)
	) name1499 (
		\u5_timer2_reg[3]/P0001 ,
		_w2397_,
		_w2457_,
		_w2458_,
		_w2459_
	);
	LUT3 #(
		.INIT('hb0)
	) name1500 (
		_w1539_,
		_w2456_,
		_w2459_,
		_w2460_
	);
	LUT3 #(
		.INIT('h54)
	) name1501 (
		_w2409_,
		_w2454_,
		_w2460_,
		_w2461_
	);
	LUT3 #(
		.INIT('h8a)
	) name1502 (
		\u5_state_reg[51]/NET0131 ,
		_w1539_,
		_w1898_,
		_w2462_
	);
	LUT4 #(
		.INIT('h040f)
	) name1503 (
		_w1539_,
		_w2160_,
		_w2389_,
		_w2409_,
		_w2463_
	);
	LUT2 #(
		.INIT('h4)
	) name1504 (
		_w2462_,
		_w2463_,
		_w2464_
	);
	LUT4 #(
		.INIT('h8000)
	) name1505 (
		_w1041_,
		_w1707_,
		_w2387_,
		_w2388_,
		_w2465_
	);
	LUT3 #(
		.INIT('h80)
	) name1506 (
		_w1540_,
		_w1541_,
		_w2465_,
		_w2466_
	);
	LUT3 #(
		.INIT('h8c)
	) name1507 (
		_w1539_,
		_w2414_,
		_w2466_,
		_w2467_
	);
	LUT4 #(
		.INIT('hefaa)
	) name1508 (
		_w2452_,
		_w2461_,
		_w2464_,
		_w2467_,
		_w2468_
	);
	LUT3 #(
		.INIT('h80)
	) name1509 (
		_w1184_,
		_w1585_,
		_w2020_,
		_w2469_
	);
	LUT4 #(
		.INIT('h153f)
	) name1510 (
		_w1059_,
		_w1100_,
		_w1108_,
		_w1189_,
		_w2470_
	);
	LUT4 #(
		.INIT('h80aa)
	) name1511 (
		_w1135_,
		_w1581_,
		_w2469_,
		_w2470_,
		_w2471_
	);
	LUT4 #(
		.INIT('h153f)
	) name1512 (
		_w1041_,
		_w1059_,
		_w1211_,
		_w1217_,
		_w2472_
	);
	LUT4 #(
		.INIT('h0100)
	) name1513 (
		_w1087_,
		_w1141_,
		_w1145_,
		_w2472_,
		_w2473_
	);
	LUT3 #(
		.INIT('h20)
	) name1514 (
		_w1314_,
		_w2471_,
		_w2473_,
		_w2474_
	);
	LUT2 #(
		.INIT('hb)
	) name1515 (
		_w1555_,
		_w2474_,
		_w2475_
	);
	LUT4 #(
		.INIT('hb8bb)
	) name1516 (
		\u5_data_oe_r2_reg/NET0131 ,
		\u5_wr_cycle_reg/NET0131 ,
		_w1555_,
		_w2474_,
		_w2476_
	);
	LUT2 #(
		.INIT('h8)
	) name1517 (
		\u5_cnt_reg/NET0131 ,
		\u5_wb_cycle_reg/NET0131 ,
		_w2477_
	);
	LUT4 #(
		.INIT('h7f00)
	) name1518 (
		_w1603_,
		_w1604_,
		_w1607_,
		_w2477_,
		_w2478_
	);
	LUT4 #(
		.INIT('h1055)
	) name1519 (
		mc_cke_pad_o__pad,
		_w1539_,
		_w1599_,
		_w2478_,
		_w2479_
	);
	LUT4 #(
		.INIT('ha800)
	) name1520 (
		_w1132_,
		_w1564_,
		_w1566_,
		_w2478_,
		_w2480_
	);
	LUT4 #(
		.INIT('h20aa)
	) name1521 (
		_w1045_,
		_w1539_,
		_w1599_,
		_w2480_,
		_w2481_
	);
	LUT3 #(
		.INIT('h20)
	) name1522 (
		\u5_cke_r_reg/NET0131 ,
		_w2479_,
		_w2481_,
		_w2482_
	);
	LUT3 #(
		.INIT('h10)
	) name1523 (
		_w1192_,
		_w1305_,
		_w2082_,
		_w2483_
	);
	LUT3 #(
		.INIT('h80)
	) name1524 (
		_w1316_,
		_w1317_,
		_w2483_,
		_w2484_
	);
	LUT4 #(
		.INIT('h135f)
	) name1525 (
		_w1035_,
		_w1068_,
		_w1264_,
		_w1288_,
		_w2485_
	);
	LUT4 #(
		.INIT('h0040)
	) name1526 (
		_w1075_,
		_w1080_,
		_w1088_,
		_w1105_,
		_w2486_
	);
	LUT2 #(
		.INIT('h8)
	) name1527 (
		_w1322_,
		_w2486_,
		_w2487_
	);
	LUT3 #(
		.INIT('h80)
	) name1528 (
		_w1322_,
		_w2485_,
		_w2486_,
		_w2488_
	);
	LUT4 #(
		.INIT('h0100)
	) name1529 (
		_w1145_,
		_w1259_,
		_w1262_,
		_w1308_,
		_w2489_
	);
	LUT3 #(
		.INIT('h57)
	) name1530 (
		_w1035_,
		_w1048_,
		_w1168_,
		_w2490_
	);
	LUT3 #(
		.INIT('h10)
	) name1531 (
		_w1045_,
		_w1141_,
		_w2490_,
		_w2491_
	);
	LUT4 #(
		.INIT('h0080)
	) name1532 (
		_w1044_,
		_w1208_,
		_w1215_,
		_w1257_,
		_w2492_
	);
	LUT4 #(
		.INIT('h8000)
	) name1533 (
		_w1254_,
		_w2489_,
		_w2491_,
		_w2492_,
		_w2493_
	);
	LUT2 #(
		.INIT('h4)
	) name1534 (
		_w1071_,
		_w1299_,
		_w2494_
	);
	LUT2 #(
		.INIT('h8)
	) name1535 (
		_w1298_,
		_w2494_,
		_w2495_
	);
	LUT4 #(
		.INIT('h8000)
	) name1536 (
		_w2484_,
		_w2488_,
		_w2493_,
		_w2495_,
		_w2496_
	);
	LUT4 #(
		.INIT('h2aaa)
	) name1537 (
		\u5_cke_r_reg/NET0131 ,
		_w1002_,
		_w1005_,
		_w1006_,
		_w2497_
	);
	LUT3 #(
		.INIT('hba)
	) name1538 (
		_w2482_,
		_w2496_,
		_w2497_,
		_w2498_
	);
	LUT2 #(
		.INIT('h2)
	) name1539 (
		\u5_state_reg[0]/NET0131 ,
		\u5_tmr_done_reg/NET0131 ,
		_w2499_
	);
	LUT3 #(
		.INIT('hb0)
	) name1540 (
		_w1207_,
		_w2490_,
		_w2499_,
		_w2500_
	);
	LUT3 #(
		.INIT('h2a)
	) name1541 (
		\wb_addr_i[21]_pad ,
		_w976_,
		_w1971_,
		_w2501_
	);
	LUT3 #(
		.INIT('h10)
	) name1542 (
		_w1970_,
		_w1976_,
		_w2501_,
		_w2502_
	);
	LUT3 #(
		.INIT('h2a)
	) name1543 (
		\wb_addr_i[20]_pad ,
		_w976_,
		_w1975_,
		_w2503_
	);
	LUT3 #(
		.INIT('h10)
	) name1544 (
		_w1972_,
		_w1974_,
		_w2503_,
		_w2504_
	);
	LUT3 #(
		.INIT('h2a)
	) name1545 (
		\wb_addr_i[19]_pad ,
		_w976_,
		_w1971_,
		_w2505_
	);
	LUT3 #(
		.INIT('h40)
	) name1546 (
		_w1970_,
		_w1976_,
		_w2505_,
		_w2506_
	);
	LUT4 #(
		.INIT('h5554)
	) name1547 (
		_w2424_,
		_w2502_,
		_w2504_,
		_w2506_,
		_w2507_
	);
	LUT3 #(
		.INIT('h02)
	) name1548 (
		\u1_acs_addr_reg[19]/P0001 ,
		\u5_cs_le_reg/P0001 ,
		wb_we_i_pad,
		_w2508_
	);
	LUT4 #(
		.INIT('h7f00)
	) name1549 (
		_w2419_,
		_w2420_,
		_w2421_,
		_w2508_,
		_w2509_
	);
	LUT3 #(
		.INIT('h01)
	) name1550 (
		\u1_acs_addr_reg[19]/P0001 ,
		\u5_cs_le_reg/P0001 ,
		wb_we_i_pad,
		_w2510_
	);
	LUT4 #(
		.INIT('h8000)
	) name1551 (
		_w2419_,
		_w2420_,
		_w2421_,
		_w2510_,
		_w2511_
	);
	LUT3 #(
		.INIT('hfe)
	) name1552 (
		_w2507_,
		_w2509_,
		_w2511_,
		_w2512_
	);
	LUT3 #(
		.INIT('h2a)
	) name1553 (
		\wb_addr_i[23]_pad ,
		_w976_,
		_w1975_,
		_w2513_
	);
	LUT3 #(
		.INIT('h10)
	) name1554 (
		_w1972_,
		_w1974_,
		_w2513_,
		_w2514_
	);
	LUT3 #(
		.INIT('h2a)
	) name1555 (
		\wb_addr_i[22]_pad ,
		_w976_,
		_w1971_,
		_w2515_
	);
	LUT3 #(
		.INIT('h40)
	) name1556 (
		_w1970_,
		_w1976_,
		_w2515_,
		_w2516_
	);
	LUT3 #(
		.INIT('h2a)
	) name1557 (
		\wb_addr_i[24]_pad ,
		_w976_,
		_w1971_,
		_w2517_
	);
	LUT4 #(
		.INIT('haebf)
	) name1558 (
		_w1970_,
		_w1976_,
		_w2515_,
		_w2517_,
		_w2518_
	);
	LUT3 #(
		.INIT('h45)
	) name1559 (
		_w2424_,
		_w2514_,
		_w2518_,
		_w2519_
	);
	LUT4 #(
		.INIT('hff60)
	) name1560 (
		\u1_acs_addr_reg[22]/P0001 ,
		_w2423_,
		_w2424_,
		_w2519_,
		_w2520_
	);
	LUT4 #(
		.INIT('h2aaa)
	) name1561 (
		_w1007_,
		_w1603_,
		_w1604_,
		_w1607_,
		_w2521_
	);
	LUT4 #(
		.INIT('h1055)
	) name1562 (
		\u5_cke_r_reg/NET0131 ,
		_w1539_,
		_w1599_,
		_w2521_,
		_w2522_
	);
	LUT4 #(
		.INIT('ha800)
	) name1563 (
		_w1132_,
		_w1564_,
		_w1566_,
		_w2521_,
		_w2523_
	);
	LUT4 #(
		.INIT('h1055)
	) name1564 (
		_w1141_,
		_w1539_,
		_w1599_,
		_w2523_,
		_w2524_
	);
	LUT2 #(
		.INIT('h4)
	) name1565 (
		\u5_cke_r_reg/NET0131 ,
		\u5_cnt_reg/NET0131 ,
		_w2525_
	);
	LUT4 #(
		.INIT('h0070)
	) name1566 (
		\u5_cke_r_reg/NET0131 ,
		\u5_cnt_reg/NET0131 ,
		wb_cyc_i_pad,
		wb_stb_i_pad,
		_w2526_
	);
	LUT4 #(
		.INIT('h010f)
	) name1567 (
		_w1564_,
		_w1566_,
		_w2525_,
		_w2526_,
		_w2527_
	);
	LUT3 #(
		.INIT('h08)
	) name1568 (
		_w1100_,
		_w1140_,
		_w2527_,
		_w2528_
	);
	LUT2 #(
		.INIT('h1)
	) name1569 (
		_w1145_,
		_w2528_,
		_w2529_
	);
	LUT3 #(
		.INIT('h0b)
	) name1570 (
		_w2522_,
		_w2524_,
		_w2529_,
		_w2530_
	);
	LUT3 #(
		.INIT('h10)
	) name1571 (
		_w1141_,
		_w1145_,
		_w1299_,
		_w2531_
	);
	LUT3 #(
		.INIT('h40)
	) name1572 (
		_w1051_,
		_w1298_,
		_w2531_,
		_w2532_
	);
	LUT4 #(
		.INIT('h8000)
	) name1573 (
		_w2484_,
		_w2488_,
		_w2493_,
		_w2532_,
		_w2533_
	);
	LUT2 #(
		.INIT('h1)
	) name1574 (
		_w2530_,
		_w2533_,
		_w2534_
	);
	LUT3 #(
		.INIT('hb0)
	) name1575 (
		_w1539_,
		_w2162_,
		_w2383_,
		_w2535_
	);
	LUT3 #(
		.INIT('h80)
	) name1576 (
		_w1540_,
		_w1541_,
		_w2117_,
		_w2536_
	);
	LUT2 #(
		.INIT('h1)
	) name1577 (
		\u5_state_reg[40]/NET0131 ,
		_w2402_,
		_w2537_
	);
	LUT4 #(
		.INIT('h7f00)
	) name1578 (
		_w2398_,
		_w2399_,
		_w2400_,
		_w2402_,
		_w2538_
	);
	LUT4 #(
		.INIT('hbeaf)
	) name1579 (
		\u5_state_reg[40]/NET0131 ,
		\u5_timer2_reg[4]/P0001 ,
		\u5_timer2_reg[5]/P0001 ,
		_w2398_,
		_w2539_
	);
	LUT3 #(
		.INIT('h51)
	) name1580 (
		\u5_state_reg[51]/NET0131 ,
		_w2538_,
		_w2539_,
		_w2540_
	);
	LUT4 #(
		.INIT('h4f00)
	) name1581 (
		_w1539_,
		_w2536_,
		_w2537_,
		_w2540_,
		_w2541_
	);
	LUT4 #(
		.INIT('h0001)
	) name1582 (
		_w1214_,
		_w2389_,
		_w2409_,
		_w2413_,
		_w2542_
	);
	LUT2 #(
		.INIT('h2)
	) name1583 (
		\u5_state_reg[51]/NET0131 ,
		_w2149_,
		_w2543_
	);
	LUT3 #(
		.INIT('h80)
	) name1584 (
		_w1540_,
		_w1541_,
		_w2543_,
		_w2544_
	);
	LUT3 #(
		.INIT('h8c)
	) name1585 (
		_w1539_,
		_w2542_,
		_w2544_,
		_w2545_
	);
	LUT3 #(
		.INIT('hba)
	) name1586 (
		_w2535_,
		_w2541_,
		_w2545_,
		_w2546_
	);
	LUT4 #(
		.INIT('h8000)
	) name1587 (
		\u1_acs_addr_reg[19]/P0001 ,
		_w2419_,
		_w2420_,
		_w2421_,
		_w2547_
	);
	LUT3 #(
		.INIT('h10)
	) name1588 (
		_w1970_,
		_w1976_,
		_w2515_,
		_w2548_
	);
	LUT4 #(
		.INIT('h0e0f)
	) name1589 (
		_w1970_,
		_w1976_,
		_w2424_,
		_w2515_,
		_w2549_
	);
	LUT3 #(
		.INIT('h2a)
	) name1590 (
		\wb_addr_i[21]_pad ,
		_w976_,
		_w1975_,
		_w2550_
	);
	LUT3 #(
		.INIT('h10)
	) name1591 (
		_w1972_,
		_w1974_,
		_w2550_,
		_w2551_
	);
	LUT3 #(
		.INIT('h2a)
	) name1592 (
		\wb_addr_i[20]_pad ,
		_w976_,
		_w1971_,
		_w2552_
	);
	LUT3 #(
		.INIT('h40)
	) name1593 (
		_w1970_,
		_w1976_,
		_w2552_,
		_w2553_
	);
	LUT3 #(
		.INIT('h02)
	) name1594 (
		_w2549_,
		_w2551_,
		_w2553_,
		_w2554_
	);
	LUT4 #(
		.INIT('h007b)
	) name1595 (
		\u1_acs_addr_reg[20]/P0001 ,
		_w2424_,
		_w2547_,
		_w2554_,
		_w2555_
	);
	LUT3 #(
		.INIT('h01)
	) name1596 (
		_w1214_,
		_w2389_,
		_w2413_,
		_w2556_
	);
	LUT3 #(
		.INIT('hb0)
	) name1597 (
		_w1539_,
		_w1697_,
		_w2409_,
		_w2557_
	);
	LUT3 #(
		.INIT('h08)
	) name1598 (
		_w1540_,
		_w1541_,
		_w2108_,
		_w2558_
	);
	LUT3 #(
		.INIT('h8a)
	) name1599 (
		\u5_state_reg[51]/NET0131 ,
		_w1539_,
		_w2558_,
		_w2559_
	);
	LUT3 #(
		.INIT('ha8)
	) name1600 (
		_w2556_,
		_w2557_,
		_w2559_,
		_w2560_
	);
	LUT3 #(
		.INIT('h8a)
	) name1601 (
		\u5_state_reg[40]/NET0131 ,
		_w1539_,
		_w1893_,
		_w2561_
	);
	LUT3 #(
		.INIT('h01)
	) name1602 (
		\u5_state_reg[36]/NET0131 ,
		\u5_state_reg[43]/NET0131 ,
		\u5_state_reg[45]/NET0131 ,
		_w2562_
	);
	LUT2 #(
		.INIT('h8)
	) name1603 (
		_w962_,
		_w2562_,
		_w2563_
	);
	LUT4 #(
		.INIT('ha600)
	) name1604 (
		\u5_timer2_reg[4]/P0001 ,
		_w2398_,
		_w2401_,
		_w2563_,
		_w2564_
	);
	LUT4 #(
		.INIT('h004f)
	) name1605 (
		_w1539_,
		_w1918_,
		_w2537_,
		_w2564_,
		_w2565_
	);
	LUT4 #(
		.INIT('h1555)
	) name1606 (
		\u5_state_reg[51]/NET0131 ,
		\u5_tmr2_done_reg/NET0131 ,
		_w1041_,
		_w1091_,
		_w2566_
	);
	LUT4 #(
		.INIT('h0100)
	) name1607 (
		_w1214_,
		_w2389_,
		_w2413_,
		_w2566_,
		_w2567_
	);
	LUT3 #(
		.INIT('hb0)
	) name1608 (
		_w2561_,
		_w2565_,
		_w2567_,
		_w2568_
	);
	LUT3 #(
		.INIT('hb0)
	) name1609 (
		_w1539_,
		_w2122_,
		_w2383_,
		_w2569_
	);
	LUT3 #(
		.INIT('hfe)
	) name1610 (
		_w2560_,
		_w2568_,
		_w2569_,
		_w2570_
	);
	LUT2 #(
		.INIT('h2)
	) name1611 (
		\u1_bank_adr_reg[0]/P0001 ,
		\u1_bank_adr_reg[1]/P0001 ,
		_w2571_
	);
	LUT3 #(
		.INIT('h80)
	) name1612 (
		\u5_state_reg[7]/NET0131 ,
		_w976_,
		_w1118_,
		_w2572_
	);
	LUT2 #(
		.INIT('h8)
	) name1613 (
		\u0_sp_csc_reg[10]/NET0131 ,
		\u5_state_reg[7]/NET0131 ,
		_w2573_
	);
	LUT3 #(
		.INIT('h70)
	) name1614 (
		_w976_,
		_w1114_,
		_w2573_,
		_w2574_
	);
	LUT3 #(
		.INIT('ha8)
	) name1615 (
		_w2571_,
		_w2572_,
		_w2574_,
		_w2575_
	);
	LUT2 #(
		.INIT('h8)
	) name1616 (
		_w1533_,
		_w2575_,
		_w2576_
	);
	LUT3 #(
		.INIT('ha8)
	) name1617 (
		\u5_state_reg[22]/NET0131 ,
		\u5_state_reg[26]/NET0131 ,
		\u5_state_reg[27]/NET0131 ,
		_w2577_
	);
	LUT3 #(
		.INIT('h01)
	) name1618 (
		\u5_state_reg[23]/NET0131 ,
		\u5_state_reg[24]/NET0131 ,
		\u5_state_reg[25]/NET0131 ,
		_w2578_
	);
	LUT3 #(
		.INIT('h20)
	) name1619 (
		_w977_,
		_w2577_,
		_w2578_,
		_w2579_
	);
	LUT3 #(
		.INIT('h41)
	) name1620 (
		\u5_state_reg[22]/NET0131 ,
		\u5_state_reg[26]/NET0131 ,
		\u5_state_reg[27]/NET0131 ,
		_w2580_
	);
	LUT3 #(
		.INIT('h01)
	) name1621 (
		\u5_state_reg[21]/NET0131 ,
		\u5_state_reg[34]/NET0131 ,
		\u5_state_reg[35]/NET0131 ,
		_w2581_
	);
	LUT3 #(
		.INIT('h20)
	) name1622 (
		_w972_,
		_w2580_,
		_w2581_,
		_w2582_
	);
	LUT4 #(
		.INIT('h0001)
	) name1623 (
		\u5_state_reg[36]/NET0131 ,
		\u5_state_reg[37]/NET0131 ,
		\u5_state_reg[44]/NET0131 ,
		\u5_state_reg[45]/NET0131 ,
		_w2583_
	);
	LUT4 #(
		.INIT('h8000)
	) name1624 (
		_w963_,
		_w970_,
		_w992_,
		_w2583_,
		_w2584_
	);
	LUT4 #(
		.INIT('h0001)
	) name1625 (
		\u5_state_reg[42]/NET0131 ,
		\u5_state_reg[43]/NET0131 ,
		\u5_state_reg[60]/NET0131 ,
		\u5_state_reg[61]/NET0131 ,
		_w2585_
	);
	LUT4 #(
		.INIT('h8000)
	) name1626 (
		_w985_,
		_w999_,
		_w1175_,
		_w2585_,
		_w2586_
	);
	LUT4 #(
		.INIT('h8000)
	) name1627 (
		_w2579_,
		_w2582_,
		_w2584_,
		_w2586_,
		_w2587_
	);
	LUT3 #(
		.INIT('h01)
	) name1628 (
		\u5_state_reg[18]/NET0131 ,
		\u5_state_reg[19]/NET0131 ,
		\u5_state_reg[20]/NET0131 ,
		_w2588_
	);
	LUT3 #(
		.INIT('h01)
	) name1629 (
		\u5_state_reg[12]/NET0131 ,
		\u5_state_reg[13]/NET0131 ,
		\u5_state_reg[7]/NET0131 ,
		_w2589_
	);
	LUT4 #(
		.INIT('h0001)
	) name1630 (
		\u5_state_reg[0]/NET0131 ,
		\u5_state_reg[1]/NET0131 ,
		\u5_state_reg[5]/NET0131 ,
		\u5_state_reg[6]/NET0131 ,
		_w2590_
	);
	LUT2 #(
		.INIT('h8)
	) name1631 (
		_w2589_,
		_w2590_,
		_w2591_
	);
	LUT3 #(
		.INIT('h80)
	) name1632 (
		_w980_,
		_w1003_,
		_w1020_,
		_w2592_
	);
	LUT2 #(
		.INIT('h8)
	) name1633 (
		_w2591_,
		_w2592_,
		_w2593_
	);
	LUT3 #(
		.INIT('h80)
	) name1634 (
		_w2587_,
		_w2588_,
		_w2593_,
		_w2594_
	);
	LUT3 #(
		.INIT('hec)
	) name1635 (
		\u5_state_reg[18]/NET0131 ,
		\u5_state_reg[19]/NET0131 ,
		\u5_state_reg[20]/NET0131 ,
		_w2595_
	);
	LUT3 #(
		.INIT('h0d)
	) name1636 (
		\u5_state_reg[18]/NET0131 ,
		\u5_state_reg[19]/NET0131 ,
		\u5_state_reg[20]/NET0131 ,
		_w2596_
	);
	LUT3 #(
		.INIT('h23)
	) name1637 (
		_w2587_,
		_w2595_,
		_w2596_,
		_w2597_
	);
	LUT3 #(
		.INIT('h01)
	) name1638 (
		\u5_state_reg[27]/NET0131 ,
		\u5_state_reg[28]/NET0131 ,
		\u5_state_reg[29]/NET0131 ,
		_w2598_
	);
	LUT2 #(
		.INIT('h8)
	) name1639 (
		_w2586_,
		_w2598_,
		_w2599_
	);
	LUT4 #(
		.INIT('h0001)
	) name1640 (
		\u5_state_reg[21]/NET0131 ,
		\u5_state_reg[22]/NET0131 ,
		\u5_state_reg[23]/NET0131 ,
		\u5_state_reg[24]/NET0131 ,
		_w2600_
	);
	LUT2 #(
		.INIT('h1)
	) name1641 (
		\u5_state_reg[25]/NET0131 ,
		\u5_state_reg[26]/NET0131 ,
		_w2601_
	);
	LUT4 #(
		.INIT('h8000)
	) name1642 (
		_w1026_,
		_w1030_,
		_w2600_,
		_w2601_,
		_w2602_
	);
	LUT4 #(
		.INIT('h8000)
	) name1643 (
		_w2584_,
		_w2586_,
		_w2598_,
		_w2602_,
		_w2603_
	);
	LUT2 #(
		.INIT('h8)
	) name1644 (
		_w2593_,
		_w2603_,
		_w2604_
	);
	LUT4 #(
		.INIT('ha888)
	) name1645 (
		_w1533_,
		_w2594_,
		_w2597_,
		_w2604_,
		_w2605_
	);
	LUT3 #(
		.INIT('h10)
	) name1646 (
		\u5_rfr_ack_r_reg/NET0131 ,
		\u5_state_reg[16]/NET0131 ,
		\u5_state_reg[4]/NET0131 ,
		_w2606_
	);
	LUT3 #(
		.INIT('h20)
	) name1647 (
		\u5_state_reg[16]/NET0131 ,
		\u5_state_reg[4]/NET0131 ,
		\u5_tmr_done_reg/NET0131 ,
		_w2607_
	);
	LUT3 #(
		.INIT('h70)
	) name1648 (
		_w976_,
		_w1118_,
		_w2607_,
		_w2608_
	);
	LUT3 #(
		.INIT('h23)
	) name1649 (
		_w1117_,
		_w2606_,
		_w2608_,
		_w2609_
	);
	LUT3 #(
		.INIT('he0)
	) name1650 (
		_w1526_,
		_w1531_,
		_w2571_,
		_w2610_
	);
	LUT3 #(
		.INIT('h10)
	) name1651 (
		_w1528_,
		_w1530_,
		_w2610_,
		_w2611_
	);
	LUT4 #(
		.INIT('h2022)
	) name1652 (
		\u2_u0_bank1_open_reg/NET0131 ,
		\u5_rfr_ack_r_reg/NET0131 ,
		_w2609_,
		_w2611_,
		_w2612_
	);
	LUT3 #(
		.INIT('hba)
	) name1653 (
		_w2576_,
		_w2605_,
		_w2612_,
		_w2613_
	);
	LUT2 #(
		.INIT('h4)
	) name1654 (
		\u1_bank_adr_reg[0]/P0001 ,
		\u1_bank_adr_reg[1]/P0001 ,
		_w2614_
	);
	LUT3 #(
		.INIT('he0)
	) name1655 (
		_w2572_,
		_w2574_,
		_w2614_,
		_w2615_
	);
	LUT2 #(
		.INIT('h8)
	) name1656 (
		_w1533_,
		_w2615_,
		_w2616_
	);
	LUT3 #(
		.INIT('he0)
	) name1657 (
		_w1526_,
		_w1531_,
		_w2614_,
		_w2617_
	);
	LUT3 #(
		.INIT('h10)
	) name1658 (
		_w1528_,
		_w1530_,
		_w2617_,
		_w2618_
	);
	LUT4 #(
		.INIT('h2022)
	) name1659 (
		\u2_u0_bank2_open_reg/NET0131 ,
		\u5_rfr_ack_r_reg/NET0131 ,
		_w2609_,
		_w2618_,
		_w2619_
	);
	LUT3 #(
		.INIT('hdc)
	) name1660 (
		_w2605_,
		_w2616_,
		_w2619_,
		_w2620_
	);
	LUT2 #(
		.INIT('h4)
	) name1661 (
		_w1579_,
		_w2615_,
		_w2621_
	);
	LUT4 #(
		.INIT('h5444)
	) name1662 (
		_w1579_,
		_w2594_,
		_w2597_,
		_w2604_,
		_w2622_
	);
	LUT4 #(
		.INIT('ha8aa)
	) name1663 (
		\u2_u1_bank2_open_reg/NET0131 ,
		_w1579_,
		_w2609_,
		_w2614_,
		_w2623_
	);
	LUT2 #(
		.INIT('h4)
	) name1664 (
		\u5_rfr_ack_r_reg/NET0131 ,
		_w2623_,
		_w2624_
	);
	LUT3 #(
		.INIT('hba)
	) name1665 (
		_w2621_,
		_w2622_,
		_w2624_,
		_w2625_
	);
	LUT2 #(
		.INIT('h4)
	) name1666 (
		_w1579_,
		_w2575_,
		_w2626_
	);
	LUT4 #(
		.INIT('haa8a)
	) name1667 (
		\u2_u1_bank1_open_reg/NET0131 ,
		_w1579_,
		_w2571_,
		_w2609_,
		_w2627_
	);
	LUT2 #(
		.INIT('h4)
	) name1668 (
		\u5_rfr_ack_r_reg/NET0131 ,
		_w2627_,
		_w2628_
	);
	LUT3 #(
		.INIT('hdc)
	) name1669 (
		_w2622_,
		_w2626_,
		_w2628_,
		_w2629_
	);
	LUT4 #(
		.INIT('h6aff)
	) name1670 (
		\u1_acs_addr_reg[16]/P0001 ,
		_w2419_,
		_w2420_,
		_w2424_,
		_w2630_
	);
	LUT3 #(
		.INIT('h2a)
	) name1671 (
		\wb_addr_i[16]_pad ,
		_w976_,
		_w1971_,
		_w2631_
	);
	LUT3 #(
		.INIT('h40)
	) name1672 (
		_w1970_,
		_w1976_,
		_w2631_,
		_w2632_
	);
	LUT4 #(
		.INIT('h0b0f)
	) name1673 (
		_w1970_,
		_w1976_,
		_w2424_,
		_w2631_,
		_w2633_
	);
	LUT3 #(
		.INIT('h2a)
	) name1674 (
		\wb_addr_i[18]_pad ,
		_w976_,
		_w1971_,
		_w2634_
	);
	LUT3 #(
		.INIT('h10)
	) name1675 (
		_w1970_,
		_w1976_,
		_w2634_,
		_w2635_
	);
	LUT3 #(
		.INIT('h2a)
	) name1676 (
		\wb_addr_i[17]_pad ,
		_w976_,
		_w1975_,
		_w2636_
	);
	LUT3 #(
		.INIT('h10)
	) name1677 (
		_w1972_,
		_w1974_,
		_w2636_,
		_w2637_
	);
	LUT3 #(
		.INIT('h02)
	) name1678 (
		_w2633_,
		_w2635_,
		_w2637_,
		_w2638_
	);
	LUT2 #(
		.INIT('h2)
	) name1679 (
		_w2630_,
		_w2638_,
		_w2639_
	);
	LUT2 #(
		.INIT('h8)
	) name1680 (
		\u1_bank_adr_reg[0]/P0001 ,
		\u1_bank_adr_reg[1]/P0001 ,
		_w2640_
	);
	LUT3 #(
		.INIT('he0)
	) name1681 (
		_w2572_,
		_w2574_,
		_w2640_,
		_w2641_
	);
	LUT2 #(
		.INIT('h8)
	) name1682 (
		_w1533_,
		_w2641_,
		_w2642_
	);
	LUT3 #(
		.INIT('he0)
	) name1683 (
		_w1526_,
		_w1531_,
		_w2640_,
		_w2643_
	);
	LUT3 #(
		.INIT('h10)
	) name1684 (
		_w1528_,
		_w1530_,
		_w2643_,
		_w2644_
	);
	LUT4 #(
		.INIT('h2022)
	) name1685 (
		\u2_u0_bank3_open_reg/NET0131 ,
		\u5_rfr_ack_r_reg/NET0131 ,
		_w2609_,
		_w2644_,
		_w2645_
	);
	LUT3 #(
		.INIT('hdc)
	) name1686 (
		_w2605_,
		_w2642_,
		_w2645_,
		_w2646_
	);
	LUT2 #(
		.INIT('h4)
	) name1687 (
		_w1579_,
		_w2641_,
		_w2647_
	);
	LUT4 #(
		.INIT('ha8aa)
	) name1688 (
		\u2_u1_bank3_open_reg/NET0131 ,
		_w1579_,
		_w2609_,
		_w2640_,
		_w2648_
	);
	LUT2 #(
		.INIT('h4)
	) name1689 (
		\u5_rfr_ack_r_reg/NET0131 ,
		_w2648_,
		_w2649_
	);
	LUT3 #(
		.INIT('hdc)
	) name1690 (
		_w2622_,
		_w2647_,
		_w2649_,
		_w2650_
	);
	LUT3 #(
		.INIT('h2a)
	) name1691 (
		\wb_addr_i[19]_pad ,
		_w976_,
		_w1975_,
		_w2651_
	);
	LUT3 #(
		.INIT('h10)
	) name1692 (
		_w1972_,
		_w1974_,
		_w2651_,
		_w2652_
	);
	LUT3 #(
		.INIT('h40)
	) name1693 (
		_w1970_,
		_w1976_,
		_w2634_,
		_w2653_
	);
	LUT3 #(
		.INIT('h10)
	) name1694 (
		_w1970_,
		_w1976_,
		_w2552_,
		_w2654_
	);
	LUT4 #(
		.INIT('habef)
	) name1695 (
		_w1970_,
		_w1976_,
		_w2552_,
		_w2634_,
		_w2655_
	);
	LUT3 #(
		.INIT('h45)
	) name1696 (
		_w2424_,
		_w2652_,
		_w2655_,
		_w2656_
	);
	LUT2 #(
		.INIT('h8)
	) name1697 (
		\u1_acs_addr_reg[16]/P0001 ,
		\u1_acs_addr_reg[17]/P0001 ,
		_w2657_
	);
	LUT4 #(
		.INIT('h1555)
	) name1698 (
		\u1_acs_addr_reg[18]/P0001 ,
		_w2419_,
		_w2420_,
		_w2657_,
		_w2658_
	);
	LUT4 #(
		.INIT('h7f00)
	) name1699 (
		_w2419_,
		_w2420_,
		_w2421_,
		_w2424_,
		_w2659_
	);
	LUT3 #(
		.INIT('hba)
	) name1700 (
		_w2656_,
		_w2658_,
		_w2659_,
		_w2660_
	);
	LUT3 #(
		.INIT('h8c)
	) name1701 (
		_w1539_,
		_w2383_,
		_w2448_,
		_w2661_
	);
	LUT2 #(
		.INIT('h8)
	) name1702 (
		\u5_state_reg[51]/NET0131 ,
		_w1709_,
		_w2662_
	);
	LUT3 #(
		.INIT('h80)
	) name1703 (
		_w1540_,
		_w1541_,
		_w2662_,
		_w2663_
	);
	LUT4 #(
		.INIT('h1555)
	) name1704 (
		\u5_timer2_reg[0]/P0001 ,
		_w2398_,
		_w2399_,
		_w2400_,
		_w2664_
	);
	LUT3 #(
		.INIT('h02)
	) name1705 (
		\u5_timer2_reg[0]/P0001 ,
		\u5_timer2_reg[7]/P0001 ,
		\u5_timer2_reg[8]/P0001 ,
		_w2665_
	);
	LUT3 #(
		.INIT('h80)
	) name1706 (
		_w2398_,
		_w2399_,
		_w2665_,
		_w2666_
	);
	LUT2 #(
		.INIT('h8)
	) name1707 (
		_w2397_,
		_w2402_,
		_w2667_
	);
	LUT3 #(
		.INIT('h10)
	) name1708 (
		_w2664_,
		_w2666_,
		_w2667_,
		_w2668_
	);
	LUT4 #(
		.INIT('h007f)
	) name1709 (
		\u5_tmr2_done_reg/NET0131 ,
		_w1041_,
		_w1091_,
		_w2668_,
		_w2669_
	);
	LUT4 #(
		.INIT('h1033)
	) name1710 (
		_w1539_,
		_w2389_,
		_w2663_,
		_w2669_,
		_w2670_
	);
	LUT4 #(
		.INIT('h8000)
	) name1711 (
		_w1041_,
		_w2137_,
		_w2387_,
		_w2388_,
		_w2671_
	);
	LUT3 #(
		.INIT('h80)
	) name1712 (
		_w1540_,
		_w1541_,
		_w2671_,
		_w2672_
	);
	LUT3 #(
		.INIT('h8c)
	) name1713 (
		_w1539_,
		_w2414_,
		_w2672_,
		_w2673_
	);
	LUT3 #(
		.INIT('hba)
	) name1714 (
		_w2661_,
		_w2670_,
		_w2673_,
		_w2674_
	);
	LUT3 #(
		.INIT('hb0)
	) name1715 (
		_w1539_,
		_w1694_,
		_w2383_,
		_w2675_
	);
	LUT2 #(
		.INIT('h2)
	) name1716 (
		_w2156_,
		_w2402_,
		_w2676_
	);
	LUT3 #(
		.INIT('h80)
	) name1717 (
		_w1540_,
		_w1541_,
		_w2676_,
		_w2677_
	);
	LUT3 #(
		.INIT('h08)
	) name1718 (
		_w2398_,
		_w2399_,
		_w2400_,
		_w2678_
	);
	LUT2 #(
		.INIT('h1)
	) name1719 (
		\u5_timer2_reg[4]/P0001 ,
		\u5_timer2_reg[5]/P0001 ,
		_w2679_
	);
	LUT4 #(
		.INIT('hd050)
	) name1720 (
		\u5_timer2_reg[6]/P0001 ,
		_w2398_,
		_w2402_,
		_w2679_,
		_w2680_
	);
	LUT3 #(
		.INIT('h8a)
	) name1721 (
		_w2397_,
		_w2678_,
		_w2680_,
		_w2681_
	);
	LUT4 #(
		.INIT('h8c00)
	) name1722 (
		_w1539_,
		_w2542_,
		_w2677_,
		_w2681_,
		_w2682_
	);
	LUT2 #(
		.INIT('he)
	) name1723 (
		_w2675_,
		_w2682_,
		_w2683_
	);
	LUT3 #(
		.INIT('h2a)
	) name1724 (
		\u0_sp_tms_reg[0]/NET0131 ,
		wb_cyc_i_pad,
		wb_stb_i_pad,
		_w2684_
	);
	LUT3 #(
		.INIT('h10)
	) name1725 (
		\u4_rfr_req_reg/NET0131 ,
		\u5_state_reg[0]/NET0131 ,
		\u5_state_reg[1]/NET0131 ,
		_w2685_
	);
	LUT2 #(
		.INIT('h8)
	) name1726 (
		_w1184_,
		_w2685_,
		_w2686_
	);
	LUT4 #(
		.INIT('h2220)
	) name1727 (
		\u5_lookup_ready2_reg/NET0131 ,
		_w1335_,
		_w1564_,
		_w1566_,
		_w2687_
	);
	LUT4 #(
		.INIT('h20aa)
	) name1728 (
		\u5_wb_stb_first_reg/NET0131 ,
		_w1533_,
		_w1579_,
		_w2687_,
		_w2688_
	);
	LUT3 #(
		.INIT('h8a)
	) name1729 (
		\u5_lookup_ready2_reg/NET0131 ,
		_w1533_,
		_w1579_,
		_w2689_
	);
	LUT3 #(
		.INIT('h54)
	) name1730 (
		_w1132_,
		_w1564_,
		_w1566_,
		_w2690_
	);
	LUT2 #(
		.INIT('h8)
	) name1731 (
		_w2020_,
		_w2690_,
		_w2691_
	);
	LUT4 #(
		.INIT('h0222)
	) name1732 (
		_w1628_,
		_w2688_,
		_w2689_,
		_w2691_,
		_w2692_
	);
	LUT2 #(
		.INIT('h2)
	) name1733 (
		_w2686_,
		_w2692_,
		_w2693_
	);
	LUT4 #(
		.INIT('h02aa)
	) name1734 (
		\u5_tmr2_done_reg/NET0131 ,
		_w1564_,
		_w1566_,
		_w2028_,
		_w2694_
	);
	LUT3 #(
		.INIT('h80)
	) name1735 (
		_w1002_,
		_w1166_,
		_w2694_,
		_w2695_
	);
	LUT4 #(
		.INIT('h222a)
	) name1736 (
		\u5_tmr_done_reg/NET0131 ,
		_w1132_,
		_w1564_,
		_w1566_,
		_w2696_
	);
	LUT3 #(
		.INIT('h80)
	) name1737 (
		_w1002_,
		_w1274_,
		_w2696_,
		_w2697_
	);
	LUT4 #(
		.INIT('haaa8)
	) name1738 (
		\u5_wb_cycle_reg/NET0131 ,
		_w1095_,
		_w2695_,
		_w2697_,
		_w2698_
	);
	LUT3 #(
		.INIT('h57)
	) name1739 (
		_w1041_,
		_w1043_,
		_w1256_,
		_w2699_
	);
	LUT2 #(
		.INIT('h4)
	) name1740 (
		_w2194_,
		_w2699_,
		_w2700_
	);
	LUT4 #(
		.INIT('h0800)
	) name1741 (
		_w1100_,
		_w1277_,
		_w1956_,
		_w2690_,
		_w2701_
	);
	LUT4 #(
		.INIT('h2000)
	) name1742 (
		\u4_rfr_req_reg/NET0131 ,
		\u5_state_reg[0]/NET0131 ,
		\u5_state_reg[1]/NET0131 ,
		\u5_wb_stb_first_reg/NET0131 ,
		_w2702_
	);
	LUT2 #(
		.INIT('h8)
	) name1743 (
		_w1184_,
		_w2702_,
		_w2703_
	);
	LUT4 #(
		.INIT('h0777)
	) name1744 (
		_w1035_,
		_w1097_,
		_w1100_,
		_w1102_,
		_w2704_
	);
	LUT3 #(
		.INIT('h10)
	) name1745 (
		_w2701_,
		_w2703_,
		_w2704_,
		_w2705_
	);
	LUT3 #(
		.INIT('h40)
	) name1746 (
		_w2698_,
		_w2700_,
		_w2705_,
		_w2706_
	);
	LUT2 #(
		.INIT('hb)
	) name1747 (
		_w2693_,
		_w2706_,
		_w2707_
	);
	LUT2 #(
		.INIT('h4)
	) name1748 (
		\u0_rf_we_reg/NET0131 ,
		\u0_sp_tms_reg[0]/NET0131 ,
		_w2708_
	);
	LUT4 #(
		.INIT('h4555)
	) name1749 (
		_w2684_,
		_w2693_,
		_w2706_,
		_w2708_,
		_w2709_
	);
	LUT2 #(
		.INIT('h4)
	) name1750 (
		\u0_spec_req_cs_reg[0]/NET0131 ,
		\u0_spec_req_cs_reg[1]/NET0131 ,
		_w2710_
	);
	LUT4 #(
		.INIT('h1b5f)
	) name1751 (
		\u0_spec_req_cs_reg[0]/NET0131 ,
		\u0_spec_req_cs_reg[1]/NET0131 ,
		\u0_u0_tms_reg[0]/P0001 ,
		\u0_u1_tms_reg[0]/P0001 ,
		_w2711_
	);
	LUT2 #(
		.INIT('h2)
	) name1752 (
		_w1013_,
		_w2711_,
		_w2712_
	);
	LUT4 #(
		.INIT('hef00)
	) name1753 (
		\u0_rf_we_reg/NET0131 ,
		_w2693_,
		_w2706_,
		_w2712_,
		_w2713_
	);
	LUT2 #(
		.INIT('hd)
	) name1754 (
		_w2709_,
		_w2713_,
		_w2714_
	);
	LUT3 #(
		.INIT('h2a)
	) name1755 (
		\u0_sp_tms_reg[10]/NET0131 ,
		wb_cyc_i_pad,
		wb_stb_i_pad,
		_w2715_
	);
	LUT2 #(
		.INIT('h4)
	) name1756 (
		\u0_rf_we_reg/NET0131 ,
		\u0_sp_tms_reg[10]/NET0131 ,
		_w2716_
	);
	LUT4 #(
		.INIT('h0b0f)
	) name1757 (
		_w2693_,
		_w2706_,
		_w2715_,
		_w2716_,
		_w2717_
	);
	LUT4 #(
		.INIT('h1b5f)
	) name1758 (
		\u0_spec_req_cs_reg[0]/NET0131 ,
		\u0_spec_req_cs_reg[1]/NET0131 ,
		\u0_u0_tms_reg[10]/P0001 ,
		\u0_u1_tms_reg[10]/P0001 ,
		_w2718_
	);
	LUT2 #(
		.INIT('h2)
	) name1759 (
		_w1013_,
		_w2718_,
		_w2719_
	);
	LUT4 #(
		.INIT('hef00)
	) name1760 (
		\u0_rf_we_reg/NET0131 ,
		_w2693_,
		_w2706_,
		_w2719_,
		_w2720_
	);
	LUT2 #(
		.INIT('hd)
	) name1761 (
		_w2717_,
		_w2720_,
		_w2721_
	);
	LUT3 #(
		.INIT('h2a)
	) name1762 (
		\u0_sp_tms_reg[11]/NET0131 ,
		wb_cyc_i_pad,
		wb_stb_i_pad,
		_w2722_
	);
	LUT2 #(
		.INIT('h4)
	) name1763 (
		\u0_rf_we_reg/NET0131 ,
		\u0_sp_tms_reg[11]/NET0131 ,
		_w2723_
	);
	LUT4 #(
		.INIT('h0b0f)
	) name1764 (
		_w2693_,
		_w2706_,
		_w2722_,
		_w2723_,
		_w2724_
	);
	LUT4 #(
		.INIT('h1b5f)
	) name1765 (
		\u0_spec_req_cs_reg[0]/NET0131 ,
		\u0_spec_req_cs_reg[1]/NET0131 ,
		\u0_u0_tms_reg[11]/P0001 ,
		\u0_u1_tms_reg[11]/P0001 ,
		_w2725_
	);
	LUT2 #(
		.INIT('h2)
	) name1766 (
		_w1013_,
		_w2725_,
		_w2726_
	);
	LUT4 #(
		.INIT('hef00)
	) name1767 (
		\u0_rf_we_reg/NET0131 ,
		_w2693_,
		_w2706_,
		_w2726_,
		_w2727_
	);
	LUT2 #(
		.INIT('hd)
	) name1768 (
		_w2724_,
		_w2727_,
		_w2728_
	);
	LUT3 #(
		.INIT('h2a)
	) name1769 (
		\u0_sp_tms_reg[12]/NET0131 ,
		wb_cyc_i_pad,
		wb_stb_i_pad,
		_w2729_
	);
	LUT2 #(
		.INIT('h4)
	) name1770 (
		\u0_rf_we_reg/NET0131 ,
		\u0_sp_tms_reg[12]/NET0131 ,
		_w2730_
	);
	LUT4 #(
		.INIT('h0b0f)
	) name1771 (
		_w2693_,
		_w2706_,
		_w2729_,
		_w2730_,
		_w2731_
	);
	LUT4 #(
		.INIT('h1b5f)
	) name1772 (
		\u0_spec_req_cs_reg[0]/NET0131 ,
		\u0_spec_req_cs_reg[1]/NET0131 ,
		\u0_u0_tms_reg[12]/P0001 ,
		\u0_u1_tms_reg[12]/P0001 ,
		_w2732_
	);
	LUT2 #(
		.INIT('h2)
	) name1773 (
		_w1013_,
		_w2732_,
		_w2733_
	);
	LUT4 #(
		.INIT('hef00)
	) name1774 (
		\u0_rf_we_reg/NET0131 ,
		_w2693_,
		_w2706_,
		_w2733_,
		_w2734_
	);
	LUT2 #(
		.INIT('hd)
	) name1775 (
		_w2731_,
		_w2734_,
		_w2735_
	);
	LUT3 #(
		.INIT('h2a)
	) name1776 (
		\u0_sp_tms_reg[14]/NET0131 ,
		wb_cyc_i_pad,
		wb_stb_i_pad,
		_w2736_
	);
	LUT2 #(
		.INIT('h4)
	) name1777 (
		\u0_rf_we_reg/NET0131 ,
		\u0_sp_tms_reg[14]/NET0131 ,
		_w2737_
	);
	LUT4 #(
		.INIT('h0b0f)
	) name1778 (
		_w2693_,
		_w2706_,
		_w2736_,
		_w2737_,
		_w2738_
	);
	LUT4 #(
		.INIT('h1b5f)
	) name1779 (
		\u0_spec_req_cs_reg[0]/NET0131 ,
		\u0_spec_req_cs_reg[1]/NET0131 ,
		\u0_u0_tms_reg[14]/P0001 ,
		\u0_u1_tms_reg[14]/P0001 ,
		_w2739_
	);
	LUT2 #(
		.INIT('h2)
	) name1780 (
		_w1013_,
		_w2739_,
		_w2740_
	);
	LUT4 #(
		.INIT('hef00)
	) name1781 (
		\u0_rf_we_reg/NET0131 ,
		_w2693_,
		_w2706_,
		_w2740_,
		_w2741_
	);
	LUT2 #(
		.INIT('hd)
	) name1782 (
		_w2738_,
		_w2741_,
		_w2742_
	);
	LUT3 #(
		.INIT('h2a)
	) name1783 (
		\u0_sp_tms_reg[13]/NET0131 ,
		wb_cyc_i_pad,
		wb_stb_i_pad,
		_w2743_
	);
	LUT2 #(
		.INIT('h4)
	) name1784 (
		\u0_rf_we_reg/NET0131 ,
		\u0_sp_tms_reg[13]/NET0131 ,
		_w2744_
	);
	LUT4 #(
		.INIT('h0b0f)
	) name1785 (
		_w2693_,
		_w2706_,
		_w2743_,
		_w2744_,
		_w2745_
	);
	LUT4 #(
		.INIT('h1b5f)
	) name1786 (
		\u0_spec_req_cs_reg[0]/NET0131 ,
		\u0_spec_req_cs_reg[1]/NET0131 ,
		\u0_u0_tms_reg[13]/P0001 ,
		\u0_u1_tms_reg[13]/P0001 ,
		_w2746_
	);
	LUT2 #(
		.INIT('h2)
	) name1787 (
		_w1013_,
		_w2746_,
		_w2747_
	);
	LUT4 #(
		.INIT('hef00)
	) name1788 (
		\u0_rf_we_reg/NET0131 ,
		_w2693_,
		_w2706_,
		_w2747_,
		_w2748_
	);
	LUT2 #(
		.INIT('hd)
	) name1789 (
		_w2745_,
		_w2748_,
		_w2749_
	);
	LUT3 #(
		.INIT('h2a)
	) name1790 (
		\u0_sp_tms_reg[16]/NET0131 ,
		wb_cyc_i_pad,
		wb_stb_i_pad,
		_w2750_
	);
	LUT2 #(
		.INIT('h4)
	) name1791 (
		\u0_rf_we_reg/NET0131 ,
		\u0_sp_tms_reg[16]/NET0131 ,
		_w2751_
	);
	LUT4 #(
		.INIT('h0b0f)
	) name1792 (
		_w2693_,
		_w2706_,
		_w2750_,
		_w2751_,
		_w2752_
	);
	LUT4 #(
		.INIT('h1b5f)
	) name1793 (
		\u0_spec_req_cs_reg[0]/NET0131 ,
		\u0_spec_req_cs_reg[1]/NET0131 ,
		\u0_u0_tms_reg[16]/P0001 ,
		\u0_u1_tms_reg[16]/P0001 ,
		_w2753_
	);
	LUT2 #(
		.INIT('h2)
	) name1794 (
		_w1013_,
		_w2753_,
		_w2754_
	);
	LUT4 #(
		.INIT('hef00)
	) name1795 (
		\u0_rf_we_reg/NET0131 ,
		_w2693_,
		_w2706_,
		_w2754_,
		_w2755_
	);
	LUT2 #(
		.INIT('hd)
	) name1796 (
		_w2752_,
		_w2755_,
		_w2756_
	);
	LUT3 #(
		.INIT('h2a)
	) name1797 (
		\u0_sp_tms_reg[17]/NET0131 ,
		wb_cyc_i_pad,
		wb_stb_i_pad,
		_w2757_
	);
	LUT2 #(
		.INIT('h4)
	) name1798 (
		\u0_rf_we_reg/NET0131 ,
		\u0_sp_tms_reg[17]/NET0131 ,
		_w2758_
	);
	LUT4 #(
		.INIT('h0b0f)
	) name1799 (
		_w2693_,
		_w2706_,
		_w2757_,
		_w2758_,
		_w2759_
	);
	LUT4 #(
		.INIT('h1b5f)
	) name1800 (
		\u0_spec_req_cs_reg[0]/NET0131 ,
		\u0_spec_req_cs_reg[1]/NET0131 ,
		\u0_u0_tms_reg[17]/P0001 ,
		\u0_u1_tms_reg[17]/P0001 ,
		_w2760_
	);
	LUT2 #(
		.INIT('h2)
	) name1801 (
		_w1013_,
		_w2760_,
		_w2761_
	);
	LUT4 #(
		.INIT('hef00)
	) name1802 (
		\u0_rf_we_reg/NET0131 ,
		_w2693_,
		_w2706_,
		_w2761_,
		_w2762_
	);
	LUT2 #(
		.INIT('hd)
	) name1803 (
		_w2759_,
		_w2762_,
		_w2763_
	);
	LUT3 #(
		.INIT('h2a)
	) name1804 (
		\u0_sp_tms_reg[18]/NET0131 ,
		wb_cyc_i_pad,
		wb_stb_i_pad,
		_w2764_
	);
	LUT2 #(
		.INIT('h4)
	) name1805 (
		\u0_rf_we_reg/NET0131 ,
		\u0_sp_tms_reg[18]/NET0131 ,
		_w2765_
	);
	LUT4 #(
		.INIT('h0b0f)
	) name1806 (
		_w2693_,
		_w2706_,
		_w2764_,
		_w2765_,
		_w2766_
	);
	LUT4 #(
		.INIT('h1b5f)
	) name1807 (
		\u0_spec_req_cs_reg[0]/NET0131 ,
		\u0_spec_req_cs_reg[1]/NET0131 ,
		\u0_u0_tms_reg[18]/P0001 ,
		\u0_u1_tms_reg[18]/P0001 ,
		_w2767_
	);
	LUT2 #(
		.INIT('h2)
	) name1808 (
		_w1013_,
		_w2767_,
		_w2768_
	);
	LUT4 #(
		.INIT('hef00)
	) name1809 (
		\u0_rf_we_reg/NET0131 ,
		_w2693_,
		_w2706_,
		_w2768_,
		_w2769_
	);
	LUT2 #(
		.INIT('hd)
	) name1810 (
		_w2766_,
		_w2769_,
		_w2770_
	);
	LUT3 #(
		.INIT('h2a)
	) name1811 (
		\u0_sp_tms_reg[19]/NET0131 ,
		wb_cyc_i_pad,
		wb_stb_i_pad,
		_w2771_
	);
	LUT2 #(
		.INIT('h4)
	) name1812 (
		\u0_rf_we_reg/NET0131 ,
		\u0_sp_tms_reg[19]/NET0131 ,
		_w2772_
	);
	LUT4 #(
		.INIT('h0b0f)
	) name1813 (
		_w2693_,
		_w2706_,
		_w2771_,
		_w2772_,
		_w2773_
	);
	LUT4 #(
		.INIT('h1b5f)
	) name1814 (
		\u0_spec_req_cs_reg[0]/NET0131 ,
		\u0_spec_req_cs_reg[1]/NET0131 ,
		\u0_u0_tms_reg[19]/P0001 ,
		\u0_u1_tms_reg[19]/P0001 ,
		_w2774_
	);
	LUT2 #(
		.INIT('h2)
	) name1815 (
		_w1013_,
		_w2774_,
		_w2775_
	);
	LUT4 #(
		.INIT('hef00)
	) name1816 (
		\u0_rf_we_reg/NET0131 ,
		_w2693_,
		_w2706_,
		_w2775_,
		_w2776_
	);
	LUT2 #(
		.INIT('hd)
	) name1817 (
		_w2773_,
		_w2776_,
		_w2777_
	);
	LUT3 #(
		.INIT('h2a)
	) name1818 (
		\u0_sp_tms_reg[15]/NET0131 ,
		wb_cyc_i_pad,
		wb_stb_i_pad,
		_w2778_
	);
	LUT2 #(
		.INIT('h4)
	) name1819 (
		\u0_rf_we_reg/NET0131 ,
		\u0_sp_tms_reg[15]/NET0131 ,
		_w2779_
	);
	LUT4 #(
		.INIT('h0b0f)
	) name1820 (
		_w2693_,
		_w2706_,
		_w2778_,
		_w2779_,
		_w2780_
	);
	LUT4 #(
		.INIT('h1b5f)
	) name1821 (
		\u0_spec_req_cs_reg[0]/NET0131 ,
		\u0_spec_req_cs_reg[1]/NET0131 ,
		\u0_u0_tms_reg[15]/P0001 ,
		\u0_u1_tms_reg[15]/P0001 ,
		_w2781_
	);
	LUT2 #(
		.INIT('h2)
	) name1822 (
		_w1013_,
		_w2781_,
		_w2782_
	);
	LUT4 #(
		.INIT('hef00)
	) name1823 (
		\u0_rf_we_reg/NET0131 ,
		_w2693_,
		_w2706_,
		_w2782_,
		_w2783_
	);
	LUT2 #(
		.INIT('hd)
	) name1824 (
		_w2780_,
		_w2783_,
		_w2784_
	);
	LUT3 #(
		.INIT('h2a)
	) name1825 (
		\u0_sp_tms_reg[1]/NET0131 ,
		wb_cyc_i_pad,
		wb_stb_i_pad,
		_w2785_
	);
	LUT2 #(
		.INIT('h4)
	) name1826 (
		\u0_rf_we_reg/NET0131 ,
		\u0_sp_tms_reg[1]/NET0131 ,
		_w2786_
	);
	LUT4 #(
		.INIT('h0b0f)
	) name1827 (
		_w2693_,
		_w2706_,
		_w2785_,
		_w2786_,
		_w2787_
	);
	LUT4 #(
		.INIT('h1b5f)
	) name1828 (
		\u0_spec_req_cs_reg[0]/NET0131 ,
		\u0_spec_req_cs_reg[1]/NET0131 ,
		\u0_u0_tms_reg[1]/P0001 ,
		\u0_u1_tms_reg[1]/P0001 ,
		_w2788_
	);
	LUT2 #(
		.INIT('h2)
	) name1829 (
		_w1013_,
		_w2788_,
		_w2789_
	);
	LUT4 #(
		.INIT('hef00)
	) name1830 (
		\u0_rf_we_reg/NET0131 ,
		_w2693_,
		_w2706_,
		_w2789_,
		_w2790_
	);
	LUT2 #(
		.INIT('hd)
	) name1831 (
		_w2787_,
		_w2790_,
		_w2791_
	);
	LUT3 #(
		.INIT('h2a)
	) name1832 (
		\u0_sp_tms_reg[21]/NET0131 ,
		wb_cyc_i_pad,
		wb_stb_i_pad,
		_w2792_
	);
	LUT2 #(
		.INIT('h4)
	) name1833 (
		\u0_rf_we_reg/NET0131 ,
		\u0_sp_tms_reg[21]/NET0131 ,
		_w2793_
	);
	LUT4 #(
		.INIT('h0b0f)
	) name1834 (
		_w2693_,
		_w2706_,
		_w2792_,
		_w2793_,
		_w2794_
	);
	LUT4 #(
		.INIT('h1b5f)
	) name1835 (
		\u0_spec_req_cs_reg[0]/NET0131 ,
		\u0_spec_req_cs_reg[1]/NET0131 ,
		\u0_u0_tms_reg[21]/P0001 ,
		\u0_u1_tms_reg[21]/P0001 ,
		_w2795_
	);
	LUT2 #(
		.INIT('h2)
	) name1836 (
		_w1013_,
		_w2795_,
		_w2796_
	);
	LUT4 #(
		.INIT('hef00)
	) name1837 (
		\u0_rf_we_reg/NET0131 ,
		_w2693_,
		_w2706_,
		_w2796_,
		_w2797_
	);
	LUT2 #(
		.INIT('hd)
	) name1838 (
		_w2794_,
		_w2797_,
		_w2798_
	);
	LUT3 #(
		.INIT('h2a)
	) name1839 (
		\u0_sp_tms_reg[20]/NET0131 ,
		wb_cyc_i_pad,
		wb_stb_i_pad,
		_w2799_
	);
	LUT2 #(
		.INIT('h4)
	) name1840 (
		\u0_rf_we_reg/NET0131 ,
		\u0_sp_tms_reg[20]/NET0131 ,
		_w2800_
	);
	LUT4 #(
		.INIT('h0b0f)
	) name1841 (
		_w2693_,
		_w2706_,
		_w2799_,
		_w2800_,
		_w2801_
	);
	LUT4 #(
		.INIT('h1b5f)
	) name1842 (
		\u0_spec_req_cs_reg[0]/NET0131 ,
		\u0_spec_req_cs_reg[1]/NET0131 ,
		\u0_u0_tms_reg[20]/P0001 ,
		\u0_u1_tms_reg[20]/P0001 ,
		_w2802_
	);
	LUT2 #(
		.INIT('h2)
	) name1843 (
		_w1013_,
		_w2802_,
		_w2803_
	);
	LUT4 #(
		.INIT('hef00)
	) name1844 (
		\u0_rf_we_reg/NET0131 ,
		_w2693_,
		_w2706_,
		_w2803_,
		_w2804_
	);
	LUT2 #(
		.INIT('hd)
	) name1845 (
		_w2801_,
		_w2804_,
		_w2805_
	);
	LUT3 #(
		.INIT('h2a)
	) name1846 (
		\u0_sp_tms_reg[22]/NET0131 ,
		wb_cyc_i_pad,
		wb_stb_i_pad,
		_w2806_
	);
	LUT2 #(
		.INIT('h4)
	) name1847 (
		\u0_rf_we_reg/NET0131 ,
		\u0_sp_tms_reg[22]/NET0131 ,
		_w2807_
	);
	LUT4 #(
		.INIT('h0b0f)
	) name1848 (
		_w2693_,
		_w2706_,
		_w2806_,
		_w2807_,
		_w2808_
	);
	LUT4 #(
		.INIT('h1b5f)
	) name1849 (
		\u0_spec_req_cs_reg[0]/NET0131 ,
		\u0_spec_req_cs_reg[1]/NET0131 ,
		\u0_u0_tms_reg[22]/P0001 ,
		\u0_u1_tms_reg[22]/P0001 ,
		_w2809_
	);
	LUT2 #(
		.INIT('h2)
	) name1850 (
		_w1013_,
		_w2809_,
		_w2810_
	);
	LUT4 #(
		.INIT('hef00)
	) name1851 (
		\u0_rf_we_reg/NET0131 ,
		_w2693_,
		_w2706_,
		_w2810_,
		_w2811_
	);
	LUT2 #(
		.INIT('hd)
	) name1852 (
		_w2808_,
		_w2811_,
		_w2812_
	);
	LUT3 #(
		.INIT('h2a)
	) name1853 (
		\u0_sp_tms_reg[23]/NET0131 ,
		wb_cyc_i_pad,
		wb_stb_i_pad,
		_w2813_
	);
	LUT2 #(
		.INIT('h4)
	) name1854 (
		\u0_rf_we_reg/NET0131 ,
		\u0_sp_tms_reg[23]/NET0131 ,
		_w2814_
	);
	LUT4 #(
		.INIT('h0b0f)
	) name1855 (
		_w2693_,
		_w2706_,
		_w2813_,
		_w2814_,
		_w2815_
	);
	LUT4 #(
		.INIT('h1b5f)
	) name1856 (
		\u0_spec_req_cs_reg[0]/NET0131 ,
		\u0_spec_req_cs_reg[1]/NET0131 ,
		\u0_u0_tms_reg[23]/P0001 ,
		\u0_u1_tms_reg[23]/P0001 ,
		_w2816_
	);
	LUT2 #(
		.INIT('h2)
	) name1857 (
		_w1013_,
		_w2816_,
		_w2817_
	);
	LUT4 #(
		.INIT('hef00)
	) name1858 (
		\u0_rf_we_reg/NET0131 ,
		_w2693_,
		_w2706_,
		_w2817_,
		_w2818_
	);
	LUT2 #(
		.INIT('hd)
	) name1859 (
		_w2815_,
		_w2818_,
		_w2819_
	);
	LUT3 #(
		.INIT('h2a)
	) name1860 (
		\u0_sp_tms_reg[24]/NET0131 ,
		wb_cyc_i_pad,
		wb_stb_i_pad,
		_w2820_
	);
	LUT2 #(
		.INIT('h4)
	) name1861 (
		\u0_rf_we_reg/NET0131 ,
		\u0_sp_tms_reg[24]/NET0131 ,
		_w2821_
	);
	LUT4 #(
		.INIT('h0b0f)
	) name1862 (
		_w2693_,
		_w2706_,
		_w2820_,
		_w2821_,
		_w2822_
	);
	LUT4 #(
		.INIT('h1b5f)
	) name1863 (
		\u0_spec_req_cs_reg[0]/NET0131 ,
		\u0_spec_req_cs_reg[1]/NET0131 ,
		\u0_u0_tms_reg[24]/P0001 ,
		\u0_u1_tms_reg[24]/P0001 ,
		_w2823_
	);
	LUT2 #(
		.INIT('h2)
	) name1864 (
		_w1013_,
		_w2823_,
		_w2824_
	);
	LUT4 #(
		.INIT('hef00)
	) name1865 (
		\u0_rf_we_reg/NET0131 ,
		_w2693_,
		_w2706_,
		_w2824_,
		_w2825_
	);
	LUT2 #(
		.INIT('hd)
	) name1866 (
		_w2822_,
		_w2825_,
		_w2826_
	);
	LUT3 #(
		.INIT('h2a)
	) name1867 (
		\u0_sp_tms_reg[25]/NET0131 ,
		wb_cyc_i_pad,
		wb_stb_i_pad,
		_w2827_
	);
	LUT2 #(
		.INIT('h4)
	) name1868 (
		\u0_rf_we_reg/NET0131 ,
		\u0_sp_tms_reg[25]/NET0131 ,
		_w2828_
	);
	LUT4 #(
		.INIT('h0b0f)
	) name1869 (
		_w2693_,
		_w2706_,
		_w2827_,
		_w2828_,
		_w2829_
	);
	LUT4 #(
		.INIT('h1b5f)
	) name1870 (
		\u0_spec_req_cs_reg[0]/NET0131 ,
		\u0_spec_req_cs_reg[1]/NET0131 ,
		\u0_u0_tms_reg[25]/P0001 ,
		\u0_u1_tms_reg[25]/P0001 ,
		_w2830_
	);
	LUT2 #(
		.INIT('h2)
	) name1871 (
		_w1013_,
		_w2830_,
		_w2831_
	);
	LUT4 #(
		.INIT('hef00)
	) name1872 (
		\u0_rf_we_reg/NET0131 ,
		_w2693_,
		_w2706_,
		_w2831_,
		_w2832_
	);
	LUT2 #(
		.INIT('hd)
	) name1873 (
		_w2829_,
		_w2832_,
		_w2833_
	);
	LUT3 #(
		.INIT('h2a)
	) name1874 (
		\u0_sp_tms_reg[26]/NET0131 ,
		wb_cyc_i_pad,
		wb_stb_i_pad,
		_w2834_
	);
	LUT2 #(
		.INIT('h4)
	) name1875 (
		\u0_rf_we_reg/NET0131 ,
		\u0_sp_tms_reg[26]/NET0131 ,
		_w2835_
	);
	LUT4 #(
		.INIT('h0b0f)
	) name1876 (
		_w2693_,
		_w2706_,
		_w2834_,
		_w2835_,
		_w2836_
	);
	LUT4 #(
		.INIT('h1b5f)
	) name1877 (
		\u0_spec_req_cs_reg[0]/NET0131 ,
		\u0_spec_req_cs_reg[1]/NET0131 ,
		\u0_u0_tms_reg[26]/P0001 ,
		\u0_u1_tms_reg[26]/P0001 ,
		_w2837_
	);
	LUT2 #(
		.INIT('h2)
	) name1878 (
		_w1013_,
		_w2837_,
		_w2838_
	);
	LUT4 #(
		.INIT('hef00)
	) name1879 (
		\u0_rf_we_reg/NET0131 ,
		_w2693_,
		_w2706_,
		_w2838_,
		_w2839_
	);
	LUT2 #(
		.INIT('hd)
	) name1880 (
		_w2836_,
		_w2839_,
		_w2840_
	);
	LUT3 #(
		.INIT('h2a)
	) name1881 (
		\u0_sp_tms_reg[27]/NET0131 ,
		wb_cyc_i_pad,
		wb_stb_i_pad,
		_w2841_
	);
	LUT2 #(
		.INIT('h4)
	) name1882 (
		\u0_rf_we_reg/NET0131 ,
		\u0_sp_tms_reg[27]/NET0131 ,
		_w2842_
	);
	LUT4 #(
		.INIT('h0b0f)
	) name1883 (
		_w2693_,
		_w2706_,
		_w2841_,
		_w2842_,
		_w2843_
	);
	LUT4 #(
		.INIT('h1b5f)
	) name1884 (
		\u0_spec_req_cs_reg[0]/NET0131 ,
		\u0_spec_req_cs_reg[1]/NET0131 ,
		\u0_u0_tms_reg[27]/P0001 ,
		\u0_u1_tms_reg[27]/P0001 ,
		_w2844_
	);
	LUT2 #(
		.INIT('h2)
	) name1885 (
		_w1013_,
		_w2844_,
		_w2845_
	);
	LUT4 #(
		.INIT('hef00)
	) name1886 (
		\u0_rf_we_reg/NET0131 ,
		_w2693_,
		_w2706_,
		_w2845_,
		_w2846_
	);
	LUT2 #(
		.INIT('hd)
	) name1887 (
		_w2843_,
		_w2846_,
		_w2847_
	);
	LUT3 #(
		.INIT('h2a)
	) name1888 (
		\u0_sp_tms_reg[2]/NET0131 ,
		wb_cyc_i_pad,
		wb_stb_i_pad,
		_w2848_
	);
	LUT2 #(
		.INIT('h4)
	) name1889 (
		\u0_rf_we_reg/NET0131 ,
		\u0_sp_tms_reg[2]/NET0131 ,
		_w2849_
	);
	LUT4 #(
		.INIT('h0b0f)
	) name1890 (
		_w2693_,
		_w2706_,
		_w2848_,
		_w2849_,
		_w2850_
	);
	LUT4 #(
		.INIT('h1b5f)
	) name1891 (
		\u0_spec_req_cs_reg[0]/NET0131 ,
		\u0_spec_req_cs_reg[1]/NET0131 ,
		\u0_u0_tms_reg[2]/P0001 ,
		\u0_u1_tms_reg[2]/P0001 ,
		_w2851_
	);
	LUT2 #(
		.INIT('h2)
	) name1892 (
		_w1013_,
		_w2851_,
		_w2852_
	);
	LUT4 #(
		.INIT('hef00)
	) name1893 (
		\u0_rf_we_reg/NET0131 ,
		_w2693_,
		_w2706_,
		_w2852_,
		_w2853_
	);
	LUT2 #(
		.INIT('hd)
	) name1894 (
		_w2850_,
		_w2853_,
		_w2854_
	);
	LUT3 #(
		.INIT('h2a)
	) name1895 (
		\u0_sp_tms_reg[3]/NET0131 ,
		wb_cyc_i_pad,
		wb_stb_i_pad,
		_w2855_
	);
	LUT2 #(
		.INIT('h4)
	) name1896 (
		\u0_rf_we_reg/NET0131 ,
		\u0_sp_tms_reg[3]/NET0131 ,
		_w2856_
	);
	LUT4 #(
		.INIT('h0b0f)
	) name1897 (
		_w2693_,
		_w2706_,
		_w2855_,
		_w2856_,
		_w2857_
	);
	LUT4 #(
		.INIT('h1b5f)
	) name1898 (
		\u0_spec_req_cs_reg[0]/NET0131 ,
		\u0_spec_req_cs_reg[1]/NET0131 ,
		\u0_u0_tms_reg[3]/P0001 ,
		\u0_u1_tms_reg[3]/P0001 ,
		_w2858_
	);
	LUT2 #(
		.INIT('h2)
	) name1899 (
		_w1013_,
		_w2858_,
		_w2859_
	);
	LUT4 #(
		.INIT('hef00)
	) name1900 (
		\u0_rf_we_reg/NET0131 ,
		_w2693_,
		_w2706_,
		_w2859_,
		_w2860_
	);
	LUT2 #(
		.INIT('hd)
	) name1901 (
		_w2857_,
		_w2860_,
		_w2861_
	);
	LUT3 #(
		.INIT('h2a)
	) name1902 (
		\u0_sp_tms_reg[4]/NET0131 ,
		wb_cyc_i_pad,
		wb_stb_i_pad,
		_w2862_
	);
	LUT2 #(
		.INIT('h4)
	) name1903 (
		\u0_rf_we_reg/NET0131 ,
		\u0_sp_tms_reg[4]/NET0131 ,
		_w2863_
	);
	LUT4 #(
		.INIT('h0b0f)
	) name1904 (
		_w2693_,
		_w2706_,
		_w2862_,
		_w2863_,
		_w2864_
	);
	LUT4 #(
		.INIT('h1b5f)
	) name1905 (
		\u0_spec_req_cs_reg[0]/NET0131 ,
		\u0_spec_req_cs_reg[1]/NET0131 ,
		\u0_u0_tms_reg[4]/P0001 ,
		\u0_u1_tms_reg[4]/P0001 ,
		_w2865_
	);
	LUT2 #(
		.INIT('h2)
	) name1906 (
		_w1013_,
		_w2865_,
		_w2866_
	);
	LUT4 #(
		.INIT('hef00)
	) name1907 (
		\u0_rf_we_reg/NET0131 ,
		_w2693_,
		_w2706_,
		_w2866_,
		_w2867_
	);
	LUT2 #(
		.INIT('hd)
	) name1908 (
		_w2864_,
		_w2867_,
		_w2868_
	);
	LUT3 #(
		.INIT('h2a)
	) name1909 (
		\u0_sp_tms_reg[5]/NET0131 ,
		wb_cyc_i_pad,
		wb_stb_i_pad,
		_w2869_
	);
	LUT2 #(
		.INIT('h4)
	) name1910 (
		\u0_rf_we_reg/NET0131 ,
		\u0_sp_tms_reg[5]/NET0131 ,
		_w2870_
	);
	LUT4 #(
		.INIT('h0b0f)
	) name1911 (
		_w2693_,
		_w2706_,
		_w2869_,
		_w2870_,
		_w2871_
	);
	LUT4 #(
		.INIT('h1b5f)
	) name1912 (
		\u0_spec_req_cs_reg[0]/NET0131 ,
		\u0_spec_req_cs_reg[1]/NET0131 ,
		\u0_u0_tms_reg[5]/P0001 ,
		\u0_u1_tms_reg[5]/P0001 ,
		_w2872_
	);
	LUT2 #(
		.INIT('h2)
	) name1913 (
		_w1013_,
		_w2872_,
		_w2873_
	);
	LUT4 #(
		.INIT('hef00)
	) name1914 (
		\u0_rf_we_reg/NET0131 ,
		_w2693_,
		_w2706_,
		_w2873_,
		_w2874_
	);
	LUT2 #(
		.INIT('hd)
	) name1915 (
		_w2871_,
		_w2874_,
		_w2875_
	);
	LUT3 #(
		.INIT('h2a)
	) name1916 (
		\u0_sp_tms_reg[7]/NET0131 ,
		wb_cyc_i_pad,
		wb_stb_i_pad,
		_w2876_
	);
	LUT2 #(
		.INIT('h4)
	) name1917 (
		\u0_rf_we_reg/NET0131 ,
		\u0_sp_tms_reg[7]/NET0131 ,
		_w2877_
	);
	LUT4 #(
		.INIT('h0b0f)
	) name1918 (
		_w2693_,
		_w2706_,
		_w2876_,
		_w2877_,
		_w2878_
	);
	LUT4 #(
		.INIT('h1b5f)
	) name1919 (
		\u0_spec_req_cs_reg[0]/NET0131 ,
		\u0_spec_req_cs_reg[1]/NET0131 ,
		\u0_u0_tms_reg[7]/P0001 ,
		\u0_u1_tms_reg[7]/P0001 ,
		_w2879_
	);
	LUT2 #(
		.INIT('h2)
	) name1920 (
		_w1013_,
		_w2879_,
		_w2880_
	);
	LUT4 #(
		.INIT('hef00)
	) name1921 (
		\u0_rf_we_reg/NET0131 ,
		_w2693_,
		_w2706_,
		_w2880_,
		_w2881_
	);
	LUT2 #(
		.INIT('hd)
	) name1922 (
		_w2878_,
		_w2881_,
		_w2882_
	);
	LUT3 #(
		.INIT('h2a)
	) name1923 (
		\u0_sp_tms_reg[6]/NET0131 ,
		wb_cyc_i_pad,
		wb_stb_i_pad,
		_w2883_
	);
	LUT2 #(
		.INIT('h4)
	) name1924 (
		\u0_rf_we_reg/NET0131 ,
		\u0_sp_tms_reg[6]/NET0131 ,
		_w2884_
	);
	LUT4 #(
		.INIT('h0b0f)
	) name1925 (
		_w2693_,
		_w2706_,
		_w2883_,
		_w2884_,
		_w2885_
	);
	LUT4 #(
		.INIT('h1b5f)
	) name1926 (
		\u0_spec_req_cs_reg[0]/NET0131 ,
		\u0_spec_req_cs_reg[1]/NET0131 ,
		\u0_u0_tms_reg[6]/P0001 ,
		\u0_u1_tms_reg[6]/P0001 ,
		_w2886_
	);
	LUT2 #(
		.INIT('h2)
	) name1927 (
		_w1013_,
		_w2886_,
		_w2887_
	);
	LUT4 #(
		.INIT('hef00)
	) name1928 (
		\u0_rf_we_reg/NET0131 ,
		_w2693_,
		_w2706_,
		_w2887_,
		_w2888_
	);
	LUT2 #(
		.INIT('hd)
	) name1929 (
		_w2885_,
		_w2888_,
		_w2889_
	);
	LUT3 #(
		.INIT('h2a)
	) name1930 (
		\u0_sp_tms_reg[8]/NET0131 ,
		wb_cyc_i_pad,
		wb_stb_i_pad,
		_w2890_
	);
	LUT2 #(
		.INIT('h4)
	) name1931 (
		\u0_rf_we_reg/NET0131 ,
		\u0_sp_tms_reg[8]/NET0131 ,
		_w2891_
	);
	LUT4 #(
		.INIT('h0b0f)
	) name1932 (
		_w2693_,
		_w2706_,
		_w2890_,
		_w2891_,
		_w2892_
	);
	LUT4 #(
		.INIT('h1b5f)
	) name1933 (
		\u0_spec_req_cs_reg[0]/NET0131 ,
		\u0_spec_req_cs_reg[1]/NET0131 ,
		\u0_u0_tms_reg[8]/P0001 ,
		\u0_u1_tms_reg[8]/P0001 ,
		_w2893_
	);
	LUT2 #(
		.INIT('h2)
	) name1934 (
		_w1013_,
		_w2893_,
		_w2894_
	);
	LUT4 #(
		.INIT('hef00)
	) name1935 (
		\u0_rf_we_reg/NET0131 ,
		_w2693_,
		_w2706_,
		_w2894_,
		_w2895_
	);
	LUT2 #(
		.INIT('hd)
	) name1936 (
		_w2892_,
		_w2895_,
		_w2896_
	);
	LUT3 #(
		.INIT('h2a)
	) name1937 (
		\u0_sp_tms_reg[9]/NET0131 ,
		wb_cyc_i_pad,
		wb_stb_i_pad,
		_w2897_
	);
	LUT2 #(
		.INIT('h4)
	) name1938 (
		\u0_rf_we_reg/NET0131 ,
		\u0_sp_tms_reg[9]/NET0131 ,
		_w2898_
	);
	LUT4 #(
		.INIT('h0b0f)
	) name1939 (
		_w2693_,
		_w2706_,
		_w2897_,
		_w2898_,
		_w2899_
	);
	LUT4 #(
		.INIT('h1b5f)
	) name1940 (
		\u0_spec_req_cs_reg[0]/NET0131 ,
		\u0_spec_req_cs_reg[1]/NET0131 ,
		\u0_u0_tms_reg[9]/P0001 ,
		\u0_u1_tms_reg[9]/P0001 ,
		_w2900_
	);
	LUT2 #(
		.INIT('h2)
	) name1941 (
		_w1013_,
		_w2900_,
		_w2901_
	);
	LUT4 #(
		.INIT('hef00)
	) name1942 (
		\u0_rf_we_reg/NET0131 ,
		_w2693_,
		_w2706_,
		_w2901_,
		_w2902_
	);
	LUT2 #(
		.INIT('hd)
	) name1943 (
		_w2899_,
		_w2902_,
		_w2903_
	);
	LUT3 #(
		.INIT('h2a)
	) name1944 (
		\u0_tms_reg[10]/NET0131 ,
		wb_cyc_i_pad,
		wb_stb_i_pad,
		_w2904_
	);
	LUT2 #(
		.INIT('h4)
	) name1945 (
		\u0_rf_we_reg/NET0131 ,
		\u0_tms_reg[10]/NET0131 ,
		_w2905_
	);
	LUT4 #(
		.INIT('h0b0f)
	) name1946 (
		_w2693_,
		_w2706_,
		_w2904_,
		_w2905_,
		_w2906_
	);
	LUT4 #(
		.INIT('hc44c)
	) name1947 (
		\u0_csc_mask_r_reg[2]/NET0131 ,
		\u0_u0_csc_reg[0]/NET0131 ,
		\u0_u0_csc_reg[18]/P0001 ,
		\wb_addr_i[23]_pad ,
		_w2907_
	);
	LUT3 #(
		.INIT('h28)
	) name1948 (
		\u0_csc_mask_r_reg[4]/NET0131 ,
		\u0_u0_csc_reg[20]/P0001 ,
		\wb_addr_i[25]_pad ,
		_w2908_
	);
	LUT3 #(
		.INIT('h28)
	) name1949 (
		\u0_csc_mask_r_reg[6]/NET0131 ,
		\u0_u0_csc_reg[22]/P0001 ,
		\wb_addr_i[27]_pad ,
		_w2909_
	);
	LUT3 #(
		.INIT('h28)
	) name1950 (
		\u0_csc_mask_r_reg[7]/NET0131 ,
		\u0_u0_csc_reg[23]/P0001 ,
		\wb_addr_i[28]_pad ,
		_w2910_
	);
	LUT3 #(
		.INIT('h28)
	) name1951 (
		\u0_csc_mask_r_reg[1]/NET0131 ,
		\u0_u0_csc_reg[17]/P0001 ,
		\wb_addr_i[22]_pad ,
		_w2911_
	);
	LUT4 #(
		.INIT('h0001)
	) name1952 (
		_w2908_,
		_w2909_,
		_w2910_,
		_w2911_,
		_w2912_
	);
	LUT2 #(
		.INIT('h8)
	) name1953 (
		\u0_u0_csc_reg[8]/P0001 ,
		wb_we_i_pad,
		_w2913_
	);
	LUT3 #(
		.INIT('h28)
	) name1954 (
		\u0_csc_mask_r_reg[5]/NET0131 ,
		\u0_u0_csc_reg[21]/P0001 ,
		\wb_addr_i[26]_pad ,
		_w2914_
	);
	LUT3 #(
		.INIT('h28)
	) name1955 (
		\u0_csc_mask_r_reg[0]/NET0131 ,
		\u0_u0_csc_reg[16]/P0001 ,
		\wb_addr_i[21]_pad ,
		_w2915_
	);
	LUT3 #(
		.INIT('h28)
	) name1956 (
		\u0_csc_mask_r_reg[3]/NET0131 ,
		\u0_u0_csc_reg[19]/P0001 ,
		\wb_addr_i[24]_pad ,
		_w2916_
	);
	LUT4 #(
		.INIT('h0001)
	) name1957 (
		_w2913_,
		_w2914_,
		_w2915_,
		_w2916_,
		_w2917_
	);
	LUT3 #(
		.INIT('h80)
	) name1958 (
		_w2907_,
		_w2912_,
		_w2917_,
		_w2918_
	);
	LUT4 #(
		.INIT('hc44c)
	) name1959 (
		\u0_csc_mask_r_reg[1]/NET0131 ,
		\u0_u1_csc_reg[0]/NET0131 ,
		\u0_u1_csc_reg[17]/P0001 ,
		\wb_addr_i[22]_pad ,
		_w2919_
	);
	LUT3 #(
		.INIT('h28)
	) name1960 (
		\u0_csc_mask_r_reg[5]/NET0131 ,
		\u0_u1_csc_reg[21]/P0001 ,
		\wb_addr_i[26]_pad ,
		_w2920_
	);
	LUT3 #(
		.INIT('h28)
	) name1961 (
		\u0_csc_mask_r_reg[6]/NET0131 ,
		\u0_u1_csc_reg[22]/P0001 ,
		\wb_addr_i[27]_pad ,
		_w2921_
	);
	LUT3 #(
		.INIT('h28)
	) name1962 (
		\u0_csc_mask_r_reg[3]/NET0131 ,
		\u0_u1_csc_reg[19]/P0001 ,
		\wb_addr_i[24]_pad ,
		_w2922_
	);
	LUT3 #(
		.INIT('h28)
	) name1963 (
		\u0_csc_mask_r_reg[0]/NET0131 ,
		\u0_u1_csc_reg[16]/P0001 ,
		\wb_addr_i[21]_pad ,
		_w2923_
	);
	LUT4 #(
		.INIT('h0001)
	) name1964 (
		_w2920_,
		_w2921_,
		_w2922_,
		_w2923_,
		_w2924_
	);
	LUT2 #(
		.INIT('h8)
	) name1965 (
		\u0_u1_csc_reg[8]/P0001 ,
		wb_we_i_pad,
		_w2925_
	);
	LUT3 #(
		.INIT('h28)
	) name1966 (
		\u0_csc_mask_r_reg[4]/NET0131 ,
		\u0_u1_csc_reg[20]/P0001 ,
		\wb_addr_i[25]_pad ,
		_w2926_
	);
	LUT3 #(
		.INIT('h28)
	) name1967 (
		\u0_csc_mask_r_reg[2]/NET0131 ,
		\u0_u1_csc_reg[18]/P0001 ,
		\wb_addr_i[23]_pad ,
		_w2927_
	);
	LUT3 #(
		.INIT('h28)
	) name1968 (
		\u0_csc_mask_r_reg[7]/NET0131 ,
		\u0_u1_csc_reg[23]/P0001 ,
		\wb_addr_i[28]_pad ,
		_w2928_
	);
	LUT4 #(
		.INIT('h0001)
	) name1969 (
		_w2925_,
		_w2926_,
		_w2927_,
		_w2928_,
		_w2929_
	);
	LUT3 #(
		.INIT('h80)
	) name1970 (
		_w2919_,
		_w2924_,
		_w2929_,
		_w2930_
	);
	LUT3 #(
		.INIT('h4c)
	) name1971 (
		\u0_u0_csc_reg[8]/P0001 ,
		\u0_u0_tms_reg[10]/P0001 ,
		wb_we_i_pad,
		_w2931_
	);
	LUT4 #(
		.INIT('h0100)
	) name1972 (
		_w2914_,
		_w2915_,
		_w2916_,
		_w2931_,
		_w2932_
	);
	LUT3 #(
		.INIT('h80)
	) name1973 (
		_w2907_,
		_w2912_,
		_w2932_,
		_w2933_
	);
	LUT4 #(
		.INIT('h00df)
	) name1974 (
		\u0_u1_tms_reg[10]/P0001 ,
		_w2918_,
		_w2930_,
		_w2933_,
		_w2934_
	);
	LUT2 #(
		.INIT('h2)
	) name1975 (
		_w1013_,
		_w2934_,
		_w2935_
	);
	LUT4 #(
		.INIT('hef00)
	) name1976 (
		\u0_rf_we_reg/NET0131 ,
		_w2693_,
		_w2706_,
		_w2935_,
		_w2936_
	);
	LUT2 #(
		.INIT('hd)
	) name1977 (
		_w2906_,
		_w2936_,
		_w2937_
	);
	LUT3 #(
		.INIT('h2a)
	) name1978 (
		\u0_tms_reg[11]/NET0131 ,
		wb_cyc_i_pad,
		wb_stb_i_pad,
		_w2938_
	);
	LUT2 #(
		.INIT('h4)
	) name1979 (
		\u0_rf_we_reg/NET0131 ,
		\u0_tms_reg[11]/NET0131 ,
		_w2939_
	);
	LUT4 #(
		.INIT('h0b0f)
	) name1980 (
		_w2693_,
		_w2706_,
		_w2938_,
		_w2939_,
		_w2940_
	);
	LUT3 #(
		.INIT('h4c)
	) name1981 (
		\u0_u0_csc_reg[8]/P0001 ,
		\u0_u0_tms_reg[11]/P0001 ,
		wb_we_i_pad,
		_w2941_
	);
	LUT4 #(
		.INIT('h0100)
	) name1982 (
		_w2914_,
		_w2915_,
		_w2916_,
		_w2941_,
		_w2942_
	);
	LUT3 #(
		.INIT('h80)
	) name1983 (
		_w2907_,
		_w2912_,
		_w2942_,
		_w2943_
	);
	LUT4 #(
		.INIT('h00df)
	) name1984 (
		\u0_u1_tms_reg[11]/P0001 ,
		_w2918_,
		_w2930_,
		_w2943_,
		_w2944_
	);
	LUT2 #(
		.INIT('h2)
	) name1985 (
		_w1013_,
		_w2944_,
		_w2945_
	);
	LUT4 #(
		.INIT('hef00)
	) name1986 (
		\u0_rf_we_reg/NET0131 ,
		_w2693_,
		_w2706_,
		_w2945_,
		_w2946_
	);
	LUT2 #(
		.INIT('hd)
	) name1987 (
		_w2940_,
		_w2946_,
		_w2947_
	);
	LUT3 #(
		.INIT('h2a)
	) name1988 (
		\u0_tms_reg[12]/NET0131 ,
		wb_cyc_i_pad,
		wb_stb_i_pad,
		_w2948_
	);
	LUT2 #(
		.INIT('h4)
	) name1989 (
		\u0_rf_we_reg/NET0131 ,
		\u0_tms_reg[12]/NET0131 ,
		_w2949_
	);
	LUT4 #(
		.INIT('h0b0f)
	) name1990 (
		_w2693_,
		_w2706_,
		_w2948_,
		_w2949_,
		_w2950_
	);
	LUT3 #(
		.INIT('h4c)
	) name1991 (
		\u0_u0_csc_reg[8]/P0001 ,
		\u0_u0_tms_reg[12]/P0001 ,
		wb_we_i_pad,
		_w2951_
	);
	LUT4 #(
		.INIT('h0100)
	) name1992 (
		_w2914_,
		_w2915_,
		_w2916_,
		_w2951_,
		_w2952_
	);
	LUT3 #(
		.INIT('h80)
	) name1993 (
		_w2907_,
		_w2912_,
		_w2952_,
		_w2953_
	);
	LUT4 #(
		.INIT('h00df)
	) name1994 (
		\u0_u1_tms_reg[12]/P0001 ,
		_w2918_,
		_w2930_,
		_w2953_,
		_w2954_
	);
	LUT2 #(
		.INIT('h2)
	) name1995 (
		_w1013_,
		_w2954_,
		_w2955_
	);
	LUT4 #(
		.INIT('hef00)
	) name1996 (
		\u0_rf_we_reg/NET0131 ,
		_w2693_,
		_w2706_,
		_w2955_,
		_w2956_
	);
	LUT2 #(
		.INIT('hd)
	) name1997 (
		_w2950_,
		_w2956_,
		_w2957_
	);
	LUT3 #(
		.INIT('h2a)
	) name1998 (
		\u0_tms_reg[13]/NET0131 ,
		wb_cyc_i_pad,
		wb_stb_i_pad,
		_w2958_
	);
	LUT2 #(
		.INIT('h4)
	) name1999 (
		\u0_rf_we_reg/NET0131 ,
		\u0_tms_reg[13]/NET0131 ,
		_w2959_
	);
	LUT4 #(
		.INIT('h0b0f)
	) name2000 (
		_w2693_,
		_w2706_,
		_w2958_,
		_w2959_,
		_w2960_
	);
	LUT3 #(
		.INIT('h4c)
	) name2001 (
		\u0_u0_csc_reg[8]/P0001 ,
		\u0_u0_tms_reg[13]/P0001 ,
		wb_we_i_pad,
		_w2961_
	);
	LUT4 #(
		.INIT('h0100)
	) name2002 (
		_w2914_,
		_w2915_,
		_w2916_,
		_w2961_,
		_w2962_
	);
	LUT3 #(
		.INIT('h80)
	) name2003 (
		_w2907_,
		_w2912_,
		_w2962_,
		_w2963_
	);
	LUT4 #(
		.INIT('h00df)
	) name2004 (
		\u0_u1_tms_reg[13]/P0001 ,
		_w2918_,
		_w2930_,
		_w2963_,
		_w2964_
	);
	LUT2 #(
		.INIT('h2)
	) name2005 (
		_w1013_,
		_w2964_,
		_w2965_
	);
	LUT4 #(
		.INIT('hef00)
	) name2006 (
		\u0_rf_we_reg/NET0131 ,
		_w2693_,
		_w2706_,
		_w2965_,
		_w2966_
	);
	LUT2 #(
		.INIT('hd)
	) name2007 (
		_w2960_,
		_w2966_,
		_w2967_
	);
	LUT3 #(
		.INIT('h2a)
	) name2008 (
		\u0_tms_reg[0]/NET0131 ,
		wb_cyc_i_pad,
		wb_stb_i_pad,
		_w2968_
	);
	LUT2 #(
		.INIT('h4)
	) name2009 (
		\u0_rf_we_reg/NET0131 ,
		\u0_tms_reg[0]/NET0131 ,
		_w2969_
	);
	LUT4 #(
		.INIT('h0b0f)
	) name2010 (
		_w2693_,
		_w2706_,
		_w2968_,
		_w2969_,
		_w2970_
	);
	LUT3 #(
		.INIT('h4c)
	) name2011 (
		\u0_u0_csc_reg[8]/P0001 ,
		\u0_u0_tms_reg[0]/P0001 ,
		wb_we_i_pad,
		_w2971_
	);
	LUT4 #(
		.INIT('h0100)
	) name2012 (
		_w2914_,
		_w2915_,
		_w2916_,
		_w2971_,
		_w2972_
	);
	LUT3 #(
		.INIT('h80)
	) name2013 (
		_w2907_,
		_w2912_,
		_w2972_,
		_w2973_
	);
	LUT4 #(
		.INIT('h00df)
	) name2014 (
		\u0_u1_tms_reg[0]/P0001 ,
		_w2918_,
		_w2930_,
		_w2973_,
		_w2974_
	);
	LUT2 #(
		.INIT('h2)
	) name2015 (
		_w1013_,
		_w2974_,
		_w2975_
	);
	LUT4 #(
		.INIT('hef00)
	) name2016 (
		\u0_rf_we_reg/NET0131 ,
		_w2693_,
		_w2706_,
		_w2975_,
		_w2976_
	);
	LUT2 #(
		.INIT('hd)
	) name2017 (
		_w2970_,
		_w2976_,
		_w2977_
	);
	LUT3 #(
		.INIT('h2a)
	) name2018 (
		\u0_tms_reg[14]/NET0131 ,
		wb_cyc_i_pad,
		wb_stb_i_pad,
		_w2978_
	);
	LUT2 #(
		.INIT('h4)
	) name2019 (
		\u0_rf_we_reg/NET0131 ,
		\u0_tms_reg[14]/NET0131 ,
		_w2979_
	);
	LUT4 #(
		.INIT('h0b0f)
	) name2020 (
		_w2693_,
		_w2706_,
		_w2978_,
		_w2979_,
		_w2980_
	);
	LUT3 #(
		.INIT('h4c)
	) name2021 (
		\u0_u0_csc_reg[8]/P0001 ,
		\u0_u0_tms_reg[14]/P0001 ,
		wb_we_i_pad,
		_w2981_
	);
	LUT4 #(
		.INIT('h0100)
	) name2022 (
		_w2914_,
		_w2915_,
		_w2916_,
		_w2981_,
		_w2982_
	);
	LUT3 #(
		.INIT('h80)
	) name2023 (
		_w2907_,
		_w2912_,
		_w2982_,
		_w2983_
	);
	LUT4 #(
		.INIT('h00df)
	) name2024 (
		\u0_u1_tms_reg[14]/P0001 ,
		_w2918_,
		_w2930_,
		_w2983_,
		_w2984_
	);
	LUT2 #(
		.INIT('h2)
	) name2025 (
		_w1013_,
		_w2984_,
		_w2985_
	);
	LUT4 #(
		.INIT('hef00)
	) name2026 (
		\u0_rf_we_reg/NET0131 ,
		_w2693_,
		_w2706_,
		_w2985_,
		_w2986_
	);
	LUT2 #(
		.INIT('hd)
	) name2027 (
		_w2980_,
		_w2986_,
		_w2987_
	);
	LUT3 #(
		.INIT('h2a)
	) name2028 (
		\u0_tms_reg[15]/NET0131 ,
		wb_cyc_i_pad,
		wb_stb_i_pad,
		_w2988_
	);
	LUT2 #(
		.INIT('h4)
	) name2029 (
		\u0_rf_we_reg/NET0131 ,
		\u0_tms_reg[15]/NET0131 ,
		_w2989_
	);
	LUT4 #(
		.INIT('h0b0f)
	) name2030 (
		_w2693_,
		_w2706_,
		_w2988_,
		_w2989_,
		_w2990_
	);
	LUT3 #(
		.INIT('h4c)
	) name2031 (
		\u0_u0_csc_reg[8]/P0001 ,
		\u0_u0_tms_reg[15]/P0001 ,
		wb_we_i_pad,
		_w2991_
	);
	LUT4 #(
		.INIT('h0100)
	) name2032 (
		_w2914_,
		_w2915_,
		_w2916_,
		_w2991_,
		_w2992_
	);
	LUT3 #(
		.INIT('h80)
	) name2033 (
		_w2907_,
		_w2912_,
		_w2992_,
		_w2993_
	);
	LUT4 #(
		.INIT('h00df)
	) name2034 (
		\u0_u1_tms_reg[15]/P0001 ,
		_w2918_,
		_w2930_,
		_w2993_,
		_w2994_
	);
	LUT2 #(
		.INIT('h2)
	) name2035 (
		_w1013_,
		_w2994_,
		_w2995_
	);
	LUT4 #(
		.INIT('hef00)
	) name2036 (
		\u0_rf_we_reg/NET0131 ,
		_w2693_,
		_w2706_,
		_w2995_,
		_w2996_
	);
	LUT2 #(
		.INIT('hd)
	) name2037 (
		_w2990_,
		_w2996_,
		_w2997_
	);
	LUT3 #(
		.INIT('h2a)
	) name2038 (
		\u0_tms_reg[16]/NET0131 ,
		wb_cyc_i_pad,
		wb_stb_i_pad,
		_w2998_
	);
	LUT2 #(
		.INIT('h4)
	) name2039 (
		\u0_rf_we_reg/NET0131 ,
		\u0_tms_reg[16]/NET0131 ,
		_w2999_
	);
	LUT4 #(
		.INIT('h0b0f)
	) name2040 (
		_w2693_,
		_w2706_,
		_w2998_,
		_w2999_,
		_w3000_
	);
	LUT3 #(
		.INIT('h4c)
	) name2041 (
		\u0_u0_csc_reg[8]/P0001 ,
		\u0_u0_tms_reg[16]/P0001 ,
		wb_we_i_pad,
		_w3001_
	);
	LUT4 #(
		.INIT('h0100)
	) name2042 (
		_w2914_,
		_w2915_,
		_w2916_,
		_w3001_,
		_w3002_
	);
	LUT3 #(
		.INIT('h80)
	) name2043 (
		_w2907_,
		_w2912_,
		_w3002_,
		_w3003_
	);
	LUT4 #(
		.INIT('h00df)
	) name2044 (
		\u0_u1_tms_reg[16]/P0001 ,
		_w2918_,
		_w2930_,
		_w3003_,
		_w3004_
	);
	LUT2 #(
		.INIT('h2)
	) name2045 (
		_w1013_,
		_w3004_,
		_w3005_
	);
	LUT4 #(
		.INIT('hef00)
	) name2046 (
		\u0_rf_we_reg/NET0131 ,
		_w2693_,
		_w2706_,
		_w3005_,
		_w3006_
	);
	LUT2 #(
		.INIT('hd)
	) name2047 (
		_w3000_,
		_w3006_,
		_w3007_
	);
	LUT3 #(
		.INIT('h2a)
	) name2048 (
		\u0_tms_reg[17]/NET0131 ,
		wb_cyc_i_pad,
		wb_stb_i_pad,
		_w3008_
	);
	LUT2 #(
		.INIT('h4)
	) name2049 (
		\u0_rf_we_reg/NET0131 ,
		\u0_tms_reg[17]/NET0131 ,
		_w3009_
	);
	LUT4 #(
		.INIT('h0b0f)
	) name2050 (
		_w2693_,
		_w2706_,
		_w3008_,
		_w3009_,
		_w3010_
	);
	LUT3 #(
		.INIT('h4c)
	) name2051 (
		\u0_u0_csc_reg[8]/P0001 ,
		\u0_u0_tms_reg[17]/P0001 ,
		wb_we_i_pad,
		_w3011_
	);
	LUT4 #(
		.INIT('h0100)
	) name2052 (
		_w2914_,
		_w2915_,
		_w2916_,
		_w3011_,
		_w3012_
	);
	LUT3 #(
		.INIT('h80)
	) name2053 (
		_w2907_,
		_w2912_,
		_w3012_,
		_w3013_
	);
	LUT4 #(
		.INIT('h00df)
	) name2054 (
		\u0_u1_tms_reg[17]/P0001 ,
		_w2918_,
		_w2930_,
		_w3013_,
		_w3014_
	);
	LUT2 #(
		.INIT('h2)
	) name2055 (
		_w1013_,
		_w3014_,
		_w3015_
	);
	LUT4 #(
		.INIT('hef00)
	) name2056 (
		\u0_rf_we_reg/NET0131 ,
		_w2693_,
		_w2706_,
		_w3015_,
		_w3016_
	);
	LUT2 #(
		.INIT('hd)
	) name2057 (
		_w3010_,
		_w3016_,
		_w3017_
	);
	LUT3 #(
		.INIT('h2a)
	) name2058 (
		\u0_tms_reg[18]/NET0131 ,
		wb_cyc_i_pad,
		wb_stb_i_pad,
		_w3018_
	);
	LUT2 #(
		.INIT('h4)
	) name2059 (
		\u0_rf_we_reg/NET0131 ,
		\u0_tms_reg[18]/NET0131 ,
		_w3019_
	);
	LUT4 #(
		.INIT('h0b0f)
	) name2060 (
		_w2693_,
		_w2706_,
		_w3018_,
		_w3019_,
		_w3020_
	);
	LUT3 #(
		.INIT('h4c)
	) name2061 (
		\u0_u0_csc_reg[8]/P0001 ,
		\u0_u0_tms_reg[18]/P0001 ,
		wb_we_i_pad,
		_w3021_
	);
	LUT4 #(
		.INIT('h0100)
	) name2062 (
		_w2914_,
		_w2915_,
		_w2916_,
		_w3021_,
		_w3022_
	);
	LUT3 #(
		.INIT('h80)
	) name2063 (
		_w2907_,
		_w2912_,
		_w3022_,
		_w3023_
	);
	LUT4 #(
		.INIT('h00df)
	) name2064 (
		\u0_u1_tms_reg[18]/P0001 ,
		_w2918_,
		_w2930_,
		_w3023_,
		_w3024_
	);
	LUT2 #(
		.INIT('h2)
	) name2065 (
		_w1013_,
		_w3024_,
		_w3025_
	);
	LUT4 #(
		.INIT('hef00)
	) name2066 (
		\u0_rf_we_reg/NET0131 ,
		_w2693_,
		_w2706_,
		_w3025_,
		_w3026_
	);
	LUT2 #(
		.INIT('hd)
	) name2067 (
		_w3020_,
		_w3026_,
		_w3027_
	);
	LUT3 #(
		.INIT('h2a)
	) name2068 (
		\u0_tms_reg[19]/NET0131 ,
		wb_cyc_i_pad,
		wb_stb_i_pad,
		_w3028_
	);
	LUT2 #(
		.INIT('h4)
	) name2069 (
		\u0_rf_we_reg/NET0131 ,
		\u0_tms_reg[19]/NET0131 ,
		_w3029_
	);
	LUT4 #(
		.INIT('h0b0f)
	) name2070 (
		_w2693_,
		_w2706_,
		_w3028_,
		_w3029_,
		_w3030_
	);
	LUT3 #(
		.INIT('h4c)
	) name2071 (
		\u0_u0_csc_reg[8]/P0001 ,
		\u0_u0_tms_reg[19]/P0001 ,
		wb_we_i_pad,
		_w3031_
	);
	LUT4 #(
		.INIT('h0100)
	) name2072 (
		_w2914_,
		_w2915_,
		_w2916_,
		_w3031_,
		_w3032_
	);
	LUT3 #(
		.INIT('h80)
	) name2073 (
		_w2907_,
		_w2912_,
		_w3032_,
		_w3033_
	);
	LUT4 #(
		.INIT('h00df)
	) name2074 (
		\u0_u1_tms_reg[19]/P0001 ,
		_w2918_,
		_w2930_,
		_w3033_,
		_w3034_
	);
	LUT2 #(
		.INIT('h2)
	) name2075 (
		_w1013_,
		_w3034_,
		_w3035_
	);
	LUT4 #(
		.INIT('hef00)
	) name2076 (
		\u0_rf_we_reg/NET0131 ,
		_w2693_,
		_w2706_,
		_w3035_,
		_w3036_
	);
	LUT2 #(
		.INIT('hd)
	) name2077 (
		_w3030_,
		_w3036_,
		_w3037_
	);
	LUT3 #(
		.INIT('h2a)
	) name2078 (
		\u0_tms_reg[1]/NET0131 ,
		wb_cyc_i_pad,
		wb_stb_i_pad,
		_w3038_
	);
	LUT2 #(
		.INIT('h4)
	) name2079 (
		\u0_rf_we_reg/NET0131 ,
		\u0_tms_reg[1]/NET0131 ,
		_w3039_
	);
	LUT4 #(
		.INIT('h0b0f)
	) name2080 (
		_w2693_,
		_w2706_,
		_w3038_,
		_w3039_,
		_w3040_
	);
	LUT3 #(
		.INIT('h4c)
	) name2081 (
		\u0_u0_csc_reg[8]/P0001 ,
		\u0_u0_tms_reg[1]/P0001 ,
		wb_we_i_pad,
		_w3041_
	);
	LUT4 #(
		.INIT('h0100)
	) name2082 (
		_w2914_,
		_w2915_,
		_w2916_,
		_w3041_,
		_w3042_
	);
	LUT3 #(
		.INIT('h80)
	) name2083 (
		_w2907_,
		_w2912_,
		_w3042_,
		_w3043_
	);
	LUT4 #(
		.INIT('h00df)
	) name2084 (
		\u0_u1_tms_reg[1]/P0001 ,
		_w2918_,
		_w2930_,
		_w3043_,
		_w3044_
	);
	LUT2 #(
		.INIT('h2)
	) name2085 (
		_w1013_,
		_w3044_,
		_w3045_
	);
	LUT4 #(
		.INIT('hef00)
	) name2086 (
		\u0_rf_we_reg/NET0131 ,
		_w2693_,
		_w2706_,
		_w3045_,
		_w3046_
	);
	LUT2 #(
		.INIT('hd)
	) name2087 (
		_w3040_,
		_w3046_,
		_w3047_
	);
	LUT3 #(
		.INIT('h2a)
	) name2088 (
		\u0_tms_reg[20]/NET0131 ,
		wb_cyc_i_pad,
		wb_stb_i_pad,
		_w3048_
	);
	LUT2 #(
		.INIT('h4)
	) name2089 (
		\u0_rf_we_reg/NET0131 ,
		\u0_tms_reg[20]/NET0131 ,
		_w3049_
	);
	LUT4 #(
		.INIT('h0b0f)
	) name2090 (
		_w2693_,
		_w2706_,
		_w3048_,
		_w3049_,
		_w3050_
	);
	LUT3 #(
		.INIT('h4c)
	) name2091 (
		\u0_u0_csc_reg[8]/P0001 ,
		\u0_u0_tms_reg[20]/P0001 ,
		wb_we_i_pad,
		_w3051_
	);
	LUT4 #(
		.INIT('h0100)
	) name2092 (
		_w2914_,
		_w2915_,
		_w2916_,
		_w3051_,
		_w3052_
	);
	LUT3 #(
		.INIT('h80)
	) name2093 (
		_w2907_,
		_w2912_,
		_w3052_,
		_w3053_
	);
	LUT4 #(
		.INIT('h00df)
	) name2094 (
		\u0_u1_tms_reg[20]/P0001 ,
		_w2918_,
		_w2930_,
		_w3053_,
		_w3054_
	);
	LUT2 #(
		.INIT('h2)
	) name2095 (
		_w1013_,
		_w3054_,
		_w3055_
	);
	LUT4 #(
		.INIT('hef00)
	) name2096 (
		\u0_rf_we_reg/NET0131 ,
		_w2693_,
		_w2706_,
		_w3055_,
		_w3056_
	);
	LUT2 #(
		.INIT('hd)
	) name2097 (
		_w3050_,
		_w3056_,
		_w3057_
	);
	LUT3 #(
		.INIT('h2a)
	) name2098 (
		\u0_tms_reg[21]/NET0131 ,
		wb_cyc_i_pad,
		wb_stb_i_pad,
		_w3058_
	);
	LUT2 #(
		.INIT('h4)
	) name2099 (
		\u0_rf_we_reg/NET0131 ,
		\u0_tms_reg[21]/NET0131 ,
		_w3059_
	);
	LUT4 #(
		.INIT('h0b0f)
	) name2100 (
		_w2693_,
		_w2706_,
		_w3058_,
		_w3059_,
		_w3060_
	);
	LUT3 #(
		.INIT('h4c)
	) name2101 (
		\u0_u0_csc_reg[8]/P0001 ,
		\u0_u0_tms_reg[21]/P0001 ,
		wb_we_i_pad,
		_w3061_
	);
	LUT4 #(
		.INIT('h0100)
	) name2102 (
		_w2914_,
		_w2915_,
		_w2916_,
		_w3061_,
		_w3062_
	);
	LUT3 #(
		.INIT('h80)
	) name2103 (
		_w2907_,
		_w2912_,
		_w3062_,
		_w3063_
	);
	LUT4 #(
		.INIT('h00df)
	) name2104 (
		\u0_u1_tms_reg[21]/P0001 ,
		_w2918_,
		_w2930_,
		_w3063_,
		_w3064_
	);
	LUT2 #(
		.INIT('h2)
	) name2105 (
		_w1013_,
		_w3064_,
		_w3065_
	);
	LUT4 #(
		.INIT('hef00)
	) name2106 (
		\u0_rf_we_reg/NET0131 ,
		_w2693_,
		_w2706_,
		_w3065_,
		_w3066_
	);
	LUT2 #(
		.INIT('hd)
	) name2107 (
		_w3060_,
		_w3066_,
		_w3067_
	);
	LUT3 #(
		.INIT('h2a)
	) name2108 (
		\u0_tms_reg[23]/NET0131 ,
		wb_cyc_i_pad,
		wb_stb_i_pad,
		_w3068_
	);
	LUT2 #(
		.INIT('h4)
	) name2109 (
		\u0_rf_we_reg/NET0131 ,
		\u0_tms_reg[23]/NET0131 ,
		_w3069_
	);
	LUT4 #(
		.INIT('h0b0f)
	) name2110 (
		_w2693_,
		_w2706_,
		_w3068_,
		_w3069_,
		_w3070_
	);
	LUT3 #(
		.INIT('h4c)
	) name2111 (
		\u0_u0_csc_reg[8]/P0001 ,
		\u0_u0_tms_reg[23]/P0001 ,
		wb_we_i_pad,
		_w3071_
	);
	LUT4 #(
		.INIT('h0100)
	) name2112 (
		_w2914_,
		_w2915_,
		_w2916_,
		_w3071_,
		_w3072_
	);
	LUT3 #(
		.INIT('h80)
	) name2113 (
		_w2907_,
		_w2912_,
		_w3072_,
		_w3073_
	);
	LUT4 #(
		.INIT('h00df)
	) name2114 (
		\u0_u1_tms_reg[23]/P0001 ,
		_w2918_,
		_w2930_,
		_w3073_,
		_w3074_
	);
	LUT2 #(
		.INIT('h2)
	) name2115 (
		_w1013_,
		_w3074_,
		_w3075_
	);
	LUT4 #(
		.INIT('hef00)
	) name2116 (
		\u0_rf_we_reg/NET0131 ,
		_w2693_,
		_w2706_,
		_w3075_,
		_w3076_
	);
	LUT2 #(
		.INIT('hd)
	) name2117 (
		_w3070_,
		_w3076_,
		_w3077_
	);
	LUT3 #(
		.INIT('h2a)
	) name2118 (
		\u0_tms_reg[24]/NET0131 ,
		wb_cyc_i_pad,
		wb_stb_i_pad,
		_w3078_
	);
	LUT2 #(
		.INIT('h4)
	) name2119 (
		\u0_rf_we_reg/NET0131 ,
		\u0_tms_reg[24]/NET0131 ,
		_w3079_
	);
	LUT4 #(
		.INIT('h0b0f)
	) name2120 (
		_w2693_,
		_w2706_,
		_w3078_,
		_w3079_,
		_w3080_
	);
	LUT3 #(
		.INIT('h4c)
	) name2121 (
		\u0_u0_csc_reg[8]/P0001 ,
		\u0_u0_tms_reg[24]/P0001 ,
		wb_we_i_pad,
		_w3081_
	);
	LUT4 #(
		.INIT('h0100)
	) name2122 (
		_w2914_,
		_w2915_,
		_w2916_,
		_w3081_,
		_w3082_
	);
	LUT3 #(
		.INIT('h80)
	) name2123 (
		_w2907_,
		_w2912_,
		_w3082_,
		_w3083_
	);
	LUT4 #(
		.INIT('h00df)
	) name2124 (
		\u0_u1_tms_reg[24]/P0001 ,
		_w2918_,
		_w2930_,
		_w3083_,
		_w3084_
	);
	LUT2 #(
		.INIT('h2)
	) name2125 (
		_w1013_,
		_w3084_,
		_w3085_
	);
	LUT4 #(
		.INIT('hef00)
	) name2126 (
		\u0_rf_we_reg/NET0131 ,
		_w2693_,
		_w2706_,
		_w3085_,
		_w3086_
	);
	LUT2 #(
		.INIT('hd)
	) name2127 (
		_w3080_,
		_w3086_,
		_w3087_
	);
	LUT3 #(
		.INIT('h2a)
	) name2128 (
		\u0_tms_reg[22]/NET0131 ,
		wb_cyc_i_pad,
		wb_stb_i_pad,
		_w3088_
	);
	LUT2 #(
		.INIT('h4)
	) name2129 (
		\u0_rf_we_reg/NET0131 ,
		\u0_tms_reg[22]/NET0131 ,
		_w3089_
	);
	LUT4 #(
		.INIT('h0b0f)
	) name2130 (
		_w2693_,
		_w2706_,
		_w3088_,
		_w3089_,
		_w3090_
	);
	LUT3 #(
		.INIT('h4c)
	) name2131 (
		\u0_u0_csc_reg[8]/P0001 ,
		\u0_u0_tms_reg[22]/P0001 ,
		wb_we_i_pad,
		_w3091_
	);
	LUT4 #(
		.INIT('h0100)
	) name2132 (
		_w2914_,
		_w2915_,
		_w2916_,
		_w3091_,
		_w3092_
	);
	LUT3 #(
		.INIT('h80)
	) name2133 (
		_w2907_,
		_w2912_,
		_w3092_,
		_w3093_
	);
	LUT4 #(
		.INIT('h00df)
	) name2134 (
		\u0_u1_tms_reg[22]/P0001 ,
		_w2918_,
		_w2930_,
		_w3093_,
		_w3094_
	);
	LUT2 #(
		.INIT('h2)
	) name2135 (
		_w1013_,
		_w3094_,
		_w3095_
	);
	LUT4 #(
		.INIT('hef00)
	) name2136 (
		\u0_rf_we_reg/NET0131 ,
		_w2693_,
		_w2706_,
		_w3095_,
		_w3096_
	);
	LUT2 #(
		.INIT('hd)
	) name2137 (
		_w3090_,
		_w3096_,
		_w3097_
	);
	LUT3 #(
		.INIT('h2a)
	) name2138 (
		\u0_tms_reg[25]/NET0131 ,
		wb_cyc_i_pad,
		wb_stb_i_pad,
		_w3098_
	);
	LUT2 #(
		.INIT('h4)
	) name2139 (
		\u0_rf_we_reg/NET0131 ,
		\u0_tms_reg[25]/NET0131 ,
		_w3099_
	);
	LUT4 #(
		.INIT('h0b0f)
	) name2140 (
		_w2693_,
		_w2706_,
		_w3098_,
		_w3099_,
		_w3100_
	);
	LUT3 #(
		.INIT('h4c)
	) name2141 (
		\u0_u0_csc_reg[8]/P0001 ,
		\u0_u0_tms_reg[25]/P0001 ,
		wb_we_i_pad,
		_w3101_
	);
	LUT4 #(
		.INIT('h0100)
	) name2142 (
		_w2914_,
		_w2915_,
		_w2916_,
		_w3101_,
		_w3102_
	);
	LUT3 #(
		.INIT('h80)
	) name2143 (
		_w2907_,
		_w2912_,
		_w3102_,
		_w3103_
	);
	LUT4 #(
		.INIT('h00df)
	) name2144 (
		\u0_u1_tms_reg[25]/P0001 ,
		_w2918_,
		_w2930_,
		_w3103_,
		_w3104_
	);
	LUT2 #(
		.INIT('h2)
	) name2145 (
		_w1013_,
		_w3104_,
		_w3105_
	);
	LUT4 #(
		.INIT('hef00)
	) name2146 (
		\u0_rf_we_reg/NET0131 ,
		_w2693_,
		_w2706_,
		_w3105_,
		_w3106_
	);
	LUT2 #(
		.INIT('hd)
	) name2147 (
		_w3100_,
		_w3106_,
		_w3107_
	);
	LUT3 #(
		.INIT('h2a)
	) name2148 (
		\u0_tms_reg[26]/NET0131 ,
		wb_cyc_i_pad,
		wb_stb_i_pad,
		_w3108_
	);
	LUT2 #(
		.INIT('h4)
	) name2149 (
		\u0_rf_we_reg/NET0131 ,
		\u0_tms_reg[26]/NET0131 ,
		_w3109_
	);
	LUT4 #(
		.INIT('h0b0f)
	) name2150 (
		_w2693_,
		_w2706_,
		_w3108_,
		_w3109_,
		_w3110_
	);
	LUT3 #(
		.INIT('h4c)
	) name2151 (
		\u0_u0_csc_reg[8]/P0001 ,
		\u0_u0_tms_reg[26]/P0001 ,
		wb_we_i_pad,
		_w3111_
	);
	LUT4 #(
		.INIT('h0100)
	) name2152 (
		_w2914_,
		_w2915_,
		_w2916_,
		_w3111_,
		_w3112_
	);
	LUT3 #(
		.INIT('h80)
	) name2153 (
		_w2907_,
		_w2912_,
		_w3112_,
		_w3113_
	);
	LUT4 #(
		.INIT('h00df)
	) name2154 (
		\u0_u1_tms_reg[26]/P0001 ,
		_w2918_,
		_w2930_,
		_w3113_,
		_w3114_
	);
	LUT2 #(
		.INIT('h2)
	) name2155 (
		_w1013_,
		_w3114_,
		_w3115_
	);
	LUT4 #(
		.INIT('hef00)
	) name2156 (
		\u0_rf_we_reg/NET0131 ,
		_w2693_,
		_w2706_,
		_w3115_,
		_w3116_
	);
	LUT2 #(
		.INIT('hd)
	) name2157 (
		_w3110_,
		_w3116_,
		_w3117_
	);
	LUT3 #(
		.INIT('h2a)
	) name2158 (
		\u0_tms_reg[27]/NET0131 ,
		wb_cyc_i_pad,
		wb_stb_i_pad,
		_w3118_
	);
	LUT2 #(
		.INIT('h4)
	) name2159 (
		\u0_rf_we_reg/NET0131 ,
		\u0_tms_reg[27]/NET0131 ,
		_w3119_
	);
	LUT4 #(
		.INIT('h0b0f)
	) name2160 (
		_w2693_,
		_w2706_,
		_w3118_,
		_w3119_,
		_w3120_
	);
	LUT3 #(
		.INIT('h4c)
	) name2161 (
		\u0_u0_csc_reg[8]/P0001 ,
		\u0_u0_tms_reg[27]/P0001 ,
		wb_we_i_pad,
		_w3121_
	);
	LUT4 #(
		.INIT('h0100)
	) name2162 (
		_w2914_,
		_w2915_,
		_w2916_,
		_w3121_,
		_w3122_
	);
	LUT3 #(
		.INIT('h80)
	) name2163 (
		_w2907_,
		_w2912_,
		_w3122_,
		_w3123_
	);
	LUT4 #(
		.INIT('h00df)
	) name2164 (
		\u0_u1_tms_reg[27]/P0001 ,
		_w2918_,
		_w2930_,
		_w3123_,
		_w3124_
	);
	LUT2 #(
		.INIT('h2)
	) name2165 (
		_w1013_,
		_w3124_,
		_w3125_
	);
	LUT4 #(
		.INIT('hef00)
	) name2166 (
		\u0_rf_we_reg/NET0131 ,
		_w2693_,
		_w2706_,
		_w3125_,
		_w3126_
	);
	LUT2 #(
		.INIT('hd)
	) name2167 (
		_w3120_,
		_w3126_,
		_w3127_
	);
	LUT3 #(
		.INIT('h2a)
	) name2168 (
		\u0_tms_reg[2]/NET0131 ,
		wb_cyc_i_pad,
		wb_stb_i_pad,
		_w3128_
	);
	LUT2 #(
		.INIT('h4)
	) name2169 (
		\u0_rf_we_reg/NET0131 ,
		\u0_tms_reg[2]/NET0131 ,
		_w3129_
	);
	LUT4 #(
		.INIT('h0b0f)
	) name2170 (
		_w2693_,
		_w2706_,
		_w3128_,
		_w3129_,
		_w3130_
	);
	LUT3 #(
		.INIT('h4c)
	) name2171 (
		\u0_u0_csc_reg[8]/P0001 ,
		\u0_u0_tms_reg[2]/P0001 ,
		wb_we_i_pad,
		_w3131_
	);
	LUT4 #(
		.INIT('h0100)
	) name2172 (
		_w2914_,
		_w2915_,
		_w2916_,
		_w3131_,
		_w3132_
	);
	LUT3 #(
		.INIT('h80)
	) name2173 (
		_w2907_,
		_w2912_,
		_w3132_,
		_w3133_
	);
	LUT4 #(
		.INIT('h00df)
	) name2174 (
		\u0_u1_tms_reg[2]/P0001 ,
		_w2918_,
		_w2930_,
		_w3133_,
		_w3134_
	);
	LUT2 #(
		.INIT('h2)
	) name2175 (
		_w1013_,
		_w3134_,
		_w3135_
	);
	LUT4 #(
		.INIT('hef00)
	) name2176 (
		\u0_rf_we_reg/NET0131 ,
		_w2693_,
		_w2706_,
		_w3135_,
		_w3136_
	);
	LUT2 #(
		.INIT('hd)
	) name2177 (
		_w3130_,
		_w3136_,
		_w3137_
	);
	LUT3 #(
		.INIT('h2a)
	) name2178 (
		\u0_tms_reg[3]/NET0131 ,
		wb_cyc_i_pad,
		wb_stb_i_pad,
		_w3138_
	);
	LUT2 #(
		.INIT('h4)
	) name2179 (
		\u0_rf_we_reg/NET0131 ,
		\u0_tms_reg[3]/NET0131 ,
		_w3139_
	);
	LUT4 #(
		.INIT('h0b0f)
	) name2180 (
		_w2693_,
		_w2706_,
		_w3138_,
		_w3139_,
		_w3140_
	);
	LUT3 #(
		.INIT('h4c)
	) name2181 (
		\u0_u0_csc_reg[8]/P0001 ,
		\u0_u0_tms_reg[3]/P0001 ,
		wb_we_i_pad,
		_w3141_
	);
	LUT4 #(
		.INIT('h0100)
	) name2182 (
		_w2914_,
		_w2915_,
		_w2916_,
		_w3141_,
		_w3142_
	);
	LUT3 #(
		.INIT('h80)
	) name2183 (
		_w2907_,
		_w2912_,
		_w3142_,
		_w3143_
	);
	LUT4 #(
		.INIT('h00df)
	) name2184 (
		\u0_u1_tms_reg[3]/P0001 ,
		_w2918_,
		_w2930_,
		_w3143_,
		_w3144_
	);
	LUT2 #(
		.INIT('h2)
	) name2185 (
		_w1013_,
		_w3144_,
		_w3145_
	);
	LUT4 #(
		.INIT('hef00)
	) name2186 (
		\u0_rf_we_reg/NET0131 ,
		_w2693_,
		_w2706_,
		_w3145_,
		_w3146_
	);
	LUT2 #(
		.INIT('hd)
	) name2187 (
		_w3140_,
		_w3146_,
		_w3147_
	);
	LUT3 #(
		.INIT('h2a)
	) name2188 (
		\u0_tms_reg[4]/NET0131 ,
		wb_cyc_i_pad,
		wb_stb_i_pad,
		_w3148_
	);
	LUT2 #(
		.INIT('h4)
	) name2189 (
		\u0_rf_we_reg/NET0131 ,
		\u0_tms_reg[4]/NET0131 ,
		_w3149_
	);
	LUT4 #(
		.INIT('h0b0f)
	) name2190 (
		_w2693_,
		_w2706_,
		_w3148_,
		_w3149_,
		_w3150_
	);
	LUT3 #(
		.INIT('h4c)
	) name2191 (
		\u0_u0_csc_reg[8]/P0001 ,
		\u0_u0_tms_reg[4]/P0001 ,
		wb_we_i_pad,
		_w3151_
	);
	LUT4 #(
		.INIT('h0100)
	) name2192 (
		_w2914_,
		_w2915_,
		_w2916_,
		_w3151_,
		_w3152_
	);
	LUT3 #(
		.INIT('h80)
	) name2193 (
		_w2907_,
		_w2912_,
		_w3152_,
		_w3153_
	);
	LUT4 #(
		.INIT('h00df)
	) name2194 (
		\u0_u1_tms_reg[4]/P0001 ,
		_w2918_,
		_w2930_,
		_w3153_,
		_w3154_
	);
	LUT2 #(
		.INIT('h2)
	) name2195 (
		_w1013_,
		_w3154_,
		_w3155_
	);
	LUT4 #(
		.INIT('hef00)
	) name2196 (
		\u0_rf_we_reg/NET0131 ,
		_w2693_,
		_w2706_,
		_w3155_,
		_w3156_
	);
	LUT2 #(
		.INIT('hd)
	) name2197 (
		_w3150_,
		_w3156_,
		_w3157_
	);
	LUT3 #(
		.INIT('h2a)
	) name2198 (
		\u0_tms_reg[5]/NET0131 ,
		wb_cyc_i_pad,
		wb_stb_i_pad,
		_w3158_
	);
	LUT2 #(
		.INIT('h4)
	) name2199 (
		\u0_rf_we_reg/NET0131 ,
		\u0_tms_reg[5]/NET0131 ,
		_w3159_
	);
	LUT4 #(
		.INIT('h0b0f)
	) name2200 (
		_w2693_,
		_w2706_,
		_w3158_,
		_w3159_,
		_w3160_
	);
	LUT3 #(
		.INIT('h4c)
	) name2201 (
		\u0_u0_csc_reg[8]/P0001 ,
		\u0_u0_tms_reg[5]/P0001 ,
		wb_we_i_pad,
		_w3161_
	);
	LUT4 #(
		.INIT('h0100)
	) name2202 (
		_w2914_,
		_w2915_,
		_w2916_,
		_w3161_,
		_w3162_
	);
	LUT3 #(
		.INIT('h80)
	) name2203 (
		_w2907_,
		_w2912_,
		_w3162_,
		_w3163_
	);
	LUT4 #(
		.INIT('h00df)
	) name2204 (
		\u0_u1_tms_reg[5]/P0001 ,
		_w2918_,
		_w2930_,
		_w3163_,
		_w3164_
	);
	LUT2 #(
		.INIT('h2)
	) name2205 (
		_w1013_,
		_w3164_,
		_w3165_
	);
	LUT4 #(
		.INIT('hef00)
	) name2206 (
		\u0_rf_we_reg/NET0131 ,
		_w2693_,
		_w2706_,
		_w3165_,
		_w3166_
	);
	LUT2 #(
		.INIT('hd)
	) name2207 (
		_w3160_,
		_w3166_,
		_w3167_
	);
	LUT3 #(
		.INIT('h2a)
	) name2208 (
		\u0_tms_reg[6]/NET0131 ,
		wb_cyc_i_pad,
		wb_stb_i_pad,
		_w3168_
	);
	LUT2 #(
		.INIT('h4)
	) name2209 (
		\u0_rf_we_reg/NET0131 ,
		\u0_tms_reg[6]/NET0131 ,
		_w3169_
	);
	LUT4 #(
		.INIT('h0b0f)
	) name2210 (
		_w2693_,
		_w2706_,
		_w3168_,
		_w3169_,
		_w3170_
	);
	LUT3 #(
		.INIT('h4c)
	) name2211 (
		\u0_u0_csc_reg[8]/P0001 ,
		\u0_u0_tms_reg[6]/P0001 ,
		wb_we_i_pad,
		_w3171_
	);
	LUT4 #(
		.INIT('h0100)
	) name2212 (
		_w2914_,
		_w2915_,
		_w2916_,
		_w3171_,
		_w3172_
	);
	LUT3 #(
		.INIT('h80)
	) name2213 (
		_w2907_,
		_w2912_,
		_w3172_,
		_w3173_
	);
	LUT4 #(
		.INIT('h00df)
	) name2214 (
		\u0_u1_tms_reg[6]/P0001 ,
		_w2918_,
		_w2930_,
		_w3173_,
		_w3174_
	);
	LUT2 #(
		.INIT('h2)
	) name2215 (
		_w1013_,
		_w3174_,
		_w3175_
	);
	LUT4 #(
		.INIT('hef00)
	) name2216 (
		\u0_rf_we_reg/NET0131 ,
		_w2693_,
		_w2706_,
		_w3175_,
		_w3176_
	);
	LUT2 #(
		.INIT('hd)
	) name2217 (
		_w3170_,
		_w3176_,
		_w3177_
	);
	LUT3 #(
		.INIT('h2a)
	) name2218 (
		\u0_tms_reg[7]/NET0131 ,
		wb_cyc_i_pad,
		wb_stb_i_pad,
		_w3178_
	);
	LUT2 #(
		.INIT('h4)
	) name2219 (
		\u0_rf_we_reg/NET0131 ,
		\u0_tms_reg[7]/NET0131 ,
		_w3179_
	);
	LUT4 #(
		.INIT('h0b0f)
	) name2220 (
		_w2693_,
		_w2706_,
		_w3178_,
		_w3179_,
		_w3180_
	);
	LUT3 #(
		.INIT('h4c)
	) name2221 (
		\u0_u0_csc_reg[8]/P0001 ,
		\u0_u0_tms_reg[7]/P0001 ,
		wb_we_i_pad,
		_w3181_
	);
	LUT4 #(
		.INIT('h0100)
	) name2222 (
		_w2914_,
		_w2915_,
		_w2916_,
		_w3181_,
		_w3182_
	);
	LUT3 #(
		.INIT('h80)
	) name2223 (
		_w2907_,
		_w2912_,
		_w3182_,
		_w3183_
	);
	LUT4 #(
		.INIT('h00df)
	) name2224 (
		\u0_u1_tms_reg[7]/P0001 ,
		_w2918_,
		_w2930_,
		_w3183_,
		_w3184_
	);
	LUT2 #(
		.INIT('h2)
	) name2225 (
		_w1013_,
		_w3184_,
		_w3185_
	);
	LUT4 #(
		.INIT('hef00)
	) name2226 (
		\u0_rf_we_reg/NET0131 ,
		_w2693_,
		_w2706_,
		_w3185_,
		_w3186_
	);
	LUT2 #(
		.INIT('hd)
	) name2227 (
		_w3180_,
		_w3186_,
		_w3187_
	);
	LUT3 #(
		.INIT('h2a)
	) name2228 (
		\u0_tms_reg[8]/NET0131 ,
		wb_cyc_i_pad,
		wb_stb_i_pad,
		_w3188_
	);
	LUT2 #(
		.INIT('h4)
	) name2229 (
		\u0_rf_we_reg/NET0131 ,
		\u0_tms_reg[8]/NET0131 ,
		_w3189_
	);
	LUT4 #(
		.INIT('h0b0f)
	) name2230 (
		_w2693_,
		_w2706_,
		_w3188_,
		_w3189_,
		_w3190_
	);
	LUT3 #(
		.INIT('h4c)
	) name2231 (
		\u0_u0_csc_reg[8]/P0001 ,
		\u0_u0_tms_reg[8]/P0001 ,
		wb_we_i_pad,
		_w3191_
	);
	LUT4 #(
		.INIT('h0100)
	) name2232 (
		_w2914_,
		_w2915_,
		_w2916_,
		_w3191_,
		_w3192_
	);
	LUT3 #(
		.INIT('h80)
	) name2233 (
		_w2907_,
		_w2912_,
		_w3192_,
		_w3193_
	);
	LUT4 #(
		.INIT('h00df)
	) name2234 (
		\u0_u1_tms_reg[8]/P0001 ,
		_w2918_,
		_w2930_,
		_w3193_,
		_w3194_
	);
	LUT2 #(
		.INIT('h2)
	) name2235 (
		_w1013_,
		_w3194_,
		_w3195_
	);
	LUT4 #(
		.INIT('hef00)
	) name2236 (
		\u0_rf_we_reg/NET0131 ,
		_w2693_,
		_w2706_,
		_w3195_,
		_w3196_
	);
	LUT2 #(
		.INIT('hd)
	) name2237 (
		_w3190_,
		_w3196_,
		_w3197_
	);
	LUT3 #(
		.INIT('h2a)
	) name2238 (
		\u0_tms_reg[9]/NET0131 ,
		wb_cyc_i_pad,
		wb_stb_i_pad,
		_w3198_
	);
	LUT2 #(
		.INIT('h4)
	) name2239 (
		\u0_rf_we_reg/NET0131 ,
		\u0_tms_reg[9]/NET0131 ,
		_w3199_
	);
	LUT4 #(
		.INIT('h0b0f)
	) name2240 (
		_w2693_,
		_w2706_,
		_w3198_,
		_w3199_,
		_w3200_
	);
	LUT3 #(
		.INIT('h4c)
	) name2241 (
		\u0_u0_csc_reg[8]/P0001 ,
		\u0_u0_tms_reg[9]/P0001 ,
		wb_we_i_pad,
		_w3201_
	);
	LUT4 #(
		.INIT('h0100)
	) name2242 (
		_w2914_,
		_w2915_,
		_w2916_,
		_w3201_,
		_w3202_
	);
	LUT3 #(
		.INIT('h80)
	) name2243 (
		_w2907_,
		_w2912_,
		_w3202_,
		_w3203_
	);
	LUT4 #(
		.INIT('h00df)
	) name2244 (
		\u0_u1_tms_reg[9]/P0001 ,
		_w2918_,
		_w2930_,
		_w3203_,
		_w3204_
	);
	LUT2 #(
		.INIT('h2)
	) name2245 (
		_w1013_,
		_w3204_,
		_w3205_
	);
	LUT4 #(
		.INIT('hef00)
	) name2246 (
		\u0_rf_we_reg/NET0131 ,
		_w2693_,
		_w2706_,
		_w3205_,
		_w3206_
	);
	LUT2 #(
		.INIT('hd)
	) name2247 (
		_w3200_,
		_w3206_,
		_w3207_
	);
	LUT3 #(
		.INIT('hb0)
	) name2248 (
		_w1539_,
		_w1898_,
		_w2383_,
		_w3208_
	);
	LUT3 #(
		.INIT('h02)
	) name2249 (
		\u0_tms_reg[6]/NET0131 ,
		\u5_lmr_ack_reg/NET0131 ,
		\u5_state_reg[26]/NET0131 ,
		_w3209_
	);
	LUT4 #(
		.INIT('h11d5)
	) name2250 (
		\u0_sp_tms_reg[6]/NET0131 ,
		_w976_,
		_w1114_,
		_w3209_,
		_w3210_
	);
	LUT2 #(
		.INIT('h4)
	) name2251 (
		_w2402_,
		_w3210_,
		_w3211_
	);
	LUT3 #(
		.INIT('h80)
	) name2252 (
		_w1540_,
		_w1541_,
		_w3211_,
		_w3212_
	);
	LUT4 #(
		.INIT('hb555)
	) name2253 (
		\u5_timer2_reg[7]/P0001 ,
		\u5_timer2_reg[8]/P0001 ,
		_w2398_,
		_w2399_,
		_w3213_
	);
	LUT3 #(
		.INIT('h2a)
	) name2254 (
		_w2397_,
		_w2402_,
		_w3213_,
		_w3214_
	);
	LUT4 #(
		.INIT('h8c00)
	) name2255 (
		_w1539_,
		_w2542_,
		_w3212_,
		_w3214_,
		_w3215_
	);
	LUT2 #(
		.INIT('he)
	) name2256 (
		_w3208_,
		_w3215_,
		_w3216_
	);
	LUT3 #(
		.INIT('h8c)
	) name2257 (
		_w1539_,
		_w2383_,
		_w2558_,
		_w3217_
	);
	LUT3 #(
		.INIT('h02)
	) name2258 (
		\u0_tms_reg[7]/NET0131 ,
		\u5_lmr_ack_reg/NET0131 ,
		\u5_state_reg[26]/NET0131 ,
		_w3218_
	);
	LUT4 #(
		.INIT('h11d5)
	) name2259 (
		\u0_sp_tms_reg[7]/NET0131 ,
		_w976_,
		_w1114_,
		_w3218_,
		_w3219_
	);
	LUT2 #(
		.INIT('h4)
	) name2260 (
		_w2402_,
		_w3219_,
		_w3220_
	);
	LUT3 #(
		.INIT('h80)
	) name2261 (
		_w1540_,
		_w1541_,
		_w3220_,
		_w3221_
	);
	LUT2 #(
		.INIT('h4)
	) name2262 (
		\u5_timer2_reg[8]/P0001 ,
		_w2402_,
		_w3222_
	);
	LUT4 #(
		.INIT('h4000)
	) name2263 (
		\u5_timer2_reg[7]/P0001 ,
		_w2398_,
		_w2399_,
		_w2402_,
		_w3223_
	);
	LUT3 #(
		.INIT('h02)
	) name2264 (
		_w2397_,
		_w3222_,
		_w3223_,
		_w3224_
	);
	LUT4 #(
		.INIT('h8c00)
	) name2265 (
		_w1539_,
		_w2542_,
		_w3221_,
		_w3224_,
		_w3225_
	);
	LUT2 #(
		.INIT('he)
	) name2266 (
		_w3217_,
		_w3225_,
		_w3226_
	);
	LUT3 #(
		.INIT('h2a)
	) name2267 (
		\wb_addr_i[16]_pad ,
		_w976_,
		_w1975_,
		_w3227_
	);
	LUT3 #(
		.INIT('h10)
	) name2268 (
		_w1972_,
		_w1974_,
		_w3227_,
		_w3228_
	);
	LUT3 #(
		.INIT('h2a)
	) name2269 (
		\wb_addr_i[15]_pad ,
		_w976_,
		_w1971_,
		_w3229_
	);
	LUT3 #(
		.INIT('h40)
	) name2270 (
		_w1970_,
		_w1976_,
		_w3229_,
		_w3230_
	);
	LUT3 #(
		.INIT('h2a)
	) name2271 (
		\wb_addr_i[17]_pad ,
		_w976_,
		_w1971_,
		_w3231_
	);
	LUT3 #(
		.INIT('h10)
	) name2272 (
		_w1970_,
		_w1976_,
		_w3231_,
		_w3232_
	);
	LUT4 #(
		.INIT('haebf)
	) name2273 (
		_w1970_,
		_w1976_,
		_w3229_,
		_w3231_,
		_w3233_
	);
	LUT3 #(
		.INIT('h45)
	) name2274 (
		_w2424_,
		_w3228_,
		_w3233_,
		_w3234_
	);
	LUT2 #(
		.INIT('h8)
	) name2275 (
		\u1_acs_addr_reg[13]/P0001 ,
		\u1_acs_addr_reg[14]/P0001 ,
		_w3235_
	);
	LUT3 #(
		.INIT('h15)
	) name2276 (
		\u1_acs_addr_reg[15]/P0001 ,
		_w2419_,
		_w3235_,
		_w3236_
	);
	LUT3 #(
		.INIT('h70)
	) name2277 (
		_w2419_,
		_w2420_,
		_w2424_,
		_w3237_
	);
	LUT3 #(
		.INIT('hba)
	) name2278 (
		_w3234_,
		_w3236_,
		_w3237_,
		_w3238_
	);
	LUT3 #(
		.INIT('h8a)
	) name2279 (
		_w1013_,
		_w2693_,
		_w2706_,
		_w3239_
	);
	LUT4 #(
		.INIT('h2a22)
	) name2280 (
		\u0_csc_reg[4]/NET0131 ,
		_w1013_,
		_w2693_,
		_w2706_,
		_w3240_
	);
	LUT3 #(
		.INIT('h80)
	) name2281 (
		\u0_u1_csc_reg[4]/P0001 ,
		wb_cyc_i_pad,
		wb_stb_i_pad,
		_w3241_
	);
	LUT3 #(
		.INIT('h40)
	) name2282 (
		_w2918_,
		_w2930_,
		_w3241_,
		_w3242_
	);
	LUT3 #(
		.INIT('h80)
	) name2283 (
		\u0_u0_csc_reg[4]/P0001 ,
		wb_cyc_i_pad,
		wb_stb_i_pad,
		_w3243_
	);
	LUT4 #(
		.INIT('h8000)
	) name2284 (
		_w2907_,
		_w2912_,
		_w2917_,
		_w3243_,
		_w3244_
	);
	LUT4 #(
		.INIT('h444f)
	) name2285 (
		_w2693_,
		_w2706_,
		_w3242_,
		_w3244_,
		_w3245_
	);
	LUT2 #(
		.INIT('hb)
	) name2286 (
		_w3240_,
		_w3245_,
		_w3246_
	);
	LUT4 #(
		.INIT('h2a22)
	) name2287 (
		\u0_csc_reg[5]/NET0131 ,
		_w1013_,
		_w2693_,
		_w2706_,
		_w3247_
	);
	LUT3 #(
		.INIT('h80)
	) name2288 (
		\u0_u1_csc_reg[5]/P0001 ,
		wb_cyc_i_pad,
		wb_stb_i_pad,
		_w3248_
	);
	LUT3 #(
		.INIT('h40)
	) name2289 (
		_w2918_,
		_w2930_,
		_w3248_,
		_w3249_
	);
	LUT3 #(
		.INIT('h80)
	) name2290 (
		\u0_u0_csc_reg[5]/P0001 ,
		wb_cyc_i_pad,
		wb_stb_i_pad,
		_w3250_
	);
	LUT4 #(
		.INIT('h8000)
	) name2291 (
		_w2907_,
		_w2912_,
		_w2917_,
		_w3250_,
		_w3251_
	);
	LUT4 #(
		.INIT('h444f)
	) name2292 (
		_w2693_,
		_w2706_,
		_w3249_,
		_w3251_,
		_w3252_
	);
	LUT2 #(
		.INIT('hb)
	) name2293 (
		_w3247_,
		_w3252_,
		_w3253_
	);
	LUT4 #(
		.INIT('h2a22)
	) name2294 (
		\u0_csc_reg[6]/NET0131 ,
		_w1013_,
		_w2693_,
		_w2706_,
		_w3254_
	);
	LUT3 #(
		.INIT('h80)
	) name2295 (
		\u0_u0_csc_reg[6]/P0001 ,
		wb_cyc_i_pad,
		wb_stb_i_pad,
		_w3255_
	);
	LUT4 #(
		.INIT('h8000)
	) name2296 (
		_w2907_,
		_w2912_,
		_w2917_,
		_w3255_,
		_w3256_
	);
	LUT3 #(
		.INIT('h80)
	) name2297 (
		\u0_u1_csc_reg[6]/P0001 ,
		wb_cyc_i_pad,
		wb_stb_i_pad,
		_w3257_
	);
	LUT3 #(
		.INIT('h40)
	) name2298 (
		_w2918_,
		_w2930_,
		_w3257_,
		_w3258_
	);
	LUT4 #(
		.INIT('h444f)
	) name2299 (
		_w2693_,
		_w2706_,
		_w3256_,
		_w3258_,
		_w3259_
	);
	LUT2 #(
		.INIT('hb)
	) name2300 (
		_w3254_,
		_w3259_,
		_w3260_
	);
	LUT4 #(
		.INIT('h2a22)
	) name2301 (
		\u0_csc_reg[9]/NET0131 ,
		_w1013_,
		_w2693_,
		_w2706_,
		_w3261_
	);
	LUT3 #(
		.INIT('h80)
	) name2302 (
		\u0_u0_csc_reg[9]/P0001 ,
		wb_cyc_i_pad,
		wb_stb_i_pad,
		_w3262_
	);
	LUT4 #(
		.INIT('h8000)
	) name2303 (
		_w2907_,
		_w2912_,
		_w2917_,
		_w3262_,
		_w3263_
	);
	LUT3 #(
		.INIT('h80)
	) name2304 (
		\u0_u1_csc_reg[9]/P0001 ,
		wb_cyc_i_pad,
		wb_stb_i_pad,
		_w3264_
	);
	LUT3 #(
		.INIT('h40)
	) name2305 (
		_w2918_,
		_w2930_,
		_w3264_,
		_w3265_
	);
	LUT4 #(
		.INIT('h444f)
	) name2306 (
		_w2693_,
		_w2706_,
		_w3263_,
		_w3265_,
		_w3266_
	);
	LUT2 #(
		.INIT('hb)
	) name2307 (
		_w3261_,
		_w3266_,
		_w3267_
	);
	LUT4 #(
		.INIT('h2a22)
	) name2308 (
		\u0_csc_reg[7]/NET0131 ,
		_w1013_,
		_w2693_,
		_w2706_,
		_w3268_
	);
	LUT3 #(
		.INIT('h80)
	) name2309 (
		\u0_u0_csc_reg[7]/P0001 ,
		wb_cyc_i_pad,
		wb_stb_i_pad,
		_w3269_
	);
	LUT4 #(
		.INIT('h8000)
	) name2310 (
		_w2907_,
		_w2912_,
		_w2917_,
		_w3269_,
		_w3270_
	);
	LUT3 #(
		.INIT('h80)
	) name2311 (
		\u0_u1_csc_reg[7]/P0001 ,
		wb_cyc_i_pad,
		wb_stb_i_pad,
		_w3271_
	);
	LUT3 #(
		.INIT('h40)
	) name2312 (
		_w2918_,
		_w2930_,
		_w3271_,
		_w3272_
	);
	LUT4 #(
		.INIT('h444f)
	) name2313 (
		_w2693_,
		_w2706_,
		_w3270_,
		_w3272_,
		_w3273_
	);
	LUT2 #(
		.INIT('hb)
	) name2314 (
		_w3268_,
		_w3273_,
		_w3274_
	);
	LUT4 #(
		.INIT('h2a22)
	) name2315 (
		\u0_sp_csc_reg[10]/NET0131 ,
		_w1013_,
		_w2693_,
		_w2706_,
		_w3275_
	);
	LUT4 #(
		.INIT('h8000)
	) name2316 (
		\u0_spec_req_cs_reg[0]/NET0131 ,
		\u0_u0_csc_reg[10]/P0001 ,
		wb_cyc_i_pad,
		wb_stb_i_pad,
		_w3276_
	);
	LUT3 #(
		.INIT('h80)
	) name2317 (
		\u0_u1_csc_reg[10]/P0001 ,
		wb_cyc_i_pad,
		wb_stb_i_pad,
		_w3277_
	);
	LUT2 #(
		.INIT('h8)
	) name2318 (
		_w2710_,
		_w3277_,
		_w3278_
	);
	LUT4 #(
		.INIT('h444f)
	) name2319 (
		_w2693_,
		_w2706_,
		_w3276_,
		_w3278_,
		_w3279_
	);
	LUT2 #(
		.INIT('hb)
	) name2320 (
		_w3275_,
		_w3279_,
		_w3280_
	);
	LUT4 #(
		.INIT('h2a22)
	) name2321 (
		\u0_sp_csc_reg[4]/NET0131 ,
		_w1013_,
		_w2693_,
		_w2706_,
		_w3281_
	);
	LUT4 #(
		.INIT('h8000)
	) name2322 (
		\u0_spec_req_cs_reg[0]/NET0131 ,
		\u0_u0_csc_reg[4]/P0001 ,
		wb_cyc_i_pad,
		wb_stb_i_pad,
		_w3282_
	);
	LUT2 #(
		.INIT('h8)
	) name2323 (
		_w2710_,
		_w3241_,
		_w3283_
	);
	LUT4 #(
		.INIT('h444f)
	) name2324 (
		_w2693_,
		_w2706_,
		_w3282_,
		_w3283_,
		_w3284_
	);
	LUT2 #(
		.INIT('hb)
	) name2325 (
		_w3281_,
		_w3284_,
		_w3285_
	);
	LUT4 #(
		.INIT('h2a22)
	) name2326 (
		\u0_sp_csc_reg[5]/NET0131 ,
		_w1013_,
		_w2693_,
		_w2706_,
		_w3286_
	);
	LUT4 #(
		.INIT('h8000)
	) name2327 (
		\u0_spec_req_cs_reg[0]/NET0131 ,
		\u0_u0_csc_reg[5]/P0001 ,
		wb_cyc_i_pad,
		wb_stb_i_pad,
		_w3287_
	);
	LUT2 #(
		.INIT('h8)
	) name2328 (
		_w2710_,
		_w3248_,
		_w3288_
	);
	LUT4 #(
		.INIT('h444f)
	) name2329 (
		_w2693_,
		_w2706_,
		_w3287_,
		_w3288_,
		_w3289_
	);
	LUT2 #(
		.INIT('hb)
	) name2330 (
		_w3286_,
		_w3289_,
		_w3290_
	);
	LUT4 #(
		.INIT('h2a22)
	) name2331 (
		\u0_sp_csc_reg[6]/NET0131 ,
		_w1013_,
		_w2693_,
		_w2706_,
		_w3291_
	);
	LUT4 #(
		.INIT('h8000)
	) name2332 (
		\u0_spec_req_cs_reg[0]/NET0131 ,
		\u0_u0_csc_reg[6]/P0001 ,
		wb_cyc_i_pad,
		wb_stb_i_pad,
		_w3292_
	);
	LUT2 #(
		.INIT('h8)
	) name2333 (
		_w2710_,
		_w3257_,
		_w3293_
	);
	LUT4 #(
		.INIT('h444f)
	) name2334 (
		_w2693_,
		_w2706_,
		_w3292_,
		_w3293_,
		_w3294_
	);
	LUT2 #(
		.INIT('hb)
	) name2335 (
		_w3291_,
		_w3294_,
		_w3295_
	);
	LUT4 #(
		.INIT('h2a22)
	) name2336 (
		\u0_sp_csc_reg[7]/NET0131 ,
		_w1013_,
		_w2693_,
		_w2706_,
		_w3296_
	);
	LUT4 #(
		.INIT('h8000)
	) name2337 (
		\u0_spec_req_cs_reg[0]/NET0131 ,
		\u0_u0_csc_reg[7]/P0001 ,
		wb_cyc_i_pad,
		wb_stb_i_pad,
		_w3297_
	);
	LUT2 #(
		.INIT('h8)
	) name2338 (
		_w2710_,
		_w3271_,
		_w3298_
	);
	LUT4 #(
		.INIT('h444f)
	) name2339 (
		_w2693_,
		_w2706_,
		_w3297_,
		_w3298_,
		_w3299_
	);
	LUT2 #(
		.INIT('hb)
	) name2340 (
		_w3296_,
		_w3299_,
		_w3300_
	);
	LUT4 #(
		.INIT('h2a22)
	) name2341 (
		\u0_sp_csc_reg[9]/NET0131 ,
		_w1013_,
		_w2693_,
		_w2706_,
		_w3301_
	);
	LUT4 #(
		.INIT('h8000)
	) name2342 (
		\u0_spec_req_cs_reg[0]/NET0131 ,
		\u0_u0_csc_reg[9]/P0001 ,
		wb_cyc_i_pad,
		wb_stb_i_pad,
		_w3302_
	);
	LUT2 #(
		.INIT('h8)
	) name2343 (
		_w2710_,
		_w3264_,
		_w3303_
	);
	LUT4 #(
		.INIT('h444f)
	) name2344 (
		_w2693_,
		_w2706_,
		_w3302_,
		_w3303_,
		_w3304_
	);
	LUT2 #(
		.INIT('hb)
	) name2345 (
		_w3301_,
		_w3304_,
		_w3305_
	);
	LUT4 #(
		.INIT('h2a22)
	) name2346 (
		\u0_csc_reg[10]/NET0131 ,
		_w1013_,
		_w2693_,
		_w2706_,
		_w3306_
	);
	LUT3 #(
		.INIT('h40)
	) name2347 (
		_w2918_,
		_w2930_,
		_w3277_,
		_w3307_
	);
	LUT3 #(
		.INIT('h80)
	) name2348 (
		\u0_u0_csc_reg[10]/P0001 ,
		wb_cyc_i_pad,
		wb_stb_i_pad,
		_w3308_
	);
	LUT4 #(
		.INIT('h8000)
	) name2349 (
		_w2907_,
		_w2912_,
		_w2917_,
		_w3308_,
		_w3309_
	);
	LUT4 #(
		.INIT('h444f)
	) name2350 (
		_w2693_,
		_w2706_,
		_w3307_,
		_w3309_,
		_w3310_
	);
	LUT2 #(
		.INIT('hb)
	) name2351 (
		_w3306_,
		_w3310_,
		_w3311_
	);
	LUT2 #(
		.INIT('h2)
	) name2352 (
		\u5_ap_en_reg/NET0131 ,
		\u5_state_reg[1]/NET0131 ,
		_w3312_
	);
	LUT3 #(
		.INIT('h80)
	) name2353 (
		_w1119_,
		_w1122_,
		_w1124_,
		_w3313_
	);
	LUT4 #(
		.INIT('hf4f0)
	) name2354 (
		_w1539_,
		_w2001_,
		_w3312_,
		_w3313_,
		_w3314_
	);
	LUT4 #(
		.INIT('h2a22)
	) name2355 (
		\u0_sp_csc_reg[2]/NET0131 ,
		_w1013_,
		_w2693_,
		_w2706_,
		_w3315_
	);
	LUT4 #(
		.INIT('h8000)
	) name2356 (
		\u0_spec_req_cs_reg[0]/NET0131 ,
		\u0_u0_csc_reg[2]/NET0131 ,
		wb_cyc_i_pad,
		wb_stb_i_pad,
		_w3316_
	);
	LUT3 #(
		.INIT('h40)
	) name2357 (
		\u0_spec_req_cs_reg[0]/NET0131 ,
		\u0_spec_req_cs_reg[1]/NET0131 ,
		\u0_u1_csc_reg[2]/NET0131 ,
		_w3317_
	);
	LUT2 #(
		.INIT('h8)
	) name2358 (
		_w1013_,
		_w3317_,
		_w3318_
	);
	LUT4 #(
		.INIT('h444f)
	) name2359 (
		_w2693_,
		_w2706_,
		_w3316_,
		_w3318_,
		_w3319_
	);
	LUT2 #(
		.INIT('hb)
	) name2360 (
		_w3315_,
		_w3319_,
		_w3320_
	);
	LUT4 #(
		.INIT('h2a22)
	) name2361 (
		\u0_sp_csc_reg[1]/NET0131 ,
		_w1013_,
		_w2693_,
		_w2706_,
		_w3321_
	);
	LUT4 #(
		.INIT('h8000)
	) name2362 (
		\u0_spec_req_cs_reg[0]/NET0131 ,
		\u0_u0_csc_reg[1]/NET0131 ,
		wb_cyc_i_pad,
		wb_stb_i_pad,
		_w3322_
	);
	LUT3 #(
		.INIT('h40)
	) name2363 (
		\u0_spec_req_cs_reg[0]/NET0131 ,
		\u0_spec_req_cs_reg[1]/NET0131 ,
		\u0_u1_csc_reg[1]/NET0131 ,
		_w3323_
	);
	LUT2 #(
		.INIT('h8)
	) name2364 (
		_w1013_,
		_w3323_,
		_w3324_
	);
	LUT4 #(
		.INIT('h444f)
	) name2365 (
		_w2693_,
		_w2706_,
		_w3322_,
		_w3324_,
		_w3325_
	);
	LUT2 #(
		.INIT('hb)
	) name2366 (
		_w3321_,
		_w3325_,
		_w3326_
	);
	LUT4 #(
		.INIT('h2a22)
	) name2367 (
		\u0_sp_csc_reg[3]/NET0131 ,
		_w1013_,
		_w2693_,
		_w2706_,
		_w3327_
	);
	LUT4 #(
		.INIT('h8000)
	) name2368 (
		\u0_spec_req_cs_reg[0]/NET0131 ,
		\u0_u0_csc_reg[3]/NET0131 ,
		wb_cyc_i_pad,
		wb_stb_i_pad,
		_w3328_
	);
	LUT3 #(
		.INIT('h40)
	) name2369 (
		\u0_spec_req_cs_reg[0]/NET0131 ,
		\u0_spec_req_cs_reg[1]/NET0131 ,
		\u0_u1_csc_reg[3]/NET0131 ,
		_w3329_
	);
	LUT2 #(
		.INIT('h8)
	) name2370 (
		_w1013_,
		_w3329_,
		_w3330_
	);
	LUT4 #(
		.INIT('h444f)
	) name2371 (
		_w2693_,
		_w2706_,
		_w3328_,
		_w3330_,
		_w3331_
	);
	LUT2 #(
		.INIT('hb)
	) name2372 (
		_w3327_,
		_w3331_,
		_w3332_
	);
	LUT3 #(
		.INIT('h57)
	) name2373 (
		_w1059_,
		_w1172_,
		_w1660_,
		_w3333_
	);
	LUT4 #(
		.INIT('h0700)
	) name2374 (
		_w1581_,
		_w1651_,
		_w1658_,
		_w3333_,
		_w3334_
	);
	LUT4 #(
		.INIT('h2300)
	) name2375 (
		_w1539_,
		_w1667_,
		_w2536_,
		_w3334_,
		_w3335_
	);
	LUT3 #(
		.INIT('h70)
	) name2376 (
		_w1059_,
		_w1083_,
		_w1901_,
		_w3336_
	);
	LUT4 #(
		.INIT('h7f00)
	) name2377 (
		_w1581_,
		_w1586_,
		_w1666_,
		_w3336_,
		_w3337_
	);
	LUT3 #(
		.INIT('h80)
	) name2378 (
		_w1591_,
		_w1908_,
		_w3337_,
		_w3338_
	);
	LUT3 #(
		.INIT('h01)
	) name2379 (
		\u5_timer_reg[2]/NET0131 ,
		\u5_timer_reg[3]/NET0131 ,
		\u5_timer_reg[4]/NET0131 ,
		_w3339_
	);
	LUT4 #(
		.INIT('h7000)
	) name2380 (
		_w1675_,
		_w1676_,
		_w1678_,
		_w3339_,
		_w3340_
	);
	LUT3 #(
		.INIT('h95)
	) name2381 (
		\u5_timer_reg[4]/NET0131 ,
		_w1674_,
		_w1679_,
		_w3341_
	);
	LUT2 #(
		.INIT('h2)
	) name2382 (
		_w3334_,
		_w3341_,
		_w3342_
	);
	LUT3 #(
		.INIT('hea)
	) name2383 (
		_w3335_,
		_w3338_,
		_w3342_,
		_w3343_
	);
	LUT3 #(
		.INIT('h80)
	) name2384 (
		_w1540_,
		_w1541_,
		_w2156_,
		_w3344_
	);
	LUT4 #(
		.INIT('h2030)
	) name2385 (
		_w1539_,
		_w1667_,
		_w3334_,
		_w3344_,
		_w3345_
	);
	LUT3 #(
		.INIT('h20)
	) name2386 (
		_w1675_,
		_w1676_,
		_w1678_,
		_w3346_
	);
	LUT3 #(
		.INIT('h0d)
	) name2387 (
		\u5_timer_reg[5]/NET0131 ,
		_w3340_,
		_w3346_,
		_w3347_
	);
	LUT2 #(
		.INIT('h2)
	) name2388 (
		_w3334_,
		_w3347_,
		_w3348_
	);
	LUT3 #(
		.INIT('hec)
	) name2389 (
		_w3338_,
		_w3345_,
		_w3348_,
		_w3349_
	);
	LUT3 #(
		.INIT('h80)
	) name2390 (
		_w1540_,
		_w1541_,
		_w3210_,
		_w3350_
	);
	LUT4 #(
		.INIT('h2030)
	) name2391 (
		_w1539_,
		_w1667_,
		_w3334_,
		_w3350_,
		_w3351_
	);
	LUT4 #(
		.INIT('ha2aa)
	) name2392 (
		\u5_timer_reg[6]/NET0131 ,
		_w1675_,
		_w1676_,
		_w1678_,
		_w3352_
	);
	LUT4 #(
		.INIT('h0001)
	) name2393 (
		\u5_mc_le_reg/NET0131 ,
		\u5_timer_reg[0]/NET0131 ,
		\u5_timer_reg[1]/NET0131 ,
		\u5_timer_reg[6]/NET0131 ,
		_w3353_
	);
	LUT3 #(
		.INIT('h20)
	) name2394 (
		_w1675_,
		_w1676_,
		_w3353_,
		_w3354_
	);
	LUT2 #(
		.INIT('h1)
	) name2395 (
		_w3352_,
		_w3354_,
		_w3355_
	);
	LUT2 #(
		.INIT('h2)
	) name2396 (
		_w3334_,
		_w3355_,
		_w3356_
	);
	LUT3 #(
		.INIT('hec)
	) name2397 (
		_w3338_,
		_w3351_,
		_w3356_,
		_w3357_
	);
	LUT3 #(
		.INIT('h80)
	) name2398 (
		_w1540_,
		_w1541_,
		_w3219_,
		_w3358_
	);
	LUT4 #(
		.INIT('h2030)
	) name2399 (
		_w1539_,
		_w1667_,
		_w3334_,
		_w3358_,
		_w3359_
	);
	LUT3 #(
		.INIT('h2a)
	) name2400 (
		\u5_timer_reg[7]/NET0131 ,
		_w1675_,
		_w3353_,
		_w3360_
	);
	LUT2 #(
		.INIT('h8)
	) name2401 (
		_w3334_,
		_w3360_,
		_w3361_
	);
	LUT3 #(
		.INIT('hec)
	) name2402 (
		_w3338_,
		_w3359_,
		_w3361_,
		_w3362_
	);
	LUT4 #(
		.INIT('h2a22)
	) name2403 (
		\u0_csc_reg[11]/NET0131 ,
		_w1013_,
		_w2693_,
		_w2706_,
		_w3363_
	);
	LUT3 #(
		.INIT('h2a)
	) name2404 (
		\u0_u0_csc_reg[11]/P0001 ,
		\u0_u0_csc_reg[8]/P0001 ,
		wb_we_i_pad,
		_w3364_
	);
	LUT4 #(
		.INIT('h0100)
	) name2405 (
		_w2914_,
		_w2915_,
		_w2916_,
		_w3364_,
		_w3365_
	);
	LUT3 #(
		.INIT('h80)
	) name2406 (
		_w2907_,
		_w2912_,
		_w3365_,
		_w3366_
	);
	LUT4 #(
		.INIT('h00df)
	) name2407 (
		\u0_u1_csc_reg[11]/P0001 ,
		_w2918_,
		_w2930_,
		_w3366_,
		_w3367_
	);
	LUT2 #(
		.INIT('h2)
	) name2408 (
		_w1013_,
		_w3367_,
		_w3368_
	);
	LUT3 #(
		.INIT('hb0)
	) name2409 (
		_w2693_,
		_w2706_,
		_w3368_,
		_w3369_
	);
	LUT2 #(
		.INIT('he)
	) name2410 (
		_w3363_,
		_w3369_,
		_w3370_
	);
	LUT3 #(
		.INIT('h2a)
	) name2411 (
		\wb_addr_i[15]_pad ,
		_w976_,
		_w1975_,
		_w3371_
	);
	LUT3 #(
		.INIT('h10)
	) name2412 (
		_w1972_,
		_w1974_,
		_w3371_,
		_w3372_
	);
	LUT3 #(
		.INIT('h2a)
	) name2413 (
		\wb_addr_i[14]_pad ,
		_w976_,
		_w1971_,
		_w3373_
	);
	LUT3 #(
		.INIT('h40)
	) name2414 (
		_w1970_,
		_w1976_,
		_w3373_,
		_w3374_
	);
	LUT3 #(
		.INIT('h10)
	) name2415 (
		_w1970_,
		_w1976_,
		_w2631_,
		_w3375_
	);
	LUT4 #(
		.INIT('habef)
	) name2416 (
		_w1970_,
		_w1976_,
		_w2631_,
		_w3373_,
		_w3376_
	);
	LUT3 #(
		.INIT('h45)
	) name2417 (
		_w2424_,
		_w3372_,
		_w3376_,
		_w3377_
	);
	LUT4 #(
		.INIT('h6c00)
	) name2418 (
		\u1_acs_addr_reg[13]/P0001 ,
		\u1_acs_addr_reg[14]/P0001 ,
		_w2419_,
		_w2424_,
		_w3378_
	);
	LUT2 #(
		.INIT('he)
	) name2419 (
		_w3377_,
		_w3378_,
		_w3379_
	);
	LUT3 #(
		.INIT('h80)
	) name2420 (
		_w1572_,
		_w1581_,
		_w1586_,
		_w3380_
	);
	LUT2 #(
		.INIT('h4)
	) name2421 (
		_w1095_,
		_w1215_,
		_w3381_
	);
	LUT4 #(
		.INIT('h00a8)
	) name2422 (
		_w991_,
		_w1077_,
		_w1250_,
		_w1566_,
		_w3382_
	);
	LUT3 #(
		.INIT('h70)
	) name2423 (
		_w991_,
		_w1250_,
		_w1571_,
		_w3383_
	);
	LUT3 #(
		.INIT('h31)
	) name2424 (
		_w1190_,
		_w3382_,
		_w3383_,
		_w3384_
	);
	LUT3 #(
		.INIT('h40)
	) name2425 (
		_w3380_,
		_w3381_,
		_w3384_,
		_w3385_
	);
	LUT3 #(
		.INIT('h80)
	) name2426 (
		\u5_wb_wait_r_reg/P0001 ,
		_w1100_,
		_w1161_,
		_w3386_
	);
	LUT2 #(
		.INIT('h1)
	) name2427 (
		_w1624_,
		_w3386_,
		_w3387_
	);
	LUT4 #(
		.INIT('h8000)
	) name2428 (
		_w1067_,
		_w1298_,
		_w1316_,
		_w3387_,
		_w3388_
	);
	LUT4 #(
		.INIT('h4000)
	) name2429 (
		_w1051_,
		_w2487_,
		_w2493_,
		_w3388_,
		_w3389_
	);
	LUT4 #(
		.INIT('hbfff)
	) name2430 (
		_w1051_,
		_w2487_,
		_w2493_,
		_w3388_,
		_w3390_
	);
	LUT3 #(
		.INIT('h8b)
	) name2431 (
		\u5_cmd_del_reg[2]/NET0131 ,
		\u5_wr_cycle_reg/NET0131 ,
		_w3389_,
		_w3391_
	);
	LUT3 #(
		.INIT('h2a)
	) name2432 (
		\wb_addr_i[22]_pad ,
		_w976_,
		_w1975_,
		_w3392_
	);
	LUT3 #(
		.INIT('h10)
	) name2433 (
		_w1972_,
		_w1974_,
		_w3392_,
		_w3393_
	);
	LUT3 #(
		.INIT('h40)
	) name2434 (
		_w1970_,
		_w1976_,
		_w2501_,
		_w3394_
	);
	LUT3 #(
		.INIT('h10)
	) name2435 (
		_w1970_,
		_w1976_,
		_w2430_,
		_w3395_
	);
	LUT4 #(
		.INIT('habef)
	) name2436 (
		_w1970_,
		_w1976_,
		_w2430_,
		_w2501_,
		_w3396_
	);
	LUT3 #(
		.INIT('h45)
	) name2437 (
		_w2424_,
		_w3393_,
		_w3396_,
		_w3397_
	);
	LUT2 #(
		.INIT('h8)
	) name2438 (
		\u1_acs_addr_reg[19]/P0001 ,
		\u1_acs_addr_reg[20]/P0001 ,
		_w3398_
	);
	LUT4 #(
		.INIT('h8000)
	) name2439 (
		_w2419_,
		_w2420_,
		_w2421_,
		_w3398_,
		_w3399_
	);
	LUT4 #(
		.INIT('h3020)
	) name2440 (
		\u1_acs_addr_reg[21]/P0001 ,
		_w2423_,
		_w2424_,
		_w3399_,
		_w3400_
	);
	LUT2 #(
		.INIT('he)
	) name2441 (
		_w3397_,
		_w3400_,
		_w3401_
	);
	LUT3 #(
		.INIT('h0e)
	) name2442 (
		\u4_rfr_clr_reg/P0001 ,
		\u4_rfr_req_reg/NET0131 ,
		\u5_rfr_ack_r_reg/NET0131 ,
		_w3402_
	);
	LUT3 #(
		.INIT('h2a)
	) name2443 (
		\wb_addr_i[14]_pad ,
		_w976_,
		_w1975_,
		_w3403_
	);
	LUT3 #(
		.INIT('h10)
	) name2444 (
		_w1972_,
		_w1974_,
		_w3403_,
		_w3404_
	);
	LUT3 #(
		.INIT('h2a)
	) name2445 (
		\wb_addr_i[13]_pad ,
		_w976_,
		_w1971_,
		_w3405_
	);
	LUT3 #(
		.INIT('h40)
	) name2446 (
		_w1970_,
		_w1976_,
		_w3405_,
		_w3406_
	);
	LUT3 #(
		.INIT('h10)
	) name2447 (
		_w1970_,
		_w1976_,
		_w3229_,
		_w3407_
	);
	LUT4 #(
		.INIT('habef)
	) name2448 (
		_w1970_,
		_w1976_,
		_w3229_,
		_w3405_,
		_w3408_
	);
	LUT3 #(
		.INIT('h45)
	) name2449 (
		_w2424_,
		_w3404_,
		_w3408_,
		_w3409_
	);
	LUT3 #(
		.INIT('h9f)
	) name2450 (
		\u1_acs_addr_reg[13]/P0001 ,
		_w2419_,
		_w2424_,
		_w3410_
	);
	LUT2 #(
		.INIT('hb)
	) name2451 (
		_w3409_,
		_w3410_,
		_w3411_
	);
	LUT2 #(
		.INIT('h4)
	) name2452 (
		\u1_u0_out_r_reg[11]/P0001 ,
		\u5_tmr2_done_reg/NET0131 ,
		_w3412_
	);
	LUT4 #(
		.INIT('h7500)
	) name2453 (
		_w964_,
		_w1974_,
		_w2417_,
		_w3412_,
		_w3413_
	);
	LUT2 #(
		.INIT('h1)
	) name2454 (
		\u1_acs_addr_reg[11]/P0001 ,
		\u5_tmr2_done_reg/NET0131 ,
		_w3414_
	);
	LUT3 #(
		.INIT('h01)
	) name2455 (
		\u1_acs_addr_reg[11]/P0001 ,
		\u5_state_reg[42]/NET0131 ,
		\u5_state_reg[44]/NET0131 ,
		_w3415_
	);
	LUT4 #(
		.INIT('h040f)
	) name2456 (
		_w1974_,
		_w2417_,
		_w3414_,
		_w3415_,
		_w3416_
	);
	LUT3 #(
		.INIT('h20)
	) name2457 (
		_w2424_,
		_w3413_,
		_w3416_,
		_w3417_
	);
	LUT3 #(
		.INIT('h10)
	) name2458 (
		_w1970_,
		_w1976_,
		_w3405_,
		_w3418_
	);
	LUT3 #(
		.INIT('h2a)
	) name2459 (
		\wb_addr_i[11]_pad ,
		_w976_,
		_w1971_,
		_w3419_
	);
	LUT3 #(
		.INIT('h40)
	) name2460 (
		_w1970_,
		_w1976_,
		_w3419_,
		_w3420_
	);
	LUT3 #(
		.INIT('h2a)
	) name2461 (
		\wb_addr_i[12]_pad ,
		_w976_,
		_w1975_,
		_w3421_
	);
	LUT3 #(
		.INIT('h10)
	) name2462 (
		_w1972_,
		_w1974_,
		_w3421_,
		_w3422_
	);
	LUT4 #(
		.INIT('h5554)
	) name2463 (
		_w2424_,
		_w3418_,
		_w3420_,
		_w3422_,
		_w3423_
	);
	LUT2 #(
		.INIT('he)
	) name2464 (
		_w3417_,
		_w3423_,
		_w3424_
	);
	LUT3 #(
		.INIT('h2a)
	) name2465 (
		\wb_addr_i[18]_pad ,
		_w976_,
		_w1975_,
		_w3425_
	);
	LUT3 #(
		.INIT('h10)
	) name2466 (
		_w1972_,
		_w1974_,
		_w3425_,
		_w3426_
	);
	LUT3 #(
		.INIT('h40)
	) name2467 (
		_w1970_,
		_w1976_,
		_w3231_,
		_w3427_
	);
	LUT3 #(
		.INIT('h10)
	) name2468 (
		_w1970_,
		_w1976_,
		_w2505_,
		_w3428_
	);
	LUT4 #(
		.INIT('habef)
	) name2469 (
		_w1970_,
		_w1976_,
		_w2505_,
		_w3231_,
		_w3429_
	);
	LUT3 #(
		.INIT('h45)
	) name2470 (
		_w2424_,
		_w3426_,
		_w3429_,
		_w3430_
	);
	LUT4 #(
		.INIT('h1333)
	) name2471 (
		\u1_acs_addr_reg[16]/P0001 ,
		\u1_acs_addr_reg[17]/P0001 ,
		_w2419_,
		_w2420_,
		_w3431_
	);
	LUT4 #(
		.INIT('h70f0)
	) name2472 (
		_w2419_,
		_w2420_,
		_w2424_,
		_w2657_,
		_w3432_
	);
	LUT3 #(
		.INIT('hba)
	) name2473 (
		_w3430_,
		_w3431_,
		_w3432_,
		_w3433_
	);
	LUT3 #(
		.INIT('h80)
	) name2474 (
		_w1582_,
		_w1584_,
		_w2022_,
		_w3434_
	);
	LUT4 #(
		.INIT('h4f00)
	) name2475 (
		_w1533_,
		_w1579_,
		_w1580_,
		_w3434_,
		_w3435_
	);
	LUT2 #(
		.INIT('h2)
	) name2476 (
		_w1186_,
		_w3435_,
		_w3436_
	);
	LUT3 #(
		.INIT('h08)
	) name2477 (
		_w1310_,
		_w2491_,
		_w3436_,
		_w3437_
	);
	LUT4 #(
		.INIT('h1000)
	) name2478 (
		_w1071_,
		_w1196_,
		_w1202_,
		_w1299_,
		_w3438_
	);
	LUT3 #(
		.INIT('h80)
	) name2479 (
		\u7_mc_br_r_reg/P0001 ,
		_w1041_,
		_w1256_,
		_w3439_
	);
	LUT4 #(
		.INIT('h0040)
	) name2480 (
		_w1051_,
		_w1625_,
		_w2485_,
		_w3439_,
		_w3440_
	);
	LUT4 #(
		.INIT('h8000)
	) name2481 (
		_w1254_,
		_w2489_,
		_w3438_,
		_w3440_,
		_w3441_
	);
	LUT4 #(
		.INIT('h7fff)
	) name2482 (
		_w2484_,
		_w2487_,
		_w3437_,
		_w3441_,
		_w3442_
	);
	LUT3 #(
		.INIT('h2a)
	) name2483 (
		\wb_addr_i[7]_pad ,
		_w976_,
		_w1971_,
		_w3443_
	);
	LUT3 #(
		.INIT('h40)
	) name2484 (
		_w1970_,
		_w1976_,
		_w3443_,
		_w3444_
	);
	LUT3 #(
		.INIT('h2a)
	) name2485 (
		\wb_addr_i[8]_pad ,
		_w976_,
		_w1975_,
		_w3445_
	);
	LUT3 #(
		.INIT('h10)
	) name2486 (
		_w1972_,
		_w1974_,
		_w3445_,
		_w3446_
	);
	LUT3 #(
		.INIT('h2a)
	) name2487 (
		\wb_addr_i[9]_pad ,
		_w976_,
		_w1971_,
		_w3447_
	);
	LUT3 #(
		.INIT('h10)
	) name2488 (
		_w1970_,
		_w1976_,
		_w3447_,
		_w3448_
	);
	LUT4 #(
		.INIT('h5554)
	) name2489 (
		_w2424_,
		_w3444_,
		_w3446_,
		_w3448_,
		_w3449_
	);
	LUT2 #(
		.INIT('h4)
	) name2490 (
		\u1_u0_out_r_reg[7]/P0001 ,
		\u5_tmr2_done_reg/NET0131 ,
		_w3450_
	);
	LUT4 #(
		.INIT('h7500)
	) name2491 (
		_w964_,
		_w1974_,
		_w2417_,
		_w3450_,
		_w3451_
	);
	LUT2 #(
		.INIT('h1)
	) name2492 (
		\u1_acs_addr_reg[7]/P0001 ,
		\u5_tmr2_done_reg/NET0131 ,
		_w3452_
	);
	LUT3 #(
		.INIT('h01)
	) name2493 (
		\u1_acs_addr_reg[7]/P0001 ,
		\u5_state_reg[42]/NET0131 ,
		\u5_state_reg[44]/NET0131 ,
		_w3453_
	);
	LUT4 #(
		.INIT('h040f)
	) name2494 (
		_w1974_,
		_w2417_,
		_w3452_,
		_w3453_,
		_w3454_
	);
	LUT3 #(
		.INIT('h20)
	) name2495 (
		_w2424_,
		_w3451_,
		_w3454_,
		_w3455_
	);
	LUT2 #(
		.INIT('he)
	) name2496 (
		_w3449_,
		_w3455_,
		_w3456_
	);
	LUT2 #(
		.INIT('h4)
	) name2497 (
		\u5_state_reg[1]/NET0131 ,
		\u5_wr_cycle_reg/NET0131 ,
		_w3457_
	);
	LUT2 #(
		.INIT('h1)
	) name2498 (
		_w1564_,
		_w1733_,
		_w3458_
	);
	LUT4 #(
		.INIT('h00a8)
	) name2499 (
		_w1100_,
		_w1108_,
		_w1110_,
		_w3458_,
		_w3459_
	);
	LUT3 #(
		.INIT('h08)
	) name2500 (
		_w1339_,
		_w2019_,
		_w3458_,
		_w3460_
	);
	LUT4 #(
		.INIT('h070f)
	) name2501 (
		_w1581_,
		_w1586_,
		_w3459_,
		_w3460_,
		_w3461_
	);
	LUT2 #(
		.INIT('hb)
	) name2502 (
		_w3457_,
		_w3461_,
		_w3462_
	);
	LUT4 #(
		.INIT('h0501)
	) name2503 (
		\u0_csr_r_reg[10]/NET0131 ,
		\u0_csr_r_reg[8]/NET0131 ,
		\u0_csr_r_reg[9]/NET0131 ,
		\u4_rfr_cnt_reg[1]/NET0131 ,
		_w3463_
	);
	LUT3 #(
		.INIT('h51)
	) name2504 (
		\u0_csr_r_reg[10]/NET0131 ,
		\u0_csr_r_reg[8]/NET0131 ,
		\u4_rfr_cnt_reg[3]/NET0131 ,
		_w3464_
	);
	LUT2 #(
		.INIT('h8)
	) name2505 (
		\u4_rfr_cnt_reg[1]/NET0131 ,
		\u4_rfr_cnt_reg[2]/NET0131 ,
		_w3465_
	);
	LUT2 #(
		.INIT('h8)
	) name2506 (
		_w3464_,
		_w3465_,
		_w3466_
	);
	LUT3 #(
		.INIT('h31)
	) name2507 (
		\u0_csr_r_reg[8]/NET0131 ,
		\u0_csr_r_reg[9]/NET0131 ,
		\u4_rfr_cnt_reg[5]/NET0131 ,
		_w3467_
	);
	LUT4 #(
		.INIT('hc040)
	) name2508 (
		\u0_csr_r_reg[8]/NET0131 ,
		\u4_rfr_cnt_reg[5]/NET0131 ,
		\u4_rfr_cnt_reg[6]/NET0131 ,
		\u4_rfr_cnt_reg[7]/NET0131 ,
		_w3468_
	);
	LUT2 #(
		.INIT('h8)
	) name2509 (
		\u4_rfr_cnt_reg[3]/NET0131 ,
		\u4_rfr_cnt_reg[4]/NET0131 ,
		_w3469_
	);
	LUT4 #(
		.INIT('h8000)
	) name2510 (
		\u4_rfr_cnt_reg[1]/NET0131 ,
		\u4_rfr_cnt_reg[2]/NET0131 ,
		\u4_rfr_cnt_reg[3]/NET0131 ,
		\u4_rfr_cnt_reg[4]/NET0131 ,
		_w3470_
	);
	LUT3 #(
		.INIT('he0)
	) name2511 (
		_w3467_,
		_w3468_,
		_w3470_,
		_w3471_
	);
	LUT2 #(
		.INIT('h8)
	) name2512 (
		\u4_rfr_cnt_reg[0]/NET0131 ,
		\u4_rfr_early_reg/NET0131 ,
		_w3472_
	);
	LUT4 #(
		.INIT('hfe00)
	) name2513 (
		_w3463_,
		_w3466_,
		_w3471_,
		_w3472_,
		_w3473_
	);
	LUT3 #(
		.INIT('h2a)
	) name2514 (
		\wb_addr_i[13]_pad ,
		_w976_,
		_w1975_,
		_w3474_
	);
	LUT3 #(
		.INIT('h10)
	) name2515 (
		_w1972_,
		_w1974_,
		_w3474_,
		_w3475_
	);
	LUT3 #(
		.INIT('h2a)
	) name2516 (
		\wb_addr_i[12]_pad ,
		_w976_,
		_w1971_,
		_w3476_
	);
	LUT3 #(
		.INIT('h40)
	) name2517 (
		_w1970_,
		_w1976_,
		_w3476_,
		_w3477_
	);
	LUT3 #(
		.INIT('h10)
	) name2518 (
		_w1970_,
		_w1976_,
		_w3373_,
		_w3478_
	);
	LUT4 #(
		.INIT('habef)
	) name2519 (
		_w1970_,
		_w1976_,
		_w3373_,
		_w3476_,
		_w3479_
	);
	LUT3 #(
		.INIT('h45)
	) name2520 (
		_w2424_,
		_w3475_,
		_w3479_,
		_w3480_
	);
	LUT2 #(
		.INIT('h8)
	) name2521 (
		\u1_u0_out_r_reg[12]/P0001 ,
		\u5_tmr2_done_reg/NET0131 ,
		_w3481_
	);
	LUT4 #(
		.INIT('h7500)
	) name2522 (
		_w964_,
		_w1974_,
		_w2417_,
		_w3481_,
		_w3482_
	);
	LUT4 #(
		.INIT('h3020)
	) name2523 (
		\u1_acs_addr_reg[12]/P0001 ,
		_w2419_,
		_w2424_,
		_w3482_,
		_w3483_
	);
	LUT2 #(
		.INIT('he)
	) name2524 (
		_w3480_,
		_w3483_,
		_w3484_
	);
	LUT2 #(
		.INIT('h1)
	) name2525 (
		\u5_ack_cnt_reg[0]/NET0131 ,
		\u5_no_wb_cycle_reg/NET0131 ,
		_w3485_
	);
	LUT3 #(
		.INIT('hb0)
	) name2526 (
		_w1568_,
		_w1737_,
		_w3485_,
		_w3486_
	);
	LUT2 #(
		.INIT('h2)
	) name2527 (
		\u5_ack_cnt_reg[0]/NET0131 ,
		\u5_no_wb_cycle_reg/NET0131 ,
		_w3487_
	);
	LUT3 #(
		.INIT('h40)
	) name2528 (
		_w1568_,
		_w1737_,
		_w3487_,
		_w3488_
	);
	LUT4 #(
		.INIT('h111f)
	) name2529 (
		_w998_,
		_w1010_,
		_w3486_,
		_w3488_,
		_w3489_
	);
	LUT3 #(
		.INIT('hb0)
	) name2530 (
		_w1568_,
		_w1737_,
		_w3487_,
		_w3490_
	);
	LUT3 #(
		.INIT('h40)
	) name2531 (
		_w1568_,
		_w1737_,
		_w3485_,
		_w3491_
	);
	LUT4 #(
		.INIT('heeef)
	) name2532 (
		_w998_,
		_w1010_,
		_w3490_,
		_w3491_,
		_w3492_
	);
	LUT2 #(
		.INIT('h7)
	) name2533 (
		_w3489_,
		_w3492_,
		_w3493_
	);
	LUT4 #(
		.INIT('h5455)
	) name2534 (
		\u5_ack_cnt_reg[0]/NET0131 ,
		_w998_,
		_w1010_,
		_w1738_,
		_w3494_
	);
	LUT2 #(
		.INIT('h6)
	) name2535 (
		\u5_ack_cnt_reg[0]/NET0131 ,
		\u5_ack_cnt_reg[1]/NET0131 ,
		_w3495_
	);
	LUT4 #(
		.INIT('hf100)
	) name2536 (
		_w998_,
		_w1010_,
		_w1738_,
		_w3495_,
		_w3496_
	);
	LUT2 #(
		.INIT('h4)
	) name2537 (
		_w3494_,
		_w3496_,
		_w3497_
	);
	LUT4 #(
		.INIT('h000e)
	) name2538 (
		_w998_,
		_w1010_,
		_w1738_,
		_w3495_,
		_w3498_
	);
	LUT4 #(
		.INIT('hef00)
	) name2539 (
		_w998_,
		_w1010_,
		_w1738_,
		_w1734_,
		_w3499_
	);
	LUT3 #(
		.INIT('h01)
	) name2540 (
		\u5_no_wb_cycle_reg/NET0131 ,
		_w3498_,
		_w3499_,
		_w3500_
	);
	LUT2 #(
		.INIT('h4)
	) name2541 (
		_w3497_,
		_w3500_,
		_w3501_
	);
	LUT3 #(
		.INIT('h40)
	) name2542 (
		_w1568_,
		_w1734_,
		_w1737_,
		_w3502_
	);
	LUT4 #(
		.INIT('ha8aa)
	) name2543 (
		\u5_ack_cnt_reg[2]/NET0131 ,
		_w998_,
		_w1010_,
		_w3502_,
		_w3503_
	);
	LUT3 #(
		.INIT('h01)
	) name2544 (
		\u5_ack_cnt_reg[0]/NET0131 ,
		\u5_ack_cnt_reg[1]/NET0131 ,
		\u5_ack_cnt_reg[2]/NET0131 ,
		_w3504_
	);
	LUT3 #(
		.INIT('h40)
	) name2545 (
		_w1568_,
		_w1737_,
		_w3504_,
		_w3505_
	);
	LUT4 #(
		.INIT('he1f1)
	) name2546 (
		_w998_,
		_w1010_,
		_w1738_,
		_w3504_,
		_w3506_
	);
	LUT3 #(
		.INIT('h78)
	) name2547 (
		\u5_ack_cnt_reg[0]/NET0131 ,
		\u5_ack_cnt_reg[1]/NET0131 ,
		\u5_ack_cnt_reg[2]/NET0131 ,
		_w3507_
	);
	LUT3 #(
		.INIT('h0b)
	) name2548 (
		_w1568_,
		_w1737_,
		_w3507_,
		_w3508_
	);
	LUT4 #(
		.INIT('h0155)
	) name2549 (
		\u5_no_wb_cycle_reg/NET0131 ,
		_w998_,
		_w1010_,
		_w3508_,
		_w3509_
	);
	LUT3 #(
		.INIT('hb0)
	) name2550 (
		_w3503_,
		_w3506_,
		_w3509_,
		_w3510_
	);
	LUT4 #(
		.INIT('ha8aa)
	) name2551 (
		\u5_ack_cnt_reg[3]/NET0131 ,
		_w998_,
		_w1010_,
		_w3505_,
		_w3511_
	);
	LUT4 #(
		.INIT('hef11)
	) name2552 (
		_w998_,
		_w1010_,
		_w1735_,
		_w1738_,
		_w3512_
	);
	LUT4 #(
		.INIT('h807f)
	) name2553 (
		\u5_ack_cnt_reg[0]/NET0131 ,
		\u5_ack_cnt_reg[1]/NET0131 ,
		\u5_ack_cnt_reg[2]/NET0131 ,
		\u5_ack_cnt_reg[3]/NET0131 ,
		_w3513_
	);
	LUT3 #(
		.INIT('hb0)
	) name2554 (
		_w1568_,
		_w1737_,
		_w3513_,
		_w3514_
	);
	LUT4 #(
		.INIT('h0155)
	) name2555 (
		\u5_no_wb_cycle_reg/NET0131 ,
		_w998_,
		_w1010_,
		_w3514_,
		_w3515_
	);
	LUT3 #(
		.INIT('hb0)
	) name2556 (
		_w3511_,
		_w3512_,
		_w3515_,
		_w3516_
	);
	LUT3 #(
		.INIT('h2a)
	) name2557 (
		\wb_addr_i[4]_pad ,
		_w976_,
		_w1971_,
		_w3517_
	);
	LUT3 #(
		.INIT('h40)
	) name2558 (
		_w1970_,
		_w1976_,
		_w3517_,
		_w3518_
	);
	LUT3 #(
		.INIT('h2a)
	) name2559 (
		\wb_addr_i[5]_pad ,
		_w976_,
		_w1975_,
		_w3519_
	);
	LUT3 #(
		.INIT('h10)
	) name2560 (
		_w1972_,
		_w1974_,
		_w3519_,
		_w3520_
	);
	LUT3 #(
		.INIT('h2a)
	) name2561 (
		\wb_addr_i[6]_pad ,
		_w976_,
		_w1971_,
		_w3521_
	);
	LUT3 #(
		.INIT('h10)
	) name2562 (
		_w1970_,
		_w1976_,
		_w3521_,
		_w3522_
	);
	LUT4 #(
		.INIT('h5554)
	) name2563 (
		_w2424_,
		_w3518_,
		_w3520_,
		_w3522_,
		_w3523_
	);
	LUT2 #(
		.INIT('h4)
	) name2564 (
		\u1_u0_out_r_reg[4]/P0001 ,
		\u5_tmr2_done_reg/NET0131 ,
		_w3524_
	);
	LUT4 #(
		.INIT('h7500)
	) name2565 (
		_w964_,
		_w1974_,
		_w2417_,
		_w3524_,
		_w3525_
	);
	LUT2 #(
		.INIT('h1)
	) name2566 (
		\u1_acs_addr_reg[4]/P0001 ,
		\u5_tmr2_done_reg/NET0131 ,
		_w3526_
	);
	LUT3 #(
		.INIT('h01)
	) name2567 (
		\u1_acs_addr_reg[4]/P0001 ,
		\u5_state_reg[42]/NET0131 ,
		\u5_state_reg[44]/NET0131 ,
		_w3527_
	);
	LUT4 #(
		.INIT('h040f)
	) name2568 (
		_w1974_,
		_w2417_,
		_w3526_,
		_w3527_,
		_w3528_
	);
	LUT3 #(
		.INIT('h20)
	) name2569 (
		_w2424_,
		_w3525_,
		_w3528_,
		_w3529_
	);
	LUT2 #(
		.INIT('he)
	) name2570 (
		_w3523_,
		_w3529_,
		_w3530_
	);
	LUT2 #(
		.INIT('h4)
	) name2571 (
		\u1_u0_out_r_reg[8]/P0001 ,
		\u5_tmr2_done_reg/NET0131 ,
		_w3531_
	);
	LUT4 #(
		.INIT('h7500)
	) name2572 (
		_w964_,
		_w1974_,
		_w2417_,
		_w3531_,
		_w3532_
	);
	LUT2 #(
		.INIT('h1)
	) name2573 (
		\u1_acs_addr_reg[8]/P0001 ,
		\u5_tmr2_done_reg/NET0131 ,
		_w3533_
	);
	LUT3 #(
		.INIT('h01)
	) name2574 (
		\u1_acs_addr_reg[8]/P0001 ,
		\u5_state_reg[42]/NET0131 ,
		\u5_state_reg[44]/NET0131 ,
		_w3534_
	);
	LUT4 #(
		.INIT('h040f)
	) name2575 (
		_w1974_,
		_w2417_,
		_w3533_,
		_w3534_,
		_w3535_
	);
	LUT3 #(
		.INIT('h20)
	) name2576 (
		_w2424_,
		_w3532_,
		_w3535_,
		_w3536_
	);
	LUT3 #(
		.INIT('h2a)
	) name2577 (
		\wb_addr_i[8]_pad ,
		_w976_,
		_w1971_,
		_w3537_
	);
	LUT3 #(
		.INIT('h40)
	) name2578 (
		_w1970_,
		_w1976_,
		_w3537_,
		_w3538_
	);
	LUT3 #(
		.INIT('h2a)
	) name2579 (
		\wb_addr_i[9]_pad ,
		_w976_,
		_w1975_,
		_w3539_
	);
	LUT3 #(
		.INIT('h10)
	) name2580 (
		_w1972_,
		_w1974_,
		_w3539_,
		_w3540_
	);
	LUT3 #(
		.INIT('h2a)
	) name2581 (
		\wb_addr_i[10]_pad ,
		_w976_,
		_w1971_,
		_w3541_
	);
	LUT3 #(
		.INIT('h10)
	) name2582 (
		_w1970_,
		_w1976_,
		_w3541_,
		_w3542_
	);
	LUT4 #(
		.INIT('h5554)
	) name2583 (
		_w2424_,
		_w3538_,
		_w3540_,
		_w3542_,
		_w3543_
	);
	LUT2 #(
		.INIT('he)
	) name2584 (
		_w3536_,
		_w3543_,
		_w3544_
	);
	LUT3 #(
		.INIT('ha8)
	) name2585 (
		_w1969_,
		_w2553_,
		_w2652_,
		_w3545_
	);
	LUT2 #(
		.INIT('h1)
	) name2586 (
		_w1966_,
		_w1968_,
		_w3546_
	);
	LUT2 #(
		.INIT('h2)
	) name2587 (
		_w3428_,
		_w3546_,
		_w3547_
	);
	LUT2 #(
		.INIT('h2)
	) name2588 (
		_w1966_,
		_w1968_,
		_w3548_
	);
	LUT2 #(
		.INIT('h4)
	) name2589 (
		_w1966_,
		_w1968_,
		_w3549_
	);
	LUT2 #(
		.INIT('h9)
	) name2590 (
		_w1966_,
		_w1968_,
		_w3550_
	);
	LUT3 #(
		.INIT('h02)
	) name2591 (
		\u0_csc_reg[9]/NET0131 ,
		\u5_lmr_ack_reg/NET0131 ,
		\u5_state_reg[26]/NET0131 ,
		_w3551_
	);
	LUT4 #(
		.INIT('h11d5)
	) name2592 (
		\u0_sp_csc_reg[9]/NET0131 ,
		_w976_,
		_w1114_,
		_w3551_,
		_w3552_
	);
	LUT4 #(
		.INIT('h00f1)
	) name2593 (
		_w2504_,
		_w3394_,
		_w3550_,
		_w3552_,
		_w3553_
	);
	LUT3 #(
		.INIT('h10)
	) name2594 (
		_w3545_,
		_w3547_,
		_w3553_,
		_w3554_
	);
	LUT3 #(
		.INIT('h2a)
	) name2595 (
		\wb_addr_i[22]_pad ,
		_w976_,
		_w1965_,
		_w3555_
	);
	LUT3 #(
		.INIT('h40)
	) name2596 (
		_w1964_,
		_w1968_,
		_w3555_,
		_w3556_
	);
	LUT4 #(
		.INIT('h33f7)
	) name2597 (
		\wb_addr_i[23]_pad ,
		_w1995_,
		_w3550_,
		_w3556_,
		_w3557_
	);
	LUT2 #(
		.INIT('h8)
	) name2598 (
		_w1969_,
		_w2551_,
		_w3558_
	);
	LUT3 #(
		.INIT('h0e)
	) name2599 (
		_w2502_,
		_w3393_,
		_w3550_,
		_w3559_
	);
	LUT3 #(
		.INIT('h70)
	) name2600 (
		_w1969_,
		_w2502_,
		_w3552_,
		_w3560_
	);
	LUT4 #(
		.INIT('h0200)
	) name2601 (
		_w3557_,
		_w3558_,
		_w3559_,
		_w3560_,
		_w3561_
	);
	LUT2 #(
		.INIT('h1)
	) name2602 (
		_w3554_,
		_w3561_,
		_w3562_
	);
	LUT4 #(
		.INIT('h8000)
	) name2603 (
		\u1_acs_addr_reg[0]/P0001 ,
		\u1_acs_addr_reg[1]/P0001 ,
		\u1_acs_addr_reg[2]/P0001 ,
		\u1_acs_addr_reg[3]/P0001 ,
		_w3563_
	);
	LUT3 #(
		.INIT('h80)
	) name2604 (
		\u1_acs_addr_reg[4]/P0001 ,
		\u1_acs_addr_reg[5]/P0001 ,
		\u1_acs_addr_reg[6]/P0001 ,
		_w3564_
	);
	LUT3 #(
		.INIT('h80)
	) name2605 (
		\u1_acs_addr_reg[7]/P0001 ,
		\u1_acs_addr_reg[8]/P0001 ,
		\u1_acs_addr_reg[9]/P0001 ,
		_w3565_
	);
	LUT3 #(
		.INIT('h80)
	) name2606 (
		_w3563_,
		_w3564_,
		_w3565_,
		_w3566_
	);
	LUT2 #(
		.INIT('h8)
	) name2607 (
		\u1_acs_addr_reg[10]/P0001 ,
		\u1_acs_addr_reg[11]/P0001 ,
		_w3567_
	);
	LUT4 #(
		.INIT('h8000)
	) name2608 (
		_w3563_,
		_w3564_,
		_w3565_,
		_w3567_,
		_w3568_
	);
	LUT3 #(
		.INIT('h6c)
	) name2609 (
		\u1_acs_addr_reg[10]/P0001 ,
		\u1_acs_addr_reg[11]/P0001 ,
		_w3566_,
		_w3569_
	);
	LUT3 #(
		.INIT('h2a)
	) name2610 (
		\wb_addr_i[10]_pad ,
		_w976_,
		_w1975_,
		_w3570_
	);
	LUT3 #(
		.INIT('h10)
	) name2611 (
		_w1972_,
		_w1974_,
		_w3570_,
		_w3571_
	);
	LUT3 #(
		.INIT('ha8)
	) name2612 (
		_w1969_,
		_w3420_,
		_w3571_,
		_w3572_
	);
	LUT2 #(
		.INIT('h2)
	) name2613 (
		_w3542_,
		_w3546_,
		_w3573_
	);
	LUT3 #(
		.INIT('h2a)
	) name2614 (
		\wb_addr_i[11]_pad ,
		_w976_,
		_w1975_,
		_w3574_
	);
	LUT3 #(
		.INIT('h10)
	) name2615 (
		_w1972_,
		_w1974_,
		_w3574_,
		_w3575_
	);
	LUT3 #(
		.INIT('h32)
	) name2616 (
		_w3477_,
		_w3550_,
		_w3575_,
		_w3576_
	);
	LUT4 #(
		.INIT('haaa8)
	) name2617 (
		_w3552_,
		_w3572_,
		_w3573_,
		_w3576_,
		_w3577_
	);
	LUT3 #(
		.INIT('h40)
	) name2618 (
		_w1970_,
		_w1976_,
		_w2426_,
		_w3578_
	);
	LUT4 #(
		.INIT('hf0e0)
	) name2619 (
		_w2429_,
		_w3395_,
		_w3549_,
		_w3578_,
		_w3579_
	);
	LUT3 #(
		.INIT('ha8)
	) name2620 (
		_w1969_,
		_w2431_,
		_w3393_,
		_w3580_
	);
	LUT3 #(
		.INIT('h40)
	) name2621 (
		_w1970_,
		_w1976_,
		_w2517_,
		_w3581_
	);
	LUT3 #(
		.INIT('hc8)
	) name2622 (
		_w2514_,
		_w3548_,
		_w3581_,
		_w3582_
	);
	LUT4 #(
		.INIT('h5d7f)
	) name2623 (
		_w1966_,
		_w1968_,
		_w2502_,
		_w2548_,
		_w3583_
	);
	LUT4 #(
		.INIT('h0100)
	) name2624 (
		_w3579_,
		_w3580_,
		_w3582_,
		_w3583_,
		_w3584_
	);
	LUT3 #(
		.INIT('hcd)
	) name2625 (
		_w3552_,
		_w3577_,
		_w3584_,
		_w3585_
	);
	LUT3 #(
		.INIT('h0e)
	) name2626 (
		_w3406_,
		_w3422_,
		_w3550_,
		_w3586_
	);
	LUT3 #(
		.INIT('ha8)
	) name2627 (
		_w1969_,
		_w3477_,
		_w3575_,
		_w3587_
	);
	LUT3 #(
		.INIT('h10)
	) name2628 (
		_w1970_,
		_w1976_,
		_w3419_,
		_w3588_
	);
	LUT2 #(
		.INIT('h4)
	) name2629 (
		_w3546_,
		_w3588_,
		_w3589_
	);
	LUT4 #(
		.INIT('haaa8)
	) name2630 (
		_w3552_,
		_w3586_,
		_w3587_,
		_w3589_,
		_w3590_
	);
	LUT2 #(
		.INIT('h8)
	) name2631 (
		_w1969_,
		_w2514_,
		_w3591_
	);
	LUT4 #(
		.INIT('hf0e0)
	) name2632 (
		_w2429_,
		_w3395_,
		_w3548_,
		_w3578_,
		_w3592_
	);
	LUT4 #(
		.INIT('habef)
	) name2633 (
		_w1970_,
		_w1976_,
		_w2515_,
		_w2517_,
		_w3593_
	);
	LUT2 #(
		.INIT('h2)
	) name2634 (
		_w1969_,
		_w3593_,
		_w3594_
	);
	LUT3 #(
		.INIT('h2a)
	) name2635 (
		\wb_addr_i[25]_pad ,
		_w976_,
		_w1975_,
		_w3595_
	);
	LUT3 #(
		.INIT('h10)
	) name2636 (
		_w1972_,
		_w1974_,
		_w3595_,
		_w3596_
	);
	LUT3 #(
		.INIT('h2a)
	) name2637 (
		\wb_addr_i[26]_pad ,
		_w976_,
		_w1971_,
		_w3597_
	);
	LUT4 #(
		.INIT('habef)
	) name2638 (
		_w1970_,
		_w1976_,
		_w2517_,
		_w3597_,
		_w3598_
	);
	LUT3 #(
		.INIT('h8a)
	) name2639 (
		_w3549_,
		_w3596_,
		_w3598_,
		_w3599_
	);
	LUT4 #(
		.INIT('h0001)
	) name2640 (
		_w3591_,
		_w3592_,
		_w3594_,
		_w3599_,
		_w3600_
	);
	LUT3 #(
		.INIT('hcd)
	) name2641 (
		_w3552_,
		_w3590_,
		_w3600_,
		_w3601_
	);
	LUT3 #(
		.INIT('h0e)
	) name2642 (
		_w3374_,
		_w3475_,
		_w3550_,
		_w3602_
	);
	LUT3 #(
		.INIT('ha8)
	) name2643 (
		_w1969_,
		_w3406_,
		_w3422_,
		_w3603_
	);
	LUT3 #(
		.INIT('h10)
	) name2644 (
		_w1970_,
		_w1976_,
		_w3476_,
		_w3604_
	);
	LUT2 #(
		.INIT('h4)
	) name2645 (
		_w3546_,
		_w3604_,
		_w3605_
	);
	LUT4 #(
		.INIT('haaa8)
	) name2646 (
		_w3552_,
		_w3602_,
		_w3603_,
		_w3605_,
		_w3606_
	);
	LUT4 #(
		.INIT('h5554)
	) name2647 (
		_w3552_,
		_w3572_,
		_w3573_,
		_w3576_,
		_w3607_
	);
	LUT2 #(
		.INIT('he)
	) name2648 (
		_w3606_,
		_w3607_,
		_w3608_
	);
	LUT3 #(
		.INIT('h0e)
	) name2649 (
		_w2516_,
		_w2551_,
		_w3550_,
		_w3609_
	);
	LUT2 #(
		.INIT('h2)
	) name2650 (
		_w2654_,
		_w3546_,
		_w3610_
	);
	LUT3 #(
		.INIT('ha8)
	) name2651 (
		_w1969_,
		_w2504_,
		_w3394_,
		_w3611_
	);
	LUT4 #(
		.INIT('h5554)
	) name2652 (
		_w3552_,
		_w3609_,
		_w3610_,
		_w3611_,
		_w3612_
	);
	LUT4 #(
		.INIT('hf0e0)
	) name2653 (
		_w2514_,
		_w2548_,
		_w3549_,
		_w3581_,
		_w3613_
	);
	LUT4 #(
		.INIT('h0200)
	) name2654 (
		_w1966_,
		_w1970_,
		_w1976_,
		_w2515_,
		_w3614_
	);
	LUT4 #(
		.INIT('h0001)
	) name2655 (
		_w3580_,
		_w3582_,
		_w3613_,
		_w3614_,
		_w3615_
	);
	LUT3 #(
		.INIT('hce)
	) name2656 (
		_w3552_,
		_w3612_,
		_w3615_,
		_w3616_
	);
	LUT3 #(
		.INIT('h0e)
	) name2657 (
		_w3230_,
		_w3404_,
		_w3550_,
		_w3617_
	);
	LUT3 #(
		.INIT('ha8)
	) name2658 (
		_w1969_,
		_w3374_,
		_w3475_,
		_w3618_
	);
	LUT2 #(
		.INIT('h2)
	) name2659 (
		_w3418_,
		_w3546_,
		_w3619_
	);
	LUT4 #(
		.INIT('haaa8)
	) name2660 (
		_w3552_,
		_w3617_,
		_w3618_,
		_w3619_,
		_w3620_
	);
	LUT4 #(
		.INIT('h5554)
	) name2661 (
		_w3552_,
		_w3586_,
		_w3587_,
		_w3589_,
		_w3621_
	);
	LUT2 #(
		.INIT('he)
	) name2662 (
		_w3620_,
		_w3621_,
		_w3622_
	);
	LUT3 #(
		.INIT('h0e)
	) name2663 (
		_w2632_,
		_w3372_,
		_w3550_,
		_w3623_
	);
	LUT3 #(
		.INIT('ha8)
	) name2664 (
		_w1969_,
		_w3230_,
		_w3404_,
		_w3624_
	);
	LUT2 #(
		.INIT('h2)
	) name2665 (
		_w3478_,
		_w3546_,
		_w3625_
	);
	LUT4 #(
		.INIT('haaa8)
	) name2666 (
		_w3552_,
		_w3623_,
		_w3624_,
		_w3625_,
		_w3626_
	);
	LUT4 #(
		.INIT('h5554)
	) name2667 (
		_w3552_,
		_w3602_,
		_w3603_,
		_w3605_,
		_w3627_
	);
	LUT2 #(
		.INIT('he)
	) name2668 (
		_w3626_,
		_w3627_,
		_w3628_
	);
	LUT3 #(
		.INIT('h0e)
	) name2669 (
		_w3228_,
		_w3427_,
		_w3550_,
		_w3629_
	);
	LUT3 #(
		.INIT('ha8)
	) name2670 (
		_w1969_,
		_w2632_,
		_w3372_,
		_w3630_
	);
	LUT2 #(
		.INIT('h2)
	) name2671 (
		_w3407_,
		_w3546_,
		_w3631_
	);
	LUT4 #(
		.INIT('haaa8)
	) name2672 (
		_w3552_,
		_w3629_,
		_w3630_,
		_w3631_,
		_w3632_
	);
	LUT4 #(
		.INIT('h5554)
	) name2673 (
		_w3552_,
		_w3617_,
		_w3618_,
		_w3619_,
		_w3633_
	);
	LUT2 #(
		.INIT('he)
	) name2674 (
		_w3632_,
		_w3633_,
		_w3634_
	);
	LUT3 #(
		.INIT('h0e)
	) name2675 (
		_w2637_,
		_w2653_,
		_w3550_,
		_w3635_
	);
	LUT3 #(
		.INIT('ha8)
	) name2676 (
		_w1969_,
		_w3228_,
		_w3427_,
		_w3636_
	);
	LUT2 #(
		.INIT('h2)
	) name2677 (
		_w3375_,
		_w3546_,
		_w3637_
	);
	LUT4 #(
		.INIT('haaa8)
	) name2678 (
		_w3552_,
		_w3635_,
		_w3636_,
		_w3637_,
		_w3638_
	);
	LUT4 #(
		.INIT('h5554)
	) name2679 (
		_w3552_,
		_w3623_,
		_w3624_,
		_w3625_,
		_w3639_
	);
	LUT2 #(
		.INIT('he)
	) name2680 (
		_w3638_,
		_w3639_,
		_w3640_
	);
	LUT3 #(
		.INIT('h0e)
	) name2681 (
		_w2506_,
		_w3426_,
		_w3550_,
		_w3641_
	);
	LUT3 #(
		.INIT('ha8)
	) name2682 (
		_w1969_,
		_w2637_,
		_w2653_,
		_w3642_
	);
	LUT2 #(
		.INIT('h2)
	) name2683 (
		_w3232_,
		_w3546_,
		_w3643_
	);
	LUT4 #(
		.INIT('haaa8)
	) name2684 (
		_w3552_,
		_w3641_,
		_w3642_,
		_w3643_,
		_w3644_
	);
	LUT4 #(
		.INIT('h5554)
	) name2685 (
		_w3552_,
		_w3629_,
		_w3630_,
		_w3631_,
		_w3645_
	);
	LUT2 #(
		.INIT('he)
	) name2686 (
		_w3644_,
		_w3645_,
		_w3646_
	);
	LUT3 #(
		.INIT('h0e)
	) name2687 (
		_w2553_,
		_w2652_,
		_w3550_,
		_w3647_
	);
	LUT3 #(
		.INIT('ha8)
	) name2688 (
		_w1969_,
		_w2506_,
		_w3426_,
		_w3648_
	);
	LUT2 #(
		.INIT('h2)
	) name2689 (
		_w2635_,
		_w3546_,
		_w3649_
	);
	LUT4 #(
		.INIT('haaa8)
	) name2690 (
		_w3552_,
		_w3647_,
		_w3648_,
		_w3649_,
		_w3650_
	);
	LUT4 #(
		.INIT('h5554)
	) name2691 (
		_w3552_,
		_w3635_,
		_w3636_,
		_w3637_,
		_w3651_
	);
	LUT2 #(
		.INIT('he)
	) name2692 (
		_w3650_,
		_w3651_,
		_w3652_
	);
	LUT4 #(
		.INIT('h00f1)
	) name2693 (
		_w2506_,
		_w3426_,
		_w3550_,
		_w3552_,
		_w3653_
	);
	LUT3 #(
		.INIT('h10)
	) name2694 (
		_w3642_,
		_w3643_,
		_w3653_,
		_w3654_
	);
	LUT4 #(
		.INIT('hf100)
	) name2695 (
		_w2504_,
		_w3394_,
		_w3550_,
		_w3552_,
		_w3655_
	);
	LUT3 #(
		.INIT('h10)
	) name2696 (
		_w3545_,
		_w3547_,
		_w3655_,
		_w3656_
	);
	LUT2 #(
		.INIT('h1)
	) name2697 (
		_w3654_,
		_w3656_,
		_w3657_
	);
	LUT4 #(
		.INIT('h5554)
	) name2698 (
		_w3552_,
		_w3647_,
		_w3648_,
		_w3649_,
		_w3658_
	);
	LUT4 #(
		.INIT('haaa8)
	) name2699 (
		_w3552_,
		_w3609_,
		_w3610_,
		_w3611_,
		_w3659_
	);
	LUT2 #(
		.INIT('he)
	) name2700 (
		_w3658_,
		_w3659_,
		_w3660_
	);
	LUT3 #(
		.INIT('h70)
	) name2701 (
		_w1187_,
		_w1292_,
		_w1540_,
		_w3661_
	);
	LUT2 #(
		.INIT('hb)
	) name2702 (
		_w1539_,
		_w3661_,
		_w3662_
	);
	LUT4 #(
		.INIT('h5551)
	) name2703 (
		_w3552_,
		_w3557_,
		_w3558_,
		_w3559_,
		_w3663_
	);
	LUT2 #(
		.INIT('h8)
	) name2704 (
		_w1969_,
		_w3581_,
		_w3664_
	);
	LUT4 #(
		.INIT('h0001)
	) name2705 (
		_w3579_,
		_w3591_,
		_w3592_,
		_w3664_,
		_w3665_
	);
	LUT3 #(
		.INIT('hce)
	) name2706 (
		_w3552_,
		_w3663_,
		_w3665_,
		_w3666_
	);
	LUT4 #(
		.INIT('h1000)
	) name2707 (
		\u0_csc_reg[4]/NET0131 ,
		\u0_csc_reg[5]/NET0131 ,
		\u5_pack_le1_reg/P0001 ,
		\u7_mc_data_ir_reg[0]/P0001 ,
		_w3667_
	);
	LUT4 #(
		.INIT('h0010)
	) name2708 (
		\u0_csc_reg[4]/NET0131 ,
		\u0_csc_reg[5]/NET0131 ,
		\u5_pack_le1_reg/P0001 ,
		\u7_mc_data_ir_reg[0]/P0001 ,
		_w3668_
	);
	LUT4 #(
		.INIT('hd0f0)
	) name2709 (
		\u0_csc_reg[4]/NET0131 ,
		\u0_csc_reg[5]/NET0131 ,
		\u3_byte1_reg[0]/P0001 ,
		\u5_pack_le0_reg/P0001 ,
		_w3669_
	);
	LUT4 #(
		.INIT('h2000)
	) name2710 (
		\u0_csc_reg[4]/NET0131 ,
		\u0_csc_reg[5]/NET0131 ,
		\u5_pack_le0_reg/P0001 ,
		\u7_mc_data_ir_reg[8]/P0001 ,
		_w3670_
	);
	LUT4 #(
		.INIT('h3332)
	) name2711 (
		_w3667_,
		_w3668_,
		_w3669_,
		_w3670_,
		_w3671_
	);
	LUT4 #(
		.INIT('h1000)
	) name2712 (
		\u0_csc_reg[4]/NET0131 ,
		\u0_csc_reg[5]/NET0131 ,
		\u5_pack_le1_reg/P0001 ,
		\u7_mc_data_ir_reg[2]/P0001 ,
		_w3672_
	);
	LUT4 #(
		.INIT('h0010)
	) name2713 (
		\u0_csc_reg[4]/NET0131 ,
		\u0_csc_reg[5]/NET0131 ,
		\u5_pack_le1_reg/P0001 ,
		\u7_mc_data_ir_reg[2]/P0001 ,
		_w3673_
	);
	LUT4 #(
		.INIT('hd0f0)
	) name2714 (
		\u0_csc_reg[4]/NET0131 ,
		\u0_csc_reg[5]/NET0131 ,
		\u3_byte1_reg[2]/P0001 ,
		\u5_pack_le0_reg/P0001 ,
		_w3674_
	);
	LUT4 #(
		.INIT('h2000)
	) name2715 (
		\u0_csc_reg[4]/NET0131 ,
		\u0_csc_reg[5]/NET0131 ,
		\u5_pack_le0_reg/P0001 ,
		\u7_mc_data_ir_reg[10]/P0001 ,
		_w3675_
	);
	LUT4 #(
		.INIT('h3332)
	) name2716 (
		_w3672_,
		_w3673_,
		_w3674_,
		_w3675_,
		_w3676_
	);
	LUT4 #(
		.INIT('h1000)
	) name2717 (
		\u0_csc_reg[4]/NET0131 ,
		\u0_csc_reg[5]/NET0131 ,
		\u5_pack_le1_reg/P0001 ,
		\u7_mc_data_ir_reg[1]/P0001 ,
		_w3677_
	);
	LUT4 #(
		.INIT('h0010)
	) name2718 (
		\u0_csc_reg[4]/NET0131 ,
		\u0_csc_reg[5]/NET0131 ,
		\u5_pack_le1_reg/P0001 ,
		\u7_mc_data_ir_reg[1]/P0001 ,
		_w3678_
	);
	LUT4 #(
		.INIT('hd0f0)
	) name2719 (
		\u0_csc_reg[4]/NET0131 ,
		\u0_csc_reg[5]/NET0131 ,
		\u3_byte1_reg[1]/P0001 ,
		\u5_pack_le0_reg/P0001 ,
		_w3679_
	);
	LUT4 #(
		.INIT('h2000)
	) name2720 (
		\u0_csc_reg[4]/NET0131 ,
		\u0_csc_reg[5]/NET0131 ,
		\u5_pack_le0_reg/P0001 ,
		\u7_mc_data_ir_reg[9]/P0001 ,
		_w3680_
	);
	LUT4 #(
		.INIT('h3332)
	) name2721 (
		_w3677_,
		_w3678_,
		_w3679_,
		_w3680_,
		_w3681_
	);
	LUT4 #(
		.INIT('h1000)
	) name2722 (
		\u0_csc_reg[4]/NET0131 ,
		\u0_csc_reg[5]/NET0131 ,
		\u5_pack_le1_reg/P0001 ,
		\u7_mc_data_ir_reg[3]/P0001 ,
		_w3682_
	);
	LUT4 #(
		.INIT('h0010)
	) name2723 (
		\u0_csc_reg[4]/NET0131 ,
		\u0_csc_reg[5]/NET0131 ,
		\u5_pack_le1_reg/P0001 ,
		\u7_mc_data_ir_reg[3]/P0001 ,
		_w3683_
	);
	LUT4 #(
		.INIT('hd0f0)
	) name2724 (
		\u0_csc_reg[4]/NET0131 ,
		\u0_csc_reg[5]/NET0131 ,
		\u3_byte1_reg[3]/P0001 ,
		\u5_pack_le0_reg/P0001 ,
		_w3684_
	);
	LUT4 #(
		.INIT('h2000)
	) name2725 (
		\u0_csc_reg[4]/NET0131 ,
		\u0_csc_reg[5]/NET0131 ,
		\u5_pack_le0_reg/P0001 ,
		\u7_mc_data_ir_reg[11]/P0001 ,
		_w3685_
	);
	LUT4 #(
		.INIT('h3332)
	) name2726 (
		_w3682_,
		_w3683_,
		_w3684_,
		_w3685_,
		_w3686_
	);
	LUT4 #(
		.INIT('h1000)
	) name2727 (
		\u0_csc_reg[4]/NET0131 ,
		\u0_csc_reg[5]/NET0131 ,
		\u5_pack_le1_reg/P0001 ,
		\u7_mc_data_ir_reg[4]/P0001 ,
		_w3687_
	);
	LUT4 #(
		.INIT('h0010)
	) name2728 (
		\u0_csc_reg[4]/NET0131 ,
		\u0_csc_reg[5]/NET0131 ,
		\u5_pack_le1_reg/P0001 ,
		\u7_mc_data_ir_reg[4]/P0001 ,
		_w3688_
	);
	LUT4 #(
		.INIT('hd0f0)
	) name2729 (
		\u0_csc_reg[4]/NET0131 ,
		\u0_csc_reg[5]/NET0131 ,
		\u3_byte1_reg[4]/P0001 ,
		\u5_pack_le0_reg/P0001 ,
		_w3689_
	);
	LUT4 #(
		.INIT('h2000)
	) name2730 (
		\u0_csc_reg[4]/NET0131 ,
		\u0_csc_reg[5]/NET0131 ,
		\u5_pack_le0_reg/P0001 ,
		\u7_mc_data_ir_reg[12]/P0001 ,
		_w3690_
	);
	LUT4 #(
		.INIT('h3332)
	) name2731 (
		_w3687_,
		_w3688_,
		_w3689_,
		_w3690_,
		_w3691_
	);
	LUT4 #(
		.INIT('h1000)
	) name2732 (
		\u0_csc_reg[4]/NET0131 ,
		\u0_csc_reg[5]/NET0131 ,
		\u5_pack_le1_reg/P0001 ,
		\u7_mc_data_ir_reg[5]/P0001 ,
		_w3692_
	);
	LUT4 #(
		.INIT('h0010)
	) name2733 (
		\u0_csc_reg[4]/NET0131 ,
		\u0_csc_reg[5]/NET0131 ,
		\u5_pack_le1_reg/P0001 ,
		\u7_mc_data_ir_reg[5]/P0001 ,
		_w3693_
	);
	LUT4 #(
		.INIT('hd0f0)
	) name2734 (
		\u0_csc_reg[4]/NET0131 ,
		\u0_csc_reg[5]/NET0131 ,
		\u3_byte1_reg[5]/P0001 ,
		\u5_pack_le0_reg/P0001 ,
		_w3694_
	);
	LUT4 #(
		.INIT('h2000)
	) name2735 (
		\u0_csc_reg[4]/NET0131 ,
		\u0_csc_reg[5]/NET0131 ,
		\u5_pack_le0_reg/P0001 ,
		\u7_mc_data_ir_reg[13]/P0001 ,
		_w3695_
	);
	LUT4 #(
		.INIT('h3332)
	) name2736 (
		_w3692_,
		_w3693_,
		_w3694_,
		_w3695_,
		_w3696_
	);
	LUT4 #(
		.INIT('h1000)
	) name2737 (
		\u0_csc_reg[4]/NET0131 ,
		\u0_csc_reg[5]/NET0131 ,
		\u5_pack_le1_reg/P0001 ,
		\u7_mc_data_ir_reg[6]/P0001 ,
		_w3697_
	);
	LUT4 #(
		.INIT('h0010)
	) name2738 (
		\u0_csc_reg[4]/NET0131 ,
		\u0_csc_reg[5]/NET0131 ,
		\u5_pack_le1_reg/P0001 ,
		\u7_mc_data_ir_reg[6]/P0001 ,
		_w3698_
	);
	LUT4 #(
		.INIT('hd0f0)
	) name2739 (
		\u0_csc_reg[4]/NET0131 ,
		\u0_csc_reg[5]/NET0131 ,
		\u3_byte1_reg[6]/P0001 ,
		\u5_pack_le0_reg/P0001 ,
		_w3699_
	);
	LUT4 #(
		.INIT('h2000)
	) name2740 (
		\u0_csc_reg[4]/NET0131 ,
		\u0_csc_reg[5]/NET0131 ,
		\u5_pack_le0_reg/P0001 ,
		\u7_mc_data_ir_reg[14]/P0001 ,
		_w3700_
	);
	LUT4 #(
		.INIT('h3332)
	) name2741 (
		_w3697_,
		_w3698_,
		_w3699_,
		_w3700_,
		_w3701_
	);
	LUT4 #(
		.INIT('h1000)
	) name2742 (
		\u0_csc_reg[4]/NET0131 ,
		\u0_csc_reg[5]/NET0131 ,
		\u5_pack_le1_reg/P0001 ,
		\u7_mc_data_ir_reg[7]/P0001 ,
		_w3702_
	);
	LUT4 #(
		.INIT('h0010)
	) name2743 (
		\u0_csc_reg[4]/NET0131 ,
		\u0_csc_reg[5]/NET0131 ,
		\u5_pack_le1_reg/P0001 ,
		\u7_mc_data_ir_reg[7]/P0001 ,
		_w3703_
	);
	LUT4 #(
		.INIT('hd0f0)
	) name2744 (
		\u0_csc_reg[4]/NET0131 ,
		\u0_csc_reg[5]/NET0131 ,
		\u3_byte1_reg[7]/P0001 ,
		\u5_pack_le0_reg/P0001 ,
		_w3704_
	);
	LUT4 #(
		.INIT('h2000)
	) name2745 (
		\u0_csc_reg[4]/NET0131 ,
		\u0_csc_reg[5]/NET0131 ,
		\u5_pack_le0_reg/P0001 ,
		\u7_mc_data_ir_reg[15]/P0001 ,
		_w3705_
	);
	LUT4 #(
		.INIT('h3332)
	) name2746 (
		_w3702_,
		_w3703_,
		_w3704_,
		_w3705_,
		_w3706_
	);
	LUT4 #(
		.INIT('h0444)
	) name2747 (
		\u3_u0_wr_adr_reg[3]/NET0131 ,
		wb_cyc_i_pad,
		wb_stb_i_pad,
		wb_we_i_pad,
		_w3707_
	);
	LUT4 #(
		.INIT('h0444)
	) name2748 (
		\u3_u0_wr_adr_reg[0]/NET0131 ,
		wb_cyc_i_pad,
		wb_stb_i_pad,
		wb_we_i_pad,
		_w3708_
	);
	LUT4 #(
		.INIT('h0e1f)
	) name2749 (
		_w998_,
		_w1010_,
		_w3707_,
		_w3708_,
		_w3709_
	);
	LUT4 #(
		.INIT('h0888)
	) name2750 (
		\u3_u0_wr_adr_reg[1]/NET0131 ,
		wb_cyc_i_pad,
		wb_stb_i_pad,
		wb_we_i_pad,
		_w3710_
	);
	LUT4 #(
		.INIT('h0888)
	) name2751 (
		\u3_u0_wr_adr_reg[2]/NET0131 ,
		wb_cyc_i_pad,
		wb_stb_i_pad,
		wb_we_i_pad,
		_w3711_
	);
	LUT4 #(
		.INIT('hf1e0)
	) name2752 (
		_w998_,
		_w1010_,
		_w3710_,
		_w3711_,
		_w3712_
	);
	LUT4 #(
		.INIT('h0888)
	) name2753 (
		\u3_u0_wr_adr_reg[3]/NET0131 ,
		wb_cyc_i_pad,
		wb_stb_i_pad,
		wb_we_i_pad,
		_w3713_
	);
	LUT4 #(
		.INIT('hf1e0)
	) name2754 (
		_w998_,
		_w1010_,
		_w3711_,
		_w3713_,
		_w3714_
	);
	LUT3 #(
		.INIT('h40)
	) name2755 (
		\u0_init_req_reg/NET0131 ,
		\u0_lmr_req_reg/NET0131 ,
		\u5_lookup_ready2_reg/NET0131 ,
		_w3715_
	);
	LUT2 #(
		.INIT('h4)
	) name2756 (
		\u4_rfr_req_reg/NET0131 ,
		\u5_state_reg[1]/NET0131 ,
		_w3716_
	);
	LUT2 #(
		.INIT('h8)
	) name2757 (
		_w3715_,
		_w3716_,
		_w3717_
	);
	LUT3 #(
		.INIT('he9)
	) name2758 (
		\u5_state_reg[18]/NET0131 ,
		\u5_state_reg[19]/NET0131 ,
		\u5_state_reg[20]/NET0131 ,
		_w3718_
	);
	LUT3 #(
		.INIT('h08)
	) name2759 (
		_w2591_,
		_w2592_,
		_w3718_,
		_w3719_
	);
	LUT3 #(
		.INIT('hec)
	) name2760 (
		_w2603_,
		_w3717_,
		_w3719_,
		_w3720_
	);
	LUT3 #(
		.INIT('h2a)
	) name2761 (
		\wb_addr_i[0]_pad ,
		_w976_,
		_w1971_,
		_w3721_
	);
	LUT3 #(
		.INIT('h40)
	) name2762 (
		_w1970_,
		_w1976_,
		_w3721_,
		_w3722_
	);
	LUT3 #(
		.INIT('h2a)
	) name2763 (
		\wb_addr_i[2]_pad ,
		_w976_,
		_w1971_,
		_w3723_
	);
	LUT3 #(
		.INIT('h10)
	) name2764 (
		_w1970_,
		_w1976_,
		_w3723_,
		_w3724_
	);
	LUT3 #(
		.INIT('h2a)
	) name2765 (
		\wb_addr_i[1]_pad ,
		_w976_,
		_w1975_,
		_w3725_
	);
	LUT3 #(
		.INIT('h10)
	) name2766 (
		_w1972_,
		_w1974_,
		_w3725_,
		_w3726_
	);
	LUT4 #(
		.INIT('h5554)
	) name2767 (
		_w2424_,
		_w3722_,
		_w3724_,
		_w3726_,
		_w3727_
	);
	LUT2 #(
		.INIT('h4)
	) name2768 (
		\u1_u0_out_r_reg[0]/P0001 ,
		\u5_tmr2_done_reg/NET0131 ,
		_w3728_
	);
	LUT4 #(
		.INIT('h7500)
	) name2769 (
		_w964_,
		_w1974_,
		_w2417_,
		_w3728_,
		_w3729_
	);
	LUT2 #(
		.INIT('h1)
	) name2770 (
		\u1_acs_addr_reg[0]/P0001 ,
		\u5_tmr2_done_reg/NET0131 ,
		_w3730_
	);
	LUT3 #(
		.INIT('h01)
	) name2771 (
		\u1_acs_addr_reg[0]/P0001 ,
		\u5_state_reg[42]/NET0131 ,
		\u5_state_reg[44]/NET0131 ,
		_w3731_
	);
	LUT4 #(
		.INIT('h040f)
	) name2772 (
		_w1974_,
		_w2417_,
		_w3730_,
		_w3731_,
		_w3732_
	);
	LUT3 #(
		.INIT('h20)
	) name2773 (
		_w2424_,
		_w3729_,
		_w3732_,
		_w3733_
	);
	LUT2 #(
		.INIT('he)
	) name2774 (
		_w3727_,
		_w3733_,
		_w3734_
	);
	LUT2 #(
		.INIT('h4)
	) name2775 (
		\u1_u0_out_r_reg[10]/P0001 ,
		\u5_tmr2_done_reg/NET0131 ,
		_w3735_
	);
	LUT4 #(
		.INIT('h7500)
	) name2776 (
		_w964_,
		_w1974_,
		_w2417_,
		_w3735_,
		_w3736_
	);
	LUT2 #(
		.INIT('h1)
	) name2777 (
		\u1_acs_addr_reg[10]/P0001 ,
		\u5_tmr2_done_reg/NET0131 ,
		_w3737_
	);
	LUT3 #(
		.INIT('h01)
	) name2778 (
		\u1_acs_addr_reg[10]/P0001 ,
		\u5_state_reg[42]/NET0131 ,
		\u5_state_reg[44]/NET0131 ,
		_w3738_
	);
	LUT4 #(
		.INIT('h040f)
	) name2779 (
		_w1974_,
		_w2417_,
		_w3737_,
		_w3738_,
		_w3739_
	);
	LUT3 #(
		.INIT('h20)
	) name2780 (
		_w2424_,
		_w3736_,
		_w3739_,
		_w3740_
	);
	LUT3 #(
		.INIT('h40)
	) name2781 (
		_w1970_,
		_w1976_,
		_w3541_,
		_w3741_
	);
	LUT4 #(
		.INIT('h5554)
	) name2782 (
		_w2424_,
		_w3575_,
		_w3604_,
		_w3741_,
		_w3742_
	);
	LUT2 #(
		.INIT('he)
	) name2783 (
		_w3740_,
		_w3742_,
		_w3743_
	);
	LUT3 #(
		.INIT('h2a)
	) name2784 (
		\wb_addr_i[2]_pad ,
		_w976_,
		_w1975_,
		_w3744_
	);
	LUT3 #(
		.INIT('h10)
	) name2785 (
		_w1972_,
		_w1974_,
		_w3744_,
		_w3745_
	);
	LUT3 #(
		.INIT('h2a)
	) name2786 (
		\wb_addr_i[3]_pad ,
		_w976_,
		_w1971_,
		_w3746_
	);
	LUT3 #(
		.INIT('h2a)
	) name2787 (
		\wb_addr_i[1]_pad ,
		_w976_,
		_w1971_,
		_w3747_
	);
	LUT4 #(
		.INIT('habef)
	) name2788 (
		_w1970_,
		_w1976_,
		_w3746_,
		_w3747_,
		_w3748_
	);
	LUT3 #(
		.INIT('h45)
	) name2789 (
		_w2424_,
		_w3745_,
		_w3748_,
		_w3749_
	);
	LUT2 #(
		.INIT('h4)
	) name2790 (
		\u1_u0_out_r_reg[1]/P0001 ,
		\u5_tmr2_done_reg/NET0131 ,
		_w3750_
	);
	LUT4 #(
		.INIT('h7500)
	) name2791 (
		_w964_,
		_w1974_,
		_w2417_,
		_w3750_,
		_w3751_
	);
	LUT2 #(
		.INIT('h1)
	) name2792 (
		\u1_acs_addr_reg[1]/P0001 ,
		\u5_tmr2_done_reg/NET0131 ,
		_w3752_
	);
	LUT3 #(
		.INIT('h01)
	) name2793 (
		\u1_acs_addr_reg[1]/P0001 ,
		\u5_state_reg[42]/NET0131 ,
		\u5_state_reg[44]/NET0131 ,
		_w3753_
	);
	LUT4 #(
		.INIT('h040f)
	) name2794 (
		_w1974_,
		_w2417_,
		_w3752_,
		_w3753_,
		_w3754_
	);
	LUT3 #(
		.INIT('h20)
	) name2795 (
		_w2424_,
		_w3751_,
		_w3754_,
		_w3755_
	);
	LUT2 #(
		.INIT('he)
	) name2796 (
		_w3749_,
		_w3755_,
		_w3756_
	);
	LUT3 #(
		.INIT('h40)
	) name2797 (
		_w1970_,
		_w1976_,
		_w3723_,
		_w3757_
	);
	LUT3 #(
		.INIT('h2a)
	) name2798 (
		\wb_addr_i[3]_pad ,
		_w976_,
		_w1975_,
		_w3758_
	);
	LUT3 #(
		.INIT('h10)
	) name2799 (
		_w1972_,
		_w1974_,
		_w3758_,
		_w3759_
	);
	LUT3 #(
		.INIT('h10)
	) name2800 (
		_w1970_,
		_w1976_,
		_w3517_,
		_w3760_
	);
	LUT4 #(
		.INIT('h5554)
	) name2801 (
		_w2424_,
		_w3757_,
		_w3759_,
		_w3760_,
		_w3761_
	);
	LUT2 #(
		.INIT('h4)
	) name2802 (
		\u1_u0_out_r_reg[2]/P0001 ,
		\u5_tmr2_done_reg/NET0131 ,
		_w3762_
	);
	LUT4 #(
		.INIT('h7500)
	) name2803 (
		_w964_,
		_w1974_,
		_w2417_,
		_w3762_,
		_w3763_
	);
	LUT2 #(
		.INIT('h1)
	) name2804 (
		\u1_acs_addr_reg[2]/P0001 ,
		\u5_tmr2_done_reg/NET0131 ,
		_w3764_
	);
	LUT3 #(
		.INIT('h01)
	) name2805 (
		\u1_acs_addr_reg[2]/P0001 ,
		\u5_state_reg[42]/NET0131 ,
		\u5_state_reg[44]/NET0131 ,
		_w3765_
	);
	LUT4 #(
		.INIT('h040f)
	) name2806 (
		_w1974_,
		_w2417_,
		_w3764_,
		_w3765_,
		_w3766_
	);
	LUT3 #(
		.INIT('h20)
	) name2807 (
		_w2424_,
		_w3763_,
		_w3766_,
		_w3767_
	);
	LUT2 #(
		.INIT('he)
	) name2808 (
		_w3761_,
		_w3767_,
		_w3768_
	);
	LUT3 #(
		.INIT('h40)
	) name2809 (
		_w1970_,
		_w1976_,
		_w3746_,
		_w3769_
	);
	LUT3 #(
		.INIT('h2a)
	) name2810 (
		\wb_addr_i[4]_pad ,
		_w976_,
		_w1975_,
		_w3770_
	);
	LUT3 #(
		.INIT('h10)
	) name2811 (
		_w1972_,
		_w1974_,
		_w3770_,
		_w3771_
	);
	LUT3 #(
		.INIT('h2a)
	) name2812 (
		\wb_addr_i[5]_pad ,
		_w976_,
		_w1971_,
		_w3772_
	);
	LUT3 #(
		.INIT('h10)
	) name2813 (
		_w1970_,
		_w1976_,
		_w3772_,
		_w3773_
	);
	LUT4 #(
		.INIT('h5554)
	) name2814 (
		_w2424_,
		_w3769_,
		_w3771_,
		_w3773_,
		_w3774_
	);
	LUT2 #(
		.INIT('h4)
	) name2815 (
		\u1_u0_out_r_reg[3]/P0001 ,
		\u5_tmr2_done_reg/NET0131 ,
		_w3775_
	);
	LUT4 #(
		.INIT('h7500)
	) name2816 (
		_w964_,
		_w1974_,
		_w2417_,
		_w3775_,
		_w3776_
	);
	LUT2 #(
		.INIT('h1)
	) name2817 (
		\u1_acs_addr_reg[3]/P0001 ,
		\u5_tmr2_done_reg/NET0131 ,
		_w3777_
	);
	LUT3 #(
		.INIT('h01)
	) name2818 (
		\u1_acs_addr_reg[3]/P0001 ,
		\u5_state_reg[42]/NET0131 ,
		\u5_state_reg[44]/NET0131 ,
		_w3778_
	);
	LUT4 #(
		.INIT('h040f)
	) name2819 (
		_w1974_,
		_w2417_,
		_w3777_,
		_w3778_,
		_w3779_
	);
	LUT3 #(
		.INIT('h20)
	) name2820 (
		_w2424_,
		_w3776_,
		_w3779_,
		_w3780_
	);
	LUT2 #(
		.INIT('he)
	) name2821 (
		_w3774_,
		_w3780_,
		_w3781_
	);
	LUT3 #(
		.INIT('h40)
	) name2822 (
		_w1970_,
		_w1976_,
		_w3772_,
		_w3782_
	);
	LUT3 #(
		.INIT('h2a)
	) name2823 (
		\wb_addr_i[6]_pad ,
		_w976_,
		_w1975_,
		_w3783_
	);
	LUT3 #(
		.INIT('h10)
	) name2824 (
		_w1972_,
		_w1974_,
		_w3783_,
		_w3784_
	);
	LUT3 #(
		.INIT('h10)
	) name2825 (
		_w1970_,
		_w1976_,
		_w3443_,
		_w3785_
	);
	LUT4 #(
		.INIT('h5554)
	) name2826 (
		_w2424_,
		_w3782_,
		_w3784_,
		_w3785_,
		_w3786_
	);
	LUT2 #(
		.INIT('h4)
	) name2827 (
		\u1_u0_out_r_reg[5]/P0001 ,
		\u5_tmr2_done_reg/NET0131 ,
		_w3787_
	);
	LUT4 #(
		.INIT('h7500)
	) name2828 (
		_w964_,
		_w1974_,
		_w2417_,
		_w3787_,
		_w3788_
	);
	LUT2 #(
		.INIT('h1)
	) name2829 (
		\u1_acs_addr_reg[5]/P0001 ,
		\u5_tmr2_done_reg/NET0131 ,
		_w3789_
	);
	LUT3 #(
		.INIT('h01)
	) name2830 (
		\u1_acs_addr_reg[5]/P0001 ,
		\u5_state_reg[42]/NET0131 ,
		\u5_state_reg[44]/NET0131 ,
		_w3790_
	);
	LUT4 #(
		.INIT('h040f)
	) name2831 (
		_w1974_,
		_w2417_,
		_w3789_,
		_w3790_,
		_w3791_
	);
	LUT3 #(
		.INIT('h20)
	) name2832 (
		_w2424_,
		_w3788_,
		_w3791_,
		_w3792_
	);
	LUT2 #(
		.INIT('he)
	) name2833 (
		_w3786_,
		_w3792_,
		_w3793_
	);
	LUT3 #(
		.INIT('h40)
	) name2834 (
		_w1970_,
		_w1976_,
		_w3521_,
		_w3794_
	);
	LUT3 #(
		.INIT('h2a)
	) name2835 (
		\wb_addr_i[7]_pad ,
		_w976_,
		_w1975_,
		_w3795_
	);
	LUT3 #(
		.INIT('h10)
	) name2836 (
		_w1972_,
		_w1974_,
		_w3795_,
		_w3796_
	);
	LUT3 #(
		.INIT('h10)
	) name2837 (
		_w1970_,
		_w1976_,
		_w3537_,
		_w3797_
	);
	LUT4 #(
		.INIT('h5554)
	) name2838 (
		_w2424_,
		_w3794_,
		_w3796_,
		_w3797_,
		_w3798_
	);
	LUT2 #(
		.INIT('h4)
	) name2839 (
		\u1_u0_out_r_reg[6]/P0001 ,
		\u5_tmr2_done_reg/NET0131 ,
		_w3799_
	);
	LUT4 #(
		.INIT('h7500)
	) name2840 (
		_w964_,
		_w1974_,
		_w2417_,
		_w3799_,
		_w3800_
	);
	LUT2 #(
		.INIT('h1)
	) name2841 (
		\u1_acs_addr_reg[6]/P0001 ,
		\u5_tmr2_done_reg/NET0131 ,
		_w3801_
	);
	LUT3 #(
		.INIT('h01)
	) name2842 (
		\u1_acs_addr_reg[6]/P0001 ,
		\u5_state_reg[42]/NET0131 ,
		\u5_state_reg[44]/NET0131 ,
		_w3802_
	);
	LUT4 #(
		.INIT('h040f)
	) name2843 (
		_w1974_,
		_w2417_,
		_w3801_,
		_w3802_,
		_w3803_
	);
	LUT3 #(
		.INIT('h20)
	) name2844 (
		_w2424_,
		_w3800_,
		_w3803_,
		_w3804_
	);
	LUT2 #(
		.INIT('he)
	) name2845 (
		_w3798_,
		_w3804_,
		_w3805_
	);
	LUT2 #(
		.INIT('h4)
	) name2846 (
		\u1_u0_out_r_reg[9]/P0001 ,
		\u5_tmr2_done_reg/NET0131 ,
		_w3806_
	);
	LUT4 #(
		.INIT('h7500)
	) name2847 (
		_w964_,
		_w1974_,
		_w2417_,
		_w3806_,
		_w3807_
	);
	LUT2 #(
		.INIT('h1)
	) name2848 (
		\u1_acs_addr_reg[9]/P0001 ,
		\u5_tmr2_done_reg/NET0131 ,
		_w3808_
	);
	LUT3 #(
		.INIT('h01)
	) name2849 (
		\u1_acs_addr_reg[9]/P0001 ,
		\u5_state_reg[42]/NET0131 ,
		\u5_state_reg[44]/NET0131 ,
		_w3809_
	);
	LUT4 #(
		.INIT('h040f)
	) name2850 (
		_w1974_,
		_w2417_,
		_w3808_,
		_w3809_,
		_w3810_
	);
	LUT3 #(
		.INIT('h20)
	) name2851 (
		_w2424_,
		_w3807_,
		_w3810_,
		_w3811_
	);
	LUT3 #(
		.INIT('h40)
	) name2852 (
		_w1970_,
		_w1976_,
		_w3447_,
		_w3812_
	);
	LUT4 #(
		.INIT('h5554)
	) name2853 (
		_w2424_,
		_w3571_,
		_w3588_,
		_w3812_,
		_w3813_
	);
	LUT2 #(
		.INIT('he)
	) name2854 (
		_w3811_,
		_w3813_,
		_w3814_
	);
	LUT4 #(
		.INIT('h5554)
	) name2855 (
		\u5_cnt_reg/NET0131 ,
		_w1045_,
		_w1141_,
		_w1145_,
		_w3815_
	);
	LUT4 #(
		.INIT('hfe00)
	) name2856 (
		\wb_addr_i[29]_pad ,
		\wb_addr_i[30]_pad ,
		\wb_addr_i[31]_pad ,
		wb_stb_i_pad,
		_w3816_
	);
	LUT2 #(
		.INIT('h8)
	) name2857 (
		\u5_wb_cycle_reg/NET0131 ,
		wb_cyc_i_pad,
		_w3817_
	);
	LUT2 #(
		.INIT('h4)
	) name2858 (
		_w3816_,
		_w3817_,
		_w3818_
	);
	LUT3 #(
		.INIT('hf8)
	) name2859 (
		_w1581_,
		_w1586_,
		_w3818_,
		_w3819_
	);
	LUT3 #(
		.INIT('h47)
	) name2860 (
		\mem_ack_r_reg/P0001 ,
		\u5_wr_cycle_reg/NET0131 ,
		wb_stb_i_pad,
		_w3820_
	);
	LUT3 #(
		.INIT('hb8)
	) name2861 (
		\mem_ack_r_reg/P0001 ,
		\u5_wr_cycle_reg/NET0131 ,
		wb_stb_i_pad,
		_w3821_
	);
	LUT4 #(
		.INIT('h404c)
	) name2862 (
		\mem_ack_r_reg/P0001 ,
		\u1_col_adr_reg[8]/P0001 ,
		\u5_wr_cycle_reg/NET0131 ,
		wb_stb_i_pad,
		_w3822_
	);
	LUT4 #(
		.INIT('hb080)
	) name2863 (
		\mem_ack_r_reg/P0001 ,
		\u5_wr_cycle_reg/NET0131 ,
		\wb_addr_i[10]_pad ,
		wb_stb_i_pad,
		_w3823_
	);
	LUT4 #(
		.INIT('he000)
	) name2864 (
		_w1966_,
		_w1968_,
		_w1976_,
		_w3823_,
		_w3824_
	);
	LUT3 #(
		.INIT('hdc)
	) name2865 (
		_w1973_,
		_w3822_,
		_w3824_,
		_w3825_
	);
	LUT3 #(
		.INIT('h6a)
	) name2866 (
		\u1_acs_addr_reg[7]/P0001 ,
		_w3563_,
		_w3564_,
		_w3826_
	);
	LUT3 #(
		.INIT('h0d)
	) name2867 (
		\u5_state_reg[61]/NET0131 ,
		\u5_tmr2_done_reg/NET0131 ,
		\u7_mc_ack_r_reg/NET0131 ,
		_w3827_
	);
	LUT4 #(
		.INIT('h0080)
	) name2868 (
		_w985_,
		_w987_,
		_w1082_,
		_w3827_,
		_w3828_
	);
	LUT2 #(
		.INIT('h2)
	) name2869 (
		\u5_state_reg[61]/NET0131 ,
		\u5_tmr_done_reg/NET0131 ,
		_w3829_
	);
	LUT3 #(
		.INIT('h07)
	) name2870 (
		_w1059_,
		_w3828_,
		_w3829_,
		_w3830_
	);
	LUT3 #(
		.INIT('h57)
	) name2871 (
		_w1059_,
		_w1086_,
		_w3828_,
		_w3831_
	);
	LUT3 #(
		.INIT('h13)
	) name2872 (
		_w1320_,
		_w3830_,
		_w3831_,
		_w3832_
	);
	LUT4 #(
		.INIT('haf23)
	) name2873 (
		\u0_csr_r2_reg[1]/NET0131 ,
		\u0_csr_r2_reg[4]/NET0131 ,
		\u4_ps_cnt_reg[1]/NET0131 ,
		\u4_ps_cnt_reg[4]/NET0131 ,
		_w3833_
	);
	LUT4 #(
		.INIT('h8caf)
	) name2874 (
		\u0_csr_r2_reg[2]/NET0131 ,
		\u0_csr_r2_reg[4]/NET0131 ,
		\u4_ps_cnt_reg[2]/NET0131 ,
		\u4_ps_cnt_reg[4]/NET0131 ,
		_w3834_
	);
	LUT4 #(
		.INIT('h8421)
	) name2875 (
		\u0_csr_r2_reg[5]/NET0131 ,
		\u0_csr_r2_reg[7]/NET0131 ,
		\u4_ps_cnt_reg[5]/NET0131 ,
		\u4_ps_cnt_reg[7]/NET0131 ,
		_w3835_
	);
	LUT3 #(
		.INIT('h80)
	) name2876 (
		_w3833_,
		_w3834_,
		_w3835_,
		_w3836_
	);
	LUT4 #(
		.INIT('hf531)
	) name2877 (
		\u0_csr_r2_reg[0]/NET0131 ,
		\u0_csr_r2_reg[3]/NET0131 ,
		\u4_ps_cnt_reg[0]/NET0131 ,
		\u4_ps_cnt_reg[3]/NET0131 ,
		_w3837_
	);
	LUT4 #(
		.INIT('haf23)
	) name2878 (
		\u0_csr_r2_reg[0]/NET0131 ,
		\u0_csr_r2_reg[1]/NET0131 ,
		\u4_ps_cnt_reg[0]/NET0131 ,
		\u4_ps_cnt_reg[1]/NET0131 ,
		_w3838_
	);
	LUT4 #(
		.INIT('hf531)
	) name2879 (
		\u0_csr_r2_reg[2]/NET0131 ,
		\u0_csr_r2_reg[6]/NET0131 ,
		\u4_ps_cnt_reg[2]/NET0131 ,
		\u4_ps_cnt_reg[6]/NET0131 ,
		_w3839_
	);
	LUT4 #(
		.INIT('h8caf)
	) name2880 (
		\u0_csr_r2_reg[3]/NET0131 ,
		\u0_csr_r2_reg[6]/NET0131 ,
		\u4_ps_cnt_reg[3]/NET0131 ,
		\u4_ps_cnt_reg[6]/NET0131 ,
		_w3840_
	);
	LUT4 #(
		.INIT('h8000)
	) name2881 (
		_w3837_,
		_w3838_,
		_w3839_,
		_w3840_,
		_w3841_
	);
	LUT2 #(
		.INIT('h8)
	) name2882 (
		_w3836_,
		_w3841_,
		_w3842_
	);
	LUT4 #(
		.INIT('h0001)
	) name2883 (
		\u0_csr_r2_reg[4]/NET0131 ,
		\u0_csr_r2_reg[5]/NET0131 ,
		\u0_csr_r2_reg[6]/NET0131 ,
		\u0_csr_r2_reg[7]/NET0131 ,
		_w3843_
	);
	LUT4 #(
		.INIT('h0001)
	) name2884 (
		\u0_csr_r2_reg[0]/NET0131 ,
		\u0_csr_r2_reg[1]/NET0131 ,
		\u0_csr_r2_reg[2]/NET0131 ,
		\u0_csr_r2_reg[3]/NET0131 ,
		_w3844_
	);
	LUT2 #(
		.INIT('h8)
	) name2885 (
		_w3843_,
		_w3844_,
		_w3845_
	);
	LUT3 #(
		.INIT('h08)
	) name2886 (
		_w3836_,
		_w3841_,
		_w3845_,
		_w3846_
	);
	LUT4 #(
		.INIT('h8000)
	) name2887 (
		\u4_ps_cnt_reg[0]/NET0131 ,
		\u4_ps_cnt_reg[1]/NET0131 ,
		\u4_ps_cnt_reg[2]/NET0131 ,
		\u4_rfr_en_reg/NET0131 ,
		_w3847_
	);
	LUT3 #(
		.INIT('h6c)
	) name2888 (
		\u4_ps_cnt_reg[3]/NET0131 ,
		\u4_ps_cnt_reg[4]/NET0131 ,
		_w3847_,
		_w3848_
	);
	LUT4 #(
		.INIT('hf700)
	) name2889 (
		_w3836_,
		_w3841_,
		_w3845_,
		_w3848_,
		_w3849_
	);
	LUT4 #(
		.INIT('h0078)
	) name2890 (
		\u4_rfr_ce_reg/NET0131 ,
		\u4_rfr_cnt_reg[0]/NET0131 ,
		\u4_rfr_cnt_reg[1]/NET0131 ,
		\u5_rfr_ack_r_reg/NET0131 ,
		_w3850_
	);
	LUT3 #(
		.INIT('h01)
	) name2891 (
		\u5_state_reg[14]/NET0131 ,
		\u5_state_reg[17]/NET0131 ,
		\u5_state_reg[7]/NET0131 ,
		_w3851_
	);
	LUT4 #(
		.INIT('h8000)
	) name2892 (
		_w1020_,
		_w1021_,
		_w2588_,
		_w3851_,
		_w3852_
	);
	LUT4 #(
		.INIT('h0014)
	) name2893 (
		\u5_state_reg[0]/NET0131 ,
		\u5_state_reg[33]/NET0131 ,
		\u5_state_reg[34]/NET0131 ,
		\u5_state_reg[35]/NET0131 ,
		_w3853_
	);
	LUT4 #(
		.INIT('h0001)
	) name2894 (
		\u5_state_reg[25]/NET0131 ,
		\u5_state_reg[26]/NET0131 ,
		\u5_state_reg[5]/NET0131 ,
		\u5_state_reg[6]/NET0131 ,
		_w3854_
	);
	LUT3 #(
		.INIT('h80)
	) name2895 (
		_w2600_,
		_w3853_,
		_w3854_,
		_w3855_
	);
	LUT4 #(
		.INIT('h8000)
	) name2896 (
		_w1029_,
		_w2584_,
		_w3852_,
		_w3855_,
		_w3856_
	);
	LUT2 #(
		.INIT('h1)
	) name2897 (
		\u0_init_req_reg/NET0131 ,
		\u0_lmr_req_reg/NET0131 ,
		_w3857_
	);
	LUT3 #(
		.INIT('h04)
	) name2898 (
		\u4_rfr_req_reg/NET0131 ,
		\u5_state_reg[35]/NET0131 ,
		\u5_susp_req_r_reg/NET0131 ,
		_w3858_
	);
	LUT2 #(
		.INIT('h8)
	) name2899 (
		_w3857_,
		_w3858_,
		_w3859_
	);
	LUT3 #(
		.INIT('h10)
	) name2900 (
		_w1564_,
		_w1566_,
		_w3859_,
		_w3860_
	);
	LUT3 #(
		.INIT('hf8)
	) name2901 (
		_w2599_,
		_w3856_,
		_w3860_,
		_w3861_
	);
	LUT3 #(
		.INIT('h06)
	) name2902 (
		\u4_rfr_ce_reg/NET0131 ,
		\u4_rfr_cnt_reg[0]/NET0131 ,
		\u5_rfr_ack_r_reg/NET0131 ,
		_w3862_
	);
	LUT4 #(
		.INIT('h8000)
	) name2903 (
		\u4_rfr_ce_reg/NET0131 ,
		\u4_rfr_cnt_reg[0]/NET0131 ,
		\u4_rfr_cnt_reg[1]/NET0131 ,
		\u4_rfr_cnt_reg[2]/NET0131 ,
		_w3863_
	);
	LUT2 #(
		.INIT('h2)
	) name2904 (
		\u4_rfr_cnt_reg[2]/NET0131 ,
		\u5_rfr_ack_r_reg/NET0131 ,
		_w3864_
	);
	LUT4 #(
		.INIT('h0080)
	) name2905 (
		\u4_rfr_ce_reg/NET0131 ,
		\u4_rfr_cnt_reg[0]/NET0131 ,
		\u4_rfr_cnt_reg[1]/NET0131 ,
		\u5_rfr_ack_r_reg/NET0131 ,
		_w3865_
	);
	LUT3 #(
		.INIT('h54)
	) name2906 (
		_w3863_,
		_w3864_,
		_w3865_,
		_w3866_
	);
	LUT3 #(
		.INIT('h12)
	) name2907 (
		\u4_rfr_cnt_reg[3]/NET0131 ,
		\u5_rfr_ack_r_reg/NET0131 ,
		_w3863_,
		_w3867_
	);
	LUT4 #(
		.INIT('h060c)
	) name2908 (
		\u4_rfr_cnt_reg[3]/NET0131 ,
		\u4_rfr_cnt_reg[4]/NET0131 ,
		\u5_rfr_ack_r_reg/NET0131 ,
		_w3863_,
		_w3868_
	);
	LUT3 #(
		.INIT('h15)
	) name2909 (
		\u4_rfr_cnt_reg[5]/NET0131 ,
		_w3469_,
		_w3863_,
		_w3869_
	);
	LUT3 #(
		.INIT('h80)
	) name2910 (
		\u4_rfr_cnt_reg[3]/NET0131 ,
		\u4_rfr_cnt_reg[4]/NET0131 ,
		\u4_rfr_cnt_reg[5]/NET0131 ,
		_w3870_
	);
	LUT3 #(
		.INIT('h15)
	) name2911 (
		\u5_rfr_ack_r_reg/NET0131 ,
		_w3863_,
		_w3870_,
		_w3871_
	);
	LUT2 #(
		.INIT('h4)
	) name2912 (
		_w3869_,
		_w3871_,
		_w3872_
	);
	LUT2 #(
		.INIT('h2)
	) name2913 (
		\u4_rfr_cnt_reg[6]/NET0131 ,
		\u5_rfr_ack_r_reg/NET0131 ,
		_w3873_
	);
	LUT4 #(
		.INIT('h1222)
	) name2914 (
		\u4_rfr_cnt_reg[6]/NET0131 ,
		\u5_rfr_ack_r_reg/NET0131 ,
		_w3863_,
		_w3870_,
		_w3874_
	);
	LUT2 #(
		.INIT('h8)
	) name2915 (
		\u4_rfr_cnt_reg[6]/NET0131 ,
		\u4_rfr_cnt_reg[7]/NET0131 ,
		_w3875_
	);
	LUT3 #(
		.INIT('h80)
	) name2916 (
		_w3863_,
		_w3870_,
		_w3875_,
		_w3876_
	);
	LUT2 #(
		.INIT('h2)
	) name2917 (
		\u4_rfr_cnt_reg[7]/NET0131 ,
		\u5_rfr_ack_r_reg/NET0131 ,
		_w3877_
	);
	LUT4 #(
		.INIT('h007f)
	) name2918 (
		_w3863_,
		_w3870_,
		_w3873_,
		_w3877_,
		_w3878_
	);
	LUT2 #(
		.INIT('h1)
	) name2919 (
		_w3876_,
		_w3878_,
		_w3879_
	);
	LUT3 #(
		.INIT('h80)
	) name2920 (
		\u5_cs_le_reg/P0001 ,
		wb_cyc_i_pad,
		wb_stb_i_pad,
		_w3880_
	);
	LUT4 #(
		.INIT('h20a0)
	) name2921 (
		\u0_wp_err_reg/NET0131 ,
		\u5_cs_le_reg/P0001 ,
		wb_cyc_i_pad,
		wb_stb_i_pad,
		_w3881_
	);
	LUT4 #(
		.INIT('h0002)
	) name2922 (
		\u0_u0_csc_reg[8]/P0001 ,
		_w2914_,
		_w2915_,
		_w2916_,
		_w3882_
	);
	LUT3 #(
		.INIT('h80)
	) name2923 (
		_w2907_,
		_w2912_,
		_w3882_,
		_w3883_
	);
	LUT4 #(
		.INIT('h0002)
	) name2924 (
		\u0_u1_csc_reg[8]/P0001 ,
		_w2926_,
		_w2927_,
		_w2928_,
		_w3884_
	);
	LUT3 #(
		.INIT('h80)
	) name2925 (
		_w2919_,
		_w2924_,
		_w3884_,
		_w3885_
	);
	LUT4 #(
		.INIT('h8000)
	) name2926 (
		\u5_cs_le_reg/P0001 ,
		wb_cyc_i_pad,
		wb_stb_i_pad,
		wb_we_i_pad,
		_w3886_
	);
	LUT4 #(
		.INIT('hfeaa)
	) name2927 (
		_w3881_,
		_w3883_,
		_w3885_,
		_w3886_,
		_w3887_
	);
	LUT2 #(
		.INIT('h8)
	) name2928 (
		\u5_mc_adv_r1_reg/NET0131 ,
		\u5_mc_le_reg/NET0131 ,
		_w3888_
	);
	LUT3 #(
		.INIT('h4c)
	) name2929 (
		_w991_,
		_w1568_,
		_w2306_,
		_w3889_
	);
	LUT4 #(
		.INIT('h1555)
	) name2930 (
		\u5_mc_le_reg/NET0131 ,
		_w991_,
		_w995_,
		_w1055_,
		_w3890_
	);
	LUT4 #(
		.INIT('hcdcc)
	) name2931 (
		_w1057_,
		_w3888_,
		_w3889_,
		_w3890_,
		_w3891_
	);
	LUT3 #(
		.INIT('hb0)
	) name2932 (
		_w1966_,
		_w1968_,
		_w3552_,
		_w3892_
	);
	LUT4 #(
		.INIT('he0f0)
	) name2933 (
		_w1972_,
		_w1974_,
		_w3552_,
		_w3595_,
		_w3893_
	);
	LUT3 #(
		.INIT('h13)
	) name2934 (
		_w3598_,
		_w3892_,
		_w3893_,
		_w3894_
	);
	LUT3 #(
		.INIT('h0b)
	) name2935 (
		_w1966_,
		_w1968_,
		_w3552_,
		_w3895_
	);
	LUT4 #(
		.INIT('h00ef)
	) name2936 (
		_w1970_,
		_w1976_,
		_w2515_,
		_w3552_,
		_w3896_
	);
	LUT4 #(
		.INIT('h0e0f)
	) name2937 (
		_w2514_,
		_w3581_,
		_w3895_,
		_w3896_,
		_w3897_
	);
	LUT2 #(
		.INIT('h8)
	) name2938 (
		_w3894_,
		_w3897_,
		_w3898_
	);
	LUT2 #(
		.INIT('h8)
	) name2939 (
		\u5_cmd_asserted_reg/NET0131 ,
		_w1263_,
		_w3899_
	);
	LUT3 #(
		.INIT('h80)
	) name2940 (
		_w984_,
		_w1046_,
		_w3899_,
		_w3900_
	);
	LUT4 #(
		.INIT('h8ccc)
	) name2941 (
		\u5_ir_cnt_reg[0]/P0001 ,
		\u5_ir_cnt_reg[1]/P0001 ,
		_w1035_,
		_w3900_,
		_w3901_
	);
	LUT2 #(
		.INIT('h1)
	) name2942 (
		\u5_ir_cnt_reg[0]/P0001 ,
		\u5_ir_cnt_reg[1]/P0001 ,
		_w3902_
	);
	LUT4 #(
		.INIT('h1555)
	) name2943 (
		\u5_state_reg[22]/NET0131 ,
		_w1035_,
		_w3900_,
		_w3902_,
		_w3903_
	);
	LUT2 #(
		.INIT('hb)
	) name2944 (
		_w3901_,
		_w3903_,
		_w3904_
	);
	LUT3 #(
		.INIT('h80)
	) name2945 (
		\u4_ps_cnt_reg[3]/NET0131 ,
		\u4_ps_cnt_reg[4]/NET0131 ,
		\u4_ps_cnt_reg[5]/NET0131 ,
		_w3905_
	);
	LUT4 #(
		.INIT('h6ccc)
	) name2946 (
		\u4_ps_cnt_reg[6]/NET0131 ,
		\u4_ps_cnt_reg[7]/NET0131 ,
		_w3847_,
		_w3905_,
		_w3906_
	);
	LUT4 #(
		.INIT('hf700)
	) name2947 (
		_w3836_,
		_w3841_,
		_w3845_,
		_w3906_,
		_w3907_
	);
	LUT4 #(
		.INIT('h0001)
	) name2948 (
		\u5_ir_cnt_reg[0]/P0001 ,
		\u5_ir_cnt_reg[1]/P0001 ,
		\u5_ir_cnt_reg[2]/P0001 ,
		\u5_ir_cnt_reg[3]/P0001 ,
		_w3908_
	);
	LUT4 #(
		.INIT('h4000)
	) name2949 (
		\u5_state_reg[22]/NET0131 ,
		_w1035_,
		_w3900_,
		_w3908_,
		_w3909_
	);
	LUT3 #(
		.INIT('h01)
	) name2950 (
		\u5_ir_cnt_reg[0]/P0001 ,
		\u5_ir_cnt_reg[1]/P0001 ,
		\u5_ir_cnt_reg[2]/P0001 ,
		_w3910_
	);
	LUT2 #(
		.INIT('h2)
	) name2951 (
		\u5_ir_cnt_reg[3]/P0001 ,
		\u5_state_reg[22]/NET0131 ,
		_w3911_
	);
	LUT4 #(
		.INIT('h7f00)
	) name2952 (
		_w1035_,
		_w3900_,
		_w3910_,
		_w3911_,
		_w3912_
	);
	LUT2 #(
		.INIT('he)
	) name2953 (
		_w3909_,
		_w3912_,
		_w3913_
	);
	LUT3 #(
		.INIT('ha8)
	) name2954 (
		\u3_u0_wr_adr_reg[1]/NET0131 ,
		_w998_,
		_w1010_,
		_w3914_
	);
	LUT3 #(
		.INIT('ha8)
	) name2955 (
		\u3_u0_wr_adr_reg[2]/NET0131 ,
		_w998_,
		_w1010_,
		_w3915_
	);
	LUT4 #(
		.INIT('h1222)
	) name2956 (
		\u5_ir_cnt_reg[0]/P0001 ,
		\u5_state_reg[22]/NET0131 ,
		_w1035_,
		_w3900_,
		_w3916_
	);
	LUT2 #(
		.INIT('h2)
	) name2957 (
		\u5_ir_cnt_reg[2]/P0001 ,
		\u5_state_reg[22]/NET0131 ,
		_w3917_
	);
	LUT4 #(
		.INIT('h7f00)
	) name2958 (
		_w1035_,
		_w3900_,
		_w3902_,
		_w3917_,
		_w3918_
	);
	LUT2 #(
		.INIT('h1)
	) name2959 (
		\u5_ir_cnt_reg[2]/P0001 ,
		\u5_state_reg[22]/NET0131 ,
		_w3919_
	);
	LUT4 #(
		.INIT('h8000)
	) name2960 (
		_w1035_,
		_w3900_,
		_w3902_,
		_w3919_,
		_w3920_
	);
	LUT2 #(
		.INIT('he)
	) name2961 (
		_w3918_,
		_w3920_,
		_w3921_
	);
	LUT4 #(
		.INIT('h8c23)
	) name2962 (
		\u1_row_adr_reg[6]/P0001 ,
		\u1_row_adr_reg[7]/P0001 ,
		\u2_u1_b3_last_row_reg[6]/P0001 ,
		\u2_u1_b3_last_row_reg[7]/P0001 ,
		_w3922_
	);
	LUT4 #(
		.INIT('hf531)
	) name2963 (
		\u1_row_adr_reg[0]/P0001 ,
		\u1_row_adr_reg[8]/P0001 ,
		\u2_u1_b3_last_row_reg[0]/P0001 ,
		\u2_u1_b3_last_row_reg[8]/P0001 ,
		_w3923_
	);
	LUT4 #(
		.INIT('h8caf)
	) name2964 (
		\u1_row_adr_reg[11]/P0001 ,
		\u1_row_adr_reg[8]/P0001 ,
		\u2_u1_b3_last_row_reg[11]/P0001 ,
		\u2_u1_b3_last_row_reg[8]/P0001 ,
		_w3924_
	);
	LUT4 #(
		.INIT('h8caf)
	) name2965 (
		\u1_row_adr_reg[12]/P0001 ,
		\u1_row_adr_reg[1]/P0001 ,
		\u2_u1_b3_last_row_reg[12]/P0001 ,
		\u2_u1_b3_last_row_reg[1]/P0001 ,
		_w3925_
	);
	LUT4 #(
		.INIT('hc4f5)
	) name2966 (
		\u1_row_adr_reg[1]/P0001 ,
		\u1_row_adr_reg[4]/P0001 ,
		\u2_u1_b3_last_row_reg[1]/P0001 ,
		\u2_u1_b3_last_row_reg[4]/P0001 ,
		_w3926_
	);
	LUT4 #(
		.INIT('h8000)
	) name2967 (
		_w3923_,
		_w3924_,
		_w3925_,
		_w3926_,
		_w3927_
	);
	LUT4 #(
		.INIT('haf23)
	) name2968 (
		\u1_row_adr_reg[0]/P0001 ,
		\u1_row_adr_reg[11]/P0001 ,
		\u2_u1_b3_last_row_reg[0]/P0001 ,
		\u2_u1_b3_last_row_reg[11]/P0001 ,
		_w3928_
	);
	LUT4 #(
		.INIT('hf531)
	) name2969 (
		\u1_row_adr_reg[12]/P0001 ,
		\u1_row_adr_reg[2]/P0001 ,
		\u2_u1_b3_last_row_reg[12]/P0001 ,
		\u2_u1_b3_last_row_reg[2]/P0001 ,
		_w3929_
	);
	LUT2 #(
		.INIT('h6)
	) name2970 (
		\u1_row_adr_reg[10]/P0001 ,
		\u2_u1_b3_last_row_reg[10]/P0001 ,
		_w3930_
	);
	LUT4 #(
		.INIT('h8808)
	) name2971 (
		\u1_bank_adr_reg[0]/P0001 ,
		\u1_bank_adr_reg[1]/P0001 ,
		\u1_row_adr_reg[3]/P0001 ,
		\u2_u1_b3_last_row_reg[3]/P0001 ,
		_w3931_
	);
	LUT4 #(
		.INIT('h0800)
	) name2972 (
		_w3928_,
		_w3929_,
		_w3930_,
		_w3931_,
		_w3932_
	);
	LUT4 #(
		.INIT('h8caf)
	) name2973 (
		\u1_row_adr_reg[5]/P0001 ,
		\u1_row_adr_reg[9]/P0001 ,
		\u2_u1_b3_last_row_reg[5]/P0001 ,
		\u2_u1_b3_last_row_reg[9]/P0001 ,
		_w3933_
	);
	LUT4 #(
		.INIT('haf23)
	) name2974 (
		\u1_row_adr_reg[2]/P0001 ,
		\u1_row_adr_reg[4]/P0001 ,
		\u2_u1_b3_last_row_reg[2]/P0001 ,
		\u2_u1_b3_last_row_reg[4]/P0001 ,
		_w3934_
	);
	LUT4 #(
		.INIT('hf531)
	) name2975 (
		\u1_row_adr_reg[5]/P0001 ,
		\u1_row_adr_reg[9]/P0001 ,
		\u2_u1_b3_last_row_reg[5]/P0001 ,
		\u2_u1_b3_last_row_reg[9]/P0001 ,
		_w3935_
	);
	LUT4 #(
		.INIT('haf23)
	) name2976 (
		\u1_row_adr_reg[3]/P0001 ,
		\u1_row_adr_reg[6]/P0001 ,
		\u2_u1_b3_last_row_reg[3]/P0001 ,
		\u2_u1_b3_last_row_reg[6]/P0001 ,
		_w3936_
	);
	LUT4 #(
		.INIT('h8000)
	) name2977 (
		_w3933_,
		_w3934_,
		_w3935_,
		_w3936_,
		_w3937_
	);
	LUT4 #(
		.INIT('h8000)
	) name2978 (
		_w3922_,
		_w3927_,
		_w3932_,
		_w3937_,
		_w3938_
	);
	LUT4 #(
		.INIT('h84a5)
	) name2979 (
		\u1_row_adr_reg[3]/P0001 ,
		\u1_row_adr_reg[8]/P0001 ,
		\u2_u1_b2_last_row_reg[3]/P0001 ,
		\u2_u1_b2_last_row_reg[8]/P0001 ,
		_w3939_
	);
	LUT4 #(
		.INIT('h8caf)
	) name2980 (
		\u1_row_adr_reg[2]/P0001 ,
		\u1_row_adr_reg[4]/P0001 ,
		\u2_u1_b2_last_row_reg[2]/P0001 ,
		\u2_u1_b2_last_row_reg[4]/P0001 ,
		_w3940_
	);
	LUT4 #(
		.INIT('haf23)
	) name2981 (
		\u1_row_adr_reg[0]/P0001 ,
		\u1_row_adr_reg[8]/P0001 ,
		\u2_u1_b2_last_row_reg[0]/P0001 ,
		\u2_u1_b2_last_row_reg[8]/P0001 ,
		_w3941_
	);
	LUT4 #(
		.INIT('hc4f5)
	) name2982 (
		\u1_row_adr_reg[2]/P0001 ,
		\u1_row_adr_reg[7]/P0001 ,
		\u2_u1_b2_last_row_reg[2]/P0001 ,
		\u2_u1_b2_last_row_reg[7]/P0001 ,
		_w3942_
	);
	LUT4 #(
		.INIT('hf531)
	) name2983 (
		\u1_row_adr_reg[0]/P0001 ,
		\u1_row_adr_reg[7]/P0001 ,
		\u2_u1_b2_last_row_reg[0]/P0001 ,
		\u2_u1_b2_last_row_reg[7]/P0001 ,
		_w3943_
	);
	LUT4 #(
		.INIT('h8000)
	) name2984 (
		_w3940_,
		_w3941_,
		_w3942_,
		_w3943_,
		_w3944_
	);
	LUT4 #(
		.INIT('haf23)
	) name2985 (
		\u1_row_adr_reg[11]/P0001 ,
		\u1_row_adr_reg[1]/P0001 ,
		\u2_u1_b2_last_row_reg[11]/P0001 ,
		\u2_u1_b2_last_row_reg[1]/P0001 ,
		_w3945_
	);
	LUT4 #(
		.INIT('hf531)
	) name2986 (
		\u1_row_adr_reg[11]/P0001 ,
		\u1_row_adr_reg[9]/P0001 ,
		\u2_u1_b2_last_row_reg[11]/P0001 ,
		\u2_u1_b2_last_row_reg[9]/P0001 ,
		_w3946_
	);
	LUT4 #(
		.INIT('h4404)
	) name2987 (
		\u1_bank_adr_reg[0]/P0001 ,
		\u1_bank_adr_reg[1]/P0001 ,
		\u1_row_adr_reg[12]/P0001 ,
		\u2_u1_b2_last_row_reg[12]/P0001 ,
		_w3947_
	);
	LUT4 #(
		.INIT('hf531)
	) name2988 (
		\u1_row_adr_reg[5]/P0001 ,
		\u1_row_adr_reg[6]/P0001 ,
		\u2_u1_b2_last_row_reg[5]/P0001 ,
		\u2_u1_b2_last_row_reg[6]/P0001 ,
		_w3948_
	);
	LUT4 #(
		.INIT('h8000)
	) name2989 (
		_w3945_,
		_w3946_,
		_w3947_,
		_w3948_,
		_w3949_
	);
	LUT4 #(
		.INIT('h8caf)
	) name2990 (
		\u1_row_adr_reg[5]/P0001 ,
		\u1_row_adr_reg[9]/P0001 ,
		\u2_u1_b2_last_row_reg[5]/P0001 ,
		\u2_u1_b2_last_row_reg[9]/P0001 ,
		_w3950_
	);
	LUT4 #(
		.INIT('hf531)
	) name2991 (
		\u1_row_adr_reg[10]/P0001 ,
		\u1_row_adr_reg[4]/P0001 ,
		\u2_u1_b2_last_row_reg[10]/P0001 ,
		\u2_u1_b2_last_row_reg[4]/P0001 ,
		_w3951_
	);
	LUT4 #(
		.INIT('h8caf)
	) name2992 (
		\u1_row_adr_reg[10]/P0001 ,
		\u1_row_adr_reg[1]/P0001 ,
		\u2_u1_b2_last_row_reg[10]/P0001 ,
		\u2_u1_b2_last_row_reg[1]/P0001 ,
		_w3952_
	);
	LUT4 #(
		.INIT('h8caf)
	) name2993 (
		\u1_row_adr_reg[12]/P0001 ,
		\u1_row_adr_reg[6]/P0001 ,
		\u2_u1_b2_last_row_reg[12]/P0001 ,
		\u2_u1_b2_last_row_reg[6]/P0001 ,
		_w3953_
	);
	LUT4 #(
		.INIT('h8000)
	) name2994 (
		_w3950_,
		_w3951_,
		_w3952_,
		_w3953_,
		_w3954_
	);
	LUT4 #(
		.INIT('h8000)
	) name2995 (
		_w3939_,
		_w3944_,
		_w3949_,
		_w3954_,
		_w3955_
	);
	LUT2 #(
		.INIT('h4)
	) name2996 (
		\u1_row_adr_reg[4]/P0001 ,
		\u2_u1_b0_last_row_reg[4]/P0001 ,
		_w3956_
	);
	LUT2 #(
		.INIT('h1)
	) name2997 (
		\u1_bank_adr_reg[0]/P0001 ,
		\u1_bank_adr_reg[1]/P0001 ,
		_w3957_
	);
	LUT4 #(
		.INIT('h1101)
	) name2998 (
		\u1_bank_adr_reg[0]/P0001 ,
		\u1_bank_adr_reg[1]/P0001 ,
		\u1_row_adr_reg[5]/P0001 ,
		\u2_u1_b0_last_row_reg[5]/P0001 ,
		_w3958_
	);
	LUT2 #(
		.INIT('h4)
	) name2999 (
		_w3956_,
		_w3958_,
		_w3959_
	);
	LUT4 #(
		.INIT('hf531)
	) name3000 (
		\u1_row_adr_reg[2]/P0001 ,
		\u1_row_adr_reg[9]/P0001 ,
		\u2_u1_b0_last_row_reg[2]/P0001 ,
		\u2_u1_b0_last_row_reg[9]/P0001 ,
		_w3960_
	);
	LUT4 #(
		.INIT('hf531)
	) name3001 (
		\u1_row_adr_reg[10]/P0001 ,
		\u1_row_adr_reg[1]/P0001 ,
		\u2_u1_b0_last_row_reg[10]/P0001 ,
		\u2_u1_b0_last_row_reg[1]/P0001 ,
		_w3961_
	);
	LUT4 #(
		.INIT('hf531)
	) name3002 (
		\u1_row_adr_reg[11]/P0001 ,
		\u1_row_adr_reg[6]/P0001 ,
		\u2_u1_b0_last_row_reg[11]/P0001 ,
		\u2_u1_b0_last_row_reg[6]/P0001 ,
		_w3962_
	);
	LUT4 #(
		.INIT('hc4f5)
	) name3003 (
		\u1_row_adr_reg[3]/P0001 ,
		\u1_row_adr_reg[9]/P0001 ,
		\u2_u1_b0_last_row_reg[3]/P0001 ,
		\u2_u1_b0_last_row_reg[9]/P0001 ,
		_w3963_
	);
	LUT4 #(
		.INIT('h8000)
	) name3004 (
		_w3960_,
		_w3961_,
		_w3962_,
		_w3963_,
		_w3964_
	);
	LUT4 #(
		.INIT('haf23)
	) name3005 (
		\u1_row_adr_reg[10]/P0001 ,
		\u1_row_adr_reg[12]/P0001 ,
		\u2_u1_b0_last_row_reg[10]/P0001 ,
		\u2_u1_b0_last_row_reg[12]/P0001 ,
		_w3965_
	);
	LUT4 #(
		.INIT('hc4f5)
	) name3006 (
		\u1_row_adr_reg[4]/P0001 ,
		\u1_row_adr_reg[8]/P0001 ,
		\u2_u1_b0_last_row_reg[4]/P0001 ,
		\u2_u1_b0_last_row_reg[8]/P0001 ,
		_w3966_
	);
	LUT4 #(
		.INIT('h8421)
	) name3007 (
		\u1_row_adr_reg[0]/P0001 ,
		\u1_row_adr_reg[7]/P0001 ,
		\u2_u1_b0_last_row_reg[0]/P0001 ,
		\u2_u1_b0_last_row_reg[7]/P0001 ,
		_w3967_
	);
	LUT3 #(
		.INIT('h80)
	) name3008 (
		_w3965_,
		_w3966_,
		_w3967_,
		_w3968_
	);
	LUT4 #(
		.INIT('h8caf)
	) name3009 (
		\u1_row_adr_reg[11]/P0001 ,
		\u1_row_adr_reg[5]/P0001 ,
		\u2_u1_b0_last_row_reg[11]/P0001 ,
		\u2_u1_b0_last_row_reg[5]/P0001 ,
		_w3969_
	);
	LUT4 #(
		.INIT('h8caf)
	) name3010 (
		\u1_row_adr_reg[1]/P0001 ,
		\u1_row_adr_reg[2]/P0001 ,
		\u2_u1_b0_last_row_reg[1]/P0001 ,
		\u2_u1_b0_last_row_reg[2]/P0001 ,
		_w3970_
	);
	LUT4 #(
		.INIT('h8caf)
	) name3011 (
		\u1_row_adr_reg[12]/P0001 ,
		\u1_row_adr_reg[3]/P0001 ,
		\u2_u1_b0_last_row_reg[12]/P0001 ,
		\u2_u1_b0_last_row_reg[3]/P0001 ,
		_w3971_
	);
	LUT4 #(
		.INIT('haf23)
	) name3012 (
		\u1_row_adr_reg[6]/P0001 ,
		\u1_row_adr_reg[8]/P0001 ,
		\u2_u1_b0_last_row_reg[6]/P0001 ,
		\u2_u1_b0_last_row_reg[8]/P0001 ,
		_w3972_
	);
	LUT4 #(
		.INIT('h8000)
	) name3013 (
		_w3969_,
		_w3970_,
		_w3971_,
		_w3972_,
		_w3973_
	);
	LUT4 #(
		.INIT('h8000)
	) name3014 (
		_w3959_,
		_w3964_,
		_w3968_,
		_w3973_,
		_w3974_
	);
	LUT4 #(
		.INIT('hc431)
	) name3015 (
		\u1_row_adr_reg[12]/P0001 ,
		\u1_row_adr_reg[3]/P0001 ,
		\u2_u1_b1_last_row_reg[12]/P0001 ,
		\u2_u1_b1_last_row_reg[3]/P0001 ,
		_w3975_
	);
	LUT4 #(
		.INIT('hc4f5)
	) name3016 (
		\u1_row_adr_reg[1]/P0001 ,
		\u1_row_adr_reg[6]/P0001 ,
		\u2_u1_b1_last_row_reg[1]/P0001 ,
		\u2_u1_b1_last_row_reg[6]/P0001 ,
		_w3976_
	);
	LUT4 #(
		.INIT('haf23)
	) name3017 (
		\u1_row_adr_reg[12]/P0001 ,
		\u1_row_adr_reg[5]/P0001 ,
		\u2_u1_b1_last_row_reg[12]/P0001 ,
		\u2_u1_b1_last_row_reg[5]/P0001 ,
		_w3977_
	);
	LUT4 #(
		.INIT('haf23)
	) name3018 (
		\u1_row_adr_reg[5]/P0001 ,
		\u1_row_adr_reg[9]/P0001 ,
		\u2_u1_b1_last_row_reg[5]/P0001 ,
		\u2_u1_b1_last_row_reg[9]/P0001 ,
		_w3978_
	);
	LUT4 #(
		.INIT('haf23)
	) name3019 (
		\u1_row_adr_reg[10]/P0001 ,
		\u1_row_adr_reg[6]/P0001 ,
		\u2_u1_b1_last_row_reg[10]/P0001 ,
		\u2_u1_b1_last_row_reg[6]/P0001 ,
		_w3979_
	);
	LUT4 #(
		.INIT('h8000)
	) name3020 (
		_w3976_,
		_w3977_,
		_w3978_,
		_w3979_,
		_w3980_
	);
	LUT4 #(
		.INIT('h8caf)
	) name3021 (
		\u1_row_adr_reg[11]/P0001 ,
		\u1_row_adr_reg[7]/P0001 ,
		\u2_u1_b1_last_row_reg[11]/P0001 ,
		\u2_u1_b1_last_row_reg[7]/P0001 ,
		_w3981_
	);
	LUT4 #(
		.INIT('hf531)
	) name3022 (
		\u1_row_adr_reg[10]/P0001 ,
		\u1_row_adr_reg[8]/P0001 ,
		\u2_u1_b1_last_row_reg[10]/P0001 ,
		\u2_u1_b1_last_row_reg[8]/P0001 ,
		_w3982_
	);
	LUT4 #(
		.INIT('h2202)
	) name3023 (
		\u1_bank_adr_reg[0]/P0001 ,
		\u1_bank_adr_reg[1]/P0001 ,
		\u1_row_adr_reg[11]/P0001 ,
		\u2_u1_b1_last_row_reg[11]/P0001 ,
		_w3983_
	);
	LUT4 #(
		.INIT('hf531)
	) name3024 (
		\u1_row_adr_reg[0]/P0001 ,
		\u1_row_adr_reg[2]/P0001 ,
		\u2_u1_b1_last_row_reg[0]/P0001 ,
		\u2_u1_b1_last_row_reg[2]/P0001 ,
		_w3984_
	);
	LUT4 #(
		.INIT('h8000)
	) name3025 (
		_w3981_,
		_w3982_,
		_w3983_,
		_w3984_,
		_w3985_
	);
	LUT4 #(
		.INIT('h8caf)
	) name3026 (
		\u1_row_adr_reg[1]/P0001 ,
		\u1_row_adr_reg[8]/P0001 ,
		\u2_u1_b1_last_row_reg[1]/P0001 ,
		\u2_u1_b1_last_row_reg[8]/P0001 ,
		_w3986_
	);
	LUT4 #(
		.INIT('h8caf)
	) name3027 (
		\u1_row_adr_reg[2]/P0001 ,
		\u1_row_adr_reg[9]/P0001 ,
		\u2_u1_b1_last_row_reg[2]/P0001 ,
		\u2_u1_b1_last_row_reg[9]/P0001 ,
		_w3987_
	);
	LUT4 #(
		.INIT('haf23)
	) name3028 (
		\u1_row_adr_reg[0]/P0001 ,
		\u1_row_adr_reg[4]/P0001 ,
		\u2_u1_b1_last_row_reg[0]/P0001 ,
		\u2_u1_b1_last_row_reg[4]/P0001 ,
		_w3988_
	);
	LUT4 #(
		.INIT('haf23)
	) name3029 (
		\u1_row_adr_reg[4]/P0001 ,
		\u1_row_adr_reg[7]/P0001 ,
		\u2_u1_b1_last_row_reg[4]/P0001 ,
		\u2_u1_b1_last_row_reg[7]/P0001 ,
		_w3989_
	);
	LUT4 #(
		.INIT('h8000)
	) name3030 (
		_w3986_,
		_w3987_,
		_w3988_,
		_w3989_,
		_w3990_
	);
	LUT4 #(
		.INIT('h8000)
	) name3031 (
		_w3975_,
		_w3980_,
		_w3985_,
		_w3990_,
		_w3991_
	);
	LUT4 #(
		.INIT('h0001)
	) name3032 (
		_w3938_,
		_w3955_,
		_w3974_,
		_w3991_,
		_w3992_
	);
	LUT4 #(
		.INIT('ha521)
	) name3033 (
		\u1_row_adr_reg[11]/P0001 ,
		\u1_row_adr_reg[5]/P0001 ,
		\u2_u0_b2_last_row_reg[11]/P0001 ,
		\u2_u0_b2_last_row_reg[5]/P0001 ,
		_w3993_
	);
	LUT4 #(
		.INIT('haf23)
	) name3034 (
		\u1_row_adr_reg[10]/P0001 ,
		\u1_row_adr_reg[9]/P0001 ,
		\u2_u0_b2_last_row_reg[10]/P0001 ,
		\u2_u0_b2_last_row_reg[9]/P0001 ,
		_w3994_
	);
	LUT2 #(
		.INIT('h9)
	) name3035 (
		\u1_row_adr_reg[8]/P0001 ,
		\u2_u0_b2_last_row_reg[8]/P0001 ,
		_w3995_
	);
	LUT4 #(
		.INIT('h8caf)
	) name3036 (
		\u1_row_adr_reg[1]/P0001 ,
		\u1_row_adr_reg[2]/P0001 ,
		\u2_u0_b2_last_row_reg[1]/P0001 ,
		\u2_u0_b2_last_row_reg[2]/P0001 ,
		_w3996_
	);
	LUT4 #(
		.INIT('hc4f5)
	) name3037 (
		\u1_row_adr_reg[3]/P0001 ,
		\u1_row_adr_reg[9]/P0001 ,
		\u2_u0_b2_last_row_reg[3]/P0001 ,
		\u2_u0_b2_last_row_reg[9]/P0001 ,
		_w3997_
	);
	LUT4 #(
		.INIT('h8000)
	) name3038 (
		_w3994_,
		_w3995_,
		_w3996_,
		_w3997_,
		_w3998_
	);
	LUT4 #(
		.INIT('h4404)
	) name3039 (
		\u1_bank_adr_reg[0]/P0001 ,
		\u1_bank_adr_reg[1]/P0001 ,
		\u1_row_adr_reg[7]/P0001 ,
		\u2_u0_b2_last_row_reg[7]/P0001 ,
		_w3999_
	);
	LUT4 #(
		.INIT('hf531)
	) name3040 (
		\u1_row_adr_reg[2]/P0001 ,
		\u1_row_adr_reg[6]/P0001 ,
		\u2_u0_b2_last_row_reg[2]/P0001 ,
		\u2_u0_b2_last_row_reg[6]/P0001 ,
		_w4000_
	);
	LUT4 #(
		.INIT('h8421)
	) name3041 (
		\u1_row_adr_reg[0]/P0001 ,
		\u1_row_adr_reg[4]/P0001 ,
		\u2_u0_b2_last_row_reg[0]/P0001 ,
		\u2_u0_b2_last_row_reg[4]/P0001 ,
		_w4001_
	);
	LUT3 #(
		.INIT('h80)
	) name3042 (
		_w3999_,
		_w4000_,
		_w4001_,
		_w4002_
	);
	LUT2 #(
		.INIT('h9)
	) name3043 (
		\u1_row_adr_reg[12]/P0001 ,
		\u2_u0_b2_last_row_reg[12]/P0001 ,
		_w4003_
	);
	LUT4 #(
		.INIT('hc4f5)
	) name3044 (
		\u1_row_adr_reg[10]/P0001 ,
		\u1_row_adr_reg[5]/P0001 ,
		\u2_u0_b2_last_row_reg[10]/P0001 ,
		\u2_u0_b2_last_row_reg[5]/P0001 ,
		_w4004_
	);
	LUT4 #(
		.INIT('h8caf)
	) name3045 (
		\u1_row_adr_reg[6]/P0001 ,
		\u1_row_adr_reg[7]/P0001 ,
		\u2_u0_b2_last_row_reg[6]/P0001 ,
		\u2_u0_b2_last_row_reg[7]/P0001 ,
		_w4005_
	);
	LUT4 #(
		.INIT('hc4f5)
	) name3046 (
		\u1_row_adr_reg[1]/P0001 ,
		\u1_row_adr_reg[3]/P0001 ,
		\u2_u0_b2_last_row_reg[1]/P0001 ,
		\u2_u0_b2_last_row_reg[3]/P0001 ,
		_w4006_
	);
	LUT4 #(
		.INIT('h8000)
	) name3047 (
		_w4003_,
		_w4004_,
		_w4005_,
		_w4006_,
		_w4007_
	);
	LUT4 #(
		.INIT('h8000)
	) name3048 (
		_w3993_,
		_w3998_,
		_w4002_,
		_w4007_,
		_w4008_
	);
	LUT2 #(
		.INIT('h2)
	) name3049 (
		\u1_row_adr_reg[3]/P0001 ,
		\u2_u0_b1_last_row_reg[3]/P0001 ,
		_w4009_
	);
	LUT4 #(
		.INIT('haf23)
	) name3050 (
		\u1_row_adr_reg[12]/P0001 ,
		\u1_row_adr_reg[6]/P0001 ,
		\u2_u0_b1_last_row_reg[12]/P0001 ,
		\u2_u0_b1_last_row_reg[6]/P0001 ,
		_w4010_
	);
	LUT2 #(
		.INIT('h4)
	) name3051 (
		_w4009_,
		_w4010_,
		_w4011_
	);
	LUT4 #(
		.INIT('hc4f5)
	) name3052 (
		\u1_row_adr_reg[1]/P0001 ,
		\u1_row_adr_reg[7]/P0001 ,
		\u2_u0_b1_last_row_reg[1]/P0001 ,
		\u2_u0_b1_last_row_reg[7]/P0001 ,
		_w4012_
	);
	LUT2 #(
		.INIT('h9)
	) name3053 (
		\u1_row_adr_reg[11]/P0001 ,
		\u2_u0_b1_last_row_reg[11]/P0001 ,
		_w4013_
	);
	LUT4 #(
		.INIT('haf23)
	) name3054 (
		\u1_row_adr_reg[3]/P0001 ,
		\u1_row_adr_reg[8]/P0001 ,
		\u2_u0_b1_last_row_reg[3]/P0001 ,
		\u2_u0_b1_last_row_reg[8]/P0001 ,
		_w4014_
	);
	LUT4 #(
		.INIT('h8caf)
	) name3055 (
		\u1_row_adr_reg[0]/P0001 ,
		\u1_row_adr_reg[10]/P0001 ,
		\u2_u0_b1_last_row_reg[0]/P0001 ,
		\u2_u0_b1_last_row_reg[10]/P0001 ,
		_w4015_
	);
	LUT4 #(
		.INIT('h8000)
	) name3056 (
		_w4012_,
		_w4013_,
		_w4014_,
		_w4015_,
		_w4016_
	);
	LUT4 #(
		.INIT('hc4f5)
	) name3057 (
		\u1_row_adr_reg[5]/P0001 ,
		\u1_row_adr_reg[9]/P0001 ,
		\u2_u0_b1_last_row_reg[5]/P0001 ,
		\u2_u0_b1_last_row_reg[9]/P0001 ,
		_w4017_
	);
	LUT4 #(
		.INIT('hc4f5)
	) name3058 (
		\u1_row_adr_reg[12]/P0001 ,
		\u1_row_adr_reg[6]/P0001 ,
		\u2_u0_b1_last_row_reg[12]/P0001 ,
		\u2_u0_b1_last_row_reg[6]/P0001 ,
		_w4018_
	);
	LUT4 #(
		.INIT('h2022)
	) name3059 (
		\u1_bank_adr_reg[0]/P0001 ,
		\u1_bank_adr_reg[1]/P0001 ,
		\u1_row_adr_reg[1]/P0001 ,
		\u2_u0_b1_last_row_reg[1]/P0001 ,
		_w4019_
	);
	LUT4 #(
		.INIT('hf531)
	) name3060 (
		\u1_row_adr_reg[4]/P0001 ,
		\u1_row_adr_reg[9]/P0001 ,
		\u2_u0_b1_last_row_reg[4]/P0001 ,
		\u2_u0_b1_last_row_reg[9]/P0001 ,
		_w4020_
	);
	LUT4 #(
		.INIT('h8000)
	) name3061 (
		_w4017_,
		_w4018_,
		_w4019_,
		_w4020_,
		_w4021_
	);
	LUT4 #(
		.INIT('hc4f5)
	) name3062 (
		\u1_row_adr_reg[10]/P0001 ,
		\u1_row_adr_reg[2]/P0001 ,
		\u2_u0_b1_last_row_reg[10]/P0001 ,
		\u2_u0_b1_last_row_reg[2]/P0001 ,
		_w4022_
	);
	LUT4 #(
		.INIT('hc4f5)
	) name3063 (
		\u1_row_adr_reg[0]/P0001 ,
		\u1_row_adr_reg[8]/P0001 ,
		\u2_u0_b1_last_row_reg[0]/P0001 ,
		\u2_u0_b1_last_row_reg[8]/P0001 ,
		_w4023_
	);
	LUT4 #(
		.INIT('haf23)
	) name3064 (
		\u1_row_adr_reg[5]/P0001 ,
		\u1_row_adr_reg[7]/P0001 ,
		\u2_u0_b1_last_row_reg[5]/P0001 ,
		\u2_u0_b1_last_row_reg[7]/P0001 ,
		_w4024_
	);
	LUT4 #(
		.INIT('hc4f5)
	) name3065 (
		\u1_row_adr_reg[2]/P0001 ,
		\u1_row_adr_reg[4]/P0001 ,
		\u2_u0_b1_last_row_reg[2]/P0001 ,
		\u2_u0_b1_last_row_reg[4]/P0001 ,
		_w4025_
	);
	LUT4 #(
		.INIT('h8000)
	) name3066 (
		_w4022_,
		_w4023_,
		_w4024_,
		_w4025_,
		_w4026_
	);
	LUT4 #(
		.INIT('h8000)
	) name3067 (
		_w4011_,
		_w4016_,
		_w4021_,
		_w4026_,
		_w4027_
	);
	LUT4 #(
		.INIT('ha521)
	) name3068 (
		\u1_row_adr_reg[12]/P0001 ,
		\u1_row_adr_reg[5]/P0001 ,
		\u2_u0_b0_last_row_reg[12]/P0001 ,
		\u2_u0_b0_last_row_reg[5]/P0001 ,
		_w4028_
	);
	LUT4 #(
		.INIT('hf531)
	) name3069 (
		\u1_row_adr_reg[10]/P0001 ,
		\u1_row_adr_reg[11]/P0001 ,
		\u2_u0_b0_last_row_reg[10]/P0001 ,
		\u2_u0_b0_last_row_reg[11]/P0001 ,
		_w4029_
	);
	LUT4 #(
		.INIT('h8caf)
	) name3070 (
		\u1_row_adr_reg[0]/P0001 ,
		\u1_row_adr_reg[6]/P0001 ,
		\u2_u0_b0_last_row_reg[0]/P0001 ,
		\u2_u0_b0_last_row_reg[6]/P0001 ,
		_w4030_
	);
	LUT4 #(
		.INIT('haf23)
	) name3071 (
		\u1_row_adr_reg[10]/P0001 ,
		\u1_row_adr_reg[6]/P0001 ,
		\u2_u0_b0_last_row_reg[10]/P0001 ,
		\u2_u0_b0_last_row_reg[6]/P0001 ,
		_w4031_
	);
	LUT4 #(
		.INIT('h8caf)
	) name3072 (
		\u1_row_adr_reg[2]/P0001 ,
		\u1_row_adr_reg[9]/P0001 ,
		\u2_u0_b0_last_row_reg[2]/P0001 ,
		\u2_u0_b0_last_row_reg[9]/P0001 ,
		_w4032_
	);
	LUT4 #(
		.INIT('h8000)
	) name3073 (
		_w4029_,
		_w4030_,
		_w4031_,
		_w4032_,
		_w4033_
	);
	LUT4 #(
		.INIT('hf531)
	) name3074 (
		\u1_row_adr_reg[1]/P0001 ,
		\u1_row_adr_reg[7]/P0001 ,
		\u2_u0_b0_last_row_reg[1]/P0001 ,
		\u2_u0_b0_last_row_reg[7]/P0001 ,
		_w4034_
	);
	LUT4 #(
		.INIT('haf23)
	) name3075 (
		\u1_row_adr_reg[11]/P0001 ,
		\u1_row_adr_reg[8]/P0001 ,
		\u2_u0_b0_last_row_reg[11]/P0001 ,
		\u2_u0_b0_last_row_reg[8]/P0001 ,
		_w4035_
	);
	LUT4 #(
		.INIT('h1011)
	) name3076 (
		\u1_bank_adr_reg[0]/P0001 ,
		\u1_bank_adr_reg[1]/P0001 ,
		\u1_row_adr_reg[5]/P0001 ,
		\u2_u0_b0_last_row_reg[5]/P0001 ,
		_w4036_
	);
	LUT4 #(
		.INIT('h8caf)
	) name3077 (
		\u1_row_adr_reg[4]/P0001 ,
		\u1_row_adr_reg[8]/P0001 ,
		\u2_u0_b0_last_row_reg[4]/P0001 ,
		\u2_u0_b0_last_row_reg[8]/P0001 ,
		_w4037_
	);
	LUT4 #(
		.INIT('h8000)
	) name3078 (
		_w4034_,
		_w4035_,
		_w4036_,
		_w4037_,
		_w4038_
	);
	LUT4 #(
		.INIT('h8caf)
	) name3079 (
		\u1_row_adr_reg[1]/P0001 ,
		\u1_row_adr_reg[3]/P0001 ,
		\u2_u0_b0_last_row_reg[1]/P0001 ,
		\u2_u0_b0_last_row_reg[3]/P0001 ,
		_w4039_
	);
	LUT4 #(
		.INIT('hf531)
	) name3080 (
		\u1_row_adr_reg[0]/P0001 ,
		\u1_row_adr_reg[2]/P0001 ,
		\u2_u0_b0_last_row_reg[0]/P0001 ,
		\u2_u0_b0_last_row_reg[2]/P0001 ,
		_w4040_
	);
	LUT4 #(
		.INIT('hf531)
	) name3081 (
		\u1_row_adr_reg[3]/P0001 ,
		\u1_row_adr_reg[4]/P0001 ,
		\u2_u0_b0_last_row_reg[3]/P0001 ,
		\u2_u0_b0_last_row_reg[4]/P0001 ,
		_w4041_
	);
	LUT4 #(
		.INIT('haf23)
	) name3082 (
		\u1_row_adr_reg[7]/P0001 ,
		\u1_row_adr_reg[9]/P0001 ,
		\u2_u0_b0_last_row_reg[7]/P0001 ,
		\u2_u0_b0_last_row_reg[9]/P0001 ,
		_w4042_
	);
	LUT4 #(
		.INIT('h8000)
	) name3083 (
		_w4039_,
		_w4040_,
		_w4041_,
		_w4042_,
		_w4043_
	);
	LUT4 #(
		.INIT('h8000)
	) name3084 (
		_w4028_,
		_w4033_,
		_w4038_,
		_w4043_,
		_w4044_
	);
	LUT4 #(
		.INIT('ha521)
	) name3085 (
		\u1_row_adr_reg[0]/P0001 ,
		\u1_row_adr_reg[11]/P0001 ,
		\u2_u0_b3_last_row_reg[0]/P0001 ,
		\u2_u0_b3_last_row_reg[11]/P0001 ,
		_w4045_
	);
	LUT4 #(
		.INIT('haf23)
	) name3086 (
		\u1_row_adr_reg[11]/P0001 ,
		\u1_row_adr_reg[7]/P0001 ,
		\u2_u0_b3_last_row_reg[11]/P0001 ,
		\u2_u0_b3_last_row_reg[7]/P0001 ,
		_w4046_
	);
	LUT4 #(
		.INIT('haf23)
	) name3087 (
		\u1_row_adr_reg[12]/P0001 ,
		\u1_row_adr_reg[1]/P0001 ,
		\u2_u0_b3_last_row_reg[12]/P0001 ,
		\u2_u0_b3_last_row_reg[1]/P0001 ,
		_w4047_
	);
	LUT4 #(
		.INIT('hc4f5)
	) name3088 (
		\u1_row_adr_reg[10]/P0001 ,
		\u1_row_adr_reg[3]/P0001 ,
		\u2_u0_b3_last_row_reg[10]/P0001 ,
		\u2_u0_b3_last_row_reg[3]/P0001 ,
		_w4048_
	);
	LUT4 #(
		.INIT('h8caf)
	) name3089 (
		\u1_row_adr_reg[5]/P0001 ,
		\u1_row_adr_reg[9]/P0001 ,
		\u2_u0_b3_last_row_reg[5]/P0001 ,
		\u2_u0_b3_last_row_reg[9]/P0001 ,
		_w4049_
	);
	LUT4 #(
		.INIT('h8000)
	) name3090 (
		_w4046_,
		_w4047_,
		_w4048_,
		_w4049_,
		_w4050_
	);
	LUT4 #(
		.INIT('haf23)
	) name3091 (
		\u1_row_adr_reg[10]/P0001 ,
		\u1_row_adr_reg[5]/P0001 ,
		\u2_u0_b3_last_row_reg[10]/P0001 ,
		\u2_u0_b3_last_row_reg[5]/P0001 ,
		_w4051_
	);
	LUT4 #(
		.INIT('hc4f5)
	) name3092 (
		\u1_row_adr_reg[2]/P0001 ,
		\u1_row_adr_reg[8]/P0001 ,
		\u2_u0_b3_last_row_reg[2]/P0001 ,
		\u2_u0_b3_last_row_reg[8]/P0001 ,
		_w4052_
	);
	LUT2 #(
		.INIT('h6)
	) name3093 (
		\u1_row_adr_reg[4]/P0001 ,
		\u2_u0_b3_last_row_reg[4]/P0001 ,
		_w4053_
	);
	LUT4 #(
		.INIT('h8808)
	) name3094 (
		\u1_bank_adr_reg[0]/P0001 ,
		\u1_bank_adr_reg[1]/P0001 ,
		\u1_row_adr_reg[6]/P0001 ,
		\u2_u0_b3_last_row_reg[6]/P0001 ,
		_w4054_
	);
	LUT4 #(
		.INIT('h0800)
	) name3095 (
		_w4051_,
		_w4052_,
		_w4053_,
		_w4054_,
		_w4055_
	);
	LUT4 #(
		.INIT('hf531)
	) name3096 (
		\u1_row_adr_reg[3]/P0001 ,
		\u1_row_adr_reg[8]/P0001 ,
		\u2_u0_b3_last_row_reg[3]/P0001 ,
		\u2_u0_b3_last_row_reg[8]/P0001 ,
		_w4056_
	);
	LUT4 #(
		.INIT('h8caf)
	) name3097 (
		\u1_row_adr_reg[2]/P0001 ,
		\u1_row_adr_reg[6]/P0001 ,
		\u2_u0_b3_last_row_reg[2]/P0001 ,
		\u2_u0_b3_last_row_reg[6]/P0001 ,
		_w4057_
	);
	LUT4 #(
		.INIT('haf23)
	) name3098 (
		\u1_row_adr_reg[7]/P0001 ,
		\u1_row_adr_reg[9]/P0001 ,
		\u2_u0_b3_last_row_reg[7]/P0001 ,
		\u2_u0_b3_last_row_reg[9]/P0001 ,
		_w4058_
	);
	LUT4 #(
		.INIT('hc4f5)
	) name3099 (
		\u1_row_adr_reg[12]/P0001 ,
		\u1_row_adr_reg[1]/P0001 ,
		\u2_u0_b3_last_row_reg[12]/P0001 ,
		\u2_u0_b3_last_row_reg[1]/P0001 ,
		_w4059_
	);
	LUT4 #(
		.INIT('h8000)
	) name3100 (
		_w4056_,
		_w4057_,
		_w4058_,
		_w4059_,
		_w4060_
	);
	LUT4 #(
		.INIT('h8000)
	) name3101 (
		_w4045_,
		_w4050_,
		_w4055_,
		_w4060_,
		_w4061_
	);
	LUT4 #(
		.INIT('h0001)
	) name3102 (
		_w4008_,
		_w4027_,
		_w4044_,
		_w4061_,
		_w4062_
	);
	LUT4 #(
		.INIT('h03ab)
	) name3103 (
		_w1533_,
		_w1579_,
		_w3992_,
		_w4062_,
		_w4063_
	);
	LUT2 #(
		.INIT('h8)
	) name3104 (
		_w2401_,
		_w2563_,
		_w4064_
	);
	LUT4 #(
		.INIT('h7f00)
	) name3105 (
		_w1184_,
		_w1185_,
		_w1569_,
		_w4064_,
		_w4065_
	);
	LUT3 #(
		.INIT('h40)
	) name3106 (
		_w2389_,
		_w2566_,
		_w4065_,
		_w4066_
	);
	LUT4 #(
		.INIT('h4ccc)
	) name3107 (
		\u5_cmd_asserted_reg/NET0131 ,
		\u5_susp_sel_r_reg/NET0131 ,
		_w1100_,
		_w1102_,
		_w4067_
	);
	LUT3 #(
		.INIT('h80)
	) name3108 (
		_w1582_,
		_w1583_,
		_w2685_,
		_w4068_
	);
	LUT2 #(
		.INIT('h8)
	) name3109 (
		_w1184_,
		_w4068_,
		_w4069_
	);
	LUT2 #(
		.INIT('he)
	) name3110 (
		_w4067_,
		_w4069_,
		_w4070_
	);
	LUT3 #(
		.INIT('h2a)
	) name3111 (
		\u0_u0_csc_reg[1]/NET0131 ,
		\u0_u0_csc_reg[8]/P0001 ,
		wb_we_i_pad,
		_w4071_
	);
	LUT4 #(
		.INIT('h0100)
	) name3112 (
		_w2914_,
		_w2915_,
		_w2916_,
		_w4071_,
		_w4072_
	);
	LUT3 #(
		.INIT('h80)
	) name3113 (
		_w2907_,
		_w2912_,
		_w4072_,
		_w4073_
	);
	LUT4 #(
		.INIT('hff20)
	) name3114 (
		\u0_u1_csc_reg[1]/NET0131 ,
		_w2918_,
		_w2930_,
		_w4073_,
		_w4074_
	);
	LUT3 #(
		.INIT('h2a)
	) name3115 (
		\u0_u0_csc_reg[2]/NET0131 ,
		\u0_u0_csc_reg[8]/P0001 ,
		wb_we_i_pad,
		_w4075_
	);
	LUT4 #(
		.INIT('h0100)
	) name3116 (
		_w2914_,
		_w2915_,
		_w2916_,
		_w4075_,
		_w4076_
	);
	LUT3 #(
		.INIT('h80)
	) name3117 (
		_w2907_,
		_w2912_,
		_w4076_,
		_w4077_
	);
	LUT4 #(
		.INIT('hff20)
	) name3118 (
		\u0_u1_csc_reg[2]/NET0131 ,
		_w2918_,
		_w2930_,
		_w4077_,
		_w4078_
	);
	LUT3 #(
		.INIT('h2a)
	) name3119 (
		\u0_u0_csc_reg[3]/NET0131 ,
		\u0_u0_csc_reg[8]/P0001 ,
		wb_we_i_pad,
		_w4079_
	);
	LUT4 #(
		.INIT('h0100)
	) name3120 (
		_w2914_,
		_w2915_,
		_w2916_,
		_w4079_,
		_w4080_
	);
	LUT3 #(
		.INIT('h80)
	) name3121 (
		_w2907_,
		_w2912_,
		_w4080_,
		_w4081_
	);
	LUT4 #(
		.INIT('hff20)
	) name3122 (
		\u0_u1_csc_reg[3]/NET0131 ,
		_w2918_,
		_w2930_,
		_w4081_,
		_w4082_
	);
	LUT2 #(
		.INIT('h6)
	) name3123 (
		\u4_ps_cnt_reg[3]/NET0131 ,
		_w3847_,
		_w4083_
	);
	LUT4 #(
		.INIT('hf700)
	) name3124 (
		_w3836_,
		_w3841_,
		_w3845_,
		_w4083_,
		_w4084_
	);
	LUT2 #(
		.INIT('h4)
	) name3125 (
		\u1_sram_addr_reg[13]/P0001 ,
		\u6_wr_hold_reg/NET0131 ,
		_w4085_
	);
	LUT4 #(
		.INIT('h3777)
	) name3126 (
		_w1333_,
		_w1335_,
		_w1338_,
		_w4085_,
		_w4086_
	);
	LUT3 #(
		.INIT('he0)
	) name3127 (
		\wb_addr_i[15]_pad ,
		_w1344_,
		_w4086_,
		_w4087_
	);
	LUT4 #(
		.INIT('h8000)
	) name3128 (
		\u1_bank_adr_reg[0]/P0001 ,
		_w1333_,
		_w1335_,
		_w1338_,
		_w4088_
	);
	LUT4 #(
		.INIT('h0080)
	) name3129 (
		\u1_acs_addr_reg[13]/P0001 ,
		_w1333_,
		_w1335_,
		_w1338_,
		_w4089_
	);
	LUT2 #(
		.INIT('h1)
	) name3130 (
		_w4088_,
		_w4089_,
		_w4090_
	);
	LUT2 #(
		.INIT('hb)
	) name3131 (
		_w4087_,
		_w4090_,
		_w4091_
	);
	LUT2 #(
		.INIT('h4)
	) name3132 (
		\u1_sram_addr_reg[14]/P0001 ,
		\u6_wr_hold_reg/NET0131 ,
		_w4092_
	);
	LUT4 #(
		.INIT('h3777)
	) name3133 (
		_w1333_,
		_w1335_,
		_w1338_,
		_w4092_,
		_w4093_
	);
	LUT3 #(
		.INIT('he0)
	) name3134 (
		\wb_addr_i[16]_pad ,
		_w1344_,
		_w4093_,
		_w4094_
	);
	LUT4 #(
		.INIT('h8000)
	) name3135 (
		\u1_bank_adr_reg[1]/P0001 ,
		_w1333_,
		_w1335_,
		_w1338_,
		_w4095_
	);
	LUT4 #(
		.INIT('h0080)
	) name3136 (
		\u1_acs_addr_reg[14]/P0001 ,
		_w1333_,
		_w1335_,
		_w1338_,
		_w4096_
	);
	LUT2 #(
		.INIT('h1)
	) name3137 (
		_w4095_,
		_w4096_,
		_w4097_
	);
	LUT2 #(
		.INIT('hb)
	) name3138 (
		_w4094_,
		_w4097_,
		_w4098_
	);
	LUT4 #(
		.INIT('h404c)
	) name3139 (
		\mem_ack_r_reg/P0001 ,
		\u1_col_adr_reg[9]/P0001 ,
		\u5_wr_cycle_reg/NET0131 ,
		wb_stb_i_pad,
		_w4099_
	);
	LUT4 #(
		.INIT('h0040)
	) name3140 (
		_w1970_,
		_w1976_,
		_w3419_,
		_w3820_,
		_w4100_
	);
	LUT3 #(
		.INIT('hdc)
	) name3141 (
		_w3550_,
		_w4099_,
		_w4100_,
		_w4101_
	);
	LUT3 #(
		.INIT('hf9)
	) name3142 (
		_w996_,
		_w1056_,
		_w3889_,
		_w4102_
	);
	LUT4 #(
		.INIT('h0080)
	) name3143 (
		\u1_acs_addr_reg[16]/P0001 ,
		_w1333_,
		_w1335_,
		_w1338_,
		_w4103_
	);
	LUT2 #(
		.INIT('h4)
	) name3144 (
		\u1_sram_addr_reg[16]/P0001 ,
		\u6_wr_hold_reg/NET0131 ,
		_w4104_
	);
	LUT4 #(
		.INIT('h3777)
	) name3145 (
		_w1333_,
		_w1335_,
		_w1338_,
		_w4104_,
		_w4105_
	);
	LUT4 #(
		.INIT('hfef0)
	) name3146 (
		\wb_addr_i[18]_pad ,
		_w1344_,
		_w4103_,
		_w4105_,
		_w4106_
	);
	LUT4 #(
		.INIT('h0080)
	) name3147 (
		\u1_acs_addr_reg[17]/P0001 ,
		_w1333_,
		_w1335_,
		_w1338_,
		_w4107_
	);
	LUT2 #(
		.INIT('h4)
	) name3148 (
		\u1_sram_addr_reg[17]/P0001 ,
		\u6_wr_hold_reg/NET0131 ,
		_w4108_
	);
	LUT4 #(
		.INIT('h3777)
	) name3149 (
		_w1333_,
		_w1335_,
		_w1338_,
		_w4108_,
		_w4109_
	);
	LUT4 #(
		.INIT('hfef0)
	) name3150 (
		\wb_addr_i[19]_pad ,
		_w1344_,
		_w4107_,
		_w4109_,
		_w4110_
	);
	LUT4 #(
		.INIT('h0080)
	) name3151 (
		\u1_acs_addr_reg[18]/P0001 ,
		_w1333_,
		_w1335_,
		_w1338_,
		_w4111_
	);
	LUT2 #(
		.INIT('h4)
	) name3152 (
		\u1_sram_addr_reg[18]/P0001 ,
		\u6_wr_hold_reg/NET0131 ,
		_w4112_
	);
	LUT4 #(
		.INIT('h3777)
	) name3153 (
		_w1333_,
		_w1335_,
		_w1338_,
		_w4112_,
		_w4113_
	);
	LUT4 #(
		.INIT('hfef0)
	) name3154 (
		\wb_addr_i[20]_pad ,
		_w1344_,
		_w4111_,
		_w4113_,
		_w4114_
	);
	LUT4 #(
		.INIT('h0080)
	) name3155 (
		\u1_acs_addr_reg[19]/P0001 ,
		_w1333_,
		_w1335_,
		_w1338_,
		_w4115_
	);
	LUT2 #(
		.INIT('h4)
	) name3156 (
		\u1_sram_addr_reg[19]/P0001 ,
		\u6_wr_hold_reg/NET0131 ,
		_w4116_
	);
	LUT4 #(
		.INIT('h3777)
	) name3157 (
		_w1333_,
		_w1335_,
		_w1338_,
		_w4116_,
		_w4117_
	);
	LUT4 #(
		.INIT('hfef0)
	) name3158 (
		\wb_addr_i[21]_pad ,
		_w1344_,
		_w4115_,
		_w4117_,
		_w4118_
	);
	LUT4 #(
		.INIT('h0080)
	) name3159 (
		\u1_acs_addr_reg[21]/P0001 ,
		_w1333_,
		_w1335_,
		_w1338_,
		_w4119_
	);
	LUT2 #(
		.INIT('h4)
	) name3160 (
		\u1_sram_addr_reg[21]/P0001 ,
		\u6_wr_hold_reg/NET0131 ,
		_w4120_
	);
	LUT4 #(
		.INIT('h3777)
	) name3161 (
		_w1333_,
		_w1335_,
		_w1338_,
		_w4120_,
		_w4121_
	);
	LUT4 #(
		.INIT('hfef0)
	) name3162 (
		\wb_addr_i[23]_pad ,
		_w1344_,
		_w4119_,
		_w4121_,
		_w4122_
	);
	LUT4 #(
		.INIT('h0080)
	) name3163 (
		\u1_acs_addr_reg[22]/P0001 ,
		_w1333_,
		_w1335_,
		_w1338_,
		_w4123_
	);
	LUT2 #(
		.INIT('h4)
	) name3164 (
		\u1_sram_addr_reg[22]/P0001 ,
		\u6_wr_hold_reg/NET0131 ,
		_w4124_
	);
	LUT4 #(
		.INIT('h3777)
	) name3165 (
		_w1333_,
		_w1335_,
		_w1338_,
		_w4124_,
		_w4125_
	);
	LUT4 #(
		.INIT('hfef0)
	) name3166 (
		\wb_addr_i[24]_pad ,
		_w1344_,
		_w4123_,
		_w4125_,
		_w4126_
	);
	LUT4 #(
		.INIT('h0080)
	) name3167 (
		\u1_acs_addr_reg[23]/P0001 ,
		_w1333_,
		_w1335_,
		_w1338_,
		_w4127_
	);
	LUT2 #(
		.INIT('h4)
	) name3168 (
		\u1_sram_addr_reg[23]/P0001 ,
		\u6_wr_hold_reg/NET0131 ,
		_w4128_
	);
	LUT4 #(
		.INIT('h3777)
	) name3169 (
		_w1333_,
		_w1335_,
		_w1338_,
		_w4128_,
		_w4129_
	);
	LUT4 #(
		.INIT('hfef0)
	) name3170 (
		\wb_addr_i[25]_pad ,
		_w1344_,
		_w4127_,
		_w4129_,
		_w4130_
	);
	LUT4 #(
		.INIT('h0080)
	) name3171 (
		\u1_acs_addr_reg[15]/P0001 ,
		_w1333_,
		_w1335_,
		_w1338_,
		_w4131_
	);
	LUT2 #(
		.INIT('h4)
	) name3172 (
		\u1_sram_addr_reg[15]/P0001 ,
		\u6_wr_hold_reg/NET0131 ,
		_w4132_
	);
	LUT4 #(
		.INIT('h3777)
	) name3173 (
		_w1333_,
		_w1335_,
		_w1338_,
		_w4132_,
		_w4133_
	);
	LUT4 #(
		.INIT('hfef0)
	) name3174 (
		\wb_addr_i[17]_pad ,
		_w1344_,
		_w4131_,
		_w4133_,
		_w4134_
	);
	LUT4 #(
		.INIT('h0080)
	) name3175 (
		\u1_acs_addr_reg[20]/P0001 ,
		_w1333_,
		_w1335_,
		_w1338_,
		_w4135_
	);
	LUT2 #(
		.INIT('h4)
	) name3176 (
		\u1_sram_addr_reg[20]/P0001 ,
		\u6_wr_hold_reg/NET0131 ,
		_w4136_
	);
	LUT4 #(
		.INIT('h3777)
	) name3177 (
		_w1333_,
		_w1335_,
		_w1338_,
		_w4136_,
		_w4137_
	);
	LUT4 #(
		.INIT('hfef0)
	) name3178 (
		\wb_addr_i[22]_pad ,
		_w1344_,
		_w4135_,
		_w4137_,
		_w4138_
	);
	LUT2 #(
		.INIT('h8)
	) name3179 (
		\u1_acs_addr_reg[7]/P0001 ,
		\u1_acs_addr_reg[8]/P0001 ,
		_w4139_
	);
	LUT4 #(
		.INIT('h6ccc)
	) name3180 (
		\u1_acs_addr_reg[7]/P0001 ,
		\u1_acs_addr_reg[8]/P0001 ,
		_w3563_,
		_w3564_,
		_w4140_
	);
	LUT4 #(
		.INIT('h78f0)
	) name3181 (
		\u4_ps_cnt_reg[0]/NET0131 ,
		\u4_ps_cnt_reg[1]/NET0131 ,
		\u4_ps_cnt_reg[2]/NET0131 ,
		\u4_rfr_en_reg/NET0131 ,
		_w4141_
	);
	LUT4 #(
		.INIT('hf700)
	) name3182 (
		_w3836_,
		_w3841_,
		_w3845_,
		_w4141_,
		_w4142_
	);
	LUT4 #(
		.INIT('h78f0)
	) name3183 (
		\u4_ps_cnt_reg[3]/NET0131 ,
		\u4_ps_cnt_reg[4]/NET0131 ,
		\u4_ps_cnt_reg[5]/NET0131 ,
		_w3847_,
		_w4143_
	);
	LUT4 #(
		.INIT('hf700)
	) name3184 (
		_w3836_,
		_w3841_,
		_w3845_,
		_w4143_,
		_w4144_
	);
	LUT3 #(
		.INIT('h6a)
	) name3185 (
		\u4_ps_cnt_reg[6]/NET0131 ,
		_w3847_,
		_w3905_,
		_w4145_
	);
	LUT4 #(
		.INIT('hf700)
	) name3186 (
		_w3836_,
		_w3841_,
		_w3845_,
		_w4145_,
		_w4146_
	);
	LUT2 #(
		.INIT('h6)
	) name3187 (
		\u4_ps_cnt_reg[0]/NET0131 ,
		\u4_rfr_en_reg/NET0131 ,
		_w4147_
	);
	LUT4 #(
		.INIT('hf700)
	) name3188 (
		_w3836_,
		_w3841_,
		_w3845_,
		_w4147_,
		_w4148_
	);
	LUT3 #(
		.INIT('h6c)
	) name3189 (
		\u4_ps_cnt_reg[0]/NET0131 ,
		\u4_ps_cnt_reg[1]/NET0131 ,
		\u4_rfr_en_reg/NET0131 ,
		_w4149_
	);
	LUT4 #(
		.INIT('hf700)
	) name3190 (
		_w3836_,
		_w3841_,
		_w3845_,
		_w4149_,
		_w4150_
	);
	LUT4 #(
		.INIT('h0200)
	) name3191 (
		\u0_init_req_reg/NET0131 ,
		\u4_rfr_req_reg/NET0131 ,
		\u5_state_reg[0]/NET0131 ,
		\u5_state_reg[1]/NET0131 ,
		_w4151_
	);
	LUT2 #(
		.INIT('h8)
	) name3192 (
		_w1184_,
		_w4151_,
		_w4152_
	);
	LUT2 #(
		.INIT('h6)
	) name3193 (
		\u1_acs_addr_reg[4]/P0001 ,
		_w3563_,
		_w4153_
	);
	LUT4 #(
		.INIT('h0800)
	) name3194 (
		\mem_ack_r_reg/P0001 ,
		\u6_read_go_r1_reg/NET0131 ,
		\u6_rmw_r_reg/NET0131 ,
		wb_cyc_i_pad,
		_w4154_
	);
	LUT4 #(
		.INIT('h0444)
	) name3195 (
		\u3_u0_rd_adr_reg[0]/NET0131 ,
		wb_cyc_i_pad,
		wb_stb_i_pad,
		wb_we_i_pad,
		_w4155_
	);
	LUT4 #(
		.INIT('h8f00)
	) name3196 (
		_w1014_,
		_w1015_,
		_w4154_,
		_w4155_,
		_w4156_
	);
	LUT4 #(
		.INIT('h0444)
	) name3197 (
		\u3_u0_rd_adr_reg[3]/NET0131 ,
		wb_cyc_i_pad,
		wb_stb_i_pad,
		wb_we_i_pad,
		_w4157_
	);
	LUT4 #(
		.INIT('h7000)
	) name3198 (
		_w1014_,
		_w1015_,
		_w4154_,
		_w4157_,
		_w4158_
	);
	LUT2 #(
		.INIT('h1)
	) name3199 (
		_w4156_,
		_w4158_,
		_w4159_
	);
	LUT4 #(
		.INIT('h0888)
	) name3200 (
		\u3_u0_rd_adr_reg[1]/NET0131 ,
		wb_cyc_i_pad,
		wb_stb_i_pad,
		wb_we_i_pad,
		_w4160_
	);
	LUT4 #(
		.INIT('h8f00)
	) name3201 (
		_w1014_,
		_w1015_,
		_w4154_,
		_w4160_,
		_w4161_
	);
	LUT4 #(
		.INIT('h0888)
	) name3202 (
		\u3_u0_rd_adr_reg[0]/NET0131 ,
		wb_cyc_i_pad,
		wb_stb_i_pad,
		wb_we_i_pad,
		_w4162_
	);
	LUT4 #(
		.INIT('h7000)
	) name3203 (
		_w1014_,
		_w1015_,
		_w4154_,
		_w4162_,
		_w4163_
	);
	LUT2 #(
		.INIT('he)
	) name3204 (
		_w4161_,
		_w4163_,
		_w4164_
	);
	LUT4 #(
		.INIT('h0888)
	) name3205 (
		\u3_u0_rd_adr_reg[2]/NET0131 ,
		wb_cyc_i_pad,
		wb_stb_i_pad,
		wb_we_i_pad,
		_w4165_
	);
	LUT4 #(
		.INIT('h8f00)
	) name3206 (
		_w1014_,
		_w1015_,
		_w4154_,
		_w4165_,
		_w4166_
	);
	LUT4 #(
		.INIT('h7000)
	) name3207 (
		_w1014_,
		_w1015_,
		_w4154_,
		_w4160_,
		_w4167_
	);
	LUT2 #(
		.INIT('he)
	) name3208 (
		_w4166_,
		_w4167_,
		_w4168_
	);
	LUT4 #(
		.INIT('h0888)
	) name3209 (
		\u3_u0_rd_adr_reg[3]/NET0131 ,
		wb_cyc_i_pad,
		wb_stb_i_pad,
		wb_we_i_pad,
		_w4169_
	);
	LUT4 #(
		.INIT('h8f00)
	) name3210 (
		_w1014_,
		_w1015_,
		_w4154_,
		_w4169_,
		_w4170_
	);
	LUT4 #(
		.INIT('h7000)
	) name3211 (
		_w1014_,
		_w1015_,
		_w4154_,
		_w4165_,
		_w4171_
	);
	LUT2 #(
		.INIT('he)
	) name3212 (
		_w4170_,
		_w4171_,
		_w4172_
	);
	LUT4 #(
		.INIT('h9bdf)
	) name3213 (
		\u1_bank_adr_reg[0]/P0001 ,
		\u1_bank_adr_reg[1]/P0001 ,
		\u2_u0_bank1_open_reg/NET0131 ,
		\u2_u0_bank2_open_reg/NET0131 ,
		_w4173_
	);
	LUT4 #(
		.INIT('h67ef)
	) name3214 (
		\u1_bank_adr_reg[0]/P0001 ,
		\u1_bank_adr_reg[1]/P0001 ,
		\u2_u0_bank0_open_reg/NET0131 ,
		\u2_u0_bank3_open_reg/NET0131 ,
		_w4174_
	);
	LUT4 #(
		.INIT('h0eee)
	) name3215 (
		_w1526_,
		_w1531_,
		_w4173_,
		_w4174_,
		_w4175_
	);
	LUT3 #(
		.INIT('h10)
	) name3216 (
		_w1528_,
		_w1530_,
		_w4175_,
		_w4176_
	);
	LUT4 #(
		.INIT('h37bf)
	) name3217 (
		\u1_bank_adr_reg[0]/P0001 ,
		\u1_bank_adr_reg[1]/P0001 ,
		\u2_u1_bank2_open_reg/NET0131 ,
		\u2_u1_bank3_open_reg/NET0131 ,
		_w4177_
	);
	LUT4 #(
		.INIT('hcdef)
	) name3218 (
		\u1_bank_adr_reg[0]/P0001 ,
		\u1_bank_adr_reg[1]/P0001 ,
		\u2_u1_bank0_open_reg/NET0131 ,
		\u2_u1_bank1_open_reg/NET0131 ,
		_w4178_
	);
	LUT2 #(
		.INIT('h8)
	) name3219 (
		_w4177_,
		_w4178_,
		_w4179_
	);
	LUT4 #(
		.INIT('h00fe)
	) name3220 (
		_w1574_,
		_w1576_,
		_w1578_,
		_w4179_,
		_w4180_
	);
	LUT2 #(
		.INIT('he)
	) name3221 (
		_w4176_,
		_w4180_,
		_w4181_
	);
	LUT3 #(
		.INIT('h01)
	) name3222 (
		\u0_u0_addr_r_reg[3]/P0001 ,
		\u0_u0_addr_r_reg[5]/P0001 ,
		\u0_u0_addr_r_reg[6]/P0001 ,
		_w4182_
	);
	LUT3 #(
		.INIT('h20)
	) name3223 (
		\u0_rf_we_reg/NET0131 ,
		\u0_u0_addr_r_reg[2]/P0001 ,
		\u0_u0_addr_r_reg[4]/P0001 ,
		_w4183_
	);
	LUT2 #(
		.INIT('h8)
	) name3224 (
		_w4182_,
		_w4183_,
		_w4184_
	);
	LUT3 #(
		.INIT('h15)
	) name3225 (
		\u0_u0_csc_reg[0]/NET0131 ,
		_w4182_,
		_w4183_,
		_w4185_
	);
	LUT4 #(
		.INIT('h0020)
	) name3226 (
		\u0_rf_we_reg/NET0131 ,
		\u0_u0_addr_r_reg[2]/P0001 ,
		\u0_u0_addr_r_reg[4]/P0001 ,
		\wb_data_i[0]_pad ,
		_w4186_
	);
	LUT3 #(
		.INIT('h15)
	) name3227 (
		\u0_rst_r2_reg/NET0131 ,
		_w4182_,
		_w4186_,
		_w4187_
	);
	LUT2 #(
		.INIT('h8)
	) name3228 (
		\poc_o[3]_pad ,
		\u0_rst_r2_reg/NET0131 ,
		_w4188_
	);
	LUT2 #(
		.INIT('h8)
	) name3229 (
		\poc_o[2]_pad ,
		\u0_rst_r2_reg/NET0131 ,
		_w4189_
	);
	LUT3 #(
		.INIT('h1f)
	) name3230 (
		\poc_o[2]_pad ,
		\poc_o[3]_pad ,
		\u0_rst_r2_reg/NET0131 ,
		_w4190_
	);
	LUT3 #(
		.INIT('h4f)
	) name3231 (
		_w4185_,
		_w4187_,
		_w4190_,
		_w4191_
	);
	LUT2 #(
		.INIT('h1)
	) name3232 (
		\u0_csc_reg[2]/NET0131 ,
		\u0_csc_reg[3]/NET0131 ,
		_w4192_
	);
	LUT2 #(
		.INIT('h8)
	) name3233 (
		_w1748_,
		_w4192_,
		_w4193_
	);
	LUT4 #(
		.INIT('h2e3f)
	) name3234 (
		\u0_csc_reg[4]/NET0131 ,
		\u0_csc_reg[5]/NET0131 ,
		\u7_mc_data_ir_reg[26]/P0001 ,
		\u7_mc_data_ir_reg[2]/P0001 ,
		_w4194_
	);
	LUT3 #(
		.INIT('h20)
	) name3235 (
		\u0_csc_reg[4]/NET0131 ,
		\u0_csc_reg[5]/NET0131 ,
		\u7_mc_data_ir_reg[10]/P0001 ,
		_w4195_
	);
	LUT4 #(
		.INIT('h7757)
	) name3236 (
		_w1748_,
		_w4192_,
		_w4194_,
		_w4195_,
		_w4196_
	);
	LUT4 #(
		.INIT('h008f)
	) name3237 (
		_w1807_,
		_w1808_,
		_w4192_,
		_w4196_,
		_w4197_
	);
	LUT2 #(
		.INIT('h1)
	) name3238 (
		\wb_addr_i[5]_pad ,
		\wb_addr_i[6]_pad ,
		_w4198_
	);
	LUT3 #(
		.INIT('h01)
	) name3239 (
		\wb_addr_i[3]_pad ,
		\wb_addr_i[5]_pad ,
		\wb_addr_i[6]_pad ,
		_w4199_
	);
	LUT3 #(
		.INIT('h02)
	) name3240 (
		\u0_csr_r2_reg[2]/NET0131 ,
		\wb_addr_i[2]_pad ,
		\wb_addr_i[4]_pad ,
		_w4200_
	);
	LUT2 #(
		.INIT('h8)
	) name3241 (
		_w4199_,
		_w4200_,
		_w4201_
	);
	LUT3 #(
		.INIT('h20)
	) name3242 (
		\u0_u0_csc_reg[26]/P0001 ,
		\wb_addr_i[2]_pad ,
		\wb_addr_i[4]_pad ,
		_w4202_
	);
	LUT3 #(
		.INIT('h02)
	) name3243 (
		\wb_addr_i[3]_pad ,
		\wb_addr_i[5]_pad ,
		\wb_addr_i[6]_pad ,
		_w4203_
	);
	LUT3 #(
		.INIT('h80)
	) name3244 (
		\u0_u1_tms_reg[26]/P0001 ,
		\wb_addr_i[2]_pad ,
		\wb_addr_i[4]_pad ,
		_w4204_
	);
	LUT4 #(
		.INIT('h37bf)
	) name3245 (
		\wb_addr_i[3]_pad ,
		_w4198_,
		_w4202_,
		_w4204_,
		_w4205_
	);
	LUT3 #(
		.INIT('h20)
	) name3246 (
		\u0_u1_csc_reg[26]/P0001 ,
		\wb_addr_i[2]_pad ,
		\wb_addr_i[4]_pad ,
		_w4206_
	);
	LUT3 #(
		.INIT('h15)
	) name3247 (
		_w1748_,
		_w4203_,
		_w4206_,
		_w4207_
	);
	LUT4 #(
		.INIT('h0002)
	) name3248 (
		\wb_addr_i[2]_pad ,
		\wb_addr_i[3]_pad ,
		\wb_addr_i[5]_pad ,
		\wb_addr_i[6]_pad ,
		_w4208_
	);
	LUT2 #(
		.INIT('h8)
	) name3249 (
		\u0_u0_tms_reg[26]/P0001 ,
		\wb_addr_i[4]_pad ,
		_w4209_
	);
	LUT2 #(
		.INIT('h2)
	) name3250 (
		\poc_o[26]_pad ,
		\wb_addr_i[4]_pad ,
		_w4210_
	);
	LUT3 #(
		.INIT('h57)
	) name3251 (
		_w4208_,
		_w4209_,
		_w4210_,
		_w4211_
	);
	LUT4 #(
		.INIT('h4000)
	) name3252 (
		_w4201_,
		_w4205_,
		_w4207_,
		_w4211_,
		_w4212_
	);
	LUT2 #(
		.INIT('h1)
	) name3253 (
		_w4197_,
		_w4212_,
		_w4213_
	);
	LUT3 #(
		.INIT('h20)
	) name3254 (
		\u0_csc_reg[4]/NET0131 ,
		\u0_csc_reg[5]/NET0131 ,
		\u7_mc_data_ir_reg[11]/P0001 ,
		_w4214_
	);
	LUT3 #(
		.INIT('h10)
	) name3255 (
		\u0_csc_reg[4]/NET0131 ,
		\u0_csc_reg[5]/NET0131 ,
		\u7_mc_data_ir_reg[3]/P0001 ,
		_w4215_
	);
	LUT4 #(
		.INIT('h0eee)
	) name3256 (
		\u0_csc_reg[2]/NET0131 ,
		\u0_csc_reg[3]/NET0131 ,
		\u0_csc_reg[5]/NET0131 ,
		\u7_mc_data_ir_reg[27]/P0001 ,
		_w4216_
	);
	LUT4 #(
		.INIT('h0200)
	) name3257 (
		_w1748_,
		_w4214_,
		_w4215_,
		_w4216_,
		_w4217_
	);
	LUT4 #(
		.INIT('h007f)
	) name3258 (
		_w1791_,
		_w1792_,
		_w4193_,
		_w4217_,
		_w4218_
	);
	LUT3 #(
		.INIT('h20)
	) name3259 (
		\u0_u1_csc_reg[27]/P0001 ,
		\wb_addr_i[2]_pad ,
		\wb_addr_i[4]_pad ,
		_w4219_
	);
	LUT2 #(
		.INIT('h8)
	) name3260 (
		_w4203_,
		_w4219_,
		_w4220_
	);
	LUT3 #(
		.INIT('h20)
	) name3261 (
		\u0_u0_csc_reg[27]/P0001 ,
		\wb_addr_i[2]_pad ,
		\wb_addr_i[4]_pad ,
		_w4221_
	);
	LUT3 #(
		.INIT('h80)
	) name3262 (
		\u0_u1_tms_reg[27]/P0001 ,
		\wb_addr_i[2]_pad ,
		\wb_addr_i[4]_pad ,
		_w4222_
	);
	LUT4 #(
		.INIT('h37bf)
	) name3263 (
		\wb_addr_i[3]_pad ,
		_w4198_,
		_w4221_,
		_w4222_,
		_w4223_
	);
	LUT3 #(
		.INIT('h02)
	) name3264 (
		\u0_csr_r2_reg[3]/NET0131 ,
		\wb_addr_i[2]_pad ,
		\wb_addr_i[4]_pad ,
		_w4224_
	);
	LUT3 #(
		.INIT('h15)
	) name3265 (
		_w1748_,
		_w4199_,
		_w4224_,
		_w4225_
	);
	LUT2 #(
		.INIT('h8)
	) name3266 (
		\u0_u0_tms_reg[27]/P0001 ,
		\wb_addr_i[4]_pad ,
		_w4226_
	);
	LUT2 #(
		.INIT('h2)
	) name3267 (
		\poc_o[27]_pad ,
		\wb_addr_i[4]_pad ,
		_w4227_
	);
	LUT3 #(
		.INIT('h57)
	) name3268 (
		_w4208_,
		_w4226_,
		_w4227_,
		_w4228_
	);
	LUT4 #(
		.INIT('h4000)
	) name3269 (
		_w4220_,
		_w4223_,
		_w4225_,
		_w4228_,
		_w4229_
	);
	LUT2 #(
		.INIT('h2)
	) name3270 (
		_w4218_,
		_w4229_,
		_w4230_
	);
	LUT3 #(
		.INIT('h20)
	) name3271 (
		\u0_csc_reg[4]/NET0131 ,
		\u0_csc_reg[5]/NET0131 ,
		\u7_mc_data_ir_reg[12]/P0001 ,
		_w4231_
	);
	LUT3 #(
		.INIT('h10)
	) name3272 (
		\u0_csc_reg[4]/NET0131 ,
		\u0_csc_reg[5]/NET0131 ,
		\u7_mc_data_ir_reg[4]/P0001 ,
		_w4232_
	);
	LUT4 #(
		.INIT('h0eee)
	) name3273 (
		\u0_csc_reg[2]/NET0131 ,
		\u0_csc_reg[3]/NET0131 ,
		\u0_csc_reg[5]/NET0131 ,
		\u7_mc_data_ir_reg[28]/P0001 ,
		_w4233_
	);
	LUT4 #(
		.INIT('h0200)
	) name3274 (
		_w1748_,
		_w4231_,
		_w4232_,
		_w4233_,
		_w4234_
	);
	LUT4 #(
		.INIT('h007f)
	) name3275 (
		_w1796_,
		_w1797_,
		_w4193_,
		_w4234_,
		_w4235_
	);
	LUT3 #(
		.INIT('h20)
	) name3276 (
		\u0_u1_csc_reg[28]/P0001 ,
		\wb_addr_i[2]_pad ,
		\wb_addr_i[4]_pad ,
		_w4236_
	);
	LUT2 #(
		.INIT('h8)
	) name3277 (
		_w4203_,
		_w4236_,
		_w4237_
	);
	LUT3 #(
		.INIT('h20)
	) name3278 (
		\u0_u0_csc_reg[28]/P0001 ,
		\wb_addr_i[2]_pad ,
		\wb_addr_i[4]_pad ,
		_w4238_
	);
	LUT3 #(
		.INIT('h80)
	) name3279 (
		\u0_u1_tms_reg[28]/P0001 ,
		\wb_addr_i[2]_pad ,
		\wb_addr_i[4]_pad ,
		_w4239_
	);
	LUT4 #(
		.INIT('h37bf)
	) name3280 (
		\wb_addr_i[3]_pad ,
		_w4198_,
		_w4238_,
		_w4239_,
		_w4240_
	);
	LUT3 #(
		.INIT('h02)
	) name3281 (
		\u0_csr_r2_reg[4]/NET0131 ,
		\wb_addr_i[2]_pad ,
		\wb_addr_i[4]_pad ,
		_w4241_
	);
	LUT3 #(
		.INIT('h15)
	) name3282 (
		_w1748_,
		_w4199_,
		_w4241_,
		_w4242_
	);
	LUT2 #(
		.INIT('h8)
	) name3283 (
		\u0_u0_tms_reg[28]/P0001 ,
		\wb_addr_i[4]_pad ,
		_w4243_
	);
	LUT2 #(
		.INIT('h2)
	) name3284 (
		\poc_o[28]_pad ,
		\wb_addr_i[4]_pad ,
		_w4244_
	);
	LUT3 #(
		.INIT('h57)
	) name3285 (
		_w4208_,
		_w4243_,
		_w4244_,
		_w4245_
	);
	LUT4 #(
		.INIT('h4000)
	) name3286 (
		_w4237_,
		_w4240_,
		_w4242_,
		_w4245_,
		_w4246_
	);
	LUT2 #(
		.INIT('h2)
	) name3287 (
		_w4235_,
		_w4246_,
		_w4247_
	);
	LUT3 #(
		.INIT('h20)
	) name3288 (
		\u0_csc_reg[4]/NET0131 ,
		\u0_csc_reg[5]/NET0131 ,
		\u7_mc_data_ir_reg[13]/P0001 ,
		_w4248_
	);
	LUT3 #(
		.INIT('h10)
	) name3289 (
		\u0_csc_reg[4]/NET0131 ,
		\u0_csc_reg[5]/NET0131 ,
		\u7_mc_data_ir_reg[5]/P0001 ,
		_w4249_
	);
	LUT4 #(
		.INIT('h0eee)
	) name3290 (
		\u0_csc_reg[2]/NET0131 ,
		\u0_csc_reg[3]/NET0131 ,
		\u0_csc_reg[5]/NET0131 ,
		\u7_mc_data_ir_reg[29]/P0001 ,
		_w4250_
	);
	LUT4 #(
		.INIT('h0200)
	) name3291 (
		_w1748_,
		_w4248_,
		_w4249_,
		_w4250_,
		_w4251_
	);
	LUT4 #(
		.INIT('h007f)
	) name3292 (
		_w1788_,
		_w1789_,
		_w4193_,
		_w4251_,
		_w4252_
	);
	LUT3 #(
		.INIT('h20)
	) name3293 (
		\u0_u1_csc_reg[29]/P0001 ,
		\wb_addr_i[2]_pad ,
		\wb_addr_i[4]_pad ,
		_w4253_
	);
	LUT2 #(
		.INIT('h8)
	) name3294 (
		_w4203_,
		_w4253_,
		_w4254_
	);
	LUT3 #(
		.INIT('h20)
	) name3295 (
		\u0_u0_csc_reg[29]/P0001 ,
		\wb_addr_i[2]_pad ,
		\wb_addr_i[4]_pad ,
		_w4255_
	);
	LUT3 #(
		.INIT('h80)
	) name3296 (
		\u0_u1_tms_reg[29]/P0001 ,
		\wb_addr_i[2]_pad ,
		\wb_addr_i[4]_pad ,
		_w4256_
	);
	LUT4 #(
		.INIT('h37bf)
	) name3297 (
		\wb_addr_i[3]_pad ,
		_w4198_,
		_w4255_,
		_w4256_,
		_w4257_
	);
	LUT3 #(
		.INIT('h02)
	) name3298 (
		\u0_csr_r2_reg[5]/NET0131 ,
		\wb_addr_i[2]_pad ,
		\wb_addr_i[4]_pad ,
		_w4258_
	);
	LUT3 #(
		.INIT('h15)
	) name3299 (
		_w1748_,
		_w4199_,
		_w4258_,
		_w4259_
	);
	LUT2 #(
		.INIT('h8)
	) name3300 (
		\u0_u0_tms_reg[29]/P0001 ,
		\wb_addr_i[4]_pad ,
		_w4260_
	);
	LUT2 #(
		.INIT('h2)
	) name3301 (
		\poc_o[29]_pad ,
		\wb_addr_i[4]_pad ,
		_w4261_
	);
	LUT3 #(
		.INIT('h57)
	) name3302 (
		_w4208_,
		_w4260_,
		_w4261_,
		_w4262_
	);
	LUT4 #(
		.INIT('h4000)
	) name3303 (
		_w4254_,
		_w4257_,
		_w4259_,
		_w4262_,
		_w4263_
	);
	LUT2 #(
		.INIT('h2)
	) name3304 (
		_w4252_,
		_w4263_,
		_w4264_
	);
	LUT3 #(
		.INIT('h20)
	) name3305 (
		\u0_csc_reg[4]/NET0131 ,
		\u0_csc_reg[5]/NET0131 ,
		\u7_mc_data_ir_reg[15]/P0001 ,
		_w4265_
	);
	LUT3 #(
		.INIT('h10)
	) name3306 (
		\u0_csc_reg[4]/NET0131 ,
		\u0_csc_reg[5]/NET0131 ,
		\u7_mc_data_ir_reg[7]/P0001 ,
		_w4266_
	);
	LUT4 #(
		.INIT('h0eee)
	) name3307 (
		\u0_csc_reg[2]/NET0131 ,
		\u0_csc_reg[3]/NET0131 ,
		\u0_csc_reg[5]/NET0131 ,
		\u7_mc_data_ir_reg[31]/P0001 ,
		_w4267_
	);
	LUT4 #(
		.INIT('h0200)
	) name3308 (
		_w1748_,
		_w4265_,
		_w4266_,
		_w4267_,
		_w4268_
	);
	LUT4 #(
		.INIT('h007f)
	) name3309 (
		_w1802_,
		_w1803_,
		_w4193_,
		_w4268_,
		_w4269_
	);
	LUT3 #(
		.INIT('h20)
	) name3310 (
		\u0_u1_csc_reg[31]/P0001 ,
		\wb_addr_i[2]_pad ,
		\wb_addr_i[4]_pad ,
		_w4270_
	);
	LUT2 #(
		.INIT('h8)
	) name3311 (
		_w4203_,
		_w4270_,
		_w4271_
	);
	LUT3 #(
		.INIT('h80)
	) name3312 (
		\u0_u1_tms_reg[31]/P0001 ,
		\wb_addr_i[2]_pad ,
		\wb_addr_i[4]_pad ,
		_w4272_
	);
	LUT3 #(
		.INIT('h02)
	) name3313 (
		\u0_csr_r2_reg[7]/NET0131 ,
		\wb_addr_i[2]_pad ,
		\wb_addr_i[4]_pad ,
		_w4273_
	);
	LUT4 #(
		.INIT('h3b7f)
	) name3314 (
		\wb_addr_i[3]_pad ,
		_w4198_,
		_w4272_,
		_w4273_,
		_w4274_
	);
	LUT3 #(
		.INIT('h20)
	) name3315 (
		\u0_u0_csc_reg[31]/P0001 ,
		\wb_addr_i[2]_pad ,
		\wb_addr_i[4]_pad ,
		_w4275_
	);
	LUT3 #(
		.INIT('h15)
	) name3316 (
		_w1748_,
		_w4199_,
		_w4275_,
		_w4276_
	);
	LUT2 #(
		.INIT('h8)
	) name3317 (
		\u0_u0_tms_reg[31]/P0001 ,
		\wb_addr_i[4]_pad ,
		_w4277_
	);
	LUT2 #(
		.INIT('h2)
	) name3318 (
		\poc_o[31]_pad ,
		\wb_addr_i[4]_pad ,
		_w4278_
	);
	LUT3 #(
		.INIT('h57)
	) name3319 (
		_w4208_,
		_w4277_,
		_w4278_,
		_w4279_
	);
	LUT4 #(
		.INIT('h4000)
	) name3320 (
		_w4271_,
		_w4274_,
		_w4276_,
		_w4279_,
		_w4280_
	);
	LUT2 #(
		.INIT('h2)
	) name3321 (
		_w4269_,
		_w4280_,
		_w4281_
	);
	LUT4 #(
		.INIT('h0100)
	) name3322 (
		\u0_u0_csc_reg[1]/NET0131 ,
		\u0_u0_csc_reg[2]/NET0131 ,
		\u0_u0_csc_reg[3]/NET0131 ,
		\u0_u0_lmr_req_we_reg/NET0131 ,
		_w4282_
	);
	LUT4 #(
		.INIT('hf070)
	) name3323 (
		\u0_lmr_ack_r_reg/P0001 ,
		\u0_spec_req_cs_reg[0]/NET0131 ,
		\u0_u0_lmr_req_reg/NET0131 ,
		\u5_lmr_ack_reg/NET0131 ,
		_w4283_
	);
	LUT3 #(
		.INIT('hb8)
	) name3324 (
		\u0_u0_inited_reg/NET0131 ,
		_w4282_,
		_w4283_,
		_w4284_
	);
	LUT4 #(
		.INIT('h0100)
	) name3325 (
		\u0_u1_csc_reg[1]/NET0131 ,
		\u0_u1_csc_reg[2]/NET0131 ,
		\u0_u1_csc_reg[3]/NET0131 ,
		\u0_u1_lmr_req_we_reg/NET0131 ,
		_w4285_
	);
	LUT4 #(
		.INIT('hf070)
	) name3326 (
		\u0_lmr_ack_r_reg/P0001 ,
		\u0_spec_req_cs_reg[1]/NET0131 ,
		\u0_u1_lmr_req_reg/NET0131 ,
		\u5_lmr_ack_reg/NET0131 ,
		_w4286_
	);
	LUT3 #(
		.INIT('hb8)
	) name3327 (
		\u0_u1_inited_reg/NET0131 ,
		_w4285_,
		_w4286_,
		_w4287_
	);
	LUT3 #(
		.INIT('h20)
	) name3328 (
		\u0_csc_reg[4]/NET0131 ,
		\u0_csc_reg[5]/NET0131 ,
		\u7_mc_data_ir_reg[14]/P0001 ,
		_w4288_
	);
	LUT3 #(
		.INIT('h10)
	) name3329 (
		\u0_csc_reg[4]/NET0131 ,
		\u0_csc_reg[5]/NET0131 ,
		\u7_mc_data_ir_reg[6]/P0001 ,
		_w4289_
	);
	LUT4 #(
		.INIT('h0eee)
	) name3330 (
		\u0_csc_reg[2]/NET0131 ,
		\u0_csc_reg[3]/NET0131 ,
		\u0_csc_reg[5]/NET0131 ,
		\u7_mc_data_ir_reg[30]/P0001 ,
		_w4290_
	);
	LUT4 #(
		.INIT('h0200)
	) name3331 (
		_w1748_,
		_w4288_,
		_w4289_,
		_w4290_,
		_w4291_
	);
	LUT4 #(
		.INIT('h007f)
	) name3332 (
		_w1786_,
		_w1787_,
		_w4193_,
		_w4291_,
		_w4292_
	);
	LUT3 #(
		.INIT('h20)
	) name3333 (
		\u0_u1_csc_reg[30]/P0001 ,
		\wb_addr_i[2]_pad ,
		\wb_addr_i[4]_pad ,
		_w4293_
	);
	LUT2 #(
		.INIT('h8)
	) name3334 (
		_w4203_,
		_w4293_,
		_w4294_
	);
	LUT3 #(
		.INIT('h20)
	) name3335 (
		\u0_u0_csc_reg[30]/P0001 ,
		\wb_addr_i[2]_pad ,
		\wb_addr_i[4]_pad ,
		_w4295_
	);
	LUT3 #(
		.INIT('h80)
	) name3336 (
		\u0_u1_tms_reg[30]/P0001 ,
		\wb_addr_i[2]_pad ,
		\wb_addr_i[4]_pad ,
		_w4296_
	);
	LUT4 #(
		.INIT('h37bf)
	) name3337 (
		\wb_addr_i[3]_pad ,
		_w4198_,
		_w4295_,
		_w4296_,
		_w4297_
	);
	LUT3 #(
		.INIT('h02)
	) name3338 (
		\u0_csr_r2_reg[6]/NET0131 ,
		\wb_addr_i[2]_pad ,
		\wb_addr_i[4]_pad ,
		_w4298_
	);
	LUT3 #(
		.INIT('h15)
	) name3339 (
		_w1748_,
		_w4199_,
		_w4298_,
		_w4299_
	);
	LUT2 #(
		.INIT('h8)
	) name3340 (
		\u0_u0_tms_reg[30]/P0001 ,
		\wb_addr_i[4]_pad ,
		_w4300_
	);
	LUT2 #(
		.INIT('h2)
	) name3341 (
		\poc_o[30]_pad ,
		\wb_addr_i[4]_pad ,
		_w4301_
	);
	LUT3 #(
		.INIT('h57)
	) name3342 (
		_w4208_,
		_w4300_,
		_w4301_,
		_w4302_
	);
	LUT4 #(
		.INIT('h4000)
	) name3343 (
		_w4294_,
		_w4297_,
		_w4299_,
		_w4302_,
		_w4303_
	);
	LUT2 #(
		.INIT('h2)
	) name3344 (
		_w4292_,
		_w4303_,
		_w4304_
	);
	LUT3 #(
		.INIT('h10)
	) name3345 (
		\u0_csc_reg[4]/NET0131 ,
		\u0_csc_reg[5]/NET0131 ,
		\u7_mc_data_ir_reg[0]/P0001 ,
		_w4305_
	);
	LUT3 #(
		.INIT('h20)
	) name3346 (
		\u0_csc_reg[4]/NET0131 ,
		\u0_csc_reg[5]/NET0131 ,
		\u7_mc_data_ir_reg[8]/P0001 ,
		_w4306_
	);
	LUT4 #(
		.INIT('h0eee)
	) name3347 (
		\u0_csc_reg[2]/NET0131 ,
		\u0_csc_reg[3]/NET0131 ,
		\u0_csc_reg[5]/NET0131 ,
		\u7_mc_data_ir_reg[24]/P0001 ,
		_w4307_
	);
	LUT4 #(
		.INIT('h0200)
	) name3348 (
		_w1748_,
		_w4305_,
		_w4306_,
		_w4307_,
		_w4308_
	);
	LUT4 #(
		.INIT('h007f)
	) name3349 (
		_w1800_,
		_w1801_,
		_w4193_,
		_w4308_,
		_w4309_
	);
	LUT3 #(
		.INIT('h20)
	) name3350 (
		\u0_u1_csc_reg[24]/P0001 ,
		\wb_addr_i[2]_pad ,
		\wb_addr_i[4]_pad ,
		_w4310_
	);
	LUT2 #(
		.INIT('h8)
	) name3351 (
		_w4203_,
		_w4310_,
		_w4311_
	);
	LUT3 #(
		.INIT('h20)
	) name3352 (
		\u0_u0_csc_reg[24]/P0001 ,
		\wb_addr_i[2]_pad ,
		\wb_addr_i[4]_pad ,
		_w4312_
	);
	LUT3 #(
		.INIT('h80)
	) name3353 (
		\u0_u1_tms_reg[24]/P0001 ,
		\wb_addr_i[2]_pad ,
		\wb_addr_i[4]_pad ,
		_w4313_
	);
	LUT4 #(
		.INIT('h37bf)
	) name3354 (
		\wb_addr_i[3]_pad ,
		_w4198_,
		_w4312_,
		_w4313_,
		_w4314_
	);
	LUT3 #(
		.INIT('h02)
	) name3355 (
		\u0_csr_r2_reg[0]/NET0131 ,
		\wb_addr_i[2]_pad ,
		\wb_addr_i[4]_pad ,
		_w4315_
	);
	LUT3 #(
		.INIT('h15)
	) name3356 (
		_w1748_,
		_w4199_,
		_w4315_,
		_w4316_
	);
	LUT2 #(
		.INIT('h8)
	) name3357 (
		\u0_u0_tms_reg[24]/P0001 ,
		\wb_addr_i[4]_pad ,
		_w4317_
	);
	LUT2 #(
		.INIT('h2)
	) name3358 (
		\poc_o[24]_pad ,
		\wb_addr_i[4]_pad ,
		_w4318_
	);
	LUT3 #(
		.INIT('h57)
	) name3359 (
		_w4208_,
		_w4317_,
		_w4318_,
		_w4319_
	);
	LUT4 #(
		.INIT('h4000)
	) name3360 (
		_w4311_,
		_w4314_,
		_w4316_,
		_w4319_,
		_w4320_
	);
	LUT2 #(
		.INIT('h2)
	) name3361 (
		_w4309_,
		_w4320_,
		_w4321_
	);
	LUT3 #(
		.INIT('h10)
	) name3362 (
		\u0_csc_reg[4]/NET0131 ,
		\u0_csc_reg[5]/NET0131 ,
		\u7_mc_data_ir_reg[1]/P0001 ,
		_w4322_
	);
	LUT3 #(
		.INIT('h20)
	) name3363 (
		\u0_csc_reg[4]/NET0131 ,
		\u0_csc_reg[5]/NET0131 ,
		\u7_mc_data_ir_reg[9]/P0001 ,
		_w4323_
	);
	LUT4 #(
		.INIT('h0eee)
	) name3364 (
		\u0_csc_reg[2]/NET0131 ,
		\u0_csc_reg[3]/NET0131 ,
		\u0_csc_reg[5]/NET0131 ,
		\u7_mc_data_ir_reg[25]/P0001 ,
		_w4324_
	);
	LUT4 #(
		.INIT('h0200)
	) name3365 (
		_w1748_,
		_w4322_,
		_w4323_,
		_w4324_,
		_w4325_
	);
	LUT4 #(
		.INIT('h007f)
	) name3366 (
		_w1794_,
		_w1795_,
		_w4193_,
		_w4325_,
		_w4326_
	);
	LUT3 #(
		.INIT('h20)
	) name3367 (
		\u0_u1_csc_reg[25]/P0001 ,
		\wb_addr_i[2]_pad ,
		\wb_addr_i[4]_pad ,
		_w4327_
	);
	LUT2 #(
		.INIT('h8)
	) name3368 (
		_w4203_,
		_w4327_,
		_w4328_
	);
	LUT3 #(
		.INIT('h20)
	) name3369 (
		\u0_u0_csc_reg[25]/P0001 ,
		\wb_addr_i[2]_pad ,
		\wb_addr_i[4]_pad ,
		_w4329_
	);
	LUT3 #(
		.INIT('h80)
	) name3370 (
		\u0_u1_tms_reg[25]/P0001 ,
		\wb_addr_i[2]_pad ,
		\wb_addr_i[4]_pad ,
		_w4330_
	);
	LUT4 #(
		.INIT('h37bf)
	) name3371 (
		\wb_addr_i[3]_pad ,
		_w4198_,
		_w4329_,
		_w4330_,
		_w4331_
	);
	LUT3 #(
		.INIT('h02)
	) name3372 (
		\u0_csr_r2_reg[1]/NET0131 ,
		\wb_addr_i[2]_pad ,
		\wb_addr_i[4]_pad ,
		_w4332_
	);
	LUT3 #(
		.INIT('h15)
	) name3373 (
		_w1748_,
		_w4199_,
		_w4332_,
		_w4333_
	);
	LUT2 #(
		.INIT('h8)
	) name3374 (
		\u0_u0_tms_reg[25]/P0001 ,
		\wb_addr_i[4]_pad ,
		_w4334_
	);
	LUT2 #(
		.INIT('h2)
	) name3375 (
		\poc_o[25]_pad ,
		\wb_addr_i[4]_pad ,
		_w4335_
	);
	LUT3 #(
		.INIT('h57)
	) name3376 (
		_w4208_,
		_w4334_,
		_w4335_,
		_w4336_
	);
	LUT4 #(
		.INIT('h4000)
	) name3377 (
		_w4328_,
		_w4331_,
		_w4333_,
		_w4336_,
		_w4337_
	);
	LUT2 #(
		.INIT('h2)
	) name3378 (
		_w4326_,
		_w4337_,
		_w4338_
	);
	LUT3 #(
		.INIT('h1b)
	) name3379 (
		\u0_csc_reg[5]/NET0131 ,
		\u3_byte0_reg[1]/P0001 ,
		\u7_mc_data_ir_reg[1]/P0001 ,
		_w4339_
	);
	LUT3 #(
		.INIT('ha8)
	) name3380 (
		_w1748_,
		_w4192_,
		_w4339_,
		_w4340_
	);
	LUT4 #(
		.INIT('h8f00)
	) name3381 (
		_w1868_,
		_w1869_,
		_w4192_,
		_w4340_,
		_w4341_
	);
	LUT3 #(
		.INIT('h20)
	) name3382 (
		\u0_u1_csc_reg[1]/NET0131 ,
		\wb_addr_i[2]_pad ,
		\wb_addr_i[4]_pad ,
		_w4342_
	);
	LUT3 #(
		.INIT('h02)
	) name3383 (
		\u0_csc_mask_r_reg[1]/NET0131 ,
		\wb_addr_i[2]_pad ,
		\wb_addr_i[4]_pad ,
		_w4343_
	);
	LUT3 #(
		.INIT('h57)
	) name3384 (
		_w4203_,
		_w4342_,
		_w4343_,
		_w4344_
	);
	LUT3 #(
		.INIT('h80)
	) name3385 (
		\u0_u1_tms_reg[1]/P0001 ,
		\wb_addr_i[2]_pad ,
		\wb_addr_i[4]_pad ,
		_w4345_
	);
	LUT3 #(
		.INIT('h02)
	) name3386 (
		mc_vpen_pad_o_pad,
		\wb_addr_i[2]_pad ,
		\wb_addr_i[4]_pad ,
		_w4346_
	);
	LUT4 #(
		.INIT('h3b7f)
	) name3387 (
		\wb_addr_i[3]_pad ,
		_w4198_,
		_w4345_,
		_w4346_,
		_w4347_
	);
	LUT3 #(
		.INIT('h20)
	) name3388 (
		\u0_u0_csc_reg[1]/NET0131 ,
		\wb_addr_i[2]_pad ,
		\wb_addr_i[4]_pad ,
		_w4348_
	);
	LUT3 #(
		.INIT('h15)
	) name3389 (
		_w1748_,
		_w4199_,
		_w4348_,
		_w4349_
	);
	LUT2 #(
		.INIT('h2)
	) name3390 (
		\poc_o[1]_pad ,
		\wb_addr_i[4]_pad ,
		_w4350_
	);
	LUT2 #(
		.INIT('h8)
	) name3391 (
		\u0_u0_tms_reg[1]/P0001 ,
		\wb_addr_i[4]_pad ,
		_w4351_
	);
	LUT3 #(
		.INIT('h57)
	) name3392 (
		_w4208_,
		_w4350_,
		_w4351_,
		_w4352_
	);
	LUT4 #(
		.INIT('h8000)
	) name3393 (
		_w4344_,
		_w4347_,
		_w4349_,
		_w4352_,
		_w4353_
	);
	LUT2 #(
		.INIT('h1)
	) name3394 (
		_w4341_,
		_w4353_,
		_w4354_
	);
	LUT3 #(
		.INIT('h1b)
	) name3395 (
		\u0_csc_reg[5]/NET0131 ,
		\u3_byte0_reg[3]/P0001 ,
		\u7_mc_data_ir_reg[3]/P0001 ,
		_w4355_
	);
	LUT3 #(
		.INIT('ha8)
	) name3396 (
		_w1748_,
		_w4192_,
		_w4355_,
		_w4356_
	);
	LUT4 #(
		.INIT('h8f00)
	) name3397 (
		_w1863_,
		_w1864_,
		_w4192_,
		_w4356_,
		_w4357_
	);
	LUT3 #(
		.INIT('h02)
	) name3398 (
		\u0_csc_mask_r_reg[3]/NET0131 ,
		\wb_addr_i[2]_pad ,
		\wb_addr_i[4]_pad ,
		_w4358_
	);
	LUT3 #(
		.INIT('h20)
	) name3399 (
		\u0_u0_csc_reg[3]/NET0131 ,
		\wb_addr_i[2]_pad ,
		\wb_addr_i[4]_pad ,
		_w4359_
	);
	LUT4 #(
		.INIT('h3b7f)
	) name3400 (
		\wb_addr_i[3]_pad ,
		_w4198_,
		_w4358_,
		_w4359_,
		_w4360_
	);
	LUT3 #(
		.INIT('h80)
	) name3401 (
		\u0_u1_tms_reg[3]/P0001 ,
		\wb_addr_i[2]_pad ,
		\wb_addr_i[4]_pad ,
		_w4361_
	);
	LUT3 #(
		.INIT('h02)
	) name3402 (
		\u0_csr_r_reg[3]/NET0131 ,
		\wb_addr_i[2]_pad ,
		\wb_addr_i[4]_pad ,
		_w4362_
	);
	LUT4 #(
		.INIT('h3b7f)
	) name3403 (
		\wb_addr_i[3]_pad ,
		_w4198_,
		_w4361_,
		_w4362_,
		_w4363_
	);
	LUT3 #(
		.INIT('h20)
	) name3404 (
		\u0_u1_csc_reg[3]/NET0131 ,
		\wb_addr_i[2]_pad ,
		\wb_addr_i[4]_pad ,
		_w4364_
	);
	LUT3 #(
		.INIT('h15)
	) name3405 (
		_w1748_,
		_w4203_,
		_w4364_,
		_w4365_
	);
	LUT2 #(
		.INIT('h2)
	) name3406 (
		\poc_o[3]_pad ,
		\wb_addr_i[4]_pad ,
		_w4366_
	);
	LUT2 #(
		.INIT('h8)
	) name3407 (
		\u0_u0_tms_reg[3]/P0001 ,
		\wb_addr_i[4]_pad ,
		_w4367_
	);
	LUT3 #(
		.INIT('h57)
	) name3408 (
		_w4208_,
		_w4366_,
		_w4367_,
		_w4368_
	);
	LUT4 #(
		.INIT('h8000)
	) name3409 (
		_w4360_,
		_w4363_,
		_w4365_,
		_w4368_,
		_w4369_
	);
	LUT2 #(
		.INIT('h1)
	) name3410 (
		_w4357_,
		_w4369_,
		_w4370_
	);
	LUT3 #(
		.INIT('h1b)
	) name3411 (
		\u0_csc_reg[5]/NET0131 ,
		\u3_byte0_reg[5]/P0001 ,
		\u7_mc_data_ir_reg[5]/P0001 ,
		_w4371_
	);
	LUT3 #(
		.INIT('ha8)
	) name3412 (
		_w1748_,
		_w4192_,
		_w4371_,
		_w4372_
	);
	LUT4 #(
		.INIT('h8f00)
	) name3413 (
		_w1861_,
		_w1862_,
		_w4192_,
		_w4372_,
		_w4373_
	);
	LUT3 #(
		.INIT('h02)
	) name3414 (
		\u0_csc_mask_r_reg[5]/NET0131 ,
		\wb_addr_i[2]_pad ,
		\wb_addr_i[4]_pad ,
		_w4374_
	);
	LUT3 #(
		.INIT('h80)
	) name3415 (
		\u0_u1_tms_reg[5]/P0001 ,
		\wb_addr_i[2]_pad ,
		\wb_addr_i[4]_pad ,
		_w4375_
	);
	LUT3 #(
		.INIT('h57)
	) name3416 (
		_w4203_,
		_w4374_,
		_w4375_,
		_w4376_
	);
	LUT3 #(
		.INIT('h20)
	) name3417 (
		\u0_u1_csc_reg[5]/P0001 ,
		\wb_addr_i[2]_pad ,
		\wb_addr_i[4]_pad ,
		_w4377_
	);
	LUT3 #(
		.INIT('h02)
	) name3418 (
		\u0_csr_r_reg[5]/NET0131 ,
		\wb_addr_i[2]_pad ,
		\wb_addr_i[4]_pad ,
		_w4378_
	);
	LUT4 #(
		.INIT('h3b7f)
	) name3419 (
		\wb_addr_i[3]_pad ,
		_w4198_,
		_w4377_,
		_w4378_,
		_w4379_
	);
	LUT3 #(
		.INIT('h20)
	) name3420 (
		\u0_u0_csc_reg[5]/P0001 ,
		\wb_addr_i[2]_pad ,
		\wb_addr_i[4]_pad ,
		_w4380_
	);
	LUT3 #(
		.INIT('h15)
	) name3421 (
		_w1748_,
		_w4199_,
		_w4380_,
		_w4381_
	);
	LUT2 #(
		.INIT('h8)
	) name3422 (
		\u0_u0_tms_reg[5]/P0001 ,
		\wb_addr_i[4]_pad ,
		_w4382_
	);
	LUT2 #(
		.INIT('h2)
	) name3423 (
		\poc_o[5]_pad ,
		\wb_addr_i[4]_pad ,
		_w4383_
	);
	LUT3 #(
		.INIT('h57)
	) name3424 (
		_w4208_,
		_w4382_,
		_w4383_,
		_w4384_
	);
	LUT4 #(
		.INIT('h8000)
	) name3425 (
		_w4376_,
		_w4379_,
		_w4381_,
		_w4384_,
		_w4385_
	);
	LUT2 #(
		.INIT('h1)
	) name3426 (
		_w4373_,
		_w4385_,
		_w4386_
	);
	LUT3 #(
		.INIT('h1b)
	) name3427 (
		\u0_csc_reg[5]/NET0131 ,
		\u3_byte1_reg[1]/P0001 ,
		\u7_mc_data_ir_reg[9]/P0001 ,
		_w4387_
	);
	LUT3 #(
		.INIT('ha8)
	) name3428 (
		_w1748_,
		_w4192_,
		_w4387_,
		_w4388_
	);
	LUT4 #(
		.INIT('h8f00)
	) name3429 (
		_w1758_,
		_w1759_,
		_w4192_,
		_w4388_,
		_w4389_
	);
	LUT3 #(
		.INIT('h20)
	) name3430 (
		\u0_u1_csc_reg[9]/P0001 ,
		\wb_addr_i[2]_pad ,
		\wb_addr_i[4]_pad ,
		_w4390_
	);
	LUT3 #(
		.INIT('h80)
	) name3431 (
		\u0_u1_tms_reg[9]/P0001 ,
		\wb_addr_i[2]_pad ,
		\wb_addr_i[4]_pad ,
		_w4391_
	);
	LUT3 #(
		.INIT('h57)
	) name3432 (
		_w4203_,
		_w4390_,
		_w4391_,
		_w4392_
	);
	LUT3 #(
		.INIT('h20)
	) name3433 (
		\u0_u0_csc_reg[9]/P0001 ,
		\wb_addr_i[2]_pad ,
		\wb_addr_i[4]_pad ,
		_w4393_
	);
	LUT3 #(
		.INIT('h02)
	) name3434 (
		\u0_csc_mask_r_reg[9]/NET0131 ,
		\wb_addr_i[2]_pad ,
		\wb_addr_i[4]_pad ,
		_w4394_
	);
	LUT4 #(
		.INIT('h37bf)
	) name3435 (
		\wb_addr_i[3]_pad ,
		_w4198_,
		_w4393_,
		_w4394_,
		_w4395_
	);
	LUT3 #(
		.INIT('h02)
	) name3436 (
		\u0_csr_r_reg[9]/NET0131 ,
		\wb_addr_i[2]_pad ,
		\wb_addr_i[4]_pad ,
		_w4396_
	);
	LUT3 #(
		.INIT('h15)
	) name3437 (
		_w1748_,
		_w4199_,
		_w4396_,
		_w4397_
	);
	LUT2 #(
		.INIT('h8)
	) name3438 (
		\u0_u0_tms_reg[9]/P0001 ,
		\wb_addr_i[4]_pad ,
		_w4398_
	);
	LUT2 #(
		.INIT('h2)
	) name3439 (
		\poc_o[9]_pad ,
		\wb_addr_i[4]_pad ,
		_w4399_
	);
	LUT3 #(
		.INIT('h57)
	) name3440 (
		_w4208_,
		_w4398_,
		_w4399_,
		_w4400_
	);
	LUT4 #(
		.INIT('h8000)
	) name3441 (
		_w4392_,
		_w4395_,
		_w4397_,
		_w4400_,
		_w4401_
	);
	LUT2 #(
		.INIT('h1)
	) name3442 (
		_w4389_,
		_w4401_,
		_w4402_
	);
	LUT3 #(
		.INIT('h1b)
	) name3443 (
		\u0_csc_reg[5]/NET0131 ,
		\u3_byte0_reg[6]/P0001 ,
		\u7_mc_data_ir_reg[6]/P0001 ,
		_w4403_
	);
	LUT3 #(
		.INIT('ha8)
	) name3444 (
		_w1748_,
		_w4192_,
		_w4403_,
		_w4404_
	);
	LUT4 #(
		.INIT('h8f00)
	) name3445 (
		_w1857_,
		_w1858_,
		_w4192_,
		_w4404_,
		_w4405_
	);
	LUT3 #(
		.INIT('h20)
	) name3446 (
		\u0_u0_csc_reg[6]/P0001 ,
		\wb_addr_i[2]_pad ,
		\wb_addr_i[4]_pad ,
		_w4406_
	);
	LUT3 #(
		.INIT('h20)
	) name3447 (
		\u0_u1_csc_reg[6]/P0001 ,
		\wb_addr_i[2]_pad ,
		\wb_addr_i[4]_pad ,
		_w4407_
	);
	LUT4 #(
		.INIT('h37bf)
	) name3448 (
		\wb_addr_i[3]_pad ,
		_w4198_,
		_w4406_,
		_w4407_,
		_w4408_
	);
	LUT3 #(
		.INIT('h02)
	) name3449 (
		\u0_csc_mask_r_reg[6]/NET0131 ,
		\wb_addr_i[2]_pad ,
		\wb_addr_i[4]_pad ,
		_w4409_
	);
	LUT3 #(
		.INIT('h02)
	) name3450 (
		\u0_csr_r_reg[6]/NET0131 ,
		\wb_addr_i[2]_pad ,
		\wb_addr_i[4]_pad ,
		_w4410_
	);
	LUT4 #(
		.INIT('h3b7f)
	) name3451 (
		\wb_addr_i[3]_pad ,
		_w4198_,
		_w4409_,
		_w4410_,
		_w4411_
	);
	LUT3 #(
		.INIT('h80)
	) name3452 (
		\u0_u1_tms_reg[6]/P0001 ,
		\wb_addr_i[2]_pad ,
		\wb_addr_i[4]_pad ,
		_w4412_
	);
	LUT3 #(
		.INIT('h15)
	) name3453 (
		_w1748_,
		_w4203_,
		_w4412_,
		_w4413_
	);
	LUT2 #(
		.INIT('h8)
	) name3454 (
		\u0_u0_tms_reg[6]/P0001 ,
		\wb_addr_i[4]_pad ,
		_w4414_
	);
	LUT2 #(
		.INIT('h2)
	) name3455 (
		\poc_o[6]_pad ,
		\wb_addr_i[4]_pad ,
		_w4415_
	);
	LUT3 #(
		.INIT('h57)
	) name3456 (
		_w4208_,
		_w4414_,
		_w4415_,
		_w4416_
	);
	LUT4 #(
		.INIT('h8000)
	) name3457 (
		_w4408_,
		_w4411_,
		_w4413_,
		_w4416_,
		_w4417_
	);
	LUT2 #(
		.INIT('h1)
	) name3458 (
		_w4405_,
		_w4417_,
		_w4418_
	);
	LUT3 #(
		.INIT('h1b)
	) name3459 (
		\u0_csc_reg[5]/NET0131 ,
		\u3_byte0_reg[4]/P0001 ,
		\u7_mc_data_ir_reg[4]/P0001 ,
		_w4419_
	);
	LUT3 #(
		.INIT('ha8)
	) name3460 (
		_w1748_,
		_w4192_,
		_w4419_,
		_w4420_
	);
	LUT4 #(
		.INIT('h8f00)
	) name3461 (
		_w1852_,
		_w1853_,
		_w4192_,
		_w4420_,
		_w4421_
	);
	LUT3 #(
		.INIT('h20)
	) name3462 (
		\u0_u0_csc_reg[4]/P0001 ,
		\wb_addr_i[2]_pad ,
		\wb_addr_i[4]_pad ,
		_w4422_
	);
	LUT3 #(
		.INIT('h20)
	) name3463 (
		\u0_u1_csc_reg[4]/P0001 ,
		\wb_addr_i[2]_pad ,
		\wb_addr_i[4]_pad ,
		_w4423_
	);
	LUT4 #(
		.INIT('h37bf)
	) name3464 (
		\wb_addr_i[3]_pad ,
		_w4198_,
		_w4422_,
		_w4423_,
		_w4424_
	);
	LUT3 #(
		.INIT('h02)
	) name3465 (
		\u0_csc_mask_r_reg[4]/NET0131 ,
		\wb_addr_i[2]_pad ,
		\wb_addr_i[4]_pad ,
		_w4425_
	);
	LUT3 #(
		.INIT('h02)
	) name3466 (
		\u0_csr_r_reg[4]/NET0131 ,
		\wb_addr_i[2]_pad ,
		\wb_addr_i[4]_pad ,
		_w4426_
	);
	LUT4 #(
		.INIT('h3b7f)
	) name3467 (
		\wb_addr_i[3]_pad ,
		_w4198_,
		_w4425_,
		_w4426_,
		_w4427_
	);
	LUT3 #(
		.INIT('h80)
	) name3468 (
		\u0_u1_tms_reg[4]/P0001 ,
		\wb_addr_i[2]_pad ,
		\wb_addr_i[4]_pad ,
		_w4428_
	);
	LUT3 #(
		.INIT('h15)
	) name3469 (
		_w1748_,
		_w4203_,
		_w4428_,
		_w4429_
	);
	LUT2 #(
		.INIT('h8)
	) name3470 (
		\u0_u0_tms_reg[4]/P0001 ,
		\wb_addr_i[4]_pad ,
		_w4430_
	);
	LUT2 #(
		.INIT('h2)
	) name3471 (
		\poc_o[4]_pad ,
		\wb_addr_i[4]_pad ,
		_w4431_
	);
	LUT3 #(
		.INIT('h57)
	) name3472 (
		_w4208_,
		_w4430_,
		_w4431_,
		_w4432_
	);
	LUT4 #(
		.INIT('h8000)
	) name3473 (
		_w4424_,
		_w4427_,
		_w4429_,
		_w4432_,
		_w4433_
	);
	LUT2 #(
		.INIT('h1)
	) name3474 (
		_w4421_,
		_w4433_,
		_w4434_
	);
	LUT3 #(
		.INIT('h20)
	) name3475 (
		\u5_state_reg[42]/NET0131 ,
		\u5_state_reg[43]/NET0131 ,
		\u5_tmr2_done_reg/NET0131 ,
		_w4435_
	);
	LUT3 #(
		.INIT('h80)
	) name3476 (
		_w963_,
		_w1238_,
		_w4435_,
		_w4436_
	);
	LUT2 #(
		.INIT('h8)
	) name3477 (
		_w1063_,
		_w4436_,
		_w4437_
	);
	LUT3 #(
		.INIT('h2a)
	) name3478 (
		\u5_state_reg[45]/NET0131 ,
		_w976_,
		_w1975_,
		_w4438_
	);
	LUT3 #(
		.INIT('h10)
	) name3479 (
		_w1972_,
		_w1974_,
		_w4438_,
		_w4439_
	);
	LUT4 #(
		.INIT('h8000)
	) name3480 (
		_w1030_,
		_w2598_,
		_w2600_,
		_w3854_,
		_w4440_
	);
	LUT3 #(
		.INIT('h80)
	) name3481 (
		_w1029_,
		_w3852_,
		_w4440_,
		_w4441_
	);
	LUT4 #(
		.INIT('h8000)
	) name3482 (
		_w965_,
		_w985_,
		_w1031_,
		_w1219_,
		_w4442_
	);
	LUT2 #(
		.INIT('h8)
	) name3483 (
		_w1018_,
		_w4442_,
		_w4443_
	);
	LUT3 #(
		.INIT('hea)
	) name3484 (
		_w4439_,
		_w4441_,
		_w4443_,
		_w4444_
	);
	LUT4 #(
		.INIT('h6aaa)
	) name3485 (
		\u1_acs_addr_reg[10]/P0001 ,
		_w3563_,
		_w3564_,
		_w3565_,
		_w4445_
	);
	LUT2 #(
		.INIT('h2)
	) name3486 (
		\u0_init_ack_r_reg/P0001 ,
		\u5_state_reg[26]/NET0131 ,
		_w4446_
	);
	LUT3 #(
		.INIT('h08)
	) name3487 (
		\u0_init_ack_r_reg/P0001 ,
		\u0_spec_req_cs_reg[0]/NET0131 ,
		\u5_state_reg[26]/NET0131 ,
		_w4447_
	);
	LUT3 #(
		.INIT('h2a)
	) name3488 (
		\u0_u0_init_req_reg/NET0131 ,
		_w976_,
		_w4447_,
		_w4448_
	);
	LUT2 #(
		.INIT('h2)
	) name3489 (
		\u0_u0_init_req_we_reg/NET0131 ,
		\u0_u0_inited_reg/NET0131 ,
		_w4449_
	);
	LUT2 #(
		.INIT('h8)
	) name3490 (
		_w1531_,
		_w4449_,
		_w4450_
	);
	LUT2 #(
		.INIT('he)
	) name3491 (
		_w4448_,
		_w4450_,
		_w4451_
	);
	LUT3 #(
		.INIT('h08)
	) name3492 (
		\u0_init_ack_r_reg/P0001 ,
		\u0_spec_req_cs_reg[1]/NET0131 ,
		\u5_state_reg[26]/NET0131 ,
		_w4452_
	);
	LUT3 #(
		.INIT('h2a)
	) name3493 (
		\u0_u1_init_req_reg/NET0131 ,
		_w976_,
		_w4452_,
		_w4453_
	);
	LUT2 #(
		.INIT('h2)
	) name3494 (
		\u0_u1_init_req_we_reg/NET0131 ,
		\u0_u1_inited_reg/NET0131 ,
		_w4454_
	);
	LUT2 #(
		.INIT('h8)
	) name3495 (
		_w1577_,
		_w4454_,
		_w4455_
	);
	LUT2 #(
		.INIT('he)
	) name3496 (
		_w4453_,
		_w4455_,
		_w4456_
	);
	LUT3 #(
		.INIT('h20)
	) name3497 (
		\u5_state_reg[50]/NET0131 ,
		\u5_state_reg[51]/NET0131 ,
		\u5_tmr2_done_reg/NET0131 ,
		_w4457_
	);
	LUT2 #(
		.INIT('h8)
	) name3498 (
		_w1176_,
		_w4457_,
		_w4458_
	);
	LUT2 #(
		.INIT('h8)
	) name3499 (
		_w1174_,
		_w4458_,
		_w4459_
	);
	LUT3 #(
		.INIT('h10)
	) name3500 (
		\u0_csc_reg[4]/NET0131 ,
		\u0_csc_reg[5]/NET0131 ,
		\u3_byte2_reg[0]/P0001 ,
		_w4460_
	);
	LUT3 #(
		.INIT('h20)
	) name3501 (
		\u0_csc_reg[4]/NET0131 ,
		\u0_csc_reg[5]/NET0131 ,
		\u7_mc_data_ir_reg[0]/P0001 ,
		_w4461_
	);
	LUT4 #(
		.INIT('h0eee)
	) name3502 (
		\u0_csc_reg[2]/NET0131 ,
		\u0_csc_reg[3]/NET0131 ,
		\u0_csc_reg[5]/NET0131 ,
		\u7_mc_data_ir_reg[16]/P0001 ,
		_w4462_
	);
	LUT4 #(
		.INIT('h0200)
	) name3503 (
		_w1748_,
		_w4460_,
		_w4461_,
		_w4462_,
		_w4463_
	);
	LUT4 #(
		.INIT('h007f)
	) name3504 (
		_w1831_,
		_w1832_,
		_w4193_,
		_w4463_,
		_w4464_
	);
	LUT3 #(
		.INIT('h20)
	) name3505 (
		\u0_u1_csc_reg[16]/P0001 ,
		\wb_addr_i[2]_pad ,
		\wb_addr_i[4]_pad ,
		_w4465_
	);
	LUT3 #(
		.INIT('h15)
	) name3506 (
		_w1748_,
		_w4203_,
		_w4465_,
		_w4466_
	);
	LUT3 #(
		.INIT('h80)
	) name3507 (
		\u0_u1_tms_reg[16]/P0001 ,
		\wb_addr_i[2]_pad ,
		\wb_addr_i[4]_pad ,
		_w4467_
	);
	LUT3 #(
		.INIT('h20)
	) name3508 (
		\u0_u0_csc_reg[16]/P0001 ,
		\wb_addr_i[2]_pad ,
		\wb_addr_i[4]_pad ,
		_w4468_
	);
	LUT4 #(
		.INIT('h3b7f)
	) name3509 (
		\wb_addr_i[3]_pad ,
		_w4198_,
		_w4467_,
		_w4468_,
		_w4469_
	);
	LUT3 #(
		.INIT('hca)
	) name3510 (
		\poc_o[16]_pad ,
		\u0_u0_tms_reg[16]/P0001 ,
		\wb_addr_i[4]_pad ,
		_w4470_
	);
	LUT2 #(
		.INIT('h8)
	) name3511 (
		_w4208_,
		_w4470_,
		_w4471_
	);
	LUT3 #(
		.INIT('h08)
	) name3512 (
		_w4466_,
		_w4469_,
		_w4471_,
		_w4472_
	);
	LUT2 #(
		.INIT('h2)
	) name3513 (
		_w4464_,
		_w4472_,
		_w4473_
	);
	LUT3 #(
		.INIT('h10)
	) name3514 (
		\u0_csc_reg[4]/NET0131 ,
		\u0_csc_reg[5]/NET0131 ,
		\u3_byte2_reg[1]/P0001 ,
		_w4474_
	);
	LUT3 #(
		.INIT('h20)
	) name3515 (
		\u0_csc_reg[4]/NET0131 ,
		\u0_csc_reg[5]/NET0131 ,
		\u7_mc_data_ir_reg[1]/P0001 ,
		_w4475_
	);
	LUT4 #(
		.INIT('h0eee)
	) name3516 (
		\u0_csc_reg[2]/NET0131 ,
		\u0_csc_reg[3]/NET0131 ,
		\u0_csc_reg[5]/NET0131 ,
		\u7_mc_data_ir_reg[17]/P0001 ,
		_w4476_
	);
	LUT4 #(
		.INIT('h0200)
	) name3517 (
		_w1748_,
		_w4474_,
		_w4475_,
		_w4476_,
		_w4477_
	);
	LUT4 #(
		.INIT('h007f)
	) name3518 (
		_w1819_,
		_w1820_,
		_w4193_,
		_w4477_,
		_w4478_
	);
	LUT3 #(
		.INIT('h20)
	) name3519 (
		\u0_u1_csc_reg[17]/P0001 ,
		\wb_addr_i[2]_pad ,
		\wb_addr_i[4]_pad ,
		_w4479_
	);
	LUT3 #(
		.INIT('h15)
	) name3520 (
		_w1748_,
		_w4203_,
		_w4479_,
		_w4480_
	);
	LUT3 #(
		.INIT('h80)
	) name3521 (
		\u0_u1_tms_reg[17]/P0001 ,
		\wb_addr_i[2]_pad ,
		\wb_addr_i[4]_pad ,
		_w4481_
	);
	LUT3 #(
		.INIT('h20)
	) name3522 (
		\u0_u0_csc_reg[17]/P0001 ,
		\wb_addr_i[2]_pad ,
		\wb_addr_i[4]_pad ,
		_w4482_
	);
	LUT4 #(
		.INIT('h3b7f)
	) name3523 (
		\wb_addr_i[3]_pad ,
		_w4198_,
		_w4481_,
		_w4482_,
		_w4483_
	);
	LUT3 #(
		.INIT('hca)
	) name3524 (
		\poc_o[17]_pad ,
		\u0_u0_tms_reg[17]/P0001 ,
		\wb_addr_i[4]_pad ,
		_w4484_
	);
	LUT2 #(
		.INIT('h8)
	) name3525 (
		_w4208_,
		_w4484_,
		_w4485_
	);
	LUT3 #(
		.INIT('h08)
	) name3526 (
		_w4480_,
		_w4483_,
		_w4485_,
		_w4486_
	);
	LUT2 #(
		.INIT('h2)
	) name3527 (
		_w4478_,
		_w4486_,
		_w4487_
	);
	LUT3 #(
		.INIT('h10)
	) name3528 (
		\u0_csc_reg[4]/NET0131 ,
		\u0_csc_reg[5]/NET0131 ,
		\u3_byte2_reg[2]/P0001 ,
		_w4488_
	);
	LUT3 #(
		.INIT('h20)
	) name3529 (
		\u0_csc_reg[4]/NET0131 ,
		\u0_csc_reg[5]/NET0131 ,
		\u7_mc_data_ir_reg[2]/P0001 ,
		_w4489_
	);
	LUT4 #(
		.INIT('h0eee)
	) name3530 (
		\u0_csc_reg[2]/NET0131 ,
		\u0_csc_reg[3]/NET0131 ,
		\u0_csc_reg[5]/NET0131 ,
		\u7_mc_data_ir_reg[18]/P0001 ,
		_w4490_
	);
	LUT4 #(
		.INIT('h0200)
	) name3531 (
		_w1748_,
		_w4488_,
		_w4489_,
		_w4490_,
		_w4491_
	);
	LUT4 #(
		.INIT('h007f)
	) name3532 (
		_w1838_,
		_w1839_,
		_w4193_,
		_w4491_,
		_w4492_
	);
	LUT3 #(
		.INIT('h20)
	) name3533 (
		\u0_u1_csc_reg[18]/P0001 ,
		\wb_addr_i[2]_pad ,
		\wb_addr_i[4]_pad ,
		_w4493_
	);
	LUT3 #(
		.INIT('h15)
	) name3534 (
		_w1748_,
		_w4203_,
		_w4493_,
		_w4494_
	);
	LUT3 #(
		.INIT('h80)
	) name3535 (
		\u0_u1_tms_reg[18]/P0001 ,
		\wb_addr_i[2]_pad ,
		\wb_addr_i[4]_pad ,
		_w4495_
	);
	LUT3 #(
		.INIT('h20)
	) name3536 (
		\u0_u0_csc_reg[18]/P0001 ,
		\wb_addr_i[2]_pad ,
		\wb_addr_i[4]_pad ,
		_w4496_
	);
	LUT4 #(
		.INIT('h3b7f)
	) name3537 (
		\wb_addr_i[3]_pad ,
		_w4198_,
		_w4495_,
		_w4496_,
		_w4497_
	);
	LUT3 #(
		.INIT('hca)
	) name3538 (
		\poc_o[18]_pad ,
		\u0_u0_tms_reg[18]/P0001 ,
		\wb_addr_i[4]_pad ,
		_w4498_
	);
	LUT2 #(
		.INIT('h8)
	) name3539 (
		_w4208_,
		_w4498_,
		_w4499_
	);
	LUT3 #(
		.INIT('h08)
	) name3540 (
		_w4494_,
		_w4497_,
		_w4499_,
		_w4500_
	);
	LUT2 #(
		.INIT('h2)
	) name3541 (
		_w4492_,
		_w4500_,
		_w4501_
	);
	LUT3 #(
		.INIT('h10)
	) name3542 (
		\u0_csc_reg[4]/NET0131 ,
		\u0_csc_reg[5]/NET0131 ,
		\u3_byte2_reg[3]/P0001 ,
		_w4502_
	);
	LUT3 #(
		.INIT('h20)
	) name3543 (
		\u0_csc_reg[4]/NET0131 ,
		\u0_csc_reg[5]/NET0131 ,
		\u7_mc_data_ir_reg[3]/P0001 ,
		_w4503_
	);
	LUT4 #(
		.INIT('h0eee)
	) name3544 (
		\u0_csc_reg[2]/NET0131 ,
		\u0_csc_reg[3]/NET0131 ,
		\u0_csc_reg[5]/NET0131 ,
		\u7_mc_data_ir_reg[19]/P0001 ,
		_w4504_
	);
	LUT4 #(
		.INIT('h0200)
	) name3545 (
		_w1748_,
		_w4502_,
		_w4503_,
		_w4504_,
		_w4505_
	);
	LUT4 #(
		.INIT('h007f)
	) name3546 (
		_w1825_,
		_w1826_,
		_w4193_,
		_w4505_,
		_w4506_
	);
	LUT3 #(
		.INIT('h20)
	) name3547 (
		\u0_u1_csc_reg[19]/P0001 ,
		\wb_addr_i[2]_pad ,
		\wb_addr_i[4]_pad ,
		_w4507_
	);
	LUT3 #(
		.INIT('h15)
	) name3548 (
		_w1748_,
		_w4203_,
		_w4507_,
		_w4508_
	);
	LUT3 #(
		.INIT('h80)
	) name3549 (
		\u0_u1_tms_reg[19]/P0001 ,
		\wb_addr_i[2]_pad ,
		\wb_addr_i[4]_pad ,
		_w4509_
	);
	LUT3 #(
		.INIT('h20)
	) name3550 (
		\u0_u0_csc_reg[19]/P0001 ,
		\wb_addr_i[2]_pad ,
		\wb_addr_i[4]_pad ,
		_w4510_
	);
	LUT4 #(
		.INIT('h3b7f)
	) name3551 (
		\wb_addr_i[3]_pad ,
		_w4198_,
		_w4509_,
		_w4510_,
		_w4511_
	);
	LUT3 #(
		.INIT('hca)
	) name3552 (
		\poc_o[19]_pad ,
		\u0_u0_tms_reg[19]/P0001 ,
		\wb_addr_i[4]_pad ,
		_w4512_
	);
	LUT2 #(
		.INIT('h8)
	) name3553 (
		_w4208_,
		_w4512_,
		_w4513_
	);
	LUT3 #(
		.INIT('h08)
	) name3554 (
		_w4508_,
		_w4511_,
		_w4513_,
		_w4514_
	);
	LUT2 #(
		.INIT('h2)
	) name3555 (
		_w4506_,
		_w4514_,
		_w4515_
	);
	LUT3 #(
		.INIT('h10)
	) name3556 (
		\u0_csc_reg[4]/NET0131 ,
		\u0_csc_reg[5]/NET0131 ,
		\u3_byte2_reg[4]/P0001 ,
		_w4516_
	);
	LUT3 #(
		.INIT('h20)
	) name3557 (
		\u0_csc_reg[4]/NET0131 ,
		\u0_csc_reg[5]/NET0131 ,
		\u7_mc_data_ir_reg[4]/P0001 ,
		_w4517_
	);
	LUT4 #(
		.INIT('h0eee)
	) name3558 (
		\u0_csc_reg[2]/NET0131 ,
		\u0_csc_reg[3]/NET0131 ,
		\u0_csc_reg[5]/NET0131 ,
		\u7_mc_data_ir_reg[20]/P0001 ,
		_w4518_
	);
	LUT4 #(
		.INIT('h0200)
	) name3559 (
		_w1748_,
		_w4516_,
		_w4517_,
		_w4518_,
		_w4519_
	);
	LUT4 #(
		.INIT('h007f)
	) name3560 (
		_w1827_,
		_w1828_,
		_w4193_,
		_w4519_,
		_w4520_
	);
	LUT3 #(
		.INIT('h20)
	) name3561 (
		\u0_u1_csc_reg[20]/P0001 ,
		\wb_addr_i[2]_pad ,
		\wb_addr_i[4]_pad ,
		_w4521_
	);
	LUT3 #(
		.INIT('h15)
	) name3562 (
		_w1748_,
		_w4203_,
		_w4521_,
		_w4522_
	);
	LUT3 #(
		.INIT('h80)
	) name3563 (
		\u0_u1_tms_reg[20]/P0001 ,
		\wb_addr_i[2]_pad ,
		\wb_addr_i[4]_pad ,
		_w4523_
	);
	LUT3 #(
		.INIT('h20)
	) name3564 (
		\u0_u0_csc_reg[20]/P0001 ,
		\wb_addr_i[2]_pad ,
		\wb_addr_i[4]_pad ,
		_w4524_
	);
	LUT4 #(
		.INIT('h3b7f)
	) name3565 (
		\wb_addr_i[3]_pad ,
		_w4198_,
		_w4523_,
		_w4524_,
		_w4525_
	);
	LUT3 #(
		.INIT('hca)
	) name3566 (
		\poc_o[20]_pad ,
		\u0_u0_tms_reg[20]/P0001 ,
		\wb_addr_i[4]_pad ,
		_w4526_
	);
	LUT2 #(
		.INIT('h8)
	) name3567 (
		_w4208_,
		_w4526_,
		_w4527_
	);
	LUT3 #(
		.INIT('h08)
	) name3568 (
		_w4522_,
		_w4525_,
		_w4527_,
		_w4528_
	);
	LUT2 #(
		.INIT('h2)
	) name3569 (
		_w4520_,
		_w4528_,
		_w4529_
	);
	LUT3 #(
		.INIT('h10)
	) name3570 (
		\u0_csc_reg[4]/NET0131 ,
		\u0_csc_reg[5]/NET0131 ,
		\u3_byte2_reg[6]/P0001 ,
		_w4530_
	);
	LUT3 #(
		.INIT('h20)
	) name3571 (
		\u0_csc_reg[4]/NET0131 ,
		\u0_csc_reg[5]/NET0131 ,
		\u7_mc_data_ir_reg[6]/P0001 ,
		_w4531_
	);
	LUT4 #(
		.INIT('h0eee)
	) name3572 (
		\u0_csc_reg[2]/NET0131 ,
		\u0_csc_reg[3]/NET0131 ,
		\u0_csc_reg[5]/NET0131 ,
		\u7_mc_data_ir_reg[22]/P0001 ,
		_w4532_
	);
	LUT4 #(
		.INIT('h0200)
	) name3573 (
		_w1748_,
		_w4530_,
		_w4531_,
		_w4532_,
		_w4533_
	);
	LUT4 #(
		.INIT('h007f)
	) name3574 (
		_w1822_,
		_w1823_,
		_w4193_,
		_w4533_,
		_w4534_
	);
	LUT3 #(
		.INIT('h20)
	) name3575 (
		\u0_u1_csc_reg[22]/P0001 ,
		\wb_addr_i[2]_pad ,
		\wb_addr_i[4]_pad ,
		_w4535_
	);
	LUT3 #(
		.INIT('h15)
	) name3576 (
		_w1748_,
		_w4203_,
		_w4535_,
		_w4536_
	);
	LUT3 #(
		.INIT('h80)
	) name3577 (
		\u0_u1_tms_reg[22]/P0001 ,
		\wb_addr_i[2]_pad ,
		\wb_addr_i[4]_pad ,
		_w4537_
	);
	LUT3 #(
		.INIT('h20)
	) name3578 (
		\u0_u0_csc_reg[22]/P0001 ,
		\wb_addr_i[2]_pad ,
		\wb_addr_i[4]_pad ,
		_w4538_
	);
	LUT4 #(
		.INIT('h3b7f)
	) name3579 (
		\wb_addr_i[3]_pad ,
		_w4198_,
		_w4537_,
		_w4538_,
		_w4539_
	);
	LUT3 #(
		.INIT('hca)
	) name3580 (
		\poc_o[22]_pad ,
		\u0_u0_tms_reg[22]/P0001 ,
		\wb_addr_i[4]_pad ,
		_w4540_
	);
	LUT2 #(
		.INIT('h8)
	) name3581 (
		_w4208_,
		_w4540_,
		_w4541_
	);
	LUT3 #(
		.INIT('h08)
	) name3582 (
		_w4536_,
		_w4539_,
		_w4541_,
		_w4542_
	);
	LUT2 #(
		.INIT('h2)
	) name3583 (
		_w4534_,
		_w4542_,
		_w4543_
	);
	LUT3 #(
		.INIT('h10)
	) name3584 (
		\u0_csc_reg[4]/NET0131 ,
		\u0_csc_reg[5]/NET0131 ,
		\u3_byte2_reg[7]/P0001 ,
		_w4544_
	);
	LUT3 #(
		.INIT('h20)
	) name3585 (
		\u0_csc_reg[4]/NET0131 ,
		\u0_csc_reg[5]/NET0131 ,
		\u7_mc_data_ir_reg[7]/P0001 ,
		_w4545_
	);
	LUT4 #(
		.INIT('h0eee)
	) name3586 (
		\u0_csc_reg[2]/NET0131 ,
		\u0_csc_reg[3]/NET0131 ,
		\u0_csc_reg[5]/NET0131 ,
		\u7_mc_data_ir_reg[23]/P0001 ,
		_w4546_
	);
	LUT4 #(
		.INIT('h0200)
	) name3587 (
		_w1748_,
		_w4544_,
		_w4545_,
		_w4546_,
		_w4547_
	);
	LUT4 #(
		.INIT('h007f)
	) name3588 (
		_w1833_,
		_w1834_,
		_w4193_,
		_w4547_,
		_w4548_
	);
	LUT3 #(
		.INIT('h20)
	) name3589 (
		\u0_u1_csc_reg[23]/P0001 ,
		\wb_addr_i[2]_pad ,
		\wb_addr_i[4]_pad ,
		_w4549_
	);
	LUT3 #(
		.INIT('h15)
	) name3590 (
		_w1748_,
		_w4203_,
		_w4549_,
		_w4550_
	);
	LUT3 #(
		.INIT('h80)
	) name3591 (
		\u0_u1_tms_reg[23]/P0001 ,
		\wb_addr_i[2]_pad ,
		\wb_addr_i[4]_pad ,
		_w4551_
	);
	LUT3 #(
		.INIT('h20)
	) name3592 (
		\u0_u0_csc_reg[23]/P0001 ,
		\wb_addr_i[2]_pad ,
		\wb_addr_i[4]_pad ,
		_w4552_
	);
	LUT4 #(
		.INIT('h3b7f)
	) name3593 (
		\wb_addr_i[3]_pad ,
		_w4198_,
		_w4551_,
		_w4552_,
		_w4553_
	);
	LUT3 #(
		.INIT('hca)
	) name3594 (
		\poc_o[23]_pad ,
		\u0_u0_tms_reg[23]/P0001 ,
		\wb_addr_i[4]_pad ,
		_w4554_
	);
	LUT2 #(
		.INIT('h8)
	) name3595 (
		_w4208_,
		_w4554_,
		_w4555_
	);
	LUT3 #(
		.INIT('h08)
	) name3596 (
		_w4550_,
		_w4553_,
		_w4555_,
		_w4556_
	);
	LUT2 #(
		.INIT('h2)
	) name3597 (
		_w4548_,
		_w4556_,
		_w4557_
	);
	LUT3 #(
		.INIT('h10)
	) name3598 (
		\u0_csc_reg[4]/NET0131 ,
		\u0_csc_reg[5]/NET0131 ,
		\u3_byte2_reg[5]/P0001 ,
		_w4558_
	);
	LUT3 #(
		.INIT('h20)
	) name3599 (
		\u0_csc_reg[4]/NET0131 ,
		\u0_csc_reg[5]/NET0131 ,
		\u7_mc_data_ir_reg[5]/P0001 ,
		_w4559_
	);
	LUT4 #(
		.INIT('h0eee)
	) name3600 (
		\u0_csc_reg[2]/NET0131 ,
		\u0_csc_reg[3]/NET0131 ,
		\u0_csc_reg[5]/NET0131 ,
		\u7_mc_data_ir_reg[21]/P0001 ,
		_w4560_
	);
	LUT4 #(
		.INIT('h0200)
	) name3601 (
		_w1748_,
		_w4558_,
		_w4559_,
		_w4560_,
		_w4561_
	);
	LUT4 #(
		.INIT('h007f)
	) name3602 (
		_w1817_,
		_w1818_,
		_w4193_,
		_w4561_,
		_w4562_
	);
	LUT3 #(
		.INIT('h20)
	) name3603 (
		\u0_u1_csc_reg[21]/P0001 ,
		\wb_addr_i[2]_pad ,
		\wb_addr_i[4]_pad ,
		_w4563_
	);
	LUT3 #(
		.INIT('h15)
	) name3604 (
		_w1748_,
		_w4203_,
		_w4563_,
		_w4564_
	);
	LUT3 #(
		.INIT('h80)
	) name3605 (
		\u0_u1_tms_reg[21]/P0001 ,
		\wb_addr_i[2]_pad ,
		\wb_addr_i[4]_pad ,
		_w4565_
	);
	LUT3 #(
		.INIT('h20)
	) name3606 (
		\u0_u0_csc_reg[21]/P0001 ,
		\wb_addr_i[2]_pad ,
		\wb_addr_i[4]_pad ,
		_w4566_
	);
	LUT4 #(
		.INIT('h3b7f)
	) name3607 (
		\wb_addr_i[3]_pad ,
		_w4198_,
		_w4565_,
		_w4566_,
		_w4567_
	);
	LUT3 #(
		.INIT('hca)
	) name3608 (
		\poc_o[21]_pad ,
		\u0_u0_tms_reg[21]/P0001 ,
		\wb_addr_i[4]_pad ,
		_w4568_
	);
	LUT2 #(
		.INIT('h8)
	) name3609 (
		_w4208_,
		_w4568_,
		_w4569_
	);
	LUT3 #(
		.INIT('h08)
	) name3610 (
		_w4564_,
		_w4567_,
		_w4569_,
		_w4570_
	);
	LUT2 #(
		.INIT('h2)
	) name3611 (
		_w4562_,
		_w4570_,
		_w4571_
	);
	LUT3 #(
		.INIT('h1b)
	) name3612 (
		\u0_csc_reg[5]/NET0131 ,
		\u3_byte1_reg[3]/P0001 ,
		\u7_mc_data_ir_reg[11]/P0001 ,
		_w4572_
	);
	LUT3 #(
		.INIT('ha8)
	) name3613 (
		_w1748_,
		_w4192_,
		_w4572_,
		_w4573_
	);
	LUT4 #(
		.INIT('h8f00)
	) name3614 (
		_w1764_,
		_w1765_,
		_w4192_,
		_w4573_,
		_w4574_
	);
	LUT3 #(
		.INIT('h20)
	) name3615 (
		\u0_u1_csc_reg[11]/P0001 ,
		\wb_addr_i[2]_pad ,
		\wb_addr_i[4]_pad ,
		_w4575_
	);
	LUT3 #(
		.INIT('h15)
	) name3616 (
		_w1748_,
		_w4203_,
		_w4575_,
		_w4576_
	);
	LUT3 #(
		.INIT('h80)
	) name3617 (
		\u0_u1_tms_reg[11]/P0001 ,
		\wb_addr_i[2]_pad ,
		\wb_addr_i[4]_pad ,
		_w4577_
	);
	LUT3 #(
		.INIT('h20)
	) name3618 (
		\u0_u0_csc_reg[11]/P0001 ,
		\wb_addr_i[2]_pad ,
		\wb_addr_i[4]_pad ,
		_w4578_
	);
	LUT4 #(
		.INIT('h3b7f)
	) name3619 (
		\wb_addr_i[3]_pad ,
		_w4198_,
		_w4577_,
		_w4578_,
		_w4579_
	);
	LUT3 #(
		.INIT('hca)
	) name3620 (
		\poc_o[11]_pad ,
		\u0_u0_tms_reg[11]/P0001 ,
		\wb_addr_i[4]_pad ,
		_w4580_
	);
	LUT2 #(
		.INIT('h8)
	) name3621 (
		_w4208_,
		_w4580_,
		_w4581_
	);
	LUT3 #(
		.INIT('h08)
	) name3622 (
		_w4576_,
		_w4579_,
		_w4581_,
		_w4582_
	);
	LUT2 #(
		.INIT('h1)
	) name3623 (
		_w4574_,
		_w4582_,
		_w4583_
	);
	LUT3 #(
		.INIT('h1b)
	) name3624 (
		\u0_csc_reg[5]/NET0131 ,
		\u3_byte1_reg[4]/P0001 ,
		\u7_mc_data_ir_reg[12]/P0001 ,
		_w4584_
	);
	LUT3 #(
		.INIT('ha8)
	) name3625 (
		_w1748_,
		_w4192_,
		_w4584_,
		_w4585_
	);
	LUT4 #(
		.INIT('h8f00)
	) name3626 (
		_w1766_,
		_w1767_,
		_w4192_,
		_w4585_,
		_w4586_
	);
	LUT3 #(
		.INIT('h20)
	) name3627 (
		\u0_u1_csc_reg[12]/P0001 ,
		\wb_addr_i[2]_pad ,
		\wb_addr_i[4]_pad ,
		_w4587_
	);
	LUT3 #(
		.INIT('h15)
	) name3628 (
		_w1748_,
		_w4203_,
		_w4587_,
		_w4588_
	);
	LUT3 #(
		.INIT('h80)
	) name3629 (
		\u0_u1_tms_reg[12]/P0001 ,
		\wb_addr_i[2]_pad ,
		\wb_addr_i[4]_pad ,
		_w4589_
	);
	LUT3 #(
		.INIT('h20)
	) name3630 (
		\u0_u0_csc_reg[12]/P0001 ,
		\wb_addr_i[2]_pad ,
		\wb_addr_i[4]_pad ,
		_w4590_
	);
	LUT4 #(
		.INIT('h3b7f)
	) name3631 (
		\wb_addr_i[3]_pad ,
		_w4198_,
		_w4589_,
		_w4590_,
		_w4591_
	);
	LUT3 #(
		.INIT('hca)
	) name3632 (
		\poc_o[12]_pad ,
		\u0_u0_tms_reg[12]/P0001 ,
		\wb_addr_i[4]_pad ,
		_w4592_
	);
	LUT2 #(
		.INIT('h8)
	) name3633 (
		_w4208_,
		_w4592_,
		_w4593_
	);
	LUT3 #(
		.INIT('h08)
	) name3634 (
		_w4588_,
		_w4591_,
		_w4593_,
		_w4594_
	);
	LUT2 #(
		.INIT('h1)
	) name3635 (
		_w4586_,
		_w4594_,
		_w4595_
	);
	LUT3 #(
		.INIT('h1b)
	) name3636 (
		\u0_csc_reg[5]/NET0131 ,
		\u3_byte1_reg[6]/P0001 ,
		\u7_mc_data_ir_reg[14]/P0001 ,
		_w4596_
	);
	LUT3 #(
		.INIT('ha8)
	) name3637 (
		_w1748_,
		_w4192_,
		_w4596_,
		_w4597_
	);
	LUT4 #(
		.INIT('h8f00)
	) name3638 (
		_w1761_,
		_w1762_,
		_w4192_,
		_w4597_,
		_w4598_
	);
	LUT3 #(
		.INIT('h20)
	) name3639 (
		\u0_u1_csc_reg[14]/P0001 ,
		\wb_addr_i[2]_pad ,
		\wb_addr_i[4]_pad ,
		_w4599_
	);
	LUT3 #(
		.INIT('h15)
	) name3640 (
		_w1748_,
		_w4203_,
		_w4599_,
		_w4600_
	);
	LUT3 #(
		.INIT('h80)
	) name3641 (
		\u0_u1_tms_reg[14]/P0001 ,
		\wb_addr_i[2]_pad ,
		\wb_addr_i[4]_pad ,
		_w4601_
	);
	LUT3 #(
		.INIT('h20)
	) name3642 (
		\u0_u0_csc_reg[14]/P0001 ,
		\wb_addr_i[2]_pad ,
		\wb_addr_i[4]_pad ,
		_w4602_
	);
	LUT4 #(
		.INIT('h3b7f)
	) name3643 (
		\wb_addr_i[3]_pad ,
		_w4198_,
		_w4601_,
		_w4602_,
		_w4603_
	);
	LUT3 #(
		.INIT('hca)
	) name3644 (
		\poc_o[14]_pad ,
		\u0_u0_tms_reg[14]/P0001 ,
		\wb_addr_i[4]_pad ,
		_w4604_
	);
	LUT2 #(
		.INIT('h8)
	) name3645 (
		_w4208_,
		_w4604_,
		_w4605_
	);
	LUT3 #(
		.INIT('h08)
	) name3646 (
		_w4600_,
		_w4603_,
		_w4605_,
		_w4606_
	);
	LUT2 #(
		.INIT('h1)
	) name3647 (
		_w4598_,
		_w4606_,
		_w4607_
	);
	LUT3 #(
		.INIT('h1b)
	) name3648 (
		\u0_csc_reg[5]/NET0131 ,
		\u3_byte1_reg[7]/P0001 ,
		\u7_mc_data_ir_reg[15]/P0001 ,
		_w4608_
	);
	LUT3 #(
		.INIT('ha8)
	) name3649 (
		_w1748_,
		_w4192_,
		_w4608_,
		_w4609_
	);
	LUT4 #(
		.INIT('h8f00)
	) name3650 (
		_w1772_,
		_w1773_,
		_w4192_,
		_w4609_,
		_w4610_
	);
	LUT3 #(
		.INIT('h20)
	) name3651 (
		\u0_u1_csc_reg[15]/P0001 ,
		\wb_addr_i[2]_pad ,
		\wb_addr_i[4]_pad ,
		_w4611_
	);
	LUT3 #(
		.INIT('h15)
	) name3652 (
		_w1748_,
		_w4203_,
		_w4611_,
		_w4612_
	);
	LUT3 #(
		.INIT('h80)
	) name3653 (
		\u0_u1_tms_reg[15]/P0001 ,
		\wb_addr_i[2]_pad ,
		\wb_addr_i[4]_pad ,
		_w4613_
	);
	LUT3 #(
		.INIT('h20)
	) name3654 (
		\u0_u0_csc_reg[15]/P0001 ,
		\wb_addr_i[2]_pad ,
		\wb_addr_i[4]_pad ,
		_w4614_
	);
	LUT4 #(
		.INIT('h3b7f)
	) name3655 (
		\wb_addr_i[3]_pad ,
		_w4198_,
		_w4613_,
		_w4614_,
		_w4615_
	);
	LUT3 #(
		.INIT('hca)
	) name3656 (
		\poc_o[15]_pad ,
		\u0_u0_tms_reg[15]/P0001 ,
		\wb_addr_i[4]_pad ,
		_w4616_
	);
	LUT2 #(
		.INIT('h8)
	) name3657 (
		_w4208_,
		_w4616_,
		_w4617_
	);
	LUT3 #(
		.INIT('h08)
	) name3658 (
		_w4612_,
		_w4615_,
		_w4617_,
		_w4618_
	);
	LUT2 #(
		.INIT('h1)
	) name3659 (
		_w4610_,
		_w4618_,
		_w4619_
	);
	LUT3 #(
		.INIT('h1b)
	) name3660 (
		\u0_csc_reg[5]/NET0131 ,
		\u3_byte1_reg[5]/P0001 ,
		\u7_mc_data_ir_reg[13]/P0001 ,
		_w4620_
	);
	LUT3 #(
		.INIT('ha8)
	) name3661 (
		_w1748_,
		_w4192_,
		_w4620_,
		_w4621_
	);
	LUT4 #(
		.INIT('h8f00)
	) name3662 (
		_w1754_,
		_w1757_,
		_w4192_,
		_w4621_,
		_w4622_
	);
	LUT3 #(
		.INIT('h20)
	) name3663 (
		\u0_u1_csc_reg[13]/P0001 ,
		\wb_addr_i[2]_pad ,
		\wb_addr_i[4]_pad ,
		_w4623_
	);
	LUT3 #(
		.INIT('h15)
	) name3664 (
		_w1748_,
		_w4203_,
		_w4623_,
		_w4624_
	);
	LUT3 #(
		.INIT('h80)
	) name3665 (
		\u0_u1_tms_reg[13]/P0001 ,
		\wb_addr_i[2]_pad ,
		\wb_addr_i[4]_pad ,
		_w4625_
	);
	LUT3 #(
		.INIT('h20)
	) name3666 (
		\u0_u0_csc_reg[13]/P0001 ,
		\wb_addr_i[2]_pad ,
		\wb_addr_i[4]_pad ,
		_w4626_
	);
	LUT4 #(
		.INIT('h3b7f)
	) name3667 (
		\wb_addr_i[3]_pad ,
		_w4198_,
		_w4625_,
		_w4626_,
		_w4627_
	);
	LUT3 #(
		.INIT('hca)
	) name3668 (
		\poc_o[13]_pad ,
		\u0_u0_tms_reg[13]/P0001 ,
		\wb_addr_i[4]_pad ,
		_w4628_
	);
	LUT2 #(
		.INIT('h8)
	) name3669 (
		_w4208_,
		_w4628_,
		_w4629_
	);
	LUT3 #(
		.INIT('h08)
	) name3670 (
		_w4624_,
		_w4627_,
		_w4629_,
		_w4630_
	);
	LUT2 #(
		.INIT('h1)
	) name3671 (
		_w4622_,
		_w4630_,
		_w4631_
	);
	LUT3 #(
		.INIT('h15)
	) name3672 (
		\u0_u0_csc_reg[1]/NET0131 ,
		_w4182_,
		_w4183_,
		_w4632_
	);
	LUT4 #(
		.INIT('h0020)
	) name3673 (
		\u0_rf_we_reg/NET0131 ,
		\u0_u0_addr_r_reg[2]/P0001 ,
		\u0_u0_addr_r_reg[4]/P0001 ,
		\wb_data_i[1]_pad ,
		_w4633_
	);
	LUT3 #(
		.INIT('h15)
	) name3674 (
		\u0_rst_r2_reg/NET0131 ,
		_w4182_,
		_w4633_,
		_w4634_
	);
	LUT3 #(
		.INIT('hba)
	) name3675 (
		_w4189_,
		_w4632_,
		_w4634_,
		_w4635_
	);
	LUT3 #(
		.INIT('h15)
	) name3676 (
		\u0_u0_csc_reg[2]/NET0131 ,
		_w4182_,
		_w4183_,
		_w4636_
	);
	LUT4 #(
		.INIT('h0020)
	) name3677 (
		\u0_rf_we_reg/NET0131 ,
		\u0_u0_addr_r_reg[2]/P0001 ,
		\u0_u0_addr_r_reg[4]/P0001 ,
		\wb_data_i[2]_pad ,
		_w4637_
	);
	LUT3 #(
		.INIT('h15)
	) name3678 (
		\u0_rst_r2_reg/NET0131 ,
		_w4182_,
		_w4637_,
		_w4638_
	);
	LUT3 #(
		.INIT('hba)
	) name3679 (
		_w4188_,
		_w4636_,
		_w4638_,
		_w4639_
	);
	LUT4 #(
		.INIT('h78f0)
	) name3680 (
		\u1_acs_addr_reg[4]/P0001 ,
		\u1_acs_addr_reg[5]/P0001 ,
		\u1_acs_addr_reg[6]/P0001 ,
		_w3563_,
		_w4640_
	);
	LUT3 #(
		.INIT('h1b)
	) name3681 (
		\u0_csc_reg[5]/NET0131 ,
		\u3_byte0_reg[0]/P0001 ,
		\u7_mc_data_ir_reg[0]/P0001 ,
		_w4641_
	);
	LUT3 #(
		.INIT('ha8)
	) name3682 (
		_w1748_,
		_w4192_,
		_w4641_,
		_w4642_
	);
	LUT4 #(
		.INIT('h8f00)
	) name3683 (
		_w1847_,
		_w1848_,
		_w4192_,
		_w4642_,
		_w4643_
	);
	LUT3 #(
		.INIT('h20)
	) name3684 (
		\u0_u0_csc_reg[0]/NET0131 ,
		\wb_addr_i[2]_pad ,
		\wb_addr_i[4]_pad ,
		_w4644_
	);
	LUT3 #(
		.INIT('h02)
	) name3685 (
		\u0_csc_mask_r_reg[0]/NET0131 ,
		\wb_addr_i[2]_pad ,
		\wb_addr_i[4]_pad ,
		_w4645_
	);
	LUT4 #(
		.INIT('h37bf)
	) name3686 (
		\wb_addr_i[3]_pad ,
		_w4198_,
		_w4644_,
		_w4645_,
		_w4646_
	);
	LUT3 #(
		.INIT('h20)
	) name3687 (
		\u0_u1_csc_reg[0]/NET0131 ,
		\wb_addr_i[2]_pad ,
		\wb_addr_i[4]_pad ,
		_w4647_
	);
	LUT3 #(
		.INIT('h02)
	) name3688 (
		\u0_csr_r_reg[0]/P0001 ,
		\wb_addr_i[2]_pad ,
		\wb_addr_i[4]_pad ,
		_w4648_
	);
	LUT4 #(
		.INIT('h3b7f)
	) name3689 (
		\wb_addr_i[3]_pad ,
		_w4198_,
		_w4647_,
		_w4648_,
		_w4649_
	);
	LUT3 #(
		.INIT('h80)
	) name3690 (
		\u0_u1_tms_reg[0]/P0001 ,
		\wb_addr_i[2]_pad ,
		\wb_addr_i[4]_pad ,
		_w4650_
	);
	LUT3 #(
		.INIT('h15)
	) name3691 (
		_w1748_,
		_w4203_,
		_w4650_,
		_w4651_
	);
	LUT2 #(
		.INIT('h8)
	) name3692 (
		\u0_u0_tms_reg[0]/P0001 ,
		\wb_addr_i[4]_pad ,
		_w4652_
	);
	LUT2 #(
		.INIT('h2)
	) name3693 (
		\poc_o[0]_pad ,
		\wb_addr_i[4]_pad ,
		_w4653_
	);
	LUT3 #(
		.INIT('h57)
	) name3694 (
		_w4208_,
		_w4652_,
		_w4653_,
		_w4654_
	);
	LUT4 #(
		.INIT('h8000)
	) name3695 (
		_w4646_,
		_w4649_,
		_w4651_,
		_w4654_,
		_w4655_
	);
	LUT2 #(
		.INIT('h1)
	) name3696 (
		_w4643_,
		_w4655_,
		_w4656_
	);
	LUT3 #(
		.INIT('h1b)
	) name3697 (
		\u0_csc_reg[5]/NET0131 ,
		\u3_byte1_reg[2]/P0001 ,
		\u7_mc_data_ir_reg[10]/P0001 ,
		_w4657_
	);
	LUT3 #(
		.INIT('ha8)
	) name3698 (
		_w1748_,
		_w4192_,
		_w4657_,
		_w4658_
	);
	LUT4 #(
		.INIT('h8f00)
	) name3699 (
		_w1777_,
		_w1778_,
		_w4192_,
		_w4658_,
		_w4659_
	);
	LUT3 #(
		.INIT('h20)
	) name3700 (
		\u0_u0_csc_reg[10]/P0001 ,
		\wb_addr_i[2]_pad ,
		\wb_addr_i[4]_pad ,
		_w4660_
	);
	LUT3 #(
		.INIT('h02)
	) name3701 (
		\u0_csr_r_reg[10]/NET0131 ,
		\wb_addr_i[2]_pad ,
		\wb_addr_i[4]_pad ,
		_w4661_
	);
	LUT3 #(
		.INIT('h57)
	) name3702 (
		_w4199_,
		_w4660_,
		_w4661_,
		_w4662_
	);
	LUT3 #(
		.INIT('h20)
	) name3703 (
		\u0_u1_csc_reg[10]/P0001 ,
		\wb_addr_i[2]_pad ,
		\wb_addr_i[4]_pad ,
		_w4663_
	);
	LUT3 #(
		.INIT('h02)
	) name3704 (
		\u0_csc_mask_r_reg[10]/NET0131 ,
		\wb_addr_i[2]_pad ,
		\wb_addr_i[4]_pad ,
		_w4664_
	);
	LUT3 #(
		.INIT('h57)
	) name3705 (
		_w4203_,
		_w4663_,
		_w4664_,
		_w4665_
	);
	LUT3 #(
		.INIT('h80)
	) name3706 (
		\u0_u1_tms_reg[10]/P0001 ,
		\wb_addr_i[2]_pad ,
		\wb_addr_i[4]_pad ,
		_w4666_
	);
	LUT3 #(
		.INIT('h15)
	) name3707 (
		_w1748_,
		_w4203_,
		_w4666_,
		_w4667_
	);
	LUT2 #(
		.INIT('h8)
	) name3708 (
		\u0_u0_tms_reg[10]/P0001 ,
		\wb_addr_i[4]_pad ,
		_w4668_
	);
	LUT2 #(
		.INIT('h2)
	) name3709 (
		\poc_o[10]_pad ,
		\wb_addr_i[4]_pad ,
		_w4669_
	);
	LUT3 #(
		.INIT('h57)
	) name3710 (
		_w4208_,
		_w4668_,
		_w4669_,
		_w4670_
	);
	LUT4 #(
		.INIT('h8000)
	) name3711 (
		_w4662_,
		_w4665_,
		_w4667_,
		_w4670_,
		_w4671_
	);
	LUT2 #(
		.INIT('h1)
	) name3712 (
		_w4659_,
		_w4671_,
		_w4672_
	);
	LUT3 #(
		.INIT('h1b)
	) name3713 (
		\u0_csc_reg[5]/NET0131 ,
		\u3_byte0_reg[2]/P0001 ,
		\u7_mc_data_ir_reg[2]/P0001 ,
		_w4673_
	);
	LUT3 #(
		.INIT('ha8)
	) name3714 (
		_w1748_,
		_w4192_,
		_w4673_,
		_w4674_
	);
	LUT4 #(
		.INIT('h8f00)
	) name3715 (
		_w1849_,
		_w1850_,
		_w4192_,
		_w4674_,
		_w4675_
	);
	LUT3 #(
		.INIT('h02)
	) name3716 (
		\u0_csr_r_reg[2]/NET0131 ,
		\wb_addr_i[2]_pad ,
		\wb_addr_i[4]_pad ,
		_w4676_
	);
	LUT3 #(
		.INIT('h20)
	) name3717 (
		\u0_u0_csc_reg[2]/NET0131 ,
		\wb_addr_i[2]_pad ,
		\wb_addr_i[4]_pad ,
		_w4677_
	);
	LUT3 #(
		.INIT('h57)
	) name3718 (
		_w4199_,
		_w4676_,
		_w4677_,
		_w4678_
	);
	LUT3 #(
		.INIT('h80)
	) name3719 (
		\u0_u1_tms_reg[2]/P0001 ,
		\wb_addr_i[2]_pad ,
		\wb_addr_i[4]_pad ,
		_w4679_
	);
	LUT3 #(
		.INIT('h02)
	) name3720 (
		\u0_csc_mask_r_reg[2]/NET0131 ,
		\wb_addr_i[2]_pad ,
		\wb_addr_i[4]_pad ,
		_w4680_
	);
	LUT3 #(
		.INIT('h57)
	) name3721 (
		_w4203_,
		_w4679_,
		_w4680_,
		_w4681_
	);
	LUT3 #(
		.INIT('h20)
	) name3722 (
		\u0_u1_csc_reg[2]/NET0131 ,
		\wb_addr_i[2]_pad ,
		\wb_addr_i[4]_pad ,
		_w4682_
	);
	LUT3 #(
		.INIT('h15)
	) name3723 (
		_w1748_,
		_w4203_,
		_w4682_,
		_w4683_
	);
	LUT2 #(
		.INIT('h8)
	) name3724 (
		\u0_u0_tms_reg[2]/P0001 ,
		\wb_addr_i[4]_pad ,
		_w4684_
	);
	LUT2 #(
		.INIT('h2)
	) name3725 (
		\poc_o[2]_pad ,
		\wb_addr_i[4]_pad ,
		_w4685_
	);
	LUT3 #(
		.INIT('h57)
	) name3726 (
		_w4208_,
		_w4684_,
		_w4685_,
		_w4686_
	);
	LUT4 #(
		.INIT('h8000)
	) name3727 (
		_w4678_,
		_w4681_,
		_w4683_,
		_w4686_,
		_w4687_
	);
	LUT2 #(
		.INIT('h1)
	) name3728 (
		_w4675_,
		_w4687_,
		_w4688_
	);
	LUT3 #(
		.INIT('h1b)
	) name3729 (
		\u0_csc_reg[5]/NET0131 ,
		\u3_byte0_reg[7]/P0001 ,
		\u7_mc_data_ir_reg[7]/P0001 ,
		_w4689_
	);
	LUT3 #(
		.INIT('ha8)
	) name3730 (
		_w1748_,
		_w4192_,
		_w4689_,
		_w4690_
	);
	LUT4 #(
		.INIT('h8f00)
	) name3731 (
		_w1855_,
		_w1856_,
		_w4192_,
		_w4690_,
		_w4691_
	);
	LUT3 #(
		.INIT('h20)
	) name3732 (
		\u0_u0_csc_reg[7]/P0001 ,
		\wb_addr_i[2]_pad ,
		\wb_addr_i[4]_pad ,
		_w4692_
	);
	LUT3 #(
		.INIT('h02)
	) name3733 (
		\u0_csc_mask_r_reg[7]/NET0131 ,
		\wb_addr_i[2]_pad ,
		\wb_addr_i[4]_pad ,
		_w4693_
	);
	LUT4 #(
		.INIT('h37bf)
	) name3734 (
		\wb_addr_i[3]_pad ,
		_w4198_,
		_w4692_,
		_w4693_,
		_w4694_
	);
	LUT3 #(
		.INIT('h20)
	) name3735 (
		\u0_u1_csc_reg[7]/P0001 ,
		\wb_addr_i[2]_pad ,
		\wb_addr_i[4]_pad ,
		_w4695_
	);
	LUT3 #(
		.INIT('h02)
	) name3736 (
		\u0_csr_r_reg[7]/NET0131 ,
		\wb_addr_i[2]_pad ,
		\wb_addr_i[4]_pad ,
		_w4696_
	);
	LUT4 #(
		.INIT('h3b7f)
	) name3737 (
		\wb_addr_i[3]_pad ,
		_w4198_,
		_w4695_,
		_w4696_,
		_w4697_
	);
	LUT3 #(
		.INIT('h80)
	) name3738 (
		\u0_u1_tms_reg[7]/P0001 ,
		\wb_addr_i[2]_pad ,
		\wb_addr_i[4]_pad ,
		_w4698_
	);
	LUT3 #(
		.INIT('h15)
	) name3739 (
		_w1748_,
		_w4203_,
		_w4698_,
		_w4699_
	);
	LUT2 #(
		.INIT('h8)
	) name3740 (
		\u0_u0_tms_reg[7]/P0001 ,
		\wb_addr_i[4]_pad ,
		_w4700_
	);
	LUT2 #(
		.INIT('h2)
	) name3741 (
		\poc_o[7]_pad ,
		\wb_addr_i[4]_pad ,
		_w4701_
	);
	LUT3 #(
		.INIT('h57)
	) name3742 (
		_w4208_,
		_w4700_,
		_w4701_,
		_w4702_
	);
	LUT4 #(
		.INIT('h8000)
	) name3743 (
		_w4694_,
		_w4697_,
		_w4699_,
		_w4702_,
		_w4703_
	);
	LUT2 #(
		.INIT('h1)
	) name3744 (
		_w4691_,
		_w4703_,
		_w4704_
	);
	LUT3 #(
		.INIT('h1b)
	) name3745 (
		\u0_csc_reg[5]/NET0131 ,
		\u3_byte1_reg[0]/P0001 ,
		\u7_mc_data_ir_reg[8]/P0001 ,
		_w4705_
	);
	LUT3 #(
		.INIT('ha8)
	) name3746 (
		_w1748_,
		_w4192_,
		_w4705_,
		_w4706_
	);
	LUT4 #(
		.INIT('h8f00)
	) name3747 (
		_w1770_,
		_w1771_,
		_w4192_,
		_w4706_,
		_w4707_
	);
	LUT3 #(
		.INIT('h20)
	) name3748 (
		\u0_u0_csc_reg[8]/P0001 ,
		\wb_addr_i[2]_pad ,
		\wb_addr_i[4]_pad ,
		_w4708_
	);
	LUT3 #(
		.INIT('h02)
	) name3749 (
		\u0_csr_r_reg[8]/NET0131 ,
		\wb_addr_i[2]_pad ,
		\wb_addr_i[4]_pad ,
		_w4709_
	);
	LUT3 #(
		.INIT('h57)
	) name3750 (
		_w4199_,
		_w4708_,
		_w4709_,
		_w4710_
	);
	LUT3 #(
		.INIT('h20)
	) name3751 (
		\u0_u1_csc_reg[8]/P0001 ,
		\wb_addr_i[2]_pad ,
		\wb_addr_i[4]_pad ,
		_w4711_
	);
	LUT3 #(
		.INIT('h02)
	) name3752 (
		\u0_csc_mask_r_reg[8]/NET0131 ,
		\wb_addr_i[2]_pad ,
		\wb_addr_i[4]_pad ,
		_w4712_
	);
	LUT3 #(
		.INIT('h57)
	) name3753 (
		_w4203_,
		_w4711_,
		_w4712_,
		_w4713_
	);
	LUT3 #(
		.INIT('h80)
	) name3754 (
		\u0_u1_tms_reg[8]/P0001 ,
		\wb_addr_i[2]_pad ,
		\wb_addr_i[4]_pad ,
		_w4714_
	);
	LUT3 #(
		.INIT('h15)
	) name3755 (
		_w1748_,
		_w4203_,
		_w4714_,
		_w4715_
	);
	LUT2 #(
		.INIT('h8)
	) name3756 (
		\u0_u0_tms_reg[8]/P0001 ,
		\wb_addr_i[4]_pad ,
		_w4716_
	);
	LUT2 #(
		.INIT('h2)
	) name3757 (
		\poc_o[8]_pad ,
		\wb_addr_i[4]_pad ,
		_w4717_
	);
	LUT3 #(
		.INIT('h57)
	) name3758 (
		_w4208_,
		_w4716_,
		_w4717_,
		_w4718_
	);
	LUT4 #(
		.INIT('h8000)
	) name3759 (
		_w4710_,
		_w4713_,
		_w4715_,
		_w4718_,
		_w4719_
	);
	LUT2 #(
		.INIT('h1)
	) name3760 (
		_w4707_,
		_w4719_,
		_w4720_
	);
	LUT4 #(
		.INIT('h2000)
	) name3761 (
		\u0_rf_we_reg/NET0131 ,
		\u0_u0_addr_r_reg[2]/P0001 ,
		\u0_u0_addr_r_reg[4]/P0001 ,
		\wb_data_i[5]_pad ,
		_w4721_
	);
	LUT3 #(
		.INIT('h40)
	) name3762 (
		\u0_rst_r2_reg/NET0131 ,
		_w4182_,
		_w4721_,
		_w4722_
	);
	LUT2 #(
		.INIT('h4)
	) name3763 (
		\u0_rst_r2_reg/NET0131 ,
		\u0_u0_csc_reg[5]/P0001 ,
		_w4723_
	);
	LUT3 #(
		.INIT('h70)
	) name3764 (
		_w4182_,
		_w4183_,
		_w4723_,
		_w4724_
	);
	LUT2 #(
		.INIT('h8)
	) name3765 (
		\poc_o[1]_pad ,
		\u0_rst_r2_reg/NET0131 ,
		_w4725_
	);
	LUT3 #(
		.INIT('hfe)
	) name3766 (
		_w4722_,
		_w4724_,
		_w4725_,
		_w4726_
	);
	LUT4 #(
		.INIT('h2000)
	) name3767 (
		\u0_rf_we_reg/NET0131 ,
		\u0_u0_addr_r_reg[2]/P0001 ,
		\u0_u0_addr_r_reg[4]/P0001 ,
		\wb_data_i[4]_pad ,
		_w4727_
	);
	LUT3 #(
		.INIT('h40)
	) name3768 (
		\u0_rst_r2_reg/NET0131 ,
		_w4182_,
		_w4727_,
		_w4728_
	);
	LUT2 #(
		.INIT('h4)
	) name3769 (
		\u0_rst_r2_reg/NET0131 ,
		\u0_u0_csc_reg[4]/P0001 ,
		_w4729_
	);
	LUT3 #(
		.INIT('h70)
	) name3770 (
		_w4182_,
		_w4183_,
		_w4729_,
		_w4730_
	);
	LUT2 #(
		.INIT('h8)
	) name3771 (
		\poc_o[0]_pad ,
		\u0_rst_r2_reg/NET0131 ,
		_w4731_
	);
	LUT3 #(
		.INIT('hfe)
	) name3772 (
		_w4728_,
		_w4730_,
		_w4731_,
		_w4732_
	);
	LUT3 #(
		.INIT('h2a)
	) name3773 (
		\u5_state_reg[45]/NET0131 ,
		_w976_,
		_w1971_,
		_w4733_
	);
	LUT3 #(
		.INIT('h40)
	) name3774 (
		_w1970_,
		_w1976_,
		_w4733_,
		_w4734_
	);
	LUT3 #(
		.INIT('h15)
	) name3775 (
		\u0_u0_csc_reg[11]/P0001 ,
		_w4182_,
		_w4183_,
		_w4735_
	);
	LUT4 #(
		.INIT('h0020)
	) name3776 (
		\u0_rf_we_reg/NET0131 ,
		\u0_u0_addr_r_reg[2]/P0001 ,
		\u0_u0_addr_r_reg[4]/P0001 ,
		\wb_data_i[11]_pad ,
		_w4736_
	);
	LUT3 #(
		.INIT('h15)
	) name3777 (
		\u0_rst_r2_reg/NET0131 ,
		_w4182_,
		_w4736_,
		_w4737_
	);
	LUT2 #(
		.INIT('h4)
	) name3778 (
		_w4735_,
		_w4737_,
		_w4738_
	);
	LUT3 #(
		.INIT('h15)
	) name3779 (
		\u0_u0_csc_reg[12]/P0001 ,
		_w4182_,
		_w4183_,
		_w4739_
	);
	LUT4 #(
		.INIT('h0020)
	) name3780 (
		\u0_rf_we_reg/NET0131 ,
		\u0_u0_addr_r_reg[2]/P0001 ,
		\u0_u0_addr_r_reg[4]/P0001 ,
		\wb_data_i[12]_pad ,
		_w4740_
	);
	LUT3 #(
		.INIT('h15)
	) name3781 (
		\u0_rst_r2_reg/NET0131 ,
		_w4182_,
		_w4740_,
		_w4741_
	);
	LUT2 #(
		.INIT('h4)
	) name3782 (
		_w4739_,
		_w4741_,
		_w4742_
	);
	LUT3 #(
		.INIT('h02)
	) name3783 (
		\u0_u0_addr_r_reg[3]/P0001 ,
		\u0_u0_addr_r_reg[5]/P0001 ,
		\u0_u0_addr_r_reg[6]/P0001 ,
		_w4743_
	);
	LUT3 #(
		.INIT('h80)
	) name3784 (
		\u0_rf_we_reg/NET0131 ,
		\u0_u0_addr_r_reg[2]/P0001 ,
		\u0_u0_addr_r_reg[4]/P0001 ,
		_w4744_
	);
	LUT2 #(
		.INIT('h8)
	) name3785 (
		_w4743_,
		_w4744_,
		_w4745_
	);
	LUT3 #(
		.INIT('h15)
	) name3786 (
		\u0_u1_tms_reg[19]/P0001 ,
		_w4743_,
		_w4744_,
		_w4746_
	);
	LUT4 #(
		.INIT('h0080)
	) name3787 (
		\u0_rf_we_reg/NET0131 ,
		\u0_u0_addr_r_reg[2]/P0001 ,
		\u0_u0_addr_r_reg[4]/P0001 ,
		\wb_data_i[19]_pad ,
		_w4747_
	);
	LUT3 #(
		.INIT('h15)
	) name3788 (
		\u0_rst_r2_reg/NET0131 ,
		_w4743_,
		_w4747_,
		_w4748_
	);
	LUT2 #(
		.INIT('h4)
	) name3789 (
		_w4746_,
		_w4748_,
		_w4749_
	);
	LUT3 #(
		.INIT('h15)
	) name3790 (
		\u0_u0_csc_reg[13]/P0001 ,
		_w4182_,
		_w4183_,
		_w4750_
	);
	LUT4 #(
		.INIT('h0020)
	) name3791 (
		\u0_rf_we_reg/NET0131 ,
		\u0_u0_addr_r_reg[2]/P0001 ,
		\u0_u0_addr_r_reg[4]/P0001 ,
		\wb_data_i[13]_pad ,
		_w4751_
	);
	LUT3 #(
		.INIT('h15)
	) name3792 (
		\u0_rst_r2_reg/NET0131 ,
		_w4182_,
		_w4751_,
		_w4752_
	);
	LUT2 #(
		.INIT('h4)
	) name3793 (
		_w4750_,
		_w4752_,
		_w4753_
	);
	LUT3 #(
		.INIT('h15)
	) name3794 (
		\u0_u0_csc_reg[14]/P0001 ,
		_w4182_,
		_w4183_,
		_w4754_
	);
	LUT4 #(
		.INIT('h0020)
	) name3795 (
		\u0_rf_we_reg/NET0131 ,
		\u0_u0_addr_r_reg[2]/P0001 ,
		\u0_u0_addr_r_reg[4]/P0001 ,
		\wb_data_i[14]_pad ,
		_w4755_
	);
	LUT3 #(
		.INIT('h15)
	) name3796 (
		\u0_rst_r2_reg/NET0131 ,
		_w4182_,
		_w4755_,
		_w4756_
	);
	LUT2 #(
		.INIT('h4)
	) name3797 (
		_w4754_,
		_w4756_,
		_w4757_
	);
	LUT3 #(
		.INIT('h15)
	) name3798 (
		\u0_u0_csc_reg[16]/P0001 ,
		_w4182_,
		_w4183_,
		_w4758_
	);
	LUT4 #(
		.INIT('h0020)
	) name3799 (
		\u0_rf_we_reg/NET0131 ,
		\u0_u0_addr_r_reg[2]/P0001 ,
		\u0_u0_addr_r_reg[4]/P0001 ,
		\wb_data_i[16]_pad ,
		_w4759_
	);
	LUT3 #(
		.INIT('h15)
	) name3800 (
		\u0_rst_r2_reg/NET0131 ,
		_w4182_,
		_w4759_,
		_w4760_
	);
	LUT2 #(
		.INIT('h4)
	) name3801 (
		_w4758_,
		_w4760_,
		_w4761_
	);
	LUT3 #(
		.INIT('h15)
	) name3802 (
		\u0_u0_csc_reg[17]/P0001 ,
		_w4182_,
		_w4183_,
		_w4762_
	);
	LUT4 #(
		.INIT('h0020)
	) name3803 (
		\u0_rf_we_reg/NET0131 ,
		\u0_u0_addr_r_reg[2]/P0001 ,
		\u0_u0_addr_r_reg[4]/P0001 ,
		\wb_data_i[17]_pad ,
		_w4763_
	);
	LUT3 #(
		.INIT('h15)
	) name3804 (
		\u0_rst_r2_reg/NET0131 ,
		_w4182_,
		_w4763_,
		_w4764_
	);
	LUT2 #(
		.INIT('h4)
	) name3805 (
		_w4762_,
		_w4764_,
		_w4765_
	);
	LUT3 #(
		.INIT('h15)
	) name3806 (
		\u0_u0_csc_reg[20]/P0001 ,
		_w4182_,
		_w4183_,
		_w4766_
	);
	LUT4 #(
		.INIT('h0020)
	) name3807 (
		\u0_rf_we_reg/NET0131 ,
		\u0_u0_addr_r_reg[2]/P0001 ,
		\u0_u0_addr_r_reg[4]/P0001 ,
		\wb_data_i[20]_pad ,
		_w4767_
	);
	LUT3 #(
		.INIT('h15)
	) name3808 (
		\u0_rst_r2_reg/NET0131 ,
		_w4182_,
		_w4767_,
		_w4768_
	);
	LUT2 #(
		.INIT('h4)
	) name3809 (
		_w4766_,
		_w4768_,
		_w4769_
	);
	LUT3 #(
		.INIT('h15)
	) name3810 (
		\u0_u0_csc_reg[21]/P0001 ,
		_w4182_,
		_w4183_,
		_w4770_
	);
	LUT4 #(
		.INIT('h0020)
	) name3811 (
		\u0_rf_we_reg/NET0131 ,
		\u0_u0_addr_r_reg[2]/P0001 ,
		\u0_u0_addr_r_reg[4]/P0001 ,
		\wb_data_i[21]_pad ,
		_w4771_
	);
	LUT3 #(
		.INIT('h15)
	) name3812 (
		\u0_rst_r2_reg/NET0131 ,
		_w4182_,
		_w4771_,
		_w4772_
	);
	LUT2 #(
		.INIT('h4)
	) name3813 (
		_w4770_,
		_w4772_,
		_w4773_
	);
	LUT3 #(
		.INIT('h15)
	) name3814 (
		\u0_u0_csc_reg[22]/P0001 ,
		_w4182_,
		_w4183_,
		_w4774_
	);
	LUT4 #(
		.INIT('h0020)
	) name3815 (
		\u0_rf_we_reg/NET0131 ,
		\u0_u0_addr_r_reg[2]/P0001 ,
		\u0_u0_addr_r_reg[4]/P0001 ,
		\wb_data_i[22]_pad ,
		_w4775_
	);
	LUT3 #(
		.INIT('h15)
	) name3816 (
		\u0_rst_r2_reg/NET0131 ,
		_w4182_,
		_w4775_,
		_w4776_
	);
	LUT2 #(
		.INIT('h4)
	) name3817 (
		_w4774_,
		_w4776_,
		_w4777_
	);
	LUT3 #(
		.INIT('h15)
	) name3818 (
		\u0_u0_csc_reg[24]/P0001 ,
		_w4182_,
		_w4183_,
		_w4778_
	);
	LUT4 #(
		.INIT('h0020)
	) name3819 (
		\u0_rf_we_reg/NET0131 ,
		\u0_u0_addr_r_reg[2]/P0001 ,
		\u0_u0_addr_r_reg[4]/P0001 ,
		\wb_data_i[24]_pad ,
		_w4779_
	);
	LUT3 #(
		.INIT('h15)
	) name3820 (
		\u0_rst_r2_reg/NET0131 ,
		_w4182_,
		_w4779_,
		_w4780_
	);
	LUT2 #(
		.INIT('h4)
	) name3821 (
		_w4778_,
		_w4780_,
		_w4781_
	);
	LUT3 #(
		.INIT('h15)
	) name3822 (
		\u0_u0_csc_reg[26]/P0001 ,
		_w4182_,
		_w4183_,
		_w4782_
	);
	LUT4 #(
		.INIT('h0020)
	) name3823 (
		\u0_rf_we_reg/NET0131 ,
		\u0_u0_addr_r_reg[2]/P0001 ,
		\u0_u0_addr_r_reg[4]/P0001 ,
		\wb_data_i[26]_pad ,
		_w4783_
	);
	LUT3 #(
		.INIT('h15)
	) name3824 (
		\u0_rst_r2_reg/NET0131 ,
		_w4182_,
		_w4783_,
		_w4784_
	);
	LUT2 #(
		.INIT('h4)
	) name3825 (
		_w4782_,
		_w4784_,
		_w4785_
	);
	LUT3 #(
		.INIT('h15)
	) name3826 (
		\u0_u0_csc_reg[27]/P0001 ,
		_w4182_,
		_w4183_,
		_w4786_
	);
	LUT4 #(
		.INIT('h0020)
	) name3827 (
		\u0_rf_we_reg/NET0131 ,
		\u0_u0_addr_r_reg[2]/P0001 ,
		\u0_u0_addr_r_reg[4]/P0001 ,
		\wb_data_i[27]_pad ,
		_w4787_
	);
	LUT3 #(
		.INIT('h15)
	) name3828 (
		\u0_rst_r2_reg/NET0131 ,
		_w4182_,
		_w4787_,
		_w4788_
	);
	LUT2 #(
		.INIT('h4)
	) name3829 (
		_w4786_,
		_w4788_,
		_w4789_
	);
	LUT3 #(
		.INIT('h15)
	) name3830 (
		\u0_u0_csc_reg[28]/P0001 ,
		_w4182_,
		_w4183_,
		_w4790_
	);
	LUT4 #(
		.INIT('h0020)
	) name3831 (
		\u0_rf_we_reg/NET0131 ,
		\u0_u0_addr_r_reg[2]/P0001 ,
		\u0_u0_addr_r_reg[4]/P0001 ,
		\wb_data_i[28]_pad ,
		_w4791_
	);
	LUT3 #(
		.INIT('h15)
	) name3832 (
		\u0_rst_r2_reg/NET0131 ,
		_w4182_,
		_w4791_,
		_w4792_
	);
	LUT2 #(
		.INIT('h4)
	) name3833 (
		_w4790_,
		_w4792_,
		_w4793_
	);
	LUT3 #(
		.INIT('h15)
	) name3834 (
		\u0_u1_tms_reg[23]/P0001 ,
		_w4743_,
		_w4744_,
		_w4794_
	);
	LUT4 #(
		.INIT('h0080)
	) name3835 (
		\u0_rf_we_reg/NET0131 ,
		\u0_u0_addr_r_reg[2]/P0001 ,
		\u0_u0_addr_r_reg[4]/P0001 ,
		\wb_data_i[23]_pad ,
		_w4795_
	);
	LUT3 #(
		.INIT('h15)
	) name3836 (
		\u0_rst_r2_reg/NET0131 ,
		_w4743_,
		_w4795_,
		_w4796_
	);
	LUT2 #(
		.INIT('h4)
	) name3837 (
		_w4794_,
		_w4796_,
		_w4797_
	);
	LUT3 #(
		.INIT('h15)
	) name3838 (
		\u0_u0_csc_reg[30]/P0001 ,
		_w4182_,
		_w4183_,
		_w4798_
	);
	LUT4 #(
		.INIT('h0020)
	) name3839 (
		\u0_rf_we_reg/NET0131 ,
		\u0_u0_addr_r_reg[2]/P0001 ,
		\u0_u0_addr_r_reg[4]/P0001 ,
		\wb_data_i[30]_pad ,
		_w4799_
	);
	LUT3 #(
		.INIT('h15)
	) name3840 (
		\u0_rst_r2_reg/NET0131 ,
		_w4182_,
		_w4799_,
		_w4800_
	);
	LUT2 #(
		.INIT('h4)
	) name3841 (
		_w4798_,
		_w4800_,
		_w4801_
	);
	LUT3 #(
		.INIT('h15)
	) name3842 (
		\u0_u0_csc_reg[3]/NET0131 ,
		_w4182_,
		_w4183_,
		_w4802_
	);
	LUT4 #(
		.INIT('h0020)
	) name3843 (
		\u0_rf_we_reg/NET0131 ,
		\u0_u0_addr_r_reg[2]/P0001 ,
		\u0_u0_addr_r_reg[4]/P0001 ,
		\wb_data_i[3]_pad ,
		_w4803_
	);
	LUT3 #(
		.INIT('h15)
	) name3844 (
		\u0_rst_r2_reg/NET0131 ,
		_w4182_,
		_w4803_,
		_w4804_
	);
	LUT2 #(
		.INIT('h4)
	) name3845 (
		_w4802_,
		_w4804_,
		_w4805_
	);
	LUT3 #(
		.INIT('h15)
	) name3846 (
		\u0_u0_csc_reg[25]/P0001 ,
		_w4182_,
		_w4183_,
		_w4806_
	);
	LUT4 #(
		.INIT('h0020)
	) name3847 (
		\u0_rf_we_reg/NET0131 ,
		\u0_u0_addr_r_reg[2]/P0001 ,
		\u0_u0_addr_r_reg[4]/P0001 ,
		\wb_data_i[25]_pad ,
		_w4807_
	);
	LUT3 #(
		.INIT('h15)
	) name3848 (
		\u0_rst_r2_reg/NET0131 ,
		_w4182_,
		_w4807_,
		_w4808_
	);
	LUT2 #(
		.INIT('h4)
	) name3849 (
		_w4806_,
		_w4808_,
		_w4809_
	);
	LUT3 #(
		.INIT('h15)
	) name3850 (
		\u0_u1_tms_reg[17]/P0001 ,
		_w4743_,
		_w4744_,
		_w4810_
	);
	LUT4 #(
		.INIT('h0080)
	) name3851 (
		\u0_rf_we_reg/NET0131 ,
		\u0_u0_addr_r_reg[2]/P0001 ,
		\u0_u0_addr_r_reg[4]/P0001 ,
		\wb_data_i[17]_pad ,
		_w4811_
	);
	LUT3 #(
		.INIT('h15)
	) name3852 (
		\u0_rst_r2_reg/NET0131 ,
		_w4743_,
		_w4811_,
		_w4812_
	);
	LUT2 #(
		.INIT('h4)
	) name3853 (
		_w4810_,
		_w4812_,
		_w4813_
	);
	LUT3 #(
		.INIT('h15)
	) name3854 (
		\u0_u1_tms_reg[16]/P0001 ,
		_w4743_,
		_w4744_,
		_w4814_
	);
	LUT4 #(
		.INIT('h0080)
	) name3855 (
		\u0_rf_we_reg/NET0131 ,
		\u0_u0_addr_r_reg[2]/P0001 ,
		\u0_u0_addr_r_reg[4]/P0001 ,
		\wb_data_i[16]_pad ,
		_w4815_
	);
	LUT3 #(
		.INIT('h15)
	) name3856 (
		\u0_rst_r2_reg/NET0131 ,
		_w4743_,
		_w4815_,
		_w4816_
	);
	LUT2 #(
		.INIT('h4)
	) name3857 (
		_w4814_,
		_w4816_,
		_w4817_
	);
	LUT2 #(
		.INIT('h8)
	) name3858 (
		_w4182_,
		_w4744_,
		_w4818_
	);
	LUT3 #(
		.INIT('h2a)
	) name3859 (
		\u0_u0_tms_reg[0]/P0001 ,
		_w4182_,
		_w4744_,
		_w4819_
	);
	LUT4 #(
		.INIT('h8000)
	) name3860 (
		\u0_rf_we_reg/NET0131 ,
		\u0_u0_addr_r_reg[2]/P0001 ,
		\u0_u0_addr_r_reg[4]/P0001 ,
		\wb_data_i[0]_pad ,
		_w4820_
	);
	LUT3 #(
		.INIT('h15)
	) name3861 (
		\u0_rst_r2_reg/NET0131 ,
		_w4182_,
		_w4820_,
		_w4821_
	);
	LUT2 #(
		.INIT('hb)
	) name3862 (
		_w4819_,
		_w4821_,
		_w4822_
	);
	LUT3 #(
		.INIT('h2a)
	) name3863 (
		\u0_u0_tms_reg[10]/P0001 ,
		_w4182_,
		_w4744_,
		_w4823_
	);
	LUT4 #(
		.INIT('h8000)
	) name3864 (
		\u0_rf_we_reg/NET0131 ,
		\u0_u0_addr_r_reg[2]/P0001 ,
		\u0_u0_addr_r_reg[4]/P0001 ,
		\wb_data_i[10]_pad ,
		_w4824_
	);
	LUT3 #(
		.INIT('h15)
	) name3865 (
		\u0_rst_r2_reg/NET0131 ,
		_w4182_,
		_w4824_,
		_w4825_
	);
	LUT2 #(
		.INIT('hb)
	) name3866 (
		_w4823_,
		_w4825_,
		_w4826_
	);
	LUT3 #(
		.INIT('h2a)
	) name3867 (
		\u0_u0_tms_reg[11]/P0001 ,
		_w4182_,
		_w4744_,
		_w4827_
	);
	LUT4 #(
		.INIT('h8000)
	) name3868 (
		\u0_rf_we_reg/NET0131 ,
		\u0_u0_addr_r_reg[2]/P0001 ,
		\u0_u0_addr_r_reg[4]/P0001 ,
		\wb_data_i[11]_pad ,
		_w4828_
	);
	LUT3 #(
		.INIT('h15)
	) name3869 (
		\u0_rst_r2_reg/NET0131 ,
		_w4182_,
		_w4828_,
		_w4829_
	);
	LUT2 #(
		.INIT('hb)
	) name3870 (
		_w4827_,
		_w4829_,
		_w4830_
	);
	LUT3 #(
		.INIT('h2a)
	) name3871 (
		\u0_u0_tms_reg[12]/P0001 ,
		_w4182_,
		_w4744_,
		_w4831_
	);
	LUT4 #(
		.INIT('h8000)
	) name3872 (
		\u0_rf_we_reg/NET0131 ,
		\u0_u0_addr_r_reg[2]/P0001 ,
		\u0_u0_addr_r_reg[4]/P0001 ,
		\wb_data_i[12]_pad ,
		_w4832_
	);
	LUT3 #(
		.INIT('h15)
	) name3873 (
		\u0_rst_r2_reg/NET0131 ,
		_w4182_,
		_w4832_,
		_w4833_
	);
	LUT2 #(
		.INIT('hb)
	) name3874 (
		_w4831_,
		_w4833_,
		_w4834_
	);
	LUT3 #(
		.INIT('h2a)
	) name3875 (
		\u0_u0_tms_reg[14]/P0001 ,
		_w4182_,
		_w4744_,
		_w4835_
	);
	LUT4 #(
		.INIT('h8000)
	) name3876 (
		\u0_rf_we_reg/NET0131 ,
		\u0_u0_addr_r_reg[2]/P0001 ,
		\u0_u0_addr_r_reg[4]/P0001 ,
		\wb_data_i[14]_pad ,
		_w4836_
	);
	LUT3 #(
		.INIT('h15)
	) name3877 (
		\u0_rst_r2_reg/NET0131 ,
		_w4182_,
		_w4836_,
		_w4837_
	);
	LUT2 #(
		.INIT('hb)
	) name3878 (
		_w4835_,
		_w4837_,
		_w4838_
	);
	LUT3 #(
		.INIT('h2a)
	) name3879 (
		\u0_u0_tms_reg[13]/P0001 ,
		_w4182_,
		_w4744_,
		_w4839_
	);
	LUT4 #(
		.INIT('h8000)
	) name3880 (
		\u0_rf_we_reg/NET0131 ,
		\u0_u0_addr_r_reg[2]/P0001 ,
		\u0_u0_addr_r_reg[4]/P0001 ,
		\wb_data_i[13]_pad ,
		_w4840_
	);
	LUT3 #(
		.INIT('h15)
	) name3881 (
		\u0_rst_r2_reg/NET0131 ,
		_w4182_,
		_w4840_,
		_w4841_
	);
	LUT2 #(
		.INIT('hb)
	) name3882 (
		_w4839_,
		_w4841_,
		_w4842_
	);
	LUT3 #(
		.INIT('h2a)
	) name3883 (
		\u0_u0_tms_reg[15]/P0001 ,
		_w4182_,
		_w4744_,
		_w4843_
	);
	LUT4 #(
		.INIT('h8000)
	) name3884 (
		\u0_rf_we_reg/NET0131 ,
		\u0_u0_addr_r_reg[2]/P0001 ,
		\u0_u0_addr_r_reg[4]/P0001 ,
		\wb_data_i[15]_pad ,
		_w4844_
	);
	LUT3 #(
		.INIT('h15)
	) name3885 (
		\u0_rst_r2_reg/NET0131 ,
		_w4182_,
		_w4844_,
		_w4845_
	);
	LUT2 #(
		.INIT('hb)
	) name3886 (
		_w4843_,
		_w4845_,
		_w4846_
	);
	LUT3 #(
		.INIT('h2a)
	) name3887 (
		\u0_u0_tms_reg[16]/P0001 ,
		_w4182_,
		_w4744_,
		_w4847_
	);
	LUT4 #(
		.INIT('h8000)
	) name3888 (
		\u0_rf_we_reg/NET0131 ,
		\u0_u0_addr_r_reg[2]/P0001 ,
		\u0_u0_addr_r_reg[4]/P0001 ,
		\wb_data_i[16]_pad ,
		_w4848_
	);
	LUT3 #(
		.INIT('h15)
	) name3889 (
		\u0_rst_r2_reg/NET0131 ,
		_w4182_,
		_w4848_,
		_w4849_
	);
	LUT2 #(
		.INIT('hb)
	) name3890 (
		_w4847_,
		_w4849_,
		_w4850_
	);
	LUT3 #(
		.INIT('h2a)
	) name3891 (
		\u0_u0_tms_reg[17]/P0001 ,
		_w4182_,
		_w4744_,
		_w4851_
	);
	LUT4 #(
		.INIT('h8000)
	) name3892 (
		\u0_rf_we_reg/NET0131 ,
		\u0_u0_addr_r_reg[2]/P0001 ,
		\u0_u0_addr_r_reg[4]/P0001 ,
		\wb_data_i[17]_pad ,
		_w4852_
	);
	LUT3 #(
		.INIT('h15)
	) name3893 (
		\u0_rst_r2_reg/NET0131 ,
		_w4182_,
		_w4852_,
		_w4853_
	);
	LUT2 #(
		.INIT('hb)
	) name3894 (
		_w4851_,
		_w4853_,
		_w4854_
	);
	LUT3 #(
		.INIT('h2a)
	) name3895 (
		\u0_u0_tms_reg[18]/P0001 ,
		_w4182_,
		_w4744_,
		_w4855_
	);
	LUT4 #(
		.INIT('h8000)
	) name3896 (
		\u0_rf_we_reg/NET0131 ,
		\u0_u0_addr_r_reg[2]/P0001 ,
		\u0_u0_addr_r_reg[4]/P0001 ,
		\wb_data_i[18]_pad ,
		_w4856_
	);
	LUT3 #(
		.INIT('h15)
	) name3897 (
		\u0_rst_r2_reg/NET0131 ,
		_w4182_,
		_w4856_,
		_w4857_
	);
	LUT2 #(
		.INIT('hb)
	) name3898 (
		_w4855_,
		_w4857_,
		_w4858_
	);
	LUT3 #(
		.INIT('h2a)
	) name3899 (
		\u0_u0_tms_reg[19]/P0001 ,
		_w4182_,
		_w4744_,
		_w4859_
	);
	LUT4 #(
		.INIT('h8000)
	) name3900 (
		\u0_rf_we_reg/NET0131 ,
		\u0_u0_addr_r_reg[2]/P0001 ,
		\u0_u0_addr_r_reg[4]/P0001 ,
		\wb_data_i[19]_pad ,
		_w4860_
	);
	LUT3 #(
		.INIT('h15)
	) name3901 (
		\u0_rst_r2_reg/NET0131 ,
		_w4182_,
		_w4860_,
		_w4861_
	);
	LUT2 #(
		.INIT('hb)
	) name3902 (
		_w4859_,
		_w4861_,
		_w4862_
	);
	LUT3 #(
		.INIT('h2a)
	) name3903 (
		\u0_u0_tms_reg[1]/P0001 ,
		_w4182_,
		_w4744_,
		_w4863_
	);
	LUT4 #(
		.INIT('h8000)
	) name3904 (
		\u0_rf_we_reg/NET0131 ,
		\u0_u0_addr_r_reg[2]/P0001 ,
		\u0_u0_addr_r_reg[4]/P0001 ,
		\wb_data_i[1]_pad ,
		_w4864_
	);
	LUT3 #(
		.INIT('h15)
	) name3905 (
		\u0_rst_r2_reg/NET0131 ,
		_w4182_,
		_w4864_,
		_w4865_
	);
	LUT2 #(
		.INIT('hb)
	) name3906 (
		_w4863_,
		_w4865_,
		_w4866_
	);
	LUT3 #(
		.INIT('h2a)
	) name3907 (
		\u0_u0_tms_reg[21]/P0001 ,
		_w4182_,
		_w4744_,
		_w4867_
	);
	LUT4 #(
		.INIT('h8000)
	) name3908 (
		\u0_rf_we_reg/NET0131 ,
		\u0_u0_addr_r_reg[2]/P0001 ,
		\u0_u0_addr_r_reg[4]/P0001 ,
		\wb_data_i[21]_pad ,
		_w4868_
	);
	LUT3 #(
		.INIT('h15)
	) name3909 (
		\u0_rst_r2_reg/NET0131 ,
		_w4182_,
		_w4868_,
		_w4869_
	);
	LUT2 #(
		.INIT('hb)
	) name3910 (
		_w4867_,
		_w4869_,
		_w4870_
	);
	LUT3 #(
		.INIT('h2a)
	) name3911 (
		\u0_u0_tms_reg[22]/P0001 ,
		_w4182_,
		_w4744_,
		_w4871_
	);
	LUT4 #(
		.INIT('h8000)
	) name3912 (
		\u0_rf_we_reg/NET0131 ,
		\u0_u0_addr_r_reg[2]/P0001 ,
		\u0_u0_addr_r_reg[4]/P0001 ,
		\wb_data_i[22]_pad ,
		_w4872_
	);
	LUT3 #(
		.INIT('h15)
	) name3913 (
		\u0_rst_r2_reg/NET0131 ,
		_w4182_,
		_w4872_,
		_w4873_
	);
	LUT2 #(
		.INIT('hb)
	) name3914 (
		_w4871_,
		_w4873_,
		_w4874_
	);
	LUT3 #(
		.INIT('h2a)
	) name3915 (
		\u0_u0_tms_reg[23]/P0001 ,
		_w4182_,
		_w4744_,
		_w4875_
	);
	LUT4 #(
		.INIT('h8000)
	) name3916 (
		\u0_rf_we_reg/NET0131 ,
		\u0_u0_addr_r_reg[2]/P0001 ,
		\u0_u0_addr_r_reg[4]/P0001 ,
		\wb_data_i[23]_pad ,
		_w4876_
	);
	LUT3 #(
		.INIT('h15)
	) name3917 (
		\u0_rst_r2_reg/NET0131 ,
		_w4182_,
		_w4876_,
		_w4877_
	);
	LUT2 #(
		.INIT('hb)
	) name3918 (
		_w4875_,
		_w4877_,
		_w4878_
	);
	LUT3 #(
		.INIT('h2a)
	) name3919 (
		\u0_u0_tms_reg[24]/P0001 ,
		_w4182_,
		_w4744_,
		_w4879_
	);
	LUT4 #(
		.INIT('h8000)
	) name3920 (
		\u0_rf_we_reg/NET0131 ,
		\u0_u0_addr_r_reg[2]/P0001 ,
		\u0_u0_addr_r_reg[4]/P0001 ,
		\wb_data_i[24]_pad ,
		_w4880_
	);
	LUT3 #(
		.INIT('h15)
	) name3921 (
		\u0_rst_r2_reg/NET0131 ,
		_w4182_,
		_w4880_,
		_w4881_
	);
	LUT2 #(
		.INIT('hb)
	) name3922 (
		_w4879_,
		_w4881_,
		_w4882_
	);
	LUT3 #(
		.INIT('h2a)
	) name3923 (
		\u0_u0_tms_reg[25]/P0001 ,
		_w4182_,
		_w4744_,
		_w4883_
	);
	LUT4 #(
		.INIT('h8000)
	) name3924 (
		\u0_rf_we_reg/NET0131 ,
		\u0_u0_addr_r_reg[2]/P0001 ,
		\u0_u0_addr_r_reg[4]/P0001 ,
		\wb_data_i[25]_pad ,
		_w4884_
	);
	LUT3 #(
		.INIT('h15)
	) name3925 (
		\u0_rst_r2_reg/NET0131 ,
		_w4182_,
		_w4884_,
		_w4885_
	);
	LUT2 #(
		.INIT('hb)
	) name3926 (
		_w4883_,
		_w4885_,
		_w4886_
	);
	LUT3 #(
		.INIT('h2a)
	) name3927 (
		\u0_u0_tms_reg[26]/P0001 ,
		_w4182_,
		_w4744_,
		_w4887_
	);
	LUT4 #(
		.INIT('h8000)
	) name3928 (
		\u0_rf_we_reg/NET0131 ,
		\u0_u0_addr_r_reg[2]/P0001 ,
		\u0_u0_addr_r_reg[4]/P0001 ,
		\wb_data_i[26]_pad ,
		_w4888_
	);
	LUT3 #(
		.INIT('h15)
	) name3929 (
		\u0_rst_r2_reg/NET0131 ,
		_w4182_,
		_w4888_,
		_w4889_
	);
	LUT2 #(
		.INIT('hb)
	) name3930 (
		_w4887_,
		_w4889_,
		_w4890_
	);
	LUT3 #(
		.INIT('h2a)
	) name3931 (
		\u0_u0_tms_reg[27]/P0001 ,
		_w4182_,
		_w4744_,
		_w4891_
	);
	LUT4 #(
		.INIT('h8000)
	) name3932 (
		\u0_rf_we_reg/NET0131 ,
		\u0_u0_addr_r_reg[2]/P0001 ,
		\u0_u0_addr_r_reg[4]/P0001 ,
		\wb_data_i[27]_pad ,
		_w4892_
	);
	LUT3 #(
		.INIT('h15)
	) name3933 (
		\u0_rst_r2_reg/NET0131 ,
		_w4182_,
		_w4892_,
		_w4893_
	);
	LUT2 #(
		.INIT('hb)
	) name3934 (
		_w4891_,
		_w4893_,
		_w4894_
	);
	LUT3 #(
		.INIT('h15)
	) name3935 (
		\u0_u1_tms_reg[22]/P0001 ,
		_w4743_,
		_w4744_,
		_w4895_
	);
	LUT4 #(
		.INIT('h0080)
	) name3936 (
		\u0_rf_we_reg/NET0131 ,
		\u0_u0_addr_r_reg[2]/P0001 ,
		\u0_u0_addr_r_reg[4]/P0001 ,
		\wb_data_i[22]_pad ,
		_w4896_
	);
	LUT3 #(
		.INIT('h15)
	) name3937 (
		\u0_rst_r2_reg/NET0131 ,
		_w4743_,
		_w4896_,
		_w4897_
	);
	LUT2 #(
		.INIT('h4)
	) name3938 (
		_w4895_,
		_w4897_,
		_w4898_
	);
	LUT3 #(
		.INIT('h2a)
	) name3939 (
		\u0_u0_tms_reg[28]/P0001 ,
		_w4182_,
		_w4744_,
		_w4899_
	);
	LUT4 #(
		.INIT('h8000)
	) name3940 (
		\u0_rf_we_reg/NET0131 ,
		\u0_u0_addr_r_reg[2]/P0001 ,
		\u0_u0_addr_r_reg[4]/P0001 ,
		\wb_data_i[28]_pad ,
		_w4900_
	);
	LUT3 #(
		.INIT('h15)
	) name3941 (
		\u0_rst_r2_reg/NET0131 ,
		_w4182_,
		_w4900_,
		_w4901_
	);
	LUT2 #(
		.INIT('hb)
	) name3942 (
		_w4899_,
		_w4901_,
		_w4902_
	);
	LUT3 #(
		.INIT('h2a)
	) name3943 (
		\u0_u0_tms_reg[29]/P0001 ,
		_w4182_,
		_w4744_,
		_w4903_
	);
	LUT4 #(
		.INIT('h8000)
	) name3944 (
		\u0_rf_we_reg/NET0131 ,
		\u0_u0_addr_r_reg[2]/P0001 ,
		\u0_u0_addr_r_reg[4]/P0001 ,
		\wb_data_i[29]_pad ,
		_w4904_
	);
	LUT3 #(
		.INIT('h15)
	) name3945 (
		\u0_rst_r2_reg/NET0131 ,
		_w4182_,
		_w4904_,
		_w4905_
	);
	LUT2 #(
		.INIT('hb)
	) name3946 (
		_w4903_,
		_w4905_,
		_w4906_
	);
	LUT3 #(
		.INIT('h2a)
	) name3947 (
		\u0_u0_tms_reg[2]/P0001 ,
		_w4182_,
		_w4744_,
		_w4907_
	);
	LUT4 #(
		.INIT('h8000)
	) name3948 (
		\u0_rf_we_reg/NET0131 ,
		\u0_u0_addr_r_reg[2]/P0001 ,
		\u0_u0_addr_r_reg[4]/P0001 ,
		\wb_data_i[2]_pad ,
		_w4908_
	);
	LUT3 #(
		.INIT('h15)
	) name3949 (
		\u0_rst_r2_reg/NET0131 ,
		_w4182_,
		_w4908_,
		_w4909_
	);
	LUT2 #(
		.INIT('hb)
	) name3950 (
		_w4907_,
		_w4909_,
		_w4910_
	);
	LUT3 #(
		.INIT('h15)
	) name3951 (
		\u0_u0_csc_reg[15]/P0001 ,
		_w4182_,
		_w4183_,
		_w4911_
	);
	LUT4 #(
		.INIT('h0020)
	) name3952 (
		\u0_rf_we_reg/NET0131 ,
		\u0_u0_addr_r_reg[2]/P0001 ,
		\u0_u0_addr_r_reg[4]/P0001 ,
		\wb_data_i[15]_pad ,
		_w4912_
	);
	LUT3 #(
		.INIT('h15)
	) name3953 (
		\u0_rst_r2_reg/NET0131 ,
		_w4182_,
		_w4912_,
		_w4913_
	);
	LUT2 #(
		.INIT('h4)
	) name3954 (
		_w4911_,
		_w4913_,
		_w4914_
	);
	LUT3 #(
		.INIT('h2a)
	) name3955 (
		\u0_u0_tms_reg[30]/P0001 ,
		_w4182_,
		_w4744_,
		_w4915_
	);
	LUT4 #(
		.INIT('h8000)
	) name3956 (
		\u0_rf_we_reg/NET0131 ,
		\u0_u0_addr_r_reg[2]/P0001 ,
		\u0_u0_addr_r_reg[4]/P0001 ,
		\wb_data_i[30]_pad ,
		_w4916_
	);
	LUT3 #(
		.INIT('h15)
	) name3957 (
		\u0_rst_r2_reg/NET0131 ,
		_w4182_,
		_w4916_,
		_w4917_
	);
	LUT2 #(
		.INIT('hb)
	) name3958 (
		_w4915_,
		_w4917_,
		_w4918_
	);
	LUT3 #(
		.INIT('h2a)
	) name3959 (
		\u0_u0_tms_reg[3]/P0001 ,
		_w4182_,
		_w4744_,
		_w4919_
	);
	LUT4 #(
		.INIT('h8000)
	) name3960 (
		\u0_rf_we_reg/NET0131 ,
		\u0_u0_addr_r_reg[2]/P0001 ,
		\u0_u0_addr_r_reg[4]/P0001 ,
		\wb_data_i[3]_pad ,
		_w4920_
	);
	LUT3 #(
		.INIT('h15)
	) name3961 (
		\u0_rst_r2_reg/NET0131 ,
		_w4182_,
		_w4920_,
		_w4921_
	);
	LUT2 #(
		.INIT('hb)
	) name3962 (
		_w4919_,
		_w4921_,
		_w4922_
	);
	LUT3 #(
		.INIT('h2a)
	) name3963 (
		\u0_u0_tms_reg[4]/P0001 ,
		_w4182_,
		_w4744_,
		_w4923_
	);
	LUT4 #(
		.INIT('h8000)
	) name3964 (
		\u0_rf_we_reg/NET0131 ,
		\u0_u0_addr_r_reg[2]/P0001 ,
		\u0_u0_addr_r_reg[4]/P0001 ,
		\wb_data_i[4]_pad ,
		_w4924_
	);
	LUT3 #(
		.INIT('h15)
	) name3965 (
		\u0_rst_r2_reg/NET0131 ,
		_w4182_,
		_w4924_,
		_w4925_
	);
	LUT2 #(
		.INIT('hb)
	) name3966 (
		_w4923_,
		_w4925_,
		_w4926_
	);
	LUT3 #(
		.INIT('h2a)
	) name3967 (
		\u0_u0_tms_reg[5]/P0001 ,
		_w4182_,
		_w4744_,
		_w4927_
	);
	LUT4 #(
		.INIT('h8000)
	) name3968 (
		\u0_rf_we_reg/NET0131 ,
		\u0_u0_addr_r_reg[2]/P0001 ,
		\u0_u0_addr_r_reg[4]/P0001 ,
		\wb_data_i[5]_pad ,
		_w4928_
	);
	LUT3 #(
		.INIT('h15)
	) name3969 (
		\u0_rst_r2_reg/NET0131 ,
		_w4182_,
		_w4928_,
		_w4929_
	);
	LUT2 #(
		.INIT('hb)
	) name3970 (
		_w4927_,
		_w4929_,
		_w4930_
	);
	LUT3 #(
		.INIT('h2a)
	) name3971 (
		\u0_u0_tms_reg[6]/P0001 ,
		_w4182_,
		_w4744_,
		_w4931_
	);
	LUT4 #(
		.INIT('h8000)
	) name3972 (
		\u0_rf_we_reg/NET0131 ,
		\u0_u0_addr_r_reg[2]/P0001 ,
		\u0_u0_addr_r_reg[4]/P0001 ,
		\wb_data_i[6]_pad ,
		_w4932_
	);
	LUT3 #(
		.INIT('h15)
	) name3973 (
		\u0_rst_r2_reg/NET0131 ,
		_w4182_,
		_w4932_,
		_w4933_
	);
	LUT2 #(
		.INIT('hb)
	) name3974 (
		_w4931_,
		_w4933_,
		_w4934_
	);
	LUT3 #(
		.INIT('h2a)
	) name3975 (
		\u0_u0_tms_reg[7]/P0001 ,
		_w4182_,
		_w4744_,
		_w4935_
	);
	LUT4 #(
		.INIT('h8000)
	) name3976 (
		\u0_rf_we_reg/NET0131 ,
		\u0_u0_addr_r_reg[2]/P0001 ,
		\u0_u0_addr_r_reg[4]/P0001 ,
		\wb_data_i[7]_pad ,
		_w4936_
	);
	LUT3 #(
		.INIT('h15)
	) name3977 (
		\u0_rst_r2_reg/NET0131 ,
		_w4182_,
		_w4936_,
		_w4937_
	);
	LUT2 #(
		.INIT('hb)
	) name3978 (
		_w4935_,
		_w4937_,
		_w4938_
	);
	LUT3 #(
		.INIT('h2a)
	) name3979 (
		\u0_u0_tms_reg[8]/P0001 ,
		_w4182_,
		_w4744_,
		_w4939_
	);
	LUT4 #(
		.INIT('h8000)
	) name3980 (
		\u0_rf_we_reg/NET0131 ,
		\u0_u0_addr_r_reg[2]/P0001 ,
		\u0_u0_addr_r_reg[4]/P0001 ,
		\wb_data_i[8]_pad ,
		_w4940_
	);
	LUT3 #(
		.INIT('h15)
	) name3981 (
		\u0_rst_r2_reg/NET0131 ,
		_w4182_,
		_w4940_,
		_w4941_
	);
	LUT2 #(
		.INIT('hb)
	) name3982 (
		_w4939_,
		_w4941_,
		_w4942_
	);
	LUT3 #(
		.INIT('h2a)
	) name3983 (
		\u0_u0_tms_reg[9]/P0001 ,
		_w4182_,
		_w4744_,
		_w4943_
	);
	LUT4 #(
		.INIT('h8000)
	) name3984 (
		\u0_rf_we_reg/NET0131 ,
		\u0_u0_addr_r_reg[2]/P0001 ,
		\u0_u0_addr_r_reg[4]/P0001 ,
		\wb_data_i[9]_pad ,
		_w4944_
	);
	LUT3 #(
		.INIT('h15)
	) name3985 (
		\u0_rst_r2_reg/NET0131 ,
		_w4182_,
		_w4944_,
		_w4945_
	);
	LUT2 #(
		.INIT('hb)
	) name3986 (
		_w4943_,
		_w4945_,
		_w4946_
	);
	LUT2 #(
		.INIT('h8)
	) name3987 (
		_w4183_,
		_w4743_,
		_w4947_
	);
	LUT3 #(
		.INIT('h15)
	) name3988 (
		\u0_u1_csc_reg[0]/NET0131 ,
		_w4183_,
		_w4743_,
		_w4948_
	);
	LUT3 #(
		.INIT('h15)
	) name3989 (
		\u0_rst_r2_reg/NET0131 ,
		_w4186_,
		_w4743_,
		_w4949_
	);
	LUT2 #(
		.INIT('h4)
	) name3990 (
		_w4948_,
		_w4949_,
		_w4950_
	);
	LUT3 #(
		.INIT('h15)
	) name3991 (
		\u0_u1_csc_reg[10]/P0001 ,
		_w4183_,
		_w4743_,
		_w4951_
	);
	LUT4 #(
		.INIT('h0020)
	) name3992 (
		\u0_rf_we_reg/NET0131 ,
		\u0_u0_addr_r_reg[2]/P0001 ,
		\u0_u0_addr_r_reg[4]/P0001 ,
		\wb_data_i[10]_pad ,
		_w4952_
	);
	LUT3 #(
		.INIT('h15)
	) name3993 (
		\u0_rst_r2_reg/NET0131 ,
		_w4743_,
		_w4952_,
		_w4953_
	);
	LUT2 #(
		.INIT('h4)
	) name3994 (
		_w4951_,
		_w4953_,
		_w4954_
	);
	LUT3 #(
		.INIT('h15)
	) name3995 (
		\u0_u1_csc_reg[11]/P0001 ,
		_w4183_,
		_w4743_,
		_w4955_
	);
	LUT3 #(
		.INIT('h15)
	) name3996 (
		\u0_rst_r2_reg/NET0131 ,
		_w4736_,
		_w4743_,
		_w4956_
	);
	LUT2 #(
		.INIT('h4)
	) name3997 (
		_w4955_,
		_w4956_,
		_w4957_
	);
	LUT3 #(
		.INIT('h15)
	) name3998 (
		\u0_u1_csc_reg[12]/P0001 ,
		_w4183_,
		_w4743_,
		_w4958_
	);
	LUT3 #(
		.INIT('h15)
	) name3999 (
		\u0_rst_r2_reg/NET0131 ,
		_w4740_,
		_w4743_,
		_w4959_
	);
	LUT2 #(
		.INIT('h4)
	) name4000 (
		_w4958_,
		_w4959_,
		_w4960_
	);
	LUT3 #(
		.INIT('h15)
	) name4001 (
		\u0_u1_csc_reg[13]/P0001 ,
		_w4183_,
		_w4743_,
		_w4961_
	);
	LUT3 #(
		.INIT('h15)
	) name4002 (
		\u0_rst_r2_reg/NET0131 ,
		_w4743_,
		_w4751_,
		_w4962_
	);
	LUT2 #(
		.INIT('h4)
	) name4003 (
		_w4961_,
		_w4962_,
		_w4963_
	);
	LUT3 #(
		.INIT('h15)
	) name4004 (
		\u0_u1_csc_reg[14]/P0001 ,
		_w4183_,
		_w4743_,
		_w4964_
	);
	LUT3 #(
		.INIT('h15)
	) name4005 (
		\u0_rst_r2_reg/NET0131 ,
		_w4743_,
		_w4755_,
		_w4965_
	);
	LUT2 #(
		.INIT('h4)
	) name4006 (
		_w4964_,
		_w4965_,
		_w4966_
	);
	LUT3 #(
		.INIT('h15)
	) name4007 (
		\u0_u1_csc_reg[15]/P0001 ,
		_w4183_,
		_w4743_,
		_w4967_
	);
	LUT3 #(
		.INIT('h15)
	) name4008 (
		\u0_rst_r2_reg/NET0131 ,
		_w4743_,
		_w4912_,
		_w4968_
	);
	LUT2 #(
		.INIT('h4)
	) name4009 (
		_w4967_,
		_w4968_,
		_w4969_
	);
	LUT3 #(
		.INIT('h15)
	) name4010 (
		\u0_u1_csc_reg[17]/P0001 ,
		_w4183_,
		_w4743_,
		_w4970_
	);
	LUT3 #(
		.INIT('h15)
	) name4011 (
		\u0_rst_r2_reg/NET0131 ,
		_w4743_,
		_w4763_,
		_w4971_
	);
	LUT2 #(
		.INIT('h4)
	) name4012 (
		_w4970_,
		_w4971_,
		_w4972_
	);
	LUT3 #(
		.INIT('h15)
	) name4013 (
		\u0_u1_csc_reg[18]/P0001 ,
		_w4183_,
		_w4743_,
		_w4973_
	);
	LUT4 #(
		.INIT('h0020)
	) name4014 (
		\u0_rf_we_reg/NET0131 ,
		\u0_u0_addr_r_reg[2]/P0001 ,
		\u0_u0_addr_r_reg[4]/P0001 ,
		\wb_data_i[18]_pad ,
		_w4974_
	);
	LUT3 #(
		.INIT('h15)
	) name4015 (
		\u0_rst_r2_reg/NET0131 ,
		_w4743_,
		_w4974_,
		_w4975_
	);
	LUT2 #(
		.INIT('h4)
	) name4016 (
		_w4973_,
		_w4975_,
		_w4976_
	);
	LUT3 #(
		.INIT('h15)
	) name4017 (
		\u0_u1_csc_reg[19]/P0001 ,
		_w4183_,
		_w4743_,
		_w4977_
	);
	LUT4 #(
		.INIT('h0020)
	) name4018 (
		\u0_rf_we_reg/NET0131 ,
		\u0_u0_addr_r_reg[2]/P0001 ,
		\u0_u0_addr_r_reg[4]/P0001 ,
		\wb_data_i[19]_pad ,
		_w4978_
	);
	LUT3 #(
		.INIT('h15)
	) name4019 (
		\u0_rst_r2_reg/NET0131 ,
		_w4743_,
		_w4978_,
		_w4979_
	);
	LUT2 #(
		.INIT('h4)
	) name4020 (
		_w4977_,
		_w4979_,
		_w4980_
	);
	LUT3 #(
		.INIT('h15)
	) name4021 (
		\u0_u1_csc_reg[1]/NET0131 ,
		_w4183_,
		_w4743_,
		_w4981_
	);
	LUT3 #(
		.INIT('h15)
	) name4022 (
		\u0_rst_r2_reg/NET0131 ,
		_w4633_,
		_w4743_,
		_w4982_
	);
	LUT2 #(
		.INIT('h4)
	) name4023 (
		_w4981_,
		_w4982_,
		_w4983_
	);
	LUT3 #(
		.INIT('h15)
	) name4024 (
		\u0_u1_csc_reg[20]/P0001 ,
		_w4183_,
		_w4743_,
		_w4984_
	);
	LUT3 #(
		.INIT('h15)
	) name4025 (
		\u0_rst_r2_reg/NET0131 ,
		_w4743_,
		_w4767_,
		_w4985_
	);
	LUT2 #(
		.INIT('h4)
	) name4026 (
		_w4984_,
		_w4985_,
		_w4986_
	);
	LUT3 #(
		.INIT('h15)
	) name4027 (
		\u0_u0_csc_reg[29]/P0001 ,
		_w4182_,
		_w4183_,
		_w4987_
	);
	LUT4 #(
		.INIT('h0020)
	) name4028 (
		\u0_rf_we_reg/NET0131 ,
		\u0_u0_addr_r_reg[2]/P0001 ,
		\u0_u0_addr_r_reg[4]/P0001 ,
		\wb_data_i[29]_pad ,
		_w4988_
	);
	LUT3 #(
		.INIT('h15)
	) name4029 (
		\u0_rst_r2_reg/NET0131 ,
		_w4182_,
		_w4988_,
		_w4989_
	);
	LUT2 #(
		.INIT('h4)
	) name4030 (
		_w4987_,
		_w4989_,
		_w4990_
	);
	LUT3 #(
		.INIT('h15)
	) name4031 (
		\u0_u1_csc_reg[22]/P0001 ,
		_w4183_,
		_w4743_,
		_w4991_
	);
	LUT3 #(
		.INIT('h15)
	) name4032 (
		\u0_rst_r2_reg/NET0131 ,
		_w4743_,
		_w4775_,
		_w4992_
	);
	LUT2 #(
		.INIT('h4)
	) name4033 (
		_w4991_,
		_w4992_,
		_w4993_
	);
	LUT3 #(
		.INIT('h15)
	) name4034 (
		\u0_u1_csc_reg[23]/P0001 ,
		_w4183_,
		_w4743_,
		_w4994_
	);
	LUT4 #(
		.INIT('h0020)
	) name4035 (
		\u0_rf_we_reg/NET0131 ,
		\u0_u0_addr_r_reg[2]/P0001 ,
		\u0_u0_addr_r_reg[4]/P0001 ,
		\wb_data_i[23]_pad ,
		_w4995_
	);
	LUT3 #(
		.INIT('h15)
	) name4036 (
		\u0_rst_r2_reg/NET0131 ,
		_w4743_,
		_w4995_,
		_w4996_
	);
	LUT2 #(
		.INIT('h4)
	) name4037 (
		_w4994_,
		_w4996_,
		_w4997_
	);
	LUT3 #(
		.INIT('h15)
	) name4038 (
		\u0_u1_csc_reg[21]/P0001 ,
		_w4183_,
		_w4743_,
		_w4998_
	);
	LUT3 #(
		.INIT('h15)
	) name4039 (
		\u0_rst_r2_reg/NET0131 ,
		_w4743_,
		_w4771_,
		_w4999_
	);
	LUT2 #(
		.INIT('h4)
	) name4040 (
		_w4998_,
		_w4999_,
		_w5000_
	);
	LUT3 #(
		.INIT('h15)
	) name4041 (
		\u0_u1_csc_reg[24]/P0001 ,
		_w4183_,
		_w4743_,
		_w5001_
	);
	LUT3 #(
		.INIT('h15)
	) name4042 (
		\u0_rst_r2_reg/NET0131 ,
		_w4743_,
		_w4779_,
		_w5002_
	);
	LUT2 #(
		.INIT('h4)
	) name4043 (
		_w5001_,
		_w5002_,
		_w5003_
	);
	LUT3 #(
		.INIT('h15)
	) name4044 (
		\u0_u1_csc_reg[25]/P0001 ,
		_w4183_,
		_w4743_,
		_w5004_
	);
	LUT3 #(
		.INIT('h15)
	) name4045 (
		\u0_rst_r2_reg/NET0131 ,
		_w4743_,
		_w4807_,
		_w5005_
	);
	LUT2 #(
		.INIT('h4)
	) name4046 (
		_w5004_,
		_w5005_,
		_w5006_
	);
	LUT3 #(
		.INIT('h15)
	) name4047 (
		\u0_u1_csc_reg[26]/P0001 ,
		_w4183_,
		_w4743_,
		_w5007_
	);
	LUT3 #(
		.INIT('h15)
	) name4048 (
		\u0_rst_r2_reg/NET0131 ,
		_w4743_,
		_w4783_,
		_w5008_
	);
	LUT2 #(
		.INIT('h4)
	) name4049 (
		_w5007_,
		_w5008_,
		_w5009_
	);
	LUT3 #(
		.INIT('h15)
	) name4050 (
		\u0_u1_csc_reg[27]/P0001 ,
		_w4183_,
		_w4743_,
		_w5010_
	);
	LUT3 #(
		.INIT('h15)
	) name4051 (
		\u0_rst_r2_reg/NET0131 ,
		_w4743_,
		_w4787_,
		_w5011_
	);
	LUT2 #(
		.INIT('h4)
	) name4052 (
		_w5010_,
		_w5011_,
		_w5012_
	);
	LUT3 #(
		.INIT('h15)
	) name4053 (
		\u0_u1_csc_reg[28]/P0001 ,
		_w4183_,
		_w4743_,
		_w5013_
	);
	LUT3 #(
		.INIT('h15)
	) name4054 (
		\u0_rst_r2_reg/NET0131 ,
		_w4743_,
		_w4791_,
		_w5014_
	);
	LUT2 #(
		.INIT('h4)
	) name4055 (
		_w5013_,
		_w5014_,
		_w5015_
	);
	LUT3 #(
		.INIT('h15)
	) name4056 (
		\u0_u0_csc_reg[7]/P0001 ,
		_w4182_,
		_w4183_,
		_w5016_
	);
	LUT4 #(
		.INIT('h0020)
	) name4057 (
		\u0_rf_we_reg/NET0131 ,
		\u0_u0_addr_r_reg[2]/P0001 ,
		\u0_u0_addr_r_reg[4]/P0001 ,
		\wb_data_i[7]_pad ,
		_w5017_
	);
	LUT3 #(
		.INIT('h15)
	) name4058 (
		\u0_rst_r2_reg/NET0131 ,
		_w4182_,
		_w5017_,
		_w5018_
	);
	LUT2 #(
		.INIT('h4)
	) name4059 (
		_w5016_,
		_w5018_,
		_w5019_
	);
	LUT3 #(
		.INIT('h15)
	) name4060 (
		\u0_u1_csc_reg[29]/P0001 ,
		_w4183_,
		_w4743_,
		_w5020_
	);
	LUT3 #(
		.INIT('h15)
	) name4061 (
		\u0_rst_r2_reg/NET0131 ,
		_w4743_,
		_w4988_,
		_w5021_
	);
	LUT2 #(
		.INIT('h4)
	) name4062 (
		_w5020_,
		_w5021_,
		_w5022_
	);
	LUT3 #(
		.INIT('h15)
	) name4063 (
		\u0_u1_csc_reg[2]/NET0131 ,
		_w4183_,
		_w4743_,
		_w5023_
	);
	LUT3 #(
		.INIT('h15)
	) name4064 (
		\u0_rst_r2_reg/NET0131 ,
		_w4637_,
		_w4743_,
		_w5024_
	);
	LUT2 #(
		.INIT('h4)
	) name4065 (
		_w5023_,
		_w5024_,
		_w5025_
	);
	LUT3 #(
		.INIT('h15)
	) name4066 (
		\u0_u1_csc_reg[30]/P0001 ,
		_w4183_,
		_w4743_,
		_w5026_
	);
	LUT3 #(
		.INIT('h15)
	) name4067 (
		\u0_rst_r2_reg/NET0131 ,
		_w4743_,
		_w4799_,
		_w5027_
	);
	LUT2 #(
		.INIT('h4)
	) name4068 (
		_w5026_,
		_w5027_,
		_w5028_
	);
	LUT3 #(
		.INIT('h15)
	) name4069 (
		\u0_u1_csc_reg[31]/P0001 ,
		_w4183_,
		_w4743_,
		_w5029_
	);
	LUT4 #(
		.INIT('h0020)
	) name4070 (
		\u0_rf_we_reg/NET0131 ,
		\u0_u0_addr_r_reg[2]/P0001 ,
		\u0_u0_addr_r_reg[4]/P0001 ,
		\wb_data_i[31]_pad ,
		_w5030_
	);
	LUT3 #(
		.INIT('h15)
	) name4071 (
		\u0_rst_r2_reg/NET0131 ,
		_w4743_,
		_w5030_,
		_w5031_
	);
	LUT2 #(
		.INIT('h4)
	) name4072 (
		_w5029_,
		_w5031_,
		_w5032_
	);
	LUT3 #(
		.INIT('h15)
	) name4073 (
		\u0_u1_csc_reg[4]/P0001 ,
		_w4183_,
		_w4743_,
		_w5033_
	);
	LUT4 #(
		.INIT('h0020)
	) name4074 (
		\u0_rf_we_reg/NET0131 ,
		\u0_u0_addr_r_reg[2]/P0001 ,
		\u0_u0_addr_r_reg[4]/P0001 ,
		\wb_data_i[4]_pad ,
		_w5034_
	);
	LUT3 #(
		.INIT('h15)
	) name4075 (
		\u0_rst_r2_reg/NET0131 ,
		_w4743_,
		_w5034_,
		_w5035_
	);
	LUT2 #(
		.INIT('h4)
	) name4076 (
		_w5033_,
		_w5035_,
		_w5036_
	);
	LUT3 #(
		.INIT('h15)
	) name4077 (
		\u0_u1_csc_reg[3]/NET0131 ,
		_w4183_,
		_w4743_,
		_w5037_
	);
	LUT3 #(
		.INIT('h15)
	) name4078 (
		\u0_rst_r2_reg/NET0131 ,
		_w4743_,
		_w4803_,
		_w5038_
	);
	LUT2 #(
		.INIT('h4)
	) name4079 (
		_w5037_,
		_w5038_,
		_w5039_
	);
	LUT3 #(
		.INIT('h15)
	) name4080 (
		\u0_u1_csc_reg[5]/P0001 ,
		_w4183_,
		_w4743_,
		_w5040_
	);
	LUT4 #(
		.INIT('h0020)
	) name4081 (
		\u0_rf_we_reg/NET0131 ,
		\u0_u0_addr_r_reg[2]/P0001 ,
		\u0_u0_addr_r_reg[4]/P0001 ,
		\wb_data_i[5]_pad ,
		_w5041_
	);
	LUT3 #(
		.INIT('h15)
	) name4082 (
		\u0_rst_r2_reg/NET0131 ,
		_w4743_,
		_w5041_,
		_w5042_
	);
	LUT2 #(
		.INIT('h4)
	) name4083 (
		_w5040_,
		_w5042_,
		_w5043_
	);
	LUT3 #(
		.INIT('h15)
	) name4084 (
		\u0_u1_csc_reg[6]/P0001 ,
		_w4183_,
		_w4743_,
		_w5044_
	);
	LUT4 #(
		.INIT('h0020)
	) name4085 (
		\u0_rf_we_reg/NET0131 ,
		\u0_u0_addr_r_reg[2]/P0001 ,
		\u0_u0_addr_r_reg[4]/P0001 ,
		\wb_data_i[6]_pad ,
		_w5045_
	);
	LUT3 #(
		.INIT('h15)
	) name4086 (
		\u0_rst_r2_reg/NET0131 ,
		_w4743_,
		_w5045_,
		_w5046_
	);
	LUT2 #(
		.INIT('h4)
	) name4087 (
		_w5044_,
		_w5046_,
		_w5047_
	);
	LUT3 #(
		.INIT('h15)
	) name4088 (
		\u0_u0_csc_reg[8]/P0001 ,
		_w4182_,
		_w4183_,
		_w5048_
	);
	LUT4 #(
		.INIT('h0020)
	) name4089 (
		\u0_rf_we_reg/NET0131 ,
		\u0_u0_addr_r_reg[2]/P0001 ,
		\u0_u0_addr_r_reg[4]/P0001 ,
		\wb_data_i[8]_pad ,
		_w5049_
	);
	LUT3 #(
		.INIT('h15)
	) name4090 (
		\u0_rst_r2_reg/NET0131 ,
		_w4182_,
		_w5049_,
		_w5050_
	);
	LUT2 #(
		.INIT('h4)
	) name4091 (
		_w5048_,
		_w5050_,
		_w5051_
	);
	LUT3 #(
		.INIT('h15)
	) name4092 (
		\u0_u1_csc_reg[8]/P0001 ,
		_w4183_,
		_w4743_,
		_w5052_
	);
	LUT3 #(
		.INIT('h15)
	) name4093 (
		\u0_rst_r2_reg/NET0131 ,
		_w4743_,
		_w5049_,
		_w5053_
	);
	LUT2 #(
		.INIT('h4)
	) name4094 (
		_w5052_,
		_w5053_,
		_w5054_
	);
	LUT3 #(
		.INIT('h15)
	) name4095 (
		\u0_u1_csc_reg[7]/P0001 ,
		_w4183_,
		_w4743_,
		_w5055_
	);
	LUT3 #(
		.INIT('h15)
	) name4096 (
		\u0_rst_r2_reg/NET0131 ,
		_w4743_,
		_w5017_,
		_w5056_
	);
	LUT2 #(
		.INIT('h4)
	) name4097 (
		_w5055_,
		_w5056_,
		_w5057_
	);
	LUT3 #(
		.INIT('h15)
	) name4098 (
		\u0_u1_csc_reg[9]/P0001 ,
		_w4183_,
		_w4743_,
		_w5058_
	);
	LUT4 #(
		.INIT('h0020)
	) name4099 (
		\u0_rf_we_reg/NET0131 ,
		\u0_u0_addr_r_reg[2]/P0001 ,
		\u0_u0_addr_r_reg[4]/P0001 ,
		\wb_data_i[9]_pad ,
		_w5059_
	);
	LUT3 #(
		.INIT('h15)
	) name4100 (
		\u0_rst_r2_reg/NET0131 ,
		_w4743_,
		_w5059_,
		_w5060_
	);
	LUT2 #(
		.INIT('h4)
	) name4101 (
		_w5058_,
		_w5060_,
		_w5061_
	);
	LUT3 #(
		.INIT('h15)
	) name4102 (
		\u0_u1_tms_reg[0]/P0001 ,
		_w4743_,
		_w4744_,
		_w5062_
	);
	LUT4 #(
		.INIT('h0080)
	) name4103 (
		\u0_rf_we_reg/NET0131 ,
		\u0_u0_addr_r_reg[2]/P0001 ,
		\u0_u0_addr_r_reg[4]/P0001 ,
		\wb_data_i[0]_pad ,
		_w5063_
	);
	LUT3 #(
		.INIT('h15)
	) name4104 (
		\u0_rst_r2_reg/NET0131 ,
		_w4743_,
		_w5063_,
		_w5064_
	);
	LUT2 #(
		.INIT('h4)
	) name4105 (
		_w5062_,
		_w5064_,
		_w5065_
	);
	LUT3 #(
		.INIT('h15)
	) name4106 (
		\u0_u1_tms_reg[30]/P0001 ,
		_w4743_,
		_w4744_,
		_w5066_
	);
	LUT4 #(
		.INIT('h0080)
	) name4107 (
		\u0_rf_we_reg/NET0131 ,
		\u0_u0_addr_r_reg[2]/P0001 ,
		\u0_u0_addr_r_reg[4]/P0001 ,
		\wb_data_i[30]_pad ,
		_w5067_
	);
	LUT3 #(
		.INIT('h15)
	) name4108 (
		\u0_rst_r2_reg/NET0131 ,
		_w4743_,
		_w5067_,
		_w5068_
	);
	LUT2 #(
		.INIT('h4)
	) name4109 (
		_w5066_,
		_w5068_,
		_w5069_
	);
	LUT3 #(
		.INIT('h15)
	) name4110 (
		\u0_u1_tms_reg[10]/P0001 ,
		_w4743_,
		_w4744_,
		_w5070_
	);
	LUT4 #(
		.INIT('h0080)
	) name4111 (
		\u0_rf_we_reg/NET0131 ,
		\u0_u0_addr_r_reg[2]/P0001 ,
		\u0_u0_addr_r_reg[4]/P0001 ,
		\wb_data_i[10]_pad ,
		_w5071_
	);
	LUT3 #(
		.INIT('h15)
	) name4112 (
		\u0_rst_r2_reg/NET0131 ,
		_w4743_,
		_w5071_,
		_w5072_
	);
	LUT2 #(
		.INIT('h4)
	) name4113 (
		_w5070_,
		_w5072_,
		_w5073_
	);
	LUT3 #(
		.INIT('h15)
	) name4114 (
		\u0_u1_tms_reg[11]/P0001 ,
		_w4743_,
		_w4744_,
		_w5074_
	);
	LUT4 #(
		.INIT('h0080)
	) name4115 (
		\u0_rf_we_reg/NET0131 ,
		\u0_u0_addr_r_reg[2]/P0001 ,
		\u0_u0_addr_r_reg[4]/P0001 ,
		\wb_data_i[11]_pad ,
		_w5075_
	);
	LUT3 #(
		.INIT('h15)
	) name4116 (
		\u0_rst_r2_reg/NET0131 ,
		_w4743_,
		_w5075_,
		_w5076_
	);
	LUT2 #(
		.INIT('h4)
	) name4117 (
		_w5074_,
		_w5076_,
		_w5077_
	);
	LUT3 #(
		.INIT('h15)
	) name4118 (
		\u0_u1_tms_reg[12]/P0001 ,
		_w4743_,
		_w4744_,
		_w5078_
	);
	LUT4 #(
		.INIT('h0080)
	) name4119 (
		\u0_rf_we_reg/NET0131 ,
		\u0_u0_addr_r_reg[2]/P0001 ,
		\u0_u0_addr_r_reg[4]/P0001 ,
		\wb_data_i[12]_pad ,
		_w5079_
	);
	LUT3 #(
		.INIT('h15)
	) name4120 (
		\u0_rst_r2_reg/NET0131 ,
		_w4743_,
		_w5079_,
		_w5080_
	);
	LUT2 #(
		.INIT('h4)
	) name4121 (
		_w5078_,
		_w5080_,
		_w5081_
	);
	LUT3 #(
		.INIT('h15)
	) name4122 (
		\u0_u1_tms_reg[13]/P0001 ,
		_w4743_,
		_w4744_,
		_w5082_
	);
	LUT4 #(
		.INIT('h0080)
	) name4123 (
		\u0_rf_we_reg/NET0131 ,
		\u0_u0_addr_r_reg[2]/P0001 ,
		\u0_u0_addr_r_reg[4]/P0001 ,
		\wb_data_i[13]_pad ,
		_w5083_
	);
	LUT3 #(
		.INIT('h15)
	) name4124 (
		\u0_rst_r2_reg/NET0131 ,
		_w4743_,
		_w5083_,
		_w5084_
	);
	LUT2 #(
		.INIT('h4)
	) name4125 (
		_w5082_,
		_w5084_,
		_w5085_
	);
	LUT3 #(
		.INIT('h15)
	) name4126 (
		\u0_u1_tms_reg[14]/P0001 ,
		_w4743_,
		_w4744_,
		_w5086_
	);
	LUT4 #(
		.INIT('h0080)
	) name4127 (
		\u0_rf_we_reg/NET0131 ,
		\u0_u0_addr_r_reg[2]/P0001 ,
		\u0_u0_addr_r_reg[4]/P0001 ,
		\wb_data_i[14]_pad ,
		_w5087_
	);
	LUT3 #(
		.INIT('h15)
	) name4128 (
		\u0_rst_r2_reg/NET0131 ,
		_w4743_,
		_w5087_,
		_w5088_
	);
	LUT2 #(
		.INIT('h4)
	) name4129 (
		_w5086_,
		_w5088_,
		_w5089_
	);
	LUT3 #(
		.INIT('h15)
	) name4130 (
		\u0_u1_tms_reg[15]/P0001 ,
		_w4743_,
		_w4744_,
		_w5090_
	);
	LUT4 #(
		.INIT('h0080)
	) name4131 (
		\u0_rf_we_reg/NET0131 ,
		\u0_u0_addr_r_reg[2]/P0001 ,
		\u0_u0_addr_r_reg[4]/P0001 ,
		\wb_data_i[15]_pad ,
		_w5091_
	);
	LUT3 #(
		.INIT('h15)
	) name4132 (
		\u0_rst_r2_reg/NET0131 ,
		_w4743_,
		_w5091_,
		_w5092_
	);
	LUT2 #(
		.INIT('h4)
	) name4133 (
		_w5090_,
		_w5092_,
		_w5093_
	);
	LUT3 #(
		.INIT('h15)
	) name4134 (
		\u0_u1_tms_reg[18]/P0001 ,
		_w4743_,
		_w4744_,
		_w5094_
	);
	LUT4 #(
		.INIT('h0080)
	) name4135 (
		\u0_rf_we_reg/NET0131 ,
		\u0_u0_addr_r_reg[2]/P0001 ,
		\u0_u0_addr_r_reg[4]/P0001 ,
		\wb_data_i[18]_pad ,
		_w5095_
	);
	LUT3 #(
		.INIT('h15)
	) name4136 (
		\u0_rst_r2_reg/NET0131 ,
		_w4743_,
		_w5095_,
		_w5096_
	);
	LUT2 #(
		.INIT('h4)
	) name4137 (
		_w5094_,
		_w5096_,
		_w5097_
	);
	LUT3 #(
		.INIT('h15)
	) name4138 (
		\u0_u1_tms_reg[20]/P0001 ,
		_w4743_,
		_w4744_,
		_w5098_
	);
	LUT4 #(
		.INIT('h0080)
	) name4139 (
		\u0_rf_we_reg/NET0131 ,
		\u0_u0_addr_r_reg[2]/P0001 ,
		\u0_u0_addr_r_reg[4]/P0001 ,
		\wb_data_i[20]_pad ,
		_w5099_
	);
	LUT3 #(
		.INIT('h15)
	) name4140 (
		\u0_rst_r2_reg/NET0131 ,
		_w4743_,
		_w5099_,
		_w5100_
	);
	LUT2 #(
		.INIT('h4)
	) name4141 (
		_w5098_,
		_w5100_,
		_w5101_
	);
	LUT3 #(
		.INIT('h15)
	) name4142 (
		\u0_u1_tms_reg[21]/P0001 ,
		_w4743_,
		_w4744_,
		_w5102_
	);
	LUT4 #(
		.INIT('h0080)
	) name4143 (
		\u0_rf_we_reg/NET0131 ,
		\u0_u0_addr_r_reg[2]/P0001 ,
		\u0_u0_addr_r_reg[4]/P0001 ,
		\wb_data_i[21]_pad ,
		_w5103_
	);
	LUT3 #(
		.INIT('h15)
	) name4144 (
		\u0_rst_r2_reg/NET0131 ,
		_w4743_,
		_w5103_,
		_w5104_
	);
	LUT2 #(
		.INIT('h4)
	) name4145 (
		_w5102_,
		_w5104_,
		_w5105_
	);
	LUT3 #(
		.INIT('h15)
	) name4146 (
		\u0_u1_tms_reg[24]/P0001 ,
		_w4743_,
		_w4744_,
		_w5106_
	);
	LUT4 #(
		.INIT('h0080)
	) name4147 (
		\u0_rf_we_reg/NET0131 ,
		\u0_u0_addr_r_reg[2]/P0001 ,
		\u0_u0_addr_r_reg[4]/P0001 ,
		\wb_data_i[24]_pad ,
		_w5107_
	);
	LUT3 #(
		.INIT('h15)
	) name4148 (
		\u0_rst_r2_reg/NET0131 ,
		_w4743_,
		_w5107_,
		_w5108_
	);
	LUT2 #(
		.INIT('h4)
	) name4149 (
		_w5106_,
		_w5108_,
		_w5109_
	);
	LUT3 #(
		.INIT('h15)
	) name4150 (
		\u0_u1_tms_reg[25]/P0001 ,
		_w4743_,
		_w4744_,
		_w5110_
	);
	LUT4 #(
		.INIT('h0080)
	) name4151 (
		\u0_rf_we_reg/NET0131 ,
		\u0_u0_addr_r_reg[2]/P0001 ,
		\u0_u0_addr_r_reg[4]/P0001 ,
		\wb_data_i[25]_pad ,
		_w5111_
	);
	LUT3 #(
		.INIT('h15)
	) name4152 (
		\u0_rst_r2_reg/NET0131 ,
		_w4743_,
		_w5111_,
		_w5112_
	);
	LUT2 #(
		.INIT('h4)
	) name4153 (
		_w5110_,
		_w5112_,
		_w5113_
	);
	LUT3 #(
		.INIT('h15)
	) name4154 (
		\u0_u1_tms_reg[27]/P0001 ,
		_w4743_,
		_w4744_,
		_w5114_
	);
	LUT4 #(
		.INIT('h0080)
	) name4155 (
		\u0_rf_we_reg/NET0131 ,
		\u0_u0_addr_r_reg[2]/P0001 ,
		\u0_u0_addr_r_reg[4]/P0001 ,
		\wb_data_i[27]_pad ,
		_w5115_
	);
	LUT3 #(
		.INIT('h15)
	) name4156 (
		\u0_rst_r2_reg/NET0131 ,
		_w4743_,
		_w5115_,
		_w5116_
	);
	LUT2 #(
		.INIT('h4)
	) name4157 (
		_w5114_,
		_w5116_,
		_w5117_
	);
	LUT3 #(
		.INIT('h15)
	) name4158 (
		\u0_u1_tms_reg[2]/P0001 ,
		_w4743_,
		_w4744_,
		_w5118_
	);
	LUT4 #(
		.INIT('h0080)
	) name4159 (
		\u0_rf_we_reg/NET0131 ,
		\u0_u0_addr_r_reg[2]/P0001 ,
		\u0_u0_addr_r_reg[4]/P0001 ,
		\wb_data_i[2]_pad ,
		_w5119_
	);
	LUT3 #(
		.INIT('h15)
	) name4160 (
		\u0_rst_r2_reg/NET0131 ,
		_w4743_,
		_w5119_,
		_w5120_
	);
	LUT2 #(
		.INIT('h4)
	) name4161 (
		_w5118_,
		_w5120_,
		_w5121_
	);
	LUT3 #(
		.INIT('h15)
	) name4162 (
		\u0_u1_tms_reg[31]/P0001 ,
		_w4743_,
		_w4744_,
		_w5122_
	);
	LUT4 #(
		.INIT('h0080)
	) name4163 (
		\u0_rf_we_reg/NET0131 ,
		\u0_u0_addr_r_reg[2]/P0001 ,
		\u0_u0_addr_r_reg[4]/P0001 ,
		\wb_data_i[31]_pad ,
		_w5123_
	);
	LUT3 #(
		.INIT('h15)
	) name4164 (
		\u0_rst_r2_reg/NET0131 ,
		_w4743_,
		_w5123_,
		_w5124_
	);
	LUT2 #(
		.INIT('h4)
	) name4165 (
		_w5122_,
		_w5124_,
		_w5125_
	);
	LUT3 #(
		.INIT('h15)
	) name4166 (
		\u0_u0_csc_reg[23]/P0001 ,
		_w4182_,
		_w4183_,
		_w5126_
	);
	LUT3 #(
		.INIT('h15)
	) name4167 (
		\u0_rst_r2_reg/NET0131 ,
		_w4182_,
		_w4995_,
		_w5127_
	);
	LUT2 #(
		.INIT('h4)
	) name4168 (
		_w5126_,
		_w5127_,
		_w5128_
	);
	LUT3 #(
		.INIT('h15)
	) name4169 (
		\u0_u1_tms_reg[3]/P0001 ,
		_w4743_,
		_w4744_,
		_w5129_
	);
	LUT4 #(
		.INIT('h0080)
	) name4170 (
		\u0_rf_we_reg/NET0131 ,
		\u0_u0_addr_r_reg[2]/P0001 ,
		\u0_u0_addr_r_reg[4]/P0001 ,
		\wb_data_i[3]_pad ,
		_w5130_
	);
	LUT3 #(
		.INIT('h15)
	) name4171 (
		\u0_rst_r2_reg/NET0131 ,
		_w4743_,
		_w5130_,
		_w5131_
	);
	LUT2 #(
		.INIT('h4)
	) name4172 (
		_w5129_,
		_w5131_,
		_w5132_
	);
	LUT3 #(
		.INIT('h15)
	) name4173 (
		\u0_u1_tms_reg[5]/P0001 ,
		_w4743_,
		_w4744_,
		_w5133_
	);
	LUT4 #(
		.INIT('h0080)
	) name4174 (
		\u0_rf_we_reg/NET0131 ,
		\u0_u0_addr_r_reg[2]/P0001 ,
		\u0_u0_addr_r_reg[4]/P0001 ,
		\wb_data_i[5]_pad ,
		_w5134_
	);
	LUT3 #(
		.INIT('h15)
	) name4175 (
		\u0_rst_r2_reg/NET0131 ,
		_w4743_,
		_w5134_,
		_w5135_
	);
	LUT2 #(
		.INIT('h4)
	) name4176 (
		_w5133_,
		_w5135_,
		_w5136_
	);
	LUT3 #(
		.INIT('h15)
	) name4177 (
		\u0_u1_tms_reg[8]/P0001 ,
		_w4743_,
		_w4744_,
		_w5137_
	);
	LUT4 #(
		.INIT('h0080)
	) name4178 (
		\u0_rf_we_reg/NET0131 ,
		\u0_u0_addr_r_reg[2]/P0001 ,
		\u0_u0_addr_r_reg[4]/P0001 ,
		\wb_data_i[8]_pad ,
		_w5138_
	);
	LUT3 #(
		.INIT('h15)
	) name4179 (
		\u0_rst_r2_reg/NET0131 ,
		_w4743_,
		_w5138_,
		_w5139_
	);
	LUT2 #(
		.INIT('h4)
	) name4180 (
		_w5137_,
		_w5139_,
		_w5140_
	);
	LUT3 #(
		.INIT('h15)
	) name4181 (
		\u0_u1_tms_reg[9]/P0001 ,
		_w4743_,
		_w4744_,
		_w5141_
	);
	LUT4 #(
		.INIT('h0080)
	) name4182 (
		\u0_rf_we_reg/NET0131 ,
		\u0_u0_addr_r_reg[2]/P0001 ,
		\u0_u0_addr_r_reg[4]/P0001 ,
		\wb_data_i[9]_pad ,
		_w5142_
	);
	LUT3 #(
		.INIT('h15)
	) name4183 (
		\u0_rst_r2_reg/NET0131 ,
		_w4743_,
		_w5142_,
		_w5143_
	);
	LUT2 #(
		.INIT('h4)
	) name4184 (
		_w5141_,
		_w5143_,
		_w5144_
	);
	LUT3 #(
		.INIT('h2a)
	) name4185 (
		\u0_u0_tms_reg[20]/P0001 ,
		_w4182_,
		_w4744_,
		_w5145_
	);
	LUT4 #(
		.INIT('h8000)
	) name4186 (
		\u0_rf_we_reg/NET0131 ,
		\u0_u0_addr_r_reg[2]/P0001 ,
		\u0_u0_addr_r_reg[4]/P0001 ,
		\wb_data_i[20]_pad ,
		_w5146_
	);
	LUT3 #(
		.INIT('h15)
	) name4187 (
		\u0_rst_r2_reg/NET0131 ,
		_w4182_,
		_w5146_,
		_w5147_
	);
	LUT2 #(
		.INIT('hb)
	) name4188 (
		_w5145_,
		_w5147_,
		_w5148_
	);
	LUT3 #(
		.INIT('h15)
	) name4189 (
		\u0_u1_tms_reg[1]/P0001 ,
		_w4743_,
		_w4744_,
		_w5149_
	);
	LUT4 #(
		.INIT('h0080)
	) name4190 (
		\u0_rf_we_reg/NET0131 ,
		\u0_u0_addr_r_reg[2]/P0001 ,
		\u0_u0_addr_r_reg[4]/P0001 ,
		\wb_data_i[1]_pad ,
		_w5150_
	);
	LUT3 #(
		.INIT('h15)
	) name4191 (
		\u0_rst_r2_reg/NET0131 ,
		_w4743_,
		_w5150_,
		_w5151_
	);
	LUT2 #(
		.INIT('h4)
	) name4192 (
		_w5149_,
		_w5151_,
		_w5152_
	);
	LUT3 #(
		.INIT('h15)
	) name4193 (
		\u0_u1_tms_reg[6]/P0001 ,
		_w4743_,
		_w4744_,
		_w5153_
	);
	LUT4 #(
		.INIT('h0080)
	) name4194 (
		\u0_rf_we_reg/NET0131 ,
		\u0_u0_addr_r_reg[2]/P0001 ,
		\u0_u0_addr_r_reg[4]/P0001 ,
		\wb_data_i[6]_pad ,
		_w5154_
	);
	LUT3 #(
		.INIT('h15)
	) name4195 (
		\u0_rst_r2_reg/NET0131 ,
		_w4743_,
		_w5154_,
		_w5155_
	);
	LUT2 #(
		.INIT('h4)
	) name4196 (
		_w5153_,
		_w5155_,
		_w5156_
	);
	LUT3 #(
		.INIT('h15)
	) name4197 (
		\u0_u1_tms_reg[29]/P0001 ,
		_w4743_,
		_w4744_,
		_w5157_
	);
	LUT4 #(
		.INIT('h0080)
	) name4198 (
		\u0_rf_we_reg/NET0131 ,
		\u0_u0_addr_r_reg[2]/P0001 ,
		\u0_u0_addr_r_reg[4]/P0001 ,
		\wb_data_i[29]_pad ,
		_w5158_
	);
	LUT3 #(
		.INIT('h15)
	) name4199 (
		\u0_rst_r2_reg/NET0131 ,
		_w4743_,
		_w5158_,
		_w5159_
	);
	LUT2 #(
		.INIT('h4)
	) name4200 (
		_w5157_,
		_w5159_,
		_w5160_
	);
	LUT3 #(
		.INIT('h15)
	) name4201 (
		\u0_u1_tms_reg[28]/P0001 ,
		_w4743_,
		_w4744_,
		_w5161_
	);
	LUT4 #(
		.INIT('h0080)
	) name4202 (
		\u0_rf_we_reg/NET0131 ,
		\u0_u0_addr_r_reg[2]/P0001 ,
		\u0_u0_addr_r_reg[4]/P0001 ,
		\wb_data_i[28]_pad ,
		_w5162_
	);
	LUT3 #(
		.INIT('h15)
	) name4203 (
		\u0_rst_r2_reg/NET0131 ,
		_w4743_,
		_w5162_,
		_w5163_
	);
	LUT2 #(
		.INIT('h4)
	) name4204 (
		_w5161_,
		_w5163_,
		_w5164_
	);
	LUT3 #(
		.INIT('h15)
	) name4205 (
		\u0_u1_tms_reg[4]/P0001 ,
		_w4743_,
		_w4744_,
		_w5165_
	);
	LUT4 #(
		.INIT('h0080)
	) name4206 (
		\u0_rf_we_reg/NET0131 ,
		\u0_u0_addr_r_reg[2]/P0001 ,
		\u0_u0_addr_r_reg[4]/P0001 ,
		\wb_data_i[4]_pad ,
		_w5166_
	);
	LUT3 #(
		.INIT('h15)
	) name4207 (
		\u0_rst_r2_reg/NET0131 ,
		_w4743_,
		_w5166_,
		_w5167_
	);
	LUT2 #(
		.INIT('h4)
	) name4208 (
		_w5165_,
		_w5167_,
		_w5168_
	);
	LUT3 #(
		.INIT('h15)
	) name4209 (
		\u0_u0_csc_reg[10]/P0001 ,
		_w4182_,
		_w4183_,
		_w5169_
	);
	LUT3 #(
		.INIT('h15)
	) name4210 (
		\u0_rst_r2_reg/NET0131 ,
		_w4182_,
		_w4952_,
		_w5170_
	);
	LUT2 #(
		.INIT('h4)
	) name4211 (
		_w5169_,
		_w5170_,
		_w5171_
	);
	LUT3 #(
		.INIT('h15)
	) name4212 (
		\u0_u1_tms_reg[26]/P0001 ,
		_w4743_,
		_w4744_,
		_w5172_
	);
	LUT4 #(
		.INIT('h0080)
	) name4213 (
		\u0_rf_we_reg/NET0131 ,
		\u0_u0_addr_r_reg[2]/P0001 ,
		\u0_u0_addr_r_reg[4]/P0001 ,
		\wb_data_i[26]_pad ,
		_w5173_
	);
	LUT3 #(
		.INIT('h15)
	) name4214 (
		\u0_rst_r2_reg/NET0131 ,
		_w4743_,
		_w5173_,
		_w5174_
	);
	LUT2 #(
		.INIT('h4)
	) name4215 (
		_w5172_,
		_w5174_,
		_w5175_
	);
	LUT3 #(
		.INIT('h15)
	) name4216 (
		\u0_u1_csc_reg[16]/P0001 ,
		_w4183_,
		_w4743_,
		_w5176_
	);
	LUT3 #(
		.INIT('h15)
	) name4217 (
		\u0_rst_r2_reg/NET0131 ,
		_w4743_,
		_w4759_,
		_w5177_
	);
	LUT2 #(
		.INIT('h4)
	) name4218 (
		_w5176_,
		_w5177_,
		_w5178_
	);
	LUT3 #(
		.INIT('h15)
	) name4219 (
		\u0_u0_csc_reg[18]/P0001 ,
		_w4182_,
		_w4183_,
		_w5179_
	);
	LUT3 #(
		.INIT('h15)
	) name4220 (
		\u0_rst_r2_reg/NET0131 ,
		_w4182_,
		_w4974_,
		_w5180_
	);
	LUT2 #(
		.INIT('h4)
	) name4221 (
		_w5179_,
		_w5180_,
		_w5181_
	);
	LUT3 #(
		.INIT('h15)
	) name4222 (
		\u0_u0_csc_reg[31]/P0001 ,
		_w4182_,
		_w4183_,
		_w5182_
	);
	LUT3 #(
		.INIT('h15)
	) name4223 (
		\u0_rst_r2_reg/NET0131 ,
		_w4182_,
		_w5030_,
		_w5183_
	);
	LUT2 #(
		.INIT('h4)
	) name4224 (
		_w5182_,
		_w5183_,
		_w5184_
	);
	LUT3 #(
		.INIT('h2a)
	) name4225 (
		\u0_u0_tms_reg[31]/P0001 ,
		_w4182_,
		_w4744_,
		_w5185_
	);
	LUT4 #(
		.INIT('h8000)
	) name4226 (
		\u0_rf_we_reg/NET0131 ,
		\u0_u0_addr_r_reg[2]/P0001 ,
		\u0_u0_addr_r_reg[4]/P0001 ,
		\wb_data_i[31]_pad ,
		_w5186_
	);
	LUT3 #(
		.INIT('h15)
	) name4227 (
		\u0_rst_r2_reg/NET0131 ,
		_w4182_,
		_w5186_,
		_w5187_
	);
	LUT2 #(
		.INIT('hb)
	) name4228 (
		_w5185_,
		_w5187_,
		_w5188_
	);
	LUT3 #(
		.INIT('h15)
	) name4229 (
		\u0_u1_tms_reg[7]/P0001 ,
		_w4743_,
		_w4744_,
		_w5189_
	);
	LUT4 #(
		.INIT('h0080)
	) name4230 (
		\u0_rf_we_reg/NET0131 ,
		\u0_u0_addr_r_reg[2]/P0001 ,
		\u0_u0_addr_r_reg[4]/P0001 ,
		\wb_data_i[7]_pad ,
		_w5190_
	);
	LUT3 #(
		.INIT('h15)
	) name4231 (
		\u0_rst_r2_reg/NET0131 ,
		_w4743_,
		_w5190_,
		_w5191_
	);
	LUT2 #(
		.INIT('h4)
	) name4232 (
		_w5189_,
		_w5191_,
		_w5192_
	);
	LUT3 #(
		.INIT('h15)
	) name4233 (
		\u0_u0_csc_reg[19]/P0001 ,
		_w4182_,
		_w4183_,
		_w5193_
	);
	LUT3 #(
		.INIT('h15)
	) name4234 (
		\u0_rst_r2_reg/NET0131 ,
		_w4182_,
		_w4978_,
		_w5194_
	);
	LUT2 #(
		.INIT('h4)
	) name4235 (
		_w5193_,
		_w5194_,
		_w5195_
	);
	LUT3 #(
		.INIT('h15)
	) name4236 (
		\u0_u0_csc_reg[6]/P0001 ,
		_w4182_,
		_w4183_,
		_w5196_
	);
	LUT3 #(
		.INIT('h15)
	) name4237 (
		\u0_rst_r2_reg/NET0131 ,
		_w4182_,
		_w5045_,
		_w5197_
	);
	LUT2 #(
		.INIT('h4)
	) name4238 (
		_w5196_,
		_w5197_,
		_w5198_
	);
	LUT3 #(
		.INIT('h15)
	) name4239 (
		\u0_u0_csc_reg[9]/P0001 ,
		_w4182_,
		_w4183_,
		_w5199_
	);
	LUT3 #(
		.INIT('h15)
	) name4240 (
		\u0_rst_r2_reg/NET0131 ,
		_w4182_,
		_w5059_,
		_w5200_
	);
	LUT2 #(
		.INIT('h4)
	) name4241 (
		_w5199_,
		_w5200_,
		_w5201_
	);
	LUT4 #(
		.INIT('h7f80)
	) name4242 (
		\u1_acs_addr_reg[0]/P0001 ,
		\u1_acs_addr_reg[1]/P0001 ,
		\u1_acs_addr_reg[2]/P0001 ,
		\u1_acs_addr_reg[3]/P0001 ,
		_w5202_
	);
	LUT3 #(
		.INIT('hea)
	) name4243 (
		\u0_u1_inited_reg/NET0131 ,
		_w976_,
		_w4452_,
		_w5203_
	);
	LUT3 #(
		.INIT('hea)
	) name4244 (
		\u0_u0_inited_reg/NET0131 ,
		_w976_,
		_w4447_,
		_w5204_
	);
	LUT4 #(
		.INIT('hfa32)
	) name4245 (
		\u0_init_req_reg/NET0131 ,
		\u0_lmr_ack_r_reg/P0001 ,
		\u0_lmr_req_reg/NET0131 ,
		\u5_lmr_ack_reg/NET0131 ,
		_w5205_
	);
	LUT3 #(
		.INIT('h8f)
	) name4246 (
		_w976_,
		_w4446_,
		_w5205_,
		_w5206_
	);
	LUT3 #(
		.INIT('h70)
	) name4247 (
		_w1014_,
		_w1015_,
		_w1133_,
		_w5207_
	);
	LUT3 #(
		.INIT('h15)
	) name4248 (
		\u6_read_go_r_reg/NET0131 ,
		_w1130_,
		_w1748_,
		_w5208_
	);
	LUT2 #(
		.INIT('h2)
	) name4249 (
		_w5207_,
		_w5208_,
		_w5209_
	);
	LUT3 #(
		.INIT('hf8)
	) name4250 (
		_w1748_,
		_w2366_,
		_w2367_,
		_w5210_
	);
	LUT4 #(
		.INIT('h1555)
	) name4251 (
		\u1_acs_addr_reg[9]/P0001 ,
		_w3563_,
		_w3564_,
		_w4139_,
		_w5211_
	);
	LUT2 #(
		.INIT('h1)
	) name4252 (
		_w3566_,
		_w5211_,
		_w5212_
	);
	LUT2 #(
		.INIT('h9)
	) name4253 (
		\wb_data_i[11]_pad ,
		\wb_data_i[13]_pad ,
		_w5213_
	);
	LUT3 #(
		.INIT('h96)
	) name4254 (
		\wb_data_i[15]_pad ,
		\wb_data_i[8]_pad ,
		\wb_data_i[9]_pad ,
		_w5214_
	);
	LUT3 #(
		.INIT('h69)
	) name4255 (
		\wb_data_i[10]_pad ,
		\wb_data_i[12]_pad ,
		\wb_data_i[14]_pad ,
		_w5215_
	);
	LUT3 #(
		.INIT('h96)
	) name4256 (
		_w5213_,
		_w5214_,
		_w5215_,
		_w5216_
	);
	LUT2 #(
		.INIT('h9)
	) name4257 (
		\wb_data_i[1]_pad ,
		\wb_data_i[6]_pad ,
		_w5217_
	);
	LUT3 #(
		.INIT('h96)
	) name4258 (
		\wb_data_i[2]_pad ,
		\wb_data_i[4]_pad ,
		\wb_data_i[5]_pad ,
		_w5218_
	);
	LUT3 #(
		.INIT('h69)
	) name4259 (
		\wb_data_i[0]_pad ,
		\wb_data_i[3]_pad ,
		\wb_data_i[7]_pad ,
		_w5219_
	);
	LUT3 #(
		.INIT('h96)
	) name4260 (
		_w5217_,
		_w5218_,
		_w5219_,
		_w5220_
	);
	LUT2 #(
		.INIT('h9)
	) name4261 (
		\wb_data_i[27]_pad ,
		\wb_data_i[29]_pad ,
		_w5221_
	);
	LUT3 #(
		.INIT('h96)
	) name4262 (
		\wb_data_i[24]_pad ,
		\wb_data_i[30]_pad ,
		\wb_data_i[31]_pad ,
		_w5222_
	);
	LUT3 #(
		.INIT('h69)
	) name4263 (
		\wb_data_i[25]_pad ,
		\wb_data_i[26]_pad ,
		\wb_data_i[28]_pad ,
		_w5223_
	);
	LUT3 #(
		.INIT('h96)
	) name4264 (
		_w5221_,
		_w5222_,
		_w5223_,
		_w5224_
	);
	LUT2 #(
		.INIT('h9)
	) name4265 (
		\wb_data_i[17]_pad ,
		\wb_data_i[22]_pad ,
		_w5225_
	);
	LUT3 #(
		.INIT('h96)
	) name4266 (
		\wb_data_i[16]_pad ,
		\wb_data_i[21]_pad ,
		\wb_data_i[23]_pad ,
		_w5226_
	);
	LUT3 #(
		.INIT('h69)
	) name4267 (
		\wb_data_i[18]_pad ,
		\wb_data_i[19]_pad ,
		\wb_data_i[20]_pad ,
		_w5227_
	);
	LUT3 #(
		.INIT('h96)
	) name4268 (
		_w5225_,
		_w5226_,
		_w5227_,
		_w5228_
	);
	LUT2 #(
		.INIT('h8)
	) name4269 (
		\u6_write_go_r_reg/NET0131 ,
		wb_cyc_i_pad,
		_w5229_
	);
	LUT3 #(
		.INIT('hec)
	) name4270 (
		_w1748_,
		_w5229_,
		_w1014_,
		_w5230_
	);
	LUT4 #(
		.INIT('h084c)
	) name4271 (
		\u0_init_req_reg/NET0131 ,
		\u0_sreq_cs_le_reg/NET0131 ,
		\u0_u1_init_req_reg/NET0131 ,
		\u0_u1_lmr_req_reg/NET0131 ,
		_w5231_
	);
	LUT2 #(
		.INIT('h1)
	) name4272 (
		\u0_spec_req_cs_reg[1]/NET0131 ,
		\u0_sreq_cs_le_reg/NET0131 ,
		_w5232_
	);
	LUT4 #(
		.INIT('hc480)
	) name4273 (
		\u0_init_req_reg/NET0131 ,
		\u0_sreq_cs_le_reg/NET0131 ,
		\u0_u0_init_req_reg/NET0131 ,
		\u0_u0_lmr_req_reg/NET0131 ,
		_w5233_
	);
	LUT3 #(
		.INIT('h01)
	) name4274 (
		_w5231_,
		_w5232_,
		_w5233_,
		_w5234_
	);
	LUT3 #(
		.INIT('h78)
	) name4275 (
		\u1_acs_addr_reg[0]/P0001 ,
		\u1_acs_addr_reg[1]/P0001 ,
		\u1_acs_addr_reg[2]/P0001 ,
		_w5235_
	);
	LUT3 #(
		.INIT('h6c)
	) name4276 (
		\u1_acs_addr_reg[4]/P0001 ,
		\u1_acs_addr_reg[5]/P0001 ,
		_w3563_,
		_w5236_
	);
	LUT2 #(
		.INIT('h1)
	) name4277 (
		suspended_o_pad,
		\u0_csr_r_reg[2]/NET0131 ,
		_w5237_
	);
	LUT4 #(
		.INIT('h4000)
	) name4278 (
		\u0_rf_we_reg/NET0131 ,
		wb_cyc_i_pad,
		wb_stb_i_pad,
		wb_we_i_pad,
		_w5238_
	);
	LUT2 #(
		.INIT('h8)
	) name4279 (
		_w1884_,
		_w5238_,
		_w5239_
	);
	LUT3 #(
		.INIT('h80)
	) name4280 (
		\u5_lookup_ready1_reg/NET0131 ,
		wb_cyc_i_pad,
		wb_stb_i_pad,
		_w5240_
	);
	LUT3 #(
		.INIT('h02)
	) name4281 (
		\u0_rf_we_reg/NET0131 ,
		\u0_u0_addr_r_reg[2]/P0001 ,
		\u0_u0_addr_r_reg[4]/P0001 ,
		_w5241_
	);
	LUT2 #(
		.INIT('h8)
	) name4282 (
		_w4182_,
		_w5241_,
		_w5242_
	);
	LUT2 #(
		.INIT('h8)
	) name4283 (
		_w4743_,
		_w5241_,
		_w5243_
	);
	LUT2 #(
		.INIT('h2)
	) name4284 (
		\u0_spec_req_cs_reg[0]/NET0131 ,
		\u0_sreq_cs_le_reg/NET0131 ,
		_w5244_
	);
	LUT2 #(
		.INIT('he)
	) name4285 (
		_w5233_,
		_w5244_,
		_w5245_
	);
	LUT4 #(
		.INIT('hfffe)
	) name4286 (
		\mem_ack_r_reg/P0001 ,
		\u0_csc_reg[1]/NET0131 ,
		\u0_csc_reg[2]/NET0131 ,
		\u0_csc_reg[3]/NET0131 ,
		_w5246_
	);
	LUT2 #(
		.INIT('hb)
	) name4287 (
		\u5_state_reg[26]/NET0131 ,
		_w976_,
		_w5247_
	);
	LUT2 #(
		.INIT('he)
	) name4288 (
		_w1531_,
		_w1577_,
		_w5248_
	);
	LUT4 #(
		.INIT('hea2a)
	) name4289 (
		\u6_wr_hold_reg/NET0131 ,
		wb_cyc_i_pad,
		wb_stb_i_pad,
		wb_we_i_pad,
		_w5249_
	);
	LUT2 #(
		.INIT('h6)
	) name4290 (
		\u1_acs_addr_reg[0]/P0001 ,
		\u1_acs_addr_reg[1]/P0001 ,
		_w5250_
	);
	LUT3 #(
		.INIT('hec)
	) name4291 (
		\u6_rmw_en_reg/NET0131 ,
		wb_ack_o_pad,
		wb_cyc_i_pad,
		_w5251_
	);
	LUT3 #(
		.INIT('hac)
	) name4292 (
		\u5_cmd_asserted2_reg/NET0131 ,
		\u5_cmd_asserted_reg/NET0131 ,
		\u5_mc_le_reg/NET0131 ,
		_w5252_
	);
	LUT2 #(
		.INIT('he)
	) name4293 (
		\u0_u0_lmr_req_reg/NET0131 ,
		\u0_u1_lmr_req_reg/NET0131 ,
		_w5253_
	);
	LUT2 #(
		.INIT('he)
	) name4294 (
		\u0_u0_init_req_reg/NET0131 ,
		\u0_u1_init_req_reg/NET0131 ,
		_w5254_
	);
	LUT2 #(
		.INIT('h6)
	) name4295 (
		\u5_state_reg[1]/NET0131 ,
		\u5_state_reg[54]/NET0131 ,
		_w5255_
	);
	LUT2 #(
		.INIT('h9)
	) name4296 (
		\u5_state_reg[36]/NET0131 ,
		\u5_state_reg[37]/NET0131 ,
		_w5256_
	);
	LUT3 #(
		.INIT('h04)
	) name4297 (
		\u5_state_reg[0]/NET0131 ,
		_w985_,
		_w5256_,
		_w5257_
	);
	LUT3 #(
		.INIT('h80)
	) name4298 (
		_w966_,
		_w1018_,
		_w5257_,
		_w5258_
	);
	LUT4 #(
		.INIT('h070f)
	) name4299 (
		_w966_,
		_w1018_,
		_w1031_,
		_w5257_,
		_w5259_
	);
	LUT3 #(
		.INIT('h09)
	) name4300 (
		\u5_state_reg[44]/NET0131 ,
		\u5_state_reg[45]/NET0131 ,
		\u5_state_reg[46]/NET0131 ,
		_w5260_
	);
	LUT3 #(
		.INIT('h01)
	) name4301 (
		\u5_state_reg[47]/NET0131 ,
		\u5_state_reg[48]/NET0131 ,
		\u5_state_reg[49]/NET0131 ,
		_w5261_
	);
	LUT3 #(
		.INIT('he0)
	) name4302 (
		\u5_state_reg[44]/NET0131 ,
		\u5_state_reg[45]/NET0131 ,
		\u5_state_reg[46]/NET0131 ,
		_w5262_
	);
	LUT3 #(
		.INIT('h04)
	) name4303 (
		_w5260_,
		_w5261_,
		_w5262_,
		_w5263_
	);
	LUT3 #(
		.INIT('h80)
	) name4304 (
		_w1183_,
		_w1235_,
		_w5263_,
		_w5264_
	);
	LUT2 #(
		.INIT('h9)
	) name4305 (
		\u5_state_reg[52]/NET0131 ,
		\u5_state_reg[53]/NET0131 ,
		_w5265_
	);
	LUT3 #(
		.INIT('h08)
	) name4306 (
		_w985_,
		_w988_,
		_w5265_,
		_w5266_
	);
	LUT2 #(
		.INIT('h9)
	) name4307 (
		\u5_state_reg[60]/NET0131 ,
		\u5_state_reg[61]/NET0131 ,
		_w5267_
	);
	LUT3 #(
		.INIT('h08)
	) name4308 (
		_w985_,
		_w1175_,
		_w5267_,
		_w5268_
	);
	LUT4 #(
		.INIT('h8000)
	) name4309 (
		_w970_,
		_w992_,
		_w999_,
		_w1238_,
		_w5269_
	);
	LUT4 #(
		.INIT('ha800)
	) name4310 (
		_w1235_,
		_w5266_,
		_w5268_,
		_w5269_,
		_w5270_
	);
	LUT4 #(
		.INIT('h9f8e)
	) name4311 (
		\u5_state_reg[42]/NET0131 ,
		\u5_state_reg[43]/NET0131 ,
		_w963_,
		_w1220_,
		_w5271_
	);
	LUT3 #(
		.INIT('h80)
	) name4312 (
		_w970_,
		_w993_,
		_w999_,
		_w5272_
	);
	LUT3 #(
		.INIT('h80)
	) name4313 (
		_w985_,
		_w988_,
		_w1238_,
		_w5273_
	);
	LUT3 #(
		.INIT('h40)
	) name4314 (
		_w5271_,
		_w5272_,
		_w5273_,
		_w5274_
	);
	LUT4 #(
		.INIT('h0001)
	) name4315 (
		_w5258_,
		_w5264_,
		_w5270_,
		_w5274_,
		_w5275_
	);
	LUT4 #(
		.INIT('h0080)
	) name4316 (
		_w1029_,
		_w3852_,
		_w4440_,
		_w5255_,
		_w5276_
	);
	LUT3 #(
		.INIT('h10)
	) name4317 (
		_w5259_,
		_w5275_,
		_w5276_,
		_w5277_
	);
	LUT4 #(
		.INIT('h5455)
	) name4318 (
		_w5255_,
		_w5259_,
		_w5275_,
		_w5276_,
		_w5278_
	);
	LUT4 #(
		.INIT('h1500)
	) name4319 (
		\u5_state_reg[1]/NET0131 ,
		_w1014_,
		_w1015_,
		_w1565_,
		_w5279_
	);
	LUT2 #(
		.INIT('h4)
	) name4320 (
		_w1608_,
		_w5279_,
		_w5280_
	);
	LUT3 #(
		.INIT('hb0)
	) name4321 (
		_w1539_,
		_w1599_,
		_w5280_,
		_w5281_
	);
	LUT2 #(
		.INIT('h1)
	) name4322 (
		\u4_rfr_req_reg/NET0131 ,
		\u5_state_reg[54]/NET0131 ,
		_w5282_
	);
	LUT3 #(
		.INIT('h20)
	) name4323 (
		_w1343_,
		_w1571_,
		_w5282_,
		_w5283_
	);
	LUT2 #(
		.INIT('h8)
	) name4324 (
		_w1631_,
		_w5283_,
		_w5284_
	);
	LUT2 #(
		.INIT('h1)
	) name4325 (
		_w5277_,
		_w5284_,
		_w5285_
	);
	LUT3 #(
		.INIT('hba)
	) name4326 (
		_w5278_,
		_w5281_,
		_w5285_,
		_w5286_
	);
	LUT2 #(
		.INIT('h1)
	) name4327 (
		\u5_cmd_asserted_reg/NET0131 ,
		\u5_state_reg[10]/NET0131 ,
		_w5287_
	);
	LUT3 #(
		.INIT('h08)
	) name4328 (
		_w1100_,
		_w1104_,
		_w5287_,
		_w5288_
	);
	LUT3 #(
		.INIT('h02)
	) name4329 (
		\u5_state_reg[10]/NET0131 ,
		\u5_state_reg[11]/NET0131 ,
		\u5_tmr_done_reg/NET0131 ,
		_w5289_
	);
	LUT3 #(
		.INIT('h80)
	) name4330 (
		_w1002_,
		_w1005_,
		_w5289_,
		_w5290_
	);
	LUT2 #(
		.INIT('he)
	) name4331 (
		_w5288_,
		_w5290_,
		_w5291_
	);
	LUT3 #(
		.INIT('h80)
	) name4332 (
		\u5_tmr_done_reg/NET0131 ,
		_w1068_,
		_w1201_,
		_w5292_
	);
	LUT3 #(
		.INIT('h40)
	) name4333 (
		\u5_cmd_asserted_reg/NET0131 ,
		_w1068_,
		_w1070_,
		_w5293_
	);
	LUT2 #(
		.INIT('he)
	) name4334 (
		_w5292_,
		_w5293_,
		_w5294_
	);
	LUT4 #(
		.INIT('hcc40)
	) name4335 (
		\u5_tmr_done_reg/NET0131 ,
		_w1035_,
		_w1228_,
		_w3900_,
		_w5295_
	);
	LUT2 #(
		.INIT('h4)
	) name4336 (
		\u5_cmd_asserted_reg/NET0131 ,
		_w1284_,
		_w5296_
	);
	LUT3 #(
		.INIT('h80)
	) name4337 (
		_w984_,
		_w1046_,
		_w5296_,
		_w5297_
	);
	LUT3 #(
		.INIT('ha8)
	) name4338 (
		_w1035_,
		_w1097_,
		_w5297_,
		_w5298_
	);
	LUT3 #(
		.INIT('h53)
	) name4339 (
		\u5_ir_cnt_done_reg/P0001 ,
		\u5_state_reg[26]/NET0131 ,
		\u5_tmr_done_reg/NET0131 ,
		_w5299_
	);
	LUT3 #(
		.INIT('h08)
	) name4340 (
		_w1035_,
		_w1228_,
		_w5299_,
		_w5300_
	);
	LUT3 #(
		.INIT('h40)
	) name4341 (
		\u5_cmd_asserted_reg/NET0131 ,
		_w1068_,
		_w1155_,
		_w5301_
	);
	LUT2 #(
		.INIT('he)
	) name4342 (
		_w5300_,
		_w5301_,
		_w5302_
	);
	LUT2 #(
		.INIT('h1)
	) name4343 (
		\u5_state_reg[38]/NET0131 ,
		\u5_tmr2_done_reg/NET0131 ,
		_w5303_
	);
	LUT3 #(
		.INIT('h2a)
	) name4344 (
		\u5_tmr2_done_reg/NET0131 ,
		_w976_,
		_w1975_,
		_w5304_
	);
	LUT3 #(
		.INIT('h23)
	) name4345 (
		_w1974_,
		_w5303_,
		_w5304_,
		_w5305_
	);
	LUT3 #(
		.INIT('h80)
	) name4346 (
		_w1041_,
		_w1195_,
		_w5305_,
		_w5306_
	);
	LUT3 #(
		.INIT('h08)
	) name4347 (
		_w1333_,
		_w1335_,
		_w1338_,
		_w5307_
	);
	LUT2 #(
		.INIT('h4)
	) name4348 (
		_w1571_,
		_w5307_,
		_w5308_
	);
	LUT4 #(
		.INIT('h33f7)
	) name4349 (
		\u5_state_reg[36]/NET0131 ,
		_w1581_,
		_w2021_,
		_w5308_,
		_w5309_
	);
	LUT3 #(
		.INIT('h8c)
	) name4350 (
		\u5_cmd_asserted2_reg/NET0131 ,
		\u5_state_reg[36]/NET0131 ,
		\u7_mc_br_r_reg/P0001 ,
		_w5310_
	);
	LUT4 #(
		.INIT('h4f00)
	) name4351 (
		_w1533_,
		_w1579_,
		_w1580_,
		_w5310_,
		_w5311_
	);
	LUT3 #(
		.INIT('ha2)
	) name4352 (
		_w1586_,
		_w5309_,
		_w5311_,
		_w5312_
	);
	LUT3 #(
		.INIT('h10)
	) name4353 (
		\u5_cmd_asserted_reg/NET0131 ,
		\u5_state_reg[12]/NET0131 ,
		\u5_state_reg[13]/NET0131 ,
		_w5313_
	);
	LUT3 #(
		.INIT('h80)
	) name4354 (
		_w1002_,
		_w1143_,
		_w5313_,
		_w5314_
	);
	LUT3 #(
		.INIT('ha2)
	) name4355 (
		\u5_state_reg[13]/NET0131 ,
		\u5_tmr_done_reg/NET0131 ,
		\u5_wb_wait_r_reg/P0001 ,
		_w5315_
	);
	LUT2 #(
		.INIT('h1)
	) name4356 (
		_w1270_,
		_w5315_,
		_w5316_
	);
	LUT3 #(
		.INIT('h08)
	) name4357 (
		_w1100_,
		_w1110_,
		_w5316_,
		_w5317_
	);
	LUT3 #(
		.INIT('hfe)
	) name4358 (
		_w1136_,
		_w5314_,
		_w5317_,
		_w5318_
	);
	LUT2 #(
		.INIT('h8)
	) name4359 (
		_w2685_,
		_w3715_,
		_w5319_
	);
	LUT2 #(
		.INIT('h8)
	) name4360 (
		_w1184_,
		_w5319_,
		_w5320_
	);
	LUT3 #(
		.INIT('h40)
	) name4361 (
		\u5_cmd_asserted_reg/NET0131 ,
		_w1035_,
		_w1283_,
		_w5321_
	);
	LUT2 #(
		.INIT('he)
	) name4362 (
		_w5320_,
		_w5321_,
		_w5322_
	);
	LUT2 #(
		.INIT('h1)
	) name4363 (
		\u5_cmd_asserted_reg/NET0131 ,
		\u5_state_reg[28]/NET0131 ,
		_w5323_
	);
	LUT3 #(
		.INIT('h08)
	) name4364 (
		_w1068_,
		_w1288_,
		_w5323_,
		_w5324_
	);
	LUT2 #(
		.INIT('h2)
	) name4365 (
		\u5_state_reg[28]/NET0131 ,
		\u5_tmr_done_reg/NET0131 ,
		_w5325_
	);
	LUT3 #(
		.INIT('hdc)
	) name4366 (
		_w2216_,
		_w5324_,
		_w5325_,
		_w5326_
	);
	LUT2 #(
		.INIT('h1)
	) name4367 (
		\u5_cmd_asserted_reg/NET0131 ,
		\u5_state_reg[30]/NET0131 ,
		_w5327_
	);
	LUT3 #(
		.INIT('h08)
	) name4368 (
		_w1068_,
		_w1070_,
		_w5327_,
		_w5328_
	);
	LUT3 #(
		.INIT('h40)
	) name4369 (
		\u5_resume_req_r_reg/NET0131 ,
		_w1035_,
		_w1050_,
		_w5329_
	);
	LUT2 #(
		.INIT('he)
	) name4370 (
		_w5328_,
		_w5329_,
		_w5330_
	);
	LUT3 #(
		.INIT('h4c)
	) name4371 (
		_w1581_,
		_w1586_,
		_w2021_,
		_w5331_
	);
	LUT2 #(
		.INIT('h1)
	) name4372 (
		\u5_state_reg[33]/NET0131 ,
		_w2023_,
		_w5332_
	);
	LUT2 #(
		.INIT('h2)
	) name4373 (
		_w5331_,
		_w5332_,
		_w5333_
	);
	LUT3 #(
		.INIT('h40)
	) name4374 (
		\u5_cmd_asserted_reg/NET0131 ,
		_w1068_,
		_w1288_,
		_w5334_
	);
	LUT2 #(
		.INIT('he)
	) name4375 (
		_w4069_,
		_w5334_,
		_w5335_
	);
	LUT2 #(
		.INIT('h2)
	) name4376 (
		\u5_state_reg[32]/NET0131 ,
		\u5_tmr_done_reg/NET0131 ,
		_w5336_
	);
	LUT4 #(
		.INIT('hefaa)
	) name4377 (
		_w1199_,
		_w1207_,
		_w2490_,
		_w5336_,
		_w5337_
	);
	LUT3 #(
		.INIT('h08)
	) name4378 (
		_w1185_,
		_w1582_,
		_w1583_,
		_w5338_
	);
	LUT2 #(
		.INIT('h8)
	) name4379 (
		_w1184_,
		_w5338_,
		_w5339_
	);
	LUT3 #(
		.INIT('h40)
	) name4380 (
		\u5_cmd_asserted_reg/NET0131 ,
		_w982_,
		_w1289_,
		_w5340_
	);
	LUT4 #(
		.INIT('h153f)
	) name4381 (
		_w1002_,
		_w1184_,
		_w1635_,
		_w5340_,
		_w5341_
	);
	LUT2 #(
		.INIT('h4)
	) name4382 (
		_w5339_,
		_w5341_,
		_w5342_
	);
	LUT3 #(
		.INIT('h54)
	) name4383 (
		\u2_row_same_reg/P0001 ,
		_w2252_,
		_w2254_,
		_w5343_
	);
	LUT3 #(
		.INIT('h80)
	) name4384 (
		_w1339_,
		_w2019_,
		_w5343_,
		_w5344_
	);
	LUT4 #(
		.INIT('h33f7)
	) name4385 (
		\u5_state_reg[4]/NET0131 ,
		_w1581_,
		_w2021_,
		_w5344_,
		_w5345_
	);
	LUT3 #(
		.INIT('h8c)
	) name4386 (
		\u5_cmd_asserted2_reg/NET0131 ,
		\u5_state_reg[4]/NET0131 ,
		\u7_mc_br_r_reg/P0001 ,
		_w5346_
	);
	LUT4 #(
		.INIT('h4f00)
	) name4387 (
		_w1533_,
		_w1579_,
		_w1580_,
		_w5346_,
		_w5347_
	);
	LUT2 #(
		.INIT('h2)
	) name4388 (
		_w5341_,
		_w5347_,
		_w5348_
	);
	LUT3 #(
		.INIT('h15)
	) name4389 (
		_w5342_,
		_w5345_,
		_w5348_,
		_w5349_
	);
	LUT2 #(
		.INIT('h1)
	) name4390 (
		\u5_cmd_asserted_reg/NET0131 ,
		\u5_state_reg[23]/NET0131 ,
		_w5350_
	);
	LUT2 #(
		.INIT('h2)
	) name4391 (
		_w1284_,
		_w5350_,
		_w5351_
	);
	LUT3 #(
		.INIT('h80)
	) name4392 (
		_w984_,
		_w1046_,
		_w5351_,
		_w5352_
	);
	LUT2 #(
		.INIT('h8)
	) name4393 (
		_w1035_,
		_w5352_,
		_w5353_
	);
	LUT2 #(
		.INIT('h2)
	) name4394 (
		\u5_state_reg[23]/NET0131 ,
		\u5_tmr_done_reg/NET0131 ,
		_w5354_
	);
	LUT4 #(
		.INIT('hfbf0)
	) name4395 (
		_w1207_,
		_w2490_,
		_w5353_,
		_w5354_,
		_w5355_
	);
	LUT4 #(
		.INIT('h8808)
	) name4396 (
		\u6_write_go_r1_reg/NET0131 ,
		wb_cyc_i_pad,
		wb_stb_i_pad,
		wb_we_i_pad,
		_w5356_
	);
	LUT2 #(
		.INIT('h2)
	) name4397 (
		\u5_state_reg[44]/NET0131 ,
		\u5_tmr2_done_reg/NET0131 ,
		_w5357_
	);
	LUT3 #(
		.INIT('hba)
	) name4398 (
		_w1247_,
		_w1557_,
		_w5357_,
		_w5358_
	);
	LUT4 #(
		.INIT('h5455)
	) name4399 (
		_w1567_,
		_w1724_,
		_w1728_,
		_w1747_,
		_w5359_
	);
	LUT2 #(
		.INIT('h8)
	) name4400 (
		\u6_read_go_r1_reg/NET0131 ,
		wb_cyc_i_pad,
		_w5360_
	);
	LUT2 #(
		.INIT('h1)
	) name4401 (
		\u5_state_reg[39]/NET0131 ,
		\u5_tmr2_done_reg/NET0131 ,
		_w5361_
	);
	LUT3 #(
		.INIT('h08)
	) name4402 (
		_w968_,
		_w1260_,
		_w5361_,
		_w5362_
	);
	LUT4 #(
		.INIT('h0002)
	) name4403 (
		\u5_state_reg[38]/NET0131 ,
		\u5_state_reg[39]/NET0131 ,
		\u5_state_reg[40]/NET0131 ,
		\u5_state_reg[41]/NET0131 ,
		_w5363_
	);
	LUT2 #(
		.INIT('h8)
	) name4404 (
		_w965_,
		_w5363_,
		_w5364_
	);
	LUT4 #(
		.INIT('heca0)
	) name4405 (
		_w1041_,
		_w1063_,
		_w5362_,
		_w5364_,
		_w5365_
	);
	LUT4 #(
		.INIT('hc4c0)
	) name4406 (
		\u5_tmr2_done_reg/NET0131 ,
		_w1041_,
		_w1079_,
		_w1195_,
		_w5366_
	);
	LUT3 #(
		.INIT('h8c)
	) name4407 (
		\u5_cs_le_r_reg/P0001 ,
		\u5_tmr2_done_reg/NET0131 ,
		\u5_wb_cycle_reg/NET0131 ,
		_w5367_
	);
	LUT4 #(
		.INIT('h1f00)
	) name4408 (
		_w1564_,
		_w1566_,
		_w2028_,
		_w5367_,
		_w5368_
	);
	LUT3 #(
		.INIT('h08)
	) name4409 (
		_w1002_,
		_w1166_,
		_w5368_,
		_w5369_
	);
	LUT3 #(
		.INIT('hfd)
	) name4410 (
		_w1066_,
		_w1231_,
		_w5369_,
		_w5370_
	);
	LUT3 #(
		.INIT('he0)
	) name4411 (
		_w2572_,
		_w2574_,
		_w3957_,
		_w5371_
	);
	LUT2 #(
		.INIT('h8)
	) name4412 (
		_w1533_,
		_w5371_,
		_w5372_
	);
	LUT3 #(
		.INIT('he0)
	) name4413 (
		_w1526_,
		_w1531_,
		_w3957_,
		_w5373_
	);
	LUT3 #(
		.INIT('h10)
	) name4414 (
		_w1528_,
		_w1530_,
		_w5373_,
		_w5374_
	);
	LUT4 #(
		.INIT('h2022)
	) name4415 (
		\u2_u0_bank0_open_reg/NET0131 ,
		\u5_rfr_ack_r_reg/NET0131 ,
		_w2609_,
		_w5374_,
		_w5375_
	);
	LUT3 #(
		.INIT('hdc)
	) name4416 (
		_w2605_,
		_w5372_,
		_w5375_,
		_w5376_
	);
	LUT2 #(
		.INIT('h4)
	) name4417 (
		_w1579_,
		_w5371_,
		_w5377_
	);
	LUT4 #(
		.INIT('ha8aa)
	) name4418 (
		\u2_u1_bank0_open_reg/NET0131 ,
		_w1579_,
		_w2609_,
		_w3957_,
		_w5378_
	);
	LUT2 #(
		.INIT('h4)
	) name4419 (
		\u5_rfr_ack_r_reg/NET0131 ,
		_w5378_,
		_w5379_
	);
	LUT3 #(
		.INIT('hdc)
	) name4420 (
		_w2622_,
		_w5377_,
		_w5379_,
		_w5380_
	);
	LUT3 #(
		.INIT('h8b)
	) name4421 (
		\u5_cmd_del_reg[1]/NET0131 ,
		\u5_wr_cycle_reg/NET0131 ,
		_w1324_,
		_w5381_
	);
	LUT3 #(
		.INIT('h10)
	) name4422 (
		\u5_cmd_asserted_reg/NET0131 ,
		\u5_state_reg[19]/NET0131 ,
		\u5_state_reg[20]/NET0131 ,
		_w5382_
	);
	LUT3 #(
		.INIT('h20)
	) name4423 (
		\u5_state_reg[19]/NET0131 ,
		\u5_state_reg[20]/NET0131 ,
		\u5_tmr_done_reg/NET0131 ,
		_w5383_
	);
	LUT4 #(
		.INIT('h8880)
	) name4424 (
		_w1035_,
		_w1148_,
		_w5382_,
		_w5383_,
		_w5384_
	);
	LUT4 #(
		.INIT('hf888)
	) name4425 (
		_w1041_,
		_w1152_,
		_w1174_,
		_w1561_,
		_w5385_
	);
	LUT4 #(
		.INIT('h1555)
	) name4426 (
		\u5_state_reg[12]/NET0131 ,
		_w1603_,
		_w1604_,
		_w1607_,
		_w5386_
	);
	LUT4 #(
		.INIT('h20aa)
	) name4427 (
		_w1045_,
		_w1539_,
		_w1599_,
		_w5386_,
		_w5387_
	);
	LUT3 #(
		.INIT('h8a)
	) name4428 (
		\u5_state_reg[12]/NET0131 ,
		_w1117_,
		_w1946_,
		_w5388_
	);
	LUT4 #(
		.INIT('hfef0)
	) name4429 (
		\u5_mem_ack_r_reg/NET0131 ,
		_w1568_,
		_w1949_,
		_w5388_,
		_w5389_
	);
	LUT2 #(
		.INIT('h8)
	) name4430 (
		_w1259_,
		_w5389_,
		_w5390_
	);
	LUT3 #(
		.INIT('hf8)
	) name4431 (
		_w2327_,
		_w5387_,
		_w5390_,
		_w5391_
	);
	LUT2 #(
		.INIT('h8)
	) name4432 (
		_w967_,
		_w970_,
		_w5392_
	);
	LUT3 #(
		.INIT('h62)
	) name4433 (
		\u5_state_reg[34]/NET0131 ,
		\u5_state_reg[35]/NET0131 ,
		\u7_mc_br_r_reg/P0001 ,
		_w5393_
	);
	LUT3 #(
		.INIT('h80)
	) name4434 (
		_w1041_,
		_w5392_,
		_w5393_,
		_w5394_
	);
	LUT3 #(
		.INIT('h80)
	) name4435 (
		_w991_,
		_w1250_,
		_w1735_,
		_w5395_
	);
	LUT3 #(
		.INIT('h80)
	) name4436 (
		_w991_,
		_w1077_,
		_w1568_,
		_w5396_
	);
	LUT3 #(
		.INIT('ha8)
	) name4437 (
		_w1566_,
		_w5395_,
		_w5396_,
		_w5397_
	);
	LUT4 #(
		.INIT('h0888)
	) name4438 (
		\u3_u0_wr_adr_reg[0]/NET0131 ,
		wb_cyc_i_pad,
		wb_stb_i_pad,
		wb_we_i_pad,
		_w5398_
	);
	LUT4 #(
		.INIT('hf1e0)
	) name4439 (
		_w998_,
		_w1010_,
		_w5398_,
		_w3710_,
		_w5399_
	);
	LUT3 #(
		.INIT('ha8)
	) name4440 (
		\u3_u0_wr_adr_reg[0]/NET0131 ,
		_w998_,
		_w1010_,
		_w5400_
	);
	LUT4 #(
		.INIT('he2aa)
	) name4441 (
		\u7_mc_dqm_r_reg[0]/P0001 ,
		wb_cyc_i_pad,
		\wb_sel_i[0]_pad ,
		wb_stb_i_pad,
		_w5401_
	);
	LUT4 #(
		.INIT('he2aa)
	) name4442 (
		\u7_mc_dqm_r_reg[1]/P0001 ,
		wb_cyc_i_pad,
		\wb_sel_i[1]_pad ,
		wb_stb_i_pad,
		_w5402_
	);
	LUT4 #(
		.INIT('he2aa)
	) name4443 (
		\u7_mc_dqm_r_reg[2]/P0001 ,
		wb_cyc_i_pad,
		\wb_sel_i[2]_pad ,
		wb_stb_i_pad,
		_w5403_
	);
	LUT4 #(
		.INIT('he2aa)
	) name4444 (
		\u7_mc_dqm_r_reg[3]/P0001 ,
		wb_cyc_i_pad,
		\wb_sel_i[3]_pad ,
		wb_stb_i_pad,
		_w5404_
	);
	LUT2 #(
		.INIT('h8)
	) name4445 (
		\u5_cmd_del_reg[0]/NET0131 ,
		\u5_wr_cycle_reg/NET0131 ,
		_w5405_
	);
	LUT2 #(
		.INIT('h4)
	) name4446 (
		\u5_cmd_del_reg[0]/NET0131 ,
		\u5_wr_cycle_reg/NET0131 ,
		_w5406_
	);
	LUT2 #(
		.INIT('h1)
	) name4447 (
		_w1623_,
		_w5405_,
		_w5407_
	);
	LUT3 #(
		.INIT('h13)
	) name4448 (
		_w1644_,
		_w5406_,
		_w5407_,
		_w5408_
	);
	assign \_al_n0  = 1'b0;
	assign \_al_n1  = 1'b1;
	assign \g22/_0_  = _w1012_ ;
	assign \g23/_0_  = _w1011_ ;
	assign \g25_dup61718/_2_  = _w1016_ ;
	assign \g43466/_0_  = _w1351_ ;
	assign \g43467/_0_  = _w1366_ ;
	assign \g43468/_0_  = _w1378_ ;
	assign \g43469/_0_  = _w1390_ ;
	assign \g43470/_0_  = _w1405_ ;
	assign \g43471/_0_  = _w1420_ ;
	assign \g43472/_0_  = _w1435_ ;
	assign \g43473/_0_  = _w1450_ ;
	assign \g43474/_0_  = _w1465_ ;
	assign \g43475/_0_  = _w1480_ ;
	assign \g43476/_0_  = _w1495_ ;
	assign \g43477/_0_  = _w1510_ ;
	assign \g43478/_0_  = _w1525_ ;
	assign \g43512/_0_  = _w1620_ ;
	assign \g43513/_0_  = _w1621_ ;
	assign \g43544/_3_  = _w1645_ ;
	assign \g43545/_0_  = _w1649_ ;
	assign \g43554/_0_  = _w1719_ ;
	assign \g43555/_0_  = _w1887_ ;
	assign \g43557/_0_  = _w1888_ ;
	assign \g43558/_0_  = _w1922_ ;
	assign \g43571/_2_  = _w1963_ ;
	assign \g43632/_0_  = _w1988_ ;
	assign \g43633/_0_  = _w1999_ ;
	assign \g43635/_0_  = _w2009_ ;
	assign \g43636/_0_  = _w2015_ ;
	assign \g43637/_0_  = _w2018_ ;
	assign \g43638/_0_  = _w2033_ ;
	assign \g43639/_0_  = _w2042_ ;
	assign \g43640/_0_  = _w2047_ ;
	assign \g43642/_0_  = _w1205_ ;
	assign \g43662/_0_  = _w2050_ ;
	assign \g43663/_0_  = _w2052_ ;
	assign \g43664/_0_  = _w2054_ ;
	assign \g43665/_0_  = _w2056_ ;
	assign \g43668/_0_  = _w2086_ ;
	assign \g43670/_0_  = _w2099_ ;
	assign \g43671/_0_  = _w2104_ ;
	assign \g43673/_0_  = _w2140_ ;
	assign \g43674/_0_  = _w2173_ ;
	assign \g43692/_0_  = _w2175_ ;
	assign \g43695/_0_  = _w2179_ ;
	assign \g43696/_0_  = _w2181_ ;
	assign \g43697/_0_  = _w2188_ ;
	assign \g43698/_0_  = _w2199_ ;
	assign \g43700/_0_  = _w2212_ ;
	assign \g43701/_0_  = _w2218_ ;
	assign \g43703/_0_  = _w2227_ ;
	assign \g43705/_0_  = _w2237_ ;
	assign \g43707/_0_  = _w2244_ ;
	assign \g43708/_0_  = _w2261_ ;
	assign \g43710/_0_  = _w2269_ ;
	assign \g43717/_0_  = _w2273_ ;
	assign \g43719/_0_  = _w2275_ ;
	assign \g43720/_0_  = _w2277_ ;
	assign \g43721/_0_  = _w2289_ ;
	assign \g43722/_1_  = _w2295_ ;
	assign \g43723/_0_  = _w2299_ ;
	assign \g43725/_0_  = _w2301_ ;
	assign \g43729/_0_  = _w2302_ ;
	assign \g43731/_0_  = _w2307_ ;
	assign \g43734/_0_  = _w2311_ ;
	assign \g43735/_0_  = _w2318_ ;
	assign \g43737/_0_  = _w2319_ ;
	assign \g43744/_0_  = _w2320_ ;
	assign \g43747/_0_  = _w2321_ ;
	assign \g43760/_2_  = _w2324_ ;
	assign \g43770/_1_  = _w2337_ ;
	assign \g43775/_2_  = _w2341_ ;
	assign \g43780/_2_  = _w2355_ ;
	assign \g43786/_0_  = _w2356_ ;
	assign \g43787/_1_  = _w2364_ ;
	assign \g43847/_0_  = _w2372_ ;
	assign \g43848/_1_  = _w2377_ ;
	assign \g43858/_1_  = _w2382_ ;
	assign \g43891/_3_  = _w2416_ ;
	assign \g43895/_0_  = _w2433_ ;
	assign \g43934/_0_  = _w2451_ ;
	assign \g43936/_3_  = _w2468_ ;
	assign \g43954/_3_  = _w2476_ ;
	assign \g43961/_0_  = _w2498_ ;
	assign \g44016/_1_  = _w2500_ ;
	assign \g44067/_0_  = _w2512_ ;
	assign \g44094/_0_  = _w2520_ ;
	assign \g44096/_0_  = _w2534_ ;
	assign \g44104/_0_  = _w2546_ ;
	assign \g44122/_0_  = _w2555_ ;
	assign \g44172/_0_  = _w2475_ ;
	assign \g44209/_0_  = _w2570_ ;
	assign \g44219/_0_  = _w2613_ ;
	assign \g44220/_0_  = _w2620_ ;
	assign \g44222/_0_  = _w2625_ ;
	assign \g44223/_0_  = _w2629_ ;
	assign \g44241/_2_  = _w2639_ ;
	assign \g44252/_0_  = _w2646_ ;
	assign \g44253/_0_  = _w2650_ ;
	assign \g44255/_2_  = _w2660_ ;
	assign \g44263/_2_  = _w2674_ ;
	assign \g44470/_0_  = _w2683_ ;
	assign \g44538/_0_  = _w2714_ ;
	assign \g44539/_0_  = _w2721_ ;
	assign \g44540/_0_  = _w2728_ ;
	assign \g44541/_0_  = _w2735_ ;
	assign \g44542/_0_  = _w2742_ ;
	assign \g44543/_0_  = _w2749_ ;
	assign \g44544/_0_  = _w2756_ ;
	assign \g44545/_0_  = _w2763_ ;
	assign \g44546/_0_  = _w2770_ ;
	assign \g44547/_0_  = _w2777_ ;
	assign \g44548/_0_  = _w2784_ ;
	assign \g44549/_0_  = _w2791_ ;
	assign \g44550/_0_  = _w2798_ ;
	assign \g44551/_0_  = _w2805_ ;
	assign \g44552/_0_  = _w2812_ ;
	assign \g44553/_0_  = _w2819_ ;
	assign \g44554/_0_  = _w2826_ ;
	assign \g44555/_0_  = _w2833_ ;
	assign \g44556/_0_  = _w2840_ ;
	assign \g44557/_0_  = _w2847_ ;
	assign \g44558/_0_  = _w2854_ ;
	assign \g44559/_0_  = _w2861_ ;
	assign \g44560/_0_  = _w2868_ ;
	assign \g44561/_0_  = _w2875_ ;
	assign \g44562/_0_  = _w2882_ ;
	assign \g44563/_0_  = _w2889_ ;
	assign \g44564/_0_  = _w2896_ ;
	assign \g44565/_0_  = _w2903_ ;
	assign \g44566/_0_  = _w2937_ ;
	assign \g44567/_0_  = _w2947_ ;
	assign \g44568/_0_  = _w2957_ ;
	assign \g44569/_0_  = _w2967_ ;
	assign \g44570/_0_  = _w2977_ ;
	assign \g44571/_0_  = _w2987_ ;
	assign \g44572/_0_  = _w2997_ ;
	assign \g44573/_0_  = _w3007_ ;
	assign \g44574/_0_  = _w3017_ ;
	assign \g44575/_0_  = _w3027_ ;
	assign \g44576/_0_  = _w3037_ ;
	assign \g44577/_0_  = _w3047_ ;
	assign \g44578/_0_  = _w3057_ ;
	assign \g44579/_0_  = _w3067_ ;
	assign \g44580/_0_  = _w3077_ ;
	assign \g44581/_0_  = _w3087_ ;
	assign \g44582/_0_  = _w3097_ ;
	assign \g44583/_0_  = _w3107_ ;
	assign \g44584/_0_  = _w3117_ ;
	assign \g44585/_0_  = _w3127_ ;
	assign \g44586/_0_  = _w3137_ ;
	assign \g44588/_0_  = _w3147_ ;
	assign \g44589/_0_  = _w3157_ ;
	assign \g44590/_0_  = _w3167_ ;
	assign \g44591/_0_  = _w3177_ ;
	assign \g44592/_0_  = _w3187_ ;
	assign \g44593/_0_  = _w3197_ ;
	assign \g44594/_0_  = _w3207_ ;
	assign \g44595/_0_  = _w3216_ ;
	assign \g44596/_0_  = _w3226_ ;
	assign \g44636/_2_  = _w3238_ ;
	assign \g44646/_0_  = _w3246_ ;
	assign \g44647/_0_  = _w3253_ ;
	assign \g44648/_0_  = _w3260_ ;
	assign \g44649/_0_  = _w3267_ ;
	assign \g44650/_0_  = _w3274_ ;
	assign \g44651/_0_  = _w3280_ ;
	assign \g44652/_0_  = _w3285_ ;
	assign \g44653/_0_  = _w3290_ ;
	assign \g44654/_0_  = _w3295_ ;
	assign \g44655/_0_  = _w3300_ ;
	assign \g44656/_0_  = _w3305_ ;
	assign \g44657/_0_  = _w3311_ ;
	assign \g44665/_0_  = _w3314_ ;
	assign \g44666/_0_  = _w3320_ ;
	assign \g44667/_0_  = _w3326_ ;
	assign \g44668/_0_  = _w3332_ ;
	assign \g44752/_0_  = _w3343_ ;
	assign \g44753/_0_  = _w3349_ ;
	assign \g44873/_0_  = _w1296_ ;
	assign \g44939/_0_  = _w3357_ ;
	assign \g44942/_0_  = _w3362_ ;
	assign \g44945/_0_  = _w3370_ ;
	assign \g45023/_2_  = _w3379_ ;
	assign \g45090/_0_  = _w3239_ ;
	assign \g45141/_0_  = _w3385_ ;
	assign \g45147/_3_  = _w3391_ ;
	assign \g45155/_0_  = _w3401_ ;
	assign \g45190/_0_  = _w3402_ ;
	assign \g45195/_2_  = _w3411_ ;
	assign \g45199/_2_  = _w3424_ ;
	assign \g45201/_2_  = _w3433_ ;
	assign \g45324/_0_  = _w3442_ ;
	assign \g45334/_2_  = _w3456_ ;
	assign \g45336/_0_  = _w3390_ ;
	assign \g45388/_0_  = _w3462_ ;
	assign \g45391/_0_  = _w3473_ ;
	assign \g45413/_2_  = _w3484_ ;
	assign \g45530/_0_  = _w3493_ ;
	assign \g45532/_0_  = _w3501_ ;
	assign \g45533/_0_  = _w3510_ ;
	assign \g45534/_0_  = _w3516_ ;
	assign \g45739/_2_  = _w3530_ ;
	assign \g45743/_2_  = _w3544_ ;
	assign \g45767/_0_  = _w3562_ ;
	assign \g45782/_0_  = _w3569_ ;
	assign \g45830/_3_  = _w3585_ ;
	assign \g45834/_3_  = _w3601_ ;
	assign \g45835/_3_  = _w3608_ ;
	assign \g45836/_3_  = _w3616_ ;
	assign \g45837/_3_  = _w3622_ ;
	assign \g45839/_3_  = _w3628_ ;
	assign \g45840/_3_  = _w3634_ ;
	assign \g45841/_3_  = _w3640_ ;
	assign \g45842/_3_  = _w3646_ ;
	assign \g45843/_3_  = _w3652_ ;
	assign \g45844/_3_  = _w3657_ ;
	assign \g45845/_3_  = _w3660_ ;
	assign \g46191/_0_  = _w3662_ ;
	assign \g46193/_3_  = _w3666_ ;
	assign \g46256/_3_  = _w3671_ ;
	assign \g46257/_3_  = _w3676_ ;
	assign \g46258/_3_  = _w3681_ ;
	assign \g46259/_3_  = _w3686_ ;
	assign \g46260/_3_  = _w3691_ ;
	assign \g46261/_3_  = _w3696_ ;
	assign \g46262/_3_  = _w3701_ ;
	assign \g46263/_3_  = _w3706_ ;
	assign \g46278/_0_  = _w3709_ ;
	assign \g46292/_0_  = _w3712_ ;
	assign \g46293/_0_  = _w3714_ ;
	assign \g46312/_0_  = _w3720_ ;
	assign \g46367/_2_  = _w3734_ ;
	assign \g46370/_2_  = _w3743_ ;
	assign \g46380/_2_  = _w3756_ ;
	assign \g46386/_2_  = _w3768_ ;
	assign \g46388/_2_  = _w3781_ ;
	assign \g46392/_2_  = _w3793_ ;
	assign \g46395/_2_  = _w3805_ ;
	assign \g46399/_2_  = _w3814_ ;
	assign \g46420/_0_  = _w3815_ ;
	assign \g46446/_0_  = _w3819_ ;
	assign \g46493/_0_  = _w3825_ ;
	assign \g46510/_0_  = _w3826_ ;
	assign \g46669/_2_  = _w3832_ ;
	assign \g46691/_0_  = _w3849_ ;
	assign \g46708/_0_  = _w3850_ ;
	assign \g46721/_00_  = _w3861_ ;
	assign \g46776/_0_  = _w3862_ ;
	assign \g46777/_0_  = _w3866_ ;
	assign \g46778/_0_  = _w3867_ ;
	assign \g46779/_0_  = _w3868_ ;
	assign \g46780/_0_  = _w3872_ ;
	assign \g46782/_0_  = _w3874_ ;
	assign \g46784/_0_  = _w3879_ ;
	assign \g46932/_0_  = _w3887_ ;
	assign \g47112/_0_  = _w3891_ ;
	assign \g47124/_0_  = _w3898_ ;
	assign \g47265/_0_  = _w3904_ ;
	assign \g47270/_0_  = _w3907_ ;
	assign \g47275/_0_  = _w3913_ ;
	assign \g47300/_1_  = _w3914_ ;
	assign \g47305/_1_  = _w3915_ ;
	assign \g47338/_0_  = _w3916_ ;
	assign \g47339/_0_  = _w3921_ ;
	assign \g47352/_0_  = _w4063_ ;
	assign \g47699/_3_  = _w4066_ ;
	assign \g47711/_0_  = _w4070_ ;
	assign \g47719/_3_  = _w4074_ ;
	assign \g47721/_3_  = _w4078_ ;
	assign \g47723/_3_  = _w4082_ ;
	assign \g47853/_0_  = _w4084_ ;
	assign \g48094/_0_  = _w4091_ ;
	assign \g48095/_0_  = _w4098_ ;
	assign \g48177/_2_  = _w4101_ ;
	assign \g48194/_0_  = _w4102_ ;
	assign \g48369/_2_  = _w4106_ ;
	assign \g48371/_2_  = _w4110_ ;
	assign \g48373/_2_  = _w4114_ ;
	assign \g48375/_2_  = _w4118_ ;
	assign \g48377/_2_  = _w4122_ ;
	assign \g48379/_2_  = _w4126_ ;
	assign \g48381/_2_  = _w4130_ ;
	assign \g48383/_2_  = _w4134_ ;
	assign \g48385/_2_  = _w4138_ ;
	assign \g48535/_0_  = _w4140_ ;
	assign \g48569/_0_  = _w4142_ ;
	assign \g48570/_0_  = _w4144_ ;
	assign \g48571/_0_  = _w4146_ ;
	assign \g48836/_0_  = _w4148_ ;
	assign \g48843/_0_  = _w4150_ ;
	assign \g49187/_3_  = _w3568_ ;
	assign \g49375/_2_  = _w4152_ ;
	assign \g49633/_0_  = _w4153_ ;
	assign \g49788/_1_  = _w2626_ ;
	assign \g49800/_1_  = _w2621_ ;
	assign \g49802/_1_  = _w2647_ ;
	assign \g49806/_1_  = _w2576_ ;
	assign \g49853/_1_  = _w2642_ ;
	assign \g49883/_0_  = _w4159_ ;
	assign \g49884/_0_  = _w4164_ ;
	assign \g49885/_0_  = _w4168_ ;
	assign \g49886/_0_  = _w4172_ ;
	assign \g49976/_1_  = _w2616_ ;
	assign \g50038/_0_  = _w4181_ ;
	assign \g50082/_0_  = _w4191_ ;
	assign \g50083/_0_  = _w3846_ ;
	assign \g50167/_3_  = _w4213_ ;
	assign \g50168/_3_  = _w4230_ ;
	assign \g50169/_3_  = _w4247_ ;
	assign \g50170/_3_  = _w4264_ ;
	assign \g50171/_3_  = _w4281_ ;
	assign \g50177/_0_  = _w4284_ ;
	assign \g50190/_0_  = _w4287_ ;
	assign \g50236/_0_  = _w2918_ ;
	assign \g50251/_3_  = _w4304_ ;
	assign \g50256/_0_  = _w2930_ ;
	assign \g50318/_3_  = _w4321_ ;
	assign \g50319/_3_  = _w4338_ ;
	assign \g50350/_3_  = _w4354_ ;
	assign \g50351/_3_  = _w4370_ ;
	assign \g50352/_3_  = _w4386_ ;
	assign \g50353/_3_  = _w4402_ ;
	assign \g50354/_3_  = _w4418_ ;
	assign \g50355/_3_  = _w4434_ ;
	assign \g50361/_2_  = _w4437_ ;
	assign \g50366/_0_  = _w4444_ ;
	assign \g50393/_0_  = _w4445_ ;
	assign \g50552/_1_  = _w1661_ ;
	assign \g51108/_0_  = _w4451_ ;
	assign \g51160/_0_  = _w4456_ ;
	assign \g51290/_1_  = _w4459_ ;
	assign \g51327/_3_  = _w4473_ ;
	assign \g51328/_3_  = _w4487_ ;
	assign \g51329/_3_  = _w4501_ ;
	assign \g51330/_3_  = _w4515_ ;
	assign \g51331/_3_  = _w4529_ ;
	assign \g51332/_3_  = _w4543_ ;
	assign \g51333/_3_  = _w4557_ ;
	assign \g51334/_3_  = _w4571_ ;
	assign \g51339/_3_  = _w4583_ ;
	assign \g51340/_3_  = _w4595_ ;
	assign \g51341/_3_  = _w4607_ ;
	assign \g51342/_3_  = _w4619_ ;
	assign \g51343/_3_  = _w4631_ ;
	assign \g51346/_0_  = _w4635_ ;
	assign \g51347/_0_  = _w4639_ ;
	assign \g51348/_0_  = _w4640_ ;
	assign \g51381/_3_  = _w4656_ ;
	assign \g51382/_3_  = _w4672_ ;
	assign \g51383/_3_  = _w4688_ ;
	assign \g51386/_3_  = _w4704_ ;
	assign \g51387/_3_  = _w4720_ ;
	assign \g51405/_3_  = _w4726_ ;
	assign \g51410/_3_  = _w4732_ ;
	assign \g51883/_0_  = _w4734_ ;
	assign \g51916/_0_  = _w3842_ ;
	assign \g51947/_0_  = _w4738_ ;
	assign \g51948/_0_  = _w4742_ ;
	assign \g51949/_0_  = _w4749_ ;
	assign \g51950/_0_  = _w4753_ ;
	assign \g51951/_0_  = _w4757_ ;
	assign \g51952/_0_  = _w4761_ ;
	assign \g51953/_0_  = _w4765_ ;
	assign \g51954/_0_  = _w4769_ ;
	assign \g51955/_0_  = _w4773_ ;
	assign \g51956/_0_  = _w4777_ ;
	assign \g51957/_0_  = _w4781_ ;
	assign \g51958/_0_  = _w4785_ ;
	assign \g51959/_0_  = _w4789_ ;
	assign \g51960/_0_  = _w4793_ ;
	assign \g51961/_0_  = _w4797_ ;
	assign \g51962/_0_  = _w4801_ ;
	assign \g51963/_0_  = _w4805_ ;
	assign \g51964/_0_  = _w4809_ ;
	assign \g51965/_0_  = _w4813_ ;
	assign \g51967/_0_  = _w4817_ ;
	assign \g51968/_0_  = _w4822_ ;
	assign \g51969/_0_  = _w4826_ ;
	assign \g51970/_0_  = _w4830_ ;
	assign \g51971/_0_  = _w4834_ ;
	assign \g51972/_0_  = _w4838_ ;
	assign \g51973/_0_  = _w4842_ ;
	assign \g51974/_0_  = _w4846_ ;
	assign \g51975/_0_  = _w4850_ ;
	assign \g51976/_0_  = _w4854_ ;
	assign \g51977/_0_  = _w4858_ ;
	assign \g51978/_0_  = _w4862_ ;
	assign \g51979/_0_  = _w4866_ ;
	assign \g51980/_0_  = _w4870_ ;
	assign \g51981/_0_  = _w4874_ ;
	assign \g51982/_0_  = _w4878_ ;
	assign \g51983/_0_  = _w4882_ ;
	assign \g51984/_0_  = _w4886_ ;
	assign \g51985/_0_  = _w4890_ ;
	assign \g51986/_0_  = _w4894_ ;
	assign \g51987/_0_  = _w4898_ ;
	assign \g51988/_0_  = _w4902_ ;
	assign \g51989/_0_  = _w4906_ ;
	assign \g51990/_0_  = _w4910_ ;
	assign \g51991/_0_  = _w4914_ ;
	assign \g51992/_0_  = _w4918_ ;
	assign \g51993/_0_  = _w4922_ ;
	assign \g51994/_0_  = _w4926_ ;
	assign \g51995/_0_  = _w4930_ ;
	assign \g51996/_0_  = _w4934_ ;
	assign \g51997/_0_  = _w4938_ ;
	assign \g51998/_0_  = _w4942_ ;
	assign \g51999/_0_  = _w4946_ ;
	assign \g52000/_0_  = _w4950_ ;
	assign \g52001/_0_  = _w4954_ ;
	assign \g52002/_0_  = _w4957_ ;
	assign \g52003/_0_  = _w4960_ ;
	assign \g52004/_0_  = _w4963_ ;
	assign \g52005/_0_  = _w4966_ ;
	assign \g52006/_0_  = _w4969_ ;
	assign \g52007/_0_  = _w4972_ ;
	assign \g52008/_0_  = _w4976_ ;
	assign \g52009/_0_  = _w4980_ ;
	assign \g52010/_0_  = _w4983_ ;
	assign \g52011/_0_  = _w4986_ ;
	assign \g52012/_0_  = _w4990_ ;
	assign \g52013/_0_  = _w4993_ ;
	assign \g52014/_0_  = _w4997_ ;
	assign \g52015/_0_  = _w5000_ ;
	assign \g52016/_0_  = _w5003_ ;
	assign \g52017/_0_  = _w5006_ ;
	assign \g52018/_0_  = _w5009_ ;
	assign \g52019/_0_  = _w5012_ ;
	assign \g52020/_0_  = _w5015_ ;
	assign \g52021/_0_  = _w5019_ ;
	assign \g52022/_0_  = _w5022_ ;
	assign \g52023/_0_  = _w5025_ ;
	assign \g52024/_0_  = _w5028_ ;
	assign \g52025/_0_  = _w5032_ ;
	assign \g52026/_0_  = _w5036_ ;
	assign \g52027/_0_  = _w5039_ ;
	assign \g52028/_0_  = _w5043_ ;
	assign \g52029/_0_  = _w5047_ ;
	assign \g52030/_0_  = _w5051_ ;
	assign \g52031/_0_  = _w5054_ ;
	assign \g52032/_0_  = _w5057_ ;
	assign \g52033/_0_  = _w5061_ ;
	assign \g52034/_0_  = _w5065_ ;
	assign \g52035/_0_  = _w5069_ ;
	assign \g52036/_0_  = _w5073_ ;
	assign \g52037/_0_  = _w5077_ ;
	assign \g52038/_0_  = _w5081_ ;
	assign \g52039/_0_  = _w5085_ ;
	assign \g52040/_0_  = _w5089_ ;
	assign \g52041/_0_  = _w5093_ ;
	assign \g52042/_0_  = _w5097_ ;
	assign \g52043/_0_  = _w5101_ ;
	assign \g52044/_0_  = _w5105_ ;
	assign \g52045/_0_  = _w5109_ ;
	assign \g52046/_0_  = _w5113_ ;
	assign \g52047/_0_  = _w5117_ ;
	assign \g52049/_0_  = _w5121_ ;
	assign \g52050/_0_  = _w5125_ ;
	assign \g52051/_0_  = _w5128_ ;
	assign \g52052/_0_  = _w5132_ ;
	assign \g52053/_0_  = _w5136_ ;
	assign \g52054/_0_  = _w5140_ ;
	assign \g52055/_0_  = _w5144_ ;
	assign \g52056/_0_  = _w5148_ ;
	assign \g52057/_0_  = _w5152_ ;
	assign \g52058/_0_  = _w5156_ ;
	assign \g52061/_0_  = _w5160_ ;
	assign \g52065/_0_  = _w5164_ ;
	assign \g52066/_0_  = _w5168_ ;
	assign \g52067/_0_  = _w5171_ ;
	assign \g52068/_0_  = _w5175_ ;
	assign \g52069/_0_  = _w5178_ ;
	assign \g52070/_0_  = _w5181_ ;
	assign \g52071/_0_  = _w5184_ ;
	assign \g52073/_0_  = _w5188_ ;
	assign \g52074/_0_  = _w5192_ ;
	assign \g52075/_0_  = _w5195_ ;
	assign \g52082/_0_  = _w5198_ ;
	assign \g52083/_0_  = _w5201_ ;
	assign \g52158/_0_  = _w5202_ ;
	assign \g52201/_0_  = _w5203_ ;
	assign \g52202/_0_  = _w5204_ ;
	assign \g52346/_0_  = _w1677_ ;
	assign \g52351/_0_  = _w5206_ ;
	assign \g52390/_0_  = _w5209_ ;
	assign \g52847/_0_  = _w5210_ ;
	assign \g52854/_0_  = _w5212_ ;
	assign \g52968/_0_  = _w5216_ ;
	assign \g52969/_0_  = _w5220_ ;
	assign \g52970/_0_  = _w5224_ ;
	assign \g52971/_0_  = _w5228_ ;
	assign \g52984/_0_  = _w5230_ ;
	assign \g52994/_0_  = _w3908_ ;
	assign \g53019/_0_  = _w4818_ ;
	assign \g53030/_0_  = _w4745_ ;
	assign \g53094/_1_  = _w4184_ ;
	assign \g53106/_0_  = _w4947_ ;
	assign \g53150/_0_  = _w5234_ ;
	assign \g53256/_0_  = _w5235_ ;
	assign \g53297/_0_  = _w5236_ ;
	assign \g53345/_0_  = _w5237_ ;
	assign \g53359/_0_  = _w5239_ ;
	assign \g53375/_0_  = _w5240_ ;
	assign \g53474/_1__syn_2  = _w5242_ ;
	assign \g53475/_2_  = _w5243_ ;
	assign \g53593/_0_  = _w5245_ ;
	assign \g53643/_1_  = _w5246_ ;
	assign \g53655/_0_  = _w5247_ ;
	assign \g53710/_0_  = _w5248_ ;
	assign \g53786/_0_  = _w5249_ ;
	assign \g53837/_0_  = _w5250_ ;
	assign \g53888/_1_  = _w3880_ ;
	assign \g53909/_0_  = _w1027_ ;
	assign \g54253/_2_  = _w5251_ ;
	assign \g54394/_3_  = _w3821_ ;
	assign \g54413/_0_  = _w5252_ ;
	assign \g55420/_0_  = _w5253_ ;
	assign \g55587/_0_  = _w5254_ ;
	assign \g55852/_0_  = _w739_ ;
	assign \g57020/_0_  = _w298_ ;
	assign \g59450/_0_  = _w5286_ ;
	assign \g59488/_2_  = _w1325_ ;
	assign \g59752/_0_  = _w5291_ ;
	assign \g59786/_0_  = _w5294_ ;
	assign \g59854/_0_  = _w5295_ ;
	assign \g59878/_0_  = _w5298_ ;
	assign \g59902/_0_  = _w5302_ ;
	assign \g59924/_0_  = _w5306_ ;
	assign \g59947/_0_  = _w5312_ ;
	assign \g59972/_0_  = _w5318_ ;
	assign \g59996/_0_  = _w5322_ ;
	assign \g60017/_0_  = _w5326_ ;
	assign \g60040/_0_  = _w5330_ ;
	assign \g60064/_0_  = _w5333_ ;
	assign \g60095/_0_  = _w5335_ ;
	assign \g60119/_0_  = _w5337_ ;
	assign \g60145/_1_  = _w5349_ ;
	assign \g60165/_0_  = _w5355_ ;
	assign \g60407/_2_  = _w1564_ ;
	assign \g60408/_0_  = _w5356_ ;
	assign \g60613/_2_  = _w5358_ ;
	assign \g60649/_0_  = _w5359_ ;
	assign \g60771/_0_  = _w5360_ ;
	assign \g60908/_1_  = _w5365_ ;
	assign \g60911/_0_  = _w5366_ ;
	assign \g60977/_0_  = _w2707_ ;
	assign \g61/_0_  = _w1039_ ;
	assign \g61002/_0_  = _w5370_ ;
	assign \g61308/_0_  = _w5376_ ;
	assign \g61312/_1_  = _w5372_ ;
	assign \g61314/_0_  = _w5380_ ;
	assign \g61319/_1_  = _w5377_ ;
	assign \g61342/_1_  = _w5381_ ;
	assign \g61360/_0_  = _w5384_ ;
	assign \g61377/_0_  = _w5385_ ;
	assign \g61423/_1_  = _w1568_ ;
	assign \g61426/_0_  = _w1567_ ;
	assign \g61479/_1_  = _w5391_ ;
	assign \g61523/_1_  = _w5394_ ;
	assign \g61558/_1_  = _w2409_ ;
	assign \g61652/_0_  = _w5397_ ;
	assign \g61866/_0_  = _w5399_ ;
	assign \g61868/_1_  = _w5400_ ;
	assign \g61887/_0_  = _w1609_ ;
	assign \u7_mc_dqm_r_reg[0]/P0001_reg_syn_3  = _w5401_ ;
	assign \u7_mc_dqm_r_reg[1]/P0001_reg_syn_3  = _w5402_ ;
	assign \u7_mc_dqm_r_reg[2]/P0001_reg_syn_3  = _w5403_ ;
	assign \u7_mc_dqm_r_reg[3]/P0001_reg_syn_3  = _w5404_ ;
	assign \u7_mc_we__reg/_05_  = _w5408_ ;
endmodule;