module top (\a0_pad , \a1_pad , \a2_pad , a_pad, \b0_pad , \b1_pad , \b2_pad , b_pad, \c0_pad , \c1_pad , \c2_pad , \d0_pad , \d1_pad , \d2_pad , \e0_pad , \e1_pad , \e2_pad , \f0_pad , \f1_pad , \f2_pad , \g0_pad , \g1_pad , \g2_pad , g_pad, \h0_pad , \h1_pad , \h2_pad , h_pad, \i0_pad , \i1_pad , \i2_pad , i_pad, \j1_pad , \j2_pad , \k0_pad , \k1_pad , \k2_pad , k_pad, \l0_pad , \l1_pad , \l2_pad , l_pad, \m0_pad , \m1_pad , \m2_pad , m_pad, \n0_pad , \n1_pad , \n2_pad , n_pad, \o0_pad , \o1_pad , \o2_pad , o_pad, \p0_pad , \p1_pad , \p2_pad , p_pad, \q0_pad , \q1_pad , \q2_pad , q_pad, \r0_pad , \r1_pad , \r2_pad , r_pad, \s0_pad , \s1_pad , \s2_pad , s_pad, \t0_pad , \t1_pad , \t2_pad , t_pad, \u0_pad , \u1_pad , \u2_pad , u_pad, \v0_pad , \v1_pad , \v2_pad , v_pad, \w0_pad , \w1_pad , w_pad, \x0_pad , \x1_pad , x_pad, \y0_pad , \y1_pad , y_pad, \z0_pad , \z1_pad , z_pad, \a3_pad , \a4_pad , \a5_pad , \b3_pad , \b4_pad , \b5_pad , \c3_pad , \c4_pad , \c5_pad , \d3_pad , \d4_pad , \d5_pad , \e3_pad , \e4_pad , \e5_pad , \f3_pad , \f4_pad , \f5_pad , \g3_pad , \g4_pad , \g5_pad , \h3_pad , \h4_pad , \h5_pad , \i3_pad , \i4_pad , \i5_pad , \j3_pad , \j4_pad , \j5_pad , \k3_pad , \k4_pad , \k5_pad , \l3_pad , \l4_pad , \l5_pad , \m3_pad , \m4_pad , \m5_pad , \n3_pad , \n4_pad , \n5_pad , \o3_pad , \o4_pad , \o5_pad , \p3_pad , \p4_pad , \q3_pad , \q4_pad , \r3_pad , \r4_pad , \s3_pad , \s4_pad , \t3_pad , \t4_pad , \u3_pad , \u4_pad , \v3_pad , \v4_pad , \w2_pad , \w3_pad , \w4_pad , \x2_pad , \x3_pad , \x4_pad , \y2_pad , \y3_pad , \y4_pad , \z2_pad , \z3_pad , \z4_pad );
	input \a0_pad  ;
	input \a1_pad  ;
	input \a2_pad  ;
	input a_pad ;
	input \b0_pad  ;
	input \b1_pad  ;
	input \b2_pad  ;
	input b_pad ;
	input \c0_pad  ;
	input \c1_pad  ;
	input \c2_pad  ;
	input \d0_pad  ;
	input \d1_pad  ;
	input \d2_pad  ;
	input \e0_pad  ;
	input \e1_pad  ;
	input \e2_pad  ;
	input \f0_pad  ;
	input \f1_pad  ;
	input \f2_pad  ;
	input \g0_pad  ;
	input \g1_pad  ;
	input \g2_pad  ;
	input g_pad ;
	input \h0_pad  ;
	input \h1_pad  ;
	input \h2_pad  ;
	input h_pad ;
	input \i0_pad  ;
	input \i1_pad  ;
	input \i2_pad  ;
	input i_pad ;
	input \j1_pad  ;
	input \j2_pad  ;
	input \k0_pad  ;
	input \k1_pad  ;
	input \k2_pad  ;
	input k_pad ;
	input \l0_pad  ;
	input \l1_pad  ;
	input \l2_pad  ;
	input l_pad ;
	input \m0_pad  ;
	input \m1_pad  ;
	input \m2_pad  ;
	input m_pad ;
	input \n0_pad  ;
	input \n1_pad  ;
	input \n2_pad  ;
	input n_pad ;
	input \o0_pad  ;
	input \o1_pad  ;
	input \o2_pad  ;
	input o_pad ;
	input \p0_pad  ;
	input \p1_pad  ;
	input \p2_pad  ;
	input p_pad ;
	input \q0_pad  ;
	input \q1_pad  ;
	input \q2_pad  ;
	input q_pad ;
	input \r0_pad  ;
	input \r1_pad  ;
	input \r2_pad  ;
	input r_pad ;
	input \s0_pad  ;
	input \s1_pad  ;
	input \s2_pad  ;
	input s_pad ;
	input \t0_pad  ;
	input \t1_pad  ;
	input \t2_pad  ;
	input t_pad ;
	input \u0_pad  ;
	input \u1_pad  ;
	input \u2_pad  ;
	input u_pad ;
	input \v0_pad  ;
	input \v1_pad  ;
	input \v2_pad  ;
	input v_pad ;
	input \w0_pad  ;
	input \w1_pad  ;
	input w_pad ;
	input \x0_pad  ;
	input \x1_pad  ;
	input x_pad ;
	input \y0_pad  ;
	input \y1_pad  ;
	input y_pad ;
	input \z0_pad  ;
	input \z1_pad  ;
	input z_pad ;
	output \a3_pad  ;
	output \a4_pad  ;
	output \a5_pad  ;
	output \b3_pad  ;
	output \b4_pad  ;
	output \b5_pad  ;
	output \c3_pad  ;
	output \c4_pad  ;
	output \c5_pad  ;
	output \d3_pad  ;
	output \d4_pad  ;
	output \d5_pad  ;
	output \e3_pad  ;
	output \e4_pad  ;
	output \e5_pad  ;
	output \f3_pad  ;
	output \f4_pad  ;
	output \f5_pad  ;
	output \g3_pad  ;
	output \g4_pad  ;
	output \g5_pad  ;
	output \h3_pad  ;
	output \h4_pad  ;
	output \h5_pad  ;
	output \i3_pad  ;
	output \i4_pad  ;
	output \i5_pad  ;
	output \j3_pad  ;
	output \j4_pad  ;
	output \j5_pad  ;
	output \k3_pad  ;
	output \k4_pad  ;
	output \k5_pad  ;
	output \l3_pad  ;
	output \l4_pad  ;
	output \l5_pad  ;
	output \m3_pad  ;
	output \m4_pad  ;
	output \m5_pad  ;
	output \n3_pad  ;
	output \n4_pad  ;
	output \n5_pad  ;
	output \o3_pad  ;
	output \o4_pad  ;
	output \o5_pad  ;
	output \p3_pad  ;
	output \p4_pad  ;
	output \q3_pad  ;
	output \q4_pad  ;
	output \r3_pad  ;
	output \r4_pad  ;
	output \s3_pad  ;
	output \s4_pad  ;
	output \t3_pad  ;
	output \t4_pad  ;
	output \u3_pad  ;
	output \u4_pad  ;
	output \v3_pad  ;
	output \v4_pad  ;
	output \w2_pad  ;
	output \w3_pad  ;
	output \w4_pad  ;
	output \x2_pad  ;
	output \x3_pad  ;
	output \x4_pad  ;
	output \y2_pad  ;
	output \y3_pad  ;
	output \y4_pad  ;
	output \z2_pad  ;
	output \z3_pad  ;
	output \z4_pad  ;
	wire _w399_ ;
	wire _w398_ ;
	wire _w397_ ;
	wire _w396_ ;
	wire _w395_ ;
	wire _w394_ ;
	wire _w393_ ;
	wire _w392_ ;
	wire _w391_ ;
	wire _w390_ ;
	wire _w389_ ;
	wire _w388_ ;
	wire _w387_ ;
	wire _w386_ ;
	wire _w385_ ;
	wire _w384_ ;
	wire _w383_ ;
	wire _w382_ ;
	wire _w381_ ;
	wire _w380_ ;
	wire _w379_ ;
	wire _w378_ ;
	wire _w377_ ;
	wire _w376_ ;
	wire _w375_ ;
	wire _w374_ ;
	wire _w373_ ;
	wire _w372_ ;
	wire _w371_ ;
	wire _w370_ ;
	wire _w369_ ;
	wire _w368_ ;
	wire _w367_ ;
	wire _w366_ ;
	wire _w365_ ;
	wire _w364_ ;
	wire _w363_ ;
	wire _w362_ ;
	wire _w361_ ;
	wire _w360_ ;
	wire _w359_ ;
	wire _w358_ ;
	wire _w357_ ;
	wire _w356_ ;
	wire _w355_ ;
	wire _w354_ ;
	wire _w353_ ;
	wire _w352_ ;
	wire _w221_ ;
	wire _w220_ ;
	wire _w219_ ;
	wire _w218_ ;
	wire _w217_ ;
	wire _w216_ ;
	wire _w215_ ;
	wire _w214_ ;
	wire _w213_ ;
	wire _w212_ ;
	wire _w211_ ;
	wire _w210_ ;
	wire _w209_ ;
	wire _w208_ ;
	wire _w207_ ;
	wire _w206_ ;
	wire _w205_ ;
	wire _w204_ ;
	wire _w203_ ;
	wire _w202_ ;
	wire _w201_ ;
	wire _w200_ ;
	wire _w199_ ;
	wire _w198_ ;
	wire _w197_ ;
	wire _w196_ ;
	wire _w195_ ;
	wire _w194_ ;
	wire _w193_ ;
	wire _w192_ ;
	wire _w191_ ;
	wire _w190_ ;
	wire _w189_ ;
	wire _w188_ ;
	wire _w187_ ;
	wire _w186_ ;
	wire _w185_ ;
	wire _w184_ ;
	wire _w183_ ;
	wire _w182_ ;
	wire _w181_ ;
	wire _w180_ ;
	wire _w179_ ;
	wire _w178_ ;
	wire _w177_ ;
	wire _w176_ ;
	wire _w175_ ;
	wire _w174_ ;
	wire _w173_ ;
	wire _w172_ ;
	wire _w171_ ;
	wire _w170_ ;
	wire _w169_ ;
	wire _w168_ ;
	wire _w167_ ;
	wire _w166_ ;
	wire _w165_ ;
	wire _w164_ ;
	wire _w163_ ;
	wire _w162_ ;
	wire _w161_ ;
	wire _w160_ ;
	wire _w159_ ;
	wire _w158_ ;
	wire _w157_ ;
	wire _w156_ ;
	wire _w155_ ;
	wire _w154_ ;
	wire _w123_ ;
	wire _w122_ ;
	wire _w121_ ;
	wire _w120_ ;
	wire _w119_ ;
	wire _w118_ ;
	wire _w117_ ;
	wire _w116_ ;
	wire _w115_ ;
	wire _w114_ ;
	wire _w113_ ;
	wire _w112_ ;
	wire _w111_ ;
	wire _w110_ ;
	wire _w109_ ;
	wire _w108_ ;
	wire _w95_ ;
	wire _w96_ ;
	wire _w97_ ;
	wire _w98_ ;
	wire _w99_ ;
	wire _w100_ ;
	wire _w101_ ;
	wire _w102_ ;
	wire _w103_ ;
	wire _w104_ ;
	wire _w105_ ;
	wire _w106_ ;
	wire _w107_ ;
	wire _w124_ ;
	wire _w125_ ;
	wire _w126_ ;
	wire _w127_ ;
	wire _w128_ ;
	wire _w129_ ;
	wire _w130_ ;
	wire _w131_ ;
	wire _w132_ ;
	wire _w133_ ;
	wire _w134_ ;
	wire _w135_ ;
	wire _w136_ ;
	wire _w137_ ;
	wire _w138_ ;
	wire _w139_ ;
	wire _w140_ ;
	wire _w141_ ;
	wire _w142_ ;
	wire _w143_ ;
	wire _w144_ ;
	wire _w145_ ;
	wire _w146_ ;
	wire _w147_ ;
	wire _w148_ ;
	wire _w149_ ;
	wire _w150_ ;
	wire _w151_ ;
	wire _w152_ ;
	wire _w153_ ;
	wire _w222_ ;
	wire _w223_ ;
	wire _w224_ ;
	wire _w225_ ;
	wire _w226_ ;
	wire _w227_ ;
	wire _w228_ ;
	wire _w229_ ;
	wire _w230_ ;
	wire _w231_ ;
	wire _w232_ ;
	wire _w233_ ;
	wire _w234_ ;
	wire _w235_ ;
	wire _w236_ ;
	wire _w237_ ;
	wire _w238_ ;
	wire _w239_ ;
	wire _w240_ ;
	wire _w241_ ;
	wire _w242_ ;
	wire _w243_ ;
	wire _w244_ ;
	wire _w245_ ;
	wire _w246_ ;
	wire _w247_ ;
	wire _w248_ ;
	wire _w249_ ;
	wire _w250_ ;
	wire _w251_ ;
	wire _w252_ ;
	wire _w253_ ;
	wire _w254_ ;
	wire _w255_ ;
	wire _w256_ ;
	wire _w257_ ;
	wire _w258_ ;
	wire _w259_ ;
	wire _w260_ ;
	wire _w261_ ;
	wire _w262_ ;
	wire _w263_ ;
	wire _w264_ ;
	wire _w265_ ;
	wire _w266_ ;
	wire _w267_ ;
	wire _w268_ ;
	wire _w269_ ;
	wire _w270_ ;
	wire _w271_ ;
	wire _w272_ ;
	wire _w273_ ;
	wire _w274_ ;
	wire _w275_ ;
	wire _w276_ ;
	wire _w277_ ;
	wire _w278_ ;
	wire _w279_ ;
	wire _w280_ ;
	wire _w281_ ;
	wire _w282_ ;
	wire _w283_ ;
	wire _w284_ ;
	wire _w285_ ;
	wire _w286_ ;
	wire _w287_ ;
	wire _w288_ ;
	wire _w289_ ;
	wire _w290_ ;
	wire _w291_ ;
	wire _w292_ ;
	wire _w293_ ;
	wire _w294_ ;
	wire _w295_ ;
	wire _w296_ ;
	wire _w297_ ;
	wire _w298_ ;
	wire _w299_ ;
	wire _w300_ ;
	wire _w301_ ;
	wire _w302_ ;
	wire _w303_ ;
	wire _w304_ ;
	wire _w305_ ;
	wire _w306_ ;
	wire _w307_ ;
	wire _w308_ ;
	wire _w309_ ;
	wire _w310_ ;
	wire _w311_ ;
	wire _w312_ ;
	wire _w313_ ;
	wire _w314_ ;
	wire _w315_ ;
	wire _w316_ ;
	wire _w317_ ;
	wire _w318_ ;
	wire _w319_ ;
	wire _w320_ ;
	wire _w321_ ;
	wire _w322_ ;
	wire _w323_ ;
	wire _w324_ ;
	wire _w325_ ;
	wire _w326_ ;
	wire _w327_ ;
	wire _w328_ ;
	wire _w329_ ;
	wire _w330_ ;
	wire _w331_ ;
	wire _w332_ ;
	wire _w333_ ;
	wire _w334_ ;
	wire _w335_ ;
	wire _w336_ ;
	wire _w337_ ;
	wire _w338_ ;
	wire _w339_ ;
	wire _w340_ ;
	wire _w341_ ;
	wire _w342_ ;
	wire _w343_ ;
	wire _w344_ ;
	wire _w345_ ;
	wire _w346_ ;
	wire _w347_ ;
	wire _w348_ ;
	wire _w349_ ;
	wire _w350_ ;
	wire _w351_ ;
	LUT2 #(
		.INIT('h1)
	) name0 (
		\p2_pad ,
		\q2_pad ,
		_w95_
	);
	LUT2 #(
		.INIT('h4)
	) name1 (
		\r2_pad ,
		_w95_,
		_w96_
	);
	LUT2 #(
		.INIT('h2)
	) name2 (
		\e1_pad ,
		\n2_pad ,
		_w97_
	);
	LUT2 #(
		.INIT('h8)
	) name3 (
		\o2_pad ,
		_w97_,
		_w98_
	);
	LUT2 #(
		.INIT('h8)
	) name4 (
		_w96_,
		_w98_,
		_w99_
	);
	LUT2 #(
		.INIT('h1)
	) name5 (
		\h1_pad ,
		_w99_,
		_w100_
	);
	LUT2 #(
		.INIT('h4)
	) name6 (
		\q0_pad ,
		_w99_,
		_w101_
	);
	LUT2 #(
		.INIT('h1)
	) name7 (
		\c1_pad ,
		_w100_,
		_w102_
	);
	LUT2 #(
		.INIT('h4)
	) name8 (
		_w101_,
		_w102_,
		_w103_
	);
	LUT2 #(
		.INIT('h1)
	) name9 (
		g_pad,
		h_pad,
		_w104_
	);
	LUT2 #(
		.INIT('h8)
	) name10 (
		\h0_pad ,
		_w104_,
		_w105_
	);
	LUT2 #(
		.INIT('h4)
	) name11 (
		i_pad,
		_w105_,
		_w106_
	);
	LUT2 #(
		.INIT('h8)
	) name12 (
		\g0_pad ,
		\v2_pad ,
		_w107_
	);
	LUT2 #(
		.INIT('h8)
	) name13 (
		\m1_pad ,
		_w107_,
		_w108_
	);
	LUT2 #(
		.INIT('h4)
	) name14 (
		_w106_,
		_w108_,
		_w109_
	);
	LUT2 #(
		.INIT('h8)
	) name15 (
		\c0_pad ,
		_w109_,
		_w110_
	);
	LUT2 #(
		.INIT('h2)
	) name16 (
		\e1_pad ,
		\m0_pad ,
		_w111_
	);
	LUT2 #(
		.INIT('h1)
	) name17 (
		\h2_pad ,
		_w111_,
		_w112_
	);
	LUT2 #(
		.INIT('h4)
	) name18 (
		\i2_pad ,
		_w111_,
		_w113_
	);
	LUT2 #(
		.INIT('h1)
	) name19 (
		_w112_,
		_w113_,
		_w114_
	);
	LUT2 #(
		.INIT('h4)
	) name20 (
		_w109_,
		_w114_,
		_w115_
	);
	LUT2 #(
		.INIT('h1)
	) name21 (
		_w110_,
		_w115_,
		_w116_
	);
	LUT2 #(
		.INIT('h1)
	) name22 (
		\i0_pad ,
		_w116_,
		_w117_
	);
	LUT2 #(
		.INIT('h1)
	) name23 (
		\i1_pad ,
		_w99_,
		_w118_
	);
	LUT2 #(
		.INIT('h4)
	) name24 (
		\r0_pad ,
		_w99_,
		_w119_
	);
	LUT2 #(
		.INIT('h1)
	) name25 (
		\c1_pad ,
		_w118_,
		_w120_
	);
	LUT2 #(
		.INIT('h4)
	) name26 (
		_w119_,
		_w120_,
		_w121_
	);
	LUT2 #(
		.INIT('h8)
	) name27 (
		\d0_pad ,
		_w109_,
		_w122_
	);
	LUT2 #(
		.INIT('h1)
	) name28 (
		\i2_pad ,
		_w111_,
		_w123_
	);
	LUT2 #(
		.INIT('h4)
	) name29 (
		\j2_pad ,
		_w111_,
		_w124_
	);
	LUT2 #(
		.INIT('h1)
	) name30 (
		_w123_,
		_w124_,
		_w125_
	);
	LUT2 #(
		.INIT('h4)
	) name31 (
		_w109_,
		_w125_,
		_w126_
	);
	LUT2 #(
		.INIT('h1)
	) name32 (
		_w122_,
		_w126_,
		_w127_
	);
	LUT2 #(
		.INIT('h1)
	) name33 (
		\i0_pad ,
		_w127_,
		_w128_
	);
	LUT2 #(
		.INIT('h8)
	) name34 (
		\e1_pad ,
		\n2_pad ,
		_w129_
	);
	LUT2 #(
		.INIT('h4)
	) name35 (
		\o2_pad ,
		_w129_,
		_w130_
	);
	LUT2 #(
		.INIT('h1)
	) name36 (
		i_pad,
		\q2_pad ,
		_w131_
	);
	LUT2 #(
		.INIT('h4)
	) name37 (
		\p2_pad ,
		\r2_pad ,
		_w132_
	);
	LUT2 #(
		.INIT('h4)
	) name38 (
		_w131_,
		_w132_,
		_w133_
	);
	LUT2 #(
		.INIT('h8)
	) name39 (
		_w130_,
		_w133_,
		_w134_
	);
	LUT2 #(
		.INIT('h1)
	) name40 (
		\s2_pad ,
		_w134_,
		_w135_
	);
	LUT2 #(
		.INIT('h2)
	) name41 (
		\h0_pad ,
		\t2_pad ,
		_w136_
	);
	LUT2 #(
		.INIT('h4)
	) name42 (
		\h0_pad ,
		\t2_pad ,
		_w137_
	);
	LUT2 #(
		.INIT('h1)
	) name43 (
		_w136_,
		_w137_,
		_w138_
	);
	LUT2 #(
		.INIT('h2)
	) name44 (
		_w134_,
		_w138_,
		_w139_
	);
	LUT2 #(
		.INIT('h1)
	) name45 (
		\i0_pad ,
		_w135_,
		_w140_
	);
	LUT2 #(
		.INIT('h4)
	) name46 (
		_w139_,
		_w140_,
		_w141_
	);
	LUT2 #(
		.INIT('h1)
	) name47 (
		\j1_pad ,
		_w99_,
		_w142_
	);
	LUT2 #(
		.INIT('h4)
	) name48 (
		\s0_pad ,
		_w99_,
		_w143_
	);
	LUT2 #(
		.INIT('h1)
	) name49 (
		\c1_pad ,
		_w142_,
		_w144_
	);
	LUT2 #(
		.INIT('h4)
	) name50 (
		_w143_,
		_w144_,
		_w145_
	);
	LUT2 #(
		.INIT('h4)
	) name51 (
		\i0_pad ,
		_w109_,
		_w146_
	);
	LUT2 #(
		.INIT('h8)
	) name52 (
		\e0_pad ,
		_w146_,
		_w147_
	);
	LUT2 #(
		.INIT('h1)
	) name53 (
		\i0_pad ,
		_w109_,
		_w148_
	);
	LUT2 #(
		.INIT('h2)
	) name54 (
		\j2_pad ,
		_w111_,
		_w149_
	);
	LUT2 #(
		.INIT('h8)
	) name55 (
		_w148_,
		_w149_,
		_w150_
	);
	LUT2 #(
		.INIT('h1)
	) name56 (
		_w147_,
		_w150_,
		_w151_
	);
	LUT2 #(
		.INIT('h2)
	) name57 (
		\m1_pad ,
		_w106_,
		_w152_
	);
	LUT2 #(
		.INIT('h2)
	) name58 (
		_w107_,
		_w152_,
		_w153_
	);
	LUT2 #(
		.INIT('h8)
	) name59 (
		\f0_pad ,
		\v2_pad ,
		_w154_
	);
	LUT2 #(
		.INIT('h1)
	) name60 (
		\k0_pad ,
		_w154_,
		_w155_
	);
	LUT2 #(
		.INIT('h4)
	) name61 (
		_w153_,
		_w155_,
		_w156_
	);
	LUT2 #(
		.INIT('h1)
	) name62 (
		\c1_pad ,
		_w156_,
		_w157_
	);
	LUT2 #(
		.INIT('h1)
	) name63 (
		\k1_pad ,
		_w99_,
		_w158_
	);
	LUT2 #(
		.INIT('h4)
	) name64 (
		\t0_pad ,
		_w99_,
		_w159_
	);
	LUT2 #(
		.INIT('h1)
	) name65 (
		\c1_pad ,
		_w158_,
		_w160_
	);
	LUT2 #(
		.INIT('h4)
	) name66 (
		_w159_,
		_w160_,
		_w161_
	);
	LUT2 #(
		.INIT('h2)
	) name67 (
		b_pad,
		\u0_pad ,
		_w162_
	);
	LUT2 #(
		.INIT('h1)
	) name68 (
		\u2_pad ,
		_w162_,
		_w163_
	);
	LUT2 #(
		.INIT('h2)
	) name69 (
		\k2_pad ,
		_w163_,
		_w164_
	);
	LUT2 #(
		.INIT('h4)
	) name70 (
		\k2_pad ,
		_w163_,
		_w165_
	);
	LUT2 #(
		.INIT('h1)
	) name71 (
		\c1_pad ,
		_w164_,
		_w166_
	);
	LUT2 #(
		.INIT('h4)
	) name72 (
		_w165_,
		_w166_,
		_w167_
	);
	LUT2 #(
		.INIT('h8)
	) name73 (
		_w96_,
		_w130_,
		_w168_
	);
	LUT2 #(
		.INIT('h1)
	) name74 (
		\l0_pad ,
		_w168_,
		_w169_
	);
	LUT2 #(
		.INIT('h1)
	) name75 (
		\c1_pad ,
		_w169_,
		_w170_
	);
	LUT2 #(
		.INIT('h1)
	) name76 (
		\l1_pad ,
		_w168_,
		_w171_
	);
	LUT2 #(
		.INIT('h1)
	) name77 (
		\c1_pad ,
		_w171_,
		_w172_
	);
	LUT2 #(
		.INIT('h4)
	) name78 (
		\k2_pad ,
		\m2_pad ,
		_w173_
	);
	LUT2 #(
		.INIT('h2)
	) name79 (
		\l2_pad ,
		_w173_,
		_w174_
	);
	LUT2 #(
		.INIT('h1)
	) name80 (
		_w164_,
		_w174_,
		_w175_
	);
	LUT2 #(
		.INIT('h2)
	) name81 (
		\l2_pad ,
		_w163_,
		_w176_
	);
	LUT2 #(
		.INIT('h8)
	) name82 (
		\k2_pad ,
		_w176_,
		_w177_
	);
	LUT2 #(
		.INIT('h1)
	) name83 (
		\c1_pad ,
		_w175_,
		_w178_
	);
	LUT2 #(
		.INIT('h4)
	) name84 (
		_w177_,
		_w178_,
		_w179_
	);
	LUT2 #(
		.INIT('h1)
	) name85 (
		\i0_pad ,
		_w153_,
		_w180_
	);
	LUT2 #(
		.INIT('h2)
	) name86 (
		\m0_pad ,
		_w107_,
		_w181_
	);
	LUT2 #(
		.INIT('h2)
	) name87 (
		_w180_,
		_w181_,
		_w182_
	);
	LUT2 #(
		.INIT('h4)
	) name88 (
		\k2_pad ,
		\l2_pad ,
		_w183_
	);
	LUT2 #(
		.INIT('h8)
	) name89 (
		\m2_pad ,
		_w183_,
		_w184_
	);
	LUT2 #(
		.INIT('h8)
	) name90 (
		_w104_,
		_w184_,
		_w185_
	);
	LUT2 #(
		.INIT('h1)
	) name91 (
		\m1_pad ,
		_w185_,
		_w186_
	);
	LUT2 #(
		.INIT('h1)
	) name92 (
		\i0_pad ,
		_w107_,
		_w187_
	);
	LUT2 #(
		.INIT('h4)
	) name93 (
		_w186_,
		_w187_,
		_w188_
	);
	LUT2 #(
		.INIT('h8)
	) name94 (
		\m2_pad ,
		_w176_,
		_w189_
	);
	LUT2 #(
		.INIT('h1)
	) name95 (
		\m2_pad ,
		_w176_,
		_w190_
	);
	LUT2 #(
		.INIT('h1)
	) name96 (
		\c1_pad ,
		_w183_,
		_w191_
	);
	LUT2 #(
		.INIT('h4)
	) name97 (
		_w189_,
		_w191_,
		_w192_
	);
	LUT2 #(
		.INIT('h4)
	) name98 (
		_w190_,
		_w192_,
		_w193_
	);
	LUT2 #(
		.INIT('h1)
	) name99 (
		\n0_pad ,
		_w168_,
		_w194_
	);
	LUT2 #(
		.INIT('h1)
	) name100 (
		\c1_pad ,
		\i0_pad ,
		_w195_
	);
	LUT2 #(
		.INIT('h4)
	) name101 (
		_w194_,
		_w195_,
		_w196_
	);
	LUT2 #(
		.INIT('h8)
	) name102 (
		i_pad,
		_w108_,
		_w197_
	);
	LUT2 #(
		.INIT('h4)
	) name103 (
		_w105_,
		_w108_,
		_w198_
	);
	LUT2 #(
		.INIT('h1)
	) name104 (
		\n1_pad ,
		_w111_,
		_w199_
	);
	LUT2 #(
		.INIT('h8)
	) name105 (
		\o1_pad ,
		_w111_,
		_w200_
	);
	LUT2 #(
		.INIT('h1)
	) name106 (
		_w199_,
		_w200_,
		_w201_
	);
	LUT2 #(
		.INIT('h4)
	) name107 (
		_w198_,
		_w201_,
		_w202_
	);
	LUT2 #(
		.INIT('h1)
	) name108 (
		_w197_,
		_w202_,
		_w203_
	);
	LUT2 #(
		.INIT('h1)
	) name109 (
		\i0_pad ,
		_w203_,
		_w204_
	);
	LUT2 #(
		.INIT('h1)
	) name110 (
		\d1_pad ,
		\e1_pad ,
		_w205_
	);
	LUT2 #(
		.INIT('h4)
	) name111 (
		_w184_,
		_w205_,
		_w206_
	);
	LUT2 #(
		.INIT('h2)
	) name112 (
		\n2_pad ,
		_w206_,
		_w207_
	);
	LUT2 #(
		.INIT('h4)
	) name113 (
		\n2_pad ,
		_w206_,
		_w208_
	);
	LUT2 #(
		.INIT('h1)
	) name114 (
		\c1_pad ,
		_w207_,
		_w209_
	);
	LUT2 #(
		.INIT('h4)
	) name115 (
		_w208_,
		_w209_,
		_w210_
	);
	LUT2 #(
		.INIT('h8)
	) name116 (
		\o0_pad ,
		_w195_,
		_w211_
	);
	LUT2 #(
		.INIT('h4)
	) name117 (
		\p1_pad ,
		_w111_,
		_w212_
	);
	LUT2 #(
		.INIT('h2)
	) name118 (
		\o1_pad ,
		_w111_,
		_w213_
	);
	LUT2 #(
		.INIT('h1)
	) name119 (
		_w212_,
		_w213_,
		_w214_
	);
	LUT2 #(
		.INIT('h8)
	) name120 (
		_w148_,
		_w214_,
		_w215_
	);
	LUT2 #(
		.INIT('h1)
	) name121 (
		\o2_pad ,
		_w207_,
		_w216_
	);
	LUT2 #(
		.INIT('h8)
	) name122 (
		\o2_pad ,
		_w207_,
		_w217_
	);
	LUT2 #(
		.INIT('h1)
	) name123 (
		\c1_pad ,
		_w216_,
		_w218_
	);
	LUT2 #(
		.INIT('h4)
	) name124 (
		_w217_,
		_w218_,
		_w219_
	);
	LUT2 #(
		.INIT('h8)
	) name125 (
		\p0_pad ,
		_w195_,
		_w220_
	);
	LUT2 #(
		.INIT('h8)
	) name126 (
		k_pad,
		_w146_,
		_w221_
	);
	LUT2 #(
		.INIT('h1)
	) name127 (
		\p1_pad ,
		_w111_,
		_w222_
	);
	LUT2 #(
		.INIT('h4)
	) name128 (
		\q1_pad ,
		_w111_,
		_w223_
	);
	LUT2 #(
		.INIT('h1)
	) name129 (
		_w222_,
		_w223_,
		_w224_
	);
	LUT2 #(
		.INIT('h8)
	) name130 (
		_w148_,
		_w224_,
		_w225_
	);
	LUT2 #(
		.INIT('h1)
	) name131 (
		_w221_,
		_w225_,
		_w226_
	);
	LUT2 #(
		.INIT('h8)
	) name132 (
		\p2_pad ,
		_w217_,
		_w227_
	);
	LUT2 #(
		.INIT('h1)
	) name133 (
		\p2_pad ,
		_w217_,
		_w228_
	);
	LUT2 #(
		.INIT('h1)
	) name134 (
		\c1_pad ,
		_w227_,
		_w229_
	);
	LUT2 #(
		.INIT('h4)
	) name135 (
		_w228_,
		_w229_,
		_w230_
	);
	LUT2 #(
		.INIT('h8)
	) name136 (
		\q0_pad ,
		_w195_,
		_w231_
	);
	LUT2 #(
		.INIT('h8)
	) name137 (
		l_pad,
		_w109_,
		_w232_
	);
	LUT2 #(
		.INIT('h1)
	) name138 (
		\q1_pad ,
		_w111_,
		_w233_
	);
	LUT2 #(
		.INIT('h4)
	) name139 (
		\r1_pad ,
		_w111_,
		_w234_
	);
	LUT2 #(
		.INIT('h1)
	) name140 (
		_w233_,
		_w234_,
		_w235_
	);
	LUT2 #(
		.INIT('h4)
	) name141 (
		_w109_,
		_w235_,
		_w236_
	);
	LUT2 #(
		.INIT('h1)
	) name142 (
		_w232_,
		_w236_,
		_w237_
	);
	LUT2 #(
		.INIT('h1)
	) name143 (
		\i0_pad ,
		_w237_,
		_w238_
	);
	LUT2 #(
		.INIT('h1)
	) name144 (
		\q2_pad ,
		_w227_,
		_w239_
	);
	LUT2 #(
		.INIT('h8)
	) name145 (
		\q2_pad ,
		_w227_,
		_w240_
	);
	LUT2 #(
		.INIT('h1)
	) name146 (
		\c1_pad ,
		_w239_,
		_w241_
	);
	LUT2 #(
		.INIT('h4)
	) name147 (
		_w240_,
		_w241_,
		_w242_
	);
	LUT2 #(
		.INIT('h8)
	) name148 (
		\r0_pad ,
		_w195_,
		_w243_
	);
	LUT2 #(
		.INIT('h8)
	) name149 (
		m_pad,
		_w109_,
		_w244_
	);
	LUT2 #(
		.INIT('h1)
	) name150 (
		\r1_pad ,
		_w111_,
		_w245_
	);
	LUT2 #(
		.INIT('h4)
	) name151 (
		\s1_pad ,
		_w111_,
		_w246_
	);
	LUT2 #(
		.INIT('h1)
	) name152 (
		_w245_,
		_w246_,
		_w247_
	);
	LUT2 #(
		.INIT('h4)
	) name153 (
		_w109_,
		_w247_,
		_w248_
	);
	LUT2 #(
		.INIT('h1)
	) name154 (
		_w244_,
		_w248_,
		_w249_
	);
	LUT2 #(
		.INIT('h1)
	) name155 (
		\i0_pad ,
		_w249_,
		_w250_
	);
	LUT2 #(
		.INIT('h1)
	) name156 (
		\r2_pad ,
		_w240_,
		_w251_
	);
	LUT2 #(
		.INIT('h8)
	) name157 (
		\r2_pad ,
		_w240_,
		_w252_
	);
	LUT2 #(
		.INIT('h1)
	) name158 (
		\c1_pad ,
		_w251_,
		_w253_
	);
	LUT2 #(
		.INIT('h4)
	) name159 (
		_w252_,
		_w253_,
		_w254_
	);
	LUT2 #(
		.INIT('h8)
	) name160 (
		\s0_pad ,
		_w195_,
		_w255_
	);
	LUT2 #(
		.INIT('h8)
	) name161 (
		n_pad,
		_w109_,
		_w256_
	);
	LUT2 #(
		.INIT('h1)
	) name162 (
		\s1_pad ,
		_w111_,
		_w257_
	);
	LUT2 #(
		.INIT('h4)
	) name163 (
		\t1_pad ,
		_w111_,
		_w258_
	);
	LUT2 #(
		.INIT('h1)
	) name164 (
		_w257_,
		_w258_,
		_w259_
	);
	LUT2 #(
		.INIT('h4)
	) name165 (
		_w109_,
		_w259_,
		_w260_
	);
	LUT2 #(
		.INIT('h1)
	) name166 (
		_w256_,
		_w260_,
		_w261_
	);
	LUT2 #(
		.INIT('h1)
	) name167 (
		\i0_pad ,
		_w261_,
		_w262_
	);
	LUT2 #(
		.INIT('h1)
	) name168 (
		\b1_pad ,
		_w111_,
		_w263_
	);
	LUT2 #(
		.INIT('h4)
	) name169 (
		\n1_pad ,
		_w111_,
		_w264_
	);
	LUT2 #(
		.INIT('h1)
	) name170 (
		\i0_pad ,
		_w263_,
		_w265_
	);
	LUT2 #(
		.INIT('h4)
	) name171 (
		_w264_,
		_w265_,
		_w266_
	);
	LUT2 #(
		.INIT('h8)
	) name172 (
		\t0_pad ,
		_w195_,
		_w267_
	);
	LUT2 #(
		.INIT('h8)
	) name173 (
		o_pad,
		_w109_,
		_w268_
	);
	LUT2 #(
		.INIT('h1)
	) name174 (
		\t1_pad ,
		_w111_,
		_w269_
	);
	LUT2 #(
		.INIT('h4)
	) name175 (
		\u1_pad ,
		_w111_,
		_w270_
	);
	LUT2 #(
		.INIT('h1)
	) name176 (
		_w269_,
		_w270_,
		_w271_
	);
	LUT2 #(
		.INIT('h4)
	) name177 (
		_w109_,
		_w271_,
		_w272_
	);
	LUT2 #(
		.INIT('h1)
	) name178 (
		_w268_,
		_w272_,
		_w273_
	);
	LUT2 #(
		.INIT('h1)
	) name179 (
		\i0_pad ,
		_w273_,
		_w274_
	);
	LUT2 #(
		.INIT('h8)
	) name180 (
		\l1_pad ,
		\s2_pad ,
		_w275_
	);
	LUT2 #(
		.INIT('h1)
	) name181 (
		\t2_pad ,
		_w275_,
		_w276_
	);
	LUT2 #(
		.INIT('h8)
	) name182 (
		\t2_pad ,
		_w275_,
		_w277_
	);
	LUT2 #(
		.INIT('h1)
	) name183 (
		\c1_pad ,
		_w276_,
		_w278_
	);
	LUT2 #(
		.INIT('h4)
	) name184 (
		_w277_,
		_w278_,
		_w279_
	);
	LUT2 #(
		.INIT('h2)
	) name185 (
		b_pad,
		\i0_pad ,
		_w280_
	);
	LUT2 #(
		.INIT('h8)
	) name186 (
		p_pad,
		_w109_,
		_w281_
	);
	LUT2 #(
		.INIT('h1)
	) name187 (
		\u1_pad ,
		_w111_,
		_w282_
	);
	LUT2 #(
		.INIT('h4)
	) name188 (
		\v1_pad ,
		_w111_,
		_w283_
	);
	LUT2 #(
		.INIT('h1)
	) name189 (
		_w282_,
		_w283_,
		_w284_
	);
	LUT2 #(
		.INIT('h4)
	) name190 (
		_w109_,
		_w284_,
		_w285_
	);
	LUT2 #(
		.INIT('h1)
	) name191 (
		_w281_,
		_w285_,
		_w286_
	);
	LUT2 #(
		.INIT('h1)
	) name192 (
		\i0_pad ,
		_w286_,
		_w287_
	);
	LUT2 #(
		.INIT('h4)
	) name193 (
		_w162_,
		_w184_,
		_w288_
	);
	LUT2 #(
		.INIT('h1)
	) name194 (
		\i0_pad ,
		_w163_,
		_w289_
	);
	LUT2 #(
		.INIT('h4)
	) name195 (
		_w288_,
		_w289_,
		_w290_
	);
	LUT2 #(
		.INIT('h2)
	) name196 (
		a_pad,
		\i0_pad ,
		_w291_
	);
	LUT2 #(
		.INIT('h8)
	) name197 (
		q_pad,
		_w109_,
		_w292_
	);
	LUT2 #(
		.INIT('h1)
	) name198 (
		\v1_pad ,
		_w111_,
		_w293_
	);
	LUT2 #(
		.INIT('h4)
	) name199 (
		\w1_pad ,
		_w111_,
		_w294_
	);
	LUT2 #(
		.INIT('h1)
	) name200 (
		_w293_,
		_w294_,
		_w295_
	);
	LUT2 #(
		.INIT('h4)
	) name201 (
		_w109_,
		_w295_,
		_w296_
	);
	LUT2 #(
		.INIT('h1)
	) name202 (
		_w292_,
		_w296_,
		_w297_
	);
	LUT2 #(
		.INIT('h1)
	) name203 (
		\i0_pad ,
		_w297_,
		_w298_
	);
	LUT2 #(
		.INIT('h4)
	) name204 (
		\f0_pad ,
		\v2_pad ,
		_w299_
	);
	LUT2 #(
		.INIT('h1)
	) name205 (
		_w134_,
		_w299_,
		_w300_
	);
	LUT2 #(
		.INIT('h2)
	) name206 (
		_w187_,
		_w300_,
		_w301_
	);
	LUT2 #(
		.INIT('h4)
	) name207 (
		\i0_pad ,
		\v0_pad ,
		_w302_
	);
	LUT2 #(
		.INIT('h8)
	) name208 (
		r_pad,
		_w109_,
		_w303_
	);
	LUT2 #(
		.INIT('h1)
	) name209 (
		\w1_pad ,
		_w111_,
		_w304_
	);
	LUT2 #(
		.INIT('h4)
	) name210 (
		\x1_pad ,
		_w111_,
		_w305_
	);
	LUT2 #(
		.INIT('h1)
	) name211 (
		_w304_,
		_w305_,
		_w306_
	);
	LUT2 #(
		.INIT('h4)
	) name212 (
		_w109_,
		_w306_,
		_w307_
	);
	LUT2 #(
		.INIT('h1)
	) name213 (
		_w303_,
		_w307_,
		_w308_
	);
	LUT2 #(
		.INIT('h1)
	) name214 (
		\i0_pad ,
		_w308_,
		_w309_
	);
	LUT2 #(
		.INIT('h4)
	) name215 (
		\i0_pad ,
		\w0_pad ,
		_w310_
	);
	LUT2 #(
		.INIT('h8)
	) name216 (
		s_pad,
		_w109_,
		_w311_
	);
	LUT2 #(
		.INIT('h1)
	) name217 (
		\x1_pad ,
		_w111_,
		_w312_
	);
	LUT2 #(
		.INIT('h4)
	) name218 (
		\y1_pad ,
		_w111_,
		_w313_
	);
	LUT2 #(
		.INIT('h1)
	) name219 (
		_w312_,
		_w313_,
		_w314_
	);
	LUT2 #(
		.INIT('h4)
	) name220 (
		_w109_,
		_w314_,
		_w315_
	);
	LUT2 #(
		.INIT('h1)
	) name221 (
		_w311_,
		_w315_,
		_w316_
	);
	LUT2 #(
		.INIT('h1)
	) name222 (
		\i0_pad ,
		_w316_,
		_w317_
	);
	LUT2 #(
		.INIT('h4)
	) name223 (
		\i0_pad ,
		\x0_pad ,
		_w318_
	);
	LUT2 #(
		.INIT('h8)
	) name224 (
		t_pad,
		_w109_,
		_w319_
	);
	LUT2 #(
		.INIT('h1)
	) name225 (
		\y1_pad ,
		_w111_,
		_w320_
	);
	LUT2 #(
		.INIT('h4)
	) name226 (
		\z1_pad ,
		_w111_,
		_w321_
	);
	LUT2 #(
		.INIT('h1)
	) name227 (
		_w320_,
		_w321_,
		_w322_
	);
	LUT2 #(
		.INIT('h4)
	) name228 (
		_w109_,
		_w322_,
		_w323_
	);
	LUT2 #(
		.INIT('h1)
	) name229 (
		_w319_,
		_w323_,
		_w324_
	);
	LUT2 #(
		.INIT('h1)
	) name230 (
		\i0_pad ,
		_w324_,
		_w325_
	);
	LUT2 #(
		.INIT('h4)
	) name231 (
		\i0_pad ,
		\y0_pad ,
		_w326_
	);
	LUT2 #(
		.INIT('h8)
	) name232 (
		u_pad,
		_w109_,
		_w327_
	);
	LUT2 #(
		.INIT('h1)
	) name233 (
		\z1_pad ,
		_w111_,
		_w328_
	);
	LUT2 #(
		.INIT('h4)
	) name234 (
		\a2_pad ,
		_w111_,
		_w329_
	);
	LUT2 #(
		.INIT('h1)
	) name235 (
		_w328_,
		_w329_,
		_w330_
	);
	LUT2 #(
		.INIT('h4)
	) name236 (
		_w109_,
		_w330_,
		_w331_
	);
	LUT2 #(
		.INIT('h1)
	) name237 (
		_w327_,
		_w331_,
		_w332_
	);
	LUT2 #(
		.INIT('h1)
	) name238 (
		\i0_pad ,
		_w332_,
		_w333_
	);
	LUT2 #(
		.INIT('h4)
	) name239 (
		\i0_pad ,
		\z0_pad ,
		_w334_
	);
	LUT2 #(
		.INIT('h8)
	) name240 (
		v_pad,
		_w109_,
		_w335_
	);
	LUT2 #(
		.INIT('h1)
	) name241 (
		\a2_pad ,
		_w111_,
		_w336_
	);
	LUT2 #(
		.INIT('h4)
	) name242 (
		\b2_pad ,
		_w111_,
		_w337_
	);
	LUT2 #(
		.INIT('h1)
	) name243 (
		_w336_,
		_w337_,
		_w338_
	);
	LUT2 #(
		.INIT('h4)
	) name244 (
		_w109_,
		_w338_,
		_w339_
	);
	LUT2 #(
		.INIT('h1)
	) name245 (
		_w335_,
		_w339_,
		_w340_
	);
	LUT2 #(
		.INIT('h1)
	) name246 (
		\i0_pad ,
		_w340_,
		_w341_
	);
	LUT2 #(
		.INIT('h2)
	) name247 (
		\a1_pad ,
		\i0_pad ,
		_w342_
	);
	LUT2 #(
		.INIT('h8)
	) name248 (
		w_pad,
		_w109_,
		_w343_
	);
	LUT2 #(
		.INIT('h1)
	) name249 (
		\b2_pad ,
		_w111_,
		_w344_
	);
	LUT2 #(
		.INIT('h4)
	) name250 (
		\c2_pad ,
		_w111_,
		_w345_
	);
	LUT2 #(
		.INIT('h1)
	) name251 (
		_w344_,
		_w345_,
		_w346_
	);
	LUT2 #(
		.INIT('h4)
	) name252 (
		_w109_,
		_w346_,
		_w347_
	);
	LUT2 #(
		.INIT('h1)
	) name253 (
		_w343_,
		_w347_,
		_w348_
	);
	LUT2 #(
		.INIT('h1)
	) name254 (
		\i0_pad ,
		_w348_,
		_w349_
	);
	LUT2 #(
		.INIT('h1)
	) name255 (
		_w134_,
		_w154_,
		_w350_
	);
	LUT2 #(
		.INIT('h8)
	) name256 (
		_w180_,
		_w350_,
		_w351_
	);
	LUT2 #(
		.INIT('h8)
	) name257 (
		x_pad,
		_w109_,
		_w352_
	);
	LUT2 #(
		.INIT('h1)
	) name258 (
		\c2_pad ,
		_w111_,
		_w353_
	);
	LUT2 #(
		.INIT('h4)
	) name259 (
		\d2_pad ,
		_w111_,
		_w354_
	);
	LUT2 #(
		.INIT('h1)
	) name260 (
		_w353_,
		_w354_,
		_w355_
	);
	LUT2 #(
		.INIT('h4)
	) name261 (
		_w109_,
		_w355_,
		_w356_
	);
	LUT2 #(
		.INIT('h1)
	) name262 (
		_w352_,
		_w356_,
		_w357_
	);
	LUT2 #(
		.INIT('h1)
	) name263 (
		\i0_pad ,
		_w357_,
		_w358_
	);
	LUT2 #(
		.INIT('h4)
	) name264 (
		\g0_pad ,
		\i0_pad ,
		_w359_
	);
	LUT2 #(
		.INIT('h4)
	) name265 (
		\m1_pad ,
		\v2_pad ,
		_w360_
	);
	LUT2 #(
		.INIT('h8)
	) name266 (
		_w359_,
		_w360_,
		_w361_
	);
	LUT2 #(
		.INIT('h4)
	) name267 (
		_w106_,
		_w361_,
		_w362_
	);
	LUT2 #(
		.INIT('h8)
	) name268 (
		y_pad,
		_w109_,
		_w363_
	);
	LUT2 #(
		.INIT('h1)
	) name269 (
		\d2_pad ,
		_w111_,
		_w364_
	);
	LUT2 #(
		.INIT('h4)
	) name270 (
		\e2_pad ,
		_w111_,
		_w365_
	);
	LUT2 #(
		.INIT('h1)
	) name271 (
		_w364_,
		_w365_,
		_w366_
	);
	LUT2 #(
		.INIT('h4)
	) name272 (
		_w109_,
		_w366_,
		_w367_
	);
	LUT2 #(
		.INIT('h1)
	) name273 (
		_w363_,
		_w367_,
		_w368_
	);
	LUT2 #(
		.INIT('h1)
	) name274 (
		\i0_pad ,
		_w368_,
		_w369_
	);
	LUT2 #(
		.INIT('h1)
	) name275 (
		\c1_pad ,
		_w206_,
		_w370_
	);
	LUT2 #(
		.INIT('h8)
	) name276 (
		z_pad,
		_w109_,
		_w371_
	);
	LUT2 #(
		.INIT('h1)
	) name277 (
		\e2_pad ,
		_w111_,
		_w372_
	);
	LUT2 #(
		.INIT('h4)
	) name278 (
		\f2_pad ,
		_w111_,
		_w373_
	);
	LUT2 #(
		.INIT('h1)
	) name279 (
		_w372_,
		_w373_,
		_w374_
	);
	LUT2 #(
		.INIT('h4)
	) name280 (
		_w109_,
		_w374_,
		_w375_
	);
	LUT2 #(
		.INIT('h1)
	) name281 (
		_w371_,
		_w375_,
		_w376_
	);
	LUT2 #(
		.INIT('h1)
	) name282 (
		\i0_pad ,
		_w376_,
		_w377_
	);
	LUT2 #(
		.INIT('h1)
	) name283 (
		\f1_pad ,
		_w99_,
		_w378_
	);
	LUT2 #(
		.INIT('h4)
	) name284 (
		\o0_pad ,
		_w99_,
		_w379_
	);
	LUT2 #(
		.INIT('h1)
	) name285 (
		\c1_pad ,
		_w378_,
		_w380_
	);
	LUT2 #(
		.INIT('h4)
	) name286 (
		_w379_,
		_w380_,
		_w381_
	);
	LUT2 #(
		.INIT('h8)
	) name287 (
		\a0_pad ,
		_w109_,
		_w382_
	);
	LUT2 #(
		.INIT('h1)
	) name288 (
		\f2_pad ,
		_w111_,
		_w383_
	);
	LUT2 #(
		.INIT('h4)
	) name289 (
		\g2_pad ,
		_w111_,
		_w384_
	);
	LUT2 #(
		.INIT('h1)
	) name290 (
		_w383_,
		_w384_,
		_w385_
	);
	LUT2 #(
		.INIT('h4)
	) name291 (
		_w109_,
		_w385_,
		_w386_
	);
	LUT2 #(
		.INIT('h1)
	) name292 (
		_w382_,
		_w386_,
		_w387_
	);
	LUT2 #(
		.INIT('h1)
	) name293 (
		\i0_pad ,
		_w387_,
		_w388_
	);
	LUT2 #(
		.INIT('h1)
	) name294 (
		\g1_pad ,
		_w99_,
		_w389_
	);
	LUT2 #(
		.INIT('h4)
	) name295 (
		\p0_pad ,
		_w99_,
		_w390_
	);
	LUT2 #(
		.INIT('h1)
	) name296 (
		\c1_pad ,
		_w389_,
		_w391_
	);
	LUT2 #(
		.INIT('h4)
	) name297 (
		_w390_,
		_w391_,
		_w392_
	);
	LUT2 #(
		.INIT('h8)
	) name298 (
		\b0_pad ,
		_w109_,
		_w393_
	);
	LUT2 #(
		.INIT('h1)
	) name299 (
		\g2_pad ,
		_w111_,
		_w394_
	);
	LUT2 #(
		.INIT('h4)
	) name300 (
		\h2_pad ,
		_w111_,
		_w395_
	);
	LUT2 #(
		.INIT('h1)
	) name301 (
		_w394_,
		_w395_,
		_w396_
	);
	LUT2 #(
		.INIT('h4)
	) name302 (
		_w109_,
		_w396_,
		_w397_
	);
	LUT2 #(
		.INIT('h1)
	) name303 (
		_w393_,
		_w397_,
		_w398_
	);
	LUT2 #(
		.INIT('h1)
	) name304 (
		\i0_pad ,
		_w398_,
		_w399_
	);
	assign \a3_pad  = \j1_pad ;
	assign \a4_pad  = _w103_ ;
	assign \a5_pad  = _w117_ ;
	assign \b3_pad  = \k1_pad ;
	assign \b4_pad  = _w121_ ;
	assign \b5_pad  = _w128_ ;
	assign \c3_pad  = _w141_ ;
	assign \c4_pad  = _w145_ ;
	assign \c5_pad  = _w151_ ;
	assign \d3_pad  = _w157_ ;
	assign \d4_pad  = _w161_ ;
	assign \d5_pad  = _w167_ ;
	assign \e3_pad  = _w170_ ;
	assign \e4_pad  = _w172_ ;
	assign \e5_pad  = _w179_ ;
	assign \f3_pad  = _w182_ ;
	assign \f4_pad  = _w188_ ;
	assign \f5_pad  = _w193_ ;
	assign \g3_pad  = _w196_ ;
	assign \g4_pad  = _w204_ ;
	assign \g5_pad  = _w210_ ;
	assign \h3_pad  = _w211_ ;
	assign \h4_pad  = _w215_ ;
	assign \h5_pad  = _w219_ ;
	assign \i3_pad  = _w220_ ;
	assign \i4_pad  = _w226_ ;
	assign \i5_pad  = _w230_ ;
	assign \j3_pad  = _w231_ ;
	assign \j4_pad  = _w238_ ;
	assign \j5_pad  = _w242_ ;
	assign \k3_pad  = _w243_ ;
	assign \k4_pad  = _w250_ ;
	assign \k5_pad  = _w254_ ;
	assign \l3_pad  = _w255_ ;
	assign \l4_pad  = _w262_ ;
	assign \l5_pad  = _w266_ ;
	assign \m3_pad  = _w267_ ;
	assign \m4_pad  = _w274_ ;
	assign \m5_pad  = _w279_ ;
	assign \n3_pad  = _w280_ ;
	assign \n4_pad  = _w287_ ;
	assign \n5_pad  = _w290_ ;
	assign \o3_pad  = _w291_ ;
	assign \o4_pad  = _w298_ ;
	assign \o5_pad  = _w301_ ;
	assign \p3_pad  = _w302_ ;
	assign \p4_pad  = _w309_ ;
	assign \q3_pad  = _w310_ ;
	assign \q4_pad  = _w317_ ;
	assign \r3_pad  = _w318_ ;
	assign \r4_pad  = _w325_ ;
	assign \s3_pad  = _w326_ ;
	assign \s4_pad  = _w333_ ;
	assign \t3_pad  = _w334_ ;
	assign \t4_pad  = _w341_ ;
	assign \u3_pad  = _w342_ ;
	assign \u4_pad  = _w349_ ;
	assign \v3_pad  = _w351_ ;
	assign \v4_pad  = _w358_ ;
	assign \w2_pad  = \f1_pad ;
	assign \w3_pad  = _w362_ ;
	assign \w4_pad  = _w369_ ;
	assign \x2_pad  = \g1_pad ;
	assign \x3_pad  = _w370_ ;
	assign \x4_pad  = _w377_ ;
	assign \y2_pad  = \h1_pad ;
	assign \y3_pad  = _w381_ ;
	assign \y4_pad  = _w388_ ;
	assign \z2_pad  = \i1_pad ;
	assign \z3_pad  = _w392_ ;
	assign \z4_pad  = _w399_ ;
endmodule;